* NGSPICE file created from opamp697.ext - technology: sky130A

.subckt opamp697 gnd CSoutput output vdd plus minus commonsourceibias outputibias
+ diffpairibias
X0 gnd.t390 commonsourceibias.t58 commonsourceibias.t59 gnd.t293 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X1 a_n2804_13878.t29 a_n2982_13878.t53 a_n2982_13878.t54 vdd.t202 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X2 a_n2804_13878.t3 a_n2982_13878.t68 vdd.t215 vdd.t214 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X3 gnd.t389 commonsourceibias.t80 CSoutput.t167 gnd.t217 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X4 gnd.t386 commonsourceibias.t81 CSoutput.t166 gnd.t247 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X5 CSoutput.t165 commonsourceibias.t82 gnd.t385 gnd.t255 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X6 vdd.t21 a_n8300_8799.t44 CSoutput.t10 vdd.t20 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X7 commonsourceibias.t57 commonsourceibias.t56 gnd.t388 gnd.t224 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X8 gnd.t387 commonsourceibias.t83 CSoutput.t164 gnd.t205 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X9 a_n8300_8799.t1 plus.t5 a_n3827_n3924.t25 gnd.t9 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.9
X10 CSoutput.t11 a_n8300_8799.t45 vdd.t23 vdd.t22 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=3.12 ps=16.78 w=8 l=0.5
X11 gnd.t384 commonsourceibias.t54 commonsourceibias.t55 gnd.t213 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X12 a_n3827_n3924.t38 diffpairibias.t20 gnd.t188 gnd.t187 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=2.73 ps=14.78 w=7 l=1
X13 CSoutput.t163 commonsourceibias.t84 gnd.t380 gnd.t333 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X14 a_n3827_n3924.t24 plus.t6 a_n8300_8799.t5 gnd.t26 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=1.155 ps=7.33 w=7 l=0.9
X15 gnd.t383 commonsourceibias.t52 commonsourceibias.t53 gnd.t191 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X16 a_n2982_8322.t37 a_n2982_13878.t69 a_n8300_8799.t25 vdd.t212 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X17 commonsourceibias.t51 commonsourceibias.t50 gnd.t382 gnd.t244 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X18 gnd.t381 commonsourceibias.t85 CSoutput.t162 gnd.t285 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X19 CSoutput.t0 a_n8300_8799.t46 vdd.t1 vdd.t0 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X20 vdd.t3 a_n8300_8799.t47 CSoutput.t1 vdd.t2 sky130_fd_pr__pfet_01v8 ad=3.12 pd=16.78 as=1.32 ps=8.33 w=8 l=0.5
X21 gnd.t176 gnd.t174 gnd.t175 gnd.t94 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=0 ps=0 w=7 l=1
X22 a_n2982_13878.t2 minus.t5 a_n3827_n3924.t4 gnd.t23 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.9
X23 a_n8300_8799.t4 plus.t7 a_n3827_n3924.t23 gnd.t20 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.9
X24 a_n8300_8799.t15 a_n2982_13878.t70 a_n2982_8322.t36 vdd.t198 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X25 CSoutput.t161 commonsourceibias.t86 gnd.t379 gnd.t262 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X26 a_n2982_13878.t10 minus.t6 a_n3827_n3924.t36 gnd.t28 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.9
X27 vdd.t150 a_n8300_8799.t48 CSoutput.t40 vdd.t128 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X28 gnd.t173 gnd.t170 gnd.t172 gnd.t171 sky130_fd_pr__nfet_01v8 ad=2.34 pd=12.78 as=0 ps=0 w=6 l=2
X29 CSoutput.t160 commonsourceibias.t87 gnd.t378 gnd.t211 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X30 vdd.t151 a_n8300_8799.t49 CSoutput.t41 vdd.t110 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X31 commonsourceibias.t25 commonsourceibias.t24 gnd.t377 gnd.t291 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X32 a_n8300_8799.t29 a_n2982_13878.t71 a_n2982_8322.t35 vdd.t161 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=3.51 ps=18.78 w=9 l=0.5
X33 gnd.t376 commonsourceibias.t88 CSoutput.t159 gnd.t193 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X34 gnd.t169 gnd.t167 gnd.t168 gnd.t83 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=0 ps=0 w=7 l=1
X35 CSoutput.t158 commonsourceibias.t89 gnd.t375 gnd.t232 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X36 CSoutput.t157 commonsourceibias.t90 gnd.t369 gnd.t333 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X37 gnd.t371 commonsourceibias.t18 commonsourceibias.t19 gnd.t285 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X38 outputibias.t7 outputibias.t6 gnd.t36 gnd.t35 sky130_fd_pr__nfet_01v8 ad=2.34 pd=12.78 as=2.34 ps=12.78 w=6 l=2
X39 gnd.t374 commonsourceibias.t22 commonsourceibias.t23 gnd.t201 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=1.155 ps=7.33 w=7 l=1
X40 CSoutput.t156 commonsourceibias.t91 gnd.t373 gnd.t295 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X41 a_n3827_n3924.t22 plus.t8 a_n8300_8799.t0 gnd.t5 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.9
X42 a_n3827_n3924.t3 diffpairibias.t21 gnd.t15 gnd.t14 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=2.73 ps=14.78 w=7 l=1
X43 commonsourceibias.t21 commonsourceibias.t20 gnd.t372 gnd.t197 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X44 a_n3827_n3924.t33 minus.t7 a_n2982_13878.t8 gnd.t179 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.9
X45 CSoutput.t26 a_n8300_8799.t50 vdd.t127 vdd.t108 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X46 vdd.t129 a_n8300_8799.t51 CSoutput.t27 vdd.t128 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X47 CSoutput.t155 commonsourceibias.t92 gnd.t370 gnd.t295 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X48 gnd.t368 commonsourceibias.t16 commonsourceibias.t17 gnd.t272 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X49 CSoutput.t154 commonsourceibias.t93 gnd.t367 gnd.t209 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=2.73 ps=14.78 w=7 l=1
X50 a_n2804_13878.t28 a_n2982_13878.t39 a_n2982_13878.t40 vdd.t171 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X51 a_n2982_13878.t12 a_n2982_13878.t11 a_n2804_13878.t27 vdd.t182 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X52 CSoutput.t170 a_n8300_8799.t52 vdd.t218 vdd.t0 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X53 vdd.t99 vdd.t97 vdd.t98 vdd.t74 sky130_fd_pr__pfet_01v8 ad=3.51 pd=18.78 as=0 ps=0 w=9 l=0.5
X54 a_n3827_n3924.t21 plus.t9 a_n8300_8799.t39 gnd.t391 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.9
X55 vdd.t219 a_n8300_8799.t53 CSoutput.t171 vdd.t2 sky130_fd_pr__pfet_01v8 ad=3.12 pd=16.78 as=1.32 ps=8.33 w=8 l=0.5
X56 CSoutput.t153 commonsourceibias.t94 gnd.t366 gnd.t226 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=2.73 ps=14.78 w=7 l=1
X57 vdd.t230 CSoutput.t192 output.t19 gnd.t401 sky130_fd_pr__nfet_01v8 ad=0.825 pd=5.33 as=0.825 ps=5.33 w=5 l=1
X58 gnd.t365 commonsourceibias.t95 CSoutput.t152 gnd.t247 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X59 plus.t4 gnd.t164 gnd.t166 gnd.t165 sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.5
X60 diffpairibias.t19 diffpairibias.t18 gnd.t47 gnd.t46 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=2.73 ps=14.78 w=7 l=1
X61 CSoutput.t151 commonsourceibias.t96 gnd.t364 gnd.t253 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X62 a_n3827_n3924.t20 plus.t10 a_n8300_8799.t11 gnd.t177 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.9
X63 gnd.t163 gnd.t161 gnd.t162 gnd.t115 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=0 ps=0 w=7 l=0.9
X64 a_n2982_13878.t32 a_n2982_13878.t31 a_n2804_13878.t26 vdd.t197 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X65 a_n8300_8799.t24 a_n2982_13878.t72 a_n2982_8322.t34 vdd.t192 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X66 CSoutput.t150 commonsourceibias.t97 gnd.t362 gnd.t304 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X67 CSoutput.t149 commonsourceibias.t98 gnd.t363 gnd.t275 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X68 CSoutput.t168 a_n8300_8799.t54 vdd.t216 vdd.t155 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X69 commonsourceibias.t15 commonsourceibias.t14 gnd.t361 gnd.t255 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X70 a_n2982_13878.t16 a_n2982_13878.t15 a_n2804_13878.t25 vdd.t213 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X71 gnd.t160 gnd.t158 gnd.t159 gnd.t62 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=0 ps=0 w=7 l=1
X72 vdd.t217 a_n8300_8799.t55 CSoutput.t169 vdd.t100 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X73 vdd.t111 a_n8300_8799.t56 CSoutput.t18 vdd.t110 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X74 CSoutput.t148 commonsourceibias.t99 gnd.t360 gnd.t333 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X75 a_n8300_8799.t22 a_n2982_13878.t73 a_n2982_8322.t33 vdd.t190 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X76 diffpairibias.t17 diffpairibias.t16 gnd.t51 gnd.t50 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=2.73 ps=14.78 w=7 l=1
X77 CSoutput.t19 a_n8300_8799.t57 vdd.t112 vdd.t103 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X78 gnd.t157 gnd.t155 gnd.t156 gnd.t62 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=0 ps=0 w=7 l=1
X79 a_n8300_8799.t26 a_n2982_13878.t74 a_n2982_8322.t32 vdd.t205 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X80 a_n2982_8322.t31 a_n2982_13878.t75 a_n8300_8799.t20 vdd.t213 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X81 CSoutput.t147 commonsourceibias.t100 gnd.t359 gnd.t226 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=2.73 ps=14.78 w=7 l=1
X82 CSoutput.t146 commonsourceibias.t101 gnd.t358 gnd.t275 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X83 vdd.t96 vdd.t94 vdd.t95 vdd.t61 sky130_fd_pr__pfet_01v8 ad=3.12 pd=16.78 as=0 ps=0 w=8 l=0.5
X84 gnd.t154 gnd.t152 gnd.t153 gnd.t98 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=0 ps=0 w=7 l=1
X85 CSoutput.t38 a_n8300_8799.t58 vdd.t148 vdd.t139 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X86 a_n3827_n3924.t44 minus.t8 a_n2982_13878.t63 gnd.t398 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.9
X87 a_n3827_n3924.t19 plus.t11 a_n8300_8799.t8 gnd.t43 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=1.155 ps=7.33 w=7 l=0.9
X88 gnd.t357 commonsourceibias.t102 CSoutput.t145 gnd.t249 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X89 CSoutput.t144 commonsourceibias.t103 gnd.t356 gnd.t270 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X90 gnd.t151 gnd.t149 gnd.t150 gnd.t70 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=0 ps=0 w=7 l=0.9
X91 a_n8300_8799.t9 plus.t12 a_n3827_n3924.t18 gnd.t2 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.9
X92 gnd.t355 commonsourceibias.t104 CSoutput.t143 gnd.t228 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=1.155 ps=7.33 w=7 l=1
X93 gnd.t148 gnd.t146 minus.t4 gnd.t147 sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.39 ps=2.78 w=1 l=0.5
X94 gnd.t145 gnd.t143 gnd.t144 gnd.t94 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=0 ps=0 w=7 l=1
X95 output.t3 outputibias.t8 gnd.t397 gnd.t396 sky130_fd_pr__nfet_01v8 ad=2.34 pd=12.78 as=2.34 ps=12.78 w=6 l=2
X96 a_n3827_n3924.t28 diffpairibias.t22 gnd.t45 gnd.t44 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=2.73 ps=14.78 w=7 l=1
X97 vdd.t149 a_n8300_8799.t59 CSoutput.t39 vdd.t106 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X98 vdd.t158 a_n8300_8799.t60 CSoutput.t46 vdd.t122 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X99 CSoutput.t142 commonsourceibias.t105 gnd.t319 gnd.t203 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X100 a_n2982_13878.t24 a_n2982_13878.t23 a_n2804_13878.t24 vdd.t212 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X101 vdd.t159 a_n8300_8799.t61 CSoutput.t47 vdd.t114 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X102 a_n3827_n3924.t17 plus.t13 a_n8300_8799.t6 gnd.t27 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.9
X103 a_n8300_8799.t27 a_n2982_13878.t76 a_n2982_8322.t30 vdd.t201 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X104 a_n2982_13878.t28 a_n2982_13878.t27 a_n2804_13878.t23 vdd.t166 sky130_fd_pr__pfet_01v8 ad=3.51 pd=18.78 as=1.485 ps=9.33 w=9 l=0.5
X105 gnd.t354 commonsourceibias.t106 CSoutput.t141 gnd.t222 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X106 vdd.t231 CSoutput.t193 output.t18 gnd.t402 sky130_fd_pr__nfet_01v8 ad=0.825 pd=5.33 as=0.825 ps=5.33 w=5 l=1
X107 commonsourceibias.t43 commonsourceibias.t42 gnd.t353 gnd.t232 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X108 gnd.t352 commonsourceibias.t107 CSoutput.t140 gnd.t195 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X109 gnd.t142 gnd.t139 gnd.t141 gnd.t140 sky130_fd_pr__nfet_01v8 ad=1.95 pd=10.78 as=0 ps=0 w=5 l=1
X110 CSoutput.t139 commonsourceibias.t108 gnd.t351 gnd.t224 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X111 CSoutput.t194 a_n2982_8322.t5 sky130_fd_pr__cap_mim_m3_1 l=12 w=12
X112 gnd.t347 commonsourceibias.t38 commonsourceibias.t39 gnd.t230 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X113 CSoutput.t138 commonsourceibias.t109 gnd.t348 gnd.t295 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X114 diffpairibias.t15 diffpairibias.t14 gnd.t411 gnd.t410 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=2.73 ps=14.78 w=7 l=1
X115 vdd.t93 vdd.t91 vdd.t92 vdd.t81 sky130_fd_pr__pfet_01v8 ad=3.51 pd=18.78 as=0 ps=0 w=9 l=0.5
X116 CSoutput.t14 a_n8300_8799.t62 vdd.t104 vdd.t103 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X117 vdd.t90 vdd.t87 vdd.t89 vdd.t88 sky130_fd_pr__pfet_01v8 ad=3.51 pd=18.78 as=0 ps=0 w=9 l=0.5
X118 gnd.t350 commonsourceibias.t110 CSoutput.t137 gnd.t237 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X119 a_n2804_13878.t22 a_n2982_13878.t21 a_n2982_13878.t22 vdd.t176 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=3.51 ps=18.78 w=9 l=0.5
X120 CSoutput.t15 a_n8300_8799.t63 vdd.t105 vdd.t8 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X121 vdd.t232 a_n8300_8799.t64 CSoutput.t182 vdd.t122 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X122 vdd.t211 a_n2982_13878.t77 a_n2982_8322.t13 vdd.t210 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X123 gnd.t349 commonsourceibias.t40 commonsourceibias.t41 gnd.t219 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X124 a_n2982_13878.t52 a_n2982_13878.t51 a_n2804_13878.t21 vdd.t174 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X125 CSoutput.t136 commonsourceibias.t111 gnd.t346 gnd.t240 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X126 vdd.t86 vdd.t84 vdd.t85 vdd.t61 sky130_fd_pr__pfet_01v8 ad=3.12 pd=16.78 as=0 ps=0 w=8 l=0.5
X127 CSoutput.t135 commonsourceibias.t112 gnd.t345 gnd.t291 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X128 a_n2982_8322.t12 a_n2982_13878.t78 vdd.t209 vdd.t208 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X129 a_n3827_n3924.t31 diffpairibias.t23 gnd.t56 gnd.t55 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=2.73 ps=14.78 w=7 l=1
X130 CSoutput.t183 a_n8300_8799.t65 vdd.t233 vdd.t139 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X131 gnd.t332 commonsourceibias.t113 CSoutput.t134 gnd.t293 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X132 commonsourceibias.t37 commonsourceibias.t36 gnd.t344 gnd.t209 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=2.73 ps=14.78 w=7 l=1
X133 vdd.t207 a_n2982_13878.t79 a_n2804_13878.t0 vdd.t206 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X134 gnd.t335 commonsourceibias.t114 CSoutput.t133 gnd.t267 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X135 commonsourceibias.t35 commonsourceibias.t34 gnd.t343 gnd.t211 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X136 vdd.t83 vdd.t80 vdd.t82 vdd.t81 sky130_fd_pr__pfet_01v8 ad=3.51 pd=18.78 as=0 ps=0 w=9 l=0.5
X137 gnd.t342 commonsourceibias.t32 commonsourceibias.t33 gnd.t193 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X138 output.t17 CSoutput.t195 vdd.t147 gnd.t54 sky130_fd_pr__nfet_01v8 ad=0.825 pd=5.33 as=0.825 ps=5.33 w=5 l=1
X139 CSoutput.t132 commonsourceibias.t115 gnd.t341 gnd.t253 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X140 gnd.t340 commonsourceibias.t116 CSoutput.t131 gnd.t205 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X141 vdd.t123 a_n8300_8799.t66 CSoutput.t24 vdd.t122 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X142 a_n2804_13878.t20 a_n2982_13878.t19 a_n2982_13878.t20 vdd.t205 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X143 plus.t3 gnd.t136 gnd.t138 gnd.t137 sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.5
X144 vdd.t124 a_n8300_8799.t67 CSoutput.t25 vdd.t114 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X145 a_n2982_8322.t29 a_n2982_13878.t80 a_n8300_8799.t33 vdd.t191 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X146 CSoutput.t130 commonsourceibias.t117 gnd.t339 gnd.t270 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X147 gnd.t135 gnd.t133 minus.t3 gnd.t134 sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.5
X148 a_n8300_8799.t40 plus.t14 a_n3827_n3924.t16 gnd.t42 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=2.73 ps=14.78 w=7 l=0.9
X149 vdd.t79 vdd.t77 vdd.t78 vdd.t43 sky130_fd_pr__pfet_01v8 ad=3.12 pd=16.78 as=0 ps=0 w=8 l=0.5
X150 commonsourceibias.t7 commonsourceibias.t6 gnd.t338 gnd.t199 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X151 a_n2982_13878.t65 minus.t9 a_n3827_n3924.t47 gnd.t405 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=2.73 ps=14.78 w=7 l=0.9
X152 vdd.t76 vdd.t73 vdd.t75 vdd.t74 sky130_fd_pr__pfet_01v8 ad=3.51 pd=18.78 as=0 ps=0 w=9 l=0.5
X153 a_n2982_8322.t11 a_n2982_13878.t81 vdd.t204 vdd.t203 sky130_fd_pr__pfet_01v8 ad=3.51 pd=18.78 as=1.485 ps=9.33 w=9 l=0.5
X154 a_n8300_8799.t18 a_n2982_13878.t82 a_n2982_8322.t28 vdd.t173 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X155 gnd.t337 commonsourceibias.t118 CSoutput.t129 gnd.t235 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X156 a_n8300_8799.t3 plus.t15 a_n3827_n3924.t15 gnd.t13 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.9
X157 CSoutput.t174 a_n8300_8799.t68 vdd.t222 vdd.t10 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X158 diffpairibias.t13 diffpairibias.t12 gnd.t39 gnd.t38 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=2.73 ps=14.78 w=7 l=1
X159 CSoutput.t196 a_n2982_8322.t4 sky130_fd_pr__cap_mim_m3_1 l=12 w=12
X160 vdd.t223 a_n8300_8799.t69 CSoutput.t175 vdd.t110 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X161 a_n2982_13878.t26 a_n2982_13878.t25 a_n2804_13878.t19 vdd.t185 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X162 a_n8300_8799.t21 a_n2982_13878.t83 a_n2982_8322.t27 vdd.t202 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X163 gnd.t336 commonsourceibias.t4 commonsourceibias.t5 gnd.t205 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X164 a_n2804_13878.t18 a_n2982_13878.t57 a_n2982_13878.t58 vdd.t201 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X165 commonsourceibias.t3 commonsourceibias.t2 gnd.t334 gnd.t333 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X166 gnd.t331 commonsourceibias.t119 CSoutput.t128 gnd.t242 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X167 gnd.t132 gnd.t130 gnd.t131 gnd.t98 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=0 ps=0 w=7 l=1
X168 output.t16 CSoutput.t197 vdd.t126 gnd.t37 sky130_fd_pr__nfet_01v8 ad=0.825 pd=5.33 as=0.825 ps=5.33 w=5 l=1
X169 gnd.t330 commonsourceibias.t120 CSoutput.t127 gnd.t219 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X170 vdd.t72 vdd.t70 vdd.t71 vdd.t29 sky130_fd_pr__pfet_01v8 ad=3.51 pd=18.78 as=0 ps=0 w=9 l=0.5
X171 CSoutput.t44 a_n8300_8799.t70 vdd.t156 vdd.t155 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X172 gnd.t129 gnd.t127 minus.t2 gnd.t128 sky130_fd_pr__nfet_01v8 ad=0.39 pd=2.78 as=0.165 ps=1.33 w=1 l=0.5
X173 vdd.t200 a_n2982_13878.t84 a_n2982_8322.t10 vdd.t199 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=3.51 ps=18.78 w=9 l=0.5
X174 a_n2804_13878.t17 a_n2982_13878.t29 a_n2982_13878.t30 vdd.t198 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X175 output.t2 outputibias.t9 gnd.t404 gnd.t403 sky130_fd_pr__nfet_01v8 ad=2.34 pd=12.78 as=2.34 ps=12.78 w=6 l=2
X176 vdd.t157 a_n8300_8799.t71 CSoutput.t45 vdd.t20 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X177 a_n2982_13878.t67 minus.t10 a_n3827_n3924.t49 gnd.t9 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.9
X178 a_n3827_n3924.t14 plus.t16 a_n8300_8799.t10 gnd.t6 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.9
X179 a_n2982_13878.t42 a_n2982_13878.t41 a_n2804_13878.t16 vdd.t170 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X180 gnd.t126 gnd.t124 gnd.t125 gnd.t94 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=0 ps=0 w=7 l=1
X181 output.t15 CSoutput.t198 vdd.t120 gnd.t31 sky130_fd_pr__nfet_01v8 ad=0.825 pd=5.33 as=0.825 ps=5.33 w=5 l=1
X182 vdd.t121 CSoutput.t199 output.t14 gnd.t32 sky130_fd_pr__nfet_01v8 ad=0.825 pd=5.33 as=0.825 ps=5.33 w=5 l=1
X183 CSoutput.t126 commonsourceibias.t121 gnd.t329 gnd.t203 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X184 gnd.t318 commonsourceibias.t122 CSoutput.t125 gnd.t249 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X185 commonsourceibias.t1 commonsourceibias.t0 gnd.t327 gnd.t262 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X186 gnd.t317 commonsourceibias.t123 CSoutput.t124 gnd.t247 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X187 vdd.t118 a_n8300_8799.t72 CSoutput.t22 vdd.t18 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X188 gnd.t328 commonsourceibias.t124 CSoutput.t123 gnd.t195 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X189 a_n3827_n3924.t29 diffpairibias.t24 gnd.t49 gnd.t48 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=2.73 ps=14.78 w=7 l=1
X190 a_n3827_n3924.t35 diffpairibias.t25 gnd.t184 gnd.t183 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=2.73 ps=14.78 w=7 l=1
X191 a_n8300_8799.t43 plus.t17 a_n3827_n3924.t13 gnd.t33 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.9
X192 vdd.t119 a_n8300_8799.t73 CSoutput.t23 vdd.t106 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X193 vdd.t69 vdd.t67 vdd.t68 vdd.t43 sky130_fd_pr__pfet_01v8 ad=3.12 pd=16.78 as=0 ps=0 w=8 l=0.5
X194 a_n8300_8799.t7 plus.t18 a_n3827_n3924.t12 gnd.t28 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.9
X195 a_n2804_13878.t15 a_n2982_13878.t55 a_n2982_13878.t56 vdd.t175 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X196 CSoutput.t200 a_n2982_8322.t3 sky130_fd_pr__cap_mim_m3_1 l=12 w=12
X197 a_n2982_8322.t26 a_n2982_13878.t85 a_n8300_8799.t32 vdd.t197 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X198 CSoutput.t190 a_n8300_8799.t74 vdd.t242 vdd.t6 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X199 CSoutput.t201 a_n2982_8322.t2 sky130_fd_pr__cap_mim_m3_1 l=12 w=12
X200 CSoutput.t122 commonsourceibias.t125 gnd.t326 gnd.t304 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X201 output.t13 CSoutput.t202 vdd.t234 gnd.t406 sky130_fd_pr__nfet_01v8 ad=0.825 pd=5.33 as=0.825 ps=5.33 w=5 l=1
X202 gnd.t123 gnd.t121 gnd.t122 gnd.t62 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=0 ps=0 w=7 l=1
X203 gnd.t325 commonsourceibias.t126 CSoutput.t121 gnd.t267 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X204 diffpairibias.t11 diffpairibias.t10 gnd.t393 gnd.t392 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=2.73 ps=14.78 w=7 l=1
X205 gnd.t120 gnd.t118 gnd.t119 gnd.t83 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=0 ps=0 w=7 l=1
X206 a_n2804_13878.t1 a_n2982_13878.t86 vdd.t196 vdd.t195 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X207 a_n2982_13878.t5 minus.t11 a_n3827_n3924.t27 gnd.t12 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.9
X208 vdd.t194 a_n2982_13878.t87 a_n2804_13878.t30 vdd.t193 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X209 gnd.t324 commonsourceibias.t127 CSoutput.t120 gnd.t222 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X210 CSoutput.t191 a_n8300_8799.t75 vdd.t243 vdd.t155 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X211 gnd.t320 commonsourceibias.t128 CSoutput.t119 gnd.t285 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X212 CSoutput.t118 commonsourceibias.t129 gnd.t323 gnd.t209 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=2.73 ps=14.78 w=7 l=1
X213 a_n3827_n3924.t11 plus.t19 a_n8300_8799.t41 gnd.t179 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.9
X214 vdd.t113 a_n8300_8799.t76 CSoutput.t20 vdd.t20 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X215 output.t12 CSoutput.t203 vdd.t235 gnd.t407 sky130_fd_pr__nfet_01v8 ad=0.825 pd=5.33 as=0.825 ps=5.33 w=5 l=1
X216 vdd.t115 a_n8300_8799.t77 CSoutput.t21 vdd.t114 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X217 CSoutput.t8 a_n8300_8799.t78 vdd.t17 vdd.t12 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X218 outputibias.t5 outputibias.t4 gnd.t17 gnd.t16 sky130_fd_pr__nfet_01v8 ad=2.34 pd=12.78 as=2.34 ps=12.78 w=6 l=2
X219 a_n2804_13878.t14 a_n2982_13878.t37 a_n2982_13878.t38 vdd.t192 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X220 diffpairibias.t9 diffpairibias.t8 gnd.t19 gnd.t18 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=2.73 ps=14.78 w=7 l=1
X221 gnd.t322 commonsourceibias.t130 CSoutput.t117 gnd.t242 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X222 gnd.t321 commonsourceibias.t131 CSoutput.t116 gnd.t217 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X223 vdd.t19 a_n8300_8799.t79 CSoutput.t9 vdd.t18 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X224 commonsourceibias.t79 commonsourceibias.t78 gnd.t316 gnd.t304 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X225 a_n3827_n3924.t32 minus.t12 a_n2982_13878.t7 gnd.t178 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.9
X226 a_n2982_8322.t25 a_n2982_13878.t88 a_n8300_8799.t35 vdd.t160 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X227 a_n2982_13878.t18 a_n2982_13878.t17 a_n2804_13878.t13 vdd.t191 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X228 CSoutput.t6 a_n8300_8799.t80 vdd.t15 vdd.t14 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=3.12 ps=16.78 w=8 l=0.5
X229 diffpairibias.t7 diffpairibias.t6 gnd.t395 gnd.t394 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=2.73 ps=14.78 w=7 l=1
X230 vdd.t16 a_n8300_8799.t81 CSoutput.t7 vdd.t2 sky130_fd_pr__pfet_01v8 ad=3.12 pd=16.78 as=1.32 ps=8.33 w=8 l=0.5
X231 a_n2804_13878.t12 a_n2982_13878.t13 a_n2982_13878.t14 vdd.t190 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X232 vdd.t66 vdd.t64 vdd.t65 vdd.t47 sky130_fd_pr__pfet_01v8 ad=3.12 pd=16.78 as=0 ps=0 w=8 l=0.5
X233 vdd.t189 a_n2982_13878.t89 a_n2982_8322.t9 vdd.t188 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=3.51 ps=18.78 w=9 l=0.5
X234 vdd.t107 a_n8300_8799.t82 CSoutput.t16 vdd.t106 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X235 a_n3827_n3924.t43 minus.t13 a_n2982_13878.t62 gnd.t177 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.9
X236 gnd.t117 gnd.t114 gnd.t116 gnd.t115 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=0 ps=0 w=7 l=0.9
X237 CSoutput.t115 commonsourceibias.t132 gnd.t315 gnd.t207 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X238 gnd.t113 gnd.t111 gnd.t112 gnd.t98 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=0 ps=0 w=7 l=1
X239 commonsourceibias.t77 commonsourceibias.t76 gnd.t314 gnd.t226 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=2.73 ps=14.78 w=7 l=1
X240 gnd.t110 gnd.t108 plus.t2 gnd.t109 sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.5
X241 commonsourceibias.t75 commonsourceibias.t74 gnd.t312 gnd.t275 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X242 a_n3827_n3924.t30 minus.t14 a_n2982_13878.t6 gnd.t26 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=1.155 ps=7.33 w=7 l=0.9
X243 CSoutput.t17 a_n8300_8799.t83 vdd.t109 vdd.t108 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X244 minus.t1 gnd.t105 gnd.t107 gnd.t106 sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.5
X245 gnd.t104 gnd.t101 gnd.t103 gnd.t102 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=0 ps=0 w=7 l=1
X246 gnd.t100 gnd.t97 gnd.t99 gnd.t98 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=0 ps=0 w=7 l=1
X247 a_n2804_13878.t4 a_n2982_13878.t90 vdd.t187 vdd.t186 sky130_fd_pr__pfet_01v8 ad=3.51 pd=18.78 as=1.485 ps=9.33 w=9 l=0.5
X248 vdd.t63 vdd.t60 vdd.t62 vdd.t61 sky130_fd_pr__pfet_01v8 ad=3.12 pd=16.78 as=0 ps=0 w=8 l=0.5
X249 vdd.t59 vdd.t57 vdd.t58 vdd.t47 sky130_fd_pr__pfet_01v8 ad=3.12 pd=16.78 as=0 ps=0 w=8 l=0.5
X250 vdd.t4 CSoutput.t204 output.t11 gnd.t3 sky130_fd_pr__nfet_01v8 ad=0.825 pd=5.33 as=0.825 ps=5.33 w=5 l=1
X251 CSoutput.t114 commonsourceibias.t133 gnd.t313 gnd.t207 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X252 gnd.t311 commonsourceibias.t134 CSoutput.t113 gnd.t293 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X253 CSoutput.t28 a_n8300_8799.t84 vdd.t130 vdd.t12 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X254 gnd.t310 commonsourceibias.t72 commonsourceibias.t73 gnd.t228 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=1.155 ps=7.33 w=7 l=1
X255 gnd.t309 commonsourceibias.t135 CSoutput.t112 gnd.t249 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X256 CSoutput.t111 commonsourceibias.t136 gnd.t308 gnd.t224 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X257 gnd.t96 gnd.t93 gnd.t95 gnd.t94 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=0 ps=0 w=7 l=1
X258 CSoutput.t110 commonsourceibias.t137 gnd.t307 gnd.t291 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X259 gnd.t306 commonsourceibias.t138 CSoutput.t109 gnd.t219 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X260 CSoutput.t108 commonsourceibias.t139 gnd.t305 gnd.t304 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X261 vdd.t132 a_n8300_8799.t85 CSoutput.t29 vdd.t131 sky130_fd_pr__pfet_01v8 ad=3.12 pd=16.78 as=1.32 ps=8.33 w=8 l=0.5
X262 vdd.t56 vdd.t54 vdd.t55 vdd.t33 sky130_fd_pr__pfet_01v8 ad=3.12 pd=16.78 as=0 ps=0 w=8 l=0.5
X263 gnd.t92 gnd.t90 gnd.t91 gnd.t83 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=0 ps=0 w=7 l=1
X264 a_n3827_n3924.t39 diffpairibias.t26 gnd.t190 gnd.t189 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=2.73 ps=14.78 w=7 l=1
X265 gnd.t303 commonsourceibias.t140 CSoutput.t107 gnd.t213 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X266 a_n2982_8322.t24 a_n2982_13878.t91 a_n8300_8799.t34 vdd.t185 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X267 commonsourceibias.t71 commonsourceibias.t70 gnd.t302 gnd.t203 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X268 vdd.t5 CSoutput.t205 output.t10 gnd.t4 sky130_fd_pr__nfet_01v8 ad=0.825 pd=5.33 as=0.825 ps=5.33 w=5 l=1
X269 vdd.t184 a_n2982_13878.t92 a_n2982_8322.t8 vdd.t183 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X270 a_n8300_8799.t37 plus.t20 a_n3827_n3924.t10 gnd.t23 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.9
X271 a_n2982_13878.t9 minus.t15 a_n3827_n3924.t34 gnd.t20 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.9
X272 CSoutput.t106 commonsourceibias.t141 gnd.t301 gnd.t244 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X273 gnd.t300 commonsourceibias.t142 CSoutput.t105 gnd.t191 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X274 a_n3827_n3924.t42 minus.t16 a_n2982_13878.t61 gnd.t43 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=1.155 ps=7.33 w=7 l=0.9
X275 CSoutput.t104 commonsourceibias.t143 gnd.t274 gnd.t244 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X276 outputibias.t3 outputibias.t2 gnd.t30 gnd.t29 sky130_fd_pr__nfet_01v8 ad=2.34 pd=12.78 as=2.34 ps=12.78 w=6 l=2
X277 gnd.t299 commonsourceibias.t144 CSoutput.t103 gnd.t272 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X278 gnd.t298 commonsourceibias.t145 CSoutput.t102 gnd.t228 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=1.155 ps=7.33 w=7 l=1
X279 CSoutput.t101 commonsourceibias.t146 gnd.t297 gnd.t199 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X280 gnd.t89 gnd.t86 gnd.t88 gnd.t87 sky130_fd_pr__nfet_01v8 ad=1.95 pd=10.78 as=0 ps=0 w=5 l=1
X281 commonsourceibias.t69 commonsourceibias.t68 gnd.t296 gnd.t295 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X282 vdd.t53 vdd.t50 vdd.t52 vdd.t51 sky130_fd_pr__pfet_01v8 ad=3.51 pd=18.78 as=0 ps=0 w=9 l=0.5
X283 a_n3827_n3924.t46 minus.t17 a_n2982_13878.t64 gnd.t27 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.9
X284 vdd.t138 a_n8300_8799.t86 CSoutput.t32 vdd.t137 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X285 CSoutput.t33 a_n8300_8799.t87 vdd.t140 vdd.t139 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X286 CSoutput.t172 a_n8300_8799.t88 vdd.t220 vdd.t14 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=3.12 ps=16.78 w=8 l=0.5
X287 a_n3827_n3924.t48 minus.t18 a_n2982_13878.t66 gnd.t5 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.9
X288 a_n2804_13878.t11 a_n2982_13878.t35 a_n2982_13878.t36 vdd.t177 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X289 vdd.t49 vdd.t46 vdd.t48 vdd.t47 sky130_fd_pr__pfet_01v8 ad=3.12 pd=16.78 as=0 ps=0 w=8 l=0.5
X290 CSoutput.t100 commonsourceibias.t147 gnd.t278 gnd.t270 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X291 a_n2982_8322.t23 a_n2982_13878.t93 a_n8300_8799.t19 vdd.t182 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X292 output.t1 outputibias.t10 gnd.t409 gnd.t408 sky130_fd_pr__nfet_01v8 ad=2.34 pd=12.78 as=2.34 ps=12.78 w=6 l=2
X293 diffpairibias.t5 diffpairibias.t4 gnd.t8 gnd.t7 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=2.73 ps=14.78 w=7 l=1
X294 gnd.t294 commonsourceibias.t148 CSoutput.t99 gnd.t293 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X295 CSoutput.t98 commonsourceibias.t149 gnd.t292 gnd.t291 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X296 gnd.t290 commonsourceibias.t66 commonsourceibias.t67 gnd.t237 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X297 gnd.t85 gnd.t82 gnd.t84 gnd.t83 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=0 ps=0 w=7 l=1
X298 outputibias.t1 outputibias.t0 gnd.t11 gnd.t10 sky130_fd_pr__nfet_01v8 ad=2.34 pd=12.78 as=2.34 ps=12.78 w=6 l=2
X299 CSoutput.t173 a_n8300_8799.t89 vdd.t221 vdd.t108 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X300 commonsourceibias.t65 commonsourceibias.t64 gnd.t289 gnd.t240 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X301 CSoutput.t4 a_n8300_8799.t90 vdd.t11 vdd.t10 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X302 gnd.t288 commonsourceibias.t150 CSoutput.t97 gnd.t272 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X303 a_n3827_n3924.t45 diffpairibias.t27 gnd.t400 gnd.t399 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=2.73 ps=14.78 w=7 l=1
X304 vdd.t45 vdd.t42 vdd.t44 vdd.t43 sky130_fd_pr__pfet_01v8 ad=3.12 pd=16.78 as=0 ps=0 w=8 l=0.5
X305 gnd.t287 commonsourceibias.t151 CSoutput.t96 gnd.t217 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X306 gnd.t286 commonsourceibias.t152 CSoutput.t95 gnd.t285 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X307 gnd.t284 commonsourceibias.t153 CSoutput.t94 gnd.t201 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=1.155 ps=7.33 w=7 l=1
X308 CSoutput.t206 a_n2982_8322.t1 sky130_fd_pr__cap_mim_m3_1 l=12 w=12
X309 gnd.t81 gnd.t79 plus.t1 gnd.t80 sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.39 ps=2.78 w=1 l=0.5
X310 a_n2982_8322.t7 a_n2982_13878.t94 vdd.t181 vdd.t180 sky130_fd_pr__pfet_01v8 ad=3.51 pd=18.78 as=1.485 ps=9.33 w=9 l=0.5
X311 CSoutput.t5 a_n8300_8799.t91 vdd.t13 vdd.t12 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X312 gnd.t283 commonsourceibias.t154 CSoutput.t93 gnd.t235 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X313 CSoutput.t92 commonsourceibias.t155 gnd.t282 gnd.t197 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X314 output.t9 CSoutput.t207 vdd.t125 gnd.t34 sky130_fd_pr__nfet_01v8 ad=0.825 pd=5.33 as=0.825 ps=5.33 w=5 l=1
X315 gnd.t281 commonsourceibias.t62 commonsourceibias.t63 gnd.t267 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X316 a_n3827_n3924.t41 minus.t19 a_n2982_13878.t60 gnd.t391 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.9
X317 vdd.t153 a_n8300_8799.t92 CSoutput.t42 vdd.t131 sky130_fd_pr__pfet_01v8 ad=3.12 pd=16.78 as=1.32 ps=8.33 w=8 l=0.5
X318 commonsourceibias.t61 commonsourceibias.t60 gnd.t280 gnd.t253 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X319 CSoutput.t43 a_n8300_8799.t93 vdd.t154 vdd.t22 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=3.12 ps=16.78 w=8 l=0.5
X320 vdd.t179 a_n2982_13878.t95 a_n2804_13878.t31 vdd.t178 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=3.51 ps=18.78 w=9 l=0.5
X321 vdd.t240 a_n8300_8799.t94 CSoutput.t188 vdd.t131 sky130_fd_pr__pfet_01v8 ad=3.12 pd=16.78 as=1.32 ps=8.33 w=8 l=0.5
X322 CSoutput.t189 a_n8300_8799.t95 vdd.t241 vdd.t0 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X323 gnd.t273 commonsourceibias.t156 CSoutput.t91 gnd.t272 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X324 CSoutput.t90 commonsourceibias.t157 gnd.t277 gnd.t197 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X325 CSoutput.t89 commonsourceibias.t158 gnd.t276 gnd.t275 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X326 gnd.t279 commonsourceibias.t159 CSoutput.t88 gnd.t193 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X327 commonsourceibias.t31 commonsourceibias.t30 gnd.t271 gnd.t270 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X328 gnd.t196 commonsourceibias.t160 CSoutput.t87 gnd.t195 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X329 gnd.t269 commonsourceibias.t28 commonsourceibias.t29 gnd.t235 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X330 a_n2982_8322.t22 a_n2982_13878.t96 a_n8300_8799.t36 vdd.t172 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X331 a_n8300_8799.t14 a_n2982_13878.t97 a_n2982_8322.t21 vdd.t177 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X332 output.t0 outputibias.t11 gnd.t41 gnd.t40 sky130_fd_pr__nfet_01v8 ad=2.34 pd=12.78 as=2.34 ps=12.78 w=6 l=2
X333 gnd.t268 commonsourceibias.t161 CSoutput.t86 gnd.t267 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X334 a_n2804_13878.t2 a_n2982_13878.t98 vdd.t165 vdd.t164 sky130_fd_pr__pfet_01v8 ad=3.51 pd=18.78 as=1.485 ps=9.33 w=9 l=0.5
X335 CSoutput.t85 commonsourceibias.t162 gnd.t266 gnd.t207 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X336 vdd.t41 vdd.t39 vdd.t40 vdd.t25 sky130_fd_pr__pfet_01v8 ad=3.51 pd=18.78 as=0 ps=0 w=9 l=0.5
X337 CSoutput.t84 commonsourceibias.t163 gnd.t265 gnd.t262 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X338 vdd.t101 a_n8300_8799.t96 CSoutput.t12 vdd.t100 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X339 gnd.t264 commonsourceibias.t164 CSoutput.t83 gnd.t237 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X340 CSoutput.t82 commonsourceibias.t165 gnd.t263 gnd.t262 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X341 CSoutput.t13 a_n8300_8799.t97 vdd.t102 vdd.t14 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=3.12 ps=16.78 w=8 l=0.5
X342 a_n2982_13878.t50 a_n2982_13878.t49 a_n2804_13878.t10 vdd.t167 sky130_fd_pr__pfet_01v8 ad=3.51 pd=18.78 as=1.485 ps=9.33 w=9 l=0.5
X343 vdd.t116 CSoutput.t208 output.t8 gnd.t21 sky130_fd_pr__nfet_01v8 ad=0.825 pd=5.33 as=0.825 ps=5.33 w=5 l=1
X344 gnd.t78 gnd.t76 plus.t0 gnd.t77 sky130_fd_pr__nfet_01v8 ad=0.39 pd=2.78 as=0.165 ps=1.33 w=1 l=0.5
X345 gnd.t261 commonsourceibias.t26 commonsourceibias.t27 gnd.t242 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X346 CSoutput.t81 commonsourceibias.t166 gnd.t260 gnd.t255 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X347 a_n8300_8799.t16 a_n2982_13878.t99 a_n2982_8322.t20 vdd.t176 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=3.51 ps=18.78 w=9 l=0.5
X348 CSoutput.t80 commonsourceibias.t167 gnd.t259 gnd.t240 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X349 a_n3827_n3924.t9 plus.t21 a_n8300_8799.t38 gnd.t398 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.9
X350 minus.t0 gnd.t73 gnd.t75 gnd.t74 sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.5
X351 a_n8300_8799.t31 a_n2982_13878.t100 a_n2982_8322.t19 vdd.t175 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X352 a_n2982_13878.t59 minus.t20 a_n3827_n3924.t40 gnd.t13 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.9
X353 CSoutput.t79 commonsourceibias.t168 gnd.t258 gnd.t199 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X354 gnd.t257 commonsourceibias.t169 CSoutput.t78 gnd.t230 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X355 a_n2982_8322.t18 a_n2982_13878.t101 a_n8300_8799.t30 vdd.t174 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X356 CSoutput.t77 commonsourceibias.t170 gnd.t256 gnd.t255 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X357 gnd.t72 gnd.t69 gnd.t71 gnd.t70 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=0 ps=0 w=7 l=0.9
X358 a_n2982_13878.t0 minus.t21 a_n3827_n3924.t1 gnd.t2 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.9
X359 vdd.t228 a_n8300_8799.t98 CSoutput.t180 vdd.t18 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X360 CSoutput.t181 a_n8300_8799.t99 vdd.t229 vdd.t10 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X361 CSoutput.t186 a_n8300_8799.t100 vdd.t238 vdd.t133 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X362 CSoutput.t76 commonsourceibias.t171 gnd.t254 gnd.t253 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X363 CSoutput.t75 commonsourceibias.t172 gnd.t252 gnd.t232 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X364 gnd.t251 commonsourceibias.t173 CSoutput.t74 gnd.t191 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X365 CSoutput.t187 a_n8300_8799.t101 vdd.t239 vdd.t133 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X366 a_n2804_13878.t9 a_n2982_13878.t47 a_n2982_13878.t48 vdd.t173 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X367 vdd.t145 a_n8300_8799.t102 CSoutput.t36 vdd.t135 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X368 output.t7 CSoutput.t209 vdd.t117 gnd.t22 sky130_fd_pr__nfet_01v8 ad=1.95 pd=10.78 as=0.825 ps=5.33 w=5 l=1
X369 gnd.t250 commonsourceibias.t48 commonsourceibias.t49 gnd.t249 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X370 CSoutput.t210 a_n2982_8322.t0 sky130_fd_pr__cap_mim_m3_1 l=12 w=12
X371 gnd.t248 commonsourceibias.t46 commonsourceibias.t47 gnd.t247 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X372 gnd.t246 commonsourceibias.t44 commonsourceibias.t45 gnd.t195 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X373 a_n3827_n3924.t2 minus.t22 a_n2982_13878.t1 gnd.t6 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.9
X374 a_n3827_n3924.t37 diffpairibias.t28 gnd.t186 gnd.t185 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=2.73 ps=14.78 w=7 l=1
X375 vdd.t146 a_n8300_8799.t103 CSoutput.t37 vdd.t137 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X376 CSoutput.t73 commonsourceibias.t174 gnd.t245 gnd.t244 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X377 gnd.t243 commonsourceibias.t175 CSoutput.t72 gnd.t242 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X378 CSoutput.t178 a_n8300_8799.t104 vdd.t226 vdd.t6 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X379 a_n2982_13878.t46 a_n2982_13878.t45 a_n2804_13878.t8 vdd.t172 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X380 a_n8300_8799.t17 a_n2982_13878.t102 a_n2982_8322.t17 vdd.t171 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X381 vdd.t227 a_n8300_8799.t105 CSoutput.t179 vdd.t135 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X382 CSoutput.t184 a_n8300_8799.t106 vdd.t236 vdd.t103 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X383 vdd.t38 vdd.t36 vdd.t37 vdd.t33 sky130_fd_pr__pfet_01v8 ad=3.12 pd=16.78 as=0 ps=0 w=8 l=0.5
X384 CSoutput.t71 commonsourceibias.t176 gnd.t241 gnd.t240 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X385 gnd.t68 gnd.t65 gnd.t67 gnd.t66 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=0 ps=0 w=7 l=1
X386 gnd.t239 commonsourceibias.t177 CSoutput.t70 gnd.t230 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X387 gnd.t238 commonsourceibias.t178 CSoutput.t69 gnd.t237 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X388 gnd.t236 commonsourceibias.t179 CSoutput.t68 gnd.t235 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X389 CSoutput.t185 a_n8300_8799.t107 vdd.t237 vdd.t8 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X390 diffpairibias.t3 diffpairibias.t2 gnd.t182 gnd.t181 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=2.73 ps=14.78 w=7 l=1
X391 gnd.t234 commonsourceibias.t180 CSoutput.t67 gnd.t222 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X392 CSoutput.t66 commonsourceibias.t181 gnd.t233 gnd.t232 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X393 output.t6 CSoutput.t211 vdd.t152 gnd.t180 sky130_fd_pr__nfet_01v8 ad=0.825 pd=5.33 as=0.825 ps=5.33 w=5 l=1
X394 a_n2982_8322.t16 a_n2982_13878.t103 a_n8300_8799.t23 vdd.t170 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X395 vdd.t141 CSoutput.t212 output.t5 gnd.t52 sky130_fd_pr__nfet_01v8 ad=0.825 pd=5.33 as=1.95 ps=10.78 w=5 l=1
X396 a_n2982_13878.t3 minus.t23 a_n3827_n3924.t5 gnd.t33 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.9
X397 gnd.t231 commonsourceibias.t182 CSoutput.t65 gnd.t230 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X398 gnd.t229 commonsourceibias.t183 CSoutput.t64 gnd.t228 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=1.155 ps=7.33 w=7 l=1
X399 vdd.t143 a_n8300_8799.t108 CSoutput.t34 vdd.t100 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X400 gnd.t64 gnd.t61 gnd.t63 gnd.t62 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=0 ps=0 w=7 l=1
X401 gnd.t60 gnd.t57 gnd.t59 gnd.t58 sky130_fd_pr__nfet_01v8 ad=2.34 pd=12.78 as=0 ps=0 w=6 l=2
X402 CSoutput.t35 a_n8300_8799.t109 vdd.t144 vdd.t22 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=3.12 ps=16.78 w=8 l=0.5
X403 diffpairibias.t1 diffpairibias.t0 gnd.t25 gnd.t24 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=2.73 ps=14.78 w=7 l=1
X404 CSoutput.t63 commonsourceibias.t184 gnd.t227 gnd.t226 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=2.73 ps=14.78 w=7 l=1
X405 CSoutput.t62 commonsourceibias.t185 gnd.t225 gnd.t224 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X406 gnd.t223 commonsourceibias.t12 commonsourceibias.t13 gnd.t222 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X407 gnd.t221 commonsourceibias.t186 CSoutput.t61 gnd.t213 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X408 vdd.t169 a_n2982_13878.t104 a_n2804_13878.t5 vdd.t168 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=3.51 ps=18.78 w=9 l=0.5
X409 CSoutput.t30 a_n8300_8799.t110 vdd.t134 vdd.t133 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X410 gnd.t220 commonsourceibias.t187 CSoutput.t60 gnd.t219 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X411 vdd.t136 a_n8300_8799.t111 CSoutput.t31 vdd.t135 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X412 gnd.t218 commonsourceibias.t10 commonsourceibias.t11 gnd.t217 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X413 gnd.t216 commonsourceibias.t188 CSoutput.t59 gnd.t201 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=1.155 ps=7.33 w=7 l=1
X414 CSoutput.t58 commonsourceibias.t189 gnd.t215 gnd.t211 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X415 a_n8300_8799.t2 plus.t22 a_n3827_n3924.t8 gnd.t12 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.9
X416 a_n2982_8322.t15 a_n2982_13878.t105 a_n8300_8799.t13 vdd.t167 sky130_fd_pr__pfet_01v8 ad=3.51 pd=18.78 as=1.485 ps=9.33 w=9 l=0.5
X417 gnd.t214 commonsourceibias.t190 CSoutput.t57 gnd.t213 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X418 a_n2982_13878.t4 minus.t24 a_n3827_n3924.t26 gnd.t42 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=2.73 ps=14.78 w=7 l=0.9
X419 a_n8300_8799.t42 plus.t23 a_n3827_n3924.t7 gnd.t405 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=2.73 ps=14.78 w=7 l=0.9
X420 a_n2982_8322.t14 a_n2982_13878.t106 a_n8300_8799.t28 vdd.t166 sky130_fd_pr__pfet_01v8 ad=3.51 pd=18.78 as=1.485 ps=9.33 w=9 l=0.5
X421 CSoutput.t56 commonsourceibias.t191 gnd.t210 gnd.t209 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=2.73 ps=14.78 w=7 l=1
X422 CSoutput.t55 commonsourceibias.t192 gnd.t212 gnd.t211 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X423 vdd.t224 a_n8300_8799.t112 CSoutput.t176 vdd.t137 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X424 vdd.t225 a_n8300_8799.t113 CSoutput.t177 vdd.t128 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X425 CSoutput.t2 a_n8300_8799.t114 vdd.t7 vdd.t6 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X426 gnd.t194 commonsourceibias.t193 CSoutput.t54 gnd.t193 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X427 commonsourceibias.t9 commonsourceibias.t8 gnd.t208 gnd.t207 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X428 gnd.t206 commonsourceibias.t194 CSoutput.t53 gnd.t205 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X429 CSoutput.t52 commonsourceibias.t195 gnd.t204 gnd.t203 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X430 vdd.t35 vdd.t32 vdd.t34 vdd.t33 sky130_fd_pr__pfet_01v8 ad=3.12 pd=16.78 as=0 ps=0 w=8 l=0.5
X431 a_n2982_8322.t6 a_n2982_13878.t107 vdd.t163 vdd.t162 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X432 gnd.t202 commonsourceibias.t196 CSoutput.t51 gnd.t201 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=1.155 ps=7.33 w=7 l=1
X433 a_n2804_13878.t7 a_n2982_13878.t43 a_n2982_13878.t44 vdd.t161 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=3.51 ps=18.78 w=9 l=0.5
X434 vdd.t142 CSoutput.t213 output.t4 gnd.t53 sky130_fd_pr__nfet_01v8 ad=0.825 pd=5.33 as=0.825 ps=5.33 w=5 l=1
X435 vdd.t31 vdd.t28 vdd.t30 vdd.t29 sky130_fd_pr__pfet_01v8 ad=3.51 pd=18.78 as=0 ps=0 w=9 l=0.5
X436 a_n3827_n3924.t6 plus.t24 a_n8300_8799.t12 gnd.t178 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.9
X437 a_n3827_n3924.t0 diffpairibias.t29 gnd.t1 gnd.t0 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=2.73 ps=14.78 w=7 l=1
X438 vdd.t27 vdd.t24 vdd.t26 vdd.t25 sky130_fd_pr__pfet_01v8 ad=3.51 pd=18.78 as=0 ps=0 w=9 l=0.5
X439 CSoutput.t3 a_n8300_8799.t115 vdd.t9 vdd.t8 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X440 CSoutput.t50 commonsourceibias.t197 gnd.t200 gnd.t199 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X441 CSoutput.t49 commonsourceibias.t198 gnd.t198 gnd.t197 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X442 a_n2982_13878.t34 a_n2982_13878.t33 a_n2804_13878.t6 vdd.t160 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X443 gnd.t192 commonsourceibias.t199 CSoutput.t48 gnd.t191 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
R0 commonsourceibias.n397 commonsourceibias.t184 222.032
R1 commonsourceibias.n281 commonsourceibias.t94 222.032
R2 commonsourceibias.n44 commonsourceibias.t76 222.032
R3 commonsourceibias.n166 commonsourceibias.t100 222.032
R4 commonsourceibias.n875 commonsourceibias.t196 222.032
R5 commonsourceibias.n759 commonsourceibias.t188 222.032
R6 commonsourceibias.n529 commonsourceibias.t22 222.032
R7 commonsourceibias.n645 commonsourceibias.t153 222.032
R8 commonsourceibias.n480 commonsourceibias.t183 207.983
R9 commonsourceibias.n364 commonsourceibias.t145 207.983
R10 commonsourceibias.n127 commonsourceibias.t72 207.983
R11 commonsourceibias.n249 commonsourceibias.t104 207.983
R12 commonsourceibias.n963 commonsourceibias.t93 207.983
R13 commonsourceibias.n847 commonsourceibias.t129 207.983
R14 commonsourceibias.n617 commonsourceibias.t36 207.983
R15 commonsourceibias.n732 commonsourceibias.t191 207.983
R16 commonsourceibias.n396 commonsourceibias.t151 168.701
R17 commonsourceibias.n402 commonsourceibias.t99 168.701
R18 commonsourceibias.n408 commonsourceibias.t81 168.701
R19 commonsourceibias.n392 commonsourceibias.t170 168.701
R20 commonsourceibias.n416 commonsourceibias.t177 168.701
R21 commonsourceibias.n422 commonsourceibias.t92 168.701
R22 commonsourceibias.n387 commonsourceibias.t186 168.701
R23 commonsourceibias.n430 commonsourceibias.t198 168.701
R24 commonsourceibias.n436 commonsourceibias.t130 168.701
R25 commonsourceibias.n382 commonsourceibias.t108 168.701
R26 commonsourceibias.n444 commonsourceibias.t88 168.701
R27 commonsourceibias.n450 commonsourceibias.t141 168.701
R28 commonsourceibias.n377 commonsourceibias.t150 168.701
R29 commonsourceibias.n458 commonsourceibias.t98 168.701
R30 commonsourceibias.n464 commonsourceibias.t199 168.701
R31 commonsourceibias.n372 commonsourceibias.t168 168.701
R32 commonsourceibias.n472 commonsourceibias.t107 168.701
R33 commonsourceibias.n478 commonsourceibias.t89 168.701
R34 commonsourceibias.n362 commonsourceibias.t172 168.701
R35 commonsourceibias.n356 commonsourceibias.t160 168.701
R36 commonsourceibias.n256 commonsourceibias.t146 168.701
R37 commonsourceibias.n348 commonsourceibias.t173 168.701
R38 commonsourceibias.n342 commonsourceibias.t158 168.701
R39 commonsourceibias.n261 commonsourceibias.t144 168.701
R40 commonsourceibias.n334 commonsourceibias.t174 168.701
R41 commonsourceibias.n328 commonsourceibias.t159 168.701
R42 commonsourceibias.n266 commonsourceibias.t185 168.701
R43 commonsourceibias.n320 commonsourceibias.t175 168.701
R44 commonsourceibias.n314 commonsourceibias.t157 168.701
R45 commonsourceibias.n271 commonsourceibias.t190 168.701
R46 commonsourceibias.n306 commonsourceibias.t91 168.701
R47 commonsourceibias.n300 commonsourceibias.t169 168.701
R48 commonsourceibias.n276 commonsourceibias.t82 168.701
R49 commonsourceibias.n292 commonsourceibias.t95 168.701
R50 commonsourceibias.n286 commonsourceibias.t90 168.701
R51 commonsourceibias.n280 commonsourceibias.t80 168.701
R52 commonsourceibias.n125 commonsourceibias.t42 168.701
R53 commonsourceibias.n119 commonsourceibias.t44 168.701
R54 commonsourceibias.n19 commonsourceibias.t6 168.701
R55 commonsourceibias.n111 commonsourceibias.t52 168.701
R56 commonsourceibias.n105 commonsourceibias.t74 168.701
R57 commonsourceibias.n24 commonsourceibias.t16 168.701
R58 commonsourceibias.n97 commonsourceibias.t50 168.701
R59 commonsourceibias.n91 commonsourceibias.t32 168.701
R60 commonsourceibias.n29 commonsourceibias.t56 168.701
R61 commonsourceibias.n83 commonsourceibias.t26 168.701
R62 commonsourceibias.n77 commonsourceibias.t20 168.701
R63 commonsourceibias.n34 commonsourceibias.t54 168.701
R64 commonsourceibias.n69 commonsourceibias.t68 168.701
R65 commonsourceibias.n63 commonsourceibias.t38 168.701
R66 commonsourceibias.n39 commonsourceibias.t14 168.701
R67 commonsourceibias.n55 commonsourceibias.t46 168.701
R68 commonsourceibias.n49 commonsourceibias.t2 168.701
R69 commonsourceibias.n43 commonsourceibias.t10 168.701
R70 commonsourceibias.n247 commonsourceibias.t181 168.701
R71 commonsourceibias.n241 commonsourceibias.t124 168.701
R72 commonsourceibias.n5 commonsourceibias.t197 168.701
R73 commonsourceibias.n233 commonsourceibias.t142 168.701
R74 commonsourceibias.n227 commonsourceibias.t101 168.701
R75 commonsourceibias.n10 commonsourceibias.t156 168.701
R76 commonsourceibias.n219 commonsourceibias.t143 168.701
R77 commonsourceibias.n213 commonsourceibias.t193 168.701
R78 commonsourceibias.n150 commonsourceibias.t136 168.701
R79 commonsourceibias.n151 commonsourceibias.t119 168.701
R80 commonsourceibias.n153 commonsourceibias.t155 168.701
R81 commonsourceibias.n155 commonsourceibias.t140 168.701
R82 commonsourceibias.n191 commonsourceibias.t109 168.701
R83 commonsourceibias.n185 commonsourceibias.t182 168.701
R84 commonsourceibias.n161 commonsourceibias.t166 168.701
R85 commonsourceibias.n177 commonsourceibias.t123 168.701
R86 commonsourceibias.n171 commonsourceibias.t84 168.701
R87 commonsourceibias.n165 commonsourceibias.t131 168.701
R88 commonsourceibias.n874 commonsourceibias.t165 168.701
R89 commonsourceibias.n880 commonsourceibias.t106 168.701
R90 commonsourceibias.n886 commonsourceibias.t87 168.701
R91 commonsourceibias.n888 commonsourceibias.t178 168.701
R92 commonsourceibias.n895 commonsourceibias.t167 168.701
R93 commonsourceibias.n901 commonsourceibias.t116 168.701
R94 commonsourceibias.n903 commonsourceibias.t96 168.701
R95 commonsourceibias.n910 commonsourceibias.t102 168.701
R96 commonsourceibias.n916 commonsourceibias.t121 168.701
R97 commonsourceibias.n918 commonsourceibias.t126 168.701
R98 commonsourceibias.n925 commonsourceibias.t112 168.701
R99 commonsourceibias.n931 commonsourceibias.t179 168.701
R100 commonsourceibias.n933 commonsourceibias.t133 168.701
R101 commonsourceibias.n940 commonsourceibias.t120 168.701
R102 commonsourceibias.n946 commonsourceibias.t103 168.701
R103 commonsourceibias.n948 commonsourceibias.t85 168.701
R104 commonsourceibias.n955 commonsourceibias.t125 168.701
R105 commonsourceibias.n961 commonsourceibias.t113 168.701
R106 commonsourceibias.n758 commonsourceibias.t163 168.701
R107 commonsourceibias.n764 commonsourceibias.t180 168.701
R108 commonsourceibias.n770 commonsourceibias.t189 168.701
R109 commonsourceibias.n772 commonsourceibias.t164 168.701
R110 commonsourceibias.n779 commonsourceibias.t176 168.701
R111 commonsourceibias.n785 commonsourceibias.t194 168.701
R112 commonsourceibias.n787 commonsourceibias.t171 168.701
R113 commonsourceibias.n794 commonsourceibias.t135 168.701
R114 commonsourceibias.n800 commonsourceibias.t195 168.701
R115 commonsourceibias.n802 commonsourceibias.t161 168.701
R116 commonsourceibias.n809 commonsourceibias.t137 168.701
R117 commonsourceibias.n815 commonsourceibias.t154 168.701
R118 commonsourceibias.n817 commonsourceibias.t162 168.701
R119 commonsourceibias.n824 commonsourceibias.t138 168.701
R120 commonsourceibias.n830 commonsourceibias.t147 168.701
R121 commonsourceibias.n832 commonsourceibias.t128 168.701
R122 commonsourceibias.n839 commonsourceibias.t139 168.701
R123 commonsourceibias.n845 commonsourceibias.t148 168.701
R124 commonsourceibias.n528 commonsourceibias.t0 168.701
R125 commonsourceibias.n534 commonsourceibias.t12 168.701
R126 commonsourceibias.n540 commonsourceibias.t34 168.701
R127 commonsourceibias.n542 commonsourceibias.t66 168.701
R128 commonsourceibias.n549 commonsourceibias.t64 168.701
R129 commonsourceibias.n555 commonsourceibias.t4 168.701
R130 commonsourceibias.n557 commonsourceibias.t60 168.701
R131 commonsourceibias.n564 commonsourceibias.t48 168.701
R132 commonsourceibias.n570 commonsourceibias.t70 168.701
R133 commonsourceibias.n572 commonsourceibias.t62 168.701
R134 commonsourceibias.n579 commonsourceibias.t24 168.701
R135 commonsourceibias.n585 commonsourceibias.t28 168.701
R136 commonsourceibias.n587 commonsourceibias.t8 168.701
R137 commonsourceibias.n594 commonsourceibias.t40 168.701
R138 commonsourceibias.n600 commonsourceibias.t30 168.701
R139 commonsourceibias.n602 commonsourceibias.t18 168.701
R140 commonsourceibias.n609 commonsourceibias.t78 168.701
R141 commonsourceibias.n615 commonsourceibias.t58 168.701
R142 commonsourceibias.n730 commonsourceibias.t134 168.701
R143 commonsourceibias.n724 commonsourceibias.t97 168.701
R144 commonsourceibias.n717 commonsourceibias.t152 168.701
R145 commonsourceibias.n715 commonsourceibias.t117 168.701
R146 commonsourceibias.n709 commonsourceibias.t187 168.701
R147 commonsourceibias.n702 commonsourceibias.t132 168.701
R148 commonsourceibias.n700 commonsourceibias.t118 168.701
R149 commonsourceibias.n694 commonsourceibias.t149 168.701
R150 commonsourceibias.n687 commonsourceibias.t114 168.701
R151 commonsourceibias.n644 commonsourceibias.t86 168.701
R152 commonsourceibias.n650 commonsourceibias.t127 168.701
R153 commonsourceibias.n656 commonsourceibias.t192 168.701
R154 commonsourceibias.n658 commonsourceibias.t110 168.701
R155 commonsourceibias.n665 commonsourceibias.t111 168.701
R156 commonsourceibias.n671 commonsourceibias.t83 168.701
R157 commonsourceibias.n635 commonsourceibias.t115 168.701
R158 commonsourceibias.n633 commonsourceibias.t122 168.701
R159 commonsourceibias.n631 commonsourceibias.t105 168.701
R160 commonsourceibias.n479 commonsourceibias.n367 161.3
R161 commonsourceibias.n477 commonsourceibias.n476 161.3
R162 commonsourceibias.n475 commonsourceibias.n368 161.3
R163 commonsourceibias.n474 commonsourceibias.n473 161.3
R164 commonsourceibias.n471 commonsourceibias.n369 161.3
R165 commonsourceibias.n470 commonsourceibias.n469 161.3
R166 commonsourceibias.n468 commonsourceibias.n370 161.3
R167 commonsourceibias.n467 commonsourceibias.n466 161.3
R168 commonsourceibias.n465 commonsourceibias.n371 161.3
R169 commonsourceibias.n463 commonsourceibias.n462 161.3
R170 commonsourceibias.n461 commonsourceibias.n373 161.3
R171 commonsourceibias.n460 commonsourceibias.n459 161.3
R172 commonsourceibias.n457 commonsourceibias.n374 161.3
R173 commonsourceibias.n456 commonsourceibias.n455 161.3
R174 commonsourceibias.n454 commonsourceibias.n375 161.3
R175 commonsourceibias.n453 commonsourceibias.n452 161.3
R176 commonsourceibias.n451 commonsourceibias.n376 161.3
R177 commonsourceibias.n449 commonsourceibias.n448 161.3
R178 commonsourceibias.n447 commonsourceibias.n378 161.3
R179 commonsourceibias.n446 commonsourceibias.n445 161.3
R180 commonsourceibias.n443 commonsourceibias.n379 161.3
R181 commonsourceibias.n442 commonsourceibias.n441 161.3
R182 commonsourceibias.n440 commonsourceibias.n380 161.3
R183 commonsourceibias.n439 commonsourceibias.n438 161.3
R184 commonsourceibias.n437 commonsourceibias.n381 161.3
R185 commonsourceibias.n435 commonsourceibias.n434 161.3
R186 commonsourceibias.n433 commonsourceibias.n383 161.3
R187 commonsourceibias.n432 commonsourceibias.n431 161.3
R188 commonsourceibias.n429 commonsourceibias.n384 161.3
R189 commonsourceibias.n428 commonsourceibias.n427 161.3
R190 commonsourceibias.n426 commonsourceibias.n385 161.3
R191 commonsourceibias.n425 commonsourceibias.n424 161.3
R192 commonsourceibias.n423 commonsourceibias.n386 161.3
R193 commonsourceibias.n421 commonsourceibias.n420 161.3
R194 commonsourceibias.n419 commonsourceibias.n388 161.3
R195 commonsourceibias.n418 commonsourceibias.n417 161.3
R196 commonsourceibias.n415 commonsourceibias.n389 161.3
R197 commonsourceibias.n414 commonsourceibias.n413 161.3
R198 commonsourceibias.n412 commonsourceibias.n390 161.3
R199 commonsourceibias.n411 commonsourceibias.n410 161.3
R200 commonsourceibias.n409 commonsourceibias.n391 161.3
R201 commonsourceibias.n407 commonsourceibias.n406 161.3
R202 commonsourceibias.n405 commonsourceibias.n393 161.3
R203 commonsourceibias.n404 commonsourceibias.n403 161.3
R204 commonsourceibias.n401 commonsourceibias.n394 161.3
R205 commonsourceibias.n400 commonsourceibias.n399 161.3
R206 commonsourceibias.n398 commonsourceibias.n395 161.3
R207 commonsourceibias.n282 commonsourceibias.n279 161.3
R208 commonsourceibias.n284 commonsourceibias.n283 161.3
R209 commonsourceibias.n285 commonsourceibias.n278 161.3
R210 commonsourceibias.n288 commonsourceibias.n287 161.3
R211 commonsourceibias.n289 commonsourceibias.n277 161.3
R212 commonsourceibias.n291 commonsourceibias.n290 161.3
R213 commonsourceibias.n293 commonsourceibias.n275 161.3
R214 commonsourceibias.n295 commonsourceibias.n294 161.3
R215 commonsourceibias.n296 commonsourceibias.n274 161.3
R216 commonsourceibias.n298 commonsourceibias.n297 161.3
R217 commonsourceibias.n299 commonsourceibias.n273 161.3
R218 commonsourceibias.n302 commonsourceibias.n301 161.3
R219 commonsourceibias.n303 commonsourceibias.n272 161.3
R220 commonsourceibias.n305 commonsourceibias.n304 161.3
R221 commonsourceibias.n307 commonsourceibias.n270 161.3
R222 commonsourceibias.n309 commonsourceibias.n308 161.3
R223 commonsourceibias.n310 commonsourceibias.n269 161.3
R224 commonsourceibias.n312 commonsourceibias.n311 161.3
R225 commonsourceibias.n313 commonsourceibias.n268 161.3
R226 commonsourceibias.n316 commonsourceibias.n315 161.3
R227 commonsourceibias.n317 commonsourceibias.n267 161.3
R228 commonsourceibias.n319 commonsourceibias.n318 161.3
R229 commonsourceibias.n321 commonsourceibias.n265 161.3
R230 commonsourceibias.n323 commonsourceibias.n322 161.3
R231 commonsourceibias.n324 commonsourceibias.n264 161.3
R232 commonsourceibias.n326 commonsourceibias.n325 161.3
R233 commonsourceibias.n327 commonsourceibias.n263 161.3
R234 commonsourceibias.n330 commonsourceibias.n329 161.3
R235 commonsourceibias.n331 commonsourceibias.n262 161.3
R236 commonsourceibias.n333 commonsourceibias.n332 161.3
R237 commonsourceibias.n335 commonsourceibias.n260 161.3
R238 commonsourceibias.n337 commonsourceibias.n336 161.3
R239 commonsourceibias.n338 commonsourceibias.n259 161.3
R240 commonsourceibias.n340 commonsourceibias.n339 161.3
R241 commonsourceibias.n341 commonsourceibias.n258 161.3
R242 commonsourceibias.n344 commonsourceibias.n343 161.3
R243 commonsourceibias.n345 commonsourceibias.n257 161.3
R244 commonsourceibias.n347 commonsourceibias.n346 161.3
R245 commonsourceibias.n349 commonsourceibias.n255 161.3
R246 commonsourceibias.n351 commonsourceibias.n350 161.3
R247 commonsourceibias.n352 commonsourceibias.n254 161.3
R248 commonsourceibias.n354 commonsourceibias.n353 161.3
R249 commonsourceibias.n355 commonsourceibias.n253 161.3
R250 commonsourceibias.n358 commonsourceibias.n357 161.3
R251 commonsourceibias.n359 commonsourceibias.n252 161.3
R252 commonsourceibias.n361 commonsourceibias.n360 161.3
R253 commonsourceibias.n363 commonsourceibias.n251 161.3
R254 commonsourceibias.n45 commonsourceibias.n42 161.3
R255 commonsourceibias.n47 commonsourceibias.n46 161.3
R256 commonsourceibias.n48 commonsourceibias.n41 161.3
R257 commonsourceibias.n51 commonsourceibias.n50 161.3
R258 commonsourceibias.n52 commonsourceibias.n40 161.3
R259 commonsourceibias.n54 commonsourceibias.n53 161.3
R260 commonsourceibias.n56 commonsourceibias.n38 161.3
R261 commonsourceibias.n58 commonsourceibias.n57 161.3
R262 commonsourceibias.n59 commonsourceibias.n37 161.3
R263 commonsourceibias.n61 commonsourceibias.n60 161.3
R264 commonsourceibias.n62 commonsourceibias.n36 161.3
R265 commonsourceibias.n65 commonsourceibias.n64 161.3
R266 commonsourceibias.n66 commonsourceibias.n35 161.3
R267 commonsourceibias.n68 commonsourceibias.n67 161.3
R268 commonsourceibias.n70 commonsourceibias.n33 161.3
R269 commonsourceibias.n72 commonsourceibias.n71 161.3
R270 commonsourceibias.n73 commonsourceibias.n32 161.3
R271 commonsourceibias.n75 commonsourceibias.n74 161.3
R272 commonsourceibias.n76 commonsourceibias.n31 161.3
R273 commonsourceibias.n79 commonsourceibias.n78 161.3
R274 commonsourceibias.n80 commonsourceibias.n30 161.3
R275 commonsourceibias.n82 commonsourceibias.n81 161.3
R276 commonsourceibias.n84 commonsourceibias.n28 161.3
R277 commonsourceibias.n86 commonsourceibias.n85 161.3
R278 commonsourceibias.n87 commonsourceibias.n27 161.3
R279 commonsourceibias.n89 commonsourceibias.n88 161.3
R280 commonsourceibias.n90 commonsourceibias.n26 161.3
R281 commonsourceibias.n93 commonsourceibias.n92 161.3
R282 commonsourceibias.n94 commonsourceibias.n25 161.3
R283 commonsourceibias.n96 commonsourceibias.n95 161.3
R284 commonsourceibias.n98 commonsourceibias.n23 161.3
R285 commonsourceibias.n100 commonsourceibias.n99 161.3
R286 commonsourceibias.n101 commonsourceibias.n22 161.3
R287 commonsourceibias.n103 commonsourceibias.n102 161.3
R288 commonsourceibias.n104 commonsourceibias.n21 161.3
R289 commonsourceibias.n107 commonsourceibias.n106 161.3
R290 commonsourceibias.n108 commonsourceibias.n20 161.3
R291 commonsourceibias.n110 commonsourceibias.n109 161.3
R292 commonsourceibias.n112 commonsourceibias.n18 161.3
R293 commonsourceibias.n114 commonsourceibias.n113 161.3
R294 commonsourceibias.n115 commonsourceibias.n17 161.3
R295 commonsourceibias.n117 commonsourceibias.n116 161.3
R296 commonsourceibias.n118 commonsourceibias.n16 161.3
R297 commonsourceibias.n121 commonsourceibias.n120 161.3
R298 commonsourceibias.n122 commonsourceibias.n15 161.3
R299 commonsourceibias.n124 commonsourceibias.n123 161.3
R300 commonsourceibias.n126 commonsourceibias.n14 161.3
R301 commonsourceibias.n167 commonsourceibias.n164 161.3
R302 commonsourceibias.n169 commonsourceibias.n168 161.3
R303 commonsourceibias.n170 commonsourceibias.n163 161.3
R304 commonsourceibias.n173 commonsourceibias.n172 161.3
R305 commonsourceibias.n174 commonsourceibias.n162 161.3
R306 commonsourceibias.n176 commonsourceibias.n175 161.3
R307 commonsourceibias.n178 commonsourceibias.n160 161.3
R308 commonsourceibias.n180 commonsourceibias.n179 161.3
R309 commonsourceibias.n181 commonsourceibias.n159 161.3
R310 commonsourceibias.n183 commonsourceibias.n182 161.3
R311 commonsourceibias.n184 commonsourceibias.n158 161.3
R312 commonsourceibias.n187 commonsourceibias.n186 161.3
R313 commonsourceibias.n188 commonsourceibias.n157 161.3
R314 commonsourceibias.n190 commonsourceibias.n189 161.3
R315 commonsourceibias.n192 commonsourceibias.n156 161.3
R316 commonsourceibias.n194 commonsourceibias.n193 161.3
R317 commonsourceibias.n196 commonsourceibias.n195 161.3
R318 commonsourceibias.n197 commonsourceibias.n154 161.3
R319 commonsourceibias.n199 commonsourceibias.n198 161.3
R320 commonsourceibias.n201 commonsourceibias.n200 161.3
R321 commonsourceibias.n202 commonsourceibias.n152 161.3
R322 commonsourceibias.n204 commonsourceibias.n203 161.3
R323 commonsourceibias.n206 commonsourceibias.n205 161.3
R324 commonsourceibias.n208 commonsourceibias.n207 161.3
R325 commonsourceibias.n209 commonsourceibias.n13 161.3
R326 commonsourceibias.n211 commonsourceibias.n210 161.3
R327 commonsourceibias.n212 commonsourceibias.n12 161.3
R328 commonsourceibias.n215 commonsourceibias.n214 161.3
R329 commonsourceibias.n216 commonsourceibias.n11 161.3
R330 commonsourceibias.n218 commonsourceibias.n217 161.3
R331 commonsourceibias.n220 commonsourceibias.n9 161.3
R332 commonsourceibias.n222 commonsourceibias.n221 161.3
R333 commonsourceibias.n223 commonsourceibias.n8 161.3
R334 commonsourceibias.n225 commonsourceibias.n224 161.3
R335 commonsourceibias.n226 commonsourceibias.n7 161.3
R336 commonsourceibias.n229 commonsourceibias.n228 161.3
R337 commonsourceibias.n230 commonsourceibias.n6 161.3
R338 commonsourceibias.n232 commonsourceibias.n231 161.3
R339 commonsourceibias.n234 commonsourceibias.n4 161.3
R340 commonsourceibias.n236 commonsourceibias.n235 161.3
R341 commonsourceibias.n237 commonsourceibias.n3 161.3
R342 commonsourceibias.n239 commonsourceibias.n238 161.3
R343 commonsourceibias.n240 commonsourceibias.n2 161.3
R344 commonsourceibias.n243 commonsourceibias.n242 161.3
R345 commonsourceibias.n244 commonsourceibias.n1 161.3
R346 commonsourceibias.n246 commonsourceibias.n245 161.3
R347 commonsourceibias.n248 commonsourceibias.n0 161.3
R348 commonsourceibias.n962 commonsourceibias.n850 161.3
R349 commonsourceibias.n960 commonsourceibias.n959 161.3
R350 commonsourceibias.n958 commonsourceibias.n851 161.3
R351 commonsourceibias.n957 commonsourceibias.n956 161.3
R352 commonsourceibias.n954 commonsourceibias.n852 161.3
R353 commonsourceibias.n953 commonsourceibias.n952 161.3
R354 commonsourceibias.n951 commonsourceibias.n853 161.3
R355 commonsourceibias.n950 commonsourceibias.n949 161.3
R356 commonsourceibias.n947 commonsourceibias.n854 161.3
R357 commonsourceibias.n945 commonsourceibias.n944 161.3
R358 commonsourceibias.n943 commonsourceibias.n855 161.3
R359 commonsourceibias.n942 commonsourceibias.n941 161.3
R360 commonsourceibias.n939 commonsourceibias.n856 161.3
R361 commonsourceibias.n938 commonsourceibias.n937 161.3
R362 commonsourceibias.n936 commonsourceibias.n857 161.3
R363 commonsourceibias.n935 commonsourceibias.n934 161.3
R364 commonsourceibias.n932 commonsourceibias.n858 161.3
R365 commonsourceibias.n930 commonsourceibias.n929 161.3
R366 commonsourceibias.n928 commonsourceibias.n859 161.3
R367 commonsourceibias.n927 commonsourceibias.n926 161.3
R368 commonsourceibias.n924 commonsourceibias.n860 161.3
R369 commonsourceibias.n923 commonsourceibias.n922 161.3
R370 commonsourceibias.n921 commonsourceibias.n861 161.3
R371 commonsourceibias.n920 commonsourceibias.n919 161.3
R372 commonsourceibias.n917 commonsourceibias.n862 161.3
R373 commonsourceibias.n915 commonsourceibias.n914 161.3
R374 commonsourceibias.n913 commonsourceibias.n863 161.3
R375 commonsourceibias.n912 commonsourceibias.n911 161.3
R376 commonsourceibias.n909 commonsourceibias.n864 161.3
R377 commonsourceibias.n908 commonsourceibias.n907 161.3
R378 commonsourceibias.n906 commonsourceibias.n865 161.3
R379 commonsourceibias.n905 commonsourceibias.n904 161.3
R380 commonsourceibias.n902 commonsourceibias.n866 161.3
R381 commonsourceibias.n900 commonsourceibias.n899 161.3
R382 commonsourceibias.n898 commonsourceibias.n867 161.3
R383 commonsourceibias.n897 commonsourceibias.n896 161.3
R384 commonsourceibias.n894 commonsourceibias.n868 161.3
R385 commonsourceibias.n893 commonsourceibias.n892 161.3
R386 commonsourceibias.n891 commonsourceibias.n869 161.3
R387 commonsourceibias.n890 commonsourceibias.n889 161.3
R388 commonsourceibias.n887 commonsourceibias.n870 161.3
R389 commonsourceibias.n885 commonsourceibias.n884 161.3
R390 commonsourceibias.n883 commonsourceibias.n871 161.3
R391 commonsourceibias.n882 commonsourceibias.n881 161.3
R392 commonsourceibias.n879 commonsourceibias.n872 161.3
R393 commonsourceibias.n878 commonsourceibias.n877 161.3
R394 commonsourceibias.n876 commonsourceibias.n873 161.3
R395 commonsourceibias.n846 commonsourceibias.n734 161.3
R396 commonsourceibias.n844 commonsourceibias.n843 161.3
R397 commonsourceibias.n842 commonsourceibias.n735 161.3
R398 commonsourceibias.n841 commonsourceibias.n840 161.3
R399 commonsourceibias.n838 commonsourceibias.n736 161.3
R400 commonsourceibias.n837 commonsourceibias.n836 161.3
R401 commonsourceibias.n835 commonsourceibias.n737 161.3
R402 commonsourceibias.n834 commonsourceibias.n833 161.3
R403 commonsourceibias.n831 commonsourceibias.n738 161.3
R404 commonsourceibias.n829 commonsourceibias.n828 161.3
R405 commonsourceibias.n827 commonsourceibias.n739 161.3
R406 commonsourceibias.n826 commonsourceibias.n825 161.3
R407 commonsourceibias.n823 commonsourceibias.n740 161.3
R408 commonsourceibias.n822 commonsourceibias.n821 161.3
R409 commonsourceibias.n820 commonsourceibias.n741 161.3
R410 commonsourceibias.n819 commonsourceibias.n818 161.3
R411 commonsourceibias.n816 commonsourceibias.n742 161.3
R412 commonsourceibias.n814 commonsourceibias.n813 161.3
R413 commonsourceibias.n812 commonsourceibias.n743 161.3
R414 commonsourceibias.n811 commonsourceibias.n810 161.3
R415 commonsourceibias.n808 commonsourceibias.n744 161.3
R416 commonsourceibias.n807 commonsourceibias.n806 161.3
R417 commonsourceibias.n805 commonsourceibias.n745 161.3
R418 commonsourceibias.n804 commonsourceibias.n803 161.3
R419 commonsourceibias.n801 commonsourceibias.n746 161.3
R420 commonsourceibias.n799 commonsourceibias.n798 161.3
R421 commonsourceibias.n797 commonsourceibias.n747 161.3
R422 commonsourceibias.n796 commonsourceibias.n795 161.3
R423 commonsourceibias.n793 commonsourceibias.n748 161.3
R424 commonsourceibias.n792 commonsourceibias.n791 161.3
R425 commonsourceibias.n790 commonsourceibias.n749 161.3
R426 commonsourceibias.n789 commonsourceibias.n788 161.3
R427 commonsourceibias.n786 commonsourceibias.n750 161.3
R428 commonsourceibias.n784 commonsourceibias.n783 161.3
R429 commonsourceibias.n782 commonsourceibias.n751 161.3
R430 commonsourceibias.n781 commonsourceibias.n780 161.3
R431 commonsourceibias.n778 commonsourceibias.n752 161.3
R432 commonsourceibias.n777 commonsourceibias.n776 161.3
R433 commonsourceibias.n775 commonsourceibias.n753 161.3
R434 commonsourceibias.n774 commonsourceibias.n773 161.3
R435 commonsourceibias.n771 commonsourceibias.n754 161.3
R436 commonsourceibias.n769 commonsourceibias.n768 161.3
R437 commonsourceibias.n767 commonsourceibias.n755 161.3
R438 commonsourceibias.n766 commonsourceibias.n765 161.3
R439 commonsourceibias.n763 commonsourceibias.n756 161.3
R440 commonsourceibias.n762 commonsourceibias.n761 161.3
R441 commonsourceibias.n760 commonsourceibias.n757 161.3
R442 commonsourceibias.n616 commonsourceibias.n504 161.3
R443 commonsourceibias.n614 commonsourceibias.n613 161.3
R444 commonsourceibias.n612 commonsourceibias.n505 161.3
R445 commonsourceibias.n611 commonsourceibias.n610 161.3
R446 commonsourceibias.n608 commonsourceibias.n506 161.3
R447 commonsourceibias.n607 commonsourceibias.n606 161.3
R448 commonsourceibias.n605 commonsourceibias.n507 161.3
R449 commonsourceibias.n604 commonsourceibias.n603 161.3
R450 commonsourceibias.n601 commonsourceibias.n508 161.3
R451 commonsourceibias.n599 commonsourceibias.n598 161.3
R452 commonsourceibias.n597 commonsourceibias.n509 161.3
R453 commonsourceibias.n596 commonsourceibias.n595 161.3
R454 commonsourceibias.n593 commonsourceibias.n510 161.3
R455 commonsourceibias.n592 commonsourceibias.n591 161.3
R456 commonsourceibias.n590 commonsourceibias.n511 161.3
R457 commonsourceibias.n589 commonsourceibias.n588 161.3
R458 commonsourceibias.n586 commonsourceibias.n512 161.3
R459 commonsourceibias.n584 commonsourceibias.n583 161.3
R460 commonsourceibias.n582 commonsourceibias.n513 161.3
R461 commonsourceibias.n581 commonsourceibias.n580 161.3
R462 commonsourceibias.n578 commonsourceibias.n514 161.3
R463 commonsourceibias.n577 commonsourceibias.n576 161.3
R464 commonsourceibias.n575 commonsourceibias.n515 161.3
R465 commonsourceibias.n574 commonsourceibias.n573 161.3
R466 commonsourceibias.n571 commonsourceibias.n516 161.3
R467 commonsourceibias.n569 commonsourceibias.n568 161.3
R468 commonsourceibias.n567 commonsourceibias.n517 161.3
R469 commonsourceibias.n566 commonsourceibias.n565 161.3
R470 commonsourceibias.n563 commonsourceibias.n518 161.3
R471 commonsourceibias.n562 commonsourceibias.n561 161.3
R472 commonsourceibias.n560 commonsourceibias.n519 161.3
R473 commonsourceibias.n559 commonsourceibias.n558 161.3
R474 commonsourceibias.n556 commonsourceibias.n520 161.3
R475 commonsourceibias.n554 commonsourceibias.n553 161.3
R476 commonsourceibias.n552 commonsourceibias.n521 161.3
R477 commonsourceibias.n551 commonsourceibias.n550 161.3
R478 commonsourceibias.n548 commonsourceibias.n522 161.3
R479 commonsourceibias.n547 commonsourceibias.n546 161.3
R480 commonsourceibias.n545 commonsourceibias.n523 161.3
R481 commonsourceibias.n544 commonsourceibias.n543 161.3
R482 commonsourceibias.n541 commonsourceibias.n524 161.3
R483 commonsourceibias.n539 commonsourceibias.n538 161.3
R484 commonsourceibias.n537 commonsourceibias.n525 161.3
R485 commonsourceibias.n536 commonsourceibias.n535 161.3
R486 commonsourceibias.n533 commonsourceibias.n526 161.3
R487 commonsourceibias.n532 commonsourceibias.n531 161.3
R488 commonsourceibias.n530 commonsourceibias.n527 161.3
R489 commonsourceibias.n686 commonsourceibias.n685 161.3
R490 commonsourceibias.n684 commonsourceibias.n683 161.3
R491 commonsourceibias.n682 commonsourceibias.n632 161.3
R492 commonsourceibias.n681 commonsourceibias.n680 161.3
R493 commonsourceibias.n679 commonsourceibias.n678 161.3
R494 commonsourceibias.n677 commonsourceibias.n634 161.3
R495 commonsourceibias.n676 commonsourceibias.n675 161.3
R496 commonsourceibias.n674 commonsourceibias.n673 161.3
R497 commonsourceibias.n672 commonsourceibias.n636 161.3
R498 commonsourceibias.n670 commonsourceibias.n669 161.3
R499 commonsourceibias.n668 commonsourceibias.n637 161.3
R500 commonsourceibias.n667 commonsourceibias.n666 161.3
R501 commonsourceibias.n664 commonsourceibias.n638 161.3
R502 commonsourceibias.n663 commonsourceibias.n662 161.3
R503 commonsourceibias.n661 commonsourceibias.n639 161.3
R504 commonsourceibias.n660 commonsourceibias.n659 161.3
R505 commonsourceibias.n657 commonsourceibias.n640 161.3
R506 commonsourceibias.n655 commonsourceibias.n654 161.3
R507 commonsourceibias.n653 commonsourceibias.n641 161.3
R508 commonsourceibias.n652 commonsourceibias.n651 161.3
R509 commonsourceibias.n649 commonsourceibias.n642 161.3
R510 commonsourceibias.n648 commonsourceibias.n647 161.3
R511 commonsourceibias.n646 commonsourceibias.n643 161.3
R512 commonsourceibias.n731 commonsourceibias.n483 161.3
R513 commonsourceibias.n729 commonsourceibias.n728 161.3
R514 commonsourceibias.n727 commonsourceibias.n484 161.3
R515 commonsourceibias.n726 commonsourceibias.n725 161.3
R516 commonsourceibias.n723 commonsourceibias.n485 161.3
R517 commonsourceibias.n722 commonsourceibias.n721 161.3
R518 commonsourceibias.n720 commonsourceibias.n486 161.3
R519 commonsourceibias.n719 commonsourceibias.n718 161.3
R520 commonsourceibias.n716 commonsourceibias.n487 161.3
R521 commonsourceibias.n714 commonsourceibias.n713 161.3
R522 commonsourceibias.n712 commonsourceibias.n488 161.3
R523 commonsourceibias.n711 commonsourceibias.n710 161.3
R524 commonsourceibias.n708 commonsourceibias.n489 161.3
R525 commonsourceibias.n707 commonsourceibias.n706 161.3
R526 commonsourceibias.n705 commonsourceibias.n490 161.3
R527 commonsourceibias.n704 commonsourceibias.n703 161.3
R528 commonsourceibias.n701 commonsourceibias.n491 161.3
R529 commonsourceibias.n699 commonsourceibias.n698 161.3
R530 commonsourceibias.n697 commonsourceibias.n492 161.3
R531 commonsourceibias.n696 commonsourceibias.n695 161.3
R532 commonsourceibias.n693 commonsourceibias.n493 161.3
R533 commonsourceibias.n692 commonsourceibias.n691 161.3
R534 commonsourceibias.n690 commonsourceibias.n494 161.3
R535 commonsourceibias.n689 commonsourceibias.n688 161.3
R536 commonsourceibias.n141 commonsourceibias.n139 81.5057
R537 commonsourceibias.n497 commonsourceibias.n495 81.5057
R538 commonsourceibias.n141 commonsourceibias.n140 80.9324
R539 commonsourceibias.n143 commonsourceibias.n142 80.9324
R540 commonsourceibias.n145 commonsourceibias.n144 80.9324
R541 commonsourceibias.n147 commonsourceibias.n146 80.9324
R542 commonsourceibias.n138 commonsourceibias.n137 80.9324
R543 commonsourceibias.n136 commonsourceibias.n135 80.9324
R544 commonsourceibias.n134 commonsourceibias.n133 80.9324
R545 commonsourceibias.n132 commonsourceibias.n131 80.9324
R546 commonsourceibias.n130 commonsourceibias.n129 80.9324
R547 commonsourceibias.n620 commonsourceibias.n619 80.9324
R548 commonsourceibias.n622 commonsourceibias.n621 80.9324
R549 commonsourceibias.n624 commonsourceibias.n623 80.9324
R550 commonsourceibias.n626 commonsourceibias.n625 80.9324
R551 commonsourceibias.n628 commonsourceibias.n627 80.9324
R552 commonsourceibias.n503 commonsourceibias.n502 80.9324
R553 commonsourceibias.n501 commonsourceibias.n500 80.9324
R554 commonsourceibias.n499 commonsourceibias.n498 80.9324
R555 commonsourceibias.n497 commonsourceibias.n496 80.9324
R556 commonsourceibias.n481 commonsourceibias.n480 80.6037
R557 commonsourceibias.n365 commonsourceibias.n364 80.6037
R558 commonsourceibias.n128 commonsourceibias.n127 80.6037
R559 commonsourceibias.n250 commonsourceibias.n249 80.6037
R560 commonsourceibias.n964 commonsourceibias.n963 80.6037
R561 commonsourceibias.n848 commonsourceibias.n847 80.6037
R562 commonsourceibias.n618 commonsourceibias.n617 80.6037
R563 commonsourceibias.n733 commonsourceibias.n732 80.6037
R564 commonsourceibias.n438 commonsourceibias.n437 56.5617
R565 commonsourceibias.n452 commonsourceibias.n451 56.5617
R566 commonsourceibias.n322 commonsourceibias.n321 56.5617
R567 commonsourceibias.n308 commonsourceibias.n307 56.5617
R568 commonsourceibias.n85 commonsourceibias.n84 56.5617
R569 commonsourceibias.n71 commonsourceibias.n70 56.5617
R570 commonsourceibias.n207 commonsourceibias.n206 56.5617
R571 commonsourceibias.n193 commonsourceibias.n192 56.5617
R572 commonsourceibias.n919 commonsourceibias.n917 56.5617
R573 commonsourceibias.n934 commonsourceibias.n932 56.5617
R574 commonsourceibias.n803 commonsourceibias.n801 56.5617
R575 commonsourceibias.n818 commonsourceibias.n816 56.5617
R576 commonsourceibias.n573 commonsourceibias.n571 56.5617
R577 commonsourceibias.n588 commonsourceibias.n586 56.5617
R578 commonsourceibias.n688 commonsourceibias.n686 56.5617
R579 commonsourceibias.n410 commonsourceibias.n409 56.5617
R580 commonsourceibias.n424 commonsourceibias.n423 56.5617
R581 commonsourceibias.n466 commonsourceibias.n465 56.5617
R582 commonsourceibias.n350 commonsourceibias.n349 56.5617
R583 commonsourceibias.n336 commonsourceibias.n335 56.5617
R584 commonsourceibias.n294 commonsourceibias.n293 56.5617
R585 commonsourceibias.n113 commonsourceibias.n112 56.5617
R586 commonsourceibias.n99 commonsourceibias.n98 56.5617
R587 commonsourceibias.n57 commonsourceibias.n56 56.5617
R588 commonsourceibias.n235 commonsourceibias.n234 56.5617
R589 commonsourceibias.n221 commonsourceibias.n220 56.5617
R590 commonsourceibias.n179 commonsourceibias.n178 56.5617
R591 commonsourceibias.n889 commonsourceibias.n887 56.5617
R592 commonsourceibias.n904 commonsourceibias.n902 56.5617
R593 commonsourceibias.n949 commonsourceibias.n947 56.5617
R594 commonsourceibias.n773 commonsourceibias.n771 56.5617
R595 commonsourceibias.n788 commonsourceibias.n786 56.5617
R596 commonsourceibias.n833 commonsourceibias.n831 56.5617
R597 commonsourceibias.n543 commonsourceibias.n541 56.5617
R598 commonsourceibias.n558 commonsourceibias.n556 56.5617
R599 commonsourceibias.n603 commonsourceibias.n601 56.5617
R600 commonsourceibias.n718 commonsourceibias.n716 56.5617
R601 commonsourceibias.n703 commonsourceibias.n701 56.5617
R602 commonsourceibias.n659 commonsourceibias.n657 56.5617
R603 commonsourceibias.n673 commonsourceibias.n672 56.5617
R604 commonsourceibias.n401 commonsourceibias.n400 51.2335
R605 commonsourceibias.n473 commonsourceibias.n368 51.2335
R606 commonsourceibias.n357 commonsourceibias.n252 51.2335
R607 commonsourceibias.n285 commonsourceibias.n284 51.2335
R608 commonsourceibias.n120 commonsourceibias.n15 51.2335
R609 commonsourceibias.n48 commonsourceibias.n47 51.2335
R610 commonsourceibias.n242 commonsourceibias.n1 51.2335
R611 commonsourceibias.n170 commonsourceibias.n169 51.2335
R612 commonsourceibias.n879 commonsourceibias.n878 51.2335
R613 commonsourceibias.n956 commonsourceibias.n851 51.2335
R614 commonsourceibias.n763 commonsourceibias.n762 51.2335
R615 commonsourceibias.n840 commonsourceibias.n735 51.2335
R616 commonsourceibias.n533 commonsourceibias.n532 51.2335
R617 commonsourceibias.n610 commonsourceibias.n505 51.2335
R618 commonsourceibias.n725 commonsourceibias.n484 51.2335
R619 commonsourceibias.n649 commonsourceibias.n648 51.2335
R620 commonsourceibias.n480 commonsourceibias.n479 50.9056
R621 commonsourceibias.n364 commonsourceibias.n363 50.9056
R622 commonsourceibias.n127 commonsourceibias.n126 50.9056
R623 commonsourceibias.n249 commonsourceibias.n248 50.9056
R624 commonsourceibias.n963 commonsourceibias.n962 50.9056
R625 commonsourceibias.n847 commonsourceibias.n846 50.9056
R626 commonsourceibias.n617 commonsourceibias.n616 50.9056
R627 commonsourceibias.n732 commonsourceibias.n731 50.9056
R628 commonsourceibias.n415 commonsourceibias.n414 50.2647
R629 commonsourceibias.n459 commonsourceibias.n373 50.2647
R630 commonsourceibias.n343 commonsourceibias.n257 50.2647
R631 commonsourceibias.n299 commonsourceibias.n298 50.2647
R632 commonsourceibias.n106 commonsourceibias.n20 50.2647
R633 commonsourceibias.n62 commonsourceibias.n61 50.2647
R634 commonsourceibias.n228 commonsourceibias.n6 50.2647
R635 commonsourceibias.n184 commonsourceibias.n183 50.2647
R636 commonsourceibias.n894 commonsourceibias.n893 50.2647
R637 commonsourceibias.n941 commonsourceibias.n855 50.2647
R638 commonsourceibias.n778 commonsourceibias.n777 50.2647
R639 commonsourceibias.n825 commonsourceibias.n739 50.2647
R640 commonsourceibias.n548 commonsourceibias.n547 50.2647
R641 commonsourceibias.n595 commonsourceibias.n509 50.2647
R642 commonsourceibias.n710 commonsourceibias.n488 50.2647
R643 commonsourceibias.n664 commonsourceibias.n663 50.2647
R644 commonsourceibias.n397 commonsourceibias.n396 49.9027
R645 commonsourceibias.n281 commonsourceibias.n280 49.9027
R646 commonsourceibias.n44 commonsourceibias.n43 49.9027
R647 commonsourceibias.n166 commonsourceibias.n165 49.9027
R648 commonsourceibias.n875 commonsourceibias.n874 49.9027
R649 commonsourceibias.n759 commonsourceibias.n758 49.9027
R650 commonsourceibias.n529 commonsourceibias.n528 49.9027
R651 commonsourceibias.n645 commonsourceibias.n644 49.9027
R652 commonsourceibias.n429 commonsourceibias.n428 49.296
R653 commonsourceibias.n445 commonsourceibias.n378 49.296
R654 commonsourceibias.n329 commonsourceibias.n262 49.296
R655 commonsourceibias.n313 commonsourceibias.n312 49.296
R656 commonsourceibias.n92 commonsourceibias.n25 49.296
R657 commonsourceibias.n76 commonsourceibias.n75 49.296
R658 commonsourceibias.n214 commonsourceibias.n11 49.296
R659 commonsourceibias.n198 commonsourceibias.n197 49.296
R660 commonsourceibias.n909 commonsourceibias.n908 49.296
R661 commonsourceibias.n926 commonsourceibias.n859 49.296
R662 commonsourceibias.n793 commonsourceibias.n792 49.296
R663 commonsourceibias.n810 commonsourceibias.n743 49.296
R664 commonsourceibias.n563 commonsourceibias.n562 49.296
R665 commonsourceibias.n580 commonsourceibias.n513 49.296
R666 commonsourceibias.n695 commonsourceibias.n492 49.296
R667 commonsourceibias.n678 commonsourceibias.n677 49.296
R668 commonsourceibias.n431 commonsourceibias.n383 48.3272
R669 commonsourceibias.n443 commonsourceibias.n442 48.3272
R670 commonsourceibias.n327 commonsourceibias.n326 48.3272
R671 commonsourceibias.n315 commonsourceibias.n267 48.3272
R672 commonsourceibias.n90 commonsourceibias.n89 48.3272
R673 commonsourceibias.n78 commonsourceibias.n30 48.3272
R674 commonsourceibias.n212 commonsourceibias.n211 48.3272
R675 commonsourceibias.n202 commonsourceibias.n201 48.3272
R676 commonsourceibias.n911 commonsourceibias.n863 48.3272
R677 commonsourceibias.n924 commonsourceibias.n923 48.3272
R678 commonsourceibias.n795 commonsourceibias.n747 48.3272
R679 commonsourceibias.n808 commonsourceibias.n807 48.3272
R680 commonsourceibias.n565 commonsourceibias.n517 48.3272
R681 commonsourceibias.n578 commonsourceibias.n577 48.3272
R682 commonsourceibias.n693 commonsourceibias.n692 48.3272
R683 commonsourceibias.n682 commonsourceibias.n681 48.3272
R684 commonsourceibias.n417 commonsourceibias.n388 47.3584
R685 commonsourceibias.n457 commonsourceibias.n456 47.3584
R686 commonsourceibias.n341 commonsourceibias.n340 47.3584
R687 commonsourceibias.n301 commonsourceibias.n272 47.3584
R688 commonsourceibias.n104 commonsourceibias.n103 47.3584
R689 commonsourceibias.n64 commonsourceibias.n35 47.3584
R690 commonsourceibias.n226 commonsourceibias.n225 47.3584
R691 commonsourceibias.n186 commonsourceibias.n157 47.3584
R692 commonsourceibias.n896 commonsourceibias.n867 47.3584
R693 commonsourceibias.n939 commonsourceibias.n938 47.3584
R694 commonsourceibias.n780 commonsourceibias.n751 47.3584
R695 commonsourceibias.n823 commonsourceibias.n822 47.3584
R696 commonsourceibias.n550 commonsourceibias.n521 47.3584
R697 commonsourceibias.n593 commonsourceibias.n592 47.3584
R698 commonsourceibias.n708 commonsourceibias.n707 47.3584
R699 commonsourceibias.n666 commonsourceibias.n637 47.3584
R700 commonsourceibias.n403 commonsourceibias.n393 46.3896
R701 commonsourceibias.n471 commonsourceibias.n470 46.3896
R702 commonsourceibias.n355 commonsourceibias.n354 46.3896
R703 commonsourceibias.n287 commonsourceibias.n277 46.3896
R704 commonsourceibias.n118 commonsourceibias.n117 46.3896
R705 commonsourceibias.n50 commonsourceibias.n40 46.3896
R706 commonsourceibias.n240 commonsourceibias.n239 46.3896
R707 commonsourceibias.n172 commonsourceibias.n162 46.3896
R708 commonsourceibias.n881 commonsourceibias.n871 46.3896
R709 commonsourceibias.n954 commonsourceibias.n953 46.3896
R710 commonsourceibias.n765 commonsourceibias.n755 46.3896
R711 commonsourceibias.n838 commonsourceibias.n837 46.3896
R712 commonsourceibias.n535 commonsourceibias.n525 46.3896
R713 commonsourceibias.n608 commonsourceibias.n607 46.3896
R714 commonsourceibias.n723 commonsourceibias.n722 46.3896
R715 commonsourceibias.n651 commonsourceibias.n641 46.3896
R716 commonsourceibias.n398 commonsourceibias.n397 44.7059
R717 commonsourceibias.n876 commonsourceibias.n875 44.7059
R718 commonsourceibias.n760 commonsourceibias.n759 44.7059
R719 commonsourceibias.n530 commonsourceibias.n529 44.7059
R720 commonsourceibias.n646 commonsourceibias.n645 44.7059
R721 commonsourceibias.n282 commonsourceibias.n281 44.7059
R722 commonsourceibias.n45 commonsourceibias.n44 44.7059
R723 commonsourceibias.n167 commonsourceibias.n166 44.7059
R724 commonsourceibias.n407 commonsourceibias.n393 34.7644
R725 commonsourceibias.n470 commonsourceibias.n370 34.7644
R726 commonsourceibias.n354 commonsourceibias.n254 34.7644
R727 commonsourceibias.n291 commonsourceibias.n277 34.7644
R728 commonsourceibias.n117 commonsourceibias.n17 34.7644
R729 commonsourceibias.n54 commonsourceibias.n40 34.7644
R730 commonsourceibias.n239 commonsourceibias.n3 34.7644
R731 commonsourceibias.n176 commonsourceibias.n162 34.7644
R732 commonsourceibias.n885 commonsourceibias.n871 34.7644
R733 commonsourceibias.n953 commonsourceibias.n853 34.7644
R734 commonsourceibias.n769 commonsourceibias.n755 34.7644
R735 commonsourceibias.n837 commonsourceibias.n737 34.7644
R736 commonsourceibias.n539 commonsourceibias.n525 34.7644
R737 commonsourceibias.n607 commonsourceibias.n507 34.7644
R738 commonsourceibias.n722 commonsourceibias.n486 34.7644
R739 commonsourceibias.n655 commonsourceibias.n641 34.7644
R740 commonsourceibias.n421 commonsourceibias.n388 33.7956
R741 commonsourceibias.n456 commonsourceibias.n375 33.7956
R742 commonsourceibias.n340 commonsourceibias.n259 33.7956
R743 commonsourceibias.n305 commonsourceibias.n272 33.7956
R744 commonsourceibias.n103 commonsourceibias.n22 33.7956
R745 commonsourceibias.n68 commonsourceibias.n35 33.7956
R746 commonsourceibias.n225 commonsourceibias.n8 33.7956
R747 commonsourceibias.n190 commonsourceibias.n157 33.7956
R748 commonsourceibias.n900 commonsourceibias.n867 33.7956
R749 commonsourceibias.n938 commonsourceibias.n857 33.7956
R750 commonsourceibias.n784 commonsourceibias.n751 33.7956
R751 commonsourceibias.n822 commonsourceibias.n741 33.7956
R752 commonsourceibias.n554 commonsourceibias.n521 33.7956
R753 commonsourceibias.n592 commonsourceibias.n511 33.7956
R754 commonsourceibias.n707 commonsourceibias.n490 33.7956
R755 commonsourceibias.n670 commonsourceibias.n637 33.7956
R756 commonsourceibias.n435 commonsourceibias.n383 32.8269
R757 commonsourceibias.n442 commonsourceibias.n380 32.8269
R758 commonsourceibias.n326 commonsourceibias.n264 32.8269
R759 commonsourceibias.n319 commonsourceibias.n267 32.8269
R760 commonsourceibias.n89 commonsourceibias.n27 32.8269
R761 commonsourceibias.n82 commonsourceibias.n30 32.8269
R762 commonsourceibias.n211 commonsourceibias.n13 32.8269
R763 commonsourceibias.n203 commonsourceibias.n202 32.8269
R764 commonsourceibias.n915 commonsourceibias.n863 32.8269
R765 commonsourceibias.n923 commonsourceibias.n861 32.8269
R766 commonsourceibias.n799 commonsourceibias.n747 32.8269
R767 commonsourceibias.n807 commonsourceibias.n745 32.8269
R768 commonsourceibias.n569 commonsourceibias.n517 32.8269
R769 commonsourceibias.n577 commonsourceibias.n515 32.8269
R770 commonsourceibias.n692 commonsourceibias.n494 32.8269
R771 commonsourceibias.n683 commonsourceibias.n682 32.8269
R772 commonsourceibias.n428 commonsourceibias.n385 31.8581
R773 commonsourceibias.n449 commonsourceibias.n378 31.8581
R774 commonsourceibias.n333 commonsourceibias.n262 31.8581
R775 commonsourceibias.n312 commonsourceibias.n269 31.8581
R776 commonsourceibias.n96 commonsourceibias.n25 31.8581
R777 commonsourceibias.n75 commonsourceibias.n32 31.8581
R778 commonsourceibias.n218 commonsourceibias.n11 31.8581
R779 commonsourceibias.n197 commonsourceibias.n196 31.8581
R780 commonsourceibias.n908 commonsourceibias.n865 31.8581
R781 commonsourceibias.n930 commonsourceibias.n859 31.8581
R782 commonsourceibias.n792 commonsourceibias.n749 31.8581
R783 commonsourceibias.n814 commonsourceibias.n743 31.8581
R784 commonsourceibias.n562 commonsourceibias.n519 31.8581
R785 commonsourceibias.n584 commonsourceibias.n513 31.8581
R786 commonsourceibias.n699 commonsourceibias.n492 31.8581
R787 commonsourceibias.n677 commonsourceibias.n676 31.8581
R788 commonsourceibias.n414 commonsourceibias.n390 30.8893
R789 commonsourceibias.n463 commonsourceibias.n373 30.8893
R790 commonsourceibias.n347 commonsourceibias.n257 30.8893
R791 commonsourceibias.n298 commonsourceibias.n274 30.8893
R792 commonsourceibias.n110 commonsourceibias.n20 30.8893
R793 commonsourceibias.n61 commonsourceibias.n37 30.8893
R794 commonsourceibias.n232 commonsourceibias.n6 30.8893
R795 commonsourceibias.n183 commonsourceibias.n159 30.8893
R796 commonsourceibias.n893 commonsourceibias.n869 30.8893
R797 commonsourceibias.n945 commonsourceibias.n855 30.8893
R798 commonsourceibias.n777 commonsourceibias.n753 30.8893
R799 commonsourceibias.n829 commonsourceibias.n739 30.8893
R800 commonsourceibias.n547 commonsourceibias.n523 30.8893
R801 commonsourceibias.n599 commonsourceibias.n509 30.8893
R802 commonsourceibias.n714 commonsourceibias.n488 30.8893
R803 commonsourceibias.n663 commonsourceibias.n639 30.8893
R804 commonsourceibias.n400 commonsourceibias.n395 29.9206
R805 commonsourceibias.n477 commonsourceibias.n368 29.9206
R806 commonsourceibias.n361 commonsourceibias.n252 29.9206
R807 commonsourceibias.n284 commonsourceibias.n279 29.9206
R808 commonsourceibias.n124 commonsourceibias.n15 29.9206
R809 commonsourceibias.n47 commonsourceibias.n42 29.9206
R810 commonsourceibias.n246 commonsourceibias.n1 29.9206
R811 commonsourceibias.n169 commonsourceibias.n164 29.9206
R812 commonsourceibias.n878 commonsourceibias.n873 29.9206
R813 commonsourceibias.n960 commonsourceibias.n851 29.9206
R814 commonsourceibias.n762 commonsourceibias.n757 29.9206
R815 commonsourceibias.n844 commonsourceibias.n735 29.9206
R816 commonsourceibias.n532 commonsourceibias.n527 29.9206
R817 commonsourceibias.n614 commonsourceibias.n505 29.9206
R818 commonsourceibias.n729 commonsourceibias.n484 29.9206
R819 commonsourceibias.n648 commonsourceibias.n643 29.9206
R820 commonsourceibias.n479 commonsourceibias.n478 21.8872
R821 commonsourceibias.n363 commonsourceibias.n362 21.8872
R822 commonsourceibias.n126 commonsourceibias.n125 21.8872
R823 commonsourceibias.n248 commonsourceibias.n247 21.8872
R824 commonsourceibias.n962 commonsourceibias.n961 21.8872
R825 commonsourceibias.n846 commonsourceibias.n845 21.8872
R826 commonsourceibias.n616 commonsourceibias.n615 21.8872
R827 commonsourceibias.n731 commonsourceibias.n730 21.8872
R828 commonsourceibias.n410 commonsourceibias.n392 21.3954
R829 commonsourceibias.n465 commonsourceibias.n464 21.3954
R830 commonsourceibias.n349 commonsourceibias.n348 21.3954
R831 commonsourceibias.n294 commonsourceibias.n276 21.3954
R832 commonsourceibias.n112 commonsourceibias.n111 21.3954
R833 commonsourceibias.n57 commonsourceibias.n39 21.3954
R834 commonsourceibias.n234 commonsourceibias.n233 21.3954
R835 commonsourceibias.n179 commonsourceibias.n161 21.3954
R836 commonsourceibias.n889 commonsourceibias.n888 21.3954
R837 commonsourceibias.n947 commonsourceibias.n946 21.3954
R838 commonsourceibias.n773 commonsourceibias.n772 21.3954
R839 commonsourceibias.n831 commonsourceibias.n830 21.3954
R840 commonsourceibias.n543 commonsourceibias.n542 21.3954
R841 commonsourceibias.n601 commonsourceibias.n600 21.3954
R842 commonsourceibias.n716 commonsourceibias.n715 21.3954
R843 commonsourceibias.n659 commonsourceibias.n658 21.3954
R844 commonsourceibias.n424 commonsourceibias.n387 20.9036
R845 commonsourceibias.n451 commonsourceibias.n450 20.9036
R846 commonsourceibias.n335 commonsourceibias.n334 20.9036
R847 commonsourceibias.n308 commonsourceibias.n271 20.9036
R848 commonsourceibias.n98 commonsourceibias.n97 20.9036
R849 commonsourceibias.n71 commonsourceibias.n34 20.9036
R850 commonsourceibias.n220 commonsourceibias.n219 20.9036
R851 commonsourceibias.n193 commonsourceibias.n155 20.9036
R852 commonsourceibias.n904 commonsourceibias.n903 20.9036
R853 commonsourceibias.n932 commonsourceibias.n931 20.9036
R854 commonsourceibias.n788 commonsourceibias.n787 20.9036
R855 commonsourceibias.n816 commonsourceibias.n815 20.9036
R856 commonsourceibias.n558 commonsourceibias.n557 20.9036
R857 commonsourceibias.n586 commonsourceibias.n585 20.9036
R858 commonsourceibias.n701 commonsourceibias.n700 20.9036
R859 commonsourceibias.n673 commonsourceibias.n635 20.9036
R860 commonsourceibias.n437 commonsourceibias.n436 20.4117
R861 commonsourceibias.n438 commonsourceibias.n382 20.4117
R862 commonsourceibias.n322 commonsourceibias.n266 20.4117
R863 commonsourceibias.n321 commonsourceibias.n320 20.4117
R864 commonsourceibias.n85 commonsourceibias.n29 20.4117
R865 commonsourceibias.n84 commonsourceibias.n83 20.4117
R866 commonsourceibias.n207 commonsourceibias.n150 20.4117
R867 commonsourceibias.n206 commonsourceibias.n151 20.4117
R868 commonsourceibias.n917 commonsourceibias.n916 20.4117
R869 commonsourceibias.n919 commonsourceibias.n918 20.4117
R870 commonsourceibias.n801 commonsourceibias.n800 20.4117
R871 commonsourceibias.n803 commonsourceibias.n802 20.4117
R872 commonsourceibias.n571 commonsourceibias.n570 20.4117
R873 commonsourceibias.n573 commonsourceibias.n572 20.4117
R874 commonsourceibias.n688 commonsourceibias.n687 20.4117
R875 commonsourceibias.n686 commonsourceibias.n631 20.4117
R876 commonsourceibias.n423 commonsourceibias.n422 19.9199
R877 commonsourceibias.n452 commonsourceibias.n377 19.9199
R878 commonsourceibias.n336 commonsourceibias.n261 19.9199
R879 commonsourceibias.n307 commonsourceibias.n306 19.9199
R880 commonsourceibias.n99 commonsourceibias.n24 19.9199
R881 commonsourceibias.n70 commonsourceibias.n69 19.9199
R882 commonsourceibias.n221 commonsourceibias.n10 19.9199
R883 commonsourceibias.n192 commonsourceibias.n191 19.9199
R884 commonsourceibias.n902 commonsourceibias.n901 19.9199
R885 commonsourceibias.n934 commonsourceibias.n933 19.9199
R886 commonsourceibias.n786 commonsourceibias.n785 19.9199
R887 commonsourceibias.n818 commonsourceibias.n817 19.9199
R888 commonsourceibias.n556 commonsourceibias.n555 19.9199
R889 commonsourceibias.n588 commonsourceibias.n587 19.9199
R890 commonsourceibias.n703 commonsourceibias.n702 19.9199
R891 commonsourceibias.n672 commonsourceibias.n671 19.9199
R892 commonsourceibias.n409 commonsourceibias.n408 19.4281
R893 commonsourceibias.n466 commonsourceibias.n372 19.4281
R894 commonsourceibias.n350 commonsourceibias.n256 19.4281
R895 commonsourceibias.n293 commonsourceibias.n292 19.4281
R896 commonsourceibias.n113 commonsourceibias.n19 19.4281
R897 commonsourceibias.n56 commonsourceibias.n55 19.4281
R898 commonsourceibias.n235 commonsourceibias.n5 19.4281
R899 commonsourceibias.n178 commonsourceibias.n177 19.4281
R900 commonsourceibias.n887 commonsourceibias.n886 19.4281
R901 commonsourceibias.n949 commonsourceibias.n948 19.4281
R902 commonsourceibias.n771 commonsourceibias.n770 19.4281
R903 commonsourceibias.n833 commonsourceibias.n832 19.4281
R904 commonsourceibias.n541 commonsourceibias.n540 19.4281
R905 commonsourceibias.n603 commonsourceibias.n602 19.4281
R906 commonsourceibias.n718 commonsourceibias.n717 19.4281
R907 commonsourceibias.n657 commonsourceibias.n656 19.4281
R908 commonsourceibias.n402 commonsourceibias.n401 13.526
R909 commonsourceibias.n473 commonsourceibias.n472 13.526
R910 commonsourceibias.n357 commonsourceibias.n356 13.526
R911 commonsourceibias.n286 commonsourceibias.n285 13.526
R912 commonsourceibias.n120 commonsourceibias.n119 13.526
R913 commonsourceibias.n49 commonsourceibias.n48 13.526
R914 commonsourceibias.n242 commonsourceibias.n241 13.526
R915 commonsourceibias.n171 commonsourceibias.n170 13.526
R916 commonsourceibias.n880 commonsourceibias.n879 13.526
R917 commonsourceibias.n956 commonsourceibias.n955 13.526
R918 commonsourceibias.n764 commonsourceibias.n763 13.526
R919 commonsourceibias.n840 commonsourceibias.n839 13.526
R920 commonsourceibias.n534 commonsourceibias.n533 13.526
R921 commonsourceibias.n610 commonsourceibias.n609 13.526
R922 commonsourceibias.n725 commonsourceibias.n724 13.526
R923 commonsourceibias.n650 commonsourceibias.n649 13.526
R924 commonsourceibias.n130 commonsourceibias.n128 13.2322
R925 commonsourceibias.n620 commonsourceibias.n618 13.2322
R926 commonsourceibias.n416 commonsourceibias.n415 13.0342
R927 commonsourceibias.n459 commonsourceibias.n458 13.0342
R928 commonsourceibias.n343 commonsourceibias.n342 13.0342
R929 commonsourceibias.n300 commonsourceibias.n299 13.0342
R930 commonsourceibias.n106 commonsourceibias.n105 13.0342
R931 commonsourceibias.n63 commonsourceibias.n62 13.0342
R932 commonsourceibias.n228 commonsourceibias.n227 13.0342
R933 commonsourceibias.n185 commonsourceibias.n184 13.0342
R934 commonsourceibias.n895 commonsourceibias.n894 13.0342
R935 commonsourceibias.n941 commonsourceibias.n940 13.0342
R936 commonsourceibias.n779 commonsourceibias.n778 13.0342
R937 commonsourceibias.n825 commonsourceibias.n824 13.0342
R938 commonsourceibias.n549 commonsourceibias.n548 13.0342
R939 commonsourceibias.n595 commonsourceibias.n594 13.0342
R940 commonsourceibias.n710 commonsourceibias.n709 13.0342
R941 commonsourceibias.n665 commonsourceibias.n664 13.0342
R942 commonsourceibias.n430 commonsourceibias.n429 12.5423
R943 commonsourceibias.n445 commonsourceibias.n444 12.5423
R944 commonsourceibias.n329 commonsourceibias.n328 12.5423
R945 commonsourceibias.n314 commonsourceibias.n313 12.5423
R946 commonsourceibias.n92 commonsourceibias.n91 12.5423
R947 commonsourceibias.n77 commonsourceibias.n76 12.5423
R948 commonsourceibias.n214 commonsourceibias.n213 12.5423
R949 commonsourceibias.n198 commonsourceibias.n153 12.5423
R950 commonsourceibias.n910 commonsourceibias.n909 12.5423
R951 commonsourceibias.n926 commonsourceibias.n925 12.5423
R952 commonsourceibias.n794 commonsourceibias.n793 12.5423
R953 commonsourceibias.n810 commonsourceibias.n809 12.5423
R954 commonsourceibias.n564 commonsourceibias.n563 12.5423
R955 commonsourceibias.n580 commonsourceibias.n579 12.5423
R956 commonsourceibias.n695 commonsourceibias.n694 12.5423
R957 commonsourceibias.n678 commonsourceibias.n633 12.5423
R958 commonsourceibias.n431 commonsourceibias.n430 12.0505
R959 commonsourceibias.n444 commonsourceibias.n443 12.0505
R960 commonsourceibias.n328 commonsourceibias.n327 12.0505
R961 commonsourceibias.n315 commonsourceibias.n314 12.0505
R962 commonsourceibias.n91 commonsourceibias.n90 12.0505
R963 commonsourceibias.n78 commonsourceibias.n77 12.0505
R964 commonsourceibias.n213 commonsourceibias.n212 12.0505
R965 commonsourceibias.n201 commonsourceibias.n153 12.0505
R966 commonsourceibias.n911 commonsourceibias.n910 12.0505
R967 commonsourceibias.n925 commonsourceibias.n924 12.0505
R968 commonsourceibias.n795 commonsourceibias.n794 12.0505
R969 commonsourceibias.n809 commonsourceibias.n808 12.0505
R970 commonsourceibias.n565 commonsourceibias.n564 12.0505
R971 commonsourceibias.n579 commonsourceibias.n578 12.0505
R972 commonsourceibias.n694 commonsourceibias.n693 12.0505
R973 commonsourceibias.n681 commonsourceibias.n633 12.0505
R974 commonsourceibias.n417 commonsourceibias.n416 11.5587
R975 commonsourceibias.n458 commonsourceibias.n457 11.5587
R976 commonsourceibias.n342 commonsourceibias.n341 11.5587
R977 commonsourceibias.n301 commonsourceibias.n300 11.5587
R978 commonsourceibias.n105 commonsourceibias.n104 11.5587
R979 commonsourceibias.n64 commonsourceibias.n63 11.5587
R980 commonsourceibias.n227 commonsourceibias.n226 11.5587
R981 commonsourceibias.n186 commonsourceibias.n185 11.5587
R982 commonsourceibias.n896 commonsourceibias.n895 11.5587
R983 commonsourceibias.n940 commonsourceibias.n939 11.5587
R984 commonsourceibias.n780 commonsourceibias.n779 11.5587
R985 commonsourceibias.n824 commonsourceibias.n823 11.5587
R986 commonsourceibias.n550 commonsourceibias.n549 11.5587
R987 commonsourceibias.n594 commonsourceibias.n593 11.5587
R988 commonsourceibias.n709 commonsourceibias.n708 11.5587
R989 commonsourceibias.n666 commonsourceibias.n665 11.5587
R990 commonsourceibias.n403 commonsourceibias.n402 11.0668
R991 commonsourceibias.n472 commonsourceibias.n471 11.0668
R992 commonsourceibias.n356 commonsourceibias.n355 11.0668
R993 commonsourceibias.n287 commonsourceibias.n286 11.0668
R994 commonsourceibias.n119 commonsourceibias.n118 11.0668
R995 commonsourceibias.n50 commonsourceibias.n49 11.0668
R996 commonsourceibias.n241 commonsourceibias.n240 11.0668
R997 commonsourceibias.n172 commonsourceibias.n171 11.0668
R998 commonsourceibias.n881 commonsourceibias.n880 11.0668
R999 commonsourceibias.n955 commonsourceibias.n954 11.0668
R1000 commonsourceibias.n765 commonsourceibias.n764 11.0668
R1001 commonsourceibias.n839 commonsourceibias.n838 11.0668
R1002 commonsourceibias.n535 commonsourceibias.n534 11.0668
R1003 commonsourceibias.n609 commonsourceibias.n608 11.0668
R1004 commonsourceibias.n724 commonsourceibias.n723 11.0668
R1005 commonsourceibias.n651 commonsourceibias.n650 11.0668
R1006 commonsourceibias.n966 commonsourceibias.n482 10.4122
R1007 commonsourceibias.n149 commonsourceibias.n148 9.50363
R1008 commonsourceibias.n630 commonsourceibias.n629 9.50363
R1009 commonsourceibias.n366 commonsourceibias.n250 8.76042
R1010 commonsourceibias.n849 commonsourceibias.n733 8.76042
R1011 commonsourceibias.n966 commonsourceibias.n965 8.46921
R1012 commonsourceibias.n408 commonsourceibias.n407 5.16479
R1013 commonsourceibias.n372 commonsourceibias.n370 5.16479
R1014 commonsourceibias.n256 commonsourceibias.n254 5.16479
R1015 commonsourceibias.n292 commonsourceibias.n291 5.16479
R1016 commonsourceibias.n19 commonsourceibias.n17 5.16479
R1017 commonsourceibias.n55 commonsourceibias.n54 5.16479
R1018 commonsourceibias.n5 commonsourceibias.n3 5.16479
R1019 commonsourceibias.n177 commonsourceibias.n176 5.16479
R1020 commonsourceibias.n886 commonsourceibias.n885 5.16479
R1021 commonsourceibias.n948 commonsourceibias.n853 5.16479
R1022 commonsourceibias.n770 commonsourceibias.n769 5.16479
R1023 commonsourceibias.n832 commonsourceibias.n737 5.16479
R1024 commonsourceibias.n540 commonsourceibias.n539 5.16479
R1025 commonsourceibias.n602 commonsourceibias.n507 5.16479
R1026 commonsourceibias.n717 commonsourceibias.n486 5.16479
R1027 commonsourceibias.n656 commonsourceibias.n655 5.16479
R1028 commonsourceibias.n482 commonsourceibias.n481 5.03125
R1029 commonsourceibias.n366 commonsourceibias.n365 5.03125
R1030 commonsourceibias.n965 commonsourceibias.n964 5.03125
R1031 commonsourceibias.n849 commonsourceibias.n848 5.03125
R1032 commonsourceibias.n422 commonsourceibias.n421 4.67295
R1033 commonsourceibias.n377 commonsourceibias.n375 4.67295
R1034 commonsourceibias.n261 commonsourceibias.n259 4.67295
R1035 commonsourceibias.n306 commonsourceibias.n305 4.67295
R1036 commonsourceibias.n24 commonsourceibias.n22 4.67295
R1037 commonsourceibias.n69 commonsourceibias.n68 4.67295
R1038 commonsourceibias.n10 commonsourceibias.n8 4.67295
R1039 commonsourceibias.n191 commonsourceibias.n190 4.67295
R1040 commonsourceibias.n901 commonsourceibias.n900 4.67295
R1041 commonsourceibias.n933 commonsourceibias.n857 4.67295
R1042 commonsourceibias.n785 commonsourceibias.n784 4.67295
R1043 commonsourceibias.n817 commonsourceibias.n741 4.67295
R1044 commonsourceibias.n555 commonsourceibias.n554 4.67295
R1045 commonsourceibias.n587 commonsourceibias.n511 4.67295
R1046 commonsourceibias.n702 commonsourceibias.n490 4.67295
R1047 commonsourceibias.n671 commonsourceibias.n670 4.67295
R1048 commonsourceibias commonsourceibias.n966 4.20978
R1049 commonsourceibias.n436 commonsourceibias.n435 4.18111
R1050 commonsourceibias.n382 commonsourceibias.n380 4.18111
R1051 commonsourceibias.n266 commonsourceibias.n264 4.18111
R1052 commonsourceibias.n320 commonsourceibias.n319 4.18111
R1053 commonsourceibias.n29 commonsourceibias.n27 4.18111
R1054 commonsourceibias.n83 commonsourceibias.n82 4.18111
R1055 commonsourceibias.n150 commonsourceibias.n13 4.18111
R1056 commonsourceibias.n203 commonsourceibias.n151 4.18111
R1057 commonsourceibias.n916 commonsourceibias.n915 4.18111
R1058 commonsourceibias.n918 commonsourceibias.n861 4.18111
R1059 commonsourceibias.n800 commonsourceibias.n799 4.18111
R1060 commonsourceibias.n802 commonsourceibias.n745 4.18111
R1061 commonsourceibias.n570 commonsourceibias.n569 4.18111
R1062 commonsourceibias.n572 commonsourceibias.n515 4.18111
R1063 commonsourceibias.n687 commonsourceibias.n494 4.18111
R1064 commonsourceibias.n683 commonsourceibias.n631 4.18111
R1065 commonsourceibias.n482 commonsourceibias.n366 3.72967
R1066 commonsourceibias.n965 commonsourceibias.n849 3.72967
R1067 commonsourceibias.n387 commonsourceibias.n385 3.68928
R1068 commonsourceibias.n450 commonsourceibias.n449 3.68928
R1069 commonsourceibias.n334 commonsourceibias.n333 3.68928
R1070 commonsourceibias.n271 commonsourceibias.n269 3.68928
R1071 commonsourceibias.n97 commonsourceibias.n96 3.68928
R1072 commonsourceibias.n34 commonsourceibias.n32 3.68928
R1073 commonsourceibias.n219 commonsourceibias.n218 3.68928
R1074 commonsourceibias.n196 commonsourceibias.n155 3.68928
R1075 commonsourceibias.n903 commonsourceibias.n865 3.68928
R1076 commonsourceibias.n931 commonsourceibias.n930 3.68928
R1077 commonsourceibias.n787 commonsourceibias.n749 3.68928
R1078 commonsourceibias.n815 commonsourceibias.n814 3.68928
R1079 commonsourceibias.n557 commonsourceibias.n519 3.68928
R1080 commonsourceibias.n585 commonsourceibias.n584 3.68928
R1081 commonsourceibias.n700 commonsourceibias.n699 3.68928
R1082 commonsourceibias.n676 commonsourceibias.n635 3.68928
R1083 commonsourceibias.n392 commonsourceibias.n390 3.19744
R1084 commonsourceibias.n464 commonsourceibias.n463 3.19744
R1085 commonsourceibias.n348 commonsourceibias.n347 3.19744
R1086 commonsourceibias.n276 commonsourceibias.n274 3.19744
R1087 commonsourceibias.n111 commonsourceibias.n110 3.19744
R1088 commonsourceibias.n39 commonsourceibias.n37 3.19744
R1089 commonsourceibias.n233 commonsourceibias.n232 3.19744
R1090 commonsourceibias.n161 commonsourceibias.n159 3.19744
R1091 commonsourceibias.n888 commonsourceibias.n869 3.19744
R1092 commonsourceibias.n946 commonsourceibias.n945 3.19744
R1093 commonsourceibias.n772 commonsourceibias.n753 3.19744
R1094 commonsourceibias.n830 commonsourceibias.n829 3.19744
R1095 commonsourceibias.n542 commonsourceibias.n523 3.19744
R1096 commonsourceibias.n600 commonsourceibias.n599 3.19744
R1097 commonsourceibias.n715 commonsourceibias.n714 3.19744
R1098 commonsourceibias.n658 commonsourceibias.n639 3.19744
R1099 commonsourceibias.n139 commonsourceibias.t11 2.82907
R1100 commonsourceibias.n139 commonsourceibias.t77 2.82907
R1101 commonsourceibias.n140 commonsourceibias.t47 2.82907
R1102 commonsourceibias.n140 commonsourceibias.t3 2.82907
R1103 commonsourceibias.n142 commonsourceibias.t39 2.82907
R1104 commonsourceibias.n142 commonsourceibias.t15 2.82907
R1105 commonsourceibias.n144 commonsourceibias.t55 2.82907
R1106 commonsourceibias.n144 commonsourceibias.t69 2.82907
R1107 commonsourceibias.n146 commonsourceibias.t27 2.82907
R1108 commonsourceibias.n146 commonsourceibias.t21 2.82907
R1109 commonsourceibias.n137 commonsourceibias.t33 2.82907
R1110 commonsourceibias.n137 commonsourceibias.t57 2.82907
R1111 commonsourceibias.n135 commonsourceibias.t17 2.82907
R1112 commonsourceibias.n135 commonsourceibias.t51 2.82907
R1113 commonsourceibias.n133 commonsourceibias.t53 2.82907
R1114 commonsourceibias.n133 commonsourceibias.t75 2.82907
R1115 commonsourceibias.n131 commonsourceibias.t45 2.82907
R1116 commonsourceibias.n131 commonsourceibias.t7 2.82907
R1117 commonsourceibias.n129 commonsourceibias.t73 2.82907
R1118 commonsourceibias.n129 commonsourceibias.t43 2.82907
R1119 commonsourceibias.n619 commonsourceibias.t59 2.82907
R1120 commonsourceibias.n619 commonsourceibias.t37 2.82907
R1121 commonsourceibias.n621 commonsourceibias.t19 2.82907
R1122 commonsourceibias.n621 commonsourceibias.t79 2.82907
R1123 commonsourceibias.n623 commonsourceibias.t41 2.82907
R1124 commonsourceibias.n623 commonsourceibias.t31 2.82907
R1125 commonsourceibias.n625 commonsourceibias.t29 2.82907
R1126 commonsourceibias.n625 commonsourceibias.t9 2.82907
R1127 commonsourceibias.n627 commonsourceibias.t63 2.82907
R1128 commonsourceibias.n627 commonsourceibias.t25 2.82907
R1129 commonsourceibias.n502 commonsourceibias.t49 2.82907
R1130 commonsourceibias.n502 commonsourceibias.t71 2.82907
R1131 commonsourceibias.n500 commonsourceibias.t5 2.82907
R1132 commonsourceibias.n500 commonsourceibias.t61 2.82907
R1133 commonsourceibias.n498 commonsourceibias.t67 2.82907
R1134 commonsourceibias.n498 commonsourceibias.t65 2.82907
R1135 commonsourceibias.n496 commonsourceibias.t13 2.82907
R1136 commonsourceibias.n496 commonsourceibias.t35 2.82907
R1137 commonsourceibias.n495 commonsourceibias.t23 2.82907
R1138 commonsourceibias.n495 commonsourceibias.t1 2.82907
R1139 commonsourceibias.n396 commonsourceibias.n395 2.7056
R1140 commonsourceibias.n478 commonsourceibias.n477 2.7056
R1141 commonsourceibias.n362 commonsourceibias.n361 2.7056
R1142 commonsourceibias.n280 commonsourceibias.n279 2.7056
R1143 commonsourceibias.n125 commonsourceibias.n124 2.7056
R1144 commonsourceibias.n43 commonsourceibias.n42 2.7056
R1145 commonsourceibias.n247 commonsourceibias.n246 2.7056
R1146 commonsourceibias.n165 commonsourceibias.n164 2.7056
R1147 commonsourceibias.n874 commonsourceibias.n873 2.7056
R1148 commonsourceibias.n961 commonsourceibias.n960 2.7056
R1149 commonsourceibias.n758 commonsourceibias.n757 2.7056
R1150 commonsourceibias.n845 commonsourceibias.n844 2.7056
R1151 commonsourceibias.n528 commonsourceibias.n527 2.7056
R1152 commonsourceibias.n615 commonsourceibias.n614 2.7056
R1153 commonsourceibias.n730 commonsourceibias.n729 2.7056
R1154 commonsourceibias.n644 commonsourceibias.n643 2.7056
R1155 commonsourceibias.n132 commonsourceibias.n130 0.573776
R1156 commonsourceibias.n134 commonsourceibias.n132 0.573776
R1157 commonsourceibias.n136 commonsourceibias.n134 0.573776
R1158 commonsourceibias.n138 commonsourceibias.n136 0.573776
R1159 commonsourceibias.n147 commonsourceibias.n145 0.573776
R1160 commonsourceibias.n145 commonsourceibias.n143 0.573776
R1161 commonsourceibias.n143 commonsourceibias.n141 0.573776
R1162 commonsourceibias.n499 commonsourceibias.n497 0.573776
R1163 commonsourceibias.n501 commonsourceibias.n499 0.573776
R1164 commonsourceibias.n503 commonsourceibias.n501 0.573776
R1165 commonsourceibias.n628 commonsourceibias.n626 0.573776
R1166 commonsourceibias.n626 commonsourceibias.n624 0.573776
R1167 commonsourceibias.n624 commonsourceibias.n622 0.573776
R1168 commonsourceibias.n622 commonsourceibias.n620 0.573776
R1169 commonsourceibias.n148 commonsourceibias.n138 0.287138
R1170 commonsourceibias.n148 commonsourceibias.n147 0.287138
R1171 commonsourceibias.n629 commonsourceibias.n503 0.287138
R1172 commonsourceibias.n629 commonsourceibias.n628 0.287138
R1173 commonsourceibias.n481 commonsourceibias.n367 0.285035
R1174 commonsourceibias.n365 commonsourceibias.n251 0.285035
R1175 commonsourceibias.n128 commonsourceibias.n14 0.285035
R1176 commonsourceibias.n250 commonsourceibias.n0 0.285035
R1177 commonsourceibias.n964 commonsourceibias.n850 0.285035
R1178 commonsourceibias.n848 commonsourceibias.n734 0.285035
R1179 commonsourceibias.n618 commonsourceibias.n504 0.285035
R1180 commonsourceibias.n733 commonsourceibias.n483 0.285035
R1181 commonsourceibias.n476 commonsourceibias.n367 0.189894
R1182 commonsourceibias.n476 commonsourceibias.n475 0.189894
R1183 commonsourceibias.n475 commonsourceibias.n474 0.189894
R1184 commonsourceibias.n474 commonsourceibias.n369 0.189894
R1185 commonsourceibias.n469 commonsourceibias.n369 0.189894
R1186 commonsourceibias.n469 commonsourceibias.n468 0.189894
R1187 commonsourceibias.n468 commonsourceibias.n467 0.189894
R1188 commonsourceibias.n467 commonsourceibias.n371 0.189894
R1189 commonsourceibias.n462 commonsourceibias.n371 0.189894
R1190 commonsourceibias.n462 commonsourceibias.n461 0.189894
R1191 commonsourceibias.n461 commonsourceibias.n460 0.189894
R1192 commonsourceibias.n460 commonsourceibias.n374 0.189894
R1193 commonsourceibias.n455 commonsourceibias.n374 0.189894
R1194 commonsourceibias.n455 commonsourceibias.n454 0.189894
R1195 commonsourceibias.n454 commonsourceibias.n453 0.189894
R1196 commonsourceibias.n453 commonsourceibias.n376 0.189894
R1197 commonsourceibias.n448 commonsourceibias.n376 0.189894
R1198 commonsourceibias.n448 commonsourceibias.n447 0.189894
R1199 commonsourceibias.n447 commonsourceibias.n446 0.189894
R1200 commonsourceibias.n446 commonsourceibias.n379 0.189894
R1201 commonsourceibias.n441 commonsourceibias.n379 0.189894
R1202 commonsourceibias.n441 commonsourceibias.n440 0.189894
R1203 commonsourceibias.n440 commonsourceibias.n439 0.189894
R1204 commonsourceibias.n439 commonsourceibias.n381 0.189894
R1205 commonsourceibias.n434 commonsourceibias.n381 0.189894
R1206 commonsourceibias.n434 commonsourceibias.n433 0.189894
R1207 commonsourceibias.n433 commonsourceibias.n432 0.189894
R1208 commonsourceibias.n432 commonsourceibias.n384 0.189894
R1209 commonsourceibias.n427 commonsourceibias.n384 0.189894
R1210 commonsourceibias.n427 commonsourceibias.n426 0.189894
R1211 commonsourceibias.n426 commonsourceibias.n425 0.189894
R1212 commonsourceibias.n425 commonsourceibias.n386 0.189894
R1213 commonsourceibias.n420 commonsourceibias.n386 0.189894
R1214 commonsourceibias.n420 commonsourceibias.n419 0.189894
R1215 commonsourceibias.n419 commonsourceibias.n418 0.189894
R1216 commonsourceibias.n418 commonsourceibias.n389 0.189894
R1217 commonsourceibias.n413 commonsourceibias.n389 0.189894
R1218 commonsourceibias.n413 commonsourceibias.n412 0.189894
R1219 commonsourceibias.n412 commonsourceibias.n411 0.189894
R1220 commonsourceibias.n411 commonsourceibias.n391 0.189894
R1221 commonsourceibias.n406 commonsourceibias.n391 0.189894
R1222 commonsourceibias.n406 commonsourceibias.n405 0.189894
R1223 commonsourceibias.n405 commonsourceibias.n404 0.189894
R1224 commonsourceibias.n404 commonsourceibias.n394 0.189894
R1225 commonsourceibias.n399 commonsourceibias.n394 0.189894
R1226 commonsourceibias.n399 commonsourceibias.n398 0.189894
R1227 commonsourceibias.n360 commonsourceibias.n251 0.189894
R1228 commonsourceibias.n360 commonsourceibias.n359 0.189894
R1229 commonsourceibias.n359 commonsourceibias.n358 0.189894
R1230 commonsourceibias.n358 commonsourceibias.n253 0.189894
R1231 commonsourceibias.n353 commonsourceibias.n253 0.189894
R1232 commonsourceibias.n353 commonsourceibias.n352 0.189894
R1233 commonsourceibias.n352 commonsourceibias.n351 0.189894
R1234 commonsourceibias.n351 commonsourceibias.n255 0.189894
R1235 commonsourceibias.n346 commonsourceibias.n255 0.189894
R1236 commonsourceibias.n346 commonsourceibias.n345 0.189894
R1237 commonsourceibias.n345 commonsourceibias.n344 0.189894
R1238 commonsourceibias.n344 commonsourceibias.n258 0.189894
R1239 commonsourceibias.n339 commonsourceibias.n258 0.189894
R1240 commonsourceibias.n339 commonsourceibias.n338 0.189894
R1241 commonsourceibias.n338 commonsourceibias.n337 0.189894
R1242 commonsourceibias.n337 commonsourceibias.n260 0.189894
R1243 commonsourceibias.n332 commonsourceibias.n260 0.189894
R1244 commonsourceibias.n332 commonsourceibias.n331 0.189894
R1245 commonsourceibias.n331 commonsourceibias.n330 0.189894
R1246 commonsourceibias.n330 commonsourceibias.n263 0.189894
R1247 commonsourceibias.n325 commonsourceibias.n263 0.189894
R1248 commonsourceibias.n325 commonsourceibias.n324 0.189894
R1249 commonsourceibias.n324 commonsourceibias.n323 0.189894
R1250 commonsourceibias.n323 commonsourceibias.n265 0.189894
R1251 commonsourceibias.n318 commonsourceibias.n265 0.189894
R1252 commonsourceibias.n318 commonsourceibias.n317 0.189894
R1253 commonsourceibias.n317 commonsourceibias.n316 0.189894
R1254 commonsourceibias.n316 commonsourceibias.n268 0.189894
R1255 commonsourceibias.n311 commonsourceibias.n268 0.189894
R1256 commonsourceibias.n311 commonsourceibias.n310 0.189894
R1257 commonsourceibias.n310 commonsourceibias.n309 0.189894
R1258 commonsourceibias.n309 commonsourceibias.n270 0.189894
R1259 commonsourceibias.n304 commonsourceibias.n270 0.189894
R1260 commonsourceibias.n304 commonsourceibias.n303 0.189894
R1261 commonsourceibias.n303 commonsourceibias.n302 0.189894
R1262 commonsourceibias.n302 commonsourceibias.n273 0.189894
R1263 commonsourceibias.n297 commonsourceibias.n273 0.189894
R1264 commonsourceibias.n297 commonsourceibias.n296 0.189894
R1265 commonsourceibias.n296 commonsourceibias.n295 0.189894
R1266 commonsourceibias.n295 commonsourceibias.n275 0.189894
R1267 commonsourceibias.n290 commonsourceibias.n275 0.189894
R1268 commonsourceibias.n290 commonsourceibias.n289 0.189894
R1269 commonsourceibias.n289 commonsourceibias.n288 0.189894
R1270 commonsourceibias.n288 commonsourceibias.n278 0.189894
R1271 commonsourceibias.n283 commonsourceibias.n278 0.189894
R1272 commonsourceibias.n283 commonsourceibias.n282 0.189894
R1273 commonsourceibias.n123 commonsourceibias.n14 0.189894
R1274 commonsourceibias.n123 commonsourceibias.n122 0.189894
R1275 commonsourceibias.n122 commonsourceibias.n121 0.189894
R1276 commonsourceibias.n121 commonsourceibias.n16 0.189894
R1277 commonsourceibias.n116 commonsourceibias.n16 0.189894
R1278 commonsourceibias.n116 commonsourceibias.n115 0.189894
R1279 commonsourceibias.n115 commonsourceibias.n114 0.189894
R1280 commonsourceibias.n114 commonsourceibias.n18 0.189894
R1281 commonsourceibias.n109 commonsourceibias.n18 0.189894
R1282 commonsourceibias.n109 commonsourceibias.n108 0.189894
R1283 commonsourceibias.n108 commonsourceibias.n107 0.189894
R1284 commonsourceibias.n107 commonsourceibias.n21 0.189894
R1285 commonsourceibias.n102 commonsourceibias.n21 0.189894
R1286 commonsourceibias.n102 commonsourceibias.n101 0.189894
R1287 commonsourceibias.n101 commonsourceibias.n100 0.189894
R1288 commonsourceibias.n100 commonsourceibias.n23 0.189894
R1289 commonsourceibias.n95 commonsourceibias.n23 0.189894
R1290 commonsourceibias.n95 commonsourceibias.n94 0.189894
R1291 commonsourceibias.n94 commonsourceibias.n93 0.189894
R1292 commonsourceibias.n93 commonsourceibias.n26 0.189894
R1293 commonsourceibias.n88 commonsourceibias.n26 0.189894
R1294 commonsourceibias.n88 commonsourceibias.n87 0.189894
R1295 commonsourceibias.n87 commonsourceibias.n86 0.189894
R1296 commonsourceibias.n86 commonsourceibias.n28 0.189894
R1297 commonsourceibias.n81 commonsourceibias.n28 0.189894
R1298 commonsourceibias.n81 commonsourceibias.n80 0.189894
R1299 commonsourceibias.n80 commonsourceibias.n79 0.189894
R1300 commonsourceibias.n79 commonsourceibias.n31 0.189894
R1301 commonsourceibias.n74 commonsourceibias.n31 0.189894
R1302 commonsourceibias.n74 commonsourceibias.n73 0.189894
R1303 commonsourceibias.n73 commonsourceibias.n72 0.189894
R1304 commonsourceibias.n72 commonsourceibias.n33 0.189894
R1305 commonsourceibias.n67 commonsourceibias.n33 0.189894
R1306 commonsourceibias.n67 commonsourceibias.n66 0.189894
R1307 commonsourceibias.n66 commonsourceibias.n65 0.189894
R1308 commonsourceibias.n65 commonsourceibias.n36 0.189894
R1309 commonsourceibias.n60 commonsourceibias.n36 0.189894
R1310 commonsourceibias.n60 commonsourceibias.n59 0.189894
R1311 commonsourceibias.n59 commonsourceibias.n58 0.189894
R1312 commonsourceibias.n58 commonsourceibias.n38 0.189894
R1313 commonsourceibias.n53 commonsourceibias.n38 0.189894
R1314 commonsourceibias.n53 commonsourceibias.n52 0.189894
R1315 commonsourceibias.n52 commonsourceibias.n51 0.189894
R1316 commonsourceibias.n51 commonsourceibias.n41 0.189894
R1317 commonsourceibias.n46 commonsourceibias.n41 0.189894
R1318 commonsourceibias.n46 commonsourceibias.n45 0.189894
R1319 commonsourceibias.n205 commonsourceibias.n204 0.189894
R1320 commonsourceibias.n204 commonsourceibias.n152 0.189894
R1321 commonsourceibias.n200 commonsourceibias.n152 0.189894
R1322 commonsourceibias.n200 commonsourceibias.n199 0.189894
R1323 commonsourceibias.n199 commonsourceibias.n154 0.189894
R1324 commonsourceibias.n195 commonsourceibias.n154 0.189894
R1325 commonsourceibias.n195 commonsourceibias.n194 0.189894
R1326 commonsourceibias.n194 commonsourceibias.n156 0.189894
R1327 commonsourceibias.n189 commonsourceibias.n156 0.189894
R1328 commonsourceibias.n189 commonsourceibias.n188 0.189894
R1329 commonsourceibias.n188 commonsourceibias.n187 0.189894
R1330 commonsourceibias.n187 commonsourceibias.n158 0.189894
R1331 commonsourceibias.n182 commonsourceibias.n158 0.189894
R1332 commonsourceibias.n182 commonsourceibias.n181 0.189894
R1333 commonsourceibias.n181 commonsourceibias.n180 0.189894
R1334 commonsourceibias.n180 commonsourceibias.n160 0.189894
R1335 commonsourceibias.n175 commonsourceibias.n160 0.189894
R1336 commonsourceibias.n175 commonsourceibias.n174 0.189894
R1337 commonsourceibias.n174 commonsourceibias.n173 0.189894
R1338 commonsourceibias.n173 commonsourceibias.n163 0.189894
R1339 commonsourceibias.n168 commonsourceibias.n163 0.189894
R1340 commonsourceibias.n168 commonsourceibias.n167 0.189894
R1341 commonsourceibias.n245 commonsourceibias.n0 0.189894
R1342 commonsourceibias.n245 commonsourceibias.n244 0.189894
R1343 commonsourceibias.n244 commonsourceibias.n243 0.189894
R1344 commonsourceibias.n243 commonsourceibias.n2 0.189894
R1345 commonsourceibias.n238 commonsourceibias.n2 0.189894
R1346 commonsourceibias.n238 commonsourceibias.n237 0.189894
R1347 commonsourceibias.n237 commonsourceibias.n236 0.189894
R1348 commonsourceibias.n236 commonsourceibias.n4 0.189894
R1349 commonsourceibias.n231 commonsourceibias.n4 0.189894
R1350 commonsourceibias.n231 commonsourceibias.n230 0.189894
R1351 commonsourceibias.n230 commonsourceibias.n229 0.189894
R1352 commonsourceibias.n229 commonsourceibias.n7 0.189894
R1353 commonsourceibias.n224 commonsourceibias.n7 0.189894
R1354 commonsourceibias.n224 commonsourceibias.n223 0.189894
R1355 commonsourceibias.n223 commonsourceibias.n222 0.189894
R1356 commonsourceibias.n222 commonsourceibias.n9 0.189894
R1357 commonsourceibias.n217 commonsourceibias.n9 0.189894
R1358 commonsourceibias.n217 commonsourceibias.n216 0.189894
R1359 commonsourceibias.n216 commonsourceibias.n215 0.189894
R1360 commonsourceibias.n215 commonsourceibias.n12 0.189894
R1361 commonsourceibias.n210 commonsourceibias.n12 0.189894
R1362 commonsourceibias.n210 commonsourceibias.n209 0.189894
R1363 commonsourceibias.n209 commonsourceibias.n208 0.189894
R1364 commonsourceibias.n877 commonsourceibias.n876 0.189894
R1365 commonsourceibias.n877 commonsourceibias.n872 0.189894
R1366 commonsourceibias.n882 commonsourceibias.n872 0.189894
R1367 commonsourceibias.n883 commonsourceibias.n882 0.189894
R1368 commonsourceibias.n884 commonsourceibias.n883 0.189894
R1369 commonsourceibias.n884 commonsourceibias.n870 0.189894
R1370 commonsourceibias.n890 commonsourceibias.n870 0.189894
R1371 commonsourceibias.n891 commonsourceibias.n890 0.189894
R1372 commonsourceibias.n892 commonsourceibias.n891 0.189894
R1373 commonsourceibias.n892 commonsourceibias.n868 0.189894
R1374 commonsourceibias.n897 commonsourceibias.n868 0.189894
R1375 commonsourceibias.n898 commonsourceibias.n897 0.189894
R1376 commonsourceibias.n899 commonsourceibias.n898 0.189894
R1377 commonsourceibias.n899 commonsourceibias.n866 0.189894
R1378 commonsourceibias.n905 commonsourceibias.n866 0.189894
R1379 commonsourceibias.n906 commonsourceibias.n905 0.189894
R1380 commonsourceibias.n907 commonsourceibias.n906 0.189894
R1381 commonsourceibias.n907 commonsourceibias.n864 0.189894
R1382 commonsourceibias.n912 commonsourceibias.n864 0.189894
R1383 commonsourceibias.n913 commonsourceibias.n912 0.189894
R1384 commonsourceibias.n914 commonsourceibias.n913 0.189894
R1385 commonsourceibias.n914 commonsourceibias.n862 0.189894
R1386 commonsourceibias.n920 commonsourceibias.n862 0.189894
R1387 commonsourceibias.n921 commonsourceibias.n920 0.189894
R1388 commonsourceibias.n922 commonsourceibias.n921 0.189894
R1389 commonsourceibias.n922 commonsourceibias.n860 0.189894
R1390 commonsourceibias.n927 commonsourceibias.n860 0.189894
R1391 commonsourceibias.n928 commonsourceibias.n927 0.189894
R1392 commonsourceibias.n929 commonsourceibias.n928 0.189894
R1393 commonsourceibias.n929 commonsourceibias.n858 0.189894
R1394 commonsourceibias.n935 commonsourceibias.n858 0.189894
R1395 commonsourceibias.n936 commonsourceibias.n935 0.189894
R1396 commonsourceibias.n937 commonsourceibias.n936 0.189894
R1397 commonsourceibias.n937 commonsourceibias.n856 0.189894
R1398 commonsourceibias.n942 commonsourceibias.n856 0.189894
R1399 commonsourceibias.n943 commonsourceibias.n942 0.189894
R1400 commonsourceibias.n944 commonsourceibias.n943 0.189894
R1401 commonsourceibias.n944 commonsourceibias.n854 0.189894
R1402 commonsourceibias.n950 commonsourceibias.n854 0.189894
R1403 commonsourceibias.n951 commonsourceibias.n950 0.189894
R1404 commonsourceibias.n952 commonsourceibias.n951 0.189894
R1405 commonsourceibias.n952 commonsourceibias.n852 0.189894
R1406 commonsourceibias.n957 commonsourceibias.n852 0.189894
R1407 commonsourceibias.n958 commonsourceibias.n957 0.189894
R1408 commonsourceibias.n959 commonsourceibias.n958 0.189894
R1409 commonsourceibias.n959 commonsourceibias.n850 0.189894
R1410 commonsourceibias.n761 commonsourceibias.n760 0.189894
R1411 commonsourceibias.n761 commonsourceibias.n756 0.189894
R1412 commonsourceibias.n766 commonsourceibias.n756 0.189894
R1413 commonsourceibias.n767 commonsourceibias.n766 0.189894
R1414 commonsourceibias.n768 commonsourceibias.n767 0.189894
R1415 commonsourceibias.n768 commonsourceibias.n754 0.189894
R1416 commonsourceibias.n774 commonsourceibias.n754 0.189894
R1417 commonsourceibias.n775 commonsourceibias.n774 0.189894
R1418 commonsourceibias.n776 commonsourceibias.n775 0.189894
R1419 commonsourceibias.n776 commonsourceibias.n752 0.189894
R1420 commonsourceibias.n781 commonsourceibias.n752 0.189894
R1421 commonsourceibias.n782 commonsourceibias.n781 0.189894
R1422 commonsourceibias.n783 commonsourceibias.n782 0.189894
R1423 commonsourceibias.n783 commonsourceibias.n750 0.189894
R1424 commonsourceibias.n789 commonsourceibias.n750 0.189894
R1425 commonsourceibias.n790 commonsourceibias.n789 0.189894
R1426 commonsourceibias.n791 commonsourceibias.n790 0.189894
R1427 commonsourceibias.n791 commonsourceibias.n748 0.189894
R1428 commonsourceibias.n796 commonsourceibias.n748 0.189894
R1429 commonsourceibias.n797 commonsourceibias.n796 0.189894
R1430 commonsourceibias.n798 commonsourceibias.n797 0.189894
R1431 commonsourceibias.n798 commonsourceibias.n746 0.189894
R1432 commonsourceibias.n804 commonsourceibias.n746 0.189894
R1433 commonsourceibias.n805 commonsourceibias.n804 0.189894
R1434 commonsourceibias.n806 commonsourceibias.n805 0.189894
R1435 commonsourceibias.n806 commonsourceibias.n744 0.189894
R1436 commonsourceibias.n811 commonsourceibias.n744 0.189894
R1437 commonsourceibias.n812 commonsourceibias.n811 0.189894
R1438 commonsourceibias.n813 commonsourceibias.n812 0.189894
R1439 commonsourceibias.n813 commonsourceibias.n742 0.189894
R1440 commonsourceibias.n819 commonsourceibias.n742 0.189894
R1441 commonsourceibias.n820 commonsourceibias.n819 0.189894
R1442 commonsourceibias.n821 commonsourceibias.n820 0.189894
R1443 commonsourceibias.n821 commonsourceibias.n740 0.189894
R1444 commonsourceibias.n826 commonsourceibias.n740 0.189894
R1445 commonsourceibias.n827 commonsourceibias.n826 0.189894
R1446 commonsourceibias.n828 commonsourceibias.n827 0.189894
R1447 commonsourceibias.n828 commonsourceibias.n738 0.189894
R1448 commonsourceibias.n834 commonsourceibias.n738 0.189894
R1449 commonsourceibias.n835 commonsourceibias.n834 0.189894
R1450 commonsourceibias.n836 commonsourceibias.n835 0.189894
R1451 commonsourceibias.n836 commonsourceibias.n736 0.189894
R1452 commonsourceibias.n841 commonsourceibias.n736 0.189894
R1453 commonsourceibias.n842 commonsourceibias.n841 0.189894
R1454 commonsourceibias.n843 commonsourceibias.n842 0.189894
R1455 commonsourceibias.n843 commonsourceibias.n734 0.189894
R1456 commonsourceibias.n531 commonsourceibias.n530 0.189894
R1457 commonsourceibias.n531 commonsourceibias.n526 0.189894
R1458 commonsourceibias.n536 commonsourceibias.n526 0.189894
R1459 commonsourceibias.n537 commonsourceibias.n536 0.189894
R1460 commonsourceibias.n538 commonsourceibias.n537 0.189894
R1461 commonsourceibias.n538 commonsourceibias.n524 0.189894
R1462 commonsourceibias.n544 commonsourceibias.n524 0.189894
R1463 commonsourceibias.n545 commonsourceibias.n544 0.189894
R1464 commonsourceibias.n546 commonsourceibias.n545 0.189894
R1465 commonsourceibias.n546 commonsourceibias.n522 0.189894
R1466 commonsourceibias.n551 commonsourceibias.n522 0.189894
R1467 commonsourceibias.n552 commonsourceibias.n551 0.189894
R1468 commonsourceibias.n553 commonsourceibias.n552 0.189894
R1469 commonsourceibias.n553 commonsourceibias.n520 0.189894
R1470 commonsourceibias.n559 commonsourceibias.n520 0.189894
R1471 commonsourceibias.n560 commonsourceibias.n559 0.189894
R1472 commonsourceibias.n561 commonsourceibias.n560 0.189894
R1473 commonsourceibias.n561 commonsourceibias.n518 0.189894
R1474 commonsourceibias.n566 commonsourceibias.n518 0.189894
R1475 commonsourceibias.n567 commonsourceibias.n566 0.189894
R1476 commonsourceibias.n568 commonsourceibias.n567 0.189894
R1477 commonsourceibias.n568 commonsourceibias.n516 0.189894
R1478 commonsourceibias.n574 commonsourceibias.n516 0.189894
R1479 commonsourceibias.n575 commonsourceibias.n574 0.189894
R1480 commonsourceibias.n576 commonsourceibias.n575 0.189894
R1481 commonsourceibias.n576 commonsourceibias.n514 0.189894
R1482 commonsourceibias.n581 commonsourceibias.n514 0.189894
R1483 commonsourceibias.n582 commonsourceibias.n581 0.189894
R1484 commonsourceibias.n583 commonsourceibias.n582 0.189894
R1485 commonsourceibias.n583 commonsourceibias.n512 0.189894
R1486 commonsourceibias.n589 commonsourceibias.n512 0.189894
R1487 commonsourceibias.n590 commonsourceibias.n589 0.189894
R1488 commonsourceibias.n591 commonsourceibias.n590 0.189894
R1489 commonsourceibias.n591 commonsourceibias.n510 0.189894
R1490 commonsourceibias.n596 commonsourceibias.n510 0.189894
R1491 commonsourceibias.n597 commonsourceibias.n596 0.189894
R1492 commonsourceibias.n598 commonsourceibias.n597 0.189894
R1493 commonsourceibias.n598 commonsourceibias.n508 0.189894
R1494 commonsourceibias.n604 commonsourceibias.n508 0.189894
R1495 commonsourceibias.n605 commonsourceibias.n604 0.189894
R1496 commonsourceibias.n606 commonsourceibias.n605 0.189894
R1497 commonsourceibias.n606 commonsourceibias.n506 0.189894
R1498 commonsourceibias.n611 commonsourceibias.n506 0.189894
R1499 commonsourceibias.n612 commonsourceibias.n611 0.189894
R1500 commonsourceibias.n613 commonsourceibias.n612 0.189894
R1501 commonsourceibias.n613 commonsourceibias.n504 0.189894
R1502 commonsourceibias.n647 commonsourceibias.n646 0.189894
R1503 commonsourceibias.n647 commonsourceibias.n642 0.189894
R1504 commonsourceibias.n652 commonsourceibias.n642 0.189894
R1505 commonsourceibias.n653 commonsourceibias.n652 0.189894
R1506 commonsourceibias.n654 commonsourceibias.n653 0.189894
R1507 commonsourceibias.n654 commonsourceibias.n640 0.189894
R1508 commonsourceibias.n660 commonsourceibias.n640 0.189894
R1509 commonsourceibias.n661 commonsourceibias.n660 0.189894
R1510 commonsourceibias.n662 commonsourceibias.n661 0.189894
R1511 commonsourceibias.n662 commonsourceibias.n638 0.189894
R1512 commonsourceibias.n667 commonsourceibias.n638 0.189894
R1513 commonsourceibias.n668 commonsourceibias.n667 0.189894
R1514 commonsourceibias.n669 commonsourceibias.n668 0.189894
R1515 commonsourceibias.n669 commonsourceibias.n636 0.189894
R1516 commonsourceibias.n674 commonsourceibias.n636 0.189894
R1517 commonsourceibias.n675 commonsourceibias.n674 0.189894
R1518 commonsourceibias.n675 commonsourceibias.n634 0.189894
R1519 commonsourceibias.n679 commonsourceibias.n634 0.189894
R1520 commonsourceibias.n680 commonsourceibias.n679 0.189894
R1521 commonsourceibias.n680 commonsourceibias.n632 0.189894
R1522 commonsourceibias.n684 commonsourceibias.n632 0.189894
R1523 commonsourceibias.n685 commonsourceibias.n684 0.189894
R1524 commonsourceibias.n690 commonsourceibias.n689 0.189894
R1525 commonsourceibias.n691 commonsourceibias.n690 0.189894
R1526 commonsourceibias.n691 commonsourceibias.n493 0.189894
R1527 commonsourceibias.n696 commonsourceibias.n493 0.189894
R1528 commonsourceibias.n697 commonsourceibias.n696 0.189894
R1529 commonsourceibias.n698 commonsourceibias.n697 0.189894
R1530 commonsourceibias.n698 commonsourceibias.n491 0.189894
R1531 commonsourceibias.n704 commonsourceibias.n491 0.189894
R1532 commonsourceibias.n705 commonsourceibias.n704 0.189894
R1533 commonsourceibias.n706 commonsourceibias.n705 0.189894
R1534 commonsourceibias.n706 commonsourceibias.n489 0.189894
R1535 commonsourceibias.n711 commonsourceibias.n489 0.189894
R1536 commonsourceibias.n712 commonsourceibias.n711 0.189894
R1537 commonsourceibias.n713 commonsourceibias.n712 0.189894
R1538 commonsourceibias.n713 commonsourceibias.n487 0.189894
R1539 commonsourceibias.n719 commonsourceibias.n487 0.189894
R1540 commonsourceibias.n720 commonsourceibias.n719 0.189894
R1541 commonsourceibias.n721 commonsourceibias.n720 0.189894
R1542 commonsourceibias.n721 commonsourceibias.n485 0.189894
R1543 commonsourceibias.n726 commonsourceibias.n485 0.189894
R1544 commonsourceibias.n727 commonsourceibias.n726 0.189894
R1545 commonsourceibias.n728 commonsourceibias.n727 0.189894
R1546 commonsourceibias.n728 commonsourceibias.n483 0.189894
R1547 commonsourceibias.n205 commonsourceibias.n149 0.0762576
R1548 commonsourceibias.n208 commonsourceibias.n149 0.0762576
R1549 commonsourceibias.n685 commonsourceibias.n630 0.0762576
R1550 commonsourceibias.n689 commonsourceibias.n630 0.0762576
R1551 gnd.n7511 gnd.n694 1008.05
R1552 gnd.n5401 gnd.n5400 939.716
R1553 gnd.n6877 gnd.n1144 766.379
R1554 gnd.n6793 gnd.n1146 766.379
R1555 gnd.n6157 gnd.n6056 766.379
R1556 gnd.n6155 gnd.n6058 766.379
R1557 gnd.n6874 gnd.n5403 756.769
R1558 gnd.n6843 gnd.n1147 756.769
R1559 gnd.n6434 gnd.n6018 756.769
R1560 gnd.n6420 gnd.n6008 756.769
R1561 gnd.n257 gnd.n247 751.963
R1562 gnd.n446 gnd.n445 751.963
R1563 gnd.n1935 gnd.n1858 751.963
R1564 gnd.n4715 gnd.n1937 751.963
R1565 gnd.n1557 gnd.n1545 751.963
R1566 gnd.n3363 gnd.n3362 751.963
R1567 gnd.n2958 gnd.n1185 751.963
R1568 gnd.n2914 gnd.n2913 751.963
R1569 gnd.n3349 gnd.n2543 711.122
R1570 gnd.n4846 gnd.n1808 711.122
R1571 gnd.n3372 gnd.n2545 711.122
R1572 gnd.n4562 gnd.n1811 711.122
R1573 gnd.n8004 gnd.n251 696.707
R1574 gnd.n7880 gnd.n7879 696.707
R1575 gnd.n4717 gnd.n1932 696.707
R1576 gnd.n4834 gnd.n1862 696.707
R1577 gnd.n5100 gnd.n1550 696.707
R1578 gnd.n2733 gnd.n2554 696.707
R1579 gnd.n5278 gnd.n1258 696.707
R1580 gnd.n5398 gnd.n1189 696.707
R1581 gnd.n7053 gnd.n967 670.282
R1582 gnd.n7510 gnd.n695 670.282
R1583 gnd.n7723 gnd.n7722 670.282
R1584 gnd.n2823 gnd.n1135 670.282
R1585 gnd.n970 gnd.n967 585
R1586 gnd.n7051 gnd.n967 585
R1587 gnd.n7049 gnd.n7048 585
R1588 gnd.n7050 gnd.n7049 585
R1589 gnd.n7047 gnd.n969 585
R1590 gnd.n969 gnd.n968 585
R1591 gnd.n7046 gnd.n7045 585
R1592 gnd.n7045 gnd.n7044 585
R1593 gnd.n975 gnd.n974 585
R1594 gnd.n7043 gnd.n975 585
R1595 gnd.n7041 gnd.n7040 585
R1596 gnd.n7042 gnd.n7041 585
R1597 gnd.n7039 gnd.n977 585
R1598 gnd.n977 gnd.n976 585
R1599 gnd.n7038 gnd.n7037 585
R1600 gnd.n7037 gnd.n7036 585
R1601 gnd.n983 gnd.n982 585
R1602 gnd.n7035 gnd.n983 585
R1603 gnd.n7033 gnd.n7032 585
R1604 gnd.n7034 gnd.n7033 585
R1605 gnd.n7031 gnd.n985 585
R1606 gnd.n985 gnd.n984 585
R1607 gnd.n7030 gnd.n7029 585
R1608 gnd.n7029 gnd.n7028 585
R1609 gnd.n991 gnd.n990 585
R1610 gnd.n7027 gnd.n991 585
R1611 gnd.n7025 gnd.n7024 585
R1612 gnd.n7026 gnd.n7025 585
R1613 gnd.n7023 gnd.n993 585
R1614 gnd.n993 gnd.n992 585
R1615 gnd.n7022 gnd.n7021 585
R1616 gnd.n7021 gnd.n7020 585
R1617 gnd.n999 gnd.n998 585
R1618 gnd.n7019 gnd.n999 585
R1619 gnd.n7017 gnd.n7016 585
R1620 gnd.n7018 gnd.n7017 585
R1621 gnd.n7015 gnd.n1001 585
R1622 gnd.n1001 gnd.n1000 585
R1623 gnd.n7014 gnd.n7013 585
R1624 gnd.n7013 gnd.n7012 585
R1625 gnd.n1007 gnd.n1006 585
R1626 gnd.n7011 gnd.n1007 585
R1627 gnd.n7009 gnd.n7008 585
R1628 gnd.n7010 gnd.n7009 585
R1629 gnd.n7007 gnd.n1009 585
R1630 gnd.n1009 gnd.n1008 585
R1631 gnd.n7006 gnd.n7005 585
R1632 gnd.n7005 gnd.n7004 585
R1633 gnd.n1015 gnd.n1014 585
R1634 gnd.n7003 gnd.n1015 585
R1635 gnd.n7001 gnd.n7000 585
R1636 gnd.n7002 gnd.n7001 585
R1637 gnd.n6999 gnd.n1017 585
R1638 gnd.n1017 gnd.n1016 585
R1639 gnd.n6998 gnd.n6997 585
R1640 gnd.n6997 gnd.n6996 585
R1641 gnd.n1023 gnd.n1022 585
R1642 gnd.n6995 gnd.n1023 585
R1643 gnd.n6993 gnd.n6992 585
R1644 gnd.n6994 gnd.n6993 585
R1645 gnd.n6991 gnd.n1025 585
R1646 gnd.n1025 gnd.n1024 585
R1647 gnd.n6990 gnd.n6989 585
R1648 gnd.n6989 gnd.n6988 585
R1649 gnd.n1031 gnd.n1030 585
R1650 gnd.n6987 gnd.n1031 585
R1651 gnd.n6985 gnd.n6984 585
R1652 gnd.n6986 gnd.n6985 585
R1653 gnd.n6983 gnd.n1033 585
R1654 gnd.n1033 gnd.n1032 585
R1655 gnd.n6982 gnd.n6981 585
R1656 gnd.n6981 gnd.n6980 585
R1657 gnd.n1039 gnd.n1038 585
R1658 gnd.n6979 gnd.n1039 585
R1659 gnd.n6977 gnd.n6976 585
R1660 gnd.n6978 gnd.n6977 585
R1661 gnd.n6975 gnd.n1041 585
R1662 gnd.n1041 gnd.n1040 585
R1663 gnd.n6974 gnd.n6973 585
R1664 gnd.n6973 gnd.n6972 585
R1665 gnd.n1047 gnd.n1046 585
R1666 gnd.n6971 gnd.n1047 585
R1667 gnd.n6969 gnd.n6968 585
R1668 gnd.n6970 gnd.n6969 585
R1669 gnd.n6967 gnd.n1049 585
R1670 gnd.n1049 gnd.n1048 585
R1671 gnd.n6966 gnd.n6965 585
R1672 gnd.n6965 gnd.n6964 585
R1673 gnd.n1055 gnd.n1054 585
R1674 gnd.n6963 gnd.n1055 585
R1675 gnd.n6961 gnd.n6960 585
R1676 gnd.n6962 gnd.n6961 585
R1677 gnd.n6959 gnd.n1057 585
R1678 gnd.n1057 gnd.n1056 585
R1679 gnd.n6958 gnd.n6957 585
R1680 gnd.n6957 gnd.n6956 585
R1681 gnd.n1063 gnd.n1062 585
R1682 gnd.n6955 gnd.n1063 585
R1683 gnd.n6953 gnd.n6952 585
R1684 gnd.n6954 gnd.n6953 585
R1685 gnd.n6951 gnd.n1065 585
R1686 gnd.n1065 gnd.n1064 585
R1687 gnd.n6950 gnd.n6949 585
R1688 gnd.n6949 gnd.n6948 585
R1689 gnd.n1071 gnd.n1070 585
R1690 gnd.n6947 gnd.n1071 585
R1691 gnd.n6945 gnd.n6944 585
R1692 gnd.n6946 gnd.n6945 585
R1693 gnd.n6943 gnd.n1073 585
R1694 gnd.n1073 gnd.n1072 585
R1695 gnd.n6942 gnd.n6941 585
R1696 gnd.n6941 gnd.n6940 585
R1697 gnd.n1079 gnd.n1078 585
R1698 gnd.n6939 gnd.n1079 585
R1699 gnd.n6937 gnd.n6936 585
R1700 gnd.n6938 gnd.n6937 585
R1701 gnd.n6935 gnd.n1081 585
R1702 gnd.n1081 gnd.n1080 585
R1703 gnd.n6934 gnd.n6933 585
R1704 gnd.n6933 gnd.n6932 585
R1705 gnd.n1087 gnd.n1086 585
R1706 gnd.n6931 gnd.n1087 585
R1707 gnd.n6929 gnd.n6928 585
R1708 gnd.n6930 gnd.n6929 585
R1709 gnd.n6927 gnd.n1089 585
R1710 gnd.n1089 gnd.n1088 585
R1711 gnd.n6926 gnd.n6925 585
R1712 gnd.n6925 gnd.n6924 585
R1713 gnd.n1095 gnd.n1094 585
R1714 gnd.n6923 gnd.n1095 585
R1715 gnd.n6921 gnd.n6920 585
R1716 gnd.n6922 gnd.n6921 585
R1717 gnd.n6919 gnd.n1097 585
R1718 gnd.n1097 gnd.n1096 585
R1719 gnd.n6918 gnd.n6917 585
R1720 gnd.n6917 gnd.n6916 585
R1721 gnd.n1103 gnd.n1102 585
R1722 gnd.n6915 gnd.n1103 585
R1723 gnd.n6913 gnd.n6912 585
R1724 gnd.n6914 gnd.n6913 585
R1725 gnd.n6911 gnd.n1105 585
R1726 gnd.n1105 gnd.n1104 585
R1727 gnd.n6910 gnd.n6909 585
R1728 gnd.n6909 gnd.n6908 585
R1729 gnd.n1111 gnd.n1110 585
R1730 gnd.n6907 gnd.n1111 585
R1731 gnd.n6905 gnd.n6904 585
R1732 gnd.n6906 gnd.n6905 585
R1733 gnd.n6903 gnd.n1113 585
R1734 gnd.n1113 gnd.n1112 585
R1735 gnd.n6902 gnd.n6901 585
R1736 gnd.n6901 gnd.n6900 585
R1737 gnd.n1119 gnd.n1118 585
R1738 gnd.n6899 gnd.n1119 585
R1739 gnd.n6897 gnd.n6896 585
R1740 gnd.n6898 gnd.n6897 585
R1741 gnd.n6895 gnd.n1121 585
R1742 gnd.n1121 gnd.n1120 585
R1743 gnd.n6894 gnd.n6893 585
R1744 gnd.n6893 gnd.n6892 585
R1745 gnd.n1127 gnd.n1126 585
R1746 gnd.n6891 gnd.n1127 585
R1747 gnd.n6889 gnd.n6888 585
R1748 gnd.n6890 gnd.n6889 585
R1749 gnd.n6887 gnd.n1129 585
R1750 gnd.n1129 gnd.n1128 585
R1751 gnd.n6886 gnd.n6885 585
R1752 gnd.n6885 gnd.n6884 585
R1753 gnd.n7054 gnd.n7053 585
R1754 gnd.n7053 gnd.n7052 585
R1755 gnd.n965 gnd.n964 585
R1756 gnd.n964 gnd.n963 585
R1757 gnd.n7059 gnd.n7058 585
R1758 gnd.n7060 gnd.n7059 585
R1759 gnd.n962 gnd.n961 585
R1760 gnd.n7061 gnd.n962 585
R1761 gnd.n7064 gnd.n7063 585
R1762 gnd.n7063 gnd.n7062 585
R1763 gnd.n959 gnd.n958 585
R1764 gnd.n958 gnd.n957 585
R1765 gnd.n7069 gnd.n7068 585
R1766 gnd.n7070 gnd.n7069 585
R1767 gnd.n956 gnd.n955 585
R1768 gnd.n7071 gnd.n956 585
R1769 gnd.n7074 gnd.n7073 585
R1770 gnd.n7073 gnd.n7072 585
R1771 gnd.n953 gnd.n952 585
R1772 gnd.n952 gnd.n951 585
R1773 gnd.n7079 gnd.n7078 585
R1774 gnd.n7080 gnd.n7079 585
R1775 gnd.n950 gnd.n949 585
R1776 gnd.n7081 gnd.n950 585
R1777 gnd.n7084 gnd.n7083 585
R1778 gnd.n7083 gnd.n7082 585
R1779 gnd.n947 gnd.n946 585
R1780 gnd.n946 gnd.n945 585
R1781 gnd.n7089 gnd.n7088 585
R1782 gnd.n7090 gnd.n7089 585
R1783 gnd.n944 gnd.n943 585
R1784 gnd.n7091 gnd.n944 585
R1785 gnd.n7094 gnd.n7093 585
R1786 gnd.n7093 gnd.n7092 585
R1787 gnd.n941 gnd.n940 585
R1788 gnd.n940 gnd.n939 585
R1789 gnd.n7099 gnd.n7098 585
R1790 gnd.n7100 gnd.n7099 585
R1791 gnd.n938 gnd.n937 585
R1792 gnd.n7101 gnd.n938 585
R1793 gnd.n7104 gnd.n7103 585
R1794 gnd.n7103 gnd.n7102 585
R1795 gnd.n935 gnd.n934 585
R1796 gnd.n934 gnd.n933 585
R1797 gnd.n7109 gnd.n7108 585
R1798 gnd.n7110 gnd.n7109 585
R1799 gnd.n932 gnd.n931 585
R1800 gnd.n7111 gnd.n932 585
R1801 gnd.n7114 gnd.n7113 585
R1802 gnd.n7113 gnd.n7112 585
R1803 gnd.n929 gnd.n928 585
R1804 gnd.n928 gnd.n927 585
R1805 gnd.n7119 gnd.n7118 585
R1806 gnd.n7120 gnd.n7119 585
R1807 gnd.n926 gnd.n925 585
R1808 gnd.n7121 gnd.n926 585
R1809 gnd.n7124 gnd.n7123 585
R1810 gnd.n7123 gnd.n7122 585
R1811 gnd.n923 gnd.n922 585
R1812 gnd.n922 gnd.n921 585
R1813 gnd.n7129 gnd.n7128 585
R1814 gnd.n7130 gnd.n7129 585
R1815 gnd.n920 gnd.n919 585
R1816 gnd.n7131 gnd.n920 585
R1817 gnd.n7134 gnd.n7133 585
R1818 gnd.n7133 gnd.n7132 585
R1819 gnd.n917 gnd.n916 585
R1820 gnd.n916 gnd.n915 585
R1821 gnd.n7139 gnd.n7138 585
R1822 gnd.n7140 gnd.n7139 585
R1823 gnd.n914 gnd.n913 585
R1824 gnd.n7141 gnd.n914 585
R1825 gnd.n7144 gnd.n7143 585
R1826 gnd.n7143 gnd.n7142 585
R1827 gnd.n911 gnd.n910 585
R1828 gnd.n910 gnd.n909 585
R1829 gnd.n7149 gnd.n7148 585
R1830 gnd.n7150 gnd.n7149 585
R1831 gnd.n908 gnd.n907 585
R1832 gnd.n7151 gnd.n908 585
R1833 gnd.n7154 gnd.n7153 585
R1834 gnd.n7153 gnd.n7152 585
R1835 gnd.n905 gnd.n904 585
R1836 gnd.n904 gnd.n903 585
R1837 gnd.n7159 gnd.n7158 585
R1838 gnd.n7160 gnd.n7159 585
R1839 gnd.n902 gnd.n901 585
R1840 gnd.n7161 gnd.n902 585
R1841 gnd.n7164 gnd.n7163 585
R1842 gnd.n7163 gnd.n7162 585
R1843 gnd.n899 gnd.n898 585
R1844 gnd.n898 gnd.n897 585
R1845 gnd.n7169 gnd.n7168 585
R1846 gnd.n7170 gnd.n7169 585
R1847 gnd.n896 gnd.n895 585
R1848 gnd.n7171 gnd.n896 585
R1849 gnd.n7174 gnd.n7173 585
R1850 gnd.n7173 gnd.n7172 585
R1851 gnd.n893 gnd.n892 585
R1852 gnd.n892 gnd.n891 585
R1853 gnd.n7179 gnd.n7178 585
R1854 gnd.n7180 gnd.n7179 585
R1855 gnd.n890 gnd.n889 585
R1856 gnd.n7181 gnd.n890 585
R1857 gnd.n7184 gnd.n7183 585
R1858 gnd.n7183 gnd.n7182 585
R1859 gnd.n887 gnd.n886 585
R1860 gnd.n886 gnd.n885 585
R1861 gnd.n7189 gnd.n7188 585
R1862 gnd.n7190 gnd.n7189 585
R1863 gnd.n884 gnd.n883 585
R1864 gnd.n7191 gnd.n884 585
R1865 gnd.n7194 gnd.n7193 585
R1866 gnd.n7193 gnd.n7192 585
R1867 gnd.n881 gnd.n880 585
R1868 gnd.n880 gnd.n879 585
R1869 gnd.n7199 gnd.n7198 585
R1870 gnd.n7200 gnd.n7199 585
R1871 gnd.n878 gnd.n877 585
R1872 gnd.n7201 gnd.n878 585
R1873 gnd.n7204 gnd.n7203 585
R1874 gnd.n7203 gnd.n7202 585
R1875 gnd.n875 gnd.n874 585
R1876 gnd.n874 gnd.n873 585
R1877 gnd.n7209 gnd.n7208 585
R1878 gnd.n7210 gnd.n7209 585
R1879 gnd.n872 gnd.n871 585
R1880 gnd.n7211 gnd.n872 585
R1881 gnd.n7214 gnd.n7213 585
R1882 gnd.n7213 gnd.n7212 585
R1883 gnd.n869 gnd.n868 585
R1884 gnd.n868 gnd.n867 585
R1885 gnd.n7219 gnd.n7218 585
R1886 gnd.n7220 gnd.n7219 585
R1887 gnd.n866 gnd.n865 585
R1888 gnd.n7221 gnd.n866 585
R1889 gnd.n7224 gnd.n7223 585
R1890 gnd.n7223 gnd.n7222 585
R1891 gnd.n863 gnd.n862 585
R1892 gnd.n862 gnd.n861 585
R1893 gnd.n7229 gnd.n7228 585
R1894 gnd.n7230 gnd.n7229 585
R1895 gnd.n860 gnd.n859 585
R1896 gnd.n7231 gnd.n860 585
R1897 gnd.n7234 gnd.n7233 585
R1898 gnd.n7233 gnd.n7232 585
R1899 gnd.n857 gnd.n856 585
R1900 gnd.n856 gnd.n855 585
R1901 gnd.n7239 gnd.n7238 585
R1902 gnd.n7240 gnd.n7239 585
R1903 gnd.n854 gnd.n853 585
R1904 gnd.n7241 gnd.n854 585
R1905 gnd.n7244 gnd.n7243 585
R1906 gnd.n7243 gnd.n7242 585
R1907 gnd.n851 gnd.n850 585
R1908 gnd.n850 gnd.n849 585
R1909 gnd.n7249 gnd.n7248 585
R1910 gnd.n7250 gnd.n7249 585
R1911 gnd.n848 gnd.n847 585
R1912 gnd.n7251 gnd.n848 585
R1913 gnd.n7254 gnd.n7253 585
R1914 gnd.n7253 gnd.n7252 585
R1915 gnd.n845 gnd.n844 585
R1916 gnd.n844 gnd.n843 585
R1917 gnd.n7259 gnd.n7258 585
R1918 gnd.n7260 gnd.n7259 585
R1919 gnd.n842 gnd.n841 585
R1920 gnd.n7261 gnd.n842 585
R1921 gnd.n7264 gnd.n7263 585
R1922 gnd.n7263 gnd.n7262 585
R1923 gnd.n839 gnd.n838 585
R1924 gnd.n838 gnd.n837 585
R1925 gnd.n7269 gnd.n7268 585
R1926 gnd.n7270 gnd.n7269 585
R1927 gnd.n836 gnd.n835 585
R1928 gnd.n7271 gnd.n836 585
R1929 gnd.n7274 gnd.n7273 585
R1930 gnd.n7273 gnd.n7272 585
R1931 gnd.n833 gnd.n832 585
R1932 gnd.n832 gnd.n831 585
R1933 gnd.n7279 gnd.n7278 585
R1934 gnd.n7280 gnd.n7279 585
R1935 gnd.n830 gnd.n829 585
R1936 gnd.n7281 gnd.n830 585
R1937 gnd.n7284 gnd.n7283 585
R1938 gnd.n7283 gnd.n7282 585
R1939 gnd.n827 gnd.n826 585
R1940 gnd.n826 gnd.n825 585
R1941 gnd.n7289 gnd.n7288 585
R1942 gnd.n7290 gnd.n7289 585
R1943 gnd.n824 gnd.n823 585
R1944 gnd.n7291 gnd.n824 585
R1945 gnd.n7294 gnd.n7293 585
R1946 gnd.n7293 gnd.n7292 585
R1947 gnd.n821 gnd.n820 585
R1948 gnd.n820 gnd.n819 585
R1949 gnd.n7299 gnd.n7298 585
R1950 gnd.n7300 gnd.n7299 585
R1951 gnd.n818 gnd.n817 585
R1952 gnd.n7301 gnd.n818 585
R1953 gnd.n7304 gnd.n7303 585
R1954 gnd.n7303 gnd.n7302 585
R1955 gnd.n815 gnd.n814 585
R1956 gnd.n814 gnd.n813 585
R1957 gnd.n7309 gnd.n7308 585
R1958 gnd.n7310 gnd.n7309 585
R1959 gnd.n812 gnd.n811 585
R1960 gnd.n7311 gnd.n812 585
R1961 gnd.n7314 gnd.n7313 585
R1962 gnd.n7313 gnd.n7312 585
R1963 gnd.n809 gnd.n808 585
R1964 gnd.n808 gnd.n807 585
R1965 gnd.n7319 gnd.n7318 585
R1966 gnd.n7320 gnd.n7319 585
R1967 gnd.n806 gnd.n805 585
R1968 gnd.n7321 gnd.n806 585
R1969 gnd.n7324 gnd.n7323 585
R1970 gnd.n7323 gnd.n7322 585
R1971 gnd.n803 gnd.n802 585
R1972 gnd.n802 gnd.n801 585
R1973 gnd.n7329 gnd.n7328 585
R1974 gnd.n7330 gnd.n7329 585
R1975 gnd.n800 gnd.n799 585
R1976 gnd.n7331 gnd.n800 585
R1977 gnd.n7334 gnd.n7333 585
R1978 gnd.n7333 gnd.n7332 585
R1979 gnd.n797 gnd.n796 585
R1980 gnd.n796 gnd.n795 585
R1981 gnd.n7339 gnd.n7338 585
R1982 gnd.n7340 gnd.n7339 585
R1983 gnd.n794 gnd.n793 585
R1984 gnd.n7341 gnd.n794 585
R1985 gnd.n7344 gnd.n7343 585
R1986 gnd.n7343 gnd.n7342 585
R1987 gnd.n791 gnd.n790 585
R1988 gnd.n790 gnd.n789 585
R1989 gnd.n7349 gnd.n7348 585
R1990 gnd.n7350 gnd.n7349 585
R1991 gnd.n788 gnd.n787 585
R1992 gnd.n7351 gnd.n788 585
R1993 gnd.n7354 gnd.n7353 585
R1994 gnd.n7353 gnd.n7352 585
R1995 gnd.n785 gnd.n784 585
R1996 gnd.n784 gnd.n783 585
R1997 gnd.n7359 gnd.n7358 585
R1998 gnd.n7360 gnd.n7359 585
R1999 gnd.n782 gnd.n781 585
R2000 gnd.n7361 gnd.n782 585
R2001 gnd.n7364 gnd.n7363 585
R2002 gnd.n7363 gnd.n7362 585
R2003 gnd.n779 gnd.n778 585
R2004 gnd.n778 gnd.n777 585
R2005 gnd.n7369 gnd.n7368 585
R2006 gnd.n7370 gnd.n7369 585
R2007 gnd.n776 gnd.n775 585
R2008 gnd.n7371 gnd.n776 585
R2009 gnd.n7374 gnd.n7373 585
R2010 gnd.n7373 gnd.n7372 585
R2011 gnd.n773 gnd.n772 585
R2012 gnd.n772 gnd.n771 585
R2013 gnd.n7379 gnd.n7378 585
R2014 gnd.n7380 gnd.n7379 585
R2015 gnd.n770 gnd.n769 585
R2016 gnd.n7381 gnd.n770 585
R2017 gnd.n7384 gnd.n7383 585
R2018 gnd.n7383 gnd.n7382 585
R2019 gnd.n767 gnd.n766 585
R2020 gnd.n766 gnd.n765 585
R2021 gnd.n7389 gnd.n7388 585
R2022 gnd.n7390 gnd.n7389 585
R2023 gnd.n764 gnd.n763 585
R2024 gnd.n7391 gnd.n764 585
R2025 gnd.n7394 gnd.n7393 585
R2026 gnd.n7393 gnd.n7392 585
R2027 gnd.n761 gnd.n760 585
R2028 gnd.n760 gnd.n759 585
R2029 gnd.n7399 gnd.n7398 585
R2030 gnd.n7400 gnd.n7399 585
R2031 gnd.n758 gnd.n757 585
R2032 gnd.n7401 gnd.n758 585
R2033 gnd.n7404 gnd.n7403 585
R2034 gnd.n7403 gnd.n7402 585
R2035 gnd.n755 gnd.n754 585
R2036 gnd.n754 gnd.n753 585
R2037 gnd.n7409 gnd.n7408 585
R2038 gnd.n7410 gnd.n7409 585
R2039 gnd.n752 gnd.n751 585
R2040 gnd.n7411 gnd.n752 585
R2041 gnd.n7414 gnd.n7413 585
R2042 gnd.n7413 gnd.n7412 585
R2043 gnd.n749 gnd.n748 585
R2044 gnd.n748 gnd.n747 585
R2045 gnd.n7419 gnd.n7418 585
R2046 gnd.n7420 gnd.n7419 585
R2047 gnd.n746 gnd.n745 585
R2048 gnd.n7421 gnd.n746 585
R2049 gnd.n7424 gnd.n7423 585
R2050 gnd.n7423 gnd.n7422 585
R2051 gnd.n743 gnd.n742 585
R2052 gnd.n742 gnd.n741 585
R2053 gnd.n7429 gnd.n7428 585
R2054 gnd.n7430 gnd.n7429 585
R2055 gnd.n740 gnd.n739 585
R2056 gnd.n7431 gnd.n740 585
R2057 gnd.n7434 gnd.n7433 585
R2058 gnd.n7433 gnd.n7432 585
R2059 gnd.n737 gnd.n736 585
R2060 gnd.n736 gnd.n735 585
R2061 gnd.n7439 gnd.n7438 585
R2062 gnd.n7440 gnd.n7439 585
R2063 gnd.n734 gnd.n733 585
R2064 gnd.n7441 gnd.n734 585
R2065 gnd.n7444 gnd.n7443 585
R2066 gnd.n7443 gnd.n7442 585
R2067 gnd.n731 gnd.n730 585
R2068 gnd.n730 gnd.n729 585
R2069 gnd.n7449 gnd.n7448 585
R2070 gnd.n7450 gnd.n7449 585
R2071 gnd.n728 gnd.n727 585
R2072 gnd.n7451 gnd.n728 585
R2073 gnd.n7454 gnd.n7453 585
R2074 gnd.n7453 gnd.n7452 585
R2075 gnd.n725 gnd.n724 585
R2076 gnd.n724 gnd.n723 585
R2077 gnd.n7459 gnd.n7458 585
R2078 gnd.n7460 gnd.n7459 585
R2079 gnd.n722 gnd.n721 585
R2080 gnd.n7461 gnd.n722 585
R2081 gnd.n7464 gnd.n7463 585
R2082 gnd.n7463 gnd.n7462 585
R2083 gnd.n719 gnd.n718 585
R2084 gnd.n718 gnd.n717 585
R2085 gnd.n7469 gnd.n7468 585
R2086 gnd.n7470 gnd.n7469 585
R2087 gnd.n716 gnd.n715 585
R2088 gnd.n7471 gnd.n716 585
R2089 gnd.n7474 gnd.n7473 585
R2090 gnd.n7473 gnd.n7472 585
R2091 gnd.n713 gnd.n712 585
R2092 gnd.n712 gnd.n711 585
R2093 gnd.n7479 gnd.n7478 585
R2094 gnd.n7480 gnd.n7479 585
R2095 gnd.n710 gnd.n709 585
R2096 gnd.n7481 gnd.n710 585
R2097 gnd.n7484 gnd.n7483 585
R2098 gnd.n7483 gnd.n7482 585
R2099 gnd.n707 gnd.n706 585
R2100 gnd.n706 gnd.n705 585
R2101 gnd.n7489 gnd.n7488 585
R2102 gnd.n7490 gnd.n7489 585
R2103 gnd.n704 gnd.n703 585
R2104 gnd.n7491 gnd.n704 585
R2105 gnd.n7494 gnd.n7493 585
R2106 gnd.n7493 gnd.n7492 585
R2107 gnd.n701 gnd.n700 585
R2108 gnd.n700 gnd.n699 585
R2109 gnd.n7500 gnd.n7499 585
R2110 gnd.n7501 gnd.n7500 585
R2111 gnd.n698 gnd.n697 585
R2112 gnd.n7502 gnd.n698 585
R2113 gnd.n7505 gnd.n7504 585
R2114 gnd.n7504 gnd.n7503 585
R2115 gnd.n7506 gnd.n695 585
R2116 gnd.n695 gnd.n694 585
R2117 gnd.n570 gnd.n569 585
R2118 gnd.n7713 gnd.n569 585
R2119 gnd.n7716 gnd.n7715 585
R2120 gnd.n7715 gnd.n7714 585
R2121 gnd.n573 gnd.n572 585
R2122 gnd.n7712 gnd.n573 585
R2123 gnd.n7710 gnd.n7709 585
R2124 gnd.n7711 gnd.n7710 585
R2125 gnd.n576 gnd.n575 585
R2126 gnd.n575 gnd.n574 585
R2127 gnd.n7705 gnd.n7704 585
R2128 gnd.n7704 gnd.n7703 585
R2129 gnd.n579 gnd.n578 585
R2130 gnd.n7702 gnd.n579 585
R2131 gnd.n7700 gnd.n7699 585
R2132 gnd.n7701 gnd.n7700 585
R2133 gnd.n582 gnd.n581 585
R2134 gnd.n581 gnd.n580 585
R2135 gnd.n7695 gnd.n7694 585
R2136 gnd.n7694 gnd.n7693 585
R2137 gnd.n585 gnd.n584 585
R2138 gnd.n7692 gnd.n585 585
R2139 gnd.n7690 gnd.n7689 585
R2140 gnd.n7691 gnd.n7690 585
R2141 gnd.n588 gnd.n587 585
R2142 gnd.n587 gnd.n586 585
R2143 gnd.n7685 gnd.n7684 585
R2144 gnd.n7684 gnd.n7683 585
R2145 gnd.n591 gnd.n590 585
R2146 gnd.n7682 gnd.n591 585
R2147 gnd.n7680 gnd.n7679 585
R2148 gnd.n7681 gnd.n7680 585
R2149 gnd.n594 gnd.n593 585
R2150 gnd.n593 gnd.n592 585
R2151 gnd.n7675 gnd.n7674 585
R2152 gnd.n7674 gnd.n7673 585
R2153 gnd.n597 gnd.n596 585
R2154 gnd.n7672 gnd.n597 585
R2155 gnd.n7670 gnd.n7669 585
R2156 gnd.n7671 gnd.n7670 585
R2157 gnd.n600 gnd.n599 585
R2158 gnd.n599 gnd.n598 585
R2159 gnd.n7665 gnd.n7664 585
R2160 gnd.n7664 gnd.n7663 585
R2161 gnd.n603 gnd.n602 585
R2162 gnd.n7662 gnd.n603 585
R2163 gnd.n7660 gnd.n7659 585
R2164 gnd.n7661 gnd.n7660 585
R2165 gnd.n606 gnd.n605 585
R2166 gnd.n605 gnd.n604 585
R2167 gnd.n7655 gnd.n7654 585
R2168 gnd.n7654 gnd.n7653 585
R2169 gnd.n609 gnd.n608 585
R2170 gnd.n7652 gnd.n609 585
R2171 gnd.n7650 gnd.n7649 585
R2172 gnd.n7651 gnd.n7650 585
R2173 gnd.n612 gnd.n611 585
R2174 gnd.n611 gnd.n610 585
R2175 gnd.n7645 gnd.n7644 585
R2176 gnd.n7644 gnd.n7643 585
R2177 gnd.n615 gnd.n614 585
R2178 gnd.n7642 gnd.n615 585
R2179 gnd.n7640 gnd.n7639 585
R2180 gnd.n7641 gnd.n7640 585
R2181 gnd.n618 gnd.n617 585
R2182 gnd.n617 gnd.n616 585
R2183 gnd.n7635 gnd.n7634 585
R2184 gnd.n7634 gnd.n7633 585
R2185 gnd.n621 gnd.n620 585
R2186 gnd.n7632 gnd.n621 585
R2187 gnd.n7630 gnd.n7629 585
R2188 gnd.n7631 gnd.n7630 585
R2189 gnd.n624 gnd.n623 585
R2190 gnd.n623 gnd.n622 585
R2191 gnd.n7625 gnd.n7624 585
R2192 gnd.n7624 gnd.n7623 585
R2193 gnd.n627 gnd.n626 585
R2194 gnd.n7622 gnd.n627 585
R2195 gnd.n7620 gnd.n7619 585
R2196 gnd.n7621 gnd.n7620 585
R2197 gnd.n630 gnd.n629 585
R2198 gnd.n629 gnd.n628 585
R2199 gnd.n7615 gnd.n7614 585
R2200 gnd.n7614 gnd.n7613 585
R2201 gnd.n633 gnd.n632 585
R2202 gnd.n7612 gnd.n633 585
R2203 gnd.n7610 gnd.n7609 585
R2204 gnd.n7611 gnd.n7610 585
R2205 gnd.n636 gnd.n635 585
R2206 gnd.n635 gnd.n634 585
R2207 gnd.n7605 gnd.n7604 585
R2208 gnd.n7604 gnd.n7603 585
R2209 gnd.n639 gnd.n638 585
R2210 gnd.n7602 gnd.n639 585
R2211 gnd.n7600 gnd.n7599 585
R2212 gnd.n7601 gnd.n7600 585
R2213 gnd.n642 gnd.n641 585
R2214 gnd.n641 gnd.n640 585
R2215 gnd.n7595 gnd.n7594 585
R2216 gnd.n7594 gnd.n7593 585
R2217 gnd.n645 gnd.n644 585
R2218 gnd.n7592 gnd.n645 585
R2219 gnd.n7590 gnd.n7589 585
R2220 gnd.n7591 gnd.n7590 585
R2221 gnd.n648 gnd.n647 585
R2222 gnd.n647 gnd.n646 585
R2223 gnd.n7585 gnd.n7584 585
R2224 gnd.n7584 gnd.n7583 585
R2225 gnd.n651 gnd.n650 585
R2226 gnd.n7582 gnd.n651 585
R2227 gnd.n7580 gnd.n7579 585
R2228 gnd.n7581 gnd.n7580 585
R2229 gnd.n654 gnd.n653 585
R2230 gnd.n653 gnd.n652 585
R2231 gnd.n7575 gnd.n7574 585
R2232 gnd.n7574 gnd.n7573 585
R2233 gnd.n657 gnd.n656 585
R2234 gnd.n7572 gnd.n657 585
R2235 gnd.n7570 gnd.n7569 585
R2236 gnd.n7571 gnd.n7570 585
R2237 gnd.n660 gnd.n659 585
R2238 gnd.n659 gnd.n658 585
R2239 gnd.n7565 gnd.n7564 585
R2240 gnd.n7564 gnd.n7563 585
R2241 gnd.n663 gnd.n662 585
R2242 gnd.n7562 gnd.n663 585
R2243 gnd.n7560 gnd.n7559 585
R2244 gnd.n7561 gnd.n7560 585
R2245 gnd.n666 gnd.n665 585
R2246 gnd.n665 gnd.n664 585
R2247 gnd.n7555 gnd.n7554 585
R2248 gnd.n7554 gnd.n7553 585
R2249 gnd.n669 gnd.n668 585
R2250 gnd.n7552 gnd.n669 585
R2251 gnd.n7550 gnd.n7549 585
R2252 gnd.n7551 gnd.n7550 585
R2253 gnd.n672 gnd.n671 585
R2254 gnd.n671 gnd.n670 585
R2255 gnd.n7545 gnd.n7544 585
R2256 gnd.n7544 gnd.n7543 585
R2257 gnd.n675 gnd.n674 585
R2258 gnd.n7542 gnd.n675 585
R2259 gnd.n7540 gnd.n7539 585
R2260 gnd.n7541 gnd.n7540 585
R2261 gnd.n678 gnd.n677 585
R2262 gnd.n677 gnd.n676 585
R2263 gnd.n7535 gnd.n7534 585
R2264 gnd.n7534 gnd.n7533 585
R2265 gnd.n681 gnd.n680 585
R2266 gnd.n7532 gnd.n681 585
R2267 gnd.n7530 gnd.n7529 585
R2268 gnd.n7531 gnd.n7530 585
R2269 gnd.n684 gnd.n683 585
R2270 gnd.n683 gnd.n682 585
R2271 gnd.n7525 gnd.n7524 585
R2272 gnd.n7524 gnd.n7523 585
R2273 gnd.n687 gnd.n686 585
R2274 gnd.n7522 gnd.n687 585
R2275 gnd.n7520 gnd.n7519 585
R2276 gnd.n7521 gnd.n7520 585
R2277 gnd.n690 gnd.n689 585
R2278 gnd.n689 gnd.n688 585
R2279 gnd.n7515 gnd.n7514 585
R2280 gnd.n7514 gnd.n7513 585
R2281 gnd.n693 gnd.n692 585
R2282 gnd.n7512 gnd.n693 585
R2283 gnd.n7510 gnd.n7509 585
R2284 gnd.n7511 gnd.n7510 585
R2285 gnd.n1545 gnd.n1544 585
R2286 gnd.n3361 gnd.n1545 585
R2287 gnd.n5109 gnd.n5108 585
R2288 gnd.n5108 gnd.n5107 585
R2289 gnd.n5110 gnd.n1540 585
R2290 gnd.n3218 gnd.n1540 585
R2291 gnd.n5112 gnd.n5111 585
R2292 gnd.n5113 gnd.n5112 585
R2293 gnd.n1524 gnd.n1523 585
R2294 gnd.n3208 gnd.n1524 585
R2295 gnd.n5121 gnd.n5120 585
R2296 gnd.n5120 gnd.n5119 585
R2297 gnd.n5122 gnd.n1519 585
R2298 gnd.n3201 gnd.n1519 585
R2299 gnd.n5124 gnd.n5123 585
R2300 gnd.n5125 gnd.n5124 585
R2301 gnd.n1504 gnd.n1503 585
R2302 gnd.n3193 gnd.n1504 585
R2303 gnd.n5133 gnd.n5132 585
R2304 gnd.n5132 gnd.n5131 585
R2305 gnd.n5134 gnd.n1499 585
R2306 gnd.n3186 gnd.n1499 585
R2307 gnd.n5136 gnd.n5135 585
R2308 gnd.n5137 gnd.n5136 585
R2309 gnd.n1483 gnd.n1482 585
R2310 gnd.n3125 gnd.n1483 585
R2311 gnd.n5145 gnd.n5144 585
R2312 gnd.n5144 gnd.n5143 585
R2313 gnd.n5146 gnd.n1478 585
R2314 gnd.n3118 gnd.n1478 585
R2315 gnd.n5148 gnd.n5147 585
R2316 gnd.n5149 gnd.n5148 585
R2317 gnd.n1463 gnd.n1462 585
R2318 gnd.n3114 gnd.n1463 585
R2319 gnd.n5157 gnd.n5156 585
R2320 gnd.n5156 gnd.n5155 585
R2321 gnd.n5158 gnd.n1458 585
R2322 gnd.n3142 gnd.n1458 585
R2323 gnd.n5160 gnd.n5159 585
R2324 gnd.n5161 gnd.n5160 585
R2325 gnd.n1442 gnd.n1441 585
R2326 gnd.n3107 gnd.n1442 585
R2327 gnd.n5169 gnd.n5168 585
R2328 gnd.n5168 gnd.n5167 585
R2329 gnd.n5170 gnd.n1437 585
R2330 gnd.n3099 gnd.n1437 585
R2331 gnd.n5172 gnd.n5171 585
R2332 gnd.n5173 gnd.n5172 585
R2333 gnd.n1423 gnd.n1422 585
R2334 gnd.n3093 gnd.n1423 585
R2335 gnd.n5181 gnd.n5180 585
R2336 gnd.n5180 gnd.n5179 585
R2337 gnd.n5182 gnd.n1417 585
R2338 gnd.n3085 gnd.n1417 585
R2339 gnd.n5184 gnd.n5183 585
R2340 gnd.n5185 gnd.n5184 585
R2341 gnd.n1418 gnd.n1416 585
R2342 gnd.n3054 gnd.n1416 585
R2343 gnd.n3036 gnd.n3035 585
R2344 gnd.n3035 gnd.n2784 585
R2345 gnd.n3037 gnd.n2793 585
R2346 gnd.n3046 gnd.n2793 585
R2347 gnd.n3039 gnd.n3038 585
R2348 gnd.n3040 gnd.n3039 585
R2349 gnd.n2801 gnd.n2800 585
R2350 gnd.n3024 gnd.n2800 585
R2351 gnd.n2878 gnd.n2877 585
R2352 gnd.n2881 gnd.n2878 585
R2353 gnd.n1395 gnd.n1394 585
R2354 gnd.n1399 gnd.n1395 585
R2355 gnd.n5194 gnd.n5193 585
R2356 gnd.n5193 gnd.n5192 585
R2357 gnd.n5195 gnd.n1390 585
R2358 gnd.n1390 gnd.n1389 585
R2359 gnd.n5197 gnd.n5196 585
R2360 gnd.n5198 gnd.n5197 585
R2361 gnd.n1377 gnd.n1376 585
R2362 gnd.n1386 gnd.n1377 585
R2363 gnd.n5206 gnd.n5205 585
R2364 gnd.n5205 gnd.n5204 585
R2365 gnd.n5207 gnd.n1372 585
R2366 gnd.n1372 gnd.n1371 585
R2367 gnd.n5209 gnd.n5208 585
R2368 gnd.n5210 gnd.n5209 585
R2369 gnd.n1358 gnd.n1357 585
R2370 gnd.n1361 gnd.n1358 585
R2371 gnd.n5218 gnd.n5217 585
R2372 gnd.n5217 gnd.n5216 585
R2373 gnd.n5219 gnd.n1353 585
R2374 gnd.n1353 gnd.n1352 585
R2375 gnd.n5221 gnd.n5220 585
R2376 gnd.n5222 gnd.n5221 585
R2377 gnd.n1339 gnd.n1338 585
R2378 gnd.n1349 gnd.n1339 585
R2379 gnd.n5230 gnd.n5229 585
R2380 gnd.n5229 gnd.n5228 585
R2381 gnd.n5231 gnd.n1334 585
R2382 gnd.n1334 gnd.n1333 585
R2383 gnd.n5233 gnd.n5232 585
R2384 gnd.n5234 gnd.n5233 585
R2385 gnd.n1320 gnd.n1319 585
R2386 gnd.n1323 gnd.n1320 585
R2387 gnd.n5242 gnd.n5241 585
R2388 gnd.n5241 gnd.n5240 585
R2389 gnd.n5243 gnd.n1315 585
R2390 gnd.n1315 gnd.n1314 585
R2391 gnd.n5245 gnd.n5244 585
R2392 gnd.n5246 gnd.n5245 585
R2393 gnd.n1301 gnd.n1300 585
R2394 gnd.n1311 gnd.n1301 585
R2395 gnd.n5254 gnd.n5253 585
R2396 gnd.n5253 gnd.n5252 585
R2397 gnd.n5255 gnd.n1296 585
R2398 gnd.n1296 gnd.n1295 585
R2399 gnd.n5257 gnd.n5256 585
R2400 gnd.n5258 gnd.n5257 585
R2401 gnd.n1282 gnd.n1281 585
R2402 gnd.n1285 gnd.n1282 585
R2403 gnd.n5266 gnd.n5265 585
R2404 gnd.n5265 gnd.n5264 585
R2405 gnd.n5267 gnd.n1275 585
R2406 gnd.n1275 gnd.n1273 585
R2407 gnd.n5269 gnd.n5268 585
R2408 gnd.n5270 gnd.n5269 585
R2409 gnd.n1277 gnd.n1274 585
R2410 gnd.n1274 gnd.n1270 585
R2411 gnd.n1276 gnd.n1261 585
R2412 gnd.n5276 gnd.n1261 585
R2413 gnd.n2913 gnd.n1255 585
R2414 gnd.n2913 gnd.n1186 585
R2415 gnd.n2915 gnd.n2914 585
R2416 gnd.n2917 gnd.n2916 585
R2417 gnd.n2919 gnd.n2918 585
R2418 gnd.n2923 gnd.n2911 585
R2419 gnd.n2925 gnd.n2924 585
R2420 gnd.n2927 gnd.n2926 585
R2421 gnd.n2929 gnd.n2928 585
R2422 gnd.n2933 gnd.n2909 585
R2423 gnd.n2935 gnd.n2934 585
R2424 gnd.n2937 gnd.n2936 585
R2425 gnd.n2939 gnd.n2938 585
R2426 gnd.n2943 gnd.n2907 585
R2427 gnd.n2945 gnd.n2944 585
R2428 gnd.n2947 gnd.n2946 585
R2429 gnd.n2949 gnd.n2948 585
R2430 gnd.n2904 gnd.n2903 585
R2431 gnd.n2953 gnd.n2905 585
R2432 gnd.n2954 gnd.n2900 585
R2433 gnd.n2955 gnd.n1185 585
R2434 gnd.n5400 gnd.n1185 585
R2435 gnd.n3364 gnd.n3363 585
R2436 gnd.n3289 gnd.n2552 585
R2437 gnd.n3291 gnd.n3290 585
R2438 gnd.n3277 gnd.n3276 585
R2439 gnd.n3298 gnd.n3275 585
R2440 gnd.n3299 gnd.n3274 585
R2441 gnd.n3273 gnd.n3267 585
R2442 gnd.n3306 gnd.n3266 585
R2443 gnd.n3307 gnd.n3265 585
R2444 gnd.n3257 gnd.n3256 585
R2445 gnd.n3314 gnd.n3255 585
R2446 gnd.n3315 gnd.n3254 585
R2447 gnd.n3253 gnd.n3247 585
R2448 gnd.n3322 gnd.n3246 585
R2449 gnd.n3323 gnd.n3245 585
R2450 gnd.n3237 gnd.n3236 585
R2451 gnd.n3330 gnd.n3235 585
R2452 gnd.n3331 gnd.n3234 585
R2453 gnd.n3233 gnd.n1557 585
R2454 gnd.n5099 gnd.n1557 585
R2455 gnd.n3362 gnd.n2553 585
R2456 gnd.n3362 gnd.n3361 585
R2457 gnd.n2738 gnd.n1548 585
R2458 gnd.n5107 gnd.n1548 585
R2459 gnd.n3217 gnd.n3216 585
R2460 gnd.n3218 gnd.n3217 585
R2461 gnd.n2737 gnd.n1538 585
R2462 gnd.n5113 gnd.n1538 585
R2463 gnd.n3210 gnd.n3209 585
R2464 gnd.n3209 gnd.n3208 585
R2465 gnd.n2740 gnd.n1527 585
R2466 gnd.n5119 gnd.n1527 585
R2467 gnd.n3200 gnd.n3199 585
R2468 gnd.n3201 gnd.n3200 585
R2469 gnd.n2742 gnd.n1517 585
R2470 gnd.n5125 gnd.n1517 585
R2471 gnd.n3195 gnd.n3194 585
R2472 gnd.n3194 gnd.n3193 585
R2473 gnd.n2744 gnd.n1506 585
R2474 gnd.n5131 gnd.n1506 585
R2475 gnd.n3128 gnd.n2746 585
R2476 gnd.n3186 gnd.n2746 585
R2477 gnd.n3129 gnd.n1497 585
R2478 gnd.n5137 gnd.n1497 585
R2479 gnd.n3130 gnd.n3126 585
R2480 gnd.n3126 gnd.n3125 585
R2481 gnd.n2765 gnd.n1486 585
R2482 gnd.n5143 gnd.n1486 585
R2483 gnd.n3134 gnd.n2764 585
R2484 gnd.n3118 gnd.n2764 585
R2485 gnd.n3135 gnd.n1476 585
R2486 gnd.n5149 gnd.n1476 585
R2487 gnd.n3136 gnd.n2763 585
R2488 gnd.n3114 gnd.n2763 585
R2489 gnd.n2760 gnd.n1465 585
R2490 gnd.n5155 gnd.n1465 585
R2491 gnd.n3141 gnd.n3140 585
R2492 gnd.n3142 gnd.n3141 585
R2493 gnd.n2759 gnd.n1456 585
R2494 gnd.n5161 gnd.n1456 585
R2495 gnd.n3106 gnd.n3105 585
R2496 gnd.n3107 gnd.n3106 585
R2497 gnd.n2769 gnd.n1445 585
R2498 gnd.n5167 gnd.n1445 585
R2499 gnd.n3101 gnd.n3100 585
R2500 gnd.n3100 gnd.n3099 585
R2501 gnd.n2771 gnd.n1435 585
R2502 gnd.n5173 gnd.n1435 585
R2503 gnd.n3092 gnd.n3091 585
R2504 gnd.n3093 gnd.n3092 585
R2505 gnd.n2774 gnd.n1425 585
R2506 gnd.n5179 gnd.n1425 585
R2507 gnd.n3087 gnd.n3086 585
R2508 gnd.n3086 gnd.n3085 585
R2509 gnd.n2776 gnd.n1414 585
R2510 gnd.n5185 gnd.n1414 585
R2511 gnd.n3053 gnd.n3052 585
R2512 gnd.n3054 gnd.n3053 585
R2513 gnd.n2787 gnd.n2786 585
R2514 gnd.n2786 gnd.n2784 585
R2515 gnd.n3048 gnd.n3047 585
R2516 gnd.n3047 gnd.n3046 585
R2517 gnd.n2790 gnd.n2789 585
R2518 gnd.n3040 gnd.n2790 585
R2519 gnd.n3023 gnd.n3022 585
R2520 gnd.n3024 gnd.n3023 585
R2521 gnd.n2883 gnd.n2882 585
R2522 gnd.n2882 gnd.n2881 585
R2523 gnd.n3018 gnd.n3017 585
R2524 gnd.n3017 gnd.n1399 585
R2525 gnd.n3016 gnd.n1398 585
R2526 gnd.n5192 gnd.n1398 585
R2527 gnd.n3015 gnd.n3014 585
R2528 gnd.n3014 gnd.n1389 585
R2529 gnd.n2885 gnd.n1388 585
R2530 gnd.n5198 gnd.n1388 585
R2531 gnd.n3010 gnd.n3009 585
R2532 gnd.n3009 gnd.n1386 585
R2533 gnd.n3008 gnd.n1379 585
R2534 gnd.n5204 gnd.n1379 585
R2535 gnd.n3007 gnd.n3006 585
R2536 gnd.n3006 gnd.n1371 585
R2537 gnd.n2887 gnd.n1370 585
R2538 gnd.n5210 gnd.n1370 585
R2539 gnd.n3002 gnd.n3001 585
R2540 gnd.n3001 gnd.n1361 585
R2541 gnd.n3000 gnd.n1360 585
R2542 gnd.n5216 gnd.n1360 585
R2543 gnd.n2999 gnd.n2998 585
R2544 gnd.n2998 gnd.n1352 585
R2545 gnd.n2889 gnd.n1351 585
R2546 gnd.n5222 gnd.n1351 585
R2547 gnd.n2994 gnd.n2993 585
R2548 gnd.n2993 gnd.n1349 585
R2549 gnd.n2992 gnd.n1341 585
R2550 gnd.n5228 gnd.n1341 585
R2551 gnd.n2991 gnd.n2990 585
R2552 gnd.n2990 gnd.n1333 585
R2553 gnd.n2891 gnd.n1332 585
R2554 gnd.n5234 gnd.n1332 585
R2555 gnd.n2986 gnd.n2985 585
R2556 gnd.n2985 gnd.n1323 585
R2557 gnd.n2984 gnd.n1322 585
R2558 gnd.n5240 gnd.n1322 585
R2559 gnd.n2983 gnd.n2982 585
R2560 gnd.n2982 gnd.n1314 585
R2561 gnd.n2893 gnd.n1313 585
R2562 gnd.n5246 gnd.n1313 585
R2563 gnd.n2978 gnd.n2977 585
R2564 gnd.n2977 gnd.n1311 585
R2565 gnd.n2976 gnd.n1303 585
R2566 gnd.n5252 gnd.n1303 585
R2567 gnd.n2975 gnd.n2974 585
R2568 gnd.n2974 gnd.n1295 585
R2569 gnd.n2895 gnd.n1294 585
R2570 gnd.n5258 gnd.n1294 585
R2571 gnd.n2970 gnd.n2969 585
R2572 gnd.n2969 gnd.n1285 585
R2573 gnd.n2968 gnd.n1284 585
R2574 gnd.n5264 gnd.n1284 585
R2575 gnd.n2967 gnd.n2966 585
R2576 gnd.n2966 gnd.n1273 585
R2577 gnd.n2897 gnd.n1272 585
R2578 gnd.n5270 gnd.n1272 585
R2579 gnd.n2962 gnd.n2961 585
R2580 gnd.n2961 gnd.n1270 585
R2581 gnd.n2960 gnd.n1260 585
R2582 gnd.n5276 gnd.n1260 585
R2583 gnd.n2959 gnd.n2958 585
R2584 gnd.n2958 gnd.n1186 585
R2585 gnd.n6878 gnd.n6877 585
R2586 gnd.n6877 gnd.n6876 585
R2587 gnd.n6879 gnd.n1139 585
R2588 gnd.n6786 gnd.n1139 585
R2589 gnd.n6881 gnd.n6880 585
R2590 gnd.n6882 gnd.n6881 585
R2591 gnd.n1140 gnd.n1138 585
R2592 gnd.n5761 gnd.n1138 585
R2593 gnd.n6778 gnd.n6777 585
R2594 gnd.n6779 gnd.n6778 585
R2595 gnd.n5492 gnd.n5491 585
R2596 gnd.n6759 gnd.n5491 585
R2597 gnd.n6752 gnd.n6751 585
R2598 gnd.n6751 gnd.n5768 585
R2599 gnd.n6750 gnd.n5772 585
R2600 gnd.n6750 gnd.n6749 585
R2601 gnd.n6735 gnd.n5773 585
R2602 gnd.n5788 gnd.n5773 585
R2603 gnd.n6737 gnd.n6736 585
R2604 gnd.n6738 gnd.n6737 585
R2605 gnd.n5782 gnd.n5781 585
R2606 gnd.n6716 gnd.n5781 585
R2607 gnd.n6707 gnd.n6706 585
R2608 gnd.n6706 gnd.n5795 585
R2609 gnd.n6705 gnd.n5799 585
R2610 gnd.n6705 gnd.n6704 585
R2611 gnd.n6690 gnd.n5800 585
R2612 gnd.n5808 gnd.n5800 585
R2613 gnd.n6692 gnd.n6691 585
R2614 gnd.n6693 gnd.n6692 585
R2615 gnd.n5811 gnd.n5810 585
R2616 gnd.n5818 gnd.n5810 585
R2617 gnd.n6668 gnd.n6667 585
R2618 gnd.n6669 gnd.n6668 585
R2619 gnd.n5829 gnd.n5828 585
R2620 gnd.n6659 gnd.n5828 585
R2621 gnd.n6646 gnd.n5845 585
R2622 gnd.n5845 gnd.n5837 585
R2623 gnd.n6648 gnd.n6647 585
R2624 gnd.n6649 gnd.n6648 585
R2625 gnd.n5846 gnd.n5844 585
R2626 gnd.n5850 gnd.n5844 585
R2627 gnd.n6627 gnd.n6626 585
R2628 gnd.n6628 gnd.n6627 585
R2629 gnd.n5862 gnd.n5861 585
R2630 gnd.n5861 gnd.n5857 585
R2631 gnd.n6617 gnd.n6616 585
R2632 gnd.n6618 gnd.n6617 585
R2633 gnd.n5870 gnd.n5869 585
R2634 gnd.n5874 gnd.n5869 585
R2635 gnd.n6595 gnd.n5886 585
R2636 gnd.n6228 gnd.n5886 585
R2637 gnd.n6597 gnd.n6596 585
R2638 gnd.n6598 gnd.n6597 585
R2639 gnd.n5887 gnd.n5885 585
R2640 gnd.n5885 gnd.n5881 585
R2641 gnd.n6586 gnd.n6585 585
R2642 gnd.n6587 gnd.n6586 585
R2643 gnd.n5895 gnd.n5894 585
R2644 gnd.n6236 gnd.n5894 585
R2645 gnd.n6564 gnd.n5911 585
R2646 gnd.n5911 gnd.n5899 585
R2647 gnd.n6566 gnd.n6565 585
R2648 gnd.n6567 gnd.n6566 585
R2649 gnd.n5912 gnd.n5910 585
R2650 gnd.n5910 gnd.n5906 585
R2651 gnd.n6555 gnd.n6554 585
R2652 gnd.n6556 gnd.n6555 585
R2653 gnd.n5920 gnd.n5919 585
R2654 gnd.n5925 gnd.n5919 585
R2655 gnd.n6533 gnd.n5937 585
R2656 gnd.n5937 gnd.n5924 585
R2657 gnd.n6535 gnd.n6534 585
R2658 gnd.n6536 gnd.n6535 585
R2659 gnd.n5938 gnd.n5936 585
R2660 gnd.n5936 gnd.n5932 585
R2661 gnd.n6524 gnd.n6523 585
R2662 gnd.n6525 gnd.n6524 585
R2663 gnd.n5945 gnd.n5944 585
R2664 gnd.n5950 gnd.n5944 585
R2665 gnd.n6502 gnd.n5963 585
R2666 gnd.n5963 gnd.n5949 585
R2667 gnd.n6504 gnd.n6503 585
R2668 gnd.n6505 gnd.n6504 585
R2669 gnd.n5964 gnd.n5962 585
R2670 gnd.n5962 gnd.n5958 585
R2671 gnd.n6493 gnd.n6492 585
R2672 gnd.n6494 gnd.n6493 585
R2673 gnd.n5971 gnd.n5970 585
R2674 gnd.n5976 gnd.n5970 585
R2675 gnd.n6471 gnd.n5989 585
R2676 gnd.n5989 gnd.n5975 585
R2677 gnd.n6473 gnd.n6472 585
R2678 gnd.n6474 gnd.n6473 585
R2679 gnd.n5990 gnd.n5988 585
R2680 gnd.n5988 gnd.n5984 585
R2681 gnd.n6462 gnd.n6461 585
R2682 gnd.n6463 gnd.n6462 585
R2683 gnd.n5998 gnd.n5997 585
R2684 gnd.n6352 gnd.n5997 585
R2685 gnd.n6440 gnd.n6014 585
R2686 gnd.n6014 gnd.n6002 585
R2687 gnd.n6442 gnd.n6441 585
R2688 gnd.n6443 gnd.n6442 585
R2689 gnd.n6015 gnd.n6013 585
R2690 gnd.n6013 gnd.n6009 585
R2691 gnd.n6431 gnd.n6430 585
R2692 gnd.n6432 gnd.n6431 585
R2693 gnd.n6022 gnd.n6021 585
R2694 gnd.n6021 gnd.n6019 585
R2695 gnd.n6425 gnd.n6424 585
R2696 gnd.n6424 gnd.n6423 585
R2697 gnd.n6026 gnd.n6025 585
R2698 gnd.n6034 gnd.n6026 585
R2699 gnd.n6187 gnd.n6186 585
R2700 gnd.n6188 gnd.n6187 585
R2701 gnd.n6036 gnd.n6035 585
R2702 gnd.n6035 gnd.n6033 585
R2703 gnd.n6182 gnd.n6181 585
R2704 gnd.n6181 gnd.n6180 585
R2705 gnd.n6039 gnd.n6038 585
R2706 gnd.n6040 gnd.n6039 585
R2707 gnd.n6171 gnd.n6170 585
R2708 gnd.n6172 gnd.n6171 585
R2709 gnd.n6048 gnd.n6047 585
R2710 gnd.n6047 gnd.n6046 585
R2711 gnd.n6166 gnd.n6165 585
R2712 gnd.n6165 gnd.n6164 585
R2713 gnd.n6051 gnd.n6050 585
R2714 gnd.n6052 gnd.n6051 585
R2715 gnd.n6155 gnd.n6154 585
R2716 gnd.n6156 gnd.n6155 585
R2717 gnd.n6151 gnd.n6058 585
R2718 gnd.n6150 gnd.n6149 585
R2719 gnd.n6147 gnd.n6060 585
R2720 gnd.n6147 gnd.n6057 585
R2721 gnd.n6146 gnd.n6145 585
R2722 gnd.n6144 gnd.n6143 585
R2723 gnd.n6142 gnd.n6065 585
R2724 gnd.n6140 gnd.n6139 585
R2725 gnd.n6138 gnd.n6066 585
R2726 gnd.n6137 gnd.n6136 585
R2727 gnd.n6134 gnd.n6071 585
R2728 gnd.n6132 gnd.n6131 585
R2729 gnd.n6130 gnd.n6072 585
R2730 gnd.n6129 gnd.n6128 585
R2731 gnd.n6126 gnd.n6077 585
R2732 gnd.n6124 gnd.n6123 585
R2733 gnd.n6122 gnd.n6078 585
R2734 gnd.n6121 gnd.n6120 585
R2735 gnd.n6118 gnd.n6083 585
R2736 gnd.n6116 gnd.n6115 585
R2737 gnd.n6114 gnd.n6084 585
R2738 gnd.n6113 gnd.n6112 585
R2739 gnd.n6110 gnd.n6089 585
R2740 gnd.n6108 gnd.n6107 585
R2741 gnd.n6105 gnd.n6090 585
R2742 gnd.n6104 gnd.n6103 585
R2743 gnd.n6101 gnd.n6099 585
R2744 gnd.n6097 gnd.n6056 585
R2745 gnd.n6794 gnd.n6793 585
R2746 gnd.n6795 gnd.n5479 585
R2747 gnd.n6797 gnd.n6796 585
R2748 gnd.n6799 gnd.n5478 585
R2749 gnd.n6801 gnd.n6800 585
R2750 gnd.n6802 gnd.n5469 585
R2751 gnd.n6804 gnd.n6803 585
R2752 gnd.n6806 gnd.n5467 585
R2753 gnd.n6808 gnd.n6807 585
R2754 gnd.n6809 gnd.n5462 585
R2755 gnd.n6811 gnd.n6810 585
R2756 gnd.n6813 gnd.n5460 585
R2757 gnd.n6815 gnd.n6814 585
R2758 gnd.n6816 gnd.n5455 585
R2759 gnd.n6818 gnd.n6817 585
R2760 gnd.n6820 gnd.n5453 585
R2761 gnd.n6822 gnd.n6821 585
R2762 gnd.n6823 gnd.n5448 585
R2763 gnd.n6825 gnd.n6824 585
R2764 gnd.n6827 gnd.n5446 585
R2765 gnd.n6829 gnd.n6828 585
R2766 gnd.n6830 gnd.n5441 585
R2767 gnd.n6832 gnd.n6831 585
R2768 gnd.n6834 gnd.n5439 585
R2769 gnd.n6836 gnd.n6835 585
R2770 gnd.n6837 gnd.n5437 585
R2771 gnd.n6838 gnd.n1144 585
R2772 gnd.n5401 gnd.n1144 585
R2773 gnd.n6789 gnd.n1146 585
R2774 gnd.n6876 gnd.n1146 585
R2775 gnd.n6788 gnd.n6787 585
R2776 gnd.n6787 gnd.n6786 585
R2777 gnd.n6785 gnd.n1136 585
R2778 gnd.n6882 gnd.n1136 585
R2779 gnd.n5488 gnd.n5484 585
R2780 gnd.n5761 gnd.n5488 585
R2781 gnd.n6781 gnd.n6780 585
R2782 gnd.n6780 gnd.n6779 585
R2783 gnd.n5487 gnd.n5486 585
R2784 gnd.n6759 gnd.n5487 585
R2785 gnd.n6745 gnd.n5776 585
R2786 gnd.n5776 gnd.n5768 585
R2787 gnd.n6747 gnd.n6746 585
R2788 gnd.n6749 gnd.n6747 585
R2789 gnd.n5777 gnd.n5775 585
R2790 gnd.n5788 gnd.n5775 585
R2791 gnd.n6740 gnd.n6739 585
R2792 gnd.n6739 gnd.n6738 585
R2793 gnd.n5780 gnd.n5779 585
R2794 gnd.n6716 gnd.n5780 585
R2795 gnd.n6700 gnd.n5803 585
R2796 gnd.n5803 gnd.n5795 585
R2797 gnd.n6702 gnd.n6701 585
R2798 gnd.n6704 gnd.n6702 585
R2799 gnd.n5804 gnd.n5802 585
R2800 gnd.n5808 gnd.n5802 585
R2801 gnd.n6695 gnd.n6694 585
R2802 gnd.n6694 gnd.n6693 585
R2803 gnd.n5807 gnd.n5806 585
R2804 gnd.n5818 gnd.n5807 585
R2805 gnd.n6656 gnd.n5826 585
R2806 gnd.n6669 gnd.n5826 585
R2807 gnd.n6658 gnd.n6657 585
R2808 gnd.n6659 gnd.n6658 585
R2809 gnd.n5839 gnd.n5838 585
R2810 gnd.n5838 gnd.n5837 585
R2811 gnd.n6651 gnd.n6650 585
R2812 gnd.n6650 gnd.n6649 585
R2813 gnd.n5842 gnd.n5841 585
R2814 gnd.n5850 gnd.n5842 585
R2815 gnd.n6222 gnd.n5859 585
R2816 gnd.n6628 gnd.n5859 585
R2817 gnd.n6224 gnd.n6223 585
R2818 gnd.n6223 gnd.n5857 585
R2819 gnd.n6225 gnd.n5868 585
R2820 gnd.n6618 gnd.n5868 585
R2821 gnd.n6227 gnd.n6226 585
R2822 gnd.n6227 gnd.n5874 585
R2823 gnd.n6230 gnd.n6229 585
R2824 gnd.n6229 gnd.n6228 585
R2825 gnd.n6231 gnd.n5883 585
R2826 gnd.n6598 gnd.n5883 585
R2827 gnd.n6233 gnd.n6232 585
R2828 gnd.n6232 gnd.n5881 585
R2829 gnd.n6234 gnd.n5893 585
R2830 gnd.n6587 gnd.n5893 585
R2831 gnd.n6237 gnd.n6235 585
R2832 gnd.n6237 gnd.n6236 585
R2833 gnd.n6239 gnd.n6238 585
R2834 gnd.n6238 gnd.n5899 585
R2835 gnd.n6240 gnd.n5908 585
R2836 gnd.n6567 gnd.n5908 585
R2837 gnd.n6243 gnd.n6242 585
R2838 gnd.n6242 gnd.n5906 585
R2839 gnd.n6244 gnd.n5918 585
R2840 gnd.n6556 gnd.n5918 585
R2841 gnd.n6247 gnd.n6246 585
R2842 gnd.n6246 gnd.n5925 585
R2843 gnd.n6245 gnd.n6212 585
R2844 gnd.n6245 gnd.n5924 585
R2845 gnd.n6331 gnd.n5934 585
R2846 gnd.n6536 gnd.n5934 585
R2847 gnd.n6333 gnd.n6332 585
R2848 gnd.n6332 gnd.n5932 585
R2849 gnd.n6334 gnd.n5943 585
R2850 gnd.n6525 gnd.n5943 585
R2851 gnd.n6336 gnd.n6335 585
R2852 gnd.n6336 gnd.n5950 585
R2853 gnd.n6338 gnd.n6337 585
R2854 gnd.n6337 gnd.n5949 585
R2855 gnd.n6339 gnd.n5960 585
R2856 gnd.n6505 gnd.n5960 585
R2857 gnd.n6341 gnd.n6340 585
R2858 gnd.n6340 gnd.n5958 585
R2859 gnd.n6342 gnd.n5969 585
R2860 gnd.n6494 gnd.n5969 585
R2861 gnd.n6344 gnd.n6343 585
R2862 gnd.n6344 gnd.n5976 585
R2863 gnd.n6346 gnd.n6345 585
R2864 gnd.n6345 gnd.n5975 585
R2865 gnd.n6347 gnd.n5986 585
R2866 gnd.n6474 gnd.n5986 585
R2867 gnd.n6349 gnd.n6348 585
R2868 gnd.n6348 gnd.n5984 585
R2869 gnd.n6350 gnd.n5996 585
R2870 gnd.n6463 gnd.n5996 585
R2871 gnd.n6353 gnd.n6351 585
R2872 gnd.n6353 gnd.n6352 585
R2873 gnd.n6355 gnd.n6354 585
R2874 gnd.n6354 gnd.n6002 585
R2875 gnd.n6356 gnd.n6011 585
R2876 gnd.n6443 gnd.n6011 585
R2877 gnd.n6358 gnd.n6357 585
R2878 gnd.n6357 gnd.n6009 585
R2879 gnd.n6359 gnd.n6020 585
R2880 gnd.n6432 gnd.n6020 585
R2881 gnd.n6360 gnd.n6028 585
R2882 gnd.n6028 gnd.n6019 585
R2883 gnd.n6362 gnd.n6361 585
R2884 gnd.n6423 gnd.n6362 585
R2885 gnd.n6029 gnd.n6027 585
R2886 gnd.n6034 gnd.n6027 585
R2887 gnd.n6190 gnd.n6189 585
R2888 gnd.n6189 gnd.n6188 585
R2889 gnd.n6032 gnd.n6031 585
R2890 gnd.n6033 gnd.n6032 585
R2891 gnd.n6179 gnd.n6178 585
R2892 gnd.n6180 gnd.n6179 585
R2893 gnd.n6042 gnd.n6041 585
R2894 gnd.n6041 gnd.n6040 585
R2895 gnd.n6174 gnd.n6173 585
R2896 gnd.n6173 gnd.n6172 585
R2897 gnd.n6045 gnd.n6044 585
R2898 gnd.n6046 gnd.n6045 585
R2899 gnd.n6163 gnd.n6162 585
R2900 gnd.n6164 gnd.n6163 585
R2901 gnd.n6054 gnd.n6053 585
R2902 gnd.n6053 gnd.n6052 585
R2903 gnd.n6158 gnd.n6157 585
R2904 gnd.n6157 gnd.n6156 585
R2905 gnd.n247 gnd.n246 585
R2906 gnd.n250 gnd.n247 585
R2907 gnd.n8013 gnd.n8012 585
R2908 gnd.n8012 gnd.n8011 585
R2909 gnd.n8014 gnd.n242 585
R2910 gnd.n242 gnd.n241 585
R2911 gnd.n8016 gnd.n8015 585
R2912 gnd.n8017 gnd.n8016 585
R2913 gnd.n227 gnd.n226 585
R2914 gnd.n231 gnd.n227 585
R2915 gnd.n8025 gnd.n8024 585
R2916 gnd.n8024 gnd.n8023 585
R2917 gnd.n8026 gnd.n222 585
R2918 gnd.n228 gnd.n222 585
R2919 gnd.n8028 gnd.n8027 585
R2920 gnd.n8029 gnd.n8028 585
R2921 gnd.n208 gnd.n207 585
R2922 gnd.n211 gnd.n208 585
R2923 gnd.n8037 gnd.n8036 585
R2924 gnd.n8036 gnd.n8035 585
R2925 gnd.n8038 gnd.n203 585
R2926 gnd.n203 gnd.n202 585
R2927 gnd.n8040 gnd.n8039 585
R2928 gnd.n8041 gnd.n8040 585
R2929 gnd.n188 gnd.n187 585
R2930 gnd.n199 gnd.n188 585
R2931 gnd.n8049 gnd.n8048 585
R2932 gnd.n8048 gnd.n8047 585
R2933 gnd.n8050 gnd.n183 585
R2934 gnd.n189 gnd.n183 585
R2935 gnd.n8052 gnd.n8051 585
R2936 gnd.n8053 gnd.n8052 585
R2937 gnd.n170 gnd.n169 585
R2938 gnd.n173 gnd.n170 585
R2939 gnd.n8061 gnd.n8060 585
R2940 gnd.n8060 gnd.n8059 585
R2941 gnd.n8062 gnd.n165 585
R2942 gnd.n165 gnd.n164 585
R2943 gnd.n8064 gnd.n8063 585
R2944 gnd.n8065 gnd.n8064 585
R2945 gnd.n150 gnd.n149 585
R2946 gnd.n161 gnd.n150 585
R2947 gnd.n8073 gnd.n8072 585
R2948 gnd.n8072 gnd.n8071 585
R2949 gnd.n8074 gnd.n145 585
R2950 gnd.n151 gnd.n145 585
R2951 gnd.n8076 gnd.n8075 585
R2952 gnd.n8077 gnd.n8076 585
R2953 gnd.n133 gnd.n132 585
R2954 gnd.n136 gnd.n133 585
R2955 gnd.n8085 gnd.n8084 585
R2956 gnd.n8084 gnd.n8083 585
R2957 gnd.n8086 gnd.n127 585
R2958 gnd.n127 gnd.n125 585
R2959 gnd.n8088 gnd.n8087 585
R2960 gnd.n8089 gnd.n8088 585
R2961 gnd.n128 gnd.n126 585
R2962 gnd.n126 gnd.n122 585
R2963 gnd.n7827 gnd.n7826 585
R2964 gnd.n7826 gnd.n107 585
R2965 gnd.n7825 gnd.n108 585
R2966 gnd.n8097 gnd.n108 585
R2967 gnd.n7824 gnd.n7823 585
R2968 gnd.n7823 gnd.n7822 585
R2969 gnd.n490 gnd.n488 585
R2970 gnd.n7808 gnd.n490 585
R2971 gnd.n7815 gnd.n7814 585
R2972 gnd.n7814 gnd.n7813 585
R2973 gnd.n496 gnd.n495 585
R2974 gnd.n7803 gnd.n496 585
R2975 gnd.n7786 gnd.n7785 585
R2976 gnd.n7785 gnd.n7784 585
R2977 gnd.n7787 gnd.n512 585
R2978 gnd.n7795 gnd.n512 585
R2979 gnd.n7789 gnd.n7788 585
R2980 gnd.n7790 gnd.n7789 585
R2981 gnd.n518 gnd.n517 585
R2982 gnd.n7776 gnd.n517 585
R2983 gnd.n7752 gnd.n7751 585
R2984 gnd.n7751 gnd.n7750 585
R2985 gnd.n7753 gnd.n535 585
R2986 gnd.n7768 gnd.n535 585
R2987 gnd.n7754 gnd.n546 585
R2988 gnd.n7744 gnd.n546 585
R2989 gnd.n7756 gnd.n7755 585
R2990 gnd.n7757 gnd.n7756 585
R2991 gnd.n547 gnd.n545 585
R2992 gnd.n2045 gnd.n545 585
R2993 gnd.n4656 gnd.n2038 585
R2994 gnd.n4652 gnd.n2038 585
R2995 gnd.n4658 gnd.n4657 585
R2996 gnd.n4659 gnd.n4658 585
R2997 gnd.n2022 gnd.n2021 585
R2998 gnd.n4640 gnd.n2022 585
R2999 gnd.n4667 gnd.n4666 585
R3000 gnd.n4666 gnd.n4665 585
R3001 gnd.n4668 gnd.n2017 585
R3002 gnd.n4624 gnd.n2017 585
R3003 gnd.n4670 gnd.n4669 585
R3004 gnd.n4671 gnd.n4670 585
R3005 gnd.n2001 gnd.n2000 585
R3006 gnd.n4615 gnd.n2001 585
R3007 gnd.n4679 gnd.n4678 585
R3008 gnd.n4678 gnd.n4677 585
R3009 gnd.n4680 gnd.n1996 585
R3010 gnd.n4607 gnd.n1996 585
R3011 gnd.n4682 gnd.n4681 585
R3012 gnd.n4683 gnd.n4682 585
R3013 gnd.n1981 gnd.n1980 585
R3014 gnd.n4601 gnd.n1981 585
R3015 gnd.n4691 gnd.n4690 585
R3016 gnd.n4690 gnd.n4689 585
R3017 gnd.n4692 gnd.n1976 585
R3018 gnd.n4593 gnd.n1976 585
R3019 gnd.n4694 gnd.n4693 585
R3020 gnd.n4695 gnd.n4694 585
R3021 gnd.n1960 gnd.n1959 585
R3022 gnd.n4587 gnd.n1960 585
R3023 gnd.n4703 gnd.n4702 585
R3024 gnd.n4702 gnd.n4701 585
R3025 gnd.n4704 gnd.n1954 585
R3026 gnd.n4579 gnd.n1954 585
R3027 gnd.n4706 gnd.n4705 585
R3028 gnd.n4707 gnd.n4706 585
R3029 gnd.n1955 gnd.n1938 585
R3030 gnd.n4573 gnd.n1938 585
R3031 gnd.n4714 gnd.n1939 585
R3032 gnd.n4714 gnd.n4713 585
R3033 gnd.n4715 gnd.n1929 585
R3034 gnd.n4716 gnd.n4715 585
R3035 gnd.n4477 gnd.n1937 585
R3036 gnd.n4480 gnd.n4479 585
R3037 gnd.n4478 gnd.n4441 585
R3038 gnd.n4494 gnd.n4493 585
R3039 gnd.n4496 gnd.n4495 585
R3040 gnd.n4499 gnd.n4498 585
R3041 gnd.n4497 gnd.n4434 585
R3042 gnd.n4513 gnd.n4512 585
R3043 gnd.n4515 gnd.n4514 585
R3044 gnd.n4518 gnd.n4517 585
R3045 gnd.n4516 gnd.n4427 585
R3046 gnd.n4532 gnd.n4531 585
R3047 gnd.n4534 gnd.n4533 585
R3048 gnd.n4537 gnd.n4536 585
R3049 gnd.n4535 gnd.n4419 585
R3050 gnd.n4550 gnd.n4549 585
R3051 gnd.n4552 gnd.n4551 585
R3052 gnd.n4553 gnd.n4416 585
R3053 gnd.n4415 gnd.n1858 585
R3054 gnd.n4836 gnd.n1858 585
R3055 gnd.n445 gnd.n371 585
R3056 gnd.n452 gnd.n451 585
R3057 gnd.n454 gnd.n453 585
R3058 gnd.n456 gnd.n455 585
R3059 gnd.n458 gnd.n457 585
R3060 gnd.n460 gnd.n459 585
R3061 gnd.n462 gnd.n461 585
R3062 gnd.n464 gnd.n463 585
R3063 gnd.n466 gnd.n465 585
R3064 gnd.n468 gnd.n467 585
R3065 gnd.n470 gnd.n469 585
R3066 gnd.n472 gnd.n471 585
R3067 gnd.n474 gnd.n473 585
R3068 gnd.n476 gnd.n475 585
R3069 gnd.n478 gnd.n477 585
R3070 gnd.n480 gnd.n479 585
R3071 gnd.n482 gnd.n481 585
R3072 gnd.n483 gnd.n355 585
R3073 gnd.n484 gnd.n257 585
R3074 gnd.n8003 gnd.n257 585
R3075 gnd.n447 gnd.n446 585
R3076 gnd.n446 gnd.n250 585
R3077 gnd.n444 gnd.n249 585
R3078 gnd.n8011 gnd.n249 585
R3079 gnd.n443 gnd.n442 585
R3080 gnd.n442 gnd.n241 585
R3081 gnd.n375 gnd.n240 585
R3082 gnd.n8017 gnd.n240 585
R3083 gnd.n438 gnd.n437 585
R3084 gnd.n437 gnd.n231 585
R3085 gnd.n436 gnd.n230 585
R3086 gnd.n8023 gnd.n230 585
R3087 gnd.n435 gnd.n434 585
R3088 gnd.n434 gnd.n228 585
R3089 gnd.n377 gnd.n221 585
R3090 gnd.n8029 gnd.n221 585
R3091 gnd.n430 gnd.n429 585
R3092 gnd.n429 gnd.n211 585
R3093 gnd.n428 gnd.n210 585
R3094 gnd.n8035 gnd.n210 585
R3095 gnd.n427 gnd.n426 585
R3096 gnd.n426 gnd.n202 585
R3097 gnd.n379 gnd.n201 585
R3098 gnd.n8041 gnd.n201 585
R3099 gnd.n422 gnd.n421 585
R3100 gnd.n421 gnd.n199 585
R3101 gnd.n420 gnd.n191 585
R3102 gnd.n8047 gnd.n191 585
R3103 gnd.n419 gnd.n418 585
R3104 gnd.n418 gnd.n189 585
R3105 gnd.n381 gnd.n182 585
R3106 gnd.n8053 gnd.n182 585
R3107 gnd.n414 gnd.n413 585
R3108 gnd.n413 gnd.n173 585
R3109 gnd.n412 gnd.n172 585
R3110 gnd.n8059 gnd.n172 585
R3111 gnd.n411 gnd.n410 585
R3112 gnd.n410 gnd.n164 585
R3113 gnd.n383 gnd.n163 585
R3114 gnd.n8065 gnd.n163 585
R3115 gnd.n406 gnd.n405 585
R3116 gnd.n405 gnd.n161 585
R3117 gnd.n404 gnd.n153 585
R3118 gnd.n8071 gnd.n153 585
R3119 gnd.n403 gnd.n402 585
R3120 gnd.n402 gnd.n151 585
R3121 gnd.n385 gnd.n144 585
R3122 gnd.n8077 gnd.n144 585
R3123 gnd.n398 gnd.n397 585
R3124 gnd.n397 gnd.n136 585
R3125 gnd.n396 gnd.n135 585
R3126 gnd.n8083 gnd.n135 585
R3127 gnd.n395 gnd.n394 585
R3128 gnd.n394 gnd.n125 585
R3129 gnd.n387 gnd.n124 585
R3130 gnd.n8089 gnd.n124 585
R3131 gnd.n390 gnd.n389 585
R3132 gnd.n389 gnd.n122 585
R3133 gnd.n104 gnd.n103 585
R3134 gnd.n107 gnd.n104 585
R3135 gnd.n8099 gnd.n8098 585
R3136 gnd.n8098 gnd.n8097 585
R3137 gnd.n8100 gnd.n102 585
R3138 gnd.n7822 gnd.n102 585
R3139 gnd.n7807 gnd.n100 585
R3140 gnd.n7808 gnd.n7807 585
R3141 gnd.n506 gnd.n499 585
R3142 gnd.n7813 gnd.n499 585
R3143 gnd.n7802 gnd.n7801 585
R3144 gnd.n7803 gnd.n7802 585
R3145 gnd.n505 gnd.n504 585
R3146 gnd.n7784 gnd.n504 585
R3147 gnd.n7797 gnd.n7796 585
R3148 gnd.n7796 gnd.n7795 585
R3149 gnd.n509 gnd.n508 585
R3150 gnd.n7790 gnd.n509 585
R3151 gnd.n7775 gnd.n7774 585
R3152 gnd.n7776 gnd.n7775 585
R3153 gnd.n528 gnd.n527 585
R3154 gnd.n7750 gnd.n527 585
R3155 gnd.n7770 gnd.n7769 585
R3156 gnd.n7769 gnd.n7768 585
R3157 gnd.n531 gnd.n530 585
R3158 gnd.n7744 gnd.n531 585
R3159 gnd.n4632 gnd.n544 585
R3160 gnd.n7757 gnd.n544 585
R3161 gnd.n4633 gnd.n4630 585
R3162 gnd.n4630 gnd.n2045 585
R3163 gnd.n4634 gnd.n2044 585
R3164 gnd.n4652 gnd.n2044 585
R3165 gnd.n2053 gnd.n2036 585
R3166 gnd.n4659 gnd.n2036 585
R3167 gnd.n4639 gnd.n4638 585
R3168 gnd.n4640 gnd.n4639 585
R3169 gnd.n2052 gnd.n2025 585
R3170 gnd.n4665 gnd.n2025 585
R3171 gnd.n4626 gnd.n4625 585
R3172 gnd.n4625 gnd.n4624 585
R3173 gnd.n2055 gnd.n2015 585
R3174 gnd.n4671 gnd.n2015 585
R3175 gnd.n4614 gnd.n4613 585
R3176 gnd.n4615 gnd.n4614 585
R3177 gnd.n2058 gnd.n2004 585
R3178 gnd.n4677 gnd.n2004 585
R3179 gnd.n4609 gnd.n4608 585
R3180 gnd.n4608 gnd.n4607 585
R3181 gnd.n2060 gnd.n1994 585
R3182 gnd.n4683 gnd.n1994 585
R3183 gnd.n4600 gnd.n4599 585
R3184 gnd.n4601 gnd.n4600 585
R3185 gnd.n2121 gnd.n1984 585
R3186 gnd.n4689 gnd.n1984 585
R3187 gnd.n4595 gnd.n4594 585
R3188 gnd.n4594 gnd.n4593 585
R3189 gnd.n2123 gnd.n1974 585
R3190 gnd.n4695 gnd.n1974 585
R3191 gnd.n4586 gnd.n4585 585
R3192 gnd.n4587 gnd.n4586 585
R3193 gnd.n2126 gnd.n1963 585
R3194 gnd.n4701 gnd.n1963 585
R3195 gnd.n4581 gnd.n4580 585
R3196 gnd.n4580 gnd.n4579 585
R3197 gnd.n2128 gnd.n1952 585
R3198 gnd.n4707 gnd.n1952 585
R3199 gnd.n4572 gnd.n4571 585
R3200 gnd.n4573 gnd.n4572 585
R3201 gnd.n2130 gnd.n1940 585
R3202 gnd.n4713 gnd.n1940 585
R3203 gnd.n4567 gnd.n1935 585
R3204 gnd.n4716 gnd.n1935 585
R3205 gnd.n6874 gnd.n6873 585
R3206 gnd.n6875 gnd.n6874 585
R3207 gnd.n5404 gnd.n5402 585
R3208 gnd.n5402 gnd.n1145 585
R3209 gnd.n6768 gnd.n5763 585
R3210 gnd.n5763 gnd.n1137 585
R3211 gnd.n6770 gnd.n6769 585
R3212 gnd.n6771 gnd.n6770 585
R3213 gnd.n5764 gnd.n5762 585
R3214 gnd.n5762 gnd.n5490 585
R3215 gnd.n6763 gnd.n6762 585
R3216 gnd.n6762 gnd.n5489 585
R3217 gnd.n6761 gnd.n5766 585
R3218 gnd.n6761 gnd.n6760 585
R3219 gnd.n6725 gnd.n5767 585
R3220 gnd.n6748 gnd.n5767 585
R3221 gnd.n6726 gnd.n5790 585
R3222 gnd.n5790 gnd.n5774 585
R3223 gnd.n6728 gnd.n6727 585
R3224 gnd.n6729 gnd.n6728 585
R3225 gnd.n5791 gnd.n5789 585
R3226 gnd.n6715 gnd.n5789 585
R3227 gnd.n6719 gnd.n6718 585
R3228 gnd.n6718 gnd.n6717 585
R3229 gnd.n5794 gnd.n5793 585
R3230 gnd.n6703 gnd.n5794 585
R3231 gnd.n6679 gnd.n6678 585
R3232 gnd.n6678 gnd.n5801 585
R3233 gnd.n6680 gnd.n5820 585
R3234 gnd.n5820 gnd.n5809 585
R3235 gnd.n6682 gnd.n6681 585
R3236 gnd.n6683 gnd.n6682 585
R3237 gnd.n5821 gnd.n5819 585
R3238 gnd.n5827 gnd.n5819 585
R3239 gnd.n6672 gnd.n6671 585
R3240 gnd.n6671 gnd.n6670 585
R3241 gnd.n5824 gnd.n5823 585
R3242 gnd.n6660 gnd.n5824 585
R3243 gnd.n6636 gnd.n5852 585
R3244 gnd.n5852 gnd.n5843 585
R3245 gnd.n6638 gnd.n6637 585
R3246 gnd.n6639 gnd.n6638 585
R3247 gnd.n5853 gnd.n5851 585
R3248 gnd.n5860 gnd.n5851 585
R3249 gnd.n6631 gnd.n6630 585
R3250 gnd.n6630 gnd.n6629 585
R3251 gnd.n5856 gnd.n5855 585
R3252 gnd.n6619 gnd.n5856 585
R3253 gnd.n6606 gnd.n5876 585
R3254 gnd.n5876 gnd.n5867 585
R3255 gnd.n6608 gnd.n6607 585
R3256 gnd.n6609 gnd.n6608 585
R3257 gnd.n5877 gnd.n5875 585
R3258 gnd.n5884 gnd.n5875 585
R3259 gnd.n6601 gnd.n6600 585
R3260 gnd.n6600 gnd.n6599 585
R3261 gnd.n5880 gnd.n5879 585
R3262 gnd.n6588 gnd.n5880 585
R3263 gnd.n6575 gnd.n5901 585
R3264 gnd.n5901 gnd.n5892 585
R3265 gnd.n6577 gnd.n6576 585
R3266 gnd.n6578 gnd.n6577 585
R3267 gnd.n5902 gnd.n5900 585
R3268 gnd.n5909 gnd.n5900 585
R3269 gnd.n6570 gnd.n6569 585
R3270 gnd.n6569 gnd.n6568 585
R3271 gnd.n5905 gnd.n5904 585
R3272 gnd.n6557 gnd.n5905 585
R3273 gnd.n6544 gnd.n5927 585
R3274 gnd.n5927 gnd.n5917 585
R3275 gnd.n6546 gnd.n6545 585
R3276 gnd.n6547 gnd.n6546 585
R3277 gnd.n5928 gnd.n5926 585
R3278 gnd.n5935 gnd.n5926 585
R3279 gnd.n6539 gnd.n6538 585
R3280 gnd.n6538 gnd.n6537 585
R3281 gnd.n5931 gnd.n5930 585
R3282 gnd.n6526 gnd.n5931 585
R3283 gnd.n6513 gnd.n5953 585
R3284 gnd.n5953 gnd.n5952 585
R3285 gnd.n6515 gnd.n6514 585
R3286 gnd.n6516 gnd.n6515 585
R3287 gnd.n5954 gnd.n5951 585
R3288 gnd.n5961 gnd.n5951 585
R3289 gnd.n6508 gnd.n6507 585
R3290 gnd.n6507 gnd.n6506 585
R3291 gnd.n5957 gnd.n5956 585
R3292 gnd.n6495 gnd.n5957 585
R3293 gnd.n6482 gnd.n5979 585
R3294 gnd.n5979 gnd.n5978 585
R3295 gnd.n6484 gnd.n6483 585
R3296 gnd.n6485 gnd.n6484 585
R3297 gnd.n5980 gnd.n5977 585
R3298 gnd.n5987 gnd.n5977 585
R3299 gnd.n6477 gnd.n6476 585
R3300 gnd.n6476 gnd.n6475 585
R3301 gnd.n5983 gnd.n5982 585
R3302 gnd.n6464 gnd.n5983 585
R3303 gnd.n6451 gnd.n6004 585
R3304 gnd.n6004 gnd.n5995 585
R3305 gnd.n6453 gnd.n6452 585
R3306 gnd.n6454 gnd.n6453 585
R3307 gnd.n6005 gnd.n6003 585
R3308 gnd.n6012 gnd.n6003 585
R3309 gnd.n6446 gnd.n6445 585
R3310 gnd.n6445 gnd.n6444 585
R3311 gnd.n6008 gnd.n6007 585
R3312 gnd.n6433 gnd.n6008 585
R3313 gnd.n6420 gnd.n6419 585
R3314 gnd.n6418 gnd.n6371 585
R3315 gnd.n6417 gnd.n6370 585
R3316 gnd.n6422 gnd.n6370 585
R3317 gnd.n6416 gnd.n6415 585
R3318 gnd.n6414 gnd.n6413 585
R3319 gnd.n6412 gnd.n6411 585
R3320 gnd.n6410 gnd.n6409 585
R3321 gnd.n6408 gnd.n6407 585
R3322 gnd.n6406 gnd.n6405 585
R3323 gnd.n6404 gnd.n6403 585
R3324 gnd.n6402 gnd.n6401 585
R3325 gnd.n6400 gnd.n6399 585
R3326 gnd.n6398 gnd.n6397 585
R3327 gnd.n6396 gnd.n6395 585
R3328 gnd.n6394 gnd.n6393 585
R3329 gnd.n6392 gnd.n6391 585
R3330 gnd.n6387 gnd.n6018 585
R3331 gnd.n6843 gnd.n6842 585
R3332 gnd.n6845 gnd.n5432 585
R3333 gnd.n6847 gnd.n6846 585
R3334 gnd.n6848 gnd.n5425 585
R3335 gnd.n6850 gnd.n6849 585
R3336 gnd.n6852 gnd.n5423 585
R3337 gnd.n6854 gnd.n6853 585
R3338 gnd.n6855 gnd.n5418 585
R3339 gnd.n6857 gnd.n6856 585
R3340 gnd.n6859 gnd.n5416 585
R3341 gnd.n6861 gnd.n6860 585
R3342 gnd.n6862 gnd.n5411 585
R3343 gnd.n6864 gnd.n6863 585
R3344 gnd.n6866 gnd.n5409 585
R3345 gnd.n6868 gnd.n6867 585
R3346 gnd.n6869 gnd.n5407 585
R3347 gnd.n6870 gnd.n5403 585
R3348 gnd.n5403 gnd.n5401 585
R3349 gnd.n5757 gnd.n1147 585
R3350 gnd.n6875 gnd.n1147 585
R3351 gnd.n5758 gnd.n5754 585
R3352 gnd.n5754 gnd.n1145 585
R3353 gnd.n5760 gnd.n5759 585
R3354 gnd.n5760 gnd.n1137 585
R3355 gnd.n6772 gnd.n5752 585
R3356 gnd.n6772 gnd.n6771 585
R3357 gnd.n6774 gnd.n6773 585
R3358 gnd.n6773 gnd.n5490 585
R3359 gnd.n5753 gnd.n5750 585
R3360 gnd.n5753 gnd.n5489 585
R3361 gnd.n6758 gnd.n6757 585
R3362 gnd.n6760 gnd.n6758 585
R3363 gnd.n5770 gnd.n5769 585
R3364 gnd.n6748 gnd.n5769 585
R3365 gnd.n6732 gnd.n6731 585
R3366 gnd.n6731 gnd.n5774 585
R3367 gnd.n6730 gnd.n5786 585
R3368 gnd.n6730 gnd.n6729 585
R3369 gnd.n6712 gnd.n5787 585
R3370 gnd.n6715 gnd.n5787 585
R3371 gnd.n6714 gnd.n6713 585
R3372 gnd.n6717 gnd.n6714 585
R3373 gnd.n5797 gnd.n5796 585
R3374 gnd.n6703 gnd.n5796 585
R3375 gnd.n6687 gnd.n6686 585
R3376 gnd.n6686 gnd.n5801 585
R3377 gnd.n6685 gnd.n5815 585
R3378 gnd.n6685 gnd.n5809 585
R3379 gnd.n6684 gnd.n5817 585
R3380 gnd.n6684 gnd.n6683 585
R3381 gnd.n6664 gnd.n5816 585
R3382 gnd.n5827 gnd.n5816 585
R3383 gnd.n6663 gnd.n5825 585
R3384 gnd.n6670 gnd.n5825 585
R3385 gnd.n6662 gnd.n6661 585
R3386 gnd.n6661 gnd.n6660 585
R3387 gnd.n5836 gnd.n5833 585
R3388 gnd.n5843 gnd.n5836 585
R3389 gnd.n6641 gnd.n6640 585
R3390 gnd.n6640 gnd.n6639 585
R3391 gnd.n5849 gnd.n5848 585
R3392 gnd.n5860 gnd.n5849 585
R3393 gnd.n6622 gnd.n5858 585
R3394 gnd.n6629 gnd.n5858 585
R3395 gnd.n6621 gnd.n6620 585
R3396 gnd.n6620 gnd.n6619 585
R3397 gnd.n5866 gnd.n5864 585
R3398 gnd.n5867 gnd.n5866 585
R3399 gnd.n6611 gnd.n6610 585
R3400 gnd.n6610 gnd.n6609 585
R3401 gnd.n5873 gnd.n5872 585
R3402 gnd.n5884 gnd.n5873 585
R3403 gnd.n6591 gnd.n5882 585
R3404 gnd.n6599 gnd.n5882 585
R3405 gnd.n6590 gnd.n6589 585
R3406 gnd.n6589 gnd.n6588 585
R3407 gnd.n5891 gnd.n5889 585
R3408 gnd.n5892 gnd.n5891 585
R3409 gnd.n6580 gnd.n6579 585
R3410 gnd.n6579 gnd.n6578 585
R3411 gnd.n5898 gnd.n5897 585
R3412 gnd.n5909 gnd.n5898 585
R3413 gnd.n6560 gnd.n5907 585
R3414 gnd.n6568 gnd.n5907 585
R3415 gnd.n6559 gnd.n6558 585
R3416 gnd.n6558 gnd.n6557 585
R3417 gnd.n5916 gnd.n5914 585
R3418 gnd.n5917 gnd.n5916 585
R3419 gnd.n6549 gnd.n6548 585
R3420 gnd.n6548 gnd.n6547 585
R3421 gnd.n5923 gnd.n5922 585
R3422 gnd.n5935 gnd.n5923 585
R3423 gnd.n6529 gnd.n5933 585
R3424 gnd.n6537 gnd.n5933 585
R3425 gnd.n6528 gnd.n6527 585
R3426 gnd.n6527 gnd.n6526 585
R3427 gnd.n5942 gnd.n5940 585
R3428 gnd.n5952 gnd.n5942 585
R3429 gnd.n6518 gnd.n6517 585
R3430 gnd.n6517 gnd.n6516 585
R3431 gnd.n5948 gnd.n5947 585
R3432 gnd.n5961 gnd.n5948 585
R3433 gnd.n6498 gnd.n5959 585
R3434 gnd.n6506 gnd.n5959 585
R3435 gnd.n6497 gnd.n6496 585
R3436 gnd.n6496 gnd.n6495 585
R3437 gnd.n5968 gnd.n5966 585
R3438 gnd.n5978 gnd.n5968 585
R3439 gnd.n6487 gnd.n6486 585
R3440 gnd.n6486 gnd.n6485 585
R3441 gnd.n5974 gnd.n5973 585
R3442 gnd.n5987 gnd.n5974 585
R3443 gnd.n6467 gnd.n5985 585
R3444 gnd.n6475 gnd.n5985 585
R3445 gnd.n6466 gnd.n6465 585
R3446 gnd.n6465 gnd.n6464 585
R3447 gnd.n5994 gnd.n5992 585
R3448 gnd.n5995 gnd.n5994 585
R3449 gnd.n6456 gnd.n6455 585
R3450 gnd.n6455 gnd.n6454 585
R3451 gnd.n6001 gnd.n6000 585
R3452 gnd.n6012 gnd.n6001 585
R3453 gnd.n6436 gnd.n6010 585
R3454 gnd.n6444 gnd.n6010 585
R3455 gnd.n6435 gnd.n6434 585
R3456 gnd.n6434 gnd.n6433 585
R3457 gnd.n3728 gnd.n3727 585
R3458 gnd.n3728 gnd.n2187 585
R3459 gnd.n3726 gnd.n3677 585
R3460 gnd.n3883 gnd.n3677 585
R3461 gnd.n3886 gnd.n3676 585
R3462 gnd.n3886 gnd.n3885 585
R3463 gnd.n3888 gnd.n3887 585
R3464 gnd.n3887 gnd.n2193 585
R3465 gnd.n3889 gnd.n3660 585
R3466 gnd.n3660 gnd.n3659 585
R3467 gnd.n3891 gnd.n3890 585
R3468 gnd.n3892 gnd.n3891 585
R3469 gnd.n3675 gnd.n3658 585
R3470 gnd.n3658 gnd.n2200 585
R3471 gnd.n3674 gnd.n3673 585
R3472 gnd.n3673 gnd.n2199 585
R3473 gnd.n3672 gnd.n3661 585
R3474 gnd.n3672 gnd.n3671 585
R3475 gnd.n3668 gnd.n3667 585
R3476 gnd.n3668 gnd.n2207 585
R3477 gnd.n3666 gnd.n3662 585
R3478 gnd.n3662 gnd.n2206 585
R3479 gnd.n3665 gnd.n3664 585
R3480 gnd.n3664 gnd.n2215 585
R3481 gnd.n3663 gnd.n3643 585
R3482 gnd.n3643 gnd.n2213 585
R3483 gnd.n3907 gnd.n3644 585
R3484 gnd.n3907 gnd.n3906 585
R3485 gnd.n3908 gnd.n3642 585
R3486 gnd.n3908 gnd.n2222 585
R3487 gnd.n3910 gnd.n3909 585
R3488 gnd.n3909 gnd.n2221 585
R3489 gnd.n3911 gnd.n3640 585
R3490 gnd.n3640 gnd.n3639 585
R3491 gnd.n3913 gnd.n3912 585
R3492 gnd.n3914 gnd.n3913 585
R3493 gnd.n3641 gnd.n3629 585
R3494 gnd.n3629 gnd.n2228 585
R3495 gnd.n3921 gnd.n3628 585
R3496 gnd.n3921 gnd.n3920 585
R3497 gnd.n3923 gnd.n3922 585
R3498 gnd.n3922 gnd.n2235 585
R3499 gnd.n3924 gnd.n3624 585
R3500 gnd.n3624 gnd.n2234 585
R3501 gnd.n3926 gnd.n3925 585
R3502 gnd.n3927 gnd.n3926 585
R3503 gnd.n3627 gnd.n3623 585
R3504 gnd.n3623 gnd.n2242 585
R3505 gnd.n3626 gnd.n3625 585
R3506 gnd.n3625 gnd.n2241 585
R3507 gnd.n3614 gnd.n3613 585
R3508 gnd.n3934 gnd.n3614 585
R3509 gnd.n3938 gnd.n3937 585
R3510 gnd.n3937 gnd.n3936 585
R3511 gnd.n3939 gnd.n3610 585
R3512 gnd.n3610 gnd.n2248 585
R3513 gnd.n3941 gnd.n3940 585
R3514 gnd.n3942 gnd.n3941 585
R3515 gnd.n3612 gnd.n3609 585
R3516 gnd.n3609 gnd.n2255 585
R3517 gnd.n3611 gnd.n3599 585
R3518 gnd.n3599 gnd.n2254 585
R3519 gnd.n3950 gnd.n3598 585
R3520 gnd.n3950 gnd.n3949 585
R3521 gnd.n3952 gnd.n3951 585
R3522 gnd.n3951 gnd.n2262 585
R3523 gnd.n3953 gnd.n3595 585
R3524 gnd.n3595 gnd.n2261 585
R3525 gnd.n3955 gnd.n3954 585
R3526 gnd.n3956 gnd.n3955 585
R3527 gnd.n3597 gnd.n3594 585
R3528 gnd.n3594 gnd.n2269 585
R3529 gnd.n3596 gnd.n3586 585
R3530 gnd.n3586 gnd.n2268 585
R3531 gnd.n3966 gnd.n3585 585
R3532 gnd.n3966 gnd.n3965 585
R3533 gnd.n3968 gnd.n3967 585
R3534 gnd.n3967 gnd.n2276 585
R3535 gnd.n3969 gnd.n3582 585
R3536 gnd.n3582 gnd.n2275 585
R3537 gnd.n3971 gnd.n3970 585
R3538 gnd.n3972 gnd.n3971 585
R3539 gnd.n3584 gnd.n3581 585
R3540 gnd.n3581 gnd.n2283 585
R3541 gnd.n3583 gnd.n3573 585
R3542 gnd.n3573 gnd.n2282 585
R3543 gnd.n3982 gnd.n3572 585
R3544 gnd.n3982 gnd.n3981 585
R3545 gnd.n3984 gnd.n3983 585
R3546 gnd.n3983 gnd.n2289 585
R3547 gnd.n3985 gnd.n3569 585
R3548 gnd.n3569 gnd.n3568 585
R3549 gnd.n3987 gnd.n3986 585
R3550 gnd.n3988 gnd.n3987 585
R3551 gnd.n3571 gnd.n3567 585
R3552 gnd.n3567 gnd.n2296 585
R3553 gnd.n3570 gnd.n3559 585
R3554 gnd.n3559 gnd.n2295 585
R3555 gnd.n3998 gnd.n3558 585
R3556 gnd.n3998 gnd.n3997 585
R3557 gnd.n4000 gnd.n3999 585
R3558 gnd.n3999 gnd.n2303 585
R3559 gnd.n4001 gnd.n3555 585
R3560 gnd.n3555 gnd.n2302 585
R3561 gnd.n4003 gnd.n4002 585
R3562 gnd.n4004 gnd.n4003 585
R3563 gnd.n3557 gnd.n3554 585
R3564 gnd.n3554 gnd.n2310 585
R3565 gnd.n3556 gnd.n3534 585
R3566 gnd.n3534 gnd.n2309 585
R3567 gnd.n4014 gnd.n3535 585
R3568 gnd.n4014 gnd.n4013 585
R3569 gnd.n4015 gnd.n3533 585
R3570 gnd.n4015 gnd.n2317 585
R3571 gnd.n4017 gnd.n4016 585
R3572 gnd.n4016 gnd.n2316 585
R3573 gnd.n4018 gnd.n3532 585
R3574 gnd.n3546 gnd.n3532 585
R3575 gnd.n4020 gnd.n4019 585
R3576 gnd.n4020 gnd.n2324 585
R3577 gnd.n4021 gnd.n3531 585
R3578 gnd.n4021 gnd.n2323 585
R3579 gnd.n4023 gnd.n4022 585
R3580 gnd.n4022 gnd.n2333 585
R3581 gnd.n4024 gnd.n3528 585
R3582 gnd.n3528 gnd.n2330 585
R3583 gnd.n4026 gnd.n4025 585
R3584 gnd.n4027 gnd.n4026 585
R3585 gnd.n3530 gnd.n3527 585
R3586 gnd.n3527 gnd.n2339 585
R3587 gnd.n3529 gnd.n3515 585
R3588 gnd.n4033 gnd.n3515 585
R3589 gnd.n4035 gnd.n3514 585
R3590 gnd.n4035 gnd.n4034 585
R3591 gnd.n4037 gnd.n4036 585
R3592 gnd.n4036 gnd.n2346 585
R3593 gnd.n4038 gnd.n3510 585
R3594 gnd.n3510 gnd.n2345 585
R3595 gnd.n4040 gnd.n4039 585
R3596 gnd.n4041 gnd.n4040 585
R3597 gnd.n3513 gnd.n3509 585
R3598 gnd.n3509 gnd.n2353 585
R3599 gnd.n3512 gnd.n3511 585
R3600 gnd.n3511 gnd.n2352 585
R3601 gnd.n3501 gnd.n3500 585
R3602 gnd.n4048 gnd.n3501 585
R3603 gnd.n4052 gnd.n4051 585
R3604 gnd.n4051 gnd.n4050 585
R3605 gnd.n4053 gnd.n3497 585
R3606 gnd.n3497 gnd.n2359 585
R3607 gnd.n4055 gnd.n4054 585
R3608 gnd.n4056 gnd.n4055 585
R3609 gnd.n3499 gnd.n3496 585
R3610 gnd.n3496 gnd.n2365 585
R3611 gnd.n3498 gnd.n3484 585
R3612 gnd.n4062 gnd.n3484 585
R3613 gnd.n4064 gnd.n3483 585
R3614 gnd.n4064 gnd.n4063 585
R3615 gnd.n4066 gnd.n4065 585
R3616 gnd.n4065 gnd.n2372 585
R3617 gnd.n4067 gnd.n3478 585
R3618 gnd.n3478 gnd.n2371 585
R3619 gnd.n4069 gnd.n4068 585
R3620 gnd.n4070 gnd.n4069 585
R3621 gnd.n3482 gnd.n3477 585
R3622 gnd.n3477 gnd.n2379 585
R3623 gnd.n3481 gnd.n3480 585
R3624 gnd.n3480 gnd.n2378 585
R3625 gnd.n3479 gnd.n2398 585
R3626 gnd.n4077 gnd.n2398 585
R3627 gnd.n4080 gnd.n2397 585
R3628 gnd.n4080 gnd.n4079 585
R3629 gnd.n4082 gnd.n4081 585
R3630 gnd.n4081 gnd.n2385 585
R3631 gnd.n4083 gnd.n2395 585
R3632 gnd.n2395 gnd.n2393 585
R3633 gnd.n4085 gnd.n4084 585
R3634 gnd.n4086 gnd.n4085 585
R3635 gnd.n2396 gnd.n2394 585
R3636 gnd.n3465 gnd.n2394 585
R3637 gnd.n3462 gnd.n3461 585
R3638 gnd.n3463 gnd.n3462 585
R3639 gnd.n3460 gnd.n2404 585
R3640 gnd.n2404 gnd.n1703 585
R3641 gnd.n3459 gnd.n3458 585
R3642 gnd.n3458 gnd.n1701 585
R3643 gnd.n3457 gnd.n2405 585
R3644 gnd.n3457 gnd.n3456 585
R3645 gnd.n1687 gnd.n1686 585
R3646 gnd.n1691 gnd.n1687 585
R3647 gnd.n4977 gnd.n4976 585
R3648 gnd.n4976 gnd.n4975 585
R3649 gnd.n4978 gnd.n1665 585
R3650 gnd.n2473 gnd.n1665 585
R3651 gnd.n5043 gnd.n5042 585
R3652 gnd.n5041 gnd.n1664 585
R3653 gnd.n5040 gnd.n1663 585
R3654 gnd.n5045 gnd.n1663 585
R3655 gnd.n5039 gnd.n5038 585
R3656 gnd.n5037 gnd.n5036 585
R3657 gnd.n5035 gnd.n5034 585
R3658 gnd.n5033 gnd.n5032 585
R3659 gnd.n5031 gnd.n5030 585
R3660 gnd.n5029 gnd.n5028 585
R3661 gnd.n5027 gnd.n5026 585
R3662 gnd.n5025 gnd.n5024 585
R3663 gnd.n5023 gnd.n5022 585
R3664 gnd.n5021 gnd.n5020 585
R3665 gnd.n5019 gnd.n5018 585
R3666 gnd.n5017 gnd.n5016 585
R3667 gnd.n5015 gnd.n5014 585
R3668 gnd.n5013 gnd.n5012 585
R3669 gnd.n5011 gnd.n5010 585
R3670 gnd.n5009 gnd.n5008 585
R3671 gnd.n5007 gnd.n5006 585
R3672 gnd.n5005 gnd.n5004 585
R3673 gnd.n5003 gnd.n5002 585
R3674 gnd.n5001 gnd.n5000 585
R3675 gnd.n4999 gnd.n4998 585
R3676 gnd.n4997 gnd.n4996 585
R3677 gnd.n4995 gnd.n4994 585
R3678 gnd.n4993 gnd.n4992 585
R3679 gnd.n4991 gnd.n4990 585
R3680 gnd.n4989 gnd.n4988 585
R3681 gnd.n4987 gnd.n4986 585
R3682 gnd.n4985 gnd.n4984 585
R3683 gnd.n4983 gnd.n1627 585
R3684 gnd.n5048 gnd.n5047 585
R3685 gnd.n1629 gnd.n1626 585
R3686 gnd.n2411 gnd.n2410 585
R3687 gnd.n2413 gnd.n2412 585
R3688 gnd.n2416 gnd.n2415 585
R3689 gnd.n2418 gnd.n2417 585
R3690 gnd.n2420 gnd.n2419 585
R3691 gnd.n2422 gnd.n2421 585
R3692 gnd.n2424 gnd.n2423 585
R3693 gnd.n2426 gnd.n2425 585
R3694 gnd.n2428 gnd.n2427 585
R3695 gnd.n2430 gnd.n2429 585
R3696 gnd.n2432 gnd.n2431 585
R3697 gnd.n2434 gnd.n2433 585
R3698 gnd.n2436 gnd.n2435 585
R3699 gnd.n2438 gnd.n2437 585
R3700 gnd.n2440 gnd.n2439 585
R3701 gnd.n2442 gnd.n2441 585
R3702 gnd.n2444 gnd.n2443 585
R3703 gnd.n2446 gnd.n2445 585
R3704 gnd.n2448 gnd.n2447 585
R3705 gnd.n2450 gnd.n2449 585
R3706 gnd.n2452 gnd.n2451 585
R3707 gnd.n2454 gnd.n2453 585
R3708 gnd.n2456 gnd.n2455 585
R3709 gnd.n2458 gnd.n2457 585
R3710 gnd.n2460 gnd.n2459 585
R3711 gnd.n2462 gnd.n2461 585
R3712 gnd.n2464 gnd.n2463 585
R3713 gnd.n2466 gnd.n2465 585
R3714 gnd.n2468 gnd.n2467 585
R3715 gnd.n2470 gnd.n2469 585
R3716 gnd.n2472 gnd.n2471 585
R3717 gnd.n3879 gnd.n3878 585
R3718 gnd.n3686 gnd.n3685 585
R3719 gnd.n3815 gnd.n3814 585
R3720 gnd.n3817 gnd.n3816 585
R3721 gnd.n3819 gnd.n3818 585
R3722 gnd.n3821 gnd.n3820 585
R3723 gnd.n3823 gnd.n3822 585
R3724 gnd.n3825 gnd.n3824 585
R3725 gnd.n3827 gnd.n3826 585
R3726 gnd.n3829 gnd.n3828 585
R3727 gnd.n3831 gnd.n3830 585
R3728 gnd.n3833 gnd.n3832 585
R3729 gnd.n3835 gnd.n3834 585
R3730 gnd.n3837 gnd.n3836 585
R3731 gnd.n3839 gnd.n3838 585
R3732 gnd.n3841 gnd.n3840 585
R3733 gnd.n3843 gnd.n3842 585
R3734 gnd.n3845 gnd.n3844 585
R3735 gnd.n3847 gnd.n3846 585
R3736 gnd.n3849 gnd.n3848 585
R3737 gnd.n3851 gnd.n3850 585
R3738 gnd.n3853 gnd.n3852 585
R3739 gnd.n3855 gnd.n3854 585
R3740 gnd.n3857 gnd.n3856 585
R3741 gnd.n3859 gnd.n3858 585
R3742 gnd.n3861 gnd.n3860 585
R3743 gnd.n3863 gnd.n3862 585
R3744 gnd.n3865 gnd.n3864 585
R3745 gnd.n3867 gnd.n3866 585
R3746 gnd.n3870 gnd.n3869 585
R3747 gnd.n3872 gnd.n3871 585
R3748 gnd.n3874 gnd.n3873 585
R3749 gnd.n3876 gnd.n3875 585
R3750 gnd.n3794 gnd.n1891 585
R3751 gnd.n3793 gnd.n3792 585
R3752 gnd.n3791 gnd.n3790 585
R3753 gnd.n3789 gnd.n3788 585
R3754 gnd.n3786 gnd.n3785 585
R3755 gnd.n3784 gnd.n3783 585
R3756 gnd.n3782 gnd.n3781 585
R3757 gnd.n3780 gnd.n3779 585
R3758 gnd.n3778 gnd.n3777 585
R3759 gnd.n3776 gnd.n3775 585
R3760 gnd.n3774 gnd.n3773 585
R3761 gnd.n3772 gnd.n3771 585
R3762 gnd.n3770 gnd.n3769 585
R3763 gnd.n3768 gnd.n3767 585
R3764 gnd.n3766 gnd.n3765 585
R3765 gnd.n3764 gnd.n3763 585
R3766 gnd.n3762 gnd.n3761 585
R3767 gnd.n3760 gnd.n3759 585
R3768 gnd.n3758 gnd.n3757 585
R3769 gnd.n3756 gnd.n3755 585
R3770 gnd.n3754 gnd.n3753 585
R3771 gnd.n3752 gnd.n3751 585
R3772 gnd.n3750 gnd.n3749 585
R3773 gnd.n3748 gnd.n3747 585
R3774 gnd.n3746 gnd.n3745 585
R3775 gnd.n3744 gnd.n3743 585
R3776 gnd.n3742 gnd.n3741 585
R3777 gnd.n3740 gnd.n3739 585
R3778 gnd.n3738 gnd.n3737 585
R3779 gnd.n3736 gnd.n3735 585
R3780 gnd.n3734 gnd.n3733 585
R3781 gnd.n3732 gnd.n3731 585
R3782 gnd.n3730 gnd.n3729 585
R3783 gnd.n3880 gnd.n3680 585
R3784 gnd.n3680 gnd.n2187 585
R3785 gnd.n3882 gnd.n3881 585
R3786 gnd.n3883 gnd.n3882 585
R3787 gnd.n3684 gnd.n3678 585
R3788 gnd.n3885 gnd.n3678 585
R3789 gnd.n3683 gnd.n3682 585
R3790 gnd.n3682 gnd.n2193 585
R3791 gnd.n3681 gnd.n3655 585
R3792 gnd.n3659 gnd.n3655 585
R3793 gnd.n3893 gnd.n3656 585
R3794 gnd.n3893 gnd.n3892 585
R3795 gnd.n3894 gnd.n3654 585
R3796 gnd.n3894 gnd.n2200 585
R3797 gnd.n3896 gnd.n3895 585
R3798 gnd.n3895 gnd.n2199 585
R3799 gnd.n3897 gnd.n3653 585
R3800 gnd.n3671 gnd.n3653 585
R3801 gnd.n3899 gnd.n3898 585
R3802 gnd.n3899 gnd.n2207 585
R3803 gnd.n3900 gnd.n3652 585
R3804 gnd.n3900 gnd.n2206 585
R3805 gnd.n3902 gnd.n3901 585
R3806 gnd.n3901 gnd.n2215 585
R3807 gnd.n3903 gnd.n3648 585
R3808 gnd.n3648 gnd.n2213 585
R3809 gnd.n3905 gnd.n3904 585
R3810 gnd.n3906 gnd.n3905 585
R3811 gnd.n3651 gnd.n3647 585
R3812 gnd.n3647 gnd.n2222 585
R3813 gnd.n3650 gnd.n3649 585
R3814 gnd.n3649 gnd.n2221 585
R3815 gnd.n3637 gnd.n3636 585
R3816 gnd.n3639 gnd.n3637 585
R3817 gnd.n3916 gnd.n3915 585
R3818 gnd.n3915 gnd.n3914 585
R3819 gnd.n3917 gnd.n3633 585
R3820 gnd.n3633 gnd.n2228 585
R3821 gnd.n3919 gnd.n3918 585
R3822 gnd.n3920 gnd.n3919 585
R3823 gnd.n3635 gnd.n3632 585
R3824 gnd.n3632 gnd.n2235 585
R3825 gnd.n3634 gnd.n3621 585
R3826 gnd.n3621 gnd.n2234 585
R3827 gnd.n3928 gnd.n3620 585
R3828 gnd.n3928 gnd.n3927 585
R3829 gnd.n3930 gnd.n3929 585
R3830 gnd.n3929 gnd.n2242 585
R3831 gnd.n3931 gnd.n3617 585
R3832 gnd.n3617 gnd.n2241 585
R3833 gnd.n3933 gnd.n3932 585
R3834 gnd.n3934 gnd.n3933 585
R3835 gnd.n3619 gnd.n3615 585
R3836 gnd.n3936 gnd.n3615 585
R3837 gnd.n3618 gnd.n3607 585
R3838 gnd.n3607 gnd.n2248 585
R3839 gnd.n3943 gnd.n3606 585
R3840 gnd.n3943 gnd.n3942 585
R3841 gnd.n3945 gnd.n3944 585
R3842 gnd.n3944 gnd.n2255 585
R3843 gnd.n3946 gnd.n3603 585
R3844 gnd.n3603 gnd.n2254 585
R3845 gnd.n3948 gnd.n3947 585
R3846 gnd.n3949 gnd.n3948 585
R3847 gnd.n3605 gnd.n3602 585
R3848 gnd.n3602 gnd.n2262 585
R3849 gnd.n3604 gnd.n3592 585
R3850 gnd.n3592 gnd.n2261 585
R3851 gnd.n3957 gnd.n3591 585
R3852 gnd.n3957 gnd.n3956 585
R3853 gnd.n3959 gnd.n3958 585
R3854 gnd.n3958 gnd.n2269 585
R3855 gnd.n3960 gnd.n3588 585
R3856 gnd.n3588 gnd.n2268 585
R3857 gnd.n3962 gnd.n3961 585
R3858 gnd.n3965 gnd.n3962 585
R3859 gnd.n3590 gnd.n3587 585
R3860 gnd.n3587 gnd.n2276 585
R3861 gnd.n3589 gnd.n3579 585
R3862 gnd.n3579 gnd.n2275 585
R3863 gnd.n3973 gnd.n3578 585
R3864 gnd.n3973 gnd.n3972 585
R3865 gnd.n3975 gnd.n3974 585
R3866 gnd.n3974 gnd.n2283 585
R3867 gnd.n3976 gnd.n3575 585
R3868 gnd.n3575 gnd.n2282 585
R3869 gnd.n3978 gnd.n3977 585
R3870 gnd.n3981 gnd.n3978 585
R3871 gnd.n3577 gnd.n3574 585
R3872 gnd.n3574 gnd.n2289 585
R3873 gnd.n3576 gnd.n3565 585
R3874 gnd.n3568 gnd.n3565 585
R3875 gnd.n3989 gnd.n3564 585
R3876 gnd.n3989 gnd.n3988 585
R3877 gnd.n3991 gnd.n3990 585
R3878 gnd.n3990 gnd.n2296 585
R3879 gnd.n3992 gnd.n3561 585
R3880 gnd.n3561 gnd.n2295 585
R3881 gnd.n3994 gnd.n3993 585
R3882 gnd.n3997 gnd.n3994 585
R3883 gnd.n3563 gnd.n3560 585
R3884 gnd.n3560 gnd.n2303 585
R3885 gnd.n3562 gnd.n3552 585
R3886 gnd.n3552 gnd.n2302 585
R3887 gnd.n4005 gnd.n3551 585
R3888 gnd.n4005 gnd.n4004 585
R3889 gnd.n4007 gnd.n4006 585
R3890 gnd.n4006 gnd.n2310 585
R3891 gnd.n4008 gnd.n3537 585
R3892 gnd.n3537 gnd.n2309 585
R3893 gnd.n4010 gnd.n4009 585
R3894 gnd.n4013 gnd.n4010 585
R3895 gnd.n3550 gnd.n3536 585
R3896 gnd.n3536 gnd.n2317 585
R3897 gnd.n3549 gnd.n3548 585
R3898 gnd.n3548 gnd.n2316 585
R3899 gnd.n3547 gnd.n3538 585
R3900 gnd.n3547 gnd.n3546 585
R3901 gnd.n3544 gnd.n3543 585
R3902 gnd.n3544 gnd.n2324 585
R3903 gnd.n3542 gnd.n3539 585
R3904 gnd.n3539 gnd.n2323 585
R3905 gnd.n3541 gnd.n3540 585
R3906 gnd.n3540 gnd.n2333 585
R3907 gnd.n3525 gnd.n3524 585
R3908 gnd.n3525 gnd.n2330 585
R3909 gnd.n4029 gnd.n4028 585
R3910 gnd.n4028 gnd.n4027 585
R3911 gnd.n4030 gnd.n3519 585
R3912 gnd.n3519 gnd.n2339 585
R3913 gnd.n4032 gnd.n4031 585
R3914 gnd.n4033 gnd.n4032 585
R3915 gnd.n3523 gnd.n3518 585
R3916 gnd.n4034 gnd.n3518 585
R3917 gnd.n3522 gnd.n3521 585
R3918 gnd.n3521 gnd.n2346 585
R3919 gnd.n3520 gnd.n3507 585
R3920 gnd.n3507 gnd.n2345 585
R3921 gnd.n4042 gnd.n3506 585
R3922 gnd.n4042 gnd.n4041 585
R3923 gnd.n4044 gnd.n4043 585
R3924 gnd.n4043 gnd.n2353 585
R3925 gnd.n4045 gnd.n3504 585
R3926 gnd.n3504 gnd.n2352 585
R3927 gnd.n4047 gnd.n4046 585
R3928 gnd.n4048 gnd.n4047 585
R3929 gnd.n3505 gnd.n3502 585
R3930 gnd.n4050 gnd.n3502 585
R3931 gnd.n3494 gnd.n3493 585
R3932 gnd.n3494 gnd.n2359 585
R3933 gnd.n4058 gnd.n4057 585
R3934 gnd.n4057 gnd.n4056 585
R3935 gnd.n4059 gnd.n3488 585
R3936 gnd.n3488 gnd.n2365 585
R3937 gnd.n4061 gnd.n4060 585
R3938 gnd.n4062 gnd.n4061 585
R3939 gnd.n3492 gnd.n3487 585
R3940 gnd.n4063 gnd.n3487 585
R3941 gnd.n3491 gnd.n3490 585
R3942 gnd.n3490 gnd.n2372 585
R3943 gnd.n3489 gnd.n3475 585
R3944 gnd.n3475 gnd.n2371 585
R3945 gnd.n4071 gnd.n3474 585
R3946 gnd.n4071 gnd.n4070 585
R3947 gnd.n4073 gnd.n4072 585
R3948 gnd.n4072 gnd.n2379 585
R3949 gnd.n4074 gnd.n2401 585
R3950 gnd.n2401 gnd.n2378 585
R3951 gnd.n4076 gnd.n4075 585
R3952 gnd.n4077 gnd.n4076 585
R3953 gnd.n3473 gnd.n2399 585
R3954 gnd.n4079 gnd.n2399 585
R3955 gnd.n3472 gnd.n3471 585
R3956 gnd.n3471 gnd.n2385 585
R3957 gnd.n3470 gnd.n3469 585
R3958 gnd.n3470 gnd.n2393 585
R3959 gnd.n3468 gnd.n2391 585
R3960 gnd.n4086 gnd.n2391 585
R3961 gnd.n3467 gnd.n3466 585
R3962 gnd.n3466 gnd.n3465 585
R3963 gnd.n2403 gnd.n2402 585
R3964 gnd.n3463 gnd.n2403 585
R3965 gnd.n2479 gnd.n2478 585
R3966 gnd.n2478 gnd.n1703 585
R3967 gnd.n2480 gnd.n2407 585
R3968 gnd.n2407 gnd.n1701 585
R3969 gnd.n2482 gnd.n2481 585
R3970 gnd.n3456 gnd.n2482 585
R3971 gnd.n2477 gnd.n2406 585
R3972 gnd.n2406 gnd.n1691 585
R3973 gnd.n2476 gnd.n1689 585
R3974 gnd.n4975 gnd.n1689 585
R3975 gnd.n2475 gnd.n2474 585
R3976 gnd.n2474 gnd.n2473 585
R3977 gnd.n5104 gnd.n1550 585
R3978 gnd.n3361 gnd.n1550 585
R3979 gnd.n5106 gnd.n5105 585
R3980 gnd.n5107 gnd.n5106 585
R3981 gnd.n1535 gnd.n1534 585
R3982 gnd.n3218 gnd.n1535 585
R3983 gnd.n5115 gnd.n5114 585
R3984 gnd.n5114 gnd.n5113 585
R3985 gnd.n5116 gnd.n1529 585
R3986 gnd.n3208 gnd.n1529 585
R3987 gnd.n5118 gnd.n5117 585
R3988 gnd.n5119 gnd.n5118 585
R3989 gnd.n1514 gnd.n1513 585
R3990 gnd.n3201 gnd.n1514 585
R3991 gnd.n5127 gnd.n5126 585
R3992 gnd.n5126 gnd.n5125 585
R3993 gnd.n5128 gnd.n1508 585
R3994 gnd.n3193 gnd.n1508 585
R3995 gnd.n5130 gnd.n5129 585
R3996 gnd.n5131 gnd.n5130 585
R3997 gnd.n1494 gnd.n1493 585
R3998 gnd.n3186 gnd.n1494 585
R3999 gnd.n5139 gnd.n5138 585
R4000 gnd.n5138 gnd.n5137 585
R4001 gnd.n5140 gnd.n1488 585
R4002 gnd.n3125 gnd.n1488 585
R4003 gnd.n5142 gnd.n5141 585
R4004 gnd.n5143 gnd.n5142 585
R4005 gnd.n1473 gnd.n1472 585
R4006 gnd.n3118 gnd.n1473 585
R4007 gnd.n5151 gnd.n5150 585
R4008 gnd.n5150 gnd.n5149 585
R4009 gnd.n5152 gnd.n1467 585
R4010 gnd.n3114 gnd.n1467 585
R4011 gnd.n5154 gnd.n5153 585
R4012 gnd.n5155 gnd.n5154 585
R4013 gnd.n1453 gnd.n1452 585
R4014 gnd.n3142 gnd.n1453 585
R4015 gnd.n5163 gnd.n5162 585
R4016 gnd.n5162 gnd.n5161 585
R4017 gnd.n5164 gnd.n1447 585
R4018 gnd.n3107 gnd.n1447 585
R4019 gnd.n5166 gnd.n5165 585
R4020 gnd.n5167 gnd.n5166 585
R4021 gnd.n1432 gnd.n1431 585
R4022 gnd.n3099 gnd.n1432 585
R4023 gnd.n5175 gnd.n5174 585
R4024 gnd.n5174 gnd.n5173 585
R4025 gnd.n5176 gnd.n1427 585
R4026 gnd.n3093 gnd.n1427 585
R4027 gnd.n5178 gnd.n5177 585
R4028 gnd.n5179 gnd.n5178 585
R4029 gnd.n1411 gnd.n1409 585
R4030 gnd.n3085 gnd.n1411 585
R4031 gnd.n5187 gnd.n5186 585
R4032 gnd.n5186 gnd.n5185 585
R4033 gnd.n1410 gnd.n1408 585
R4034 gnd.n3054 gnd.n1410 585
R4035 gnd.n3043 gnd.n3042 585
R4036 gnd.n3042 gnd.n2784 585
R4037 gnd.n3045 gnd.n3044 585
R4038 gnd.n3046 gnd.n3045 585
R4039 gnd.n3041 gnd.n2796 585
R4040 gnd.n3041 gnd.n3040 585
R4041 gnd.n2795 gnd.n2794 585
R4042 gnd.n3024 gnd.n2794 585
R4043 gnd.n2880 gnd.n2879 585
R4044 gnd.n2881 gnd.n2880 585
R4045 gnd.n1402 gnd.n1400 585
R4046 gnd.n1400 gnd.n1399 585
R4047 gnd.n5191 gnd.n5190 585
R4048 gnd.n5192 gnd.n5191 585
R4049 gnd.n1401 gnd.n1385 585
R4050 gnd.n1389 gnd.n1385 585
R4051 gnd.n5200 gnd.n5199 585
R4052 gnd.n5199 gnd.n5198 585
R4053 gnd.n5201 gnd.n1380 585
R4054 gnd.n1386 gnd.n1380 585
R4055 gnd.n5203 gnd.n5202 585
R4056 gnd.n5204 gnd.n5203 585
R4057 gnd.n1368 gnd.n1367 585
R4058 gnd.n1371 gnd.n1368 585
R4059 gnd.n5212 gnd.n5211 585
R4060 gnd.n5211 gnd.n5210 585
R4061 gnd.n5213 gnd.n1362 585
R4062 gnd.n1362 gnd.n1361 585
R4063 gnd.n5215 gnd.n5214 585
R4064 gnd.n5216 gnd.n5215 585
R4065 gnd.n1348 gnd.n1347 585
R4066 gnd.n1352 gnd.n1348 585
R4067 gnd.n5224 gnd.n5223 585
R4068 gnd.n5223 gnd.n5222 585
R4069 gnd.n5225 gnd.n1342 585
R4070 gnd.n1349 gnd.n1342 585
R4071 gnd.n5227 gnd.n5226 585
R4072 gnd.n5228 gnd.n5227 585
R4073 gnd.n1330 gnd.n1329 585
R4074 gnd.n1333 gnd.n1330 585
R4075 gnd.n5236 gnd.n5235 585
R4076 gnd.n5235 gnd.n5234 585
R4077 gnd.n5237 gnd.n1324 585
R4078 gnd.n1324 gnd.n1323 585
R4079 gnd.n5239 gnd.n5238 585
R4080 gnd.n5240 gnd.n5239 585
R4081 gnd.n1310 gnd.n1309 585
R4082 gnd.n1314 gnd.n1310 585
R4083 gnd.n5248 gnd.n5247 585
R4084 gnd.n5247 gnd.n5246 585
R4085 gnd.n5249 gnd.n1304 585
R4086 gnd.n1311 gnd.n1304 585
R4087 gnd.n5251 gnd.n5250 585
R4088 gnd.n5252 gnd.n5251 585
R4089 gnd.n1292 gnd.n1291 585
R4090 gnd.n1295 gnd.n1292 585
R4091 gnd.n5260 gnd.n5259 585
R4092 gnd.n5259 gnd.n5258 585
R4093 gnd.n5261 gnd.n1286 585
R4094 gnd.n1286 gnd.n1285 585
R4095 gnd.n5263 gnd.n5262 585
R4096 gnd.n5264 gnd.n5263 585
R4097 gnd.n1269 gnd.n1268 585
R4098 gnd.n1273 gnd.n1269 585
R4099 gnd.n5272 gnd.n5271 585
R4100 gnd.n5271 gnd.n5270 585
R4101 gnd.n5273 gnd.n1262 585
R4102 gnd.n1270 gnd.n1262 585
R4103 gnd.n5275 gnd.n5274 585
R4104 gnd.n5276 gnd.n5275 585
R4105 gnd.n1263 gnd.n1189 585
R4106 gnd.n1189 gnd.n1186 585
R4107 gnd.n5398 gnd.n5397 585
R4108 gnd.n5396 gnd.n1188 585
R4109 gnd.n5395 gnd.n1187 585
R4110 gnd.n5400 gnd.n1187 585
R4111 gnd.n5394 gnd.n5393 585
R4112 gnd.n5392 gnd.n5391 585
R4113 gnd.n5390 gnd.n5389 585
R4114 gnd.n5388 gnd.n5387 585
R4115 gnd.n5386 gnd.n5385 585
R4116 gnd.n5384 gnd.n5383 585
R4117 gnd.n5382 gnd.n5381 585
R4118 gnd.n5380 gnd.n5379 585
R4119 gnd.n5378 gnd.n5377 585
R4120 gnd.n5376 gnd.n5375 585
R4121 gnd.n5374 gnd.n5373 585
R4122 gnd.n5372 gnd.n5371 585
R4123 gnd.n5370 gnd.n5369 585
R4124 gnd.n5368 gnd.n5367 585
R4125 gnd.n5366 gnd.n5365 585
R4126 gnd.n5363 gnd.n5362 585
R4127 gnd.n5361 gnd.n5360 585
R4128 gnd.n5359 gnd.n5358 585
R4129 gnd.n5357 gnd.n5356 585
R4130 gnd.n5355 gnd.n5354 585
R4131 gnd.n5353 gnd.n5352 585
R4132 gnd.n5351 gnd.n5350 585
R4133 gnd.n5349 gnd.n5348 585
R4134 gnd.n5347 gnd.n5346 585
R4135 gnd.n5345 gnd.n5344 585
R4136 gnd.n5343 gnd.n5342 585
R4137 gnd.n5341 gnd.n5340 585
R4138 gnd.n5339 gnd.n5338 585
R4139 gnd.n5337 gnd.n5336 585
R4140 gnd.n5335 gnd.n5334 585
R4141 gnd.n5333 gnd.n5332 585
R4142 gnd.n5331 gnd.n5330 585
R4143 gnd.n5329 gnd.n5328 585
R4144 gnd.n5327 gnd.n5326 585
R4145 gnd.n5325 gnd.n5324 585
R4146 gnd.n5323 gnd.n5322 585
R4147 gnd.n5321 gnd.n5320 585
R4148 gnd.n5319 gnd.n5318 585
R4149 gnd.n5317 gnd.n5316 585
R4150 gnd.n5315 gnd.n5314 585
R4151 gnd.n5313 gnd.n5312 585
R4152 gnd.n5311 gnd.n5310 585
R4153 gnd.n5309 gnd.n5308 585
R4154 gnd.n5307 gnd.n5306 585
R4155 gnd.n5305 gnd.n5304 585
R4156 gnd.n5303 gnd.n5302 585
R4157 gnd.n5301 gnd.n5300 585
R4158 gnd.n5299 gnd.n5298 585
R4159 gnd.n5297 gnd.n5296 585
R4160 gnd.n5295 gnd.n5294 585
R4161 gnd.n5293 gnd.n5292 585
R4162 gnd.n5291 gnd.n5290 585
R4163 gnd.n5289 gnd.n5288 585
R4164 gnd.n5287 gnd.n5286 585
R4165 gnd.n5285 gnd.n5284 585
R4166 gnd.n1258 gnd.n1251 585
R4167 gnd.n2734 gnd.n2733 585
R4168 gnd.n2732 gnd.n2643 585
R4169 gnd.n2731 gnd.n2730 585
R4170 gnd.n2724 gnd.n2644 585
R4171 gnd.n2726 gnd.n2725 585
R4172 gnd.n2723 gnd.n2722 585
R4173 gnd.n2721 gnd.n2720 585
R4174 gnd.n2714 gnd.n2646 585
R4175 gnd.n2716 gnd.n2715 585
R4176 gnd.n2713 gnd.n2712 585
R4177 gnd.n2711 gnd.n2710 585
R4178 gnd.n2704 gnd.n2648 585
R4179 gnd.n2706 gnd.n2705 585
R4180 gnd.n2703 gnd.n2702 585
R4181 gnd.n2701 gnd.n2700 585
R4182 gnd.n2694 gnd.n2650 585
R4183 gnd.n2696 gnd.n2695 585
R4184 gnd.n2693 gnd.n2692 585
R4185 gnd.n2691 gnd.n2690 585
R4186 gnd.n2684 gnd.n2652 585
R4187 gnd.n2686 gnd.n2685 585
R4188 gnd.n2683 gnd.n2656 585
R4189 gnd.n2682 gnd.n2681 585
R4190 gnd.n2675 gnd.n2657 585
R4191 gnd.n2677 gnd.n2676 585
R4192 gnd.n2674 gnd.n2673 585
R4193 gnd.n2672 gnd.n2671 585
R4194 gnd.n2665 gnd.n2659 585
R4195 gnd.n2667 gnd.n2666 585
R4196 gnd.n2664 gnd.n2663 585
R4197 gnd.n2662 gnd.n1623 585
R4198 gnd.n5051 gnd.n5050 585
R4199 gnd.n5053 gnd.n5052 585
R4200 gnd.n5055 gnd.n5054 585
R4201 gnd.n5057 gnd.n5056 585
R4202 gnd.n5059 gnd.n5058 585
R4203 gnd.n5061 gnd.n5060 585
R4204 gnd.n5063 gnd.n5062 585
R4205 gnd.n5065 gnd.n5064 585
R4206 gnd.n5068 gnd.n5067 585
R4207 gnd.n5070 gnd.n5069 585
R4208 gnd.n5072 gnd.n5071 585
R4209 gnd.n5074 gnd.n5073 585
R4210 gnd.n5076 gnd.n5075 585
R4211 gnd.n5078 gnd.n5077 585
R4212 gnd.n5080 gnd.n5079 585
R4213 gnd.n5082 gnd.n5081 585
R4214 gnd.n5084 gnd.n5083 585
R4215 gnd.n5086 gnd.n5085 585
R4216 gnd.n5088 gnd.n5087 585
R4217 gnd.n5090 gnd.n5089 585
R4218 gnd.n5092 gnd.n5091 585
R4219 gnd.n5094 gnd.n5093 585
R4220 gnd.n5095 gnd.n1596 585
R4221 gnd.n5097 gnd.n5096 585
R4222 gnd.n1555 gnd.n1554 585
R4223 gnd.n5101 gnd.n5100 585
R4224 gnd.n5100 gnd.n5099 585
R4225 gnd.n3222 gnd.n2554 585
R4226 gnd.n3361 gnd.n2554 585
R4227 gnd.n3221 gnd.n1547 585
R4228 gnd.n5107 gnd.n1547 585
R4229 gnd.n3220 gnd.n3219 585
R4230 gnd.n3219 gnd.n3218 585
R4231 gnd.n2736 gnd.n1537 585
R4232 gnd.n5113 gnd.n1537 585
R4233 gnd.n3207 gnd.n3206 585
R4234 gnd.n3208 gnd.n3207 585
R4235 gnd.n3204 gnd.n1526 585
R4236 gnd.n5119 gnd.n1526 585
R4237 gnd.n3203 gnd.n3202 585
R4238 gnd.n3202 gnd.n3201 585
R4239 gnd.n2741 gnd.n1516 585
R4240 gnd.n5125 gnd.n1516 585
R4241 gnd.n3192 gnd.n3191 585
R4242 gnd.n3193 gnd.n3192 585
R4243 gnd.n3189 gnd.n1505 585
R4244 gnd.n5131 gnd.n1505 585
R4245 gnd.n3188 gnd.n3187 585
R4246 gnd.n3187 gnd.n3186 585
R4247 gnd.n2745 gnd.n1496 585
R4248 gnd.n5137 gnd.n1496 585
R4249 gnd.n3124 gnd.n3123 585
R4250 gnd.n3125 gnd.n3124 585
R4251 gnd.n3121 gnd.n1485 585
R4252 gnd.n5143 gnd.n1485 585
R4253 gnd.n3120 gnd.n3119 585
R4254 gnd.n3119 gnd.n3118 585
R4255 gnd.n3117 gnd.n1475 585
R4256 gnd.n5149 gnd.n1475 585
R4257 gnd.n3116 gnd.n3115 585
R4258 gnd.n3115 gnd.n3114 585
R4259 gnd.n3112 gnd.n1464 585
R4260 gnd.n5155 gnd.n1464 585
R4261 gnd.n3111 gnd.n2758 585
R4262 gnd.n3142 gnd.n2758 585
R4263 gnd.n3110 gnd.n1455 585
R4264 gnd.n5161 gnd.n1455 585
R4265 gnd.n3109 gnd.n3108 585
R4266 gnd.n3108 gnd.n3107 585
R4267 gnd.n2767 gnd.n1444 585
R4268 gnd.n5167 gnd.n1444 585
R4269 gnd.n3098 gnd.n3097 585
R4270 gnd.n3099 gnd.n3098 585
R4271 gnd.n3096 gnd.n1434 585
R4272 gnd.n5173 gnd.n1434 585
R4273 gnd.n3095 gnd.n3094 585
R4274 gnd.n3094 gnd.n3093 585
R4275 gnd.n2772 gnd.n1424 585
R4276 gnd.n5179 gnd.n1424 585
R4277 gnd.n3029 gnd.n2777 585
R4278 gnd.n3085 gnd.n2777 585
R4279 gnd.n3030 gnd.n1413 585
R4280 gnd.n5185 gnd.n1413 585
R4281 gnd.n3031 gnd.n2785 585
R4282 gnd.n3054 gnd.n2785 585
R4283 gnd.n3033 gnd.n3032 585
R4284 gnd.n3032 gnd.n2784 585
R4285 gnd.n3028 gnd.n2791 585
R4286 gnd.n3046 gnd.n2791 585
R4287 gnd.n3027 gnd.n2798 585
R4288 gnd.n3040 gnd.n2798 585
R4289 gnd.n3026 gnd.n3025 585
R4290 gnd.n3025 gnd.n3024 585
R4291 gnd.n2807 gnd.n2805 585
R4292 gnd.n2881 gnd.n2807 585
R4293 gnd.n2874 gnd.n2873 585
R4294 gnd.n2873 gnd.n1399 585
R4295 gnd.n2872 gnd.n1397 585
R4296 gnd.n5192 gnd.n1397 585
R4297 gnd.n2871 gnd.n2870 585
R4298 gnd.n2870 gnd.n1389 585
R4299 gnd.n2869 gnd.n1387 585
R4300 gnd.n5198 gnd.n1387 585
R4301 gnd.n2868 gnd.n2867 585
R4302 gnd.n2867 gnd.n1386 585
R4303 gnd.n2865 gnd.n1378 585
R4304 gnd.n5204 gnd.n1378 585
R4305 gnd.n2864 gnd.n2863 585
R4306 gnd.n2863 gnd.n1371 585
R4307 gnd.n2862 gnd.n1369 585
R4308 gnd.n5210 gnd.n1369 585
R4309 gnd.n2861 gnd.n2860 585
R4310 gnd.n2860 gnd.n1361 585
R4311 gnd.n2858 gnd.n1359 585
R4312 gnd.n5216 gnd.n1359 585
R4313 gnd.n2857 gnd.n2856 585
R4314 gnd.n2856 gnd.n1352 585
R4315 gnd.n2855 gnd.n1350 585
R4316 gnd.n5222 gnd.n1350 585
R4317 gnd.n2854 gnd.n2853 585
R4318 gnd.n2853 gnd.n1349 585
R4319 gnd.n2851 gnd.n1340 585
R4320 gnd.n5228 gnd.n1340 585
R4321 gnd.n2850 gnd.n2849 585
R4322 gnd.n2849 gnd.n1333 585
R4323 gnd.n2848 gnd.n1331 585
R4324 gnd.n5234 gnd.n1331 585
R4325 gnd.n2847 gnd.n2846 585
R4326 gnd.n2846 gnd.n1323 585
R4327 gnd.n2844 gnd.n1321 585
R4328 gnd.n5240 gnd.n1321 585
R4329 gnd.n2843 gnd.n2842 585
R4330 gnd.n2842 gnd.n1314 585
R4331 gnd.n2841 gnd.n1312 585
R4332 gnd.n5246 gnd.n1312 585
R4333 gnd.n2840 gnd.n2839 585
R4334 gnd.n2839 gnd.n1311 585
R4335 gnd.n2837 gnd.n1302 585
R4336 gnd.n5252 gnd.n1302 585
R4337 gnd.n2836 gnd.n2835 585
R4338 gnd.n2835 gnd.n1295 585
R4339 gnd.n2834 gnd.n1293 585
R4340 gnd.n5258 gnd.n1293 585
R4341 gnd.n2833 gnd.n2832 585
R4342 gnd.n2832 gnd.n1285 585
R4343 gnd.n2830 gnd.n1283 585
R4344 gnd.n5264 gnd.n1283 585
R4345 gnd.n2829 gnd.n2828 585
R4346 gnd.n2828 gnd.n1273 585
R4347 gnd.n2827 gnd.n1271 585
R4348 gnd.n5270 gnd.n1271 585
R4349 gnd.n2826 gnd.n1259 585
R4350 gnd.n1270 gnd.n1259 585
R4351 gnd.n5277 gnd.n1257 585
R4352 gnd.n5277 gnd.n5276 585
R4353 gnd.n5279 gnd.n5278 585
R4354 gnd.n5278 gnd.n1186 585
R4355 gnd.n8008 gnd.n251 585
R4356 gnd.n251 gnd.n250 585
R4357 gnd.n8010 gnd.n8009 585
R4358 gnd.n8011 gnd.n8010 585
R4359 gnd.n238 gnd.n237 585
R4360 gnd.n241 gnd.n238 585
R4361 gnd.n8019 gnd.n8018 585
R4362 gnd.n8018 gnd.n8017 585
R4363 gnd.n8020 gnd.n232 585
R4364 gnd.n232 gnd.n231 585
R4365 gnd.n8022 gnd.n8021 585
R4366 gnd.n8023 gnd.n8022 585
R4367 gnd.n218 gnd.n217 585
R4368 gnd.n228 gnd.n218 585
R4369 gnd.n8031 gnd.n8030 585
R4370 gnd.n8030 gnd.n8029 585
R4371 gnd.n8032 gnd.n212 585
R4372 gnd.n212 gnd.n211 585
R4373 gnd.n8034 gnd.n8033 585
R4374 gnd.n8035 gnd.n8034 585
R4375 gnd.n198 gnd.n197 585
R4376 gnd.n202 gnd.n198 585
R4377 gnd.n8043 gnd.n8042 585
R4378 gnd.n8042 gnd.n8041 585
R4379 gnd.n8044 gnd.n192 585
R4380 gnd.n199 gnd.n192 585
R4381 gnd.n8046 gnd.n8045 585
R4382 gnd.n8047 gnd.n8046 585
R4383 gnd.n180 gnd.n179 585
R4384 gnd.n189 gnd.n180 585
R4385 gnd.n8055 gnd.n8054 585
R4386 gnd.n8054 gnd.n8053 585
R4387 gnd.n8056 gnd.n174 585
R4388 gnd.n174 gnd.n173 585
R4389 gnd.n8058 gnd.n8057 585
R4390 gnd.n8059 gnd.n8058 585
R4391 gnd.n160 gnd.n159 585
R4392 gnd.n164 gnd.n160 585
R4393 gnd.n8067 gnd.n8066 585
R4394 gnd.n8066 gnd.n8065 585
R4395 gnd.n8068 gnd.n154 585
R4396 gnd.n161 gnd.n154 585
R4397 gnd.n8070 gnd.n8069 585
R4398 gnd.n8071 gnd.n8070 585
R4399 gnd.n142 gnd.n141 585
R4400 gnd.n151 gnd.n142 585
R4401 gnd.n8079 gnd.n8078 585
R4402 gnd.n8078 gnd.n8077 585
R4403 gnd.n8080 gnd.n137 585
R4404 gnd.n137 gnd.n136 585
R4405 gnd.n8082 gnd.n8081 585
R4406 gnd.n8083 gnd.n8082 585
R4407 gnd.n121 gnd.n119 585
R4408 gnd.n125 gnd.n121 585
R4409 gnd.n8091 gnd.n8090 585
R4410 gnd.n8090 gnd.n8089 585
R4411 gnd.n120 gnd.n112 585
R4412 gnd.n122 gnd.n120 585
R4413 gnd.n8094 gnd.n110 585
R4414 gnd.n110 gnd.n107 585
R4415 gnd.n8096 gnd.n8095 585
R4416 gnd.n8097 gnd.n8096 585
R4417 gnd.n7805 gnd.n109 585
R4418 gnd.n7822 gnd.n109 585
R4419 gnd.n7809 gnd.n7806 585
R4420 gnd.n7809 gnd.n7808 585
R4421 gnd.n7812 gnd.n7811 585
R4422 gnd.n7813 gnd.n7812 585
R4423 gnd.n7810 gnd.n7804 585
R4424 gnd.n7804 gnd.n7803 585
R4425 gnd.n7792 gnd.n501 585
R4426 gnd.n7784 gnd.n501 585
R4427 gnd.n7794 gnd.n7793 585
R4428 gnd.n7795 gnd.n7794 585
R4429 gnd.n7791 gnd.n514 585
R4430 gnd.n7791 gnd.n7790 585
R4431 gnd.n7764 gnd.n513 585
R4432 gnd.n7776 gnd.n513 585
R4433 gnd.n7765 gnd.n537 585
R4434 gnd.n7750 gnd.n537 585
R4435 gnd.n7767 gnd.n7766 585
R4436 gnd.n7768 gnd.n7767 585
R4437 gnd.n538 gnd.n536 585
R4438 gnd.n7744 gnd.n536 585
R4439 gnd.n7759 gnd.n7758 585
R4440 gnd.n7758 gnd.n7757 585
R4441 gnd.n541 gnd.n540 585
R4442 gnd.n2045 gnd.n541 585
R4443 gnd.n2033 gnd.n2032 585
R4444 gnd.n4652 gnd.n2033 585
R4445 gnd.n4661 gnd.n4660 585
R4446 gnd.n4660 gnd.n4659 585
R4447 gnd.n4662 gnd.n2026 585
R4448 gnd.n4640 gnd.n2026 585
R4449 gnd.n4664 gnd.n4663 585
R4450 gnd.n4665 gnd.n4664 585
R4451 gnd.n2012 gnd.n2011 585
R4452 gnd.n4624 gnd.n2012 585
R4453 gnd.n4673 gnd.n4672 585
R4454 gnd.n4672 gnd.n4671 585
R4455 gnd.n4674 gnd.n2006 585
R4456 gnd.n4615 gnd.n2006 585
R4457 gnd.n4676 gnd.n4675 585
R4458 gnd.n4677 gnd.n4676 585
R4459 gnd.n1991 gnd.n1990 585
R4460 gnd.n4607 gnd.n1991 585
R4461 gnd.n4685 gnd.n4684 585
R4462 gnd.n4684 gnd.n4683 585
R4463 gnd.n4686 gnd.n1985 585
R4464 gnd.n4601 gnd.n1985 585
R4465 gnd.n4688 gnd.n4687 585
R4466 gnd.n4689 gnd.n4688 585
R4467 gnd.n1971 gnd.n1970 585
R4468 gnd.n4593 gnd.n1971 585
R4469 gnd.n4697 gnd.n4696 585
R4470 gnd.n4696 gnd.n4695 585
R4471 gnd.n4698 gnd.n1965 585
R4472 gnd.n4587 gnd.n1965 585
R4473 gnd.n4700 gnd.n4699 585
R4474 gnd.n4701 gnd.n4700 585
R4475 gnd.n1949 gnd.n1948 585
R4476 gnd.n4579 gnd.n1949 585
R4477 gnd.n4709 gnd.n4708 585
R4478 gnd.n4708 gnd.n4707 585
R4479 gnd.n4710 gnd.n1942 585
R4480 gnd.n4573 gnd.n1942 585
R4481 gnd.n4712 gnd.n4711 585
R4482 gnd.n4713 gnd.n4712 585
R4483 gnd.n1943 gnd.n1862 585
R4484 gnd.n4716 gnd.n1862 585
R4485 gnd.n4834 gnd.n4833 585
R4486 gnd.n4832 gnd.n1861 585
R4487 gnd.n4831 gnd.n1860 585
R4488 gnd.n4836 gnd.n1860 585
R4489 gnd.n4830 gnd.n4829 585
R4490 gnd.n4828 gnd.n4827 585
R4491 gnd.n4826 gnd.n4825 585
R4492 gnd.n4824 gnd.n4823 585
R4493 gnd.n4822 gnd.n4821 585
R4494 gnd.n4820 gnd.n4819 585
R4495 gnd.n4818 gnd.n4817 585
R4496 gnd.n4816 gnd.n4815 585
R4497 gnd.n4814 gnd.n4813 585
R4498 gnd.n4812 gnd.n4811 585
R4499 gnd.n4810 gnd.n4809 585
R4500 gnd.n4808 gnd.n4807 585
R4501 gnd.n4806 gnd.n4805 585
R4502 gnd.n4804 gnd.n4803 585
R4503 gnd.n4802 gnd.n4801 585
R4504 gnd.n4799 gnd.n4798 585
R4505 gnd.n4797 gnd.n4796 585
R4506 gnd.n4795 gnd.n4794 585
R4507 gnd.n4793 gnd.n4792 585
R4508 gnd.n4791 gnd.n4790 585
R4509 gnd.n4789 gnd.n4788 585
R4510 gnd.n4787 gnd.n4786 585
R4511 gnd.n4785 gnd.n4784 585
R4512 gnd.n4782 gnd.n4781 585
R4513 gnd.n4780 gnd.n4779 585
R4514 gnd.n4778 gnd.n4777 585
R4515 gnd.n4776 gnd.n4775 585
R4516 gnd.n4774 gnd.n4773 585
R4517 gnd.n4772 gnd.n4771 585
R4518 gnd.n4770 gnd.n4769 585
R4519 gnd.n4768 gnd.n4767 585
R4520 gnd.n4766 gnd.n4765 585
R4521 gnd.n4764 gnd.n4763 585
R4522 gnd.n4762 gnd.n4761 585
R4523 gnd.n4760 gnd.n4759 585
R4524 gnd.n4758 gnd.n4757 585
R4525 gnd.n4756 gnd.n4755 585
R4526 gnd.n4754 gnd.n4753 585
R4527 gnd.n4752 gnd.n4751 585
R4528 gnd.n4750 gnd.n4749 585
R4529 gnd.n4748 gnd.n4747 585
R4530 gnd.n4746 gnd.n4745 585
R4531 gnd.n4744 gnd.n4743 585
R4532 gnd.n4742 gnd.n4741 585
R4533 gnd.n4740 gnd.n4739 585
R4534 gnd.n4738 gnd.n4737 585
R4535 gnd.n4736 gnd.n4735 585
R4536 gnd.n4734 gnd.n4733 585
R4537 gnd.n4732 gnd.n4731 585
R4538 gnd.n4730 gnd.n4729 585
R4539 gnd.n4728 gnd.n4727 585
R4540 gnd.n4726 gnd.n4725 585
R4541 gnd.n4724 gnd.n4723 585
R4542 gnd.n1932 gnd.n1925 585
R4543 gnd.n7879 gnd.n351 585
R4544 gnd.n7887 gnd.n7886 585
R4545 gnd.n7889 gnd.n7888 585
R4546 gnd.n7891 gnd.n7890 585
R4547 gnd.n7893 gnd.n7892 585
R4548 gnd.n7895 gnd.n7894 585
R4549 gnd.n7897 gnd.n7896 585
R4550 gnd.n7899 gnd.n7898 585
R4551 gnd.n7901 gnd.n7900 585
R4552 gnd.n7903 gnd.n7902 585
R4553 gnd.n7905 gnd.n7904 585
R4554 gnd.n7907 gnd.n7906 585
R4555 gnd.n7909 gnd.n7908 585
R4556 gnd.n7911 gnd.n7910 585
R4557 gnd.n7913 gnd.n7912 585
R4558 gnd.n7915 gnd.n7914 585
R4559 gnd.n7917 gnd.n7916 585
R4560 gnd.n7919 gnd.n7918 585
R4561 gnd.n7921 gnd.n7920 585
R4562 gnd.n7924 gnd.n7923 585
R4563 gnd.n7922 gnd.n331 585
R4564 gnd.n7929 gnd.n7928 585
R4565 gnd.n7931 gnd.n7930 585
R4566 gnd.n7933 gnd.n7932 585
R4567 gnd.n7935 gnd.n7934 585
R4568 gnd.n7937 gnd.n7936 585
R4569 gnd.n7939 gnd.n7938 585
R4570 gnd.n7941 gnd.n7940 585
R4571 gnd.n7943 gnd.n7942 585
R4572 gnd.n7945 gnd.n7944 585
R4573 gnd.n7947 gnd.n7946 585
R4574 gnd.n7949 gnd.n7948 585
R4575 gnd.n7951 gnd.n7950 585
R4576 gnd.n7953 gnd.n7952 585
R4577 gnd.n7955 gnd.n7954 585
R4578 gnd.n7957 gnd.n7956 585
R4579 gnd.n7959 gnd.n7958 585
R4580 gnd.n7961 gnd.n7960 585
R4581 gnd.n7963 gnd.n7962 585
R4582 gnd.n7965 gnd.n7964 585
R4583 gnd.n7967 gnd.n7966 585
R4584 gnd.n7972 gnd.n7971 585
R4585 gnd.n7974 gnd.n7973 585
R4586 gnd.n7976 gnd.n7975 585
R4587 gnd.n7978 gnd.n7977 585
R4588 gnd.n7980 gnd.n7979 585
R4589 gnd.n7982 gnd.n7981 585
R4590 gnd.n7984 gnd.n7983 585
R4591 gnd.n7986 gnd.n7985 585
R4592 gnd.n7988 gnd.n7987 585
R4593 gnd.n7990 gnd.n7989 585
R4594 gnd.n7992 gnd.n7991 585
R4595 gnd.n7994 gnd.n7993 585
R4596 gnd.n7996 gnd.n7995 585
R4597 gnd.n7998 gnd.n7997 585
R4598 gnd.n7999 gnd.n295 585
R4599 gnd.n8001 gnd.n8000 585
R4600 gnd.n256 gnd.n255 585
R4601 gnd.n8005 gnd.n8004 585
R4602 gnd.n8004 gnd.n8003 585
R4603 gnd.n7881 gnd.n7880 585
R4604 gnd.n7880 gnd.n250 585
R4605 gnd.n7878 gnd.n248 585
R4606 gnd.n8011 gnd.n248 585
R4607 gnd.n7877 gnd.n7876 585
R4608 gnd.n7876 gnd.n241 585
R4609 gnd.n7875 gnd.n239 585
R4610 gnd.n8017 gnd.n239 585
R4611 gnd.n7874 gnd.n7873 585
R4612 gnd.n7873 gnd.n231 585
R4613 gnd.n7871 gnd.n229 585
R4614 gnd.n8023 gnd.n229 585
R4615 gnd.n7870 gnd.n7869 585
R4616 gnd.n7869 gnd.n228 585
R4617 gnd.n7868 gnd.n220 585
R4618 gnd.n8029 gnd.n220 585
R4619 gnd.n7867 gnd.n7866 585
R4620 gnd.n7866 gnd.n211 585
R4621 gnd.n7864 gnd.n209 585
R4622 gnd.n8035 gnd.n209 585
R4623 gnd.n7863 gnd.n7862 585
R4624 gnd.n7862 gnd.n202 585
R4625 gnd.n7861 gnd.n200 585
R4626 gnd.n8041 gnd.n200 585
R4627 gnd.n7860 gnd.n7859 585
R4628 gnd.n7859 gnd.n199 585
R4629 gnd.n7857 gnd.n190 585
R4630 gnd.n8047 gnd.n190 585
R4631 gnd.n7856 gnd.n7855 585
R4632 gnd.n7855 gnd.n189 585
R4633 gnd.n7854 gnd.n181 585
R4634 gnd.n8053 gnd.n181 585
R4635 gnd.n7853 gnd.n7852 585
R4636 gnd.n7852 gnd.n173 585
R4637 gnd.n7850 gnd.n171 585
R4638 gnd.n8059 gnd.n171 585
R4639 gnd.n7849 gnd.n7848 585
R4640 gnd.n7848 gnd.n164 585
R4641 gnd.n7847 gnd.n162 585
R4642 gnd.n8065 gnd.n162 585
R4643 gnd.n7846 gnd.n7845 585
R4644 gnd.n7845 gnd.n161 585
R4645 gnd.n7843 gnd.n152 585
R4646 gnd.n8071 gnd.n152 585
R4647 gnd.n7842 gnd.n7841 585
R4648 gnd.n7841 gnd.n151 585
R4649 gnd.n7840 gnd.n143 585
R4650 gnd.n8077 gnd.n143 585
R4651 gnd.n7839 gnd.n7838 585
R4652 gnd.n7838 gnd.n136 585
R4653 gnd.n7836 gnd.n134 585
R4654 gnd.n8083 gnd.n134 585
R4655 gnd.n7835 gnd.n7834 585
R4656 gnd.n7834 gnd.n125 585
R4657 gnd.n7833 gnd.n123 585
R4658 gnd.n8089 gnd.n123 585
R4659 gnd.n7832 gnd.n7831 585
R4660 gnd.n7831 gnd.n122 585
R4661 gnd.n7830 gnd.n486 585
R4662 gnd.n7830 gnd.n107 585
R4663 gnd.n7819 gnd.n106 585
R4664 gnd.n8097 gnd.n106 585
R4665 gnd.n7821 gnd.n7820 585
R4666 gnd.n7822 gnd.n7821 585
R4667 gnd.n7818 gnd.n492 585
R4668 gnd.n7808 gnd.n492 585
R4669 gnd.n498 gnd.n493 585
R4670 gnd.n7813 gnd.n498 585
R4671 gnd.n7781 gnd.n503 585
R4672 gnd.n7803 gnd.n503 585
R4673 gnd.n7783 gnd.n7782 585
R4674 gnd.n7784 gnd.n7783 585
R4675 gnd.n7780 gnd.n511 585
R4676 gnd.n7795 gnd.n511 585
R4677 gnd.n7779 gnd.n516 585
R4678 gnd.n7790 gnd.n516 585
R4679 gnd.n7778 gnd.n7777 585
R4680 gnd.n7777 gnd.n7776 585
R4681 gnd.n525 gnd.n523 585
R4682 gnd.n7750 gnd.n525 585
R4683 gnd.n7747 gnd.n533 585
R4684 gnd.n7768 gnd.n533 585
R4685 gnd.n7746 gnd.n7745 585
R4686 gnd.n7745 gnd.n7744 585
R4687 gnd.n550 gnd.n543 585
R4688 gnd.n7757 gnd.n543 585
R4689 gnd.n2043 gnd.n2042 585
R4690 gnd.n2045 gnd.n2043 585
R4691 gnd.n4654 gnd.n4653 585
R4692 gnd.n4653 gnd.n4652 585
R4693 gnd.n2041 gnd.n2035 585
R4694 gnd.n4659 gnd.n2035 585
R4695 gnd.n4620 gnd.n2051 585
R4696 gnd.n4640 gnd.n2051 585
R4697 gnd.n4621 gnd.n2024 585
R4698 gnd.n4665 gnd.n2024 585
R4699 gnd.n4623 gnd.n4622 585
R4700 gnd.n4624 gnd.n4623 585
R4701 gnd.n4618 gnd.n2014 585
R4702 gnd.n4671 gnd.n2014 585
R4703 gnd.n4617 gnd.n4616 585
R4704 gnd.n4616 gnd.n4615 585
R4705 gnd.n2056 gnd.n2003 585
R4706 gnd.n4677 gnd.n2003 585
R4707 gnd.n4606 gnd.n4605 585
R4708 gnd.n4607 gnd.n4606 585
R4709 gnd.n4604 gnd.n1993 585
R4710 gnd.n4683 gnd.n1993 585
R4711 gnd.n4603 gnd.n4602 585
R4712 gnd.n4602 gnd.n4601 585
R4713 gnd.n2061 gnd.n1983 585
R4714 gnd.n4689 gnd.n1983 585
R4715 gnd.n4592 gnd.n4591 585
R4716 gnd.n4593 gnd.n4592 585
R4717 gnd.n4590 gnd.n1973 585
R4718 gnd.n4695 gnd.n1973 585
R4719 gnd.n4589 gnd.n4588 585
R4720 gnd.n4588 gnd.n4587 585
R4721 gnd.n2124 gnd.n1962 585
R4722 gnd.n4701 gnd.n1962 585
R4723 gnd.n4578 gnd.n4577 585
R4724 gnd.n4579 gnd.n4578 585
R4725 gnd.n4576 gnd.n1951 585
R4726 gnd.n4707 gnd.n1951 585
R4727 gnd.n4575 gnd.n4574 585
R4728 gnd.n4574 gnd.n4573 585
R4729 gnd.n1933 gnd.n1931 585
R4730 gnd.n4713 gnd.n1933 585
R4731 gnd.n4718 gnd.n4717 585
R4732 gnd.n4717 gnd.n4716 585
R4733 gnd.n1135 gnd.n1134 585
R4734 gnd.n1396 gnd.n1135 585
R4735 gnd.n7722 gnd.n7720 585
R4736 gnd.n7722 gnd.n7721 585
R4737 gnd.n7724 gnd.n7723 585
R4738 gnd.n7723 gnd.n105 585
R4739 gnd.n7725 gnd.n565 585
R4740 gnd.n565 gnd.n491 585
R4741 gnd.n7727 gnd.n7726 585
R4742 gnd.n7727 gnd.n500 585
R4743 gnd.n7728 gnd.n563 585
R4744 gnd.n7728 gnd.n497 585
R4745 gnd.n7730 gnd.n7729 585
R4746 gnd.n7729 gnd.n502 585
R4747 gnd.n564 gnd.n561 585
R4748 gnd.n564 gnd.n522 585
R4749 gnd.n7734 gnd.n558 585
R4750 gnd.n558 gnd.n510 585
R4751 gnd.n7736 gnd.n7735 585
R4752 gnd.n7736 gnd.n515 585
R4753 gnd.n7737 gnd.n557 585
R4754 gnd.n7737 gnd.n526 585
R4755 gnd.n7739 gnd.n7738 585
R4756 gnd.n7738 gnd.n534 585
R4757 gnd.n7740 gnd.n552 585
R4758 gnd.n552 gnd.n532 585
R4759 gnd.n7742 gnd.n7741 585
R4760 gnd.n7743 gnd.n7742 585
R4761 gnd.n553 gnd.n551 585
R4762 gnd.n551 gnd.n542 585
R4763 gnd.n4650 gnd.n4649 585
R4764 gnd.n4651 gnd.n4650 585
R4765 gnd.n2047 gnd.n2046 585
R4766 gnd.n2046 gnd.n2037 585
R4767 gnd.n4644 gnd.n4643 585
R4768 gnd.n4643 gnd.n2034 585
R4769 gnd.n4642 gnd.n2049 585
R4770 gnd.n4642 gnd.n4641 585
R4771 gnd.n2108 gnd.n2050 585
R4772 gnd.n2050 gnd.n2023 585
R4773 gnd.n2110 gnd.n2109 585
R4774 gnd.n2109 gnd.n2016 585
R4775 gnd.n2111 gnd.n2102 585
R4776 gnd.n2102 gnd.n2013 585
R4777 gnd.n2113 gnd.n2112 585
R4778 gnd.n2113 gnd.n2005 585
R4779 gnd.n2114 gnd.n2101 585
R4780 gnd.n2114 gnd.n2002 585
R4781 gnd.n2116 gnd.n2115 585
R4782 gnd.n2115 gnd.n1995 585
R4783 gnd.n2117 gnd.n2064 585
R4784 gnd.n2064 gnd.n1992 585
R4785 gnd.n2119 gnd.n2118 585
R4786 gnd.n2120 gnd.n2119 585
R4787 gnd.n2065 gnd.n2063 585
R4788 gnd.n2063 gnd.n1982 585
R4789 gnd.n2095 gnd.n2094 585
R4790 gnd.n2094 gnd.n1975 585
R4791 gnd.n2093 gnd.n2067 585
R4792 gnd.n2093 gnd.n1972 585
R4793 gnd.n2092 gnd.n2091 585
R4794 gnd.n2092 gnd.n1964 585
R4795 gnd.n2069 gnd.n2068 585
R4796 gnd.n2068 gnd.n1961 585
R4797 gnd.n2087 gnd.n2086 585
R4798 gnd.n2086 gnd.n1953 585
R4799 gnd.n2085 gnd.n2071 585
R4800 gnd.n2085 gnd.n1950 585
R4801 gnd.n2084 gnd.n2083 585
R4802 gnd.n2084 gnd.n1941 585
R4803 gnd.n2073 gnd.n2072 585
R4804 gnd.n2072 gnd.n1936 585
R4805 gnd.n2079 gnd.n2078 585
R4806 gnd.n2078 gnd.n1934 585
R4807 gnd.n2077 gnd.n2076 585
R4808 gnd.n2077 gnd.n1859 585
R4809 gnd.n1819 gnd.n1818 585
R4810 gnd.n4837 gnd.n1819 585
R4811 gnd.n4840 gnd.n4839 585
R4812 gnd.n4839 gnd.n4838 585
R4813 gnd.n4841 gnd.n1813 585
R4814 gnd.n1820 gnd.n1813 585
R4815 gnd.n4843 gnd.n4842 585
R4816 gnd.n4844 gnd.n4843 585
R4817 gnd.n1814 gnd.n1810 585
R4818 gnd.n4845 gnd.n1810 585
R4819 gnd.n4397 gnd.n2137 585
R4820 gnd.n2137 gnd.n1809 585
R4821 gnd.n4399 gnd.n4398 585
R4822 gnd.n4400 gnd.n4399 585
R4823 gnd.n2138 gnd.n2136 585
R4824 gnd.n2136 gnd.n2135 585
R4825 gnd.n4391 gnd.n4390 585
R4826 gnd.n4390 gnd.n4389 585
R4827 gnd.n2141 gnd.n2140 585
R4828 gnd.n2142 gnd.n2141 585
R4829 gnd.n4378 gnd.n4377 585
R4830 gnd.n4379 gnd.n4378 585
R4831 gnd.n2150 gnd.n2149 585
R4832 gnd.n2156 gnd.n2149 585
R4833 gnd.n4373 gnd.n4372 585
R4834 gnd.n4372 gnd.n4371 585
R4835 gnd.n2153 gnd.n2152 585
R4836 gnd.n2154 gnd.n2153 585
R4837 gnd.n4362 gnd.n4361 585
R4838 gnd.n4363 gnd.n4362 585
R4839 gnd.n2165 gnd.n2164 585
R4840 gnd.n2164 gnd.n2163 585
R4841 gnd.n4357 gnd.n4356 585
R4842 gnd.n4356 gnd.n4355 585
R4843 gnd.n2168 gnd.n2167 585
R4844 gnd.n2169 gnd.n2168 585
R4845 gnd.n4346 gnd.n4345 585
R4846 gnd.n4347 gnd.n4346 585
R4847 gnd.n2178 gnd.n2177 585
R4848 gnd.n2177 gnd.n2176 585
R4849 gnd.n4341 gnd.n4340 585
R4850 gnd.n4340 gnd.n4339 585
R4851 gnd.n2181 gnd.n2180 585
R4852 gnd.n3687 gnd.n2181 585
R4853 gnd.n4330 gnd.n4329 585
R4854 gnd.n4331 gnd.n4330 585
R4855 gnd.n2189 gnd.n2188 585
R4856 gnd.n3884 gnd.n2188 585
R4857 gnd.n4325 gnd.n4324 585
R4858 gnd.n4324 gnd.n4323 585
R4859 gnd.n2192 gnd.n2191 585
R4860 gnd.n3657 gnd.n2192 585
R4861 gnd.n4314 gnd.n4313 585
R4862 gnd.n4315 gnd.n4314 585
R4863 gnd.n2202 gnd.n2201 585
R4864 gnd.n3670 gnd.n2201 585
R4865 gnd.n4309 gnd.n4308 585
R4866 gnd.n4308 gnd.n4307 585
R4867 gnd.n2205 gnd.n2204 585
R4868 gnd.n2214 gnd.n2205 585
R4869 gnd.n4298 gnd.n4297 585
R4870 gnd.n4299 gnd.n4298 585
R4871 gnd.n2217 gnd.n2216 585
R4872 gnd.n3646 gnd.n2216 585
R4873 gnd.n4293 gnd.n4292 585
R4874 gnd.n4292 gnd.n4291 585
R4875 gnd.n2220 gnd.n2219 585
R4876 gnd.n3638 gnd.n2220 585
R4877 gnd.n4282 gnd.n4281 585
R4878 gnd.n4283 gnd.n4282 585
R4879 gnd.n2230 gnd.n2229 585
R4880 gnd.n3631 gnd.n2229 585
R4881 gnd.n4277 gnd.n4276 585
R4882 gnd.n4276 gnd.n4275 585
R4883 gnd.n2233 gnd.n2232 585
R4884 gnd.n3622 gnd.n2233 585
R4885 gnd.n4266 gnd.n4265 585
R4886 gnd.n4267 gnd.n4266 585
R4887 gnd.n2244 gnd.n2243 585
R4888 gnd.n3935 gnd.n2243 585
R4889 gnd.n4261 gnd.n4260 585
R4890 gnd.n4260 gnd.n4259 585
R4891 gnd.n2247 gnd.n2246 585
R4892 gnd.n3608 gnd.n2247 585
R4893 gnd.n4250 gnd.n4249 585
R4894 gnd.n4251 gnd.n4250 585
R4895 gnd.n2257 gnd.n2256 585
R4896 gnd.n3601 gnd.n2256 585
R4897 gnd.n4245 gnd.n4244 585
R4898 gnd.n4244 gnd.n4243 585
R4899 gnd.n2260 gnd.n2259 585
R4900 gnd.n3593 gnd.n2260 585
R4901 gnd.n4234 gnd.n4233 585
R4902 gnd.n4235 gnd.n4234 585
R4903 gnd.n2271 gnd.n2270 585
R4904 gnd.n3964 gnd.n2270 585
R4905 gnd.n4229 gnd.n4228 585
R4906 gnd.n4228 gnd.n4227 585
R4907 gnd.n2274 gnd.n2273 585
R4908 gnd.n3580 gnd.n2274 585
R4909 gnd.n4218 gnd.n4217 585
R4910 gnd.n4219 gnd.n4218 585
R4911 gnd.n2285 gnd.n2284 585
R4912 gnd.n3980 gnd.n2284 585
R4913 gnd.n4213 gnd.n4212 585
R4914 gnd.n4212 gnd.n4211 585
R4915 gnd.n2288 gnd.n2287 585
R4916 gnd.n3566 gnd.n2288 585
R4917 gnd.n4202 gnd.n4201 585
R4918 gnd.n4203 gnd.n4202 585
R4919 gnd.n2298 gnd.n2297 585
R4920 gnd.n3996 gnd.n2297 585
R4921 gnd.n4197 gnd.n4196 585
R4922 gnd.n4196 gnd.n4195 585
R4923 gnd.n2301 gnd.n2300 585
R4924 gnd.n3553 gnd.n2301 585
R4925 gnd.n4186 gnd.n4185 585
R4926 gnd.n4187 gnd.n4186 585
R4927 gnd.n2312 gnd.n2311 585
R4928 gnd.n4012 gnd.n2311 585
R4929 gnd.n4181 gnd.n4180 585
R4930 gnd.n4180 gnd.n4179 585
R4931 gnd.n2315 gnd.n2314 585
R4932 gnd.n3545 gnd.n2315 585
R4933 gnd.n4170 gnd.n4169 585
R4934 gnd.n4171 gnd.n4170 585
R4935 gnd.n2326 gnd.n2325 585
R4936 gnd.n2332 gnd.n2325 585
R4937 gnd.n4165 gnd.n4164 585
R4938 gnd.n4164 gnd.n4163 585
R4939 gnd.n2329 gnd.n2328 585
R4940 gnd.n3526 gnd.n2329 585
R4941 gnd.n4154 gnd.n4153 585
R4942 gnd.n4155 gnd.n4154 585
R4943 gnd.n2341 gnd.n2340 585
R4944 gnd.n3517 gnd.n2340 585
R4945 gnd.n4149 gnd.n4148 585
R4946 gnd.n4148 gnd.n4147 585
R4947 gnd.n2344 gnd.n2343 585
R4948 gnd.n3508 gnd.n2344 585
R4949 gnd.n4138 gnd.n4137 585
R4950 gnd.n4139 gnd.n4138 585
R4951 gnd.n2355 gnd.n2354 585
R4952 gnd.n4049 gnd.n2354 585
R4953 gnd.n4133 gnd.n4132 585
R4954 gnd.n4132 gnd.n4131 585
R4955 gnd.n2358 gnd.n2357 585
R4956 gnd.n3495 gnd.n2358 585
R4957 gnd.n4122 gnd.n4121 585
R4958 gnd.n4123 gnd.n4122 585
R4959 gnd.n2367 gnd.n2366 585
R4960 gnd.n3486 gnd.n2366 585
R4961 gnd.n4117 gnd.n4116 585
R4962 gnd.n4116 gnd.n4115 585
R4963 gnd.n2370 gnd.n2369 585
R4964 gnd.n3476 gnd.n2370 585
R4965 gnd.n4106 gnd.n4105 585
R4966 gnd.n4107 gnd.n4106 585
R4967 gnd.n2381 gnd.n2380 585
R4968 gnd.n4078 gnd.n2380 585
R4969 gnd.n4101 gnd.n4100 585
R4970 gnd.n4100 gnd.n4099 585
R4971 gnd.n2384 gnd.n2383 585
R4972 gnd.n2392 gnd.n2384 585
R4973 gnd.n4090 gnd.n4089 585
R4974 gnd.n4091 gnd.n4090 585
R4975 gnd.n1700 gnd.n1699 585
R4976 gnd.n3464 gnd.n1700 585
R4977 gnd.n4970 gnd.n4969 585
R4978 gnd.n4969 gnd.t109 585
R4979 gnd.n4971 gnd.n1694 585
R4980 gnd.n3455 gnd.n1694 585
R4981 gnd.n4973 gnd.n4972 585
R4982 gnd.n4974 gnd.n4973 585
R4983 gnd.n1695 gnd.n1693 585
R4984 gnd.n1693 gnd.n1688 585
R4985 gnd.n3432 gnd.n3431 585
R4986 gnd.n3432 gnd.n1662 585
R4987 gnd.n3434 gnd.n3433 585
R4988 gnd.n3433 gnd.n1630 585
R4989 gnd.n3435 gnd.n2496 585
R4990 gnd.n2496 gnd.n2494 585
R4991 gnd.n3437 gnd.n3436 585
R4992 gnd.n3438 gnd.n3437 585
R4993 gnd.n2497 gnd.n2495 585
R4994 gnd.n2495 gnd.n2492 585
R4995 gnd.n3423 gnd.n3422 585
R4996 gnd.n3422 gnd.n3421 585
R4997 gnd.n2500 gnd.n2499 585
R4998 gnd.n2509 gnd.n2500 585
R4999 gnd.n3412 gnd.n3411 585
R5000 gnd.n3413 gnd.n3412 585
R5001 gnd.n2511 gnd.n2510 585
R5002 gnd.n2510 gnd.n2507 585
R5003 gnd.n3407 gnd.n3406 585
R5004 gnd.n3406 gnd.n3405 585
R5005 gnd.n2514 gnd.n2513 585
R5006 gnd.n2515 gnd.n2514 585
R5007 gnd.n3396 gnd.n3395 585
R5008 gnd.n3397 gnd.n3396 585
R5009 gnd.n2525 gnd.n2524 585
R5010 gnd.n2524 gnd.n2522 585
R5011 gnd.n3391 gnd.n3390 585
R5012 gnd.n3390 gnd.n3389 585
R5013 gnd.n2528 gnd.n2527 585
R5014 gnd.n2529 gnd.n2528 585
R5015 gnd.n3380 gnd.n3379 585
R5016 gnd.n3381 gnd.n3380 585
R5017 gnd.n2538 gnd.n2537 585
R5018 gnd.n2544 gnd.n2537 585
R5019 gnd.n3375 gnd.n3374 585
R5020 gnd.n3374 gnd.n3373 585
R5021 gnd.n2541 gnd.n2540 585
R5022 gnd.n2542 gnd.n2541 585
R5023 gnd.n2565 gnd.n2564 585
R5024 gnd.n3352 gnd.n2565 585
R5025 gnd.n3354 gnd.n2561 585
R5026 gnd.n3354 gnd.n3353 585
R5027 gnd.n3356 gnd.n3355 585
R5028 gnd.n3355 gnd.n1567 585
R5029 gnd.n3357 gnd.n2556 585
R5030 gnd.n2556 gnd.n1556 585
R5031 gnd.n3359 gnd.n3358 585
R5032 gnd.n3360 gnd.n3359 585
R5033 gnd.n2557 gnd.n2555 585
R5034 gnd.n2555 gnd.n1549 585
R5035 gnd.n3172 gnd.n3171 585
R5036 gnd.n3172 gnd.n1546 585
R5037 gnd.n3173 gnd.n3167 585
R5038 gnd.n3173 gnd.n1539 585
R5039 gnd.n3175 gnd.n3174 585
R5040 gnd.n3174 gnd.n1536 585
R5041 gnd.n3176 gnd.n3162 585
R5042 gnd.n3162 gnd.n1528 585
R5043 gnd.n3178 gnd.n3177 585
R5044 gnd.n3178 gnd.n1525 585
R5045 gnd.n3179 gnd.n3161 585
R5046 gnd.n3179 gnd.n1518 585
R5047 gnd.n3181 gnd.n3180 585
R5048 gnd.n3180 gnd.n1515 585
R5049 gnd.n3182 gnd.n2748 585
R5050 gnd.n2748 gnd.n1507 585
R5051 gnd.n3184 gnd.n3183 585
R5052 gnd.n3185 gnd.n3184 585
R5053 gnd.n2749 gnd.n2747 585
R5054 gnd.n2747 gnd.n1498 585
R5055 gnd.n3155 gnd.n3154 585
R5056 gnd.n3154 gnd.n1495 585
R5057 gnd.n3153 gnd.n2751 585
R5058 gnd.n3153 gnd.n1487 585
R5059 gnd.n3152 gnd.n3151 585
R5060 gnd.n3152 gnd.n1484 585
R5061 gnd.n2753 gnd.n2752 585
R5062 gnd.n2752 gnd.n1477 585
R5063 gnd.n3147 gnd.n3146 585
R5064 gnd.n3146 gnd.n1474 585
R5065 gnd.n3145 gnd.n2755 585
R5066 gnd.n3145 gnd.n1466 585
R5067 gnd.n3144 gnd.n2757 585
R5068 gnd.n3144 gnd.n3143 585
R5069 gnd.n3072 gnd.n2756 585
R5070 gnd.n2756 gnd.n1457 585
R5071 gnd.n3074 gnd.n3073 585
R5072 gnd.n3073 gnd.n1454 585
R5073 gnd.n3075 gnd.n3065 585
R5074 gnd.n3065 gnd.n1446 585
R5075 gnd.n3077 gnd.n3076 585
R5076 gnd.n3077 gnd.n1443 585
R5077 gnd.n3078 gnd.n3064 585
R5078 gnd.n3078 gnd.n1436 585
R5079 gnd.n3080 gnd.n3079 585
R5080 gnd.n3079 gnd.n1433 585
R5081 gnd.n3081 gnd.n2779 585
R5082 gnd.n2779 gnd.n1426 585
R5083 gnd.n3083 gnd.n3082 585
R5084 gnd.n3084 gnd.n3083 585
R5085 gnd.n2780 gnd.n2778 585
R5086 gnd.n2778 gnd.n1415 585
R5087 gnd.n3058 gnd.n3057 585
R5088 gnd.n3057 gnd.n1412 585
R5089 gnd.n3056 gnd.n2782 585
R5090 gnd.n3056 gnd.n3055 585
R5091 gnd.n2816 gnd.n2783 585
R5092 gnd.n2792 gnd.n2783 585
R5093 gnd.n2818 gnd.n2817 585
R5094 gnd.n2818 gnd.n2799 585
R5095 gnd.n2820 gnd.n2819 585
R5096 gnd.n2819 gnd.n2797 585
R5097 gnd.n2821 gnd.n2809 585
R5098 gnd.n2809 gnd.n2808 585
R5099 gnd.n2823 gnd.n2822 585
R5100 gnd.n2824 gnd.n2823 585
R5101 gnd.n4847 gnd.n4846 585
R5102 gnd.n4846 gnd.n4845 585
R5103 gnd.n4848 gnd.n1806 585
R5104 gnd.n1809 gnd.n1806 585
R5105 gnd.n4849 gnd.n1805 585
R5106 gnd.n4400 gnd.n1805 585
R5107 gnd.n2134 gnd.n1803 585
R5108 gnd.n2135 gnd.n2134 585
R5109 gnd.n4853 gnd.n1802 585
R5110 gnd.n4389 gnd.n1802 585
R5111 gnd.n4854 gnd.n1801 585
R5112 gnd.n2142 gnd.n1801 585
R5113 gnd.n4855 gnd.n1800 585
R5114 gnd.n4379 gnd.n1800 585
R5115 gnd.n2155 gnd.n1798 585
R5116 gnd.n2156 gnd.n2155 585
R5117 gnd.n4859 gnd.n1797 585
R5118 gnd.n4371 gnd.n1797 585
R5119 gnd.n4860 gnd.n1796 585
R5120 gnd.n2154 gnd.n1796 585
R5121 gnd.n4861 gnd.n1795 585
R5122 gnd.n4363 gnd.n1795 585
R5123 gnd.n2162 gnd.n1793 585
R5124 gnd.n2163 gnd.n2162 585
R5125 gnd.n4865 gnd.n1792 585
R5126 gnd.n4355 gnd.n1792 585
R5127 gnd.n4866 gnd.n1791 585
R5128 gnd.n2169 gnd.n1791 585
R5129 gnd.n4867 gnd.n1790 585
R5130 gnd.n4347 gnd.n1790 585
R5131 gnd.n2175 gnd.n1788 585
R5132 gnd.n2176 gnd.n2175 585
R5133 gnd.n4871 gnd.n1787 585
R5134 gnd.n4339 gnd.n1787 585
R5135 gnd.n4872 gnd.n1786 585
R5136 gnd.n3687 gnd.n1786 585
R5137 gnd.n4873 gnd.n1785 585
R5138 gnd.n4331 gnd.n1785 585
R5139 gnd.n3679 gnd.n1783 585
R5140 gnd.n3884 gnd.n3679 585
R5141 gnd.n4877 gnd.n1782 585
R5142 gnd.n4323 gnd.n1782 585
R5143 gnd.n4878 gnd.n1781 585
R5144 gnd.n3657 gnd.n1781 585
R5145 gnd.n4879 gnd.n1780 585
R5146 gnd.n4315 gnd.n1780 585
R5147 gnd.n3669 gnd.n1778 585
R5148 gnd.n3670 gnd.n3669 585
R5149 gnd.n4883 gnd.n1777 585
R5150 gnd.n4307 gnd.n1777 585
R5151 gnd.n4884 gnd.n1776 585
R5152 gnd.n2214 gnd.n1776 585
R5153 gnd.n4885 gnd.n1775 585
R5154 gnd.n4299 gnd.n1775 585
R5155 gnd.n3645 gnd.n1773 585
R5156 gnd.n3646 gnd.n3645 585
R5157 gnd.n4889 gnd.n1772 585
R5158 gnd.n4291 gnd.n1772 585
R5159 gnd.n4890 gnd.n1771 585
R5160 gnd.n3638 gnd.n1771 585
R5161 gnd.n4891 gnd.n1770 585
R5162 gnd.n4283 gnd.n1770 585
R5163 gnd.n3630 gnd.n1768 585
R5164 gnd.n3631 gnd.n3630 585
R5165 gnd.n4895 gnd.n1767 585
R5166 gnd.n4275 gnd.n1767 585
R5167 gnd.n4896 gnd.n1766 585
R5168 gnd.n3622 gnd.n1766 585
R5169 gnd.n4897 gnd.n1765 585
R5170 gnd.n4267 gnd.n1765 585
R5171 gnd.n3616 gnd.n1763 585
R5172 gnd.n3935 gnd.n3616 585
R5173 gnd.n4901 gnd.n1762 585
R5174 gnd.n4259 gnd.n1762 585
R5175 gnd.n4902 gnd.n1761 585
R5176 gnd.n3608 gnd.n1761 585
R5177 gnd.n4903 gnd.n1760 585
R5178 gnd.n4251 gnd.n1760 585
R5179 gnd.n3600 gnd.n1758 585
R5180 gnd.n3601 gnd.n3600 585
R5181 gnd.n4907 gnd.n1757 585
R5182 gnd.n4243 gnd.n1757 585
R5183 gnd.n4908 gnd.n1756 585
R5184 gnd.n3593 gnd.n1756 585
R5185 gnd.n4909 gnd.n1755 585
R5186 gnd.n4235 gnd.n1755 585
R5187 gnd.n3963 gnd.n1753 585
R5188 gnd.n3964 gnd.n3963 585
R5189 gnd.n4913 gnd.n1752 585
R5190 gnd.n4227 gnd.n1752 585
R5191 gnd.n4914 gnd.n1751 585
R5192 gnd.n3580 gnd.n1751 585
R5193 gnd.n4915 gnd.n1750 585
R5194 gnd.n4219 gnd.n1750 585
R5195 gnd.n3979 gnd.n1748 585
R5196 gnd.n3980 gnd.n3979 585
R5197 gnd.n4919 gnd.n1747 585
R5198 gnd.n4211 gnd.n1747 585
R5199 gnd.n4920 gnd.n1746 585
R5200 gnd.n3566 gnd.n1746 585
R5201 gnd.n4921 gnd.n1745 585
R5202 gnd.n4203 gnd.n1745 585
R5203 gnd.n3995 gnd.n1743 585
R5204 gnd.n3996 gnd.n3995 585
R5205 gnd.n4925 gnd.n1742 585
R5206 gnd.n4195 gnd.n1742 585
R5207 gnd.n4926 gnd.n1741 585
R5208 gnd.n3553 gnd.n1741 585
R5209 gnd.n4927 gnd.n1740 585
R5210 gnd.n4187 gnd.n1740 585
R5211 gnd.n4011 gnd.n1738 585
R5212 gnd.n4012 gnd.n4011 585
R5213 gnd.n4931 gnd.n1737 585
R5214 gnd.n4179 gnd.n1737 585
R5215 gnd.n4932 gnd.n1736 585
R5216 gnd.n3545 gnd.n1736 585
R5217 gnd.n4933 gnd.n1735 585
R5218 gnd.n4171 gnd.n1735 585
R5219 gnd.n2331 gnd.n1733 585
R5220 gnd.n2332 gnd.n2331 585
R5221 gnd.n4937 gnd.n1732 585
R5222 gnd.n4163 gnd.n1732 585
R5223 gnd.n4938 gnd.n1731 585
R5224 gnd.n3526 gnd.n1731 585
R5225 gnd.n4939 gnd.n1730 585
R5226 gnd.n4155 gnd.n1730 585
R5227 gnd.n3516 gnd.n1728 585
R5228 gnd.n3517 gnd.n3516 585
R5229 gnd.n4943 gnd.n1727 585
R5230 gnd.n4147 gnd.n1727 585
R5231 gnd.n4944 gnd.n1726 585
R5232 gnd.n3508 gnd.n1726 585
R5233 gnd.n4945 gnd.n1725 585
R5234 gnd.n4139 gnd.n1725 585
R5235 gnd.n3503 gnd.n1723 585
R5236 gnd.n4049 gnd.n3503 585
R5237 gnd.n4949 gnd.n1722 585
R5238 gnd.n4131 gnd.n1722 585
R5239 gnd.n4950 gnd.n1721 585
R5240 gnd.n3495 gnd.n1721 585
R5241 gnd.n4951 gnd.n1720 585
R5242 gnd.n4123 gnd.n1720 585
R5243 gnd.n3485 gnd.n1718 585
R5244 gnd.n3486 gnd.n3485 585
R5245 gnd.n4955 gnd.n1717 585
R5246 gnd.n4115 gnd.n1717 585
R5247 gnd.n4956 gnd.n1716 585
R5248 gnd.n3476 gnd.n1716 585
R5249 gnd.n4957 gnd.n1715 585
R5250 gnd.n4107 gnd.n1715 585
R5251 gnd.n2400 gnd.n1713 585
R5252 gnd.n4078 gnd.n2400 585
R5253 gnd.n4961 gnd.n1712 585
R5254 gnd.n4099 gnd.n1712 585
R5255 gnd.n4962 gnd.n1711 585
R5256 gnd.n2392 gnd.n1711 585
R5257 gnd.n4963 gnd.n1710 585
R5258 gnd.n4091 gnd.n1710 585
R5259 gnd.n1707 gnd.n1705 585
R5260 gnd.n3464 gnd.n1705 585
R5261 gnd.n4968 gnd.n4967 585
R5262 gnd.t109 gnd.n4968 585
R5263 gnd.n1706 gnd.n1704 585
R5264 gnd.n3455 gnd.n1704 585
R5265 gnd.n2602 gnd.n1690 585
R5266 gnd.n4974 gnd.n1690 585
R5267 gnd.n2605 gnd.n2601 585
R5268 gnd.n2601 gnd.n1688 585
R5269 gnd.n2606 gnd.n2600 585
R5270 gnd.n2600 gnd.n1662 585
R5271 gnd.n2607 gnd.n2599 585
R5272 gnd.n2599 gnd.n1630 585
R5273 gnd.n2598 gnd.n2596 585
R5274 gnd.n2598 gnd.n2494 585
R5275 gnd.n2611 gnd.n2493 585
R5276 gnd.n3438 gnd.n2493 585
R5277 gnd.n2612 gnd.n2595 585
R5278 gnd.n2595 gnd.n2492 585
R5279 gnd.n2613 gnd.n2501 585
R5280 gnd.n3421 gnd.n2501 585
R5281 gnd.n2593 gnd.n2592 585
R5282 gnd.n2592 gnd.n2509 585
R5283 gnd.n2617 gnd.n2508 585
R5284 gnd.n3413 gnd.n2508 585
R5285 gnd.n2618 gnd.n2591 585
R5286 gnd.n2591 gnd.n2507 585
R5287 gnd.n2619 gnd.n2516 585
R5288 gnd.n3405 gnd.n2516 585
R5289 gnd.n2589 gnd.n2588 585
R5290 gnd.n2588 gnd.n2515 585
R5291 gnd.n2623 gnd.n2523 585
R5292 gnd.n3397 gnd.n2523 585
R5293 gnd.n2624 gnd.n2587 585
R5294 gnd.n2587 gnd.n2522 585
R5295 gnd.n2625 gnd.n2530 585
R5296 gnd.n3389 gnd.n2530 585
R5297 gnd.n2585 gnd.n2584 585
R5298 gnd.n2584 gnd.n2529 585
R5299 gnd.n2629 gnd.n2536 585
R5300 gnd.n3381 gnd.n2536 585
R5301 gnd.n2630 gnd.n2583 585
R5302 gnd.n2583 gnd.n2544 585
R5303 gnd.n2631 gnd.n2543 585
R5304 gnd.n3373 gnd.n2543 585
R5305 gnd.n3349 gnd.n3348 585
R5306 gnd.n3347 gnd.n2581 585
R5307 gnd.n2634 gnd.n2580 585
R5308 gnd.n3351 gnd.n2580 585
R5309 gnd.n3343 gnd.n2636 585
R5310 gnd.n3342 gnd.n2637 585
R5311 gnd.n3341 gnd.n2638 585
R5312 gnd.n3226 gnd.n2639 585
R5313 gnd.n3336 gnd.n3227 585
R5314 gnd.n3335 gnd.n3228 585
R5315 gnd.n3334 gnd.n3229 585
R5316 gnd.n3239 gnd.n3230 585
R5317 gnd.n3327 gnd.n3240 585
R5318 gnd.n3326 gnd.n3241 585
R5319 gnd.n3243 gnd.n3242 585
R5320 gnd.n3319 gnd.n3249 585
R5321 gnd.n3318 gnd.n3250 585
R5322 gnd.n3259 gnd.n3251 585
R5323 gnd.n3311 gnd.n3260 585
R5324 gnd.n3310 gnd.n3261 585
R5325 gnd.n3263 gnd.n3262 585
R5326 gnd.n3303 gnd.n3269 585
R5327 gnd.n3302 gnd.n3270 585
R5328 gnd.n3279 gnd.n3271 585
R5329 gnd.n3295 gnd.n3280 585
R5330 gnd.n3294 gnd.n3281 585
R5331 gnd.n3287 gnd.n3286 585
R5332 gnd.n2577 gnd.n2547 585
R5333 gnd.n3367 gnd.n2548 585
R5334 gnd.n3368 gnd.n2545 585
R5335 gnd.n4404 gnd.n1811 585
R5336 gnd.n4845 gnd.n1811 585
R5337 gnd.n4403 gnd.n4402 585
R5338 gnd.n4402 gnd.n1809 585
R5339 gnd.n4401 gnd.n2132 585
R5340 gnd.n4401 gnd.n4400 585
R5341 gnd.n2145 gnd.n2133 585
R5342 gnd.n2135 gnd.n2133 585
R5343 gnd.n4388 gnd.n4387 585
R5344 gnd.n4389 gnd.n4388 585
R5345 gnd.n2144 gnd.n2143 585
R5346 gnd.n2143 gnd.n2142 585
R5347 gnd.n4381 gnd.n4380 585
R5348 gnd.n4380 gnd.n4379 585
R5349 gnd.n2148 gnd.n2147 585
R5350 gnd.n2156 gnd.n2148 585
R5351 gnd.n4370 gnd.n4369 585
R5352 gnd.n4371 gnd.n4370 585
R5353 gnd.n2158 gnd.n2157 585
R5354 gnd.n2157 gnd.n2154 585
R5355 gnd.n4365 gnd.n4364 585
R5356 gnd.n4364 gnd.n4363 585
R5357 gnd.n2161 gnd.n2160 585
R5358 gnd.n2163 gnd.n2161 585
R5359 gnd.n4354 gnd.n4353 585
R5360 gnd.n4355 gnd.n4354 585
R5361 gnd.n2171 gnd.n2170 585
R5362 gnd.n2170 gnd.n2169 585
R5363 gnd.n4349 gnd.n4348 585
R5364 gnd.n4348 gnd.n4347 585
R5365 gnd.n2174 gnd.n2173 585
R5366 gnd.n2176 gnd.n2174 585
R5367 gnd.n4338 gnd.n4337 585
R5368 gnd.n4339 gnd.n4338 585
R5369 gnd.n2183 gnd.n2182 585
R5370 gnd.n3687 gnd.n2182 585
R5371 gnd.n4333 gnd.n4332 585
R5372 gnd.n4332 gnd.n4331 585
R5373 gnd.n2186 gnd.n2185 585
R5374 gnd.n3884 gnd.n2186 585
R5375 gnd.n4322 gnd.n4321 585
R5376 gnd.n4323 gnd.n4322 585
R5377 gnd.n2195 gnd.n2194 585
R5378 gnd.n3657 gnd.n2194 585
R5379 gnd.n4317 gnd.n4316 585
R5380 gnd.n4316 gnd.n4315 585
R5381 gnd.n2198 gnd.n2197 585
R5382 gnd.n3670 gnd.n2198 585
R5383 gnd.n4306 gnd.n4305 585
R5384 gnd.n4307 gnd.n4306 585
R5385 gnd.n2209 gnd.n2208 585
R5386 gnd.n2214 gnd.n2208 585
R5387 gnd.n4301 gnd.n4300 585
R5388 gnd.n4300 gnd.n4299 585
R5389 gnd.n2212 gnd.n2211 585
R5390 gnd.n3646 gnd.n2212 585
R5391 gnd.n4290 gnd.n4289 585
R5392 gnd.n4291 gnd.n4290 585
R5393 gnd.n2224 gnd.n2223 585
R5394 gnd.n3638 gnd.n2223 585
R5395 gnd.n4285 gnd.n4284 585
R5396 gnd.n4284 gnd.n4283 585
R5397 gnd.n2227 gnd.n2226 585
R5398 gnd.n3631 gnd.n2227 585
R5399 gnd.n4274 gnd.n4273 585
R5400 gnd.n4275 gnd.n4274 585
R5401 gnd.n2237 gnd.n2236 585
R5402 gnd.n3622 gnd.n2236 585
R5403 gnd.n4269 gnd.n4268 585
R5404 gnd.n4268 gnd.n4267 585
R5405 gnd.n2240 gnd.n2239 585
R5406 gnd.n3935 gnd.n2240 585
R5407 gnd.n4258 gnd.n4257 585
R5408 gnd.n4259 gnd.n4258 585
R5409 gnd.n2250 gnd.n2249 585
R5410 gnd.n3608 gnd.n2249 585
R5411 gnd.n4253 gnd.n4252 585
R5412 gnd.n4252 gnd.n4251 585
R5413 gnd.n2253 gnd.n2252 585
R5414 gnd.n3601 gnd.n2253 585
R5415 gnd.n4242 gnd.n4241 585
R5416 gnd.n4243 gnd.n4242 585
R5417 gnd.n2264 gnd.n2263 585
R5418 gnd.n3593 gnd.n2263 585
R5419 gnd.n4237 gnd.n4236 585
R5420 gnd.n4236 gnd.n4235 585
R5421 gnd.n2267 gnd.n2266 585
R5422 gnd.n3964 gnd.n2267 585
R5423 gnd.n4226 gnd.n4225 585
R5424 gnd.n4227 gnd.n4226 585
R5425 gnd.n2278 gnd.n2277 585
R5426 gnd.n3580 gnd.n2277 585
R5427 gnd.n4221 gnd.n4220 585
R5428 gnd.n4220 gnd.n4219 585
R5429 gnd.n2281 gnd.n2280 585
R5430 gnd.n3980 gnd.n2281 585
R5431 gnd.n4210 gnd.n4209 585
R5432 gnd.n4211 gnd.n4210 585
R5433 gnd.n2291 gnd.n2290 585
R5434 gnd.n3566 gnd.n2290 585
R5435 gnd.n4205 gnd.n4204 585
R5436 gnd.n4204 gnd.n4203 585
R5437 gnd.n2294 gnd.n2293 585
R5438 gnd.n3996 gnd.n2294 585
R5439 gnd.n4194 gnd.n4193 585
R5440 gnd.n4195 gnd.n4194 585
R5441 gnd.n2305 gnd.n2304 585
R5442 gnd.n3553 gnd.n2304 585
R5443 gnd.n4189 gnd.n4188 585
R5444 gnd.n4188 gnd.n4187 585
R5445 gnd.n2308 gnd.n2307 585
R5446 gnd.n4012 gnd.n2308 585
R5447 gnd.n4178 gnd.n4177 585
R5448 gnd.n4179 gnd.n4178 585
R5449 gnd.n2319 gnd.n2318 585
R5450 gnd.n3545 gnd.n2318 585
R5451 gnd.n4173 gnd.n4172 585
R5452 gnd.n4172 gnd.n4171 585
R5453 gnd.n2322 gnd.n2321 585
R5454 gnd.n2332 gnd.n2322 585
R5455 gnd.n4162 gnd.n4161 585
R5456 gnd.n4163 gnd.n4162 585
R5457 gnd.n2335 gnd.n2334 585
R5458 gnd.n3526 gnd.n2334 585
R5459 gnd.n4157 gnd.n4156 585
R5460 gnd.n4156 gnd.n4155 585
R5461 gnd.n2338 gnd.n2337 585
R5462 gnd.n3517 gnd.n2338 585
R5463 gnd.n4146 gnd.n4145 585
R5464 gnd.n4147 gnd.n4146 585
R5465 gnd.n2348 gnd.n2347 585
R5466 gnd.n3508 gnd.n2347 585
R5467 gnd.n4141 gnd.n4140 585
R5468 gnd.n4140 gnd.n4139 585
R5469 gnd.n2351 gnd.n2350 585
R5470 gnd.n4049 gnd.n2351 585
R5471 gnd.n4130 gnd.n4129 585
R5472 gnd.n4131 gnd.n4130 585
R5473 gnd.n2361 gnd.n2360 585
R5474 gnd.n3495 gnd.n2360 585
R5475 gnd.n4125 gnd.n4124 585
R5476 gnd.n4124 gnd.n4123 585
R5477 gnd.n2364 gnd.n2363 585
R5478 gnd.n3486 gnd.n2364 585
R5479 gnd.n4114 gnd.n4113 585
R5480 gnd.n4115 gnd.n4114 585
R5481 gnd.n2374 gnd.n2373 585
R5482 gnd.n3476 gnd.n2373 585
R5483 gnd.n4109 gnd.n4108 585
R5484 gnd.n4108 gnd.n4107 585
R5485 gnd.n2377 gnd.n2376 585
R5486 gnd.n4078 gnd.n2377 585
R5487 gnd.n4098 gnd.n4097 585
R5488 gnd.n4099 gnd.n4098 585
R5489 gnd.n2387 gnd.n2386 585
R5490 gnd.n2392 gnd.n2386 585
R5491 gnd.n4093 gnd.n4092 585
R5492 gnd.n4092 gnd.n4091 585
R5493 gnd.n2390 gnd.n2389 585
R5494 gnd.n3464 gnd.n2390 585
R5495 gnd.n2484 gnd.n1702 585
R5496 gnd.t109 gnd.n1702 585
R5497 gnd.n3454 gnd.n3453 585
R5498 gnd.n3455 gnd.n3454 585
R5499 gnd.n2483 gnd.n1692 585
R5500 gnd.n4974 gnd.n1692 585
R5501 gnd.n3448 gnd.n3447 585
R5502 gnd.n3447 gnd.n1688 585
R5503 gnd.n3446 gnd.n2486 585
R5504 gnd.n3446 gnd.n1662 585
R5505 gnd.n3445 gnd.n3444 585
R5506 gnd.n3445 gnd.n1630 585
R5507 gnd.n2488 gnd.n2487 585
R5508 gnd.n2494 gnd.n2487 585
R5509 gnd.n3440 gnd.n3439 585
R5510 gnd.n3439 gnd.n3438 585
R5511 gnd.n2491 gnd.n2490 585
R5512 gnd.n2492 gnd.n2491 585
R5513 gnd.n3420 gnd.n3419 585
R5514 gnd.n3421 gnd.n3420 585
R5515 gnd.n2503 gnd.n2502 585
R5516 gnd.n2509 gnd.n2502 585
R5517 gnd.n3415 gnd.n3414 585
R5518 gnd.n3414 gnd.n3413 585
R5519 gnd.n2506 gnd.n2505 585
R5520 gnd.n2507 gnd.n2506 585
R5521 gnd.n3404 gnd.n3403 585
R5522 gnd.n3405 gnd.n3404 585
R5523 gnd.n2518 gnd.n2517 585
R5524 gnd.n2517 gnd.n2515 585
R5525 gnd.n3399 gnd.n3398 585
R5526 gnd.n3398 gnd.n3397 585
R5527 gnd.n2521 gnd.n2520 585
R5528 gnd.n2522 gnd.n2521 585
R5529 gnd.n3388 gnd.n3387 585
R5530 gnd.n3389 gnd.n3388 585
R5531 gnd.n2532 gnd.n2531 585
R5532 gnd.n2531 gnd.n2529 585
R5533 gnd.n3383 gnd.n3382 585
R5534 gnd.n3382 gnd.n3381 585
R5535 gnd.n2535 gnd.n2534 585
R5536 gnd.n2544 gnd.n2535 585
R5537 gnd.n3372 gnd.n3371 585
R5538 gnd.n3373 gnd.n3372 585
R5539 gnd.n4546 gnd.n4409 585
R5540 gnd.n4409 gnd.n1812 585
R5541 gnd.n4545 gnd.n4544 585
R5542 gnd.n4542 gnd.n4421 585
R5543 gnd.n4541 gnd.n4540 585
R5544 gnd.n4525 gnd.n4423 585
R5545 gnd.n4527 gnd.n4526 585
R5546 gnd.n4523 gnd.n4429 585
R5547 gnd.n4522 gnd.n4521 585
R5548 gnd.n4506 gnd.n4431 585
R5549 gnd.n4508 gnd.n4507 585
R5550 gnd.n4504 gnd.n4436 585
R5551 gnd.n4503 gnd.n4502 585
R5552 gnd.n4487 gnd.n4438 585
R5553 gnd.n4489 gnd.n4488 585
R5554 gnd.n4485 gnd.n4443 585
R5555 gnd.n4484 gnd.n4483 585
R5556 gnd.n4470 gnd.n4445 585
R5557 gnd.n4472 gnd.n4471 585
R5558 gnd.n4468 gnd.n4446 585
R5559 gnd.n4467 gnd.n4466 585
R5560 gnd.n4459 gnd.n4448 585
R5561 gnd.n4461 gnd.n4460 585
R5562 gnd.n4457 gnd.n4450 585
R5563 gnd.n4456 gnd.n4455 585
R5564 gnd.n4452 gnd.n1808 585
R5565 gnd.n4563 gnd.n4562 585
R5566 gnd.n4564 gnd.n4560 585
R5567 gnd.n4559 gnd.n4408 585
R5568 gnd.n4557 gnd.n4556 585
R5569 gnd.n3729 gnd.n3728 468.476
R5570 gnd.n3878 gnd.n3680 468.476
R5571 gnd.n2474 gnd.n2472 468.476
R5572 gnd.n5043 gnd.n1665 468.476
R5573 gnd.n2408 gnd.t149 389.64
R5574 gnd.n3812 gnd.t114 389.64
R5575 gnd.n4980 gnd.t69 389.64
R5576 gnd.n3704 gnd.t161 389.64
R5577 gnd.n7052 gnd.n7051 374.827
R5578 gnd.n3282 gnd.t101 371.625
R5579 gnd.n4417 gnd.t61 371.625
R5580 gnd.n2550 gnd.t93 371.625
R5581 gnd.n1881 gnd.t155 371.625
R5582 gnd.n1904 gnd.t158 371.625
R5583 gnd.n1926 gnd.t121 371.625
R5584 gnd.n352 gnd.t82 371.625
R5585 gnd.n332 gnd.t90 371.625
R5586 gnd.n7968 gnd.t118 371.625
R5587 gnd.n372 gnd.t167 371.625
R5588 gnd.n1208 gnd.t111 371.625
R5589 gnd.n1230 gnd.t130 371.625
R5590 gnd.n1252 gnd.t152 371.625
R5591 gnd.n2901 gnd.t97 371.625
R5592 gnd.n1613 gnd.t124 371.625
R5593 gnd.n2641 gnd.t143 371.625
R5594 gnd.n2654 gnd.t174 371.625
R5595 gnd.n4410 gnd.t65 371.625
R5596 gnd.n6388 gnd.t86 323.425
R5597 gnd.n5430 gnd.t139 323.425
R5598 gnd.n5741 gnd.n5715 289.615
R5599 gnd.n5709 gnd.n5683 289.615
R5600 gnd.n5677 gnd.n5651 289.615
R5601 gnd.n5646 gnd.n5620 289.615
R5602 gnd.n5614 gnd.n5588 289.615
R5603 gnd.n5582 gnd.n5556 289.615
R5604 gnd.n5550 gnd.n5524 289.615
R5605 gnd.n5519 gnd.n5493 289.615
R5606 gnd.n6093 gnd.t57 279.217
R5607 gnd.n5474 gnd.t170 279.217
R5608 gnd.n1672 gnd.t78 260.649
R5609 gnd.n3717 gnd.t129 260.649
R5610 gnd.n5045 gnd.n5044 256.663
R5611 gnd.n5045 gnd.n1631 256.663
R5612 gnd.n5045 gnd.n1632 256.663
R5613 gnd.n5045 gnd.n1633 256.663
R5614 gnd.n5045 gnd.n1634 256.663
R5615 gnd.n5045 gnd.n1635 256.663
R5616 gnd.n5045 gnd.n1636 256.663
R5617 gnd.n5045 gnd.n1637 256.663
R5618 gnd.n5045 gnd.n1638 256.663
R5619 gnd.n5045 gnd.n1639 256.663
R5620 gnd.n5045 gnd.n1640 256.663
R5621 gnd.n5045 gnd.n1641 256.663
R5622 gnd.n5045 gnd.n1642 256.663
R5623 gnd.n5045 gnd.n1643 256.663
R5624 gnd.n5045 gnd.n1644 256.663
R5625 gnd.n5045 gnd.n1645 256.663
R5626 gnd.n5048 gnd.n1628 256.663
R5627 gnd.n5046 gnd.n5045 256.663
R5628 gnd.n5045 gnd.n1646 256.663
R5629 gnd.n5045 gnd.n1647 256.663
R5630 gnd.n5045 gnd.n1648 256.663
R5631 gnd.n5045 gnd.n1649 256.663
R5632 gnd.n5045 gnd.n1650 256.663
R5633 gnd.n5045 gnd.n1651 256.663
R5634 gnd.n5045 gnd.n1652 256.663
R5635 gnd.n5045 gnd.n1653 256.663
R5636 gnd.n5045 gnd.n1654 256.663
R5637 gnd.n5045 gnd.n1655 256.663
R5638 gnd.n5045 gnd.n1656 256.663
R5639 gnd.n5045 gnd.n1657 256.663
R5640 gnd.n5045 gnd.n1658 256.663
R5641 gnd.n5045 gnd.n1659 256.663
R5642 gnd.n5045 gnd.n1660 256.663
R5643 gnd.n5045 gnd.n1661 256.663
R5644 gnd.n3877 gnd.n3876 256.663
R5645 gnd.n3876 gnd.n3796 256.663
R5646 gnd.n3876 gnd.n3797 256.663
R5647 gnd.n3876 gnd.n3798 256.663
R5648 gnd.n3876 gnd.n3799 256.663
R5649 gnd.n3876 gnd.n3800 256.663
R5650 gnd.n3876 gnd.n3801 256.663
R5651 gnd.n3876 gnd.n3802 256.663
R5652 gnd.n3876 gnd.n3803 256.663
R5653 gnd.n3876 gnd.n3804 256.663
R5654 gnd.n3876 gnd.n3805 256.663
R5655 gnd.n3876 gnd.n3806 256.663
R5656 gnd.n3876 gnd.n3807 256.663
R5657 gnd.n3876 gnd.n3808 256.663
R5658 gnd.n3876 gnd.n3809 256.663
R5659 gnd.n3876 gnd.n3810 256.663
R5660 gnd.n3811 gnd.n1891 256.663
R5661 gnd.n3876 gnd.n3795 256.663
R5662 gnd.n3876 gnd.n3703 256.663
R5663 gnd.n3876 gnd.n3702 256.663
R5664 gnd.n3876 gnd.n3701 256.663
R5665 gnd.n3876 gnd.n3700 256.663
R5666 gnd.n3876 gnd.n3699 256.663
R5667 gnd.n3876 gnd.n3698 256.663
R5668 gnd.n3876 gnd.n3697 256.663
R5669 gnd.n3876 gnd.n3696 256.663
R5670 gnd.n3876 gnd.n3695 256.663
R5671 gnd.n3876 gnd.n3694 256.663
R5672 gnd.n3876 gnd.n3693 256.663
R5673 gnd.n3876 gnd.n3692 256.663
R5674 gnd.n3876 gnd.n3691 256.663
R5675 gnd.n3876 gnd.n3690 256.663
R5676 gnd.n3876 gnd.n3689 256.663
R5677 gnd.n3876 gnd.n3688 256.663
R5678 gnd.n5400 gnd.n1176 242.672
R5679 gnd.n5400 gnd.n1177 242.672
R5680 gnd.n5400 gnd.n1178 242.672
R5681 gnd.n5400 gnd.n1179 242.672
R5682 gnd.n5400 gnd.n1180 242.672
R5683 gnd.n5400 gnd.n1181 242.672
R5684 gnd.n5400 gnd.n1182 242.672
R5685 gnd.n5400 gnd.n1183 242.672
R5686 gnd.n5400 gnd.n1184 242.672
R5687 gnd.n5099 gnd.n1566 242.672
R5688 gnd.n5099 gnd.n1565 242.672
R5689 gnd.n5099 gnd.n1564 242.672
R5690 gnd.n5099 gnd.n1563 242.672
R5691 gnd.n5099 gnd.n1562 242.672
R5692 gnd.n5099 gnd.n1561 242.672
R5693 gnd.n5099 gnd.n1560 242.672
R5694 gnd.n5099 gnd.n1559 242.672
R5695 gnd.n5099 gnd.n1558 242.672
R5696 gnd.n6148 gnd.n6057 242.672
R5697 gnd.n6061 gnd.n6057 242.672
R5698 gnd.n6141 gnd.n6057 242.672
R5699 gnd.n6135 gnd.n6057 242.672
R5700 gnd.n6133 gnd.n6057 242.672
R5701 gnd.n6127 gnd.n6057 242.672
R5702 gnd.n6125 gnd.n6057 242.672
R5703 gnd.n6119 gnd.n6057 242.672
R5704 gnd.n6117 gnd.n6057 242.672
R5705 gnd.n6111 gnd.n6057 242.672
R5706 gnd.n6109 gnd.n6057 242.672
R5707 gnd.n6102 gnd.n6057 242.672
R5708 gnd.n6100 gnd.n6057 242.672
R5709 gnd.n6792 gnd.n5401 242.672
R5710 gnd.n6798 gnd.n5401 242.672
R5711 gnd.n5477 gnd.n5401 242.672
R5712 gnd.n6805 gnd.n5401 242.672
R5713 gnd.n5468 gnd.n5401 242.672
R5714 gnd.n6812 gnd.n5401 242.672
R5715 gnd.n5461 gnd.n5401 242.672
R5716 gnd.n6819 gnd.n5401 242.672
R5717 gnd.n5454 gnd.n5401 242.672
R5718 gnd.n6826 gnd.n5401 242.672
R5719 gnd.n5447 gnd.n5401 242.672
R5720 gnd.n6833 gnd.n5401 242.672
R5721 gnd.n5440 gnd.n5401 242.672
R5722 gnd.n4836 gnd.n1849 242.672
R5723 gnd.n4836 gnd.n1850 242.672
R5724 gnd.n4836 gnd.n1851 242.672
R5725 gnd.n4836 gnd.n1852 242.672
R5726 gnd.n4836 gnd.n1853 242.672
R5727 gnd.n4836 gnd.n1854 242.672
R5728 gnd.n4836 gnd.n1855 242.672
R5729 gnd.n4836 gnd.n1856 242.672
R5730 gnd.n4836 gnd.n1857 242.672
R5731 gnd.n8003 gnd.n266 242.672
R5732 gnd.n8003 gnd.n265 242.672
R5733 gnd.n8003 gnd.n264 242.672
R5734 gnd.n8003 gnd.n263 242.672
R5735 gnd.n8003 gnd.n262 242.672
R5736 gnd.n8003 gnd.n261 242.672
R5737 gnd.n8003 gnd.n260 242.672
R5738 gnd.n8003 gnd.n259 242.672
R5739 gnd.n8003 gnd.n258 242.672
R5740 gnd.n6422 gnd.n6421 242.672
R5741 gnd.n6422 gnd.n6363 242.672
R5742 gnd.n6422 gnd.n6364 242.672
R5743 gnd.n6422 gnd.n6365 242.672
R5744 gnd.n6422 gnd.n6366 242.672
R5745 gnd.n6422 gnd.n6367 242.672
R5746 gnd.n6422 gnd.n6368 242.672
R5747 gnd.n6422 gnd.n6369 242.672
R5748 gnd.n6844 gnd.n5401 242.672
R5749 gnd.n5433 gnd.n5401 242.672
R5750 gnd.n6851 gnd.n5401 242.672
R5751 gnd.n5424 gnd.n5401 242.672
R5752 gnd.n6858 gnd.n5401 242.672
R5753 gnd.n5417 gnd.n5401 242.672
R5754 gnd.n6865 gnd.n5401 242.672
R5755 gnd.n5410 gnd.n5401 242.672
R5756 gnd.n5400 gnd.n5399 242.672
R5757 gnd.n5400 gnd.n1148 242.672
R5758 gnd.n5400 gnd.n1149 242.672
R5759 gnd.n5400 gnd.n1150 242.672
R5760 gnd.n5400 gnd.n1151 242.672
R5761 gnd.n5400 gnd.n1152 242.672
R5762 gnd.n5400 gnd.n1153 242.672
R5763 gnd.n5400 gnd.n1154 242.672
R5764 gnd.n5400 gnd.n1155 242.672
R5765 gnd.n5400 gnd.n1156 242.672
R5766 gnd.n5400 gnd.n1157 242.672
R5767 gnd.n5400 gnd.n1158 242.672
R5768 gnd.n5400 gnd.n1159 242.672
R5769 gnd.n5400 gnd.n1160 242.672
R5770 gnd.n5400 gnd.n1161 242.672
R5771 gnd.n5400 gnd.n1162 242.672
R5772 gnd.n5400 gnd.n1163 242.672
R5773 gnd.n5400 gnd.n1164 242.672
R5774 gnd.n5400 gnd.n1165 242.672
R5775 gnd.n5400 gnd.n1166 242.672
R5776 gnd.n5400 gnd.n1167 242.672
R5777 gnd.n5400 gnd.n1168 242.672
R5778 gnd.n5400 gnd.n1169 242.672
R5779 gnd.n5400 gnd.n1170 242.672
R5780 gnd.n5400 gnd.n1171 242.672
R5781 gnd.n5400 gnd.n1172 242.672
R5782 gnd.n5400 gnd.n1173 242.672
R5783 gnd.n5400 gnd.n1174 242.672
R5784 gnd.n5400 gnd.n1175 242.672
R5785 gnd.n5099 gnd.n1568 242.672
R5786 gnd.n5099 gnd.n1569 242.672
R5787 gnd.n5099 gnd.n1570 242.672
R5788 gnd.n5099 gnd.n1571 242.672
R5789 gnd.n5099 gnd.n1572 242.672
R5790 gnd.n5099 gnd.n1573 242.672
R5791 gnd.n5099 gnd.n1574 242.672
R5792 gnd.n5099 gnd.n1575 242.672
R5793 gnd.n5099 gnd.n1576 242.672
R5794 gnd.n5099 gnd.n1577 242.672
R5795 gnd.n5099 gnd.n1578 242.672
R5796 gnd.n5099 gnd.n1579 242.672
R5797 gnd.n5099 gnd.n1580 242.672
R5798 gnd.n5099 gnd.n1581 242.672
R5799 gnd.n5099 gnd.n1582 242.672
R5800 gnd.n5099 gnd.n1583 242.672
R5801 gnd.n5049 gnd.n1624 242.672
R5802 gnd.n5099 gnd.n1584 242.672
R5803 gnd.n5099 gnd.n1585 242.672
R5804 gnd.n5099 gnd.n1586 242.672
R5805 gnd.n5099 gnd.n1587 242.672
R5806 gnd.n5099 gnd.n1588 242.672
R5807 gnd.n5099 gnd.n1589 242.672
R5808 gnd.n5099 gnd.n1590 242.672
R5809 gnd.n5099 gnd.n1591 242.672
R5810 gnd.n5099 gnd.n1592 242.672
R5811 gnd.n5099 gnd.n1593 242.672
R5812 gnd.n5099 gnd.n1594 242.672
R5813 gnd.n5099 gnd.n1595 242.672
R5814 gnd.n5099 gnd.n5098 242.672
R5815 gnd.n4836 gnd.n4835 242.672
R5816 gnd.n4836 gnd.n1821 242.672
R5817 gnd.n4836 gnd.n1822 242.672
R5818 gnd.n4836 gnd.n1823 242.672
R5819 gnd.n4836 gnd.n1824 242.672
R5820 gnd.n4836 gnd.n1825 242.672
R5821 gnd.n4836 gnd.n1826 242.672
R5822 gnd.n4836 gnd.n1827 242.672
R5823 gnd.n4836 gnd.n1828 242.672
R5824 gnd.n4836 gnd.n1829 242.672
R5825 gnd.n4836 gnd.n1830 242.672
R5826 gnd.n4836 gnd.n1831 242.672
R5827 gnd.n4836 gnd.n1832 242.672
R5828 gnd.n4783 gnd.n1892 242.672
R5829 gnd.n4836 gnd.n1833 242.672
R5830 gnd.n4836 gnd.n1834 242.672
R5831 gnd.n4836 gnd.n1835 242.672
R5832 gnd.n4836 gnd.n1836 242.672
R5833 gnd.n4836 gnd.n1837 242.672
R5834 gnd.n4836 gnd.n1838 242.672
R5835 gnd.n4836 gnd.n1839 242.672
R5836 gnd.n4836 gnd.n1840 242.672
R5837 gnd.n4836 gnd.n1841 242.672
R5838 gnd.n4836 gnd.n1842 242.672
R5839 gnd.n4836 gnd.n1843 242.672
R5840 gnd.n4836 gnd.n1844 242.672
R5841 gnd.n4836 gnd.n1845 242.672
R5842 gnd.n4836 gnd.n1846 242.672
R5843 gnd.n4836 gnd.n1847 242.672
R5844 gnd.n4836 gnd.n1848 242.672
R5845 gnd.n8003 gnd.n267 242.672
R5846 gnd.n8003 gnd.n268 242.672
R5847 gnd.n8003 gnd.n269 242.672
R5848 gnd.n8003 gnd.n270 242.672
R5849 gnd.n8003 gnd.n271 242.672
R5850 gnd.n8003 gnd.n272 242.672
R5851 gnd.n8003 gnd.n273 242.672
R5852 gnd.n8003 gnd.n274 242.672
R5853 gnd.n8003 gnd.n275 242.672
R5854 gnd.n8003 gnd.n276 242.672
R5855 gnd.n8003 gnd.n277 242.672
R5856 gnd.n8003 gnd.n278 242.672
R5857 gnd.n8003 gnd.n279 242.672
R5858 gnd.n8003 gnd.n280 242.672
R5859 gnd.n8003 gnd.n281 242.672
R5860 gnd.n8003 gnd.n282 242.672
R5861 gnd.n8003 gnd.n283 242.672
R5862 gnd.n8003 gnd.n284 242.672
R5863 gnd.n8003 gnd.n285 242.672
R5864 gnd.n8003 gnd.n286 242.672
R5865 gnd.n8003 gnd.n287 242.672
R5866 gnd.n8003 gnd.n288 242.672
R5867 gnd.n8003 gnd.n289 242.672
R5868 gnd.n8003 gnd.n290 242.672
R5869 gnd.n8003 gnd.n291 242.672
R5870 gnd.n8003 gnd.n292 242.672
R5871 gnd.n8003 gnd.n293 242.672
R5872 gnd.n8003 gnd.n294 242.672
R5873 gnd.n8003 gnd.n8002 242.672
R5874 gnd.n3351 gnd.n3350 242.672
R5875 gnd.n3351 gnd.n2566 242.672
R5876 gnd.n3351 gnd.n2567 242.672
R5877 gnd.n3351 gnd.n2568 242.672
R5878 gnd.n3351 gnd.n2569 242.672
R5879 gnd.n3351 gnd.n2570 242.672
R5880 gnd.n3351 gnd.n2571 242.672
R5881 gnd.n3351 gnd.n2572 242.672
R5882 gnd.n3351 gnd.n2573 242.672
R5883 gnd.n3351 gnd.n2574 242.672
R5884 gnd.n3351 gnd.n2575 242.672
R5885 gnd.n3351 gnd.n2576 242.672
R5886 gnd.n3351 gnd.n2578 242.672
R5887 gnd.n3351 gnd.n2579 242.672
R5888 gnd.n4543 gnd.n1812 242.672
R5889 gnd.n4422 gnd.n1812 242.672
R5890 gnd.n4524 gnd.n1812 242.672
R5891 gnd.n4430 gnd.n1812 242.672
R5892 gnd.n4505 gnd.n1812 242.672
R5893 gnd.n4437 gnd.n1812 242.672
R5894 gnd.n4486 gnd.n1812 242.672
R5895 gnd.n4444 gnd.n1812 242.672
R5896 gnd.n4469 gnd.n1812 242.672
R5897 gnd.n4447 gnd.n1812 242.672
R5898 gnd.n4458 gnd.n1812 242.672
R5899 gnd.n4451 gnd.n1812 242.672
R5900 gnd.n4561 gnd.n1812 242.672
R5901 gnd.n4558 gnd.n1812 242.672
R5902 gnd.n8004 gnd.n256 240.244
R5903 gnd.n8001 gnd.n295 240.244
R5904 gnd.n7997 gnd.n7996 240.244
R5905 gnd.n7993 gnd.n7992 240.244
R5906 gnd.n7989 gnd.n7988 240.244
R5907 gnd.n7985 gnd.n7984 240.244
R5908 gnd.n7981 gnd.n7980 240.244
R5909 gnd.n7977 gnd.n7976 240.244
R5910 gnd.n7973 gnd.n7972 240.244
R5911 gnd.n7966 gnd.n7965 240.244
R5912 gnd.n7962 gnd.n7961 240.244
R5913 gnd.n7958 gnd.n7957 240.244
R5914 gnd.n7954 gnd.n7953 240.244
R5915 gnd.n7950 gnd.n7949 240.244
R5916 gnd.n7946 gnd.n7945 240.244
R5917 gnd.n7942 gnd.n7941 240.244
R5918 gnd.n7938 gnd.n7937 240.244
R5919 gnd.n7934 gnd.n7933 240.244
R5920 gnd.n7930 gnd.n7929 240.244
R5921 gnd.n7923 gnd.n7922 240.244
R5922 gnd.n7920 gnd.n7919 240.244
R5923 gnd.n7916 gnd.n7915 240.244
R5924 gnd.n7912 gnd.n7911 240.244
R5925 gnd.n7908 gnd.n7907 240.244
R5926 gnd.n7904 gnd.n7903 240.244
R5927 gnd.n7900 gnd.n7899 240.244
R5928 gnd.n7896 gnd.n7895 240.244
R5929 gnd.n7892 gnd.n7891 240.244
R5930 gnd.n7888 gnd.n7887 240.244
R5931 gnd.n4717 gnd.n1933 240.244
R5932 gnd.n4574 gnd.n1933 240.244
R5933 gnd.n4574 gnd.n1951 240.244
R5934 gnd.n4578 gnd.n1951 240.244
R5935 gnd.n4578 gnd.n1962 240.244
R5936 gnd.n4588 gnd.n1962 240.244
R5937 gnd.n4588 gnd.n1973 240.244
R5938 gnd.n4592 gnd.n1973 240.244
R5939 gnd.n4592 gnd.n1983 240.244
R5940 gnd.n4602 gnd.n1983 240.244
R5941 gnd.n4602 gnd.n1993 240.244
R5942 gnd.n4606 gnd.n1993 240.244
R5943 gnd.n4606 gnd.n2003 240.244
R5944 gnd.n4616 gnd.n2003 240.244
R5945 gnd.n4616 gnd.n2014 240.244
R5946 gnd.n4623 gnd.n2014 240.244
R5947 gnd.n4623 gnd.n2024 240.244
R5948 gnd.n2051 gnd.n2024 240.244
R5949 gnd.n2051 gnd.n2035 240.244
R5950 gnd.n4653 gnd.n2035 240.244
R5951 gnd.n4653 gnd.n2043 240.244
R5952 gnd.n2043 gnd.n543 240.244
R5953 gnd.n7745 gnd.n543 240.244
R5954 gnd.n7745 gnd.n533 240.244
R5955 gnd.n533 gnd.n525 240.244
R5956 gnd.n7777 gnd.n525 240.244
R5957 gnd.n7777 gnd.n516 240.244
R5958 gnd.n516 gnd.n511 240.244
R5959 gnd.n7783 gnd.n511 240.244
R5960 gnd.n7783 gnd.n503 240.244
R5961 gnd.n503 gnd.n498 240.244
R5962 gnd.n498 gnd.n492 240.244
R5963 gnd.n7821 gnd.n492 240.244
R5964 gnd.n7821 gnd.n106 240.244
R5965 gnd.n7830 gnd.n106 240.244
R5966 gnd.n7831 gnd.n7830 240.244
R5967 gnd.n7831 gnd.n123 240.244
R5968 gnd.n7834 gnd.n123 240.244
R5969 gnd.n7834 gnd.n134 240.244
R5970 gnd.n7838 gnd.n134 240.244
R5971 gnd.n7838 gnd.n143 240.244
R5972 gnd.n7841 gnd.n143 240.244
R5973 gnd.n7841 gnd.n152 240.244
R5974 gnd.n7845 gnd.n152 240.244
R5975 gnd.n7845 gnd.n162 240.244
R5976 gnd.n7848 gnd.n162 240.244
R5977 gnd.n7848 gnd.n171 240.244
R5978 gnd.n7852 gnd.n171 240.244
R5979 gnd.n7852 gnd.n181 240.244
R5980 gnd.n7855 gnd.n181 240.244
R5981 gnd.n7855 gnd.n190 240.244
R5982 gnd.n7859 gnd.n190 240.244
R5983 gnd.n7859 gnd.n200 240.244
R5984 gnd.n7862 gnd.n200 240.244
R5985 gnd.n7862 gnd.n209 240.244
R5986 gnd.n7866 gnd.n209 240.244
R5987 gnd.n7866 gnd.n220 240.244
R5988 gnd.n7869 gnd.n220 240.244
R5989 gnd.n7869 gnd.n229 240.244
R5990 gnd.n7873 gnd.n229 240.244
R5991 gnd.n7873 gnd.n239 240.244
R5992 gnd.n7876 gnd.n239 240.244
R5993 gnd.n7876 gnd.n248 240.244
R5994 gnd.n7880 gnd.n248 240.244
R5995 gnd.n1861 gnd.n1860 240.244
R5996 gnd.n4829 gnd.n1860 240.244
R5997 gnd.n4827 gnd.n4826 240.244
R5998 gnd.n4823 gnd.n4822 240.244
R5999 gnd.n4819 gnd.n4818 240.244
R6000 gnd.n4815 gnd.n4814 240.244
R6001 gnd.n4811 gnd.n4810 240.244
R6002 gnd.n4807 gnd.n4806 240.244
R6003 gnd.n4803 gnd.n4802 240.244
R6004 gnd.n4798 gnd.n4797 240.244
R6005 gnd.n4794 gnd.n4793 240.244
R6006 gnd.n4790 gnd.n4789 240.244
R6007 gnd.n4786 gnd.n4785 240.244
R6008 gnd.n4781 gnd.n4780 240.244
R6009 gnd.n4777 gnd.n4776 240.244
R6010 gnd.n4773 gnd.n4772 240.244
R6011 gnd.n4769 gnd.n4768 240.244
R6012 gnd.n4765 gnd.n4764 240.244
R6013 gnd.n4761 gnd.n4760 240.244
R6014 gnd.n4757 gnd.n4756 240.244
R6015 gnd.n4753 gnd.n4752 240.244
R6016 gnd.n4749 gnd.n4748 240.244
R6017 gnd.n4745 gnd.n4744 240.244
R6018 gnd.n4741 gnd.n4740 240.244
R6019 gnd.n4737 gnd.n4736 240.244
R6020 gnd.n4733 gnd.n4732 240.244
R6021 gnd.n4729 gnd.n4728 240.244
R6022 gnd.n4725 gnd.n4724 240.244
R6023 gnd.n4712 gnd.n1862 240.244
R6024 gnd.n4712 gnd.n1942 240.244
R6025 gnd.n4708 gnd.n1942 240.244
R6026 gnd.n4708 gnd.n1949 240.244
R6027 gnd.n4700 gnd.n1949 240.244
R6028 gnd.n4700 gnd.n1965 240.244
R6029 gnd.n4696 gnd.n1965 240.244
R6030 gnd.n4696 gnd.n1971 240.244
R6031 gnd.n4688 gnd.n1971 240.244
R6032 gnd.n4688 gnd.n1985 240.244
R6033 gnd.n4684 gnd.n1985 240.244
R6034 gnd.n4684 gnd.n1991 240.244
R6035 gnd.n4676 gnd.n1991 240.244
R6036 gnd.n4676 gnd.n2006 240.244
R6037 gnd.n4672 gnd.n2006 240.244
R6038 gnd.n4672 gnd.n2012 240.244
R6039 gnd.n4664 gnd.n2012 240.244
R6040 gnd.n4664 gnd.n2026 240.244
R6041 gnd.n4660 gnd.n2026 240.244
R6042 gnd.n4660 gnd.n2033 240.244
R6043 gnd.n2033 gnd.n541 240.244
R6044 gnd.n7758 gnd.n541 240.244
R6045 gnd.n7758 gnd.n536 240.244
R6046 gnd.n7767 gnd.n536 240.244
R6047 gnd.n7767 gnd.n537 240.244
R6048 gnd.n537 gnd.n513 240.244
R6049 gnd.n7791 gnd.n513 240.244
R6050 gnd.n7794 gnd.n7791 240.244
R6051 gnd.n7794 gnd.n501 240.244
R6052 gnd.n7804 gnd.n501 240.244
R6053 gnd.n7812 gnd.n7804 240.244
R6054 gnd.n7812 gnd.n7809 240.244
R6055 gnd.n7809 gnd.n109 240.244
R6056 gnd.n8096 gnd.n109 240.244
R6057 gnd.n8096 gnd.n110 240.244
R6058 gnd.n120 gnd.n110 240.244
R6059 gnd.n8090 gnd.n120 240.244
R6060 gnd.n8090 gnd.n121 240.244
R6061 gnd.n8082 gnd.n121 240.244
R6062 gnd.n8082 gnd.n137 240.244
R6063 gnd.n8078 gnd.n137 240.244
R6064 gnd.n8078 gnd.n142 240.244
R6065 gnd.n8070 gnd.n142 240.244
R6066 gnd.n8070 gnd.n154 240.244
R6067 gnd.n8066 gnd.n154 240.244
R6068 gnd.n8066 gnd.n160 240.244
R6069 gnd.n8058 gnd.n160 240.244
R6070 gnd.n8058 gnd.n174 240.244
R6071 gnd.n8054 gnd.n174 240.244
R6072 gnd.n8054 gnd.n180 240.244
R6073 gnd.n8046 gnd.n180 240.244
R6074 gnd.n8046 gnd.n192 240.244
R6075 gnd.n8042 gnd.n192 240.244
R6076 gnd.n8042 gnd.n198 240.244
R6077 gnd.n8034 gnd.n198 240.244
R6078 gnd.n8034 gnd.n212 240.244
R6079 gnd.n8030 gnd.n212 240.244
R6080 gnd.n8030 gnd.n218 240.244
R6081 gnd.n8022 gnd.n218 240.244
R6082 gnd.n8022 gnd.n232 240.244
R6083 gnd.n8018 gnd.n232 240.244
R6084 gnd.n8018 gnd.n238 240.244
R6085 gnd.n8010 gnd.n238 240.244
R6086 gnd.n8010 gnd.n251 240.244
R6087 gnd.n5100 gnd.n1555 240.244
R6088 gnd.n5097 gnd.n1596 240.244
R6089 gnd.n5093 gnd.n5092 240.244
R6090 gnd.n5089 gnd.n5088 240.244
R6091 gnd.n5085 gnd.n5084 240.244
R6092 gnd.n5081 gnd.n5080 240.244
R6093 gnd.n5077 gnd.n5076 240.244
R6094 gnd.n5073 gnd.n5072 240.244
R6095 gnd.n5069 gnd.n5068 240.244
R6096 gnd.n5064 gnd.n5063 240.244
R6097 gnd.n5060 gnd.n5059 240.244
R6098 gnd.n5056 gnd.n5055 240.244
R6099 gnd.n5052 gnd.n5051 240.244
R6100 gnd.n2663 gnd.n2662 240.244
R6101 gnd.n2666 gnd.n2665 240.244
R6102 gnd.n2673 gnd.n2672 240.244
R6103 gnd.n2676 gnd.n2675 240.244
R6104 gnd.n2681 gnd.n2656 240.244
R6105 gnd.n2685 gnd.n2684 240.244
R6106 gnd.n2692 gnd.n2691 240.244
R6107 gnd.n2695 gnd.n2694 240.244
R6108 gnd.n2702 gnd.n2701 240.244
R6109 gnd.n2705 gnd.n2704 240.244
R6110 gnd.n2712 gnd.n2711 240.244
R6111 gnd.n2715 gnd.n2714 240.244
R6112 gnd.n2722 gnd.n2721 240.244
R6113 gnd.n2725 gnd.n2724 240.244
R6114 gnd.n2730 gnd.n2643 240.244
R6115 gnd.n5278 gnd.n5277 240.244
R6116 gnd.n5277 gnd.n1259 240.244
R6117 gnd.n1271 gnd.n1259 240.244
R6118 gnd.n2828 gnd.n1271 240.244
R6119 gnd.n2828 gnd.n1283 240.244
R6120 gnd.n2832 gnd.n1283 240.244
R6121 gnd.n2832 gnd.n1293 240.244
R6122 gnd.n2835 gnd.n1293 240.244
R6123 gnd.n2835 gnd.n1302 240.244
R6124 gnd.n2839 gnd.n1302 240.244
R6125 gnd.n2839 gnd.n1312 240.244
R6126 gnd.n2842 gnd.n1312 240.244
R6127 gnd.n2842 gnd.n1321 240.244
R6128 gnd.n2846 gnd.n1321 240.244
R6129 gnd.n2846 gnd.n1331 240.244
R6130 gnd.n2849 gnd.n1331 240.244
R6131 gnd.n2849 gnd.n1340 240.244
R6132 gnd.n2853 gnd.n1340 240.244
R6133 gnd.n2853 gnd.n1350 240.244
R6134 gnd.n2856 gnd.n1350 240.244
R6135 gnd.n2856 gnd.n1359 240.244
R6136 gnd.n2860 gnd.n1359 240.244
R6137 gnd.n2860 gnd.n1369 240.244
R6138 gnd.n2863 gnd.n1369 240.244
R6139 gnd.n2863 gnd.n1378 240.244
R6140 gnd.n2867 gnd.n1378 240.244
R6141 gnd.n2867 gnd.n1387 240.244
R6142 gnd.n2870 gnd.n1387 240.244
R6143 gnd.n2870 gnd.n1397 240.244
R6144 gnd.n2873 gnd.n1397 240.244
R6145 gnd.n2873 gnd.n2807 240.244
R6146 gnd.n3025 gnd.n2807 240.244
R6147 gnd.n3025 gnd.n2798 240.244
R6148 gnd.n2798 gnd.n2791 240.244
R6149 gnd.n3032 gnd.n2791 240.244
R6150 gnd.n3032 gnd.n2785 240.244
R6151 gnd.n2785 gnd.n1413 240.244
R6152 gnd.n2777 gnd.n1413 240.244
R6153 gnd.n2777 gnd.n1424 240.244
R6154 gnd.n3094 gnd.n1424 240.244
R6155 gnd.n3094 gnd.n1434 240.244
R6156 gnd.n3098 gnd.n1434 240.244
R6157 gnd.n3098 gnd.n1444 240.244
R6158 gnd.n3108 gnd.n1444 240.244
R6159 gnd.n3108 gnd.n1455 240.244
R6160 gnd.n2758 gnd.n1455 240.244
R6161 gnd.n2758 gnd.n1464 240.244
R6162 gnd.n3115 gnd.n1464 240.244
R6163 gnd.n3115 gnd.n1475 240.244
R6164 gnd.n3119 gnd.n1475 240.244
R6165 gnd.n3119 gnd.n1485 240.244
R6166 gnd.n3124 gnd.n1485 240.244
R6167 gnd.n3124 gnd.n1496 240.244
R6168 gnd.n3187 gnd.n1496 240.244
R6169 gnd.n3187 gnd.n1505 240.244
R6170 gnd.n3192 gnd.n1505 240.244
R6171 gnd.n3192 gnd.n1516 240.244
R6172 gnd.n3202 gnd.n1516 240.244
R6173 gnd.n3202 gnd.n1526 240.244
R6174 gnd.n3207 gnd.n1526 240.244
R6175 gnd.n3207 gnd.n1537 240.244
R6176 gnd.n3219 gnd.n1537 240.244
R6177 gnd.n3219 gnd.n1547 240.244
R6178 gnd.n2554 gnd.n1547 240.244
R6179 gnd.n1188 gnd.n1187 240.244
R6180 gnd.n5393 gnd.n1187 240.244
R6181 gnd.n5391 gnd.n5390 240.244
R6182 gnd.n5387 gnd.n5386 240.244
R6183 gnd.n5383 gnd.n5382 240.244
R6184 gnd.n5379 gnd.n5378 240.244
R6185 gnd.n5375 gnd.n5374 240.244
R6186 gnd.n5371 gnd.n5370 240.244
R6187 gnd.n5367 gnd.n5366 240.244
R6188 gnd.n5362 gnd.n5361 240.244
R6189 gnd.n5358 gnd.n5357 240.244
R6190 gnd.n5354 gnd.n5353 240.244
R6191 gnd.n5350 gnd.n5349 240.244
R6192 gnd.n5346 gnd.n5345 240.244
R6193 gnd.n5342 gnd.n5341 240.244
R6194 gnd.n5338 gnd.n5337 240.244
R6195 gnd.n5334 gnd.n5333 240.244
R6196 gnd.n5330 gnd.n5329 240.244
R6197 gnd.n5326 gnd.n5325 240.244
R6198 gnd.n5322 gnd.n5321 240.244
R6199 gnd.n5318 gnd.n5317 240.244
R6200 gnd.n5314 gnd.n5313 240.244
R6201 gnd.n5310 gnd.n5309 240.244
R6202 gnd.n5306 gnd.n5305 240.244
R6203 gnd.n5302 gnd.n5301 240.244
R6204 gnd.n5298 gnd.n5297 240.244
R6205 gnd.n5294 gnd.n5293 240.244
R6206 gnd.n5290 gnd.n5289 240.244
R6207 gnd.n5286 gnd.n5285 240.244
R6208 gnd.n5275 gnd.n1189 240.244
R6209 gnd.n5275 gnd.n1262 240.244
R6210 gnd.n5271 gnd.n1262 240.244
R6211 gnd.n5271 gnd.n1269 240.244
R6212 gnd.n5263 gnd.n1269 240.244
R6213 gnd.n5263 gnd.n1286 240.244
R6214 gnd.n5259 gnd.n1286 240.244
R6215 gnd.n5259 gnd.n1292 240.244
R6216 gnd.n5251 gnd.n1292 240.244
R6217 gnd.n5251 gnd.n1304 240.244
R6218 gnd.n5247 gnd.n1304 240.244
R6219 gnd.n5247 gnd.n1310 240.244
R6220 gnd.n5239 gnd.n1310 240.244
R6221 gnd.n5239 gnd.n1324 240.244
R6222 gnd.n5235 gnd.n1324 240.244
R6223 gnd.n5235 gnd.n1330 240.244
R6224 gnd.n5227 gnd.n1330 240.244
R6225 gnd.n5227 gnd.n1342 240.244
R6226 gnd.n5223 gnd.n1342 240.244
R6227 gnd.n5223 gnd.n1348 240.244
R6228 gnd.n5215 gnd.n1348 240.244
R6229 gnd.n5215 gnd.n1362 240.244
R6230 gnd.n5211 gnd.n1362 240.244
R6231 gnd.n5211 gnd.n1368 240.244
R6232 gnd.n5203 gnd.n1368 240.244
R6233 gnd.n5203 gnd.n1380 240.244
R6234 gnd.n5199 gnd.n1380 240.244
R6235 gnd.n5199 gnd.n1385 240.244
R6236 gnd.n5191 gnd.n1385 240.244
R6237 gnd.n5191 gnd.n1400 240.244
R6238 gnd.n2880 gnd.n1400 240.244
R6239 gnd.n2880 gnd.n2794 240.244
R6240 gnd.n3041 gnd.n2794 240.244
R6241 gnd.n3045 gnd.n3041 240.244
R6242 gnd.n3045 gnd.n3042 240.244
R6243 gnd.n3042 gnd.n1410 240.244
R6244 gnd.n5186 gnd.n1410 240.244
R6245 gnd.n5186 gnd.n1411 240.244
R6246 gnd.n5178 gnd.n1411 240.244
R6247 gnd.n5178 gnd.n1427 240.244
R6248 gnd.n5174 gnd.n1427 240.244
R6249 gnd.n5174 gnd.n1432 240.244
R6250 gnd.n5166 gnd.n1432 240.244
R6251 gnd.n5166 gnd.n1447 240.244
R6252 gnd.n5162 gnd.n1447 240.244
R6253 gnd.n5162 gnd.n1453 240.244
R6254 gnd.n5154 gnd.n1453 240.244
R6255 gnd.n5154 gnd.n1467 240.244
R6256 gnd.n5150 gnd.n1467 240.244
R6257 gnd.n5150 gnd.n1473 240.244
R6258 gnd.n5142 gnd.n1473 240.244
R6259 gnd.n5142 gnd.n1488 240.244
R6260 gnd.n5138 gnd.n1488 240.244
R6261 gnd.n5138 gnd.n1494 240.244
R6262 gnd.n5130 gnd.n1494 240.244
R6263 gnd.n5130 gnd.n1508 240.244
R6264 gnd.n5126 gnd.n1508 240.244
R6265 gnd.n5126 gnd.n1514 240.244
R6266 gnd.n5118 gnd.n1514 240.244
R6267 gnd.n5118 gnd.n1529 240.244
R6268 gnd.n5114 gnd.n1529 240.244
R6269 gnd.n5114 gnd.n1535 240.244
R6270 gnd.n5106 gnd.n1535 240.244
R6271 gnd.n5106 gnd.n1550 240.244
R6272 gnd.n5407 gnd.n5403 240.244
R6273 gnd.n6867 gnd.n6866 240.244
R6274 gnd.n6864 gnd.n5411 240.244
R6275 gnd.n6860 gnd.n6859 240.244
R6276 gnd.n6857 gnd.n5418 240.244
R6277 gnd.n6853 gnd.n6852 240.244
R6278 gnd.n6850 gnd.n5425 240.244
R6279 gnd.n6846 gnd.n6845 240.244
R6280 gnd.n6434 gnd.n6010 240.244
R6281 gnd.n6010 gnd.n6001 240.244
R6282 gnd.n6455 gnd.n6001 240.244
R6283 gnd.n6455 gnd.n5994 240.244
R6284 gnd.n6465 gnd.n5994 240.244
R6285 gnd.n6465 gnd.n5985 240.244
R6286 gnd.n5985 gnd.n5974 240.244
R6287 gnd.n6486 gnd.n5974 240.244
R6288 gnd.n6486 gnd.n5968 240.244
R6289 gnd.n6496 gnd.n5968 240.244
R6290 gnd.n6496 gnd.n5959 240.244
R6291 gnd.n5959 gnd.n5948 240.244
R6292 gnd.n6517 gnd.n5948 240.244
R6293 gnd.n6517 gnd.n5942 240.244
R6294 gnd.n6527 gnd.n5942 240.244
R6295 gnd.n6527 gnd.n5933 240.244
R6296 gnd.n5933 gnd.n5923 240.244
R6297 gnd.n6548 gnd.n5923 240.244
R6298 gnd.n6548 gnd.n5916 240.244
R6299 gnd.n6558 gnd.n5916 240.244
R6300 gnd.n6558 gnd.n5907 240.244
R6301 gnd.n5907 gnd.n5898 240.244
R6302 gnd.n6579 gnd.n5898 240.244
R6303 gnd.n6579 gnd.n5891 240.244
R6304 gnd.n6589 gnd.n5891 240.244
R6305 gnd.n6589 gnd.n5882 240.244
R6306 gnd.n5882 gnd.n5873 240.244
R6307 gnd.n6610 gnd.n5873 240.244
R6308 gnd.n6610 gnd.n5866 240.244
R6309 gnd.n6620 gnd.n5866 240.244
R6310 gnd.n6620 gnd.n5858 240.244
R6311 gnd.n5858 gnd.n5849 240.244
R6312 gnd.n6640 gnd.n5849 240.244
R6313 gnd.n6640 gnd.n5836 240.244
R6314 gnd.n6661 gnd.n5836 240.244
R6315 gnd.n6661 gnd.n5825 240.244
R6316 gnd.n5825 gnd.n5816 240.244
R6317 gnd.n6684 gnd.n5816 240.244
R6318 gnd.n6685 gnd.n6684 240.244
R6319 gnd.n6686 gnd.n6685 240.244
R6320 gnd.n6686 gnd.n5796 240.244
R6321 gnd.n6714 gnd.n5796 240.244
R6322 gnd.n6714 gnd.n5787 240.244
R6323 gnd.n6730 gnd.n5787 240.244
R6324 gnd.n6731 gnd.n6730 240.244
R6325 gnd.n6731 gnd.n5769 240.244
R6326 gnd.n6758 gnd.n5769 240.244
R6327 gnd.n6758 gnd.n5753 240.244
R6328 gnd.n6773 gnd.n5753 240.244
R6329 gnd.n6773 gnd.n6772 240.244
R6330 gnd.n6772 gnd.n5760 240.244
R6331 gnd.n5760 gnd.n5754 240.244
R6332 gnd.n5754 gnd.n1147 240.244
R6333 gnd.n6371 gnd.n6370 240.244
R6334 gnd.n6415 gnd.n6370 240.244
R6335 gnd.n6413 gnd.n6412 240.244
R6336 gnd.n6409 gnd.n6408 240.244
R6337 gnd.n6405 gnd.n6404 240.244
R6338 gnd.n6401 gnd.n6400 240.244
R6339 gnd.n6397 gnd.n6396 240.244
R6340 gnd.n6393 gnd.n6392 240.244
R6341 gnd.n6445 gnd.n6008 240.244
R6342 gnd.n6445 gnd.n6003 240.244
R6343 gnd.n6453 gnd.n6003 240.244
R6344 gnd.n6453 gnd.n6004 240.244
R6345 gnd.n6004 gnd.n5983 240.244
R6346 gnd.n6476 gnd.n5983 240.244
R6347 gnd.n6476 gnd.n5977 240.244
R6348 gnd.n6484 gnd.n5977 240.244
R6349 gnd.n6484 gnd.n5979 240.244
R6350 gnd.n5979 gnd.n5957 240.244
R6351 gnd.n6507 gnd.n5957 240.244
R6352 gnd.n6507 gnd.n5951 240.244
R6353 gnd.n6515 gnd.n5951 240.244
R6354 gnd.n6515 gnd.n5953 240.244
R6355 gnd.n5953 gnd.n5931 240.244
R6356 gnd.n6538 gnd.n5931 240.244
R6357 gnd.n6538 gnd.n5926 240.244
R6358 gnd.n6546 gnd.n5926 240.244
R6359 gnd.n6546 gnd.n5927 240.244
R6360 gnd.n5927 gnd.n5905 240.244
R6361 gnd.n6569 gnd.n5905 240.244
R6362 gnd.n6569 gnd.n5900 240.244
R6363 gnd.n6577 gnd.n5900 240.244
R6364 gnd.n6577 gnd.n5901 240.244
R6365 gnd.n5901 gnd.n5880 240.244
R6366 gnd.n6600 gnd.n5880 240.244
R6367 gnd.n6600 gnd.n5875 240.244
R6368 gnd.n6608 gnd.n5875 240.244
R6369 gnd.n6608 gnd.n5876 240.244
R6370 gnd.n5876 gnd.n5856 240.244
R6371 gnd.n6630 gnd.n5856 240.244
R6372 gnd.n6630 gnd.n5851 240.244
R6373 gnd.n6638 gnd.n5851 240.244
R6374 gnd.n6638 gnd.n5852 240.244
R6375 gnd.n5852 gnd.n5824 240.244
R6376 gnd.n6671 gnd.n5824 240.244
R6377 gnd.n6671 gnd.n5819 240.244
R6378 gnd.n6682 gnd.n5819 240.244
R6379 gnd.n6682 gnd.n5820 240.244
R6380 gnd.n6678 gnd.n5820 240.244
R6381 gnd.n6678 gnd.n5794 240.244
R6382 gnd.n6718 gnd.n5794 240.244
R6383 gnd.n6718 gnd.n5789 240.244
R6384 gnd.n6728 gnd.n5789 240.244
R6385 gnd.n6728 gnd.n5790 240.244
R6386 gnd.n5790 gnd.n5767 240.244
R6387 gnd.n6761 gnd.n5767 240.244
R6388 gnd.n6762 gnd.n6761 240.244
R6389 gnd.n6762 gnd.n5762 240.244
R6390 gnd.n6770 gnd.n5762 240.244
R6391 gnd.n6770 gnd.n5763 240.244
R6392 gnd.n5763 gnd.n5402 240.244
R6393 gnd.n6874 gnd.n5402 240.244
R6394 gnd.n355 gnd.n257 240.244
R6395 gnd.n481 gnd.n480 240.244
R6396 gnd.n477 gnd.n476 240.244
R6397 gnd.n473 gnd.n472 240.244
R6398 gnd.n469 gnd.n468 240.244
R6399 gnd.n465 gnd.n464 240.244
R6400 gnd.n461 gnd.n460 240.244
R6401 gnd.n457 gnd.n456 240.244
R6402 gnd.n453 gnd.n452 240.244
R6403 gnd.n1940 gnd.n1935 240.244
R6404 gnd.n4572 gnd.n1940 240.244
R6405 gnd.n4572 gnd.n1952 240.244
R6406 gnd.n4580 gnd.n1952 240.244
R6407 gnd.n4580 gnd.n1963 240.244
R6408 gnd.n4586 gnd.n1963 240.244
R6409 gnd.n4586 gnd.n1974 240.244
R6410 gnd.n4594 gnd.n1974 240.244
R6411 gnd.n4594 gnd.n1984 240.244
R6412 gnd.n4600 gnd.n1984 240.244
R6413 gnd.n4600 gnd.n1994 240.244
R6414 gnd.n4608 gnd.n1994 240.244
R6415 gnd.n4608 gnd.n2004 240.244
R6416 gnd.n4614 gnd.n2004 240.244
R6417 gnd.n4614 gnd.n2015 240.244
R6418 gnd.n4625 gnd.n2015 240.244
R6419 gnd.n4625 gnd.n2025 240.244
R6420 gnd.n4639 gnd.n2025 240.244
R6421 gnd.n4639 gnd.n2036 240.244
R6422 gnd.n2044 gnd.n2036 240.244
R6423 gnd.n4630 gnd.n2044 240.244
R6424 gnd.n4630 gnd.n544 240.244
R6425 gnd.n544 gnd.n531 240.244
R6426 gnd.n7769 gnd.n531 240.244
R6427 gnd.n7769 gnd.n527 240.244
R6428 gnd.n7775 gnd.n527 240.244
R6429 gnd.n7775 gnd.n509 240.244
R6430 gnd.n7796 gnd.n509 240.244
R6431 gnd.n7796 gnd.n504 240.244
R6432 gnd.n7802 gnd.n504 240.244
R6433 gnd.n7802 gnd.n499 240.244
R6434 gnd.n7807 gnd.n499 240.244
R6435 gnd.n7807 gnd.n102 240.244
R6436 gnd.n8098 gnd.n102 240.244
R6437 gnd.n8098 gnd.n104 240.244
R6438 gnd.n389 gnd.n104 240.244
R6439 gnd.n389 gnd.n124 240.244
R6440 gnd.n394 gnd.n124 240.244
R6441 gnd.n394 gnd.n135 240.244
R6442 gnd.n397 gnd.n135 240.244
R6443 gnd.n397 gnd.n144 240.244
R6444 gnd.n402 gnd.n144 240.244
R6445 gnd.n402 gnd.n153 240.244
R6446 gnd.n405 gnd.n153 240.244
R6447 gnd.n405 gnd.n163 240.244
R6448 gnd.n410 gnd.n163 240.244
R6449 gnd.n410 gnd.n172 240.244
R6450 gnd.n413 gnd.n172 240.244
R6451 gnd.n413 gnd.n182 240.244
R6452 gnd.n418 gnd.n182 240.244
R6453 gnd.n418 gnd.n191 240.244
R6454 gnd.n421 gnd.n191 240.244
R6455 gnd.n421 gnd.n201 240.244
R6456 gnd.n426 gnd.n201 240.244
R6457 gnd.n426 gnd.n210 240.244
R6458 gnd.n429 gnd.n210 240.244
R6459 gnd.n429 gnd.n221 240.244
R6460 gnd.n434 gnd.n221 240.244
R6461 gnd.n434 gnd.n230 240.244
R6462 gnd.n437 gnd.n230 240.244
R6463 gnd.n437 gnd.n240 240.244
R6464 gnd.n442 gnd.n240 240.244
R6465 gnd.n442 gnd.n249 240.244
R6466 gnd.n446 gnd.n249 240.244
R6467 gnd.n4479 gnd.n4478 240.244
R6468 gnd.n4495 gnd.n4494 240.244
R6469 gnd.n4498 gnd.n4497 240.244
R6470 gnd.n4514 gnd.n4513 240.244
R6471 gnd.n4517 gnd.n4516 240.244
R6472 gnd.n4533 gnd.n4532 240.244
R6473 gnd.n4536 gnd.n4535 240.244
R6474 gnd.n4551 gnd.n4550 240.244
R6475 gnd.n4416 gnd.n1858 240.244
R6476 gnd.n4715 gnd.n4714 240.244
R6477 gnd.n4714 gnd.n1938 240.244
R6478 gnd.n4706 gnd.n1938 240.244
R6479 gnd.n4706 gnd.n1954 240.244
R6480 gnd.n4702 gnd.n1954 240.244
R6481 gnd.n4702 gnd.n1960 240.244
R6482 gnd.n4694 gnd.n1960 240.244
R6483 gnd.n4694 gnd.n1976 240.244
R6484 gnd.n4690 gnd.n1976 240.244
R6485 gnd.n4690 gnd.n1981 240.244
R6486 gnd.n4682 gnd.n1981 240.244
R6487 gnd.n4682 gnd.n1996 240.244
R6488 gnd.n4678 gnd.n1996 240.244
R6489 gnd.n4678 gnd.n2001 240.244
R6490 gnd.n4670 gnd.n2001 240.244
R6491 gnd.n4670 gnd.n2017 240.244
R6492 gnd.n4666 gnd.n2017 240.244
R6493 gnd.n4666 gnd.n2022 240.244
R6494 gnd.n4658 gnd.n2022 240.244
R6495 gnd.n4658 gnd.n2038 240.244
R6496 gnd.n2038 gnd.n545 240.244
R6497 gnd.n7756 gnd.n545 240.244
R6498 gnd.n7756 gnd.n546 240.244
R6499 gnd.n546 gnd.n535 240.244
R6500 gnd.n7751 gnd.n535 240.244
R6501 gnd.n7751 gnd.n517 240.244
R6502 gnd.n7789 gnd.n517 240.244
R6503 gnd.n7789 gnd.n512 240.244
R6504 gnd.n7785 gnd.n512 240.244
R6505 gnd.n7785 gnd.n496 240.244
R6506 gnd.n7814 gnd.n496 240.244
R6507 gnd.n7814 gnd.n490 240.244
R6508 gnd.n7823 gnd.n490 240.244
R6509 gnd.n7823 gnd.n108 240.244
R6510 gnd.n7826 gnd.n108 240.244
R6511 gnd.n7826 gnd.n126 240.244
R6512 gnd.n8088 gnd.n126 240.244
R6513 gnd.n8088 gnd.n127 240.244
R6514 gnd.n8084 gnd.n127 240.244
R6515 gnd.n8084 gnd.n133 240.244
R6516 gnd.n8076 gnd.n133 240.244
R6517 gnd.n8076 gnd.n145 240.244
R6518 gnd.n8072 gnd.n145 240.244
R6519 gnd.n8072 gnd.n150 240.244
R6520 gnd.n8064 gnd.n150 240.244
R6521 gnd.n8064 gnd.n165 240.244
R6522 gnd.n8060 gnd.n165 240.244
R6523 gnd.n8060 gnd.n170 240.244
R6524 gnd.n8052 gnd.n170 240.244
R6525 gnd.n8052 gnd.n183 240.244
R6526 gnd.n8048 gnd.n183 240.244
R6527 gnd.n8048 gnd.n188 240.244
R6528 gnd.n8040 gnd.n188 240.244
R6529 gnd.n8040 gnd.n203 240.244
R6530 gnd.n8036 gnd.n203 240.244
R6531 gnd.n8036 gnd.n208 240.244
R6532 gnd.n8028 gnd.n208 240.244
R6533 gnd.n8028 gnd.n222 240.244
R6534 gnd.n8024 gnd.n222 240.244
R6535 gnd.n8024 gnd.n227 240.244
R6536 gnd.n8016 gnd.n227 240.244
R6537 gnd.n8016 gnd.n242 240.244
R6538 gnd.n8012 gnd.n242 240.244
R6539 gnd.n8012 gnd.n247 240.244
R6540 gnd.n5437 gnd.n1144 240.244
R6541 gnd.n6835 gnd.n6834 240.244
R6542 gnd.n6832 gnd.n5441 240.244
R6543 gnd.n6828 gnd.n6827 240.244
R6544 gnd.n6825 gnd.n5448 240.244
R6545 gnd.n6821 gnd.n6820 240.244
R6546 gnd.n6818 gnd.n5455 240.244
R6547 gnd.n6814 gnd.n6813 240.244
R6548 gnd.n6811 gnd.n5462 240.244
R6549 gnd.n6807 gnd.n6806 240.244
R6550 gnd.n6804 gnd.n5469 240.244
R6551 gnd.n6800 gnd.n6799 240.244
R6552 gnd.n6797 gnd.n5479 240.244
R6553 gnd.n6157 gnd.n6053 240.244
R6554 gnd.n6163 gnd.n6053 240.244
R6555 gnd.n6163 gnd.n6045 240.244
R6556 gnd.n6173 gnd.n6045 240.244
R6557 gnd.n6173 gnd.n6041 240.244
R6558 gnd.n6179 gnd.n6041 240.244
R6559 gnd.n6179 gnd.n6032 240.244
R6560 gnd.n6189 gnd.n6032 240.244
R6561 gnd.n6189 gnd.n6027 240.244
R6562 gnd.n6362 gnd.n6027 240.244
R6563 gnd.n6362 gnd.n6028 240.244
R6564 gnd.n6028 gnd.n6020 240.244
R6565 gnd.n6357 gnd.n6020 240.244
R6566 gnd.n6357 gnd.n6011 240.244
R6567 gnd.n6354 gnd.n6011 240.244
R6568 gnd.n6354 gnd.n6353 240.244
R6569 gnd.n6353 gnd.n5996 240.244
R6570 gnd.n6348 gnd.n5996 240.244
R6571 gnd.n6348 gnd.n5986 240.244
R6572 gnd.n6345 gnd.n5986 240.244
R6573 gnd.n6345 gnd.n6344 240.244
R6574 gnd.n6344 gnd.n5969 240.244
R6575 gnd.n6340 gnd.n5969 240.244
R6576 gnd.n6340 gnd.n5960 240.244
R6577 gnd.n6337 gnd.n5960 240.244
R6578 gnd.n6337 gnd.n6336 240.244
R6579 gnd.n6336 gnd.n5943 240.244
R6580 gnd.n6332 gnd.n5943 240.244
R6581 gnd.n6332 gnd.n5934 240.244
R6582 gnd.n6245 gnd.n5934 240.244
R6583 gnd.n6246 gnd.n6245 240.244
R6584 gnd.n6246 gnd.n5918 240.244
R6585 gnd.n6242 gnd.n5918 240.244
R6586 gnd.n6242 gnd.n5908 240.244
R6587 gnd.n6238 gnd.n5908 240.244
R6588 gnd.n6238 gnd.n6237 240.244
R6589 gnd.n6237 gnd.n5893 240.244
R6590 gnd.n6232 gnd.n5893 240.244
R6591 gnd.n6232 gnd.n5883 240.244
R6592 gnd.n6229 gnd.n5883 240.244
R6593 gnd.n6229 gnd.n6227 240.244
R6594 gnd.n6227 gnd.n5868 240.244
R6595 gnd.n6223 gnd.n5868 240.244
R6596 gnd.n6223 gnd.n5859 240.244
R6597 gnd.n5859 gnd.n5842 240.244
R6598 gnd.n6650 gnd.n5842 240.244
R6599 gnd.n6650 gnd.n5838 240.244
R6600 gnd.n6658 gnd.n5838 240.244
R6601 gnd.n6658 gnd.n5826 240.244
R6602 gnd.n5826 gnd.n5807 240.244
R6603 gnd.n6694 gnd.n5807 240.244
R6604 gnd.n6694 gnd.n5802 240.244
R6605 gnd.n6702 gnd.n5802 240.244
R6606 gnd.n6702 gnd.n5803 240.244
R6607 gnd.n5803 gnd.n5780 240.244
R6608 gnd.n6739 gnd.n5780 240.244
R6609 gnd.n6739 gnd.n5775 240.244
R6610 gnd.n6747 gnd.n5775 240.244
R6611 gnd.n6747 gnd.n5776 240.244
R6612 gnd.n5776 gnd.n5487 240.244
R6613 gnd.n6780 gnd.n5487 240.244
R6614 gnd.n6780 gnd.n5488 240.244
R6615 gnd.n5488 gnd.n1136 240.244
R6616 gnd.n6787 gnd.n1136 240.244
R6617 gnd.n6787 gnd.n1146 240.244
R6618 gnd.n6149 gnd.n6147 240.244
R6619 gnd.n6147 gnd.n6146 240.244
R6620 gnd.n6143 gnd.n6142 240.244
R6621 gnd.n6140 gnd.n6066 240.244
R6622 gnd.n6136 gnd.n6134 240.244
R6623 gnd.n6132 gnd.n6072 240.244
R6624 gnd.n6128 gnd.n6126 240.244
R6625 gnd.n6124 gnd.n6078 240.244
R6626 gnd.n6120 gnd.n6118 240.244
R6627 gnd.n6116 gnd.n6084 240.244
R6628 gnd.n6112 gnd.n6110 240.244
R6629 gnd.n6108 gnd.n6090 240.244
R6630 gnd.n6103 gnd.n6101 240.244
R6631 gnd.n6155 gnd.n6051 240.244
R6632 gnd.n6165 gnd.n6051 240.244
R6633 gnd.n6165 gnd.n6047 240.244
R6634 gnd.n6171 gnd.n6047 240.244
R6635 gnd.n6171 gnd.n6039 240.244
R6636 gnd.n6181 gnd.n6039 240.244
R6637 gnd.n6181 gnd.n6035 240.244
R6638 gnd.n6187 gnd.n6035 240.244
R6639 gnd.n6187 gnd.n6026 240.244
R6640 gnd.n6424 gnd.n6026 240.244
R6641 gnd.n6424 gnd.n6021 240.244
R6642 gnd.n6431 gnd.n6021 240.244
R6643 gnd.n6431 gnd.n6013 240.244
R6644 gnd.n6442 gnd.n6013 240.244
R6645 gnd.n6442 gnd.n6014 240.244
R6646 gnd.n6014 gnd.n5997 240.244
R6647 gnd.n6462 gnd.n5997 240.244
R6648 gnd.n6462 gnd.n5988 240.244
R6649 gnd.n6473 gnd.n5988 240.244
R6650 gnd.n6473 gnd.n5989 240.244
R6651 gnd.n5989 gnd.n5970 240.244
R6652 gnd.n6493 gnd.n5970 240.244
R6653 gnd.n6493 gnd.n5962 240.244
R6654 gnd.n6504 gnd.n5962 240.244
R6655 gnd.n6504 gnd.n5963 240.244
R6656 gnd.n5963 gnd.n5944 240.244
R6657 gnd.n6524 gnd.n5944 240.244
R6658 gnd.n6524 gnd.n5936 240.244
R6659 gnd.n6535 gnd.n5936 240.244
R6660 gnd.n6535 gnd.n5937 240.244
R6661 gnd.n5937 gnd.n5919 240.244
R6662 gnd.n6555 gnd.n5919 240.244
R6663 gnd.n6555 gnd.n5910 240.244
R6664 gnd.n6566 gnd.n5910 240.244
R6665 gnd.n6566 gnd.n5911 240.244
R6666 gnd.n5911 gnd.n5894 240.244
R6667 gnd.n6586 gnd.n5894 240.244
R6668 gnd.n6586 gnd.n5885 240.244
R6669 gnd.n6597 gnd.n5885 240.244
R6670 gnd.n6597 gnd.n5886 240.244
R6671 gnd.n5886 gnd.n5869 240.244
R6672 gnd.n6617 gnd.n5869 240.244
R6673 gnd.n6617 gnd.n5861 240.244
R6674 gnd.n6627 gnd.n5861 240.244
R6675 gnd.n6627 gnd.n5844 240.244
R6676 gnd.n6648 gnd.n5844 240.244
R6677 gnd.n6648 gnd.n5845 240.244
R6678 gnd.n5845 gnd.n5828 240.244
R6679 gnd.n6668 gnd.n5828 240.244
R6680 gnd.n6668 gnd.n5810 240.244
R6681 gnd.n6692 gnd.n5810 240.244
R6682 gnd.n6692 gnd.n5800 240.244
R6683 gnd.n6705 gnd.n5800 240.244
R6684 gnd.n6706 gnd.n6705 240.244
R6685 gnd.n6706 gnd.n5781 240.244
R6686 gnd.n6737 gnd.n5781 240.244
R6687 gnd.n6737 gnd.n5773 240.244
R6688 gnd.n6750 gnd.n5773 240.244
R6689 gnd.n6751 gnd.n6750 240.244
R6690 gnd.n6751 gnd.n5491 240.244
R6691 gnd.n6778 gnd.n5491 240.244
R6692 gnd.n6778 gnd.n1138 240.244
R6693 gnd.n6881 gnd.n1138 240.244
R6694 gnd.n6881 gnd.n1139 240.244
R6695 gnd.n6877 gnd.n1139 240.244
R6696 gnd.n3234 gnd.n1557 240.244
R6697 gnd.n3236 gnd.n3235 240.244
R6698 gnd.n3246 gnd.n3245 240.244
R6699 gnd.n3254 gnd.n3253 240.244
R6700 gnd.n3256 gnd.n3255 240.244
R6701 gnd.n3266 gnd.n3265 240.244
R6702 gnd.n3274 gnd.n3273 240.244
R6703 gnd.n3276 gnd.n3275 240.244
R6704 gnd.n3290 gnd.n3289 240.244
R6705 gnd.n2958 gnd.n1260 240.244
R6706 gnd.n2961 gnd.n1260 240.244
R6707 gnd.n2961 gnd.n1272 240.244
R6708 gnd.n2966 gnd.n1272 240.244
R6709 gnd.n2966 gnd.n1284 240.244
R6710 gnd.n2969 gnd.n1284 240.244
R6711 gnd.n2969 gnd.n1294 240.244
R6712 gnd.n2974 gnd.n1294 240.244
R6713 gnd.n2974 gnd.n1303 240.244
R6714 gnd.n2977 gnd.n1303 240.244
R6715 gnd.n2977 gnd.n1313 240.244
R6716 gnd.n2982 gnd.n1313 240.244
R6717 gnd.n2982 gnd.n1322 240.244
R6718 gnd.n2985 gnd.n1322 240.244
R6719 gnd.n2985 gnd.n1332 240.244
R6720 gnd.n2990 gnd.n1332 240.244
R6721 gnd.n2990 gnd.n1341 240.244
R6722 gnd.n2993 gnd.n1341 240.244
R6723 gnd.n2993 gnd.n1351 240.244
R6724 gnd.n2998 gnd.n1351 240.244
R6725 gnd.n2998 gnd.n1360 240.244
R6726 gnd.n3001 gnd.n1360 240.244
R6727 gnd.n3001 gnd.n1370 240.244
R6728 gnd.n3006 gnd.n1370 240.244
R6729 gnd.n3006 gnd.n1379 240.244
R6730 gnd.n3009 gnd.n1379 240.244
R6731 gnd.n3009 gnd.n1388 240.244
R6732 gnd.n3014 gnd.n1388 240.244
R6733 gnd.n3014 gnd.n1398 240.244
R6734 gnd.n3017 gnd.n1398 240.244
R6735 gnd.n3017 gnd.n2882 240.244
R6736 gnd.n3023 gnd.n2882 240.244
R6737 gnd.n3023 gnd.n2790 240.244
R6738 gnd.n3047 gnd.n2790 240.244
R6739 gnd.n3047 gnd.n2786 240.244
R6740 gnd.n3053 gnd.n2786 240.244
R6741 gnd.n3053 gnd.n1414 240.244
R6742 gnd.n3086 gnd.n1414 240.244
R6743 gnd.n3086 gnd.n1425 240.244
R6744 gnd.n3092 gnd.n1425 240.244
R6745 gnd.n3092 gnd.n1435 240.244
R6746 gnd.n3100 gnd.n1435 240.244
R6747 gnd.n3100 gnd.n1445 240.244
R6748 gnd.n3106 gnd.n1445 240.244
R6749 gnd.n3106 gnd.n1456 240.244
R6750 gnd.n3141 gnd.n1456 240.244
R6751 gnd.n3141 gnd.n1465 240.244
R6752 gnd.n2763 gnd.n1465 240.244
R6753 gnd.n2763 gnd.n1476 240.244
R6754 gnd.n2764 gnd.n1476 240.244
R6755 gnd.n2764 gnd.n1486 240.244
R6756 gnd.n3126 gnd.n1486 240.244
R6757 gnd.n3126 gnd.n1497 240.244
R6758 gnd.n2746 gnd.n1497 240.244
R6759 gnd.n2746 gnd.n1506 240.244
R6760 gnd.n3194 gnd.n1506 240.244
R6761 gnd.n3194 gnd.n1517 240.244
R6762 gnd.n3200 gnd.n1517 240.244
R6763 gnd.n3200 gnd.n1527 240.244
R6764 gnd.n3209 gnd.n1527 240.244
R6765 gnd.n3209 gnd.n1538 240.244
R6766 gnd.n3217 gnd.n1538 240.244
R6767 gnd.n3217 gnd.n1548 240.244
R6768 gnd.n3362 gnd.n1548 240.244
R6769 gnd.n2918 gnd.n2917 240.244
R6770 gnd.n2924 gnd.n2923 240.244
R6771 gnd.n2928 gnd.n2927 240.244
R6772 gnd.n2934 gnd.n2933 240.244
R6773 gnd.n2938 gnd.n2937 240.244
R6774 gnd.n2944 gnd.n2943 240.244
R6775 gnd.n2948 gnd.n2947 240.244
R6776 gnd.n2905 gnd.n2904 240.244
R6777 gnd.n2900 gnd.n1185 240.244
R6778 gnd.n2913 gnd.n1261 240.244
R6779 gnd.n1274 gnd.n1261 240.244
R6780 gnd.n5269 gnd.n1274 240.244
R6781 gnd.n5269 gnd.n1275 240.244
R6782 gnd.n5265 gnd.n1275 240.244
R6783 gnd.n5265 gnd.n1282 240.244
R6784 gnd.n5257 gnd.n1282 240.244
R6785 gnd.n5257 gnd.n1296 240.244
R6786 gnd.n5253 gnd.n1296 240.244
R6787 gnd.n5253 gnd.n1301 240.244
R6788 gnd.n5245 gnd.n1301 240.244
R6789 gnd.n5245 gnd.n1315 240.244
R6790 gnd.n5241 gnd.n1315 240.244
R6791 gnd.n5241 gnd.n1320 240.244
R6792 gnd.n5233 gnd.n1320 240.244
R6793 gnd.n5233 gnd.n1334 240.244
R6794 gnd.n5229 gnd.n1334 240.244
R6795 gnd.n5229 gnd.n1339 240.244
R6796 gnd.n5221 gnd.n1339 240.244
R6797 gnd.n5221 gnd.n1353 240.244
R6798 gnd.n5217 gnd.n1353 240.244
R6799 gnd.n5217 gnd.n1358 240.244
R6800 gnd.n5209 gnd.n1358 240.244
R6801 gnd.n5209 gnd.n1372 240.244
R6802 gnd.n5205 gnd.n1372 240.244
R6803 gnd.n5205 gnd.n1377 240.244
R6804 gnd.n5197 gnd.n1377 240.244
R6805 gnd.n5197 gnd.n1390 240.244
R6806 gnd.n5193 gnd.n1390 240.244
R6807 gnd.n5193 gnd.n1395 240.244
R6808 gnd.n2878 gnd.n1395 240.244
R6809 gnd.n2878 gnd.n2800 240.244
R6810 gnd.n3039 gnd.n2800 240.244
R6811 gnd.n3039 gnd.n2793 240.244
R6812 gnd.n3035 gnd.n2793 240.244
R6813 gnd.n3035 gnd.n1416 240.244
R6814 gnd.n5184 gnd.n1416 240.244
R6815 gnd.n5184 gnd.n1417 240.244
R6816 gnd.n5180 gnd.n1417 240.244
R6817 gnd.n5180 gnd.n1423 240.244
R6818 gnd.n5172 gnd.n1423 240.244
R6819 gnd.n5172 gnd.n1437 240.244
R6820 gnd.n5168 gnd.n1437 240.244
R6821 gnd.n5168 gnd.n1442 240.244
R6822 gnd.n5160 gnd.n1442 240.244
R6823 gnd.n5160 gnd.n1458 240.244
R6824 gnd.n5156 gnd.n1458 240.244
R6825 gnd.n5156 gnd.n1463 240.244
R6826 gnd.n5148 gnd.n1463 240.244
R6827 gnd.n5148 gnd.n1478 240.244
R6828 gnd.n5144 gnd.n1478 240.244
R6829 gnd.n5144 gnd.n1483 240.244
R6830 gnd.n5136 gnd.n1483 240.244
R6831 gnd.n5136 gnd.n1499 240.244
R6832 gnd.n5132 gnd.n1499 240.244
R6833 gnd.n5132 gnd.n1504 240.244
R6834 gnd.n5124 gnd.n1504 240.244
R6835 gnd.n5124 gnd.n1519 240.244
R6836 gnd.n5120 gnd.n1519 240.244
R6837 gnd.n5120 gnd.n1524 240.244
R6838 gnd.n5112 gnd.n1524 240.244
R6839 gnd.n5112 gnd.n1540 240.244
R6840 gnd.n5108 gnd.n1540 240.244
R6841 gnd.n5108 gnd.n1545 240.244
R6842 gnd.n7053 gnd.n964 240.244
R6843 gnd.n7059 gnd.n964 240.244
R6844 gnd.n7059 gnd.n962 240.244
R6845 gnd.n7063 gnd.n962 240.244
R6846 gnd.n7063 gnd.n958 240.244
R6847 gnd.n7069 gnd.n958 240.244
R6848 gnd.n7069 gnd.n956 240.244
R6849 gnd.n7073 gnd.n956 240.244
R6850 gnd.n7073 gnd.n952 240.244
R6851 gnd.n7079 gnd.n952 240.244
R6852 gnd.n7079 gnd.n950 240.244
R6853 gnd.n7083 gnd.n950 240.244
R6854 gnd.n7083 gnd.n946 240.244
R6855 gnd.n7089 gnd.n946 240.244
R6856 gnd.n7089 gnd.n944 240.244
R6857 gnd.n7093 gnd.n944 240.244
R6858 gnd.n7093 gnd.n940 240.244
R6859 gnd.n7099 gnd.n940 240.244
R6860 gnd.n7099 gnd.n938 240.244
R6861 gnd.n7103 gnd.n938 240.244
R6862 gnd.n7103 gnd.n934 240.244
R6863 gnd.n7109 gnd.n934 240.244
R6864 gnd.n7109 gnd.n932 240.244
R6865 gnd.n7113 gnd.n932 240.244
R6866 gnd.n7113 gnd.n928 240.244
R6867 gnd.n7119 gnd.n928 240.244
R6868 gnd.n7119 gnd.n926 240.244
R6869 gnd.n7123 gnd.n926 240.244
R6870 gnd.n7123 gnd.n922 240.244
R6871 gnd.n7129 gnd.n922 240.244
R6872 gnd.n7129 gnd.n920 240.244
R6873 gnd.n7133 gnd.n920 240.244
R6874 gnd.n7133 gnd.n916 240.244
R6875 gnd.n7139 gnd.n916 240.244
R6876 gnd.n7139 gnd.n914 240.244
R6877 gnd.n7143 gnd.n914 240.244
R6878 gnd.n7143 gnd.n910 240.244
R6879 gnd.n7149 gnd.n910 240.244
R6880 gnd.n7149 gnd.n908 240.244
R6881 gnd.n7153 gnd.n908 240.244
R6882 gnd.n7153 gnd.n904 240.244
R6883 gnd.n7159 gnd.n904 240.244
R6884 gnd.n7159 gnd.n902 240.244
R6885 gnd.n7163 gnd.n902 240.244
R6886 gnd.n7163 gnd.n898 240.244
R6887 gnd.n7169 gnd.n898 240.244
R6888 gnd.n7169 gnd.n896 240.244
R6889 gnd.n7173 gnd.n896 240.244
R6890 gnd.n7173 gnd.n892 240.244
R6891 gnd.n7179 gnd.n892 240.244
R6892 gnd.n7179 gnd.n890 240.244
R6893 gnd.n7183 gnd.n890 240.244
R6894 gnd.n7183 gnd.n886 240.244
R6895 gnd.n7189 gnd.n886 240.244
R6896 gnd.n7189 gnd.n884 240.244
R6897 gnd.n7193 gnd.n884 240.244
R6898 gnd.n7193 gnd.n880 240.244
R6899 gnd.n7199 gnd.n880 240.244
R6900 gnd.n7199 gnd.n878 240.244
R6901 gnd.n7203 gnd.n878 240.244
R6902 gnd.n7203 gnd.n874 240.244
R6903 gnd.n7209 gnd.n874 240.244
R6904 gnd.n7209 gnd.n872 240.244
R6905 gnd.n7213 gnd.n872 240.244
R6906 gnd.n7213 gnd.n868 240.244
R6907 gnd.n7219 gnd.n868 240.244
R6908 gnd.n7219 gnd.n866 240.244
R6909 gnd.n7223 gnd.n866 240.244
R6910 gnd.n7223 gnd.n862 240.244
R6911 gnd.n7229 gnd.n862 240.244
R6912 gnd.n7229 gnd.n860 240.244
R6913 gnd.n7233 gnd.n860 240.244
R6914 gnd.n7233 gnd.n856 240.244
R6915 gnd.n7239 gnd.n856 240.244
R6916 gnd.n7239 gnd.n854 240.244
R6917 gnd.n7243 gnd.n854 240.244
R6918 gnd.n7243 gnd.n850 240.244
R6919 gnd.n7249 gnd.n850 240.244
R6920 gnd.n7249 gnd.n848 240.244
R6921 gnd.n7253 gnd.n848 240.244
R6922 gnd.n7253 gnd.n844 240.244
R6923 gnd.n7259 gnd.n844 240.244
R6924 gnd.n7259 gnd.n842 240.244
R6925 gnd.n7263 gnd.n842 240.244
R6926 gnd.n7263 gnd.n838 240.244
R6927 gnd.n7269 gnd.n838 240.244
R6928 gnd.n7269 gnd.n836 240.244
R6929 gnd.n7273 gnd.n836 240.244
R6930 gnd.n7273 gnd.n832 240.244
R6931 gnd.n7279 gnd.n832 240.244
R6932 gnd.n7279 gnd.n830 240.244
R6933 gnd.n7283 gnd.n830 240.244
R6934 gnd.n7283 gnd.n826 240.244
R6935 gnd.n7289 gnd.n826 240.244
R6936 gnd.n7289 gnd.n824 240.244
R6937 gnd.n7293 gnd.n824 240.244
R6938 gnd.n7293 gnd.n820 240.244
R6939 gnd.n7299 gnd.n820 240.244
R6940 gnd.n7299 gnd.n818 240.244
R6941 gnd.n7303 gnd.n818 240.244
R6942 gnd.n7303 gnd.n814 240.244
R6943 gnd.n7309 gnd.n814 240.244
R6944 gnd.n7309 gnd.n812 240.244
R6945 gnd.n7313 gnd.n812 240.244
R6946 gnd.n7313 gnd.n808 240.244
R6947 gnd.n7319 gnd.n808 240.244
R6948 gnd.n7319 gnd.n806 240.244
R6949 gnd.n7323 gnd.n806 240.244
R6950 gnd.n7323 gnd.n802 240.244
R6951 gnd.n7329 gnd.n802 240.244
R6952 gnd.n7329 gnd.n800 240.244
R6953 gnd.n7333 gnd.n800 240.244
R6954 gnd.n7333 gnd.n796 240.244
R6955 gnd.n7339 gnd.n796 240.244
R6956 gnd.n7339 gnd.n794 240.244
R6957 gnd.n7343 gnd.n794 240.244
R6958 gnd.n7343 gnd.n790 240.244
R6959 gnd.n7349 gnd.n790 240.244
R6960 gnd.n7349 gnd.n788 240.244
R6961 gnd.n7353 gnd.n788 240.244
R6962 gnd.n7353 gnd.n784 240.244
R6963 gnd.n7359 gnd.n784 240.244
R6964 gnd.n7359 gnd.n782 240.244
R6965 gnd.n7363 gnd.n782 240.244
R6966 gnd.n7363 gnd.n778 240.244
R6967 gnd.n7369 gnd.n778 240.244
R6968 gnd.n7369 gnd.n776 240.244
R6969 gnd.n7373 gnd.n776 240.244
R6970 gnd.n7373 gnd.n772 240.244
R6971 gnd.n7379 gnd.n772 240.244
R6972 gnd.n7379 gnd.n770 240.244
R6973 gnd.n7383 gnd.n770 240.244
R6974 gnd.n7383 gnd.n766 240.244
R6975 gnd.n7389 gnd.n766 240.244
R6976 gnd.n7389 gnd.n764 240.244
R6977 gnd.n7393 gnd.n764 240.244
R6978 gnd.n7393 gnd.n760 240.244
R6979 gnd.n7399 gnd.n760 240.244
R6980 gnd.n7399 gnd.n758 240.244
R6981 gnd.n7403 gnd.n758 240.244
R6982 gnd.n7403 gnd.n754 240.244
R6983 gnd.n7409 gnd.n754 240.244
R6984 gnd.n7409 gnd.n752 240.244
R6985 gnd.n7413 gnd.n752 240.244
R6986 gnd.n7413 gnd.n748 240.244
R6987 gnd.n7419 gnd.n748 240.244
R6988 gnd.n7419 gnd.n746 240.244
R6989 gnd.n7423 gnd.n746 240.244
R6990 gnd.n7423 gnd.n742 240.244
R6991 gnd.n7429 gnd.n742 240.244
R6992 gnd.n7429 gnd.n740 240.244
R6993 gnd.n7433 gnd.n740 240.244
R6994 gnd.n7433 gnd.n736 240.244
R6995 gnd.n7439 gnd.n736 240.244
R6996 gnd.n7439 gnd.n734 240.244
R6997 gnd.n7443 gnd.n734 240.244
R6998 gnd.n7443 gnd.n730 240.244
R6999 gnd.n7449 gnd.n730 240.244
R7000 gnd.n7449 gnd.n728 240.244
R7001 gnd.n7453 gnd.n728 240.244
R7002 gnd.n7453 gnd.n724 240.244
R7003 gnd.n7459 gnd.n724 240.244
R7004 gnd.n7459 gnd.n722 240.244
R7005 gnd.n7463 gnd.n722 240.244
R7006 gnd.n7463 gnd.n718 240.244
R7007 gnd.n7469 gnd.n718 240.244
R7008 gnd.n7469 gnd.n716 240.244
R7009 gnd.n7473 gnd.n716 240.244
R7010 gnd.n7473 gnd.n712 240.244
R7011 gnd.n7479 gnd.n712 240.244
R7012 gnd.n7479 gnd.n710 240.244
R7013 gnd.n7483 gnd.n710 240.244
R7014 gnd.n7483 gnd.n706 240.244
R7015 gnd.n7489 gnd.n706 240.244
R7016 gnd.n7489 gnd.n704 240.244
R7017 gnd.n7493 gnd.n704 240.244
R7018 gnd.n7493 gnd.n700 240.244
R7019 gnd.n7500 gnd.n700 240.244
R7020 gnd.n7500 gnd.n698 240.244
R7021 gnd.n7504 gnd.n698 240.244
R7022 gnd.n7504 gnd.n695 240.244
R7023 gnd.n7510 gnd.n693 240.244
R7024 gnd.n7514 gnd.n693 240.244
R7025 gnd.n7514 gnd.n689 240.244
R7026 gnd.n7520 gnd.n689 240.244
R7027 gnd.n7520 gnd.n687 240.244
R7028 gnd.n7524 gnd.n687 240.244
R7029 gnd.n7524 gnd.n683 240.244
R7030 gnd.n7530 gnd.n683 240.244
R7031 gnd.n7530 gnd.n681 240.244
R7032 gnd.n7534 gnd.n681 240.244
R7033 gnd.n7534 gnd.n677 240.244
R7034 gnd.n7540 gnd.n677 240.244
R7035 gnd.n7540 gnd.n675 240.244
R7036 gnd.n7544 gnd.n675 240.244
R7037 gnd.n7544 gnd.n671 240.244
R7038 gnd.n7550 gnd.n671 240.244
R7039 gnd.n7550 gnd.n669 240.244
R7040 gnd.n7554 gnd.n669 240.244
R7041 gnd.n7554 gnd.n665 240.244
R7042 gnd.n7560 gnd.n665 240.244
R7043 gnd.n7560 gnd.n663 240.244
R7044 gnd.n7564 gnd.n663 240.244
R7045 gnd.n7564 gnd.n659 240.244
R7046 gnd.n7570 gnd.n659 240.244
R7047 gnd.n7570 gnd.n657 240.244
R7048 gnd.n7574 gnd.n657 240.244
R7049 gnd.n7574 gnd.n653 240.244
R7050 gnd.n7580 gnd.n653 240.244
R7051 gnd.n7580 gnd.n651 240.244
R7052 gnd.n7584 gnd.n651 240.244
R7053 gnd.n7584 gnd.n647 240.244
R7054 gnd.n7590 gnd.n647 240.244
R7055 gnd.n7590 gnd.n645 240.244
R7056 gnd.n7594 gnd.n645 240.244
R7057 gnd.n7594 gnd.n641 240.244
R7058 gnd.n7600 gnd.n641 240.244
R7059 gnd.n7600 gnd.n639 240.244
R7060 gnd.n7604 gnd.n639 240.244
R7061 gnd.n7604 gnd.n635 240.244
R7062 gnd.n7610 gnd.n635 240.244
R7063 gnd.n7610 gnd.n633 240.244
R7064 gnd.n7614 gnd.n633 240.244
R7065 gnd.n7614 gnd.n629 240.244
R7066 gnd.n7620 gnd.n629 240.244
R7067 gnd.n7620 gnd.n627 240.244
R7068 gnd.n7624 gnd.n627 240.244
R7069 gnd.n7624 gnd.n623 240.244
R7070 gnd.n7630 gnd.n623 240.244
R7071 gnd.n7630 gnd.n621 240.244
R7072 gnd.n7634 gnd.n621 240.244
R7073 gnd.n7634 gnd.n617 240.244
R7074 gnd.n7640 gnd.n617 240.244
R7075 gnd.n7640 gnd.n615 240.244
R7076 gnd.n7644 gnd.n615 240.244
R7077 gnd.n7644 gnd.n611 240.244
R7078 gnd.n7650 gnd.n611 240.244
R7079 gnd.n7650 gnd.n609 240.244
R7080 gnd.n7654 gnd.n609 240.244
R7081 gnd.n7654 gnd.n605 240.244
R7082 gnd.n7660 gnd.n605 240.244
R7083 gnd.n7660 gnd.n603 240.244
R7084 gnd.n7664 gnd.n603 240.244
R7085 gnd.n7664 gnd.n599 240.244
R7086 gnd.n7670 gnd.n599 240.244
R7087 gnd.n7670 gnd.n597 240.244
R7088 gnd.n7674 gnd.n597 240.244
R7089 gnd.n7674 gnd.n593 240.244
R7090 gnd.n7680 gnd.n593 240.244
R7091 gnd.n7680 gnd.n591 240.244
R7092 gnd.n7684 gnd.n591 240.244
R7093 gnd.n7684 gnd.n587 240.244
R7094 gnd.n7690 gnd.n587 240.244
R7095 gnd.n7690 gnd.n585 240.244
R7096 gnd.n7694 gnd.n585 240.244
R7097 gnd.n7694 gnd.n581 240.244
R7098 gnd.n7700 gnd.n581 240.244
R7099 gnd.n7700 gnd.n579 240.244
R7100 gnd.n7704 gnd.n579 240.244
R7101 gnd.n7704 gnd.n575 240.244
R7102 gnd.n7710 gnd.n575 240.244
R7103 gnd.n7710 gnd.n573 240.244
R7104 gnd.n7715 gnd.n573 240.244
R7105 gnd.n7715 gnd.n569 240.244
R7106 gnd.n7722 gnd.n569 240.244
R7107 gnd.n2823 gnd.n2809 240.244
R7108 gnd.n2819 gnd.n2809 240.244
R7109 gnd.n2819 gnd.n2818 240.244
R7110 gnd.n2818 gnd.n2783 240.244
R7111 gnd.n3056 gnd.n2783 240.244
R7112 gnd.n3057 gnd.n3056 240.244
R7113 gnd.n3057 gnd.n2778 240.244
R7114 gnd.n3083 gnd.n2778 240.244
R7115 gnd.n3083 gnd.n2779 240.244
R7116 gnd.n3079 gnd.n2779 240.244
R7117 gnd.n3079 gnd.n3078 240.244
R7118 gnd.n3078 gnd.n3077 240.244
R7119 gnd.n3077 gnd.n3065 240.244
R7120 gnd.n3073 gnd.n3065 240.244
R7121 gnd.n3073 gnd.n2756 240.244
R7122 gnd.n3144 gnd.n2756 240.244
R7123 gnd.n3145 gnd.n3144 240.244
R7124 gnd.n3146 gnd.n3145 240.244
R7125 gnd.n3146 gnd.n2752 240.244
R7126 gnd.n3152 gnd.n2752 240.244
R7127 gnd.n3153 gnd.n3152 240.244
R7128 gnd.n3154 gnd.n3153 240.244
R7129 gnd.n3154 gnd.n2747 240.244
R7130 gnd.n3184 gnd.n2747 240.244
R7131 gnd.n3184 gnd.n2748 240.244
R7132 gnd.n3180 gnd.n2748 240.244
R7133 gnd.n3180 gnd.n3179 240.244
R7134 gnd.n3179 gnd.n3178 240.244
R7135 gnd.n3178 gnd.n3162 240.244
R7136 gnd.n3174 gnd.n3162 240.244
R7137 gnd.n3174 gnd.n3173 240.244
R7138 gnd.n3173 gnd.n3172 240.244
R7139 gnd.n3172 gnd.n2555 240.244
R7140 gnd.n3359 gnd.n2555 240.244
R7141 gnd.n3359 gnd.n2556 240.244
R7142 gnd.n3355 gnd.n2556 240.244
R7143 gnd.n3355 gnd.n3354 240.244
R7144 gnd.n3354 gnd.n2565 240.244
R7145 gnd.n2565 gnd.n2541 240.244
R7146 gnd.n3374 gnd.n2541 240.244
R7147 gnd.n3374 gnd.n2537 240.244
R7148 gnd.n3380 gnd.n2537 240.244
R7149 gnd.n3380 gnd.n2528 240.244
R7150 gnd.n3390 gnd.n2528 240.244
R7151 gnd.n3390 gnd.n2524 240.244
R7152 gnd.n3396 gnd.n2524 240.244
R7153 gnd.n3396 gnd.n2514 240.244
R7154 gnd.n3406 gnd.n2514 240.244
R7155 gnd.n3406 gnd.n2510 240.244
R7156 gnd.n3412 gnd.n2510 240.244
R7157 gnd.n3412 gnd.n2500 240.244
R7158 gnd.n3422 gnd.n2500 240.244
R7159 gnd.n3422 gnd.n2495 240.244
R7160 gnd.n3437 gnd.n2495 240.244
R7161 gnd.n3437 gnd.n2496 240.244
R7162 gnd.n3433 gnd.n2496 240.244
R7163 gnd.n3433 gnd.n3432 240.244
R7164 gnd.n3432 gnd.n1693 240.244
R7165 gnd.n4973 gnd.n1693 240.244
R7166 gnd.n4973 gnd.n1694 240.244
R7167 gnd.n4969 gnd.n1694 240.244
R7168 gnd.n4969 gnd.n1700 240.244
R7169 gnd.n4090 gnd.n1700 240.244
R7170 gnd.n4090 gnd.n2384 240.244
R7171 gnd.n4100 gnd.n2384 240.244
R7172 gnd.n4100 gnd.n2380 240.244
R7173 gnd.n4106 gnd.n2380 240.244
R7174 gnd.n4106 gnd.n2370 240.244
R7175 gnd.n4116 gnd.n2370 240.244
R7176 gnd.n4116 gnd.n2366 240.244
R7177 gnd.n4122 gnd.n2366 240.244
R7178 gnd.n4122 gnd.n2358 240.244
R7179 gnd.n4132 gnd.n2358 240.244
R7180 gnd.n4132 gnd.n2354 240.244
R7181 gnd.n4138 gnd.n2354 240.244
R7182 gnd.n4138 gnd.n2344 240.244
R7183 gnd.n4148 gnd.n2344 240.244
R7184 gnd.n4148 gnd.n2340 240.244
R7185 gnd.n4154 gnd.n2340 240.244
R7186 gnd.n4154 gnd.n2329 240.244
R7187 gnd.n4164 gnd.n2329 240.244
R7188 gnd.n4164 gnd.n2325 240.244
R7189 gnd.n4170 gnd.n2325 240.244
R7190 gnd.n4170 gnd.n2315 240.244
R7191 gnd.n4180 gnd.n2315 240.244
R7192 gnd.n4180 gnd.n2311 240.244
R7193 gnd.n4186 gnd.n2311 240.244
R7194 gnd.n4186 gnd.n2301 240.244
R7195 gnd.n4196 gnd.n2301 240.244
R7196 gnd.n4196 gnd.n2297 240.244
R7197 gnd.n4202 gnd.n2297 240.244
R7198 gnd.n4202 gnd.n2288 240.244
R7199 gnd.n4212 gnd.n2288 240.244
R7200 gnd.n4212 gnd.n2284 240.244
R7201 gnd.n4218 gnd.n2284 240.244
R7202 gnd.n4218 gnd.n2274 240.244
R7203 gnd.n4228 gnd.n2274 240.244
R7204 gnd.n4228 gnd.n2270 240.244
R7205 gnd.n4234 gnd.n2270 240.244
R7206 gnd.n4234 gnd.n2260 240.244
R7207 gnd.n4244 gnd.n2260 240.244
R7208 gnd.n4244 gnd.n2256 240.244
R7209 gnd.n4250 gnd.n2256 240.244
R7210 gnd.n4250 gnd.n2247 240.244
R7211 gnd.n4260 gnd.n2247 240.244
R7212 gnd.n4260 gnd.n2243 240.244
R7213 gnd.n4266 gnd.n2243 240.244
R7214 gnd.n4266 gnd.n2233 240.244
R7215 gnd.n4276 gnd.n2233 240.244
R7216 gnd.n4276 gnd.n2229 240.244
R7217 gnd.n4282 gnd.n2229 240.244
R7218 gnd.n4282 gnd.n2220 240.244
R7219 gnd.n4292 gnd.n2220 240.244
R7220 gnd.n4292 gnd.n2216 240.244
R7221 gnd.n4298 gnd.n2216 240.244
R7222 gnd.n4298 gnd.n2205 240.244
R7223 gnd.n4308 gnd.n2205 240.244
R7224 gnd.n4308 gnd.n2201 240.244
R7225 gnd.n4314 gnd.n2201 240.244
R7226 gnd.n4314 gnd.n2192 240.244
R7227 gnd.n4324 gnd.n2192 240.244
R7228 gnd.n4324 gnd.n2188 240.244
R7229 gnd.n4330 gnd.n2188 240.244
R7230 gnd.n4330 gnd.n2181 240.244
R7231 gnd.n4340 gnd.n2181 240.244
R7232 gnd.n4340 gnd.n2177 240.244
R7233 gnd.n4346 gnd.n2177 240.244
R7234 gnd.n4346 gnd.n2168 240.244
R7235 gnd.n4356 gnd.n2168 240.244
R7236 gnd.n4356 gnd.n2164 240.244
R7237 gnd.n4362 gnd.n2164 240.244
R7238 gnd.n4362 gnd.n2153 240.244
R7239 gnd.n4372 gnd.n2153 240.244
R7240 gnd.n4372 gnd.n2149 240.244
R7241 gnd.n4378 gnd.n2149 240.244
R7242 gnd.n4378 gnd.n2141 240.244
R7243 gnd.n4390 gnd.n2141 240.244
R7244 gnd.n4390 gnd.n2136 240.244
R7245 gnd.n4399 gnd.n2136 240.244
R7246 gnd.n4399 gnd.n2137 240.244
R7247 gnd.n2137 gnd.n1810 240.244
R7248 gnd.n4843 gnd.n1810 240.244
R7249 gnd.n4843 gnd.n1813 240.244
R7250 gnd.n4839 gnd.n1813 240.244
R7251 gnd.n4839 gnd.n1819 240.244
R7252 gnd.n2077 gnd.n1819 240.244
R7253 gnd.n2078 gnd.n2077 240.244
R7254 gnd.n2078 gnd.n2072 240.244
R7255 gnd.n2084 gnd.n2072 240.244
R7256 gnd.n2085 gnd.n2084 240.244
R7257 gnd.n2086 gnd.n2085 240.244
R7258 gnd.n2086 gnd.n2068 240.244
R7259 gnd.n2092 gnd.n2068 240.244
R7260 gnd.n2093 gnd.n2092 240.244
R7261 gnd.n2094 gnd.n2093 240.244
R7262 gnd.n2094 gnd.n2063 240.244
R7263 gnd.n2119 gnd.n2063 240.244
R7264 gnd.n2119 gnd.n2064 240.244
R7265 gnd.n2115 gnd.n2064 240.244
R7266 gnd.n2115 gnd.n2114 240.244
R7267 gnd.n2114 gnd.n2113 240.244
R7268 gnd.n2113 gnd.n2102 240.244
R7269 gnd.n2109 gnd.n2102 240.244
R7270 gnd.n2109 gnd.n2050 240.244
R7271 gnd.n4642 gnd.n2050 240.244
R7272 gnd.n4643 gnd.n4642 240.244
R7273 gnd.n4643 gnd.n2046 240.244
R7274 gnd.n4650 gnd.n2046 240.244
R7275 gnd.n4650 gnd.n551 240.244
R7276 gnd.n7742 gnd.n551 240.244
R7277 gnd.n7742 gnd.n552 240.244
R7278 gnd.n7738 gnd.n552 240.244
R7279 gnd.n7738 gnd.n7737 240.244
R7280 gnd.n7737 gnd.n7736 240.244
R7281 gnd.n7736 gnd.n558 240.244
R7282 gnd.n564 gnd.n558 240.244
R7283 gnd.n7729 gnd.n564 240.244
R7284 gnd.n7729 gnd.n7728 240.244
R7285 gnd.n7728 gnd.n7727 240.244
R7286 gnd.n7727 gnd.n565 240.244
R7287 gnd.n7723 gnd.n565 240.244
R7288 gnd.n7049 gnd.n967 240.244
R7289 gnd.n7049 gnd.n969 240.244
R7290 gnd.n7045 gnd.n969 240.244
R7291 gnd.n7045 gnd.n975 240.244
R7292 gnd.n7041 gnd.n975 240.244
R7293 gnd.n7041 gnd.n977 240.244
R7294 gnd.n7037 gnd.n977 240.244
R7295 gnd.n7037 gnd.n983 240.244
R7296 gnd.n7033 gnd.n983 240.244
R7297 gnd.n7033 gnd.n985 240.244
R7298 gnd.n7029 gnd.n985 240.244
R7299 gnd.n7029 gnd.n991 240.244
R7300 gnd.n7025 gnd.n991 240.244
R7301 gnd.n7025 gnd.n993 240.244
R7302 gnd.n7021 gnd.n993 240.244
R7303 gnd.n7021 gnd.n999 240.244
R7304 gnd.n7017 gnd.n999 240.244
R7305 gnd.n7017 gnd.n1001 240.244
R7306 gnd.n7013 gnd.n1001 240.244
R7307 gnd.n7013 gnd.n1007 240.244
R7308 gnd.n7009 gnd.n1007 240.244
R7309 gnd.n7009 gnd.n1009 240.244
R7310 gnd.n7005 gnd.n1009 240.244
R7311 gnd.n7005 gnd.n1015 240.244
R7312 gnd.n7001 gnd.n1015 240.244
R7313 gnd.n7001 gnd.n1017 240.244
R7314 gnd.n6997 gnd.n1017 240.244
R7315 gnd.n6997 gnd.n1023 240.244
R7316 gnd.n6993 gnd.n1023 240.244
R7317 gnd.n6993 gnd.n1025 240.244
R7318 gnd.n6989 gnd.n1025 240.244
R7319 gnd.n6989 gnd.n1031 240.244
R7320 gnd.n6985 gnd.n1031 240.244
R7321 gnd.n6985 gnd.n1033 240.244
R7322 gnd.n6981 gnd.n1033 240.244
R7323 gnd.n6981 gnd.n1039 240.244
R7324 gnd.n6977 gnd.n1039 240.244
R7325 gnd.n6977 gnd.n1041 240.244
R7326 gnd.n6973 gnd.n1041 240.244
R7327 gnd.n6973 gnd.n1047 240.244
R7328 gnd.n6969 gnd.n1047 240.244
R7329 gnd.n6969 gnd.n1049 240.244
R7330 gnd.n6965 gnd.n1049 240.244
R7331 gnd.n6965 gnd.n1055 240.244
R7332 gnd.n6961 gnd.n1055 240.244
R7333 gnd.n6961 gnd.n1057 240.244
R7334 gnd.n6957 gnd.n1057 240.244
R7335 gnd.n6957 gnd.n1063 240.244
R7336 gnd.n6953 gnd.n1063 240.244
R7337 gnd.n6953 gnd.n1065 240.244
R7338 gnd.n6949 gnd.n1065 240.244
R7339 gnd.n6949 gnd.n1071 240.244
R7340 gnd.n6945 gnd.n1071 240.244
R7341 gnd.n6945 gnd.n1073 240.244
R7342 gnd.n6941 gnd.n1073 240.244
R7343 gnd.n6941 gnd.n1079 240.244
R7344 gnd.n6937 gnd.n1079 240.244
R7345 gnd.n6937 gnd.n1081 240.244
R7346 gnd.n6933 gnd.n1081 240.244
R7347 gnd.n6933 gnd.n1087 240.244
R7348 gnd.n6929 gnd.n1087 240.244
R7349 gnd.n6929 gnd.n1089 240.244
R7350 gnd.n6925 gnd.n1089 240.244
R7351 gnd.n6925 gnd.n1095 240.244
R7352 gnd.n6921 gnd.n1095 240.244
R7353 gnd.n6921 gnd.n1097 240.244
R7354 gnd.n6917 gnd.n1097 240.244
R7355 gnd.n6917 gnd.n1103 240.244
R7356 gnd.n6913 gnd.n1103 240.244
R7357 gnd.n6913 gnd.n1105 240.244
R7358 gnd.n6909 gnd.n1105 240.244
R7359 gnd.n6909 gnd.n1111 240.244
R7360 gnd.n6905 gnd.n1111 240.244
R7361 gnd.n6905 gnd.n1113 240.244
R7362 gnd.n6901 gnd.n1113 240.244
R7363 gnd.n6901 gnd.n1119 240.244
R7364 gnd.n6897 gnd.n1119 240.244
R7365 gnd.n6897 gnd.n1121 240.244
R7366 gnd.n6893 gnd.n1121 240.244
R7367 gnd.n6893 gnd.n1127 240.244
R7368 gnd.n6889 gnd.n1127 240.244
R7369 gnd.n6889 gnd.n1129 240.244
R7370 gnd.n6885 gnd.n1129 240.244
R7371 gnd.n6885 gnd.n1135 240.244
R7372 gnd.n2583 gnd.n2543 240.244
R7373 gnd.n2583 gnd.n2536 240.244
R7374 gnd.n2584 gnd.n2536 240.244
R7375 gnd.n2584 gnd.n2530 240.244
R7376 gnd.n2587 gnd.n2530 240.244
R7377 gnd.n2587 gnd.n2523 240.244
R7378 gnd.n2588 gnd.n2523 240.244
R7379 gnd.n2588 gnd.n2516 240.244
R7380 gnd.n2591 gnd.n2516 240.244
R7381 gnd.n2591 gnd.n2508 240.244
R7382 gnd.n2592 gnd.n2508 240.244
R7383 gnd.n2592 gnd.n2501 240.244
R7384 gnd.n2595 gnd.n2501 240.244
R7385 gnd.n2595 gnd.n2493 240.244
R7386 gnd.n2598 gnd.n2493 240.244
R7387 gnd.n2599 gnd.n2598 240.244
R7388 gnd.n2600 gnd.n2599 240.244
R7389 gnd.n2601 gnd.n2600 240.244
R7390 gnd.n2601 gnd.n1690 240.244
R7391 gnd.n1704 gnd.n1690 240.244
R7392 gnd.n4968 gnd.n1704 240.244
R7393 gnd.n4968 gnd.n1705 240.244
R7394 gnd.n1710 gnd.n1705 240.244
R7395 gnd.n1711 gnd.n1710 240.244
R7396 gnd.n1712 gnd.n1711 240.244
R7397 gnd.n2400 gnd.n1712 240.244
R7398 gnd.n2400 gnd.n1715 240.244
R7399 gnd.n1716 gnd.n1715 240.244
R7400 gnd.n1717 gnd.n1716 240.244
R7401 gnd.n3485 gnd.n1717 240.244
R7402 gnd.n3485 gnd.n1720 240.244
R7403 gnd.n1721 gnd.n1720 240.244
R7404 gnd.n1722 gnd.n1721 240.244
R7405 gnd.n3503 gnd.n1722 240.244
R7406 gnd.n3503 gnd.n1725 240.244
R7407 gnd.n1726 gnd.n1725 240.244
R7408 gnd.n1727 gnd.n1726 240.244
R7409 gnd.n3516 gnd.n1727 240.244
R7410 gnd.n3516 gnd.n1730 240.244
R7411 gnd.n1731 gnd.n1730 240.244
R7412 gnd.n1732 gnd.n1731 240.244
R7413 gnd.n2331 gnd.n1732 240.244
R7414 gnd.n2331 gnd.n1735 240.244
R7415 gnd.n1736 gnd.n1735 240.244
R7416 gnd.n1737 gnd.n1736 240.244
R7417 gnd.n4011 gnd.n1737 240.244
R7418 gnd.n4011 gnd.n1740 240.244
R7419 gnd.n1741 gnd.n1740 240.244
R7420 gnd.n1742 gnd.n1741 240.244
R7421 gnd.n3995 gnd.n1742 240.244
R7422 gnd.n3995 gnd.n1745 240.244
R7423 gnd.n1746 gnd.n1745 240.244
R7424 gnd.n1747 gnd.n1746 240.244
R7425 gnd.n3979 gnd.n1747 240.244
R7426 gnd.n3979 gnd.n1750 240.244
R7427 gnd.n1751 gnd.n1750 240.244
R7428 gnd.n1752 gnd.n1751 240.244
R7429 gnd.n3963 gnd.n1752 240.244
R7430 gnd.n3963 gnd.n1755 240.244
R7431 gnd.n1756 gnd.n1755 240.244
R7432 gnd.n1757 gnd.n1756 240.244
R7433 gnd.n3600 gnd.n1757 240.244
R7434 gnd.n3600 gnd.n1760 240.244
R7435 gnd.n1761 gnd.n1760 240.244
R7436 gnd.n1762 gnd.n1761 240.244
R7437 gnd.n3616 gnd.n1762 240.244
R7438 gnd.n3616 gnd.n1765 240.244
R7439 gnd.n1766 gnd.n1765 240.244
R7440 gnd.n1767 gnd.n1766 240.244
R7441 gnd.n3630 gnd.n1767 240.244
R7442 gnd.n3630 gnd.n1770 240.244
R7443 gnd.n1771 gnd.n1770 240.244
R7444 gnd.n1772 gnd.n1771 240.244
R7445 gnd.n3645 gnd.n1772 240.244
R7446 gnd.n3645 gnd.n1775 240.244
R7447 gnd.n1776 gnd.n1775 240.244
R7448 gnd.n1777 gnd.n1776 240.244
R7449 gnd.n3669 gnd.n1777 240.244
R7450 gnd.n3669 gnd.n1780 240.244
R7451 gnd.n1781 gnd.n1780 240.244
R7452 gnd.n1782 gnd.n1781 240.244
R7453 gnd.n3679 gnd.n1782 240.244
R7454 gnd.n3679 gnd.n1785 240.244
R7455 gnd.n1786 gnd.n1785 240.244
R7456 gnd.n1787 gnd.n1786 240.244
R7457 gnd.n2175 gnd.n1787 240.244
R7458 gnd.n2175 gnd.n1790 240.244
R7459 gnd.n1791 gnd.n1790 240.244
R7460 gnd.n1792 gnd.n1791 240.244
R7461 gnd.n2162 gnd.n1792 240.244
R7462 gnd.n2162 gnd.n1795 240.244
R7463 gnd.n1796 gnd.n1795 240.244
R7464 gnd.n1797 gnd.n1796 240.244
R7465 gnd.n2155 gnd.n1797 240.244
R7466 gnd.n2155 gnd.n1800 240.244
R7467 gnd.n1801 gnd.n1800 240.244
R7468 gnd.n1802 gnd.n1801 240.244
R7469 gnd.n2134 gnd.n1802 240.244
R7470 gnd.n2134 gnd.n1805 240.244
R7471 gnd.n1806 gnd.n1805 240.244
R7472 gnd.n4846 gnd.n1806 240.244
R7473 gnd.n2581 gnd.n2580 240.244
R7474 gnd.n2636 gnd.n2580 240.244
R7475 gnd.n2638 gnd.n2637 240.244
R7476 gnd.n3227 gnd.n3226 240.244
R7477 gnd.n3229 gnd.n3228 240.244
R7478 gnd.n3240 gnd.n3239 240.244
R7479 gnd.n3242 gnd.n3241 240.244
R7480 gnd.n3250 gnd.n3249 240.244
R7481 gnd.n3260 gnd.n3259 240.244
R7482 gnd.n3262 gnd.n3261 240.244
R7483 gnd.n3270 gnd.n3269 240.244
R7484 gnd.n3280 gnd.n3279 240.244
R7485 gnd.n3286 gnd.n3281 240.244
R7486 gnd.n2577 gnd.n2548 240.244
R7487 gnd.n3372 gnd.n2535 240.244
R7488 gnd.n3382 gnd.n2535 240.244
R7489 gnd.n3382 gnd.n2531 240.244
R7490 gnd.n3388 gnd.n2531 240.244
R7491 gnd.n3388 gnd.n2521 240.244
R7492 gnd.n3398 gnd.n2521 240.244
R7493 gnd.n3398 gnd.n2517 240.244
R7494 gnd.n3404 gnd.n2517 240.244
R7495 gnd.n3404 gnd.n2506 240.244
R7496 gnd.n3414 gnd.n2506 240.244
R7497 gnd.n3414 gnd.n2502 240.244
R7498 gnd.n3420 gnd.n2502 240.244
R7499 gnd.n3420 gnd.n2491 240.244
R7500 gnd.n3439 gnd.n2491 240.244
R7501 gnd.n3439 gnd.n2487 240.244
R7502 gnd.n3445 gnd.n2487 240.244
R7503 gnd.n3446 gnd.n3445 240.244
R7504 gnd.n3447 gnd.n3446 240.244
R7505 gnd.n3447 gnd.n1692 240.244
R7506 gnd.n3454 gnd.n1692 240.244
R7507 gnd.n3454 gnd.n1702 240.244
R7508 gnd.n2390 gnd.n1702 240.244
R7509 gnd.n4092 gnd.n2390 240.244
R7510 gnd.n4092 gnd.n2386 240.244
R7511 gnd.n4098 gnd.n2386 240.244
R7512 gnd.n4098 gnd.n2377 240.244
R7513 gnd.n4108 gnd.n2377 240.244
R7514 gnd.n4108 gnd.n2373 240.244
R7515 gnd.n4114 gnd.n2373 240.244
R7516 gnd.n4114 gnd.n2364 240.244
R7517 gnd.n4124 gnd.n2364 240.244
R7518 gnd.n4124 gnd.n2360 240.244
R7519 gnd.n4130 gnd.n2360 240.244
R7520 gnd.n4130 gnd.n2351 240.244
R7521 gnd.n4140 gnd.n2351 240.244
R7522 gnd.n4140 gnd.n2347 240.244
R7523 gnd.n4146 gnd.n2347 240.244
R7524 gnd.n4146 gnd.n2338 240.244
R7525 gnd.n4156 gnd.n2338 240.244
R7526 gnd.n4156 gnd.n2334 240.244
R7527 gnd.n4162 gnd.n2334 240.244
R7528 gnd.n4162 gnd.n2322 240.244
R7529 gnd.n4172 gnd.n2322 240.244
R7530 gnd.n4172 gnd.n2318 240.244
R7531 gnd.n4178 gnd.n2318 240.244
R7532 gnd.n4178 gnd.n2308 240.244
R7533 gnd.n4188 gnd.n2308 240.244
R7534 gnd.n4188 gnd.n2304 240.244
R7535 gnd.n4194 gnd.n2304 240.244
R7536 gnd.n4194 gnd.n2294 240.244
R7537 gnd.n4204 gnd.n2294 240.244
R7538 gnd.n4204 gnd.n2290 240.244
R7539 gnd.n4210 gnd.n2290 240.244
R7540 gnd.n4210 gnd.n2281 240.244
R7541 gnd.n4220 gnd.n2281 240.244
R7542 gnd.n4220 gnd.n2277 240.244
R7543 gnd.n4226 gnd.n2277 240.244
R7544 gnd.n4226 gnd.n2267 240.244
R7545 gnd.n4236 gnd.n2267 240.244
R7546 gnd.n4236 gnd.n2263 240.244
R7547 gnd.n4242 gnd.n2263 240.244
R7548 gnd.n4242 gnd.n2253 240.244
R7549 gnd.n4252 gnd.n2253 240.244
R7550 gnd.n4252 gnd.n2249 240.244
R7551 gnd.n4258 gnd.n2249 240.244
R7552 gnd.n4258 gnd.n2240 240.244
R7553 gnd.n4268 gnd.n2240 240.244
R7554 gnd.n4268 gnd.n2236 240.244
R7555 gnd.n4274 gnd.n2236 240.244
R7556 gnd.n4274 gnd.n2227 240.244
R7557 gnd.n4284 gnd.n2227 240.244
R7558 gnd.n4284 gnd.n2223 240.244
R7559 gnd.n4290 gnd.n2223 240.244
R7560 gnd.n4290 gnd.n2212 240.244
R7561 gnd.n4300 gnd.n2212 240.244
R7562 gnd.n4300 gnd.n2208 240.244
R7563 gnd.n4306 gnd.n2208 240.244
R7564 gnd.n4306 gnd.n2198 240.244
R7565 gnd.n4316 gnd.n2198 240.244
R7566 gnd.n4316 gnd.n2194 240.244
R7567 gnd.n4322 gnd.n2194 240.244
R7568 gnd.n4322 gnd.n2186 240.244
R7569 gnd.n4332 gnd.n2186 240.244
R7570 gnd.n4332 gnd.n2182 240.244
R7571 gnd.n4338 gnd.n2182 240.244
R7572 gnd.n4338 gnd.n2174 240.244
R7573 gnd.n4348 gnd.n2174 240.244
R7574 gnd.n4348 gnd.n2170 240.244
R7575 gnd.n4354 gnd.n2170 240.244
R7576 gnd.n4354 gnd.n2161 240.244
R7577 gnd.n4364 gnd.n2161 240.244
R7578 gnd.n4364 gnd.n2157 240.244
R7579 gnd.n4370 gnd.n2157 240.244
R7580 gnd.n4370 gnd.n2148 240.244
R7581 gnd.n4380 gnd.n2148 240.244
R7582 gnd.n4380 gnd.n2143 240.244
R7583 gnd.n4388 gnd.n2143 240.244
R7584 gnd.n4388 gnd.n2133 240.244
R7585 gnd.n4401 gnd.n2133 240.244
R7586 gnd.n4402 gnd.n4401 240.244
R7587 gnd.n4402 gnd.n1811 240.244
R7588 gnd.n4457 gnd.n4456 240.244
R7589 gnd.n4460 gnd.n4459 240.244
R7590 gnd.n4468 gnd.n4467 240.244
R7591 gnd.n4471 gnd.n4470 240.244
R7592 gnd.n4485 gnd.n4484 240.244
R7593 gnd.n4488 gnd.n4487 240.244
R7594 gnd.n4504 gnd.n4503 240.244
R7595 gnd.n4507 gnd.n4506 240.244
R7596 gnd.n4523 gnd.n4522 240.244
R7597 gnd.n4526 gnd.n4525 240.244
R7598 gnd.n4542 gnd.n4541 240.244
R7599 gnd.n4544 gnd.n4409 240.244
R7600 gnd.n4557 gnd.n4409 240.244
R7601 gnd.n4560 gnd.n4559 240.244
R7602 gnd.n1672 gnd.n1671 240.132
R7603 gnd.n3717 gnd.n3716 240.132
R7604 gnd.n7052 gnd.n963 225.874
R7605 gnd.n7060 gnd.n963 225.874
R7606 gnd.n7061 gnd.n7060 225.874
R7607 gnd.n7062 gnd.n7061 225.874
R7608 gnd.n7062 gnd.n957 225.874
R7609 gnd.n7070 gnd.n957 225.874
R7610 gnd.n7071 gnd.n7070 225.874
R7611 gnd.n7072 gnd.n7071 225.874
R7612 gnd.n7072 gnd.n951 225.874
R7613 gnd.n7080 gnd.n951 225.874
R7614 gnd.n7081 gnd.n7080 225.874
R7615 gnd.n7082 gnd.n7081 225.874
R7616 gnd.n7082 gnd.n945 225.874
R7617 gnd.n7090 gnd.n945 225.874
R7618 gnd.n7091 gnd.n7090 225.874
R7619 gnd.n7092 gnd.n7091 225.874
R7620 gnd.n7092 gnd.n939 225.874
R7621 gnd.n7100 gnd.n939 225.874
R7622 gnd.n7101 gnd.n7100 225.874
R7623 gnd.n7102 gnd.n7101 225.874
R7624 gnd.n7102 gnd.n933 225.874
R7625 gnd.n7110 gnd.n933 225.874
R7626 gnd.n7111 gnd.n7110 225.874
R7627 gnd.n7112 gnd.n7111 225.874
R7628 gnd.n7112 gnd.n927 225.874
R7629 gnd.n7120 gnd.n927 225.874
R7630 gnd.n7121 gnd.n7120 225.874
R7631 gnd.n7122 gnd.n7121 225.874
R7632 gnd.n7122 gnd.n921 225.874
R7633 gnd.n7130 gnd.n921 225.874
R7634 gnd.n7131 gnd.n7130 225.874
R7635 gnd.n7132 gnd.n7131 225.874
R7636 gnd.n7132 gnd.n915 225.874
R7637 gnd.n7140 gnd.n915 225.874
R7638 gnd.n7141 gnd.n7140 225.874
R7639 gnd.n7142 gnd.n7141 225.874
R7640 gnd.n7142 gnd.n909 225.874
R7641 gnd.n7150 gnd.n909 225.874
R7642 gnd.n7151 gnd.n7150 225.874
R7643 gnd.n7152 gnd.n7151 225.874
R7644 gnd.n7152 gnd.n903 225.874
R7645 gnd.n7160 gnd.n903 225.874
R7646 gnd.n7161 gnd.n7160 225.874
R7647 gnd.n7162 gnd.n7161 225.874
R7648 gnd.n7162 gnd.n897 225.874
R7649 gnd.n7170 gnd.n897 225.874
R7650 gnd.n7171 gnd.n7170 225.874
R7651 gnd.n7172 gnd.n7171 225.874
R7652 gnd.n7172 gnd.n891 225.874
R7653 gnd.n7180 gnd.n891 225.874
R7654 gnd.n7181 gnd.n7180 225.874
R7655 gnd.n7182 gnd.n7181 225.874
R7656 gnd.n7182 gnd.n885 225.874
R7657 gnd.n7190 gnd.n885 225.874
R7658 gnd.n7191 gnd.n7190 225.874
R7659 gnd.n7192 gnd.n7191 225.874
R7660 gnd.n7192 gnd.n879 225.874
R7661 gnd.n7200 gnd.n879 225.874
R7662 gnd.n7201 gnd.n7200 225.874
R7663 gnd.n7202 gnd.n7201 225.874
R7664 gnd.n7202 gnd.n873 225.874
R7665 gnd.n7210 gnd.n873 225.874
R7666 gnd.n7211 gnd.n7210 225.874
R7667 gnd.n7212 gnd.n7211 225.874
R7668 gnd.n7212 gnd.n867 225.874
R7669 gnd.n7220 gnd.n867 225.874
R7670 gnd.n7221 gnd.n7220 225.874
R7671 gnd.n7222 gnd.n7221 225.874
R7672 gnd.n7222 gnd.n861 225.874
R7673 gnd.n7230 gnd.n861 225.874
R7674 gnd.n7231 gnd.n7230 225.874
R7675 gnd.n7232 gnd.n7231 225.874
R7676 gnd.n7232 gnd.n855 225.874
R7677 gnd.n7240 gnd.n855 225.874
R7678 gnd.n7241 gnd.n7240 225.874
R7679 gnd.n7242 gnd.n7241 225.874
R7680 gnd.n7242 gnd.n849 225.874
R7681 gnd.n7250 gnd.n849 225.874
R7682 gnd.n7251 gnd.n7250 225.874
R7683 gnd.n7252 gnd.n7251 225.874
R7684 gnd.n7252 gnd.n843 225.874
R7685 gnd.n7260 gnd.n843 225.874
R7686 gnd.n7261 gnd.n7260 225.874
R7687 gnd.n7262 gnd.n7261 225.874
R7688 gnd.n7262 gnd.n837 225.874
R7689 gnd.n7270 gnd.n837 225.874
R7690 gnd.n7271 gnd.n7270 225.874
R7691 gnd.n7272 gnd.n7271 225.874
R7692 gnd.n7272 gnd.n831 225.874
R7693 gnd.n7280 gnd.n831 225.874
R7694 gnd.n7281 gnd.n7280 225.874
R7695 gnd.n7282 gnd.n7281 225.874
R7696 gnd.n7282 gnd.n825 225.874
R7697 gnd.n7290 gnd.n825 225.874
R7698 gnd.n7291 gnd.n7290 225.874
R7699 gnd.n7292 gnd.n7291 225.874
R7700 gnd.n7292 gnd.n819 225.874
R7701 gnd.n7300 gnd.n819 225.874
R7702 gnd.n7301 gnd.n7300 225.874
R7703 gnd.n7302 gnd.n7301 225.874
R7704 gnd.n7302 gnd.n813 225.874
R7705 gnd.n7310 gnd.n813 225.874
R7706 gnd.n7311 gnd.n7310 225.874
R7707 gnd.n7312 gnd.n7311 225.874
R7708 gnd.n7312 gnd.n807 225.874
R7709 gnd.n7320 gnd.n807 225.874
R7710 gnd.n7321 gnd.n7320 225.874
R7711 gnd.n7322 gnd.n7321 225.874
R7712 gnd.n7322 gnd.n801 225.874
R7713 gnd.n7330 gnd.n801 225.874
R7714 gnd.n7331 gnd.n7330 225.874
R7715 gnd.n7332 gnd.n7331 225.874
R7716 gnd.n7332 gnd.n795 225.874
R7717 gnd.n7340 gnd.n795 225.874
R7718 gnd.n7341 gnd.n7340 225.874
R7719 gnd.n7342 gnd.n7341 225.874
R7720 gnd.n7342 gnd.n789 225.874
R7721 gnd.n7350 gnd.n789 225.874
R7722 gnd.n7351 gnd.n7350 225.874
R7723 gnd.n7352 gnd.n7351 225.874
R7724 gnd.n7352 gnd.n783 225.874
R7725 gnd.n7360 gnd.n783 225.874
R7726 gnd.n7361 gnd.n7360 225.874
R7727 gnd.n7362 gnd.n7361 225.874
R7728 gnd.n7362 gnd.n777 225.874
R7729 gnd.n7370 gnd.n777 225.874
R7730 gnd.n7371 gnd.n7370 225.874
R7731 gnd.n7372 gnd.n7371 225.874
R7732 gnd.n7372 gnd.n771 225.874
R7733 gnd.n7380 gnd.n771 225.874
R7734 gnd.n7381 gnd.n7380 225.874
R7735 gnd.n7382 gnd.n7381 225.874
R7736 gnd.n7382 gnd.n765 225.874
R7737 gnd.n7390 gnd.n765 225.874
R7738 gnd.n7391 gnd.n7390 225.874
R7739 gnd.n7392 gnd.n7391 225.874
R7740 gnd.n7392 gnd.n759 225.874
R7741 gnd.n7400 gnd.n759 225.874
R7742 gnd.n7401 gnd.n7400 225.874
R7743 gnd.n7402 gnd.n7401 225.874
R7744 gnd.n7402 gnd.n753 225.874
R7745 gnd.n7410 gnd.n753 225.874
R7746 gnd.n7411 gnd.n7410 225.874
R7747 gnd.n7412 gnd.n7411 225.874
R7748 gnd.n7412 gnd.n747 225.874
R7749 gnd.n7420 gnd.n747 225.874
R7750 gnd.n7421 gnd.n7420 225.874
R7751 gnd.n7422 gnd.n7421 225.874
R7752 gnd.n7422 gnd.n741 225.874
R7753 gnd.n7430 gnd.n741 225.874
R7754 gnd.n7431 gnd.n7430 225.874
R7755 gnd.n7432 gnd.n7431 225.874
R7756 gnd.n7432 gnd.n735 225.874
R7757 gnd.n7440 gnd.n735 225.874
R7758 gnd.n7441 gnd.n7440 225.874
R7759 gnd.n7442 gnd.n7441 225.874
R7760 gnd.n7442 gnd.n729 225.874
R7761 gnd.n7450 gnd.n729 225.874
R7762 gnd.n7451 gnd.n7450 225.874
R7763 gnd.n7452 gnd.n7451 225.874
R7764 gnd.n7452 gnd.n723 225.874
R7765 gnd.n7460 gnd.n723 225.874
R7766 gnd.n7461 gnd.n7460 225.874
R7767 gnd.n7462 gnd.n7461 225.874
R7768 gnd.n7462 gnd.n717 225.874
R7769 gnd.n7470 gnd.n717 225.874
R7770 gnd.n7471 gnd.n7470 225.874
R7771 gnd.n7472 gnd.n7471 225.874
R7772 gnd.n7472 gnd.n711 225.874
R7773 gnd.n7480 gnd.n711 225.874
R7774 gnd.n7481 gnd.n7480 225.874
R7775 gnd.n7482 gnd.n7481 225.874
R7776 gnd.n7482 gnd.n705 225.874
R7777 gnd.n7490 gnd.n705 225.874
R7778 gnd.n7491 gnd.n7490 225.874
R7779 gnd.n7492 gnd.n7491 225.874
R7780 gnd.n7492 gnd.n699 225.874
R7781 gnd.n7501 gnd.n699 225.874
R7782 gnd.n7502 gnd.n7501 225.874
R7783 gnd.n7503 gnd.n7502 225.874
R7784 gnd.n7503 gnd.n694 225.874
R7785 gnd.n6093 gnd.t60 224.174
R7786 gnd.n5474 gnd.t172 224.174
R7787 gnd.n1892 gnd.n1832 199.319
R7788 gnd.n1892 gnd.n1833 199.319
R7789 gnd.n1624 gnd.n1584 199.319
R7790 gnd.n1624 gnd.n1583 199.319
R7791 gnd.n1673 gnd.n1670 186.49
R7792 gnd.n3718 gnd.n3715 186.49
R7793 gnd.n5742 gnd.n5741 185
R7794 gnd.n5740 gnd.n5739 185
R7795 gnd.n5719 gnd.n5718 185
R7796 gnd.n5734 gnd.n5733 185
R7797 gnd.n5732 gnd.n5731 185
R7798 gnd.n5723 gnd.n5722 185
R7799 gnd.n5726 gnd.n5725 185
R7800 gnd.n5710 gnd.n5709 185
R7801 gnd.n5708 gnd.n5707 185
R7802 gnd.n5687 gnd.n5686 185
R7803 gnd.n5702 gnd.n5701 185
R7804 gnd.n5700 gnd.n5699 185
R7805 gnd.n5691 gnd.n5690 185
R7806 gnd.n5694 gnd.n5693 185
R7807 gnd.n5678 gnd.n5677 185
R7808 gnd.n5676 gnd.n5675 185
R7809 gnd.n5655 gnd.n5654 185
R7810 gnd.n5670 gnd.n5669 185
R7811 gnd.n5668 gnd.n5667 185
R7812 gnd.n5659 gnd.n5658 185
R7813 gnd.n5662 gnd.n5661 185
R7814 gnd.n5647 gnd.n5646 185
R7815 gnd.n5645 gnd.n5644 185
R7816 gnd.n5624 gnd.n5623 185
R7817 gnd.n5639 gnd.n5638 185
R7818 gnd.n5637 gnd.n5636 185
R7819 gnd.n5628 gnd.n5627 185
R7820 gnd.n5631 gnd.n5630 185
R7821 gnd.n5615 gnd.n5614 185
R7822 gnd.n5613 gnd.n5612 185
R7823 gnd.n5592 gnd.n5591 185
R7824 gnd.n5607 gnd.n5606 185
R7825 gnd.n5605 gnd.n5604 185
R7826 gnd.n5596 gnd.n5595 185
R7827 gnd.n5599 gnd.n5598 185
R7828 gnd.n5583 gnd.n5582 185
R7829 gnd.n5581 gnd.n5580 185
R7830 gnd.n5560 gnd.n5559 185
R7831 gnd.n5575 gnd.n5574 185
R7832 gnd.n5573 gnd.n5572 185
R7833 gnd.n5564 gnd.n5563 185
R7834 gnd.n5567 gnd.n5566 185
R7835 gnd.n5551 gnd.n5550 185
R7836 gnd.n5549 gnd.n5548 185
R7837 gnd.n5528 gnd.n5527 185
R7838 gnd.n5543 gnd.n5542 185
R7839 gnd.n5541 gnd.n5540 185
R7840 gnd.n5532 gnd.n5531 185
R7841 gnd.n5535 gnd.n5534 185
R7842 gnd.n5520 gnd.n5519 185
R7843 gnd.n5518 gnd.n5517 185
R7844 gnd.n5497 gnd.n5496 185
R7845 gnd.n5512 gnd.n5511 185
R7846 gnd.n5510 gnd.n5509 185
R7847 gnd.n5501 gnd.n5500 185
R7848 gnd.n5504 gnd.n5503 185
R7849 gnd.n6094 gnd.t59 178.987
R7850 gnd.n5475 gnd.t173 178.987
R7851 gnd.n1 gnd.t188 170.774
R7852 gnd.n9 gnd.t400 170.103
R7853 gnd.n8 gnd.t56 170.103
R7854 gnd.n7 gnd.t186 170.103
R7855 gnd.n6 gnd.t184 170.103
R7856 gnd.n5 gnd.t1 170.103
R7857 gnd.n4 gnd.t49 170.103
R7858 gnd.n3 gnd.t15 170.103
R7859 gnd.n2 gnd.t45 170.103
R7860 gnd.n1 gnd.t190 170.103
R7861 gnd.n3733 gnd.n3732 163.367
R7862 gnd.n3737 gnd.n3736 163.367
R7863 gnd.n3741 gnd.n3740 163.367
R7864 gnd.n3745 gnd.n3744 163.367
R7865 gnd.n3749 gnd.n3748 163.367
R7866 gnd.n3753 gnd.n3752 163.367
R7867 gnd.n3757 gnd.n3756 163.367
R7868 gnd.n3761 gnd.n3760 163.367
R7869 gnd.n3765 gnd.n3764 163.367
R7870 gnd.n3769 gnd.n3768 163.367
R7871 gnd.n3773 gnd.n3772 163.367
R7872 gnd.n3777 gnd.n3776 163.367
R7873 gnd.n3781 gnd.n3780 163.367
R7874 gnd.n3785 gnd.n3784 163.367
R7875 gnd.n3790 gnd.n3789 163.367
R7876 gnd.n3794 gnd.n3793 163.367
R7877 gnd.n3875 gnd.n3874 163.367
R7878 gnd.n3871 gnd.n3870 163.367
R7879 gnd.n3866 gnd.n3865 163.367
R7880 gnd.n3862 gnd.n3861 163.367
R7881 gnd.n3858 gnd.n3857 163.367
R7882 gnd.n3854 gnd.n3853 163.367
R7883 gnd.n3850 gnd.n3849 163.367
R7884 gnd.n3846 gnd.n3845 163.367
R7885 gnd.n3842 gnd.n3841 163.367
R7886 gnd.n3838 gnd.n3837 163.367
R7887 gnd.n3834 gnd.n3833 163.367
R7888 gnd.n3830 gnd.n3829 163.367
R7889 gnd.n3826 gnd.n3825 163.367
R7890 gnd.n3822 gnd.n3821 163.367
R7891 gnd.n3818 gnd.n3817 163.367
R7892 gnd.n3814 gnd.n3686 163.367
R7893 gnd.n2474 gnd.n1689 163.367
R7894 gnd.n2406 gnd.n1689 163.367
R7895 gnd.n2482 gnd.n2406 163.367
R7896 gnd.n2482 gnd.n2407 163.367
R7897 gnd.n2478 gnd.n2407 163.367
R7898 gnd.n2478 gnd.n2403 163.367
R7899 gnd.n3466 gnd.n2403 163.367
R7900 gnd.n3466 gnd.n2391 163.367
R7901 gnd.n3470 gnd.n2391 163.367
R7902 gnd.n3471 gnd.n3470 163.367
R7903 gnd.n3471 gnd.n2399 163.367
R7904 gnd.n4076 gnd.n2399 163.367
R7905 gnd.n4076 gnd.n2401 163.367
R7906 gnd.n4072 gnd.n2401 163.367
R7907 gnd.n4072 gnd.n4071 163.367
R7908 gnd.n4071 gnd.n3475 163.367
R7909 gnd.n3490 gnd.n3475 163.367
R7910 gnd.n3490 gnd.n3487 163.367
R7911 gnd.n4061 gnd.n3487 163.367
R7912 gnd.n4061 gnd.n3488 163.367
R7913 gnd.n4057 gnd.n3488 163.367
R7914 gnd.n4057 gnd.n3494 163.367
R7915 gnd.n3502 gnd.n3494 163.367
R7916 gnd.n4047 gnd.n3502 163.367
R7917 gnd.n4047 gnd.n3504 163.367
R7918 gnd.n4043 gnd.n3504 163.367
R7919 gnd.n4043 gnd.n4042 163.367
R7920 gnd.n4042 gnd.n3507 163.367
R7921 gnd.n3521 gnd.n3507 163.367
R7922 gnd.n3521 gnd.n3518 163.367
R7923 gnd.n4032 gnd.n3518 163.367
R7924 gnd.n4032 gnd.n3519 163.367
R7925 gnd.n4028 gnd.n3519 163.367
R7926 gnd.n4028 gnd.n3525 163.367
R7927 gnd.n3540 gnd.n3525 163.367
R7928 gnd.n3540 gnd.n3539 163.367
R7929 gnd.n3544 gnd.n3539 163.367
R7930 gnd.n3547 gnd.n3544 163.367
R7931 gnd.n3548 gnd.n3547 163.367
R7932 gnd.n3548 gnd.n3536 163.367
R7933 gnd.n4010 gnd.n3536 163.367
R7934 gnd.n4010 gnd.n3537 163.367
R7935 gnd.n4006 gnd.n3537 163.367
R7936 gnd.n4006 gnd.n4005 163.367
R7937 gnd.n4005 gnd.n3552 163.367
R7938 gnd.n3560 gnd.n3552 163.367
R7939 gnd.n3994 gnd.n3560 163.367
R7940 gnd.n3994 gnd.n3561 163.367
R7941 gnd.n3990 gnd.n3561 163.367
R7942 gnd.n3990 gnd.n3989 163.367
R7943 gnd.n3989 gnd.n3565 163.367
R7944 gnd.n3574 gnd.n3565 163.367
R7945 gnd.n3978 gnd.n3574 163.367
R7946 gnd.n3978 gnd.n3575 163.367
R7947 gnd.n3974 gnd.n3575 163.367
R7948 gnd.n3974 gnd.n3973 163.367
R7949 gnd.n3973 gnd.n3579 163.367
R7950 gnd.n3587 gnd.n3579 163.367
R7951 gnd.n3962 gnd.n3587 163.367
R7952 gnd.n3962 gnd.n3588 163.367
R7953 gnd.n3958 gnd.n3588 163.367
R7954 gnd.n3958 gnd.n3957 163.367
R7955 gnd.n3957 gnd.n3592 163.367
R7956 gnd.n3602 gnd.n3592 163.367
R7957 gnd.n3948 gnd.n3602 163.367
R7958 gnd.n3948 gnd.n3603 163.367
R7959 gnd.n3944 gnd.n3603 163.367
R7960 gnd.n3944 gnd.n3943 163.367
R7961 gnd.n3943 gnd.n3607 163.367
R7962 gnd.n3615 gnd.n3607 163.367
R7963 gnd.n3933 gnd.n3615 163.367
R7964 gnd.n3933 gnd.n3617 163.367
R7965 gnd.n3929 gnd.n3617 163.367
R7966 gnd.n3929 gnd.n3928 163.367
R7967 gnd.n3928 gnd.n3621 163.367
R7968 gnd.n3632 gnd.n3621 163.367
R7969 gnd.n3919 gnd.n3632 163.367
R7970 gnd.n3919 gnd.n3633 163.367
R7971 gnd.n3915 gnd.n3633 163.367
R7972 gnd.n3915 gnd.n3637 163.367
R7973 gnd.n3649 gnd.n3637 163.367
R7974 gnd.n3649 gnd.n3647 163.367
R7975 gnd.n3905 gnd.n3647 163.367
R7976 gnd.n3905 gnd.n3648 163.367
R7977 gnd.n3901 gnd.n3648 163.367
R7978 gnd.n3901 gnd.n3900 163.367
R7979 gnd.n3900 gnd.n3899 163.367
R7980 gnd.n3899 gnd.n3653 163.367
R7981 gnd.n3895 gnd.n3653 163.367
R7982 gnd.n3895 gnd.n3894 163.367
R7983 gnd.n3894 gnd.n3893 163.367
R7984 gnd.n3893 gnd.n3655 163.367
R7985 gnd.n3682 gnd.n3655 163.367
R7986 gnd.n3682 gnd.n3678 163.367
R7987 gnd.n3882 gnd.n3678 163.367
R7988 gnd.n3882 gnd.n3680 163.367
R7989 gnd.n1664 gnd.n1663 163.367
R7990 gnd.n5038 gnd.n1663 163.367
R7991 gnd.n5036 gnd.n5035 163.367
R7992 gnd.n5032 gnd.n5031 163.367
R7993 gnd.n5028 gnd.n5027 163.367
R7994 gnd.n5024 gnd.n5023 163.367
R7995 gnd.n5020 gnd.n5019 163.367
R7996 gnd.n5016 gnd.n5015 163.367
R7997 gnd.n5012 gnd.n5011 163.367
R7998 gnd.n5008 gnd.n5007 163.367
R7999 gnd.n5004 gnd.n5003 163.367
R8000 gnd.n5000 gnd.n4999 163.367
R8001 gnd.n4996 gnd.n4995 163.367
R8002 gnd.n4992 gnd.n4991 163.367
R8003 gnd.n4988 gnd.n4987 163.367
R8004 gnd.n4984 gnd.n4983 163.367
R8005 gnd.n5047 gnd.n1629 163.367
R8006 gnd.n2412 gnd.n2411 163.367
R8007 gnd.n2417 gnd.n2416 163.367
R8008 gnd.n2421 gnd.n2420 163.367
R8009 gnd.n2425 gnd.n2424 163.367
R8010 gnd.n2429 gnd.n2428 163.367
R8011 gnd.n2433 gnd.n2432 163.367
R8012 gnd.n2437 gnd.n2436 163.367
R8013 gnd.n2441 gnd.n2440 163.367
R8014 gnd.n2445 gnd.n2444 163.367
R8015 gnd.n2449 gnd.n2448 163.367
R8016 gnd.n2453 gnd.n2452 163.367
R8017 gnd.n2457 gnd.n2456 163.367
R8018 gnd.n2461 gnd.n2460 163.367
R8019 gnd.n2465 gnd.n2464 163.367
R8020 gnd.n2469 gnd.n2468 163.367
R8021 gnd.n4976 gnd.n1665 163.367
R8022 gnd.n4976 gnd.n1687 163.367
R8023 gnd.n3457 gnd.n1687 163.367
R8024 gnd.n3458 gnd.n3457 163.367
R8025 gnd.n3458 gnd.n2404 163.367
R8026 gnd.n3462 gnd.n2404 163.367
R8027 gnd.n3462 gnd.n2394 163.367
R8028 gnd.n4085 gnd.n2394 163.367
R8029 gnd.n4085 gnd.n2395 163.367
R8030 gnd.n4081 gnd.n2395 163.367
R8031 gnd.n4081 gnd.n4080 163.367
R8032 gnd.n4080 gnd.n2398 163.367
R8033 gnd.n3480 gnd.n2398 163.367
R8034 gnd.n3480 gnd.n3477 163.367
R8035 gnd.n4069 gnd.n3477 163.367
R8036 gnd.n4069 gnd.n3478 163.367
R8037 gnd.n4065 gnd.n3478 163.367
R8038 gnd.n4065 gnd.n4064 163.367
R8039 gnd.n4064 gnd.n3484 163.367
R8040 gnd.n3496 gnd.n3484 163.367
R8041 gnd.n4055 gnd.n3496 163.367
R8042 gnd.n4055 gnd.n3497 163.367
R8043 gnd.n4051 gnd.n3497 163.367
R8044 gnd.n4051 gnd.n3501 163.367
R8045 gnd.n3511 gnd.n3501 163.367
R8046 gnd.n3511 gnd.n3509 163.367
R8047 gnd.n4040 gnd.n3509 163.367
R8048 gnd.n4040 gnd.n3510 163.367
R8049 gnd.n4036 gnd.n3510 163.367
R8050 gnd.n4036 gnd.n4035 163.367
R8051 gnd.n4035 gnd.n3515 163.367
R8052 gnd.n3527 gnd.n3515 163.367
R8053 gnd.n4026 gnd.n3527 163.367
R8054 gnd.n4026 gnd.n3528 163.367
R8055 gnd.n4022 gnd.n3528 163.367
R8056 gnd.n4022 gnd.n4021 163.367
R8057 gnd.n4021 gnd.n4020 163.367
R8058 gnd.n4020 gnd.n3532 163.367
R8059 gnd.n4016 gnd.n3532 163.367
R8060 gnd.n4016 gnd.n4015 163.367
R8061 gnd.n4015 gnd.n4014 163.367
R8062 gnd.n4014 gnd.n3534 163.367
R8063 gnd.n3554 gnd.n3534 163.367
R8064 gnd.n4003 gnd.n3554 163.367
R8065 gnd.n4003 gnd.n3555 163.367
R8066 gnd.n3999 gnd.n3555 163.367
R8067 gnd.n3999 gnd.n3998 163.367
R8068 gnd.n3998 gnd.n3559 163.367
R8069 gnd.n3567 gnd.n3559 163.367
R8070 gnd.n3987 gnd.n3567 163.367
R8071 gnd.n3987 gnd.n3569 163.367
R8072 gnd.n3983 gnd.n3569 163.367
R8073 gnd.n3983 gnd.n3982 163.367
R8074 gnd.n3982 gnd.n3573 163.367
R8075 gnd.n3581 gnd.n3573 163.367
R8076 gnd.n3971 gnd.n3581 163.367
R8077 gnd.n3971 gnd.n3582 163.367
R8078 gnd.n3967 gnd.n3582 163.367
R8079 gnd.n3967 gnd.n3966 163.367
R8080 gnd.n3966 gnd.n3586 163.367
R8081 gnd.n3594 gnd.n3586 163.367
R8082 gnd.n3955 gnd.n3594 163.367
R8083 gnd.n3955 gnd.n3595 163.367
R8084 gnd.n3951 gnd.n3595 163.367
R8085 gnd.n3951 gnd.n3950 163.367
R8086 gnd.n3950 gnd.n3599 163.367
R8087 gnd.n3609 gnd.n3599 163.367
R8088 gnd.n3941 gnd.n3609 163.367
R8089 gnd.n3941 gnd.n3610 163.367
R8090 gnd.n3937 gnd.n3610 163.367
R8091 gnd.n3937 gnd.n3614 163.367
R8092 gnd.n3625 gnd.n3614 163.367
R8093 gnd.n3625 gnd.n3623 163.367
R8094 gnd.n3926 gnd.n3623 163.367
R8095 gnd.n3926 gnd.n3624 163.367
R8096 gnd.n3922 gnd.n3624 163.367
R8097 gnd.n3922 gnd.n3921 163.367
R8098 gnd.n3921 gnd.n3629 163.367
R8099 gnd.n3913 gnd.n3629 163.367
R8100 gnd.n3913 gnd.n3640 163.367
R8101 gnd.n3909 gnd.n3640 163.367
R8102 gnd.n3909 gnd.n3908 163.367
R8103 gnd.n3908 gnd.n3907 163.367
R8104 gnd.n3907 gnd.n3643 163.367
R8105 gnd.n3664 gnd.n3643 163.367
R8106 gnd.n3664 gnd.n3662 163.367
R8107 gnd.n3668 gnd.n3662 163.367
R8108 gnd.n3672 gnd.n3668 163.367
R8109 gnd.n3673 gnd.n3672 163.367
R8110 gnd.n3673 gnd.n3658 163.367
R8111 gnd.n3891 gnd.n3658 163.367
R8112 gnd.n3891 gnd.n3660 163.367
R8113 gnd.n3887 gnd.n3660 163.367
R8114 gnd.n3887 gnd.n3886 163.367
R8115 gnd.n3886 gnd.n3677 163.367
R8116 gnd.n3728 gnd.n3677 163.367
R8117 gnd.n3724 gnd.n3723 156.462
R8118 gnd.n5682 gnd.n5650 153.042
R8119 gnd.n5746 gnd.n5745 152.079
R8120 gnd.n5714 gnd.n5713 152.079
R8121 gnd.n5682 gnd.n5681 152.079
R8122 gnd.n1678 gnd.n1677 152
R8123 gnd.n1679 gnd.n1668 152
R8124 gnd.n1681 gnd.n1680 152
R8125 gnd.n1683 gnd.n1666 152
R8126 gnd.n1685 gnd.n1684 152
R8127 gnd.n3722 gnd.n3706 152
R8128 gnd.n3714 gnd.n3707 152
R8129 gnd.n3713 gnd.n3712 152
R8130 gnd.n3711 gnd.n3708 152
R8131 gnd.n3709 gnd.t127 150.546
R8132 gnd.t41 gnd.n5724 147.661
R8133 gnd.t404 gnd.n5692 147.661
R8134 gnd.t397 gnd.n5660 147.661
R8135 gnd.t409 gnd.n5629 147.661
R8136 gnd.t17 gnd.n5597 147.661
R8137 gnd.t36 gnd.n5565 147.661
R8138 gnd.t30 gnd.n5533 147.661
R8139 gnd.t11 gnd.n5502 147.661
R8140 gnd.n3811 gnd.n3795 143.351
R8141 gnd.n1645 gnd.n1628 143.351
R8142 gnd.n5046 gnd.n1628 143.351
R8143 gnd.n4783 gnd.n1891 136.385
R8144 gnd.n5049 gnd.n5048 136.385
R8145 gnd.n1675 gnd.t79 130.484
R8146 gnd.n1684 gnd.t76 126.766
R8147 gnd.n1682 gnd.t136 126.766
R8148 gnd.n1668 gnd.t108 126.766
R8149 gnd.n1676 gnd.t164 126.766
R8150 gnd.n3710 gnd.t105 126.766
R8151 gnd.n3712 gnd.t133 126.766
R8152 gnd.n3721 gnd.t73 126.766
R8153 gnd.n3723 gnd.t146 126.766
R8154 gnd.n5741 gnd.n5740 104.615
R8155 gnd.n5740 gnd.n5718 104.615
R8156 gnd.n5733 gnd.n5718 104.615
R8157 gnd.n5733 gnd.n5732 104.615
R8158 gnd.n5732 gnd.n5722 104.615
R8159 gnd.n5725 gnd.n5722 104.615
R8160 gnd.n5709 gnd.n5708 104.615
R8161 gnd.n5708 gnd.n5686 104.615
R8162 gnd.n5701 gnd.n5686 104.615
R8163 gnd.n5701 gnd.n5700 104.615
R8164 gnd.n5700 gnd.n5690 104.615
R8165 gnd.n5693 gnd.n5690 104.615
R8166 gnd.n5677 gnd.n5676 104.615
R8167 gnd.n5676 gnd.n5654 104.615
R8168 gnd.n5669 gnd.n5654 104.615
R8169 gnd.n5669 gnd.n5668 104.615
R8170 gnd.n5668 gnd.n5658 104.615
R8171 gnd.n5661 gnd.n5658 104.615
R8172 gnd.n5646 gnd.n5645 104.615
R8173 gnd.n5645 gnd.n5623 104.615
R8174 gnd.n5638 gnd.n5623 104.615
R8175 gnd.n5638 gnd.n5637 104.615
R8176 gnd.n5637 gnd.n5627 104.615
R8177 gnd.n5630 gnd.n5627 104.615
R8178 gnd.n5614 gnd.n5613 104.615
R8179 gnd.n5613 gnd.n5591 104.615
R8180 gnd.n5606 gnd.n5591 104.615
R8181 gnd.n5606 gnd.n5605 104.615
R8182 gnd.n5605 gnd.n5595 104.615
R8183 gnd.n5598 gnd.n5595 104.615
R8184 gnd.n5582 gnd.n5581 104.615
R8185 gnd.n5581 gnd.n5559 104.615
R8186 gnd.n5574 gnd.n5559 104.615
R8187 gnd.n5574 gnd.n5573 104.615
R8188 gnd.n5573 gnd.n5563 104.615
R8189 gnd.n5566 gnd.n5563 104.615
R8190 gnd.n5550 gnd.n5549 104.615
R8191 gnd.n5549 gnd.n5527 104.615
R8192 gnd.n5542 gnd.n5527 104.615
R8193 gnd.n5542 gnd.n5541 104.615
R8194 gnd.n5541 gnd.n5531 104.615
R8195 gnd.n5534 gnd.n5531 104.615
R8196 gnd.n5519 gnd.n5518 104.615
R8197 gnd.n5518 gnd.n5496 104.615
R8198 gnd.n5511 gnd.n5496 104.615
R8199 gnd.n5511 gnd.n5510 104.615
R8200 gnd.n5510 gnd.n5500 104.615
R8201 gnd.n5503 gnd.n5500 104.615
R8202 gnd.n6388 gnd.t89 100.632
R8203 gnd.n5430 gnd.t141 100.632
R8204 gnd.n8002 gnd.n8001 99.6594
R8205 gnd.n7997 gnd.n294 99.6594
R8206 gnd.n7993 gnd.n293 99.6594
R8207 gnd.n7989 gnd.n292 99.6594
R8208 gnd.n7985 gnd.n291 99.6594
R8209 gnd.n7981 gnd.n290 99.6594
R8210 gnd.n7977 gnd.n289 99.6594
R8211 gnd.n7973 gnd.n288 99.6594
R8212 gnd.n7966 gnd.n287 99.6594
R8213 gnd.n7962 gnd.n286 99.6594
R8214 gnd.n7958 gnd.n285 99.6594
R8215 gnd.n7954 gnd.n284 99.6594
R8216 gnd.n7950 gnd.n283 99.6594
R8217 gnd.n7946 gnd.n282 99.6594
R8218 gnd.n7942 gnd.n281 99.6594
R8219 gnd.n7938 gnd.n280 99.6594
R8220 gnd.n7934 gnd.n279 99.6594
R8221 gnd.n7930 gnd.n278 99.6594
R8222 gnd.n7922 gnd.n277 99.6594
R8223 gnd.n7920 gnd.n276 99.6594
R8224 gnd.n7916 gnd.n275 99.6594
R8225 gnd.n7912 gnd.n274 99.6594
R8226 gnd.n7908 gnd.n273 99.6594
R8227 gnd.n7904 gnd.n272 99.6594
R8228 gnd.n7900 gnd.n271 99.6594
R8229 gnd.n7896 gnd.n270 99.6594
R8230 gnd.n7892 gnd.n269 99.6594
R8231 gnd.n7888 gnd.n268 99.6594
R8232 gnd.n7879 gnd.n267 99.6594
R8233 gnd.n4835 gnd.n4834 99.6594
R8234 gnd.n4829 gnd.n1821 99.6594
R8235 gnd.n4826 gnd.n1822 99.6594
R8236 gnd.n4822 gnd.n1823 99.6594
R8237 gnd.n4818 gnd.n1824 99.6594
R8238 gnd.n4814 gnd.n1825 99.6594
R8239 gnd.n4810 gnd.n1826 99.6594
R8240 gnd.n4806 gnd.n1827 99.6594
R8241 gnd.n4802 gnd.n1828 99.6594
R8242 gnd.n4797 gnd.n1829 99.6594
R8243 gnd.n4793 gnd.n1830 99.6594
R8244 gnd.n4789 gnd.n1831 99.6594
R8245 gnd.n4785 gnd.n1832 99.6594
R8246 gnd.n4780 gnd.n1834 99.6594
R8247 gnd.n4776 gnd.n1835 99.6594
R8248 gnd.n4772 gnd.n1836 99.6594
R8249 gnd.n4768 gnd.n1837 99.6594
R8250 gnd.n4764 gnd.n1838 99.6594
R8251 gnd.n4760 gnd.n1839 99.6594
R8252 gnd.n4756 gnd.n1840 99.6594
R8253 gnd.n4752 gnd.n1841 99.6594
R8254 gnd.n4748 gnd.n1842 99.6594
R8255 gnd.n4744 gnd.n1843 99.6594
R8256 gnd.n4740 gnd.n1844 99.6594
R8257 gnd.n4736 gnd.n1845 99.6594
R8258 gnd.n4732 gnd.n1846 99.6594
R8259 gnd.n4728 gnd.n1847 99.6594
R8260 gnd.n4724 gnd.n1848 99.6594
R8261 gnd.n5098 gnd.n5097 99.6594
R8262 gnd.n5093 gnd.n1595 99.6594
R8263 gnd.n5089 gnd.n1594 99.6594
R8264 gnd.n5085 gnd.n1593 99.6594
R8265 gnd.n5081 gnd.n1592 99.6594
R8266 gnd.n5077 gnd.n1591 99.6594
R8267 gnd.n5073 gnd.n1590 99.6594
R8268 gnd.n5069 gnd.n1589 99.6594
R8269 gnd.n5064 gnd.n1588 99.6594
R8270 gnd.n5060 gnd.n1587 99.6594
R8271 gnd.n5056 gnd.n1586 99.6594
R8272 gnd.n5052 gnd.n1585 99.6594
R8273 gnd.n2662 gnd.n1583 99.6594
R8274 gnd.n2666 gnd.n1582 99.6594
R8275 gnd.n2672 gnd.n1581 99.6594
R8276 gnd.n2676 gnd.n1580 99.6594
R8277 gnd.n2681 gnd.n1579 99.6594
R8278 gnd.n2685 gnd.n1578 99.6594
R8279 gnd.n2691 gnd.n1577 99.6594
R8280 gnd.n2695 gnd.n1576 99.6594
R8281 gnd.n2701 gnd.n1575 99.6594
R8282 gnd.n2705 gnd.n1574 99.6594
R8283 gnd.n2711 gnd.n1573 99.6594
R8284 gnd.n2715 gnd.n1572 99.6594
R8285 gnd.n2721 gnd.n1571 99.6594
R8286 gnd.n2725 gnd.n1570 99.6594
R8287 gnd.n2730 gnd.n1569 99.6594
R8288 gnd.n2733 gnd.n1568 99.6594
R8289 gnd.n5399 gnd.n5398 99.6594
R8290 gnd.n5393 gnd.n1148 99.6594
R8291 gnd.n5390 gnd.n1149 99.6594
R8292 gnd.n5386 gnd.n1150 99.6594
R8293 gnd.n5382 gnd.n1151 99.6594
R8294 gnd.n5378 gnd.n1152 99.6594
R8295 gnd.n5374 gnd.n1153 99.6594
R8296 gnd.n5370 gnd.n1154 99.6594
R8297 gnd.n5366 gnd.n1155 99.6594
R8298 gnd.n5361 gnd.n1156 99.6594
R8299 gnd.n5357 gnd.n1157 99.6594
R8300 gnd.n5353 gnd.n1158 99.6594
R8301 gnd.n5349 gnd.n1159 99.6594
R8302 gnd.n5345 gnd.n1160 99.6594
R8303 gnd.n5341 gnd.n1161 99.6594
R8304 gnd.n5337 gnd.n1162 99.6594
R8305 gnd.n5333 gnd.n1163 99.6594
R8306 gnd.n5329 gnd.n1164 99.6594
R8307 gnd.n5325 gnd.n1165 99.6594
R8308 gnd.n5321 gnd.n1166 99.6594
R8309 gnd.n5317 gnd.n1167 99.6594
R8310 gnd.n5313 gnd.n1168 99.6594
R8311 gnd.n5309 gnd.n1169 99.6594
R8312 gnd.n5305 gnd.n1170 99.6594
R8313 gnd.n5301 gnd.n1171 99.6594
R8314 gnd.n5297 gnd.n1172 99.6594
R8315 gnd.n5293 gnd.n1173 99.6594
R8316 gnd.n5289 gnd.n1174 99.6594
R8317 gnd.n5285 gnd.n1175 99.6594
R8318 gnd.n6867 gnd.n5410 99.6594
R8319 gnd.n6865 gnd.n6864 99.6594
R8320 gnd.n6860 gnd.n5417 99.6594
R8321 gnd.n6858 gnd.n6857 99.6594
R8322 gnd.n6853 gnd.n5424 99.6594
R8323 gnd.n6851 gnd.n6850 99.6594
R8324 gnd.n6846 gnd.n5433 99.6594
R8325 gnd.n6844 gnd.n6843 99.6594
R8326 gnd.n6421 gnd.n6420 99.6594
R8327 gnd.n6415 gnd.n6363 99.6594
R8328 gnd.n6412 gnd.n6364 99.6594
R8329 gnd.n6408 gnd.n6365 99.6594
R8330 gnd.n6404 gnd.n6366 99.6594
R8331 gnd.n6400 gnd.n6367 99.6594
R8332 gnd.n6396 gnd.n6368 99.6594
R8333 gnd.n6392 gnd.n6369 99.6594
R8334 gnd.n481 gnd.n258 99.6594
R8335 gnd.n477 gnd.n259 99.6594
R8336 gnd.n473 gnd.n260 99.6594
R8337 gnd.n469 gnd.n261 99.6594
R8338 gnd.n465 gnd.n262 99.6594
R8339 gnd.n461 gnd.n263 99.6594
R8340 gnd.n457 gnd.n264 99.6594
R8341 gnd.n453 gnd.n265 99.6594
R8342 gnd.n445 gnd.n266 99.6594
R8343 gnd.n1937 gnd.n1849 99.6594
R8344 gnd.n4478 gnd.n1850 99.6594
R8345 gnd.n4495 gnd.n1851 99.6594
R8346 gnd.n4497 gnd.n1852 99.6594
R8347 gnd.n4514 gnd.n1853 99.6594
R8348 gnd.n4516 gnd.n1854 99.6594
R8349 gnd.n4533 gnd.n1855 99.6594
R8350 gnd.n4535 gnd.n1856 99.6594
R8351 gnd.n4551 gnd.n1857 99.6594
R8352 gnd.n6835 gnd.n5440 99.6594
R8353 gnd.n6833 gnd.n6832 99.6594
R8354 gnd.n6828 gnd.n5447 99.6594
R8355 gnd.n6826 gnd.n6825 99.6594
R8356 gnd.n6821 gnd.n5454 99.6594
R8357 gnd.n6819 gnd.n6818 99.6594
R8358 gnd.n6814 gnd.n5461 99.6594
R8359 gnd.n6812 gnd.n6811 99.6594
R8360 gnd.n6807 gnd.n5468 99.6594
R8361 gnd.n6805 gnd.n6804 99.6594
R8362 gnd.n6800 gnd.n5477 99.6594
R8363 gnd.n6798 gnd.n6797 99.6594
R8364 gnd.n6793 gnd.n6792 99.6594
R8365 gnd.n6148 gnd.n6058 99.6594
R8366 gnd.n6146 gnd.n6061 99.6594
R8367 gnd.n6142 gnd.n6141 99.6594
R8368 gnd.n6135 gnd.n6066 99.6594
R8369 gnd.n6134 gnd.n6133 99.6594
R8370 gnd.n6127 gnd.n6072 99.6594
R8371 gnd.n6126 gnd.n6125 99.6594
R8372 gnd.n6119 gnd.n6078 99.6594
R8373 gnd.n6118 gnd.n6117 99.6594
R8374 gnd.n6111 gnd.n6084 99.6594
R8375 gnd.n6110 gnd.n6109 99.6594
R8376 gnd.n6102 gnd.n6090 99.6594
R8377 gnd.n6101 gnd.n6100 99.6594
R8378 gnd.n3235 gnd.n1558 99.6594
R8379 gnd.n3245 gnd.n1559 99.6594
R8380 gnd.n3253 gnd.n1560 99.6594
R8381 gnd.n3255 gnd.n1561 99.6594
R8382 gnd.n3265 gnd.n1562 99.6594
R8383 gnd.n3273 gnd.n1563 99.6594
R8384 gnd.n3275 gnd.n1564 99.6594
R8385 gnd.n3290 gnd.n1565 99.6594
R8386 gnd.n3363 gnd.n1566 99.6594
R8387 gnd.n2914 gnd.n1176 99.6594
R8388 gnd.n2918 gnd.n1177 99.6594
R8389 gnd.n2924 gnd.n1178 99.6594
R8390 gnd.n2928 gnd.n1179 99.6594
R8391 gnd.n2934 gnd.n1180 99.6594
R8392 gnd.n2938 gnd.n1181 99.6594
R8393 gnd.n2944 gnd.n1182 99.6594
R8394 gnd.n2948 gnd.n1183 99.6594
R8395 gnd.n2905 gnd.n1184 99.6594
R8396 gnd.n2917 gnd.n1176 99.6594
R8397 gnd.n2923 gnd.n1177 99.6594
R8398 gnd.n2927 gnd.n1178 99.6594
R8399 gnd.n2933 gnd.n1179 99.6594
R8400 gnd.n2937 gnd.n1180 99.6594
R8401 gnd.n2943 gnd.n1181 99.6594
R8402 gnd.n2947 gnd.n1182 99.6594
R8403 gnd.n2904 gnd.n1183 99.6594
R8404 gnd.n2900 gnd.n1184 99.6594
R8405 gnd.n3289 gnd.n1566 99.6594
R8406 gnd.n3276 gnd.n1565 99.6594
R8407 gnd.n3274 gnd.n1564 99.6594
R8408 gnd.n3266 gnd.n1563 99.6594
R8409 gnd.n3256 gnd.n1562 99.6594
R8410 gnd.n3254 gnd.n1561 99.6594
R8411 gnd.n3246 gnd.n1560 99.6594
R8412 gnd.n3236 gnd.n1559 99.6594
R8413 gnd.n3234 gnd.n1558 99.6594
R8414 gnd.n6149 gnd.n6148 99.6594
R8415 gnd.n6143 gnd.n6061 99.6594
R8416 gnd.n6141 gnd.n6140 99.6594
R8417 gnd.n6136 gnd.n6135 99.6594
R8418 gnd.n6133 gnd.n6132 99.6594
R8419 gnd.n6128 gnd.n6127 99.6594
R8420 gnd.n6125 gnd.n6124 99.6594
R8421 gnd.n6120 gnd.n6119 99.6594
R8422 gnd.n6117 gnd.n6116 99.6594
R8423 gnd.n6112 gnd.n6111 99.6594
R8424 gnd.n6109 gnd.n6108 99.6594
R8425 gnd.n6103 gnd.n6102 99.6594
R8426 gnd.n6100 gnd.n6056 99.6594
R8427 gnd.n6792 gnd.n5479 99.6594
R8428 gnd.n6799 gnd.n6798 99.6594
R8429 gnd.n5477 gnd.n5469 99.6594
R8430 gnd.n6806 gnd.n6805 99.6594
R8431 gnd.n5468 gnd.n5462 99.6594
R8432 gnd.n6813 gnd.n6812 99.6594
R8433 gnd.n5461 gnd.n5455 99.6594
R8434 gnd.n6820 gnd.n6819 99.6594
R8435 gnd.n5454 gnd.n5448 99.6594
R8436 gnd.n6827 gnd.n6826 99.6594
R8437 gnd.n5447 gnd.n5441 99.6594
R8438 gnd.n6834 gnd.n6833 99.6594
R8439 gnd.n5440 gnd.n5437 99.6594
R8440 gnd.n4479 gnd.n1849 99.6594
R8441 gnd.n4494 gnd.n1850 99.6594
R8442 gnd.n4498 gnd.n1851 99.6594
R8443 gnd.n4513 gnd.n1852 99.6594
R8444 gnd.n4517 gnd.n1853 99.6594
R8445 gnd.n4532 gnd.n1854 99.6594
R8446 gnd.n4536 gnd.n1855 99.6594
R8447 gnd.n4550 gnd.n1856 99.6594
R8448 gnd.n4416 gnd.n1857 99.6594
R8449 gnd.n452 gnd.n266 99.6594
R8450 gnd.n456 gnd.n265 99.6594
R8451 gnd.n460 gnd.n264 99.6594
R8452 gnd.n464 gnd.n263 99.6594
R8453 gnd.n468 gnd.n262 99.6594
R8454 gnd.n472 gnd.n261 99.6594
R8455 gnd.n476 gnd.n260 99.6594
R8456 gnd.n480 gnd.n259 99.6594
R8457 gnd.n355 gnd.n258 99.6594
R8458 gnd.n6421 gnd.n6371 99.6594
R8459 gnd.n6413 gnd.n6363 99.6594
R8460 gnd.n6409 gnd.n6364 99.6594
R8461 gnd.n6405 gnd.n6365 99.6594
R8462 gnd.n6401 gnd.n6366 99.6594
R8463 gnd.n6397 gnd.n6367 99.6594
R8464 gnd.n6393 gnd.n6368 99.6594
R8465 gnd.n6369 gnd.n6018 99.6594
R8466 gnd.n6845 gnd.n6844 99.6594
R8467 gnd.n5433 gnd.n5425 99.6594
R8468 gnd.n6852 gnd.n6851 99.6594
R8469 gnd.n5424 gnd.n5418 99.6594
R8470 gnd.n6859 gnd.n6858 99.6594
R8471 gnd.n5417 gnd.n5411 99.6594
R8472 gnd.n6866 gnd.n6865 99.6594
R8473 gnd.n5410 gnd.n5407 99.6594
R8474 gnd.n5399 gnd.n1188 99.6594
R8475 gnd.n5391 gnd.n1148 99.6594
R8476 gnd.n5387 gnd.n1149 99.6594
R8477 gnd.n5383 gnd.n1150 99.6594
R8478 gnd.n5379 gnd.n1151 99.6594
R8479 gnd.n5375 gnd.n1152 99.6594
R8480 gnd.n5371 gnd.n1153 99.6594
R8481 gnd.n5367 gnd.n1154 99.6594
R8482 gnd.n5362 gnd.n1155 99.6594
R8483 gnd.n5358 gnd.n1156 99.6594
R8484 gnd.n5354 gnd.n1157 99.6594
R8485 gnd.n5350 gnd.n1158 99.6594
R8486 gnd.n5346 gnd.n1159 99.6594
R8487 gnd.n5342 gnd.n1160 99.6594
R8488 gnd.n5338 gnd.n1161 99.6594
R8489 gnd.n5334 gnd.n1162 99.6594
R8490 gnd.n5330 gnd.n1163 99.6594
R8491 gnd.n5326 gnd.n1164 99.6594
R8492 gnd.n5322 gnd.n1165 99.6594
R8493 gnd.n5318 gnd.n1166 99.6594
R8494 gnd.n5314 gnd.n1167 99.6594
R8495 gnd.n5310 gnd.n1168 99.6594
R8496 gnd.n5306 gnd.n1169 99.6594
R8497 gnd.n5302 gnd.n1170 99.6594
R8498 gnd.n5298 gnd.n1171 99.6594
R8499 gnd.n5294 gnd.n1172 99.6594
R8500 gnd.n5290 gnd.n1173 99.6594
R8501 gnd.n5286 gnd.n1174 99.6594
R8502 gnd.n1258 gnd.n1175 99.6594
R8503 gnd.n2643 gnd.n1568 99.6594
R8504 gnd.n2724 gnd.n1569 99.6594
R8505 gnd.n2722 gnd.n1570 99.6594
R8506 gnd.n2714 gnd.n1571 99.6594
R8507 gnd.n2712 gnd.n1572 99.6594
R8508 gnd.n2704 gnd.n1573 99.6594
R8509 gnd.n2702 gnd.n1574 99.6594
R8510 gnd.n2694 gnd.n1575 99.6594
R8511 gnd.n2692 gnd.n1576 99.6594
R8512 gnd.n2684 gnd.n1577 99.6594
R8513 gnd.n2656 gnd.n1578 99.6594
R8514 gnd.n2675 gnd.n1579 99.6594
R8515 gnd.n2673 gnd.n1580 99.6594
R8516 gnd.n2665 gnd.n1581 99.6594
R8517 gnd.n2663 gnd.n1582 99.6594
R8518 gnd.n5051 gnd.n1584 99.6594
R8519 gnd.n5055 gnd.n1585 99.6594
R8520 gnd.n5059 gnd.n1586 99.6594
R8521 gnd.n5063 gnd.n1587 99.6594
R8522 gnd.n5068 gnd.n1588 99.6594
R8523 gnd.n5072 gnd.n1589 99.6594
R8524 gnd.n5076 gnd.n1590 99.6594
R8525 gnd.n5080 gnd.n1591 99.6594
R8526 gnd.n5084 gnd.n1592 99.6594
R8527 gnd.n5088 gnd.n1593 99.6594
R8528 gnd.n5092 gnd.n1594 99.6594
R8529 gnd.n1596 gnd.n1595 99.6594
R8530 gnd.n5098 gnd.n1555 99.6594
R8531 gnd.n4835 gnd.n1861 99.6594
R8532 gnd.n4827 gnd.n1821 99.6594
R8533 gnd.n4823 gnd.n1822 99.6594
R8534 gnd.n4819 gnd.n1823 99.6594
R8535 gnd.n4815 gnd.n1824 99.6594
R8536 gnd.n4811 gnd.n1825 99.6594
R8537 gnd.n4807 gnd.n1826 99.6594
R8538 gnd.n4803 gnd.n1827 99.6594
R8539 gnd.n4798 gnd.n1828 99.6594
R8540 gnd.n4794 gnd.n1829 99.6594
R8541 gnd.n4790 gnd.n1830 99.6594
R8542 gnd.n4786 gnd.n1831 99.6594
R8543 gnd.n4781 gnd.n1833 99.6594
R8544 gnd.n4777 gnd.n1834 99.6594
R8545 gnd.n4773 gnd.n1835 99.6594
R8546 gnd.n4769 gnd.n1836 99.6594
R8547 gnd.n4765 gnd.n1837 99.6594
R8548 gnd.n4761 gnd.n1838 99.6594
R8549 gnd.n4757 gnd.n1839 99.6594
R8550 gnd.n4753 gnd.n1840 99.6594
R8551 gnd.n4749 gnd.n1841 99.6594
R8552 gnd.n4745 gnd.n1842 99.6594
R8553 gnd.n4741 gnd.n1843 99.6594
R8554 gnd.n4737 gnd.n1844 99.6594
R8555 gnd.n4733 gnd.n1845 99.6594
R8556 gnd.n4729 gnd.n1846 99.6594
R8557 gnd.n4725 gnd.n1847 99.6594
R8558 gnd.n1932 gnd.n1848 99.6594
R8559 gnd.n7887 gnd.n267 99.6594
R8560 gnd.n7891 gnd.n268 99.6594
R8561 gnd.n7895 gnd.n269 99.6594
R8562 gnd.n7899 gnd.n270 99.6594
R8563 gnd.n7903 gnd.n271 99.6594
R8564 gnd.n7907 gnd.n272 99.6594
R8565 gnd.n7911 gnd.n273 99.6594
R8566 gnd.n7915 gnd.n274 99.6594
R8567 gnd.n7919 gnd.n275 99.6594
R8568 gnd.n7923 gnd.n276 99.6594
R8569 gnd.n7929 gnd.n277 99.6594
R8570 gnd.n7933 gnd.n278 99.6594
R8571 gnd.n7937 gnd.n279 99.6594
R8572 gnd.n7941 gnd.n280 99.6594
R8573 gnd.n7945 gnd.n281 99.6594
R8574 gnd.n7949 gnd.n282 99.6594
R8575 gnd.n7953 gnd.n283 99.6594
R8576 gnd.n7957 gnd.n284 99.6594
R8577 gnd.n7961 gnd.n285 99.6594
R8578 gnd.n7965 gnd.n286 99.6594
R8579 gnd.n7972 gnd.n287 99.6594
R8580 gnd.n7976 gnd.n288 99.6594
R8581 gnd.n7980 gnd.n289 99.6594
R8582 gnd.n7984 gnd.n290 99.6594
R8583 gnd.n7988 gnd.n291 99.6594
R8584 gnd.n7992 gnd.n292 99.6594
R8585 gnd.n7996 gnd.n293 99.6594
R8586 gnd.n295 gnd.n294 99.6594
R8587 gnd.n8002 gnd.n256 99.6594
R8588 gnd.n3350 gnd.n3349 99.6594
R8589 gnd.n2636 gnd.n2566 99.6594
R8590 gnd.n2638 gnd.n2567 99.6594
R8591 gnd.n3227 gnd.n2568 99.6594
R8592 gnd.n3229 gnd.n2569 99.6594
R8593 gnd.n3240 gnd.n2570 99.6594
R8594 gnd.n3242 gnd.n2571 99.6594
R8595 gnd.n3250 gnd.n2572 99.6594
R8596 gnd.n3260 gnd.n2573 99.6594
R8597 gnd.n3262 gnd.n2574 99.6594
R8598 gnd.n3270 gnd.n2575 99.6594
R8599 gnd.n3280 gnd.n2576 99.6594
R8600 gnd.n3286 gnd.n2578 99.6594
R8601 gnd.n2579 gnd.n2548 99.6594
R8602 gnd.n3350 gnd.n2581 99.6594
R8603 gnd.n2637 gnd.n2566 99.6594
R8604 gnd.n3226 gnd.n2567 99.6594
R8605 gnd.n3228 gnd.n2568 99.6594
R8606 gnd.n3239 gnd.n2569 99.6594
R8607 gnd.n3241 gnd.n2570 99.6594
R8608 gnd.n3249 gnd.n2571 99.6594
R8609 gnd.n3259 gnd.n2572 99.6594
R8610 gnd.n3261 gnd.n2573 99.6594
R8611 gnd.n3269 gnd.n2574 99.6594
R8612 gnd.n3279 gnd.n2575 99.6594
R8613 gnd.n3281 gnd.n2576 99.6594
R8614 gnd.n2578 gnd.n2577 99.6594
R8615 gnd.n2579 gnd.n2545 99.6594
R8616 gnd.n4456 gnd.n4451 99.6594
R8617 gnd.n4460 gnd.n4458 99.6594
R8618 gnd.n4467 gnd.n4447 99.6594
R8619 gnd.n4471 gnd.n4469 99.6594
R8620 gnd.n4484 gnd.n4444 99.6594
R8621 gnd.n4488 gnd.n4486 99.6594
R8622 gnd.n4503 gnd.n4437 99.6594
R8623 gnd.n4507 gnd.n4505 99.6594
R8624 gnd.n4522 gnd.n4430 99.6594
R8625 gnd.n4526 gnd.n4524 99.6594
R8626 gnd.n4541 gnd.n4422 99.6594
R8627 gnd.n4544 gnd.n4543 99.6594
R8628 gnd.n4558 gnd.n4557 99.6594
R8629 gnd.n4561 gnd.n4560 99.6594
R8630 gnd.n4543 gnd.n4542 99.6594
R8631 gnd.n4525 gnd.n4422 99.6594
R8632 gnd.n4524 gnd.n4523 99.6594
R8633 gnd.n4506 gnd.n4430 99.6594
R8634 gnd.n4505 gnd.n4504 99.6594
R8635 gnd.n4487 gnd.n4437 99.6594
R8636 gnd.n4486 gnd.n4485 99.6594
R8637 gnd.n4470 gnd.n4444 99.6594
R8638 gnd.n4469 gnd.n4468 99.6594
R8639 gnd.n4459 gnd.n4447 99.6594
R8640 gnd.n4458 gnd.n4457 99.6594
R8641 gnd.n4451 gnd.n1808 99.6594
R8642 gnd.n4562 gnd.n4561 99.6594
R8643 gnd.n4559 gnd.n4558 99.6594
R8644 gnd.n3282 gnd.t104 98.63
R8645 gnd.n4417 gnd.t64 98.63
R8646 gnd.n2550 gnd.t95 98.63
R8647 gnd.n1881 gnd.t157 98.63
R8648 gnd.n1904 gnd.t160 98.63
R8649 gnd.n1926 gnd.t123 98.63
R8650 gnd.n352 gnd.t84 98.63
R8651 gnd.n332 gnd.t91 98.63
R8652 gnd.n7968 gnd.t119 98.63
R8653 gnd.n372 gnd.t168 98.63
R8654 gnd.n1208 gnd.t113 98.63
R8655 gnd.n1230 gnd.t132 98.63
R8656 gnd.n1252 gnd.t154 98.63
R8657 gnd.n2901 gnd.t100 98.63
R8658 gnd.n1613 gnd.t125 98.63
R8659 gnd.n2641 gnd.t144 98.63
R8660 gnd.n2654 gnd.t175 98.63
R8661 gnd.n4410 gnd.t67 98.63
R8662 gnd.n7512 gnd.n7511 97.3241
R8663 gnd.n7513 gnd.n7512 97.3241
R8664 gnd.n7513 gnd.n688 97.3241
R8665 gnd.n7521 gnd.n688 97.3241
R8666 gnd.n7522 gnd.n7521 97.3241
R8667 gnd.n7523 gnd.n7522 97.3241
R8668 gnd.n7523 gnd.n682 97.3241
R8669 gnd.n7531 gnd.n682 97.3241
R8670 gnd.n7532 gnd.n7531 97.3241
R8671 gnd.n7533 gnd.n7532 97.3241
R8672 gnd.n7533 gnd.n676 97.3241
R8673 gnd.n7541 gnd.n676 97.3241
R8674 gnd.n7542 gnd.n7541 97.3241
R8675 gnd.n7543 gnd.n7542 97.3241
R8676 gnd.n7543 gnd.n670 97.3241
R8677 gnd.n7551 gnd.n670 97.3241
R8678 gnd.n7552 gnd.n7551 97.3241
R8679 gnd.n7553 gnd.n7552 97.3241
R8680 gnd.n7553 gnd.n664 97.3241
R8681 gnd.n7561 gnd.n664 97.3241
R8682 gnd.n7562 gnd.n7561 97.3241
R8683 gnd.n7563 gnd.n7562 97.3241
R8684 gnd.n7563 gnd.n658 97.3241
R8685 gnd.n7571 gnd.n658 97.3241
R8686 gnd.n7572 gnd.n7571 97.3241
R8687 gnd.n7573 gnd.n7572 97.3241
R8688 gnd.n7573 gnd.n652 97.3241
R8689 gnd.n7581 gnd.n652 97.3241
R8690 gnd.n7582 gnd.n7581 97.3241
R8691 gnd.n7583 gnd.n7582 97.3241
R8692 gnd.n7583 gnd.n646 97.3241
R8693 gnd.n7591 gnd.n646 97.3241
R8694 gnd.n7592 gnd.n7591 97.3241
R8695 gnd.n7593 gnd.n7592 97.3241
R8696 gnd.n7593 gnd.n640 97.3241
R8697 gnd.n7601 gnd.n640 97.3241
R8698 gnd.n7602 gnd.n7601 97.3241
R8699 gnd.n7603 gnd.n7602 97.3241
R8700 gnd.n7603 gnd.n634 97.3241
R8701 gnd.n7611 gnd.n634 97.3241
R8702 gnd.n7612 gnd.n7611 97.3241
R8703 gnd.n7613 gnd.n7612 97.3241
R8704 gnd.n7613 gnd.n628 97.3241
R8705 gnd.n7621 gnd.n628 97.3241
R8706 gnd.n7622 gnd.n7621 97.3241
R8707 gnd.n7623 gnd.n7622 97.3241
R8708 gnd.n7623 gnd.n622 97.3241
R8709 gnd.n7631 gnd.n622 97.3241
R8710 gnd.n7632 gnd.n7631 97.3241
R8711 gnd.n7633 gnd.n7632 97.3241
R8712 gnd.n7633 gnd.n616 97.3241
R8713 gnd.n7641 gnd.n616 97.3241
R8714 gnd.n7642 gnd.n7641 97.3241
R8715 gnd.n7643 gnd.n7642 97.3241
R8716 gnd.n7643 gnd.n610 97.3241
R8717 gnd.n7651 gnd.n610 97.3241
R8718 gnd.n7652 gnd.n7651 97.3241
R8719 gnd.n7653 gnd.n7652 97.3241
R8720 gnd.n7653 gnd.n604 97.3241
R8721 gnd.n7661 gnd.n604 97.3241
R8722 gnd.n7662 gnd.n7661 97.3241
R8723 gnd.n7663 gnd.n7662 97.3241
R8724 gnd.n7663 gnd.n598 97.3241
R8725 gnd.n7671 gnd.n598 97.3241
R8726 gnd.n7672 gnd.n7671 97.3241
R8727 gnd.n7673 gnd.n7672 97.3241
R8728 gnd.n7673 gnd.n592 97.3241
R8729 gnd.n7681 gnd.n592 97.3241
R8730 gnd.n7682 gnd.n7681 97.3241
R8731 gnd.n7683 gnd.n7682 97.3241
R8732 gnd.n7683 gnd.n586 97.3241
R8733 gnd.n7691 gnd.n586 97.3241
R8734 gnd.n7692 gnd.n7691 97.3241
R8735 gnd.n7693 gnd.n7692 97.3241
R8736 gnd.n7693 gnd.n580 97.3241
R8737 gnd.n7701 gnd.n580 97.3241
R8738 gnd.n7702 gnd.n7701 97.3241
R8739 gnd.n7703 gnd.n7702 97.3241
R8740 gnd.n7703 gnd.n574 97.3241
R8741 gnd.n7711 gnd.n574 97.3241
R8742 gnd.n7712 gnd.n7711 97.3241
R8743 gnd.n7714 gnd.n7712 97.3241
R8744 gnd.n7714 gnd.n7713 97.3241
R8745 gnd.n2408 gnd.t151 96.6984
R8746 gnd.n3812 gnd.t116 96.6984
R8747 gnd.n4980 gnd.t72 96.6906
R8748 gnd.n3704 gnd.t162 96.6906
R8749 gnd.n1675 gnd.n1674 81.8399
R8750 gnd.n6389 gnd.t88 74.8376
R8751 gnd.n5431 gnd.t142 74.8376
R8752 gnd.n2409 gnd.t150 72.8438
R8753 gnd.n3813 gnd.t117 72.8438
R8754 gnd.n1676 gnd.n1669 72.8411
R8755 gnd.n1682 gnd.n1667 72.8411
R8756 gnd.n3721 gnd.n3720 72.8411
R8757 gnd.n3283 gnd.t103 72.836
R8758 gnd.n4981 gnd.t71 72.836
R8759 gnd.n3705 gnd.t163 72.836
R8760 gnd.n4418 gnd.t63 72.836
R8761 gnd.n2551 gnd.t96 72.836
R8762 gnd.n1882 gnd.t156 72.836
R8763 gnd.n1905 gnd.t159 72.836
R8764 gnd.n1927 gnd.t122 72.836
R8765 gnd.n353 gnd.t85 72.836
R8766 gnd.n333 gnd.t92 72.836
R8767 gnd.n7969 gnd.t120 72.836
R8768 gnd.n373 gnd.t169 72.836
R8769 gnd.n1209 gnd.t112 72.836
R8770 gnd.n1231 gnd.t131 72.836
R8771 gnd.n1253 gnd.t153 72.836
R8772 gnd.n2902 gnd.t99 72.836
R8773 gnd.n1614 gnd.t126 72.836
R8774 gnd.n2642 gnd.t145 72.836
R8775 gnd.n2655 gnd.t176 72.836
R8776 gnd.n4411 gnd.t68 72.836
R8777 gnd.n3732 gnd.n3688 71.676
R8778 gnd.n3736 gnd.n3689 71.676
R8779 gnd.n3740 gnd.n3690 71.676
R8780 gnd.n3744 gnd.n3691 71.676
R8781 gnd.n3748 gnd.n3692 71.676
R8782 gnd.n3752 gnd.n3693 71.676
R8783 gnd.n3756 gnd.n3694 71.676
R8784 gnd.n3760 gnd.n3695 71.676
R8785 gnd.n3764 gnd.n3696 71.676
R8786 gnd.n3768 gnd.n3697 71.676
R8787 gnd.n3772 gnd.n3698 71.676
R8788 gnd.n3776 gnd.n3699 71.676
R8789 gnd.n3780 gnd.n3700 71.676
R8790 gnd.n3784 gnd.n3701 71.676
R8791 gnd.n3789 gnd.n3702 71.676
R8792 gnd.n3793 gnd.n3703 71.676
R8793 gnd.n3875 gnd.n3811 71.676
R8794 gnd.n3871 gnd.n3810 71.676
R8795 gnd.n3866 gnd.n3809 71.676
R8796 gnd.n3862 gnd.n3808 71.676
R8797 gnd.n3858 gnd.n3807 71.676
R8798 gnd.n3854 gnd.n3806 71.676
R8799 gnd.n3850 gnd.n3805 71.676
R8800 gnd.n3846 gnd.n3804 71.676
R8801 gnd.n3842 gnd.n3803 71.676
R8802 gnd.n3838 gnd.n3802 71.676
R8803 gnd.n3834 gnd.n3801 71.676
R8804 gnd.n3830 gnd.n3800 71.676
R8805 gnd.n3826 gnd.n3799 71.676
R8806 gnd.n3822 gnd.n3798 71.676
R8807 gnd.n3818 gnd.n3797 71.676
R8808 gnd.n3814 gnd.n3796 71.676
R8809 gnd.n3878 gnd.n3877 71.676
R8810 gnd.n5044 gnd.n5043 71.676
R8811 gnd.n5038 gnd.n1631 71.676
R8812 gnd.n5035 gnd.n1632 71.676
R8813 gnd.n5031 gnd.n1633 71.676
R8814 gnd.n5027 gnd.n1634 71.676
R8815 gnd.n5023 gnd.n1635 71.676
R8816 gnd.n5019 gnd.n1636 71.676
R8817 gnd.n5015 gnd.n1637 71.676
R8818 gnd.n5011 gnd.n1638 71.676
R8819 gnd.n5007 gnd.n1639 71.676
R8820 gnd.n5003 gnd.n1640 71.676
R8821 gnd.n4999 gnd.n1641 71.676
R8822 gnd.n4995 gnd.n1642 71.676
R8823 gnd.n4991 gnd.n1643 71.676
R8824 gnd.n4987 gnd.n1644 71.676
R8825 gnd.n4983 gnd.n1645 71.676
R8826 gnd.n1646 gnd.n1629 71.676
R8827 gnd.n2412 gnd.n1647 71.676
R8828 gnd.n2417 gnd.n1648 71.676
R8829 gnd.n2421 gnd.n1649 71.676
R8830 gnd.n2425 gnd.n1650 71.676
R8831 gnd.n2429 gnd.n1651 71.676
R8832 gnd.n2433 gnd.n1652 71.676
R8833 gnd.n2437 gnd.n1653 71.676
R8834 gnd.n2441 gnd.n1654 71.676
R8835 gnd.n2445 gnd.n1655 71.676
R8836 gnd.n2449 gnd.n1656 71.676
R8837 gnd.n2453 gnd.n1657 71.676
R8838 gnd.n2457 gnd.n1658 71.676
R8839 gnd.n2461 gnd.n1659 71.676
R8840 gnd.n2465 gnd.n1660 71.676
R8841 gnd.n2469 gnd.n1661 71.676
R8842 gnd.n5044 gnd.n1664 71.676
R8843 gnd.n5036 gnd.n1631 71.676
R8844 gnd.n5032 gnd.n1632 71.676
R8845 gnd.n5028 gnd.n1633 71.676
R8846 gnd.n5024 gnd.n1634 71.676
R8847 gnd.n5020 gnd.n1635 71.676
R8848 gnd.n5016 gnd.n1636 71.676
R8849 gnd.n5012 gnd.n1637 71.676
R8850 gnd.n5008 gnd.n1638 71.676
R8851 gnd.n5004 gnd.n1639 71.676
R8852 gnd.n5000 gnd.n1640 71.676
R8853 gnd.n4996 gnd.n1641 71.676
R8854 gnd.n4992 gnd.n1642 71.676
R8855 gnd.n4988 gnd.n1643 71.676
R8856 gnd.n4984 gnd.n1644 71.676
R8857 gnd.n5047 gnd.n5046 71.676
R8858 gnd.n2411 gnd.n1646 71.676
R8859 gnd.n2416 gnd.n1647 71.676
R8860 gnd.n2420 gnd.n1648 71.676
R8861 gnd.n2424 gnd.n1649 71.676
R8862 gnd.n2428 gnd.n1650 71.676
R8863 gnd.n2432 gnd.n1651 71.676
R8864 gnd.n2436 gnd.n1652 71.676
R8865 gnd.n2440 gnd.n1653 71.676
R8866 gnd.n2444 gnd.n1654 71.676
R8867 gnd.n2448 gnd.n1655 71.676
R8868 gnd.n2452 gnd.n1656 71.676
R8869 gnd.n2456 gnd.n1657 71.676
R8870 gnd.n2460 gnd.n1658 71.676
R8871 gnd.n2464 gnd.n1659 71.676
R8872 gnd.n2468 gnd.n1660 71.676
R8873 gnd.n2472 gnd.n1661 71.676
R8874 gnd.n3877 gnd.n3686 71.676
R8875 gnd.n3817 gnd.n3796 71.676
R8876 gnd.n3821 gnd.n3797 71.676
R8877 gnd.n3825 gnd.n3798 71.676
R8878 gnd.n3829 gnd.n3799 71.676
R8879 gnd.n3833 gnd.n3800 71.676
R8880 gnd.n3837 gnd.n3801 71.676
R8881 gnd.n3841 gnd.n3802 71.676
R8882 gnd.n3845 gnd.n3803 71.676
R8883 gnd.n3849 gnd.n3804 71.676
R8884 gnd.n3853 gnd.n3805 71.676
R8885 gnd.n3857 gnd.n3806 71.676
R8886 gnd.n3861 gnd.n3807 71.676
R8887 gnd.n3865 gnd.n3808 71.676
R8888 gnd.n3870 gnd.n3809 71.676
R8889 gnd.n3874 gnd.n3810 71.676
R8890 gnd.n3795 gnd.n3794 71.676
R8891 gnd.n3790 gnd.n3703 71.676
R8892 gnd.n3785 gnd.n3702 71.676
R8893 gnd.n3781 gnd.n3701 71.676
R8894 gnd.n3777 gnd.n3700 71.676
R8895 gnd.n3773 gnd.n3699 71.676
R8896 gnd.n3769 gnd.n3698 71.676
R8897 gnd.n3765 gnd.n3697 71.676
R8898 gnd.n3761 gnd.n3696 71.676
R8899 gnd.n3757 gnd.n3695 71.676
R8900 gnd.n3753 gnd.n3694 71.676
R8901 gnd.n3749 gnd.n3693 71.676
R8902 gnd.n3745 gnd.n3692 71.676
R8903 gnd.n3741 gnd.n3691 71.676
R8904 gnd.n3737 gnd.n3690 71.676
R8905 gnd.n3733 gnd.n3689 71.676
R8906 gnd.n3729 gnd.n3688 71.676
R8907 gnd.n10 gnd.t19 69.1507
R8908 gnd.n18 gnd.t411 68.4792
R8909 gnd.n17 gnd.t25 68.4792
R8910 gnd.n16 gnd.t393 68.4792
R8911 gnd.n15 gnd.t39 68.4792
R8912 gnd.n14 gnd.t395 68.4792
R8913 gnd.n13 gnd.t182 68.4792
R8914 gnd.n12 gnd.t51 68.4792
R8915 gnd.n11 gnd.t8 68.4792
R8916 gnd.n10 gnd.t47 68.4792
R8917 gnd.n6156 gnd.n6057 64.369
R8918 gnd.n2414 gnd.n2409 59.5399
R8919 gnd.n3868 gnd.n3813 59.5399
R8920 gnd.n4982 gnd.n4981 59.5399
R8921 gnd.n3787 gnd.n3705 59.5399
R8922 gnd.n4979 gnd.n1685 59.1804
R8923 gnd.n7713 gnd.n219 58.3947
R8924 gnd.n6875 gnd.n5401 57.3586
R8925 gnd.n6309 gnd.t344 56.407
R8926 gnd.n6250 gnd.t367 56.407
R8927 gnd.n6269 gnd.t323 56.407
R8928 gnd.n6289 gnd.t210 56.407
R8929 gnd.n80 gnd.t310 56.407
R8930 gnd.n21 gnd.t229 56.407
R8931 gnd.n40 gnd.t298 56.407
R8932 gnd.n60 gnd.t355 56.407
R8933 gnd.n6326 gnd.t374 55.8337
R8934 gnd.n6267 gnd.t202 55.8337
R8935 gnd.n6286 gnd.t216 55.8337
R8936 gnd.n6306 gnd.t284 55.8337
R8937 gnd.n97 gnd.t314 55.8337
R8938 gnd.n38 gnd.t227 55.8337
R8939 gnd.n57 gnd.t366 55.8337
R8940 gnd.n77 gnd.t359 55.8337
R8941 gnd.n1673 gnd.n1672 54.358
R8942 gnd.n3718 gnd.n3717 54.358
R8943 gnd.n6309 gnd.n6308 53.0052
R8944 gnd.n6311 gnd.n6310 53.0052
R8945 gnd.n6313 gnd.n6312 53.0052
R8946 gnd.n6315 gnd.n6314 53.0052
R8947 gnd.n6317 gnd.n6316 53.0052
R8948 gnd.n6319 gnd.n6318 53.0052
R8949 gnd.n6321 gnd.n6320 53.0052
R8950 gnd.n6323 gnd.n6322 53.0052
R8951 gnd.n6325 gnd.n6324 53.0052
R8952 gnd.n6250 gnd.n6249 53.0052
R8953 gnd.n6252 gnd.n6251 53.0052
R8954 gnd.n6254 gnd.n6253 53.0052
R8955 gnd.n6256 gnd.n6255 53.0052
R8956 gnd.n6258 gnd.n6257 53.0052
R8957 gnd.n6260 gnd.n6259 53.0052
R8958 gnd.n6262 gnd.n6261 53.0052
R8959 gnd.n6264 gnd.n6263 53.0052
R8960 gnd.n6266 gnd.n6265 53.0052
R8961 gnd.n6269 gnd.n6268 53.0052
R8962 gnd.n6271 gnd.n6270 53.0052
R8963 gnd.n6273 gnd.n6272 53.0052
R8964 gnd.n6275 gnd.n6274 53.0052
R8965 gnd.n6277 gnd.n6276 53.0052
R8966 gnd.n6279 gnd.n6278 53.0052
R8967 gnd.n6281 gnd.n6280 53.0052
R8968 gnd.n6283 gnd.n6282 53.0052
R8969 gnd.n6285 gnd.n6284 53.0052
R8970 gnd.n6289 gnd.n6288 53.0052
R8971 gnd.n6291 gnd.n6290 53.0052
R8972 gnd.n6293 gnd.n6292 53.0052
R8973 gnd.n6295 gnd.n6294 53.0052
R8974 gnd.n6297 gnd.n6296 53.0052
R8975 gnd.n6299 gnd.n6298 53.0052
R8976 gnd.n6301 gnd.n6300 53.0052
R8977 gnd.n6303 gnd.n6302 53.0052
R8978 gnd.n6305 gnd.n6304 53.0052
R8979 gnd.n96 gnd.n95 53.0052
R8980 gnd.n94 gnd.n93 53.0052
R8981 gnd.n92 gnd.n91 53.0052
R8982 gnd.n90 gnd.n89 53.0052
R8983 gnd.n88 gnd.n87 53.0052
R8984 gnd.n86 gnd.n85 53.0052
R8985 gnd.n84 gnd.n83 53.0052
R8986 gnd.n82 gnd.n81 53.0052
R8987 gnd.n80 gnd.n79 53.0052
R8988 gnd.n37 gnd.n36 53.0052
R8989 gnd.n35 gnd.n34 53.0052
R8990 gnd.n33 gnd.n32 53.0052
R8991 gnd.n31 gnd.n30 53.0052
R8992 gnd.n29 gnd.n28 53.0052
R8993 gnd.n27 gnd.n26 53.0052
R8994 gnd.n25 gnd.n24 53.0052
R8995 gnd.n23 gnd.n22 53.0052
R8996 gnd.n21 gnd.n20 53.0052
R8997 gnd.n56 gnd.n55 53.0052
R8998 gnd.n54 gnd.n53 53.0052
R8999 gnd.n52 gnd.n51 53.0052
R9000 gnd.n50 gnd.n49 53.0052
R9001 gnd.n48 gnd.n47 53.0052
R9002 gnd.n46 gnd.n45 53.0052
R9003 gnd.n44 gnd.n43 53.0052
R9004 gnd.n42 gnd.n41 53.0052
R9005 gnd.n40 gnd.n39 53.0052
R9006 gnd.n76 gnd.n75 53.0052
R9007 gnd.n74 gnd.n73 53.0052
R9008 gnd.n72 gnd.n71 53.0052
R9009 gnd.n70 gnd.n69 53.0052
R9010 gnd.n68 gnd.n67 53.0052
R9011 gnd.n66 gnd.n65 53.0052
R9012 gnd.n64 gnd.n63 53.0052
R9013 gnd.n62 gnd.n61 53.0052
R9014 gnd.n60 gnd.n59 53.0052
R9015 gnd.n3709 gnd.n3708 52.4801
R9016 gnd.n5725 gnd.t41 52.3082
R9017 gnd.n5693 gnd.t404 52.3082
R9018 gnd.n5661 gnd.t397 52.3082
R9019 gnd.n5630 gnd.t409 52.3082
R9020 gnd.n5598 gnd.t17 52.3082
R9021 gnd.n5566 gnd.t36 52.3082
R9022 gnd.n5534 gnd.t30 52.3082
R9023 gnd.n5503 gnd.t11 52.3082
R9024 gnd.n5400 gnd.n1186 51.6227
R9025 gnd.n8003 gnd.n250 51.6227
R9026 gnd.n5555 gnd.n5523 51.4173
R9027 gnd.n5619 gnd.n5618 50.455
R9028 gnd.n5587 gnd.n5586 50.455
R9029 gnd.n5555 gnd.n5554 50.455
R9030 gnd.n6094 gnd.n6093 45.1884
R9031 gnd.n5475 gnd.n5474 45.1884
R9032 gnd.n3725 gnd.n3724 44.3322
R9033 gnd.n1676 gnd.n1675 44.3189
R9034 gnd.n3284 gnd.n3283 42.4732
R9035 gnd.n4412 gnd.n4411 42.4732
R9036 gnd.n4553 gnd.n4418 42.2793
R9037 gnd.n6106 gnd.n6094 42.2793
R9038 gnd.n5476 gnd.n5475 42.2793
R9039 gnd.n6391 gnd.n6389 42.2793
R9040 gnd.n5432 gnd.n5431 42.2793
R9041 gnd.n2552 gnd.n2551 42.2793
R9042 gnd.n4800 gnd.n1882 42.2793
R9043 gnd.n4763 gnd.n1905 42.2793
R9044 gnd.n4723 gnd.n1927 42.2793
R9045 gnd.n7886 gnd.n353 42.2793
R9046 gnd.n7928 gnd.n333 42.2793
R9047 gnd.n7970 gnd.n7969 42.2793
R9048 gnd.n451 gnd.n373 42.2793
R9049 gnd.n5364 gnd.n1209 42.2793
R9050 gnd.n5324 gnd.n1231 42.2793
R9051 gnd.n5284 gnd.n1253 42.2793
R9052 gnd.n2954 gnd.n2902 42.2793
R9053 gnd.n5066 gnd.n1614 42.2793
R9054 gnd.n2732 gnd.n2642 42.2793
R9055 gnd.n2683 gnd.n2655 42.2793
R9056 gnd.n1674 gnd.n1673 41.6274
R9057 gnd.n3719 gnd.n3718 41.6274
R9058 gnd.n1683 gnd.n1682 40.8975
R9059 gnd.n3722 gnd.n3721 40.8975
R9060 gnd.n1682 gnd.n1681 35.055
R9061 gnd.n1677 gnd.n1676 35.055
R9062 gnd.n3711 gnd.n3710 35.055
R9063 gnd.n3721 gnd.n3707 35.055
R9064 gnd.n7051 gnd.n7050 33.6191
R9065 gnd.n7050 gnd.n968 33.6191
R9066 gnd.n7044 gnd.n968 33.6191
R9067 gnd.n7044 gnd.n7043 33.6191
R9068 gnd.n7043 gnd.n7042 33.6191
R9069 gnd.n7042 gnd.n976 33.6191
R9070 gnd.n7036 gnd.n976 33.6191
R9071 gnd.n7036 gnd.n7035 33.6191
R9072 gnd.n7035 gnd.n7034 33.6191
R9073 gnd.n7034 gnd.n984 33.6191
R9074 gnd.n7028 gnd.n984 33.6191
R9075 gnd.n7028 gnd.n7027 33.6191
R9076 gnd.n7027 gnd.n7026 33.6191
R9077 gnd.n7026 gnd.n992 33.6191
R9078 gnd.n7020 gnd.n992 33.6191
R9079 gnd.n7020 gnd.n7019 33.6191
R9080 gnd.n7019 gnd.n7018 33.6191
R9081 gnd.n7018 gnd.n1000 33.6191
R9082 gnd.n7012 gnd.n1000 33.6191
R9083 gnd.n7012 gnd.n7011 33.6191
R9084 gnd.n7011 gnd.n7010 33.6191
R9085 gnd.n7010 gnd.n1008 33.6191
R9086 gnd.n7004 gnd.n1008 33.6191
R9087 gnd.n7004 gnd.n7003 33.6191
R9088 gnd.n7003 gnd.n7002 33.6191
R9089 gnd.n7002 gnd.n1016 33.6191
R9090 gnd.n6996 gnd.n1016 33.6191
R9091 gnd.n6996 gnd.n6995 33.6191
R9092 gnd.n6995 gnd.n6994 33.6191
R9093 gnd.n6994 gnd.n1024 33.6191
R9094 gnd.n6988 gnd.n1024 33.6191
R9095 gnd.n6988 gnd.n6987 33.6191
R9096 gnd.n6987 gnd.n6986 33.6191
R9097 gnd.n6986 gnd.n1032 33.6191
R9098 gnd.n6980 gnd.n1032 33.6191
R9099 gnd.n6980 gnd.n6979 33.6191
R9100 gnd.n6979 gnd.n6978 33.6191
R9101 gnd.n6978 gnd.n1040 33.6191
R9102 gnd.n6972 gnd.n1040 33.6191
R9103 gnd.n6972 gnd.n6971 33.6191
R9104 gnd.n6971 gnd.n6970 33.6191
R9105 gnd.n6970 gnd.n1048 33.6191
R9106 gnd.n6964 gnd.n1048 33.6191
R9107 gnd.n6964 gnd.n6963 33.6191
R9108 gnd.n6963 gnd.n6962 33.6191
R9109 gnd.n6962 gnd.n1056 33.6191
R9110 gnd.n6956 gnd.n1056 33.6191
R9111 gnd.n6956 gnd.n6955 33.6191
R9112 gnd.n6955 gnd.n6954 33.6191
R9113 gnd.n6954 gnd.n1064 33.6191
R9114 gnd.n6948 gnd.n1064 33.6191
R9115 gnd.n6948 gnd.n6947 33.6191
R9116 gnd.n6947 gnd.n6946 33.6191
R9117 gnd.n6946 gnd.n1072 33.6191
R9118 gnd.n6940 gnd.n1072 33.6191
R9119 gnd.n6940 gnd.n6939 33.6191
R9120 gnd.n6939 gnd.n6938 33.6191
R9121 gnd.n6938 gnd.n1080 33.6191
R9122 gnd.n6932 gnd.n1080 33.6191
R9123 gnd.n6932 gnd.n6931 33.6191
R9124 gnd.n6931 gnd.n6930 33.6191
R9125 gnd.n6930 gnd.n1088 33.6191
R9126 gnd.n6924 gnd.n1088 33.6191
R9127 gnd.n6924 gnd.n6923 33.6191
R9128 gnd.n6923 gnd.n6922 33.6191
R9129 gnd.n6922 gnd.n1096 33.6191
R9130 gnd.n6916 gnd.n1096 33.6191
R9131 gnd.n6916 gnd.n6915 33.6191
R9132 gnd.n6915 gnd.n6914 33.6191
R9133 gnd.n6914 gnd.n1104 33.6191
R9134 gnd.n6908 gnd.n1104 33.6191
R9135 gnd.n6908 gnd.n6907 33.6191
R9136 gnd.n6907 gnd.n6906 33.6191
R9137 gnd.n6906 gnd.n1112 33.6191
R9138 gnd.n6900 gnd.n1112 33.6191
R9139 gnd.n6900 gnd.n6899 33.6191
R9140 gnd.n6899 gnd.n6898 33.6191
R9141 gnd.n6898 gnd.n1120 33.6191
R9142 gnd.n6892 gnd.n1120 33.6191
R9143 gnd.n6892 gnd.n6891 33.6191
R9144 gnd.n6891 gnd.n6890 33.6191
R9145 gnd.n6890 gnd.n1128 33.6191
R9146 gnd.n6884 gnd.n1128 33.6191
R9147 gnd.n6156 gnd.n6052 31.8661
R9148 gnd.n6164 gnd.n6052 31.8661
R9149 gnd.n6172 gnd.n6046 31.8661
R9150 gnd.n6172 gnd.n6040 31.8661
R9151 gnd.n6180 gnd.n6040 31.8661
R9152 gnd.n6180 gnd.n6033 31.8661
R9153 gnd.n6188 gnd.n6033 31.8661
R9154 gnd.n6188 gnd.n6034 31.8661
R9155 gnd.n6432 gnd.n6019 31.8661
R9156 gnd.n5276 gnd.n1186 31.8661
R9157 gnd.n5270 gnd.n1270 31.8661
R9158 gnd.n5270 gnd.n1273 31.8661
R9159 gnd.n5264 gnd.n1273 31.8661
R9160 gnd.n5264 gnd.n1285 31.8661
R9161 gnd.n5258 gnd.n1295 31.8661
R9162 gnd.n5252 gnd.n1295 31.8661
R9163 gnd.n5246 gnd.n1311 31.8661
R9164 gnd.n5246 gnd.n1314 31.8661
R9165 gnd.n5240 gnd.n1323 31.8661
R9166 gnd.n5234 gnd.n1333 31.8661
R9167 gnd.n5228 gnd.n1333 31.8661
R9168 gnd.n5222 gnd.n1349 31.8661
R9169 gnd.n5222 gnd.n1352 31.8661
R9170 gnd.n5216 gnd.n1361 31.8661
R9171 gnd.n5210 gnd.n1371 31.8661
R9172 gnd.n5204 gnd.n1371 31.8661
R9173 gnd.n5198 gnd.n1386 31.8661
R9174 gnd.n5198 gnd.n1389 31.8661
R9175 gnd.n5192 gnd.n1399 31.8661
R9176 gnd.n3360 gnd.n1556 31.8661
R9177 gnd.n3353 gnd.n1567 31.8661
R9178 gnd.n3353 gnd.n3352 31.8661
R9179 gnd.n3373 gnd.n2542 31.8661
R9180 gnd.n3373 gnd.n2544 31.8661
R9181 gnd.n3381 gnd.n2529 31.8661
R9182 gnd.n3389 gnd.n2529 31.8661
R9183 gnd.n3389 gnd.n2522 31.8661
R9184 gnd.n3397 gnd.n2522 31.8661
R9185 gnd.n3405 gnd.n2515 31.8661
R9186 gnd.n3405 gnd.n2507 31.8661
R9187 gnd.n3413 gnd.n2507 31.8661
R9188 gnd.n3413 gnd.n2509 31.8661
R9189 gnd.n3421 gnd.n2492 31.8661
R9190 gnd.n3438 gnd.n2492 31.8661
R9191 gnd.n3438 gnd.n2494 31.8661
R9192 gnd.n4347 gnd.n2176 31.8661
R9193 gnd.n4347 gnd.n2169 31.8661
R9194 gnd.n4355 gnd.n2169 31.8661
R9195 gnd.n4363 gnd.n2163 31.8661
R9196 gnd.n4363 gnd.n2154 31.8661
R9197 gnd.n4371 gnd.n2154 31.8661
R9198 gnd.n4371 gnd.n2156 31.8661
R9199 gnd.n4379 gnd.n2142 31.8661
R9200 gnd.n4389 gnd.n2142 31.8661
R9201 gnd.n4389 gnd.n2135 31.8661
R9202 gnd.n4400 gnd.n2135 31.8661
R9203 gnd.n4845 gnd.n1809 31.8661
R9204 gnd.n4845 gnd.n4844 31.8661
R9205 gnd.n4838 gnd.n1820 31.8661
R9206 gnd.n4838 gnd.n4837 31.8661
R9207 gnd.n1934 gnd.n1859 31.8661
R9208 gnd.n8097 gnd.n107 31.8661
R9209 gnd.n8089 gnd.n122 31.8661
R9210 gnd.n8089 gnd.n125 31.8661
R9211 gnd.n8083 gnd.n136 31.8661
R9212 gnd.n8077 gnd.n136 31.8661
R9213 gnd.n8071 gnd.n151 31.8661
R9214 gnd.n8065 gnd.n161 31.8661
R9215 gnd.n8065 gnd.n164 31.8661
R9216 gnd.n8059 gnd.n173 31.8661
R9217 gnd.n8053 gnd.n173 31.8661
R9218 gnd.n8047 gnd.n189 31.8661
R9219 gnd.n8041 gnd.n199 31.8661
R9220 gnd.n8041 gnd.n202 31.8661
R9221 gnd.n8035 gnd.n211 31.8661
R9222 gnd.n8023 gnd.n228 31.8661
R9223 gnd.n8023 gnd.n231 31.8661
R9224 gnd.n8017 gnd.n231 31.8661
R9225 gnd.n8017 gnd.n241 31.8661
R9226 gnd.n8011 gnd.n250 31.8661
R9227 gnd.n5216 gnd.t240 30.9101
R9228 gnd.n8071 gnd.t230 30.9101
R9229 gnd.n3880 gnd.n3879 30.4395
R9230 gnd.n2475 gnd.n2471 30.4395
R9231 gnd.n5240 gnd.t222 30.2728
R9232 gnd.n8047 gnd.t333 30.2728
R9233 gnd.n5276 gnd.t98 28.3609
R9234 gnd.n8011 gnd.t83 28.3609
R9235 gnd.n3687 gnd.n2187 27.4049
R9236 gnd.n2494 gnd.t189 27.0862
R9237 gnd.t24 gnd.n2176 27.0862
R9238 gnd.n3283 gnd.n3282 25.7944
R9239 gnd.n4418 gnd.n4417 25.7944
R9240 gnd.n6389 gnd.n6388 25.7944
R9241 gnd.n5431 gnd.n5430 25.7944
R9242 gnd.n2551 gnd.n2550 25.7944
R9243 gnd.n1882 gnd.n1881 25.7944
R9244 gnd.n1905 gnd.n1904 25.7944
R9245 gnd.n1927 gnd.n1926 25.7944
R9246 gnd.n353 gnd.n352 25.7944
R9247 gnd.n333 gnd.n332 25.7944
R9248 gnd.n7969 gnd.n7968 25.7944
R9249 gnd.n373 gnd.n372 25.7944
R9250 gnd.n1209 gnd.n1208 25.7944
R9251 gnd.n1231 gnd.n1230 25.7944
R9252 gnd.n1253 gnd.n1252 25.7944
R9253 gnd.n2902 gnd.n2901 25.7944
R9254 gnd.n1614 gnd.n1613 25.7944
R9255 gnd.n2642 gnd.n2641 25.7944
R9256 gnd.n2655 gnd.n2654 25.7944
R9257 gnd.n4411 gnd.n4410 25.7944
R9258 gnd.n6433 gnd.n6009 24.8557
R9259 gnd.n6012 gnd.n6002 24.8557
R9260 gnd.n6463 gnd.n5995 24.8557
R9261 gnd.n6464 gnd.n5984 24.8557
R9262 gnd.n5987 gnd.n5975 24.8557
R9263 gnd.n6485 gnd.n5976 24.8557
R9264 gnd.n6506 gnd.n6505 24.8557
R9265 gnd.n5961 gnd.n5949 24.8557
R9266 gnd.n6516 gnd.n5950 24.8557
R9267 gnd.n6526 gnd.n5932 24.8557
R9268 gnd.n6537 gnd.n6536 24.8557
R9269 gnd.n6547 gnd.n5925 24.8557
R9270 gnd.n6556 gnd.n5917 24.8557
R9271 gnd.n6557 gnd.n5906 24.8557
R9272 gnd.n6568 gnd.n6567 24.8557
R9273 gnd.n6587 gnd.n5892 24.8557
R9274 gnd.n6599 gnd.n6598 24.8557
R9275 gnd.n6228 gnd.n5884 24.8557
R9276 gnd.n6609 gnd.n5874 24.8557
R9277 gnd.n6618 gnd.n5867 24.8557
R9278 gnd.n6629 gnd.n6628 24.8557
R9279 gnd.n5860 gnd.n5850 24.8557
R9280 gnd.n5843 gnd.n5837 24.8557
R9281 gnd.n6660 gnd.n6659 24.8557
R9282 gnd.n6670 gnd.n6669 24.8557
R9283 gnd.n5827 gnd.n5818 24.8557
R9284 gnd.n5809 gnd.n5808 24.8557
R9285 gnd.n6704 gnd.n5801 24.8557
R9286 gnd.n6717 gnd.n6716 24.8557
R9287 gnd.n6729 gnd.n5788 24.8557
R9288 gnd.n6749 gnd.n5774 24.8557
R9289 gnd.n6760 gnd.n6759 24.8557
R9290 gnd.n6779 gnd.n5489 24.8557
R9291 gnd.n5761 gnd.n5490 24.8557
R9292 gnd.n6876 gnd.n1145 24.8557
R9293 gnd.n2544 gnd.t102 24.537
R9294 gnd.n3421 gnd.t18 24.537
R9295 gnd.n4355 gnd.t399 24.537
R9296 gnd.t66 gnd.n1809 24.537
R9297 gnd.n3024 gnd.n2808 24.2183
R9298 gnd.n3040 gnd.n2797 24.2183
R9299 gnd.n2792 gnd.n2784 24.2183
R9300 gnd.n5185 gnd.n1412 24.2183
R9301 gnd.n3085 gnd.n1415 24.2183
R9302 gnd.n3093 gnd.n1426 24.2183
R9303 gnd.n5173 gnd.n1433 24.2183
R9304 gnd.n5167 gnd.n1443 24.2183
R9305 gnd.n5161 gnd.n1454 24.2183
R9306 gnd.n3142 gnd.n1457 24.2183
R9307 gnd.n3114 gnd.n1466 24.2183
R9308 gnd.n5149 gnd.n1474 24.2183
R9309 gnd.n5143 gnd.n1484 24.2183
R9310 gnd.n5137 gnd.n1495 24.2183
R9311 gnd.n3186 gnd.n1498 24.2183
R9312 gnd.n3193 gnd.n1507 24.2183
R9313 gnd.n5125 gnd.n1515 24.2183
R9314 gnd.n5119 gnd.n1525 24.2183
R9315 gnd.n3208 gnd.n1528 24.2183
R9316 gnd.n5113 gnd.n1536 24.2183
R9317 gnd.n3218 gnd.n1539 24.2183
R9318 gnd.n5107 gnd.n1546 24.2183
R9319 gnd.n3361 gnd.n1549 24.2183
R9320 gnd.n4716 gnd.n1936 24.2183
R9321 gnd.n4713 gnd.n1941 24.2183
R9322 gnd.n4573 gnd.n1950 24.2183
R9323 gnd.n4707 gnd.n1953 24.2183
R9324 gnd.n4579 gnd.n1961 24.2183
R9325 gnd.n4701 gnd.n1964 24.2183
R9326 gnd.n4695 gnd.n1975 24.2183
R9327 gnd.n4593 gnd.n1982 24.2183
R9328 gnd.n4601 gnd.n1992 24.2183
R9329 gnd.n4683 gnd.n1995 24.2183
R9330 gnd.n4677 gnd.n2005 24.2183
R9331 gnd.n4671 gnd.n2016 24.2183
R9332 gnd.n4624 gnd.n2023 24.2183
R9333 gnd.n4640 gnd.n2034 24.2183
R9334 gnd.n4659 gnd.n2037 24.2183
R9335 gnd.n2045 gnd.n542 24.2183
R9336 gnd.n7744 gnd.n532 24.2183
R9337 gnd.n7768 gnd.n534 24.2183
R9338 gnd.n7776 gnd.n515 24.2183
R9339 gnd.n7790 gnd.n510 24.2183
R9340 gnd.n7784 gnd.n502 24.2183
R9341 gnd.n7813 gnd.n500 24.2183
R9342 gnd.n7808 gnd.n491 24.2183
R9343 gnd.n3055 gnd.t291 23.8997
R9344 gnd.n3351 gnd.n2542 23.8997
R9345 gnd.n4844 gnd.n1812 23.8997
R9346 gnd.n522 gnd.t193 23.8997
R9347 gnd.n2409 gnd.n2408 23.855
R9348 gnd.n3813 gnd.n3812 23.855
R9349 gnd.n4981 gnd.n4980 23.855
R9350 gnd.n3705 gnd.n3704 23.855
R9351 gnd.n6454 gnd.t10 23.2624
R9352 gnd.t201 gnd.n1285 23.2624
R9353 gnd.t219 gnd.n1446 23.2624
R9354 gnd.n3201 gnd.t209 23.2624
R9355 gnd.n4587 gnd.t228 23.2624
R9356 gnd.t275 gnd.n4651 23.2624
R9357 gnd.n228 gnd.t226 23.2624
R9358 gnd.n6444 gnd.t87 22.6251
R9359 gnd.t211 gnd.n1323 22.6251
R9360 gnd.n3118 gnd.t285 22.6251
R9361 gnd.t304 gnd.n1487 22.6251
R9362 gnd.t195 gnd.n2002 22.6251
R9363 gnd.n4615 gnd.t199 22.6251
R9364 gnd.n189 gnd.t247 22.6251
R9365 gnd.t205 gnd.n1361 21.9878
R9366 gnd.n3099 gnd.t207 21.9878
R9367 gnd.n5045 gnd.n1630 21.9878
R9368 gnd.n7757 gnd.t272 21.9878
R9369 gnd.n151 gnd.t295 21.9878
R9370 gnd.t77 gnd.n1662 21.6691
R9371 gnd.n4086 gnd.n2393 21.6691
R9372 gnd.n4063 gnd.n4062 21.6691
R9373 gnd.n4056 gnd.n2359 21.6691
R9374 gnd.n4041 gnd.n2345 21.6691
R9375 gnd.n4004 gnd.n2310 21.6691
R9376 gnd.n3997 gnd.n2303 21.6691
R9377 gnd.n3988 gnd.n2296 21.6691
R9378 gnd.n3981 gnd.n2289 21.6691
R9379 gnd.n3942 gnd.n2248 21.6691
R9380 gnd.n3927 gnd.n2234 21.6691
R9381 gnd.n3920 gnd.n2228 21.6691
R9382 gnd.n3671 gnd.n2207 21.6691
R9383 gnd.n6423 gnd.t408 21.3504
R9384 gnd.n3046 gnd.t267 21.3504
R9385 gnd.n7803 gnd.t224 21.3504
R9386 gnd.n4079 gnd.n4078 21.0318
R9387 gnd.t26 gnd.n2378 21.0318
R9388 gnd.n4163 gnd.n2333 21.0318
R9389 gnd.n4171 gnd.n2323 21.0318
R9390 gnd.t391 gnd.n2317 21.0318
R9391 gnd.n3972 gnd.t9 21.0318
R9392 gnd.n3964 gnd.n2268 21.0318
R9393 gnd.n3593 gnd.n2269 21.0318
R9394 gnd.n3906 gnd.t405 21.0318
R9395 gnd.n4299 gnd.n2215 21.0318
R9396 gnd.n4307 gnd.n2206 21.0318
R9397 gnd.t3 gnd.n5795 20.7131
R9398 gnd.n1386 gnd.t253 20.7131
R9399 gnd.t213 gnd.n125 20.7131
R9400 gnd.n1396 gnd.t249 20.3945
R9401 gnd.n3885 gnd.t134 20.3945
R9402 gnd.n7721 gnd.t197 20.3945
R9403 gnd.n6884 gnd.n6883 20.1716
R9404 gnd.n6649 gnd.t406 20.0758
R9405 gnd.n1349 gnd.t237 20.0758
R9406 gnd.t255 gnd.n164 20.0758
R9407 gnd.n1671 gnd.t138 19.8005
R9408 gnd.n1671 gnd.t110 19.8005
R9409 gnd.n1670 gnd.t166 19.8005
R9410 gnd.n1670 gnd.t81 19.8005
R9411 gnd.n3716 gnd.t107 19.8005
R9412 gnd.n3716 gnd.t135 19.8005
R9413 gnd.n3715 gnd.t75 19.8005
R9414 gnd.n3715 gnd.t148 19.8005
R9415 gnd.n5099 gnd.n1567 19.7572
R9416 gnd.n3465 gnd.n3464 19.7572
R9417 gnd.n3476 gnd.n2379 19.7572
R9418 gnd.n4155 gnd.n2339 19.7572
R9419 gnd.n4179 gnd.n2316 19.7572
R9420 gnd.n3580 gnd.n2275 19.7572
R9421 gnd.n3601 gnd.n2262 19.7572
R9422 gnd.n4291 gnd.n2222 19.7572
R9423 gnd.n4315 gnd.n2199 19.7572
R9424 gnd.n4837 gnd.n4836 19.7572
R9425 gnd.n1667 gnd.n1666 19.5087
R9426 gnd.n1680 gnd.n1667 19.5087
R9427 gnd.n1678 gnd.n1669 19.5087
R9428 gnd.n3720 gnd.n3714 19.5087
R9429 gnd.t401 gnd.n5881 19.4385
R9430 gnd.n1311 gnd.t262 19.4385
R9431 gnd.n3397 gnd.t187 19.4385
R9432 gnd.n4379 gnd.t410 19.4385
R9433 gnd.t217 gnd.n202 19.4385
R9434 gnd.n3371 gnd.n2534 19.3944
R9435 gnd.n3383 gnd.n2534 19.3944
R9436 gnd.n3383 gnd.n2532 19.3944
R9437 gnd.n3387 gnd.n2532 19.3944
R9438 gnd.n3387 gnd.n2520 19.3944
R9439 gnd.n3399 gnd.n2520 19.3944
R9440 gnd.n3399 gnd.n2518 19.3944
R9441 gnd.n3403 gnd.n2518 19.3944
R9442 gnd.n3403 gnd.n2505 19.3944
R9443 gnd.n3415 gnd.n2505 19.3944
R9444 gnd.n3415 gnd.n2503 19.3944
R9445 gnd.n3419 gnd.n2503 19.3944
R9446 gnd.n3419 gnd.n2490 19.3944
R9447 gnd.n3440 gnd.n2490 19.3944
R9448 gnd.n3440 gnd.n2488 19.3944
R9449 gnd.n3444 gnd.n2488 19.3944
R9450 gnd.n3444 gnd.n2486 19.3944
R9451 gnd.n3448 gnd.n2486 19.3944
R9452 gnd.n3448 gnd.n2483 19.3944
R9453 gnd.n3453 gnd.n2483 19.3944
R9454 gnd.n3453 gnd.n2484 19.3944
R9455 gnd.n2484 gnd.n2389 19.3944
R9456 gnd.n4093 gnd.n2389 19.3944
R9457 gnd.n4093 gnd.n2387 19.3944
R9458 gnd.n4097 gnd.n2387 19.3944
R9459 gnd.n4097 gnd.n2376 19.3944
R9460 gnd.n4109 gnd.n2376 19.3944
R9461 gnd.n4109 gnd.n2374 19.3944
R9462 gnd.n4113 gnd.n2374 19.3944
R9463 gnd.n4113 gnd.n2363 19.3944
R9464 gnd.n4125 gnd.n2363 19.3944
R9465 gnd.n4125 gnd.n2361 19.3944
R9466 gnd.n4129 gnd.n2361 19.3944
R9467 gnd.n4129 gnd.n2350 19.3944
R9468 gnd.n4141 gnd.n2350 19.3944
R9469 gnd.n4141 gnd.n2348 19.3944
R9470 gnd.n4145 gnd.n2348 19.3944
R9471 gnd.n4145 gnd.n2337 19.3944
R9472 gnd.n4157 gnd.n2337 19.3944
R9473 gnd.n4157 gnd.n2335 19.3944
R9474 gnd.n4161 gnd.n2335 19.3944
R9475 gnd.n4161 gnd.n2321 19.3944
R9476 gnd.n4173 gnd.n2321 19.3944
R9477 gnd.n4173 gnd.n2319 19.3944
R9478 gnd.n4177 gnd.n2319 19.3944
R9479 gnd.n4177 gnd.n2307 19.3944
R9480 gnd.n4189 gnd.n2307 19.3944
R9481 gnd.n4189 gnd.n2305 19.3944
R9482 gnd.n4193 gnd.n2305 19.3944
R9483 gnd.n4193 gnd.n2293 19.3944
R9484 gnd.n4205 gnd.n2293 19.3944
R9485 gnd.n4205 gnd.n2291 19.3944
R9486 gnd.n4209 gnd.n2291 19.3944
R9487 gnd.n4209 gnd.n2280 19.3944
R9488 gnd.n4221 gnd.n2280 19.3944
R9489 gnd.n4221 gnd.n2278 19.3944
R9490 gnd.n4225 gnd.n2278 19.3944
R9491 gnd.n4225 gnd.n2266 19.3944
R9492 gnd.n4237 gnd.n2266 19.3944
R9493 gnd.n4237 gnd.n2264 19.3944
R9494 gnd.n4241 gnd.n2264 19.3944
R9495 gnd.n4241 gnd.n2252 19.3944
R9496 gnd.n4253 gnd.n2252 19.3944
R9497 gnd.n4253 gnd.n2250 19.3944
R9498 gnd.n4257 gnd.n2250 19.3944
R9499 gnd.n4257 gnd.n2239 19.3944
R9500 gnd.n4269 gnd.n2239 19.3944
R9501 gnd.n4269 gnd.n2237 19.3944
R9502 gnd.n4273 gnd.n2237 19.3944
R9503 gnd.n4273 gnd.n2226 19.3944
R9504 gnd.n4285 gnd.n2226 19.3944
R9505 gnd.n4285 gnd.n2224 19.3944
R9506 gnd.n4289 gnd.n2224 19.3944
R9507 gnd.n4289 gnd.n2211 19.3944
R9508 gnd.n4301 gnd.n2211 19.3944
R9509 gnd.n4301 gnd.n2209 19.3944
R9510 gnd.n4305 gnd.n2209 19.3944
R9511 gnd.n4305 gnd.n2197 19.3944
R9512 gnd.n4317 gnd.n2197 19.3944
R9513 gnd.n4317 gnd.n2195 19.3944
R9514 gnd.n4321 gnd.n2195 19.3944
R9515 gnd.n4321 gnd.n2185 19.3944
R9516 gnd.n4333 gnd.n2185 19.3944
R9517 gnd.n4333 gnd.n2183 19.3944
R9518 gnd.n4337 gnd.n2183 19.3944
R9519 gnd.n4337 gnd.n2173 19.3944
R9520 gnd.n4349 gnd.n2173 19.3944
R9521 gnd.n4349 gnd.n2171 19.3944
R9522 gnd.n4353 gnd.n2171 19.3944
R9523 gnd.n4353 gnd.n2160 19.3944
R9524 gnd.n4365 gnd.n2160 19.3944
R9525 gnd.n4365 gnd.n2158 19.3944
R9526 gnd.n4369 gnd.n2158 19.3944
R9527 gnd.n4369 gnd.n2147 19.3944
R9528 gnd.n4381 gnd.n2147 19.3944
R9529 gnd.n4381 gnd.n2144 19.3944
R9530 gnd.n4387 gnd.n2144 19.3944
R9531 gnd.n4387 gnd.n2145 19.3944
R9532 gnd.n2145 gnd.n2132 19.3944
R9533 gnd.n4403 gnd.n2132 19.3944
R9534 gnd.n4404 gnd.n4403 19.3944
R9535 gnd.n3287 gnd.n2547 19.3944
R9536 gnd.n3367 gnd.n2547 19.3944
R9537 gnd.n3368 gnd.n3367 19.3944
R9538 gnd.n3348 gnd.n3347 19.3944
R9539 gnd.n3347 gnd.n2634 19.3944
R9540 gnd.n3343 gnd.n2634 19.3944
R9541 gnd.n3343 gnd.n3342 19.3944
R9542 gnd.n3342 gnd.n3341 19.3944
R9543 gnd.n3341 gnd.n2639 19.3944
R9544 gnd.n3336 gnd.n2639 19.3944
R9545 gnd.n3336 gnd.n3335 19.3944
R9546 gnd.n3335 gnd.n3334 19.3944
R9547 gnd.n3334 gnd.n3230 19.3944
R9548 gnd.n3327 gnd.n3230 19.3944
R9549 gnd.n3327 gnd.n3326 19.3944
R9550 gnd.n3326 gnd.n3243 19.3944
R9551 gnd.n3319 gnd.n3243 19.3944
R9552 gnd.n3319 gnd.n3318 19.3944
R9553 gnd.n3318 gnd.n3251 19.3944
R9554 gnd.n3311 gnd.n3251 19.3944
R9555 gnd.n3311 gnd.n3310 19.3944
R9556 gnd.n3310 gnd.n3263 19.3944
R9557 gnd.n3303 gnd.n3263 19.3944
R9558 gnd.n3303 gnd.n3302 19.3944
R9559 gnd.n3302 gnd.n3271 19.3944
R9560 gnd.n3295 gnd.n3271 19.3944
R9561 gnd.n3295 gnd.n3294 19.3944
R9562 gnd.n4480 gnd.n4477 19.3944
R9563 gnd.n4480 gnd.n4441 19.3944
R9564 gnd.n4493 gnd.n4441 19.3944
R9565 gnd.n4496 gnd.n4493 19.3944
R9566 gnd.n4499 gnd.n4496 19.3944
R9567 gnd.n4499 gnd.n4434 19.3944
R9568 gnd.n4512 gnd.n4434 19.3944
R9569 gnd.n4515 gnd.n4512 19.3944
R9570 gnd.n4518 gnd.n4515 19.3944
R9571 gnd.n4518 gnd.n4427 19.3944
R9572 gnd.n4531 gnd.n4427 19.3944
R9573 gnd.n4534 gnd.n4531 19.3944
R9574 gnd.n4537 gnd.n4534 19.3944
R9575 gnd.n4537 gnd.n4419 19.3944
R9576 gnd.n4549 gnd.n4419 19.3944
R9577 gnd.n4552 gnd.n4549 19.3944
R9578 gnd.n6151 gnd.n6150 19.3944
R9579 gnd.n6150 gnd.n6060 19.3944
R9580 gnd.n6145 gnd.n6060 19.3944
R9581 gnd.n6145 gnd.n6144 19.3944
R9582 gnd.n6144 gnd.n6065 19.3944
R9583 gnd.n6139 gnd.n6065 19.3944
R9584 gnd.n6139 gnd.n6138 19.3944
R9585 gnd.n6138 gnd.n6137 19.3944
R9586 gnd.n6137 gnd.n6071 19.3944
R9587 gnd.n6131 gnd.n6071 19.3944
R9588 gnd.n6131 gnd.n6130 19.3944
R9589 gnd.n6130 gnd.n6129 19.3944
R9590 gnd.n6129 gnd.n6077 19.3944
R9591 gnd.n6123 gnd.n6077 19.3944
R9592 gnd.n6123 gnd.n6122 19.3944
R9593 gnd.n6122 gnd.n6121 19.3944
R9594 gnd.n6121 gnd.n6083 19.3944
R9595 gnd.n6115 gnd.n6083 19.3944
R9596 gnd.n6115 gnd.n6114 19.3944
R9597 gnd.n6114 gnd.n6113 19.3944
R9598 gnd.n6113 gnd.n6089 19.3944
R9599 gnd.n6107 gnd.n6089 19.3944
R9600 gnd.n6105 gnd.n6104 19.3944
R9601 gnd.n6104 gnd.n6099 19.3944
R9602 gnd.n6099 gnd.n6097 19.3944
R9603 gnd.n6796 gnd.n5478 19.3944
R9604 gnd.n6796 gnd.n6795 19.3944
R9605 gnd.n6795 gnd.n6794 19.3944
R9606 gnd.n6838 gnd.n6837 19.3944
R9607 gnd.n6837 gnd.n6836 19.3944
R9608 gnd.n6836 gnd.n5439 19.3944
R9609 gnd.n6831 gnd.n5439 19.3944
R9610 gnd.n6831 gnd.n6830 19.3944
R9611 gnd.n6830 gnd.n6829 19.3944
R9612 gnd.n6829 gnd.n5446 19.3944
R9613 gnd.n6824 gnd.n5446 19.3944
R9614 gnd.n6824 gnd.n6823 19.3944
R9615 gnd.n6823 gnd.n6822 19.3944
R9616 gnd.n6822 gnd.n5453 19.3944
R9617 gnd.n6817 gnd.n5453 19.3944
R9618 gnd.n6817 gnd.n6816 19.3944
R9619 gnd.n6816 gnd.n6815 19.3944
R9620 gnd.n6815 gnd.n5460 19.3944
R9621 gnd.n6810 gnd.n5460 19.3944
R9622 gnd.n6810 gnd.n6809 19.3944
R9623 gnd.n6809 gnd.n6808 19.3944
R9624 gnd.n6808 gnd.n5467 19.3944
R9625 gnd.n6803 gnd.n5467 19.3944
R9626 gnd.n6803 gnd.n6802 19.3944
R9627 gnd.n6802 gnd.n6801 19.3944
R9628 gnd.n6436 gnd.n6435 19.3944
R9629 gnd.n6436 gnd.n6000 19.3944
R9630 gnd.n6456 gnd.n6000 19.3944
R9631 gnd.n6456 gnd.n5992 19.3944
R9632 gnd.n6466 gnd.n5992 19.3944
R9633 gnd.n6467 gnd.n6466 19.3944
R9634 gnd.n6467 gnd.n5973 19.3944
R9635 gnd.n6487 gnd.n5973 19.3944
R9636 gnd.n6487 gnd.n5966 19.3944
R9637 gnd.n6497 gnd.n5966 19.3944
R9638 gnd.n6498 gnd.n6497 19.3944
R9639 gnd.n6498 gnd.n5947 19.3944
R9640 gnd.n6518 gnd.n5947 19.3944
R9641 gnd.n6518 gnd.n5940 19.3944
R9642 gnd.n6528 gnd.n5940 19.3944
R9643 gnd.n6529 gnd.n6528 19.3944
R9644 gnd.n6529 gnd.n5922 19.3944
R9645 gnd.n6549 gnd.n5922 19.3944
R9646 gnd.n6549 gnd.n5914 19.3944
R9647 gnd.n6559 gnd.n5914 19.3944
R9648 gnd.n6560 gnd.n6559 19.3944
R9649 gnd.n6560 gnd.n5897 19.3944
R9650 gnd.n6580 gnd.n5897 19.3944
R9651 gnd.n6580 gnd.n5889 19.3944
R9652 gnd.n6590 gnd.n5889 19.3944
R9653 gnd.n6591 gnd.n6590 19.3944
R9654 gnd.n6591 gnd.n5872 19.3944
R9655 gnd.n6611 gnd.n5872 19.3944
R9656 gnd.n6611 gnd.n5864 19.3944
R9657 gnd.n6621 gnd.n5864 19.3944
R9658 gnd.n6622 gnd.n6621 19.3944
R9659 gnd.n6622 gnd.n5848 19.3944
R9660 gnd.n6641 gnd.n5848 19.3944
R9661 gnd.n6641 gnd.n5833 19.3944
R9662 gnd.n6662 gnd.n5833 19.3944
R9663 gnd.n6663 gnd.n6662 19.3944
R9664 gnd.n6664 gnd.n6663 19.3944
R9665 gnd.n6664 gnd.n5817 19.3944
R9666 gnd.n5817 gnd.n5815 19.3944
R9667 gnd.n6687 gnd.n5815 19.3944
R9668 gnd.n6687 gnd.n5797 19.3944
R9669 gnd.n6713 gnd.n5797 19.3944
R9670 gnd.n6713 gnd.n6712 19.3944
R9671 gnd.n6712 gnd.n5786 19.3944
R9672 gnd.n6732 gnd.n5786 19.3944
R9673 gnd.n6732 gnd.n5770 19.3944
R9674 gnd.n6757 gnd.n5770 19.3944
R9675 gnd.n6757 gnd.n5750 19.3944
R9676 gnd.n6774 gnd.n5750 19.3944
R9677 gnd.n6774 gnd.n5752 19.3944
R9678 gnd.n5759 gnd.n5752 19.3944
R9679 gnd.n5759 gnd.n5758 19.3944
R9680 gnd.n5758 gnd.n5757 19.3944
R9681 gnd.n6419 gnd.n6418 19.3944
R9682 gnd.n6418 gnd.n6417 19.3944
R9683 gnd.n6417 gnd.n6416 19.3944
R9684 gnd.n6416 gnd.n6414 19.3944
R9685 gnd.n6414 gnd.n6411 19.3944
R9686 gnd.n6411 gnd.n6410 19.3944
R9687 gnd.n6410 gnd.n6407 19.3944
R9688 gnd.n6407 gnd.n6406 19.3944
R9689 gnd.n6406 gnd.n6403 19.3944
R9690 gnd.n6403 gnd.n6402 19.3944
R9691 gnd.n6402 gnd.n6399 19.3944
R9692 gnd.n6399 gnd.n6398 19.3944
R9693 gnd.n6398 gnd.n6395 19.3944
R9694 gnd.n6395 gnd.n6394 19.3944
R9695 gnd.n6446 gnd.n6007 19.3944
R9696 gnd.n6446 gnd.n6005 19.3944
R9697 gnd.n6452 gnd.n6005 19.3944
R9698 gnd.n6452 gnd.n6451 19.3944
R9699 gnd.n6451 gnd.n5982 19.3944
R9700 gnd.n6477 gnd.n5982 19.3944
R9701 gnd.n6477 gnd.n5980 19.3944
R9702 gnd.n6483 gnd.n5980 19.3944
R9703 gnd.n6483 gnd.n6482 19.3944
R9704 gnd.n6482 gnd.n5956 19.3944
R9705 gnd.n6508 gnd.n5956 19.3944
R9706 gnd.n6508 gnd.n5954 19.3944
R9707 gnd.n6514 gnd.n5954 19.3944
R9708 gnd.n6514 gnd.n6513 19.3944
R9709 gnd.n6513 gnd.n5930 19.3944
R9710 gnd.n6539 gnd.n5930 19.3944
R9711 gnd.n6539 gnd.n5928 19.3944
R9712 gnd.n6545 gnd.n5928 19.3944
R9713 gnd.n6545 gnd.n6544 19.3944
R9714 gnd.n6544 gnd.n5904 19.3944
R9715 gnd.n6570 gnd.n5904 19.3944
R9716 gnd.n6570 gnd.n5902 19.3944
R9717 gnd.n6576 gnd.n5902 19.3944
R9718 gnd.n6576 gnd.n6575 19.3944
R9719 gnd.n6575 gnd.n5879 19.3944
R9720 gnd.n6601 gnd.n5879 19.3944
R9721 gnd.n6601 gnd.n5877 19.3944
R9722 gnd.n6607 gnd.n5877 19.3944
R9723 gnd.n6607 gnd.n6606 19.3944
R9724 gnd.n6606 gnd.n5855 19.3944
R9725 gnd.n6631 gnd.n5855 19.3944
R9726 gnd.n6631 gnd.n5853 19.3944
R9727 gnd.n6637 gnd.n5853 19.3944
R9728 gnd.n6637 gnd.n6636 19.3944
R9729 gnd.n6636 gnd.n5823 19.3944
R9730 gnd.n6672 gnd.n5823 19.3944
R9731 gnd.n6672 gnd.n5821 19.3944
R9732 gnd.n6681 gnd.n5821 19.3944
R9733 gnd.n6681 gnd.n6680 19.3944
R9734 gnd.n6680 gnd.n6679 19.3944
R9735 gnd.n6679 gnd.n5793 19.3944
R9736 gnd.n6719 gnd.n5793 19.3944
R9737 gnd.n6719 gnd.n5791 19.3944
R9738 gnd.n6727 gnd.n5791 19.3944
R9739 gnd.n6727 gnd.n6726 19.3944
R9740 gnd.n6726 gnd.n6725 19.3944
R9741 gnd.n6725 gnd.n5766 19.3944
R9742 gnd.n6763 gnd.n5766 19.3944
R9743 gnd.n6763 gnd.n5764 19.3944
R9744 gnd.n6769 gnd.n5764 19.3944
R9745 gnd.n6769 gnd.n6768 19.3944
R9746 gnd.n6768 gnd.n5404 19.3944
R9747 gnd.n6873 gnd.n5404 19.3944
R9748 gnd.n6870 gnd.n6869 19.3944
R9749 gnd.n6869 gnd.n6868 19.3944
R9750 gnd.n6868 gnd.n5409 19.3944
R9751 gnd.n6863 gnd.n5409 19.3944
R9752 gnd.n6863 gnd.n6862 19.3944
R9753 gnd.n6862 gnd.n6861 19.3944
R9754 gnd.n6861 gnd.n5416 19.3944
R9755 gnd.n6856 gnd.n5416 19.3944
R9756 gnd.n6856 gnd.n6855 19.3944
R9757 gnd.n6855 gnd.n6854 19.3944
R9758 gnd.n6854 gnd.n5423 19.3944
R9759 gnd.n6849 gnd.n5423 19.3944
R9760 gnd.n6849 gnd.n6848 19.3944
R9761 gnd.n6848 gnd.n6847 19.3944
R9762 gnd.n6158 gnd.n6054 19.3944
R9763 gnd.n6162 gnd.n6054 19.3944
R9764 gnd.n6162 gnd.n6044 19.3944
R9765 gnd.n6174 gnd.n6044 19.3944
R9766 gnd.n6174 gnd.n6042 19.3944
R9767 gnd.n6178 gnd.n6042 19.3944
R9768 gnd.n6178 gnd.n6031 19.3944
R9769 gnd.n6190 gnd.n6031 19.3944
R9770 gnd.n6190 gnd.n6029 19.3944
R9771 gnd.n6361 gnd.n6029 19.3944
R9772 gnd.n6361 gnd.n6360 19.3944
R9773 gnd.n6360 gnd.n6359 19.3944
R9774 gnd.n6359 gnd.n6358 19.3944
R9775 gnd.n6358 gnd.n6356 19.3944
R9776 gnd.n6356 gnd.n6355 19.3944
R9777 gnd.n6355 gnd.n6351 19.3944
R9778 gnd.n6351 gnd.n6350 19.3944
R9779 gnd.n6350 gnd.n6349 19.3944
R9780 gnd.n6349 gnd.n6347 19.3944
R9781 gnd.n6347 gnd.n6346 19.3944
R9782 gnd.n6346 gnd.n6343 19.3944
R9783 gnd.n6343 gnd.n6342 19.3944
R9784 gnd.n6342 gnd.n6341 19.3944
R9785 gnd.n6341 gnd.n6339 19.3944
R9786 gnd.n6339 gnd.n6338 19.3944
R9787 gnd.n6338 gnd.n6335 19.3944
R9788 gnd.n6335 gnd.n6334 19.3944
R9789 gnd.n6334 gnd.n6333 19.3944
R9790 gnd.n6333 gnd.n6331 19.3944
R9791 gnd.n6247 gnd.n6212 19.3944
R9792 gnd.n6244 gnd.n6243 19.3944
R9793 gnd.n6240 gnd.n6239 19.3944
R9794 gnd.n6235 gnd.n6234 19.3944
R9795 gnd.n6234 gnd.n6233 19.3944
R9796 gnd.n6233 gnd.n6231 19.3944
R9797 gnd.n6231 gnd.n6230 19.3944
R9798 gnd.n6230 gnd.n6226 19.3944
R9799 gnd.n6226 gnd.n6225 19.3944
R9800 gnd.n6225 gnd.n6224 19.3944
R9801 gnd.n6224 gnd.n6222 19.3944
R9802 gnd.n6222 gnd.n5841 19.3944
R9803 gnd.n6651 gnd.n5841 19.3944
R9804 gnd.n6651 gnd.n5839 19.3944
R9805 gnd.n6657 gnd.n5839 19.3944
R9806 gnd.n6657 gnd.n6656 19.3944
R9807 gnd.n6656 gnd.n5806 19.3944
R9808 gnd.n6695 gnd.n5806 19.3944
R9809 gnd.n6695 gnd.n5804 19.3944
R9810 gnd.n6701 gnd.n5804 19.3944
R9811 gnd.n6701 gnd.n6700 19.3944
R9812 gnd.n6700 gnd.n5779 19.3944
R9813 gnd.n6740 gnd.n5779 19.3944
R9814 gnd.n6740 gnd.n5777 19.3944
R9815 gnd.n6746 gnd.n5777 19.3944
R9816 gnd.n6746 gnd.n6745 19.3944
R9817 gnd.n6745 gnd.n5486 19.3944
R9818 gnd.n6781 gnd.n5486 19.3944
R9819 gnd.n6781 gnd.n5484 19.3944
R9820 gnd.n6785 gnd.n5484 19.3944
R9821 gnd.n6788 gnd.n6785 19.3944
R9822 gnd.n6789 gnd.n6788 19.3944
R9823 gnd.n6154 gnd.n6050 19.3944
R9824 gnd.n6166 gnd.n6050 19.3944
R9825 gnd.n6166 gnd.n6048 19.3944
R9826 gnd.n6170 gnd.n6048 19.3944
R9827 gnd.n6170 gnd.n6038 19.3944
R9828 gnd.n6182 gnd.n6038 19.3944
R9829 gnd.n6182 gnd.n6036 19.3944
R9830 gnd.n6186 gnd.n6036 19.3944
R9831 gnd.n6186 gnd.n6025 19.3944
R9832 gnd.n6425 gnd.n6025 19.3944
R9833 gnd.n6425 gnd.n6022 19.3944
R9834 gnd.n6430 gnd.n6022 19.3944
R9835 gnd.n6430 gnd.n6015 19.3944
R9836 gnd.n6441 gnd.n6015 19.3944
R9837 gnd.n6441 gnd.n6440 19.3944
R9838 gnd.n6440 gnd.n5998 19.3944
R9839 gnd.n6461 gnd.n5998 19.3944
R9840 gnd.n6461 gnd.n5990 19.3944
R9841 gnd.n6472 gnd.n5990 19.3944
R9842 gnd.n6472 gnd.n6471 19.3944
R9843 gnd.n6471 gnd.n5971 19.3944
R9844 gnd.n6492 gnd.n5971 19.3944
R9845 gnd.n6492 gnd.n5964 19.3944
R9846 gnd.n6503 gnd.n5964 19.3944
R9847 gnd.n6503 gnd.n6502 19.3944
R9848 gnd.n6502 gnd.n5945 19.3944
R9849 gnd.n6523 gnd.n5945 19.3944
R9850 gnd.n6523 gnd.n5938 19.3944
R9851 gnd.n6534 gnd.n5938 19.3944
R9852 gnd.n6534 gnd.n6533 19.3944
R9853 gnd.n6533 gnd.n5920 19.3944
R9854 gnd.n6554 gnd.n5920 19.3944
R9855 gnd.n6554 gnd.n5912 19.3944
R9856 gnd.n6565 gnd.n5912 19.3944
R9857 gnd.n6565 gnd.n6564 19.3944
R9858 gnd.n6564 gnd.n5895 19.3944
R9859 gnd.n6585 gnd.n5895 19.3944
R9860 gnd.n6585 gnd.n5887 19.3944
R9861 gnd.n6596 gnd.n5887 19.3944
R9862 gnd.n6596 gnd.n6595 19.3944
R9863 gnd.n6595 gnd.n5870 19.3944
R9864 gnd.n6616 gnd.n5870 19.3944
R9865 gnd.n6616 gnd.n5862 19.3944
R9866 gnd.n6626 gnd.n5862 19.3944
R9867 gnd.n6626 gnd.n5846 19.3944
R9868 gnd.n6647 gnd.n5846 19.3944
R9869 gnd.n6647 gnd.n6646 19.3944
R9870 gnd.n6646 gnd.n5829 19.3944
R9871 gnd.n6667 gnd.n5829 19.3944
R9872 gnd.n6667 gnd.n5811 19.3944
R9873 gnd.n6691 gnd.n5811 19.3944
R9874 gnd.n6691 gnd.n6690 19.3944
R9875 gnd.n6690 gnd.n5799 19.3944
R9876 gnd.n6707 gnd.n5799 19.3944
R9877 gnd.n6707 gnd.n5782 19.3944
R9878 gnd.n6736 gnd.n5782 19.3944
R9879 gnd.n6736 gnd.n6735 19.3944
R9880 gnd.n6735 gnd.n5772 19.3944
R9881 gnd.n6752 gnd.n5772 19.3944
R9882 gnd.n6752 gnd.n5492 19.3944
R9883 gnd.n6777 gnd.n5492 19.3944
R9884 gnd.n6777 gnd.n1140 19.3944
R9885 gnd.n6880 gnd.n1140 19.3944
R9886 gnd.n6880 gnd.n6879 19.3944
R9887 gnd.n6879 gnd.n6878 19.3944
R9888 gnd.n3331 gnd.n3233 19.3944
R9889 gnd.n3331 gnd.n3330 19.3944
R9890 gnd.n3330 gnd.n3237 19.3944
R9891 gnd.n3323 gnd.n3237 19.3944
R9892 gnd.n3323 gnd.n3322 19.3944
R9893 gnd.n3322 gnd.n3247 19.3944
R9894 gnd.n3315 gnd.n3247 19.3944
R9895 gnd.n3315 gnd.n3314 19.3944
R9896 gnd.n3314 gnd.n3257 19.3944
R9897 gnd.n3307 gnd.n3257 19.3944
R9898 gnd.n3307 gnd.n3306 19.3944
R9899 gnd.n3306 gnd.n3267 19.3944
R9900 gnd.n3299 gnd.n3267 19.3944
R9901 gnd.n3299 gnd.n3298 19.3944
R9902 gnd.n3298 gnd.n3277 19.3944
R9903 gnd.n3291 gnd.n3277 19.3944
R9904 gnd.n2822 gnd.n2821 19.3944
R9905 gnd.n2821 gnd.n2820 19.3944
R9906 gnd.n2820 gnd.n2817 19.3944
R9907 gnd.n2817 gnd.n2816 19.3944
R9908 gnd.n2816 gnd.n2782 19.3944
R9909 gnd.n3058 gnd.n2782 19.3944
R9910 gnd.n3058 gnd.n2780 19.3944
R9911 gnd.n3082 gnd.n2780 19.3944
R9912 gnd.n3082 gnd.n3081 19.3944
R9913 gnd.n3081 gnd.n3080 19.3944
R9914 gnd.n3080 gnd.n3064 19.3944
R9915 gnd.n3076 gnd.n3064 19.3944
R9916 gnd.n3076 gnd.n3075 19.3944
R9917 gnd.n3075 gnd.n3074 19.3944
R9918 gnd.n3074 gnd.n3072 19.3944
R9919 gnd.n3072 gnd.n2757 19.3944
R9920 gnd.n2757 gnd.n2755 19.3944
R9921 gnd.n3147 gnd.n2755 19.3944
R9922 gnd.n3147 gnd.n2753 19.3944
R9923 gnd.n3151 gnd.n2753 19.3944
R9924 gnd.n3151 gnd.n2751 19.3944
R9925 gnd.n3155 gnd.n2751 19.3944
R9926 gnd.n3155 gnd.n2749 19.3944
R9927 gnd.n3183 gnd.n2749 19.3944
R9928 gnd.n3183 gnd.n3182 19.3944
R9929 gnd.n3182 gnd.n3181 19.3944
R9930 gnd.n3181 gnd.n3161 19.3944
R9931 gnd.n3177 gnd.n3161 19.3944
R9932 gnd.n3177 gnd.n3176 19.3944
R9933 gnd.n3176 gnd.n3175 19.3944
R9934 gnd.n3175 gnd.n3167 19.3944
R9935 gnd.n3171 gnd.n3167 19.3944
R9936 gnd.n3171 gnd.n2557 19.3944
R9937 gnd.n3358 gnd.n2557 19.3944
R9938 gnd.n3358 gnd.n3357 19.3944
R9939 gnd.n3357 gnd.n3356 19.3944
R9940 gnd.n3356 gnd.n2561 19.3944
R9941 gnd.n2564 gnd.n2561 19.3944
R9942 gnd.n2564 gnd.n2540 19.3944
R9943 gnd.n3375 gnd.n2540 19.3944
R9944 gnd.n3375 gnd.n2538 19.3944
R9945 gnd.n3379 gnd.n2538 19.3944
R9946 gnd.n3379 gnd.n2527 19.3944
R9947 gnd.n3391 gnd.n2527 19.3944
R9948 gnd.n3391 gnd.n2525 19.3944
R9949 gnd.n3395 gnd.n2525 19.3944
R9950 gnd.n3395 gnd.n2513 19.3944
R9951 gnd.n3407 gnd.n2513 19.3944
R9952 gnd.n3407 gnd.n2511 19.3944
R9953 gnd.n3411 gnd.n2511 19.3944
R9954 gnd.n3411 gnd.n2499 19.3944
R9955 gnd.n3423 gnd.n2499 19.3944
R9956 gnd.n3423 gnd.n2497 19.3944
R9957 gnd.n3436 gnd.n2497 19.3944
R9958 gnd.n3436 gnd.n3435 19.3944
R9959 gnd.n3435 gnd.n3434 19.3944
R9960 gnd.n3434 gnd.n3431 19.3944
R9961 gnd.n3431 gnd.n1695 19.3944
R9962 gnd.n4972 gnd.n1695 19.3944
R9963 gnd.n4972 gnd.n4971 19.3944
R9964 gnd.n4971 gnd.n4970 19.3944
R9965 gnd.n4970 gnd.n1699 19.3944
R9966 gnd.n4089 gnd.n1699 19.3944
R9967 gnd.n4089 gnd.n2383 19.3944
R9968 gnd.n4101 gnd.n2383 19.3944
R9969 gnd.n4101 gnd.n2381 19.3944
R9970 gnd.n4105 gnd.n2381 19.3944
R9971 gnd.n4105 gnd.n2369 19.3944
R9972 gnd.n4117 gnd.n2369 19.3944
R9973 gnd.n4117 gnd.n2367 19.3944
R9974 gnd.n4121 gnd.n2367 19.3944
R9975 gnd.n4121 gnd.n2357 19.3944
R9976 gnd.n4133 gnd.n2357 19.3944
R9977 gnd.n4133 gnd.n2355 19.3944
R9978 gnd.n4137 gnd.n2355 19.3944
R9979 gnd.n4137 gnd.n2343 19.3944
R9980 gnd.n4149 gnd.n2343 19.3944
R9981 gnd.n4149 gnd.n2341 19.3944
R9982 gnd.n4153 gnd.n2341 19.3944
R9983 gnd.n4153 gnd.n2328 19.3944
R9984 gnd.n4165 gnd.n2328 19.3944
R9985 gnd.n4165 gnd.n2326 19.3944
R9986 gnd.n4169 gnd.n2326 19.3944
R9987 gnd.n4169 gnd.n2314 19.3944
R9988 gnd.n4181 gnd.n2314 19.3944
R9989 gnd.n4181 gnd.n2312 19.3944
R9990 gnd.n4185 gnd.n2312 19.3944
R9991 gnd.n4185 gnd.n2300 19.3944
R9992 gnd.n4197 gnd.n2300 19.3944
R9993 gnd.n4197 gnd.n2298 19.3944
R9994 gnd.n4201 gnd.n2298 19.3944
R9995 gnd.n4201 gnd.n2287 19.3944
R9996 gnd.n4213 gnd.n2287 19.3944
R9997 gnd.n4213 gnd.n2285 19.3944
R9998 gnd.n4217 gnd.n2285 19.3944
R9999 gnd.n4217 gnd.n2273 19.3944
R10000 gnd.n4229 gnd.n2273 19.3944
R10001 gnd.n4229 gnd.n2271 19.3944
R10002 gnd.n4233 gnd.n2271 19.3944
R10003 gnd.n4233 gnd.n2259 19.3944
R10004 gnd.n4245 gnd.n2259 19.3944
R10005 gnd.n4245 gnd.n2257 19.3944
R10006 gnd.n4249 gnd.n2257 19.3944
R10007 gnd.n4249 gnd.n2246 19.3944
R10008 gnd.n4261 gnd.n2246 19.3944
R10009 gnd.n4261 gnd.n2244 19.3944
R10010 gnd.n4265 gnd.n2244 19.3944
R10011 gnd.n4265 gnd.n2232 19.3944
R10012 gnd.n4277 gnd.n2232 19.3944
R10013 gnd.n4277 gnd.n2230 19.3944
R10014 gnd.n4281 gnd.n2230 19.3944
R10015 gnd.n4281 gnd.n2219 19.3944
R10016 gnd.n4293 gnd.n2219 19.3944
R10017 gnd.n4293 gnd.n2217 19.3944
R10018 gnd.n4297 gnd.n2217 19.3944
R10019 gnd.n4297 gnd.n2204 19.3944
R10020 gnd.n4309 gnd.n2204 19.3944
R10021 gnd.n4309 gnd.n2202 19.3944
R10022 gnd.n4313 gnd.n2202 19.3944
R10023 gnd.n4313 gnd.n2191 19.3944
R10024 gnd.n4325 gnd.n2191 19.3944
R10025 gnd.n4325 gnd.n2189 19.3944
R10026 gnd.n4329 gnd.n2189 19.3944
R10027 gnd.n4329 gnd.n2180 19.3944
R10028 gnd.n4341 gnd.n2180 19.3944
R10029 gnd.n4341 gnd.n2178 19.3944
R10030 gnd.n4345 gnd.n2178 19.3944
R10031 gnd.n4345 gnd.n2167 19.3944
R10032 gnd.n4357 gnd.n2167 19.3944
R10033 gnd.n4357 gnd.n2165 19.3944
R10034 gnd.n4361 gnd.n2165 19.3944
R10035 gnd.n4361 gnd.n2152 19.3944
R10036 gnd.n4373 gnd.n2152 19.3944
R10037 gnd.n4373 gnd.n2150 19.3944
R10038 gnd.n4377 gnd.n2150 19.3944
R10039 gnd.n4377 gnd.n2140 19.3944
R10040 gnd.n4391 gnd.n2140 19.3944
R10041 gnd.n4391 gnd.n2138 19.3944
R10042 gnd.n4398 gnd.n2138 19.3944
R10043 gnd.n4398 gnd.n4397 19.3944
R10044 gnd.n4397 gnd.n1814 19.3944
R10045 gnd.n4842 gnd.n1814 19.3944
R10046 gnd.n4842 gnd.n4841 19.3944
R10047 gnd.n4841 gnd.n4840 19.3944
R10048 gnd.n4840 gnd.n1818 19.3944
R10049 gnd.n2076 gnd.n1818 19.3944
R10050 gnd.n2079 gnd.n2076 19.3944
R10051 gnd.n2079 gnd.n2073 19.3944
R10052 gnd.n2083 gnd.n2073 19.3944
R10053 gnd.n2083 gnd.n2071 19.3944
R10054 gnd.n2087 gnd.n2071 19.3944
R10055 gnd.n2087 gnd.n2069 19.3944
R10056 gnd.n2091 gnd.n2069 19.3944
R10057 gnd.n2091 gnd.n2067 19.3944
R10058 gnd.n2095 gnd.n2067 19.3944
R10059 gnd.n2095 gnd.n2065 19.3944
R10060 gnd.n2118 gnd.n2065 19.3944
R10061 gnd.n2118 gnd.n2117 19.3944
R10062 gnd.n2117 gnd.n2116 19.3944
R10063 gnd.n2116 gnd.n2101 19.3944
R10064 gnd.n2112 gnd.n2101 19.3944
R10065 gnd.n2112 gnd.n2111 19.3944
R10066 gnd.n2111 gnd.n2110 19.3944
R10067 gnd.n2110 gnd.n2108 19.3944
R10068 gnd.n2108 gnd.n2049 19.3944
R10069 gnd.n4644 gnd.n2049 19.3944
R10070 gnd.n4644 gnd.n2047 19.3944
R10071 gnd.n4649 gnd.n2047 19.3944
R10072 gnd.n4649 gnd.n553 19.3944
R10073 gnd.n7741 gnd.n553 19.3944
R10074 gnd.n7741 gnd.n7740 19.3944
R10075 gnd.n7740 gnd.n7739 19.3944
R10076 gnd.n7739 gnd.n557 19.3944
R10077 gnd.n7735 gnd.n557 19.3944
R10078 gnd.n7735 gnd.n7734 19.3944
R10079 gnd.n7734 gnd.n561 19.3944
R10080 gnd.n7730 gnd.n561 19.3944
R10081 gnd.n7730 gnd.n563 19.3944
R10082 gnd.n7726 gnd.n563 19.3944
R10083 gnd.n7726 gnd.n7725 19.3944
R10084 gnd.n7725 gnd.n7724 19.3944
R10085 gnd.n7509 gnd.n692 19.3944
R10086 gnd.n7515 gnd.n692 19.3944
R10087 gnd.n7515 gnd.n690 19.3944
R10088 gnd.n7519 gnd.n690 19.3944
R10089 gnd.n7519 gnd.n686 19.3944
R10090 gnd.n7525 gnd.n686 19.3944
R10091 gnd.n7525 gnd.n684 19.3944
R10092 gnd.n7529 gnd.n684 19.3944
R10093 gnd.n7529 gnd.n680 19.3944
R10094 gnd.n7535 gnd.n680 19.3944
R10095 gnd.n7535 gnd.n678 19.3944
R10096 gnd.n7539 gnd.n678 19.3944
R10097 gnd.n7539 gnd.n674 19.3944
R10098 gnd.n7545 gnd.n674 19.3944
R10099 gnd.n7545 gnd.n672 19.3944
R10100 gnd.n7549 gnd.n672 19.3944
R10101 gnd.n7549 gnd.n668 19.3944
R10102 gnd.n7555 gnd.n668 19.3944
R10103 gnd.n7555 gnd.n666 19.3944
R10104 gnd.n7559 gnd.n666 19.3944
R10105 gnd.n7559 gnd.n662 19.3944
R10106 gnd.n7565 gnd.n662 19.3944
R10107 gnd.n7565 gnd.n660 19.3944
R10108 gnd.n7569 gnd.n660 19.3944
R10109 gnd.n7569 gnd.n656 19.3944
R10110 gnd.n7575 gnd.n656 19.3944
R10111 gnd.n7575 gnd.n654 19.3944
R10112 gnd.n7579 gnd.n654 19.3944
R10113 gnd.n7579 gnd.n650 19.3944
R10114 gnd.n7585 gnd.n650 19.3944
R10115 gnd.n7585 gnd.n648 19.3944
R10116 gnd.n7589 gnd.n648 19.3944
R10117 gnd.n7589 gnd.n644 19.3944
R10118 gnd.n7595 gnd.n644 19.3944
R10119 gnd.n7595 gnd.n642 19.3944
R10120 gnd.n7599 gnd.n642 19.3944
R10121 gnd.n7599 gnd.n638 19.3944
R10122 gnd.n7605 gnd.n638 19.3944
R10123 gnd.n7605 gnd.n636 19.3944
R10124 gnd.n7609 gnd.n636 19.3944
R10125 gnd.n7609 gnd.n632 19.3944
R10126 gnd.n7615 gnd.n632 19.3944
R10127 gnd.n7615 gnd.n630 19.3944
R10128 gnd.n7619 gnd.n630 19.3944
R10129 gnd.n7619 gnd.n626 19.3944
R10130 gnd.n7625 gnd.n626 19.3944
R10131 gnd.n7625 gnd.n624 19.3944
R10132 gnd.n7629 gnd.n624 19.3944
R10133 gnd.n7629 gnd.n620 19.3944
R10134 gnd.n7635 gnd.n620 19.3944
R10135 gnd.n7635 gnd.n618 19.3944
R10136 gnd.n7639 gnd.n618 19.3944
R10137 gnd.n7639 gnd.n614 19.3944
R10138 gnd.n7645 gnd.n614 19.3944
R10139 gnd.n7645 gnd.n612 19.3944
R10140 gnd.n7649 gnd.n612 19.3944
R10141 gnd.n7649 gnd.n608 19.3944
R10142 gnd.n7655 gnd.n608 19.3944
R10143 gnd.n7655 gnd.n606 19.3944
R10144 gnd.n7659 gnd.n606 19.3944
R10145 gnd.n7659 gnd.n602 19.3944
R10146 gnd.n7665 gnd.n602 19.3944
R10147 gnd.n7665 gnd.n600 19.3944
R10148 gnd.n7669 gnd.n600 19.3944
R10149 gnd.n7669 gnd.n596 19.3944
R10150 gnd.n7675 gnd.n596 19.3944
R10151 gnd.n7675 gnd.n594 19.3944
R10152 gnd.n7679 gnd.n594 19.3944
R10153 gnd.n7679 gnd.n590 19.3944
R10154 gnd.n7685 gnd.n590 19.3944
R10155 gnd.n7685 gnd.n588 19.3944
R10156 gnd.n7689 gnd.n588 19.3944
R10157 gnd.n7689 gnd.n584 19.3944
R10158 gnd.n7695 gnd.n584 19.3944
R10159 gnd.n7695 gnd.n582 19.3944
R10160 gnd.n7699 gnd.n582 19.3944
R10161 gnd.n7699 gnd.n578 19.3944
R10162 gnd.n7705 gnd.n578 19.3944
R10163 gnd.n7705 gnd.n576 19.3944
R10164 gnd.n7709 gnd.n576 19.3944
R10165 gnd.n7709 gnd.n572 19.3944
R10166 gnd.n7716 gnd.n572 19.3944
R10167 gnd.n7716 gnd.n570 19.3944
R10168 gnd.n7720 gnd.n570 19.3944
R10169 gnd.n7054 gnd.n965 19.3944
R10170 gnd.n7058 gnd.n965 19.3944
R10171 gnd.n7058 gnd.n961 19.3944
R10172 gnd.n7064 gnd.n961 19.3944
R10173 gnd.n7064 gnd.n959 19.3944
R10174 gnd.n7068 gnd.n959 19.3944
R10175 gnd.n7068 gnd.n955 19.3944
R10176 gnd.n7074 gnd.n955 19.3944
R10177 gnd.n7074 gnd.n953 19.3944
R10178 gnd.n7078 gnd.n953 19.3944
R10179 gnd.n7078 gnd.n949 19.3944
R10180 gnd.n7084 gnd.n949 19.3944
R10181 gnd.n7084 gnd.n947 19.3944
R10182 gnd.n7088 gnd.n947 19.3944
R10183 gnd.n7088 gnd.n943 19.3944
R10184 gnd.n7094 gnd.n943 19.3944
R10185 gnd.n7094 gnd.n941 19.3944
R10186 gnd.n7098 gnd.n941 19.3944
R10187 gnd.n7098 gnd.n937 19.3944
R10188 gnd.n7104 gnd.n937 19.3944
R10189 gnd.n7104 gnd.n935 19.3944
R10190 gnd.n7108 gnd.n935 19.3944
R10191 gnd.n7108 gnd.n931 19.3944
R10192 gnd.n7114 gnd.n931 19.3944
R10193 gnd.n7114 gnd.n929 19.3944
R10194 gnd.n7118 gnd.n929 19.3944
R10195 gnd.n7118 gnd.n925 19.3944
R10196 gnd.n7124 gnd.n925 19.3944
R10197 gnd.n7124 gnd.n923 19.3944
R10198 gnd.n7128 gnd.n923 19.3944
R10199 gnd.n7128 gnd.n919 19.3944
R10200 gnd.n7134 gnd.n919 19.3944
R10201 gnd.n7134 gnd.n917 19.3944
R10202 gnd.n7138 gnd.n917 19.3944
R10203 gnd.n7138 gnd.n913 19.3944
R10204 gnd.n7144 gnd.n913 19.3944
R10205 gnd.n7144 gnd.n911 19.3944
R10206 gnd.n7148 gnd.n911 19.3944
R10207 gnd.n7148 gnd.n907 19.3944
R10208 gnd.n7154 gnd.n907 19.3944
R10209 gnd.n7154 gnd.n905 19.3944
R10210 gnd.n7158 gnd.n905 19.3944
R10211 gnd.n7158 gnd.n901 19.3944
R10212 gnd.n7164 gnd.n901 19.3944
R10213 gnd.n7164 gnd.n899 19.3944
R10214 gnd.n7168 gnd.n899 19.3944
R10215 gnd.n7168 gnd.n895 19.3944
R10216 gnd.n7174 gnd.n895 19.3944
R10217 gnd.n7174 gnd.n893 19.3944
R10218 gnd.n7178 gnd.n893 19.3944
R10219 gnd.n7178 gnd.n889 19.3944
R10220 gnd.n7184 gnd.n889 19.3944
R10221 gnd.n7184 gnd.n887 19.3944
R10222 gnd.n7188 gnd.n887 19.3944
R10223 gnd.n7188 gnd.n883 19.3944
R10224 gnd.n7194 gnd.n883 19.3944
R10225 gnd.n7194 gnd.n881 19.3944
R10226 gnd.n7198 gnd.n881 19.3944
R10227 gnd.n7198 gnd.n877 19.3944
R10228 gnd.n7204 gnd.n877 19.3944
R10229 gnd.n7204 gnd.n875 19.3944
R10230 gnd.n7208 gnd.n875 19.3944
R10231 gnd.n7208 gnd.n871 19.3944
R10232 gnd.n7214 gnd.n871 19.3944
R10233 gnd.n7214 gnd.n869 19.3944
R10234 gnd.n7218 gnd.n869 19.3944
R10235 gnd.n7218 gnd.n865 19.3944
R10236 gnd.n7224 gnd.n865 19.3944
R10237 gnd.n7224 gnd.n863 19.3944
R10238 gnd.n7228 gnd.n863 19.3944
R10239 gnd.n7228 gnd.n859 19.3944
R10240 gnd.n7234 gnd.n859 19.3944
R10241 gnd.n7234 gnd.n857 19.3944
R10242 gnd.n7238 gnd.n857 19.3944
R10243 gnd.n7238 gnd.n853 19.3944
R10244 gnd.n7244 gnd.n853 19.3944
R10245 gnd.n7244 gnd.n851 19.3944
R10246 gnd.n7248 gnd.n851 19.3944
R10247 gnd.n7248 gnd.n847 19.3944
R10248 gnd.n7254 gnd.n847 19.3944
R10249 gnd.n7254 gnd.n845 19.3944
R10250 gnd.n7258 gnd.n845 19.3944
R10251 gnd.n7258 gnd.n841 19.3944
R10252 gnd.n7264 gnd.n841 19.3944
R10253 gnd.n7264 gnd.n839 19.3944
R10254 gnd.n7268 gnd.n839 19.3944
R10255 gnd.n7268 gnd.n835 19.3944
R10256 gnd.n7274 gnd.n835 19.3944
R10257 gnd.n7274 gnd.n833 19.3944
R10258 gnd.n7278 gnd.n833 19.3944
R10259 gnd.n7278 gnd.n829 19.3944
R10260 gnd.n7284 gnd.n829 19.3944
R10261 gnd.n7284 gnd.n827 19.3944
R10262 gnd.n7288 gnd.n827 19.3944
R10263 gnd.n7288 gnd.n823 19.3944
R10264 gnd.n7294 gnd.n823 19.3944
R10265 gnd.n7294 gnd.n821 19.3944
R10266 gnd.n7298 gnd.n821 19.3944
R10267 gnd.n7298 gnd.n817 19.3944
R10268 gnd.n7304 gnd.n817 19.3944
R10269 gnd.n7304 gnd.n815 19.3944
R10270 gnd.n7308 gnd.n815 19.3944
R10271 gnd.n7308 gnd.n811 19.3944
R10272 gnd.n7314 gnd.n811 19.3944
R10273 gnd.n7314 gnd.n809 19.3944
R10274 gnd.n7318 gnd.n809 19.3944
R10275 gnd.n7318 gnd.n805 19.3944
R10276 gnd.n7324 gnd.n805 19.3944
R10277 gnd.n7324 gnd.n803 19.3944
R10278 gnd.n7328 gnd.n803 19.3944
R10279 gnd.n7328 gnd.n799 19.3944
R10280 gnd.n7334 gnd.n799 19.3944
R10281 gnd.n7334 gnd.n797 19.3944
R10282 gnd.n7338 gnd.n797 19.3944
R10283 gnd.n7338 gnd.n793 19.3944
R10284 gnd.n7344 gnd.n793 19.3944
R10285 gnd.n7344 gnd.n791 19.3944
R10286 gnd.n7348 gnd.n791 19.3944
R10287 gnd.n7348 gnd.n787 19.3944
R10288 gnd.n7354 gnd.n787 19.3944
R10289 gnd.n7354 gnd.n785 19.3944
R10290 gnd.n7358 gnd.n785 19.3944
R10291 gnd.n7358 gnd.n781 19.3944
R10292 gnd.n7364 gnd.n781 19.3944
R10293 gnd.n7364 gnd.n779 19.3944
R10294 gnd.n7368 gnd.n779 19.3944
R10295 gnd.n7368 gnd.n775 19.3944
R10296 gnd.n7374 gnd.n775 19.3944
R10297 gnd.n7374 gnd.n773 19.3944
R10298 gnd.n7378 gnd.n773 19.3944
R10299 gnd.n7378 gnd.n769 19.3944
R10300 gnd.n7384 gnd.n769 19.3944
R10301 gnd.n7384 gnd.n767 19.3944
R10302 gnd.n7388 gnd.n767 19.3944
R10303 gnd.n7388 gnd.n763 19.3944
R10304 gnd.n7394 gnd.n763 19.3944
R10305 gnd.n7394 gnd.n761 19.3944
R10306 gnd.n7398 gnd.n761 19.3944
R10307 gnd.n7398 gnd.n757 19.3944
R10308 gnd.n7404 gnd.n757 19.3944
R10309 gnd.n7404 gnd.n755 19.3944
R10310 gnd.n7408 gnd.n755 19.3944
R10311 gnd.n7408 gnd.n751 19.3944
R10312 gnd.n7414 gnd.n751 19.3944
R10313 gnd.n7414 gnd.n749 19.3944
R10314 gnd.n7418 gnd.n749 19.3944
R10315 gnd.n7418 gnd.n745 19.3944
R10316 gnd.n7424 gnd.n745 19.3944
R10317 gnd.n7424 gnd.n743 19.3944
R10318 gnd.n7428 gnd.n743 19.3944
R10319 gnd.n7428 gnd.n739 19.3944
R10320 gnd.n7434 gnd.n739 19.3944
R10321 gnd.n7434 gnd.n737 19.3944
R10322 gnd.n7438 gnd.n737 19.3944
R10323 gnd.n7438 gnd.n733 19.3944
R10324 gnd.n7444 gnd.n733 19.3944
R10325 gnd.n7444 gnd.n731 19.3944
R10326 gnd.n7448 gnd.n731 19.3944
R10327 gnd.n7448 gnd.n727 19.3944
R10328 gnd.n7454 gnd.n727 19.3944
R10329 gnd.n7454 gnd.n725 19.3944
R10330 gnd.n7458 gnd.n725 19.3944
R10331 gnd.n7458 gnd.n721 19.3944
R10332 gnd.n7464 gnd.n721 19.3944
R10333 gnd.n7464 gnd.n719 19.3944
R10334 gnd.n7468 gnd.n719 19.3944
R10335 gnd.n7468 gnd.n715 19.3944
R10336 gnd.n7474 gnd.n715 19.3944
R10337 gnd.n7474 gnd.n713 19.3944
R10338 gnd.n7478 gnd.n713 19.3944
R10339 gnd.n7478 gnd.n709 19.3944
R10340 gnd.n7484 gnd.n709 19.3944
R10341 gnd.n7484 gnd.n707 19.3944
R10342 gnd.n7488 gnd.n707 19.3944
R10343 gnd.n7488 gnd.n703 19.3944
R10344 gnd.n7494 gnd.n703 19.3944
R10345 gnd.n7494 gnd.n701 19.3944
R10346 gnd.n7499 gnd.n701 19.3944
R10347 gnd.n7499 gnd.n697 19.3944
R10348 gnd.n7505 gnd.n697 19.3944
R10349 gnd.n7506 gnd.n7505 19.3944
R10350 gnd.n4833 gnd.n4832 19.3944
R10351 gnd.n4832 gnd.n4831 19.3944
R10352 gnd.n4831 gnd.n4830 19.3944
R10353 gnd.n4830 gnd.n4828 19.3944
R10354 gnd.n4828 gnd.n4825 19.3944
R10355 gnd.n4825 gnd.n4824 19.3944
R10356 gnd.n4824 gnd.n4821 19.3944
R10357 gnd.n4821 gnd.n4820 19.3944
R10358 gnd.n4820 gnd.n4817 19.3944
R10359 gnd.n4817 gnd.n4816 19.3944
R10360 gnd.n4816 gnd.n4813 19.3944
R10361 gnd.n4813 gnd.n4812 19.3944
R10362 gnd.n4812 gnd.n4809 19.3944
R10363 gnd.n4809 gnd.n4808 19.3944
R10364 gnd.n4808 gnd.n4805 19.3944
R10365 gnd.n4805 gnd.n4804 19.3944
R10366 gnd.n4804 gnd.n4801 19.3944
R10367 gnd.n4799 gnd.n4796 19.3944
R10368 gnd.n4796 gnd.n4795 19.3944
R10369 gnd.n4795 gnd.n4792 19.3944
R10370 gnd.n4792 gnd.n4791 19.3944
R10371 gnd.n4791 gnd.n4788 19.3944
R10372 gnd.n4788 gnd.n4787 19.3944
R10373 gnd.n4787 gnd.n4784 19.3944
R10374 gnd.n4782 gnd.n4779 19.3944
R10375 gnd.n4779 gnd.n4778 19.3944
R10376 gnd.n4778 gnd.n4775 19.3944
R10377 gnd.n4775 gnd.n4774 19.3944
R10378 gnd.n4774 gnd.n4771 19.3944
R10379 gnd.n4771 gnd.n4770 19.3944
R10380 gnd.n4770 gnd.n4767 19.3944
R10381 gnd.n4767 gnd.n4766 19.3944
R10382 gnd.n4762 gnd.n4759 19.3944
R10383 gnd.n4759 gnd.n4758 19.3944
R10384 gnd.n4758 gnd.n4755 19.3944
R10385 gnd.n4755 gnd.n4754 19.3944
R10386 gnd.n4754 gnd.n4751 19.3944
R10387 gnd.n4751 gnd.n4750 19.3944
R10388 gnd.n4750 gnd.n4747 19.3944
R10389 gnd.n4747 gnd.n4746 19.3944
R10390 gnd.n4746 gnd.n4743 19.3944
R10391 gnd.n4743 gnd.n4742 19.3944
R10392 gnd.n4742 gnd.n4739 19.3944
R10393 gnd.n4739 gnd.n4738 19.3944
R10394 gnd.n4738 gnd.n4735 19.3944
R10395 gnd.n4735 gnd.n4734 19.3944
R10396 gnd.n4734 gnd.n4731 19.3944
R10397 gnd.n4731 gnd.n4730 19.3944
R10398 gnd.n4730 gnd.n4727 19.3944
R10399 gnd.n4727 gnd.n4726 19.3944
R10400 gnd.n4718 gnd.n1931 19.3944
R10401 gnd.n4575 gnd.n1931 19.3944
R10402 gnd.n4576 gnd.n4575 19.3944
R10403 gnd.n4577 gnd.n4576 19.3944
R10404 gnd.n4577 gnd.n2124 19.3944
R10405 gnd.n4589 gnd.n2124 19.3944
R10406 gnd.n4590 gnd.n4589 19.3944
R10407 gnd.n4591 gnd.n4590 19.3944
R10408 gnd.n4591 gnd.n2061 19.3944
R10409 gnd.n4603 gnd.n2061 19.3944
R10410 gnd.n4604 gnd.n4603 19.3944
R10411 gnd.n4605 gnd.n4604 19.3944
R10412 gnd.n4605 gnd.n2056 19.3944
R10413 gnd.n4617 gnd.n2056 19.3944
R10414 gnd.n4618 gnd.n4617 19.3944
R10415 gnd.n4622 gnd.n4618 19.3944
R10416 gnd.n4622 gnd.n4621 19.3944
R10417 gnd.n4621 gnd.n4620 19.3944
R10418 gnd.n4620 gnd.n2041 19.3944
R10419 gnd.n4654 gnd.n2041 19.3944
R10420 gnd.n4654 gnd.n2042 19.3944
R10421 gnd.n2042 gnd.n550 19.3944
R10422 gnd.n7746 gnd.n550 19.3944
R10423 gnd.n7747 gnd.n7746 19.3944
R10424 gnd.n7747 gnd.n523 19.3944
R10425 gnd.n7778 gnd.n523 19.3944
R10426 gnd.n7779 gnd.n7778 19.3944
R10427 gnd.n7780 gnd.n7779 19.3944
R10428 gnd.n7782 gnd.n7780 19.3944
R10429 gnd.n7782 gnd.n7781 19.3944
R10430 gnd.n7781 gnd.n493 19.3944
R10431 gnd.n7818 gnd.n493 19.3944
R10432 gnd.n7820 gnd.n7818 19.3944
R10433 gnd.n7820 gnd.n7819 19.3944
R10434 gnd.n7819 gnd.n486 19.3944
R10435 gnd.n7832 gnd.n486 19.3944
R10436 gnd.n7833 gnd.n7832 19.3944
R10437 gnd.n7835 gnd.n7833 19.3944
R10438 gnd.n7836 gnd.n7835 19.3944
R10439 gnd.n7839 gnd.n7836 19.3944
R10440 gnd.n7840 gnd.n7839 19.3944
R10441 gnd.n7842 gnd.n7840 19.3944
R10442 gnd.n7843 gnd.n7842 19.3944
R10443 gnd.n7846 gnd.n7843 19.3944
R10444 gnd.n7847 gnd.n7846 19.3944
R10445 gnd.n7849 gnd.n7847 19.3944
R10446 gnd.n7850 gnd.n7849 19.3944
R10447 gnd.n7853 gnd.n7850 19.3944
R10448 gnd.n7854 gnd.n7853 19.3944
R10449 gnd.n7856 gnd.n7854 19.3944
R10450 gnd.n7857 gnd.n7856 19.3944
R10451 gnd.n7860 gnd.n7857 19.3944
R10452 gnd.n7861 gnd.n7860 19.3944
R10453 gnd.n7863 gnd.n7861 19.3944
R10454 gnd.n7864 gnd.n7863 19.3944
R10455 gnd.n7867 gnd.n7864 19.3944
R10456 gnd.n7868 gnd.n7867 19.3944
R10457 gnd.n7870 gnd.n7868 19.3944
R10458 gnd.n7871 gnd.n7870 19.3944
R10459 gnd.n7874 gnd.n7871 19.3944
R10460 gnd.n7875 gnd.n7874 19.3944
R10461 gnd.n7877 gnd.n7875 19.3944
R10462 gnd.n7878 gnd.n7877 19.3944
R10463 gnd.n7881 gnd.n7878 19.3944
R10464 gnd.n1939 gnd.n1929 19.3944
R10465 gnd.n1955 gnd.n1939 19.3944
R10466 gnd.n4705 gnd.n1955 19.3944
R10467 gnd.n4705 gnd.n4704 19.3944
R10468 gnd.n4704 gnd.n4703 19.3944
R10469 gnd.n4703 gnd.n1959 19.3944
R10470 gnd.n4693 gnd.n1959 19.3944
R10471 gnd.n4693 gnd.n4692 19.3944
R10472 gnd.n4692 gnd.n4691 19.3944
R10473 gnd.n4691 gnd.n1980 19.3944
R10474 gnd.n4681 gnd.n1980 19.3944
R10475 gnd.n4681 gnd.n4680 19.3944
R10476 gnd.n4680 gnd.n4679 19.3944
R10477 gnd.n4679 gnd.n2000 19.3944
R10478 gnd.n4669 gnd.n2000 19.3944
R10479 gnd.n4669 gnd.n4668 19.3944
R10480 gnd.n4668 gnd.n4667 19.3944
R10481 gnd.n4667 gnd.n2021 19.3944
R10482 gnd.n4657 gnd.n2021 19.3944
R10483 gnd.n4657 gnd.n4656 19.3944
R10484 gnd.n4656 gnd.n547 19.3944
R10485 gnd.n7755 gnd.n547 19.3944
R10486 gnd.n7755 gnd.n7754 19.3944
R10487 gnd.n7754 gnd.n7753 19.3944
R10488 gnd.n7753 gnd.n7752 19.3944
R10489 gnd.n7752 gnd.n518 19.3944
R10490 gnd.n7788 gnd.n518 19.3944
R10491 gnd.n7788 gnd.n7787 19.3944
R10492 gnd.n7787 gnd.n7786 19.3944
R10493 gnd.n7786 gnd.n495 19.3944
R10494 gnd.n7815 gnd.n495 19.3944
R10495 gnd.n7815 gnd.n488 19.3944
R10496 gnd.n7824 gnd.n488 19.3944
R10497 gnd.n7825 gnd.n7824 19.3944
R10498 gnd.n7827 gnd.n7825 19.3944
R10499 gnd.n7827 gnd.n128 19.3944
R10500 gnd.n8087 gnd.n128 19.3944
R10501 gnd.n8087 gnd.n8086 19.3944
R10502 gnd.n8086 gnd.n8085 19.3944
R10503 gnd.n8085 gnd.n132 19.3944
R10504 gnd.n8075 gnd.n132 19.3944
R10505 gnd.n8075 gnd.n8074 19.3944
R10506 gnd.n8074 gnd.n8073 19.3944
R10507 gnd.n8073 gnd.n149 19.3944
R10508 gnd.n8063 gnd.n149 19.3944
R10509 gnd.n8063 gnd.n8062 19.3944
R10510 gnd.n8062 gnd.n8061 19.3944
R10511 gnd.n8061 gnd.n169 19.3944
R10512 gnd.n8051 gnd.n169 19.3944
R10513 gnd.n8051 gnd.n8050 19.3944
R10514 gnd.n8050 gnd.n8049 19.3944
R10515 gnd.n8049 gnd.n187 19.3944
R10516 gnd.n8039 gnd.n187 19.3944
R10517 gnd.n8039 gnd.n8038 19.3944
R10518 gnd.n8038 gnd.n8037 19.3944
R10519 gnd.n8037 gnd.n207 19.3944
R10520 gnd.n8027 gnd.n207 19.3944
R10521 gnd.n8027 gnd.n8026 19.3944
R10522 gnd.n8026 gnd.n8025 19.3944
R10523 gnd.n8025 gnd.n226 19.3944
R10524 gnd.n8015 gnd.n226 19.3944
R10525 gnd.n8015 gnd.n8014 19.3944
R10526 gnd.n8014 gnd.n8013 19.3944
R10527 gnd.n8013 gnd.n246 19.3944
R10528 gnd.n7924 gnd.n331 19.3944
R10529 gnd.n7924 gnd.n7921 19.3944
R10530 gnd.n7921 gnd.n7918 19.3944
R10531 gnd.n7918 gnd.n7917 19.3944
R10532 gnd.n7917 gnd.n7914 19.3944
R10533 gnd.n7914 gnd.n7913 19.3944
R10534 gnd.n7913 gnd.n7910 19.3944
R10535 gnd.n7910 gnd.n7909 19.3944
R10536 gnd.n7909 gnd.n7906 19.3944
R10537 gnd.n7906 gnd.n7905 19.3944
R10538 gnd.n7905 gnd.n7902 19.3944
R10539 gnd.n7902 gnd.n7901 19.3944
R10540 gnd.n7901 gnd.n7898 19.3944
R10541 gnd.n7898 gnd.n7897 19.3944
R10542 gnd.n7897 gnd.n7894 19.3944
R10543 gnd.n7894 gnd.n7893 19.3944
R10544 gnd.n7893 gnd.n7890 19.3944
R10545 gnd.n7890 gnd.n7889 19.3944
R10546 gnd.n7967 gnd.n7964 19.3944
R10547 gnd.n7964 gnd.n7963 19.3944
R10548 gnd.n7963 gnd.n7960 19.3944
R10549 gnd.n7960 gnd.n7959 19.3944
R10550 gnd.n7959 gnd.n7956 19.3944
R10551 gnd.n7956 gnd.n7955 19.3944
R10552 gnd.n7955 gnd.n7952 19.3944
R10553 gnd.n7952 gnd.n7951 19.3944
R10554 gnd.n7951 gnd.n7948 19.3944
R10555 gnd.n7948 gnd.n7947 19.3944
R10556 gnd.n7947 gnd.n7944 19.3944
R10557 gnd.n7944 gnd.n7943 19.3944
R10558 gnd.n7943 gnd.n7940 19.3944
R10559 gnd.n7940 gnd.n7939 19.3944
R10560 gnd.n7939 gnd.n7936 19.3944
R10561 gnd.n7936 gnd.n7935 19.3944
R10562 gnd.n7935 gnd.n7932 19.3944
R10563 gnd.n7932 gnd.n7931 19.3944
R10564 gnd.n8005 gnd.n255 19.3944
R10565 gnd.n8000 gnd.n255 19.3944
R10566 gnd.n8000 gnd.n7999 19.3944
R10567 gnd.n7999 gnd.n7998 19.3944
R10568 gnd.n7998 gnd.n7995 19.3944
R10569 gnd.n7995 gnd.n7994 19.3944
R10570 gnd.n7994 gnd.n7991 19.3944
R10571 gnd.n7991 gnd.n7990 19.3944
R10572 gnd.n7990 gnd.n7987 19.3944
R10573 gnd.n7987 gnd.n7986 19.3944
R10574 gnd.n7986 gnd.n7983 19.3944
R10575 gnd.n7983 gnd.n7982 19.3944
R10576 gnd.n7982 gnd.n7979 19.3944
R10577 gnd.n7979 gnd.n7978 19.3944
R10578 gnd.n7978 gnd.n7975 19.3944
R10579 gnd.n7975 gnd.n7974 19.3944
R10580 gnd.n7974 gnd.n7971 19.3944
R10581 gnd.n484 gnd.n483 19.3944
R10582 gnd.n483 gnd.n482 19.3944
R10583 gnd.n482 gnd.n479 19.3944
R10584 gnd.n479 gnd.n478 19.3944
R10585 gnd.n478 gnd.n475 19.3944
R10586 gnd.n475 gnd.n474 19.3944
R10587 gnd.n474 gnd.n471 19.3944
R10588 gnd.n471 gnd.n470 19.3944
R10589 gnd.n470 gnd.n467 19.3944
R10590 gnd.n467 gnd.n466 19.3944
R10591 gnd.n466 gnd.n463 19.3944
R10592 gnd.n463 gnd.n462 19.3944
R10593 gnd.n462 gnd.n459 19.3944
R10594 gnd.n459 gnd.n458 19.3944
R10595 gnd.n458 gnd.n455 19.3944
R10596 gnd.n455 gnd.n454 19.3944
R10597 gnd.n4567 gnd.n2130 19.3944
R10598 gnd.n4571 gnd.n2130 19.3944
R10599 gnd.n4571 gnd.n2128 19.3944
R10600 gnd.n4581 gnd.n2128 19.3944
R10601 gnd.n4581 gnd.n2126 19.3944
R10602 gnd.n4585 gnd.n2126 19.3944
R10603 gnd.n4585 gnd.n2123 19.3944
R10604 gnd.n4595 gnd.n2123 19.3944
R10605 gnd.n4595 gnd.n2121 19.3944
R10606 gnd.n4599 gnd.n2121 19.3944
R10607 gnd.n4599 gnd.n2060 19.3944
R10608 gnd.n4609 gnd.n2060 19.3944
R10609 gnd.n4609 gnd.n2058 19.3944
R10610 gnd.n4613 gnd.n2058 19.3944
R10611 gnd.n4613 gnd.n2055 19.3944
R10612 gnd.n4626 gnd.n2055 19.3944
R10613 gnd.n4626 gnd.n2052 19.3944
R10614 gnd.n4638 gnd.n2052 19.3944
R10615 gnd.n4638 gnd.n2053 19.3944
R10616 gnd.n4634 gnd.n2053 19.3944
R10617 gnd.n4634 gnd.n4633 19.3944
R10618 gnd.n4633 gnd.n4632 19.3944
R10619 gnd.n4632 gnd.n530 19.3944
R10620 gnd.n7770 gnd.n530 19.3944
R10621 gnd.n7770 gnd.n528 19.3944
R10622 gnd.n7774 gnd.n528 19.3944
R10623 gnd.n7774 gnd.n508 19.3944
R10624 gnd.n7797 gnd.n508 19.3944
R10625 gnd.n7797 gnd.n505 19.3944
R10626 gnd.n7801 gnd.n505 19.3944
R10627 gnd.n7801 gnd.n506 19.3944
R10628 gnd.n506 gnd.n100 19.3944
R10629 gnd.n8100 gnd.n100 19.3944
R10630 gnd.n8100 gnd.n8099 19.3944
R10631 gnd.n8099 gnd.n103 19.3944
R10632 gnd.n390 gnd.n103 19.3944
R10633 gnd.n390 gnd.n387 19.3944
R10634 gnd.n395 gnd.n387 19.3944
R10635 gnd.n396 gnd.n395 19.3944
R10636 gnd.n398 gnd.n396 19.3944
R10637 gnd.n398 gnd.n385 19.3944
R10638 gnd.n403 gnd.n385 19.3944
R10639 gnd.n404 gnd.n403 19.3944
R10640 gnd.n406 gnd.n404 19.3944
R10641 gnd.n406 gnd.n383 19.3944
R10642 gnd.n411 gnd.n383 19.3944
R10643 gnd.n412 gnd.n411 19.3944
R10644 gnd.n414 gnd.n412 19.3944
R10645 gnd.n414 gnd.n381 19.3944
R10646 gnd.n419 gnd.n381 19.3944
R10647 gnd.n420 gnd.n419 19.3944
R10648 gnd.n422 gnd.n420 19.3944
R10649 gnd.n422 gnd.n379 19.3944
R10650 gnd.n427 gnd.n379 19.3944
R10651 gnd.n428 gnd.n427 19.3944
R10652 gnd.n430 gnd.n428 19.3944
R10653 gnd.n430 gnd.n377 19.3944
R10654 gnd.n435 gnd.n377 19.3944
R10655 gnd.n436 gnd.n435 19.3944
R10656 gnd.n438 gnd.n436 19.3944
R10657 gnd.n438 gnd.n375 19.3944
R10658 gnd.n443 gnd.n375 19.3944
R10659 gnd.n444 gnd.n443 19.3944
R10660 gnd.n447 gnd.n444 19.3944
R10661 gnd.n4711 gnd.n1943 19.3944
R10662 gnd.n4711 gnd.n4710 19.3944
R10663 gnd.n4710 gnd.n4709 19.3944
R10664 gnd.n4709 gnd.n1948 19.3944
R10665 gnd.n4699 gnd.n1948 19.3944
R10666 gnd.n4699 gnd.n4698 19.3944
R10667 gnd.n4698 gnd.n4697 19.3944
R10668 gnd.n4697 gnd.n1970 19.3944
R10669 gnd.n4687 gnd.n1970 19.3944
R10670 gnd.n4687 gnd.n4686 19.3944
R10671 gnd.n4686 gnd.n4685 19.3944
R10672 gnd.n4685 gnd.n1990 19.3944
R10673 gnd.n4675 gnd.n1990 19.3944
R10674 gnd.n4675 gnd.n4674 19.3944
R10675 gnd.n4674 gnd.n4673 19.3944
R10676 gnd.n4673 gnd.n2011 19.3944
R10677 gnd.n4663 gnd.n2011 19.3944
R10678 gnd.n4663 gnd.n4662 19.3944
R10679 gnd.n4662 gnd.n4661 19.3944
R10680 gnd.n4661 gnd.n2032 19.3944
R10681 gnd.n2032 gnd.n540 19.3944
R10682 gnd.n7759 gnd.n540 19.3944
R10683 gnd.n7759 gnd.n538 19.3944
R10684 gnd.n7766 gnd.n538 19.3944
R10685 gnd.n7766 gnd.n7765 19.3944
R10686 gnd.n7765 gnd.n7764 19.3944
R10687 gnd.n7764 gnd.n514 19.3944
R10688 gnd.n7793 gnd.n7792 19.3944
R10689 gnd.n7811 gnd.n7810 19.3944
R10690 gnd.n7806 gnd.n7805 19.3944
R10691 gnd.n8095 gnd.n8094 19.3944
R10692 gnd.n8091 gnd.n112 19.3944
R10693 gnd.n8091 gnd.n119 19.3944
R10694 gnd.n8081 gnd.n119 19.3944
R10695 gnd.n8081 gnd.n8080 19.3944
R10696 gnd.n8080 gnd.n8079 19.3944
R10697 gnd.n8079 gnd.n141 19.3944
R10698 gnd.n8069 gnd.n141 19.3944
R10699 gnd.n8069 gnd.n8068 19.3944
R10700 gnd.n8068 gnd.n8067 19.3944
R10701 gnd.n8067 gnd.n159 19.3944
R10702 gnd.n8057 gnd.n159 19.3944
R10703 gnd.n8057 gnd.n8056 19.3944
R10704 gnd.n8056 gnd.n8055 19.3944
R10705 gnd.n8055 gnd.n179 19.3944
R10706 gnd.n8045 gnd.n179 19.3944
R10707 gnd.n8045 gnd.n8044 19.3944
R10708 gnd.n8044 gnd.n8043 19.3944
R10709 gnd.n8043 gnd.n197 19.3944
R10710 gnd.n8033 gnd.n197 19.3944
R10711 gnd.n8033 gnd.n8032 19.3944
R10712 gnd.n8032 gnd.n8031 19.3944
R10713 gnd.n8031 gnd.n217 19.3944
R10714 gnd.n8021 gnd.n217 19.3944
R10715 gnd.n8021 gnd.n8020 19.3944
R10716 gnd.n8020 gnd.n8019 19.3944
R10717 gnd.n8019 gnd.n237 19.3944
R10718 gnd.n8009 gnd.n237 19.3944
R10719 gnd.n8009 gnd.n8008 19.3944
R10720 gnd.n5397 gnd.n5396 19.3944
R10721 gnd.n5396 gnd.n5395 19.3944
R10722 gnd.n5395 gnd.n5394 19.3944
R10723 gnd.n5394 gnd.n5392 19.3944
R10724 gnd.n5392 gnd.n5389 19.3944
R10725 gnd.n5389 gnd.n5388 19.3944
R10726 gnd.n5388 gnd.n5385 19.3944
R10727 gnd.n5385 gnd.n5384 19.3944
R10728 gnd.n5384 gnd.n5381 19.3944
R10729 gnd.n5381 gnd.n5380 19.3944
R10730 gnd.n5380 gnd.n5377 19.3944
R10731 gnd.n5377 gnd.n5376 19.3944
R10732 gnd.n5376 gnd.n5373 19.3944
R10733 gnd.n5373 gnd.n5372 19.3944
R10734 gnd.n5372 gnd.n5369 19.3944
R10735 gnd.n5369 gnd.n5368 19.3944
R10736 gnd.n5368 gnd.n5365 19.3944
R10737 gnd.n5363 gnd.n5360 19.3944
R10738 gnd.n5360 gnd.n5359 19.3944
R10739 gnd.n5359 gnd.n5356 19.3944
R10740 gnd.n5356 gnd.n5355 19.3944
R10741 gnd.n5355 gnd.n5352 19.3944
R10742 gnd.n5352 gnd.n5351 19.3944
R10743 gnd.n5351 gnd.n5348 19.3944
R10744 gnd.n5348 gnd.n5347 19.3944
R10745 gnd.n5347 gnd.n5344 19.3944
R10746 gnd.n5344 gnd.n5343 19.3944
R10747 gnd.n5343 gnd.n5340 19.3944
R10748 gnd.n5340 gnd.n5339 19.3944
R10749 gnd.n5339 gnd.n5336 19.3944
R10750 gnd.n5336 gnd.n5335 19.3944
R10751 gnd.n5335 gnd.n5332 19.3944
R10752 gnd.n5332 gnd.n5331 19.3944
R10753 gnd.n5331 gnd.n5328 19.3944
R10754 gnd.n5328 gnd.n5327 19.3944
R10755 gnd.n5323 gnd.n5320 19.3944
R10756 gnd.n5320 gnd.n5319 19.3944
R10757 gnd.n5319 gnd.n5316 19.3944
R10758 gnd.n5316 gnd.n5315 19.3944
R10759 gnd.n5315 gnd.n5312 19.3944
R10760 gnd.n5312 gnd.n5311 19.3944
R10761 gnd.n5311 gnd.n5308 19.3944
R10762 gnd.n5308 gnd.n5307 19.3944
R10763 gnd.n5307 gnd.n5304 19.3944
R10764 gnd.n5304 gnd.n5303 19.3944
R10765 gnd.n5303 gnd.n5300 19.3944
R10766 gnd.n5300 gnd.n5299 19.3944
R10767 gnd.n5299 gnd.n5296 19.3944
R10768 gnd.n5296 gnd.n5295 19.3944
R10769 gnd.n5295 gnd.n5292 19.3944
R10770 gnd.n5292 gnd.n5291 19.3944
R10771 gnd.n5291 gnd.n5288 19.3944
R10772 gnd.n5288 gnd.n5287 19.3944
R10773 gnd.n2916 gnd.n2915 19.3944
R10774 gnd.n2919 gnd.n2916 19.3944
R10775 gnd.n2919 gnd.n2911 19.3944
R10776 gnd.n2925 gnd.n2911 19.3944
R10777 gnd.n2926 gnd.n2925 19.3944
R10778 gnd.n2929 gnd.n2926 19.3944
R10779 gnd.n2929 gnd.n2909 19.3944
R10780 gnd.n2935 gnd.n2909 19.3944
R10781 gnd.n2936 gnd.n2935 19.3944
R10782 gnd.n2939 gnd.n2936 19.3944
R10783 gnd.n2939 gnd.n2907 19.3944
R10784 gnd.n2945 gnd.n2907 19.3944
R10785 gnd.n2946 gnd.n2945 19.3944
R10786 gnd.n2949 gnd.n2946 19.3944
R10787 gnd.n2949 gnd.n2903 19.3944
R10788 gnd.n2953 gnd.n2903 19.3944
R10789 gnd.n2960 gnd.n2959 19.3944
R10790 gnd.n2962 gnd.n2960 19.3944
R10791 gnd.n2962 gnd.n2897 19.3944
R10792 gnd.n2967 gnd.n2897 19.3944
R10793 gnd.n2968 gnd.n2967 19.3944
R10794 gnd.n2970 gnd.n2968 19.3944
R10795 gnd.n2970 gnd.n2895 19.3944
R10796 gnd.n2975 gnd.n2895 19.3944
R10797 gnd.n2976 gnd.n2975 19.3944
R10798 gnd.n2978 gnd.n2976 19.3944
R10799 gnd.n2978 gnd.n2893 19.3944
R10800 gnd.n2983 gnd.n2893 19.3944
R10801 gnd.n2984 gnd.n2983 19.3944
R10802 gnd.n2986 gnd.n2984 19.3944
R10803 gnd.n2986 gnd.n2891 19.3944
R10804 gnd.n2991 gnd.n2891 19.3944
R10805 gnd.n2992 gnd.n2991 19.3944
R10806 gnd.n2994 gnd.n2992 19.3944
R10807 gnd.n2994 gnd.n2889 19.3944
R10808 gnd.n2999 gnd.n2889 19.3944
R10809 gnd.n3000 gnd.n2999 19.3944
R10810 gnd.n3002 gnd.n3000 19.3944
R10811 gnd.n3002 gnd.n2887 19.3944
R10812 gnd.n3007 gnd.n2887 19.3944
R10813 gnd.n3008 gnd.n3007 19.3944
R10814 gnd.n3010 gnd.n3008 19.3944
R10815 gnd.n3010 gnd.n2885 19.3944
R10816 gnd.n3015 gnd.n2885 19.3944
R10817 gnd.n3016 gnd.n3015 19.3944
R10818 gnd.n3018 gnd.n3016 19.3944
R10819 gnd.n3018 gnd.n2883 19.3944
R10820 gnd.n3022 gnd.n2883 19.3944
R10821 gnd.n3022 gnd.n2789 19.3944
R10822 gnd.n3048 gnd.n2789 19.3944
R10823 gnd.n3048 gnd.n2787 19.3944
R10824 gnd.n3052 gnd.n2787 19.3944
R10825 gnd.n3052 gnd.n2776 19.3944
R10826 gnd.n3087 gnd.n2776 19.3944
R10827 gnd.n3087 gnd.n2774 19.3944
R10828 gnd.n3091 gnd.n2774 19.3944
R10829 gnd.n3091 gnd.n2771 19.3944
R10830 gnd.n3101 gnd.n2771 19.3944
R10831 gnd.n3101 gnd.n2769 19.3944
R10832 gnd.n3105 gnd.n2769 19.3944
R10833 gnd.n3105 gnd.n2759 19.3944
R10834 gnd.n3140 gnd.n2759 19.3944
R10835 gnd.n3140 gnd.n2760 19.3944
R10836 gnd.n3136 gnd.n2760 19.3944
R10837 gnd.n3136 gnd.n3135 19.3944
R10838 gnd.n3135 gnd.n3134 19.3944
R10839 gnd.n3134 gnd.n2765 19.3944
R10840 gnd.n3130 gnd.n2765 19.3944
R10841 gnd.n3130 gnd.n3129 19.3944
R10842 gnd.n3129 gnd.n3128 19.3944
R10843 gnd.n3128 gnd.n2744 19.3944
R10844 gnd.n3195 gnd.n2744 19.3944
R10845 gnd.n3195 gnd.n2742 19.3944
R10846 gnd.n3199 gnd.n2742 19.3944
R10847 gnd.n3199 gnd.n2740 19.3944
R10848 gnd.n3210 gnd.n2740 19.3944
R10849 gnd.n3210 gnd.n2737 19.3944
R10850 gnd.n3216 gnd.n2737 19.3944
R10851 gnd.n3216 gnd.n2738 19.3944
R10852 gnd.n2738 gnd.n2553 19.3944
R10853 gnd.n5279 gnd.n1257 19.3944
R10854 gnd.n2826 gnd.n1257 19.3944
R10855 gnd.n2827 gnd.n2826 19.3944
R10856 gnd.n2829 gnd.n2827 19.3944
R10857 gnd.n2830 gnd.n2829 19.3944
R10858 gnd.n2833 gnd.n2830 19.3944
R10859 gnd.n2834 gnd.n2833 19.3944
R10860 gnd.n2836 gnd.n2834 19.3944
R10861 gnd.n2837 gnd.n2836 19.3944
R10862 gnd.n2840 gnd.n2837 19.3944
R10863 gnd.n2841 gnd.n2840 19.3944
R10864 gnd.n2843 gnd.n2841 19.3944
R10865 gnd.n2844 gnd.n2843 19.3944
R10866 gnd.n2847 gnd.n2844 19.3944
R10867 gnd.n2848 gnd.n2847 19.3944
R10868 gnd.n2850 gnd.n2848 19.3944
R10869 gnd.n2851 gnd.n2850 19.3944
R10870 gnd.n2854 gnd.n2851 19.3944
R10871 gnd.n2855 gnd.n2854 19.3944
R10872 gnd.n2857 gnd.n2855 19.3944
R10873 gnd.n2858 gnd.n2857 19.3944
R10874 gnd.n2861 gnd.n2858 19.3944
R10875 gnd.n2862 gnd.n2861 19.3944
R10876 gnd.n2864 gnd.n2862 19.3944
R10877 gnd.n2865 gnd.n2864 19.3944
R10878 gnd.n2868 gnd.n2865 19.3944
R10879 gnd.n2869 gnd.n2868 19.3944
R10880 gnd.n2871 gnd.n2869 19.3944
R10881 gnd.n2872 gnd.n2871 19.3944
R10882 gnd.n2874 gnd.n2872 19.3944
R10883 gnd.n2874 gnd.n2805 19.3944
R10884 gnd.n3026 gnd.n2805 19.3944
R10885 gnd.n3027 gnd.n3026 19.3944
R10886 gnd.n3028 gnd.n3027 19.3944
R10887 gnd.n3033 gnd.n3028 19.3944
R10888 gnd.n3033 gnd.n3031 19.3944
R10889 gnd.n3031 gnd.n3030 19.3944
R10890 gnd.n3030 gnd.n3029 19.3944
R10891 gnd.n3029 gnd.n2772 19.3944
R10892 gnd.n3095 gnd.n2772 19.3944
R10893 gnd.n3096 gnd.n3095 19.3944
R10894 gnd.n3097 gnd.n3096 19.3944
R10895 gnd.n3097 gnd.n2767 19.3944
R10896 gnd.n3109 gnd.n2767 19.3944
R10897 gnd.n3110 gnd.n3109 19.3944
R10898 gnd.n3111 gnd.n3110 19.3944
R10899 gnd.n3112 gnd.n3111 19.3944
R10900 gnd.n3116 gnd.n3112 19.3944
R10901 gnd.n3117 gnd.n3116 19.3944
R10902 gnd.n3120 gnd.n3117 19.3944
R10903 gnd.n3121 gnd.n3120 19.3944
R10904 gnd.n3123 gnd.n3121 19.3944
R10905 gnd.n3123 gnd.n2745 19.3944
R10906 gnd.n3188 gnd.n2745 19.3944
R10907 gnd.n3189 gnd.n3188 19.3944
R10908 gnd.n3191 gnd.n3189 19.3944
R10909 gnd.n3191 gnd.n2741 19.3944
R10910 gnd.n3203 gnd.n2741 19.3944
R10911 gnd.n3204 gnd.n3203 19.3944
R10912 gnd.n3206 gnd.n3204 19.3944
R10913 gnd.n3206 gnd.n2736 19.3944
R10914 gnd.n3220 gnd.n2736 19.3944
R10915 gnd.n3221 gnd.n3220 19.3944
R10916 gnd.n3222 gnd.n3221 19.3944
R10917 gnd.n1276 gnd.n1255 19.3944
R10918 gnd.n1277 gnd.n1276 19.3944
R10919 gnd.n5268 gnd.n1277 19.3944
R10920 gnd.n5268 gnd.n5267 19.3944
R10921 gnd.n5267 gnd.n5266 19.3944
R10922 gnd.n5266 gnd.n1281 19.3944
R10923 gnd.n5256 gnd.n1281 19.3944
R10924 gnd.n5256 gnd.n5255 19.3944
R10925 gnd.n5255 gnd.n5254 19.3944
R10926 gnd.n5254 gnd.n1300 19.3944
R10927 gnd.n5244 gnd.n1300 19.3944
R10928 gnd.n5244 gnd.n5243 19.3944
R10929 gnd.n5243 gnd.n5242 19.3944
R10930 gnd.n5242 gnd.n1319 19.3944
R10931 gnd.n5232 gnd.n1319 19.3944
R10932 gnd.n5232 gnd.n5231 19.3944
R10933 gnd.n5231 gnd.n5230 19.3944
R10934 gnd.n5230 gnd.n1338 19.3944
R10935 gnd.n5220 gnd.n1338 19.3944
R10936 gnd.n5220 gnd.n5219 19.3944
R10937 gnd.n5219 gnd.n5218 19.3944
R10938 gnd.n5218 gnd.n1357 19.3944
R10939 gnd.n5208 gnd.n1357 19.3944
R10940 gnd.n5208 gnd.n5207 19.3944
R10941 gnd.n5207 gnd.n5206 19.3944
R10942 gnd.n5206 gnd.n1376 19.3944
R10943 gnd.n5196 gnd.n1376 19.3944
R10944 gnd.n5196 gnd.n5195 19.3944
R10945 gnd.n5195 gnd.n5194 19.3944
R10946 gnd.n5194 gnd.n1394 19.3944
R10947 gnd.n2877 gnd.n1394 19.3944
R10948 gnd.n2877 gnd.n2801 19.3944
R10949 gnd.n3038 gnd.n2801 19.3944
R10950 gnd.n3038 gnd.n3037 19.3944
R10951 gnd.n3037 gnd.n3036 19.3944
R10952 gnd.n3036 gnd.n1418 19.3944
R10953 gnd.n5183 gnd.n1418 19.3944
R10954 gnd.n5183 gnd.n5182 19.3944
R10955 gnd.n5182 gnd.n5181 19.3944
R10956 gnd.n5181 gnd.n1422 19.3944
R10957 gnd.n5171 gnd.n1422 19.3944
R10958 gnd.n5171 gnd.n5170 19.3944
R10959 gnd.n5170 gnd.n5169 19.3944
R10960 gnd.n5169 gnd.n1441 19.3944
R10961 gnd.n5159 gnd.n1441 19.3944
R10962 gnd.n5159 gnd.n5158 19.3944
R10963 gnd.n5158 gnd.n5157 19.3944
R10964 gnd.n5157 gnd.n1462 19.3944
R10965 gnd.n5147 gnd.n1462 19.3944
R10966 gnd.n5147 gnd.n5146 19.3944
R10967 gnd.n5146 gnd.n5145 19.3944
R10968 gnd.n5145 gnd.n1482 19.3944
R10969 gnd.n5135 gnd.n1482 19.3944
R10970 gnd.n5135 gnd.n5134 19.3944
R10971 gnd.n5134 gnd.n5133 19.3944
R10972 gnd.n5133 gnd.n1503 19.3944
R10973 gnd.n5123 gnd.n1503 19.3944
R10974 gnd.n5123 gnd.n5122 19.3944
R10975 gnd.n5122 gnd.n5121 19.3944
R10976 gnd.n5121 gnd.n1523 19.3944
R10977 gnd.n5111 gnd.n1523 19.3944
R10978 gnd.n5111 gnd.n5110 19.3944
R10979 gnd.n5110 gnd.n5109 19.3944
R10980 gnd.n5109 gnd.n1544 19.3944
R10981 gnd.n5101 gnd.n1554 19.3944
R10982 gnd.n5096 gnd.n1554 19.3944
R10983 gnd.n5096 gnd.n5095 19.3944
R10984 gnd.n5095 gnd.n5094 19.3944
R10985 gnd.n5094 gnd.n5091 19.3944
R10986 gnd.n5091 gnd.n5090 19.3944
R10987 gnd.n5090 gnd.n5087 19.3944
R10988 gnd.n5087 gnd.n5086 19.3944
R10989 gnd.n5086 gnd.n5083 19.3944
R10990 gnd.n5083 gnd.n5082 19.3944
R10991 gnd.n5082 gnd.n5079 19.3944
R10992 gnd.n5079 gnd.n5078 19.3944
R10993 gnd.n5078 gnd.n5075 19.3944
R10994 gnd.n5075 gnd.n5074 19.3944
R10995 gnd.n5074 gnd.n5071 19.3944
R10996 gnd.n5071 gnd.n5070 19.3944
R10997 gnd.n5070 gnd.n5067 19.3944
R10998 gnd.n2686 gnd.n2652 19.3944
R10999 gnd.n2690 gnd.n2652 19.3944
R11000 gnd.n2693 gnd.n2690 19.3944
R11001 gnd.n2696 gnd.n2693 19.3944
R11002 gnd.n2696 gnd.n2650 19.3944
R11003 gnd.n2700 gnd.n2650 19.3944
R11004 gnd.n2703 gnd.n2700 19.3944
R11005 gnd.n2706 gnd.n2703 19.3944
R11006 gnd.n2706 gnd.n2648 19.3944
R11007 gnd.n2710 gnd.n2648 19.3944
R11008 gnd.n2713 gnd.n2710 19.3944
R11009 gnd.n2716 gnd.n2713 19.3944
R11010 gnd.n2716 gnd.n2646 19.3944
R11011 gnd.n2720 gnd.n2646 19.3944
R11012 gnd.n2723 gnd.n2720 19.3944
R11013 gnd.n2726 gnd.n2723 19.3944
R11014 gnd.n2726 gnd.n2644 19.3944
R11015 gnd.n2731 gnd.n2644 19.3944
R11016 gnd.n2664 gnd.n1623 19.3944
R11017 gnd.n2667 gnd.n2664 19.3944
R11018 gnd.n2667 gnd.n2659 19.3944
R11019 gnd.n2671 gnd.n2659 19.3944
R11020 gnd.n2674 gnd.n2671 19.3944
R11021 gnd.n2677 gnd.n2674 19.3944
R11022 gnd.n2677 gnd.n2657 19.3944
R11023 gnd.n2682 gnd.n2657 19.3944
R11024 gnd.n5065 gnd.n5062 19.3944
R11025 gnd.n5062 gnd.n5061 19.3944
R11026 gnd.n5061 gnd.n5058 19.3944
R11027 gnd.n5058 gnd.n5057 19.3944
R11028 gnd.n5057 gnd.n5054 19.3944
R11029 gnd.n5054 gnd.n5053 19.3944
R11030 gnd.n5053 gnd.n5050 19.3944
R11031 gnd.n5274 gnd.n1263 19.3944
R11032 gnd.n5274 gnd.n5273 19.3944
R11033 gnd.n5273 gnd.n5272 19.3944
R11034 gnd.n5272 gnd.n1268 19.3944
R11035 gnd.n5262 gnd.n1268 19.3944
R11036 gnd.n5262 gnd.n5261 19.3944
R11037 gnd.n5261 gnd.n5260 19.3944
R11038 gnd.n5260 gnd.n1291 19.3944
R11039 gnd.n5250 gnd.n1291 19.3944
R11040 gnd.n5250 gnd.n5249 19.3944
R11041 gnd.n5249 gnd.n5248 19.3944
R11042 gnd.n5248 gnd.n1309 19.3944
R11043 gnd.n5238 gnd.n1309 19.3944
R11044 gnd.n5238 gnd.n5237 19.3944
R11045 gnd.n5237 gnd.n5236 19.3944
R11046 gnd.n5236 gnd.n1329 19.3944
R11047 gnd.n5226 gnd.n1329 19.3944
R11048 gnd.n5226 gnd.n5225 19.3944
R11049 gnd.n5225 gnd.n5224 19.3944
R11050 gnd.n5224 gnd.n1347 19.3944
R11051 gnd.n5214 gnd.n1347 19.3944
R11052 gnd.n5214 gnd.n5213 19.3944
R11053 gnd.n5213 gnd.n5212 19.3944
R11054 gnd.n5212 gnd.n1367 19.3944
R11055 gnd.n5202 gnd.n1367 19.3944
R11056 gnd.n5202 gnd.n5201 19.3944
R11057 gnd.n5201 gnd.n5200 19.3944
R11058 gnd.n5190 gnd.n1401 19.3944
R11059 gnd.n2879 gnd.n1402 19.3944
R11060 gnd.n2796 gnd.n2795 19.3944
R11061 gnd.n3044 gnd.n3043 19.3944
R11062 gnd.n5187 gnd.n1408 19.3944
R11063 gnd.n5187 gnd.n1409 19.3944
R11064 gnd.n5177 gnd.n1409 19.3944
R11065 gnd.n5177 gnd.n5176 19.3944
R11066 gnd.n5176 gnd.n5175 19.3944
R11067 gnd.n5175 gnd.n1431 19.3944
R11068 gnd.n5165 gnd.n1431 19.3944
R11069 gnd.n5165 gnd.n5164 19.3944
R11070 gnd.n5164 gnd.n5163 19.3944
R11071 gnd.n5163 gnd.n1452 19.3944
R11072 gnd.n5153 gnd.n1452 19.3944
R11073 gnd.n5153 gnd.n5152 19.3944
R11074 gnd.n5152 gnd.n5151 19.3944
R11075 gnd.n5151 gnd.n1472 19.3944
R11076 gnd.n5141 gnd.n1472 19.3944
R11077 gnd.n5141 gnd.n5140 19.3944
R11078 gnd.n5140 gnd.n5139 19.3944
R11079 gnd.n5139 gnd.n1493 19.3944
R11080 gnd.n5129 gnd.n1493 19.3944
R11081 gnd.n5129 gnd.n5128 19.3944
R11082 gnd.n5128 gnd.n5127 19.3944
R11083 gnd.n5127 gnd.n1513 19.3944
R11084 gnd.n5117 gnd.n1513 19.3944
R11085 gnd.n5117 gnd.n5116 19.3944
R11086 gnd.n5116 gnd.n5115 19.3944
R11087 gnd.n5115 gnd.n1534 19.3944
R11088 gnd.n5105 gnd.n1534 19.3944
R11089 gnd.n5105 gnd.n5104 19.3944
R11090 gnd.n7048 gnd.n970 19.3944
R11091 gnd.n7048 gnd.n7047 19.3944
R11092 gnd.n7047 gnd.n7046 19.3944
R11093 gnd.n7046 gnd.n974 19.3944
R11094 gnd.n7040 gnd.n974 19.3944
R11095 gnd.n7040 gnd.n7039 19.3944
R11096 gnd.n7039 gnd.n7038 19.3944
R11097 gnd.n7038 gnd.n982 19.3944
R11098 gnd.n7032 gnd.n982 19.3944
R11099 gnd.n7032 gnd.n7031 19.3944
R11100 gnd.n7031 gnd.n7030 19.3944
R11101 gnd.n7030 gnd.n990 19.3944
R11102 gnd.n7024 gnd.n990 19.3944
R11103 gnd.n7024 gnd.n7023 19.3944
R11104 gnd.n7023 gnd.n7022 19.3944
R11105 gnd.n7022 gnd.n998 19.3944
R11106 gnd.n7016 gnd.n998 19.3944
R11107 gnd.n7016 gnd.n7015 19.3944
R11108 gnd.n7015 gnd.n7014 19.3944
R11109 gnd.n7014 gnd.n1006 19.3944
R11110 gnd.n7008 gnd.n1006 19.3944
R11111 gnd.n7008 gnd.n7007 19.3944
R11112 gnd.n7007 gnd.n7006 19.3944
R11113 gnd.n7006 gnd.n1014 19.3944
R11114 gnd.n7000 gnd.n1014 19.3944
R11115 gnd.n7000 gnd.n6999 19.3944
R11116 gnd.n6999 gnd.n6998 19.3944
R11117 gnd.n6998 gnd.n1022 19.3944
R11118 gnd.n6992 gnd.n1022 19.3944
R11119 gnd.n6992 gnd.n6991 19.3944
R11120 gnd.n6991 gnd.n6990 19.3944
R11121 gnd.n6990 gnd.n1030 19.3944
R11122 gnd.n6984 gnd.n1030 19.3944
R11123 gnd.n6984 gnd.n6983 19.3944
R11124 gnd.n6983 gnd.n6982 19.3944
R11125 gnd.n6982 gnd.n1038 19.3944
R11126 gnd.n6976 gnd.n1038 19.3944
R11127 gnd.n6976 gnd.n6975 19.3944
R11128 gnd.n6975 gnd.n6974 19.3944
R11129 gnd.n6974 gnd.n1046 19.3944
R11130 gnd.n6968 gnd.n1046 19.3944
R11131 gnd.n6968 gnd.n6967 19.3944
R11132 gnd.n6967 gnd.n6966 19.3944
R11133 gnd.n6966 gnd.n1054 19.3944
R11134 gnd.n6960 gnd.n1054 19.3944
R11135 gnd.n6960 gnd.n6959 19.3944
R11136 gnd.n6959 gnd.n6958 19.3944
R11137 gnd.n6958 gnd.n1062 19.3944
R11138 gnd.n6952 gnd.n1062 19.3944
R11139 gnd.n6952 gnd.n6951 19.3944
R11140 gnd.n6951 gnd.n6950 19.3944
R11141 gnd.n6950 gnd.n1070 19.3944
R11142 gnd.n6944 gnd.n1070 19.3944
R11143 gnd.n6944 gnd.n6943 19.3944
R11144 gnd.n6943 gnd.n6942 19.3944
R11145 gnd.n6942 gnd.n1078 19.3944
R11146 gnd.n6936 gnd.n1078 19.3944
R11147 gnd.n6936 gnd.n6935 19.3944
R11148 gnd.n6935 gnd.n6934 19.3944
R11149 gnd.n6934 gnd.n1086 19.3944
R11150 gnd.n6928 gnd.n1086 19.3944
R11151 gnd.n6928 gnd.n6927 19.3944
R11152 gnd.n6927 gnd.n6926 19.3944
R11153 gnd.n6926 gnd.n1094 19.3944
R11154 gnd.n6920 gnd.n1094 19.3944
R11155 gnd.n6920 gnd.n6919 19.3944
R11156 gnd.n6919 gnd.n6918 19.3944
R11157 gnd.n6918 gnd.n1102 19.3944
R11158 gnd.n6912 gnd.n1102 19.3944
R11159 gnd.n6912 gnd.n6911 19.3944
R11160 gnd.n6911 gnd.n6910 19.3944
R11161 gnd.n6910 gnd.n1110 19.3944
R11162 gnd.n6904 gnd.n1110 19.3944
R11163 gnd.n6904 gnd.n6903 19.3944
R11164 gnd.n6903 gnd.n6902 19.3944
R11165 gnd.n6902 gnd.n1118 19.3944
R11166 gnd.n6896 gnd.n1118 19.3944
R11167 gnd.n6896 gnd.n6895 19.3944
R11168 gnd.n6895 gnd.n6894 19.3944
R11169 gnd.n6894 gnd.n1126 19.3944
R11170 gnd.n6888 gnd.n1126 19.3944
R11171 gnd.n6888 gnd.n6887 19.3944
R11172 gnd.n6887 gnd.n6886 19.3944
R11173 gnd.n6886 gnd.n1134 19.3944
R11174 gnd.n2631 gnd.n2630 19.3944
R11175 gnd.n2630 gnd.n2629 19.3944
R11176 gnd.n2629 gnd.n2585 19.3944
R11177 gnd.n2625 gnd.n2585 19.3944
R11178 gnd.n2625 gnd.n2624 19.3944
R11179 gnd.n2624 gnd.n2623 19.3944
R11180 gnd.n2623 gnd.n2589 19.3944
R11181 gnd.n2619 gnd.n2589 19.3944
R11182 gnd.n2619 gnd.n2618 19.3944
R11183 gnd.n2618 gnd.n2617 19.3944
R11184 gnd.n2617 gnd.n2593 19.3944
R11185 gnd.n2613 gnd.n2593 19.3944
R11186 gnd.n2613 gnd.n2612 19.3944
R11187 gnd.n2612 gnd.n2611 19.3944
R11188 gnd.n2611 gnd.n2596 19.3944
R11189 gnd.n2607 gnd.n2596 19.3944
R11190 gnd.n2607 gnd.n2606 19.3944
R11191 gnd.n2606 gnd.n2605 19.3944
R11192 gnd.n2605 gnd.n2602 19.3944
R11193 gnd.n2602 gnd.n1706 19.3944
R11194 gnd.n4967 gnd.n1706 19.3944
R11195 gnd.n4967 gnd.n1707 19.3944
R11196 gnd.n4963 gnd.n1707 19.3944
R11197 gnd.n4963 gnd.n4962 19.3944
R11198 gnd.n4962 gnd.n4961 19.3944
R11199 gnd.n4961 gnd.n1713 19.3944
R11200 gnd.n4957 gnd.n1713 19.3944
R11201 gnd.n4957 gnd.n4956 19.3944
R11202 gnd.n4956 gnd.n4955 19.3944
R11203 gnd.n4955 gnd.n1718 19.3944
R11204 gnd.n4951 gnd.n1718 19.3944
R11205 gnd.n4951 gnd.n4950 19.3944
R11206 gnd.n4950 gnd.n4949 19.3944
R11207 gnd.n4949 gnd.n1723 19.3944
R11208 gnd.n4945 gnd.n1723 19.3944
R11209 gnd.n4945 gnd.n4944 19.3944
R11210 gnd.n4944 gnd.n4943 19.3944
R11211 gnd.n4943 gnd.n1728 19.3944
R11212 gnd.n4939 gnd.n1728 19.3944
R11213 gnd.n4939 gnd.n4938 19.3944
R11214 gnd.n4938 gnd.n4937 19.3944
R11215 gnd.n4937 gnd.n1733 19.3944
R11216 gnd.n4933 gnd.n1733 19.3944
R11217 gnd.n4933 gnd.n4932 19.3944
R11218 gnd.n4932 gnd.n4931 19.3944
R11219 gnd.n4931 gnd.n1738 19.3944
R11220 gnd.n4927 gnd.n1738 19.3944
R11221 gnd.n4927 gnd.n4926 19.3944
R11222 gnd.n4926 gnd.n4925 19.3944
R11223 gnd.n4925 gnd.n1743 19.3944
R11224 gnd.n4921 gnd.n1743 19.3944
R11225 gnd.n4921 gnd.n4920 19.3944
R11226 gnd.n4920 gnd.n4919 19.3944
R11227 gnd.n4919 gnd.n1748 19.3944
R11228 gnd.n4915 gnd.n1748 19.3944
R11229 gnd.n4915 gnd.n4914 19.3944
R11230 gnd.n4914 gnd.n4913 19.3944
R11231 gnd.n4913 gnd.n1753 19.3944
R11232 gnd.n4909 gnd.n1753 19.3944
R11233 gnd.n4909 gnd.n4908 19.3944
R11234 gnd.n4908 gnd.n4907 19.3944
R11235 gnd.n4907 gnd.n1758 19.3944
R11236 gnd.n4903 gnd.n1758 19.3944
R11237 gnd.n4903 gnd.n4902 19.3944
R11238 gnd.n4902 gnd.n4901 19.3944
R11239 gnd.n4901 gnd.n1763 19.3944
R11240 gnd.n4897 gnd.n1763 19.3944
R11241 gnd.n4897 gnd.n4896 19.3944
R11242 gnd.n4896 gnd.n4895 19.3944
R11243 gnd.n4895 gnd.n1768 19.3944
R11244 gnd.n4891 gnd.n1768 19.3944
R11245 gnd.n4891 gnd.n4890 19.3944
R11246 gnd.n4890 gnd.n4889 19.3944
R11247 gnd.n4889 gnd.n1773 19.3944
R11248 gnd.n4885 gnd.n1773 19.3944
R11249 gnd.n4885 gnd.n4884 19.3944
R11250 gnd.n4884 gnd.n4883 19.3944
R11251 gnd.n4883 gnd.n1778 19.3944
R11252 gnd.n4879 gnd.n1778 19.3944
R11253 gnd.n4879 gnd.n4878 19.3944
R11254 gnd.n4878 gnd.n4877 19.3944
R11255 gnd.n4877 gnd.n1783 19.3944
R11256 gnd.n4873 gnd.n1783 19.3944
R11257 gnd.n4873 gnd.n4872 19.3944
R11258 gnd.n4872 gnd.n4871 19.3944
R11259 gnd.n4871 gnd.n1788 19.3944
R11260 gnd.n4867 gnd.n1788 19.3944
R11261 gnd.n4867 gnd.n4866 19.3944
R11262 gnd.n4866 gnd.n4865 19.3944
R11263 gnd.n4865 gnd.n1793 19.3944
R11264 gnd.n4861 gnd.n1793 19.3944
R11265 gnd.n4861 gnd.n4860 19.3944
R11266 gnd.n4860 gnd.n4859 19.3944
R11267 gnd.n4859 gnd.n1798 19.3944
R11268 gnd.n4855 gnd.n1798 19.3944
R11269 gnd.n4855 gnd.n4854 19.3944
R11270 gnd.n4854 gnd.n4853 19.3944
R11271 gnd.n4853 gnd.n1803 19.3944
R11272 gnd.n4849 gnd.n1803 19.3944
R11273 gnd.n4849 gnd.n4848 19.3944
R11274 gnd.n4848 gnd.n4847 19.3944
R11275 gnd.n4455 gnd.n4452 19.3944
R11276 gnd.n4455 gnd.n4450 19.3944
R11277 gnd.n4461 gnd.n4450 19.3944
R11278 gnd.n4461 gnd.n4448 19.3944
R11279 gnd.n4466 gnd.n4448 19.3944
R11280 gnd.n4466 gnd.n4446 19.3944
R11281 gnd.n4472 gnd.n4446 19.3944
R11282 gnd.n4472 gnd.n4445 19.3944
R11283 gnd.n4483 gnd.n4445 19.3944
R11284 gnd.n4483 gnd.n4443 19.3944
R11285 gnd.n4489 gnd.n4443 19.3944
R11286 gnd.n4489 gnd.n4438 19.3944
R11287 gnd.n4502 gnd.n4438 19.3944
R11288 gnd.n4502 gnd.n4436 19.3944
R11289 gnd.n4508 gnd.n4436 19.3944
R11290 gnd.n4508 gnd.n4431 19.3944
R11291 gnd.n4521 gnd.n4431 19.3944
R11292 gnd.n4521 gnd.n4429 19.3944
R11293 gnd.n4527 gnd.n4429 19.3944
R11294 gnd.n4527 gnd.n4423 19.3944
R11295 gnd.n4540 gnd.n4423 19.3944
R11296 gnd.n4540 gnd.n4421 19.3944
R11297 gnd.n4545 gnd.n4421 19.3944
R11298 gnd.n4546 gnd.n4545 19.3944
R11299 gnd.n4556 gnd.n4408 19.3944
R11300 gnd.n4564 gnd.n4408 19.3944
R11301 gnd.n4564 gnd.n4563 19.3944
R11302 gnd.t28 gnd.n4033 19.1199
R11303 gnd.n3949 gnd.t6 19.1199
R11304 gnd.t34 gnd.n5924 18.8012
R11305 gnd.n6578 gnd.t403 18.8012
R11306 gnd.n6422 gnd.n6019 18.4825
R11307 gnd.n4147 gnd.n2346 18.4825
R11308 gnd.n4187 gnd.n2309 18.4825
R11309 gnd.n3980 gnd.n2282 18.4825
R11310 gnd.n3608 gnd.n2255 18.4825
R11311 gnd.n4784 gnd.n4783 18.4247
R11312 gnd.n5050 gnd.n5049 18.4247
R11313 gnd.n4979 gnd.n4978 18.2639
R11314 gnd.n3727 gnd.n3725 18.2639
R11315 gnd.n4553 gnd.n4552 18.2308
R11316 gnd.n3291 gnd.n2552 18.2308
R11317 gnd.n454 gnd.n451 18.2308
R11318 gnd.n2954 gnd.n2953 18.2308
R11319 gnd.n6494 gnd.t4 18.1639
R11320 gnd.n3456 gnd.t137 17.8452
R11321 gnd.n6475 gnd.t22 17.5266
R11322 gnd.n219 gnd.n211 17.5266
R11323 gnd.n4975 gnd.n1688 17.2079
R11324 gnd.n3463 gnd.t70 17.2079
R11325 gnd.n3495 gnd.n2365 17.2079
R11326 gnd.n4139 gnd.n2353 17.2079
R11327 gnd.n4195 gnd.n2302 17.2079
R11328 gnd.n3568 gnd.n3566 17.2079
R11329 gnd.n3936 gnd.n3935 17.2079
R11330 gnd.n4275 gnd.n2235 17.2079
R11331 gnd.n4339 gnd.t147 17.2079
R11332 gnd.n5952 gnd.t402 16.8893
R11333 gnd.t14 gnd.n2352 16.8893
R11334 gnd.n3934 gnd.t38 16.8893
R11335 gnd.n4766 gnd.n4763 16.6793
R11336 gnd.n7931 gnd.n7928 16.6793
R11337 gnd.n5327 gnd.n5324 16.6793
R11338 gnd.n2683 gnd.n2682 16.6793
R11339 gnd.t58 gnd.n6046 16.2519
R11340 gnd.n5909 gnd.t54 16.2519
R11341 gnd.n4050 gnd.n4049 15.9333
R11342 gnd.n4027 gnd.t178 15.9333
R11343 gnd.n3996 gnd.n2295 15.9333
R11344 gnd.n4203 gnd.n2295 15.9333
R11345 gnd.t23 gnd.n2261 15.9333
R11346 gnd.n4267 gnd.n2242 15.9333
R11347 gnd.n5726 gnd.n5724 15.6674
R11348 gnd.n5694 gnd.n5692 15.6674
R11349 gnd.n5662 gnd.n5660 15.6674
R11350 gnd.n5631 gnd.n5629 15.6674
R11351 gnd.n5599 gnd.n5597 15.6674
R11352 gnd.n5567 gnd.n5565 15.6674
R11353 gnd.n5535 gnd.n5533 15.6674
R11354 gnd.n5504 gnd.n5502 15.6674
R11355 gnd.n6164 gnd.t58 15.6146
R11356 gnd.n6786 gnd.t140 15.6146
R11357 gnd.n4723 gnd.n1925 15.3217
R11358 gnd.n7886 gnd.n351 15.3217
R11359 gnd.n5284 gnd.n1251 15.3217
R11360 gnd.n2734 gnd.n2732 15.3217
R11361 gnd.n3710 gnd.n3709 15.0827
R11362 gnd.n1674 gnd.n1669 15.0481
R11363 gnd.n3720 gnd.n3719 15.0481
R11364 gnd.n6683 gnd.t407 14.9773
R11365 gnd.n3455 gnd.t46 14.9773
R11366 gnd.n4323 gnd.t55 14.9773
R11367 gnd.n4975 gnd.n4974 14.6587
R11368 gnd.n4123 gnd.n2365 14.6587
R11369 gnd.n3631 gnd.n2235 14.6587
R11370 gnd.n3884 gnd.n3883 14.6587
R11371 gnd.n6715 gnd.t16 14.34
R11372 gnd.n6748 gnd.t52 14.34
R11373 gnd.n8029 gnd.n219 14.34
R11374 gnd.n4070 gnd.t2 14.0214
R11375 gnd.t177 gnd.n2221 14.0214
R11376 gnd.t396 gnd.n5958 13.7027
R11377 gnd.t203 gnd.n2824 13.7027
R11378 gnd.t242 gnd.n105 13.7027
R11379 gnd.n6391 gnd.n6387 13.5763
R11380 gnd.n6842 gnd.n5432 13.5763
R11381 gnd.n6423 gnd.n6422 13.384
R11382 gnd.t109 gnd.n1701 13.384
R11383 gnd.n4115 gnd.n2372 13.384
R11384 gnd.n4131 gnd.t20 13.384
R11385 gnd.n3517 gnd.n2346 13.384
R11386 gnd.n4012 gnd.n2309 13.384
R11387 gnd.n4219 gnd.n2282 13.384
R11388 gnd.n4251 gnd.n2255 13.384
R11389 gnd.n3622 gnd.t27 13.384
R11390 gnd.n3914 gnd.n3638 13.384
R11391 gnd.t106 gnd.n2200 13.384
R11392 gnd.n3659 gnd.n3657 13.384
R11393 gnd.n1685 gnd.n1666 13.1884
R11394 gnd.n1680 gnd.n1679 13.1884
R11395 gnd.n1679 gnd.n1678 13.1884
R11396 gnd.n3713 gnd.n3708 13.1884
R11397 gnd.n3714 gnd.n3713 13.1884
R11398 gnd.n1681 gnd.n1668 13.146
R11399 gnd.n1677 gnd.n1668 13.146
R11400 gnd.n3712 gnd.n3711 13.146
R11401 gnd.n3712 gnd.n3707 13.146
R11402 gnd.n3084 gnd.t235 13.0654
R11403 gnd.t244 gnd.n526 13.0654
R11404 gnd.n5727 gnd.n5723 12.8005
R11405 gnd.n5695 gnd.n5691 12.8005
R11406 gnd.n5663 gnd.n5659 12.8005
R11407 gnd.n5632 gnd.n5628 12.8005
R11408 gnd.n5600 gnd.n5596 12.8005
R11409 gnd.n5568 gnd.n5564 12.8005
R11410 gnd.n5536 gnd.n5532 12.8005
R11411 gnd.n5505 gnd.n5501 12.8005
R11412 gnd.n5252 gnd.t262 12.4281
R11413 gnd.n3143 gnd.t270 12.4281
R11414 gnd.n5131 gnd.t293 12.4281
R11415 gnd.t187 gnd.n2515 12.4281
R11416 gnd.n2156 gnd.t410 12.4281
R11417 gnd.n4689 gnd.t232 12.4281
R11418 gnd.n4641 gnd.t191 12.4281
R11419 gnd.n8035 gnd.t217 12.4281
R11420 gnd.n6394 gnd.n6391 12.4126
R11421 gnd.n6847 gnd.n5432 12.4126
R11422 gnd.n5042 gnd.n4979 12.1761
R11423 gnd.n3730 gnd.n3725 12.1761
R11424 gnd.n5099 gnd.n1556 12.1094
R11425 gnd.n4107 gnd.n2379 12.1094
R11426 gnd.n3526 gnd.n2339 12.1094
R11427 gnd.n3545 gnd.n2316 12.1094
R11428 gnd.n4227 gnd.n2275 12.1094
R11429 gnd.n4243 gnd.n2262 12.1094
R11430 gnd.n3646 gnd.n2222 12.1094
R11431 gnd.n3670 gnd.n2199 12.1094
R11432 gnd.n4836 gnd.n1859 12.1094
R11433 gnd.n5731 gnd.n5730 12.0247
R11434 gnd.n5699 gnd.n5698 12.0247
R11435 gnd.n5667 gnd.n5666 12.0247
R11436 gnd.n5636 gnd.n5635 12.0247
R11437 gnd.n5604 gnd.n5603 12.0247
R11438 gnd.n5572 gnd.n5571 12.0247
R11439 gnd.n5540 gnd.n5539 12.0247
R11440 gnd.n5509 gnd.n5508 12.0247
R11441 gnd.n5228 gnd.t237 11.7908
R11442 gnd.n5155 gnd.t270 11.7908
R11443 gnd.n3185 gnd.t293 11.7908
R11444 gnd.n2120 gnd.t232 11.7908
R11445 gnd.n4665 gnd.t191 11.7908
R11446 gnd.n8059 gnd.t255 11.7908
R11447 gnd.n5734 gnd.n5721 11.249
R11448 gnd.n5702 gnd.n5689 11.249
R11449 gnd.n5670 gnd.n5657 11.249
R11450 gnd.n5639 gnd.n5626 11.249
R11451 gnd.n5607 gnd.n5594 11.249
R11452 gnd.n5575 gnd.n5562 11.249
R11453 gnd.n5543 gnd.n5530 11.249
R11454 gnd.n5512 gnd.n5499 11.249
R11455 gnd.n6495 gnd.t396 11.1535
R11456 gnd.n5204 gnd.t253 11.1535
R11457 gnd.n5192 gnd.n1396 11.1535
R11458 gnd.n5179 gnd.t235 11.1535
R11459 gnd.n7750 gnd.t244 11.1535
R11460 gnd.n7721 gnd.n107 11.1535
R11461 gnd.n8083 gnd.t213 11.1535
R11462 gnd.n4091 gnd.t165 10.8348
R11463 gnd.t80 gnd.n2385 10.8348
R11464 gnd.n4099 gnd.n2385 10.8348
R11465 gnd.t179 gnd.n2353 10.8348
R11466 gnd.n2333 gnd.n2332 10.8348
R11467 gnd.n2332 gnd.n2323 10.8348
R11468 gnd.n4235 gnd.n2268 10.8348
R11469 gnd.n4235 gnd.n2269 10.8348
R11470 gnd.n3936 gnd.t33 10.8348
R11471 gnd.n2214 gnd.n2206 10.8348
R11472 gnd.n3883 gnd.t74 10.8348
R11473 gnd.n4726 gnd.n4723 10.6672
R11474 gnd.n7889 gnd.n7886 10.6672
R11475 gnd.n5287 gnd.n5284 10.6672
R11476 gnd.n2732 gnd.n2731 10.6672
R11477 gnd.n3873 gnd.n3872 10.6151
R11478 gnd.n3872 gnd.n3869 10.6151
R11479 gnd.n3867 gnd.n3864 10.6151
R11480 gnd.n3864 gnd.n3863 10.6151
R11481 gnd.n3863 gnd.n3860 10.6151
R11482 gnd.n3860 gnd.n3859 10.6151
R11483 gnd.n3859 gnd.n3856 10.6151
R11484 gnd.n3856 gnd.n3855 10.6151
R11485 gnd.n3855 gnd.n3852 10.6151
R11486 gnd.n3852 gnd.n3851 10.6151
R11487 gnd.n3851 gnd.n3848 10.6151
R11488 gnd.n3848 gnd.n3847 10.6151
R11489 gnd.n3847 gnd.n3844 10.6151
R11490 gnd.n3844 gnd.n3843 10.6151
R11491 gnd.n3843 gnd.n3840 10.6151
R11492 gnd.n3840 gnd.n3839 10.6151
R11493 gnd.n3839 gnd.n3836 10.6151
R11494 gnd.n3836 gnd.n3835 10.6151
R11495 gnd.n3835 gnd.n3832 10.6151
R11496 gnd.n3832 gnd.n3831 10.6151
R11497 gnd.n3831 gnd.n3828 10.6151
R11498 gnd.n3828 gnd.n3827 10.6151
R11499 gnd.n3827 gnd.n3824 10.6151
R11500 gnd.n3824 gnd.n3823 10.6151
R11501 gnd.n3823 gnd.n3820 10.6151
R11502 gnd.n3820 gnd.n3819 10.6151
R11503 gnd.n3819 gnd.n3816 10.6151
R11504 gnd.n3816 gnd.n3815 10.6151
R11505 gnd.n3815 gnd.n3685 10.6151
R11506 gnd.n3879 gnd.n3685 10.6151
R11507 gnd.n2476 gnd.n2475 10.6151
R11508 gnd.n2477 gnd.n2476 10.6151
R11509 gnd.n2481 gnd.n2477 10.6151
R11510 gnd.n2481 gnd.n2480 10.6151
R11511 gnd.n2480 gnd.n2479 10.6151
R11512 gnd.n2479 gnd.n2402 10.6151
R11513 gnd.n3467 gnd.n2402 10.6151
R11514 gnd.n3468 gnd.n3467 10.6151
R11515 gnd.n3469 gnd.n3468 10.6151
R11516 gnd.n3472 gnd.n3469 10.6151
R11517 gnd.n3473 gnd.n3472 10.6151
R11518 gnd.n4075 gnd.n3473 10.6151
R11519 gnd.n4075 gnd.n4074 10.6151
R11520 gnd.n4074 gnd.n4073 10.6151
R11521 gnd.n4073 gnd.n3474 10.6151
R11522 gnd.n3489 gnd.n3474 10.6151
R11523 gnd.n3491 gnd.n3489 10.6151
R11524 gnd.n3492 gnd.n3491 10.6151
R11525 gnd.n4060 gnd.n3492 10.6151
R11526 gnd.n4060 gnd.n4059 10.6151
R11527 gnd.n4059 gnd.n4058 10.6151
R11528 gnd.n4058 gnd.n3493 10.6151
R11529 gnd.n3505 gnd.n3493 10.6151
R11530 gnd.n4046 gnd.n3505 10.6151
R11531 gnd.n4046 gnd.n4045 10.6151
R11532 gnd.n4045 gnd.n4044 10.6151
R11533 gnd.n4044 gnd.n3506 10.6151
R11534 gnd.n3520 gnd.n3506 10.6151
R11535 gnd.n3522 gnd.n3520 10.6151
R11536 gnd.n3523 gnd.n3522 10.6151
R11537 gnd.n4031 gnd.n3523 10.6151
R11538 gnd.n4031 gnd.n4030 10.6151
R11539 gnd.n4030 gnd.n4029 10.6151
R11540 gnd.n4029 gnd.n3524 10.6151
R11541 gnd.n3541 gnd.n3524 10.6151
R11542 gnd.n3542 gnd.n3541 10.6151
R11543 gnd.n3543 gnd.n3542 10.6151
R11544 gnd.n3543 gnd.n3538 10.6151
R11545 gnd.n3549 gnd.n3538 10.6151
R11546 gnd.n3550 gnd.n3549 10.6151
R11547 gnd.n4009 gnd.n3550 10.6151
R11548 gnd.n4009 gnd.n4008 10.6151
R11549 gnd.n4008 gnd.n4007 10.6151
R11550 gnd.n4007 gnd.n3551 10.6151
R11551 gnd.n3562 gnd.n3551 10.6151
R11552 gnd.n3563 gnd.n3562 10.6151
R11553 gnd.n3993 gnd.n3563 10.6151
R11554 gnd.n3993 gnd.n3992 10.6151
R11555 gnd.n3992 gnd.n3991 10.6151
R11556 gnd.n3991 gnd.n3564 10.6151
R11557 gnd.n3576 gnd.n3564 10.6151
R11558 gnd.n3577 gnd.n3576 10.6151
R11559 gnd.n3977 gnd.n3577 10.6151
R11560 gnd.n3977 gnd.n3976 10.6151
R11561 gnd.n3976 gnd.n3975 10.6151
R11562 gnd.n3975 gnd.n3578 10.6151
R11563 gnd.n3589 gnd.n3578 10.6151
R11564 gnd.n3590 gnd.n3589 10.6151
R11565 gnd.n3961 gnd.n3590 10.6151
R11566 gnd.n3961 gnd.n3960 10.6151
R11567 gnd.n3960 gnd.n3959 10.6151
R11568 gnd.n3959 gnd.n3591 10.6151
R11569 gnd.n3604 gnd.n3591 10.6151
R11570 gnd.n3605 gnd.n3604 10.6151
R11571 gnd.n3947 gnd.n3605 10.6151
R11572 gnd.n3947 gnd.n3946 10.6151
R11573 gnd.n3946 gnd.n3945 10.6151
R11574 gnd.n3945 gnd.n3606 10.6151
R11575 gnd.n3618 gnd.n3606 10.6151
R11576 gnd.n3619 gnd.n3618 10.6151
R11577 gnd.n3932 gnd.n3619 10.6151
R11578 gnd.n3932 gnd.n3931 10.6151
R11579 gnd.n3931 gnd.n3930 10.6151
R11580 gnd.n3930 gnd.n3620 10.6151
R11581 gnd.n3634 gnd.n3620 10.6151
R11582 gnd.n3635 gnd.n3634 10.6151
R11583 gnd.n3918 gnd.n3635 10.6151
R11584 gnd.n3918 gnd.n3917 10.6151
R11585 gnd.n3917 gnd.n3916 10.6151
R11586 gnd.n3916 gnd.n3636 10.6151
R11587 gnd.n3650 gnd.n3636 10.6151
R11588 gnd.n3651 gnd.n3650 10.6151
R11589 gnd.n3904 gnd.n3651 10.6151
R11590 gnd.n3904 gnd.n3903 10.6151
R11591 gnd.n3903 gnd.n3902 10.6151
R11592 gnd.n3902 gnd.n3652 10.6151
R11593 gnd.n3898 gnd.n3652 10.6151
R11594 gnd.n3898 gnd.n3897 10.6151
R11595 gnd.n3897 gnd.n3896 10.6151
R11596 gnd.n3896 gnd.n3654 10.6151
R11597 gnd.n3656 gnd.n3654 10.6151
R11598 gnd.n3681 gnd.n3656 10.6151
R11599 gnd.n3683 gnd.n3681 10.6151
R11600 gnd.n3684 gnd.n3683 10.6151
R11601 gnd.n3881 gnd.n3684 10.6151
R11602 gnd.n3881 gnd.n3880 10.6151
R11603 gnd.n2410 gnd.n1626 10.6151
R11604 gnd.n2413 gnd.n2410 10.6151
R11605 gnd.n2418 gnd.n2415 10.6151
R11606 gnd.n2419 gnd.n2418 10.6151
R11607 gnd.n2422 gnd.n2419 10.6151
R11608 gnd.n2423 gnd.n2422 10.6151
R11609 gnd.n2426 gnd.n2423 10.6151
R11610 gnd.n2427 gnd.n2426 10.6151
R11611 gnd.n2430 gnd.n2427 10.6151
R11612 gnd.n2431 gnd.n2430 10.6151
R11613 gnd.n2434 gnd.n2431 10.6151
R11614 gnd.n2435 gnd.n2434 10.6151
R11615 gnd.n2438 gnd.n2435 10.6151
R11616 gnd.n2439 gnd.n2438 10.6151
R11617 gnd.n2442 gnd.n2439 10.6151
R11618 gnd.n2443 gnd.n2442 10.6151
R11619 gnd.n2446 gnd.n2443 10.6151
R11620 gnd.n2447 gnd.n2446 10.6151
R11621 gnd.n2450 gnd.n2447 10.6151
R11622 gnd.n2451 gnd.n2450 10.6151
R11623 gnd.n2454 gnd.n2451 10.6151
R11624 gnd.n2455 gnd.n2454 10.6151
R11625 gnd.n2458 gnd.n2455 10.6151
R11626 gnd.n2459 gnd.n2458 10.6151
R11627 gnd.n2462 gnd.n2459 10.6151
R11628 gnd.n2463 gnd.n2462 10.6151
R11629 gnd.n2466 gnd.n2463 10.6151
R11630 gnd.n2467 gnd.n2466 10.6151
R11631 gnd.n2470 gnd.n2467 10.6151
R11632 gnd.n2471 gnd.n2470 10.6151
R11633 gnd.n5042 gnd.n5041 10.6151
R11634 gnd.n5041 gnd.n5040 10.6151
R11635 gnd.n5040 gnd.n5039 10.6151
R11636 gnd.n5039 gnd.n5037 10.6151
R11637 gnd.n5037 gnd.n5034 10.6151
R11638 gnd.n5034 gnd.n5033 10.6151
R11639 gnd.n5033 gnd.n5030 10.6151
R11640 gnd.n5030 gnd.n5029 10.6151
R11641 gnd.n5029 gnd.n5026 10.6151
R11642 gnd.n5026 gnd.n5025 10.6151
R11643 gnd.n5025 gnd.n5022 10.6151
R11644 gnd.n5022 gnd.n5021 10.6151
R11645 gnd.n5021 gnd.n5018 10.6151
R11646 gnd.n5018 gnd.n5017 10.6151
R11647 gnd.n5017 gnd.n5014 10.6151
R11648 gnd.n5014 gnd.n5013 10.6151
R11649 gnd.n5013 gnd.n5010 10.6151
R11650 gnd.n5010 gnd.n5009 10.6151
R11651 gnd.n5009 gnd.n5006 10.6151
R11652 gnd.n5006 gnd.n5005 10.6151
R11653 gnd.n5005 gnd.n5002 10.6151
R11654 gnd.n5002 gnd.n5001 10.6151
R11655 gnd.n5001 gnd.n4998 10.6151
R11656 gnd.n4998 gnd.n4997 10.6151
R11657 gnd.n4997 gnd.n4994 10.6151
R11658 gnd.n4994 gnd.n4993 10.6151
R11659 gnd.n4993 gnd.n4990 10.6151
R11660 gnd.n4990 gnd.n4989 10.6151
R11661 gnd.n4986 gnd.n4985 10.6151
R11662 gnd.n4985 gnd.n1627 10.6151
R11663 gnd.n3731 gnd.n3730 10.6151
R11664 gnd.n3734 gnd.n3731 10.6151
R11665 gnd.n3735 gnd.n3734 10.6151
R11666 gnd.n3738 gnd.n3735 10.6151
R11667 gnd.n3739 gnd.n3738 10.6151
R11668 gnd.n3742 gnd.n3739 10.6151
R11669 gnd.n3743 gnd.n3742 10.6151
R11670 gnd.n3746 gnd.n3743 10.6151
R11671 gnd.n3747 gnd.n3746 10.6151
R11672 gnd.n3750 gnd.n3747 10.6151
R11673 gnd.n3751 gnd.n3750 10.6151
R11674 gnd.n3754 gnd.n3751 10.6151
R11675 gnd.n3755 gnd.n3754 10.6151
R11676 gnd.n3758 gnd.n3755 10.6151
R11677 gnd.n3759 gnd.n3758 10.6151
R11678 gnd.n3762 gnd.n3759 10.6151
R11679 gnd.n3763 gnd.n3762 10.6151
R11680 gnd.n3766 gnd.n3763 10.6151
R11681 gnd.n3767 gnd.n3766 10.6151
R11682 gnd.n3770 gnd.n3767 10.6151
R11683 gnd.n3771 gnd.n3770 10.6151
R11684 gnd.n3774 gnd.n3771 10.6151
R11685 gnd.n3775 gnd.n3774 10.6151
R11686 gnd.n3778 gnd.n3775 10.6151
R11687 gnd.n3779 gnd.n3778 10.6151
R11688 gnd.n3782 gnd.n3779 10.6151
R11689 gnd.n3783 gnd.n3782 10.6151
R11690 gnd.n3786 gnd.n3783 10.6151
R11691 gnd.n3791 gnd.n3788 10.6151
R11692 gnd.n3792 gnd.n3791 10.6151
R11693 gnd.n4978 gnd.n4977 10.6151
R11694 gnd.n4977 gnd.n1686 10.6151
R11695 gnd.n2405 gnd.n1686 10.6151
R11696 gnd.n3459 gnd.n2405 10.6151
R11697 gnd.n3460 gnd.n3459 10.6151
R11698 gnd.n3461 gnd.n3460 10.6151
R11699 gnd.n3461 gnd.n2396 10.6151
R11700 gnd.n4084 gnd.n2396 10.6151
R11701 gnd.n4084 gnd.n4083 10.6151
R11702 gnd.n4083 gnd.n4082 10.6151
R11703 gnd.n4082 gnd.n2397 10.6151
R11704 gnd.n3479 gnd.n2397 10.6151
R11705 gnd.n3481 gnd.n3479 10.6151
R11706 gnd.n3482 gnd.n3481 10.6151
R11707 gnd.n4068 gnd.n3482 10.6151
R11708 gnd.n4068 gnd.n4067 10.6151
R11709 gnd.n4067 gnd.n4066 10.6151
R11710 gnd.n4066 gnd.n3483 10.6151
R11711 gnd.n3498 gnd.n3483 10.6151
R11712 gnd.n3499 gnd.n3498 10.6151
R11713 gnd.n4054 gnd.n3499 10.6151
R11714 gnd.n4054 gnd.n4053 10.6151
R11715 gnd.n4053 gnd.n4052 10.6151
R11716 gnd.n4052 gnd.n3500 10.6151
R11717 gnd.n3512 gnd.n3500 10.6151
R11718 gnd.n3513 gnd.n3512 10.6151
R11719 gnd.n4039 gnd.n3513 10.6151
R11720 gnd.n4039 gnd.n4038 10.6151
R11721 gnd.n4038 gnd.n4037 10.6151
R11722 gnd.n4037 gnd.n3514 10.6151
R11723 gnd.n3529 gnd.n3514 10.6151
R11724 gnd.n3530 gnd.n3529 10.6151
R11725 gnd.n4025 gnd.n3530 10.6151
R11726 gnd.n4025 gnd.n4024 10.6151
R11727 gnd.n4024 gnd.n4023 10.6151
R11728 gnd.n4023 gnd.n3531 10.6151
R11729 gnd.n4019 gnd.n3531 10.6151
R11730 gnd.n4019 gnd.n4018 10.6151
R11731 gnd.n4018 gnd.n4017 10.6151
R11732 gnd.n4017 gnd.n3533 10.6151
R11733 gnd.n3535 gnd.n3533 10.6151
R11734 gnd.n3556 gnd.n3535 10.6151
R11735 gnd.n3557 gnd.n3556 10.6151
R11736 gnd.n4002 gnd.n3557 10.6151
R11737 gnd.n4002 gnd.n4001 10.6151
R11738 gnd.n4001 gnd.n4000 10.6151
R11739 gnd.n4000 gnd.n3558 10.6151
R11740 gnd.n3570 gnd.n3558 10.6151
R11741 gnd.n3571 gnd.n3570 10.6151
R11742 gnd.n3986 gnd.n3571 10.6151
R11743 gnd.n3986 gnd.n3985 10.6151
R11744 gnd.n3985 gnd.n3984 10.6151
R11745 gnd.n3984 gnd.n3572 10.6151
R11746 gnd.n3583 gnd.n3572 10.6151
R11747 gnd.n3584 gnd.n3583 10.6151
R11748 gnd.n3970 gnd.n3584 10.6151
R11749 gnd.n3970 gnd.n3969 10.6151
R11750 gnd.n3969 gnd.n3968 10.6151
R11751 gnd.n3968 gnd.n3585 10.6151
R11752 gnd.n3596 gnd.n3585 10.6151
R11753 gnd.n3597 gnd.n3596 10.6151
R11754 gnd.n3954 gnd.n3597 10.6151
R11755 gnd.n3954 gnd.n3953 10.6151
R11756 gnd.n3953 gnd.n3952 10.6151
R11757 gnd.n3952 gnd.n3598 10.6151
R11758 gnd.n3611 gnd.n3598 10.6151
R11759 gnd.n3612 gnd.n3611 10.6151
R11760 gnd.n3940 gnd.n3612 10.6151
R11761 gnd.n3940 gnd.n3939 10.6151
R11762 gnd.n3939 gnd.n3938 10.6151
R11763 gnd.n3938 gnd.n3613 10.6151
R11764 gnd.n3626 gnd.n3613 10.6151
R11765 gnd.n3627 gnd.n3626 10.6151
R11766 gnd.n3925 gnd.n3627 10.6151
R11767 gnd.n3925 gnd.n3924 10.6151
R11768 gnd.n3924 gnd.n3923 10.6151
R11769 gnd.n3923 gnd.n3628 10.6151
R11770 gnd.n3641 gnd.n3628 10.6151
R11771 gnd.n3912 gnd.n3641 10.6151
R11772 gnd.n3912 gnd.n3911 10.6151
R11773 gnd.n3911 gnd.n3910 10.6151
R11774 gnd.n3910 gnd.n3642 10.6151
R11775 gnd.n3644 gnd.n3642 10.6151
R11776 gnd.n3663 gnd.n3644 10.6151
R11777 gnd.n3665 gnd.n3663 10.6151
R11778 gnd.n3666 gnd.n3665 10.6151
R11779 gnd.n3667 gnd.n3666 10.6151
R11780 gnd.n3667 gnd.n3661 10.6151
R11781 gnd.n3674 gnd.n3661 10.6151
R11782 gnd.n3675 gnd.n3674 10.6151
R11783 gnd.n3890 gnd.n3675 10.6151
R11784 gnd.n3890 gnd.n3889 10.6151
R11785 gnd.n3889 gnd.n3888 10.6151
R11786 gnd.n3888 gnd.n3676 10.6151
R11787 gnd.n3726 gnd.n3676 10.6151
R11788 gnd.n3727 gnd.n3726 10.6151
R11789 gnd.n6034 gnd.t408 10.5161
R11790 gnd.n6738 gnd.t16 10.5161
R11791 gnd.t52 gnd.n5768 10.5161
R11792 gnd.n2881 gnd.t203 10.5161
R11793 gnd.n7822 gnd.t242 10.5161
R11794 gnd.n5735 gnd.n5719 10.4732
R11795 gnd.n5703 gnd.n5687 10.4732
R11796 gnd.n5671 gnd.n5655 10.4732
R11797 gnd.n5640 gnd.n5624 10.4732
R11798 gnd.n5608 gnd.n5592 10.4732
R11799 gnd.n5576 gnd.n5560 10.4732
R11800 gnd.n5544 gnd.n5528 10.4732
R11801 gnd.n5513 gnd.n5497 10.4732
R11802 gnd.n2392 gnd.t80 10.1975
R11803 gnd.n6693 gnd.t407 9.87883
R11804 gnd.n5210 gnd.t205 9.87883
R11805 gnd.n5045 gnd.n1662 9.87883
R11806 gnd.t48 gnd.t12 9.87883
R11807 gnd.t398 gnd.t394 9.87883
R11808 gnd.n3876 gnd.n3687 9.87883
R11809 gnd.n8077 gnd.t295 9.87883
R11810 gnd.n5739 gnd.n5738 9.69747
R11811 gnd.n5707 gnd.n5706 9.69747
R11812 gnd.n5675 gnd.n5674 9.69747
R11813 gnd.n5644 gnd.n5643 9.69747
R11814 gnd.n5612 gnd.n5611 9.69747
R11815 gnd.n5580 gnd.n5579 9.69747
R11816 gnd.n5548 gnd.n5547 9.69747
R11817 gnd.n5517 gnd.n5516 9.69747
R11818 gnd.n4091 gnd.n4086 9.56018
R11819 gnd.n4107 gnd.n2378 9.56018
R11820 gnd.n4027 gnd.n3526 9.56018
R11821 gnd.n3546 gnd.n3545 9.56018
R11822 gnd.n4227 gnd.n2276 9.56018
R11823 gnd.n4243 gnd.n2261 9.56018
R11824 gnd.n3906 gnd.n3646 9.56018
R11825 gnd.n5745 gnd.n5744 9.45567
R11826 gnd.n5713 gnd.n5712 9.45567
R11827 gnd.n5681 gnd.n5680 9.45567
R11828 gnd.n5650 gnd.n5649 9.45567
R11829 gnd.n5618 gnd.n5617 9.45567
R11830 gnd.n5586 gnd.n5585 9.45567
R11831 gnd.n5554 gnd.n5553 9.45567
R11832 gnd.n5523 gnd.n5522 9.45567
R11833 gnd.n4763 gnd.n4762 9.30959
R11834 gnd.n7928 gnd.n331 9.30959
R11835 gnd.n5324 gnd.n5323 9.30959
R11836 gnd.n2686 gnd.n2683 9.30959
R11837 gnd.n5744 gnd.n5743 9.3005
R11838 gnd.n5717 gnd.n5716 9.3005
R11839 gnd.n5738 gnd.n5737 9.3005
R11840 gnd.n5736 gnd.n5735 9.3005
R11841 gnd.n5721 gnd.n5720 9.3005
R11842 gnd.n5730 gnd.n5729 9.3005
R11843 gnd.n5728 gnd.n5727 9.3005
R11844 gnd.n5712 gnd.n5711 9.3005
R11845 gnd.n5685 gnd.n5684 9.3005
R11846 gnd.n5706 gnd.n5705 9.3005
R11847 gnd.n5704 gnd.n5703 9.3005
R11848 gnd.n5689 gnd.n5688 9.3005
R11849 gnd.n5698 gnd.n5697 9.3005
R11850 gnd.n5696 gnd.n5695 9.3005
R11851 gnd.n5680 gnd.n5679 9.3005
R11852 gnd.n5653 gnd.n5652 9.3005
R11853 gnd.n5674 gnd.n5673 9.3005
R11854 gnd.n5672 gnd.n5671 9.3005
R11855 gnd.n5657 gnd.n5656 9.3005
R11856 gnd.n5666 gnd.n5665 9.3005
R11857 gnd.n5664 gnd.n5663 9.3005
R11858 gnd.n5649 gnd.n5648 9.3005
R11859 gnd.n5622 gnd.n5621 9.3005
R11860 gnd.n5643 gnd.n5642 9.3005
R11861 gnd.n5641 gnd.n5640 9.3005
R11862 gnd.n5626 gnd.n5625 9.3005
R11863 gnd.n5635 gnd.n5634 9.3005
R11864 gnd.n5633 gnd.n5632 9.3005
R11865 gnd.n5617 gnd.n5616 9.3005
R11866 gnd.n5590 gnd.n5589 9.3005
R11867 gnd.n5611 gnd.n5610 9.3005
R11868 gnd.n5609 gnd.n5608 9.3005
R11869 gnd.n5594 gnd.n5593 9.3005
R11870 gnd.n5603 gnd.n5602 9.3005
R11871 gnd.n5601 gnd.n5600 9.3005
R11872 gnd.n5585 gnd.n5584 9.3005
R11873 gnd.n5558 gnd.n5557 9.3005
R11874 gnd.n5579 gnd.n5578 9.3005
R11875 gnd.n5577 gnd.n5576 9.3005
R11876 gnd.n5562 gnd.n5561 9.3005
R11877 gnd.n5571 gnd.n5570 9.3005
R11878 gnd.n5569 gnd.n5568 9.3005
R11879 gnd.n5553 gnd.n5552 9.3005
R11880 gnd.n5526 gnd.n5525 9.3005
R11881 gnd.n5547 gnd.n5546 9.3005
R11882 gnd.n5545 gnd.n5544 9.3005
R11883 gnd.n5530 gnd.n5529 9.3005
R11884 gnd.n5539 gnd.n5538 9.3005
R11885 gnd.n5537 gnd.n5536 9.3005
R11886 gnd.n5522 gnd.n5521 9.3005
R11887 gnd.n5495 gnd.n5494 9.3005
R11888 gnd.n5516 gnd.n5515 9.3005
R11889 gnd.n5514 gnd.n5513 9.3005
R11890 gnd.n5499 gnd.n5498 9.3005
R11891 gnd.n5508 gnd.n5507 9.3005
R11892 gnd.n5506 gnd.n5505 9.3005
R11893 gnd.n6869 gnd.n5406 9.3005
R11894 gnd.n6868 gnd.n5408 9.3005
R11895 gnd.n5412 gnd.n5409 9.3005
R11896 gnd.n6863 gnd.n5413 9.3005
R11897 gnd.n6862 gnd.n5414 9.3005
R11898 gnd.n6861 gnd.n5415 9.3005
R11899 gnd.n5419 gnd.n5416 9.3005
R11900 gnd.n6856 gnd.n5420 9.3005
R11901 gnd.n6855 gnd.n5421 9.3005
R11902 gnd.n6854 gnd.n5422 9.3005
R11903 gnd.n5426 gnd.n5423 9.3005
R11904 gnd.n6849 gnd.n5427 9.3005
R11905 gnd.n6848 gnd.n5428 9.3005
R11906 gnd.n6847 gnd.n5429 9.3005
R11907 gnd.n5434 gnd.n5432 9.3005
R11908 gnd.n6842 gnd.n6841 9.3005
R11909 gnd.n6871 gnd.n6870 9.3005
R11910 gnd.n6447 gnd.n6446 9.3005
R11911 gnd.n6448 gnd.n6005 9.3005
R11912 gnd.n6452 gnd.n6449 9.3005
R11913 gnd.n6451 gnd.n6450 9.3005
R11914 gnd.n5982 gnd.n5981 9.3005
R11915 gnd.n6478 gnd.n6477 9.3005
R11916 gnd.n6479 gnd.n5980 9.3005
R11917 gnd.n6483 gnd.n6480 9.3005
R11918 gnd.n6482 gnd.n6481 9.3005
R11919 gnd.n5956 gnd.n5955 9.3005
R11920 gnd.n6509 gnd.n6508 9.3005
R11921 gnd.n6510 gnd.n5954 9.3005
R11922 gnd.n6514 gnd.n6511 9.3005
R11923 gnd.n6513 gnd.n6512 9.3005
R11924 gnd.n5930 gnd.n5929 9.3005
R11925 gnd.n6540 gnd.n6539 9.3005
R11926 gnd.n6541 gnd.n5928 9.3005
R11927 gnd.n6545 gnd.n6542 9.3005
R11928 gnd.n6544 gnd.n6543 9.3005
R11929 gnd.n5904 gnd.n5903 9.3005
R11930 gnd.n6571 gnd.n6570 9.3005
R11931 gnd.n6572 gnd.n5902 9.3005
R11932 gnd.n6576 gnd.n6573 9.3005
R11933 gnd.n6575 gnd.n6574 9.3005
R11934 gnd.n5879 gnd.n5878 9.3005
R11935 gnd.n6602 gnd.n6601 9.3005
R11936 gnd.n6603 gnd.n5877 9.3005
R11937 gnd.n6607 gnd.n6604 9.3005
R11938 gnd.n6606 gnd.n6605 9.3005
R11939 gnd.n5855 gnd.n5854 9.3005
R11940 gnd.n6632 gnd.n6631 9.3005
R11941 gnd.n6633 gnd.n5853 9.3005
R11942 gnd.n6637 gnd.n6634 9.3005
R11943 gnd.n6636 gnd.n6635 9.3005
R11944 gnd.n5823 gnd.n5822 9.3005
R11945 gnd.n6673 gnd.n6672 9.3005
R11946 gnd.n6674 gnd.n5821 9.3005
R11947 gnd.n6681 gnd.n6675 9.3005
R11948 gnd.n6680 gnd.n6676 9.3005
R11949 gnd.n6679 gnd.n6677 9.3005
R11950 gnd.n5793 gnd.n5792 9.3005
R11951 gnd.n6720 gnd.n6719 9.3005
R11952 gnd.n6721 gnd.n5791 9.3005
R11953 gnd.n6727 gnd.n6722 9.3005
R11954 gnd.n6726 gnd.n6723 9.3005
R11955 gnd.n6725 gnd.n6724 9.3005
R11956 gnd.n5766 gnd.n5765 9.3005
R11957 gnd.n6764 gnd.n6763 9.3005
R11958 gnd.n6765 gnd.n5764 9.3005
R11959 gnd.n6769 gnd.n6766 9.3005
R11960 gnd.n6768 gnd.n6767 9.3005
R11961 gnd.n5405 gnd.n5404 9.3005
R11962 gnd.n6873 gnd.n6872 9.3005
R11963 gnd.n6007 gnd.n6006 9.3005
R11964 gnd.n6391 gnd.n6390 9.3005
R11965 gnd.n6394 gnd.n6386 9.3005
R11966 gnd.n6395 gnd.n6385 9.3005
R11967 gnd.n6398 gnd.n6384 9.3005
R11968 gnd.n6399 gnd.n6383 9.3005
R11969 gnd.n6402 gnd.n6382 9.3005
R11970 gnd.n6403 gnd.n6381 9.3005
R11971 gnd.n6406 gnd.n6380 9.3005
R11972 gnd.n6407 gnd.n6379 9.3005
R11973 gnd.n6410 gnd.n6378 9.3005
R11974 gnd.n6411 gnd.n6377 9.3005
R11975 gnd.n6414 gnd.n6376 9.3005
R11976 gnd.n6416 gnd.n6375 9.3005
R11977 gnd.n6417 gnd.n6374 9.3005
R11978 gnd.n6418 gnd.n6373 9.3005
R11979 gnd.n6419 gnd.n6372 9.3005
R11980 gnd.n6387 gnd.n6023 9.3005
R11981 gnd.n6437 gnd.n6436 9.3005
R11982 gnd.n6438 gnd.n6000 9.3005
R11983 gnd.n6457 gnd.n6456 9.3005
R11984 gnd.n6459 gnd.n5992 9.3005
R11985 gnd.n6466 gnd.n5993 9.3005
R11986 gnd.n6468 gnd.n6467 9.3005
R11987 gnd.n6469 gnd.n5973 9.3005
R11988 gnd.n6488 gnd.n6487 9.3005
R11989 gnd.n6490 gnd.n5966 9.3005
R11990 gnd.n6497 gnd.n5967 9.3005
R11991 gnd.n6499 gnd.n6498 9.3005
R11992 gnd.n6500 gnd.n5947 9.3005
R11993 gnd.n6519 gnd.n6518 9.3005
R11994 gnd.n6521 gnd.n5940 9.3005
R11995 gnd.n6528 gnd.n5941 9.3005
R11996 gnd.n6530 gnd.n6529 9.3005
R11997 gnd.n6531 gnd.n5922 9.3005
R11998 gnd.n6550 gnd.n6549 9.3005
R11999 gnd.n6552 gnd.n5914 9.3005
R12000 gnd.n6559 gnd.n5915 9.3005
R12001 gnd.n6561 gnd.n6560 9.3005
R12002 gnd.n6562 gnd.n5897 9.3005
R12003 gnd.n6581 gnd.n6580 9.3005
R12004 gnd.n6583 gnd.n5889 9.3005
R12005 gnd.n6590 gnd.n5890 9.3005
R12006 gnd.n6592 gnd.n6591 9.3005
R12007 gnd.n6593 gnd.n5872 9.3005
R12008 gnd.n6612 gnd.n6611 9.3005
R12009 gnd.n6614 gnd.n5864 9.3005
R12010 gnd.n6621 gnd.n5865 9.3005
R12011 gnd.n6623 gnd.n6622 9.3005
R12012 gnd.n6624 gnd.n5848 9.3005
R12013 gnd.n6642 gnd.n6641 9.3005
R12014 gnd.n6644 gnd.n5833 9.3005
R12015 gnd.n6662 gnd.n5835 9.3005
R12016 gnd.n6663 gnd.n5830 9.3005
R12017 gnd.n6665 gnd.n6664 9.3005
R12018 gnd.n5831 gnd.n5817 9.3005
R12019 gnd.n5815 gnd.n5813 9.3005
R12020 gnd.n6688 gnd.n6687 9.3005
R12021 gnd.n5798 gnd.n5797 9.3005
R12022 gnd.n6713 gnd.n6709 9.3005
R12023 gnd.n6712 gnd.n6711 9.3005
R12024 gnd.n5786 gnd.n5784 9.3005
R12025 gnd.n6733 gnd.n6732 9.3005
R12026 gnd.n5771 gnd.n5770 9.3005
R12027 gnd.n6757 gnd.n6756 9.3005
R12028 gnd.n6754 gnd.n5750 9.3005
R12029 gnd.n6775 gnd.n6774 9.3005
R12030 gnd.n5752 gnd.n5751 9.3005
R12031 gnd.n5759 gnd.n5755 9.3005
R12032 gnd.n5758 gnd.n5756 9.3005
R12033 gnd.n5757 gnd.n5435 9.3005
R12034 gnd.n6435 gnd.n6017 9.3005
R12035 gnd.n6837 gnd.n5436 9.3005
R12036 gnd.n6836 gnd.n5438 9.3005
R12037 gnd.n5442 gnd.n5439 9.3005
R12038 gnd.n6831 gnd.n5443 9.3005
R12039 gnd.n6830 gnd.n5444 9.3005
R12040 gnd.n6829 gnd.n5445 9.3005
R12041 gnd.n5449 gnd.n5446 9.3005
R12042 gnd.n6824 gnd.n5450 9.3005
R12043 gnd.n6823 gnd.n5451 9.3005
R12044 gnd.n6822 gnd.n5452 9.3005
R12045 gnd.n5456 gnd.n5453 9.3005
R12046 gnd.n6817 gnd.n5457 9.3005
R12047 gnd.n6816 gnd.n5458 9.3005
R12048 gnd.n6815 gnd.n5459 9.3005
R12049 gnd.n5463 gnd.n5460 9.3005
R12050 gnd.n6810 gnd.n5464 9.3005
R12051 gnd.n6809 gnd.n5465 9.3005
R12052 gnd.n6808 gnd.n5466 9.3005
R12053 gnd.n5470 gnd.n5467 9.3005
R12054 gnd.n6803 gnd.n5471 9.3005
R12055 gnd.n6802 gnd.n5472 9.3005
R12056 gnd.n6801 gnd.n5473 9.3005
R12057 gnd.n5480 gnd.n5478 9.3005
R12058 gnd.n6796 gnd.n5481 9.3005
R12059 gnd.n6795 gnd.n5482 9.3005
R12060 gnd.n6794 gnd.n6791 9.3005
R12061 gnd.n6839 gnd.n6838 9.3005
R12062 gnd.n6234 gnd.n6213 9.3005
R12063 gnd.n6233 gnd.n6215 9.3005
R12064 gnd.n6231 gnd.n6216 9.3005
R12065 gnd.n6230 gnd.n6217 9.3005
R12066 gnd.n6226 gnd.n6218 9.3005
R12067 gnd.n6225 gnd.n6219 9.3005
R12068 gnd.n6224 gnd.n6220 9.3005
R12069 gnd.n6222 gnd.n6221 9.3005
R12070 gnd.n5841 gnd.n5840 9.3005
R12071 gnd.n6652 gnd.n6651 9.3005
R12072 gnd.n6653 gnd.n5839 9.3005
R12073 gnd.n6657 gnd.n6654 9.3005
R12074 gnd.n6656 gnd.n6655 9.3005
R12075 gnd.n5806 gnd.n5805 9.3005
R12076 gnd.n6696 gnd.n6695 9.3005
R12077 gnd.n6697 gnd.n5804 9.3005
R12078 gnd.n6701 gnd.n6698 9.3005
R12079 gnd.n6700 gnd.n6699 9.3005
R12080 gnd.n5779 gnd.n5778 9.3005
R12081 gnd.n6741 gnd.n6740 9.3005
R12082 gnd.n6742 gnd.n5777 9.3005
R12083 gnd.n6746 gnd.n6743 9.3005
R12084 gnd.n6745 gnd.n6744 9.3005
R12085 gnd.n5486 gnd.n5485 9.3005
R12086 gnd.n6782 gnd.n6781 9.3005
R12087 gnd.n6783 gnd.n5484 9.3005
R12088 gnd.n6785 gnd.n6784 9.3005
R12089 gnd.n6788 gnd.n5483 9.3005
R12090 gnd.n6790 gnd.n6789 9.3005
R12091 gnd.n6160 gnd.n6054 9.3005
R12092 gnd.n6162 gnd.n6161 9.3005
R12093 gnd.n6044 gnd.n6043 9.3005
R12094 gnd.n6175 gnd.n6174 9.3005
R12095 gnd.n6176 gnd.n6042 9.3005
R12096 gnd.n6178 gnd.n6177 9.3005
R12097 gnd.n6031 gnd.n6030 9.3005
R12098 gnd.n6191 gnd.n6190 9.3005
R12099 gnd.n6192 gnd.n6029 9.3005
R12100 gnd.n6361 gnd.n6193 9.3005
R12101 gnd.n6360 gnd.n6194 9.3005
R12102 gnd.n6359 gnd.n6195 9.3005
R12103 gnd.n6358 gnd.n6196 9.3005
R12104 gnd.n6356 gnd.n6197 9.3005
R12105 gnd.n6355 gnd.n6198 9.3005
R12106 gnd.n6351 gnd.n6199 9.3005
R12107 gnd.n6350 gnd.n6200 9.3005
R12108 gnd.n6349 gnd.n6201 9.3005
R12109 gnd.n6347 gnd.n6202 9.3005
R12110 gnd.n6346 gnd.n6203 9.3005
R12111 gnd.n6343 gnd.n6204 9.3005
R12112 gnd.n6342 gnd.n6205 9.3005
R12113 gnd.n6341 gnd.n6206 9.3005
R12114 gnd.n6339 gnd.n6207 9.3005
R12115 gnd.n6338 gnd.n6208 9.3005
R12116 gnd.n6335 gnd.n6209 9.3005
R12117 gnd.n6334 gnd.n6210 9.3005
R12118 gnd.n6333 gnd.n6211 9.3005
R12119 gnd.n6159 gnd.n6158 9.3005
R12120 gnd.n6099 gnd.n6098 9.3005
R12121 gnd.n6104 gnd.n6096 9.3005
R12122 gnd.n6105 gnd.n6095 9.3005
R12123 gnd.n6107 gnd.n6092 9.3005
R12124 gnd.n6091 gnd.n6089 9.3005
R12125 gnd.n6113 gnd.n6088 9.3005
R12126 gnd.n6114 gnd.n6087 9.3005
R12127 gnd.n6115 gnd.n6086 9.3005
R12128 gnd.n6085 gnd.n6083 9.3005
R12129 gnd.n6121 gnd.n6082 9.3005
R12130 gnd.n6122 gnd.n6081 9.3005
R12131 gnd.n6123 gnd.n6080 9.3005
R12132 gnd.n6079 gnd.n6077 9.3005
R12133 gnd.n6129 gnd.n6076 9.3005
R12134 gnd.n6130 gnd.n6075 9.3005
R12135 gnd.n6131 gnd.n6074 9.3005
R12136 gnd.n6073 gnd.n6071 9.3005
R12137 gnd.n6137 gnd.n6070 9.3005
R12138 gnd.n6138 gnd.n6069 9.3005
R12139 gnd.n6139 gnd.n6068 9.3005
R12140 gnd.n6067 gnd.n6065 9.3005
R12141 gnd.n6144 gnd.n6064 9.3005
R12142 gnd.n6145 gnd.n6063 9.3005
R12143 gnd.n6062 gnd.n6060 9.3005
R12144 gnd.n6150 gnd.n6059 9.3005
R12145 gnd.n6152 gnd.n6151 9.3005
R12146 gnd.n6097 gnd.n6055 9.3005
R12147 gnd.n6050 gnd.n6049 9.3005
R12148 gnd.n6167 gnd.n6166 9.3005
R12149 gnd.n6168 gnd.n6048 9.3005
R12150 gnd.n6170 gnd.n6169 9.3005
R12151 gnd.n6038 gnd.n6037 9.3005
R12152 gnd.n6183 gnd.n6182 9.3005
R12153 gnd.n6184 gnd.n6036 9.3005
R12154 gnd.n6186 gnd.n6185 9.3005
R12155 gnd.n6025 gnd.n6024 9.3005
R12156 gnd.n6426 gnd.n6425 9.3005
R12157 gnd.n6428 gnd.n6022 9.3005
R12158 gnd.n6430 gnd.n6429 9.3005
R12159 gnd.n6016 gnd.n6015 9.3005
R12160 gnd.n6441 gnd.n6439 9.3005
R12161 gnd.n6440 gnd.n5999 9.3005
R12162 gnd.n6458 gnd.n5998 9.3005
R12163 gnd.n6461 gnd.n6460 9.3005
R12164 gnd.n5991 gnd.n5990 9.3005
R12165 gnd.n6472 gnd.n6470 9.3005
R12166 gnd.n6471 gnd.n5972 9.3005
R12167 gnd.n6489 gnd.n5971 9.3005
R12168 gnd.n6492 gnd.n6491 9.3005
R12169 gnd.n5965 gnd.n5964 9.3005
R12170 gnd.n6503 gnd.n6501 9.3005
R12171 gnd.n6502 gnd.n5946 9.3005
R12172 gnd.n6520 gnd.n5945 9.3005
R12173 gnd.n6523 gnd.n6522 9.3005
R12174 gnd.n5939 gnd.n5938 9.3005
R12175 gnd.n6534 gnd.n6532 9.3005
R12176 gnd.n6533 gnd.n5921 9.3005
R12177 gnd.n6551 gnd.n5920 9.3005
R12178 gnd.n6554 gnd.n6553 9.3005
R12179 gnd.n5913 gnd.n5912 9.3005
R12180 gnd.n6565 gnd.n6563 9.3005
R12181 gnd.n6564 gnd.n5896 9.3005
R12182 gnd.n6582 gnd.n5895 9.3005
R12183 gnd.n6585 gnd.n6584 9.3005
R12184 gnd.n5888 gnd.n5887 9.3005
R12185 gnd.n6596 gnd.n6594 9.3005
R12186 gnd.n6595 gnd.n5871 9.3005
R12187 gnd.n6613 gnd.n5870 9.3005
R12188 gnd.n6616 gnd.n6615 9.3005
R12189 gnd.n5863 gnd.n5862 9.3005
R12190 gnd.n6626 gnd.n6625 9.3005
R12191 gnd.n5847 gnd.n5846 9.3005
R12192 gnd.n6647 gnd.n6643 9.3005
R12193 gnd.n6646 gnd.n6645 9.3005
R12194 gnd.n5834 gnd.n5829 9.3005
R12195 gnd.n6667 gnd.n6666 9.3005
R12196 gnd.n5832 gnd.n5811 9.3005
R12197 gnd.n6691 gnd.n5812 9.3005
R12198 gnd.n6690 gnd.n6689 9.3005
R12199 gnd.n5814 gnd.n5799 9.3005
R12200 gnd.n6708 gnd.n6707 9.3005
R12201 gnd.n6710 gnd.n5782 9.3005
R12202 gnd.n6736 gnd.n5783 9.3005
R12203 gnd.n6735 gnd.n6734 9.3005
R12204 gnd.n5785 gnd.n5772 9.3005
R12205 gnd.n6753 gnd.n6752 9.3005
R12206 gnd.n6755 gnd.n5492 9.3005
R12207 gnd.n6777 gnd.n6776 9.3005
R12208 gnd.n5749 gnd.n1140 9.3005
R12209 gnd.n6880 gnd.n1141 9.3005
R12210 gnd.n6879 gnd.n1142 9.3005
R12211 gnd.n6878 gnd.n1143 9.3005
R12212 gnd.n6154 gnd.n6153 9.3005
R12213 gnd.n7055 gnd.n7054 9.3005
R12214 gnd.n7056 gnd.n965 9.3005
R12215 gnd.n7058 gnd.n7057 9.3005
R12216 gnd.n961 gnd.n960 9.3005
R12217 gnd.n7065 gnd.n7064 9.3005
R12218 gnd.n7066 gnd.n959 9.3005
R12219 gnd.n7068 gnd.n7067 9.3005
R12220 gnd.n955 gnd.n954 9.3005
R12221 gnd.n7075 gnd.n7074 9.3005
R12222 gnd.n7076 gnd.n953 9.3005
R12223 gnd.n7078 gnd.n7077 9.3005
R12224 gnd.n949 gnd.n948 9.3005
R12225 gnd.n7085 gnd.n7084 9.3005
R12226 gnd.n7086 gnd.n947 9.3005
R12227 gnd.n7088 gnd.n7087 9.3005
R12228 gnd.n943 gnd.n942 9.3005
R12229 gnd.n7095 gnd.n7094 9.3005
R12230 gnd.n7096 gnd.n941 9.3005
R12231 gnd.n7098 gnd.n7097 9.3005
R12232 gnd.n937 gnd.n936 9.3005
R12233 gnd.n7105 gnd.n7104 9.3005
R12234 gnd.n7106 gnd.n935 9.3005
R12235 gnd.n7108 gnd.n7107 9.3005
R12236 gnd.n931 gnd.n930 9.3005
R12237 gnd.n7115 gnd.n7114 9.3005
R12238 gnd.n7116 gnd.n929 9.3005
R12239 gnd.n7118 gnd.n7117 9.3005
R12240 gnd.n925 gnd.n924 9.3005
R12241 gnd.n7125 gnd.n7124 9.3005
R12242 gnd.n7126 gnd.n923 9.3005
R12243 gnd.n7128 gnd.n7127 9.3005
R12244 gnd.n919 gnd.n918 9.3005
R12245 gnd.n7135 gnd.n7134 9.3005
R12246 gnd.n7136 gnd.n917 9.3005
R12247 gnd.n7138 gnd.n7137 9.3005
R12248 gnd.n913 gnd.n912 9.3005
R12249 gnd.n7145 gnd.n7144 9.3005
R12250 gnd.n7146 gnd.n911 9.3005
R12251 gnd.n7148 gnd.n7147 9.3005
R12252 gnd.n907 gnd.n906 9.3005
R12253 gnd.n7155 gnd.n7154 9.3005
R12254 gnd.n7156 gnd.n905 9.3005
R12255 gnd.n7158 gnd.n7157 9.3005
R12256 gnd.n901 gnd.n900 9.3005
R12257 gnd.n7165 gnd.n7164 9.3005
R12258 gnd.n7166 gnd.n899 9.3005
R12259 gnd.n7168 gnd.n7167 9.3005
R12260 gnd.n895 gnd.n894 9.3005
R12261 gnd.n7175 gnd.n7174 9.3005
R12262 gnd.n7176 gnd.n893 9.3005
R12263 gnd.n7178 gnd.n7177 9.3005
R12264 gnd.n889 gnd.n888 9.3005
R12265 gnd.n7185 gnd.n7184 9.3005
R12266 gnd.n7186 gnd.n887 9.3005
R12267 gnd.n7188 gnd.n7187 9.3005
R12268 gnd.n883 gnd.n882 9.3005
R12269 gnd.n7195 gnd.n7194 9.3005
R12270 gnd.n7196 gnd.n881 9.3005
R12271 gnd.n7198 gnd.n7197 9.3005
R12272 gnd.n877 gnd.n876 9.3005
R12273 gnd.n7205 gnd.n7204 9.3005
R12274 gnd.n7206 gnd.n875 9.3005
R12275 gnd.n7208 gnd.n7207 9.3005
R12276 gnd.n871 gnd.n870 9.3005
R12277 gnd.n7215 gnd.n7214 9.3005
R12278 gnd.n7216 gnd.n869 9.3005
R12279 gnd.n7218 gnd.n7217 9.3005
R12280 gnd.n865 gnd.n864 9.3005
R12281 gnd.n7225 gnd.n7224 9.3005
R12282 gnd.n7226 gnd.n863 9.3005
R12283 gnd.n7228 gnd.n7227 9.3005
R12284 gnd.n859 gnd.n858 9.3005
R12285 gnd.n7235 gnd.n7234 9.3005
R12286 gnd.n7236 gnd.n857 9.3005
R12287 gnd.n7238 gnd.n7237 9.3005
R12288 gnd.n853 gnd.n852 9.3005
R12289 gnd.n7245 gnd.n7244 9.3005
R12290 gnd.n7246 gnd.n851 9.3005
R12291 gnd.n7248 gnd.n7247 9.3005
R12292 gnd.n847 gnd.n846 9.3005
R12293 gnd.n7255 gnd.n7254 9.3005
R12294 gnd.n7256 gnd.n845 9.3005
R12295 gnd.n7258 gnd.n7257 9.3005
R12296 gnd.n841 gnd.n840 9.3005
R12297 gnd.n7265 gnd.n7264 9.3005
R12298 gnd.n7266 gnd.n839 9.3005
R12299 gnd.n7268 gnd.n7267 9.3005
R12300 gnd.n835 gnd.n834 9.3005
R12301 gnd.n7275 gnd.n7274 9.3005
R12302 gnd.n7276 gnd.n833 9.3005
R12303 gnd.n7278 gnd.n7277 9.3005
R12304 gnd.n829 gnd.n828 9.3005
R12305 gnd.n7285 gnd.n7284 9.3005
R12306 gnd.n7286 gnd.n827 9.3005
R12307 gnd.n7288 gnd.n7287 9.3005
R12308 gnd.n823 gnd.n822 9.3005
R12309 gnd.n7295 gnd.n7294 9.3005
R12310 gnd.n7296 gnd.n821 9.3005
R12311 gnd.n7298 gnd.n7297 9.3005
R12312 gnd.n817 gnd.n816 9.3005
R12313 gnd.n7305 gnd.n7304 9.3005
R12314 gnd.n7306 gnd.n815 9.3005
R12315 gnd.n7308 gnd.n7307 9.3005
R12316 gnd.n811 gnd.n810 9.3005
R12317 gnd.n7315 gnd.n7314 9.3005
R12318 gnd.n7316 gnd.n809 9.3005
R12319 gnd.n7318 gnd.n7317 9.3005
R12320 gnd.n805 gnd.n804 9.3005
R12321 gnd.n7325 gnd.n7324 9.3005
R12322 gnd.n7326 gnd.n803 9.3005
R12323 gnd.n7328 gnd.n7327 9.3005
R12324 gnd.n799 gnd.n798 9.3005
R12325 gnd.n7335 gnd.n7334 9.3005
R12326 gnd.n7336 gnd.n797 9.3005
R12327 gnd.n7338 gnd.n7337 9.3005
R12328 gnd.n793 gnd.n792 9.3005
R12329 gnd.n7345 gnd.n7344 9.3005
R12330 gnd.n7346 gnd.n791 9.3005
R12331 gnd.n7348 gnd.n7347 9.3005
R12332 gnd.n787 gnd.n786 9.3005
R12333 gnd.n7355 gnd.n7354 9.3005
R12334 gnd.n7356 gnd.n785 9.3005
R12335 gnd.n7358 gnd.n7357 9.3005
R12336 gnd.n781 gnd.n780 9.3005
R12337 gnd.n7365 gnd.n7364 9.3005
R12338 gnd.n7366 gnd.n779 9.3005
R12339 gnd.n7368 gnd.n7367 9.3005
R12340 gnd.n775 gnd.n774 9.3005
R12341 gnd.n7375 gnd.n7374 9.3005
R12342 gnd.n7376 gnd.n773 9.3005
R12343 gnd.n7378 gnd.n7377 9.3005
R12344 gnd.n769 gnd.n768 9.3005
R12345 gnd.n7385 gnd.n7384 9.3005
R12346 gnd.n7386 gnd.n767 9.3005
R12347 gnd.n7388 gnd.n7387 9.3005
R12348 gnd.n763 gnd.n762 9.3005
R12349 gnd.n7395 gnd.n7394 9.3005
R12350 gnd.n7396 gnd.n761 9.3005
R12351 gnd.n7398 gnd.n7397 9.3005
R12352 gnd.n757 gnd.n756 9.3005
R12353 gnd.n7405 gnd.n7404 9.3005
R12354 gnd.n7406 gnd.n755 9.3005
R12355 gnd.n7408 gnd.n7407 9.3005
R12356 gnd.n751 gnd.n750 9.3005
R12357 gnd.n7415 gnd.n7414 9.3005
R12358 gnd.n7416 gnd.n749 9.3005
R12359 gnd.n7418 gnd.n7417 9.3005
R12360 gnd.n745 gnd.n744 9.3005
R12361 gnd.n7425 gnd.n7424 9.3005
R12362 gnd.n7426 gnd.n743 9.3005
R12363 gnd.n7428 gnd.n7427 9.3005
R12364 gnd.n739 gnd.n738 9.3005
R12365 gnd.n7435 gnd.n7434 9.3005
R12366 gnd.n7436 gnd.n737 9.3005
R12367 gnd.n7438 gnd.n7437 9.3005
R12368 gnd.n733 gnd.n732 9.3005
R12369 gnd.n7445 gnd.n7444 9.3005
R12370 gnd.n7446 gnd.n731 9.3005
R12371 gnd.n7448 gnd.n7447 9.3005
R12372 gnd.n727 gnd.n726 9.3005
R12373 gnd.n7455 gnd.n7454 9.3005
R12374 gnd.n7456 gnd.n725 9.3005
R12375 gnd.n7458 gnd.n7457 9.3005
R12376 gnd.n721 gnd.n720 9.3005
R12377 gnd.n7465 gnd.n7464 9.3005
R12378 gnd.n7466 gnd.n719 9.3005
R12379 gnd.n7468 gnd.n7467 9.3005
R12380 gnd.n715 gnd.n714 9.3005
R12381 gnd.n7475 gnd.n7474 9.3005
R12382 gnd.n7476 gnd.n713 9.3005
R12383 gnd.n7478 gnd.n7477 9.3005
R12384 gnd.n709 gnd.n708 9.3005
R12385 gnd.n7485 gnd.n7484 9.3005
R12386 gnd.n7486 gnd.n707 9.3005
R12387 gnd.n7488 gnd.n7487 9.3005
R12388 gnd.n703 gnd.n702 9.3005
R12389 gnd.n7495 gnd.n7494 9.3005
R12390 gnd.n7496 gnd.n701 9.3005
R12391 gnd.n7499 gnd.n7498 9.3005
R12392 gnd.n7497 gnd.n697 9.3005
R12393 gnd.n7505 gnd.n696 9.3005
R12394 gnd.n7507 gnd.n7506 9.3005
R12395 gnd.n692 gnd.n691 9.3005
R12396 gnd.n7516 gnd.n7515 9.3005
R12397 gnd.n7517 gnd.n690 9.3005
R12398 gnd.n7519 gnd.n7518 9.3005
R12399 gnd.n686 gnd.n685 9.3005
R12400 gnd.n7526 gnd.n7525 9.3005
R12401 gnd.n7527 gnd.n684 9.3005
R12402 gnd.n7529 gnd.n7528 9.3005
R12403 gnd.n680 gnd.n679 9.3005
R12404 gnd.n7536 gnd.n7535 9.3005
R12405 gnd.n7537 gnd.n678 9.3005
R12406 gnd.n7539 gnd.n7538 9.3005
R12407 gnd.n674 gnd.n673 9.3005
R12408 gnd.n7546 gnd.n7545 9.3005
R12409 gnd.n7547 gnd.n672 9.3005
R12410 gnd.n7549 gnd.n7548 9.3005
R12411 gnd.n668 gnd.n667 9.3005
R12412 gnd.n7556 gnd.n7555 9.3005
R12413 gnd.n7557 gnd.n666 9.3005
R12414 gnd.n7559 gnd.n7558 9.3005
R12415 gnd.n662 gnd.n661 9.3005
R12416 gnd.n7566 gnd.n7565 9.3005
R12417 gnd.n7567 gnd.n660 9.3005
R12418 gnd.n7569 gnd.n7568 9.3005
R12419 gnd.n656 gnd.n655 9.3005
R12420 gnd.n7576 gnd.n7575 9.3005
R12421 gnd.n7577 gnd.n654 9.3005
R12422 gnd.n7579 gnd.n7578 9.3005
R12423 gnd.n650 gnd.n649 9.3005
R12424 gnd.n7586 gnd.n7585 9.3005
R12425 gnd.n7587 gnd.n648 9.3005
R12426 gnd.n7589 gnd.n7588 9.3005
R12427 gnd.n644 gnd.n643 9.3005
R12428 gnd.n7596 gnd.n7595 9.3005
R12429 gnd.n7597 gnd.n642 9.3005
R12430 gnd.n7599 gnd.n7598 9.3005
R12431 gnd.n638 gnd.n637 9.3005
R12432 gnd.n7606 gnd.n7605 9.3005
R12433 gnd.n7607 gnd.n636 9.3005
R12434 gnd.n7609 gnd.n7608 9.3005
R12435 gnd.n632 gnd.n631 9.3005
R12436 gnd.n7616 gnd.n7615 9.3005
R12437 gnd.n7617 gnd.n630 9.3005
R12438 gnd.n7619 gnd.n7618 9.3005
R12439 gnd.n626 gnd.n625 9.3005
R12440 gnd.n7626 gnd.n7625 9.3005
R12441 gnd.n7627 gnd.n624 9.3005
R12442 gnd.n7629 gnd.n7628 9.3005
R12443 gnd.n620 gnd.n619 9.3005
R12444 gnd.n7636 gnd.n7635 9.3005
R12445 gnd.n7637 gnd.n618 9.3005
R12446 gnd.n7639 gnd.n7638 9.3005
R12447 gnd.n614 gnd.n613 9.3005
R12448 gnd.n7646 gnd.n7645 9.3005
R12449 gnd.n7647 gnd.n612 9.3005
R12450 gnd.n7649 gnd.n7648 9.3005
R12451 gnd.n608 gnd.n607 9.3005
R12452 gnd.n7656 gnd.n7655 9.3005
R12453 gnd.n7657 gnd.n606 9.3005
R12454 gnd.n7659 gnd.n7658 9.3005
R12455 gnd.n602 gnd.n601 9.3005
R12456 gnd.n7666 gnd.n7665 9.3005
R12457 gnd.n7667 gnd.n600 9.3005
R12458 gnd.n7669 gnd.n7668 9.3005
R12459 gnd.n596 gnd.n595 9.3005
R12460 gnd.n7676 gnd.n7675 9.3005
R12461 gnd.n7677 gnd.n594 9.3005
R12462 gnd.n7679 gnd.n7678 9.3005
R12463 gnd.n590 gnd.n589 9.3005
R12464 gnd.n7686 gnd.n7685 9.3005
R12465 gnd.n7687 gnd.n588 9.3005
R12466 gnd.n7689 gnd.n7688 9.3005
R12467 gnd.n584 gnd.n583 9.3005
R12468 gnd.n7696 gnd.n7695 9.3005
R12469 gnd.n7697 gnd.n582 9.3005
R12470 gnd.n7699 gnd.n7698 9.3005
R12471 gnd.n578 gnd.n577 9.3005
R12472 gnd.n7706 gnd.n7705 9.3005
R12473 gnd.n7707 gnd.n576 9.3005
R12474 gnd.n7709 gnd.n7708 9.3005
R12475 gnd.n572 gnd.n571 9.3005
R12476 gnd.n7717 gnd.n7716 9.3005
R12477 gnd.n7718 gnd.n570 9.3005
R12478 gnd.n7720 gnd.n7719 9.3005
R12479 gnd.n7509 gnd.n7508 9.3005
R12480 gnd.n8101 gnd.n8100 9.3005
R12481 gnd.n8099 gnd.n101 9.3005
R12482 gnd.n388 gnd.n103 9.3005
R12483 gnd.n391 gnd.n390 9.3005
R12484 gnd.n392 gnd.n387 9.3005
R12485 gnd.n395 gnd.n393 9.3005
R12486 gnd.n396 gnd.n386 9.3005
R12487 gnd.n399 gnd.n398 9.3005
R12488 gnd.n400 gnd.n385 9.3005
R12489 gnd.n403 gnd.n401 9.3005
R12490 gnd.n404 gnd.n384 9.3005
R12491 gnd.n407 gnd.n406 9.3005
R12492 gnd.n408 gnd.n383 9.3005
R12493 gnd.n411 gnd.n409 9.3005
R12494 gnd.n412 gnd.n382 9.3005
R12495 gnd.n415 gnd.n414 9.3005
R12496 gnd.n416 gnd.n381 9.3005
R12497 gnd.n419 gnd.n417 9.3005
R12498 gnd.n420 gnd.n380 9.3005
R12499 gnd.n423 gnd.n422 9.3005
R12500 gnd.n424 gnd.n379 9.3005
R12501 gnd.n427 gnd.n425 9.3005
R12502 gnd.n428 gnd.n378 9.3005
R12503 gnd.n431 gnd.n430 9.3005
R12504 gnd.n432 gnd.n377 9.3005
R12505 gnd.n435 gnd.n433 9.3005
R12506 gnd.n436 gnd.n376 9.3005
R12507 gnd.n439 gnd.n438 9.3005
R12508 gnd.n440 gnd.n375 9.3005
R12509 gnd.n443 gnd.n441 9.3005
R12510 gnd.n444 gnd.n374 9.3005
R12511 gnd.n448 gnd.n447 9.3005
R12512 gnd.n483 gnd.n354 9.3005
R12513 gnd.n482 gnd.n356 9.3005
R12514 gnd.n479 gnd.n357 9.3005
R12515 gnd.n478 gnd.n358 9.3005
R12516 gnd.n475 gnd.n359 9.3005
R12517 gnd.n474 gnd.n360 9.3005
R12518 gnd.n471 gnd.n361 9.3005
R12519 gnd.n470 gnd.n362 9.3005
R12520 gnd.n467 gnd.n363 9.3005
R12521 gnd.n466 gnd.n364 9.3005
R12522 gnd.n463 gnd.n365 9.3005
R12523 gnd.n462 gnd.n366 9.3005
R12524 gnd.n459 gnd.n367 9.3005
R12525 gnd.n458 gnd.n368 9.3005
R12526 gnd.n455 gnd.n369 9.3005
R12527 gnd.n454 gnd.n370 9.3005
R12528 gnd.n451 gnd.n450 9.3005
R12529 gnd.n449 gnd.n371 9.3005
R12530 gnd.n485 gnd.n484 9.3005
R12531 gnd.n255 gnd.n254 9.3005
R12532 gnd.n8000 gnd.n296 9.3005
R12533 gnd.n7999 gnd.n297 9.3005
R12534 gnd.n7998 gnd.n298 9.3005
R12535 gnd.n7995 gnd.n299 9.3005
R12536 gnd.n7994 gnd.n300 9.3005
R12537 gnd.n7991 gnd.n301 9.3005
R12538 gnd.n7990 gnd.n302 9.3005
R12539 gnd.n7987 gnd.n303 9.3005
R12540 gnd.n7986 gnd.n304 9.3005
R12541 gnd.n7983 gnd.n305 9.3005
R12542 gnd.n7982 gnd.n306 9.3005
R12543 gnd.n7979 gnd.n307 9.3005
R12544 gnd.n7978 gnd.n308 9.3005
R12545 gnd.n7975 gnd.n309 9.3005
R12546 gnd.n7974 gnd.n310 9.3005
R12547 gnd.n7971 gnd.n311 9.3005
R12548 gnd.n7967 gnd.n312 9.3005
R12549 gnd.n7964 gnd.n313 9.3005
R12550 gnd.n7963 gnd.n314 9.3005
R12551 gnd.n7960 gnd.n315 9.3005
R12552 gnd.n7959 gnd.n316 9.3005
R12553 gnd.n7956 gnd.n317 9.3005
R12554 gnd.n7955 gnd.n318 9.3005
R12555 gnd.n7952 gnd.n319 9.3005
R12556 gnd.n7951 gnd.n320 9.3005
R12557 gnd.n7948 gnd.n321 9.3005
R12558 gnd.n7947 gnd.n322 9.3005
R12559 gnd.n7944 gnd.n323 9.3005
R12560 gnd.n7943 gnd.n324 9.3005
R12561 gnd.n7940 gnd.n325 9.3005
R12562 gnd.n7939 gnd.n326 9.3005
R12563 gnd.n7936 gnd.n327 9.3005
R12564 gnd.n7935 gnd.n328 9.3005
R12565 gnd.n7932 gnd.n329 9.3005
R12566 gnd.n7931 gnd.n330 9.3005
R12567 gnd.n7928 gnd.n7927 9.3005
R12568 gnd.n7926 gnd.n331 9.3005
R12569 gnd.n7925 gnd.n7924 9.3005
R12570 gnd.n7921 gnd.n334 9.3005
R12571 gnd.n7918 gnd.n335 9.3005
R12572 gnd.n7917 gnd.n336 9.3005
R12573 gnd.n7914 gnd.n337 9.3005
R12574 gnd.n7913 gnd.n338 9.3005
R12575 gnd.n7910 gnd.n339 9.3005
R12576 gnd.n7909 gnd.n340 9.3005
R12577 gnd.n7906 gnd.n341 9.3005
R12578 gnd.n7905 gnd.n342 9.3005
R12579 gnd.n7902 gnd.n343 9.3005
R12580 gnd.n7901 gnd.n344 9.3005
R12581 gnd.n7898 gnd.n345 9.3005
R12582 gnd.n7897 gnd.n346 9.3005
R12583 gnd.n7894 gnd.n347 9.3005
R12584 gnd.n7893 gnd.n348 9.3005
R12585 gnd.n7890 gnd.n349 9.3005
R12586 gnd.n7889 gnd.n350 9.3005
R12587 gnd.n7886 gnd.n7885 9.3005
R12588 gnd.n7884 gnd.n351 9.3005
R12589 gnd.n8006 gnd.n8005 9.3005
R12590 gnd.n1939 gnd.n1930 9.3005
R12591 gnd.n2129 gnd.n1955 9.3005
R12592 gnd.n4705 gnd.n1956 9.3005
R12593 gnd.n4704 gnd.n1957 9.3005
R12594 gnd.n4703 gnd.n1958 9.3005
R12595 gnd.n2125 gnd.n1959 9.3005
R12596 gnd.n4693 gnd.n1977 9.3005
R12597 gnd.n4692 gnd.n1978 9.3005
R12598 gnd.n4691 gnd.n1979 9.3005
R12599 gnd.n2062 gnd.n1980 9.3005
R12600 gnd.n4681 gnd.n1997 9.3005
R12601 gnd.n4680 gnd.n1998 9.3005
R12602 gnd.n4679 gnd.n1999 9.3005
R12603 gnd.n2057 gnd.n2000 9.3005
R12604 gnd.n4669 gnd.n2018 9.3005
R12605 gnd.n4668 gnd.n2019 9.3005
R12606 gnd.n4667 gnd.n2020 9.3005
R12607 gnd.n4619 gnd.n2021 9.3005
R12608 gnd.n4657 gnd.n2039 9.3005
R12609 gnd.n4656 gnd.n4655 9.3005
R12610 gnd.n2040 gnd.n547 9.3005
R12611 gnd.n7755 gnd.n548 9.3005
R12612 gnd.n7754 gnd.n549 9.3005
R12613 gnd.n7753 gnd.n7748 9.3005
R12614 gnd.n7752 gnd.n7749 9.3005
R12615 gnd.n524 gnd.n518 9.3005
R12616 gnd.n7788 gnd.n519 9.3005
R12617 gnd.n7787 gnd.n520 9.3005
R12618 gnd.n7786 gnd.n521 9.3005
R12619 gnd.n495 gnd.n494 9.3005
R12620 gnd.n7816 gnd.n7815 9.3005
R12621 gnd.n7817 gnd.n488 9.3005
R12622 gnd.n7824 gnd.n489 9.3005
R12623 gnd.n7825 gnd.n487 9.3005
R12624 gnd.n7828 gnd.n7827 9.3005
R12625 gnd.n7829 gnd.n128 9.3005
R12626 gnd.n8087 gnd.n129 9.3005
R12627 gnd.n8086 gnd.n130 9.3005
R12628 gnd.n8085 gnd.n131 9.3005
R12629 gnd.n7837 gnd.n132 9.3005
R12630 gnd.n8075 gnd.n146 9.3005
R12631 gnd.n8074 gnd.n147 9.3005
R12632 gnd.n8073 gnd.n148 9.3005
R12633 gnd.n7844 gnd.n149 9.3005
R12634 gnd.n8063 gnd.n166 9.3005
R12635 gnd.n8062 gnd.n167 9.3005
R12636 gnd.n8061 gnd.n168 9.3005
R12637 gnd.n7851 gnd.n169 9.3005
R12638 gnd.n8051 gnd.n184 9.3005
R12639 gnd.n8050 gnd.n185 9.3005
R12640 gnd.n8049 gnd.n186 9.3005
R12641 gnd.n7858 gnd.n187 9.3005
R12642 gnd.n8039 gnd.n204 9.3005
R12643 gnd.n8038 gnd.n205 9.3005
R12644 gnd.n8037 gnd.n206 9.3005
R12645 gnd.n7865 gnd.n207 9.3005
R12646 gnd.n8027 gnd.n223 9.3005
R12647 gnd.n8026 gnd.n224 9.3005
R12648 gnd.n8025 gnd.n225 9.3005
R12649 gnd.n7872 gnd.n226 9.3005
R12650 gnd.n8015 gnd.n243 9.3005
R12651 gnd.n8014 gnd.n244 9.3005
R12652 gnd.n8013 gnd.n245 9.3005
R12653 gnd.n7882 gnd.n246 9.3005
R12654 gnd.n4719 gnd.n1929 9.3005
R12655 gnd.n1931 gnd.n1930 9.3005
R12656 gnd.n4575 gnd.n2129 9.3005
R12657 gnd.n4576 gnd.n1956 9.3005
R12658 gnd.n4577 gnd.n1957 9.3005
R12659 gnd.n2124 gnd.n1958 9.3005
R12660 gnd.n4589 gnd.n2125 9.3005
R12661 gnd.n4590 gnd.n1977 9.3005
R12662 gnd.n4591 gnd.n1978 9.3005
R12663 gnd.n2061 gnd.n1979 9.3005
R12664 gnd.n4603 gnd.n2062 9.3005
R12665 gnd.n4604 gnd.n1997 9.3005
R12666 gnd.n4605 gnd.n1998 9.3005
R12667 gnd.n2056 gnd.n1999 9.3005
R12668 gnd.n4617 gnd.n2057 9.3005
R12669 gnd.n4618 gnd.n2018 9.3005
R12670 gnd.n4622 gnd.n2019 9.3005
R12671 gnd.n4621 gnd.n2020 9.3005
R12672 gnd.n4620 gnd.n4619 9.3005
R12673 gnd.n2041 gnd.n2039 9.3005
R12674 gnd.n4655 gnd.n4654 9.3005
R12675 gnd.n2042 gnd.n2040 9.3005
R12676 gnd.n550 gnd.n548 9.3005
R12677 gnd.n7746 gnd.n549 9.3005
R12678 gnd.n7748 gnd.n7747 9.3005
R12679 gnd.n7749 gnd.n523 9.3005
R12680 gnd.n7778 gnd.n524 9.3005
R12681 gnd.n7779 gnd.n519 9.3005
R12682 gnd.n7780 gnd.n520 9.3005
R12683 gnd.n7782 gnd.n521 9.3005
R12684 gnd.n7781 gnd.n494 9.3005
R12685 gnd.n7816 gnd.n493 9.3005
R12686 gnd.n7818 gnd.n7817 9.3005
R12687 gnd.n7820 gnd.n489 9.3005
R12688 gnd.n7819 gnd.n487 9.3005
R12689 gnd.n7828 gnd.n486 9.3005
R12690 gnd.n7832 gnd.n7829 9.3005
R12691 gnd.n7833 gnd.n129 9.3005
R12692 gnd.n7835 gnd.n130 9.3005
R12693 gnd.n7836 gnd.n131 9.3005
R12694 gnd.n7839 gnd.n7837 9.3005
R12695 gnd.n7840 gnd.n146 9.3005
R12696 gnd.n7842 gnd.n147 9.3005
R12697 gnd.n7843 gnd.n148 9.3005
R12698 gnd.n7846 gnd.n7844 9.3005
R12699 gnd.n7847 gnd.n166 9.3005
R12700 gnd.n7849 gnd.n167 9.3005
R12701 gnd.n7850 gnd.n168 9.3005
R12702 gnd.n7853 gnd.n7851 9.3005
R12703 gnd.n7854 gnd.n184 9.3005
R12704 gnd.n7856 gnd.n185 9.3005
R12705 gnd.n7857 gnd.n186 9.3005
R12706 gnd.n7860 gnd.n7858 9.3005
R12707 gnd.n7861 gnd.n204 9.3005
R12708 gnd.n7863 gnd.n205 9.3005
R12709 gnd.n7864 gnd.n206 9.3005
R12710 gnd.n7867 gnd.n7865 9.3005
R12711 gnd.n7868 gnd.n223 9.3005
R12712 gnd.n7870 gnd.n224 9.3005
R12713 gnd.n7871 gnd.n225 9.3005
R12714 gnd.n7874 gnd.n7872 9.3005
R12715 gnd.n7875 gnd.n243 9.3005
R12716 gnd.n7877 gnd.n244 9.3005
R12717 gnd.n7878 gnd.n245 9.3005
R12718 gnd.n7882 gnd.n7881 9.3005
R12719 gnd.n4719 gnd.n4718 9.3005
R12720 gnd.n4723 gnd.n4722 9.3005
R12721 gnd.n4726 gnd.n1924 9.3005
R12722 gnd.n4727 gnd.n1923 9.3005
R12723 gnd.n4730 gnd.n1922 9.3005
R12724 gnd.n4731 gnd.n1921 9.3005
R12725 gnd.n4734 gnd.n1920 9.3005
R12726 gnd.n4735 gnd.n1919 9.3005
R12727 gnd.n4738 gnd.n1918 9.3005
R12728 gnd.n4739 gnd.n1917 9.3005
R12729 gnd.n4742 gnd.n1916 9.3005
R12730 gnd.n4743 gnd.n1915 9.3005
R12731 gnd.n4746 gnd.n1914 9.3005
R12732 gnd.n4747 gnd.n1913 9.3005
R12733 gnd.n4750 gnd.n1912 9.3005
R12734 gnd.n4751 gnd.n1911 9.3005
R12735 gnd.n4754 gnd.n1910 9.3005
R12736 gnd.n4755 gnd.n1909 9.3005
R12737 gnd.n4758 gnd.n1908 9.3005
R12738 gnd.n4759 gnd.n1907 9.3005
R12739 gnd.n4762 gnd.n1906 9.3005
R12740 gnd.n4766 gnd.n1902 9.3005
R12741 gnd.n4767 gnd.n1901 9.3005
R12742 gnd.n4770 gnd.n1900 9.3005
R12743 gnd.n4771 gnd.n1899 9.3005
R12744 gnd.n4774 gnd.n1898 9.3005
R12745 gnd.n4775 gnd.n1897 9.3005
R12746 gnd.n4778 gnd.n1896 9.3005
R12747 gnd.n4779 gnd.n1895 9.3005
R12748 gnd.n4782 gnd.n1894 9.3005
R12749 gnd.n4784 gnd.n1890 9.3005
R12750 gnd.n4787 gnd.n1889 9.3005
R12751 gnd.n4788 gnd.n1888 9.3005
R12752 gnd.n4791 gnd.n1887 9.3005
R12753 gnd.n4792 gnd.n1886 9.3005
R12754 gnd.n4795 gnd.n1885 9.3005
R12755 gnd.n4796 gnd.n1884 9.3005
R12756 gnd.n4799 gnd.n1883 9.3005
R12757 gnd.n4801 gnd.n1880 9.3005
R12758 gnd.n4804 gnd.n1879 9.3005
R12759 gnd.n4805 gnd.n1878 9.3005
R12760 gnd.n4808 gnd.n1877 9.3005
R12761 gnd.n4809 gnd.n1876 9.3005
R12762 gnd.n4812 gnd.n1875 9.3005
R12763 gnd.n4813 gnd.n1874 9.3005
R12764 gnd.n4816 gnd.n1873 9.3005
R12765 gnd.n4817 gnd.n1872 9.3005
R12766 gnd.n4820 gnd.n1871 9.3005
R12767 gnd.n4821 gnd.n1870 9.3005
R12768 gnd.n4824 gnd.n1869 9.3005
R12769 gnd.n4825 gnd.n1868 9.3005
R12770 gnd.n4828 gnd.n1867 9.3005
R12771 gnd.n4830 gnd.n1866 9.3005
R12772 gnd.n4831 gnd.n1865 9.3005
R12773 gnd.n4832 gnd.n1864 9.3005
R12774 gnd.n4833 gnd.n1863 9.3005
R12775 gnd.n4763 gnd.n1903 9.3005
R12776 gnd.n4721 gnd.n1925 9.3005
R12777 gnd.n4711 gnd.n1945 9.3005
R12778 gnd.n4710 gnd.n1946 9.3005
R12779 gnd.n4709 gnd.n1947 9.3005
R12780 gnd.n1966 gnd.n1948 9.3005
R12781 gnd.n4699 gnd.n1967 9.3005
R12782 gnd.n4698 gnd.n1968 9.3005
R12783 gnd.n4697 gnd.n1969 9.3005
R12784 gnd.n1986 gnd.n1970 9.3005
R12785 gnd.n4687 gnd.n1987 9.3005
R12786 gnd.n4686 gnd.n1988 9.3005
R12787 gnd.n4685 gnd.n1989 9.3005
R12788 gnd.n2007 gnd.n1990 9.3005
R12789 gnd.n4675 gnd.n2008 9.3005
R12790 gnd.n4674 gnd.n2009 9.3005
R12791 gnd.n4673 gnd.n2010 9.3005
R12792 gnd.n2027 gnd.n2011 9.3005
R12793 gnd.n4663 gnd.n2028 9.3005
R12794 gnd.n4662 gnd.n2029 9.3005
R12795 gnd.n4661 gnd.n2030 9.3005
R12796 gnd.n2032 gnd.n2031 9.3005
R12797 gnd.n540 gnd.n539 9.3005
R12798 gnd.n7760 gnd.n7759 9.3005
R12799 gnd.n7761 gnd.n538 9.3005
R12800 gnd.n7766 gnd.n7762 9.3005
R12801 gnd.n7765 gnd.n7763 9.3005
R12802 gnd.n7764 gnd.n114 9.3005
R12803 gnd.n119 gnd.n113 9.3005
R12804 gnd.n8081 gnd.n138 9.3005
R12805 gnd.n8080 gnd.n139 9.3005
R12806 gnd.n8079 gnd.n140 9.3005
R12807 gnd.n155 gnd.n141 9.3005
R12808 gnd.n8069 gnd.n156 9.3005
R12809 gnd.n8068 gnd.n157 9.3005
R12810 gnd.n8067 gnd.n158 9.3005
R12811 gnd.n175 gnd.n159 9.3005
R12812 gnd.n8057 gnd.n176 9.3005
R12813 gnd.n8056 gnd.n177 9.3005
R12814 gnd.n8055 gnd.n178 9.3005
R12815 gnd.n193 gnd.n179 9.3005
R12816 gnd.n8045 gnd.n194 9.3005
R12817 gnd.n8044 gnd.n195 9.3005
R12818 gnd.n8043 gnd.n196 9.3005
R12819 gnd.n213 gnd.n197 9.3005
R12820 gnd.n8033 gnd.n214 9.3005
R12821 gnd.n8032 gnd.n215 9.3005
R12822 gnd.n8031 gnd.n216 9.3005
R12823 gnd.n233 gnd.n217 9.3005
R12824 gnd.n8021 gnd.n234 9.3005
R12825 gnd.n8020 gnd.n235 9.3005
R12826 gnd.n8019 gnd.n236 9.3005
R12827 gnd.n252 gnd.n237 9.3005
R12828 gnd.n8009 gnd.n253 9.3005
R12829 gnd.n8008 gnd.n8007 9.3005
R12830 gnd.n1944 gnd.n1943 9.3005
R12831 gnd.n8092 gnd.n8091 9.3005
R12832 gnd.n7734 gnd.n7733 9.3005
R12833 gnd.n7732 gnd.n561 9.3005
R12834 gnd.n7731 gnd.n7730 9.3005
R12835 gnd.n563 gnd.n562 9.3005
R12836 gnd.n7726 gnd.n566 9.3005
R12837 gnd.n7725 gnd.n567 9.3005
R12838 gnd.n7724 gnd.n568 9.3005
R12839 gnd.n3060 gnd.n2780 9.3005
R12840 gnd.n3082 gnd.n3061 9.3005
R12841 gnd.n3081 gnd.n3062 9.3005
R12842 gnd.n3080 gnd.n3063 9.3005
R12843 gnd.n3066 gnd.n3064 9.3005
R12844 gnd.n3076 gnd.n3067 9.3005
R12845 gnd.n3075 gnd.n3068 9.3005
R12846 gnd.n3074 gnd.n3069 9.3005
R12847 gnd.n3072 gnd.n3071 9.3005
R12848 gnd.n3070 gnd.n2757 9.3005
R12849 gnd.n2755 gnd.n2754 9.3005
R12850 gnd.n3148 gnd.n3147 9.3005
R12851 gnd.n3149 gnd.n2753 9.3005
R12852 gnd.n3151 gnd.n3150 9.3005
R12853 gnd.n2751 gnd.n2750 9.3005
R12854 gnd.n3156 gnd.n3155 9.3005
R12855 gnd.n3157 gnd.n2749 9.3005
R12856 gnd.n3183 gnd.n3158 9.3005
R12857 gnd.n3182 gnd.n3159 9.3005
R12858 gnd.n3181 gnd.n3160 9.3005
R12859 gnd.n3163 gnd.n3161 9.3005
R12860 gnd.n3177 gnd.n3164 9.3005
R12861 gnd.n3176 gnd.n3165 9.3005
R12862 gnd.n3175 gnd.n3166 9.3005
R12863 gnd.n3168 gnd.n3167 9.3005
R12864 gnd.n3171 gnd.n3170 9.3005
R12865 gnd.n3169 gnd.n2557 9.3005
R12866 gnd.n3358 gnd.n2558 9.3005
R12867 gnd.n3357 gnd.n2559 9.3005
R12868 gnd.n3356 gnd.n2560 9.3005
R12869 gnd.n2562 gnd.n2561 9.3005
R12870 gnd.n2564 gnd.n2563 9.3005
R12871 gnd.n2540 gnd.n2539 9.3005
R12872 gnd.n3376 gnd.n3375 9.3005
R12873 gnd.n3377 gnd.n2538 9.3005
R12874 gnd.n3379 gnd.n3378 9.3005
R12875 gnd.n2527 gnd.n2526 9.3005
R12876 gnd.n3392 gnd.n3391 9.3005
R12877 gnd.n3393 gnd.n2525 9.3005
R12878 gnd.n3395 gnd.n3394 9.3005
R12879 gnd.n2513 gnd.n2512 9.3005
R12880 gnd.n3408 gnd.n3407 9.3005
R12881 gnd.n3409 gnd.n2511 9.3005
R12882 gnd.n3411 gnd.n3410 9.3005
R12883 gnd.n2499 gnd.n2498 9.3005
R12884 gnd.n3424 gnd.n3423 9.3005
R12885 gnd.n3425 gnd.n2497 9.3005
R12886 gnd.n3436 gnd.n3426 9.3005
R12887 gnd.n3435 gnd.n3427 9.3005
R12888 gnd.n3434 gnd.n3428 9.3005
R12889 gnd.n3431 gnd.n3430 9.3005
R12890 gnd.n3429 gnd.n1695 9.3005
R12891 gnd.n4972 gnd.n1696 9.3005
R12892 gnd.n4971 gnd.n1697 9.3005
R12893 gnd.n4970 gnd.n1698 9.3005
R12894 gnd.n4087 gnd.n1699 9.3005
R12895 gnd.n4089 gnd.n4088 9.3005
R12896 gnd.n2383 gnd.n2382 9.3005
R12897 gnd.n4102 gnd.n4101 9.3005
R12898 gnd.n4103 gnd.n2381 9.3005
R12899 gnd.n4105 gnd.n4104 9.3005
R12900 gnd.n2369 gnd.n2368 9.3005
R12901 gnd.n4118 gnd.n4117 9.3005
R12902 gnd.n4119 gnd.n2367 9.3005
R12903 gnd.n4121 gnd.n4120 9.3005
R12904 gnd.n2357 gnd.n2356 9.3005
R12905 gnd.n4134 gnd.n4133 9.3005
R12906 gnd.n4135 gnd.n2355 9.3005
R12907 gnd.n4137 gnd.n4136 9.3005
R12908 gnd.n2343 gnd.n2342 9.3005
R12909 gnd.n4150 gnd.n4149 9.3005
R12910 gnd.n4151 gnd.n2341 9.3005
R12911 gnd.n4153 gnd.n4152 9.3005
R12912 gnd.n2328 gnd.n2327 9.3005
R12913 gnd.n4166 gnd.n4165 9.3005
R12914 gnd.n4167 gnd.n2326 9.3005
R12915 gnd.n4169 gnd.n4168 9.3005
R12916 gnd.n2314 gnd.n2313 9.3005
R12917 gnd.n4182 gnd.n4181 9.3005
R12918 gnd.n4183 gnd.n2312 9.3005
R12919 gnd.n4185 gnd.n4184 9.3005
R12920 gnd.n2300 gnd.n2299 9.3005
R12921 gnd.n4198 gnd.n4197 9.3005
R12922 gnd.n4199 gnd.n2298 9.3005
R12923 gnd.n4201 gnd.n4200 9.3005
R12924 gnd.n2287 gnd.n2286 9.3005
R12925 gnd.n4214 gnd.n4213 9.3005
R12926 gnd.n4215 gnd.n2285 9.3005
R12927 gnd.n4217 gnd.n4216 9.3005
R12928 gnd.n2273 gnd.n2272 9.3005
R12929 gnd.n4230 gnd.n4229 9.3005
R12930 gnd.n4231 gnd.n2271 9.3005
R12931 gnd.n4233 gnd.n4232 9.3005
R12932 gnd.n2259 gnd.n2258 9.3005
R12933 gnd.n4246 gnd.n4245 9.3005
R12934 gnd.n4247 gnd.n2257 9.3005
R12935 gnd.n4249 gnd.n4248 9.3005
R12936 gnd.n2246 gnd.n2245 9.3005
R12937 gnd.n4262 gnd.n4261 9.3005
R12938 gnd.n4263 gnd.n2244 9.3005
R12939 gnd.n4265 gnd.n4264 9.3005
R12940 gnd.n2232 gnd.n2231 9.3005
R12941 gnd.n4278 gnd.n4277 9.3005
R12942 gnd.n4279 gnd.n2230 9.3005
R12943 gnd.n4281 gnd.n4280 9.3005
R12944 gnd.n2219 gnd.n2218 9.3005
R12945 gnd.n4294 gnd.n4293 9.3005
R12946 gnd.n4295 gnd.n2217 9.3005
R12947 gnd.n4297 gnd.n4296 9.3005
R12948 gnd.n2204 gnd.n2203 9.3005
R12949 gnd.n4310 gnd.n4309 9.3005
R12950 gnd.n4311 gnd.n2202 9.3005
R12951 gnd.n4313 gnd.n4312 9.3005
R12952 gnd.n2191 gnd.n2190 9.3005
R12953 gnd.n4326 gnd.n4325 9.3005
R12954 gnd.n4327 gnd.n2189 9.3005
R12955 gnd.n4329 gnd.n4328 9.3005
R12956 gnd.n2180 gnd.n2179 9.3005
R12957 gnd.n4342 gnd.n4341 9.3005
R12958 gnd.n4343 gnd.n2178 9.3005
R12959 gnd.n4345 gnd.n4344 9.3005
R12960 gnd.n2167 gnd.n2166 9.3005
R12961 gnd.n4358 gnd.n4357 9.3005
R12962 gnd.n4359 gnd.n2165 9.3005
R12963 gnd.n4361 gnd.n4360 9.3005
R12964 gnd.n2152 gnd.n2151 9.3005
R12965 gnd.n4374 gnd.n4373 9.3005
R12966 gnd.n4375 gnd.n2150 9.3005
R12967 gnd.n4377 gnd.n4376 9.3005
R12968 gnd.n2140 gnd.n2139 9.3005
R12969 gnd.n4392 gnd.n4391 9.3005
R12970 gnd.n4393 gnd.n2138 9.3005
R12971 gnd.n4398 gnd.n4394 9.3005
R12972 gnd.n4397 gnd.n4396 9.3005
R12973 gnd.n4395 gnd.n1814 9.3005
R12974 gnd.n4842 gnd.n1815 9.3005
R12975 gnd.n4841 gnd.n1816 9.3005
R12976 gnd.n4840 gnd.n1817 9.3005
R12977 gnd.n2074 gnd.n1818 9.3005
R12978 gnd.n2076 gnd.n2075 9.3005
R12979 gnd.n2080 gnd.n2079 9.3005
R12980 gnd.n2081 gnd.n2073 9.3005
R12981 gnd.n2083 gnd.n2082 9.3005
R12982 gnd.n2071 gnd.n2070 9.3005
R12983 gnd.n2088 gnd.n2087 9.3005
R12984 gnd.n2089 gnd.n2069 9.3005
R12985 gnd.n2091 gnd.n2090 9.3005
R12986 gnd.n2067 gnd.n2066 9.3005
R12987 gnd.n2096 gnd.n2095 9.3005
R12988 gnd.n2097 gnd.n2065 9.3005
R12989 gnd.n2118 gnd.n2098 9.3005
R12990 gnd.n2117 gnd.n2099 9.3005
R12991 gnd.n2116 gnd.n2100 9.3005
R12992 gnd.n2103 gnd.n2101 9.3005
R12993 gnd.n2112 gnd.n2104 9.3005
R12994 gnd.n2111 gnd.n2105 9.3005
R12995 gnd.n2110 gnd.n2106 9.3005
R12996 gnd.n2108 gnd.n2107 9.3005
R12997 gnd.n2049 gnd.n2048 9.3005
R12998 gnd.n4645 gnd.n4644 9.3005
R12999 gnd.n4646 gnd.n2047 9.3005
R13000 gnd.n4649 gnd.n4648 9.3005
R13001 gnd.n4647 gnd.n553 9.3005
R13002 gnd.n7741 gnd.n554 9.3005
R13003 gnd.n7740 gnd.n555 9.3005
R13004 gnd.n7739 gnd.n556 9.3005
R13005 gnd.n559 gnd.n557 9.3005
R13006 gnd.n7735 gnd.n560 9.3005
R13007 gnd.n3022 gnd.n3021 9.3005
R13008 gnd.n2960 gnd.n2898 9.3005
R13009 gnd.n2963 gnd.n2962 9.3005
R13010 gnd.n2964 gnd.n2897 9.3005
R13011 gnd.n2967 gnd.n2965 9.3005
R13012 gnd.n2968 gnd.n2896 9.3005
R13013 gnd.n2971 gnd.n2970 9.3005
R13014 gnd.n2972 gnd.n2895 9.3005
R13015 gnd.n2975 gnd.n2973 9.3005
R13016 gnd.n2976 gnd.n2894 9.3005
R13017 gnd.n2979 gnd.n2978 9.3005
R13018 gnd.n2980 gnd.n2893 9.3005
R13019 gnd.n2983 gnd.n2981 9.3005
R13020 gnd.n2984 gnd.n2892 9.3005
R13021 gnd.n2987 gnd.n2986 9.3005
R13022 gnd.n2988 gnd.n2891 9.3005
R13023 gnd.n2991 gnd.n2989 9.3005
R13024 gnd.n2992 gnd.n2890 9.3005
R13025 gnd.n2995 gnd.n2994 9.3005
R13026 gnd.n2996 gnd.n2889 9.3005
R13027 gnd.n2999 gnd.n2997 9.3005
R13028 gnd.n3000 gnd.n2888 9.3005
R13029 gnd.n3003 gnd.n3002 9.3005
R13030 gnd.n3004 gnd.n2887 9.3005
R13031 gnd.n3007 gnd.n3005 9.3005
R13032 gnd.n3008 gnd.n2886 9.3005
R13033 gnd.n3011 gnd.n3010 9.3005
R13034 gnd.n3012 gnd.n2885 9.3005
R13035 gnd.n3015 gnd.n3013 9.3005
R13036 gnd.n3016 gnd.n2884 9.3005
R13037 gnd.n3019 gnd.n3018 9.3005
R13038 gnd.n3020 gnd.n2883 9.3005
R13039 gnd.n2959 gnd.n2957 9.3005
R13040 gnd.n2953 gnd.n2952 9.3005
R13041 gnd.n2951 gnd.n2903 9.3005
R13042 gnd.n2950 gnd.n2949 9.3005
R13043 gnd.n2946 gnd.n2906 9.3005
R13044 gnd.n2945 gnd.n2942 9.3005
R13045 gnd.n2941 gnd.n2907 9.3005
R13046 gnd.n2940 gnd.n2939 9.3005
R13047 gnd.n2936 gnd.n2908 9.3005
R13048 gnd.n2935 gnd.n2932 9.3005
R13049 gnd.n2931 gnd.n2909 9.3005
R13050 gnd.n2930 gnd.n2929 9.3005
R13051 gnd.n2926 gnd.n2910 9.3005
R13052 gnd.n2925 gnd.n2922 9.3005
R13053 gnd.n2921 gnd.n2911 9.3005
R13054 gnd.n2920 gnd.n2919 9.3005
R13055 gnd.n2916 gnd.n2912 9.3005
R13056 gnd.n2915 gnd.n1254 9.3005
R13057 gnd.n2954 gnd.n2899 9.3005
R13058 gnd.n2956 gnd.n2955 9.3005
R13059 gnd.n5050 gnd.n1622 9.3005
R13060 gnd.n5053 gnd.n1621 9.3005
R13061 gnd.n5054 gnd.n1620 9.3005
R13062 gnd.n5057 gnd.n1619 9.3005
R13063 gnd.n5058 gnd.n1618 9.3005
R13064 gnd.n5061 gnd.n1617 9.3005
R13065 gnd.n5062 gnd.n1616 9.3005
R13066 gnd.n5065 gnd.n1615 9.3005
R13067 gnd.n5067 gnd.n1612 9.3005
R13068 gnd.n5070 gnd.n1611 9.3005
R13069 gnd.n5071 gnd.n1610 9.3005
R13070 gnd.n5074 gnd.n1609 9.3005
R13071 gnd.n5075 gnd.n1608 9.3005
R13072 gnd.n5078 gnd.n1607 9.3005
R13073 gnd.n5079 gnd.n1606 9.3005
R13074 gnd.n5082 gnd.n1605 9.3005
R13075 gnd.n5083 gnd.n1604 9.3005
R13076 gnd.n5086 gnd.n1603 9.3005
R13077 gnd.n5087 gnd.n1602 9.3005
R13078 gnd.n5090 gnd.n1601 9.3005
R13079 gnd.n5091 gnd.n1600 9.3005
R13080 gnd.n5094 gnd.n1599 9.3005
R13081 gnd.n5095 gnd.n1598 9.3005
R13082 gnd.n5096 gnd.n1597 9.3005
R13083 gnd.n1554 gnd.n1553 9.3005
R13084 gnd.n5102 gnd.n5101 9.3005
R13085 gnd.n2664 gnd.n2661 9.3005
R13086 gnd.n2668 gnd.n2667 9.3005
R13087 gnd.n2669 gnd.n2659 9.3005
R13088 gnd.n2671 gnd.n2670 9.3005
R13089 gnd.n2674 gnd.n2658 9.3005
R13090 gnd.n2678 gnd.n2677 9.3005
R13091 gnd.n2679 gnd.n2657 9.3005
R13092 gnd.n2682 gnd.n2680 9.3005
R13093 gnd.n2683 gnd.n2653 9.3005
R13094 gnd.n2687 gnd.n2686 9.3005
R13095 gnd.n2688 gnd.n2652 9.3005
R13096 gnd.n2690 gnd.n2689 9.3005
R13097 gnd.n2693 gnd.n2651 9.3005
R13098 gnd.n2697 gnd.n2696 9.3005
R13099 gnd.n2698 gnd.n2650 9.3005
R13100 gnd.n2700 gnd.n2699 9.3005
R13101 gnd.n2703 gnd.n2649 9.3005
R13102 gnd.n2707 gnd.n2706 9.3005
R13103 gnd.n2708 gnd.n2648 9.3005
R13104 gnd.n2710 gnd.n2709 9.3005
R13105 gnd.n2713 gnd.n2647 9.3005
R13106 gnd.n2717 gnd.n2716 9.3005
R13107 gnd.n2718 gnd.n2646 9.3005
R13108 gnd.n2720 gnd.n2719 9.3005
R13109 gnd.n2723 gnd.n2645 9.3005
R13110 gnd.n2727 gnd.n2726 9.3005
R13111 gnd.n2728 gnd.n2644 9.3005
R13112 gnd.n2731 gnd.n2729 9.3005
R13113 gnd.n2732 gnd.n2640 9.3005
R13114 gnd.n2735 gnd.n2734 9.3005
R13115 gnd.n2660 gnd.n1623 9.3005
R13116 gnd.n1276 gnd.n1256 9.3005
R13117 gnd.n2825 gnd.n1277 9.3005
R13118 gnd.n5268 gnd.n1278 9.3005
R13119 gnd.n5267 gnd.n1279 9.3005
R13120 gnd.n5266 gnd.n1280 9.3005
R13121 gnd.n2831 gnd.n1281 9.3005
R13122 gnd.n5256 gnd.n1297 9.3005
R13123 gnd.n5255 gnd.n1298 9.3005
R13124 gnd.n5254 gnd.n1299 9.3005
R13125 gnd.n2838 gnd.n1300 9.3005
R13126 gnd.n5244 gnd.n1316 9.3005
R13127 gnd.n5243 gnd.n1317 9.3005
R13128 gnd.n5242 gnd.n1318 9.3005
R13129 gnd.n2845 gnd.n1319 9.3005
R13130 gnd.n5232 gnd.n1335 9.3005
R13131 gnd.n5231 gnd.n1336 9.3005
R13132 gnd.n5230 gnd.n1337 9.3005
R13133 gnd.n2852 gnd.n1338 9.3005
R13134 gnd.n5220 gnd.n1354 9.3005
R13135 gnd.n5219 gnd.n1355 9.3005
R13136 gnd.n5218 gnd.n1356 9.3005
R13137 gnd.n2859 gnd.n1357 9.3005
R13138 gnd.n5208 gnd.n1373 9.3005
R13139 gnd.n5207 gnd.n1374 9.3005
R13140 gnd.n5206 gnd.n1375 9.3005
R13141 gnd.n2866 gnd.n1376 9.3005
R13142 gnd.n5196 gnd.n1391 9.3005
R13143 gnd.n5195 gnd.n1392 9.3005
R13144 gnd.n5194 gnd.n1393 9.3005
R13145 gnd.n2875 gnd.n1394 9.3005
R13146 gnd.n2877 gnd.n2876 9.3005
R13147 gnd.n2806 gnd.n2801 9.3005
R13148 gnd.n3038 gnd.n2802 9.3005
R13149 gnd.n3037 gnd.n2803 9.3005
R13150 gnd.n3036 gnd.n3034 9.3005
R13151 gnd.n2804 gnd.n1418 9.3005
R13152 gnd.n5183 gnd.n1419 9.3005
R13153 gnd.n5182 gnd.n1420 9.3005
R13154 gnd.n5181 gnd.n1421 9.3005
R13155 gnd.n2773 gnd.n1422 9.3005
R13156 gnd.n5171 gnd.n1438 9.3005
R13157 gnd.n5170 gnd.n1439 9.3005
R13158 gnd.n5169 gnd.n1440 9.3005
R13159 gnd.n2768 gnd.n1441 9.3005
R13160 gnd.n5159 gnd.n1459 9.3005
R13161 gnd.n5158 gnd.n1460 9.3005
R13162 gnd.n5157 gnd.n1461 9.3005
R13163 gnd.n3113 gnd.n1462 9.3005
R13164 gnd.n5147 gnd.n1479 9.3005
R13165 gnd.n5146 gnd.n1480 9.3005
R13166 gnd.n5145 gnd.n1481 9.3005
R13167 gnd.n3122 gnd.n1482 9.3005
R13168 gnd.n5135 gnd.n1500 9.3005
R13169 gnd.n5134 gnd.n1501 9.3005
R13170 gnd.n5133 gnd.n1502 9.3005
R13171 gnd.n3190 gnd.n1503 9.3005
R13172 gnd.n5123 gnd.n1520 9.3005
R13173 gnd.n5122 gnd.n1521 9.3005
R13174 gnd.n5121 gnd.n1522 9.3005
R13175 gnd.n3205 gnd.n1523 9.3005
R13176 gnd.n5111 gnd.n1541 9.3005
R13177 gnd.n5110 gnd.n1542 9.3005
R13178 gnd.n5109 gnd.n1543 9.3005
R13179 gnd.n3223 gnd.n1544 9.3005
R13180 gnd.n5280 gnd.n1255 9.3005
R13181 gnd.n1257 gnd.n1256 9.3005
R13182 gnd.n2826 gnd.n2825 9.3005
R13183 gnd.n2827 gnd.n1278 9.3005
R13184 gnd.n2829 gnd.n1279 9.3005
R13185 gnd.n2830 gnd.n1280 9.3005
R13186 gnd.n2833 gnd.n2831 9.3005
R13187 gnd.n2834 gnd.n1297 9.3005
R13188 gnd.n2836 gnd.n1298 9.3005
R13189 gnd.n2837 gnd.n1299 9.3005
R13190 gnd.n2840 gnd.n2838 9.3005
R13191 gnd.n2841 gnd.n1316 9.3005
R13192 gnd.n2843 gnd.n1317 9.3005
R13193 gnd.n2844 gnd.n1318 9.3005
R13194 gnd.n2847 gnd.n2845 9.3005
R13195 gnd.n2848 gnd.n1335 9.3005
R13196 gnd.n2850 gnd.n1336 9.3005
R13197 gnd.n2851 gnd.n1337 9.3005
R13198 gnd.n2854 gnd.n2852 9.3005
R13199 gnd.n2855 gnd.n1354 9.3005
R13200 gnd.n2857 gnd.n1355 9.3005
R13201 gnd.n2858 gnd.n1356 9.3005
R13202 gnd.n2861 gnd.n2859 9.3005
R13203 gnd.n2862 gnd.n1373 9.3005
R13204 gnd.n2864 gnd.n1374 9.3005
R13205 gnd.n2865 gnd.n1375 9.3005
R13206 gnd.n2868 gnd.n2866 9.3005
R13207 gnd.n2869 gnd.n1391 9.3005
R13208 gnd.n2871 gnd.n1392 9.3005
R13209 gnd.n2872 gnd.n1393 9.3005
R13210 gnd.n2875 gnd.n2874 9.3005
R13211 gnd.n2876 gnd.n2805 9.3005
R13212 gnd.n3026 gnd.n2806 9.3005
R13213 gnd.n3027 gnd.n2802 9.3005
R13214 gnd.n3028 gnd.n2803 9.3005
R13215 gnd.n3034 gnd.n3033 9.3005
R13216 gnd.n3031 gnd.n2804 9.3005
R13217 gnd.n3030 gnd.n1419 9.3005
R13218 gnd.n3029 gnd.n1420 9.3005
R13219 gnd.n2772 gnd.n1421 9.3005
R13220 gnd.n3095 gnd.n2773 9.3005
R13221 gnd.n3096 gnd.n1438 9.3005
R13222 gnd.n3097 gnd.n1439 9.3005
R13223 gnd.n2767 gnd.n1440 9.3005
R13224 gnd.n3109 gnd.n2768 9.3005
R13225 gnd.n3110 gnd.n1459 9.3005
R13226 gnd.n3111 gnd.n1460 9.3005
R13227 gnd.n3112 gnd.n1461 9.3005
R13228 gnd.n3116 gnd.n3113 9.3005
R13229 gnd.n3117 gnd.n1479 9.3005
R13230 gnd.n3120 gnd.n1480 9.3005
R13231 gnd.n3121 gnd.n1481 9.3005
R13232 gnd.n3123 gnd.n3122 9.3005
R13233 gnd.n2745 gnd.n1500 9.3005
R13234 gnd.n3188 gnd.n1501 9.3005
R13235 gnd.n3189 gnd.n1502 9.3005
R13236 gnd.n3191 gnd.n3190 9.3005
R13237 gnd.n2741 gnd.n1520 9.3005
R13238 gnd.n3203 gnd.n1521 9.3005
R13239 gnd.n3204 gnd.n1522 9.3005
R13240 gnd.n3206 gnd.n3205 9.3005
R13241 gnd.n2736 gnd.n1541 9.3005
R13242 gnd.n3220 gnd.n1542 9.3005
R13243 gnd.n3221 gnd.n1543 9.3005
R13244 gnd.n3223 gnd.n3222 9.3005
R13245 gnd.n5280 gnd.n5279 9.3005
R13246 gnd.n5284 gnd.n5283 9.3005
R13247 gnd.n5287 gnd.n1250 9.3005
R13248 gnd.n5288 gnd.n1249 9.3005
R13249 gnd.n5291 gnd.n1248 9.3005
R13250 gnd.n5292 gnd.n1247 9.3005
R13251 gnd.n5295 gnd.n1246 9.3005
R13252 gnd.n5296 gnd.n1245 9.3005
R13253 gnd.n5299 gnd.n1244 9.3005
R13254 gnd.n5300 gnd.n1243 9.3005
R13255 gnd.n5303 gnd.n1242 9.3005
R13256 gnd.n5304 gnd.n1241 9.3005
R13257 gnd.n5307 gnd.n1240 9.3005
R13258 gnd.n5308 gnd.n1239 9.3005
R13259 gnd.n5311 gnd.n1238 9.3005
R13260 gnd.n5312 gnd.n1237 9.3005
R13261 gnd.n5315 gnd.n1236 9.3005
R13262 gnd.n5316 gnd.n1235 9.3005
R13263 gnd.n5319 gnd.n1234 9.3005
R13264 gnd.n5320 gnd.n1233 9.3005
R13265 gnd.n5323 gnd.n1232 9.3005
R13266 gnd.n5327 gnd.n1228 9.3005
R13267 gnd.n5328 gnd.n1227 9.3005
R13268 gnd.n5331 gnd.n1226 9.3005
R13269 gnd.n5332 gnd.n1225 9.3005
R13270 gnd.n5335 gnd.n1224 9.3005
R13271 gnd.n5336 gnd.n1223 9.3005
R13272 gnd.n5339 gnd.n1222 9.3005
R13273 gnd.n5340 gnd.n1221 9.3005
R13274 gnd.n5343 gnd.n1220 9.3005
R13275 gnd.n5344 gnd.n1219 9.3005
R13276 gnd.n5347 gnd.n1218 9.3005
R13277 gnd.n5348 gnd.n1217 9.3005
R13278 gnd.n5351 gnd.n1216 9.3005
R13279 gnd.n5352 gnd.n1215 9.3005
R13280 gnd.n5355 gnd.n1214 9.3005
R13281 gnd.n5356 gnd.n1213 9.3005
R13282 gnd.n5359 gnd.n1212 9.3005
R13283 gnd.n5360 gnd.n1211 9.3005
R13284 gnd.n5363 gnd.n1210 9.3005
R13285 gnd.n5365 gnd.n1207 9.3005
R13286 gnd.n5368 gnd.n1206 9.3005
R13287 gnd.n5369 gnd.n1205 9.3005
R13288 gnd.n5372 gnd.n1204 9.3005
R13289 gnd.n5373 gnd.n1203 9.3005
R13290 gnd.n5376 gnd.n1202 9.3005
R13291 gnd.n5377 gnd.n1201 9.3005
R13292 gnd.n5380 gnd.n1200 9.3005
R13293 gnd.n5381 gnd.n1199 9.3005
R13294 gnd.n5384 gnd.n1198 9.3005
R13295 gnd.n5385 gnd.n1197 9.3005
R13296 gnd.n5388 gnd.n1196 9.3005
R13297 gnd.n5389 gnd.n1195 9.3005
R13298 gnd.n5392 gnd.n1194 9.3005
R13299 gnd.n5394 gnd.n1193 9.3005
R13300 gnd.n5395 gnd.n1192 9.3005
R13301 gnd.n5396 gnd.n1191 9.3005
R13302 gnd.n5397 gnd.n1190 9.3005
R13303 gnd.n5324 gnd.n1229 9.3005
R13304 gnd.n5282 gnd.n1251 9.3005
R13305 gnd.n5274 gnd.n1265 9.3005
R13306 gnd.n5273 gnd.n1266 9.3005
R13307 gnd.n5272 gnd.n1267 9.3005
R13308 gnd.n1287 gnd.n1268 9.3005
R13309 gnd.n5262 gnd.n1288 9.3005
R13310 gnd.n5261 gnd.n1289 9.3005
R13311 gnd.n5260 gnd.n1290 9.3005
R13312 gnd.n1305 gnd.n1291 9.3005
R13313 gnd.n5250 gnd.n1306 9.3005
R13314 gnd.n5249 gnd.n1307 9.3005
R13315 gnd.n5248 gnd.n1308 9.3005
R13316 gnd.n1325 gnd.n1309 9.3005
R13317 gnd.n5238 gnd.n1326 9.3005
R13318 gnd.n5237 gnd.n1327 9.3005
R13319 gnd.n5236 gnd.n1328 9.3005
R13320 gnd.n1343 gnd.n1329 9.3005
R13321 gnd.n5226 gnd.n1344 9.3005
R13322 gnd.n5225 gnd.n1345 9.3005
R13323 gnd.n5224 gnd.n1346 9.3005
R13324 gnd.n1363 gnd.n1347 9.3005
R13325 gnd.n5214 gnd.n1364 9.3005
R13326 gnd.n5213 gnd.n1365 9.3005
R13327 gnd.n5212 gnd.n1366 9.3005
R13328 gnd.n1381 gnd.n1367 9.3005
R13329 gnd.n5202 gnd.n1382 9.3005
R13330 gnd.n5201 gnd.n1383 9.3005
R13331 gnd.n1409 gnd.n1403 9.3005
R13332 gnd.n5177 gnd.n1428 9.3005
R13333 gnd.n5176 gnd.n1429 9.3005
R13334 gnd.n5175 gnd.n1430 9.3005
R13335 gnd.n1448 gnd.n1431 9.3005
R13336 gnd.n5165 gnd.n1449 9.3005
R13337 gnd.n5164 gnd.n1450 9.3005
R13338 gnd.n5163 gnd.n1451 9.3005
R13339 gnd.n1468 gnd.n1452 9.3005
R13340 gnd.n5153 gnd.n1469 9.3005
R13341 gnd.n5152 gnd.n1470 9.3005
R13342 gnd.n5151 gnd.n1471 9.3005
R13343 gnd.n1489 gnd.n1472 9.3005
R13344 gnd.n5141 gnd.n1490 9.3005
R13345 gnd.n5140 gnd.n1491 9.3005
R13346 gnd.n5139 gnd.n1492 9.3005
R13347 gnd.n1509 gnd.n1493 9.3005
R13348 gnd.n5129 gnd.n1510 9.3005
R13349 gnd.n5128 gnd.n1511 9.3005
R13350 gnd.n5127 gnd.n1512 9.3005
R13351 gnd.n1530 gnd.n1513 9.3005
R13352 gnd.n5117 gnd.n1531 9.3005
R13353 gnd.n5116 gnd.n1532 9.3005
R13354 gnd.n5115 gnd.n1533 9.3005
R13355 gnd.n1551 gnd.n1534 9.3005
R13356 gnd.n5105 gnd.n1552 9.3005
R13357 gnd.n5104 gnd.n5103 9.3005
R13358 gnd.n1264 gnd.n1263 9.3005
R13359 gnd.n5188 gnd.n5187 9.3005
R13360 gnd.n2821 gnd.n2812 9.3005
R13361 gnd.n2820 gnd.n2813 9.3005
R13362 gnd.n2817 gnd.n2814 9.3005
R13363 gnd.n2816 gnd.n2815 9.3005
R13364 gnd.n2782 gnd.n2781 9.3005
R13365 gnd.n3059 gnd.n3058 9.3005
R13366 gnd.n2822 gnd.n2811 9.3005
R13367 gnd.n6886 gnd.n1133 9.3005
R13368 gnd.n6887 gnd.n1132 9.3005
R13369 gnd.n6888 gnd.n1131 9.3005
R13370 gnd.n1130 gnd.n1126 9.3005
R13371 gnd.n6894 gnd.n1125 9.3005
R13372 gnd.n6895 gnd.n1124 9.3005
R13373 gnd.n6896 gnd.n1123 9.3005
R13374 gnd.n1122 gnd.n1118 9.3005
R13375 gnd.n6902 gnd.n1117 9.3005
R13376 gnd.n6903 gnd.n1116 9.3005
R13377 gnd.n6904 gnd.n1115 9.3005
R13378 gnd.n1114 gnd.n1110 9.3005
R13379 gnd.n6910 gnd.n1109 9.3005
R13380 gnd.n6911 gnd.n1108 9.3005
R13381 gnd.n6912 gnd.n1107 9.3005
R13382 gnd.n1106 gnd.n1102 9.3005
R13383 gnd.n6918 gnd.n1101 9.3005
R13384 gnd.n6919 gnd.n1100 9.3005
R13385 gnd.n6920 gnd.n1099 9.3005
R13386 gnd.n1098 gnd.n1094 9.3005
R13387 gnd.n6926 gnd.n1093 9.3005
R13388 gnd.n6927 gnd.n1092 9.3005
R13389 gnd.n6928 gnd.n1091 9.3005
R13390 gnd.n1090 gnd.n1086 9.3005
R13391 gnd.n6934 gnd.n1085 9.3005
R13392 gnd.n6935 gnd.n1084 9.3005
R13393 gnd.n6936 gnd.n1083 9.3005
R13394 gnd.n1082 gnd.n1078 9.3005
R13395 gnd.n6942 gnd.n1077 9.3005
R13396 gnd.n6943 gnd.n1076 9.3005
R13397 gnd.n6944 gnd.n1075 9.3005
R13398 gnd.n1074 gnd.n1070 9.3005
R13399 gnd.n6950 gnd.n1069 9.3005
R13400 gnd.n6951 gnd.n1068 9.3005
R13401 gnd.n6952 gnd.n1067 9.3005
R13402 gnd.n1066 gnd.n1062 9.3005
R13403 gnd.n6958 gnd.n1061 9.3005
R13404 gnd.n6959 gnd.n1060 9.3005
R13405 gnd.n6960 gnd.n1059 9.3005
R13406 gnd.n1058 gnd.n1054 9.3005
R13407 gnd.n6966 gnd.n1053 9.3005
R13408 gnd.n6967 gnd.n1052 9.3005
R13409 gnd.n6968 gnd.n1051 9.3005
R13410 gnd.n1050 gnd.n1046 9.3005
R13411 gnd.n6974 gnd.n1045 9.3005
R13412 gnd.n6975 gnd.n1044 9.3005
R13413 gnd.n6976 gnd.n1043 9.3005
R13414 gnd.n1042 gnd.n1038 9.3005
R13415 gnd.n6982 gnd.n1037 9.3005
R13416 gnd.n6983 gnd.n1036 9.3005
R13417 gnd.n6984 gnd.n1035 9.3005
R13418 gnd.n1034 gnd.n1030 9.3005
R13419 gnd.n6990 gnd.n1029 9.3005
R13420 gnd.n6991 gnd.n1028 9.3005
R13421 gnd.n6992 gnd.n1027 9.3005
R13422 gnd.n1026 gnd.n1022 9.3005
R13423 gnd.n6998 gnd.n1021 9.3005
R13424 gnd.n6999 gnd.n1020 9.3005
R13425 gnd.n7000 gnd.n1019 9.3005
R13426 gnd.n1018 gnd.n1014 9.3005
R13427 gnd.n7006 gnd.n1013 9.3005
R13428 gnd.n7007 gnd.n1012 9.3005
R13429 gnd.n7008 gnd.n1011 9.3005
R13430 gnd.n1010 gnd.n1006 9.3005
R13431 gnd.n7014 gnd.n1005 9.3005
R13432 gnd.n7015 gnd.n1004 9.3005
R13433 gnd.n7016 gnd.n1003 9.3005
R13434 gnd.n1002 gnd.n998 9.3005
R13435 gnd.n7022 gnd.n997 9.3005
R13436 gnd.n7023 gnd.n996 9.3005
R13437 gnd.n7024 gnd.n995 9.3005
R13438 gnd.n994 gnd.n990 9.3005
R13439 gnd.n7030 gnd.n989 9.3005
R13440 gnd.n7031 gnd.n988 9.3005
R13441 gnd.n7032 gnd.n987 9.3005
R13442 gnd.n986 gnd.n982 9.3005
R13443 gnd.n7038 gnd.n981 9.3005
R13444 gnd.n7039 gnd.n980 9.3005
R13445 gnd.n7040 gnd.n979 9.3005
R13446 gnd.n978 gnd.n974 9.3005
R13447 gnd.n7046 gnd.n973 9.3005
R13448 gnd.n7047 gnd.n972 9.3005
R13449 gnd.n7048 gnd.n971 9.3005
R13450 gnd.n970 gnd.n966 9.3005
R13451 gnd.n2810 gnd.n1134 9.3005
R13452 gnd.n4563 gnd.n4406 9.3005
R13453 gnd.n2534 gnd.n2533 9.3005
R13454 gnd.n3384 gnd.n3383 9.3005
R13455 gnd.n3385 gnd.n2532 9.3005
R13456 gnd.n3387 gnd.n3386 9.3005
R13457 gnd.n2520 gnd.n2519 9.3005
R13458 gnd.n3400 gnd.n3399 9.3005
R13459 gnd.n3401 gnd.n2518 9.3005
R13460 gnd.n3403 gnd.n3402 9.3005
R13461 gnd.n2505 gnd.n2504 9.3005
R13462 gnd.n3416 gnd.n3415 9.3005
R13463 gnd.n3417 gnd.n2503 9.3005
R13464 gnd.n3419 gnd.n3418 9.3005
R13465 gnd.n2490 gnd.n2489 9.3005
R13466 gnd.n3441 gnd.n3440 9.3005
R13467 gnd.n3442 gnd.n2488 9.3005
R13468 gnd.n3444 gnd.n3443 9.3005
R13469 gnd.n2486 gnd.n2485 9.3005
R13470 gnd.n3449 gnd.n3448 9.3005
R13471 gnd.n3450 gnd.n2483 9.3005
R13472 gnd.n3453 gnd.n3452 9.3005
R13473 gnd.n3451 gnd.n2484 9.3005
R13474 gnd.n2389 gnd.n2388 9.3005
R13475 gnd.n4094 gnd.n4093 9.3005
R13476 gnd.n4095 gnd.n2387 9.3005
R13477 gnd.n4097 gnd.n4096 9.3005
R13478 gnd.n2376 gnd.n2375 9.3005
R13479 gnd.n4110 gnd.n4109 9.3005
R13480 gnd.n4111 gnd.n2374 9.3005
R13481 gnd.n4113 gnd.n4112 9.3005
R13482 gnd.n2363 gnd.n2362 9.3005
R13483 gnd.n4126 gnd.n4125 9.3005
R13484 gnd.n4127 gnd.n2361 9.3005
R13485 gnd.n4129 gnd.n4128 9.3005
R13486 gnd.n2350 gnd.n2349 9.3005
R13487 gnd.n4142 gnd.n4141 9.3005
R13488 gnd.n4143 gnd.n2348 9.3005
R13489 gnd.n4145 gnd.n4144 9.3005
R13490 gnd.n2337 gnd.n2336 9.3005
R13491 gnd.n4158 gnd.n4157 9.3005
R13492 gnd.n4159 gnd.n2335 9.3005
R13493 gnd.n4161 gnd.n4160 9.3005
R13494 gnd.n2321 gnd.n2320 9.3005
R13495 gnd.n4174 gnd.n4173 9.3005
R13496 gnd.n4175 gnd.n2319 9.3005
R13497 gnd.n4177 gnd.n4176 9.3005
R13498 gnd.n2307 gnd.n2306 9.3005
R13499 gnd.n4190 gnd.n4189 9.3005
R13500 gnd.n4191 gnd.n2305 9.3005
R13501 gnd.n4193 gnd.n4192 9.3005
R13502 gnd.n2293 gnd.n2292 9.3005
R13503 gnd.n4206 gnd.n4205 9.3005
R13504 gnd.n4207 gnd.n2291 9.3005
R13505 gnd.n4209 gnd.n4208 9.3005
R13506 gnd.n2280 gnd.n2279 9.3005
R13507 gnd.n4222 gnd.n4221 9.3005
R13508 gnd.n4223 gnd.n2278 9.3005
R13509 gnd.n4225 gnd.n4224 9.3005
R13510 gnd.n2266 gnd.n2265 9.3005
R13511 gnd.n4238 gnd.n4237 9.3005
R13512 gnd.n4239 gnd.n2264 9.3005
R13513 gnd.n4241 gnd.n4240 9.3005
R13514 gnd.n2252 gnd.n2251 9.3005
R13515 gnd.n4254 gnd.n4253 9.3005
R13516 gnd.n4255 gnd.n2250 9.3005
R13517 gnd.n4257 gnd.n4256 9.3005
R13518 gnd.n2239 gnd.n2238 9.3005
R13519 gnd.n4270 gnd.n4269 9.3005
R13520 gnd.n4271 gnd.n2237 9.3005
R13521 gnd.n4273 gnd.n4272 9.3005
R13522 gnd.n2226 gnd.n2225 9.3005
R13523 gnd.n4286 gnd.n4285 9.3005
R13524 gnd.n4287 gnd.n2224 9.3005
R13525 gnd.n4289 gnd.n4288 9.3005
R13526 gnd.n2211 gnd.n2210 9.3005
R13527 gnd.n4302 gnd.n4301 9.3005
R13528 gnd.n4303 gnd.n2209 9.3005
R13529 gnd.n4305 gnd.n4304 9.3005
R13530 gnd.n2197 gnd.n2196 9.3005
R13531 gnd.n4318 gnd.n4317 9.3005
R13532 gnd.n4319 gnd.n2195 9.3005
R13533 gnd.n4321 gnd.n4320 9.3005
R13534 gnd.n2185 gnd.n2184 9.3005
R13535 gnd.n4334 gnd.n4333 9.3005
R13536 gnd.n4335 gnd.n2183 9.3005
R13537 gnd.n4337 gnd.n4336 9.3005
R13538 gnd.n2173 gnd.n2172 9.3005
R13539 gnd.n4350 gnd.n4349 9.3005
R13540 gnd.n4351 gnd.n2171 9.3005
R13541 gnd.n4353 gnd.n4352 9.3005
R13542 gnd.n2160 gnd.n2159 9.3005
R13543 gnd.n4366 gnd.n4365 9.3005
R13544 gnd.n4367 gnd.n2158 9.3005
R13545 gnd.n4369 gnd.n4368 9.3005
R13546 gnd.n2147 gnd.n2146 9.3005
R13547 gnd.n4382 gnd.n4381 9.3005
R13548 gnd.n4383 gnd.n2144 9.3005
R13549 gnd.n4387 gnd.n4386 9.3005
R13550 gnd.n4385 gnd.n2145 9.3005
R13551 gnd.n4384 gnd.n2132 9.3005
R13552 gnd.n4403 gnd.n2131 9.3005
R13553 gnd.n4405 gnd.n4404 9.3005
R13554 gnd.n3371 gnd.n3370 9.3005
R13555 gnd.n3369 gnd.n3368 9.3005
R13556 gnd.n2789 gnd.n2788 9.3005
R13557 gnd.n3049 gnd.n3048 9.3005
R13558 gnd.n3050 gnd.n2787 9.3005
R13559 gnd.n3052 gnd.n3051 9.3005
R13560 gnd.n2776 gnd.n2775 9.3005
R13561 gnd.n3088 gnd.n3087 9.3005
R13562 gnd.n3089 gnd.n2774 9.3005
R13563 gnd.n3091 gnd.n3090 9.3005
R13564 gnd.n2771 gnd.n2770 9.3005
R13565 gnd.n3102 gnd.n3101 9.3005
R13566 gnd.n3103 gnd.n2769 9.3005
R13567 gnd.n3105 gnd.n3104 9.3005
R13568 gnd.n2761 gnd.n2759 9.3005
R13569 gnd.n3140 gnd.n3139 9.3005
R13570 gnd.n3138 gnd.n2760 9.3005
R13571 gnd.n3137 gnd.n3136 9.3005
R13572 gnd.n3135 gnd.n2762 9.3005
R13573 gnd.n3134 gnd.n3133 9.3005
R13574 gnd.n3132 gnd.n2765 9.3005
R13575 gnd.n3131 gnd.n3130 9.3005
R13576 gnd.n3129 gnd.n2766 9.3005
R13577 gnd.n3128 gnd.n3127 9.3005
R13578 gnd.n2744 gnd.n2743 9.3005
R13579 gnd.n3196 gnd.n3195 9.3005
R13580 gnd.n3197 gnd.n2742 9.3005
R13581 gnd.n3199 gnd.n3198 9.3005
R13582 gnd.n2740 gnd.n2739 9.3005
R13583 gnd.n3211 gnd.n3210 9.3005
R13584 gnd.n3212 gnd.n2737 9.3005
R13585 gnd.n3216 gnd.n3215 9.3005
R13586 gnd.n3214 gnd.n2738 9.3005
R13587 gnd.n3213 gnd.n2553 9.3005
R13588 gnd.n3332 gnd.n3331 9.3005
R13589 gnd.n3330 gnd.n3329 9.3005
R13590 gnd.n3238 gnd.n3237 9.3005
R13591 gnd.n3324 gnd.n3323 9.3005
R13592 gnd.n3322 gnd.n3321 9.3005
R13593 gnd.n3248 gnd.n3247 9.3005
R13594 gnd.n3316 gnd.n3315 9.3005
R13595 gnd.n3314 gnd.n3313 9.3005
R13596 gnd.n3258 gnd.n3257 9.3005
R13597 gnd.n3308 gnd.n3307 9.3005
R13598 gnd.n3306 gnd.n3305 9.3005
R13599 gnd.n3268 gnd.n3267 9.3005
R13600 gnd.n3300 gnd.n3299 9.3005
R13601 gnd.n3298 gnd.n3297 9.3005
R13602 gnd.n3278 gnd.n3277 9.3005
R13603 gnd.n3292 gnd.n3291 9.3005
R13604 gnd.n3285 gnd.n2552 9.3005
R13605 gnd.n3365 gnd.n3364 9.3005
R13606 gnd.n3233 gnd.n3231 9.3005
R13607 gnd.n3367 gnd.n3366 9.3005
R13608 gnd.n2549 gnd.n2547 9.3005
R13609 gnd.n3288 gnd.n3287 9.3005
R13610 gnd.n3294 gnd.n3293 9.3005
R13611 gnd.n3296 gnd.n3295 9.3005
R13612 gnd.n3272 gnd.n3271 9.3005
R13613 gnd.n3302 gnd.n3301 9.3005
R13614 gnd.n3304 gnd.n3303 9.3005
R13615 gnd.n3264 gnd.n3263 9.3005
R13616 gnd.n3310 gnd.n3309 9.3005
R13617 gnd.n3312 gnd.n3311 9.3005
R13618 gnd.n3252 gnd.n3251 9.3005
R13619 gnd.n3318 gnd.n3317 9.3005
R13620 gnd.n3320 gnd.n3319 9.3005
R13621 gnd.n3244 gnd.n3243 9.3005
R13622 gnd.n3326 gnd.n3325 9.3005
R13623 gnd.n3328 gnd.n3327 9.3005
R13624 gnd.n3232 gnd.n3230 9.3005
R13625 gnd.n3334 gnd.n3333 9.3005
R13626 gnd.n3335 gnd.n3225 9.3005
R13627 gnd.n3337 gnd.n3336 9.3005
R13628 gnd.n3339 gnd.n2639 9.3005
R13629 gnd.n3341 gnd.n3340 9.3005
R13630 gnd.n3342 gnd.n2635 9.3005
R13631 gnd.n3344 gnd.n3343 9.3005
R13632 gnd.n3345 gnd.n2634 9.3005
R13633 gnd.n3347 gnd.n3346 9.3005
R13634 gnd.n3348 gnd.n2633 9.3005
R13635 gnd.n2630 gnd.n2582 9.3005
R13636 gnd.n2629 gnd.n2628 9.3005
R13637 gnd.n2627 gnd.n2585 9.3005
R13638 gnd.n2626 gnd.n2625 9.3005
R13639 gnd.n2624 gnd.n2586 9.3005
R13640 gnd.n2623 gnd.n2622 9.3005
R13641 gnd.n2621 gnd.n2589 9.3005
R13642 gnd.n2620 gnd.n2619 9.3005
R13643 gnd.n2618 gnd.n2590 9.3005
R13644 gnd.n2617 gnd.n2616 9.3005
R13645 gnd.n2615 gnd.n2593 9.3005
R13646 gnd.n2614 gnd.n2613 9.3005
R13647 gnd.n2612 gnd.n2594 9.3005
R13648 gnd.n2611 gnd.n2610 9.3005
R13649 gnd.n2609 gnd.n2596 9.3005
R13650 gnd.n2608 gnd.n2607 9.3005
R13651 gnd.n2606 gnd.n2597 9.3005
R13652 gnd.n2605 gnd.n2604 9.3005
R13653 gnd.n2603 gnd.n2602 9.3005
R13654 gnd.n1708 gnd.n1706 9.3005
R13655 gnd.n4967 gnd.n4966 9.3005
R13656 gnd.n4965 gnd.n1707 9.3005
R13657 gnd.n4964 gnd.n4963 9.3005
R13658 gnd.n4962 gnd.n1709 9.3005
R13659 gnd.n4961 gnd.n4960 9.3005
R13660 gnd.n4959 gnd.n1713 9.3005
R13661 gnd.n4958 gnd.n4957 9.3005
R13662 gnd.n4956 gnd.n1714 9.3005
R13663 gnd.n4955 gnd.n4954 9.3005
R13664 gnd.n4953 gnd.n1718 9.3005
R13665 gnd.n4952 gnd.n4951 9.3005
R13666 gnd.n4950 gnd.n1719 9.3005
R13667 gnd.n4949 gnd.n4948 9.3005
R13668 gnd.n4947 gnd.n1723 9.3005
R13669 gnd.n4946 gnd.n4945 9.3005
R13670 gnd.n4944 gnd.n1724 9.3005
R13671 gnd.n4943 gnd.n4942 9.3005
R13672 gnd.n4941 gnd.n1728 9.3005
R13673 gnd.n4940 gnd.n4939 9.3005
R13674 gnd.n4938 gnd.n1729 9.3005
R13675 gnd.n4937 gnd.n4936 9.3005
R13676 gnd.n4935 gnd.n1733 9.3005
R13677 gnd.n4934 gnd.n4933 9.3005
R13678 gnd.n4932 gnd.n1734 9.3005
R13679 gnd.n4931 gnd.n4930 9.3005
R13680 gnd.n4929 gnd.n1738 9.3005
R13681 gnd.n4928 gnd.n4927 9.3005
R13682 gnd.n4926 gnd.n1739 9.3005
R13683 gnd.n4925 gnd.n4924 9.3005
R13684 gnd.n4923 gnd.n1743 9.3005
R13685 gnd.n4922 gnd.n4921 9.3005
R13686 gnd.n4920 gnd.n1744 9.3005
R13687 gnd.n4919 gnd.n4918 9.3005
R13688 gnd.n4917 gnd.n1748 9.3005
R13689 gnd.n4916 gnd.n4915 9.3005
R13690 gnd.n4914 gnd.n1749 9.3005
R13691 gnd.n4913 gnd.n4912 9.3005
R13692 gnd.n4911 gnd.n1753 9.3005
R13693 gnd.n4910 gnd.n4909 9.3005
R13694 gnd.n4908 gnd.n1754 9.3005
R13695 gnd.n4907 gnd.n4906 9.3005
R13696 gnd.n4905 gnd.n1758 9.3005
R13697 gnd.n4904 gnd.n4903 9.3005
R13698 gnd.n4902 gnd.n1759 9.3005
R13699 gnd.n4901 gnd.n4900 9.3005
R13700 gnd.n4899 gnd.n1763 9.3005
R13701 gnd.n4898 gnd.n4897 9.3005
R13702 gnd.n4896 gnd.n1764 9.3005
R13703 gnd.n4895 gnd.n4894 9.3005
R13704 gnd.n4893 gnd.n1768 9.3005
R13705 gnd.n4892 gnd.n4891 9.3005
R13706 gnd.n4890 gnd.n1769 9.3005
R13707 gnd.n4889 gnd.n4888 9.3005
R13708 gnd.n4887 gnd.n1773 9.3005
R13709 gnd.n4886 gnd.n4885 9.3005
R13710 gnd.n4884 gnd.n1774 9.3005
R13711 gnd.n4883 gnd.n4882 9.3005
R13712 gnd.n4881 gnd.n1778 9.3005
R13713 gnd.n4880 gnd.n4879 9.3005
R13714 gnd.n4878 gnd.n1779 9.3005
R13715 gnd.n4877 gnd.n4876 9.3005
R13716 gnd.n4875 gnd.n1783 9.3005
R13717 gnd.n4874 gnd.n4873 9.3005
R13718 gnd.n4872 gnd.n1784 9.3005
R13719 gnd.n4871 gnd.n4870 9.3005
R13720 gnd.n4869 gnd.n1788 9.3005
R13721 gnd.n4868 gnd.n4867 9.3005
R13722 gnd.n4866 gnd.n1789 9.3005
R13723 gnd.n4865 gnd.n4864 9.3005
R13724 gnd.n4863 gnd.n1793 9.3005
R13725 gnd.n4862 gnd.n4861 9.3005
R13726 gnd.n4860 gnd.n1794 9.3005
R13727 gnd.n4859 gnd.n4858 9.3005
R13728 gnd.n4857 gnd.n1798 9.3005
R13729 gnd.n4856 gnd.n4855 9.3005
R13730 gnd.n4854 gnd.n1799 9.3005
R13731 gnd.n4853 gnd.n4852 9.3005
R13732 gnd.n4851 gnd.n1803 9.3005
R13733 gnd.n4850 gnd.n4849 9.3005
R13734 gnd.n4848 gnd.n1804 9.3005
R13735 gnd.n4847 gnd.n1807 9.3005
R13736 gnd.n2632 gnd.n2631 9.3005
R13737 gnd.n4455 gnd.n4454 9.3005
R13738 gnd.n4450 gnd.n4449 9.3005
R13739 gnd.n4462 gnd.n4461 9.3005
R13740 gnd.n4463 gnd.n4448 9.3005
R13741 gnd.n4466 gnd.n4465 9.3005
R13742 gnd.n4464 gnd.n4446 9.3005
R13743 gnd.n4453 gnd.n4452 9.3005
R13744 gnd.n4552 gnd.n4413 9.3005
R13745 gnd.n4549 gnd.n4548 9.3005
R13746 gnd.n4425 gnd.n4419 9.3005
R13747 gnd.n4538 gnd.n4537 9.3005
R13748 gnd.n4534 gnd.n4424 9.3005
R13749 gnd.n4531 gnd.n4530 9.3005
R13750 gnd.n4428 gnd.n4427 9.3005
R13751 gnd.n4519 gnd.n4518 9.3005
R13752 gnd.n4515 gnd.n4432 9.3005
R13753 gnd.n4512 gnd.n4511 9.3005
R13754 gnd.n4435 gnd.n4434 9.3005
R13755 gnd.n4500 gnd.n4499 9.3005
R13756 gnd.n4496 gnd.n4439 9.3005
R13757 gnd.n4493 gnd.n4492 9.3005
R13758 gnd.n4442 gnd.n4441 9.3005
R13759 gnd.n4481 gnd.n4480 9.3005
R13760 gnd.n4477 gnd.n4475 9.3005
R13761 gnd.n4554 gnd.n4553 9.3005
R13762 gnd.n4415 gnd.n4407 9.3005
R13763 gnd.n4473 gnd.n4472 9.3005
R13764 gnd.n4474 gnd.n4445 9.3005
R13765 gnd.n4483 gnd.n4482 9.3005
R13766 gnd.n4476 gnd.n4443 9.3005
R13767 gnd.n4490 gnd.n4489 9.3005
R13768 gnd.n4491 gnd.n4438 9.3005
R13769 gnd.n4502 gnd.n4501 9.3005
R13770 gnd.n4440 gnd.n4436 9.3005
R13771 gnd.n4509 gnd.n4508 9.3005
R13772 gnd.n4510 gnd.n4431 9.3005
R13773 gnd.n4521 gnd.n4520 9.3005
R13774 gnd.n4433 gnd.n4429 9.3005
R13775 gnd.n4528 gnd.n4527 9.3005
R13776 gnd.n4529 gnd.n4423 9.3005
R13777 gnd.n4540 gnd.n4539 9.3005
R13778 gnd.n4426 gnd.n4421 9.3005
R13779 gnd.n4545 gnd.n4420 9.3005
R13780 gnd.n4547 gnd.n4546 9.3005
R13781 gnd.n4556 gnd.n4555 9.3005
R13782 gnd.n4414 gnd.n4408 9.3005
R13783 gnd.n4565 gnd.n4564 9.3005
R13784 gnd.n4569 gnd.n2130 9.3005
R13785 gnd.n4571 gnd.n4570 9.3005
R13786 gnd.n2128 gnd.n2127 9.3005
R13787 gnd.n4582 gnd.n4581 9.3005
R13788 gnd.n4583 gnd.n2126 9.3005
R13789 gnd.n4585 gnd.n4584 9.3005
R13790 gnd.n2123 gnd.n2122 9.3005
R13791 gnd.n4596 gnd.n4595 9.3005
R13792 gnd.n4597 gnd.n2121 9.3005
R13793 gnd.n4599 gnd.n4598 9.3005
R13794 gnd.n2060 gnd.n2059 9.3005
R13795 gnd.n4610 gnd.n4609 9.3005
R13796 gnd.n4611 gnd.n2058 9.3005
R13797 gnd.n4613 gnd.n4612 9.3005
R13798 gnd.n2055 gnd.n2054 9.3005
R13799 gnd.n4627 gnd.n4626 9.3005
R13800 gnd.n4628 gnd.n2052 9.3005
R13801 gnd.n4638 gnd.n4637 9.3005
R13802 gnd.n4636 gnd.n2053 9.3005
R13803 gnd.n4635 gnd.n4634 9.3005
R13804 gnd.n4633 gnd.n4629 9.3005
R13805 gnd.n4632 gnd.n4631 9.3005
R13806 gnd.n530 gnd.n529 9.3005
R13807 gnd.n7771 gnd.n7770 9.3005
R13808 gnd.n7772 gnd.n528 9.3005
R13809 gnd.n7774 gnd.n7773 9.3005
R13810 gnd.n508 gnd.n507 9.3005
R13811 gnd.n7798 gnd.n7797 9.3005
R13812 gnd.n7799 gnd.n505 9.3005
R13813 gnd.n7801 gnd.n7800 9.3005
R13814 gnd.n506 gnd.n99 9.3005
R13815 gnd.n4568 gnd.n4567 9.3005
R13816 gnd.n8102 gnd.n100 9.3005
R13817 gnd.t32 gnd.n5857 9.24152
R13818 gnd.n6771 gnd.t171 9.24152
R13819 gnd.t140 gnd.n1137 9.24152
R13820 gnd.n5234 gnd.t211 9.24152
R13821 gnd.t7 gnd.n2372 9.24152
R13822 gnd.n3486 gnd.t7 9.24152
R13823 gnd.n4283 gnd.t185 9.24152
R13824 gnd.n3914 gnd.t185 9.24152
R13825 gnd.n8053 gnd.t247 9.24152
R13826 gnd.t35 gnd.t32 8.92286
R13827 gnd.n5742 gnd.n5717 8.92171
R13828 gnd.n5710 gnd.n5685 8.92171
R13829 gnd.n5678 gnd.n5653 8.92171
R13830 gnd.n5647 gnd.n5622 8.92171
R13831 gnd.n5615 gnd.n5590 8.92171
R13832 gnd.n5583 gnd.n5558 8.92171
R13833 gnd.n5551 gnd.n5526 8.92171
R13834 gnd.n5520 gnd.n5495 8.92171
R13835 gnd.n3724 gnd.n3706 8.72777
R13836 gnd.t54 gnd.n5899 8.60421
R13837 gnd.n5258 gnd.t201 8.60421
R13838 gnd.t181 gnd.n2302 8.60421
R13839 gnd.n3568 gnd.t0 8.60421
R13840 gnd.n8029 gnd.t226 8.60421
R13841 gnd.n6287 gnd.n6267 8.43656
R13842 gnd.n58 gnd.n38 8.43656
R13843 gnd.t109 gnd.n1703 8.28555
R13844 gnd.n4115 gnd.n2371 8.28555
R13845 gnd.n4034 gnd.n3517 8.28555
R13846 gnd.n4013 gnd.n4012 8.28555
R13847 gnd.n4219 gnd.n2283 8.28555
R13848 gnd.n4251 gnd.n2254 8.28555
R13849 gnd.n3639 gnd.n3638 8.28555
R13850 gnd.n3892 gnd.n3657 8.28555
R13851 gnd.n5743 gnd.n5715 8.14595
R13852 gnd.n5711 gnd.n5683 8.14595
R13853 gnd.n5679 gnd.n5651 8.14595
R13854 gnd.n5648 gnd.n5620 8.14595
R13855 gnd.n5616 gnd.n5588 8.14595
R13856 gnd.n5584 gnd.n5556 8.14595
R13857 gnd.n5552 gnd.n5524 8.14595
R13858 gnd.n5521 gnd.n5493 8.14595
R13859 gnd.n3021 gnd.n0 8.10675
R13860 gnd.n8103 gnd.n8102 8.10675
R13861 gnd.n5748 gnd.n5747 7.97301
R13862 gnd.n6525 gnd.t402 7.9669
R13863 gnd.n6883 gnd.n6882 7.9669
R13864 gnd.n3352 gnd.n3351 7.9669
R13865 gnd.n4079 gnd.t44 7.9669
R13866 gnd.n2215 gnd.t392 7.9669
R13867 gnd.n1820 gnd.n1812 7.9669
R13868 gnd.n8103 gnd.n98 7.95236
R13869 gnd.n4553 gnd.n4415 7.75808
R13870 gnd.n3364 gnd.n2552 7.75808
R13871 gnd.n451 gnd.n371 7.75808
R13872 gnd.n2955 gnd.n2954 7.75808
R13873 gnd.n6883 gnd.t171 7.64824
R13874 gnd.n2824 gnd.n1399 7.64824
R13875 gnd.n2881 gnd.n2808 7.64824
R13876 gnd.n3024 gnd.n2797 7.64824
R13877 gnd.n3040 gnd.n2799 7.64824
R13878 gnd.n3046 gnd.n2792 7.64824
R13879 gnd.n3055 gnd.n2784 7.64824
R13880 gnd.n3054 gnd.n1412 7.64824
R13881 gnd.n5185 gnd.n1415 7.64824
R13882 gnd.n3085 gnd.n3084 7.64824
R13883 gnd.n5179 gnd.n1426 7.64824
R13884 gnd.n3093 gnd.n1433 7.64824
R13885 gnd.n5173 gnd.n1436 7.64824
R13886 gnd.n3099 gnd.n1443 7.64824
R13887 gnd.n5167 gnd.n1446 7.64824
R13888 gnd.n3107 gnd.n1454 7.64824
R13889 gnd.n5161 gnd.n1457 7.64824
R13890 gnd.n3143 gnd.n3142 7.64824
R13891 gnd.n5155 gnd.n1466 7.64824
R13892 gnd.n3114 gnd.n1474 7.64824
R13893 gnd.n5149 gnd.n1477 7.64824
R13894 gnd.n3118 gnd.n1484 7.64824
R13895 gnd.n5143 gnd.n1487 7.64824
R13896 gnd.n3125 gnd.n1495 7.64824
R13897 gnd.n5137 gnd.n1498 7.64824
R13898 gnd.n3186 gnd.n3185 7.64824
R13899 gnd.n5131 gnd.n1507 7.64824
R13900 gnd.n3193 gnd.n1515 7.64824
R13901 gnd.n5125 gnd.n1518 7.64824
R13902 gnd.n3201 gnd.n1525 7.64824
R13903 gnd.n5119 gnd.n1528 7.64824
R13904 gnd.n3208 gnd.n1536 7.64824
R13905 gnd.n5113 gnd.n1539 7.64824
R13906 gnd.n5107 gnd.n1549 7.64824
R13907 gnd.n3361 gnd.n3360 7.64824
R13908 gnd.t2 gnd.n2371 7.64824
R13909 gnd.t12 gnd.n2324 7.64824
R13910 gnd.n3965 gnd.t398 7.64824
R13911 gnd.n3639 gnd.t177 7.64824
R13912 gnd.n4716 gnd.n1934 7.64824
R13913 gnd.n4713 gnd.n1936 7.64824
R13914 gnd.n4707 gnd.n1950 7.64824
R13915 gnd.n4579 gnd.n1953 7.64824
R13916 gnd.n4701 gnd.n1961 7.64824
R13917 gnd.n4587 gnd.n1964 7.64824
R13918 gnd.n4695 gnd.n1972 7.64824
R13919 gnd.n4593 gnd.n1975 7.64824
R13920 gnd.n4689 gnd.n1982 7.64824
R13921 gnd.n4601 gnd.n2120 7.64824
R13922 gnd.n4683 gnd.n1992 7.64824
R13923 gnd.n4607 gnd.n1995 7.64824
R13924 gnd.n4677 gnd.n2002 7.64824
R13925 gnd.n4615 gnd.n2005 7.64824
R13926 gnd.n4671 gnd.n2013 7.64824
R13927 gnd.n4624 gnd.n2016 7.64824
R13928 gnd.n4665 gnd.n2023 7.64824
R13929 gnd.n4641 gnd.n4640 7.64824
R13930 gnd.n4659 gnd.n2034 7.64824
R13931 gnd.n4652 gnd.n2037 7.64824
R13932 gnd.n4651 gnd.n2045 7.64824
R13933 gnd.n7757 gnd.n542 7.64824
R13934 gnd.n7744 gnd.n7743 7.64824
R13935 gnd.n7768 gnd.n532 7.64824
R13936 gnd.n7750 gnd.n534 7.64824
R13937 gnd.n7776 gnd.n526 7.64824
R13938 gnd.n7790 gnd.n515 7.64824
R13939 gnd.n7795 gnd.n510 7.64824
R13940 gnd.n7784 gnd.n522 7.64824
R13941 gnd.n7803 gnd.n502 7.64824
R13942 gnd.n7813 gnd.n497 7.64824
R13943 gnd.n7808 gnd.n500 7.64824
R13944 gnd.n7822 gnd.n491 7.64824
R13945 gnd.n8097 gnd.n105 7.64824
R13946 gnd.n6328 gnd.n6327 7.53171
R13947 gnd.t22 gnd.n6474 7.32958
R13948 gnd.n3381 gnd.t102 7.32958
R13949 gnd.n2509 gnd.t18 7.32958
R13950 gnd.t399 gnd.n2163 7.32958
R13951 gnd.n4400 gnd.t66 7.32958
R13952 gnd.n1684 gnd.n1683 7.30353
R13953 gnd.n3723 gnd.n3722 7.30353
R13954 gnd.n6433 gnd.n6432 7.01093
R13955 gnd.n6444 gnd.n6009 7.01093
R13956 gnd.n6443 gnd.n6012 7.01093
R13957 gnd.n6454 gnd.n6002 7.01093
R13958 gnd.n6352 gnd.n5995 7.01093
R13959 gnd.n6464 gnd.n6463 7.01093
R13960 gnd.n6475 gnd.n5984 7.01093
R13961 gnd.n6474 gnd.n5987 7.01093
R13962 gnd.n6485 gnd.n5975 7.01093
R13963 gnd.n5978 gnd.n5976 7.01093
R13964 gnd.n6495 gnd.n6494 7.01093
R13965 gnd.n6506 gnd.n5958 7.01093
R13966 gnd.n6516 gnd.n5949 7.01093
R13967 gnd.n5952 gnd.n5950 7.01093
R13968 gnd.n6526 gnd.n6525 7.01093
R13969 gnd.n6537 gnd.n5932 7.01093
R13970 gnd.n6547 gnd.n5924 7.01093
R13971 gnd.n5925 gnd.n5917 7.01093
R13972 gnd.n6568 gnd.n5906 7.01093
R13973 gnd.n6567 gnd.n5909 7.01093
R13974 gnd.n6578 gnd.n5899 7.01093
R13975 gnd.n6236 gnd.n5892 7.01093
R13976 gnd.n6588 gnd.n6587 7.01093
R13977 gnd.n6599 gnd.n5881 7.01093
R13978 gnd.n6598 gnd.n5884 7.01093
R13979 gnd.n5874 gnd.n5867 7.01093
R13980 gnd.n6619 gnd.n6618 7.01093
R13981 gnd.n6629 gnd.n5857 7.01093
R13982 gnd.n6628 gnd.n5860 7.01093
R13983 gnd.n6639 gnd.n5850 7.01093
R13984 gnd.n6649 gnd.n5843 7.01093
R13985 gnd.n6660 gnd.n5837 7.01093
R13986 gnd.n6683 gnd.n5818 7.01093
R13987 gnd.n6693 gnd.n5809 7.01093
R13988 gnd.n5808 gnd.n5801 7.01093
R13989 gnd.n6704 gnd.n6703 7.01093
R13990 gnd.n6717 gnd.n5795 7.01093
R13991 gnd.n6716 gnd.n6715 7.01093
R13992 gnd.n5788 gnd.n5774 7.01093
R13993 gnd.n6749 gnd.n6748 7.01093
R13994 gnd.n6760 gnd.n5768 7.01093
R13995 gnd.n6759 gnd.n5489 7.01093
R13996 gnd.n6779 gnd.n5490 7.01093
R13997 gnd.n6771 gnd.n5761 7.01093
R13998 gnd.n6882 gnd.n1137 7.01093
R13999 gnd.n6786 gnd.n1145 7.01093
R14000 gnd.n6876 gnd.n6875 7.01093
R14001 gnd.n4974 gnd.n1691 7.01093
R14002 gnd.n4041 gnd.n3508 7.01093
R14003 gnd.n4004 gnd.n3553 7.01093
R14004 gnd.n4211 gnd.n2289 7.01093
R14005 gnd.n4259 gnd.n2248 7.01093
R14006 gnd.n3885 gnd.n3884 7.01093
R14007 gnd.n5978 gnd.t4 6.69227
R14008 gnd.n6619 gnd.t35 6.69227
R14009 gnd.n6729 gnd.t37 6.69227
R14010 gnd.n3869 gnd.n3868 6.5566
R14011 gnd.n2414 gnd.n2413 6.5566
R14012 gnd.n4986 gnd.n4982 6.5566
R14013 gnd.n3788 gnd.n3787 6.5566
R14014 gnd.n4331 gnd.t74 6.37362
R14015 gnd.n3287 gnd.n3284 6.20656
R14016 gnd.n4556 gnd.n4412 6.20656
R14017 gnd.n6536 gnd.t29 6.05496
R14018 gnd.n5935 gnd.t34 6.05496
R14019 gnd.n6236 gnd.t403 6.05496
R14020 gnd.n6670 gnd.t53 6.05496
R14021 gnd.n5745 gnd.n5715 5.81868
R14022 gnd.n5713 gnd.n5683 5.81868
R14023 gnd.n5681 gnd.n5651 5.81868
R14024 gnd.n5650 gnd.n5620 5.81868
R14025 gnd.n5618 gnd.n5588 5.81868
R14026 gnd.n5586 gnd.n5556 5.81868
R14027 gnd.n5554 gnd.n5524 5.81868
R14028 gnd.n5523 gnd.n5493 5.81868
R14029 gnd.n2473 gnd.t77 5.73631
R14030 gnd.n4062 gnd.t5 5.73631
R14031 gnd.n4131 gnd.n2359 5.73631
R14032 gnd.n4049 gnd.n4048 5.73631
R14033 gnd.t178 gnd.n2330 5.73631
R14034 gnd.n3553 gnd.t42 5.73631
R14035 gnd.n3997 gnd.n3996 5.73631
R14036 gnd.n4203 gnd.n2296 5.73631
R14037 gnd.n4211 gnd.t43 5.73631
R14038 gnd.n3956 gnd.t23 5.73631
R14039 gnd.n4267 gnd.n2241 5.73631
R14040 gnd.n3927 gnd.n3622 5.73631
R14041 gnd.n3920 gnd.t13 5.73631
R14042 gnd.t128 gnd.n3670 5.73631
R14043 gnd.n3873 gnd.n1891 5.62001
R14044 gnd.n5048 gnd.n1626 5.62001
R14045 gnd.n5048 gnd.n1627 5.62001
R14046 gnd.n3792 gnd.n1891 5.62001
R14047 gnd.n6106 gnd.n6105 5.4308
R14048 gnd.n5478 gnd.n5476 5.4308
R14049 gnd.n6588 gnd.t401 5.41765
R14050 gnd.n6609 gnd.t180 5.41765
R14051 gnd.t40 gnd.n5827 5.41765
R14052 gnd.n5743 gnd.n5742 5.04292
R14053 gnd.n5711 gnd.n5710 5.04292
R14054 gnd.n5679 gnd.n5678 5.04292
R14055 gnd.n5648 gnd.n5647 5.04292
R14056 gnd.n5616 gnd.n5615 5.04292
R14057 gnd.n5584 gnd.n5583 5.04292
R14058 gnd.n5552 gnd.n5551 5.04292
R14059 gnd.n5521 gnd.n5520 5.04292
R14060 gnd.n6557 gnd.t21 4.78034
R14061 gnd.n6639 gnd.t406 4.78034
R14062 gnd.t189 gnd.n1630 4.78034
R14063 gnd.n4048 gnd.t14 4.78034
R14064 gnd.t38 gnd.n2241 4.78034
R14065 gnd.n3876 gnd.t147 4.78034
R14066 gnd.n4339 gnd.t24 4.78034
R14067 gnd.n6331 gnd.n6330 4.74817
R14068 gnd.n6248 gnd.n6244 4.74817
R14069 gnd.n6241 gnd.n6240 4.74817
R14070 gnd.n6235 gnd.n6214 4.74817
R14071 gnd.n6330 gnd.n6212 4.74817
R14072 gnd.n6248 gnd.n6247 4.74817
R14073 gnd.n6243 gnd.n6241 4.74817
R14074 gnd.n6239 gnd.n6214 4.74817
R14075 gnd.n7793 gnd.n118 4.74817
R14076 gnd.n7810 gnd.n117 4.74817
R14077 gnd.n7806 gnd.n116 4.74817
R14078 gnd.n8095 gnd.n111 4.74817
R14079 gnd.n8093 gnd.n112 4.74817
R14080 gnd.n514 gnd.n118 4.74817
R14081 gnd.n7792 gnd.n117 4.74817
R14082 gnd.n7811 gnd.n116 4.74817
R14083 gnd.n7805 gnd.n111 4.74817
R14084 gnd.n8094 gnd.n8093 4.74817
R14085 gnd.n1401 gnd.n1384 4.74817
R14086 gnd.n5189 gnd.n1402 4.74817
R14087 gnd.n2795 gnd.n1407 4.74817
R14088 gnd.n3044 gnd.n1406 4.74817
R14089 gnd.n1408 gnd.n1405 4.74817
R14090 gnd.n5200 gnd.n1384 4.74817
R14091 gnd.n5190 gnd.n5189 4.74817
R14092 gnd.n2879 gnd.n1407 4.74817
R14093 gnd.n2796 gnd.n1406 4.74817
R14094 gnd.n3043 gnd.n1405 4.74817
R14095 gnd.n6327 gnd.n6326 4.74296
R14096 gnd.n98 gnd.n97 4.74296
R14097 gnd.n6287 gnd.n6286 4.7074
R14098 gnd.n6307 gnd.n6306 4.7074
R14099 gnd.n58 gnd.n57 4.7074
R14100 gnd.n78 gnd.n77 4.7074
R14101 gnd.n6327 gnd.n6307 4.65959
R14102 gnd.n98 gnd.n78 4.65959
R14103 gnd.n4783 gnd.n1893 4.6132
R14104 gnd.n5049 gnd.n1625 4.6132
R14105 gnd.n2473 gnd.n1688 4.46168
R14106 gnd.t70 gnd.n1703 4.46168
R14107 gnd.n4056 gnd.n3495 4.46168
R14108 gnd.n4139 gnd.n2352 4.46168
R14109 gnd.n4195 gnd.n2303 4.46168
R14110 gnd.n3988 gnd.n3566 4.46168
R14111 gnd.n3935 gnd.n3934 4.46168
R14112 gnd.n4275 gnd.n2234 4.46168
R14113 gnd.n3892 gnd.t115 4.46168
R14114 gnd.n4331 gnd.n2187 4.46168
R14115 gnd.n3719 gnd.n3706 4.46111
R14116 gnd.n5728 gnd.n5724 4.38594
R14117 gnd.n5696 gnd.n5692 4.38594
R14118 gnd.n5664 gnd.n5660 4.38594
R14119 gnd.n5633 gnd.n5629 4.38594
R14120 gnd.n5601 gnd.n5597 4.38594
R14121 gnd.n5569 gnd.n5565 4.38594
R14122 gnd.n5537 gnd.n5533 4.38594
R14123 gnd.n5506 gnd.n5502 4.38594
R14124 gnd.n5739 gnd.n5717 4.26717
R14125 gnd.n5707 gnd.n5685 4.26717
R14126 gnd.n5675 gnd.n5653 4.26717
R14127 gnd.n5644 gnd.n5622 4.26717
R14128 gnd.n5612 gnd.n5590 4.26717
R14129 gnd.n5580 gnd.n5558 4.26717
R14130 gnd.n5548 gnd.n5526 4.26717
R14131 gnd.n5517 gnd.n5495 4.26717
R14132 gnd.t31 gnd.n5961 4.14303
R14133 gnd.n6703 gnd.t3 4.14303
R14134 gnd.t94 gnd.n1546 4.14303
R14135 gnd.n3546 gnd.t48 4.14303
R14136 gnd.t394 gnd.n2276 4.14303
R14137 gnd.t62 gnd.n1941 4.14303
R14138 gnd.n5747 gnd.n5746 4.08274
R14139 gnd.n3868 gnd.n3867 4.05904
R14140 gnd.n2415 gnd.n2414 4.05904
R14141 gnd.n4989 gnd.n4982 4.05904
R14142 gnd.n3787 gnd.n3786 4.05904
R14143 gnd.n19 gnd.n9 3.99943
R14144 gnd.t137 gnd.n1691 3.82437
R14145 gnd.n3508 gnd.t179 3.82437
R14146 gnd.n4259 gnd.t33 3.82437
R14147 gnd.n3671 gnd.t128 3.82437
R14148 gnd.t115 gnd.t106 3.82437
R14149 gnd.n6329 gnd.n6328 3.81325
R14150 gnd.n6307 gnd.n6287 3.72967
R14151 gnd.n78 gnd.n58 3.72967
R14152 gnd.n5747 gnd.n5619 3.70378
R14153 gnd.n19 gnd.n18 3.60163
R14154 gnd.n1270 gnd.t98 3.50571
R14155 gnd.n3218 gnd.t94 3.50571
R14156 gnd.t46 gnd.n1701 3.50571
R14157 gnd.n3659 gnd.t55 3.50571
R14158 gnd.n4573 gnd.t62 3.50571
R14159 gnd.t83 gnd.n241 3.50571
R14160 gnd.n5738 gnd.n5719 3.49141
R14161 gnd.n5706 gnd.n5687 3.49141
R14162 gnd.n5674 gnd.n5655 3.49141
R14163 gnd.n5643 gnd.n5624 3.49141
R14164 gnd.n5611 gnd.n5592 3.49141
R14165 gnd.n5579 gnd.n5560 3.49141
R14166 gnd.n5547 gnd.n5528 3.49141
R14167 gnd.n5516 gnd.n5497 3.49141
R14168 gnd.n4801 gnd.n4800 3.29747
R14169 gnd.n4800 gnd.n4799 3.29747
R14170 gnd.n7970 gnd.n7967 3.29747
R14171 gnd.n7971 gnd.n7970 3.29747
R14172 gnd.n5365 gnd.n5364 3.29747
R14173 gnd.n5364 gnd.n5363 3.29747
R14174 gnd.n5067 gnd.n5066 3.29747
R14175 gnd.n5066 gnd.n5065 3.29747
R14176 gnd.n3456 gnd.n3455 3.18706
R14177 gnd.n4063 gnd.n3486 3.18706
R14178 gnd.n4147 gnd.n2345 3.18706
R14179 gnd.n4187 gnd.n2310 3.18706
R14180 gnd.n3981 gnd.n3980 3.18706
R14181 gnd.n3942 gnd.n3608 3.18706
R14182 gnd.n4283 gnd.n2228 3.18706
R14183 gnd.n4323 gnd.n2193 3.18706
R14184 gnd.n6505 gnd.t31 2.8684
R14185 gnd.n2799 gnd.t267 2.8684
R14186 gnd.n4099 gnd.t44 2.8684
R14187 gnd.t392 gnd.n2214 2.8684
R14188 gnd.t224 gnd.n497 2.8684
R14189 gnd.n6308 gnd.t316 2.82907
R14190 gnd.n6308 gnd.t390 2.82907
R14191 gnd.n6310 gnd.t271 2.82907
R14192 gnd.n6310 gnd.t371 2.82907
R14193 gnd.n6312 gnd.t208 2.82907
R14194 gnd.n6312 gnd.t349 2.82907
R14195 gnd.n6314 gnd.t377 2.82907
R14196 gnd.n6314 gnd.t269 2.82907
R14197 gnd.n6316 gnd.t302 2.82907
R14198 gnd.n6316 gnd.t281 2.82907
R14199 gnd.n6318 gnd.t280 2.82907
R14200 gnd.n6318 gnd.t250 2.82907
R14201 gnd.n6320 gnd.t289 2.82907
R14202 gnd.n6320 gnd.t336 2.82907
R14203 gnd.n6322 gnd.t343 2.82907
R14204 gnd.n6322 gnd.t290 2.82907
R14205 gnd.n6324 gnd.t327 2.82907
R14206 gnd.n6324 gnd.t223 2.82907
R14207 gnd.n6249 gnd.t326 2.82907
R14208 gnd.n6249 gnd.t332 2.82907
R14209 gnd.n6251 gnd.t356 2.82907
R14210 gnd.n6251 gnd.t381 2.82907
R14211 gnd.n6253 gnd.t313 2.82907
R14212 gnd.n6253 gnd.t330 2.82907
R14213 gnd.n6255 gnd.t345 2.82907
R14214 gnd.n6255 gnd.t236 2.82907
R14215 gnd.n6257 gnd.t329 2.82907
R14216 gnd.n6257 gnd.t325 2.82907
R14217 gnd.n6259 gnd.t364 2.82907
R14218 gnd.n6259 gnd.t357 2.82907
R14219 gnd.n6261 gnd.t259 2.82907
R14220 gnd.n6261 gnd.t340 2.82907
R14221 gnd.n6263 gnd.t378 2.82907
R14222 gnd.n6263 gnd.t238 2.82907
R14223 gnd.n6265 gnd.t263 2.82907
R14224 gnd.n6265 gnd.t354 2.82907
R14225 gnd.n6268 gnd.t305 2.82907
R14226 gnd.n6268 gnd.t294 2.82907
R14227 gnd.n6270 gnd.t278 2.82907
R14228 gnd.n6270 gnd.t320 2.82907
R14229 gnd.n6272 gnd.t266 2.82907
R14230 gnd.n6272 gnd.t306 2.82907
R14231 gnd.n6274 gnd.t307 2.82907
R14232 gnd.n6274 gnd.t283 2.82907
R14233 gnd.n6276 gnd.t204 2.82907
R14234 gnd.n6276 gnd.t268 2.82907
R14235 gnd.n6278 gnd.t254 2.82907
R14236 gnd.n6278 gnd.t309 2.82907
R14237 gnd.n6280 gnd.t241 2.82907
R14238 gnd.n6280 gnd.t206 2.82907
R14239 gnd.n6282 gnd.t215 2.82907
R14240 gnd.n6282 gnd.t264 2.82907
R14241 gnd.n6284 gnd.t265 2.82907
R14242 gnd.n6284 gnd.t234 2.82907
R14243 gnd.n6288 gnd.t362 2.82907
R14244 gnd.n6288 gnd.t311 2.82907
R14245 gnd.n6290 gnd.t339 2.82907
R14246 gnd.n6290 gnd.t286 2.82907
R14247 gnd.n6292 gnd.t315 2.82907
R14248 gnd.n6292 gnd.t220 2.82907
R14249 gnd.n6294 gnd.t292 2.82907
R14250 gnd.n6294 gnd.t337 2.82907
R14251 gnd.n6296 gnd.t319 2.82907
R14252 gnd.n6296 gnd.t335 2.82907
R14253 gnd.n6298 gnd.t341 2.82907
R14254 gnd.n6298 gnd.t318 2.82907
R14255 gnd.n6300 gnd.t346 2.82907
R14256 gnd.n6300 gnd.t387 2.82907
R14257 gnd.n6302 gnd.t212 2.82907
R14258 gnd.n6302 gnd.t350 2.82907
R14259 gnd.n6304 gnd.t379 2.82907
R14260 gnd.n6304 gnd.t324 2.82907
R14261 gnd.n95 gnd.t334 2.82907
R14262 gnd.n95 gnd.t218 2.82907
R14263 gnd.n93 gnd.t361 2.82907
R14264 gnd.n93 gnd.t248 2.82907
R14265 gnd.n91 gnd.t296 2.82907
R14266 gnd.n91 gnd.t347 2.82907
R14267 gnd.n89 gnd.t372 2.82907
R14268 gnd.n89 gnd.t384 2.82907
R14269 gnd.n87 gnd.t388 2.82907
R14270 gnd.n87 gnd.t261 2.82907
R14271 gnd.n85 gnd.t382 2.82907
R14272 gnd.n85 gnd.t342 2.82907
R14273 gnd.n83 gnd.t312 2.82907
R14274 gnd.n83 gnd.t368 2.82907
R14275 gnd.n81 gnd.t338 2.82907
R14276 gnd.n81 gnd.t383 2.82907
R14277 gnd.n79 gnd.t353 2.82907
R14278 gnd.n79 gnd.t246 2.82907
R14279 gnd.n36 gnd.t360 2.82907
R14280 gnd.n36 gnd.t287 2.82907
R14281 gnd.n34 gnd.t256 2.82907
R14282 gnd.n34 gnd.t386 2.82907
R14283 gnd.n32 gnd.t370 2.82907
R14284 gnd.n32 gnd.t239 2.82907
R14285 gnd.n30 gnd.t198 2.82907
R14286 gnd.n30 gnd.t221 2.82907
R14287 gnd.n28 gnd.t351 2.82907
R14288 gnd.n28 gnd.t322 2.82907
R14289 gnd.n26 gnd.t301 2.82907
R14290 gnd.n26 gnd.t376 2.82907
R14291 gnd.n24 gnd.t363 2.82907
R14292 gnd.n24 gnd.t288 2.82907
R14293 gnd.n22 gnd.t258 2.82907
R14294 gnd.n22 gnd.t192 2.82907
R14295 gnd.n20 gnd.t375 2.82907
R14296 gnd.n20 gnd.t352 2.82907
R14297 gnd.n55 gnd.t369 2.82907
R14298 gnd.n55 gnd.t389 2.82907
R14299 gnd.n53 gnd.t385 2.82907
R14300 gnd.n53 gnd.t365 2.82907
R14301 gnd.n51 gnd.t373 2.82907
R14302 gnd.n51 gnd.t257 2.82907
R14303 gnd.n49 gnd.t277 2.82907
R14304 gnd.n49 gnd.t214 2.82907
R14305 gnd.n47 gnd.t225 2.82907
R14306 gnd.n47 gnd.t243 2.82907
R14307 gnd.n45 gnd.t245 2.82907
R14308 gnd.n45 gnd.t279 2.82907
R14309 gnd.n43 gnd.t276 2.82907
R14310 gnd.n43 gnd.t299 2.82907
R14311 gnd.n41 gnd.t297 2.82907
R14312 gnd.n41 gnd.t251 2.82907
R14313 gnd.n39 gnd.t252 2.82907
R14314 gnd.n39 gnd.t196 2.82907
R14315 gnd.n75 gnd.t380 2.82907
R14316 gnd.n75 gnd.t321 2.82907
R14317 gnd.n73 gnd.t260 2.82907
R14318 gnd.n73 gnd.t317 2.82907
R14319 gnd.n71 gnd.t348 2.82907
R14320 gnd.n71 gnd.t231 2.82907
R14321 gnd.n69 gnd.t282 2.82907
R14322 gnd.n69 gnd.t303 2.82907
R14323 gnd.n67 gnd.t308 2.82907
R14324 gnd.n67 gnd.t331 2.82907
R14325 gnd.n65 gnd.t274 2.82907
R14326 gnd.n65 gnd.t194 2.82907
R14327 gnd.n63 gnd.t358 2.82907
R14328 gnd.n63 gnd.t273 2.82907
R14329 gnd.n61 gnd.t200 2.82907
R14330 gnd.n61 gnd.t300 2.82907
R14331 gnd.n59 gnd.t233 2.82907
R14332 gnd.n59 gnd.t328 2.82907
R14333 gnd.n5735 gnd.n5734 2.71565
R14334 gnd.n5703 gnd.n5702 2.71565
R14335 gnd.n5671 gnd.n5670 2.71565
R14336 gnd.n5640 gnd.n5639 2.71565
R14337 gnd.n5608 gnd.n5607 2.71565
R14338 gnd.n5576 gnd.n5575 2.71565
R14339 gnd.n5544 gnd.n5543 2.71565
R14340 gnd.n5513 gnd.n5512 2.71565
R14341 gnd.n4050 gnd.t20 2.54975
R14342 gnd.n4034 gnd.t28 2.54975
R14343 gnd.t6 gnd.n2254 2.54975
R14344 gnd.t27 gnd.n2242 2.54975
R14345 gnd.n6330 gnd.n6329 2.27742
R14346 gnd.n6329 gnd.n6248 2.27742
R14347 gnd.n6329 gnd.n6241 2.27742
R14348 gnd.n6329 gnd.n6214 2.27742
R14349 gnd.n8092 gnd.n118 2.27742
R14350 gnd.n8092 gnd.n117 2.27742
R14351 gnd.n8092 gnd.n116 2.27742
R14352 gnd.n8092 gnd.n111 2.27742
R14353 gnd.n8093 gnd.n8092 2.27742
R14354 gnd.n5188 gnd.n1384 2.27742
R14355 gnd.n5189 gnd.n5188 2.27742
R14356 gnd.n5188 gnd.n1407 2.27742
R14357 gnd.n5188 gnd.n1406 2.27742
R14358 gnd.n5188 gnd.n1405 2.27742
R14359 gnd.t87 gnd.n6443 2.23109
R14360 gnd.t21 gnd.n6556 2.23109
R14361 gnd.t207 gnd.n1436 2.23109
R14362 gnd.n7743 gnd.t272 2.23109
R14363 gnd.n5731 gnd.n5721 1.93989
R14364 gnd.n5699 gnd.n5689 1.93989
R14365 gnd.n5667 gnd.n5657 1.93989
R14366 gnd.n5636 gnd.n5626 1.93989
R14367 gnd.n5604 gnd.n5594 1.93989
R14368 gnd.n5572 gnd.n5562 1.93989
R14369 gnd.n5540 gnd.n5530 1.93989
R14370 gnd.n5509 gnd.n5499 1.93989
R14371 gnd.n3464 gnd.n3463 1.91244
R14372 gnd.n4070 gnd.n3476 1.91244
R14373 gnd.n4179 gnd.n2317 1.91244
R14374 gnd.n3972 gnd.n3580 1.91244
R14375 gnd.n4291 gnd.n2221 1.91244
R14376 gnd.n4315 gnd.n2200 1.91244
R14377 gnd.n6352 gnd.t10 1.59378
R14378 gnd.n6228 gnd.t180 1.59378
R14379 gnd.n6669 gnd.t40 1.59378
R14380 gnd.t222 gnd.n1314 1.59378
R14381 gnd.t285 gnd.n1477 1.59378
R14382 gnd.n3125 gnd.t304 1.59378
R14383 gnd.n4155 gnd.t50 1.59378
R14384 gnd.t183 gnd.n3601 1.59378
R14385 gnd.n4607 gnd.t195 1.59378
R14386 gnd.t199 gnd.n2013 1.59378
R14387 gnd.n199 gnd.t333 1.59378
R14388 gnd.n3465 gnd.t165 1.27512
R14389 gnd.n4123 gnd.t5 1.27512
R14390 gnd.t13 gnd.n3631 1.27512
R14391 gnd.t134 gnd.n2193 1.27512
R14392 gnd.n6107 gnd.n6106 1.16414
R14393 gnd.n6801 gnd.n5476 1.16414
R14394 gnd.n5730 gnd.n5723 1.16414
R14395 gnd.n5698 gnd.n5691 1.16414
R14396 gnd.n5666 gnd.n5659 1.16414
R14397 gnd.n5635 gnd.n5628 1.16414
R14398 gnd.n5603 gnd.n5596 1.16414
R14399 gnd.n5571 gnd.n5564 1.16414
R14400 gnd.n5539 gnd.n5532 1.16414
R14401 gnd.n5508 gnd.n5501 1.16414
R14402 gnd.n4783 gnd.n4782 0.970197
R14403 gnd.n5049 gnd.n1623 0.970197
R14404 gnd.n5714 gnd.n5682 0.962709
R14405 gnd.n5746 gnd.n5714 0.962709
R14406 gnd.n5587 gnd.n5555 0.962709
R14407 gnd.n5619 gnd.n5587 0.962709
R14408 gnd.t29 gnd.n5935 0.956468
R14409 gnd.n6659 gnd.t53 0.956468
R14410 gnd.t240 gnd.n1352 0.956468
R14411 gnd.n3107 gnd.t219 0.956468
R14412 gnd.t209 gnd.n1518 0.956468
R14413 gnd.t228 gnd.n1972 0.956468
R14414 gnd.n4652 gnd.t275 0.956468
R14415 gnd.n161 gnd.t230 0.956468
R14416 gnd gnd.n0 0.70738
R14417 gnd.n2 gnd.n1 0.672012
R14418 gnd.n3 gnd.n2 0.672012
R14419 gnd.n4 gnd.n3 0.672012
R14420 gnd.n5 gnd.n4 0.672012
R14421 gnd.n6 gnd.n5 0.672012
R14422 gnd.n7 gnd.n6 0.672012
R14423 gnd.n8 gnd.n7 0.672012
R14424 gnd.n9 gnd.n8 0.672012
R14425 gnd.n11 gnd.n10 0.672012
R14426 gnd.n12 gnd.n11 0.672012
R14427 gnd.n13 gnd.n12 0.672012
R14428 gnd.n14 gnd.n13 0.672012
R14429 gnd.n15 gnd.n14 0.672012
R14430 gnd.n16 gnd.n15 0.672012
R14431 gnd.n17 gnd.n16 0.672012
R14432 gnd.n18 gnd.n17 0.672012
R14433 gnd.n2393 gnd.n2392 0.637812
R14434 gnd.n4078 gnd.n4077 0.637812
R14435 gnd.n4077 gnd.t26 0.637812
R14436 gnd.n4163 gnd.n2330 0.637812
R14437 gnd.n4171 gnd.n2324 0.637812
R14438 gnd.n4013 gnd.t391 0.637812
R14439 gnd.t9 gnd.n2283 0.637812
R14440 gnd.n3965 gnd.n3964 0.637812
R14441 gnd.n3956 gnd.n3593 0.637812
R14442 gnd.t405 gnd.n2213 0.637812
R14443 gnd.n4299 gnd.n2213 0.637812
R14444 gnd.n4307 gnd.n2207 0.637812
R14445 gnd.n8104 gnd.n8103 0.637193
R14446 gnd.n6326 gnd.n6325 0.573776
R14447 gnd.n6325 gnd.n6323 0.573776
R14448 gnd.n6323 gnd.n6321 0.573776
R14449 gnd.n6321 gnd.n6319 0.573776
R14450 gnd.n6319 gnd.n6317 0.573776
R14451 gnd.n6317 gnd.n6315 0.573776
R14452 gnd.n6315 gnd.n6313 0.573776
R14453 gnd.n6313 gnd.n6311 0.573776
R14454 gnd.n6311 gnd.n6309 0.573776
R14455 gnd.n6267 gnd.n6266 0.573776
R14456 gnd.n6266 gnd.n6264 0.573776
R14457 gnd.n6264 gnd.n6262 0.573776
R14458 gnd.n6262 gnd.n6260 0.573776
R14459 gnd.n6260 gnd.n6258 0.573776
R14460 gnd.n6258 gnd.n6256 0.573776
R14461 gnd.n6256 gnd.n6254 0.573776
R14462 gnd.n6254 gnd.n6252 0.573776
R14463 gnd.n6252 gnd.n6250 0.573776
R14464 gnd.n6286 gnd.n6285 0.573776
R14465 gnd.n6285 gnd.n6283 0.573776
R14466 gnd.n6283 gnd.n6281 0.573776
R14467 gnd.n6281 gnd.n6279 0.573776
R14468 gnd.n6279 gnd.n6277 0.573776
R14469 gnd.n6277 gnd.n6275 0.573776
R14470 gnd.n6275 gnd.n6273 0.573776
R14471 gnd.n6273 gnd.n6271 0.573776
R14472 gnd.n6271 gnd.n6269 0.573776
R14473 gnd.n6306 gnd.n6305 0.573776
R14474 gnd.n6305 gnd.n6303 0.573776
R14475 gnd.n6303 gnd.n6301 0.573776
R14476 gnd.n6301 gnd.n6299 0.573776
R14477 gnd.n6299 gnd.n6297 0.573776
R14478 gnd.n6297 gnd.n6295 0.573776
R14479 gnd.n6295 gnd.n6293 0.573776
R14480 gnd.n6293 gnd.n6291 0.573776
R14481 gnd.n6291 gnd.n6289 0.573776
R14482 gnd.n82 gnd.n80 0.573776
R14483 gnd.n84 gnd.n82 0.573776
R14484 gnd.n86 gnd.n84 0.573776
R14485 gnd.n88 gnd.n86 0.573776
R14486 gnd.n90 gnd.n88 0.573776
R14487 gnd.n92 gnd.n90 0.573776
R14488 gnd.n94 gnd.n92 0.573776
R14489 gnd.n96 gnd.n94 0.573776
R14490 gnd.n97 gnd.n96 0.573776
R14491 gnd.n23 gnd.n21 0.573776
R14492 gnd.n25 gnd.n23 0.573776
R14493 gnd.n27 gnd.n25 0.573776
R14494 gnd.n29 gnd.n27 0.573776
R14495 gnd.n31 gnd.n29 0.573776
R14496 gnd.n33 gnd.n31 0.573776
R14497 gnd.n35 gnd.n33 0.573776
R14498 gnd.n37 gnd.n35 0.573776
R14499 gnd.n38 gnd.n37 0.573776
R14500 gnd.n42 gnd.n40 0.573776
R14501 gnd.n44 gnd.n42 0.573776
R14502 gnd.n46 gnd.n44 0.573776
R14503 gnd.n48 gnd.n46 0.573776
R14504 gnd.n50 gnd.n48 0.573776
R14505 gnd.n52 gnd.n50 0.573776
R14506 gnd.n54 gnd.n52 0.573776
R14507 gnd.n56 gnd.n54 0.573776
R14508 gnd.n57 gnd.n56 0.573776
R14509 gnd.n62 gnd.n60 0.573776
R14510 gnd.n64 gnd.n62 0.573776
R14511 gnd.n66 gnd.n64 0.573776
R14512 gnd.n68 gnd.n66 0.573776
R14513 gnd.n70 gnd.n68 0.573776
R14514 gnd.n72 gnd.n70 0.573776
R14515 gnd.n74 gnd.n72 0.573776
R14516 gnd.n76 gnd.n74 0.573776
R14517 gnd.n77 gnd.n76 0.573776
R14518 gnd.n6791 gnd.n6790 0.486781
R14519 gnd.n6159 gnd.n6055 0.48678
R14520 gnd.n6872 gnd.n6871 0.480683
R14521 gnd.n6372 gnd.n6006 0.480683
R14522 gnd.n449 gnd.n448 0.477634
R14523 gnd.n2957 gnd.n2956 0.477634
R14524 gnd.n4406 gnd.n4405 0.451719
R14525 gnd.n3370 gnd.n3369 0.451719
R14526 gnd.n2633 gnd.n2632 0.451719
R14527 gnd.n4453 gnd.n1807 0.451719
R14528 gnd.n8007 gnd.n8006 0.442573
R14529 gnd.n1944 gnd.n1863 0.442573
R14530 gnd.n5103 gnd.n5102 0.442573
R14531 gnd.n1264 gnd.n1190 0.442573
R14532 gnd.n7055 gnd.n966 0.425805
R14533 gnd.n7508 gnd.n7507 0.425805
R14534 gnd.n7719 gnd.n568 0.425805
R14535 gnd.n2811 gnd.n2810 0.425805
R14536 gnd.n8092 gnd.n115 0.420375
R14537 gnd.n5188 gnd.n1404 0.420375
R14538 gnd.n3294 gnd.n3284 0.388379
R14539 gnd.n5727 gnd.n5726 0.388379
R14540 gnd.n5695 gnd.n5694 0.388379
R14541 gnd.n5663 gnd.n5662 0.388379
R14542 gnd.n5632 gnd.n5631 0.388379
R14543 gnd.n5600 gnd.n5599 0.388379
R14544 gnd.n5568 gnd.n5567 0.388379
R14545 gnd.n5536 gnd.n5535 0.388379
R14546 gnd.n5505 gnd.n5504 0.388379
R14547 gnd.n4546 gnd.n4412 0.388379
R14548 gnd.n8104 gnd.n19 0.374463
R14549 gnd gnd.n8104 0.367492
R14550 gnd.n6738 gnd.t37 0.319156
R14551 gnd.t249 gnd.n1389 0.319156
R14552 gnd.t291 gnd.n3054 0.319156
R14553 gnd.n4033 gnd.t50 0.319156
R14554 gnd.t42 gnd.t181 0.319156
R14555 gnd.t0 gnd.t43 0.319156
R14556 gnd.n3949 gnd.t183 0.319156
R14557 gnd.n7795 gnd.t193 0.319156
R14558 gnd.t197 gnd.n122 0.319156
R14559 gnd.n6153 gnd.n6152 0.311721
R14560 gnd.n7883 gnd.n485 0.293183
R14561 gnd.n5281 gnd.n1254 0.293183
R14562 gnd.n6841 gnd.n6840 0.268793
R14563 gnd.n7884 gnd.n7883 0.258122
R14564 gnd.n4721 gnd.n4720 0.258122
R14565 gnd.n3224 gnd.n2735 0.258122
R14566 gnd.n5282 gnd.n5281 0.258122
R14567 gnd.n3213 gnd.n2546 0.247451
R14568 gnd.n4568 gnd.n4566 0.247451
R14569 gnd.n6840 gnd.n6839 0.241354
R14570 gnd.n1893 gnd.n1890 0.229039
R14571 gnd.n1894 gnd.n1893 0.229039
R14572 gnd.n1625 gnd.n1622 0.229039
R14573 gnd.n2660 gnd.n1625 0.229039
R14574 gnd.n6328 gnd.n0 0.210825
R14575 gnd.n6427 gnd.n6023 0.206293
R14576 gnd.n5744 gnd.n5716 0.155672
R14577 gnd.n5737 gnd.n5716 0.155672
R14578 gnd.n5737 gnd.n5736 0.155672
R14579 gnd.n5736 gnd.n5720 0.155672
R14580 gnd.n5729 gnd.n5720 0.155672
R14581 gnd.n5729 gnd.n5728 0.155672
R14582 gnd.n5712 gnd.n5684 0.155672
R14583 gnd.n5705 gnd.n5684 0.155672
R14584 gnd.n5705 gnd.n5704 0.155672
R14585 gnd.n5704 gnd.n5688 0.155672
R14586 gnd.n5697 gnd.n5688 0.155672
R14587 gnd.n5697 gnd.n5696 0.155672
R14588 gnd.n5680 gnd.n5652 0.155672
R14589 gnd.n5673 gnd.n5652 0.155672
R14590 gnd.n5673 gnd.n5672 0.155672
R14591 gnd.n5672 gnd.n5656 0.155672
R14592 gnd.n5665 gnd.n5656 0.155672
R14593 gnd.n5665 gnd.n5664 0.155672
R14594 gnd.n5649 gnd.n5621 0.155672
R14595 gnd.n5642 gnd.n5621 0.155672
R14596 gnd.n5642 gnd.n5641 0.155672
R14597 gnd.n5641 gnd.n5625 0.155672
R14598 gnd.n5634 gnd.n5625 0.155672
R14599 gnd.n5634 gnd.n5633 0.155672
R14600 gnd.n5617 gnd.n5589 0.155672
R14601 gnd.n5610 gnd.n5589 0.155672
R14602 gnd.n5610 gnd.n5609 0.155672
R14603 gnd.n5609 gnd.n5593 0.155672
R14604 gnd.n5602 gnd.n5593 0.155672
R14605 gnd.n5602 gnd.n5601 0.155672
R14606 gnd.n5585 gnd.n5557 0.155672
R14607 gnd.n5578 gnd.n5557 0.155672
R14608 gnd.n5578 gnd.n5577 0.155672
R14609 gnd.n5577 gnd.n5561 0.155672
R14610 gnd.n5570 gnd.n5561 0.155672
R14611 gnd.n5570 gnd.n5569 0.155672
R14612 gnd.n5553 gnd.n5525 0.155672
R14613 gnd.n5546 gnd.n5525 0.155672
R14614 gnd.n5546 gnd.n5545 0.155672
R14615 gnd.n5545 gnd.n5529 0.155672
R14616 gnd.n5538 gnd.n5529 0.155672
R14617 gnd.n5538 gnd.n5537 0.155672
R14618 gnd.n5522 gnd.n5494 0.155672
R14619 gnd.n5515 gnd.n5494 0.155672
R14620 gnd.n5515 gnd.n5514 0.155672
R14621 gnd.n5514 gnd.n5498 0.155672
R14622 gnd.n5507 gnd.n5498 0.155672
R14623 gnd.n5507 gnd.n5506 0.155672
R14624 gnd.n6871 gnd.n5406 0.152939
R14625 gnd.n5408 gnd.n5406 0.152939
R14626 gnd.n5412 gnd.n5408 0.152939
R14627 gnd.n5413 gnd.n5412 0.152939
R14628 gnd.n5414 gnd.n5413 0.152939
R14629 gnd.n5415 gnd.n5414 0.152939
R14630 gnd.n5419 gnd.n5415 0.152939
R14631 gnd.n5420 gnd.n5419 0.152939
R14632 gnd.n5421 gnd.n5420 0.152939
R14633 gnd.n5422 gnd.n5421 0.152939
R14634 gnd.n5426 gnd.n5422 0.152939
R14635 gnd.n5427 gnd.n5426 0.152939
R14636 gnd.n5428 gnd.n5427 0.152939
R14637 gnd.n5429 gnd.n5428 0.152939
R14638 gnd.n5434 gnd.n5429 0.152939
R14639 gnd.n6841 gnd.n5434 0.152939
R14640 gnd.n6447 gnd.n6006 0.152939
R14641 gnd.n6448 gnd.n6447 0.152939
R14642 gnd.n6449 gnd.n6448 0.152939
R14643 gnd.n6450 gnd.n6449 0.152939
R14644 gnd.n6450 gnd.n5981 0.152939
R14645 gnd.n6478 gnd.n5981 0.152939
R14646 gnd.n6479 gnd.n6478 0.152939
R14647 gnd.n6480 gnd.n6479 0.152939
R14648 gnd.n6481 gnd.n6480 0.152939
R14649 gnd.n6481 gnd.n5955 0.152939
R14650 gnd.n6509 gnd.n5955 0.152939
R14651 gnd.n6510 gnd.n6509 0.152939
R14652 gnd.n6511 gnd.n6510 0.152939
R14653 gnd.n6512 gnd.n6511 0.152939
R14654 gnd.n6512 gnd.n5929 0.152939
R14655 gnd.n6540 gnd.n5929 0.152939
R14656 gnd.n6541 gnd.n6540 0.152939
R14657 gnd.n6542 gnd.n6541 0.152939
R14658 gnd.n6543 gnd.n6542 0.152939
R14659 gnd.n6543 gnd.n5903 0.152939
R14660 gnd.n6571 gnd.n5903 0.152939
R14661 gnd.n6572 gnd.n6571 0.152939
R14662 gnd.n6573 gnd.n6572 0.152939
R14663 gnd.n6574 gnd.n6573 0.152939
R14664 gnd.n6574 gnd.n5878 0.152939
R14665 gnd.n6602 gnd.n5878 0.152939
R14666 gnd.n6603 gnd.n6602 0.152939
R14667 gnd.n6604 gnd.n6603 0.152939
R14668 gnd.n6605 gnd.n6604 0.152939
R14669 gnd.n6605 gnd.n5854 0.152939
R14670 gnd.n6632 gnd.n5854 0.152939
R14671 gnd.n6633 gnd.n6632 0.152939
R14672 gnd.n6634 gnd.n6633 0.152939
R14673 gnd.n6635 gnd.n6634 0.152939
R14674 gnd.n6635 gnd.n5822 0.152939
R14675 gnd.n6673 gnd.n5822 0.152939
R14676 gnd.n6674 gnd.n6673 0.152939
R14677 gnd.n6675 gnd.n6674 0.152939
R14678 gnd.n6676 gnd.n6675 0.152939
R14679 gnd.n6677 gnd.n6676 0.152939
R14680 gnd.n6677 gnd.n5792 0.152939
R14681 gnd.n6720 gnd.n5792 0.152939
R14682 gnd.n6721 gnd.n6720 0.152939
R14683 gnd.n6722 gnd.n6721 0.152939
R14684 gnd.n6723 gnd.n6722 0.152939
R14685 gnd.n6724 gnd.n6723 0.152939
R14686 gnd.n6724 gnd.n5765 0.152939
R14687 gnd.n6764 gnd.n5765 0.152939
R14688 gnd.n6765 gnd.n6764 0.152939
R14689 gnd.n6766 gnd.n6765 0.152939
R14690 gnd.n6767 gnd.n6766 0.152939
R14691 gnd.n6767 gnd.n5405 0.152939
R14692 gnd.n6872 gnd.n5405 0.152939
R14693 gnd.n6373 gnd.n6372 0.152939
R14694 gnd.n6374 gnd.n6373 0.152939
R14695 gnd.n6375 gnd.n6374 0.152939
R14696 gnd.n6376 gnd.n6375 0.152939
R14697 gnd.n6377 gnd.n6376 0.152939
R14698 gnd.n6378 gnd.n6377 0.152939
R14699 gnd.n6379 gnd.n6378 0.152939
R14700 gnd.n6380 gnd.n6379 0.152939
R14701 gnd.n6381 gnd.n6380 0.152939
R14702 gnd.n6382 gnd.n6381 0.152939
R14703 gnd.n6383 gnd.n6382 0.152939
R14704 gnd.n6384 gnd.n6383 0.152939
R14705 gnd.n6385 gnd.n6384 0.152939
R14706 gnd.n6386 gnd.n6385 0.152939
R14707 gnd.n6390 gnd.n6386 0.152939
R14708 gnd.n6390 gnd.n6023 0.152939
R14709 gnd.n6839 gnd.n5436 0.152939
R14710 gnd.n5438 gnd.n5436 0.152939
R14711 gnd.n5442 gnd.n5438 0.152939
R14712 gnd.n5443 gnd.n5442 0.152939
R14713 gnd.n5444 gnd.n5443 0.152939
R14714 gnd.n5445 gnd.n5444 0.152939
R14715 gnd.n5449 gnd.n5445 0.152939
R14716 gnd.n5450 gnd.n5449 0.152939
R14717 gnd.n5451 gnd.n5450 0.152939
R14718 gnd.n5452 gnd.n5451 0.152939
R14719 gnd.n5456 gnd.n5452 0.152939
R14720 gnd.n5457 gnd.n5456 0.152939
R14721 gnd.n5458 gnd.n5457 0.152939
R14722 gnd.n5459 gnd.n5458 0.152939
R14723 gnd.n5463 gnd.n5459 0.152939
R14724 gnd.n5464 gnd.n5463 0.152939
R14725 gnd.n5465 gnd.n5464 0.152939
R14726 gnd.n5466 gnd.n5465 0.152939
R14727 gnd.n5470 gnd.n5466 0.152939
R14728 gnd.n5471 gnd.n5470 0.152939
R14729 gnd.n5472 gnd.n5471 0.152939
R14730 gnd.n5473 gnd.n5472 0.152939
R14731 gnd.n5480 gnd.n5473 0.152939
R14732 gnd.n5481 gnd.n5480 0.152939
R14733 gnd.n5482 gnd.n5481 0.152939
R14734 gnd.n6791 gnd.n5482 0.152939
R14735 gnd.n6215 gnd.n6213 0.152939
R14736 gnd.n6216 gnd.n6215 0.152939
R14737 gnd.n6217 gnd.n6216 0.152939
R14738 gnd.n6218 gnd.n6217 0.152939
R14739 gnd.n6219 gnd.n6218 0.152939
R14740 gnd.n6220 gnd.n6219 0.152939
R14741 gnd.n6221 gnd.n6220 0.152939
R14742 gnd.n6221 gnd.n5840 0.152939
R14743 gnd.n6652 gnd.n5840 0.152939
R14744 gnd.n6653 gnd.n6652 0.152939
R14745 gnd.n6654 gnd.n6653 0.152939
R14746 gnd.n6655 gnd.n6654 0.152939
R14747 gnd.n6655 gnd.n5805 0.152939
R14748 gnd.n6696 gnd.n5805 0.152939
R14749 gnd.n6697 gnd.n6696 0.152939
R14750 gnd.n6698 gnd.n6697 0.152939
R14751 gnd.n6699 gnd.n6698 0.152939
R14752 gnd.n6699 gnd.n5778 0.152939
R14753 gnd.n6741 gnd.n5778 0.152939
R14754 gnd.n6742 gnd.n6741 0.152939
R14755 gnd.n6743 gnd.n6742 0.152939
R14756 gnd.n6744 gnd.n6743 0.152939
R14757 gnd.n6744 gnd.n5485 0.152939
R14758 gnd.n6782 gnd.n5485 0.152939
R14759 gnd.n6783 gnd.n6782 0.152939
R14760 gnd.n6784 gnd.n6783 0.152939
R14761 gnd.n6784 gnd.n5483 0.152939
R14762 gnd.n6790 gnd.n5483 0.152939
R14763 gnd.n6160 gnd.n6159 0.152939
R14764 gnd.n6161 gnd.n6160 0.152939
R14765 gnd.n6161 gnd.n6043 0.152939
R14766 gnd.n6175 gnd.n6043 0.152939
R14767 gnd.n6176 gnd.n6175 0.152939
R14768 gnd.n6177 gnd.n6176 0.152939
R14769 gnd.n6177 gnd.n6030 0.152939
R14770 gnd.n6191 gnd.n6030 0.152939
R14771 gnd.n6192 gnd.n6191 0.152939
R14772 gnd.n6193 gnd.n6192 0.152939
R14773 gnd.n6194 gnd.n6193 0.152939
R14774 gnd.n6195 gnd.n6194 0.152939
R14775 gnd.n6196 gnd.n6195 0.152939
R14776 gnd.n6197 gnd.n6196 0.152939
R14777 gnd.n6198 gnd.n6197 0.152939
R14778 gnd.n6199 gnd.n6198 0.152939
R14779 gnd.n6200 gnd.n6199 0.152939
R14780 gnd.n6201 gnd.n6200 0.152939
R14781 gnd.n6202 gnd.n6201 0.152939
R14782 gnd.n6203 gnd.n6202 0.152939
R14783 gnd.n6204 gnd.n6203 0.152939
R14784 gnd.n6205 gnd.n6204 0.152939
R14785 gnd.n6206 gnd.n6205 0.152939
R14786 gnd.n6207 gnd.n6206 0.152939
R14787 gnd.n6208 gnd.n6207 0.152939
R14788 gnd.n6209 gnd.n6208 0.152939
R14789 gnd.n6210 gnd.n6209 0.152939
R14790 gnd.n6211 gnd.n6210 0.152939
R14791 gnd.n6152 gnd.n6059 0.152939
R14792 gnd.n6062 gnd.n6059 0.152939
R14793 gnd.n6063 gnd.n6062 0.152939
R14794 gnd.n6064 gnd.n6063 0.152939
R14795 gnd.n6067 gnd.n6064 0.152939
R14796 gnd.n6068 gnd.n6067 0.152939
R14797 gnd.n6069 gnd.n6068 0.152939
R14798 gnd.n6070 gnd.n6069 0.152939
R14799 gnd.n6073 gnd.n6070 0.152939
R14800 gnd.n6074 gnd.n6073 0.152939
R14801 gnd.n6075 gnd.n6074 0.152939
R14802 gnd.n6076 gnd.n6075 0.152939
R14803 gnd.n6079 gnd.n6076 0.152939
R14804 gnd.n6080 gnd.n6079 0.152939
R14805 gnd.n6081 gnd.n6080 0.152939
R14806 gnd.n6082 gnd.n6081 0.152939
R14807 gnd.n6085 gnd.n6082 0.152939
R14808 gnd.n6086 gnd.n6085 0.152939
R14809 gnd.n6087 gnd.n6086 0.152939
R14810 gnd.n6088 gnd.n6087 0.152939
R14811 gnd.n6091 gnd.n6088 0.152939
R14812 gnd.n6092 gnd.n6091 0.152939
R14813 gnd.n6095 gnd.n6092 0.152939
R14814 gnd.n6096 gnd.n6095 0.152939
R14815 gnd.n6098 gnd.n6096 0.152939
R14816 gnd.n6098 gnd.n6055 0.152939
R14817 gnd.n7056 gnd.n7055 0.152939
R14818 gnd.n7057 gnd.n7056 0.152939
R14819 gnd.n7057 gnd.n960 0.152939
R14820 gnd.n7065 gnd.n960 0.152939
R14821 gnd.n7066 gnd.n7065 0.152939
R14822 gnd.n7067 gnd.n7066 0.152939
R14823 gnd.n7067 gnd.n954 0.152939
R14824 gnd.n7075 gnd.n954 0.152939
R14825 gnd.n7076 gnd.n7075 0.152939
R14826 gnd.n7077 gnd.n7076 0.152939
R14827 gnd.n7077 gnd.n948 0.152939
R14828 gnd.n7085 gnd.n948 0.152939
R14829 gnd.n7086 gnd.n7085 0.152939
R14830 gnd.n7087 gnd.n7086 0.152939
R14831 gnd.n7087 gnd.n942 0.152939
R14832 gnd.n7095 gnd.n942 0.152939
R14833 gnd.n7096 gnd.n7095 0.152939
R14834 gnd.n7097 gnd.n7096 0.152939
R14835 gnd.n7097 gnd.n936 0.152939
R14836 gnd.n7105 gnd.n936 0.152939
R14837 gnd.n7106 gnd.n7105 0.152939
R14838 gnd.n7107 gnd.n7106 0.152939
R14839 gnd.n7107 gnd.n930 0.152939
R14840 gnd.n7115 gnd.n930 0.152939
R14841 gnd.n7116 gnd.n7115 0.152939
R14842 gnd.n7117 gnd.n7116 0.152939
R14843 gnd.n7117 gnd.n924 0.152939
R14844 gnd.n7125 gnd.n924 0.152939
R14845 gnd.n7126 gnd.n7125 0.152939
R14846 gnd.n7127 gnd.n7126 0.152939
R14847 gnd.n7127 gnd.n918 0.152939
R14848 gnd.n7135 gnd.n918 0.152939
R14849 gnd.n7136 gnd.n7135 0.152939
R14850 gnd.n7137 gnd.n7136 0.152939
R14851 gnd.n7137 gnd.n912 0.152939
R14852 gnd.n7145 gnd.n912 0.152939
R14853 gnd.n7146 gnd.n7145 0.152939
R14854 gnd.n7147 gnd.n7146 0.152939
R14855 gnd.n7147 gnd.n906 0.152939
R14856 gnd.n7155 gnd.n906 0.152939
R14857 gnd.n7156 gnd.n7155 0.152939
R14858 gnd.n7157 gnd.n7156 0.152939
R14859 gnd.n7157 gnd.n900 0.152939
R14860 gnd.n7165 gnd.n900 0.152939
R14861 gnd.n7166 gnd.n7165 0.152939
R14862 gnd.n7167 gnd.n7166 0.152939
R14863 gnd.n7167 gnd.n894 0.152939
R14864 gnd.n7175 gnd.n894 0.152939
R14865 gnd.n7176 gnd.n7175 0.152939
R14866 gnd.n7177 gnd.n7176 0.152939
R14867 gnd.n7177 gnd.n888 0.152939
R14868 gnd.n7185 gnd.n888 0.152939
R14869 gnd.n7186 gnd.n7185 0.152939
R14870 gnd.n7187 gnd.n7186 0.152939
R14871 gnd.n7187 gnd.n882 0.152939
R14872 gnd.n7195 gnd.n882 0.152939
R14873 gnd.n7196 gnd.n7195 0.152939
R14874 gnd.n7197 gnd.n7196 0.152939
R14875 gnd.n7197 gnd.n876 0.152939
R14876 gnd.n7205 gnd.n876 0.152939
R14877 gnd.n7206 gnd.n7205 0.152939
R14878 gnd.n7207 gnd.n7206 0.152939
R14879 gnd.n7207 gnd.n870 0.152939
R14880 gnd.n7215 gnd.n870 0.152939
R14881 gnd.n7216 gnd.n7215 0.152939
R14882 gnd.n7217 gnd.n7216 0.152939
R14883 gnd.n7217 gnd.n864 0.152939
R14884 gnd.n7225 gnd.n864 0.152939
R14885 gnd.n7226 gnd.n7225 0.152939
R14886 gnd.n7227 gnd.n7226 0.152939
R14887 gnd.n7227 gnd.n858 0.152939
R14888 gnd.n7235 gnd.n858 0.152939
R14889 gnd.n7236 gnd.n7235 0.152939
R14890 gnd.n7237 gnd.n7236 0.152939
R14891 gnd.n7237 gnd.n852 0.152939
R14892 gnd.n7245 gnd.n852 0.152939
R14893 gnd.n7246 gnd.n7245 0.152939
R14894 gnd.n7247 gnd.n7246 0.152939
R14895 gnd.n7247 gnd.n846 0.152939
R14896 gnd.n7255 gnd.n846 0.152939
R14897 gnd.n7256 gnd.n7255 0.152939
R14898 gnd.n7257 gnd.n7256 0.152939
R14899 gnd.n7257 gnd.n840 0.152939
R14900 gnd.n7265 gnd.n840 0.152939
R14901 gnd.n7266 gnd.n7265 0.152939
R14902 gnd.n7267 gnd.n7266 0.152939
R14903 gnd.n7267 gnd.n834 0.152939
R14904 gnd.n7275 gnd.n834 0.152939
R14905 gnd.n7276 gnd.n7275 0.152939
R14906 gnd.n7277 gnd.n7276 0.152939
R14907 gnd.n7277 gnd.n828 0.152939
R14908 gnd.n7285 gnd.n828 0.152939
R14909 gnd.n7286 gnd.n7285 0.152939
R14910 gnd.n7287 gnd.n7286 0.152939
R14911 gnd.n7287 gnd.n822 0.152939
R14912 gnd.n7295 gnd.n822 0.152939
R14913 gnd.n7296 gnd.n7295 0.152939
R14914 gnd.n7297 gnd.n7296 0.152939
R14915 gnd.n7297 gnd.n816 0.152939
R14916 gnd.n7305 gnd.n816 0.152939
R14917 gnd.n7306 gnd.n7305 0.152939
R14918 gnd.n7307 gnd.n7306 0.152939
R14919 gnd.n7307 gnd.n810 0.152939
R14920 gnd.n7315 gnd.n810 0.152939
R14921 gnd.n7316 gnd.n7315 0.152939
R14922 gnd.n7317 gnd.n7316 0.152939
R14923 gnd.n7317 gnd.n804 0.152939
R14924 gnd.n7325 gnd.n804 0.152939
R14925 gnd.n7326 gnd.n7325 0.152939
R14926 gnd.n7327 gnd.n7326 0.152939
R14927 gnd.n7327 gnd.n798 0.152939
R14928 gnd.n7335 gnd.n798 0.152939
R14929 gnd.n7336 gnd.n7335 0.152939
R14930 gnd.n7337 gnd.n7336 0.152939
R14931 gnd.n7337 gnd.n792 0.152939
R14932 gnd.n7345 gnd.n792 0.152939
R14933 gnd.n7346 gnd.n7345 0.152939
R14934 gnd.n7347 gnd.n7346 0.152939
R14935 gnd.n7347 gnd.n786 0.152939
R14936 gnd.n7355 gnd.n786 0.152939
R14937 gnd.n7356 gnd.n7355 0.152939
R14938 gnd.n7357 gnd.n7356 0.152939
R14939 gnd.n7357 gnd.n780 0.152939
R14940 gnd.n7365 gnd.n780 0.152939
R14941 gnd.n7366 gnd.n7365 0.152939
R14942 gnd.n7367 gnd.n7366 0.152939
R14943 gnd.n7367 gnd.n774 0.152939
R14944 gnd.n7375 gnd.n774 0.152939
R14945 gnd.n7376 gnd.n7375 0.152939
R14946 gnd.n7377 gnd.n7376 0.152939
R14947 gnd.n7377 gnd.n768 0.152939
R14948 gnd.n7385 gnd.n768 0.152939
R14949 gnd.n7386 gnd.n7385 0.152939
R14950 gnd.n7387 gnd.n7386 0.152939
R14951 gnd.n7387 gnd.n762 0.152939
R14952 gnd.n7395 gnd.n762 0.152939
R14953 gnd.n7396 gnd.n7395 0.152939
R14954 gnd.n7397 gnd.n7396 0.152939
R14955 gnd.n7397 gnd.n756 0.152939
R14956 gnd.n7405 gnd.n756 0.152939
R14957 gnd.n7406 gnd.n7405 0.152939
R14958 gnd.n7407 gnd.n7406 0.152939
R14959 gnd.n7407 gnd.n750 0.152939
R14960 gnd.n7415 gnd.n750 0.152939
R14961 gnd.n7416 gnd.n7415 0.152939
R14962 gnd.n7417 gnd.n7416 0.152939
R14963 gnd.n7417 gnd.n744 0.152939
R14964 gnd.n7425 gnd.n744 0.152939
R14965 gnd.n7426 gnd.n7425 0.152939
R14966 gnd.n7427 gnd.n7426 0.152939
R14967 gnd.n7427 gnd.n738 0.152939
R14968 gnd.n7435 gnd.n738 0.152939
R14969 gnd.n7436 gnd.n7435 0.152939
R14970 gnd.n7437 gnd.n7436 0.152939
R14971 gnd.n7437 gnd.n732 0.152939
R14972 gnd.n7445 gnd.n732 0.152939
R14973 gnd.n7446 gnd.n7445 0.152939
R14974 gnd.n7447 gnd.n7446 0.152939
R14975 gnd.n7447 gnd.n726 0.152939
R14976 gnd.n7455 gnd.n726 0.152939
R14977 gnd.n7456 gnd.n7455 0.152939
R14978 gnd.n7457 gnd.n7456 0.152939
R14979 gnd.n7457 gnd.n720 0.152939
R14980 gnd.n7465 gnd.n720 0.152939
R14981 gnd.n7466 gnd.n7465 0.152939
R14982 gnd.n7467 gnd.n7466 0.152939
R14983 gnd.n7467 gnd.n714 0.152939
R14984 gnd.n7475 gnd.n714 0.152939
R14985 gnd.n7476 gnd.n7475 0.152939
R14986 gnd.n7477 gnd.n7476 0.152939
R14987 gnd.n7477 gnd.n708 0.152939
R14988 gnd.n7485 gnd.n708 0.152939
R14989 gnd.n7486 gnd.n7485 0.152939
R14990 gnd.n7487 gnd.n7486 0.152939
R14991 gnd.n7487 gnd.n702 0.152939
R14992 gnd.n7495 gnd.n702 0.152939
R14993 gnd.n7496 gnd.n7495 0.152939
R14994 gnd.n7498 gnd.n7496 0.152939
R14995 gnd.n7498 gnd.n7497 0.152939
R14996 gnd.n7497 gnd.n696 0.152939
R14997 gnd.n7507 gnd.n696 0.152939
R14998 gnd.n7508 gnd.n691 0.152939
R14999 gnd.n7516 gnd.n691 0.152939
R15000 gnd.n7517 gnd.n7516 0.152939
R15001 gnd.n7518 gnd.n7517 0.152939
R15002 gnd.n7518 gnd.n685 0.152939
R15003 gnd.n7526 gnd.n685 0.152939
R15004 gnd.n7527 gnd.n7526 0.152939
R15005 gnd.n7528 gnd.n7527 0.152939
R15006 gnd.n7528 gnd.n679 0.152939
R15007 gnd.n7536 gnd.n679 0.152939
R15008 gnd.n7537 gnd.n7536 0.152939
R15009 gnd.n7538 gnd.n7537 0.152939
R15010 gnd.n7538 gnd.n673 0.152939
R15011 gnd.n7546 gnd.n673 0.152939
R15012 gnd.n7547 gnd.n7546 0.152939
R15013 gnd.n7548 gnd.n7547 0.152939
R15014 gnd.n7548 gnd.n667 0.152939
R15015 gnd.n7556 gnd.n667 0.152939
R15016 gnd.n7557 gnd.n7556 0.152939
R15017 gnd.n7558 gnd.n7557 0.152939
R15018 gnd.n7558 gnd.n661 0.152939
R15019 gnd.n7566 gnd.n661 0.152939
R15020 gnd.n7567 gnd.n7566 0.152939
R15021 gnd.n7568 gnd.n7567 0.152939
R15022 gnd.n7568 gnd.n655 0.152939
R15023 gnd.n7576 gnd.n655 0.152939
R15024 gnd.n7577 gnd.n7576 0.152939
R15025 gnd.n7578 gnd.n7577 0.152939
R15026 gnd.n7578 gnd.n649 0.152939
R15027 gnd.n7586 gnd.n649 0.152939
R15028 gnd.n7587 gnd.n7586 0.152939
R15029 gnd.n7588 gnd.n7587 0.152939
R15030 gnd.n7588 gnd.n643 0.152939
R15031 gnd.n7596 gnd.n643 0.152939
R15032 gnd.n7597 gnd.n7596 0.152939
R15033 gnd.n7598 gnd.n7597 0.152939
R15034 gnd.n7598 gnd.n637 0.152939
R15035 gnd.n7606 gnd.n637 0.152939
R15036 gnd.n7607 gnd.n7606 0.152939
R15037 gnd.n7608 gnd.n7607 0.152939
R15038 gnd.n7608 gnd.n631 0.152939
R15039 gnd.n7616 gnd.n631 0.152939
R15040 gnd.n7617 gnd.n7616 0.152939
R15041 gnd.n7618 gnd.n7617 0.152939
R15042 gnd.n7618 gnd.n625 0.152939
R15043 gnd.n7626 gnd.n625 0.152939
R15044 gnd.n7627 gnd.n7626 0.152939
R15045 gnd.n7628 gnd.n7627 0.152939
R15046 gnd.n7628 gnd.n619 0.152939
R15047 gnd.n7636 gnd.n619 0.152939
R15048 gnd.n7637 gnd.n7636 0.152939
R15049 gnd.n7638 gnd.n7637 0.152939
R15050 gnd.n7638 gnd.n613 0.152939
R15051 gnd.n7646 gnd.n613 0.152939
R15052 gnd.n7647 gnd.n7646 0.152939
R15053 gnd.n7648 gnd.n7647 0.152939
R15054 gnd.n7648 gnd.n607 0.152939
R15055 gnd.n7656 gnd.n607 0.152939
R15056 gnd.n7657 gnd.n7656 0.152939
R15057 gnd.n7658 gnd.n7657 0.152939
R15058 gnd.n7658 gnd.n601 0.152939
R15059 gnd.n7666 gnd.n601 0.152939
R15060 gnd.n7667 gnd.n7666 0.152939
R15061 gnd.n7668 gnd.n7667 0.152939
R15062 gnd.n7668 gnd.n595 0.152939
R15063 gnd.n7676 gnd.n595 0.152939
R15064 gnd.n7677 gnd.n7676 0.152939
R15065 gnd.n7678 gnd.n7677 0.152939
R15066 gnd.n7678 gnd.n589 0.152939
R15067 gnd.n7686 gnd.n589 0.152939
R15068 gnd.n7687 gnd.n7686 0.152939
R15069 gnd.n7688 gnd.n7687 0.152939
R15070 gnd.n7688 gnd.n583 0.152939
R15071 gnd.n7696 gnd.n583 0.152939
R15072 gnd.n7697 gnd.n7696 0.152939
R15073 gnd.n7698 gnd.n7697 0.152939
R15074 gnd.n7698 gnd.n577 0.152939
R15075 gnd.n7706 gnd.n577 0.152939
R15076 gnd.n7707 gnd.n7706 0.152939
R15077 gnd.n7708 gnd.n7707 0.152939
R15078 gnd.n7708 gnd.n571 0.152939
R15079 gnd.n7717 gnd.n571 0.152939
R15080 gnd.n7718 gnd.n7717 0.152939
R15081 gnd.n7719 gnd.n7718 0.152939
R15082 gnd.n8092 gnd.n113 0.152939
R15083 gnd.n138 gnd.n113 0.152939
R15084 gnd.n139 gnd.n138 0.152939
R15085 gnd.n140 gnd.n139 0.152939
R15086 gnd.n155 gnd.n140 0.152939
R15087 gnd.n156 gnd.n155 0.152939
R15088 gnd.n157 gnd.n156 0.152939
R15089 gnd.n158 gnd.n157 0.152939
R15090 gnd.n175 gnd.n158 0.152939
R15091 gnd.n176 gnd.n175 0.152939
R15092 gnd.n177 gnd.n176 0.152939
R15093 gnd.n178 gnd.n177 0.152939
R15094 gnd.n193 gnd.n178 0.152939
R15095 gnd.n194 gnd.n193 0.152939
R15096 gnd.n195 gnd.n194 0.152939
R15097 gnd.n196 gnd.n195 0.152939
R15098 gnd.n213 gnd.n196 0.152939
R15099 gnd.n214 gnd.n213 0.152939
R15100 gnd.n215 gnd.n214 0.152939
R15101 gnd.n216 gnd.n215 0.152939
R15102 gnd.n233 gnd.n216 0.152939
R15103 gnd.n234 gnd.n233 0.152939
R15104 gnd.n235 gnd.n234 0.152939
R15105 gnd.n236 gnd.n235 0.152939
R15106 gnd.n252 gnd.n236 0.152939
R15107 gnd.n253 gnd.n252 0.152939
R15108 gnd.n8007 gnd.n253 0.152939
R15109 gnd.n8101 gnd.n101 0.152939
R15110 gnd.n388 gnd.n101 0.152939
R15111 gnd.n391 gnd.n388 0.152939
R15112 gnd.n392 gnd.n391 0.152939
R15113 gnd.n393 gnd.n392 0.152939
R15114 gnd.n393 gnd.n386 0.152939
R15115 gnd.n399 gnd.n386 0.152939
R15116 gnd.n400 gnd.n399 0.152939
R15117 gnd.n401 gnd.n400 0.152939
R15118 gnd.n401 gnd.n384 0.152939
R15119 gnd.n407 gnd.n384 0.152939
R15120 gnd.n408 gnd.n407 0.152939
R15121 gnd.n409 gnd.n408 0.152939
R15122 gnd.n409 gnd.n382 0.152939
R15123 gnd.n415 gnd.n382 0.152939
R15124 gnd.n416 gnd.n415 0.152939
R15125 gnd.n417 gnd.n416 0.152939
R15126 gnd.n417 gnd.n380 0.152939
R15127 gnd.n423 gnd.n380 0.152939
R15128 gnd.n424 gnd.n423 0.152939
R15129 gnd.n425 gnd.n424 0.152939
R15130 gnd.n425 gnd.n378 0.152939
R15131 gnd.n431 gnd.n378 0.152939
R15132 gnd.n432 gnd.n431 0.152939
R15133 gnd.n433 gnd.n432 0.152939
R15134 gnd.n433 gnd.n376 0.152939
R15135 gnd.n439 gnd.n376 0.152939
R15136 gnd.n440 gnd.n439 0.152939
R15137 gnd.n441 gnd.n440 0.152939
R15138 gnd.n441 gnd.n374 0.152939
R15139 gnd.n448 gnd.n374 0.152939
R15140 gnd.n485 gnd.n354 0.152939
R15141 gnd.n356 gnd.n354 0.152939
R15142 gnd.n357 gnd.n356 0.152939
R15143 gnd.n358 gnd.n357 0.152939
R15144 gnd.n359 gnd.n358 0.152939
R15145 gnd.n360 gnd.n359 0.152939
R15146 gnd.n361 gnd.n360 0.152939
R15147 gnd.n362 gnd.n361 0.152939
R15148 gnd.n363 gnd.n362 0.152939
R15149 gnd.n364 gnd.n363 0.152939
R15150 gnd.n365 gnd.n364 0.152939
R15151 gnd.n366 gnd.n365 0.152939
R15152 gnd.n367 gnd.n366 0.152939
R15153 gnd.n368 gnd.n367 0.152939
R15154 gnd.n369 gnd.n368 0.152939
R15155 gnd.n370 gnd.n369 0.152939
R15156 gnd.n450 gnd.n370 0.152939
R15157 gnd.n450 gnd.n449 0.152939
R15158 gnd.n8006 gnd.n254 0.152939
R15159 gnd.n296 gnd.n254 0.152939
R15160 gnd.n297 gnd.n296 0.152939
R15161 gnd.n298 gnd.n297 0.152939
R15162 gnd.n299 gnd.n298 0.152939
R15163 gnd.n300 gnd.n299 0.152939
R15164 gnd.n301 gnd.n300 0.152939
R15165 gnd.n302 gnd.n301 0.152939
R15166 gnd.n303 gnd.n302 0.152939
R15167 gnd.n304 gnd.n303 0.152939
R15168 gnd.n305 gnd.n304 0.152939
R15169 gnd.n306 gnd.n305 0.152939
R15170 gnd.n307 gnd.n306 0.152939
R15171 gnd.n308 gnd.n307 0.152939
R15172 gnd.n309 gnd.n308 0.152939
R15173 gnd.n310 gnd.n309 0.152939
R15174 gnd.n311 gnd.n310 0.152939
R15175 gnd.n312 gnd.n311 0.152939
R15176 gnd.n313 gnd.n312 0.152939
R15177 gnd.n314 gnd.n313 0.152939
R15178 gnd.n315 gnd.n314 0.152939
R15179 gnd.n316 gnd.n315 0.152939
R15180 gnd.n317 gnd.n316 0.152939
R15181 gnd.n318 gnd.n317 0.152939
R15182 gnd.n319 gnd.n318 0.152939
R15183 gnd.n320 gnd.n319 0.152939
R15184 gnd.n321 gnd.n320 0.152939
R15185 gnd.n322 gnd.n321 0.152939
R15186 gnd.n323 gnd.n322 0.152939
R15187 gnd.n324 gnd.n323 0.152939
R15188 gnd.n325 gnd.n324 0.152939
R15189 gnd.n326 gnd.n325 0.152939
R15190 gnd.n327 gnd.n326 0.152939
R15191 gnd.n328 gnd.n327 0.152939
R15192 gnd.n329 gnd.n328 0.152939
R15193 gnd.n330 gnd.n329 0.152939
R15194 gnd.n7927 gnd.n330 0.152939
R15195 gnd.n7927 gnd.n7926 0.152939
R15196 gnd.n7926 gnd.n7925 0.152939
R15197 gnd.n7925 gnd.n334 0.152939
R15198 gnd.n335 gnd.n334 0.152939
R15199 gnd.n336 gnd.n335 0.152939
R15200 gnd.n337 gnd.n336 0.152939
R15201 gnd.n338 gnd.n337 0.152939
R15202 gnd.n339 gnd.n338 0.152939
R15203 gnd.n340 gnd.n339 0.152939
R15204 gnd.n341 gnd.n340 0.152939
R15205 gnd.n342 gnd.n341 0.152939
R15206 gnd.n343 gnd.n342 0.152939
R15207 gnd.n344 gnd.n343 0.152939
R15208 gnd.n345 gnd.n344 0.152939
R15209 gnd.n346 gnd.n345 0.152939
R15210 gnd.n347 gnd.n346 0.152939
R15211 gnd.n348 gnd.n347 0.152939
R15212 gnd.n349 gnd.n348 0.152939
R15213 gnd.n350 gnd.n349 0.152939
R15214 gnd.n7885 gnd.n350 0.152939
R15215 gnd.n7885 gnd.n7884 0.152939
R15216 gnd.n1864 gnd.n1863 0.152939
R15217 gnd.n1865 gnd.n1864 0.152939
R15218 gnd.n1866 gnd.n1865 0.152939
R15219 gnd.n1867 gnd.n1866 0.152939
R15220 gnd.n1868 gnd.n1867 0.152939
R15221 gnd.n1869 gnd.n1868 0.152939
R15222 gnd.n1870 gnd.n1869 0.152939
R15223 gnd.n1871 gnd.n1870 0.152939
R15224 gnd.n1872 gnd.n1871 0.152939
R15225 gnd.n1873 gnd.n1872 0.152939
R15226 gnd.n1874 gnd.n1873 0.152939
R15227 gnd.n1875 gnd.n1874 0.152939
R15228 gnd.n1876 gnd.n1875 0.152939
R15229 gnd.n1877 gnd.n1876 0.152939
R15230 gnd.n1878 gnd.n1877 0.152939
R15231 gnd.n1879 gnd.n1878 0.152939
R15232 gnd.n1880 gnd.n1879 0.152939
R15233 gnd.n1883 gnd.n1880 0.152939
R15234 gnd.n1884 gnd.n1883 0.152939
R15235 gnd.n1885 gnd.n1884 0.152939
R15236 gnd.n1886 gnd.n1885 0.152939
R15237 gnd.n1887 gnd.n1886 0.152939
R15238 gnd.n1888 gnd.n1887 0.152939
R15239 gnd.n1889 gnd.n1888 0.152939
R15240 gnd.n1890 gnd.n1889 0.152939
R15241 gnd.n1895 gnd.n1894 0.152939
R15242 gnd.n1896 gnd.n1895 0.152939
R15243 gnd.n1897 gnd.n1896 0.152939
R15244 gnd.n1898 gnd.n1897 0.152939
R15245 gnd.n1899 gnd.n1898 0.152939
R15246 gnd.n1900 gnd.n1899 0.152939
R15247 gnd.n1901 gnd.n1900 0.152939
R15248 gnd.n1902 gnd.n1901 0.152939
R15249 gnd.n1903 gnd.n1902 0.152939
R15250 gnd.n1906 gnd.n1903 0.152939
R15251 gnd.n1907 gnd.n1906 0.152939
R15252 gnd.n1908 gnd.n1907 0.152939
R15253 gnd.n1909 gnd.n1908 0.152939
R15254 gnd.n1910 gnd.n1909 0.152939
R15255 gnd.n1911 gnd.n1910 0.152939
R15256 gnd.n1912 gnd.n1911 0.152939
R15257 gnd.n1913 gnd.n1912 0.152939
R15258 gnd.n1914 gnd.n1913 0.152939
R15259 gnd.n1915 gnd.n1914 0.152939
R15260 gnd.n1916 gnd.n1915 0.152939
R15261 gnd.n1917 gnd.n1916 0.152939
R15262 gnd.n1918 gnd.n1917 0.152939
R15263 gnd.n1919 gnd.n1918 0.152939
R15264 gnd.n1920 gnd.n1919 0.152939
R15265 gnd.n1921 gnd.n1920 0.152939
R15266 gnd.n1922 gnd.n1921 0.152939
R15267 gnd.n1923 gnd.n1922 0.152939
R15268 gnd.n1924 gnd.n1923 0.152939
R15269 gnd.n4722 gnd.n1924 0.152939
R15270 gnd.n4722 gnd.n4721 0.152939
R15271 gnd.n1945 gnd.n1944 0.152939
R15272 gnd.n1946 gnd.n1945 0.152939
R15273 gnd.n1947 gnd.n1946 0.152939
R15274 gnd.n1966 gnd.n1947 0.152939
R15275 gnd.n1967 gnd.n1966 0.152939
R15276 gnd.n1968 gnd.n1967 0.152939
R15277 gnd.n1969 gnd.n1968 0.152939
R15278 gnd.n1986 gnd.n1969 0.152939
R15279 gnd.n1987 gnd.n1986 0.152939
R15280 gnd.n1988 gnd.n1987 0.152939
R15281 gnd.n1989 gnd.n1988 0.152939
R15282 gnd.n2007 gnd.n1989 0.152939
R15283 gnd.n2008 gnd.n2007 0.152939
R15284 gnd.n2009 gnd.n2008 0.152939
R15285 gnd.n2010 gnd.n2009 0.152939
R15286 gnd.n2027 gnd.n2010 0.152939
R15287 gnd.n2028 gnd.n2027 0.152939
R15288 gnd.n2029 gnd.n2028 0.152939
R15289 gnd.n2030 gnd.n2029 0.152939
R15290 gnd.n2031 gnd.n2030 0.152939
R15291 gnd.n2031 gnd.n539 0.152939
R15292 gnd.n7760 gnd.n539 0.152939
R15293 gnd.n7761 gnd.n7760 0.152939
R15294 gnd.n7762 gnd.n7761 0.152939
R15295 gnd.n7763 gnd.n7762 0.152939
R15296 gnd.n7763 gnd.n114 0.152939
R15297 gnd.n8092 gnd.n114 0.152939
R15298 gnd.n7733 gnd.n560 0.152939
R15299 gnd.n7733 gnd.n7732 0.152939
R15300 gnd.n7732 gnd.n7731 0.152939
R15301 gnd.n7731 gnd.n562 0.152939
R15302 gnd.n567 gnd.n566 0.152939
R15303 gnd.n568 gnd.n567 0.152939
R15304 gnd.n3060 gnd.n3059 0.152939
R15305 gnd.n3061 gnd.n3060 0.152939
R15306 gnd.n3062 gnd.n3061 0.152939
R15307 gnd.n3063 gnd.n3062 0.152939
R15308 gnd.n3066 gnd.n3063 0.152939
R15309 gnd.n3067 gnd.n3066 0.152939
R15310 gnd.n3068 gnd.n3067 0.152939
R15311 gnd.n3069 gnd.n3068 0.152939
R15312 gnd.n3071 gnd.n3069 0.152939
R15313 gnd.n3071 gnd.n3070 0.152939
R15314 gnd.n3070 gnd.n2754 0.152939
R15315 gnd.n3148 gnd.n2754 0.152939
R15316 gnd.n3149 gnd.n3148 0.152939
R15317 gnd.n3150 gnd.n3149 0.152939
R15318 gnd.n3150 gnd.n2750 0.152939
R15319 gnd.n3156 gnd.n2750 0.152939
R15320 gnd.n3157 gnd.n3156 0.152939
R15321 gnd.n3158 gnd.n3157 0.152939
R15322 gnd.n3159 gnd.n3158 0.152939
R15323 gnd.n3160 gnd.n3159 0.152939
R15324 gnd.n3163 gnd.n3160 0.152939
R15325 gnd.n3164 gnd.n3163 0.152939
R15326 gnd.n3165 gnd.n3164 0.152939
R15327 gnd.n3166 gnd.n3165 0.152939
R15328 gnd.n3168 gnd.n3166 0.152939
R15329 gnd.n3170 gnd.n3168 0.152939
R15330 gnd.n3170 gnd.n3169 0.152939
R15331 gnd.n3169 gnd.n2558 0.152939
R15332 gnd.n2559 gnd.n2558 0.152939
R15333 gnd.n2560 gnd.n2559 0.152939
R15334 gnd.n2562 gnd.n2560 0.152939
R15335 gnd.n2563 gnd.n2562 0.152939
R15336 gnd.n2563 gnd.n2539 0.152939
R15337 gnd.n3376 gnd.n2539 0.152939
R15338 gnd.n3377 gnd.n3376 0.152939
R15339 gnd.n3378 gnd.n3377 0.152939
R15340 gnd.n3378 gnd.n2526 0.152939
R15341 gnd.n3392 gnd.n2526 0.152939
R15342 gnd.n3393 gnd.n3392 0.152939
R15343 gnd.n3394 gnd.n3393 0.152939
R15344 gnd.n3394 gnd.n2512 0.152939
R15345 gnd.n3408 gnd.n2512 0.152939
R15346 gnd.n3409 gnd.n3408 0.152939
R15347 gnd.n3410 gnd.n3409 0.152939
R15348 gnd.n3410 gnd.n2498 0.152939
R15349 gnd.n3424 gnd.n2498 0.152939
R15350 gnd.n3425 gnd.n3424 0.152939
R15351 gnd.n3426 gnd.n3425 0.152939
R15352 gnd.n3427 gnd.n3426 0.152939
R15353 gnd.n3428 gnd.n3427 0.152939
R15354 gnd.n3430 gnd.n3428 0.152939
R15355 gnd.n3430 gnd.n3429 0.152939
R15356 gnd.n3429 gnd.n1696 0.152939
R15357 gnd.n1697 gnd.n1696 0.152939
R15358 gnd.n1698 gnd.n1697 0.152939
R15359 gnd.n4087 gnd.n1698 0.152939
R15360 gnd.n4088 gnd.n4087 0.152939
R15361 gnd.n4088 gnd.n2382 0.152939
R15362 gnd.n4102 gnd.n2382 0.152939
R15363 gnd.n4103 gnd.n4102 0.152939
R15364 gnd.n4104 gnd.n4103 0.152939
R15365 gnd.n4104 gnd.n2368 0.152939
R15366 gnd.n4118 gnd.n2368 0.152939
R15367 gnd.n4119 gnd.n4118 0.152939
R15368 gnd.n4120 gnd.n4119 0.152939
R15369 gnd.n4120 gnd.n2356 0.152939
R15370 gnd.n4134 gnd.n2356 0.152939
R15371 gnd.n4135 gnd.n4134 0.152939
R15372 gnd.n4136 gnd.n4135 0.152939
R15373 gnd.n4136 gnd.n2342 0.152939
R15374 gnd.n4150 gnd.n2342 0.152939
R15375 gnd.n4151 gnd.n4150 0.152939
R15376 gnd.n4152 gnd.n4151 0.152939
R15377 gnd.n4152 gnd.n2327 0.152939
R15378 gnd.n4166 gnd.n2327 0.152939
R15379 gnd.n4167 gnd.n4166 0.152939
R15380 gnd.n4168 gnd.n4167 0.152939
R15381 gnd.n4168 gnd.n2313 0.152939
R15382 gnd.n4182 gnd.n2313 0.152939
R15383 gnd.n4183 gnd.n4182 0.152939
R15384 gnd.n4184 gnd.n4183 0.152939
R15385 gnd.n4184 gnd.n2299 0.152939
R15386 gnd.n4198 gnd.n2299 0.152939
R15387 gnd.n4199 gnd.n4198 0.152939
R15388 gnd.n4200 gnd.n4199 0.152939
R15389 gnd.n4200 gnd.n2286 0.152939
R15390 gnd.n4214 gnd.n2286 0.152939
R15391 gnd.n4215 gnd.n4214 0.152939
R15392 gnd.n4216 gnd.n4215 0.152939
R15393 gnd.n4216 gnd.n2272 0.152939
R15394 gnd.n4230 gnd.n2272 0.152939
R15395 gnd.n4231 gnd.n4230 0.152939
R15396 gnd.n4232 gnd.n4231 0.152939
R15397 gnd.n4232 gnd.n2258 0.152939
R15398 gnd.n4246 gnd.n2258 0.152939
R15399 gnd.n4247 gnd.n4246 0.152939
R15400 gnd.n4248 gnd.n4247 0.152939
R15401 gnd.n4248 gnd.n2245 0.152939
R15402 gnd.n4262 gnd.n2245 0.152939
R15403 gnd.n4263 gnd.n4262 0.152939
R15404 gnd.n4264 gnd.n4263 0.152939
R15405 gnd.n4264 gnd.n2231 0.152939
R15406 gnd.n4278 gnd.n2231 0.152939
R15407 gnd.n4279 gnd.n4278 0.152939
R15408 gnd.n4280 gnd.n4279 0.152939
R15409 gnd.n4280 gnd.n2218 0.152939
R15410 gnd.n4294 gnd.n2218 0.152939
R15411 gnd.n4295 gnd.n4294 0.152939
R15412 gnd.n4296 gnd.n4295 0.152939
R15413 gnd.n4296 gnd.n2203 0.152939
R15414 gnd.n4310 gnd.n2203 0.152939
R15415 gnd.n4311 gnd.n4310 0.152939
R15416 gnd.n4312 gnd.n4311 0.152939
R15417 gnd.n4312 gnd.n2190 0.152939
R15418 gnd.n4326 gnd.n2190 0.152939
R15419 gnd.n4327 gnd.n4326 0.152939
R15420 gnd.n4328 gnd.n4327 0.152939
R15421 gnd.n4328 gnd.n2179 0.152939
R15422 gnd.n4342 gnd.n2179 0.152939
R15423 gnd.n4343 gnd.n4342 0.152939
R15424 gnd.n4344 gnd.n4343 0.152939
R15425 gnd.n4344 gnd.n2166 0.152939
R15426 gnd.n4358 gnd.n2166 0.152939
R15427 gnd.n4359 gnd.n4358 0.152939
R15428 gnd.n4360 gnd.n4359 0.152939
R15429 gnd.n4360 gnd.n2151 0.152939
R15430 gnd.n4374 gnd.n2151 0.152939
R15431 gnd.n4375 gnd.n4374 0.152939
R15432 gnd.n4376 gnd.n4375 0.152939
R15433 gnd.n4376 gnd.n2139 0.152939
R15434 gnd.n4392 gnd.n2139 0.152939
R15435 gnd.n4393 gnd.n4392 0.152939
R15436 gnd.n4394 gnd.n4393 0.152939
R15437 gnd.n4396 gnd.n4394 0.152939
R15438 gnd.n4396 gnd.n4395 0.152939
R15439 gnd.n4395 gnd.n1815 0.152939
R15440 gnd.n1816 gnd.n1815 0.152939
R15441 gnd.n1817 gnd.n1816 0.152939
R15442 gnd.n2074 gnd.n1817 0.152939
R15443 gnd.n2075 gnd.n2074 0.152939
R15444 gnd.n2080 gnd.n2075 0.152939
R15445 gnd.n2081 gnd.n2080 0.152939
R15446 gnd.n2082 gnd.n2081 0.152939
R15447 gnd.n2082 gnd.n2070 0.152939
R15448 gnd.n2088 gnd.n2070 0.152939
R15449 gnd.n2089 gnd.n2088 0.152939
R15450 gnd.n2090 gnd.n2089 0.152939
R15451 gnd.n2090 gnd.n2066 0.152939
R15452 gnd.n2096 gnd.n2066 0.152939
R15453 gnd.n2097 gnd.n2096 0.152939
R15454 gnd.n2098 gnd.n2097 0.152939
R15455 gnd.n2099 gnd.n2098 0.152939
R15456 gnd.n2100 gnd.n2099 0.152939
R15457 gnd.n2103 gnd.n2100 0.152939
R15458 gnd.n2104 gnd.n2103 0.152939
R15459 gnd.n2105 gnd.n2104 0.152939
R15460 gnd.n2106 gnd.n2105 0.152939
R15461 gnd.n2107 gnd.n2106 0.152939
R15462 gnd.n2107 gnd.n2048 0.152939
R15463 gnd.n4645 gnd.n2048 0.152939
R15464 gnd.n4646 gnd.n4645 0.152939
R15465 gnd.n4648 gnd.n4646 0.152939
R15466 gnd.n4648 gnd.n4647 0.152939
R15467 gnd.n4647 gnd.n554 0.152939
R15468 gnd.n555 gnd.n554 0.152939
R15469 gnd.n556 gnd.n555 0.152939
R15470 gnd.n559 gnd.n556 0.152939
R15471 gnd.n560 gnd.n559 0.152939
R15472 gnd.n2957 gnd.n2898 0.152939
R15473 gnd.n2963 gnd.n2898 0.152939
R15474 gnd.n2964 gnd.n2963 0.152939
R15475 gnd.n2965 gnd.n2964 0.152939
R15476 gnd.n2965 gnd.n2896 0.152939
R15477 gnd.n2971 gnd.n2896 0.152939
R15478 gnd.n2972 gnd.n2971 0.152939
R15479 gnd.n2973 gnd.n2972 0.152939
R15480 gnd.n2973 gnd.n2894 0.152939
R15481 gnd.n2979 gnd.n2894 0.152939
R15482 gnd.n2980 gnd.n2979 0.152939
R15483 gnd.n2981 gnd.n2980 0.152939
R15484 gnd.n2981 gnd.n2892 0.152939
R15485 gnd.n2987 gnd.n2892 0.152939
R15486 gnd.n2988 gnd.n2987 0.152939
R15487 gnd.n2989 gnd.n2988 0.152939
R15488 gnd.n2989 gnd.n2890 0.152939
R15489 gnd.n2995 gnd.n2890 0.152939
R15490 gnd.n2996 gnd.n2995 0.152939
R15491 gnd.n2997 gnd.n2996 0.152939
R15492 gnd.n2997 gnd.n2888 0.152939
R15493 gnd.n3003 gnd.n2888 0.152939
R15494 gnd.n3004 gnd.n3003 0.152939
R15495 gnd.n3005 gnd.n3004 0.152939
R15496 gnd.n3005 gnd.n2886 0.152939
R15497 gnd.n3011 gnd.n2886 0.152939
R15498 gnd.n3012 gnd.n3011 0.152939
R15499 gnd.n3013 gnd.n3012 0.152939
R15500 gnd.n3013 gnd.n2884 0.152939
R15501 gnd.n3019 gnd.n2884 0.152939
R15502 gnd.n3020 gnd.n3019 0.152939
R15503 gnd.n2912 gnd.n1254 0.152939
R15504 gnd.n2920 gnd.n2912 0.152939
R15505 gnd.n2921 gnd.n2920 0.152939
R15506 gnd.n2922 gnd.n2921 0.152939
R15507 gnd.n2922 gnd.n2910 0.152939
R15508 gnd.n2930 gnd.n2910 0.152939
R15509 gnd.n2931 gnd.n2930 0.152939
R15510 gnd.n2932 gnd.n2931 0.152939
R15511 gnd.n2932 gnd.n2908 0.152939
R15512 gnd.n2940 gnd.n2908 0.152939
R15513 gnd.n2941 gnd.n2940 0.152939
R15514 gnd.n2942 gnd.n2941 0.152939
R15515 gnd.n2942 gnd.n2906 0.152939
R15516 gnd.n2950 gnd.n2906 0.152939
R15517 gnd.n2951 gnd.n2950 0.152939
R15518 gnd.n2952 gnd.n2951 0.152939
R15519 gnd.n2952 gnd.n2899 0.152939
R15520 gnd.n2956 gnd.n2899 0.152939
R15521 gnd.n5188 gnd.n1403 0.152939
R15522 gnd.n1428 gnd.n1403 0.152939
R15523 gnd.n1429 gnd.n1428 0.152939
R15524 gnd.n1430 gnd.n1429 0.152939
R15525 gnd.n1448 gnd.n1430 0.152939
R15526 gnd.n1449 gnd.n1448 0.152939
R15527 gnd.n1450 gnd.n1449 0.152939
R15528 gnd.n1451 gnd.n1450 0.152939
R15529 gnd.n1468 gnd.n1451 0.152939
R15530 gnd.n1469 gnd.n1468 0.152939
R15531 gnd.n1470 gnd.n1469 0.152939
R15532 gnd.n1471 gnd.n1470 0.152939
R15533 gnd.n1489 gnd.n1471 0.152939
R15534 gnd.n1490 gnd.n1489 0.152939
R15535 gnd.n1491 gnd.n1490 0.152939
R15536 gnd.n1492 gnd.n1491 0.152939
R15537 gnd.n1509 gnd.n1492 0.152939
R15538 gnd.n1510 gnd.n1509 0.152939
R15539 gnd.n1511 gnd.n1510 0.152939
R15540 gnd.n1512 gnd.n1511 0.152939
R15541 gnd.n1530 gnd.n1512 0.152939
R15542 gnd.n1531 gnd.n1530 0.152939
R15543 gnd.n1532 gnd.n1531 0.152939
R15544 gnd.n1533 gnd.n1532 0.152939
R15545 gnd.n1551 gnd.n1533 0.152939
R15546 gnd.n1552 gnd.n1551 0.152939
R15547 gnd.n5103 gnd.n1552 0.152939
R15548 gnd.n5102 gnd.n1553 0.152939
R15549 gnd.n1597 gnd.n1553 0.152939
R15550 gnd.n1598 gnd.n1597 0.152939
R15551 gnd.n1599 gnd.n1598 0.152939
R15552 gnd.n1600 gnd.n1599 0.152939
R15553 gnd.n1601 gnd.n1600 0.152939
R15554 gnd.n1602 gnd.n1601 0.152939
R15555 gnd.n1603 gnd.n1602 0.152939
R15556 gnd.n1604 gnd.n1603 0.152939
R15557 gnd.n1605 gnd.n1604 0.152939
R15558 gnd.n1606 gnd.n1605 0.152939
R15559 gnd.n1607 gnd.n1606 0.152939
R15560 gnd.n1608 gnd.n1607 0.152939
R15561 gnd.n1609 gnd.n1608 0.152939
R15562 gnd.n1610 gnd.n1609 0.152939
R15563 gnd.n1611 gnd.n1610 0.152939
R15564 gnd.n1612 gnd.n1611 0.152939
R15565 gnd.n1615 gnd.n1612 0.152939
R15566 gnd.n1616 gnd.n1615 0.152939
R15567 gnd.n1617 gnd.n1616 0.152939
R15568 gnd.n1618 gnd.n1617 0.152939
R15569 gnd.n1619 gnd.n1618 0.152939
R15570 gnd.n1620 gnd.n1619 0.152939
R15571 gnd.n1621 gnd.n1620 0.152939
R15572 gnd.n1622 gnd.n1621 0.152939
R15573 gnd.n2661 gnd.n2660 0.152939
R15574 gnd.n2668 gnd.n2661 0.152939
R15575 gnd.n2669 gnd.n2668 0.152939
R15576 gnd.n2670 gnd.n2669 0.152939
R15577 gnd.n2670 gnd.n2658 0.152939
R15578 gnd.n2678 gnd.n2658 0.152939
R15579 gnd.n2679 gnd.n2678 0.152939
R15580 gnd.n2680 gnd.n2679 0.152939
R15581 gnd.n2680 gnd.n2653 0.152939
R15582 gnd.n2687 gnd.n2653 0.152939
R15583 gnd.n2688 gnd.n2687 0.152939
R15584 gnd.n2689 gnd.n2688 0.152939
R15585 gnd.n2689 gnd.n2651 0.152939
R15586 gnd.n2697 gnd.n2651 0.152939
R15587 gnd.n2698 gnd.n2697 0.152939
R15588 gnd.n2699 gnd.n2698 0.152939
R15589 gnd.n2699 gnd.n2649 0.152939
R15590 gnd.n2707 gnd.n2649 0.152939
R15591 gnd.n2708 gnd.n2707 0.152939
R15592 gnd.n2709 gnd.n2708 0.152939
R15593 gnd.n2709 gnd.n2647 0.152939
R15594 gnd.n2717 gnd.n2647 0.152939
R15595 gnd.n2718 gnd.n2717 0.152939
R15596 gnd.n2719 gnd.n2718 0.152939
R15597 gnd.n2719 gnd.n2645 0.152939
R15598 gnd.n2727 gnd.n2645 0.152939
R15599 gnd.n2728 gnd.n2727 0.152939
R15600 gnd.n2729 gnd.n2728 0.152939
R15601 gnd.n2729 gnd.n2640 0.152939
R15602 gnd.n2735 gnd.n2640 0.152939
R15603 gnd.n1191 gnd.n1190 0.152939
R15604 gnd.n1192 gnd.n1191 0.152939
R15605 gnd.n1193 gnd.n1192 0.152939
R15606 gnd.n1194 gnd.n1193 0.152939
R15607 gnd.n1195 gnd.n1194 0.152939
R15608 gnd.n1196 gnd.n1195 0.152939
R15609 gnd.n1197 gnd.n1196 0.152939
R15610 gnd.n1198 gnd.n1197 0.152939
R15611 gnd.n1199 gnd.n1198 0.152939
R15612 gnd.n1200 gnd.n1199 0.152939
R15613 gnd.n1201 gnd.n1200 0.152939
R15614 gnd.n1202 gnd.n1201 0.152939
R15615 gnd.n1203 gnd.n1202 0.152939
R15616 gnd.n1204 gnd.n1203 0.152939
R15617 gnd.n1205 gnd.n1204 0.152939
R15618 gnd.n1206 gnd.n1205 0.152939
R15619 gnd.n1207 gnd.n1206 0.152939
R15620 gnd.n1210 gnd.n1207 0.152939
R15621 gnd.n1211 gnd.n1210 0.152939
R15622 gnd.n1212 gnd.n1211 0.152939
R15623 gnd.n1213 gnd.n1212 0.152939
R15624 gnd.n1214 gnd.n1213 0.152939
R15625 gnd.n1215 gnd.n1214 0.152939
R15626 gnd.n1216 gnd.n1215 0.152939
R15627 gnd.n1217 gnd.n1216 0.152939
R15628 gnd.n1218 gnd.n1217 0.152939
R15629 gnd.n1219 gnd.n1218 0.152939
R15630 gnd.n1220 gnd.n1219 0.152939
R15631 gnd.n1221 gnd.n1220 0.152939
R15632 gnd.n1222 gnd.n1221 0.152939
R15633 gnd.n1223 gnd.n1222 0.152939
R15634 gnd.n1224 gnd.n1223 0.152939
R15635 gnd.n1225 gnd.n1224 0.152939
R15636 gnd.n1226 gnd.n1225 0.152939
R15637 gnd.n1227 gnd.n1226 0.152939
R15638 gnd.n1228 gnd.n1227 0.152939
R15639 gnd.n1229 gnd.n1228 0.152939
R15640 gnd.n1232 gnd.n1229 0.152939
R15641 gnd.n1233 gnd.n1232 0.152939
R15642 gnd.n1234 gnd.n1233 0.152939
R15643 gnd.n1235 gnd.n1234 0.152939
R15644 gnd.n1236 gnd.n1235 0.152939
R15645 gnd.n1237 gnd.n1236 0.152939
R15646 gnd.n1238 gnd.n1237 0.152939
R15647 gnd.n1239 gnd.n1238 0.152939
R15648 gnd.n1240 gnd.n1239 0.152939
R15649 gnd.n1241 gnd.n1240 0.152939
R15650 gnd.n1242 gnd.n1241 0.152939
R15651 gnd.n1243 gnd.n1242 0.152939
R15652 gnd.n1244 gnd.n1243 0.152939
R15653 gnd.n1245 gnd.n1244 0.152939
R15654 gnd.n1246 gnd.n1245 0.152939
R15655 gnd.n1247 gnd.n1246 0.152939
R15656 gnd.n1248 gnd.n1247 0.152939
R15657 gnd.n1249 gnd.n1248 0.152939
R15658 gnd.n1250 gnd.n1249 0.152939
R15659 gnd.n5283 gnd.n1250 0.152939
R15660 gnd.n5283 gnd.n5282 0.152939
R15661 gnd.n1265 gnd.n1264 0.152939
R15662 gnd.n1266 gnd.n1265 0.152939
R15663 gnd.n1267 gnd.n1266 0.152939
R15664 gnd.n1287 gnd.n1267 0.152939
R15665 gnd.n1288 gnd.n1287 0.152939
R15666 gnd.n1289 gnd.n1288 0.152939
R15667 gnd.n1290 gnd.n1289 0.152939
R15668 gnd.n1305 gnd.n1290 0.152939
R15669 gnd.n1306 gnd.n1305 0.152939
R15670 gnd.n1307 gnd.n1306 0.152939
R15671 gnd.n1308 gnd.n1307 0.152939
R15672 gnd.n1325 gnd.n1308 0.152939
R15673 gnd.n1326 gnd.n1325 0.152939
R15674 gnd.n1327 gnd.n1326 0.152939
R15675 gnd.n1328 gnd.n1327 0.152939
R15676 gnd.n1343 gnd.n1328 0.152939
R15677 gnd.n1344 gnd.n1343 0.152939
R15678 gnd.n1345 gnd.n1344 0.152939
R15679 gnd.n1346 gnd.n1345 0.152939
R15680 gnd.n1363 gnd.n1346 0.152939
R15681 gnd.n1364 gnd.n1363 0.152939
R15682 gnd.n1365 gnd.n1364 0.152939
R15683 gnd.n1366 gnd.n1365 0.152939
R15684 gnd.n1381 gnd.n1366 0.152939
R15685 gnd.n1382 gnd.n1381 0.152939
R15686 gnd.n1383 gnd.n1382 0.152939
R15687 gnd.n5188 gnd.n1383 0.152939
R15688 gnd.n2812 gnd.n2811 0.152939
R15689 gnd.n2813 gnd.n2812 0.152939
R15690 gnd.n2815 gnd.n2814 0.152939
R15691 gnd.n2815 gnd.n2781 0.152939
R15692 gnd.n3059 gnd.n2781 0.152939
R15693 gnd.n971 gnd.n966 0.152939
R15694 gnd.n972 gnd.n971 0.152939
R15695 gnd.n973 gnd.n972 0.152939
R15696 gnd.n978 gnd.n973 0.152939
R15697 gnd.n979 gnd.n978 0.152939
R15698 gnd.n980 gnd.n979 0.152939
R15699 gnd.n981 gnd.n980 0.152939
R15700 gnd.n986 gnd.n981 0.152939
R15701 gnd.n987 gnd.n986 0.152939
R15702 gnd.n988 gnd.n987 0.152939
R15703 gnd.n989 gnd.n988 0.152939
R15704 gnd.n994 gnd.n989 0.152939
R15705 gnd.n995 gnd.n994 0.152939
R15706 gnd.n996 gnd.n995 0.152939
R15707 gnd.n997 gnd.n996 0.152939
R15708 gnd.n1002 gnd.n997 0.152939
R15709 gnd.n1003 gnd.n1002 0.152939
R15710 gnd.n1004 gnd.n1003 0.152939
R15711 gnd.n1005 gnd.n1004 0.152939
R15712 gnd.n1010 gnd.n1005 0.152939
R15713 gnd.n1011 gnd.n1010 0.152939
R15714 gnd.n1012 gnd.n1011 0.152939
R15715 gnd.n1013 gnd.n1012 0.152939
R15716 gnd.n1018 gnd.n1013 0.152939
R15717 gnd.n1019 gnd.n1018 0.152939
R15718 gnd.n1020 gnd.n1019 0.152939
R15719 gnd.n1021 gnd.n1020 0.152939
R15720 gnd.n1026 gnd.n1021 0.152939
R15721 gnd.n1027 gnd.n1026 0.152939
R15722 gnd.n1028 gnd.n1027 0.152939
R15723 gnd.n1029 gnd.n1028 0.152939
R15724 gnd.n1034 gnd.n1029 0.152939
R15725 gnd.n1035 gnd.n1034 0.152939
R15726 gnd.n1036 gnd.n1035 0.152939
R15727 gnd.n1037 gnd.n1036 0.152939
R15728 gnd.n1042 gnd.n1037 0.152939
R15729 gnd.n1043 gnd.n1042 0.152939
R15730 gnd.n1044 gnd.n1043 0.152939
R15731 gnd.n1045 gnd.n1044 0.152939
R15732 gnd.n1050 gnd.n1045 0.152939
R15733 gnd.n1051 gnd.n1050 0.152939
R15734 gnd.n1052 gnd.n1051 0.152939
R15735 gnd.n1053 gnd.n1052 0.152939
R15736 gnd.n1058 gnd.n1053 0.152939
R15737 gnd.n1059 gnd.n1058 0.152939
R15738 gnd.n1060 gnd.n1059 0.152939
R15739 gnd.n1061 gnd.n1060 0.152939
R15740 gnd.n1066 gnd.n1061 0.152939
R15741 gnd.n1067 gnd.n1066 0.152939
R15742 gnd.n1068 gnd.n1067 0.152939
R15743 gnd.n1069 gnd.n1068 0.152939
R15744 gnd.n1074 gnd.n1069 0.152939
R15745 gnd.n1075 gnd.n1074 0.152939
R15746 gnd.n1076 gnd.n1075 0.152939
R15747 gnd.n1077 gnd.n1076 0.152939
R15748 gnd.n1082 gnd.n1077 0.152939
R15749 gnd.n1083 gnd.n1082 0.152939
R15750 gnd.n1084 gnd.n1083 0.152939
R15751 gnd.n1085 gnd.n1084 0.152939
R15752 gnd.n1090 gnd.n1085 0.152939
R15753 gnd.n1091 gnd.n1090 0.152939
R15754 gnd.n1092 gnd.n1091 0.152939
R15755 gnd.n1093 gnd.n1092 0.152939
R15756 gnd.n1098 gnd.n1093 0.152939
R15757 gnd.n1099 gnd.n1098 0.152939
R15758 gnd.n1100 gnd.n1099 0.152939
R15759 gnd.n1101 gnd.n1100 0.152939
R15760 gnd.n1106 gnd.n1101 0.152939
R15761 gnd.n1107 gnd.n1106 0.152939
R15762 gnd.n1108 gnd.n1107 0.152939
R15763 gnd.n1109 gnd.n1108 0.152939
R15764 gnd.n1114 gnd.n1109 0.152939
R15765 gnd.n1115 gnd.n1114 0.152939
R15766 gnd.n1116 gnd.n1115 0.152939
R15767 gnd.n1117 gnd.n1116 0.152939
R15768 gnd.n1122 gnd.n1117 0.152939
R15769 gnd.n1123 gnd.n1122 0.152939
R15770 gnd.n1124 gnd.n1123 0.152939
R15771 gnd.n1125 gnd.n1124 0.152939
R15772 gnd.n1130 gnd.n1125 0.152939
R15773 gnd.n1131 gnd.n1130 0.152939
R15774 gnd.n1132 gnd.n1131 0.152939
R15775 gnd.n1133 gnd.n1132 0.152939
R15776 gnd.n2810 gnd.n1133 0.152939
R15777 gnd.n3370 gnd.n2533 0.152939
R15778 gnd.n3384 gnd.n2533 0.152939
R15779 gnd.n3385 gnd.n3384 0.152939
R15780 gnd.n3386 gnd.n3385 0.152939
R15781 gnd.n3386 gnd.n2519 0.152939
R15782 gnd.n3400 gnd.n2519 0.152939
R15783 gnd.n3401 gnd.n3400 0.152939
R15784 gnd.n3402 gnd.n3401 0.152939
R15785 gnd.n3402 gnd.n2504 0.152939
R15786 gnd.n3416 gnd.n2504 0.152939
R15787 gnd.n3417 gnd.n3416 0.152939
R15788 gnd.n3418 gnd.n3417 0.152939
R15789 gnd.n3418 gnd.n2489 0.152939
R15790 gnd.n3441 gnd.n2489 0.152939
R15791 gnd.n3442 gnd.n3441 0.152939
R15792 gnd.n3443 gnd.n3442 0.152939
R15793 gnd.n3443 gnd.n2485 0.152939
R15794 gnd.n3449 gnd.n2485 0.152939
R15795 gnd.n3450 gnd.n3449 0.152939
R15796 gnd.n3452 gnd.n3450 0.152939
R15797 gnd.n3452 gnd.n3451 0.152939
R15798 gnd.n3451 gnd.n2388 0.152939
R15799 gnd.n4094 gnd.n2388 0.152939
R15800 gnd.n4095 gnd.n4094 0.152939
R15801 gnd.n4096 gnd.n4095 0.152939
R15802 gnd.n4096 gnd.n2375 0.152939
R15803 gnd.n4110 gnd.n2375 0.152939
R15804 gnd.n4111 gnd.n4110 0.152939
R15805 gnd.n4112 gnd.n4111 0.152939
R15806 gnd.n4112 gnd.n2362 0.152939
R15807 gnd.n4126 gnd.n2362 0.152939
R15808 gnd.n4127 gnd.n4126 0.152939
R15809 gnd.n4128 gnd.n4127 0.152939
R15810 gnd.n4128 gnd.n2349 0.152939
R15811 gnd.n4142 gnd.n2349 0.152939
R15812 gnd.n4143 gnd.n4142 0.152939
R15813 gnd.n4144 gnd.n4143 0.152939
R15814 gnd.n4144 gnd.n2336 0.152939
R15815 gnd.n4158 gnd.n2336 0.152939
R15816 gnd.n4159 gnd.n4158 0.152939
R15817 gnd.n4160 gnd.n4159 0.152939
R15818 gnd.n4160 gnd.n2320 0.152939
R15819 gnd.n4174 gnd.n2320 0.152939
R15820 gnd.n4175 gnd.n4174 0.152939
R15821 gnd.n4176 gnd.n4175 0.152939
R15822 gnd.n4176 gnd.n2306 0.152939
R15823 gnd.n4190 gnd.n2306 0.152939
R15824 gnd.n4191 gnd.n4190 0.152939
R15825 gnd.n4192 gnd.n4191 0.152939
R15826 gnd.n4192 gnd.n2292 0.152939
R15827 gnd.n4206 gnd.n2292 0.152939
R15828 gnd.n4207 gnd.n4206 0.152939
R15829 gnd.n4208 gnd.n4207 0.152939
R15830 gnd.n4208 gnd.n2279 0.152939
R15831 gnd.n4222 gnd.n2279 0.152939
R15832 gnd.n4223 gnd.n4222 0.152939
R15833 gnd.n4224 gnd.n4223 0.152939
R15834 gnd.n4224 gnd.n2265 0.152939
R15835 gnd.n4238 gnd.n2265 0.152939
R15836 gnd.n4239 gnd.n4238 0.152939
R15837 gnd.n4240 gnd.n4239 0.152939
R15838 gnd.n4240 gnd.n2251 0.152939
R15839 gnd.n4254 gnd.n2251 0.152939
R15840 gnd.n4255 gnd.n4254 0.152939
R15841 gnd.n4256 gnd.n4255 0.152939
R15842 gnd.n4256 gnd.n2238 0.152939
R15843 gnd.n4270 gnd.n2238 0.152939
R15844 gnd.n4271 gnd.n4270 0.152939
R15845 gnd.n4272 gnd.n4271 0.152939
R15846 gnd.n4272 gnd.n2225 0.152939
R15847 gnd.n4286 gnd.n2225 0.152939
R15848 gnd.n4287 gnd.n4286 0.152939
R15849 gnd.n4288 gnd.n4287 0.152939
R15850 gnd.n4288 gnd.n2210 0.152939
R15851 gnd.n4302 gnd.n2210 0.152939
R15852 gnd.n4303 gnd.n4302 0.152939
R15853 gnd.n4304 gnd.n4303 0.152939
R15854 gnd.n4304 gnd.n2196 0.152939
R15855 gnd.n4318 gnd.n2196 0.152939
R15856 gnd.n4319 gnd.n4318 0.152939
R15857 gnd.n4320 gnd.n4319 0.152939
R15858 gnd.n4320 gnd.n2184 0.152939
R15859 gnd.n4334 gnd.n2184 0.152939
R15860 gnd.n4335 gnd.n4334 0.152939
R15861 gnd.n4336 gnd.n4335 0.152939
R15862 gnd.n4336 gnd.n2172 0.152939
R15863 gnd.n4350 gnd.n2172 0.152939
R15864 gnd.n4351 gnd.n4350 0.152939
R15865 gnd.n4352 gnd.n4351 0.152939
R15866 gnd.n4352 gnd.n2159 0.152939
R15867 gnd.n4366 gnd.n2159 0.152939
R15868 gnd.n4367 gnd.n4366 0.152939
R15869 gnd.n4368 gnd.n4367 0.152939
R15870 gnd.n4368 gnd.n2146 0.152939
R15871 gnd.n4382 gnd.n2146 0.152939
R15872 gnd.n4383 gnd.n4382 0.152939
R15873 gnd.n4386 gnd.n4383 0.152939
R15874 gnd.n4386 gnd.n4385 0.152939
R15875 gnd.n4385 gnd.n4384 0.152939
R15876 gnd.n4384 gnd.n2131 0.152939
R15877 gnd.n4405 gnd.n2131 0.152939
R15878 gnd.n3049 gnd.n2788 0.152939
R15879 gnd.n3050 gnd.n3049 0.152939
R15880 gnd.n3051 gnd.n3050 0.152939
R15881 gnd.n3051 gnd.n2775 0.152939
R15882 gnd.n3088 gnd.n2775 0.152939
R15883 gnd.n3089 gnd.n3088 0.152939
R15884 gnd.n3090 gnd.n3089 0.152939
R15885 gnd.n3090 gnd.n2770 0.152939
R15886 gnd.n3102 gnd.n2770 0.152939
R15887 gnd.n3103 gnd.n3102 0.152939
R15888 gnd.n3104 gnd.n3103 0.152939
R15889 gnd.n3104 gnd.n2761 0.152939
R15890 gnd.n3139 gnd.n2761 0.152939
R15891 gnd.n3139 gnd.n3138 0.152939
R15892 gnd.n3138 gnd.n3137 0.152939
R15893 gnd.n3137 gnd.n2762 0.152939
R15894 gnd.n3133 gnd.n2762 0.152939
R15895 gnd.n3133 gnd.n3132 0.152939
R15896 gnd.n3132 gnd.n3131 0.152939
R15897 gnd.n3131 gnd.n2766 0.152939
R15898 gnd.n3127 gnd.n2766 0.152939
R15899 gnd.n3127 gnd.n2743 0.152939
R15900 gnd.n3196 gnd.n2743 0.152939
R15901 gnd.n3197 gnd.n3196 0.152939
R15902 gnd.n3198 gnd.n3197 0.152939
R15903 gnd.n3198 gnd.n2739 0.152939
R15904 gnd.n3211 gnd.n2739 0.152939
R15905 gnd.n3212 gnd.n3211 0.152939
R15906 gnd.n3215 gnd.n3212 0.152939
R15907 gnd.n3215 gnd.n3214 0.152939
R15908 gnd.n3214 gnd.n3213 0.152939
R15909 gnd.n3346 gnd.n2633 0.152939
R15910 gnd.n3346 gnd.n3345 0.152939
R15911 gnd.n3345 gnd.n3344 0.152939
R15912 gnd.n3344 gnd.n2635 0.152939
R15913 gnd.n3340 gnd.n2635 0.152939
R15914 gnd.n3340 gnd.n3339 0.152939
R15915 gnd.n2632 gnd.n2582 0.152939
R15916 gnd.n2628 gnd.n2582 0.152939
R15917 gnd.n2628 gnd.n2627 0.152939
R15918 gnd.n2627 gnd.n2626 0.152939
R15919 gnd.n2626 gnd.n2586 0.152939
R15920 gnd.n2622 gnd.n2586 0.152939
R15921 gnd.n2622 gnd.n2621 0.152939
R15922 gnd.n2621 gnd.n2620 0.152939
R15923 gnd.n2620 gnd.n2590 0.152939
R15924 gnd.n2616 gnd.n2590 0.152939
R15925 gnd.n2616 gnd.n2615 0.152939
R15926 gnd.n2615 gnd.n2614 0.152939
R15927 gnd.n2614 gnd.n2594 0.152939
R15928 gnd.n2610 gnd.n2594 0.152939
R15929 gnd.n2610 gnd.n2609 0.152939
R15930 gnd.n2609 gnd.n2608 0.152939
R15931 gnd.n2608 gnd.n2597 0.152939
R15932 gnd.n2604 gnd.n2597 0.152939
R15933 gnd.n2604 gnd.n2603 0.152939
R15934 gnd.n2603 gnd.n1708 0.152939
R15935 gnd.n4966 gnd.n1708 0.152939
R15936 gnd.n4966 gnd.n4965 0.152939
R15937 gnd.n4965 gnd.n4964 0.152939
R15938 gnd.n4964 gnd.n1709 0.152939
R15939 gnd.n4960 gnd.n1709 0.152939
R15940 gnd.n4960 gnd.n4959 0.152939
R15941 gnd.n4959 gnd.n4958 0.152939
R15942 gnd.n4958 gnd.n1714 0.152939
R15943 gnd.n4954 gnd.n1714 0.152939
R15944 gnd.n4954 gnd.n4953 0.152939
R15945 gnd.n4953 gnd.n4952 0.152939
R15946 gnd.n4952 gnd.n1719 0.152939
R15947 gnd.n4948 gnd.n1719 0.152939
R15948 gnd.n4948 gnd.n4947 0.152939
R15949 gnd.n4947 gnd.n4946 0.152939
R15950 gnd.n4946 gnd.n1724 0.152939
R15951 gnd.n4942 gnd.n1724 0.152939
R15952 gnd.n4942 gnd.n4941 0.152939
R15953 gnd.n4941 gnd.n4940 0.152939
R15954 gnd.n4940 gnd.n1729 0.152939
R15955 gnd.n4936 gnd.n1729 0.152939
R15956 gnd.n4936 gnd.n4935 0.152939
R15957 gnd.n4935 gnd.n4934 0.152939
R15958 gnd.n4934 gnd.n1734 0.152939
R15959 gnd.n4930 gnd.n1734 0.152939
R15960 gnd.n4930 gnd.n4929 0.152939
R15961 gnd.n4929 gnd.n4928 0.152939
R15962 gnd.n4928 gnd.n1739 0.152939
R15963 gnd.n4924 gnd.n1739 0.152939
R15964 gnd.n4924 gnd.n4923 0.152939
R15965 gnd.n4923 gnd.n4922 0.152939
R15966 gnd.n4922 gnd.n1744 0.152939
R15967 gnd.n4918 gnd.n1744 0.152939
R15968 gnd.n4918 gnd.n4917 0.152939
R15969 gnd.n4917 gnd.n4916 0.152939
R15970 gnd.n4916 gnd.n1749 0.152939
R15971 gnd.n4912 gnd.n1749 0.152939
R15972 gnd.n4912 gnd.n4911 0.152939
R15973 gnd.n4911 gnd.n4910 0.152939
R15974 gnd.n4910 gnd.n1754 0.152939
R15975 gnd.n4906 gnd.n1754 0.152939
R15976 gnd.n4906 gnd.n4905 0.152939
R15977 gnd.n4905 gnd.n4904 0.152939
R15978 gnd.n4904 gnd.n1759 0.152939
R15979 gnd.n4900 gnd.n1759 0.152939
R15980 gnd.n4900 gnd.n4899 0.152939
R15981 gnd.n4899 gnd.n4898 0.152939
R15982 gnd.n4898 gnd.n1764 0.152939
R15983 gnd.n4894 gnd.n1764 0.152939
R15984 gnd.n4894 gnd.n4893 0.152939
R15985 gnd.n4893 gnd.n4892 0.152939
R15986 gnd.n4892 gnd.n1769 0.152939
R15987 gnd.n4888 gnd.n1769 0.152939
R15988 gnd.n4888 gnd.n4887 0.152939
R15989 gnd.n4887 gnd.n4886 0.152939
R15990 gnd.n4886 gnd.n1774 0.152939
R15991 gnd.n4882 gnd.n1774 0.152939
R15992 gnd.n4882 gnd.n4881 0.152939
R15993 gnd.n4881 gnd.n4880 0.152939
R15994 gnd.n4880 gnd.n1779 0.152939
R15995 gnd.n4876 gnd.n1779 0.152939
R15996 gnd.n4876 gnd.n4875 0.152939
R15997 gnd.n4875 gnd.n4874 0.152939
R15998 gnd.n4874 gnd.n1784 0.152939
R15999 gnd.n4870 gnd.n1784 0.152939
R16000 gnd.n4870 gnd.n4869 0.152939
R16001 gnd.n4869 gnd.n4868 0.152939
R16002 gnd.n4868 gnd.n1789 0.152939
R16003 gnd.n4864 gnd.n1789 0.152939
R16004 gnd.n4864 gnd.n4863 0.152939
R16005 gnd.n4863 gnd.n4862 0.152939
R16006 gnd.n4862 gnd.n1794 0.152939
R16007 gnd.n4858 gnd.n1794 0.152939
R16008 gnd.n4858 gnd.n4857 0.152939
R16009 gnd.n4857 gnd.n4856 0.152939
R16010 gnd.n4856 gnd.n1799 0.152939
R16011 gnd.n4852 gnd.n1799 0.152939
R16012 gnd.n4852 gnd.n4851 0.152939
R16013 gnd.n4851 gnd.n4850 0.152939
R16014 gnd.n4850 gnd.n1804 0.152939
R16015 gnd.n1807 gnd.n1804 0.152939
R16016 gnd.n4454 gnd.n4453 0.152939
R16017 gnd.n4454 gnd.n4449 0.152939
R16018 gnd.n4462 gnd.n4449 0.152939
R16019 gnd.n4463 gnd.n4462 0.152939
R16020 gnd.n4465 gnd.n4463 0.152939
R16021 gnd.n4465 gnd.n4464 0.152939
R16022 gnd.n4569 gnd.n4568 0.152939
R16023 gnd.n4570 gnd.n4569 0.152939
R16024 gnd.n4570 gnd.n2127 0.152939
R16025 gnd.n4582 gnd.n2127 0.152939
R16026 gnd.n4583 gnd.n4582 0.152939
R16027 gnd.n4584 gnd.n4583 0.152939
R16028 gnd.n4584 gnd.n2122 0.152939
R16029 gnd.n4596 gnd.n2122 0.152939
R16030 gnd.n4597 gnd.n4596 0.152939
R16031 gnd.n4598 gnd.n4597 0.152939
R16032 gnd.n4598 gnd.n2059 0.152939
R16033 gnd.n4610 gnd.n2059 0.152939
R16034 gnd.n4611 gnd.n4610 0.152939
R16035 gnd.n4612 gnd.n4611 0.152939
R16036 gnd.n4612 gnd.n2054 0.152939
R16037 gnd.n4627 gnd.n2054 0.152939
R16038 gnd.n4628 gnd.n4627 0.152939
R16039 gnd.n4637 gnd.n4628 0.152939
R16040 gnd.n4637 gnd.n4636 0.152939
R16041 gnd.n4636 gnd.n4635 0.152939
R16042 gnd.n4635 gnd.n4629 0.152939
R16043 gnd.n4631 gnd.n4629 0.152939
R16044 gnd.n4631 gnd.n529 0.152939
R16045 gnd.n7771 gnd.n529 0.152939
R16046 gnd.n7772 gnd.n7771 0.152939
R16047 gnd.n7773 gnd.n7772 0.152939
R16048 gnd.n7773 gnd.n507 0.152939
R16049 gnd.n7798 gnd.n507 0.152939
R16050 gnd.n7799 gnd.n7798 0.152939
R16051 gnd.n7800 gnd.n7799 0.152939
R16052 gnd.n7800 gnd.n99 0.152939
R16053 gnd.n8102 gnd.n8101 0.145814
R16054 gnd.n3021 gnd.n3020 0.145814
R16055 gnd.n3021 gnd.n2788 0.145814
R16056 gnd.n8102 gnd.n99 0.145814
R16057 gnd.n3339 gnd.n3338 0.128549
R16058 gnd.n4464 gnd.n1928 0.128549
R16059 gnd.n562 gnd.n115 0.0950122
R16060 gnd.n2814 gnd.n1404 0.0950122
R16061 gnd.n6329 gnd.n6213 0.0767195
R16062 gnd.n6329 gnd.n6211 0.0767195
R16063 gnd.n3338 gnd.n3224 0.063
R16064 gnd.n4720 gnd.n1928 0.063
R16065 gnd.n566 gnd.n115 0.0584268
R16066 gnd.n2813 gnd.n1404 0.0584268
R16067 gnd.n6840 gnd.n5435 0.0477147
R16068 gnd.n6153 gnd.n6049 0.0442063
R16069 gnd.n6167 gnd.n6049 0.0442063
R16070 gnd.n6168 gnd.n6167 0.0442063
R16071 gnd.n6169 gnd.n6168 0.0442063
R16072 gnd.n6169 gnd.n6037 0.0442063
R16073 gnd.n6183 gnd.n6037 0.0442063
R16074 gnd.n6184 gnd.n6183 0.0442063
R16075 gnd.n6185 gnd.n6184 0.0442063
R16076 gnd.n6185 gnd.n6024 0.0442063
R16077 gnd.n6426 gnd.n6024 0.0442063
R16078 gnd.n4720 gnd.n4719 0.0416005
R16079 gnd.n7883 gnd.n7882 0.0416005
R16080 gnd.n5281 gnd.n5280 0.0416005
R16081 gnd.n3224 gnd.n3223 0.0416005
R16082 gnd.n6429 gnd.n6428 0.0344674
R16083 gnd.n4719 gnd.n1930 0.0344674
R16084 gnd.n2129 gnd.n1930 0.0344674
R16085 gnd.n2129 gnd.n1956 0.0344674
R16086 gnd.n1957 gnd.n1956 0.0344674
R16087 gnd.n1958 gnd.n1957 0.0344674
R16088 gnd.n2125 gnd.n1958 0.0344674
R16089 gnd.n2125 gnd.n1977 0.0344674
R16090 gnd.n1978 gnd.n1977 0.0344674
R16091 gnd.n1979 gnd.n1978 0.0344674
R16092 gnd.n2062 gnd.n1979 0.0344674
R16093 gnd.n2062 gnd.n1997 0.0344674
R16094 gnd.n1998 gnd.n1997 0.0344674
R16095 gnd.n1999 gnd.n1998 0.0344674
R16096 gnd.n2057 gnd.n1999 0.0344674
R16097 gnd.n2057 gnd.n2018 0.0344674
R16098 gnd.n2019 gnd.n2018 0.0344674
R16099 gnd.n2020 gnd.n2019 0.0344674
R16100 gnd.n4619 gnd.n2020 0.0344674
R16101 gnd.n4619 gnd.n2039 0.0344674
R16102 gnd.n4655 gnd.n2039 0.0344674
R16103 gnd.n4655 gnd.n2040 0.0344674
R16104 gnd.n2040 gnd.n548 0.0344674
R16105 gnd.n549 gnd.n548 0.0344674
R16106 gnd.n7748 gnd.n549 0.0344674
R16107 gnd.n7749 gnd.n7748 0.0344674
R16108 gnd.n7749 gnd.n524 0.0344674
R16109 gnd.n524 gnd.n519 0.0344674
R16110 gnd.n520 gnd.n519 0.0344674
R16111 gnd.n521 gnd.n520 0.0344674
R16112 gnd.n521 gnd.n494 0.0344674
R16113 gnd.n7816 gnd.n494 0.0344674
R16114 gnd.n7817 gnd.n7816 0.0344674
R16115 gnd.n7817 gnd.n489 0.0344674
R16116 gnd.n489 gnd.n487 0.0344674
R16117 gnd.n7828 gnd.n487 0.0344674
R16118 gnd.n7829 gnd.n7828 0.0344674
R16119 gnd.n7829 gnd.n129 0.0344674
R16120 gnd.n130 gnd.n129 0.0344674
R16121 gnd.n131 gnd.n130 0.0344674
R16122 gnd.n7837 gnd.n131 0.0344674
R16123 gnd.n7837 gnd.n146 0.0344674
R16124 gnd.n147 gnd.n146 0.0344674
R16125 gnd.n148 gnd.n147 0.0344674
R16126 gnd.n7844 gnd.n148 0.0344674
R16127 gnd.n7844 gnd.n166 0.0344674
R16128 gnd.n167 gnd.n166 0.0344674
R16129 gnd.n168 gnd.n167 0.0344674
R16130 gnd.n7851 gnd.n168 0.0344674
R16131 gnd.n7851 gnd.n184 0.0344674
R16132 gnd.n185 gnd.n184 0.0344674
R16133 gnd.n186 gnd.n185 0.0344674
R16134 gnd.n7858 gnd.n186 0.0344674
R16135 gnd.n7858 gnd.n204 0.0344674
R16136 gnd.n205 gnd.n204 0.0344674
R16137 gnd.n206 gnd.n205 0.0344674
R16138 gnd.n7865 gnd.n206 0.0344674
R16139 gnd.n7865 gnd.n223 0.0344674
R16140 gnd.n224 gnd.n223 0.0344674
R16141 gnd.n225 gnd.n224 0.0344674
R16142 gnd.n7872 gnd.n225 0.0344674
R16143 gnd.n7872 gnd.n243 0.0344674
R16144 gnd.n244 gnd.n243 0.0344674
R16145 gnd.n245 gnd.n244 0.0344674
R16146 gnd.n7882 gnd.n245 0.0344674
R16147 gnd.n5280 gnd.n1256 0.0344674
R16148 gnd.n2825 gnd.n1256 0.0344674
R16149 gnd.n2825 gnd.n1278 0.0344674
R16150 gnd.n1279 gnd.n1278 0.0344674
R16151 gnd.n1280 gnd.n1279 0.0344674
R16152 gnd.n2831 gnd.n1280 0.0344674
R16153 gnd.n2831 gnd.n1297 0.0344674
R16154 gnd.n1298 gnd.n1297 0.0344674
R16155 gnd.n1299 gnd.n1298 0.0344674
R16156 gnd.n2838 gnd.n1299 0.0344674
R16157 gnd.n2838 gnd.n1316 0.0344674
R16158 gnd.n1317 gnd.n1316 0.0344674
R16159 gnd.n1318 gnd.n1317 0.0344674
R16160 gnd.n2845 gnd.n1318 0.0344674
R16161 gnd.n2845 gnd.n1335 0.0344674
R16162 gnd.n1336 gnd.n1335 0.0344674
R16163 gnd.n1337 gnd.n1336 0.0344674
R16164 gnd.n2852 gnd.n1337 0.0344674
R16165 gnd.n2852 gnd.n1354 0.0344674
R16166 gnd.n1355 gnd.n1354 0.0344674
R16167 gnd.n1356 gnd.n1355 0.0344674
R16168 gnd.n2859 gnd.n1356 0.0344674
R16169 gnd.n2859 gnd.n1373 0.0344674
R16170 gnd.n1374 gnd.n1373 0.0344674
R16171 gnd.n1375 gnd.n1374 0.0344674
R16172 gnd.n2866 gnd.n1375 0.0344674
R16173 gnd.n2866 gnd.n1391 0.0344674
R16174 gnd.n1392 gnd.n1391 0.0344674
R16175 gnd.n1393 gnd.n1392 0.0344674
R16176 gnd.n2875 gnd.n1393 0.0344674
R16177 gnd.n2876 gnd.n2875 0.0344674
R16178 gnd.n2876 gnd.n2806 0.0344674
R16179 gnd.n2806 gnd.n2802 0.0344674
R16180 gnd.n2803 gnd.n2802 0.0344674
R16181 gnd.n3034 gnd.n2803 0.0344674
R16182 gnd.n3034 gnd.n2804 0.0344674
R16183 gnd.n2804 gnd.n1419 0.0344674
R16184 gnd.n1420 gnd.n1419 0.0344674
R16185 gnd.n1421 gnd.n1420 0.0344674
R16186 gnd.n2773 gnd.n1421 0.0344674
R16187 gnd.n2773 gnd.n1438 0.0344674
R16188 gnd.n1439 gnd.n1438 0.0344674
R16189 gnd.n1440 gnd.n1439 0.0344674
R16190 gnd.n2768 gnd.n1440 0.0344674
R16191 gnd.n2768 gnd.n1459 0.0344674
R16192 gnd.n1460 gnd.n1459 0.0344674
R16193 gnd.n1461 gnd.n1460 0.0344674
R16194 gnd.n3113 gnd.n1461 0.0344674
R16195 gnd.n3113 gnd.n1479 0.0344674
R16196 gnd.n1480 gnd.n1479 0.0344674
R16197 gnd.n1481 gnd.n1480 0.0344674
R16198 gnd.n3122 gnd.n1481 0.0344674
R16199 gnd.n3122 gnd.n1500 0.0344674
R16200 gnd.n1501 gnd.n1500 0.0344674
R16201 gnd.n1502 gnd.n1501 0.0344674
R16202 gnd.n3190 gnd.n1502 0.0344674
R16203 gnd.n3190 gnd.n1520 0.0344674
R16204 gnd.n1521 gnd.n1520 0.0344674
R16205 gnd.n1522 gnd.n1521 0.0344674
R16206 gnd.n3205 gnd.n1522 0.0344674
R16207 gnd.n3205 gnd.n1541 0.0344674
R16208 gnd.n1542 gnd.n1541 0.0344674
R16209 gnd.n1543 gnd.n1542 0.0344674
R16210 gnd.n3223 gnd.n1543 0.0344674
R16211 gnd.n3337 gnd.n3225 0.0343753
R16212 gnd.n4474 gnd.n4473 0.0343753
R16213 gnd.n3366 gnd.n2546 0.0296328
R16214 gnd.n4566 gnd.n4565 0.0296328
R16215 gnd.n6017 gnd.n6016 0.0269946
R16216 gnd.n6439 gnd.n6437 0.0269946
R16217 gnd.n6438 gnd.n5999 0.0269946
R16218 gnd.n6458 gnd.n6457 0.0269946
R16219 gnd.n6460 gnd.n6459 0.0269946
R16220 gnd.n5993 gnd.n5991 0.0269946
R16221 gnd.n6470 gnd.n6468 0.0269946
R16222 gnd.n6469 gnd.n5972 0.0269946
R16223 gnd.n6489 gnd.n6488 0.0269946
R16224 gnd.n6491 gnd.n6490 0.0269946
R16225 gnd.n5967 gnd.n5965 0.0269946
R16226 gnd.n6501 gnd.n6499 0.0269946
R16227 gnd.n6500 gnd.n5946 0.0269946
R16228 gnd.n6520 gnd.n6519 0.0269946
R16229 gnd.n6522 gnd.n6521 0.0269946
R16230 gnd.n5941 gnd.n5939 0.0269946
R16231 gnd.n6532 gnd.n6530 0.0269946
R16232 gnd.n6531 gnd.n5921 0.0269946
R16233 gnd.n6551 gnd.n6550 0.0269946
R16234 gnd.n6553 gnd.n6552 0.0269946
R16235 gnd.n5915 gnd.n5913 0.0269946
R16236 gnd.n6563 gnd.n6561 0.0269946
R16237 gnd.n6562 gnd.n5896 0.0269946
R16238 gnd.n6582 gnd.n6581 0.0269946
R16239 gnd.n6584 gnd.n6583 0.0269946
R16240 gnd.n5890 gnd.n5888 0.0269946
R16241 gnd.n6594 gnd.n6592 0.0269946
R16242 gnd.n6593 gnd.n5871 0.0269946
R16243 gnd.n6613 gnd.n6612 0.0269946
R16244 gnd.n6615 gnd.n6614 0.0269946
R16245 gnd.n5865 gnd.n5863 0.0269946
R16246 gnd.n6625 gnd.n6623 0.0269946
R16247 gnd.n6624 gnd.n5847 0.0269946
R16248 gnd.n6643 gnd.n6642 0.0269946
R16249 gnd.n6645 gnd.n6644 0.0269946
R16250 gnd.n5835 gnd.n5834 0.0269946
R16251 gnd.n6666 gnd.n5830 0.0269946
R16252 gnd.n6665 gnd.n5832 0.0269946
R16253 gnd.n5831 gnd.n5812 0.0269946
R16254 gnd.n6689 gnd.n5813 0.0269946
R16255 gnd.n6688 gnd.n5814 0.0269946
R16256 gnd.n6708 gnd.n5798 0.0269946
R16257 gnd.n6710 gnd.n6709 0.0269946
R16258 gnd.n6711 gnd.n5783 0.0269946
R16259 gnd.n6734 gnd.n5784 0.0269946
R16260 gnd.n6733 gnd.n5785 0.0269946
R16261 gnd.n6753 gnd.n5771 0.0269946
R16262 gnd.n6756 gnd.n6755 0.0269946
R16263 gnd.n6775 gnd.n5749 0.0269946
R16264 gnd.n5751 gnd.n1141 0.0269946
R16265 gnd.n5755 gnd.n1142 0.0269946
R16266 gnd.n5756 gnd.n1143 0.0269946
R16267 gnd.n3333 gnd.n3231 0.022519
R16268 gnd.n3332 gnd.n3232 0.022519
R16269 gnd.n3329 gnd.n3328 0.022519
R16270 gnd.n3325 gnd.n3238 0.022519
R16271 gnd.n3324 gnd.n3244 0.022519
R16272 gnd.n3321 gnd.n3320 0.022519
R16273 gnd.n3317 gnd.n3248 0.022519
R16274 gnd.n3316 gnd.n3252 0.022519
R16275 gnd.n3313 gnd.n3312 0.022519
R16276 gnd.n3309 gnd.n3258 0.022519
R16277 gnd.n3308 gnd.n3264 0.022519
R16278 gnd.n3305 gnd.n3304 0.022519
R16279 gnd.n3301 gnd.n3268 0.022519
R16280 gnd.n3300 gnd.n3272 0.022519
R16281 gnd.n3297 gnd.n3296 0.022519
R16282 gnd.n3293 gnd.n3278 0.022519
R16283 gnd.n3292 gnd.n3288 0.022519
R16284 gnd.n3285 gnd.n2549 0.022519
R16285 gnd.n3366 gnd.n3365 0.022519
R16286 gnd.n4482 gnd.n4475 0.022519
R16287 gnd.n4481 gnd.n4476 0.022519
R16288 gnd.n4490 gnd.n4442 0.022519
R16289 gnd.n4492 gnd.n4491 0.022519
R16290 gnd.n4501 gnd.n4439 0.022519
R16291 gnd.n4500 gnd.n4440 0.022519
R16292 gnd.n4509 gnd.n4435 0.022519
R16293 gnd.n4511 gnd.n4510 0.022519
R16294 gnd.n4520 gnd.n4432 0.022519
R16295 gnd.n4519 gnd.n4433 0.022519
R16296 gnd.n4528 gnd.n4428 0.022519
R16297 gnd.n4530 gnd.n4529 0.022519
R16298 gnd.n4539 gnd.n4424 0.022519
R16299 gnd.n4538 gnd.n4426 0.022519
R16300 gnd.n4425 gnd.n4420 0.022519
R16301 gnd.n4548 gnd.n4547 0.022519
R16302 gnd.n4555 gnd.n4413 0.022519
R16303 gnd.n4554 gnd.n4414 0.022519
R16304 gnd.n4565 gnd.n4407 0.022519
R16305 gnd.n4566 gnd.n4406 0.0218415
R16306 gnd.n3369 gnd.n2546 0.0218415
R16307 gnd.n6428 gnd.n6427 0.0202011
R16308 gnd.n6427 gnd.n6426 0.0148637
R16309 gnd.n6754 gnd.n5748 0.0144266
R16310 gnd.n6776 gnd.n5748 0.0130679
R16311 gnd.n3231 gnd.n3225 0.0123564
R16312 gnd.n3333 gnd.n3332 0.0123564
R16313 gnd.n3329 gnd.n3232 0.0123564
R16314 gnd.n3328 gnd.n3238 0.0123564
R16315 gnd.n3325 gnd.n3324 0.0123564
R16316 gnd.n3321 gnd.n3244 0.0123564
R16317 gnd.n3320 gnd.n3248 0.0123564
R16318 gnd.n3317 gnd.n3316 0.0123564
R16319 gnd.n3313 gnd.n3252 0.0123564
R16320 gnd.n3312 gnd.n3258 0.0123564
R16321 gnd.n3309 gnd.n3308 0.0123564
R16322 gnd.n3305 gnd.n3264 0.0123564
R16323 gnd.n3304 gnd.n3268 0.0123564
R16324 gnd.n3301 gnd.n3300 0.0123564
R16325 gnd.n3297 gnd.n3272 0.0123564
R16326 gnd.n3296 gnd.n3278 0.0123564
R16327 gnd.n3293 gnd.n3292 0.0123564
R16328 gnd.n3288 gnd.n3285 0.0123564
R16329 gnd.n3365 gnd.n2549 0.0123564
R16330 gnd.n4475 gnd.n4474 0.0123564
R16331 gnd.n4482 gnd.n4481 0.0123564
R16332 gnd.n4476 gnd.n4442 0.0123564
R16333 gnd.n4492 gnd.n4490 0.0123564
R16334 gnd.n4491 gnd.n4439 0.0123564
R16335 gnd.n4501 gnd.n4500 0.0123564
R16336 gnd.n4440 gnd.n4435 0.0123564
R16337 gnd.n4511 gnd.n4509 0.0123564
R16338 gnd.n4510 gnd.n4432 0.0123564
R16339 gnd.n4520 gnd.n4519 0.0123564
R16340 gnd.n4433 gnd.n4428 0.0123564
R16341 gnd.n4530 gnd.n4528 0.0123564
R16342 gnd.n4529 gnd.n4424 0.0123564
R16343 gnd.n4539 gnd.n4538 0.0123564
R16344 gnd.n4426 gnd.n4425 0.0123564
R16345 gnd.n4548 gnd.n4420 0.0123564
R16346 gnd.n4547 gnd.n4413 0.0123564
R16347 gnd.n4555 gnd.n4554 0.0123564
R16348 gnd.n4414 gnd.n4407 0.0123564
R16349 gnd.n6429 gnd.n6017 0.00797283
R16350 gnd.n6437 gnd.n6016 0.00797283
R16351 gnd.n6439 gnd.n6438 0.00797283
R16352 gnd.n6457 gnd.n5999 0.00797283
R16353 gnd.n6459 gnd.n6458 0.00797283
R16354 gnd.n6460 gnd.n5993 0.00797283
R16355 gnd.n6468 gnd.n5991 0.00797283
R16356 gnd.n6470 gnd.n6469 0.00797283
R16357 gnd.n6488 gnd.n5972 0.00797283
R16358 gnd.n6490 gnd.n6489 0.00797283
R16359 gnd.n6491 gnd.n5967 0.00797283
R16360 gnd.n6499 gnd.n5965 0.00797283
R16361 gnd.n6501 gnd.n6500 0.00797283
R16362 gnd.n6519 gnd.n5946 0.00797283
R16363 gnd.n6521 gnd.n6520 0.00797283
R16364 gnd.n6522 gnd.n5941 0.00797283
R16365 gnd.n6530 gnd.n5939 0.00797283
R16366 gnd.n6532 gnd.n6531 0.00797283
R16367 gnd.n6550 gnd.n5921 0.00797283
R16368 gnd.n6552 gnd.n6551 0.00797283
R16369 gnd.n6553 gnd.n5915 0.00797283
R16370 gnd.n6561 gnd.n5913 0.00797283
R16371 gnd.n6563 gnd.n6562 0.00797283
R16372 gnd.n6581 gnd.n5896 0.00797283
R16373 gnd.n6583 gnd.n6582 0.00797283
R16374 gnd.n6584 gnd.n5890 0.00797283
R16375 gnd.n6592 gnd.n5888 0.00797283
R16376 gnd.n6594 gnd.n6593 0.00797283
R16377 gnd.n6612 gnd.n5871 0.00797283
R16378 gnd.n6614 gnd.n6613 0.00797283
R16379 gnd.n6615 gnd.n5865 0.00797283
R16380 gnd.n6623 gnd.n5863 0.00797283
R16381 gnd.n6625 gnd.n6624 0.00797283
R16382 gnd.n6642 gnd.n5847 0.00797283
R16383 gnd.n6644 gnd.n6643 0.00797283
R16384 gnd.n6645 gnd.n5835 0.00797283
R16385 gnd.n5834 gnd.n5830 0.00797283
R16386 gnd.n6666 gnd.n6665 0.00797283
R16387 gnd.n5832 gnd.n5831 0.00797283
R16388 gnd.n5813 gnd.n5812 0.00797283
R16389 gnd.n6689 gnd.n6688 0.00797283
R16390 gnd.n5814 gnd.n5798 0.00797283
R16391 gnd.n6709 gnd.n6708 0.00797283
R16392 gnd.n6711 gnd.n6710 0.00797283
R16393 gnd.n5784 gnd.n5783 0.00797283
R16394 gnd.n6734 gnd.n6733 0.00797283
R16395 gnd.n5785 gnd.n5771 0.00797283
R16396 gnd.n6756 gnd.n6753 0.00797283
R16397 gnd.n6755 gnd.n6754 0.00797283
R16398 gnd.n6776 gnd.n6775 0.00797283
R16399 gnd.n5751 gnd.n5749 0.00797283
R16400 gnd.n5755 gnd.n1141 0.00797283
R16401 gnd.n5756 gnd.n1142 0.00797283
R16402 gnd.n5435 gnd.n1143 0.00797283
R16403 gnd.n3338 gnd.n3337 0.00592005
R16404 gnd.n4473 gnd.n1928 0.00592005
R16405 a_n2982_13878.n133 a_n2982_13878.t90 512.366
R16406 a_n2982_13878.n132 a_n2982_13878.t79 512.366
R16407 a_n2982_13878.n131 a_n2982_13878.t68 512.366
R16408 a_n2982_13878.n135 a_n2982_13878.t98 512.366
R16409 a_n2982_13878.n134 a_n2982_13878.t87 512.366
R16410 a_n2982_13878.n130 a_n2982_13878.t86 512.366
R16411 a_n2982_13878.n137 a_n2982_13878.t94 512.366
R16412 a_n2982_13878.n136 a_n2982_13878.t77 512.366
R16413 a_n2982_13878.n129 a_n2982_13878.t78 512.366
R16414 a_n2982_13878.n139 a_n2982_13878.t81 512.366
R16415 a_n2982_13878.n138 a_n2982_13878.t92 512.366
R16416 a_n2982_13878.n128 a_n2982_13878.t107 512.366
R16417 a_n2982_13878.n34 a_n2982_13878.t106 538.698
R16418 a_n2982_13878.n104 a_n2982_13878.t83 512.366
R16419 a_n2982_13878.n103 a_n2982_13878.t88 512.366
R16420 a_n2982_13878.n95 a_n2982_13878.t76 512.366
R16421 a_n2982_13878.n102 a_n2982_13878.t93 512.366
R16422 a_n2982_13878.n101 a_n2982_13878.t102 512.366
R16423 a_n2982_13878.n96 a_n2982_13878.t103 512.366
R16424 a_n2982_13878.n100 a_n2982_13878.t70 512.366
R16425 a_n2982_13878.n99 a_n2982_13878.t85 512.366
R16426 a_n2982_13878.n97 a_n2982_13878.t73 512.366
R16427 a_n2982_13878.n98 a_n2982_13878.t80 512.366
R16428 a_n2982_13878.n28 a_n2982_13878.t49 538.698
R16429 a_n2982_13878.n121 a_n2982_13878.t19 512.366
R16430 a_n2982_13878.n120 a_n2982_13878.t15 512.366
R16431 a_n2982_13878.n93 a_n2982_13878.t55 512.366
R16432 a_n2982_13878.n119 a_n2982_13878.t51 512.366
R16433 a_n2982_13878.n118 a_n2982_13878.t37 512.366
R16434 a_n2982_13878.n94 a_n2982_13878.t45 512.366
R16435 a_n2982_13878.n117 a_n2982_13878.t35 512.366
R16436 a_n2982_13878.n116 a_n2982_13878.t23 512.366
R16437 a_n2982_13878.n83 a_n2982_13878.t47 512.366
R16438 a_n2982_13878.n105 a_n2982_13878.t25 512.366
R16439 a_n2982_13878.n17 a_n2982_13878.t27 538.698
R16440 a_n2982_13878.n147 a_n2982_13878.t53 512.366
R16441 a_n2982_13878.n88 a_n2982_13878.t33 512.366
R16442 a_n2982_13878.n148 a_n2982_13878.t57 512.366
R16443 a_n2982_13878.n87 a_n2982_13878.t11 512.366
R16444 a_n2982_13878.n149 a_n2982_13878.t39 512.366
R16445 a_n2982_13878.n150 a_n2982_13878.t41 512.366
R16446 a_n2982_13878.n86 a_n2982_13878.t29 512.366
R16447 a_n2982_13878.n151 a_n2982_13878.t31 512.366
R16448 a_n2982_13878.n85 a_n2982_13878.t13 512.366
R16449 a_n2982_13878.n152 a_n2982_13878.t17 512.366
R16450 a_n2982_13878.n23 a_n2982_13878.t105 538.698
R16451 a_n2982_13878.n141 a_n2982_13878.t74 512.366
R16452 a_n2982_13878.n92 a_n2982_13878.t75 512.366
R16453 a_n2982_13878.n142 a_n2982_13878.t100 512.366
R16454 a_n2982_13878.n91 a_n2982_13878.t101 512.366
R16455 a_n2982_13878.n143 a_n2982_13878.t72 512.366
R16456 a_n2982_13878.n144 a_n2982_13878.t96 512.366
R16457 a_n2982_13878.n90 a_n2982_13878.t97 512.366
R16458 a_n2982_13878.n145 a_n2982_13878.t69 512.366
R16459 a_n2982_13878.n89 a_n2982_13878.t82 512.366
R16460 a_n2982_13878.n146 a_n2982_13878.t91 512.366
R16461 a_n2982_13878.n4 a_n2982_13878.n81 70.1674
R16462 a_n2982_13878.n6 a_n2982_13878.n79 70.1674
R16463 a_n2982_13878.n8 a_n2982_13878.n77 70.1674
R16464 a_n2982_13878.n10 a_n2982_13878.n75 70.1674
R16465 a_n2982_13878.n51 a_n2982_13878.n29 70.5844
R16466 a_n2982_13878.n42 a_n2982_13878.n35 70.5844
R16467 a_n2982_13878.n35 a_n2982_13878.n82 70.1674
R16468 a_n2982_13878.n29 a_n2982_13878.n49 70.1674
R16469 a_n2982_13878.n49 a_n2982_13878.n97 20.9683
R16470 a_n2982_13878.n48 a_n2982_13878.n30 74.73
R16471 a_n2982_13878.n99 a_n2982_13878.n48 11.843
R16472 a_n2982_13878.n47 a_n2982_13878.n30 80.4688
R16473 a_n2982_13878.n47 a_n2982_13878.n100 0.365327
R16474 a_n2982_13878.n31 a_n2982_13878.n46 75.0448
R16475 a_n2982_13878.n45 a_n2982_13878.n31 70.1674
R16476 a_n2982_13878.n102 a_n2982_13878.n45 20.9683
R16477 a_n2982_13878.n33 a_n2982_13878.n44 70.3058
R16478 a_n2982_13878.n44 a_n2982_13878.n95 20.6913
R16479 a_n2982_13878.n43 a_n2982_13878.n33 75.3623
R16480 a_n2982_13878.n103 a_n2982_13878.n43 10.5784
R16481 a_n2982_13878.n32 a_n2982_13878.n34 44.7878
R16482 a_n2982_13878.n82 a_n2982_13878.n83 20.9683
R16483 a_n2982_13878.n57 a_n2982_13878.n35 74.73
R16484 a_n2982_13878.n116 a_n2982_13878.n57 11.843
R16485 a_n2982_13878.n56 a_n2982_13878.n24 80.4688
R16486 a_n2982_13878.n56 a_n2982_13878.n117 0.365327
R16487 a_n2982_13878.n25 a_n2982_13878.n55 75.0448
R16488 a_n2982_13878.n54 a_n2982_13878.n25 70.1674
R16489 a_n2982_13878.n119 a_n2982_13878.n54 20.9683
R16490 a_n2982_13878.n27 a_n2982_13878.n53 70.3058
R16491 a_n2982_13878.n53 a_n2982_13878.n93 20.6913
R16492 a_n2982_13878.n52 a_n2982_13878.n27 75.3623
R16493 a_n2982_13878.n120 a_n2982_13878.n52 10.5784
R16494 a_n2982_13878.n26 a_n2982_13878.n28 44.7878
R16495 a_n2982_13878.n13 a_n2982_13878.n73 70.5844
R16496 a_n2982_13878.n19 a_n2982_13878.n65 70.5844
R16497 a_n2982_13878.n64 a_n2982_13878.n19 70.1674
R16498 a_n2982_13878.n64 a_n2982_13878.n89 20.9683
R16499 a_n2982_13878.n18 a_n2982_13878.n63 74.73
R16500 a_n2982_13878.n145 a_n2982_13878.n63 11.843
R16501 a_n2982_13878.n62 a_n2982_13878.n18 80.4688
R16502 a_n2982_13878.n62 a_n2982_13878.n90 0.365327
R16503 a_n2982_13878.n20 a_n2982_13878.n61 75.0448
R16504 a_n2982_13878.n60 a_n2982_13878.n20 70.1674
R16505 a_n2982_13878.n60 a_n2982_13878.n91 20.9683
R16506 a_n2982_13878.n21 a_n2982_13878.n59 70.3058
R16507 a_n2982_13878.n142 a_n2982_13878.n59 20.6913
R16508 a_n2982_13878.n58 a_n2982_13878.n21 75.3623
R16509 a_n2982_13878.n58 a_n2982_13878.n92 10.5784
R16510 a_n2982_13878.n23 a_n2982_13878.n22 44.7878
R16511 a_n2982_13878.n72 a_n2982_13878.n13 70.1674
R16512 a_n2982_13878.n72 a_n2982_13878.n85 20.9683
R16513 a_n2982_13878.n12 a_n2982_13878.n71 74.73
R16514 a_n2982_13878.n151 a_n2982_13878.n71 11.843
R16515 a_n2982_13878.n70 a_n2982_13878.n12 80.4688
R16516 a_n2982_13878.n70 a_n2982_13878.n86 0.365327
R16517 a_n2982_13878.n14 a_n2982_13878.n69 75.0448
R16518 a_n2982_13878.n68 a_n2982_13878.n14 70.1674
R16519 a_n2982_13878.n68 a_n2982_13878.n87 20.9683
R16520 a_n2982_13878.n15 a_n2982_13878.n67 70.3058
R16521 a_n2982_13878.n148 a_n2982_13878.n67 20.6913
R16522 a_n2982_13878.n66 a_n2982_13878.n15 75.3623
R16523 a_n2982_13878.n66 a_n2982_13878.n88 10.5784
R16524 a_n2982_13878.n17 a_n2982_13878.n16 44.7878
R16525 a_n2982_13878.n75 a_n2982_13878.n128 20.9683
R16526 a_n2982_13878.n74 a_n2982_13878.n11 75.0448
R16527 a_n2982_13878.n138 a_n2982_13878.n74 11.2134
R16528 a_n2982_13878.n11 a_n2982_13878.n139 161.3
R16529 a_n2982_13878.n77 a_n2982_13878.n129 20.9683
R16530 a_n2982_13878.n76 a_n2982_13878.n9 75.0448
R16531 a_n2982_13878.n136 a_n2982_13878.n76 11.2134
R16532 a_n2982_13878.n9 a_n2982_13878.n137 161.3
R16533 a_n2982_13878.n79 a_n2982_13878.n130 20.9683
R16534 a_n2982_13878.n78 a_n2982_13878.n7 75.0448
R16535 a_n2982_13878.n134 a_n2982_13878.n78 11.2134
R16536 a_n2982_13878.n7 a_n2982_13878.n135 161.3
R16537 a_n2982_13878.n81 a_n2982_13878.n131 20.9683
R16538 a_n2982_13878.n80 a_n2982_13878.n5 75.0448
R16539 a_n2982_13878.n132 a_n2982_13878.n80 11.2134
R16540 a_n2982_13878.n5 a_n2982_13878.n133 161.3
R16541 a_n2982_13878.n3 a_n2982_13878.n114 81.4626
R16542 a_n2982_13878.n1 a_n2982_13878.n109 81.4626
R16543 a_n2982_13878.n0 a_n2982_13878.n106 81.4626
R16544 a_n2982_13878.n3 a_n2982_13878.n115 80.9324
R16545 a_n2982_13878.n3 a_n2982_13878.n113 80.9324
R16546 a_n2982_13878.n2 a_n2982_13878.n112 80.9324
R16547 a_n2982_13878.n2 a_n2982_13878.n111 80.9324
R16548 a_n2982_13878.n1 a_n2982_13878.n110 80.9324
R16549 a_n2982_13878.n1 a_n2982_13878.n108 80.9324
R16550 a_n2982_13878.n0 a_n2982_13878.n107 80.9324
R16551 a_n2982_13878.n40 a_n2982_13878.t28 74.6477
R16552 a_n2982_13878.n38 a_n2982_13878.t44 74.6477
R16553 a_n2982_13878.n37 a_n2982_13878.t50 74.2899
R16554 a_n2982_13878.n41 a_n2982_13878.t22 74.2897
R16555 a_n2982_13878.n41 a_n2982_13878.n154 70.6783
R16556 a_n2982_13878.n39 a_n2982_13878.n155 70.6783
R16557 a_n2982_13878.n39 a_n2982_13878.n156 70.6783
R16558 a_n2982_13878.n40 a_n2982_13878.n84 70.6783
R16559 a_n2982_13878.n38 a_n2982_13878.n122 70.6783
R16560 a_n2982_13878.n38 a_n2982_13878.n123 70.6783
R16561 a_n2982_13878.n36 a_n2982_13878.n124 70.6783
R16562 a_n2982_13878.n36 a_n2982_13878.n125 70.6783
R16563 a_n2982_13878.n37 a_n2982_13878.n126 70.6783
R16564 a_n2982_13878.n157 a_n2982_13878.n40 70.6782
R16565 a_n2982_13878.n133 a_n2982_13878.n132 48.2005
R16566 a_n2982_13878.t95 a_n2982_13878.n81 533.335
R16567 a_n2982_13878.n135 a_n2982_13878.n134 48.2005
R16568 a_n2982_13878.t104 a_n2982_13878.n79 533.335
R16569 a_n2982_13878.n137 a_n2982_13878.n136 48.2005
R16570 a_n2982_13878.t89 a_n2982_13878.n77 533.335
R16571 a_n2982_13878.n139 a_n2982_13878.n138 48.2005
R16572 a_n2982_13878.t84 a_n2982_13878.n75 533.335
R16573 a_n2982_13878.n104 a_n2982_13878.n103 48.2005
R16574 a_n2982_13878.n45 a_n2982_13878.n101 20.9683
R16575 a_n2982_13878.n100 a_n2982_13878.n96 48.2005
R16576 a_n2982_13878.n98 a_n2982_13878.n49 20.9683
R16577 a_n2982_13878.n121 a_n2982_13878.n120 48.2005
R16578 a_n2982_13878.n54 a_n2982_13878.n118 20.9683
R16579 a_n2982_13878.n117 a_n2982_13878.n94 48.2005
R16580 a_n2982_13878.n105 a_n2982_13878.n82 20.9683
R16581 a_n2982_13878.n147 a_n2982_13878.n88 48.2005
R16582 a_n2982_13878.n149 a_n2982_13878.n68 20.9683
R16583 a_n2982_13878.n150 a_n2982_13878.n86 48.2005
R16584 a_n2982_13878.n152 a_n2982_13878.n72 20.9683
R16585 a_n2982_13878.n141 a_n2982_13878.n92 48.2005
R16586 a_n2982_13878.n143 a_n2982_13878.n60 20.9683
R16587 a_n2982_13878.n144 a_n2982_13878.n90 48.2005
R16588 a_n2982_13878.n146 a_n2982_13878.n64 20.9683
R16589 a_n2982_13878.n102 a_n2982_13878.n44 21.4216
R16590 a_n2982_13878.n119 a_n2982_13878.n53 21.4216
R16591 a_n2982_13878.n87 a_n2982_13878.n67 21.4216
R16592 a_n2982_13878.n91 a_n2982_13878.n59 21.4216
R16593 a_n2982_13878.n51 a_n2982_13878.t99 532.5
R16594 a_n2982_13878.n42 a_n2982_13878.t43 532.5
R16595 a_n2982_13878.t21 a_n2982_13878.n73 532.5
R16596 a_n2982_13878.t71 a_n2982_13878.n65 532.5
R16597 a_n2982_13878.n2 a_n2982_13878.n1 32.7898
R16598 a_n2982_13878.n48 a_n2982_13878.n97 34.4824
R16599 a_n2982_13878.n57 a_n2982_13878.n83 34.4824
R16600 a_n2982_13878.n85 a_n2982_13878.n71 34.4824
R16601 a_n2982_13878.n89 a_n2982_13878.n63 34.4824
R16602 a_n2982_13878.n80 a_n2982_13878.n131 35.3134
R16603 a_n2982_13878.n78 a_n2982_13878.n130 35.3134
R16604 a_n2982_13878.n76 a_n2982_13878.n129 35.3134
R16605 a_n2982_13878.n74 a_n2982_13878.n128 35.3134
R16606 a_n2982_13878.n101 a_n2982_13878.n46 35.3134
R16607 a_n2982_13878.n46 a_n2982_13878.n96 11.2134
R16608 a_n2982_13878.n118 a_n2982_13878.n55 35.3134
R16609 a_n2982_13878.n55 a_n2982_13878.n94 11.2134
R16610 a_n2982_13878.n69 a_n2982_13878.n149 35.3134
R16611 a_n2982_13878.n150 a_n2982_13878.n69 11.2134
R16612 a_n2982_13878.n61 a_n2982_13878.n143 35.3134
R16613 a_n2982_13878.n144 a_n2982_13878.n61 11.2134
R16614 a_n2982_13878.n35 a_n2982_13878.n3 23.891
R16615 a_n2982_13878.n43 a_n2982_13878.n95 36.139
R16616 a_n2982_13878.n52 a_n2982_13878.n93 36.139
R16617 a_n2982_13878.n148 a_n2982_13878.n66 36.139
R16618 a_n2982_13878.n142 a_n2982_13878.n58 36.139
R16619 a_n2982_13878.n22 a_n2982_13878.n140 13.9285
R16620 a_n2982_13878.n29 a_n2982_13878.n50 13.724
R16621 a_n2982_13878.n127 a_n2982_13878.n26 12.4191
R16622 a_n2982_13878.n140 a_n2982_13878.n11 11.2486
R16623 a_n2982_13878.n4 a_n2982_13878.n50 11.2486
R16624 a_n2982_13878.n41 a_n2982_13878.n153 10.5745
R16625 a_n2982_13878.n153 a_n2982_13878.n13 8.58383
R16626 a_n2982_13878.n127 a_n2982_13878.n37 6.7311
R16627 a_n2982_13878.n153 a_n2982_13878.n50 5.3452
R16628 a_n2982_13878.n35 a_n2982_13878.n32 3.94368
R16629 a_n2982_13878.n16 a_n2982_13878.n19 3.94368
R16630 a_n2982_13878.n154 a_n2982_13878.t14 3.61217
R16631 a_n2982_13878.n154 a_n2982_13878.t18 3.61217
R16632 a_n2982_13878.n155 a_n2982_13878.t30 3.61217
R16633 a_n2982_13878.n155 a_n2982_13878.t32 3.61217
R16634 a_n2982_13878.n156 a_n2982_13878.t40 3.61217
R16635 a_n2982_13878.n156 a_n2982_13878.t42 3.61217
R16636 a_n2982_13878.n84 a_n2982_13878.t54 3.61217
R16637 a_n2982_13878.n84 a_n2982_13878.t34 3.61217
R16638 a_n2982_13878.n122 a_n2982_13878.t48 3.61217
R16639 a_n2982_13878.n122 a_n2982_13878.t26 3.61217
R16640 a_n2982_13878.n123 a_n2982_13878.t36 3.61217
R16641 a_n2982_13878.n123 a_n2982_13878.t24 3.61217
R16642 a_n2982_13878.n124 a_n2982_13878.t38 3.61217
R16643 a_n2982_13878.n124 a_n2982_13878.t46 3.61217
R16644 a_n2982_13878.n125 a_n2982_13878.t56 3.61217
R16645 a_n2982_13878.n125 a_n2982_13878.t52 3.61217
R16646 a_n2982_13878.n126 a_n2982_13878.t20 3.61217
R16647 a_n2982_13878.n126 a_n2982_13878.t16 3.61217
R16648 a_n2982_13878.n157 a_n2982_13878.t58 3.61217
R16649 a_n2982_13878.t12 a_n2982_13878.n157 3.61217
R16650 a_n2982_13878.n114 a_n2982_13878.t60 2.82907
R16651 a_n2982_13878.n114 a_n2982_13878.t4 2.82907
R16652 a_n2982_13878.n115 a_n2982_13878.t7 2.82907
R16653 a_n2982_13878.n115 a_n2982_13878.t5 2.82907
R16654 a_n2982_13878.n113 a_n2982_13878.t8 2.82907
R16655 a_n2982_13878.n113 a_n2982_13878.t10 2.82907
R16656 a_n2982_13878.n112 a_n2982_13878.t66 2.82907
R16657 a_n2982_13878.n112 a_n2982_13878.t9 2.82907
R16658 a_n2982_13878.n111 a_n2982_13878.t6 2.82907
R16659 a_n2982_13878.n111 a_n2982_13878.t0 2.82907
R16660 a_n2982_13878.n109 a_n2982_13878.t62 2.82907
R16661 a_n2982_13878.n109 a_n2982_13878.t65 2.82907
R16662 a_n2982_13878.n110 a_n2982_13878.t64 2.82907
R16663 a_n2982_13878.n110 a_n2982_13878.t59 2.82907
R16664 a_n2982_13878.n108 a_n2982_13878.t1 2.82907
R16665 a_n2982_13878.n108 a_n2982_13878.t3 2.82907
R16666 a_n2982_13878.n107 a_n2982_13878.t63 2.82907
R16667 a_n2982_13878.n107 a_n2982_13878.t2 2.82907
R16668 a_n2982_13878.n106 a_n2982_13878.t61 2.82907
R16669 a_n2982_13878.n106 a_n2982_13878.t67 2.82907
R16670 a_n2982_13878.n34 a_n2982_13878.n104 14.1668
R16671 a_n2982_13878.n98 a_n2982_13878.n51 22.3251
R16672 a_n2982_13878.n28 a_n2982_13878.n121 14.1668
R16673 a_n2982_13878.n105 a_n2982_13878.n42 22.3251
R16674 a_n2982_13878.n147 a_n2982_13878.n17 14.1668
R16675 a_n2982_13878.n73 a_n2982_13878.n152 22.3251
R16676 a_n2982_13878.n141 a_n2982_13878.n23 14.1668
R16677 a_n2982_13878.n65 a_n2982_13878.n146 22.3251
R16678 a_n2982_13878.n140 a_n2982_13878.n127 1.30542
R16679 a_n2982_13878.n8 a_n2982_13878.n7 1.04595
R16680 a_n2982_13878.n47 a_n2982_13878.n99 47.835
R16681 a_n2982_13878.n56 a_n2982_13878.n116 47.835
R16682 a_n2982_13878.n151 a_n2982_13878.n70 47.835
R16683 a_n2982_13878.n145 a_n2982_13878.n62 47.835
R16684 a_n2982_13878.n3 a_n2982_13878.n2 1.59102
R16685 a_n2982_13878.n30 a_n2982_13878.n29 1.13686
R16686 a_n2982_13878.n19 a_n2982_13878.n18 1.13686
R16687 a_n2982_13878.n13 a_n2982_13878.n12 1.13686
R16688 a_n2982_13878.n35 a_n2982_13878.n24 1.09898
R16689 a_n2982_13878.n40 a_n2982_13878.n39 1.07378
R16690 a_n2982_13878.n37 a_n2982_13878.n36 1.07378
R16691 a_n2982_13878.n1 a_n2982_13878.n0 1.06084
R16692 a_n2982_13878.n33 a_n2982_13878.n32 0.758076
R16693 a_n2982_13878.n33 a_n2982_13878.n31 0.758076
R16694 a_n2982_13878.n31 a_n2982_13878.n30 0.758076
R16695 a_n2982_13878.n27 a_n2982_13878.n26 0.758076
R16696 a_n2982_13878.n27 a_n2982_13878.n25 0.758076
R16697 a_n2982_13878.n25 a_n2982_13878.n24 0.758076
R16698 a_n2982_13878.n21 a_n2982_13878.n22 0.758076
R16699 a_n2982_13878.n20 a_n2982_13878.n21 0.758076
R16700 a_n2982_13878.n18 a_n2982_13878.n20 0.758076
R16701 a_n2982_13878.n15 a_n2982_13878.n16 0.758076
R16702 a_n2982_13878.n14 a_n2982_13878.n15 0.758076
R16703 a_n2982_13878.n12 a_n2982_13878.n14 0.758076
R16704 a_n2982_13878.n11 a_n2982_13878.n10 0.758076
R16705 a_n2982_13878.n9 a_n2982_13878.n8 0.758076
R16706 a_n2982_13878.n7 a_n2982_13878.n6 0.758076
R16707 a_n2982_13878.n5 a_n2982_13878.n4 0.758076
R16708 a_n2982_13878.n39 a_n2982_13878.n41 0.716017
R16709 a_n2982_13878.n36 a_n2982_13878.n38 0.716017
R16710 a_n2982_13878.n10 a_n2982_13878.n9 0.67853
R16711 a_n2982_13878.n6 a_n2982_13878.n5 0.67853
R16712 a_n2804_13878.n29 a_n2804_13878.n28 98.9632
R16713 a_n2804_13878.n2 a_n2804_13878.n0 98.7517
R16714 a_n2804_13878.n22 a_n2804_13878.n21 98.6055
R16715 a_n2804_13878.n24 a_n2804_13878.n23 98.6055
R16716 a_n2804_13878.n26 a_n2804_13878.n25 98.6055
R16717 a_n2804_13878.n28 a_n2804_13878.n27 98.6055
R16718 a_n2804_13878.n10 a_n2804_13878.n9 98.6055
R16719 a_n2804_13878.n8 a_n2804_13878.n7 98.6055
R16720 a_n2804_13878.n6 a_n2804_13878.n5 98.6055
R16721 a_n2804_13878.n4 a_n2804_13878.n3 98.6055
R16722 a_n2804_13878.n2 a_n2804_13878.n1 98.6055
R16723 a_n2804_13878.n20 a_n2804_13878.n19 98.6054
R16724 a_n2804_13878.n12 a_n2804_13878.t2 74.6477
R16725 a_n2804_13878.n17 a_n2804_13878.t31 74.2899
R16726 a_n2804_13878.n14 a_n2804_13878.t4 74.2899
R16727 a_n2804_13878.n13 a_n2804_13878.t5 74.2899
R16728 a_n2804_13878.n16 a_n2804_13878.n15 70.6783
R16729 a_n2804_13878.n12 a_n2804_13878.n11 70.6783
R16730 a_n2804_13878.n18 a_n2804_13878.n10 15.7159
R16731 a_n2804_13878.n20 a_n2804_13878.n18 12.6495
R16732 a_n2804_13878.n18 a_n2804_13878.n17 8.38735
R16733 a_n2804_13878.n19 a_n2804_13878.t13 3.61217
R16734 a_n2804_13878.n19 a_n2804_13878.t22 3.61217
R16735 a_n2804_13878.n21 a_n2804_13878.t26 3.61217
R16736 a_n2804_13878.n21 a_n2804_13878.t12 3.61217
R16737 a_n2804_13878.n23 a_n2804_13878.t16 3.61217
R16738 a_n2804_13878.n23 a_n2804_13878.t17 3.61217
R16739 a_n2804_13878.n25 a_n2804_13878.t27 3.61217
R16740 a_n2804_13878.n25 a_n2804_13878.t28 3.61217
R16741 a_n2804_13878.n27 a_n2804_13878.t6 3.61217
R16742 a_n2804_13878.n27 a_n2804_13878.t18 3.61217
R16743 a_n2804_13878.n15 a_n2804_13878.t0 3.61217
R16744 a_n2804_13878.n15 a_n2804_13878.t3 3.61217
R16745 a_n2804_13878.n11 a_n2804_13878.t30 3.61217
R16746 a_n2804_13878.n11 a_n2804_13878.t1 3.61217
R16747 a_n2804_13878.n9 a_n2804_13878.t19 3.61217
R16748 a_n2804_13878.n9 a_n2804_13878.t7 3.61217
R16749 a_n2804_13878.n7 a_n2804_13878.t24 3.61217
R16750 a_n2804_13878.n7 a_n2804_13878.t9 3.61217
R16751 a_n2804_13878.n5 a_n2804_13878.t8 3.61217
R16752 a_n2804_13878.n5 a_n2804_13878.t11 3.61217
R16753 a_n2804_13878.n3 a_n2804_13878.t21 3.61217
R16754 a_n2804_13878.n3 a_n2804_13878.t14 3.61217
R16755 a_n2804_13878.n1 a_n2804_13878.t25 3.61217
R16756 a_n2804_13878.n1 a_n2804_13878.t15 3.61217
R16757 a_n2804_13878.n0 a_n2804_13878.t10 3.61217
R16758 a_n2804_13878.n0 a_n2804_13878.t20 3.61217
R16759 a_n2804_13878.n29 a_n2804_13878.t23 3.61217
R16760 a_n2804_13878.t29 a_n2804_13878.n29 3.61217
R16761 a_n2804_13878.n13 a_n2804_13878.n12 0.358259
R16762 a_n2804_13878.n16 a_n2804_13878.n14 0.358259
R16763 a_n2804_13878.n17 a_n2804_13878.n16 0.358259
R16764 a_n2804_13878.n28 a_n2804_13878.n26 0.358259
R16765 a_n2804_13878.n26 a_n2804_13878.n24 0.358259
R16766 a_n2804_13878.n24 a_n2804_13878.n22 0.358259
R16767 a_n2804_13878.n22 a_n2804_13878.n20 0.358259
R16768 a_n2804_13878.n4 a_n2804_13878.n2 0.146627
R16769 a_n2804_13878.n6 a_n2804_13878.n4 0.146627
R16770 a_n2804_13878.n8 a_n2804_13878.n6 0.146627
R16771 a_n2804_13878.n10 a_n2804_13878.n8 0.146627
R16772 a_n2804_13878.n14 a_n2804_13878.n13 0.101793
R16773 vdd.n303 vdd.n267 756.745
R16774 vdd.n252 vdd.n216 756.745
R16775 vdd.n209 vdd.n173 756.745
R16776 vdd.n158 vdd.n122 756.745
R16777 vdd.n116 vdd.n80 756.745
R16778 vdd.n65 vdd.n29 756.745
R16779 vdd.n1953 vdd.n1917 756.745
R16780 vdd.n2004 vdd.n1968 756.745
R16781 vdd.n1859 vdd.n1823 756.745
R16782 vdd.n1910 vdd.n1874 756.745
R16783 vdd.n1766 vdd.n1730 756.745
R16784 vdd.n1817 vdd.n1781 756.745
R16785 vdd.n1143 vdd.t28 640.208
R16786 vdd.n838 vdd.t73 640.208
R16787 vdd.n1147 vdd.t70 640.208
R16788 vdd.n829 vdd.t97 640.208
R16789 vdd.n724 vdd.t50 640.208
R16790 vdd.n2535 vdd.t91 640.208
R16791 vdd.n661 vdd.t39 640.208
R16792 vdd.n2532 vdd.t80 640.208
R16793 vdd.n625 vdd.t24 640.208
R16794 vdd.n899 vdd.t87 640.208
R16795 vdd.n1565 vdd.t60 592.009
R16796 vdd.n1602 vdd.t84 592.009
R16797 vdd.n1476 vdd.t94 592.009
R16798 vdd.n2074 vdd.t54 592.009
R16799 vdd.n1076 vdd.t32 592.009
R16800 vdd.n1036 vdd.t36 592.009
R16801 vdd.n3293 vdd.t57 592.009
R16802 vdd.n427 vdd.t46 592.009
R16803 vdd.n387 vdd.t64 592.009
R16804 vdd.n580 vdd.t67 592.009
R16805 vdd.n543 vdd.t77 592.009
R16806 vdd.n3080 vdd.t42 592.009
R16807 vdd.n304 vdd.n303 585
R16808 vdd.n302 vdd.n269 585
R16809 vdd.n301 vdd.n300 585
R16810 vdd.n272 vdd.n270 585
R16811 vdd.n295 vdd.n294 585
R16812 vdd.n293 vdd.n292 585
R16813 vdd.n276 vdd.n275 585
R16814 vdd.n287 vdd.n286 585
R16815 vdd.n285 vdd.n284 585
R16816 vdd.n280 vdd.n279 585
R16817 vdd.n253 vdd.n252 585
R16818 vdd.n251 vdd.n218 585
R16819 vdd.n250 vdd.n249 585
R16820 vdd.n221 vdd.n219 585
R16821 vdd.n244 vdd.n243 585
R16822 vdd.n242 vdd.n241 585
R16823 vdd.n225 vdd.n224 585
R16824 vdd.n236 vdd.n235 585
R16825 vdd.n234 vdd.n233 585
R16826 vdd.n229 vdd.n228 585
R16827 vdd.n210 vdd.n209 585
R16828 vdd.n208 vdd.n175 585
R16829 vdd.n207 vdd.n206 585
R16830 vdd.n178 vdd.n176 585
R16831 vdd.n201 vdd.n200 585
R16832 vdd.n199 vdd.n198 585
R16833 vdd.n182 vdd.n181 585
R16834 vdd.n193 vdd.n192 585
R16835 vdd.n191 vdd.n190 585
R16836 vdd.n186 vdd.n185 585
R16837 vdd.n159 vdd.n158 585
R16838 vdd.n157 vdd.n124 585
R16839 vdd.n156 vdd.n155 585
R16840 vdd.n127 vdd.n125 585
R16841 vdd.n150 vdd.n149 585
R16842 vdd.n148 vdd.n147 585
R16843 vdd.n131 vdd.n130 585
R16844 vdd.n142 vdd.n141 585
R16845 vdd.n140 vdd.n139 585
R16846 vdd.n135 vdd.n134 585
R16847 vdd.n117 vdd.n116 585
R16848 vdd.n115 vdd.n82 585
R16849 vdd.n114 vdd.n113 585
R16850 vdd.n85 vdd.n83 585
R16851 vdd.n108 vdd.n107 585
R16852 vdd.n106 vdd.n105 585
R16853 vdd.n89 vdd.n88 585
R16854 vdd.n100 vdd.n99 585
R16855 vdd.n98 vdd.n97 585
R16856 vdd.n93 vdd.n92 585
R16857 vdd.n66 vdd.n65 585
R16858 vdd.n64 vdd.n31 585
R16859 vdd.n63 vdd.n62 585
R16860 vdd.n34 vdd.n32 585
R16861 vdd.n57 vdd.n56 585
R16862 vdd.n55 vdd.n54 585
R16863 vdd.n38 vdd.n37 585
R16864 vdd.n49 vdd.n48 585
R16865 vdd.n47 vdd.n46 585
R16866 vdd.n42 vdd.n41 585
R16867 vdd.n1954 vdd.n1953 585
R16868 vdd.n1952 vdd.n1919 585
R16869 vdd.n1951 vdd.n1950 585
R16870 vdd.n1922 vdd.n1920 585
R16871 vdd.n1945 vdd.n1944 585
R16872 vdd.n1943 vdd.n1942 585
R16873 vdd.n1926 vdd.n1925 585
R16874 vdd.n1937 vdd.n1936 585
R16875 vdd.n1935 vdd.n1934 585
R16876 vdd.n1930 vdd.n1929 585
R16877 vdd.n2005 vdd.n2004 585
R16878 vdd.n2003 vdd.n1970 585
R16879 vdd.n2002 vdd.n2001 585
R16880 vdd.n1973 vdd.n1971 585
R16881 vdd.n1996 vdd.n1995 585
R16882 vdd.n1994 vdd.n1993 585
R16883 vdd.n1977 vdd.n1976 585
R16884 vdd.n1988 vdd.n1987 585
R16885 vdd.n1986 vdd.n1985 585
R16886 vdd.n1981 vdd.n1980 585
R16887 vdd.n1860 vdd.n1859 585
R16888 vdd.n1858 vdd.n1825 585
R16889 vdd.n1857 vdd.n1856 585
R16890 vdd.n1828 vdd.n1826 585
R16891 vdd.n1851 vdd.n1850 585
R16892 vdd.n1849 vdd.n1848 585
R16893 vdd.n1832 vdd.n1831 585
R16894 vdd.n1843 vdd.n1842 585
R16895 vdd.n1841 vdd.n1840 585
R16896 vdd.n1836 vdd.n1835 585
R16897 vdd.n1911 vdd.n1910 585
R16898 vdd.n1909 vdd.n1876 585
R16899 vdd.n1908 vdd.n1907 585
R16900 vdd.n1879 vdd.n1877 585
R16901 vdd.n1902 vdd.n1901 585
R16902 vdd.n1900 vdd.n1899 585
R16903 vdd.n1883 vdd.n1882 585
R16904 vdd.n1894 vdd.n1893 585
R16905 vdd.n1892 vdd.n1891 585
R16906 vdd.n1887 vdd.n1886 585
R16907 vdd.n1767 vdd.n1766 585
R16908 vdd.n1765 vdd.n1732 585
R16909 vdd.n1764 vdd.n1763 585
R16910 vdd.n1735 vdd.n1733 585
R16911 vdd.n1758 vdd.n1757 585
R16912 vdd.n1756 vdd.n1755 585
R16913 vdd.n1739 vdd.n1738 585
R16914 vdd.n1750 vdd.n1749 585
R16915 vdd.n1748 vdd.n1747 585
R16916 vdd.n1743 vdd.n1742 585
R16917 vdd.n1818 vdd.n1817 585
R16918 vdd.n1816 vdd.n1783 585
R16919 vdd.n1815 vdd.n1814 585
R16920 vdd.n1786 vdd.n1784 585
R16921 vdd.n1809 vdd.n1808 585
R16922 vdd.n1807 vdd.n1806 585
R16923 vdd.n1790 vdd.n1789 585
R16924 vdd.n1801 vdd.n1800 585
R16925 vdd.n1799 vdd.n1798 585
R16926 vdd.n1794 vdd.n1793 585
R16927 vdd.n3409 vdd.n352 488.781
R16928 vdd.n3291 vdd.n350 488.781
R16929 vdd.n3213 vdd.n515 488.781
R16930 vdd.n3211 vdd.n517 488.781
R16931 vdd.n2069 vdd.n1358 488.781
R16932 vdd.n2072 vdd.n2071 488.781
R16933 vdd.n1671 vdd.n1436 488.781
R16934 vdd.n1669 vdd.n1439 488.781
R16935 vdd.n281 vdd.t144 329.043
R16936 vdd.n230 vdd.t3 329.043
R16937 vdd.n187 vdd.t23 329.043
R16938 vdd.n136 vdd.t219 329.043
R16939 vdd.n94 vdd.t154 329.043
R16940 vdd.n43 vdd.t16 329.043
R16941 vdd.n1931 vdd.t220 329.043
R16942 vdd.n1982 vdd.t132 329.043
R16943 vdd.n1837 vdd.t102 329.043
R16944 vdd.n1888 vdd.t153 329.043
R16945 vdd.n1744 vdd.t15 329.043
R16946 vdd.n1795 vdd.t240 329.043
R16947 vdd.n1565 vdd.t63 319.788
R16948 vdd.n1602 vdd.t86 319.788
R16949 vdd.n1476 vdd.t96 319.788
R16950 vdd.n2074 vdd.t55 319.788
R16951 vdd.n1076 vdd.t34 319.788
R16952 vdd.n1036 vdd.t37 319.788
R16953 vdd.n3293 vdd.t58 319.788
R16954 vdd.n427 vdd.t48 319.788
R16955 vdd.n387 vdd.t65 319.788
R16956 vdd.n580 vdd.t69 319.788
R16957 vdd.n543 vdd.t79 319.788
R16958 vdd.n3080 vdd.t45 319.788
R16959 vdd.n1566 vdd.t62 303.69
R16960 vdd.n1603 vdd.t85 303.69
R16961 vdd.n1477 vdd.t95 303.69
R16962 vdd.n2075 vdd.t56 303.69
R16963 vdd.n1077 vdd.t35 303.69
R16964 vdd.n1037 vdd.t38 303.69
R16965 vdd.n3294 vdd.t59 303.69
R16966 vdd.n428 vdd.t49 303.69
R16967 vdd.n388 vdd.t66 303.69
R16968 vdd.n581 vdd.t68 303.69
R16969 vdd.n544 vdd.t78 303.69
R16970 vdd.n3081 vdd.t44 303.69
R16971 vdd.n2802 vdd.n788 279.512
R16972 vdd.n3042 vdd.n635 279.512
R16973 vdd.n2979 vdd.n632 279.512
R16974 vdd.n2734 vdd.n2733 279.512
R16975 vdd.n2495 vdd.n826 279.512
R16976 vdd.n2426 vdd.n2425 279.512
R16977 vdd.n1183 vdd.n1182 279.512
R16978 vdd.n2220 vdd.n966 279.512
R16979 vdd.n2958 vdd.n633 279.512
R16980 vdd.n3045 vdd.n3044 279.512
R16981 vdd.n2607 vdd.n2530 279.512
R16982 vdd.n2538 vdd.n784 279.512
R16983 vdd.n2423 vdd.n836 279.512
R16984 vdd.n834 vdd.n808 279.512
R16985 vdd.n1308 vdd.n1003 279.512
R16986 vdd.n1108 vdd.n961 279.512
R16987 vdd.n2218 vdd.n969 254.619
R16988 vdd.n613 vdd.n516 254.619
R16989 vdd.n2960 vdd.n633 185
R16990 vdd.n3043 vdd.n633 185
R16991 vdd.n2962 vdd.n2961 185
R16992 vdd.n2961 vdd.n631 185
R16993 vdd.n2963 vdd.n667 185
R16994 vdd.n2973 vdd.n667 185
R16995 vdd.n2964 vdd.n676 185
R16996 vdd.n676 vdd.n674 185
R16997 vdd.n2966 vdd.n2965 185
R16998 vdd.n2967 vdd.n2966 185
R16999 vdd.n2919 vdd.n675 185
R17000 vdd.n675 vdd.n671 185
R17001 vdd.n2918 vdd.n2917 185
R17002 vdd.n2917 vdd.n2916 185
R17003 vdd.n678 vdd.n677 185
R17004 vdd.n679 vdd.n678 185
R17005 vdd.n2909 vdd.n2908 185
R17006 vdd.n2910 vdd.n2909 185
R17007 vdd.n2907 vdd.n687 185
R17008 vdd.n692 vdd.n687 185
R17009 vdd.n2906 vdd.n2905 185
R17010 vdd.n2905 vdd.n2904 185
R17011 vdd.n689 vdd.n688 185
R17012 vdd.n698 vdd.n689 185
R17013 vdd.n2897 vdd.n2896 185
R17014 vdd.n2898 vdd.n2897 185
R17015 vdd.n2895 vdd.n699 185
R17016 vdd.n705 vdd.n699 185
R17017 vdd.n2894 vdd.n2893 185
R17018 vdd.n2893 vdd.n2892 185
R17019 vdd.n701 vdd.n700 185
R17020 vdd.n702 vdd.n701 185
R17021 vdd.n2885 vdd.n2884 185
R17022 vdd.n2886 vdd.n2885 185
R17023 vdd.n2883 vdd.n712 185
R17024 vdd.n712 vdd.n709 185
R17025 vdd.n2882 vdd.n2881 185
R17026 vdd.n2881 vdd.n2880 185
R17027 vdd.n714 vdd.n713 185
R17028 vdd.n715 vdd.n714 185
R17029 vdd.n2873 vdd.n2872 185
R17030 vdd.n2874 vdd.n2873 185
R17031 vdd.n2871 vdd.n723 185
R17032 vdd.n729 vdd.n723 185
R17033 vdd.n2870 vdd.n2869 185
R17034 vdd.n2869 vdd.n2868 185
R17035 vdd.n2859 vdd.n726 185
R17036 vdd.n736 vdd.n726 185
R17037 vdd.n2861 vdd.n2860 185
R17038 vdd.n2862 vdd.n2861 185
R17039 vdd.n2858 vdd.n737 185
R17040 vdd.n737 vdd.n733 185
R17041 vdd.n2857 vdd.n2856 185
R17042 vdd.n2856 vdd.n2855 185
R17043 vdd.n739 vdd.n738 185
R17044 vdd.n740 vdd.n739 185
R17045 vdd.n2848 vdd.n2847 185
R17046 vdd.n2849 vdd.n2848 185
R17047 vdd.n2846 vdd.n748 185
R17048 vdd.n753 vdd.n748 185
R17049 vdd.n2845 vdd.n2844 185
R17050 vdd.n2844 vdd.n2843 185
R17051 vdd.n750 vdd.n749 185
R17052 vdd.n759 vdd.n750 185
R17053 vdd.n2836 vdd.n2835 185
R17054 vdd.n2837 vdd.n2836 185
R17055 vdd.n2834 vdd.n760 185
R17056 vdd.n2710 vdd.n760 185
R17057 vdd.n2833 vdd.n2832 185
R17058 vdd.n2832 vdd.n2831 185
R17059 vdd.n762 vdd.n761 185
R17060 vdd.n2716 vdd.n762 185
R17061 vdd.n2824 vdd.n2823 185
R17062 vdd.n2825 vdd.n2824 185
R17063 vdd.n2822 vdd.n771 185
R17064 vdd.n771 vdd.n768 185
R17065 vdd.n2821 vdd.n2820 185
R17066 vdd.n2820 vdd.n2819 185
R17067 vdd.n773 vdd.n772 185
R17068 vdd.n774 vdd.n773 185
R17069 vdd.n2812 vdd.n2811 185
R17070 vdd.n2813 vdd.n2812 185
R17071 vdd.n2810 vdd.n782 185
R17072 vdd.n2728 vdd.n782 185
R17073 vdd.n2809 vdd.n2808 185
R17074 vdd.n2808 vdd.n2807 185
R17075 vdd.n784 vdd.n783 185
R17076 vdd.n785 vdd.n784 185
R17077 vdd.n2539 vdd.n2538 185
R17078 vdd.n2541 vdd.n2540 185
R17079 vdd.n2543 vdd.n2542 185
R17080 vdd.n2545 vdd.n2544 185
R17081 vdd.n2547 vdd.n2546 185
R17082 vdd.n2549 vdd.n2548 185
R17083 vdd.n2551 vdd.n2550 185
R17084 vdd.n2553 vdd.n2552 185
R17085 vdd.n2555 vdd.n2554 185
R17086 vdd.n2557 vdd.n2556 185
R17087 vdd.n2559 vdd.n2558 185
R17088 vdd.n2561 vdd.n2560 185
R17089 vdd.n2563 vdd.n2562 185
R17090 vdd.n2565 vdd.n2564 185
R17091 vdd.n2567 vdd.n2566 185
R17092 vdd.n2569 vdd.n2568 185
R17093 vdd.n2571 vdd.n2570 185
R17094 vdd.n2573 vdd.n2572 185
R17095 vdd.n2575 vdd.n2574 185
R17096 vdd.n2577 vdd.n2576 185
R17097 vdd.n2579 vdd.n2578 185
R17098 vdd.n2581 vdd.n2580 185
R17099 vdd.n2583 vdd.n2582 185
R17100 vdd.n2585 vdd.n2584 185
R17101 vdd.n2587 vdd.n2586 185
R17102 vdd.n2589 vdd.n2588 185
R17103 vdd.n2591 vdd.n2590 185
R17104 vdd.n2593 vdd.n2592 185
R17105 vdd.n2595 vdd.n2594 185
R17106 vdd.n2597 vdd.n2596 185
R17107 vdd.n2599 vdd.n2598 185
R17108 vdd.n2601 vdd.n2600 185
R17109 vdd.n2603 vdd.n2602 185
R17110 vdd.n2605 vdd.n2604 185
R17111 vdd.n2606 vdd.n2530 185
R17112 vdd.n2800 vdd.n2530 185
R17113 vdd.n3046 vdd.n3045 185
R17114 vdd.n3047 vdd.n624 185
R17115 vdd.n3049 vdd.n3048 185
R17116 vdd.n3051 vdd.n622 185
R17117 vdd.n3053 vdd.n3052 185
R17118 vdd.n3054 vdd.n621 185
R17119 vdd.n3056 vdd.n3055 185
R17120 vdd.n3058 vdd.n619 185
R17121 vdd.n3060 vdd.n3059 185
R17122 vdd.n3061 vdd.n618 185
R17123 vdd.n3063 vdd.n3062 185
R17124 vdd.n3065 vdd.n616 185
R17125 vdd.n3067 vdd.n3066 185
R17126 vdd.n3068 vdd.n615 185
R17127 vdd.n3070 vdd.n3069 185
R17128 vdd.n3072 vdd.n614 185
R17129 vdd.n3073 vdd.n611 185
R17130 vdd.n3076 vdd.n3075 185
R17131 vdd.n612 vdd.n610 185
R17132 vdd.n2932 vdd.n2931 185
R17133 vdd.n2934 vdd.n2933 185
R17134 vdd.n2936 vdd.n2928 185
R17135 vdd.n2938 vdd.n2937 185
R17136 vdd.n2939 vdd.n2927 185
R17137 vdd.n2941 vdd.n2940 185
R17138 vdd.n2943 vdd.n2925 185
R17139 vdd.n2945 vdd.n2944 185
R17140 vdd.n2946 vdd.n2924 185
R17141 vdd.n2948 vdd.n2947 185
R17142 vdd.n2950 vdd.n2922 185
R17143 vdd.n2952 vdd.n2951 185
R17144 vdd.n2953 vdd.n2921 185
R17145 vdd.n2955 vdd.n2954 185
R17146 vdd.n2957 vdd.n2920 185
R17147 vdd.n2959 vdd.n2958 185
R17148 vdd.n2958 vdd.n613 185
R17149 vdd.n3044 vdd.n628 185
R17150 vdd.n3044 vdd.n3043 185
R17151 vdd.n2661 vdd.n630 185
R17152 vdd.n631 vdd.n630 185
R17153 vdd.n2662 vdd.n666 185
R17154 vdd.n2973 vdd.n666 185
R17155 vdd.n2664 vdd.n2663 185
R17156 vdd.n2663 vdd.n674 185
R17157 vdd.n2665 vdd.n673 185
R17158 vdd.n2967 vdd.n673 185
R17159 vdd.n2667 vdd.n2666 185
R17160 vdd.n2666 vdd.n671 185
R17161 vdd.n2668 vdd.n681 185
R17162 vdd.n2916 vdd.n681 185
R17163 vdd.n2670 vdd.n2669 185
R17164 vdd.n2669 vdd.n679 185
R17165 vdd.n2671 vdd.n686 185
R17166 vdd.n2910 vdd.n686 185
R17167 vdd.n2673 vdd.n2672 185
R17168 vdd.n2672 vdd.n692 185
R17169 vdd.n2674 vdd.n691 185
R17170 vdd.n2904 vdd.n691 185
R17171 vdd.n2676 vdd.n2675 185
R17172 vdd.n2675 vdd.n698 185
R17173 vdd.n2677 vdd.n697 185
R17174 vdd.n2898 vdd.n697 185
R17175 vdd.n2679 vdd.n2678 185
R17176 vdd.n2678 vdd.n705 185
R17177 vdd.n2680 vdd.n704 185
R17178 vdd.n2892 vdd.n704 185
R17179 vdd.n2682 vdd.n2681 185
R17180 vdd.n2681 vdd.n702 185
R17181 vdd.n2683 vdd.n711 185
R17182 vdd.n2886 vdd.n711 185
R17183 vdd.n2685 vdd.n2684 185
R17184 vdd.n2684 vdd.n709 185
R17185 vdd.n2686 vdd.n717 185
R17186 vdd.n2880 vdd.n717 185
R17187 vdd.n2688 vdd.n2687 185
R17188 vdd.n2687 vdd.n715 185
R17189 vdd.n2689 vdd.n722 185
R17190 vdd.n2874 vdd.n722 185
R17191 vdd.n2691 vdd.n2690 185
R17192 vdd.n2690 vdd.n729 185
R17193 vdd.n2692 vdd.n728 185
R17194 vdd.n2868 vdd.n728 185
R17195 vdd.n2694 vdd.n2693 185
R17196 vdd.n2693 vdd.n736 185
R17197 vdd.n2695 vdd.n735 185
R17198 vdd.n2862 vdd.n735 185
R17199 vdd.n2697 vdd.n2696 185
R17200 vdd.n2696 vdd.n733 185
R17201 vdd.n2698 vdd.n742 185
R17202 vdd.n2855 vdd.n742 185
R17203 vdd.n2700 vdd.n2699 185
R17204 vdd.n2699 vdd.n740 185
R17205 vdd.n2701 vdd.n747 185
R17206 vdd.n2849 vdd.n747 185
R17207 vdd.n2703 vdd.n2702 185
R17208 vdd.n2702 vdd.n753 185
R17209 vdd.n2704 vdd.n752 185
R17210 vdd.n2843 vdd.n752 185
R17211 vdd.n2706 vdd.n2705 185
R17212 vdd.n2705 vdd.n759 185
R17213 vdd.n2707 vdd.n758 185
R17214 vdd.n2837 vdd.n758 185
R17215 vdd.n2709 vdd.n2708 185
R17216 vdd.n2710 vdd.n2709 185
R17217 vdd.n2610 vdd.n764 185
R17218 vdd.n2831 vdd.n764 185
R17219 vdd.n2718 vdd.n2717 185
R17220 vdd.n2717 vdd.n2716 185
R17221 vdd.n2719 vdd.n770 185
R17222 vdd.n2825 vdd.n770 185
R17223 vdd.n2721 vdd.n2720 185
R17224 vdd.n2720 vdd.n768 185
R17225 vdd.n2722 vdd.n776 185
R17226 vdd.n2819 vdd.n776 185
R17227 vdd.n2724 vdd.n2723 185
R17228 vdd.n2723 vdd.n774 185
R17229 vdd.n2725 vdd.n781 185
R17230 vdd.n2813 vdd.n781 185
R17231 vdd.n2727 vdd.n2726 185
R17232 vdd.n2728 vdd.n2727 185
R17233 vdd.n2609 vdd.n787 185
R17234 vdd.n2807 vdd.n787 185
R17235 vdd.n2608 vdd.n2607 185
R17236 vdd.n2607 vdd.n785 185
R17237 vdd.n2069 vdd.n2068 185
R17238 vdd.n2070 vdd.n2069 185
R17239 vdd.n1359 vdd.n1357 185
R17240 vdd.n2061 vdd.n1357 185
R17241 vdd.n2064 vdd.n2063 185
R17242 vdd.n2063 vdd.n2062 185
R17243 vdd.n1362 vdd.n1361 185
R17244 vdd.n1363 vdd.n1362 185
R17245 vdd.n2050 vdd.n2049 185
R17246 vdd.n2051 vdd.n2050 185
R17247 vdd.n1371 vdd.n1370 185
R17248 vdd.n2042 vdd.n1370 185
R17249 vdd.n2045 vdd.n2044 185
R17250 vdd.n2044 vdd.n2043 185
R17251 vdd.n1374 vdd.n1373 185
R17252 vdd.n1380 vdd.n1374 185
R17253 vdd.n2033 vdd.n2032 185
R17254 vdd.n2034 vdd.n2033 185
R17255 vdd.n1382 vdd.n1381 185
R17256 vdd.n2025 vdd.n1381 185
R17257 vdd.n2028 vdd.n2027 185
R17258 vdd.n2027 vdd.n2026 185
R17259 vdd.n1385 vdd.n1384 185
R17260 vdd.n1386 vdd.n1385 185
R17261 vdd.n2016 vdd.n2015 185
R17262 vdd.n2017 vdd.n2016 185
R17263 vdd.n1394 vdd.n1393 185
R17264 vdd.n1393 vdd.n1392 185
R17265 vdd.n1729 vdd.n1728 185
R17266 vdd.n1728 vdd.n1727 185
R17267 vdd.n1397 vdd.n1396 185
R17268 vdd.n1403 vdd.n1397 185
R17269 vdd.n1718 vdd.n1717 185
R17270 vdd.n1719 vdd.n1718 185
R17271 vdd.n1405 vdd.n1404 185
R17272 vdd.n1710 vdd.n1404 185
R17273 vdd.n1713 vdd.n1712 185
R17274 vdd.n1712 vdd.n1711 185
R17275 vdd.n1408 vdd.n1407 185
R17276 vdd.n1415 vdd.n1408 185
R17277 vdd.n1701 vdd.n1700 185
R17278 vdd.n1702 vdd.n1701 185
R17279 vdd.n1417 vdd.n1416 185
R17280 vdd.n1416 vdd.n1414 185
R17281 vdd.n1696 vdd.n1695 185
R17282 vdd.n1695 vdd.n1694 185
R17283 vdd.n1420 vdd.n1419 185
R17284 vdd.n1421 vdd.n1420 185
R17285 vdd.n1685 vdd.n1684 185
R17286 vdd.n1686 vdd.n1685 185
R17287 vdd.n1429 vdd.n1428 185
R17288 vdd.n1428 vdd.n1427 185
R17289 vdd.n1680 vdd.n1679 185
R17290 vdd.n1679 vdd.n1678 185
R17291 vdd.n1432 vdd.n1431 185
R17292 vdd.n1438 vdd.n1432 185
R17293 vdd.n1669 vdd.n1668 185
R17294 vdd.n1670 vdd.n1669 185
R17295 vdd.n1665 vdd.n1439 185
R17296 vdd.n1664 vdd.n1442 185
R17297 vdd.n1663 vdd.n1443 185
R17298 vdd.n1443 vdd.n1437 185
R17299 vdd.n1446 vdd.n1444 185
R17300 vdd.n1659 vdd.n1448 185
R17301 vdd.n1658 vdd.n1449 185
R17302 vdd.n1657 vdd.n1451 185
R17303 vdd.n1454 vdd.n1452 185
R17304 vdd.n1653 vdd.n1456 185
R17305 vdd.n1652 vdd.n1457 185
R17306 vdd.n1651 vdd.n1459 185
R17307 vdd.n1462 vdd.n1460 185
R17308 vdd.n1647 vdd.n1464 185
R17309 vdd.n1646 vdd.n1465 185
R17310 vdd.n1645 vdd.n1467 185
R17311 vdd.n1470 vdd.n1468 185
R17312 vdd.n1641 vdd.n1472 185
R17313 vdd.n1640 vdd.n1473 185
R17314 vdd.n1639 vdd.n1475 185
R17315 vdd.n1480 vdd.n1478 185
R17316 vdd.n1635 vdd.n1482 185
R17317 vdd.n1634 vdd.n1483 185
R17318 vdd.n1633 vdd.n1485 185
R17319 vdd.n1488 vdd.n1486 185
R17320 vdd.n1629 vdd.n1490 185
R17321 vdd.n1628 vdd.n1491 185
R17322 vdd.n1627 vdd.n1493 185
R17323 vdd.n1496 vdd.n1494 185
R17324 vdd.n1623 vdd.n1498 185
R17325 vdd.n1622 vdd.n1499 185
R17326 vdd.n1621 vdd.n1501 185
R17327 vdd.n1504 vdd.n1502 185
R17328 vdd.n1617 vdd.n1506 185
R17329 vdd.n1616 vdd.n1507 185
R17330 vdd.n1615 vdd.n1509 185
R17331 vdd.n1512 vdd.n1510 185
R17332 vdd.n1611 vdd.n1514 185
R17333 vdd.n1610 vdd.n1515 185
R17334 vdd.n1609 vdd.n1517 185
R17335 vdd.n1520 vdd.n1518 185
R17336 vdd.n1605 vdd.n1522 185
R17337 vdd.n1604 vdd.n1601 185
R17338 vdd.n1599 vdd.n1523 185
R17339 vdd.n1598 vdd.n1597 185
R17340 vdd.n1528 vdd.n1525 185
R17341 vdd.n1593 vdd.n1529 185
R17342 vdd.n1592 vdd.n1531 185
R17343 vdd.n1591 vdd.n1532 185
R17344 vdd.n1536 vdd.n1533 185
R17345 vdd.n1587 vdd.n1537 185
R17346 vdd.n1586 vdd.n1539 185
R17347 vdd.n1585 vdd.n1540 185
R17348 vdd.n1544 vdd.n1541 185
R17349 vdd.n1581 vdd.n1545 185
R17350 vdd.n1580 vdd.n1547 185
R17351 vdd.n1579 vdd.n1548 185
R17352 vdd.n1552 vdd.n1549 185
R17353 vdd.n1575 vdd.n1553 185
R17354 vdd.n1574 vdd.n1555 185
R17355 vdd.n1573 vdd.n1556 185
R17356 vdd.n1560 vdd.n1557 185
R17357 vdd.n1569 vdd.n1561 185
R17358 vdd.n1568 vdd.n1563 185
R17359 vdd.n1564 vdd.n1436 185
R17360 vdd.n1437 vdd.n1436 185
R17361 vdd.n2073 vdd.n2072 185
R17362 vdd.n2077 vdd.n1353 185
R17363 vdd.n1352 vdd.n1346 185
R17364 vdd.n1350 vdd.n1349 185
R17365 vdd.n1348 vdd.n1107 185
R17366 vdd.n2081 vdd.n1104 185
R17367 vdd.n2083 vdd.n2082 185
R17368 vdd.n2085 vdd.n1102 185
R17369 vdd.n2087 vdd.n2086 185
R17370 vdd.n2088 vdd.n1097 185
R17371 vdd.n2090 vdd.n2089 185
R17372 vdd.n2092 vdd.n1095 185
R17373 vdd.n2094 vdd.n2093 185
R17374 vdd.n2095 vdd.n1090 185
R17375 vdd.n2097 vdd.n2096 185
R17376 vdd.n2099 vdd.n1088 185
R17377 vdd.n2101 vdd.n2100 185
R17378 vdd.n2102 vdd.n1084 185
R17379 vdd.n2104 vdd.n2103 185
R17380 vdd.n2106 vdd.n1081 185
R17381 vdd.n2108 vdd.n2107 185
R17382 vdd.n1082 vdd.n1075 185
R17383 vdd.n2112 vdd.n1079 185
R17384 vdd.n2113 vdd.n1071 185
R17385 vdd.n2115 vdd.n2114 185
R17386 vdd.n2117 vdd.n1069 185
R17387 vdd.n2119 vdd.n2118 185
R17388 vdd.n2120 vdd.n1064 185
R17389 vdd.n2122 vdd.n2121 185
R17390 vdd.n2124 vdd.n1062 185
R17391 vdd.n2126 vdd.n2125 185
R17392 vdd.n2127 vdd.n1057 185
R17393 vdd.n2129 vdd.n2128 185
R17394 vdd.n2131 vdd.n1055 185
R17395 vdd.n2133 vdd.n2132 185
R17396 vdd.n2134 vdd.n1050 185
R17397 vdd.n2136 vdd.n2135 185
R17398 vdd.n2138 vdd.n1048 185
R17399 vdd.n2140 vdd.n2139 185
R17400 vdd.n2141 vdd.n1044 185
R17401 vdd.n2143 vdd.n2142 185
R17402 vdd.n2145 vdd.n1041 185
R17403 vdd.n2147 vdd.n2146 185
R17404 vdd.n1042 vdd.n1035 185
R17405 vdd.n2151 vdd.n1039 185
R17406 vdd.n2152 vdd.n1031 185
R17407 vdd.n2154 vdd.n2153 185
R17408 vdd.n2156 vdd.n1029 185
R17409 vdd.n2158 vdd.n2157 185
R17410 vdd.n2159 vdd.n1024 185
R17411 vdd.n2161 vdd.n2160 185
R17412 vdd.n2163 vdd.n1022 185
R17413 vdd.n2165 vdd.n2164 185
R17414 vdd.n2166 vdd.n1017 185
R17415 vdd.n2168 vdd.n2167 185
R17416 vdd.n2170 vdd.n1015 185
R17417 vdd.n2172 vdd.n2171 185
R17418 vdd.n2173 vdd.n1013 185
R17419 vdd.n2175 vdd.n2174 185
R17420 vdd.n2178 vdd.n2177 185
R17421 vdd.n2180 vdd.n2179 185
R17422 vdd.n2182 vdd.n1011 185
R17423 vdd.n2184 vdd.n2183 185
R17424 vdd.n1358 vdd.n1010 185
R17425 vdd.n2071 vdd.n1356 185
R17426 vdd.n2071 vdd.n2070 185
R17427 vdd.n1366 vdd.n1355 185
R17428 vdd.n2061 vdd.n1355 185
R17429 vdd.n2060 vdd.n2059 185
R17430 vdd.n2062 vdd.n2060 185
R17431 vdd.n1365 vdd.n1364 185
R17432 vdd.n1364 vdd.n1363 185
R17433 vdd.n2053 vdd.n2052 185
R17434 vdd.n2052 vdd.n2051 185
R17435 vdd.n1369 vdd.n1368 185
R17436 vdd.n2042 vdd.n1369 185
R17437 vdd.n2041 vdd.n2040 185
R17438 vdd.n2043 vdd.n2041 185
R17439 vdd.n1376 vdd.n1375 185
R17440 vdd.n1380 vdd.n1375 185
R17441 vdd.n2036 vdd.n2035 185
R17442 vdd.n2035 vdd.n2034 185
R17443 vdd.n1379 vdd.n1378 185
R17444 vdd.n2025 vdd.n1379 185
R17445 vdd.n2024 vdd.n2023 185
R17446 vdd.n2026 vdd.n2024 185
R17447 vdd.n1388 vdd.n1387 185
R17448 vdd.n1387 vdd.n1386 185
R17449 vdd.n2019 vdd.n2018 185
R17450 vdd.n2018 vdd.n2017 185
R17451 vdd.n1391 vdd.n1390 185
R17452 vdd.n1392 vdd.n1391 185
R17453 vdd.n1726 vdd.n1725 185
R17454 vdd.n1727 vdd.n1726 185
R17455 vdd.n1399 vdd.n1398 185
R17456 vdd.n1403 vdd.n1398 185
R17457 vdd.n1721 vdd.n1720 185
R17458 vdd.n1720 vdd.n1719 185
R17459 vdd.n1402 vdd.n1401 185
R17460 vdd.n1710 vdd.n1402 185
R17461 vdd.n1709 vdd.n1708 185
R17462 vdd.n1711 vdd.n1709 185
R17463 vdd.n1410 vdd.n1409 185
R17464 vdd.n1415 vdd.n1409 185
R17465 vdd.n1704 vdd.n1703 185
R17466 vdd.n1703 vdd.n1702 185
R17467 vdd.n1413 vdd.n1412 185
R17468 vdd.n1414 vdd.n1413 185
R17469 vdd.n1693 vdd.n1692 185
R17470 vdd.n1694 vdd.n1693 185
R17471 vdd.n1423 vdd.n1422 185
R17472 vdd.n1422 vdd.n1421 185
R17473 vdd.n1688 vdd.n1687 185
R17474 vdd.n1687 vdd.n1686 185
R17475 vdd.n1426 vdd.n1425 185
R17476 vdd.n1427 vdd.n1426 185
R17477 vdd.n1677 vdd.n1676 185
R17478 vdd.n1678 vdd.n1677 185
R17479 vdd.n1434 vdd.n1433 185
R17480 vdd.n1438 vdd.n1433 185
R17481 vdd.n1672 vdd.n1671 185
R17482 vdd.n1671 vdd.n1670 185
R17483 vdd.n828 vdd.n826 185
R17484 vdd.n2424 vdd.n826 185
R17485 vdd.n2346 vdd.n846 185
R17486 vdd.n846 vdd.n833 185
R17487 vdd.n2348 vdd.n2347 185
R17488 vdd.n2349 vdd.n2348 185
R17489 vdd.n2345 vdd.n845 185
R17490 vdd.n1227 vdd.n845 185
R17491 vdd.n2344 vdd.n2343 185
R17492 vdd.n2343 vdd.n2342 185
R17493 vdd.n848 vdd.n847 185
R17494 vdd.n849 vdd.n848 185
R17495 vdd.n2333 vdd.n2332 185
R17496 vdd.n2334 vdd.n2333 185
R17497 vdd.n2331 vdd.n859 185
R17498 vdd.n859 vdd.n856 185
R17499 vdd.n2330 vdd.n2329 185
R17500 vdd.n2329 vdd.n2328 185
R17501 vdd.n861 vdd.n860 185
R17502 vdd.n1253 vdd.n861 185
R17503 vdd.n2321 vdd.n2320 185
R17504 vdd.n2322 vdd.n2321 185
R17505 vdd.n2319 vdd.n869 185
R17506 vdd.n874 vdd.n869 185
R17507 vdd.n2318 vdd.n2317 185
R17508 vdd.n2317 vdd.n2316 185
R17509 vdd.n871 vdd.n870 185
R17510 vdd.n880 vdd.n871 185
R17511 vdd.n2309 vdd.n2308 185
R17512 vdd.n2310 vdd.n2309 185
R17513 vdd.n2307 vdd.n881 185
R17514 vdd.n1265 vdd.n881 185
R17515 vdd.n2306 vdd.n2305 185
R17516 vdd.n2305 vdd.n2304 185
R17517 vdd.n883 vdd.n882 185
R17518 vdd.n884 vdd.n883 185
R17519 vdd.n2297 vdd.n2296 185
R17520 vdd.n2298 vdd.n2297 185
R17521 vdd.n2295 vdd.n893 185
R17522 vdd.n893 vdd.n890 185
R17523 vdd.n2294 vdd.n2293 185
R17524 vdd.n2293 vdd.n2292 185
R17525 vdd.n895 vdd.n894 185
R17526 vdd.n904 vdd.n895 185
R17527 vdd.n2284 vdd.n2283 185
R17528 vdd.n2285 vdd.n2284 185
R17529 vdd.n2282 vdd.n905 185
R17530 vdd.n911 vdd.n905 185
R17531 vdd.n2281 vdd.n2280 185
R17532 vdd.n2280 vdd.n2279 185
R17533 vdd.n907 vdd.n906 185
R17534 vdd.n908 vdd.n907 185
R17535 vdd.n2272 vdd.n2271 185
R17536 vdd.n2273 vdd.n2272 185
R17537 vdd.n2270 vdd.n918 185
R17538 vdd.n918 vdd.n915 185
R17539 vdd.n2269 vdd.n2268 185
R17540 vdd.n2268 vdd.n2267 185
R17541 vdd.n920 vdd.n919 185
R17542 vdd.n921 vdd.n920 185
R17543 vdd.n2260 vdd.n2259 185
R17544 vdd.n2261 vdd.n2260 185
R17545 vdd.n2258 vdd.n929 185
R17546 vdd.n934 vdd.n929 185
R17547 vdd.n2257 vdd.n2256 185
R17548 vdd.n2256 vdd.n2255 185
R17549 vdd.n931 vdd.n930 185
R17550 vdd.n940 vdd.n931 185
R17551 vdd.n2248 vdd.n2247 185
R17552 vdd.n2249 vdd.n2248 185
R17553 vdd.n2246 vdd.n941 185
R17554 vdd.n947 vdd.n941 185
R17555 vdd.n2245 vdd.n2244 185
R17556 vdd.n2244 vdd.n2243 185
R17557 vdd.n943 vdd.n942 185
R17558 vdd.n944 vdd.n943 185
R17559 vdd.n2236 vdd.n2235 185
R17560 vdd.n2237 vdd.n2236 185
R17561 vdd.n2234 vdd.n954 185
R17562 vdd.n954 vdd.n951 185
R17563 vdd.n2233 vdd.n2232 185
R17564 vdd.n2232 vdd.n2231 185
R17565 vdd.n956 vdd.n955 185
R17566 vdd.n965 vdd.n956 185
R17567 vdd.n2224 vdd.n2223 185
R17568 vdd.n2225 vdd.n2224 185
R17569 vdd.n2222 vdd.n966 185
R17570 vdd.n966 vdd.n962 185
R17571 vdd.n2221 vdd.n2220 185
R17572 vdd.n968 vdd.n967 185
R17573 vdd.n2217 vdd.n2216 185
R17574 vdd.n2218 vdd.n2217 185
R17575 vdd.n2215 vdd.n1004 185
R17576 vdd.n2214 vdd.n2213 185
R17577 vdd.n2212 vdd.n2211 185
R17578 vdd.n2210 vdd.n2209 185
R17579 vdd.n2208 vdd.n2207 185
R17580 vdd.n2206 vdd.n2205 185
R17581 vdd.n2204 vdd.n2203 185
R17582 vdd.n2202 vdd.n2201 185
R17583 vdd.n2200 vdd.n2199 185
R17584 vdd.n2198 vdd.n2197 185
R17585 vdd.n2196 vdd.n2195 185
R17586 vdd.n2194 vdd.n2193 185
R17587 vdd.n2192 vdd.n2191 185
R17588 vdd.n2190 vdd.n2189 185
R17589 vdd.n2188 vdd.n2187 185
R17590 vdd.n1149 vdd.n1005 185
R17591 vdd.n1151 vdd.n1150 185
R17592 vdd.n1153 vdd.n1152 185
R17593 vdd.n1155 vdd.n1154 185
R17594 vdd.n1157 vdd.n1156 185
R17595 vdd.n1159 vdd.n1158 185
R17596 vdd.n1161 vdd.n1160 185
R17597 vdd.n1163 vdd.n1162 185
R17598 vdd.n1165 vdd.n1164 185
R17599 vdd.n1167 vdd.n1166 185
R17600 vdd.n1169 vdd.n1168 185
R17601 vdd.n1171 vdd.n1170 185
R17602 vdd.n1173 vdd.n1172 185
R17603 vdd.n1175 vdd.n1174 185
R17604 vdd.n1178 vdd.n1177 185
R17605 vdd.n1180 vdd.n1179 185
R17606 vdd.n1182 vdd.n1181 185
R17607 vdd.n2427 vdd.n2426 185
R17608 vdd.n2429 vdd.n2428 185
R17609 vdd.n2431 vdd.n2430 185
R17610 vdd.n2434 vdd.n2433 185
R17611 vdd.n2436 vdd.n2435 185
R17612 vdd.n2438 vdd.n2437 185
R17613 vdd.n2440 vdd.n2439 185
R17614 vdd.n2442 vdd.n2441 185
R17615 vdd.n2444 vdd.n2443 185
R17616 vdd.n2446 vdd.n2445 185
R17617 vdd.n2448 vdd.n2447 185
R17618 vdd.n2450 vdd.n2449 185
R17619 vdd.n2452 vdd.n2451 185
R17620 vdd.n2454 vdd.n2453 185
R17621 vdd.n2456 vdd.n2455 185
R17622 vdd.n2458 vdd.n2457 185
R17623 vdd.n2460 vdd.n2459 185
R17624 vdd.n2462 vdd.n2461 185
R17625 vdd.n2464 vdd.n2463 185
R17626 vdd.n2466 vdd.n2465 185
R17627 vdd.n2468 vdd.n2467 185
R17628 vdd.n2470 vdd.n2469 185
R17629 vdd.n2472 vdd.n2471 185
R17630 vdd.n2474 vdd.n2473 185
R17631 vdd.n2476 vdd.n2475 185
R17632 vdd.n2478 vdd.n2477 185
R17633 vdd.n2480 vdd.n2479 185
R17634 vdd.n2482 vdd.n2481 185
R17635 vdd.n2484 vdd.n2483 185
R17636 vdd.n2486 vdd.n2485 185
R17637 vdd.n2488 vdd.n2487 185
R17638 vdd.n2490 vdd.n2489 185
R17639 vdd.n2492 vdd.n2491 185
R17640 vdd.n2493 vdd.n827 185
R17641 vdd.n2495 vdd.n2494 185
R17642 vdd.n2496 vdd.n2495 185
R17643 vdd.n2425 vdd.n831 185
R17644 vdd.n2425 vdd.n2424 185
R17645 vdd.n1225 vdd.n832 185
R17646 vdd.n833 vdd.n832 185
R17647 vdd.n1226 vdd.n843 185
R17648 vdd.n2349 vdd.n843 185
R17649 vdd.n1229 vdd.n1228 185
R17650 vdd.n1228 vdd.n1227 185
R17651 vdd.n1230 vdd.n850 185
R17652 vdd.n2342 vdd.n850 185
R17653 vdd.n1232 vdd.n1231 185
R17654 vdd.n1231 vdd.n849 185
R17655 vdd.n1233 vdd.n857 185
R17656 vdd.n2334 vdd.n857 185
R17657 vdd.n1235 vdd.n1234 185
R17658 vdd.n1234 vdd.n856 185
R17659 vdd.n1236 vdd.n862 185
R17660 vdd.n2328 vdd.n862 185
R17661 vdd.n1255 vdd.n1254 185
R17662 vdd.n1254 vdd.n1253 185
R17663 vdd.n1256 vdd.n867 185
R17664 vdd.n2322 vdd.n867 185
R17665 vdd.n1258 vdd.n1257 185
R17666 vdd.n1257 vdd.n874 185
R17667 vdd.n1259 vdd.n872 185
R17668 vdd.n2316 vdd.n872 185
R17669 vdd.n1261 vdd.n1260 185
R17670 vdd.n1260 vdd.n880 185
R17671 vdd.n1262 vdd.n878 185
R17672 vdd.n2310 vdd.n878 185
R17673 vdd.n1264 vdd.n1263 185
R17674 vdd.n1265 vdd.n1264 185
R17675 vdd.n1224 vdd.n885 185
R17676 vdd.n2304 vdd.n885 185
R17677 vdd.n1223 vdd.n1222 185
R17678 vdd.n1222 vdd.n884 185
R17679 vdd.n1221 vdd.n891 185
R17680 vdd.n2298 vdd.n891 185
R17681 vdd.n1220 vdd.n1219 185
R17682 vdd.n1219 vdd.n890 185
R17683 vdd.n1218 vdd.n896 185
R17684 vdd.n2292 vdd.n896 185
R17685 vdd.n1217 vdd.n1216 185
R17686 vdd.n1216 vdd.n904 185
R17687 vdd.n1215 vdd.n902 185
R17688 vdd.n2285 vdd.n902 185
R17689 vdd.n1214 vdd.n1213 185
R17690 vdd.n1213 vdd.n911 185
R17691 vdd.n1212 vdd.n909 185
R17692 vdd.n2279 vdd.n909 185
R17693 vdd.n1211 vdd.n1210 185
R17694 vdd.n1210 vdd.n908 185
R17695 vdd.n1209 vdd.n916 185
R17696 vdd.n2273 vdd.n916 185
R17697 vdd.n1208 vdd.n1207 185
R17698 vdd.n1207 vdd.n915 185
R17699 vdd.n1206 vdd.n922 185
R17700 vdd.n2267 vdd.n922 185
R17701 vdd.n1205 vdd.n1204 185
R17702 vdd.n1204 vdd.n921 185
R17703 vdd.n1203 vdd.n927 185
R17704 vdd.n2261 vdd.n927 185
R17705 vdd.n1202 vdd.n1201 185
R17706 vdd.n1201 vdd.n934 185
R17707 vdd.n1200 vdd.n932 185
R17708 vdd.n2255 vdd.n932 185
R17709 vdd.n1199 vdd.n1198 185
R17710 vdd.n1198 vdd.n940 185
R17711 vdd.n1197 vdd.n938 185
R17712 vdd.n2249 vdd.n938 185
R17713 vdd.n1196 vdd.n1195 185
R17714 vdd.n1195 vdd.n947 185
R17715 vdd.n1194 vdd.n945 185
R17716 vdd.n2243 vdd.n945 185
R17717 vdd.n1193 vdd.n1192 185
R17718 vdd.n1192 vdd.n944 185
R17719 vdd.n1191 vdd.n952 185
R17720 vdd.n2237 vdd.n952 185
R17721 vdd.n1190 vdd.n1189 185
R17722 vdd.n1189 vdd.n951 185
R17723 vdd.n1188 vdd.n957 185
R17724 vdd.n2231 vdd.n957 185
R17725 vdd.n1187 vdd.n1186 185
R17726 vdd.n1186 vdd.n965 185
R17727 vdd.n1185 vdd.n963 185
R17728 vdd.n2225 vdd.n963 185
R17729 vdd.n1184 vdd.n1183 185
R17730 vdd.n1183 vdd.n962 185
R17731 vdd.n3409 vdd.n3408 185
R17732 vdd.n3410 vdd.n3409 185
R17733 vdd.n347 vdd.n346 185
R17734 vdd.n3411 vdd.n347 185
R17735 vdd.n3414 vdd.n3413 185
R17736 vdd.n3413 vdd.n3412 185
R17737 vdd.n3415 vdd.n341 185
R17738 vdd.n341 vdd.n340 185
R17739 vdd.n3417 vdd.n3416 185
R17740 vdd.n3418 vdd.n3417 185
R17741 vdd.n336 vdd.n335 185
R17742 vdd.n3419 vdd.n336 185
R17743 vdd.n3422 vdd.n3421 185
R17744 vdd.n3421 vdd.n3420 185
R17745 vdd.n3423 vdd.n330 185
R17746 vdd.n330 vdd.n329 185
R17747 vdd.n3425 vdd.n3424 185
R17748 vdd.n3426 vdd.n3425 185
R17749 vdd.n324 vdd.n323 185
R17750 vdd.n3427 vdd.n324 185
R17751 vdd.n3430 vdd.n3429 185
R17752 vdd.n3429 vdd.n3428 185
R17753 vdd.n3431 vdd.n319 185
R17754 vdd.n325 vdd.n319 185
R17755 vdd.n3433 vdd.n3432 185
R17756 vdd.n3434 vdd.n3433 185
R17757 vdd.n315 vdd.n313 185
R17758 vdd.n3435 vdd.n315 185
R17759 vdd.n3438 vdd.n3437 185
R17760 vdd.n3437 vdd.n3436 185
R17761 vdd.n314 vdd.n312 185
R17762 vdd.n481 vdd.n314 185
R17763 vdd.n3260 vdd.n3259 185
R17764 vdd.n3261 vdd.n3260 185
R17765 vdd.n483 vdd.n482 185
R17766 vdd.n3252 vdd.n482 185
R17767 vdd.n3255 vdd.n3254 185
R17768 vdd.n3254 vdd.n3253 185
R17769 vdd.n486 vdd.n485 185
R17770 vdd.n493 vdd.n486 185
R17771 vdd.n3243 vdd.n3242 185
R17772 vdd.n3244 vdd.n3243 185
R17773 vdd.n495 vdd.n494 185
R17774 vdd.n494 vdd.n492 185
R17775 vdd.n3238 vdd.n3237 185
R17776 vdd.n3237 vdd.n3236 185
R17777 vdd.n498 vdd.n497 185
R17778 vdd.n499 vdd.n498 185
R17779 vdd.n3227 vdd.n3226 185
R17780 vdd.n3228 vdd.n3227 185
R17781 vdd.n507 vdd.n506 185
R17782 vdd.n506 vdd.n505 185
R17783 vdd.n3222 vdd.n3221 185
R17784 vdd.n3221 vdd.n3220 185
R17785 vdd.n510 vdd.n509 185
R17786 vdd.n511 vdd.n510 185
R17787 vdd.n3211 vdd.n3210 185
R17788 vdd.n3212 vdd.n3211 185
R17789 vdd.n3207 vdd.n517 185
R17790 vdd.n3206 vdd.n3205 185
R17791 vdd.n3203 vdd.n519 185
R17792 vdd.n3203 vdd.n516 185
R17793 vdd.n3202 vdd.n3201 185
R17794 vdd.n3200 vdd.n3199 185
R17795 vdd.n3198 vdd.n3197 185
R17796 vdd.n3196 vdd.n3195 185
R17797 vdd.n3194 vdd.n525 185
R17798 vdd.n3192 vdd.n3191 185
R17799 vdd.n3190 vdd.n526 185
R17800 vdd.n3189 vdd.n3188 185
R17801 vdd.n3186 vdd.n531 185
R17802 vdd.n3184 vdd.n3183 185
R17803 vdd.n3182 vdd.n532 185
R17804 vdd.n3181 vdd.n3180 185
R17805 vdd.n3178 vdd.n537 185
R17806 vdd.n3176 vdd.n3175 185
R17807 vdd.n3174 vdd.n538 185
R17808 vdd.n3173 vdd.n3172 185
R17809 vdd.n3170 vdd.n545 185
R17810 vdd.n3168 vdd.n3167 185
R17811 vdd.n3166 vdd.n546 185
R17812 vdd.n3165 vdd.n3164 185
R17813 vdd.n3162 vdd.n551 185
R17814 vdd.n3160 vdd.n3159 185
R17815 vdd.n3158 vdd.n552 185
R17816 vdd.n3157 vdd.n3156 185
R17817 vdd.n3154 vdd.n557 185
R17818 vdd.n3152 vdd.n3151 185
R17819 vdd.n3150 vdd.n558 185
R17820 vdd.n3149 vdd.n3148 185
R17821 vdd.n3146 vdd.n563 185
R17822 vdd.n3144 vdd.n3143 185
R17823 vdd.n3142 vdd.n564 185
R17824 vdd.n3141 vdd.n3140 185
R17825 vdd.n3138 vdd.n569 185
R17826 vdd.n3136 vdd.n3135 185
R17827 vdd.n3134 vdd.n570 185
R17828 vdd.n3133 vdd.n3132 185
R17829 vdd.n3130 vdd.n575 185
R17830 vdd.n3128 vdd.n3127 185
R17831 vdd.n3126 vdd.n576 185
R17832 vdd.n585 vdd.n579 185
R17833 vdd.n3122 vdd.n3121 185
R17834 vdd.n3119 vdd.n583 185
R17835 vdd.n3118 vdd.n3117 185
R17836 vdd.n3116 vdd.n3115 185
R17837 vdd.n3114 vdd.n589 185
R17838 vdd.n3112 vdd.n3111 185
R17839 vdd.n3110 vdd.n590 185
R17840 vdd.n3109 vdd.n3108 185
R17841 vdd.n3106 vdd.n595 185
R17842 vdd.n3104 vdd.n3103 185
R17843 vdd.n3102 vdd.n596 185
R17844 vdd.n3101 vdd.n3100 185
R17845 vdd.n3098 vdd.n601 185
R17846 vdd.n3096 vdd.n3095 185
R17847 vdd.n3094 vdd.n602 185
R17848 vdd.n3093 vdd.n3092 185
R17849 vdd.n3090 vdd.n3089 185
R17850 vdd.n3088 vdd.n3087 185
R17851 vdd.n3086 vdd.n3085 185
R17852 vdd.n3084 vdd.n3083 185
R17853 vdd.n3079 vdd.n515 185
R17854 vdd.n516 vdd.n515 185
R17855 vdd.n3292 vdd.n3291 185
R17856 vdd.n3296 vdd.n462 185
R17857 vdd.n3298 vdd.n3297 185
R17858 vdd.n3300 vdd.n460 185
R17859 vdd.n3302 vdd.n3301 185
R17860 vdd.n3303 vdd.n455 185
R17861 vdd.n3305 vdd.n3304 185
R17862 vdd.n3307 vdd.n453 185
R17863 vdd.n3309 vdd.n3308 185
R17864 vdd.n3310 vdd.n448 185
R17865 vdd.n3312 vdd.n3311 185
R17866 vdd.n3314 vdd.n446 185
R17867 vdd.n3316 vdd.n3315 185
R17868 vdd.n3317 vdd.n441 185
R17869 vdd.n3319 vdd.n3318 185
R17870 vdd.n3321 vdd.n439 185
R17871 vdd.n3323 vdd.n3322 185
R17872 vdd.n3324 vdd.n435 185
R17873 vdd.n3326 vdd.n3325 185
R17874 vdd.n3328 vdd.n432 185
R17875 vdd.n3330 vdd.n3329 185
R17876 vdd.n433 vdd.n426 185
R17877 vdd.n3334 vdd.n430 185
R17878 vdd.n3335 vdd.n422 185
R17879 vdd.n3337 vdd.n3336 185
R17880 vdd.n3339 vdd.n420 185
R17881 vdd.n3341 vdd.n3340 185
R17882 vdd.n3342 vdd.n415 185
R17883 vdd.n3344 vdd.n3343 185
R17884 vdd.n3346 vdd.n413 185
R17885 vdd.n3348 vdd.n3347 185
R17886 vdd.n3349 vdd.n408 185
R17887 vdd.n3351 vdd.n3350 185
R17888 vdd.n3353 vdd.n406 185
R17889 vdd.n3355 vdd.n3354 185
R17890 vdd.n3356 vdd.n401 185
R17891 vdd.n3358 vdd.n3357 185
R17892 vdd.n3360 vdd.n399 185
R17893 vdd.n3362 vdd.n3361 185
R17894 vdd.n3363 vdd.n395 185
R17895 vdd.n3365 vdd.n3364 185
R17896 vdd.n3367 vdd.n392 185
R17897 vdd.n3369 vdd.n3368 185
R17898 vdd.n393 vdd.n386 185
R17899 vdd.n3373 vdd.n390 185
R17900 vdd.n3374 vdd.n382 185
R17901 vdd.n3376 vdd.n3375 185
R17902 vdd.n3378 vdd.n380 185
R17903 vdd.n3380 vdd.n3379 185
R17904 vdd.n3381 vdd.n375 185
R17905 vdd.n3383 vdd.n3382 185
R17906 vdd.n3385 vdd.n373 185
R17907 vdd.n3387 vdd.n3386 185
R17908 vdd.n3388 vdd.n368 185
R17909 vdd.n3390 vdd.n3389 185
R17910 vdd.n3392 vdd.n366 185
R17911 vdd.n3394 vdd.n3393 185
R17912 vdd.n3395 vdd.n360 185
R17913 vdd.n3397 vdd.n3396 185
R17914 vdd.n3399 vdd.n359 185
R17915 vdd.n3400 vdd.n358 185
R17916 vdd.n3403 vdd.n3402 185
R17917 vdd.n3404 vdd.n356 185
R17918 vdd.n3405 vdd.n352 185
R17919 vdd.n3287 vdd.n350 185
R17920 vdd.n3410 vdd.n350 185
R17921 vdd.n3286 vdd.n349 185
R17922 vdd.n3411 vdd.n349 185
R17923 vdd.n3285 vdd.n348 185
R17924 vdd.n3412 vdd.n348 185
R17925 vdd.n468 vdd.n467 185
R17926 vdd.n467 vdd.n340 185
R17927 vdd.n3281 vdd.n339 185
R17928 vdd.n3418 vdd.n339 185
R17929 vdd.n3280 vdd.n338 185
R17930 vdd.n3419 vdd.n338 185
R17931 vdd.n3279 vdd.n337 185
R17932 vdd.n3420 vdd.n337 185
R17933 vdd.n471 vdd.n470 185
R17934 vdd.n470 vdd.n329 185
R17935 vdd.n3275 vdd.n328 185
R17936 vdd.n3426 vdd.n328 185
R17937 vdd.n3274 vdd.n327 185
R17938 vdd.n3427 vdd.n327 185
R17939 vdd.n3273 vdd.n326 185
R17940 vdd.n3428 vdd.n326 185
R17941 vdd.n474 vdd.n473 185
R17942 vdd.n473 vdd.n325 185
R17943 vdd.n3269 vdd.n318 185
R17944 vdd.n3434 vdd.n318 185
R17945 vdd.n3268 vdd.n317 185
R17946 vdd.n3435 vdd.n317 185
R17947 vdd.n3267 vdd.n316 185
R17948 vdd.n3436 vdd.n316 185
R17949 vdd.n480 vdd.n476 185
R17950 vdd.n481 vdd.n480 185
R17951 vdd.n3263 vdd.n3262 185
R17952 vdd.n3262 vdd.n3261 185
R17953 vdd.n479 vdd.n478 185
R17954 vdd.n3252 vdd.n479 185
R17955 vdd.n3251 vdd.n3250 185
R17956 vdd.n3253 vdd.n3251 185
R17957 vdd.n488 vdd.n487 185
R17958 vdd.n493 vdd.n487 185
R17959 vdd.n3246 vdd.n3245 185
R17960 vdd.n3245 vdd.n3244 185
R17961 vdd.n491 vdd.n490 185
R17962 vdd.n492 vdd.n491 185
R17963 vdd.n3235 vdd.n3234 185
R17964 vdd.n3236 vdd.n3235 185
R17965 vdd.n501 vdd.n500 185
R17966 vdd.n500 vdd.n499 185
R17967 vdd.n3230 vdd.n3229 185
R17968 vdd.n3229 vdd.n3228 185
R17969 vdd.n504 vdd.n503 185
R17970 vdd.n505 vdd.n504 185
R17971 vdd.n3219 vdd.n3218 185
R17972 vdd.n3220 vdd.n3219 185
R17973 vdd.n513 vdd.n512 185
R17974 vdd.n512 vdd.n511 185
R17975 vdd.n3214 vdd.n3213 185
R17976 vdd.n3213 vdd.n3212 185
R17977 vdd.n2803 vdd.n2802 185
R17978 vdd.n790 vdd.n789 185
R17979 vdd.n2799 vdd.n2798 185
R17980 vdd.n2800 vdd.n2799 185
R17981 vdd.n2797 vdd.n2531 185
R17982 vdd.n2796 vdd.n2795 185
R17983 vdd.n2794 vdd.n2793 185
R17984 vdd.n2792 vdd.n2791 185
R17985 vdd.n2790 vdd.n2789 185
R17986 vdd.n2788 vdd.n2787 185
R17987 vdd.n2786 vdd.n2785 185
R17988 vdd.n2784 vdd.n2783 185
R17989 vdd.n2782 vdd.n2781 185
R17990 vdd.n2780 vdd.n2779 185
R17991 vdd.n2778 vdd.n2777 185
R17992 vdd.n2776 vdd.n2775 185
R17993 vdd.n2774 vdd.n2773 185
R17994 vdd.n2772 vdd.n2771 185
R17995 vdd.n2770 vdd.n2769 185
R17996 vdd.n2768 vdd.n2767 185
R17997 vdd.n2766 vdd.n2765 185
R17998 vdd.n2764 vdd.n2763 185
R17999 vdd.n2762 vdd.n2761 185
R18000 vdd.n2760 vdd.n2759 185
R18001 vdd.n2758 vdd.n2757 185
R18002 vdd.n2756 vdd.n2755 185
R18003 vdd.n2754 vdd.n2753 185
R18004 vdd.n2752 vdd.n2751 185
R18005 vdd.n2750 vdd.n2749 185
R18006 vdd.n2748 vdd.n2747 185
R18007 vdd.n2746 vdd.n2745 185
R18008 vdd.n2744 vdd.n2743 185
R18009 vdd.n2742 vdd.n2741 185
R18010 vdd.n2739 vdd.n2738 185
R18011 vdd.n2737 vdd.n2736 185
R18012 vdd.n2735 vdd.n2734 185
R18013 vdd.n2980 vdd.n2979 185
R18014 vdd.n2981 vdd.n660 185
R18015 vdd.n2983 vdd.n2982 185
R18016 vdd.n2985 vdd.n658 185
R18017 vdd.n2987 vdd.n2986 185
R18018 vdd.n2988 vdd.n657 185
R18019 vdd.n2990 vdd.n2989 185
R18020 vdd.n2992 vdd.n655 185
R18021 vdd.n2994 vdd.n2993 185
R18022 vdd.n2995 vdd.n654 185
R18023 vdd.n2997 vdd.n2996 185
R18024 vdd.n2999 vdd.n652 185
R18025 vdd.n3001 vdd.n3000 185
R18026 vdd.n3002 vdd.n651 185
R18027 vdd.n3004 vdd.n3003 185
R18028 vdd.n3006 vdd.n649 185
R18029 vdd.n3008 vdd.n3007 185
R18030 vdd.n3010 vdd.n648 185
R18031 vdd.n3012 vdd.n3011 185
R18032 vdd.n3014 vdd.n646 185
R18033 vdd.n3016 vdd.n3015 185
R18034 vdd.n3017 vdd.n645 185
R18035 vdd.n3019 vdd.n3018 185
R18036 vdd.n3021 vdd.n643 185
R18037 vdd.n3023 vdd.n3022 185
R18038 vdd.n3024 vdd.n642 185
R18039 vdd.n3026 vdd.n3025 185
R18040 vdd.n3028 vdd.n640 185
R18041 vdd.n3030 vdd.n3029 185
R18042 vdd.n3031 vdd.n639 185
R18043 vdd.n3033 vdd.n3032 185
R18044 vdd.n3035 vdd.n638 185
R18045 vdd.n3036 vdd.n637 185
R18046 vdd.n3039 vdd.n3038 185
R18047 vdd.n3040 vdd.n635 185
R18048 vdd.n635 vdd.n613 185
R18049 vdd.n2977 vdd.n632 185
R18050 vdd.n3043 vdd.n632 185
R18051 vdd.n2976 vdd.n2975 185
R18052 vdd.n2975 vdd.n631 185
R18053 vdd.n2974 vdd.n664 185
R18054 vdd.n2974 vdd.n2973 185
R18055 vdd.n2617 vdd.n665 185
R18056 vdd.n674 vdd.n665 185
R18057 vdd.n2618 vdd.n672 185
R18058 vdd.n2967 vdd.n672 185
R18059 vdd.n2620 vdd.n2619 185
R18060 vdd.n2619 vdd.n671 185
R18061 vdd.n2621 vdd.n680 185
R18062 vdd.n2916 vdd.n680 185
R18063 vdd.n2623 vdd.n2622 185
R18064 vdd.n2622 vdd.n679 185
R18065 vdd.n2624 vdd.n685 185
R18066 vdd.n2910 vdd.n685 185
R18067 vdd.n2626 vdd.n2625 185
R18068 vdd.n2625 vdd.n692 185
R18069 vdd.n2627 vdd.n690 185
R18070 vdd.n2904 vdd.n690 185
R18071 vdd.n2629 vdd.n2628 185
R18072 vdd.n2628 vdd.n698 185
R18073 vdd.n2630 vdd.n696 185
R18074 vdd.n2898 vdd.n696 185
R18075 vdd.n2632 vdd.n2631 185
R18076 vdd.n2631 vdd.n705 185
R18077 vdd.n2633 vdd.n703 185
R18078 vdd.n2892 vdd.n703 185
R18079 vdd.n2635 vdd.n2634 185
R18080 vdd.n2634 vdd.n702 185
R18081 vdd.n2636 vdd.n710 185
R18082 vdd.n2886 vdd.n710 185
R18083 vdd.n2638 vdd.n2637 185
R18084 vdd.n2637 vdd.n709 185
R18085 vdd.n2639 vdd.n716 185
R18086 vdd.n2880 vdd.n716 185
R18087 vdd.n2641 vdd.n2640 185
R18088 vdd.n2640 vdd.n715 185
R18089 vdd.n2642 vdd.n721 185
R18090 vdd.n2874 vdd.n721 185
R18091 vdd.n2644 vdd.n2643 185
R18092 vdd.n2643 vdd.n729 185
R18093 vdd.n2645 vdd.n727 185
R18094 vdd.n2868 vdd.n727 185
R18095 vdd.n2647 vdd.n2646 185
R18096 vdd.n2646 vdd.n736 185
R18097 vdd.n2648 vdd.n734 185
R18098 vdd.n2862 vdd.n734 185
R18099 vdd.n2650 vdd.n2649 185
R18100 vdd.n2649 vdd.n733 185
R18101 vdd.n2651 vdd.n741 185
R18102 vdd.n2855 vdd.n741 185
R18103 vdd.n2653 vdd.n2652 185
R18104 vdd.n2652 vdd.n740 185
R18105 vdd.n2654 vdd.n746 185
R18106 vdd.n2849 vdd.n746 185
R18107 vdd.n2656 vdd.n2655 185
R18108 vdd.n2655 vdd.n753 185
R18109 vdd.n2657 vdd.n751 185
R18110 vdd.n2843 vdd.n751 185
R18111 vdd.n2659 vdd.n2658 185
R18112 vdd.n2658 vdd.n759 185
R18113 vdd.n2660 vdd.n757 185
R18114 vdd.n2837 vdd.n757 185
R18115 vdd.n2712 vdd.n2711 185
R18116 vdd.n2711 vdd.n2710 185
R18117 vdd.n2713 vdd.n763 185
R18118 vdd.n2831 vdd.n763 185
R18119 vdd.n2715 vdd.n2714 185
R18120 vdd.n2716 vdd.n2715 185
R18121 vdd.n2616 vdd.n769 185
R18122 vdd.n2825 vdd.n769 185
R18123 vdd.n2615 vdd.n2614 185
R18124 vdd.n2614 vdd.n768 185
R18125 vdd.n2613 vdd.n775 185
R18126 vdd.n2819 vdd.n775 185
R18127 vdd.n2612 vdd.n2611 185
R18128 vdd.n2611 vdd.n774 185
R18129 vdd.n2534 vdd.n780 185
R18130 vdd.n2813 vdd.n780 185
R18131 vdd.n2730 vdd.n2729 185
R18132 vdd.n2729 vdd.n2728 185
R18133 vdd.n2731 vdd.n786 185
R18134 vdd.n2807 vdd.n786 185
R18135 vdd.n2733 vdd.n2732 185
R18136 vdd.n2733 vdd.n785 185
R18137 vdd.n2804 vdd.n788 185
R18138 vdd.n788 vdd.n785 185
R18139 vdd.n2806 vdd.n2805 185
R18140 vdd.n2807 vdd.n2806 185
R18141 vdd.n779 vdd.n778 185
R18142 vdd.n2728 vdd.n779 185
R18143 vdd.n2815 vdd.n2814 185
R18144 vdd.n2814 vdd.n2813 185
R18145 vdd.n2816 vdd.n777 185
R18146 vdd.n777 vdd.n774 185
R18147 vdd.n2818 vdd.n2817 185
R18148 vdd.n2819 vdd.n2818 185
R18149 vdd.n767 vdd.n766 185
R18150 vdd.n768 vdd.n767 185
R18151 vdd.n2827 vdd.n2826 185
R18152 vdd.n2826 vdd.n2825 185
R18153 vdd.n2828 vdd.n765 185
R18154 vdd.n2716 vdd.n765 185
R18155 vdd.n2830 vdd.n2829 185
R18156 vdd.n2831 vdd.n2830 185
R18157 vdd.n756 vdd.n755 185
R18158 vdd.n2710 vdd.n756 185
R18159 vdd.n2839 vdd.n2838 185
R18160 vdd.n2838 vdd.n2837 185
R18161 vdd.n2840 vdd.n754 185
R18162 vdd.n759 vdd.n754 185
R18163 vdd.n2842 vdd.n2841 185
R18164 vdd.n2843 vdd.n2842 185
R18165 vdd.n745 vdd.n744 185
R18166 vdd.n753 vdd.n745 185
R18167 vdd.n2851 vdd.n2850 185
R18168 vdd.n2850 vdd.n2849 185
R18169 vdd.n2852 vdd.n743 185
R18170 vdd.n743 vdd.n740 185
R18171 vdd.n2854 vdd.n2853 185
R18172 vdd.n2855 vdd.n2854 185
R18173 vdd.n732 vdd.n731 185
R18174 vdd.n733 vdd.n732 185
R18175 vdd.n2864 vdd.n2863 185
R18176 vdd.n2863 vdd.n2862 185
R18177 vdd.n2865 vdd.n730 185
R18178 vdd.n736 vdd.n730 185
R18179 vdd.n2867 vdd.n2866 185
R18180 vdd.n2868 vdd.n2867 185
R18181 vdd.n720 vdd.n719 185
R18182 vdd.n729 vdd.n720 185
R18183 vdd.n2876 vdd.n2875 185
R18184 vdd.n2875 vdd.n2874 185
R18185 vdd.n2877 vdd.n718 185
R18186 vdd.n718 vdd.n715 185
R18187 vdd.n2879 vdd.n2878 185
R18188 vdd.n2880 vdd.n2879 185
R18189 vdd.n708 vdd.n707 185
R18190 vdd.n709 vdd.n708 185
R18191 vdd.n2888 vdd.n2887 185
R18192 vdd.n2887 vdd.n2886 185
R18193 vdd.n2889 vdd.n706 185
R18194 vdd.n706 vdd.n702 185
R18195 vdd.n2891 vdd.n2890 185
R18196 vdd.n2892 vdd.n2891 185
R18197 vdd.n695 vdd.n694 185
R18198 vdd.n705 vdd.n695 185
R18199 vdd.n2900 vdd.n2899 185
R18200 vdd.n2899 vdd.n2898 185
R18201 vdd.n2901 vdd.n693 185
R18202 vdd.n698 vdd.n693 185
R18203 vdd.n2903 vdd.n2902 185
R18204 vdd.n2904 vdd.n2903 185
R18205 vdd.n684 vdd.n683 185
R18206 vdd.n692 vdd.n684 185
R18207 vdd.n2912 vdd.n2911 185
R18208 vdd.n2911 vdd.n2910 185
R18209 vdd.n2913 vdd.n682 185
R18210 vdd.n682 vdd.n679 185
R18211 vdd.n2915 vdd.n2914 185
R18212 vdd.n2916 vdd.n2915 185
R18213 vdd.n670 vdd.n669 185
R18214 vdd.n671 vdd.n670 185
R18215 vdd.n2969 vdd.n2968 185
R18216 vdd.n2968 vdd.n2967 185
R18217 vdd.n2970 vdd.n668 185
R18218 vdd.n674 vdd.n668 185
R18219 vdd.n2972 vdd.n2971 185
R18220 vdd.n2973 vdd.n2972 185
R18221 vdd.n636 vdd.n634 185
R18222 vdd.n634 vdd.n631 185
R18223 vdd.n3042 vdd.n3041 185
R18224 vdd.n3043 vdd.n3042 185
R18225 vdd.n2423 vdd.n2422 185
R18226 vdd.n2424 vdd.n2423 185
R18227 vdd.n837 vdd.n835 185
R18228 vdd.n835 vdd.n833 185
R18229 vdd.n2338 vdd.n844 185
R18230 vdd.n2349 vdd.n844 185
R18231 vdd.n2339 vdd.n853 185
R18232 vdd.n1227 vdd.n853 185
R18233 vdd.n2341 vdd.n2340 185
R18234 vdd.n2342 vdd.n2341 185
R18235 vdd.n2337 vdd.n852 185
R18236 vdd.n852 vdd.n849 185
R18237 vdd.n2336 vdd.n2335 185
R18238 vdd.n2335 vdd.n2334 185
R18239 vdd.n855 vdd.n854 185
R18240 vdd.n856 vdd.n855 185
R18241 vdd.n2327 vdd.n2326 185
R18242 vdd.n2328 vdd.n2327 185
R18243 vdd.n2325 vdd.n864 185
R18244 vdd.n1253 vdd.n864 185
R18245 vdd.n2324 vdd.n2323 185
R18246 vdd.n2323 vdd.n2322 185
R18247 vdd.n866 vdd.n865 185
R18248 vdd.n874 vdd.n866 185
R18249 vdd.n2315 vdd.n2314 185
R18250 vdd.n2316 vdd.n2315 185
R18251 vdd.n2313 vdd.n875 185
R18252 vdd.n880 vdd.n875 185
R18253 vdd.n2312 vdd.n2311 185
R18254 vdd.n2311 vdd.n2310 185
R18255 vdd.n877 vdd.n876 185
R18256 vdd.n1265 vdd.n877 185
R18257 vdd.n2303 vdd.n2302 185
R18258 vdd.n2304 vdd.n2303 185
R18259 vdd.n2301 vdd.n887 185
R18260 vdd.n887 vdd.n884 185
R18261 vdd.n2300 vdd.n2299 185
R18262 vdd.n2299 vdd.n2298 185
R18263 vdd.n889 vdd.n888 185
R18264 vdd.n890 vdd.n889 185
R18265 vdd.n2291 vdd.n2290 185
R18266 vdd.n2292 vdd.n2291 185
R18267 vdd.n2288 vdd.n898 185
R18268 vdd.n904 vdd.n898 185
R18269 vdd.n2287 vdd.n2286 185
R18270 vdd.n2286 vdd.n2285 185
R18271 vdd.n901 vdd.n900 185
R18272 vdd.n911 vdd.n901 185
R18273 vdd.n2278 vdd.n2277 185
R18274 vdd.n2279 vdd.n2278 185
R18275 vdd.n2276 vdd.n912 185
R18276 vdd.n912 vdd.n908 185
R18277 vdd.n2275 vdd.n2274 185
R18278 vdd.n2274 vdd.n2273 185
R18279 vdd.n914 vdd.n913 185
R18280 vdd.n915 vdd.n914 185
R18281 vdd.n2266 vdd.n2265 185
R18282 vdd.n2267 vdd.n2266 185
R18283 vdd.n2264 vdd.n924 185
R18284 vdd.n924 vdd.n921 185
R18285 vdd.n2263 vdd.n2262 185
R18286 vdd.n2262 vdd.n2261 185
R18287 vdd.n926 vdd.n925 185
R18288 vdd.n934 vdd.n926 185
R18289 vdd.n2254 vdd.n2253 185
R18290 vdd.n2255 vdd.n2254 185
R18291 vdd.n2252 vdd.n935 185
R18292 vdd.n940 vdd.n935 185
R18293 vdd.n2251 vdd.n2250 185
R18294 vdd.n2250 vdd.n2249 185
R18295 vdd.n937 vdd.n936 185
R18296 vdd.n947 vdd.n937 185
R18297 vdd.n2242 vdd.n2241 185
R18298 vdd.n2243 vdd.n2242 185
R18299 vdd.n2240 vdd.n948 185
R18300 vdd.n948 vdd.n944 185
R18301 vdd.n2239 vdd.n2238 185
R18302 vdd.n2238 vdd.n2237 185
R18303 vdd.n950 vdd.n949 185
R18304 vdd.n951 vdd.n950 185
R18305 vdd.n2230 vdd.n2229 185
R18306 vdd.n2231 vdd.n2230 185
R18307 vdd.n2228 vdd.n959 185
R18308 vdd.n965 vdd.n959 185
R18309 vdd.n2227 vdd.n2226 185
R18310 vdd.n2226 vdd.n2225 185
R18311 vdd.n961 vdd.n960 185
R18312 vdd.n962 vdd.n961 185
R18313 vdd.n2354 vdd.n808 185
R18314 vdd.n2496 vdd.n808 185
R18315 vdd.n2356 vdd.n2355 185
R18316 vdd.n2358 vdd.n2357 185
R18317 vdd.n2360 vdd.n2359 185
R18318 vdd.n2362 vdd.n2361 185
R18319 vdd.n2364 vdd.n2363 185
R18320 vdd.n2366 vdd.n2365 185
R18321 vdd.n2368 vdd.n2367 185
R18322 vdd.n2370 vdd.n2369 185
R18323 vdd.n2372 vdd.n2371 185
R18324 vdd.n2374 vdd.n2373 185
R18325 vdd.n2376 vdd.n2375 185
R18326 vdd.n2378 vdd.n2377 185
R18327 vdd.n2380 vdd.n2379 185
R18328 vdd.n2382 vdd.n2381 185
R18329 vdd.n2384 vdd.n2383 185
R18330 vdd.n2386 vdd.n2385 185
R18331 vdd.n2388 vdd.n2387 185
R18332 vdd.n2390 vdd.n2389 185
R18333 vdd.n2392 vdd.n2391 185
R18334 vdd.n2394 vdd.n2393 185
R18335 vdd.n2396 vdd.n2395 185
R18336 vdd.n2398 vdd.n2397 185
R18337 vdd.n2400 vdd.n2399 185
R18338 vdd.n2402 vdd.n2401 185
R18339 vdd.n2404 vdd.n2403 185
R18340 vdd.n2406 vdd.n2405 185
R18341 vdd.n2408 vdd.n2407 185
R18342 vdd.n2410 vdd.n2409 185
R18343 vdd.n2412 vdd.n2411 185
R18344 vdd.n2414 vdd.n2413 185
R18345 vdd.n2416 vdd.n2415 185
R18346 vdd.n2418 vdd.n2417 185
R18347 vdd.n2420 vdd.n2419 185
R18348 vdd.n2421 vdd.n836 185
R18349 vdd.n2353 vdd.n834 185
R18350 vdd.n2424 vdd.n834 185
R18351 vdd.n2352 vdd.n2351 185
R18352 vdd.n2351 vdd.n833 185
R18353 vdd.n2350 vdd.n841 185
R18354 vdd.n2350 vdd.n2349 185
R18355 vdd.n1243 vdd.n842 185
R18356 vdd.n1227 vdd.n842 185
R18357 vdd.n1244 vdd.n851 185
R18358 vdd.n2342 vdd.n851 185
R18359 vdd.n1246 vdd.n1245 185
R18360 vdd.n1245 vdd.n849 185
R18361 vdd.n1247 vdd.n858 185
R18362 vdd.n2334 vdd.n858 185
R18363 vdd.n1249 vdd.n1248 185
R18364 vdd.n1248 vdd.n856 185
R18365 vdd.n1250 vdd.n863 185
R18366 vdd.n2328 vdd.n863 185
R18367 vdd.n1252 vdd.n1251 185
R18368 vdd.n1253 vdd.n1252 185
R18369 vdd.n1242 vdd.n868 185
R18370 vdd.n2322 vdd.n868 185
R18371 vdd.n1241 vdd.n1240 185
R18372 vdd.n1240 vdd.n874 185
R18373 vdd.n1239 vdd.n873 185
R18374 vdd.n2316 vdd.n873 185
R18375 vdd.n1238 vdd.n1237 185
R18376 vdd.n1237 vdd.n880 185
R18377 vdd.n1146 vdd.n879 185
R18378 vdd.n2310 vdd.n879 185
R18379 vdd.n1267 vdd.n1266 185
R18380 vdd.n1266 vdd.n1265 185
R18381 vdd.n1268 vdd.n886 185
R18382 vdd.n2304 vdd.n886 185
R18383 vdd.n1270 vdd.n1269 185
R18384 vdd.n1269 vdd.n884 185
R18385 vdd.n1271 vdd.n892 185
R18386 vdd.n2298 vdd.n892 185
R18387 vdd.n1273 vdd.n1272 185
R18388 vdd.n1272 vdd.n890 185
R18389 vdd.n1274 vdd.n897 185
R18390 vdd.n2292 vdd.n897 185
R18391 vdd.n1276 vdd.n1275 185
R18392 vdd.n1275 vdd.n904 185
R18393 vdd.n1277 vdd.n903 185
R18394 vdd.n2285 vdd.n903 185
R18395 vdd.n1279 vdd.n1278 185
R18396 vdd.n1278 vdd.n911 185
R18397 vdd.n1280 vdd.n910 185
R18398 vdd.n2279 vdd.n910 185
R18399 vdd.n1282 vdd.n1281 185
R18400 vdd.n1281 vdd.n908 185
R18401 vdd.n1283 vdd.n917 185
R18402 vdd.n2273 vdd.n917 185
R18403 vdd.n1285 vdd.n1284 185
R18404 vdd.n1284 vdd.n915 185
R18405 vdd.n1286 vdd.n923 185
R18406 vdd.n2267 vdd.n923 185
R18407 vdd.n1288 vdd.n1287 185
R18408 vdd.n1287 vdd.n921 185
R18409 vdd.n1289 vdd.n928 185
R18410 vdd.n2261 vdd.n928 185
R18411 vdd.n1291 vdd.n1290 185
R18412 vdd.n1290 vdd.n934 185
R18413 vdd.n1292 vdd.n933 185
R18414 vdd.n2255 vdd.n933 185
R18415 vdd.n1294 vdd.n1293 185
R18416 vdd.n1293 vdd.n940 185
R18417 vdd.n1295 vdd.n939 185
R18418 vdd.n2249 vdd.n939 185
R18419 vdd.n1297 vdd.n1296 185
R18420 vdd.n1296 vdd.n947 185
R18421 vdd.n1298 vdd.n946 185
R18422 vdd.n2243 vdd.n946 185
R18423 vdd.n1300 vdd.n1299 185
R18424 vdd.n1299 vdd.n944 185
R18425 vdd.n1301 vdd.n953 185
R18426 vdd.n2237 vdd.n953 185
R18427 vdd.n1303 vdd.n1302 185
R18428 vdd.n1302 vdd.n951 185
R18429 vdd.n1304 vdd.n958 185
R18430 vdd.n2231 vdd.n958 185
R18431 vdd.n1306 vdd.n1305 185
R18432 vdd.n1305 vdd.n965 185
R18433 vdd.n1307 vdd.n964 185
R18434 vdd.n2225 vdd.n964 185
R18435 vdd.n1309 vdd.n1308 185
R18436 vdd.n1308 vdd.n962 185
R18437 vdd.n1109 vdd.n1108 185
R18438 vdd.n1111 vdd.n1110 185
R18439 vdd.n1113 vdd.n1112 185
R18440 vdd.n1115 vdd.n1114 185
R18441 vdd.n1117 vdd.n1116 185
R18442 vdd.n1119 vdd.n1118 185
R18443 vdd.n1121 vdd.n1120 185
R18444 vdd.n1123 vdd.n1122 185
R18445 vdd.n1125 vdd.n1124 185
R18446 vdd.n1127 vdd.n1126 185
R18447 vdd.n1129 vdd.n1128 185
R18448 vdd.n1131 vdd.n1130 185
R18449 vdd.n1133 vdd.n1132 185
R18450 vdd.n1135 vdd.n1134 185
R18451 vdd.n1137 vdd.n1136 185
R18452 vdd.n1139 vdd.n1138 185
R18453 vdd.n1141 vdd.n1140 185
R18454 vdd.n1343 vdd.n1142 185
R18455 vdd.n1342 vdd.n1341 185
R18456 vdd.n1340 vdd.n1339 185
R18457 vdd.n1338 vdd.n1337 185
R18458 vdd.n1336 vdd.n1335 185
R18459 vdd.n1334 vdd.n1333 185
R18460 vdd.n1332 vdd.n1331 185
R18461 vdd.n1330 vdd.n1329 185
R18462 vdd.n1328 vdd.n1327 185
R18463 vdd.n1326 vdd.n1325 185
R18464 vdd.n1324 vdd.n1323 185
R18465 vdd.n1322 vdd.n1321 185
R18466 vdd.n1320 vdd.n1319 185
R18467 vdd.n1318 vdd.n1317 185
R18468 vdd.n1316 vdd.n1315 185
R18469 vdd.n1314 vdd.n1313 185
R18470 vdd.n1312 vdd.n1311 185
R18471 vdd.n1310 vdd.n1003 185
R18472 vdd.n2218 vdd.n1003 185
R18473 vdd.n303 vdd.n302 171.744
R18474 vdd.n302 vdd.n301 171.744
R18475 vdd.n301 vdd.n270 171.744
R18476 vdd.n294 vdd.n270 171.744
R18477 vdd.n294 vdd.n293 171.744
R18478 vdd.n293 vdd.n275 171.744
R18479 vdd.n286 vdd.n275 171.744
R18480 vdd.n286 vdd.n285 171.744
R18481 vdd.n285 vdd.n279 171.744
R18482 vdd.n252 vdd.n251 171.744
R18483 vdd.n251 vdd.n250 171.744
R18484 vdd.n250 vdd.n219 171.744
R18485 vdd.n243 vdd.n219 171.744
R18486 vdd.n243 vdd.n242 171.744
R18487 vdd.n242 vdd.n224 171.744
R18488 vdd.n235 vdd.n224 171.744
R18489 vdd.n235 vdd.n234 171.744
R18490 vdd.n234 vdd.n228 171.744
R18491 vdd.n209 vdd.n208 171.744
R18492 vdd.n208 vdd.n207 171.744
R18493 vdd.n207 vdd.n176 171.744
R18494 vdd.n200 vdd.n176 171.744
R18495 vdd.n200 vdd.n199 171.744
R18496 vdd.n199 vdd.n181 171.744
R18497 vdd.n192 vdd.n181 171.744
R18498 vdd.n192 vdd.n191 171.744
R18499 vdd.n191 vdd.n185 171.744
R18500 vdd.n158 vdd.n157 171.744
R18501 vdd.n157 vdd.n156 171.744
R18502 vdd.n156 vdd.n125 171.744
R18503 vdd.n149 vdd.n125 171.744
R18504 vdd.n149 vdd.n148 171.744
R18505 vdd.n148 vdd.n130 171.744
R18506 vdd.n141 vdd.n130 171.744
R18507 vdd.n141 vdd.n140 171.744
R18508 vdd.n140 vdd.n134 171.744
R18509 vdd.n116 vdd.n115 171.744
R18510 vdd.n115 vdd.n114 171.744
R18511 vdd.n114 vdd.n83 171.744
R18512 vdd.n107 vdd.n83 171.744
R18513 vdd.n107 vdd.n106 171.744
R18514 vdd.n106 vdd.n88 171.744
R18515 vdd.n99 vdd.n88 171.744
R18516 vdd.n99 vdd.n98 171.744
R18517 vdd.n98 vdd.n92 171.744
R18518 vdd.n65 vdd.n64 171.744
R18519 vdd.n64 vdd.n63 171.744
R18520 vdd.n63 vdd.n32 171.744
R18521 vdd.n56 vdd.n32 171.744
R18522 vdd.n56 vdd.n55 171.744
R18523 vdd.n55 vdd.n37 171.744
R18524 vdd.n48 vdd.n37 171.744
R18525 vdd.n48 vdd.n47 171.744
R18526 vdd.n47 vdd.n41 171.744
R18527 vdd.n1953 vdd.n1952 171.744
R18528 vdd.n1952 vdd.n1951 171.744
R18529 vdd.n1951 vdd.n1920 171.744
R18530 vdd.n1944 vdd.n1920 171.744
R18531 vdd.n1944 vdd.n1943 171.744
R18532 vdd.n1943 vdd.n1925 171.744
R18533 vdd.n1936 vdd.n1925 171.744
R18534 vdd.n1936 vdd.n1935 171.744
R18535 vdd.n1935 vdd.n1929 171.744
R18536 vdd.n2004 vdd.n2003 171.744
R18537 vdd.n2003 vdd.n2002 171.744
R18538 vdd.n2002 vdd.n1971 171.744
R18539 vdd.n1995 vdd.n1971 171.744
R18540 vdd.n1995 vdd.n1994 171.744
R18541 vdd.n1994 vdd.n1976 171.744
R18542 vdd.n1987 vdd.n1976 171.744
R18543 vdd.n1987 vdd.n1986 171.744
R18544 vdd.n1986 vdd.n1980 171.744
R18545 vdd.n1859 vdd.n1858 171.744
R18546 vdd.n1858 vdd.n1857 171.744
R18547 vdd.n1857 vdd.n1826 171.744
R18548 vdd.n1850 vdd.n1826 171.744
R18549 vdd.n1850 vdd.n1849 171.744
R18550 vdd.n1849 vdd.n1831 171.744
R18551 vdd.n1842 vdd.n1831 171.744
R18552 vdd.n1842 vdd.n1841 171.744
R18553 vdd.n1841 vdd.n1835 171.744
R18554 vdd.n1910 vdd.n1909 171.744
R18555 vdd.n1909 vdd.n1908 171.744
R18556 vdd.n1908 vdd.n1877 171.744
R18557 vdd.n1901 vdd.n1877 171.744
R18558 vdd.n1901 vdd.n1900 171.744
R18559 vdd.n1900 vdd.n1882 171.744
R18560 vdd.n1893 vdd.n1882 171.744
R18561 vdd.n1893 vdd.n1892 171.744
R18562 vdd.n1892 vdd.n1886 171.744
R18563 vdd.n1766 vdd.n1765 171.744
R18564 vdd.n1765 vdd.n1764 171.744
R18565 vdd.n1764 vdd.n1733 171.744
R18566 vdd.n1757 vdd.n1733 171.744
R18567 vdd.n1757 vdd.n1756 171.744
R18568 vdd.n1756 vdd.n1738 171.744
R18569 vdd.n1749 vdd.n1738 171.744
R18570 vdd.n1749 vdd.n1748 171.744
R18571 vdd.n1748 vdd.n1742 171.744
R18572 vdd.n1817 vdd.n1816 171.744
R18573 vdd.n1816 vdd.n1815 171.744
R18574 vdd.n1815 vdd.n1784 171.744
R18575 vdd.n1808 vdd.n1784 171.744
R18576 vdd.n1808 vdd.n1807 171.744
R18577 vdd.n1807 vdd.n1789 171.744
R18578 vdd.n1800 vdd.n1789 171.744
R18579 vdd.n1800 vdd.n1799 171.744
R18580 vdd.n1799 vdd.n1793 171.744
R18581 vdd.n3402 vdd.n356 146.341
R18582 vdd.n3400 vdd.n3399 146.341
R18583 vdd.n3397 vdd.n360 146.341
R18584 vdd.n3393 vdd.n3392 146.341
R18585 vdd.n3390 vdd.n368 146.341
R18586 vdd.n3386 vdd.n3385 146.341
R18587 vdd.n3383 vdd.n375 146.341
R18588 vdd.n3379 vdd.n3378 146.341
R18589 vdd.n3376 vdd.n382 146.341
R18590 vdd.n393 vdd.n390 146.341
R18591 vdd.n3368 vdd.n3367 146.341
R18592 vdd.n3365 vdd.n395 146.341
R18593 vdd.n3361 vdd.n3360 146.341
R18594 vdd.n3358 vdd.n401 146.341
R18595 vdd.n3354 vdd.n3353 146.341
R18596 vdd.n3351 vdd.n408 146.341
R18597 vdd.n3347 vdd.n3346 146.341
R18598 vdd.n3344 vdd.n415 146.341
R18599 vdd.n3340 vdd.n3339 146.341
R18600 vdd.n3337 vdd.n422 146.341
R18601 vdd.n433 vdd.n430 146.341
R18602 vdd.n3329 vdd.n3328 146.341
R18603 vdd.n3326 vdd.n435 146.341
R18604 vdd.n3322 vdd.n3321 146.341
R18605 vdd.n3319 vdd.n441 146.341
R18606 vdd.n3315 vdd.n3314 146.341
R18607 vdd.n3312 vdd.n448 146.341
R18608 vdd.n3308 vdd.n3307 146.341
R18609 vdd.n3305 vdd.n455 146.341
R18610 vdd.n3301 vdd.n3300 146.341
R18611 vdd.n3298 vdd.n462 146.341
R18612 vdd.n3213 vdd.n512 146.341
R18613 vdd.n3219 vdd.n512 146.341
R18614 vdd.n3219 vdd.n504 146.341
R18615 vdd.n3229 vdd.n504 146.341
R18616 vdd.n3229 vdd.n500 146.341
R18617 vdd.n3235 vdd.n500 146.341
R18618 vdd.n3235 vdd.n491 146.341
R18619 vdd.n3245 vdd.n491 146.341
R18620 vdd.n3245 vdd.n487 146.341
R18621 vdd.n3251 vdd.n487 146.341
R18622 vdd.n3251 vdd.n479 146.341
R18623 vdd.n3262 vdd.n479 146.341
R18624 vdd.n3262 vdd.n480 146.341
R18625 vdd.n480 vdd.n316 146.341
R18626 vdd.n317 vdd.n316 146.341
R18627 vdd.n318 vdd.n317 146.341
R18628 vdd.n473 vdd.n318 146.341
R18629 vdd.n473 vdd.n326 146.341
R18630 vdd.n327 vdd.n326 146.341
R18631 vdd.n328 vdd.n327 146.341
R18632 vdd.n470 vdd.n328 146.341
R18633 vdd.n470 vdd.n337 146.341
R18634 vdd.n338 vdd.n337 146.341
R18635 vdd.n339 vdd.n338 146.341
R18636 vdd.n467 vdd.n339 146.341
R18637 vdd.n467 vdd.n348 146.341
R18638 vdd.n349 vdd.n348 146.341
R18639 vdd.n350 vdd.n349 146.341
R18640 vdd.n3205 vdd.n3203 146.341
R18641 vdd.n3203 vdd.n3202 146.341
R18642 vdd.n3199 vdd.n3198 146.341
R18643 vdd.n3195 vdd.n3194 146.341
R18644 vdd.n3192 vdd.n526 146.341
R18645 vdd.n3188 vdd.n3186 146.341
R18646 vdd.n3184 vdd.n532 146.341
R18647 vdd.n3180 vdd.n3178 146.341
R18648 vdd.n3176 vdd.n538 146.341
R18649 vdd.n3172 vdd.n3170 146.341
R18650 vdd.n3168 vdd.n546 146.341
R18651 vdd.n3164 vdd.n3162 146.341
R18652 vdd.n3160 vdd.n552 146.341
R18653 vdd.n3156 vdd.n3154 146.341
R18654 vdd.n3152 vdd.n558 146.341
R18655 vdd.n3148 vdd.n3146 146.341
R18656 vdd.n3144 vdd.n564 146.341
R18657 vdd.n3140 vdd.n3138 146.341
R18658 vdd.n3136 vdd.n570 146.341
R18659 vdd.n3132 vdd.n3130 146.341
R18660 vdd.n3128 vdd.n576 146.341
R18661 vdd.n3121 vdd.n585 146.341
R18662 vdd.n3119 vdd.n3118 146.341
R18663 vdd.n3115 vdd.n3114 146.341
R18664 vdd.n3112 vdd.n590 146.341
R18665 vdd.n3108 vdd.n3106 146.341
R18666 vdd.n3104 vdd.n596 146.341
R18667 vdd.n3100 vdd.n3098 146.341
R18668 vdd.n3096 vdd.n602 146.341
R18669 vdd.n3092 vdd.n3090 146.341
R18670 vdd.n3087 vdd.n3086 146.341
R18671 vdd.n3083 vdd.n515 146.341
R18672 vdd.n3211 vdd.n510 146.341
R18673 vdd.n3221 vdd.n510 146.341
R18674 vdd.n3221 vdd.n506 146.341
R18675 vdd.n3227 vdd.n506 146.341
R18676 vdd.n3227 vdd.n498 146.341
R18677 vdd.n3237 vdd.n498 146.341
R18678 vdd.n3237 vdd.n494 146.341
R18679 vdd.n3243 vdd.n494 146.341
R18680 vdd.n3243 vdd.n486 146.341
R18681 vdd.n3254 vdd.n486 146.341
R18682 vdd.n3254 vdd.n482 146.341
R18683 vdd.n3260 vdd.n482 146.341
R18684 vdd.n3260 vdd.n314 146.341
R18685 vdd.n3437 vdd.n314 146.341
R18686 vdd.n3437 vdd.n315 146.341
R18687 vdd.n3433 vdd.n315 146.341
R18688 vdd.n3433 vdd.n319 146.341
R18689 vdd.n3429 vdd.n319 146.341
R18690 vdd.n3429 vdd.n324 146.341
R18691 vdd.n3425 vdd.n324 146.341
R18692 vdd.n3425 vdd.n330 146.341
R18693 vdd.n3421 vdd.n330 146.341
R18694 vdd.n3421 vdd.n336 146.341
R18695 vdd.n3417 vdd.n336 146.341
R18696 vdd.n3417 vdd.n341 146.341
R18697 vdd.n3413 vdd.n341 146.341
R18698 vdd.n3413 vdd.n347 146.341
R18699 vdd.n3409 vdd.n347 146.341
R18700 vdd.n2183 vdd.n2182 146.341
R18701 vdd.n2180 vdd.n2177 146.341
R18702 vdd.n2175 vdd.n1013 146.341
R18703 vdd.n2171 vdd.n2170 146.341
R18704 vdd.n2168 vdd.n1017 146.341
R18705 vdd.n2164 vdd.n2163 146.341
R18706 vdd.n2161 vdd.n1024 146.341
R18707 vdd.n2157 vdd.n2156 146.341
R18708 vdd.n2154 vdd.n1031 146.341
R18709 vdd.n1042 vdd.n1039 146.341
R18710 vdd.n2146 vdd.n2145 146.341
R18711 vdd.n2143 vdd.n1044 146.341
R18712 vdd.n2139 vdd.n2138 146.341
R18713 vdd.n2136 vdd.n1050 146.341
R18714 vdd.n2132 vdd.n2131 146.341
R18715 vdd.n2129 vdd.n1057 146.341
R18716 vdd.n2125 vdd.n2124 146.341
R18717 vdd.n2122 vdd.n1064 146.341
R18718 vdd.n2118 vdd.n2117 146.341
R18719 vdd.n2115 vdd.n1071 146.341
R18720 vdd.n1082 vdd.n1079 146.341
R18721 vdd.n2107 vdd.n2106 146.341
R18722 vdd.n2104 vdd.n1084 146.341
R18723 vdd.n2100 vdd.n2099 146.341
R18724 vdd.n2097 vdd.n1090 146.341
R18725 vdd.n2093 vdd.n2092 146.341
R18726 vdd.n2090 vdd.n1097 146.341
R18727 vdd.n2086 vdd.n2085 146.341
R18728 vdd.n2083 vdd.n1104 146.341
R18729 vdd.n1350 vdd.n1348 146.341
R18730 vdd.n1353 vdd.n1352 146.341
R18731 vdd.n1671 vdd.n1433 146.341
R18732 vdd.n1677 vdd.n1433 146.341
R18733 vdd.n1677 vdd.n1426 146.341
R18734 vdd.n1687 vdd.n1426 146.341
R18735 vdd.n1687 vdd.n1422 146.341
R18736 vdd.n1693 vdd.n1422 146.341
R18737 vdd.n1693 vdd.n1413 146.341
R18738 vdd.n1703 vdd.n1413 146.341
R18739 vdd.n1703 vdd.n1409 146.341
R18740 vdd.n1709 vdd.n1409 146.341
R18741 vdd.n1709 vdd.n1402 146.341
R18742 vdd.n1720 vdd.n1402 146.341
R18743 vdd.n1720 vdd.n1398 146.341
R18744 vdd.n1726 vdd.n1398 146.341
R18745 vdd.n1726 vdd.n1391 146.341
R18746 vdd.n2018 vdd.n1391 146.341
R18747 vdd.n2018 vdd.n1387 146.341
R18748 vdd.n2024 vdd.n1387 146.341
R18749 vdd.n2024 vdd.n1379 146.341
R18750 vdd.n2035 vdd.n1379 146.341
R18751 vdd.n2035 vdd.n1375 146.341
R18752 vdd.n2041 vdd.n1375 146.341
R18753 vdd.n2041 vdd.n1369 146.341
R18754 vdd.n2052 vdd.n1369 146.341
R18755 vdd.n2052 vdd.n1364 146.341
R18756 vdd.n2060 vdd.n1364 146.341
R18757 vdd.n2060 vdd.n1355 146.341
R18758 vdd.n2071 vdd.n1355 146.341
R18759 vdd.n1443 vdd.n1442 146.341
R18760 vdd.n1446 vdd.n1443 146.341
R18761 vdd.n1449 vdd.n1448 146.341
R18762 vdd.n1454 vdd.n1451 146.341
R18763 vdd.n1457 vdd.n1456 146.341
R18764 vdd.n1462 vdd.n1459 146.341
R18765 vdd.n1465 vdd.n1464 146.341
R18766 vdd.n1470 vdd.n1467 146.341
R18767 vdd.n1473 vdd.n1472 146.341
R18768 vdd.n1480 vdd.n1475 146.341
R18769 vdd.n1483 vdd.n1482 146.341
R18770 vdd.n1488 vdd.n1485 146.341
R18771 vdd.n1491 vdd.n1490 146.341
R18772 vdd.n1496 vdd.n1493 146.341
R18773 vdd.n1499 vdd.n1498 146.341
R18774 vdd.n1504 vdd.n1501 146.341
R18775 vdd.n1507 vdd.n1506 146.341
R18776 vdd.n1512 vdd.n1509 146.341
R18777 vdd.n1515 vdd.n1514 146.341
R18778 vdd.n1520 vdd.n1517 146.341
R18779 vdd.n1601 vdd.n1522 146.341
R18780 vdd.n1599 vdd.n1598 146.341
R18781 vdd.n1529 vdd.n1528 146.341
R18782 vdd.n1532 vdd.n1531 146.341
R18783 vdd.n1537 vdd.n1536 146.341
R18784 vdd.n1540 vdd.n1539 146.341
R18785 vdd.n1545 vdd.n1544 146.341
R18786 vdd.n1548 vdd.n1547 146.341
R18787 vdd.n1553 vdd.n1552 146.341
R18788 vdd.n1556 vdd.n1555 146.341
R18789 vdd.n1561 vdd.n1560 146.341
R18790 vdd.n1563 vdd.n1436 146.341
R18791 vdd.n1669 vdd.n1432 146.341
R18792 vdd.n1679 vdd.n1432 146.341
R18793 vdd.n1679 vdd.n1428 146.341
R18794 vdd.n1685 vdd.n1428 146.341
R18795 vdd.n1685 vdd.n1420 146.341
R18796 vdd.n1695 vdd.n1420 146.341
R18797 vdd.n1695 vdd.n1416 146.341
R18798 vdd.n1701 vdd.n1416 146.341
R18799 vdd.n1701 vdd.n1408 146.341
R18800 vdd.n1712 vdd.n1408 146.341
R18801 vdd.n1712 vdd.n1404 146.341
R18802 vdd.n1718 vdd.n1404 146.341
R18803 vdd.n1718 vdd.n1397 146.341
R18804 vdd.n1728 vdd.n1397 146.341
R18805 vdd.n1728 vdd.n1393 146.341
R18806 vdd.n2016 vdd.n1393 146.341
R18807 vdd.n2016 vdd.n1385 146.341
R18808 vdd.n2027 vdd.n1385 146.341
R18809 vdd.n2027 vdd.n1381 146.341
R18810 vdd.n2033 vdd.n1381 146.341
R18811 vdd.n2033 vdd.n1374 146.341
R18812 vdd.n2044 vdd.n1374 146.341
R18813 vdd.n2044 vdd.n1370 146.341
R18814 vdd.n2050 vdd.n1370 146.341
R18815 vdd.n2050 vdd.n1362 146.341
R18816 vdd.n2063 vdd.n1362 146.341
R18817 vdd.n2063 vdd.n1357 146.341
R18818 vdd.n2069 vdd.n1357 146.341
R18819 vdd.n1143 vdd.t31 127.284
R18820 vdd.n838 vdd.t75 127.284
R18821 vdd.n1147 vdd.t72 127.284
R18822 vdd.n829 vdd.t98 127.284
R18823 vdd.n724 vdd.t52 127.284
R18824 vdd.n724 vdd.t53 127.284
R18825 vdd.n2535 vdd.t93 127.284
R18826 vdd.n661 vdd.t40 127.284
R18827 vdd.n2532 vdd.t83 127.284
R18828 vdd.n625 vdd.t26 127.284
R18829 vdd.n899 vdd.t89 127.284
R18830 vdd.n899 vdd.t90 127.284
R18831 vdd.n22 vdd.n20 117.314
R18832 vdd.n17 vdd.n15 117.314
R18833 vdd.n27 vdd.n26 116.927
R18834 vdd.n24 vdd.n23 116.927
R18835 vdd.n22 vdd.n21 116.927
R18836 vdd.n17 vdd.n16 116.927
R18837 vdd.n19 vdd.n18 116.927
R18838 vdd.n27 vdd.n25 116.927
R18839 vdd.n1144 vdd.t30 111.188
R18840 vdd.n839 vdd.t76 111.188
R18841 vdd.n1148 vdd.t71 111.188
R18842 vdd.n830 vdd.t99 111.188
R18843 vdd.n2536 vdd.t92 111.188
R18844 vdd.n662 vdd.t41 111.188
R18845 vdd.n2533 vdd.t82 111.188
R18846 vdd.n626 vdd.t27 111.188
R18847 vdd.n2806 vdd.n788 99.5127
R18848 vdd.n2806 vdd.n779 99.5127
R18849 vdd.n2814 vdd.n779 99.5127
R18850 vdd.n2814 vdd.n777 99.5127
R18851 vdd.n2818 vdd.n777 99.5127
R18852 vdd.n2818 vdd.n767 99.5127
R18853 vdd.n2826 vdd.n767 99.5127
R18854 vdd.n2826 vdd.n765 99.5127
R18855 vdd.n2830 vdd.n765 99.5127
R18856 vdd.n2830 vdd.n756 99.5127
R18857 vdd.n2838 vdd.n756 99.5127
R18858 vdd.n2838 vdd.n754 99.5127
R18859 vdd.n2842 vdd.n754 99.5127
R18860 vdd.n2842 vdd.n745 99.5127
R18861 vdd.n2850 vdd.n745 99.5127
R18862 vdd.n2850 vdd.n743 99.5127
R18863 vdd.n2854 vdd.n743 99.5127
R18864 vdd.n2854 vdd.n732 99.5127
R18865 vdd.n2863 vdd.n732 99.5127
R18866 vdd.n2863 vdd.n730 99.5127
R18867 vdd.n2867 vdd.n730 99.5127
R18868 vdd.n2867 vdd.n720 99.5127
R18869 vdd.n2875 vdd.n720 99.5127
R18870 vdd.n2875 vdd.n718 99.5127
R18871 vdd.n2879 vdd.n718 99.5127
R18872 vdd.n2879 vdd.n708 99.5127
R18873 vdd.n2887 vdd.n708 99.5127
R18874 vdd.n2887 vdd.n706 99.5127
R18875 vdd.n2891 vdd.n706 99.5127
R18876 vdd.n2891 vdd.n695 99.5127
R18877 vdd.n2899 vdd.n695 99.5127
R18878 vdd.n2899 vdd.n693 99.5127
R18879 vdd.n2903 vdd.n693 99.5127
R18880 vdd.n2903 vdd.n684 99.5127
R18881 vdd.n2911 vdd.n684 99.5127
R18882 vdd.n2911 vdd.n682 99.5127
R18883 vdd.n2915 vdd.n682 99.5127
R18884 vdd.n2915 vdd.n670 99.5127
R18885 vdd.n2968 vdd.n670 99.5127
R18886 vdd.n2968 vdd.n668 99.5127
R18887 vdd.n2972 vdd.n668 99.5127
R18888 vdd.n2972 vdd.n634 99.5127
R18889 vdd.n3042 vdd.n634 99.5127
R18890 vdd.n3038 vdd.n635 99.5127
R18891 vdd.n3036 vdd.n3035 99.5127
R18892 vdd.n3033 vdd.n639 99.5127
R18893 vdd.n3029 vdd.n3028 99.5127
R18894 vdd.n3026 vdd.n642 99.5127
R18895 vdd.n3022 vdd.n3021 99.5127
R18896 vdd.n3019 vdd.n645 99.5127
R18897 vdd.n3015 vdd.n3014 99.5127
R18898 vdd.n3012 vdd.n648 99.5127
R18899 vdd.n3007 vdd.n3006 99.5127
R18900 vdd.n3004 vdd.n651 99.5127
R18901 vdd.n3000 vdd.n2999 99.5127
R18902 vdd.n2997 vdd.n654 99.5127
R18903 vdd.n2993 vdd.n2992 99.5127
R18904 vdd.n2990 vdd.n657 99.5127
R18905 vdd.n2986 vdd.n2985 99.5127
R18906 vdd.n2983 vdd.n660 99.5127
R18907 vdd.n2733 vdd.n786 99.5127
R18908 vdd.n2729 vdd.n786 99.5127
R18909 vdd.n2729 vdd.n780 99.5127
R18910 vdd.n2611 vdd.n780 99.5127
R18911 vdd.n2611 vdd.n775 99.5127
R18912 vdd.n2614 vdd.n775 99.5127
R18913 vdd.n2614 vdd.n769 99.5127
R18914 vdd.n2715 vdd.n769 99.5127
R18915 vdd.n2715 vdd.n763 99.5127
R18916 vdd.n2711 vdd.n763 99.5127
R18917 vdd.n2711 vdd.n757 99.5127
R18918 vdd.n2658 vdd.n757 99.5127
R18919 vdd.n2658 vdd.n751 99.5127
R18920 vdd.n2655 vdd.n751 99.5127
R18921 vdd.n2655 vdd.n746 99.5127
R18922 vdd.n2652 vdd.n746 99.5127
R18923 vdd.n2652 vdd.n741 99.5127
R18924 vdd.n2649 vdd.n741 99.5127
R18925 vdd.n2649 vdd.n734 99.5127
R18926 vdd.n2646 vdd.n734 99.5127
R18927 vdd.n2646 vdd.n727 99.5127
R18928 vdd.n2643 vdd.n727 99.5127
R18929 vdd.n2643 vdd.n721 99.5127
R18930 vdd.n2640 vdd.n721 99.5127
R18931 vdd.n2640 vdd.n716 99.5127
R18932 vdd.n2637 vdd.n716 99.5127
R18933 vdd.n2637 vdd.n710 99.5127
R18934 vdd.n2634 vdd.n710 99.5127
R18935 vdd.n2634 vdd.n703 99.5127
R18936 vdd.n2631 vdd.n703 99.5127
R18937 vdd.n2631 vdd.n696 99.5127
R18938 vdd.n2628 vdd.n696 99.5127
R18939 vdd.n2628 vdd.n690 99.5127
R18940 vdd.n2625 vdd.n690 99.5127
R18941 vdd.n2625 vdd.n685 99.5127
R18942 vdd.n2622 vdd.n685 99.5127
R18943 vdd.n2622 vdd.n680 99.5127
R18944 vdd.n2619 vdd.n680 99.5127
R18945 vdd.n2619 vdd.n672 99.5127
R18946 vdd.n672 vdd.n665 99.5127
R18947 vdd.n2974 vdd.n665 99.5127
R18948 vdd.n2975 vdd.n2974 99.5127
R18949 vdd.n2975 vdd.n632 99.5127
R18950 vdd.n2799 vdd.n790 99.5127
R18951 vdd.n2799 vdd.n2531 99.5127
R18952 vdd.n2795 vdd.n2794 99.5127
R18953 vdd.n2791 vdd.n2790 99.5127
R18954 vdd.n2787 vdd.n2786 99.5127
R18955 vdd.n2783 vdd.n2782 99.5127
R18956 vdd.n2779 vdd.n2778 99.5127
R18957 vdd.n2775 vdd.n2774 99.5127
R18958 vdd.n2771 vdd.n2770 99.5127
R18959 vdd.n2767 vdd.n2766 99.5127
R18960 vdd.n2763 vdd.n2762 99.5127
R18961 vdd.n2759 vdd.n2758 99.5127
R18962 vdd.n2755 vdd.n2754 99.5127
R18963 vdd.n2751 vdd.n2750 99.5127
R18964 vdd.n2747 vdd.n2746 99.5127
R18965 vdd.n2743 vdd.n2742 99.5127
R18966 vdd.n2738 vdd.n2737 99.5127
R18967 vdd.n2495 vdd.n827 99.5127
R18968 vdd.n2491 vdd.n2490 99.5127
R18969 vdd.n2487 vdd.n2486 99.5127
R18970 vdd.n2483 vdd.n2482 99.5127
R18971 vdd.n2479 vdd.n2478 99.5127
R18972 vdd.n2475 vdd.n2474 99.5127
R18973 vdd.n2471 vdd.n2470 99.5127
R18974 vdd.n2467 vdd.n2466 99.5127
R18975 vdd.n2463 vdd.n2462 99.5127
R18976 vdd.n2459 vdd.n2458 99.5127
R18977 vdd.n2455 vdd.n2454 99.5127
R18978 vdd.n2451 vdd.n2450 99.5127
R18979 vdd.n2447 vdd.n2446 99.5127
R18980 vdd.n2443 vdd.n2442 99.5127
R18981 vdd.n2439 vdd.n2438 99.5127
R18982 vdd.n2435 vdd.n2434 99.5127
R18983 vdd.n2430 vdd.n2429 99.5127
R18984 vdd.n1183 vdd.n963 99.5127
R18985 vdd.n1186 vdd.n963 99.5127
R18986 vdd.n1186 vdd.n957 99.5127
R18987 vdd.n1189 vdd.n957 99.5127
R18988 vdd.n1189 vdd.n952 99.5127
R18989 vdd.n1192 vdd.n952 99.5127
R18990 vdd.n1192 vdd.n945 99.5127
R18991 vdd.n1195 vdd.n945 99.5127
R18992 vdd.n1195 vdd.n938 99.5127
R18993 vdd.n1198 vdd.n938 99.5127
R18994 vdd.n1198 vdd.n932 99.5127
R18995 vdd.n1201 vdd.n932 99.5127
R18996 vdd.n1201 vdd.n927 99.5127
R18997 vdd.n1204 vdd.n927 99.5127
R18998 vdd.n1204 vdd.n922 99.5127
R18999 vdd.n1207 vdd.n922 99.5127
R19000 vdd.n1207 vdd.n916 99.5127
R19001 vdd.n1210 vdd.n916 99.5127
R19002 vdd.n1210 vdd.n909 99.5127
R19003 vdd.n1213 vdd.n909 99.5127
R19004 vdd.n1213 vdd.n902 99.5127
R19005 vdd.n1216 vdd.n902 99.5127
R19006 vdd.n1216 vdd.n896 99.5127
R19007 vdd.n1219 vdd.n896 99.5127
R19008 vdd.n1219 vdd.n891 99.5127
R19009 vdd.n1222 vdd.n891 99.5127
R19010 vdd.n1222 vdd.n885 99.5127
R19011 vdd.n1264 vdd.n885 99.5127
R19012 vdd.n1264 vdd.n878 99.5127
R19013 vdd.n1260 vdd.n878 99.5127
R19014 vdd.n1260 vdd.n872 99.5127
R19015 vdd.n1257 vdd.n872 99.5127
R19016 vdd.n1257 vdd.n867 99.5127
R19017 vdd.n1254 vdd.n867 99.5127
R19018 vdd.n1254 vdd.n862 99.5127
R19019 vdd.n1234 vdd.n862 99.5127
R19020 vdd.n1234 vdd.n857 99.5127
R19021 vdd.n1231 vdd.n857 99.5127
R19022 vdd.n1231 vdd.n850 99.5127
R19023 vdd.n1228 vdd.n850 99.5127
R19024 vdd.n1228 vdd.n843 99.5127
R19025 vdd.n843 vdd.n832 99.5127
R19026 vdd.n2425 vdd.n832 99.5127
R19027 vdd.n2217 vdd.n968 99.5127
R19028 vdd.n2217 vdd.n1004 99.5127
R19029 vdd.n2213 vdd.n2212 99.5127
R19030 vdd.n2209 vdd.n2208 99.5127
R19031 vdd.n2205 vdd.n2204 99.5127
R19032 vdd.n2201 vdd.n2200 99.5127
R19033 vdd.n2197 vdd.n2196 99.5127
R19034 vdd.n2193 vdd.n2192 99.5127
R19035 vdd.n2189 vdd.n2188 99.5127
R19036 vdd.n1150 vdd.n1149 99.5127
R19037 vdd.n1154 vdd.n1153 99.5127
R19038 vdd.n1158 vdd.n1157 99.5127
R19039 vdd.n1162 vdd.n1161 99.5127
R19040 vdd.n1166 vdd.n1165 99.5127
R19041 vdd.n1170 vdd.n1169 99.5127
R19042 vdd.n1174 vdd.n1173 99.5127
R19043 vdd.n1179 vdd.n1178 99.5127
R19044 vdd.n2224 vdd.n966 99.5127
R19045 vdd.n2224 vdd.n956 99.5127
R19046 vdd.n2232 vdd.n956 99.5127
R19047 vdd.n2232 vdd.n954 99.5127
R19048 vdd.n2236 vdd.n954 99.5127
R19049 vdd.n2236 vdd.n943 99.5127
R19050 vdd.n2244 vdd.n943 99.5127
R19051 vdd.n2244 vdd.n941 99.5127
R19052 vdd.n2248 vdd.n941 99.5127
R19053 vdd.n2248 vdd.n931 99.5127
R19054 vdd.n2256 vdd.n931 99.5127
R19055 vdd.n2256 vdd.n929 99.5127
R19056 vdd.n2260 vdd.n929 99.5127
R19057 vdd.n2260 vdd.n920 99.5127
R19058 vdd.n2268 vdd.n920 99.5127
R19059 vdd.n2268 vdd.n918 99.5127
R19060 vdd.n2272 vdd.n918 99.5127
R19061 vdd.n2272 vdd.n907 99.5127
R19062 vdd.n2280 vdd.n907 99.5127
R19063 vdd.n2280 vdd.n905 99.5127
R19064 vdd.n2284 vdd.n905 99.5127
R19065 vdd.n2284 vdd.n895 99.5127
R19066 vdd.n2293 vdd.n895 99.5127
R19067 vdd.n2293 vdd.n893 99.5127
R19068 vdd.n2297 vdd.n893 99.5127
R19069 vdd.n2297 vdd.n883 99.5127
R19070 vdd.n2305 vdd.n883 99.5127
R19071 vdd.n2305 vdd.n881 99.5127
R19072 vdd.n2309 vdd.n881 99.5127
R19073 vdd.n2309 vdd.n871 99.5127
R19074 vdd.n2317 vdd.n871 99.5127
R19075 vdd.n2317 vdd.n869 99.5127
R19076 vdd.n2321 vdd.n869 99.5127
R19077 vdd.n2321 vdd.n861 99.5127
R19078 vdd.n2329 vdd.n861 99.5127
R19079 vdd.n2329 vdd.n859 99.5127
R19080 vdd.n2333 vdd.n859 99.5127
R19081 vdd.n2333 vdd.n848 99.5127
R19082 vdd.n2343 vdd.n848 99.5127
R19083 vdd.n2343 vdd.n845 99.5127
R19084 vdd.n2348 vdd.n845 99.5127
R19085 vdd.n2348 vdd.n846 99.5127
R19086 vdd.n846 vdd.n826 99.5127
R19087 vdd.n2958 vdd.n2957 99.5127
R19088 vdd.n2955 vdd.n2921 99.5127
R19089 vdd.n2951 vdd.n2950 99.5127
R19090 vdd.n2948 vdd.n2924 99.5127
R19091 vdd.n2944 vdd.n2943 99.5127
R19092 vdd.n2941 vdd.n2927 99.5127
R19093 vdd.n2937 vdd.n2936 99.5127
R19094 vdd.n2934 vdd.n2931 99.5127
R19095 vdd.n3075 vdd.n612 99.5127
R19096 vdd.n3073 vdd.n3072 99.5127
R19097 vdd.n3070 vdd.n615 99.5127
R19098 vdd.n3066 vdd.n3065 99.5127
R19099 vdd.n3063 vdd.n618 99.5127
R19100 vdd.n3059 vdd.n3058 99.5127
R19101 vdd.n3056 vdd.n621 99.5127
R19102 vdd.n3052 vdd.n3051 99.5127
R19103 vdd.n3049 vdd.n624 99.5127
R19104 vdd.n2607 vdd.n787 99.5127
R19105 vdd.n2727 vdd.n787 99.5127
R19106 vdd.n2727 vdd.n781 99.5127
R19107 vdd.n2723 vdd.n781 99.5127
R19108 vdd.n2723 vdd.n776 99.5127
R19109 vdd.n2720 vdd.n776 99.5127
R19110 vdd.n2720 vdd.n770 99.5127
R19111 vdd.n2717 vdd.n770 99.5127
R19112 vdd.n2717 vdd.n764 99.5127
R19113 vdd.n2709 vdd.n764 99.5127
R19114 vdd.n2709 vdd.n758 99.5127
R19115 vdd.n2705 vdd.n758 99.5127
R19116 vdd.n2705 vdd.n752 99.5127
R19117 vdd.n2702 vdd.n752 99.5127
R19118 vdd.n2702 vdd.n747 99.5127
R19119 vdd.n2699 vdd.n747 99.5127
R19120 vdd.n2699 vdd.n742 99.5127
R19121 vdd.n2696 vdd.n742 99.5127
R19122 vdd.n2696 vdd.n735 99.5127
R19123 vdd.n2693 vdd.n735 99.5127
R19124 vdd.n2693 vdd.n728 99.5127
R19125 vdd.n2690 vdd.n728 99.5127
R19126 vdd.n2690 vdd.n722 99.5127
R19127 vdd.n2687 vdd.n722 99.5127
R19128 vdd.n2687 vdd.n717 99.5127
R19129 vdd.n2684 vdd.n717 99.5127
R19130 vdd.n2684 vdd.n711 99.5127
R19131 vdd.n2681 vdd.n711 99.5127
R19132 vdd.n2681 vdd.n704 99.5127
R19133 vdd.n2678 vdd.n704 99.5127
R19134 vdd.n2678 vdd.n697 99.5127
R19135 vdd.n2675 vdd.n697 99.5127
R19136 vdd.n2675 vdd.n691 99.5127
R19137 vdd.n2672 vdd.n691 99.5127
R19138 vdd.n2672 vdd.n686 99.5127
R19139 vdd.n2669 vdd.n686 99.5127
R19140 vdd.n2669 vdd.n681 99.5127
R19141 vdd.n2666 vdd.n681 99.5127
R19142 vdd.n2666 vdd.n673 99.5127
R19143 vdd.n2663 vdd.n673 99.5127
R19144 vdd.n2663 vdd.n666 99.5127
R19145 vdd.n666 vdd.n630 99.5127
R19146 vdd.n3044 vdd.n630 99.5127
R19147 vdd.n2542 vdd.n2541 99.5127
R19148 vdd.n2546 vdd.n2545 99.5127
R19149 vdd.n2550 vdd.n2549 99.5127
R19150 vdd.n2554 vdd.n2553 99.5127
R19151 vdd.n2558 vdd.n2557 99.5127
R19152 vdd.n2562 vdd.n2561 99.5127
R19153 vdd.n2566 vdd.n2565 99.5127
R19154 vdd.n2570 vdd.n2569 99.5127
R19155 vdd.n2574 vdd.n2573 99.5127
R19156 vdd.n2578 vdd.n2577 99.5127
R19157 vdd.n2582 vdd.n2581 99.5127
R19158 vdd.n2586 vdd.n2585 99.5127
R19159 vdd.n2590 vdd.n2589 99.5127
R19160 vdd.n2594 vdd.n2593 99.5127
R19161 vdd.n2598 vdd.n2597 99.5127
R19162 vdd.n2602 vdd.n2601 99.5127
R19163 vdd.n2604 vdd.n2530 99.5127
R19164 vdd.n2808 vdd.n784 99.5127
R19165 vdd.n2808 vdd.n782 99.5127
R19166 vdd.n2812 vdd.n782 99.5127
R19167 vdd.n2812 vdd.n773 99.5127
R19168 vdd.n2820 vdd.n773 99.5127
R19169 vdd.n2820 vdd.n771 99.5127
R19170 vdd.n2824 vdd.n771 99.5127
R19171 vdd.n2824 vdd.n762 99.5127
R19172 vdd.n2832 vdd.n762 99.5127
R19173 vdd.n2832 vdd.n760 99.5127
R19174 vdd.n2836 vdd.n760 99.5127
R19175 vdd.n2836 vdd.n750 99.5127
R19176 vdd.n2844 vdd.n750 99.5127
R19177 vdd.n2844 vdd.n748 99.5127
R19178 vdd.n2848 vdd.n748 99.5127
R19179 vdd.n2848 vdd.n739 99.5127
R19180 vdd.n2856 vdd.n739 99.5127
R19181 vdd.n2856 vdd.n737 99.5127
R19182 vdd.n2861 vdd.n737 99.5127
R19183 vdd.n2861 vdd.n726 99.5127
R19184 vdd.n2869 vdd.n726 99.5127
R19185 vdd.n2869 vdd.n723 99.5127
R19186 vdd.n2873 vdd.n723 99.5127
R19187 vdd.n2873 vdd.n714 99.5127
R19188 vdd.n2881 vdd.n714 99.5127
R19189 vdd.n2881 vdd.n712 99.5127
R19190 vdd.n2885 vdd.n712 99.5127
R19191 vdd.n2885 vdd.n701 99.5127
R19192 vdd.n2893 vdd.n701 99.5127
R19193 vdd.n2893 vdd.n699 99.5127
R19194 vdd.n2897 vdd.n699 99.5127
R19195 vdd.n2897 vdd.n689 99.5127
R19196 vdd.n2905 vdd.n689 99.5127
R19197 vdd.n2905 vdd.n687 99.5127
R19198 vdd.n2909 vdd.n687 99.5127
R19199 vdd.n2909 vdd.n678 99.5127
R19200 vdd.n2917 vdd.n678 99.5127
R19201 vdd.n2917 vdd.n675 99.5127
R19202 vdd.n2966 vdd.n675 99.5127
R19203 vdd.n2966 vdd.n676 99.5127
R19204 vdd.n676 vdd.n667 99.5127
R19205 vdd.n2961 vdd.n667 99.5127
R19206 vdd.n2961 vdd.n633 99.5127
R19207 vdd.n2419 vdd.n2418 99.5127
R19208 vdd.n2415 vdd.n2414 99.5127
R19209 vdd.n2411 vdd.n2410 99.5127
R19210 vdd.n2407 vdd.n2406 99.5127
R19211 vdd.n2403 vdd.n2402 99.5127
R19212 vdd.n2399 vdd.n2398 99.5127
R19213 vdd.n2395 vdd.n2394 99.5127
R19214 vdd.n2391 vdd.n2390 99.5127
R19215 vdd.n2387 vdd.n2386 99.5127
R19216 vdd.n2383 vdd.n2382 99.5127
R19217 vdd.n2379 vdd.n2378 99.5127
R19218 vdd.n2375 vdd.n2374 99.5127
R19219 vdd.n2371 vdd.n2370 99.5127
R19220 vdd.n2367 vdd.n2366 99.5127
R19221 vdd.n2363 vdd.n2362 99.5127
R19222 vdd.n2359 vdd.n2358 99.5127
R19223 vdd.n2355 vdd.n808 99.5127
R19224 vdd.n1308 vdd.n964 99.5127
R19225 vdd.n1305 vdd.n964 99.5127
R19226 vdd.n1305 vdd.n958 99.5127
R19227 vdd.n1302 vdd.n958 99.5127
R19228 vdd.n1302 vdd.n953 99.5127
R19229 vdd.n1299 vdd.n953 99.5127
R19230 vdd.n1299 vdd.n946 99.5127
R19231 vdd.n1296 vdd.n946 99.5127
R19232 vdd.n1296 vdd.n939 99.5127
R19233 vdd.n1293 vdd.n939 99.5127
R19234 vdd.n1293 vdd.n933 99.5127
R19235 vdd.n1290 vdd.n933 99.5127
R19236 vdd.n1290 vdd.n928 99.5127
R19237 vdd.n1287 vdd.n928 99.5127
R19238 vdd.n1287 vdd.n923 99.5127
R19239 vdd.n1284 vdd.n923 99.5127
R19240 vdd.n1284 vdd.n917 99.5127
R19241 vdd.n1281 vdd.n917 99.5127
R19242 vdd.n1281 vdd.n910 99.5127
R19243 vdd.n1278 vdd.n910 99.5127
R19244 vdd.n1278 vdd.n903 99.5127
R19245 vdd.n1275 vdd.n903 99.5127
R19246 vdd.n1275 vdd.n897 99.5127
R19247 vdd.n1272 vdd.n897 99.5127
R19248 vdd.n1272 vdd.n892 99.5127
R19249 vdd.n1269 vdd.n892 99.5127
R19250 vdd.n1269 vdd.n886 99.5127
R19251 vdd.n1266 vdd.n886 99.5127
R19252 vdd.n1266 vdd.n879 99.5127
R19253 vdd.n1237 vdd.n879 99.5127
R19254 vdd.n1237 vdd.n873 99.5127
R19255 vdd.n1240 vdd.n873 99.5127
R19256 vdd.n1240 vdd.n868 99.5127
R19257 vdd.n1252 vdd.n868 99.5127
R19258 vdd.n1252 vdd.n863 99.5127
R19259 vdd.n1248 vdd.n863 99.5127
R19260 vdd.n1248 vdd.n858 99.5127
R19261 vdd.n1245 vdd.n858 99.5127
R19262 vdd.n1245 vdd.n851 99.5127
R19263 vdd.n851 vdd.n842 99.5127
R19264 vdd.n2350 vdd.n842 99.5127
R19265 vdd.n2351 vdd.n2350 99.5127
R19266 vdd.n2351 vdd.n834 99.5127
R19267 vdd.n1112 vdd.n1111 99.5127
R19268 vdd.n1116 vdd.n1115 99.5127
R19269 vdd.n1120 vdd.n1119 99.5127
R19270 vdd.n1124 vdd.n1123 99.5127
R19271 vdd.n1128 vdd.n1127 99.5127
R19272 vdd.n1132 vdd.n1131 99.5127
R19273 vdd.n1136 vdd.n1135 99.5127
R19274 vdd.n1140 vdd.n1139 99.5127
R19275 vdd.n1341 vdd.n1142 99.5127
R19276 vdd.n1339 vdd.n1338 99.5127
R19277 vdd.n1335 vdd.n1334 99.5127
R19278 vdd.n1331 vdd.n1330 99.5127
R19279 vdd.n1327 vdd.n1326 99.5127
R19280 vdd.n1323 vdd.n1322 99.5127
R19281 vdd.n1319 vdd.n1318 99.5127
R19282 vdd.n1315 vdd.n1314 99.5127
R19283 vdd.n1311 vdd.n1003 99.5127
R19284 vdd.n2226 vdd.n961 99.5127
R19285 vdd.n2226 vdd.n959 99.5127
R19286 vdd.n2230 vdd.n959 99.5127
R19287 vdd.n2230 vdd.n950 99.5127
R19288 vdd.n2238 vdd.n950 99.5127
R19289 vdd.n2238 vdd.n948 99.5127
R19290 vdd.n2242 vdd.n948 99.5127
R19291 vdd.n2242 vdd.n937 99.5127
R19292 vdd.n2250 vdd.n937 99.5127
R19293 vdd.n2250 vdd.n935 99.5127
R19294 vdd.n2254 vdd.n935 99.5127
R19295 vdd.n2254 vdd.n926 99.5127
R19296 vdd.n2262 vdd.n926 99.5127
R19297 vdd.n2262 vdd.n924 99.5127
R19298 vdd.n2266 vdd.n924 99.5127
R19299 vdd.n2266 vdd.n914 99.5127
R19300 vdd.n2274 vdd.n914 99.5127
R19301 vdd.n2274 vdd.n912 99.5127
R19302 vdd.n2278 vdd.n912 99.5127
R19303 vdd.n2278 vdd.n901 99.5127
R19304 vdd.n2286 vdd.n901 99.5127
R19305 vdd.n2286 vdd.n898 99.5127
R19306 vdd.n2291 vdd.n898 99.5127
R19307 vdd.n2291 vdd.n889 99.5127
R19308 vdd.n2299 vdd.n889 99.5127
R19309 vdd.n2299 vdd.n887 99.5127
R19310 vdd.n2303 vdd.n887 99.5127
R19311 vdd.n2303 vdd.n877 99.5127
R19312 vdd.n2311 vdd.n877 99.5127
R19313 vdd.n2311 vdd.n875 99.5127
R19314 vdd.n2315 vdd.n875 99.5127
R19315 vdd.n2315 vdd.n866 99.5127
R19316 vdd.n2323 vdd.n866 99.5127
R19317 vdd.n2323 vdd.n864 99.5127
R19318 vdd.n2327 vdd.n864 99.5127
R19319 vdd.n2327 vdd.n855 99.5127
R19320 vdd.n2335 vdd.n855 99.5127
R19321 vdd.n2335 vdd.n852 99.5127
R19322 vdd.n2341 vdd.n852 99.5127
R19323 vdd.n2341 vdd.n853 99.5127
R19324 vdd.n853 vdd.n844 99.5127
R19325 vdd.n844 vdd.n835 99.5127
R19326 vdd.n2423 vdd.n835 99.5127
R19327 vdd.n9 vdd.n7 98.9633
R19328 vdd.n2 vdd.n0 98.9633
R19329 vdd.n9 vdd.n8 98.6055
R19330 vdd.n11 vdd.n10 98.6055
R19331 vdd.n13 vdd.n12 98.6055
R19332 vdd.n6 vdd.n5 98.6055
R19333 vdd.n4 vdd.n3 98.6055
R19334 vdd.n2 vdd.n1 98.6055
R19335 vdd.t144 vdd.n279 85.8723
R19336 vdd.t3 vdd.n228 85.8723
R19337 vdd.t23 vdd.n185 85.8723
R19338 vdd.t219 vdd.n134 85.8723
R19339 vdd.t154 vdd.n92 85.8723
R19340 vdd.t16 vdd.n41 85.8723
R19341 vdd.t220 vdd.n1929 85.8723
R19342 vdd.t132 vdd.n1980 85.8723
R19343 vdd.t102 vdd.n1835 85.8723
R19344 vdd.t153 vdd.n1886 85.8723
R19345 vdd.t15 vdd.n1742 85.8723
R19346 vdd.t240 vdd.n1793 85.8723
R19347 vdd.n725 vdd.n724 78.546
R19348 vdd.n2289 vdd.n899 78.546
R19349 vdd.n266 vdd.n265 75.1835
R19350 vdd.n264 vdd.n263 75.1835
R19351 vdd.n262 vdd.n261 75.1835
R19352 vdd.n260 vdd.n259 75.1835
R19353 vdd.n258 vdd.n257 75.1835
R19354 vdd.n172 vdd.n171 75.1835
R19355 vdd.n170 vdd.n169 75.1835
R19356 vdd.n168 vdd.n167 75.1835
R19357 vdd.n166 vdd.n165 75.1835
R19358 vdd.n164 vdd.n163 75.1835
R19359 vdd.n79 vdd.n78 75.1835
R19360 vdd.n77 vdd.n76 75.1835
R19361 vdd.n75 vdd.n74 75.1835
R19362 vdd.n73 vdd.n72 75.1835
R19363 vdd.n71 vdd.n70 75.1835
R19364 vdd.n1959 vdd.n1958 75.1835
R19365 vdd.n1961 vdd.n1960 75.1835
R19366 vdd.n1963 vdd.n1962 75.1835
R19367 vdd.n1965 vdd.n1964 75.1835
R19368 vdd.n1967 vdd.n1966 75.1835
R19369 vdd.n1865 vdd.n1864 75.1835
R19370 vdd.n1867 vdd.n1866 75.1835
R19371 vdd.n1869 vdd.n1868 75.1835
R19372 vdd.n1871 vdd.n1870 75.1835
R19373 vdd.n1873 vdd.n1872 75.1835
R19374 vdd.n1772 vdd.n1771 75.1835
R19375 vdd.n1774 vdd.n1773 75.1835
R19376 vdd.n1776 vdd.n1775 75.1835
R19377 vdd.n1778 vdd.n1777 75.1835
R19378 vdd.n1780 vdd.n1779 75.1835
R19379 vdd.n2800 vdd.n2513 72.8958
R19380 vdd.n2800 vdd.n2514 72.8958
R19381 vdd.n2800 vdd.n2515 72.8958
R19382 vdd.n2800 vdd.n2516 72.8958
R19383 vdd.n2800 vdd.n2517 72.8958
R19384 vdd.n2800 vdd.n2518 72.8958
R19385 vdd.n2800 vdd.n2519 72.8958
R19386 vdd.n2800 vdd.n2520 72.8958
R19387 vdd.n2800 vdd.n2521 72.8958
R19388 vdd.n2800 vdd.n2522 72.8958
R19389 vdd.n2800 vdd.n2523 72.8958
R19390 vdd.n2800 vdd.n2524 72.8958
R19391 vdd.n2800 vdd.n2525 72.8958
R19392 vdd.n2800 vdd.n2526 72.8958
R19393 vdd.n2800 vdd.n2527 72.8958
R19394 vdd.n2800 vdd.n2528 72.8958
R19395 vdd.n2800 vdd.n2529 72.8958
R19396 vdd.n629 vdd.n613 72.8958
R19397 vdd.n3050 vdd.n613 72.8958
R19398 vdd.n623 vdd.n613 72.8958
R19399 vdd.n3057 vdd.n613 72.8958
R19400 vdd.n620 vdd.n613 72.8958
R19401 vdd.n3064 vdd.n613 72.8958
R19402 vdd.n617 vdd.n613 72.8958
R19403 vdd.n3071 vdd.n613 72.8958
R19404 vdd.n3074 vdd.n613 72.8958
R19405 vdd.n2930 vdd.n613 72.8958
R19406 vdd.n2935 vdd.n613 72.8958
R19407 vdd.n2929 vdd.n613 72.8958
R19408 vdd.n2942 vdd.n613 72.8958
R19409 vdd.n2926 vdd.n613 72.8958
R19410 vdd.n2949 vdd.n613 72.8958
R19411 vdd.n2923 vdd.n613 72.8958
R19412 vdd.n2956 vdd.n613 72.8958
R19413 vdd.n2219 vdd.n2218 72.8958
R19414 vdd.n2218 vdd.n970 72.8958
R19415 vdd.n2218 vdd.n971 72.8958
R19416 vdd.n2218 vdd.n972 72.8958
R19417 vdd.n2218 vdd.n973 72.8958
R19418 vdd.n2218 vdd.n974 72.8958
R19419 vdd.n2218 vdd.n975 72.8958
R19420 vdd.n2218 vdd.n976 72.8958
R19421 vdd.n2218 vdd.n977 72.8958
R19422 vdd.n2218 vdd.n978 72.8958
R19423 vdd.n2218 vdd.n979 72.8958
R19424 vdd.n2218 vdd.n980 72.8958
R19425 vdd.n2218 vdd.n981 72.8958
R19426 vdd.n2218 vdd.n982 72.8958
R19427 vdd.n2218 vdd.n983 72.8958
R19428 vdd.n2218 vdd.n984 72.8958
R19429 vdd.n2218 vdd.n985 72.8958
R19430 vdd.n2496 vdd.n809 72.8958
R19431 vdd.n2496 vdd.n810 72.8958
R19432 vdd.n2496 vdd.n811 72.8958
R19433 vdd.n2496 vdd.n812 72.8958
R19434 vdd.n2496 vdd.n813 72.8958
R19435 vdd.n2496 vdd.n814 72.8958
R19436 vdd.n2496 vdd.n815 72.8958
R19437 vdd.n2496 vdd.n816 72.8958
R19438 vdd.n2496 vdd.n817 72.8958
R19439 vdd.n2496 vdd.n818 72.8958
R19440 vdd.n2496 vdd.n819 72.8958
R19441 vdd.n2496 vdd.n820 72.8958
R19442 vdd.n2496 vdd.n821 72.8958
R19443 vdd.n2496 vdd.n822 72.8958
R19444 vdd.n2496 vdd.n823 72.8958
R19445 vdd.n2496 vdd.n824 72.8958
R19446 vdd.n2496 vdd.n825 72.8958
R19447 vdd.n2801 vdd.n2800 72.8958
R19448 vdd.n2800 vdd.n2497 72.8958
R19449 vdd.n2800 vdd.n2498 72.8958
R19450 vdd.n2800 vdd.n2499 72.8958
R19451 vdd.n2800 vdd.n2500 72.8958
R19452 vdd.n2800 vdd.n2501 72.8958
R19453 vdd.n2800 vdd.n2502 72.8958
R19454 vdd.n2800 vdd.n2503 72.8958
R19455 vdd.n2800 vdd.n2504 72.8958
R19456 vdd.n2800 vdd.n2505 72.8958
R19457 vdd.n2800 vdd.n2506 72.8958
R19458 vdd.n2800 vdd.n2507 72.8958
R19459 vdd.n2800 vdd.n2508 72.8958
R19460 vdd.n2800 vdd.n2509 72.8958
R19461 vdd.n2800 vdd.n2510 72.8958
R19462 vdd.n2800 vdd.n2511 72.8958
R19463 vdd.n2800 vdd.n2512 72.8958
R19464 vdd.n2978 vdd.n613 72.8958
R19465 vdd.n2984 vdd.n613 72.8958
R19466 vdd.n659 vdd.n613 72.8958
R19467 vdd.n2991 vdd.n613 72.8958
R19468 vdd.n656 vdd.n613 72.8958
R19469 vdd.n2998 vdd.n613 72.8958
R19470 vdd.n653 vdd.n613 72.8958
R19471 vdd.n3005 vdd.n613 72.8958
R19472 vdd.n650 vdd.n613 72.8958
R19473 vdd.n3013 vdd.n613 72.8958
R19474 vdd.n647 vdd.n613 72.8958
R19475 vdd.n3020 vdd.n613 72.8958
R19476 vdd.n644 vdd.n613 72.8958
R19477 vdd.n3027 vdd.n613 72.8958
R19478 vdd.n641 vdd.n613 72.8958
R19479 vdd.n3034 vdd.n613 72.8958
R19480 vdd.n3037 vdd.n613 72.8958
R19481 vdd.n2496 vdd.n807 72.8958
R19482 vdd.n2496 vdd.n806 72.8958
R19483 vdd.n2496 vdd.n805 72.8958
R19484 vdd.n2496 vdd.n804 72.8958
R19485 vdd.n2496 vdd.n803 72.8958
R19486 vdd.n2496 vdd.n802 72.8958
R19487 vdd.n2496 vdd.n801 72.8958
R19488 vdd.n2496 vdd.n800 72.8958
R19489 vdd.n2496 vdd.n799 72.8958
R19490 vdd.n2496 vdd.n798 72.8958
R19491 vdd.n2496 vdd.n797 72.8958
R19492 vdd.n2496 vdd.n796 72.8958
R19493 vdd.n2496 vdd.n795 72.8958
R19494 vdd.n2496 vdd.n794 72.8958
R19495 vdd.n2496 vdd.n793 72.8958
R19496 vdd.n2496 vdd.n792 72.8958
R19497 vdd.n2496 vdd.n791 72.8958
R19498 vdd.n2218 vdd.n986 72.8958
R19499 vdd.n2218 vdd.n987 72.8958
R19500 vdd.n2218 vdd.n988 72.8958
R19501 vdd.n2218 vdd.n989 72.8958
R19502 vdd.n2218 vdd.n990 72.8958
R19503 vdd.n2218 vdd.n991 72.8958
R19504 vdd.n2218 vdd.n992 72.8958
R19505 vdd.n2218 vdd.n993 72.8958
R19506 vdd.n2218 vdd.n994 72.8958
R19507 vdd.n2218 vdd.n995 72.8958
R19508 vdd.n2218 vdd.n996 72.8958
R19509 vdd.n2218 vdd.n997 72.8958
R19510 vdd.n2218 vdd.n998 72.8958
R19511 vdd.n2218 vdd.n999 72.8958
R19512 vdd.n2218 vdd.n1000 72.8958
R19513 vdd.n2218 vdd.n1001 72.8958
R19514 vdd.n2218 vdd.n1002 72.8958
R19515 vdd.n1441 vdd.n1437 66.2847
R19516 vdd.n1447 vdd.n1437 66.2847
R19517 vdd.n1450 vdd.n1437 66.2847
R19518 vdd.n1455 vdd.n1437 66.2847
R19519 vdd.n1458 vdd.n1437 66.2847
R19520 vdd.n1463 vdd.n1437 66.2847
R19521 vdd.n1466 vdd.n1437 66.2847
R19522 vdd.n1471 vdd.n1437 66.2847
R19523 vdd.n1474 vdd.n1437 66.2847
R19524 vdd.n1481 vdd.n1437 66.2847
R19525 vdd.n1484 vdd.n1437 66.2847
R19526 vdd.n1489 vdd.n1437 66.2847
R19527 vdd.n1492 vdd.n1437 66.2847
R19528 vdd.n1497 vdd.n1437 66.2847
R19529 vdd.n1500 vdd.n1437 66.2847
R19530 vdd.n1505 vdd.n1437 66.2847
R19531 vdd.n1508 vdd.n1437 66.2847
R19532 vdd.n1513 vdd.n1437 66.2847
R19533 vdd.n1516 vdd.n1437 66.2847
R19534 vdd.n1521 vdd.n1437 66.2847
R19535 vdd.n1600 vdd.n1437 66.2847
R19536 vdd.n1524 vdd.n1437 66.2847
R19537 vdd.n1530 vdd.n1437 66.2847
R19538 vdd.n1535 vdd.n1437 66.2847
R19539 vdd.n1538 vdd.n1437 66.2847
R19540 vdd.n1543 vdd.n1437 66.2847
R19541 vdd.n1546 vdd.n1437 66.2847
R19542 vdd.n1551 vdd.n1437 66.2847
R19543 vdd.n1554 vdd.n1437 66.2847
R19544 vdd.n1559 vdd.n1437 66.2847
R19545 vdd.n1562 vdd.n1437 66.2847
R19546 vdd.n1354 vdd.n969 66.2847
R19547 vdd.n1351 vdd.n969 66.2847
R19548 vdd.n1347 vdd.n969 66.2847
R19549 vdd.n2084 vdd.n969 66.2847
R19550 vdd.n1103 vdd.n969 66.2847
R19551 vdd.n2091 vdd.n969 66.2847
R19552 vdd.n1096 vdd.n969 66.2847
R19553 vdd.n2098 vdd.n969 66.2847
R19554 vdd.n1089 vdd.n969 66.2847
R19555 vdd.n2105 vdd.n969 66.2847
R19556 vdd.n1083 vdd.n969 66.2847
R19557 vdd.n1078 vdd.n969 66.2847
R19558 vdd.n2116 vdd.n969 66.2847
R19559 vdd.n1070 vdd.n969 66.2847
R19560 vdd.n2123 vdd.n969 66.2847
R19561 vdd.n1063 vdd.n969 66.2847
R19562 vdd.n2130 vdd.n969 66.2847
R19563 vdd.n1056 vdd.n969 66.2847
R19564 vdd.n2137 vdd.n969 66.2847
R19565 vdd.n1049 vdd.n969 66.2847
R19566 vdd.n2144 vdd.n969 66.2847
R19567 vdd.n1043 vdd.n969 66.2847
R19568 vdd.n1038 vdd.n969 66.2847
R19569 vdd.n2155 vdd.n969 66.2847
R19570 vdd.n1030 vdd.n969 66.2847
R19571 vdd.n2162 vdd.n969 66.2847
R19572 vdd.n1023 vdd.n969 66.2847
R19573 vdd.n2169 vdd.n969 66.2847
R19574 vdd.n1016 vdd.n969 66.2847
R19575 vdd.n2176 vdd.n969 66.2847
R19576 vdd.n2181 vdd.n969 66.2847
R19577 vdd.n1012 vdd.n969 66.2847
R19578 vdd.n3204 vdd.n516 66.2847
R19579 vdd.n520 vdd.n516 66.2847
R19580 vdd.n523 vdd.n516 66.2847
R19581 vdd.n3193 vdd.n516 66.2847
R19582 vdd.n3187 vdd.n516 66.2847
R19583 vdd.n3185 vdd.n516 66.2847
R19584 vdd.n3179 vdd.n516 66.2847
R19585 vdd.n3177 vdd.n516 66.2847
R19586 vdd.n3171 vdd.n516 66.2847
R19587 vdd.n3169 vdd.n516 66.2847
R19588 vdd.n3163 vdd.n516 66.2847
R19589 vdd.n3161 vdd.n516 66.2847
R19590 vdd.n3155 vdd.n516 66.2847
R19591 vdd.n3153 vdd.n516 66.2847
R19592 vdd.n3147 vdd.n516 66.2847
R19593 vdd.n3145 vdd.n516 66.2847
R19594 vdd.n3139 vdd.n516 66.2847
R19595 vdd.n3137 vdd.n516 66.2847
R19596 vdd.n3131 vdd.n516 66.2847
R19597 vdd.n3129 vdd.n516 66.2847
R19598 vdd.n584 vdd.n516 66.2847
R19599 vdd.n3120 vdd.n516 66.2847
R19600 vdd.n586 vdd.n516 66.2847
R19601 vdd.n3113 vdd.n516 66.2847
R19602 vdd.n3107 vdd.n516 66.2847
R19603 vdd.n3105 vdd.n516 66.2847
R19604 vdd.n3099 vdd.n516 66.2847
R19605 vdd.n3097 vdd.n516 66.2847
R19606 vdd.n3091 vdd.n516 66.2847
R19607 vdd.n607 vdd.n516 66.2847
R19608 vdd.n609 vdd.n516 66.2847
R19609 vdd.n3290 vdd.n351 66.2847
R19610 vdd.n3299 vdd.n351 66.2847
R19611 vdd.n461 vdd.n351 66.2847
R19612 vdd.n3306 vdd.n351 66.2847
R19613 vdd.n454 vdd.n351 66.2847
R19614 vdd.n3313 vdd.n351 66.2847
R19615 vdd.n447 vdd.n351 66.2847
R19616 vdd.n3320 vdd.n351 66.2847
R19617 vdd.n440 vdd.n351 66.2847
R19618 vdd.n3327 vdd.n351 66.2847
R19619 vdd.n434 vdd.n351 66.2847
R19620 vdd.n429 vdd.n351 66.2847
R19621 vdd.n3338 vdd.n351 66.2847
R19622 vdd.n421 vdd.n351 66.2847
R19623 vdd.n3345 vdd.n351 66.2847
R19624 vdd.n414 vdd.n351 66.2847
R19625 vdd.n3352 vdd.n351 66.2847
R19626 vdd.n407 vdd.n351 66.2847
R19627 vdd.n3359 vdd.n351 66.2847
R19628 vdd.n400 vdd.n351 66.2847
R19629 vdd.n3366 vdd.n351 66.2847
R19630 vdd.n394 vdd.n351 66.2847
R19631 vdd.n389 vdd.n351 66.2847
R19632 vdd.n3377 vdd.n351 66.2847
R19633 vdd.n381 vdd.n351 66.2847
R19634 vdd.n3384 vdd.n351 66.2847
R19635 vdd.n374 vdd.n351 66.2847
R19636 vdd.n3391 vdd.n351 66.2847
R19637 vdd.n367 vdd.n351 66.2847
R19638 vdd.n3398 vdd.n351 66.2847
R19639 vdd.n3401 vdd.n351 66.2847
R19640 vdd.n355 vdd.n351 66.2847
R19641 vdd.n356 vdd.n355 52.4337
R19642 vdd.n3401 vdd.n3400 52.4337
R19643 vdd.n3398 vdd.n3397 52.4337
R19644 vdd.n3393 vdd.n367 52.4337
R19645 vdd.n3391 vdd.n3390 52.4337
R19646 vdd.n3386 vdd.n374 52.4337
R19647 vdd.n3384 vdd.n3383 52.4337
R19648 vdd.n3379 vdd.n381 52.4337
R19649 vdd.n3377 vdd.n3376 52.4337
R19650 vdd.n390 vdd.n389 52.4337
R19651 vdd.n3368 vdd.n394 52.4337
R19652 vdd.n3366 vdd.n3365 52.4337
R19653 vdd.n3361 vdd.n400 52.4337
R19654 vdd.n3359 vdd.n3358 52.4337
R19655 vdd.n3354 vdd.n407 52.4337
R19656 vdd.n3352 vdd.n3351 52.4337
R19657 vdd.n3347 vdd.n414 52.4337
R19658 vdd.n3345 vdd.n3344 52.4337
R19659 vdd.n3340 vdd.n421 52.4337
R19660 vdd.n3338 vdd.n3337 52.4337
R19661 vdd.n430 vdd.n429 52.4337
R19662 vdd.n3329 vdd.n434 52.4337
R19663 vdd.n3327 vdd.n3326 52.4337
R19664 vdd.n3322 vdd.n440 52.4337
R19665 vdd.n3320 vdd.n3319 52.4337
R19666 vdd.n3315 vdd.n447 52.4337
R19667 vdd.n3313 vdd.n3312 52.4337
R19668 vdd.n3308 vdd.n454 52.4337
R19669 vdd.n3306 vdd.n3305 52.4337
R19670 vdd.n3301 vdd.n461 52.4337
R19671 vdd.n3299 vdd.n3298 52.4337
R19672 vdd.n3291 vdd.n3290 52.4337
R19673 vdd.n3204 vdd.n517 52.4337
R19674 vdd.n3202 vdd.n520 52.4337
R19675 vdd.n3198 vdd.n523 52.4337
R19676 vdd.n3194 vdd.n3193 52.4337
R19677 vdd.n3187 vdd.n526 52.4337
R19678 vdd.n3186 vdd.n3185 52.4337
R19679 vdd.n3179 vdd.n532 52.4337
R19680 vdd.n3178 vdd.n3177 52.4337
R19681 vdd.n3171 vdd.n538 52.4337
R19682 vdd.n3170 vdd.n3169 52.4337
R19683 vdd.n3163 vdd.n546 52.4337
R19684 vdd.n3162 vdd.n3161 52.4337
R19685 vdd.n3155 vdd.n552 52.4337
R19686 vdd.n3154 vdd.n3153 52.4337
R19687 vdd.n3147 vdd.n558 52.4337
R19688 vdd.n3146 vdd.n3145 52.4337
R19689 vdd.n3139 vdd.n564 52.4337
R19690 vdd.n3138 vdd.n3137 52.4337
R19691 vdd.n3131 vdd.n570 52.4337
R19692 vdd.n3130 vdd.n3129 52.4337
R19693 vdd.n584 vdd.n576 52.4337
R19694 vdd.n3121 vdd.n3120 52.4337
R19695 vdd.n3118 vdd.n586 52.4337
R19696 vdd.n3114 vdd.n3113 52.4337
R19697 vdd.n3107 vdd.n590 52.4337
R19698 vdd.n3106 vdd.n3105 52.4337
R19699 vdd.n3099 vdd.n596 52.4337
R19700 vdd.n3098 vdd.n3097 52.4337
R19701 vdd.n3091 vdd.n602 52.4337
R19702 vdd.n3090 vdd.n607 52.4337
R19703 vdd.n3086 vdd.n609 52.4337
R19704 vdd.n2183 vdd.n1012 52.4337
R19705 vdd.n2181 vdd.n2180 52.4337
R19706 vdd.n2176 vdd.n2175 52.4337
R19707 vdd.n2171 vdd.n1016 52.4337
R19708 vdd.n2169 vdd.n2168 52.4337
R19709 vdd.n2164 vdd.n1023 52.4337
R19710 vdd.n2162 vdd.n2161 52.4337
R19711 vdd.n2157 vdd.n1030 52.4337
R19712 vdd.n2155 vdd.n2154 52.4337
R19713 vdd.n1039 vdd.n1038 52.4337
R19714 vdd.n2146 vdd.n1043 52.4337
R19715 vdd.n2144 vdd.n2143 52.4337
R19716 vdd.n2139 vdd.n1049 52.4337
R19717 vdd.n2137 vdd.n2136 52.4337
R19718 vdd.n2132 vdd.n1056 52.4337
R19719 vdd.n2130 vdd.n2129 52.4337
R19720 vdd.n2125 vdd.n1063 52.4337
R19721 vdd.n2123 vdd.n2122 52.4337
R19722 vdd.n2118 vdd.n1070 52.4337
R19723 vdd.n2116 vdd.n2115 52.4337
R19724 vdd.n1079 vdd.n1078 52.4337
R19725 vdd.n2107 vdd.n1083 52.4337
R19726 vdd.n2105 vdd.n2104 52.4337
R19727 vdd.n2100 vdd.n1089 52.4337
R19728 vdd.n2098 vdd.n2097 52.4337
R19729 vdd.n2093 vdd.n1096 52.4337
R19730 vdd.n2091 vdd.n2090 52.4337
R19731 vdd.n2086 vdd.n1103 52.4337
R19732 vdd.n2084 vdd.n2083 52.4337
R19733 vdd.n1348 vdd.n1347 52.4337
R19734 vdd.n1352 vdd.n1351 52.4337
R19735 vdd.n2072 vdd.n1354 52.4337
R19736 vdd.n1441 vdd.n1439 52.4337
R19737 vdd.n1447 vdd.n1446 52.4337
R19738 vdd.n1450 vdd.n1449 52.4337
R19739 vdd.n1455 vdd.n1454 52.4337
R19740 vdd.n1458 vdd.n1457 52.4337
R19741 vdd.n1463 vdd.n1462 52.4337
R19742 vdd.n1466 vdd.n1465 52.4337
R19743 vdd.n1471 vdd.n1470 52.4337
R19744 vdd.n1474 vdd.n1473 52.4337
R19745 vdd.n1481 vdd.n1480 52.4337
R19746 vdd.n1484 vdd.n1483 52.4337
R19747 vdd.n1489 vdd.n1488 52.4337
R19748 vdd.n1492 vdd.n1491 52.4337
R19749 vdd.n1497 vdd.n1496 52.4337
R19750 vdd.n1500 vdd.n1499 52.4337
R19751 vdd.n1505 vdd.n1504 52.4337
R19752 vdd.n1508 vdd.n1507 52.4337
R19753 vdd.n1513 vdd.n1512 52.4337
R19754 vdd.n1516 vdd.n1515 52.4337
R19755 vdd.n1521 vdd.n1520 52.4337
R19756 vdd.n1601 vdd.n1600 52.4337
R19757 vdd.n1598 vdd.n1524 52.4337
R19758 vdd.n1530 vdd.n1529 52.4337
R19759 vdd.n1535 vdd.n1532 52.4337
R19760 vdd.n1538 vdd.n1537 52.4337
R19761 vdd.n1543 vdd.n1540 52.4337
R19762 vdd.n1546 vdd.n1545 52.4337
R19763 vdd.n1551 vdd.n1548 52.4337
R19764 vdd.n1554 vdd.n1553 52.4337
R19765 vdd.n1559 vdd.n1556 52.4337
R19766 vdd.n1562 vdd.n1561 52.4337
R19767 vdd.n1442 vdd.n1441 52.4337
R19768 vdd.n1448 vdd.n1447 52.4337
R19769 vdd.n1451 vdd.n1450 52.4337
R19770 vdd.n1456 vdd.n1455 52.4337
R19771 vdd.n1459 vdd.n1458 52.4337
R19772 vdd.n1464 vdd.n1463 52.4337
R19773 vdd.n1467 vdd.n1466 52.4337
R19774 vdd.n1472 vdd.n1471 52.4337
R19775 vdd.n1475 vdd.n1474 52.4337
R19776 vdd.n1482 vdd.n1481 52.4337
R19777 vdd.n1485 vdd.n1484 52.4337
R19778 vdd.n1490 vdd.n1489 52.4337
R19779 vdd.n1493 vdd.n1492 52.4337
R19780 vdd.n1498 vdd.n1497 52.4337
R19781 vdd.n1501 vdd.n1500 52.4337
R19782 vdd.n1506 vdd.n1505 52.4337
R19783 vdd.n1509 vdd.n1508 52.4337
R19784 vdd.n1514 vdd.n1513 52.4337
R19785 vdd.n1517 vdd.n1516 52.4337
R19786 vdd.n1522 vdd.n1521 52.4337
R19787 vdd.n1600 vdd.n1599 52.4337
R19788 vdd.n1528 vdd.n1524 52.4337
R19789 vdd.n1531 vdd.n1530 52.4337
R19790 vdd.n1536 vdd.n1535 52.4337
R19791 vdd.n1539 vdd.n1538 52.4337
R19792 vdd.n1544 vdd.n1543 52.4337
R19793 vdd.n1547 vdd.n1546 52.4337
R19794 vdd.n1552 vdd.n1551 52.4337
R19795 vdd.n1555 vdd.n1554 52.4337
R19796 vdd.n1560 vdd.n1559 52.4337
R19797 vdd.n1563 vdd.n1562 52.4337
R19798 vdd.n1354 vdd.n1353 52.4337
R19799 vdd.n1351 vdd.n1350 52.4337
R19800 vdd.n1347 vdd.n1104 52.4337
R19801 vdd.n2085 vdd.n2084 52.4337
R19802 vdd.n1103 vdd.n1097 52.4337
R19803 vdd.n2092 vdd.n2091 52.4337
R19804 vdd.n1096 vdd.n1090 52.4337
R19805 vdd.n2099 vdd.n2098 52.4337
R19806 vdd.n1089 vdd.n1084 52.4337
R19807 vdd.n2106 vdd.n2105 52.4337
R19808 vdd.n1083 vdd.n1082 52.4337
R19809 vdd.n1078 vdd.n1071 52.4337
R19810 vdd.n2117 vdd.n2116 52.4337
R19811 vdd.n1070 vdd.n1064 52.4337
R19812 vdd.n2124 vdd.n2123 52.4337
R19813 vdd.n1063 vdd.n1057 52.4337
R19814 vdd.n2131 vdd.n2130 52.4337
R19815 vdd.n1056 vdd.n1050 52.4337
R19816 vdd.n2138 vdd.n2137 52.4337
R19817 vdd.n1049 vdd.n1044 52.4337
R19818 vdd.n2145 vdd.n2144 52.4337
R19819 vdd.n1043 vdd.n1042 52.4337
R19820 vdd.n1038 vdd.n1031 52.4337
R19821 vdd.n2156 vdd.n2155 52.4337
R19822 vdd.n1030 vdd.n1024 52.4337
R19823 vdd.n2163 vdd.n2162 52.4337
R19824 vdd.n1023 vdd.n1017 52.4337
R19825 vdd.n2170 vdd.n2169 52.4337
R19826 vdd.n1016 vdd.n1013 52.4337
R19827 vdd.n2177 vdd.n2176 52.4337
R19828 vdd.n2182 vdd.n2181 52.4337
R19829 vdd.n1358 vdd.n1012 52.4337
R19830 vdd.n3205 vdd.n3204 52.4337
R19831 vdd.n3199 vdd.n520 52.4337
R19832 vdd.n3195 vdd.n523 52.4337
R19833 vdd.n3193 vdd.n3192 52.4337
R19834 vdd.n3188 vdd.n3187 52.4337
R19835 vdd.n3185 vdd.n3184 52.4337
R19836 vdd.n3180 vdd.n3179 52.4337
R19837 vdd.n3177 vdd.n3176 52.4337
R19838 vdd.n3172 vdd.n3171 52.4337
R19839 vdd.n3169 vdd.n3168 52.4337
R19840 vdd.n3164 vdd.n3163 52.4337
R19841 vdd.n3161 vdd.n3160 52.4337
R19842 vdd.n3156 vdd.n3155 52.4337
R19843 vdd.n3153 vdd.n3152 52.4337
R19844 vdd.n3148 vdd.n3147 52.4337
R19845 vdd.n3145 vdd.n3144 52.4337
R19846 vdd.n3140 vdd.n3139 52.4337
R19847 vdd.n3137 vdd.n3136 52.4337
R19848 vdd.n3132 vdd.n3131 52.4337
R19849 vdd.n3129 vdd.n3128 52.4337
R19850 vdd.n585 vdd.n584 52.4337
R19851 vdd.n3120 vdd.n3119 52.4337
R19852 vdd.n3115 vdd.n586 52.4337
R19853 vdd.n3113 vdd.n3112 52.4337
R19854 vdd.n3108 vdd.n3107 52.4337
R19855 vdd.n3105 vdd.n3104 52.4337
R19856 vdd.n3100 vdd.n3099 52.4337
R19857 vdd.n3097 vdd.n3096 52.4337
R19858 vdd.n3092 vdd.n3091 52.4337
R19859 vdd.n3087 vdd.n607 52.4337
R19860 vdd.n3083 vdd.n609 52.4337
R19861 vdd.n3290 vdd.n462 52.4337
R19862 vdd.n3300 vdd.n3299 52.4337
R19863 vdd.n461 vdd.n455 52.4337
R19864 vdd.n3307 vdd.n3306 52.4337
R19865 vdd.n454 vdd.n448 52.4337
R19866 vdd.n3314 vdd.n3313 52.4337
R19867 vdd.n447 vdd.n441 52.4337
R19868 vdd.n3321 vdd.n3320 52.4337
R19869 vdd.n440 vdd.n435 52.4337
R19870 vdd.n3328 vdd.n3327 52.4337
R19871 vdd.n434 vdd.n433 52.4337
R19872 vdd.n429 vdd.n422 52.4337
R19873 vdd.n3339 vdd.n3338 52.4337
R19874 vdd.n421 vdd.n415 52.4337
R19875 vdd.n3346 vdd.n3345 52.4337
R19876 vdd.n414 vdd.n408 52.4337
R19877 vdd.n3353 vdd.n3352 52.4337
R19878 vdd.n407 vdd.n401 52.4337
R19879 vdd.n3360 vdd.n3359 52.4337
R19880 vdd.n400 vdd.n395 52.4337
R19881 vdd.n3367 vdd.n3366 52.4337
R19882 vdd.n394 vdd.n393 52.4337
R19883 vdd.n389 vdd.n382 52.4337
R19884 vdd.n3378 vdd.n3377 52.4337
R19885 vdd.n381 vdd.n375 52.4337
R19886 vdd.n3385 vdd.n3384 52.4337
R19887 vdd.n374 vdd.n368 52.4337
R19888 vdd.n3392 vdd.n3391 52.4337
R19889 vdd.n367 vdd.n360 52.4337
R19890 vdd.n3399 vdd.n3398 52.4337
R19891 vdd.n3402 vdd.n3401 52.4337
R19892 vdd.n355 vdd.n352 52.4337
R19893 vdd.t164 vdd.t188 51.4683
R19894 vdd.n258 vdd.n256 42.0461
R19895 vdd.n164 vdd.n162 42.0461
R19896 vdd.n71 vdd.n69 42.0461
R19897 vdd.n1959 vdd.n1957 42.0461
R19898 vdd.n1865 vdd.n1863 42.0461
R19899 vdd.n1772 vdd.n1770 42.0461
R19900 vdd.n308 vdd.n307 41.6884
R19901 vdd.n214 vdd.n213 41.6884
R19902 vdd.n121 vdd.n120 41.6884
R19903 vdd.n2009 vdd.n2008 41.6884
R19904 vdd.n1915 vdd.n1914 41.6884
R19905 vdd.n1822 vdd.n1821 41.6884
R19906 vdd.n1567 vdd.n1566 41.1157
R19907 vdd.n1604 vdd.n1603 41.1157
R19908 vdd.n1478 vdd.n1477 41.1157
R19909 vdd.n3295 vdd.n3294 41.1157
R19910 vdd.n3334 vdd.n428 41.1157
R19911 vdd.n3373 vdd.n388 41.1157
R19912 vdd.n3037 vdd.n3036 39.2114
R19913 vdd.n3034 vdd.n3033 39.2114
R19914 vdd.n3029 vdd.n641 39.2114
R19915 vdd.n3027 vdd.n3026 39.2114
R19916 vdd.n3022 vdd.n644 39.2114
R19917 vdd.n3020 vdd.n3019 39.2114
R19918 vdd.n3015 vdd.n647 39.2114
R19919 vdd.n3013 vdd.n3012 39.2114
R19920 vdd.n3007 vdd.n650 39.2114
R19921 vdd.n3005 vdd.n3004 39.2114
R19922 vdd.n3000 vdd.n653 39.2114
R19923 vdd.n2998 vdd.n2997 39.2114
R19924 vdd.n2993 vdd.n656 39.2114
R19925 vdd.n2991 vdd.n2990 39.2114
R19926 vdd.n2986 vdd.n659 39.2114
R19927 vdd.n2984 vdd.n2983 39.2114
R19928 vdd.n2979 vdd.n2978 39.2114
R19929 vdd.n2802 vdd.n2801 39.2114
R19930 vdd.n2531 vdd.n2497 39.2114
R19931 vdd.n2794 vdd.n2498 39.2114
R19932 vdd.n2790 vdd.n2499 39.2114
R19933 vdd.n2786 vdd.n2500 39.2114
R19934 vdd.n2782 vdd.n2501 39.2114
R19935 vdd.n2778 vdd.n2502 39.2114
R19936 vdd.n2774 vdd.n2503 39.2114
R19937 vdd.n2770 vdd.n2504 39.2114
R19938 vdd.n2766 vdd.n2505 39.2114
R19939 vdd.n2762 vdd.n2506 39.2114
R19940 vdd.n2758 vdd.n2507 39.2114
R19941 vdd.n2754 vdd.n2508 39.2114
R19942 vdd.n2750 vdd.n2509 39.2114
R19943 vdd.n2746 vdd.n2510 39.2114
R19944 vdd.n2742 vdd.n2511 39.2114
R19945 vdd.n2737 vdd.n2512 39.2114
R19946 vdd.n2491 vdd.n825 39.2114
R19947 vdd.n2487 vdd.n824 39.2114
R19948 vdd.n2483 vdd.n823 39.2114
R19949 vdd.n2479 vdd.n822 39.2114
R19950 vdd.n2475 vdd.n821 39.2114
R19951 vdd.n2471 vdd.n820 39.2114
R19952 vdd.n2467 vdd.n819 39.2114
R19953 vdd.n2463 vdd.n818 39.2114
R19954 vdd.n2459 vdd.n817 39.2114
R19955 vdd.n2455 vdd.n816 39.2114
R19956 vdd.n2451 vdd.n815 39.2114
R19957 vdd.n2447 vdd.n814 39.2114
R19958 vdd.n2443 vdd.n813 39.2114
R19959 vdd.n2439 vdd.n812 39.2114
R19960 vdd.n2435 vdd.n811 39.2114
R19961 vdd.n2430 vdd.n810 39.2114
R19962 vdd.n2426 vdd.n809 39.2114
R19963 vdd.n2220 vdd.n2219 39.2114
R19964 vdd.n1004 vdd.n970 39.2114
R19965 vdd.n2212 vdd.n971 39.2114
R19966 vdd.n2208 vdd.n972 39.2114
R19967 vdd.n2204 vdd.n973 39.2114
R19968 vdd.n2200 vdd.n974 39.2114
R19969 vdd.n2196 vdd.n975 39.2114
R19970 vdd.n2192 vdd.n976 39.2114
R19971 vdd.n2188 vdd.n977 39.2114
R19972 vdd.n1150 vdd.n978 39.2114
R19973 vdd.n1154 vdd.n979 39.2114
R19974 vdd.n1158 vdd.n980 39.2114
R19975 vdd.n1162 vdd.n981 39.2114
R19976 vdd.n1166 vdd.n982 39.2114
R19977 vdd.n1170 vdd.n983 39.2114
R19978 vdd.n1174 vdd.n984 39.2114
R19979 vdd.n1179 vdd.n985 39.2114
R19980 vdd.n2956 vdd.n2955 39.2114
R19981 vdd.n2951 vdd.n2923 39.2114
R19982 vdd.n2949 vdd.n2948 39.2114
R19983 vdd.n2944 vdd.n2926 39.2114
R19984 vdd.n2942 vdd.n2941 39.2114
R19985 vdd.n2937 vdd.n2929 39.2114
R19986 vdd.n2935 vdd.n2934 39.2114
R19987 vdd.n2930 vdd.n612 39.2114
R19988 vdd.n3074 vdd.n3073 39.2114
R19989 vdd.n3071 vdd.n3070 39.2114
R19990 vdd.n3066 vdd.n617 39.2114
R19991 vdd.n3064 vdd.n3063 39.2114
R19992 vdd.n3059 vdd.n620 39.2114
R19993 vdd.n3057 vdd.n3056 39.2114
R19994 vdd.n3052 vdd.n623 39.2114
R19995 vdd.n3050 vdd.n3049 39.2114
R19996 vdd.n3045 vdd.n629 39.2114
R19997 vdd.n2538 vdd.n2513 39.2114
R19998 vdd.n2542 vdd.n2514 39.2114
R19999 vdd.n2546 vdd.n2515 39.2114
R20000 vdd.n2550 vdd.n2516 39.2114
R20001 vdd.n2554 vdd.n2517 39.2114
R20002 vdd.n2558 vdd.n2518 39.2114
R20003 vdd.n2562 vdd.n2519 39.2114
R20004 vdd.n2566 vdd.n2520 39.2114
R20005 vdd.n2570 vdd.n2521 39.2114
R20006 vdd.n2574 vdd.n2522 39.2114
R20007 vdd.n2578 vdd.n2523 39.2114
R20008 vdd.n2582 vdd.n2524 39.2114
R20009 vdd.n2586 vdd.n2525 39.2114
R20010 vdd.n2590 vdd.n2526 39.2114
R20011 vdd.n2594 vdd.n2527 39.2114
R20012 vdd.n2598 vdd.n2528 39.2114
R20013 vdd.n2602 vdd.n2529 39.2114
R20014 vdd.n2541 vdd.n2513 39.2114
R20015 vdd.n2545 vdd.n2514 39.2114
R20016 vdd.n2549 vdd.n2515 39.2114
R20017 vdd.n2553 vdd.n2516 39.2114
R20018 vdd.n2557 vdd.n2517 39.2114
R20019 vdd.n2561 vdd.n2518 39.2114
R20020 vdd.n2565 vdd.n2519 39.2114
R20021 vdd.n2569 vdd.n2520 39.2114
R20022 vdd.n2573 vdd.n2521 39.2114
R20023 vdd.n2577 vdd.n2522 39.2114
R20024 vdd.n2581 vdd.n2523 39.2114
R20025 vdd.n2585 vdd.n2524 39.2114
R20026 vdd.n2589 vdd.n2525 39.2114
R20027 vdd.n2593 vdd.n2526 39.2114
R20028 vdd.n2597 vdd.n2527 39.2114
R20029 vdd.n2601 vdd.n2528 39.2114
R20030 vdd.n2604 vdd.n2529 39.2114
R20031 vdd.n629 vdd.n624 39.2114
R20032 vdd.n3051 vdd.n3050 39.2114
R20033 vdd.n623 vdd.n621 39.2114
R20034 vdd.n3058 vdd.n3057 39.2114
R20035 vdd.n620 vdd.n618 39.2114
R20036 vdd.n3065 vdd.n3064 39.2114
R20037 vdd.n617 vdd.n615 39.2114
R20038 vdd.n3072 vdd.n3071 39.2114
R20039 vdd.n3075 vdd.n3074 39.2114
R20040 vdd.n2931 vdd.n2930 39.2114
R20041 vdd.n2936 vdd.n2935 39.2114
R20042 vdd.n2929 vdd.n2927 39.2114
R20043 vdd.n2943 vdd.n2942 39.2114
R20044 vdd.n2926 vdd.n2924 39.2114
R20045 vdd.n2950 vdd.n2949 39.2114
R20046 vdd.n2923 vdd.n2921 39.2114
R20047 vdd.n2957 vdd.n2956 39.2114
R20048 vdd.n2219 vdd.n968 39.2114
R20049 vdd.n2213 vdd.n970 39.2114
R20050 vdd.n2209 vdd.n971 39.2114
R20051 vdd.n2205 vdd.n972 39.2114
R20052 vdd.n2201 vdd.n973 39.2114
R20053 vdd.n2197 vdd.n974 39.2114
R20054 vdd.n2193 vdd.n975 39.2114
R20055 vdd.n2189 vdd.n976 39.2114
R20056 vdd.n1149 vdd.n977 39.2114
R20057 vdd.n1153 vdd.n978 39.2114
R20058 vdd.n1157 vdd.n979 39.2114
R20059 vdd.n1161 vdd.n980 39.2114
R20060 vdd.n1165 vdd.n981 39.2114
R20061 vdd.n1169 vdd.n982 39.2114
R20062 vdd.n1173 vdd.n983 39.2114
R20063 vdd.n1178 vdd.n984 39.2114
R20064 vdd.n1182 vdd.n985 39.2114
R20065 vdd.n2429 vdd.n809 39.2114
R20066 vdd.n2434 vdd.n810 39.2114
R20067 vdd.n2438 vdd.n811 39.2114
R20068 vdd.n2442 vdd.n812 39.2114
R20069 vdd.n2446 vdd.n813 39.2114
R20070 vdd.n2450 vdd.n814 39.2114
R20071 vdd.n2454 vdd.n815 39.2114
R20072 vdd.n2458 vdd.n816 39.2114
R20073 vdd.n2462 vdd.n817 39.2114
R20074 vdd.n2466 vdd.n818 39.2114
R20075 vdd.n2470 vdd.n819 39.2114
R20076 vdd.n2474 vdd.n820 39.2114
R20077 vdd.n2478 vdd.n821 39.2114
R20078 vdd.n2482 vdd.n822 39.2114
R20079 vdd.n2486 vdd.n823 39.2114
R20080 vdd.n2490 vdd.n824 39.2114
R20081 vdd.n827 vdd.n825 39.2114
R20082 vdd.n2801 vdd.n790 39.2114
R20083 vdd.n2795 vdd.n2497 39.2114
R20084 vdd.n2791 vdd.n2498 39.2114
R20085 vdd.n2787 vdd.n2499 39.2114
R20086 vdd.n2783 vdd.n2500 39.2114
R20087 vdd.n2779 vdd.n2501 39.2114
R20088 vdd.n2775 vdd.n2502 39.2114
R20089 vdd.n2771 vdd.n2503 39.2114
R20090 vdd.n2767 vdd.n2504 39.2114
R20091 vdd.n2763 vdd.n2505 39.2114
R20092 vdd.n2759 vdd.n2506 39.2114
R20093 vdd.n2755 vdd.n2507 39.2114
R20094 vdd.n2751 vdd.n2508 39.2114
R20095 vdd.n2747 vdd.n2509 39.2114
R20096 vdd.n2743 vdd.n2510 39.2114
R20097 vdd.n2738 vdd.n2511 39.2114
R20098 vdd.n2734 vdd.n2512 39.2114
R20099 vdd.n2978 vdd.n660 39.2114
R20100 vdd.n2985 vdd.n2984 39.2114
R20101 vdd.n659 vdd.n657 39.2114
R20102 vdd.n2992 vdd.n2991 39.2114
R20103 vdd.n656 vdd.n654 39.2114
R20104 vdd.n2999 vdd.n2998 39.2114
R20105 vdd.n653 vdd.n651 39.2114
R20106 vdd.n3006 vdd.n3005 39.2114
R20107 vdd.n650 vdd.n648 39.2114
R20108 vdd.n3014 vdd.n3013 39.2114
R20109 vdd.n647 vdd.n645 39.2114
R20110 vdd.n3021 vdd.n3020 39.2114
R20111 vdd.n644 vdd.n642 39.2114
R20112 vdd.n3028 vdd.n3027 39.2114
R20113 vdd.n641 vdd.n639 39.2114
R20114 vdd.n3035 vdd.n3034 39.2114
R20115 vdd.n3038 vdd.n3037 39.2114
R20116 vdd.n836 vdd.n791 39.2114
R20117 vdd.n2418 vdd.n792 39.2114
R20118 vdd.n2414 vdd.n793 39.2114
R20119 vdd.n2410 vdd.n794 39.2114
R20120 vdd.n2406 vdd.n795 39.2114
R20121 vdd.n2402 vdd.n796 39.2114
R20122 vdd.n2398 vdd.n797 39.2114
R20123 vdd.n2394 vdd.n798 39.2114
R20124 vdd.n2390 vdd.n799 39.2114
R20125 vdd.n2386 vdd.n800 39.2114
R20126 vdd.n2382 vdd.n801 39.2114
R20127 vdd.n2378 vdd.n802 39.2114
R20128 vdd.n2374 vdd.n803 39.2114
R20129 vdd.n2370 vdd.n804 39.2114
R20130 vdd.n2366 vdd.n805 39.2114
R20131 vdd.n2362 vdd.n806 39.2114
R20132 vdd.n2358 vdd.n807 39.2114
R20133 vdd.n1108 vdd.n986 39.2114
R20134 vdd.n1112 vdd.n987 39.2114
R20135 vdd.n1116 vdd.n988 39.2114
R20136 vdd.n1120 vdd.n989 39.2114
R20137 vdd.n1124 vdd.n990 39.2114
R20138 vdd.n1128 vdd.n991 39.2114
R20139 vdd.n1132 vdd.n992 39.2114
R20140 vdd.n1136 vdd.n993 39.2114
R20141 vdd.n1140 vdd.n994 39.2114
R20142 vdd.n1341 vdd.n995 39.2114
R20143 vdd.n1338 vdd.n996 39.2114
R20144 vdd.n1334 vdd.n997 39.2114
R20145 vdd.n1330 vdd.n998 39.2114
R20146 vdd.n1326 vdd.n999 39.2114
R20147 vdd.n1322 vdd.n1000 39.2114
R20148 vdd.n1318 vdd.n1001 39.2114
R20149 vdd.n1314 vdd.n1002 39.2114
R20150 vdd.n2355 vdd.n807 39.2114
R20151 vdd.n2359 vdd.n806 39.2114
R20152 vdd.n2363 vdd.n805 39.2114
R20153 vdd.n2367 vdd.n804 39.2114
R20154 vdd.n2371 vdd.n803 39.2114
R20155 vdd.n2375 vdd.n802 39.2114
R20156 vdd.n2379 vdd.n801 39.2114
R20157 vdd.n2383 vdd.n800 39.2114
R20158 vdd.n2387 vdd.n799 39.2114
R20159 vdd.n2391 vdd.n798 39.2114
R20160 vdd.n2395 vdd.n797 39.2114
R20161 vdd.n2399 vdd.n796 39.2114
R20162 vdd.n2403 vdd.n795 39.2114
R20163 vdd.n2407 vdd.n794 39.2114
R20164 vdd.n2411 vdd.n793 39.2114
R20165 vdd.n2415 vdd.n792 39.2114
R20166 vdd.n2419 vdd.n791 39.2114
R20167 vdd.n1111 vdd.n986 39.2114
R20168 vdd.n1115 vdd.n987 39.2114
R20169 vdd.n1119 vdd.n988 39.2114
R20170 vdd.n1123 vdd.n989 39.2114
R20171 vdd.n1127 vdd.n990 39.2114
R20172 vdd.n1131 vdd.n991 39.2114
R20173 vdd.n1135 vdd.n992 39.2114
R20174 vdd.n1139 vdd.n993 39.2114
R20175 vdd.n1142 vdd.n994 39.2114
R20176 vdd.n1339 vdd.n995 39.2114
R20177 vdd.n1335 vdd.n996 39.2114
R20178 vdd.n1331 vdd.n997 39.2114
R20179 vdd.n1327 vdd.n998 39.2114
R20180 vdd.n1323 vdd.n999 39.2114
R20181 vdd.n1319 vdd.n1000 39.2114
R20182 vdd.n1315 vdd.n1001 39.2114
R20183 vdd.n1311 vdd.n1002 39.2114
R20184 vdd.n2076 vdd.n2075 37.2369
R20185 vdd.n2112 vdd.n1077 37.2369
R20186 vdd.n2151 vdd.n1037 37.2369
R20187 vdd.n3126 vdd.n581 37.2369
R20188 vdd.n545 vdd.n544 37.2369
R20189 vdd.n3082 vdd.n3081 37.2369
R20190 vdd.n1145 vdd.n1144 30.449
R20191 vdd.n840 vdd.n839 30.449
R20192 vdd.n1176 vdd.n1148 30.449
R20193 vdd.n2432 vdd.n830 30.449
R20194 vdd.n2537 vdd.n2536 30.449
R20195 vdd.n663 vdd.n662 30.449
R20196 vdd.n2740 vdd.n2533 30.449
R20197 vdd.n627 vdd.n626 30.449
R20198 vdd.n2222 vdd.n2221 29.8151
R20199 vdd.n2494 vdd.n828 29.8151
R20200 vdd.n2427 vdd.n831 29.8151
R20201 vdd.n1184 vdd.n1181 29.8151
R20202 vdd.n2735 vdd.n2732 29.8151
R20203 vdd.n2980 vdd.n2977 29.8151
R20204 vdd.n2804 vdd.n2803 29.8151
R20205 vdd.n3041 vdd.n3040 29.8151
R20206 vdd.n2960 vdd.n2959 29.8151
R20207 vdd.n3046 vdd.n628 29.8151
R20208 vdd.n2608 vdd.n2606 29.8151
R20209 vdd.n2539 vdd.n783 29.8151
R20210 vdd.n1109 vdd.n960 29.8151
R20211 vdd.n2422 vdd.n2421 29.8151
R20212 vdd.n2354 vdd.n2353 29.8151
R20213 vdd.n1310 vdd.n1309 29.8151
R20214 vdd.n1670 vdd.n1437 20.633
R20215 vdd.n2070 vdd.n969 20.633
R20216 vdd.n3212 vdd.n516 20.633
R20217 vdd.n3410 vdd.n351 20.633
R20218 vdd.n1672 vdd.n1434 19.3944
R20219 vdd.n1676 vdd.n1434 19.3944
R20220 vdd.n1676 vdd.n1425 19.3944
R20221 vdd.n1688 vdd.n1425 19.3944
R20222 vdd.n1688 vdd.n1423 19.3944
R20223 vdd.n1692 vdd.n1423 19.3944
R20224 vdd.n1692 vdd.n1412 19.3944
R20225 vdd.n1704 vdd.n1412 19.3944
R20226 vdd.n1704 vdd.n1410 19.3944
R20227 vdd.n1708 vdd.n1410 19.3944
R20228 vdd.n1708 vdd.n1401 19.3944
R20229 vdd.n1721 vdd.n1401 19.3944
R20230 vdd.n1721 vdd.n1399 19.3944
R20231 vdd.n1725 vdd.n1399 19.3944
R20232 vdd.n1725 vdd.n1390 19.3944
R20233 vdd.n2019 vdd.n1390 19.3944
R20234 vdd.n2019 vdd.n1388 19.3944
R20235 vdd.n2023 vdd.n1388 19.3944
R20236 vdd.n2023 vdd.n1378 19.3944
R20237 vdd.n2036 vdd.n1378 19.3944
R20238 vdd.n2036 vdd.n1376 19.3944
R20239 vdd.n2040 vdd.n1376 19.3944
R20240 vdd.n2040 vdd.n1368 19.3944
R20241 vdd.n2053 vdd.n1368 19.3944
R20242 vdd.n2053 vdd.n1365 19.3944
R20243 vdd.n2059 vdd.n1365 19.3944
R20244 vdd.n2059 vdd.n1366 19.3944
R20245 vdd.n1366 vdd.n1356 19.3944
R20246 vdd.n1597 vdd.n1523 19.3944
R20247 vdd.n1597 vdd.n1525 19.3944
R20248 vdd.n1593 vdd.n1525 19.3944
R20249 vdd.n1593 vdd.n1592 19.3944
R20250 vdd.n1592 vdd.n1591 19.3944
R20251 vdd.n1591 vdd.n1533 19.3944
R20252 vdd.n1587 vdd.n1533 19.3944
R20253 vdd.n1587 vdd.n1586 19.3944
R20254 vdd.n1586 vdd.n1585 19.3944
R20255 vdd.n1585 vdd.n1541 19.3944
R20256 vdd.n1581 vdd.n1541 19.3944
R20257 vdd.n1581 vdd.n1580 19.3944
R20258 vdd.n1580 vdd.n1579 19.3944
R20259 vdd.n1579 vdd.n1549 19.3944
R20260 vdd.n1575 vdd.n1549 19.3944
R20261 vdd.n1575 vdd.n1574 19.3944
R20262 vdd.n1574 vdd.n1573 19.3944
R20263 vdd.n1573 vdd.n1557 19.3944
R20264 vdd.n1569 vdd.n1557 19.3944
R20265 vdd.n1569 vdd.n1568 19.3944
R20266 vdd.n1635 vdd.n1634 19.3944
R20267 vdd.n1634 vdd.n1633 19.3944
R20268 vdd.n1633 vdd.n1486 19.3944
R20269 vdd.n1629 vdd.n1486 19.3944
R20270 vdd.n1629 vdd.n1628 19.3944
R20271 vdd.n1628 vdd.n1627 19.3944
R20272 vdd.n1627 vdd.n1494 19.3944
R20273 vdd.n1623 vdd.n1494 19.3944
R20274 vdd.n1623 vdd.n1622 19.3944
R20275 vdd.n1622 vdd.n1621 19.3944
R20276 vdd.n1621 vdd.n1502 19.3944
R20277 vdd.n1617 vdd.n1502 19.3944
R20278 vdd.n1617 vdd.n1616 19.3944
R20279 vdd.n1616 vdd.n1615 19.3944
R20280 vdd.n1615 vdd.n1510 19.3944
R20281 vdd.n1611 vdd.n1510 19.3944
R20282 vdd.n1611 vdd.n1610 19.3944
R20283 vdd.n1610 vdd.n1609 19.3944
R20284 vdd.n1609 vdd.n1518 19.3944
R20285 vdd.n1605 vdd.n1518 19.3944
R20286 vdd.n1665 vdd.n1664 19.3944
R20287 vdd.n1664 vdd.n1663 19.3944
R20288 vdd.n1663 vdd.n1444 19.3944
R20289 vdd.n1659 vdd.n1444 19.3944
R20290 vdd.n1659 vdd.n1658 19.3944
R20291 vdd.n1658 vdd.n1657 19.3944
R20292 vdd.n1657 vdd.n1452 19.3944
R20293 vdd.n1653 vdd.n1452 19.3944
R20294 vdd.n1653 vdd.n1652 19.3944
R20295 vdd.n1652 vdd.n1651 19.3944
R20296 vdd.n1651 vdd.n1460 19.3944
R20297 vdd.n1647 vdd.n1460 19.3944
R20298 vdd.n1647 vdd.n1646 19.3944
R20299 vdd.n1646 vdd.n1645 19.3944
R20300 vdd.n1645 vdd.n1468 19.3944
R20301 vdd.n1641 vdd.n1468 19.3944
R20302 vdd.n1641 vdd.n1640 19.3944
R20303 vdd.n1640 vdd.n1639 19.3944
R20304 vdd.n2108 vdd.n1075 19.3944
R20305 vdd.n2108 vdd.n1081 19.3944
R20306 vdd.n2103 vdd.n1081 19.3944
R20307 vdd.n2103 vdd.n2102 19.3944
R20308 vdd.n2102 vdd.n2101 19.3944
R20309 vdd.n2101 vdd.n1088 19.3944
R20310 vdd.n2096 vdd.n1088 19.3944
R20311 vdd.n2096 vdd.n2095 19.3944
R20312 vdd.n2095 vdd.n2094 19.3944
R20313 vdd.n2094 vdd.n1095 19.3944
R20314 vdd.n2089 vdd.n1095 19.3944
R20315 vdd.n2089 vdd.n2088 19.3944
R20316 vdd.n2088 vdd.n2087 19.3944
R20317 vdd.n2087 vdd.n1102 19.3944
R20318 vdd.n2082 vdd.n1102 19.3944
R20319 vdd.n2082 vdd.n2081 19.3944
R20320 vdd.n1349 vdd.n1107 19.3944
R20321 vdd.n2077 vdd.n1346 19.3944
R20322 vdd.n2147 vdd.n1035 19.3944
R20323 vdd.n2147 vdd.n1041 19.3944
R20324 vdd.n2142 vdd.n1041 19.3944
R20325 vdd.n2142 vdd.n2141 19.3944
R20326 vdd.n2141 vdd.n2140 19.3944
R20327 vdd.n2140 vdd.n1048 19.3944
R20328 vdd.n2135 vdd.n1048 19.3944
R20329 vdd.n2135 vdd.n2134 19.3944
R20330 vdd.n2134 vdd.n2133 19.3944
R20331 vdd.n2133 vdd.n1055 19.3944
R20332 vdd.n2128 vdd.n1055 19.3944
R20333 vdd.n2128 vdd.n2127 19.3944
R20334 vdd.n2127 vdd.n2126 19.3944
R20335 vdd.n2126 vdd.n1062 19.3944
R20336 vdd.n2121 vdd.n1062 19.3944
R20337 vdd.n2121 vdd.n2120 19.3944
R20338 vdd.n2120 vdd.n2119 19.3944
R20339 vdd.n2119 vdd.n1069 19.3944
R20340 vdd.n2114 vdd.n1069 19.3944
R20341 vdd.n2114 vdd.n2113 19.3944
R20342 vdd.n2184 vdd.n1010 19.3944
R20343 vdd.n2184 vdd.n1011 19.3944
R20344 vdd.n2179 vdd.n2178 19.3944
R20345 vdd.n2174 vdd.n2173 19.3944
R20346 vdd.n2173 vdd.n2172 19.3944
R20347 vdd.n2172 vdd.n1015 19.3944
R20348 vdd.n2167 vdd.n1015 19.3944
R20349 vdd.n2167 vdd.n2166 19.3944
R20350 vdd.n2166 vdd.n2165 19.3944
R20351 vdd.n2165 vdd.n1022 19.3944
R20352 vdd.n2160 vdd.n1022 19.3944
R20353 vdd.n2160 vdd.n2159 19.3944
R20354 vdd.n2159 vdd.n2158 19.3944
R20355 vdd.n2158 vdd.n1029 19.3944
R20356 vdd.n2153 vdd.n1029 19.3944
R20357 vdd.n2153 vdd.n2152 19.3944
R20358 vdd.n1668 vdd.n1431 19.3944
R20359 vdd.n1680 vdd.n1431 19.3944
R20360 vdd.n1680 vdd.n1429 19.3944
R20361 vdd.n1684 vdd.n1429 19.3944
R20362 vdd.n1684 vdd.n1419 19.3944
R20363 vdd.n1696 vdd.n1419 19.3944
R20364 vdd.n1696 vdd.n1417 19.3944
R20365 vdd.n1700 vdd.n1417 19.3944
R20366 vdd.n1700 vdd.n1407 19.3944
R20367 vdd.n1713 vdd.n1407 19.3944
R20368 vdd.n1713 vdd.n1405 19.3944
R20369 vdd.n1717 vdd.n1405 19.3944
R20370 vdd.n1717 vdd.n1396 19.3944
R20371 vdd.n1729 vdd.n1396 19.3944
R20372 vdd.n1729 vdd.n1394 19.3944
R20373 vdd.n2015 vdd.n1394 19.3944
R20374 vdd.n2015 vdd.n1384 19.3944
R20375 vdd.n2028 vdd.n1384 19.3944
R20376 vdd.n2028 vdd.n1382 19.3944
R20377 vdd.n2032 vdd.n1382 19.3944
R20378 vdd.n2032 vdd.n1373 19.3944
R20379 vdd.n2045 vdd.n1373 19.3944
R20380 vdd.n2045 vdd.n1371 19.3944
R20381 vdd.n2049 vdd.n1371 19.3944
R20382 vdd.n2049 vdd.n1361 19.3944
R20383 vdd.n2064 vdd.n1361 19.3944
R20384 vdd.n2064 vdd.n1359 19.3944
R20385 vdd.n2068 vdd.n1359 19.3944
R20386 vdd.n3214 vdd.n513 19.3944
R20387 vdd.n3218 vdd.n513 19.3944
R20388 vdd.n3218 vdd.n503 19.3944
R20389 vdd.n3230 vdd.n503 19.3944
R20390 vdd.n3230 vdd.n501 19.3944
R20391 vdd.n3234 vdd.n501 19.3944
R20392 vdd.n3234 vdd.n490 19.3944
R20393 vdd.n3246 vdd.n490 19.3944
R20394 vdd.n3246 vdd.n488 19.3944
R20395 vdd.n3250 vdd.n488 19.3944
R20396 vdd.n3250 vdd.n478 19.3944
R20397 vdd.n3263 vdd.n478 19.3944
R20398 vdd.n3263 vdd.n476 19.3944
R20399 vdd.n3267 vdd.n476 19.3944
R20400 vdd.n3268 vdd.n3267 19.3944
R20401 vdd.n3269 vdd.n3268 19.3944
R20402 vdd.n3269 vdd.n474 19.3944
R20403 vdd.n3273 vdd.n474 19.3944
R20404 vdd.n3274 vdd.n3273 19.3944
R20405 vdd.n3275 vdd.n3274 19.3944
R20406 vdd.n3275 vdd.n471 19.3944
R20407 vdd.n3279 vdd.n471 19.3944
R20408 vdd.n3280 vdd.n3279 19.3944
R20409 vdd.n3281 vdd.n3280 19.3944
R20410 vdd.n3281 vdd.n468 19.3944
R20411 vdd.n3285 vdd.n468 19.3944
R20412 vdd.n3286 vdd.n3285 19.3944
R20413 vdd.n3287 vdd.n3286 19.3944
R20414 vdd.n3330 vdd.n426 19.3944
R20415 vdd.n3330 vdd.n432 19.3944
R20416 vdd.n3325 vdd.n432 19.3944
R20417 vdd.n3325 vdd.n3324 19.3944
R20418 vdd.n3324 vdd.n3323 19.3944
R20419 vdd.n3323 vdd.n439 19.3944
R20420 vdd.n3318 vdd.n439 19.3944
R20421 vdd.n3318 vdd.n3317 19.3944
R20422 vdd.n3317 vdd.n3316 19.3944
R20423 vdd.n3316 vdd.n446 19.3944
R20424 vdd.n3311 vdd.n446 19.3944
R20425 vdd.n3311 vdd.n3310 19.3944
R20426 vdd.n3310 vdd.n3309 19.3944
R20427 vdd.n3309 vdd.n453 19.3944
R20428 vdd.n3304 vdd.n453 19.3944
R20429 vdd.n3304 vdd.n3303 19.3944
R20430 vdd.n3303 vdd.n3302 19.3944
R20431 vdd.n3302 vdd.n460 19.3944
R20432 vdd.n3297 vdd.n460 19.3944
R20433 vdd.n3297 vdd.n3296 19.3944
R20434 vdd.n3369 vdd.n386 19.3944
R20435 vdd.n3369 vdd.n392 19.3944
R20436 vdd.n3364 vdd.n392 19.3944
R20437 vdd.n3364 vdd.n3363 19.3944
R20438 vdd.n3363 vdd.n3362 19.3944
R20439 vdd.n3362 vdd.n399 19.3944
R20440 vdd.n3357 vdd.n399 19.3944
R20441 vdd.n3357 vdd.n3356 19.3944
R20442 vdd.n3356 vdd.n3355 19.3944
R20443 vdd.n3355 vdd.n406 19.3944
R20444 vdd.n3350 vdd.n406 19.3944
R20445 vdd.n3350 vdd.n3349 19.3944
R20446 vdd.n3349 vdd.n3348 19.3944
R20447 vdd.n3348 vdd.n413 19.3944
R20448 vdd.n3343 vdd.n413 19.3944
R20449 vdd.n3343 vdd.n3342 19.3944
R20450 vdd.n3342 vdd.n3341 19.3944
R20451 vdd.n3341 vdd.n420 19.3944
R20452 vdd.n3336 vdd.n420 19.3944
R20453 vdd.n3336 vdd.n3335 19.3944
R20454 vdd.n3405 vdd.n3404 19.3944
R20455 vdd.n3404 vdd.n3403 19.3944
R20456 vdd.n3403 vdd.n358 19.3944
R20457 vdd.n359 vdd.n358 19.3944
R20458 vdd.n3396 vdd.n359 19.3944
R20459 vdd.n3396 vdd.n3395 19.3944
R20460 vdd.n3395 vdd.n3394 19.3944
R20461 vdd.n3394 vdd.n366 19.3944
R20462 vdd.n3389 vdd.n366 19.3944
R20463 vdd.n3389 vdd.n3388 19.3944
R20464 vdd.n3388 vdd.n3387 19.3944
R20465 vdd.n3387 vdd.n373 19.3944
R20466 vdd.n3382 vdd.n373 19.3944
R20467 vdd.n3382 vdd.n3381 19.3944
R20468 vdd.n3381 vdd.n3380 19.3944
R20469 vdd.n3380 vdd.n380 19.3944
R20470 vdd.n3375 vdd.n380 19.3944
R20471 vdd.n3375 vdd.n3374 19.3944
R20472 vdd.n3210 vdd.n509 19.3944
R20473 vdd.n3222 vdd.n509 19.3944
R20474 vdd.n3222 vdd.n507 19.3944
R20475 vdd.n3226 vdd.n507 19.3944
R20476 vdd.n3226 vdd.n497 19.3944
R20477 vdd.n3238 vdd.n497 19.3944
R20478 vdd.n3238 vdd.n495 19.3944
R20479 vdd.n3242 vdd.n495 19.3944
R20480 vdd.n3242 vdd.n485 19.3944
R20481 vdd.n3255 vdd.n485 19.3944
R20482 vdd.n3255 vdd.n483 19.3944
R20483 vdd.n3259 vdd.n483 19.3944
R20484 vdd.n3259 vdd.n312 19.3944
R20485 vdd.n3438 vdd.n312 19.3944
R20486 vdd.n3438 vdd.n313 19.3944
R20487 vdd.n3432 vdd.n313 19.3944
R20488 vdd.n3432 vdd.n3431 19.3944
R20489 vdd.n3431 vdd.n3430 19.3944
R20490 vdd.n3430 vdd.n323 19.3944
R20491 vdd.n3424 vdd.n323 19.3944
R20492 vdd.n3424 vdd.n3423 19.3944
R20493 vdd.n3423 vdd.n3422 19.3944
R20494 vdd.n3422 vdd.n335 19.3944
R20495 vdd.n3416 vdd.n335 19.3944
R20496 vdd.n3416 vdd.n3415 19.3944
R20497 vdd.n3415 vdd.n3414 19.3944
R20498 vdd.n3414 vdd.n346 19.3944
R20499 vdd.n3408 vdd.n346 19.3944
R20500 vdd.n3167 vdd.n3166 19.3944
R20501 vdd.n3166 vdd.n3165 19.3944
R20502 vdd.n3165 vdd.n551 19.3944
R20503 vdd.n3159 vdd.n551 19.3944
R20504 vdd.n3159 vdd.n3158 19.3944
R20505 vdd.n3158 vdd.n3157 19.3944
R20506 vdd.n3157 vdd.n557 19.3944
R20507 vdd.n3151 vdd.n557 19.3944
R20508 vdd.n3151 vdd.n3150 19.3944
R20509 vdd.n3150 vdd.n3149 19.3944
R20510 vdd.n3149 vdd.n563 19.3944
R20511 vdd.n3143 vdd.n563 19.3944
R20512 vdd.n3143 vdd.n3142 19.3944
R20513 vdd.n3142 vdd.n3141 19.3944
R20514 vdd.n3141 vdd.n569 19.3944
R20515 vdd.n3135 vdd.n569 19.3944
R20516 vdd.n3135 vdd.n3134 19.3944
R20517 vdd.n3134 vdd.n3133 19.3944
R20518 vdd.n3133 vdd.n575 19.3944
R20519 vdd.n3127 vdd.n575 19.3944
R20520 vdd.n3207 vdd.n3206 19.3944
R20521 vdd.n3206 vdd.n519 19.3944
R20522 vdd.n3201 vdd.n3200 19.3944
R20523 vdd.n3197 vdd.n3196 19.3944
R20524 vdd.n3196 vdd.n525 19.3944
R20525 vdd.n3191 vdd.n525 19.3944
R20526 vdd.n3191 vdd.n3190 19.3944
R20527 vdd.n3190 vdd.n3189 19.3944
R20528 vdd.n3189 vdd.n531 19.3944
R20529 vdd.n3183 vdd.n531 19.3944
R20530 vdd.n3183 vdd.n3182 19.3944
R20531 vdd.n3182 vdd.n3181 19.3944
R20532 vdd.n3181 vdd.n537 19.3944
R20533 vdd.n3175 vdd.n537 19.3944
R20534 vdd.n3175 vdd.n3174 19.3944
R20535 vdd.n3174 vdd.n3173 19.3944
R20536 vdd.n3122 vdd.n579 19.3944
R20537 vdd.n3122 vdd.n583 19.3944
R20538 vdd.n3117 vdd.n583 19.3944
R20539 vdd.n3117 vdd.n3116 19.3944
R20540 vdd.n3116 vdd.n589 19.3944
R20541 vdd.n3111 vdd.n589 19.3944
R20542 vdd.n3111 vdd.n3110 19.3944
R20543 vdd.n3110 vdd.n3109 19.3944
R20544 vdd.n3109 vdd.n595 19.3944
R20545 vdd.n3103 vdd.n595 19.3944
R20546 vdd.n3103 vdd.n3102 19.3944
R20547 vdd.n3102 vdd.n3101 19.3944
R20548 vdd.n3101 vdd.n601 19.3944
R20549 vdd.n3095 vdd.n601 19.3944
R20550 vdd.n3095 vdd.n3094 19.3944
R20551 vdd.n3094 vdd.n3093 19.3944
R20552 vdd.n3089 vdd.n3088 19.3944
R20553 vdd.n3085 vdd.n3084 19.3944
R20554 vdd.n1604 vdd.n1523 19.0066
R20555 vdd.n2112 vdd.n1075 19.0066
R20556 vdd.n3334 vdd.n426 19.0066
R20557 vdd.n3126 vdd.n579 19.0066
R20558 vdd.n1144 vdd.n1143 16.0975
R20559 vdd.n839 vdd.n838 16.0975
R20560 vdd.n1566 vdd.n1565 16.0975
R20561 vdd.n1603 vdd.n1602 16.0975
R20562 vdd.n1477 vdd.n1476 16.0975
R20563 vdd.n2075 vdd.n2074 16.0975
R20564 vdd.n1077 vdd.n1076 16.0975
R20565 vdd.n1037 vdd.n1036 16.0975
R20566 vdd.n1148 vdd.n1147 16.0975
R20567 vdd.n830 vdd.n829 16.0975
R20568 vdd.n2536 vdd.n2535 16.0975
R20569 vdd.n3294 vdd.n3293 16.0975
R20570 vdd.n428 vdd.n427 16.0975
R20571 vdd.n388 vdd.n387 16.0975
R20572 vdd.n581 vdd.n580 16.0975
R20573 vdd.n544 vdd.n543 16.0975
R20574 vdd.n662 vdd.n661 16.0975
R20575 vdd.n2533 vdd.n2532 16.0975
R20576 vdd.n3081 vdd.n3080 16.0975
R20577 vdd.n626 vdd.n625 16.0975
R20578 vdd.t188 vdd.n2496 15.4182
R20579 vdd.n2800 vdd.t164 15.4182
R20580 vdd.n28 vdd.n27 14.8792
R20581 vdd.n304 vdd.n269 13.1884
R20582 vdd.n253 vdd.n218 13.1884
R20583 vdd.n210 vdd.n175 13.1884
R20584 vdd.n159 vdd.n124 13.1884
R20585 vdd.n117 vdd.n82 13.1884
R20586 vdd.n66 vdd.n31 13.1884
R20587 vdd.n1954 vdd.n1919 13.1884
R20588 vdd.n2005 vdd.n1970 13.1884
R20589 vdd.n1860 vdd.n1825 13.1884
R20590 vdd.n1911 vdd.n1876 13.1884
R20591 vdd.n1767 vdd.n1732 13.1884
R20592 vdd.n1818 vdd.n1783 13.1884
R20593 vdd.n2218 vdd.n962 13.1509
R20594 vdd.n3043 vdd.n613 13.1509
R20595 vdd.n1635 vdd.n1478 12.9944
R20596 vdd.n1639 vdd.n1478 12.9944
R20597 vdd.n2151 vdd.n1035 12.9944
R20598 vdd.n2152 vdd.n2151 12.9944
R20599 vdd.n3373 vdd.n386 12.9944
R20600 vdd.n3374 vdd.n3373 12.9944
R20601 vdd.n3167 vdd.n545 12.9944
R20602 vdd.n3173 vdd.n545 12.9944
R20603 vdd.n305 vdd.n267 12.8005
R20604 vdd.n300 vdd.n271 12.8005
R20605 vdd.n254 vdd.n216 12.8005
R20606 vdd.n249 vdd.n220 12.8005
R20607 vdd.n211 vdd.n173 12.8005
R20608 vdd.n206 vdd.n177 12.8005
R20609 vdd.n160 vdd.n122 12.8005
R20610 vdd.n155 vdd.n126 12.8005
R20611 vdd.n118 vdd.n80 12.8005
R20612 vdd.n113 vdd.n84 12.8005
R20613 vdd.n67 vdd.n29 12.8005
R20614 vdd.n62 vdd.n33 12.8005
R20615 vdd.n1955 vdd.n1917 12.8005
R20616 vdd.n1950 vdd.n1921 12.8005
R20617 vdd.n2006 vdd.n1968 12.8005
R20618 vdd.n2001 vdd.n1972 12.8005
R20619 vdd.n1861 vdd.n1823 12.8005
R20620 vdd.n1856 vdd.n1827 12.8005
R20621 vdd.n1912 vdd.n1874 12.8005
R20622 vdd.n1907 vdd.n1878 12.8005
R20623 vdd.n1768 vdd.n1730 12.8005
R20624 vdd.n1763 vdd.n1734 12.8005
R20625 vdd.n1819 vdd.n1781 12.8005
R20626 vdd.n1814 vdd.n1785 12.8005
R20627 vdd.n299 vdd.n272 12.0247
R20628 vdd.n248 vdd.n221 12.0247
R20629 vdd.n205 vdd.n178 12.0247
R20630 vdd.n154 vdd.n127 12.0247
R20631 vdd.n112 vdd.n85 12.0247
R20632 vdd.n61 vdd.n34 12.0247
R20633 vdd.n1949 vdd.n1922 12.0247
R20634 vdd.n2000 vdd.n1973 12.0247
R20635 vdd.n1855 vdd.n1828 12.0247
R20636 vdd.n1906 vdd.n1879 12.0247
R20637 vdd.n1762 vdd.n1735 12.0247
R20638 vdd.n1813 vdd.n1786 12.0247
R20639 vdd.n1670 vdd.n1438 11.337
R20640 vdd.n1678 vdd.n1427 11.337
R20641 vdd.n1686 vdd.n1427 11.337
R20642 vdd.n1694 vdd.n1421 11.337
R20643 vdd.n1702 vdd.n1414 11.337
R20644 vdd.n1711 vdd.n1710 11.337
R20645 vdd.n1719 vdd.n1403 11.337
R20646 vdd.n2017 vdd.n1392 11.337
R20647 vdd.n2026 vdd.n1386 11.337
R20648 vdd.n2034 vdd.n1380 11.337
R20649 vdd.n2043 vdd.n2042 11.337
R20650 vdd.n2051 vdd.n1363 11.337
R20651 vdd.n2062 vdd.n1363 11.337
R20652 vdd.n2062 vdd.n2061 11.337
R20653 vdd.n3220 vdd.n511 11.337
R20654 vdd.n3220 vdd.n505 11.337
R20655 vdd.n3228 vdd.n505 11.337
R20656 vdd.n3236 vdd.n499 11.337
R20657 vdd.n3244 vdd.n492 11.337
R20658 vdd.n3253 vdd.n3252 11.337
R20659 vdd.n3261 vdd.n481 11.337
R20660 vdd.n3435 vdd.n3434 11.337
R20661 vdd.n3428 vdd.n325 11.337
R20662 vdd.n3426 vdd.n329 11.337
R20663 vdd.n3420 vdd.n3419 11.337
R20664 vdd.n3418 vdd.n340 11.337
R20665 vdd.n3412 vdd.n340 11.337
R20666 vdd.n3411 vdd.n3410 11.337
R20667 vdd.n296 vdd.n295 11.249
R20668 vdd.n245 vdd.n244 11.249
R20669 vdd.n202 vdd.n201 11.249
R20670 vdd.n151 vdd.n150 11.249
R20671 vdd.n109 vdd.n108 11.249
R20672 vdd.n58 vdd.n57 11.249
R20673 vdd.n1946 vdd.n1945 11.249
R20674 vdd.n1997 vdd.n1996 11.249
R20675 vdd.n1852 vdd.n1851 11.249
R20676 vdd.n1903 vdd.n1902 11.249
R20677 vdd.n1759 vdd.n1758 11.249
R20678 vdd.n1810 vdd.n1809 11.249
R20679 vdd.n1686 vdd.t131 10.9969
R20680 vdd.t22 vdd.n3418 10.9969
R20681 vdd.n1415 vdd.t108 10.7702
R20682 vdd.t128 vdd.n3427 10.7702
R20683 vdd.n281 vdd.n280 10.7238
R20684 vdd.n230 vdd.n229 10.7238
R20685 vdd.n187 vdd.n186 10.7238
R20686 vdd.n136 vdd.n135 10.7238
R20687 vdd.n94 vdd.n93 10.7238
R20688 vdd.n43 vdd.n42 10.7238
R20689 vdd.n1931 vdd.n1930 10.7238
R20690 vdd.n1982 vdd.n1981 10.7238
R20691 vdd.n1837 vdd.n1836 10.7238
R20692 vdd.n1888 vdd.n1887 10.7238
R20693 vdd.n1744 vdd.n1743 10.7238
R20694 vdd.n1795 vdd.n1794 10.7238
R20695 vdd.n2223 vdd.n2222 10.6151
R20696 vdd.n2223 vdd.n955 10.6151
R20697 vdd.n2233 vdd.n955 10.6151
R20698 vdd.n2234 vdd.n2233 10.6151
R20699 vdd.n2235 vdd.n2234 10.6151
R20700 vdd.n2235 vdd.n942 10.6151
R20701 vdd.n2245 vdd.n942 10.6151
R20702 vdd.n2246 vdd.n2245 10.6151
R20703 vdd.n2247 vdd.n2246 10.6151
R20704 vdd.n2247 vdd.n930 10.6151
R20705 vdd.n2257 vdd.n930 10.6151
R20706 vdd.n2258 vdd.n2257 10.6151
R20707 vdd.n2259 vdd.n2258 10.6151
R20708 vdd.n2259 vdd.n919 10.6151
R20709 vdd.n2269 vdd.n919 10.6151
R20710 vdd.n2270 vdd.n2269 10.6151
R20711 vdd.n2271 vdd.n2270 10.6151
R20712 vdd.n2271 vdd.n906 10.6151
R20713 vdd.n2281 vdd.n906 10.6151
R20714 vdd.n2282 vdd.n2281 10.6151
R20715 vdd.n2283 vdd.n2282 10.6151
R20716 vdd.n2283 vdd.n894 10.6151
R20717 vdd.n2294 vdd.n894 10.6151
R20718 vdd.n2295 vdd.n2294 10.6151
R20719 vdd.n2296 vdd.n2295 10.6151
R20720 vdd.n2296 vdd.n882 10.6151
R20721 vdd.n2306 vdd.n882 10.6151
R20722 vdd.n2307 vdd.n2306 10.6151
R20723 vdd.n2308 vdd.n2307 10.6151
R20724 vdd.n2308 vdd.n870 10.6151
R20725 vdd.n2318 vdd.n870 10.6151
R20726 vdd.n2319 vdd.n2318 10.6151
R20727 vdd.n2320 vdd.n2319 10.6151
R20728 vdd.n2320 vdd.n860 10.6151
R20729 vdd.n2330 vdd.n860 10.6151
R20730 vdd.n2331 vdd.n2330 10.6151
R20731 vdd.n2332 vdd.n2331 10.6151
R20732 vdd.n2332 vdd.n847 10.6151
R20733 vdd.n2344 vdd.n847 10.6151
R20734 vdd.n2345 vdd.n2344 10.6151
R20735 vdd.n2347 vdd.n2345 10.6151
R20736 vdd.n2347 vdd.n2346 10.6151
R20737 vdd.n2346 vdd.n828 10.6151
R20738 vdd.n2494 vdd.n2493 10.6151
R20739 vdd.n2493 vdd.n2492 10.6151
R20740 vdd.n2492 vdd.n2489 10.6151
R20741 vdd.n2489 vdd.n2488 10.6151
R20742 vdd.n2488 vdd.n2485 10.6151
R20743 vdd.n2485 vdd.n2484 10.6151
R20744 vdd.n2484 vdd.n2481 10.6151
R20745 vdd.n2481 vdd.n2480 10.6151
R20746 vdd.n2480 vdd.n2477 10.6151
R20747 vdd.n2477 vdd.n2476 10.6151
R20748 vdd.n2476 vdd.n2473 10.6151
R20749 vdd.n2473 vdd.n2472 10.6151
R20750 vdd.n2472 vdd.n2469 10.6151
R20751 vdd.n2469 vdd.n2468 10.6151
R20752 vdd.n2468 vdd.n2465 10.6151
R20753 vdd.n2465 vdd.n2464 10.6151
R20754 vdd.n2464 vdd.n2461 10.6151
R20755 vdd.n2461 vdd.n2460 10.6151
R20756 vdd.n2460 vdd.n2457 10.6151
R20757 vdd.n2457 vdd.n2456 10.6151
R20758 vdd.n2456 vdd.n2453 10.6151
R20759 vdd.n2453 vdd.n2452 10.6151
R20760 vdd.n2452 vdd.n2449 10.6151
R20761 vdd.n2449 vdd.n2448 10.6151
R20762 vdd.n2448 vdd.n2445 10.6151
R20763 vdd.n2445 vdd.n2444 10.6151
R20764 vdd.n2444 vdd.n2441 10.6151
R20765 vdd.n2441 vdd.n2440 10.6151
R20766 vdd.n2440 vdd.n2437 10.6151
R20767 vdd.n2437 vdd.n2436 10.6151
R20768 vdd.n2436 vdd.n2433 10.6151
R20769 vdd.n2431 vdd.n2428 10.6151
R20770 vdd.n2428 vdd.n2427 10.6151
R20771 vdd.n1185 vdd.n1184 10.6151
R20772 vdd.n1187 vdd.n1185 10.6151
R20773 vdd.n1188 vdd.n1187 10.6151
R20774 vdd.n1190 vdd.n1188 10.6151
R20775 vdd.n1191 vdd.n1190 10.6151
R20776 vdd.n1193 vdd.n1191 10.6151
R20777 vdd.n1194 vdd.n1193 10.6151
R20778 vdd.n1196 vdd.n1194 10.6151
R20779 vdd.n1197 vdd.n1196 10.6151
R20780 vdd.n1199 vdd.n1197 10.6151
R20781 vdd.n1200 vdd.n1199 10.6151
R20782 vdd.n1202 vdd.n1200 10.6151
R20783 vdd.n1203 vdd.n1202 10.6151
R20784 vdd.n1205 vdd.n1203 10.6151
R20785 vdd.n1206 vdd.n1205 10.6151
R20786 vdd.n1208 vdd.n1206 10.6151
R20787 vdd.n1209 vdd.n1208 10.6151
R20788 vdd.n1211 vdd.n1209 10.6151
R20789 vdd.n1212 vdd.n1211 10.6151
R20790 vdd.n1214 vdd.n1212 10.6151
R20791 vdd.n1215 vdd.n1214 10.6151
R20792 vdd.n1217 vdd.n1215 10.6151
R20793 vdd.n1218 vdd.n1217 10.6151
R20794 vdd.n1220 vdd.n1218 10.6151
R20795 vdd.n1221 vdd.n1220 10.6151
R20796 vdd.n1223 vdd.n1221 10.6151
R20797 vdd.n1224 vdd.n1223 10.6151
R20798 vdd.n1263 vdd.n1224 10.6151
R20799 vdd.n1263 vdd.n1262 10.6151
R20800 vdd.n1262 vdd.n1261 10.6151
R20801 vdd.n1261 vdd.n1259 10.6151
R20802 vdd.n1259 vdd.n1258 10.6151
R20803 vdd.n1258 vdd.n1256 10.6151
R20804 vdd.n1256 vdd.n1255 10.6151
R20805 vdd.n1255 vdd.n1236 10.6151
R20806 vdd.n1236 vdd.n1235 10.6151
R20807 vdd.n1235 vdd.n1233 10.6151
R20808 vdd.n1233 vdd.n1232 10.6151
R20809 vdd.n1232 vdd.n1230 10.6151
R20810 vdd.n1230 vdd.n1229 10.6151
R20811 vdd.n1229 vdd.n1226 10.6151
R20812 vdd.n1226 vdd.n1225 10.6151
R20813 vdd.n1225 vdd.n831 10.6151
R20814 vdd.n2221 vdd.n967 10.6151
R20815 vdd.n2216 vdd.n967 10.6151
R20816 vdd.n2216 vdd.n2215 10.6151
R20817 vdd.n2215 vdd.n2214 10.6151
R20818 vdd.n2214 vdd.n2211 10.6151
R20819 vdd.n2211 vdd.n2210 10.6151
R20820 vdd.n2210 vdd.n2207 10.6151
R20821 vdd.n2207 vdd.n2206 10.6151
R20822 vdd.n2206 vdd.n2203 10.6151
R20823 vdd.n2203 vdd.n2202 10.6151
R20824 vdd.n2202 vdd.n2199 10.6151
R20825 vdd.n2199 vdd.n2198 10.6151
R20826 vdd.n2198 vdd.n2195 10.6151
R20827 vdd.n2195 vdd.n2194 10.6151
R20828 vdd.n2194 vdd.n2191 10.6151
R20829 vdd.n2191 vdd.n2190 10.6151
R20830 vdd.n2190 vdd.n2187 10.6151
R20831 vdd.n2187 vdd.n1005 10.6151
R20832 vdd.n1151 vdd.n1005 10.6151
R20833 vdd.n1152 vdd.n1151 10.6151
R20834 vdd.n1155 vdd.n1152 10.6151
R20835 vdd.n1156 vdd.n1155 10.6151
R20836 vdd.n1159 vdd.n1156 10.6151
R20837 vdd.n1160 vdd.n1159 10.6151
R20838 vdd.n1163 vdd.n1160 10.6151
R20839 vdd.n1164 vdd.n1163 10.6151
R20840 vdd.n1167 vdd.n1164 10.6151
R20841 vdd.n1168 vdd.n1167 10.6151
R20842 vdd.n1171 vdd.n1168 10.6151
R20843 vdd.n1172 vdd.n1171 10.6151
R20844 vdd.n1175 vdd.n1172 10.6151
R20845 vdd.n1180 vdd.n1177 10.6151
R20846 vdd.n1181 vdd.n1180 10.6151
R20847 vdd.n2732 vdd.n2731 10.6151
R20848 vdd.n2731 vdd.n2730 10.6151
R20849 vdd.n2730 vdd.n2534 10.6151
R20850 vdd.n2612 vdd.n2534 10.6151
R20851 vdd.n2613 vdd.n2612 10.6151
R20852 vdd.n2615 vdd.n2613 10.6151
R20853 vdd.n2616 vdd.n2615 10.6151
R20854 vdd.n2714 vdd.n2616 10.6151
R20855 vdd.n2714 vdd.n2713 10.6151
R20856 vdd.n2713 vdd.n2712 10.6151
R20857 vdd.n2712 vdd.n2660 10.6151
R20858 vdd.n2660 vdd.n2659 10.6151
R20859 vdd.n2659 vdd.n2657 10.6151
R20860 vdd.n2657 vdd.n2656 10.6151
R20861 vdd.n2656 vdd.n2654 10.6151
R20862 vdd.n2654 vdd.n2653 10.6151
R20863 vdd.n2653 vdd.n2651 10.6151
R20864 vdd.n2651 vdd.n2650 10.6151
R20865 vdd.n2650 vdd.n2648 10.6151
R20866 vdd.n2648 vdd.n2647 10.6151
R20867 vdd.n2647 vdd.n2645 10.6151
R20868 vdd.n2645 vdd.n2644 10.6151
R20869 vdd.n2644 vdd.n2642 10.6151
R20870 vdd.n2642 vdd.n2641 10.6151
R20871 vdd.n2641 vdd.n2639 10.6151
R20872 vdd.n2639 vdd.n2638 10.6151
R20873 vdd.n2638 vdd.n2636 10.6151
R20874 vdd.n2636 vdd.n2635 10.6151
R20875 vdd.n2635 vdd.n2633 10.6151
R20876 vdd.n2633 vdd.n2632 10.6151
R20877 vdd.n2632 vdd.n2630 10.6151
R20878 vdd.n2630 vdd.n2629 10.6151
R20879 vdd.n2629 vdd.n2627 10.6151
R20880 vdd.n2627 vdd.n2626 10.6151
R20881 vdd.n2626 vdd.n2624 10.6151
R20882 vdd.n2624 vdd.n2623 10.6151
R20883 vdd.n2623 vdd.n2621 10.6151
R20884 vdd.n2621 vdd.n2620 10.6151
R20885 vdd.n2620 vdd.n2618 10.6151
R20886 vdd.n2618 vdd.n2617 10.6151
R20887 vdd.n2617 vdd.n664 10.6151
R20888 vdd.n2976 vdd.n664 10.6151
R20889 vdd.n2977 vdd.n2976 10.6151
R20890 vdd.n2803 vdd.n789 10.6151
R20891 vdd.n2798 vdd.n789 10.6151
R20892 vdd.n2798 vdd.n2797 10.6151
R20893 vdd.n2797 vdd.n2796 10.6151
R20894 vdd.n2796 vdd.n2793 10.6151
R20895 vdd.n2793 vdd.n2792 10.6151
R20896 vdd.n2792 vdd.n2789 10.6151
R20897 vdd.n2789 vdd.n2788 10.6151
R20898 vdd.n2788 vdd.n2785 10.6151
R20899 vdd.n2785 vdd.n2784 10.6151
R20900 vdd.n2784 vdd.n2781 10.6151
R20901 vdd.n2781 vdd.n2780 10.6151
R20902 vdd.n2780 vdd.n2777 10.6151
R20903 vdd.n2777 vdd.n2776 10.6151
R20904 vdd.n2776 vdd.n2773 10.6151
R20905 vdd.n2773 vdd.n2772 10.6151
R20906 vdd.n2772 vdd.n2769 10.6151
R20907 vdd.n2769 vdd.n2768 10.6151
R20908 vdd.n2768 vdd.n2765 10.6151
R20909 vdd.n2765 vdd.n2764 10.6151
R20910 vdd.n2764 vdd.n2761 10.6151
R20911 vdd.n2761 vdd.n2760 10.6151
R20912 vdd.n2760 vdd.n2757 10.6151
R20913 vdd.n2757 vdd.n2756 10.6151
R20914 vdd.n2756 vdd.n2753 10.6151
R20915 vdd.n2753 vdd.n2752 10.6151
R20916 vdd.n2752 vdd.n2749 10.6151
R20917 vdd.n2749 vdd.n2748 10.6151
R20918 vdd.n2748 vdd.n2745 10.6151
R20919 vdd.n2745 vdd.n2744 10.6151
R20920 vdd.n2744 vdd.n2741 10.6151
R20921 vdd.n2739 vdd.n2736 10.6151
R20922 vdd.n2736 vdd.n2735 10.6151
R20923 vdd.n2805 vdd.n2804 10.6151
R20924 vdd.n2805 vdd.n778 10.6151
R20925 vdd.n2815 vdd.n778 10.6151
R20926 vdd.n2816 vdd.n2815 10.6151
R20927 vdd.n2817 vdd.n2816 10.6151
R20928 vdd.n2817 vdd.n766 10.6151
R20929 vdd.n2827 vdd.n766 10.6151
R20930 vdd.n2828 vdd.n2827 10.6151
R20931 vdd.n2829 vdd.n2828 10.6151
R20932 vdd.n2829 vdd.n755 10.6151
R20933 vdd.n2839 vdd.n755 10.6151
R20934 vdd.n2840 vdd.n2839 10.6151
R20935 vdd.n2841 vdd.n2840 10.6151
R20936 vdd.n2841 vdd.n744 10.6151
R20937 vdd.n2851 vdd.n744 10.6151
R20938 vdd.n2852 vdd.n2851 10.6151
R20939 vdd.n2853 vdd.n2852 10.6151
R20940 vdd.n2853 vdd.n731 10.6151
R20941 vdd.n2864 vdd.n731 10.6151
R20942 vdd.n2865 vdd.n2864 10.6151
R20943 vdd.n2866 vdd.n2865 10.6151
R20944 vdd.n2866 vdd.n719 10.6151
R20945 vdd.n2876 vdd.n719 10.6151
R20946 vdd.n2877 vdd.n2876 10.6151
R20947 vdd.n2878 vdd.n2877 10.6151
R20948 vdd.n2878 vdd.n707 10.6151
R20949 vdd.n2888 vdd.n707 10.6151
R20950 vdd.n2889 vdd.n2888 10.6151
R20951 vdd.n2890 vdd.n2889 10.6151
R20952 vdd.n2890 vdd.n694 10.6151
R20953 vdd.n2900 vdd.n694 10.6151
R20954 vdd.n2901 vdd.n2900 10.6151
R20955 vdd.n2902 vdd.n2901 10.6151
R20956 vdd.n2902 vdd.n683 10.6151
R20957 vdd.n2912 vdd.n683 10.6151
R20958 vdd.n2913 vdd.n2912 10.6151
R20959 vdd.n2914 vdd.n2913 10.6151
R20960 vdd.n2914 vdd.n669 10.6151
R20961 vdd.n2969 vdd.n669 10.6151
R20962 vdd.n2970 vdd.n2969 10.6151
R20963 vdd.n2971 vdd.n2970 10.6151
R20964 vdd.n2971 vdd.n636 10.6151
R20965 vdd.n3041 vdd.n636 10.6151
R20966 vdd.n3040 vdd.n3039 10.6151
R20967 vdd.n3039 vdd.n637 10.6151
R20968 vdd.n638 vdd.n637 10.6151
R20969 vdd.n3032 vdd.n638 10.6151
R20970 vdd.n3032 vdd.n3031 10.6151
R20971 vdd.n3031 vdd.n3030 10.6151
R20972 vdd.n3030 vdd.n640 10.6151
R20973 vdd.n3025 vdd.n640 10.6151
R20974 vdd.n3025 vdd.n3024 10.6151
R20975 vdd.n3024 vdd.n3023 10.6151
R20976 vdd.n3023 vdd.n643 10.6151
R20977 vdd.n3018 vdd.n643 10.6151
R20978 vdd.n3018 vdd.n3017 10.6151
R20979 vdd.n3017 vdd.n3016 10.6151
R20980 vdd.n3016 vdd.n646 10.6151
R20981 vdd.n3011 vdd.n646 10.6151
R20982 vdd.n3011 vdd.n3010 10.6151
R20983 vdd.n3010 vdd.n3008 10.6151
R20984 vdd.n3008 vdd.n649 10.6151
R20985 vdd.n3003 vdd.n649 10.6151
R20986 vdd.n3003 vdd.n3002 10.6151
R20987 vdd.n3002 vdd.n3001 10.6151
R20988 vdd.n3001 vdd.n652 10.6151
R20989 vdd.n2996 vdd.n652 10.6151
R20990 vdd.n2996 vdd.n2995 10.6151
R20991 vdd.n2995 vdd.n2994 10.6151
R20992 vdd.n2994 vdd.n655 10.6151
R20993 vdd.n2989 vdd.n655 10.6151
R20994 vdd.n2989 vdd.n2988 10.6151
R20995 vdd.n2988 vdd.n2987 10.6151
R20996 vdd.n2987 vdd.n658 10.6151
R20997 vdd.n2982 vdd.n2981 10.6151
R20998 vdd.n2981 vdd.n2980 10.6151
R20999 vdd.n2959 vdd.n2920 10.6151
R21000 vdd.n2954 vdd.n2920 10.6151
R21001 vdd.n2954 vdd.n2953 10.6151
R21002 vdd.n2953 vdd.n2952 10.6151
R21003 vdd.n2952 vdd.n2922 10.6151
R21004 vdd.n2947 vdd.n2922 10.6151
R21005 vdd.n2947 vdd.n2946 10.6151
R21006 vdd.n2946 vdd.n2945 10.6151
R21007 vdd.n2945 vdd.n2925 10.6151
R21008 vdd.n2940 vdd.n2925 10.6151
R21009 vdd.n2940 vdd.n2939 10.6151
R21010 vdd.n2939 vdd.n2938 10.6151
R21011 vdd.n2938 vdd.n2928 10.6151
R21012 vdd.n2933 vdd.n2928 10.6151
R21013 vdd.n2933 vdd.n2932 10.6151
R21014 vdd.n2932 vdd.n610 10.6151
R21015 vdd.n3076 vdd.n610 10.6151
R21016 vdd.n3076 vdd.n611 10.6151
R21017 vdd.n614 vdd.n611 10.6151
R21018 vdd.n3069 vdd.n614 10.6151
R21019 vdd.n3069 vdd.n3068 10.6151
R21020 vdd.n3068 vdd.n3067 10.6151
R21021 vdd.n3067 vdd.n616 10.6151
R21022 vdd.n3062 vdd.n616 10.6151
R21023 vdd.n3062 vdd.n3061 10.6151
R21024 vdd.n3061 vdd.n3060 10.6151
R21025 vdd.n3060 vdd.n619 10.6151
R21026 vdd.n3055 vdd.n619 10.6151
R21027 vdd.n3055 vdd.n3054 10.6151
R21028 vdd.n3054 vdd.n3053 10.6151
R21029 vdd.n3053 vdd.n622 10.6151
R21030 vdd.n3048 vdd.n3047 10.6151
R21031 vdd.n3047 vdd.n3046 10.6151
R21032 vdd.n2609 vdd.n2608 10.6151
R21033 vdd.n2726 vdd.n2609 10.6151
R21034 vdd.n2726 vdd.n2725 10.6151
R21035 vdd.n2725 vdd.n2724 10.6151
R21036 vdd.n2724 vdd.n2722 10.6151
R21037 vdd.n2722 vdd.n2721 10.6151
R21038 vdd.n2721 vdd.n2719 10.6151
R21039 vdd.n2719 vdd.n2718 10.6151
R21040 vdd.n2718 vdd.n2610 10.6151
R21041 vdd.n2708 vdd.n2610 10.6151
R21042 vdd.n2708 vdd.n2707 10.6151
R21043 vdd.n2707 vdd.n2706 10.6151
R21044 vdd.n2706 vdd.n2704 10.6151
R21045 vdd.n2704 vdd.n2703 10.6151
R21046 vdd.n2703 vdd.n2701 10.6151
R21047 vdd.n2701 vdd.n2700 10.6151
R21048 vdd.n2700 vdd.n2698 10.6151
R21049 vdd.n2698 vdd.n2697 10.6151
R21050 vdd.n2697 vdd.n2695 10.6151
R21051 vdd.n2695 vdd.n2694 10.6151
R21052 vdd.n2694 vdd.n2692 10.6151
R21053 vdd.n2692 vdd.n2691 10.6151
R21054 vdd.n2691 vdd.n2689 10.6151
R21055 vdd.n2689 vdd.n2688 10.6151
R21056 vdd.n2688 vdd.n2686 10.6151
R21057 vdd.n2686 vdd.n2685 10.6151
R21058 vdd.n2685 vdd.n2683 10.6151
R21059 vdd.n2683 vdd.n2682 10.6151
R21060 vdd.n2682 vdd.n2680 10.6151
R21061 vdd.n2680 vdd.n2679 10.6151
R21062 vdd.n2679 vdd.n2677 10.6151
R21063 vdd.n2677 vdd.n2676 10.6151
R21064 vdd.n2676 vdd.n2674 10.6151
R21065 vdd.n2674 vdd.n2673 10.6151
R21066 vdd.n2673 vdd.n2671 10.6151
R21067 vdd.n2671 vdd.n2670 10.6151
R21068 vdd.n2670 vdd.n2668 10.6151
R21069 vdd.n2668 vdd.n2667 10.6151
R21070 vdd.n2667 vdd.n2665 10.6151
R21071 vdd.n2665 vdd.n2664 10.6151
R21072 vdd.n2664 vdd.n2662 10.6151
R21073 vdd.n2662 vdd.n2661 10.6151
R21074 vdd.n2661 vdd.n628 10.6151
R21075 vdd.n2540 vdd.n2539 10.6151
R21076 vdd.n2543 vdd.n2540 10.6151
R21077 vdd.n2544 vdd.n2543 10.6151
R21078 vdd.n2547 vdd.n2544 10.6151
R21079 vdd.n2548 vdd.n2547 10.6151
R21080 vdd.n2551 vdd.n2548 10.6151
R21081 vdd.n2552 vdd.n2551 10.6151
R21082 vdd.n2555 vdd.n2552 10.6151
R21083 vdd.n2556 vdd.n2555 10.6151
R21084 vdd.n2559 vdd.n2556 10.6151
R21085 vdd.n2560 vdd.n2559 10.6151
R21086 vdd.n2563 vdd.n2560 10.6151
R21087 vdd.n2564 vdd.n2563 10.6151
R21088 vdd.n2567 vdd.n2564 10.6151
R21089 vdd.n2568 vdd.n2567 10.6151
R21090 vdd.n2571 vdd.n2568 10.6151
R21091 vdd.n2572 vdd.n2571 10.6151
R21092 vdd.n2575 vdd.n2572 10.6151
R21093 vdd.n2576 vdd.n2575 10.6151
R21094 vdd.n2579 vdd.n2576 10.6151
R21095 vdd.n2580 vdd.n2579 10.6151
R21096 vdd.n2583 vdd.n2580 10.6151
R21097 vdd.n2584 vdd.n2583 10.6151
R21098 vdd.n2587 vdd.n2584 10.6151
R21099 vdd.n2588 vdd.n2587 10.6151
R21100 vdd.n2591 vdd.n2588 10.6151
R21101 vdd.n2592 vdd.n2591 10.6151
R21102 vdd.n2595 vdd.n2592 10.6151
R21103 vdd.n2596 vdd.n2595 10.6151
R21104 vdd.n2599 vdd.n2596 10.6151
R21105 vdd.n2600 vdd.n2599 10.6151
R21106 vdd.n2605 vdd.n2603 10.6151
R21107 vdd.n2606 vdd.n2605 10.6151
R21108 vdd.n2809 vdd.n783 10.6151
R21109 vdd.n2810 vdd.n2809 10.6151
R21110 vdd.n2811 vdd.n2810 10.6151
R21111 vdd.n2811 vdd.n772 10.6151
R21112 vdd.n2821 vdd.n772 10.6151
R21113 vdd.n2822 vdd.n2821 10.6151
R21114 vdd.n2823 vdd.n2822 10.6151
R21115 vdd.n2823 vdd.n761 10.6151
R21116 vdd.n2833 vdd.n761 10.6151
R21117 vdd.n2834 vdd.n2833 10.6151
R21118 vdd.n2835 vdd.n2834 10.6151
R21119 vdd.n2835 vdd.n749 10.6151
R21120 vdd.n2845 vdd.n749 10.6151
R21121 vdd.n2846 vdd.n2845 10.6151
R21122 vdd.n2847 vdd.n2846 10.6151
R21123 vdd.n2847 vdd.n738 10.6151
R21124 vdd.n2857 vdd.n738 10.6151
R21125 vdd.n2858 vdd.n2857 10.6151
R21126 vdd.n2860 vdd.n2858 10.6151
R21127 vdd.n2860 vdd.n2859 10.6151
R21128 vdd.n2871 vdd.n2870 10.6151
R21129 vdd.n2872 vdd.n2871 10.6151
R21130 vdd.n2872 vdd.n713 10.6151
R21131 vdd.n2882 vdd.n713 10.6151
R21132 vdd.n2883 vdd.n2882 10.6151
R21133 vdd.n2884 vdd.n2883 10.6151
R21134 vdd.n2884 vdd.n700 10.6151
R21135 vdd.n2894 vdd.n700 10.6151
R21136 vdd.n2895 vdd.n2894 10.6151
R21137 vdd.n2896 vdd.n2895 10.6151
R21138 vdd.n2896 vdd.n688 10.6151
R21139 vdd.n2906 vdd.n688 10.6151
R21140 vdd.n2907 vdd.n2906 10.6151
R21141 vdd.n2908 vdd.n2907 10.6151
R21142 vdd.n2908 vdd.n677 10.6151
R21143 vdd.n2918 vdd.n677 10.6151
R21144 vdd.n2919 vdd.n2918 10.6151
R21145 vdd.n2965 vdd.n2919 10.6151
R21146 vdd.n2965 vdd.n2964 10.6151
R21147 vdd.n2964 vdd.n2963 10.6151
R21148 vdd.n2963 vdd.n2962 10.6151
R21149 vdd.n2962 vdd.n2960 10.6151
R21150 vdd.n2227 vdd.n960 10.6151
R21151 vdd.n2228 vdd.n2227 10.6151
R21152 vdd.n2229 vdd.n2228 10.6151
R21153 vdd.n2229 vdd.n949 10.6151
R21154 vdd.n2239 vdd.n949 10.6151
R21155 vdd.n2240 vdd.n2239 10.6151
R21156 vdd.n2241 vdd.n2240 10.6151
R21157 vdd.n2241 vdd.n936 10.6151
R21158 vdd.n2251 vdd.n936 10.6151
R21159 vdd.n2252 vdd.n2251 10.6151
R21160 vdd.n2253 vdd.n2252 10.6151
R21161 vdd.n2253 vdd.n925 10.6151
R21162 vdd.n2263 vdd.n925 10.6151
R21163 vdd.n2264 vdd.n2263 10.6151
R21164 vdd.n2265 vdd.n2264 10.6151
R21165 vdd.n2265 vdd.n913 10.6151
R21166 vdd.n2275 vdd.n913 10.6151
R21167 vdd.n2276 vdd.n2275 10.6151
R21168 vdd.n2277 vdd.n2276 10.6151
R21169 vdd.n2277 vdd.n900 10.6151
R21170 vdd.n2287 vdd.n900 10.6151
R21171 vdd.n2288 vdd.n2287 10.6151
R21172 vdd.n2290 vdd.n888 10.6151
R21173 vdd.n2300 vdd.n888 10.6151
R21174 vdd.n2301 vdd.n2300 10.6151
R21175 vdd.n2302 vdd.n2301 10.6151
R21176 vdd.n2302 vdd.n876 10.6151
R21177 vdd.n2312 vdd.n876 10.6151
R21178 vdd.n2313 vdd.n2312 10.6151
R21179 vdd.n2314 vdd.n2313 10.6151
R21180 vdd.n2314 vdd.n865 10.6151
R21181 vdd.n2324 vdd.n865 10.6151
R21182 vdd.n2325 vdd.n2324 10.6151
R21183 vdd.n2326 vdd.n2325 10.6151
R21184 vdd.n2326 vdd.n854 10.6151
R21185 vdd.n2336 vdd.n854 10.6151
R21186 vdd.n2337 vdd.n2336 10.6151
R21187 vdd.n2340 vdd.n2337 10.6151
R21188 vdd.n2340 vdd.n2339 10.6151
R21189 vdd.n2339 vdd.n2338 10.6151
R21190 vdd.n2338 vdd.n837 10.6151
R21191 vdd.n2422 vdd.n837 10.6151
R21192 vdd.n2421 vdd.n2420 10.6151
R21193 vdd.n2420 vdd.n2417 10.6151
R21194 vdd.n2417 vdd.n2416 10.6151
R21195 vdd.n2416 vdd.n2413 10.6151
R21196 vdd.n2413 vdd.n2412 10.6151
R21197 vdd.n2412 vdd.n2409 10.6151
R21198 vdd.n2409 vdd.n2408 10.6151
R21199 vdd.n2408 vdd.n2405 10.6151
R21200 vdd.n2405 vdd.n2404 10.6151
R21201 vdd.n2404 vdd.n2401 10.6151
R21202 vdd.n2401 vdd.n2400 10.6151
R21203 vdd.n2400 vdd.n2397 10.6151
R21204 vdd.n2397 vdd.n2396 10.6151
R21205 vdd.n2396 vdd.n2393 10.6151
R21206 vdd.n2393 vdd.n2392 10.6151
R21207 vdd.n2392 vdd.n2389 10.6151
R21208 vdd.n2389 vdd.n2388 10.6151
R21209 vdd.n2388 vdd.n2385 10.6151
R21210 vdd.n2385 vdd.n2384 10.6151
R21211 vdd.n2384 vdd.n2381 10.6151
R21212 vdd.n2381 vdd.n2380 10.6151
R21213 vdd.n2380 vdd.n2377 10.6151
R21214 vdd.n2377 vdd.n2376 10.6151
R21215 vdd.n2376 vdd.n2373 10.6151
R21216 vdd.n2373 vdd.n2372 10.6151
R21217 vdd.n2372 vdd.n2369 10.6151
R21218 vdd.n2369 vdd.n2368 10.6151
R21219 vdd.n2368 vdd.n2365 10.6151
R21220 vdd.n2365 vdd.n2364 10.6151
R21221 vdd.n2364 vdd.n2361 10.6151
R21222 vdd.n2361 vdd.n2360 10.6151
R21223 vdd.n2357 vdd.n2356 10.6151
R21224 vdd.n2356 vdd.n2354 10.6151
R21225 vdd.n1309 vdd.n1307 10.6151
R21226 vdd.n1307 vdd.n1306 10.6151
R21227 vdd.n1306 vdd.n1304 10.6151
R21228 vdd.n1304 vdd.n1303 10.6151
R21229 vdd.n1303 vdd.n1301 10.6151
R21230 vdd.n1301 vdd.n1300 10.6151
R21231 vdd.n1300 vdd.n1298 10.6151
R21232 vdd.n1298 vdd.n1297 10.6151
R21233 vdd.n1297 vdd.n1295 10.6151
R21234 vdd.n1295 vdd.n1294 10.6151
R21235 vdd.n1294 vdd.n1292 10.6151
R21236 vdd.n1292 vdd.n1291 10.6151
R21237 vdd.n1291 vdd.n1289 10.6151
R21238 vdd.n1289 vdd.n1288 10.6151
R21239 vdd.n1288 vdd.n1286 10.6151
R21240 vdd.n1286 vdd.n1285 10.6151
R21241 vdd.n1285 vdd.n1283 10.6151
R21242 vdd.n1283 vdd.n1282 10.6151
R21243 vdd.n1282 vdd.n1280 10.6151
R21244 vdd.n1280 vdd.n1279 10.6151
R21245 vdd.n1279 vdd.n1277 10.6151
R21246 vdd.n1277 vdd.n1276 10.6151
R21247 vdd.n1276 vdd.n1274 10.6151
R21248 vdd.n1274 vdd.n1273 10.6151
R21249 vdd.n1273 vdd.n1271 10.6151
R21250 vdd.n1271 vdd.n1270 10.6151
R21251 vdd.n1270 vdd.n1268 10.6151
R21252 vdd.n1268 vdd.n1267 10.6151
R21253 vdd.n1267 vdd.n1146 10.6151
R21254 vdd.n1238 vdd.n1146 10.6151
R21255 vdd.n1239 vdd.n1238 10.6151
R21256 vdd.n1241 vdd.n1239 10.6151
R21257 vdd.n1242 vdd.n1241 10.6151
R21258 vdd.n1251 vdd.n1242 10.6151
R21259 vdd.n1251 vdd.n1250 10.6151
R21260 vdd.n1250 vdd.n1249 10.6151
R21261 vdd.n1249 vdd.n1247 10.6151
R21262 vdd.n1247 vdd.n1246 10.6151
R21263 vdd.n1246 vdd.n1244 10.6151
R21264 vdd.n1244 vdd.n1243 10.6151
R21265 vdd.n1243 vdd.n841 10.6151
R21266 vdd.n2352 vdd.n841 10.6151
R21267 vdd.n2353 vdd.n2352 10.6151
R21268 vdd.n1110 vdd.n1109 10.6151
R21269 vdd.n1113 vdd.n1110 10.6151
R21270 vdd.n1114 vdd.n1113 10.6151
R21271 vdd.n1117 vdd.n1114 10.6151
R21272 vdd.n1118 vdd.n1117 10.6151
R21273 vdd.n1121 vdd.n1118 10.6151
R21274 vdd.n1122 vdd.n1121 10.6151
R21275 vdd.n1125 vdd.n1122 10.6151
R21276 vdd.n1126 vdd.n1125 10.6151
R21277 vdd.n1129 vdd.n1126 10.6151
R21278 vdd.n1130 vdd.n1129 10.6151
R21279 vdd.n1133 vdd.n1130 10.6151
R21280 vdd.n1134 vdd.n1133 10.6151
R21281 vdd.n1137 vdd.n1134 10.6151
R21282 vdd.n1138 vdd.n1137 10.6151
R21283 vdd.n1141 vdd.n1138 10.6151
R21284 vdd.n1343 vdd.n1141 10.6151
R21285 vdd.n1343 vdd.n1342 10.6151
R21286 vdd.n1342 vdd.n1340 10.6151
R21287 vdd.n1340 vdd.n1337 10.6151
R21288 vdd.n1337 vdd.n1336 10.6151
R21289 vdd.n1336 vdd.n1333 10.6151
R21290 vdd.n1333 vdd.n1332 10.6151
R21291 vdd.n1332 vdd.n1329 10.6151
R21292 vdd.n1329 vdd.n1328 10.6151
R21293 vdd.n1328 vdd.n1325 10.6151
R21294 vdd.n1325 vdd.n1324 10.6151
R21295 vdd.n1324 vdd.n1321 10.6151
R21296 vdd.n1321 vdd.n1320 10.6151
R21297 vdd.n1320 vdd.n1317 10.6151
R21298 vdd.n1317 vdd.n1316 10.6151
R21299 vdd.n1313 vdd.n1312 10.6151
R21300 vdd.n1312 vdd.n1310 10.6151
R21301 vdd.n1727 vdd.t18 10.5435
R21302 vdd.n2070 vdd.t33 10.5435
R21303 vdd.n3212 vdd.t43 10.5435
R21304 vdd.n3436 vdd.t133 10.5435
R21305 vdd.n292 vdd.n274 10.4732
R21306 vdd.n241 vdd.n223 10.4732
R21307 vdd.n198 vdd.n180 10.4732
R21308 vdd.n147 vdd.n129 10.4732
R21309 vdd.n105 vdd.n87 10.4732
R21310 vdd.n54 vdd.n36 10.4732
R21311 vdd.n1942 vdd.n1924 10.4732
R21312 vdd.n1993 vdd.n1975 10.4732
R21313 vdd.n1848 vdd.n1830 10.4732
R21314 vdd.n1899 vdd.n1881 10.4732
R21315 vdd.n1755 vdd.n1737 10.4732
R21316 vdd.n1806 vdd.n1788 10.4732
R21317 vdd.n2025 vdd.t155 10.3167
R21318 vdd.t100 vdd.n493 10.3167
R21319 vdd.n2187 vdd.n2186 9.98956
R21320 vdd.n3010 vdd.n3009 9.98956
R21321 vdd.n3077 vdd.n3076 9.98956
R21322 vdd.n2079 vdd.n1343 9.98956
R21323 vdd.n1678 vdd.t61 9.86327
R21324 vdd.n3412 vdd.t47 9.86327
R21325 vdd.n2424 vdd.t208 9.7499
R21326 vdd.t193 vdd.n785 9.7499
R21327 vdd.n291 vdd.n276 9.69747
R21328 vdd.n240 vdd.n225 9.69747
R21329 vdd.n197 vdd.n182 9.69747
R21330 vdd.n146 vdd.n131 9.69747
R21331 vdd.n104 vdd.n89 9.69747
R21332 vdd.n53 vdd.n38 9.69747
R21333 vdd.n1941 vdd.n1926 9.69747
R21334 vdd.n1992 vdd.n1977 9.69747
R21335 vdd.n1847 vdd.n1832 9.69747
R21336 vdd.n1898 vdd.n1883 9.69747
R21337 vdd.n1754 vdd.n1739 9.69747
R21338 vdd.n1805 vdd.n1790 9.69747
R21339 vdd.n307 vdd.n306 9.45567
R21340 vdd.n256 vdd.n255 9.45567
R21341 vdd.n213 vdd.n212 9.45567
R21342 vdd.n162 vdd.n161 9.45567
R21343 vdd.n120 vdd.n119 9.45567
R21344 vdd.n69 vdd.n68 9.45567
R21345 vdd.n1957 vdd.n1956 9.45567
R21346 vdd.n2008 vdd.n2007 9.45567
R21347 vdd.n1863 vdd.n1862 9.45567
R21348 vdd.n1914 vdd.n1913 9.45567
R21349 vdd.n1770 vdd.n1769 9.45567
R21350 vdd.n1821 vdd.n1820 9.45567
R21351 vdd.n2149 vdd.n1035 9.3005
R21352 vdd.n2148 vdd.n2147 9.3005
R21353 vdd.n1041 vdd.n1040 9.3005
R21354 vdd.n2142 vdd.n1045 9.3005
R21355 vdd.n2141 vdd.n1046 9.3005
R21356 vdd.n2140 vdd.n1047 9.3005
R21357 vdd.n1051 vdd.n1048 9.3005
R21358 vdd.n2135 vdd.n1052 9.3005
R21359 vdd.n2134 vdd.n1053 9.3005
R21360 vdd.n2133 vdd.n1054 9.3005
R21361 vdd.n1058 vdd.n1055 9.3005
R21362 vdd.n2128 vdd.n1059 9.3005
R21363 vdd.n2127 vdd.n1060 9.3005
R21364 vdd.n2126 vdd.n1061 9.3005
R21365 vdd.n1065 vdd.n1062 9.3005
R21366 vdd.n2121 vdd.n1066 9.3005
R21367 vdd.n2120 vdd.n1067 9.3005
R21368 vdd.n2119 vdd.n1068 9.3005
R21369 vdd.n1072 vdd.n1069 9.3005
R21370 vdd.n2114 vdd.n1073 9.3005
R21371 vdd.n2113 vdd.n1074 9.3005
R21372 vdd.n2112 vdd.n2111 9.3005
R21373 vdd.n2110 vdd.n1075 9.3005
R21374 vdd.n2109 vdd.n2108 9.3005
R21375 vdd.n1081 vdd.n1080 9.3005
R21376 vdd.n2103 vdd.n1085 9.3005
R21377 vdd.n2102 vdd.n1086 9.3005
R21378 vdd.n2101 vdd.n1087 9.3005
R21379 vdd.n1091 vdd.n1088 9.3005
R21380 vdd.n2096 vdd.n1092 9.3005
R21381 vdd.n2095 vdd.n1093 9.3005
R21382 vdd.n2094 vdd.n1094 9.3005
R21383 vdd.n1098 vdd.n1095 9.3005
R21384 vdd.n2089 vdd.n1099 9.3005
R21385 vdd.n2088 vdd.n1100 9.3005
R21386 vdd.n2087 vdd.n1101 9.3005
R21387 vdd.n1105 vdd.n1102 9.3005
R21388 vdd.n2082 vdd.n1106 9.3005
R21389 vdd.n2151 vdd.n2150 9.3005
R21390 vdd.n2173 vdd.n1006 9.3005
R21391 vdd.n2172 vdd.n1014 9.3005
R21392 vdd.n1018 vdd.n1015 9.3005
R21393 vdd.n2167 vdd.n1019 9.3005
R21394 vdd.n2166 vdd.n1020 9.3005
R21395 vdd.n2165 vdd.n1021 9.3005
R21396 vdd.n1025 vdd.n1022 9.3005
R21397 vdd.n2160 vdd.n1026 9.3005
R21398 vdd.n2159 vdd.n1027 9.3005
R21399 vdd.n2158 vdd.n1028 9.3005
R21400 vdd.n1032 vdd.n1029 9.3005
R21401 vdd.n2153 vdd.n1033 9.3005
R21402 vdd.n2152 vdd.n1034 9.3005
R21403 vdd.n2185 vdd.n2184 9.3005
R21404 vdd.n1010 vdd.n1009 9.3005
R21405 vdd.n2013 vdd.n1394 9.3005
R21406 vdd.n2015 vdd.n2014 9.3005
R21407 vdd.n1384 vdd.n1383 9.3005
R21408 vdd.n2029 vdd.n2028 9.3005
R21409 vdd.n2030 vdd.n1382 9.3005
R21410 vdd.n2032 vdd.n2031 9.3005
R21411 vdd.n1373 vdd.n1372 9.3005
R21412 vdd.n2046 vdd.n2045 9.3005
R21413 vdd.n2047 vdd.n1371 9.3005
R21414 vdd.n2049 vdd.n2048 9.3005
R21415 vdd.n1361 vdd.n1360 9.3005
R21416 vdd.n2065 vdd.n2064 9.3005
R21417 vdd.n2066 vdd.n1359 9.3005
R21418 vdd.n2068 vdd.n2067 9.3005
R21419 vdd.n283 vdd.n282 9.3005
R21420 vdd.n278 vdd.n277 9.3005
R21421 vdd.n289 vdd.n288 9.3005
R21422 vdd.n291 vdd.n290 9.3005
R21423 vdd.n274 vdd.n273 9.3005
R21424 vdd.n297 vdd.n296 9.3005
R21425 vdd.n299 vdd.n298 9.3005
R21426 vdd.n271 vdd.n268 9.3005
R21427 vdd.n306 vdd.n305 9.3005
R21428 vdd.n232 vdd.n231 9.3005
R21429 vdd.n227 vdd.n226 9.3005
R21430 vdd.n238 vdd.n237 9.3005
R21431 vdd.n240 vdd.n239 9.3005
R21432 vdd.n223 vdd.n222 9.3005
R21433 vdd.n246 vdd.n245 9.3005
R21434 vdd.n248 vdd.n247 9.3005
R21435 vdd.n220 vdd.n217 9.3005
R21436 vdd.n255 vdd.n254 9.3005
R21437 vdd.n189 vdd.n188 9.3005
R21438 vdd.n184 vdd.n183 9.3005
R21439 vdd.n195 vdd.n194 9.3005
R21440 vdd.n197 vdd.n196 9.3005
R21441 vdd.n180 vdd.n179 9.3005
R21442 vdd.n203 vdd.n202 9.3005
R21443 vdd.n205 vdd.n204 9.3005
R21444 vdd.n177 vdd.n174 9.3005
R21445 vdd.n212 vdd.n211 9.3005
R21446 vdd.n138 vdd.n137 9.3005
R21447 vdd.n133 vdd.n132 9.3005
R21448 vdd.n144 vdd.n143 9.3005
R21449 vdd.n146 vdd.n145 9.3005
R21450 vdd.n129 vdd.n128 9.3005
R21451 vdd.n152 vdd.n151 9.3005
R21452 vdd.n154 vdd.n153 9.3005
R21453 vdd.n126 vdd.n123 9.3005
R21454 vdd.n161 vdd.n160 9.3005
R21455 vdd.n96 vdd.n95 9.3005
R21456 vdd.n91 vdd.n90 9.3005
R21457 vdd.n102 vdd.n101 9.3005
R21458 vdd.n104 vdd.n103 9.3005
R21459 vdd.n87 vdd.n86 9.3005
R21460 vdd.n110 vdd.n109 9.3005
R21461 vdd.n112 vdd.n111 9.3005
R21462 vdd.n84 vdd.n81 9.3005
R21463 vdd.n119 vdd.n118 9.3005
R21464 vdd.n45 vdd.n44 9.3005
R21465 vdd.n40 vdd.n39 9.3005
R21466 vdd.n51 vdd.n50 9.3005
R21467 vdd.n53 vdd.n52 9.3005
R21468 vdd.n36 vdd.n35 9.3005
R21469 vdd.n59 vdd.n58 9.3005
R21470 vdd.n61 vdd.n60 9.3005
R21471 vdd.n33 vdd.n30 9.3005
R21472 vdd.n68 vdd.n67 9.3005
R21473 vdd.n3126 vdd.n3125 9.3005
R21474 vdd.n3127 vdd.n578 9.3005
R21475 vdd.n577 vdd.n575 9.3005
R21476 vdd.n3133 vdd.n574 9.3005
R21477 vdd.n3134 vdd.n573 9.3005
R21478 vdd.n3135 vdd.n572 9.3005
R21479 vdd.n571 vdd.n569 9.3005
R21480 vdd.n3141 vdd.n568 9.3005
R21481 vdd.n3142 vdd.n567 9.3005
R21482 vdd.n3143 vdd.n566 9.3005
R21483 vdd.n565 vdd.n563 9.3005
R21484 vdd.n3149 vdd.n562 9.3005
R21485 vdd.n3150 vdd.n561 9.3005
R21486 vdd.n3151 vdd.n560 9.3005
R21487 vdd.n559 vdd.n557 9.3005
R21488 vdd.n3157 vdd.n556 9.3005
R21489 vdd.n3158 vdd.n555 9.3005
R21490 vdd.n3159 vdd.n554 9.3005
R21491 vdd.n553 vdd.n551 9.3005
R21492 vdd.n3165 vdd.n550 9.3005
R21493 vdd.n3166 vdd.n549 9.3005
R21494 vdd.n3167 vdd.n548 9.3005
R21495 vdd.n547 vdd.n545 9.3005
R21496 vdd.n3173 vdd.n542 9.3005
R21497 vdd.n3174 vdd.n541 9.3005
R21498 vdd.n3175 vdd.n540 9.3005
R21499 vdd.n539 vdd.n537 9.3005
R21500 vdd.n3181 vdd.n536 9.3005
R21501 vdd.n3182 vdd.n535 9.3005
R21502 vdd.n3183 vdd.n534 9.3005
R21503 vdd.n533 vdd.n531 9.3005
R21504 vdd.n3189 vdd.n530 9.3005
R21505 vdd.n3190 vdd.n529 9.3005
R21506 vdd.n3191 vdd.n528 9.3005
R21507 vdd.n527 vdd.n525 9.3005
R21508 vdd.n3196 vdd.n524 9.3005
R21509 vdd.n3206 vdd.n518 9.3005
R21510 vdd.n3208 vdd.n3207 9.3005
R21511 vdd.n509 vdd.n508 9.3005
R21512 vdd.n3223 vdd.n3222 9.3005
R21513 vdd.n3224 vdd.n507 9.3005
R21514 vdd.n3226 vdd.n3225 9.3005
R21515 vdd.n497 vdd.n496 9.3005
R21516 vdd.n3239 vdd.n3238 9.3005
R21517 vdd.n3240 vdd.n495 9.3005
R21518 vdd.n3242 vdd.n3241 9.3005
R21519 vdd.n485 vdd.n484 9.3005
R21520 vdd.n3256 vdd.n3255 9.3005
R21521 vdd.n3257 vdd.n483 9.3005
R21522 vdd.n3259 vdd.n3258 9.3005
R21523 vdd.n312 vdd.n310 9.3005
R21524 vdd.n3210 vdd.n3209 9.3005
R21525 vdd.n3439 vdd.n3438 9.3005
R21526 vdd.n313 vdd.n311 9.3005
R21527 vdd.n3432 vdd.n320 9.3005
R21528 vdd.n3431 vdd.n321 9.3005
R21529 vdd.n3430 vdd.n322 9.3005
R21530 vdd.n331 vdd.n323 9.3005
R21531 vdd.n3424 vdd.n332 9.3005
R21532 vdd.n3423 vdd.n333 9.3005
R21533 vdd.n3422 vdd.n334 9.3005
R21534 vdd.n342 vdd.n335 9.3005
R21535 vdd.n3416 vdd.n343 9.3005
R21536 vdd.n3415 vdd.n344 9.3005
R21537 vdd.n3414 vdd.n345 9.3005
R21538 vdd.n353 vdd.n346 9.3005
R21539 vdd.n3408 vdd.n3407 9.3005
R21540 vdd.n3404 vdd.n354 9.3005
R21541 vdd.n3403 vdd.n357 9.3005
R21542 vdd.n361 vdd.n358 9.3005
R21543 vdd.n362 vdd.n359 9.3005
R21544 vdd.n3396 vdd.n363 9.3005
R21545 vdd.n3395 vdd.n364 9.3005
R21546 vdd.n3394 vdd.n365 9.3005
R21547 vdd.n369 vdd.n366 9.3005
R21548 vdd.n3389 vdd.n370 9.3005
R21549 vdd.n3388 vdd.n371 9.3005
R21550 vdd.n3387 vdd.n372 9.3005
R21551 vdd.n376 vdd.n373 9.3005
R21552 vdd.n3382 vdd.n377 9.3005
R21553 vdd.n3381 vdd.n378 9.3005
R21554 vdd.n3380 vdd.n379 9.3005
R21555 vdd.n383 vdd.n380 9.3005
R21556 vdd.n3375 vdd.n384 9.3005
R21557 vdd.n3374 vdd.n385 9.3005
R21558 vdd.n3373 vdd.n3372 9.3005
R21559 vdd.n3371 vdd.n386 9.3005
R21560 vdd.n3370 vdd.n3369 9.3005
R21561 vdd.n392 vdd.n391 9.3005
R21562 vdd.n3364 vdd.n396 9.3005
R21563 vdd.n3363 vdd.n397 9.3005
R21564 vdd.n3362 vdd.n398 9.3005
R21565 vdd.n402 vdd.n399 9.3005
R21566 vdd.n3357 vdd.n403 9.3005
R21567 vdd.n3356 vdd.n404 9.3005
R21568 vdd.n3355 vdd.n405 9.3005
R21569 vdd.n409 vdd.n406 9.3005
R21570 vdd.n3350 vdd.n410 9.3005
R21571 vdd.n3349 vdd.n411 9.3005
R21572 vdd.n3348 vdd.n412 9.3005
R21573 vdd.n416 vdd.n413 9.3005
R21574 vdd.n3343 vdd.n417 9.3005
R21575 vdd.n3342 vdd.n418 9.3005
R21576 vdd.n3341 vdd.n419 9.3005
R21577 vdd.n423 vdd.n420 9.3005
R21578 vdd.n3336 vdd.n424 9.3005
R21579 vdd.n3335 vdd.n425 9.3005
R21580 vdd.n3334 vdd.n3333 9.3005
R21581 vdd.n3332 vdd.n426 9.3005
R21582 vdd.n3331 vdd.n3330 9.3005
R21583 vdd.n432 vdd.n431 9.3005
R21584 vdd.n3325 vdd.n436 9.3005
R21585 vdd.n3324 vdd.n437 9.3005
R21586 vdd.n3323 vdd.n438 9.3005
R21587 vdd.n442 vdd.n439 9.3005
R21588 vdd.n3318 vdd.n443 9.3005
R21589 vdd.n3317 vdd.n444 9.3005
R21590 vdd.n3316 vdd.n445 9.3005
R21591 vdd.n449 vdd.n446 9.3005
R21592 vdd.n3311 vdd.n450 9.3005
R21593 vdd.n3310 vdd.n451 9.3005
R21594 vdd.n3309 vdd.n452 9.3005
R21595 vdd.n456 vdd.n453 9.3005
R21596 vdd.n3304 vdd.n457 9.3005
R21597 vdd.n3303 vdd.n458 9.3005
R21598 vdd.n3302 vdd.n459 9.3005
R21599 vdd.n463 vdd.n460 9.3005
R21600 vdd.n3297 vdd.n464 9.3005
R21601 vdd.n3296 vdd.n465 9.3005
R21602 vdd.n3292 vdd.n3289 9.3005
R21603 vdd.n3406 vdd.n3405 9.3005
R21604 vdd.n3216 vdd.n513 9.3005
R21605 vdd.n3218 vdd.n3217 9.3005
R21606 vdd.n503 vdd.n502 9.3005
R21607 vdd.n3231 vdd.n3230 9.3005
R21608 vdd.n3232 vdd.n501 9.3005
R21609 vdd.n3234 vdd.n3233 9.3005
R21610 vdd.n490 vdd.n489 9.3005
R21611 vdd.n3247 vdd.n3246 9.3005
R21612 vdd.n3248 vdd.n488 9.3005
R21613 vdd.n3250 vdd.n3249 9.3005
R21614 vdd.n478 vdd.n477 9.3005
R21615 vdd.n3264 vdd.n3263 9.3005
R21616 vdd.n3265 vdd.n476 9.3005
R21617 vdd.n3267 vdd.n3266 9.3005
R21618 vdd.n3268 vdd.n475 9.3005
R21619 vdd.n3270 vdd.n3269 9.3005
R21620 vdd.n3271 vdd.n474 9.3005
R21621 vdd.n3273 vdd.n3272 9.3005
R21622 vdd.n3274 vdd.n472 9.3005
R21623 vdd.n3276 vdd.n3275 9.3005
R21624 vdd.n3277 vdd.n471 9.3005
R21625 vdd.n3279 vdd.n3278 9.3005
R21626 vdd.n3280 vdd.n469 9.3005
R21627 vdd.n3282 vdd.n3281 9.3005
R21628 vdd.n3283 vdd.n468 9.3005
R21629 vdd.n3285 vdd.n3284 9.3005
R21630 vdd.n3286 vdd.n466 9.3005
R21631 vdd.n3288 vdd.n3287 9.3005
R21632 vdd.n3215 vdd.n3214 9.3005
R21633 vdd.n3079 vdd.n514 9.3005
R21634 vdd.n3084 vdd.n3078 9.3005
R21635 vdd.n3094 vdd.n605 9.3005
R21636 vdd.n3095 vdd.n604 9.3005
R21637 vdd.n603 vdd.n601 9.3005
R21638 vdd.n3101 vdd.n600 9.3005
R21639 vdd.n3102 vdd.n599 9.3005
R21640 vdd.n3103 vdd.n598 9.3005
R21641 vdd.n597 vdd.n595 9.3005
R21642 vdd.n3109 vdd.n594 9.3005
R21643 vdd.n3110 vdd.n593 9.3005
R21644 vdd.n3111 vdd.n592 9.3005
R21645 vdd.n591 vdd.n589 9.3005
R21646 vdd.n3116 vdd.n588 9.3005
R21647 vdd.n3117 vdd.n587 9.3005
R21648 vdd.n583 vdd.n582 9.3005
R21649 vdd.n3123 vdd.n3122 9.3005
R21650 vdd.n3124 vdd.n579 9.3005
R21651 vdd.n2078 vdd.n2077 9.3005
R21652 vdd.n2073 vdd.n1345 9.3005
R21653 vdd.n1674 vdd.n1434 9.3005
R21654 vdd.n1676 vdd.n1675 9.3005
R21655 vdd.n1425 vdd.n1424 9.3005
R21656 vdd.n1689 vdd.n1688 9.3005
R21657 vdd.n1690 vdd.n1423 9.3005
R21658 vdd.n1692 vdd.n1691 9.3005
R21659 vdd.n1412 vdd.n1411 9.3005
R21660 vdd.n1705 vdd.n1704 9.3005
R21661 vdd.n1706 vdd.n1410 9.3005
R21662 vdd.n1708 vdd.n1707 9.3005
R21663 vdd.n1401 vdd.n1400 9.3005
R21664 vdd.n1722 vdd.n1721 9.3005
R21665 vdd.n1723 vdd.n1399 9.3005
R21666 vdd.n1725 vdd.n1724 9.3005
R21667 vdd.n1390 vdd.n1389 9.3005
R21668 vdd.n2020 vdd.n2019 9.3005
R21669 vdd.n2021 vdd.n1388 9.3005
R21670 vdd.n2023 vdd.n2022 9.3005
R21671 vdd.n1378 vdd.n1377 9.3005
R21672 vdd.n2037 vdd.n2036 9.3005
R21673 vdd.n2038 vdd.n1376 9.3005
R21674 vdd.n2040 vdd.n2039 9.3005
R21675 vdd.n1368 vdd.n1367 9.3005
R21676 vdd.n2054 vdd.n2053 9.3005
R21677 vdd.n2055 vdd.n1365 9.3005
R21678 vdd.n2059 vdd.n2058 9.3005
R21679 vdd.n2057 vdd.n1366 9.3005
R21680 vdd.n2056 vdd.n1356 9.3005
R21681 vdd.n1673 vdd.n1672 9.3005
R21682 vdd.n1568 vdd.n1558 9.3005
R21683 vdd.n1570 vdd.n1569 9.3005
R21684 vdd.n1571 vdd.n1557 9.3005
R21685 vdd.n1573 vdd.n1572 9.3005
R21686 vdd.n1574 vdd.n1550 9.3005
R21687 vdd.n1576 vdd.n1575 9.3005
R21688 vdd.n1577 vdd.n1549 9.3005
R21689 vdd.n1579 vdd.n1578 9.3005
R21690 vdd.n1580 vdd.n1542 9.3005
R21691 vdd.n1582 vdd.n1581 9.3005
R21692 vdd.n1583 vdd.n1541 9.3005
R21693 vdd.n1585 vdd.n1584 9.3005
R21694 vdd.n1586 vdd.n1534 9.3005
R21695 vdd.n1588 vdd.n1587 9.3005
R21696 vdd.n1589 vdd.n1533 9.3005
R21697 vdd.n1591 vdd.n1590 9.3005
R21698 vdd.n1592 vdd.n1527 9.3005
R21699 vdd.n1594 vdd.n1593 9.3005
R21700 vdd.n1595 vdd.n1525 9.3005
R21701 vdd.n1597 vdd.n1596 9.3005
R21702 vdd.n1526 vdd.n1523 9.3005
R21703 vdd.n1604 vdd.n1519 9.3005
R21704 vdd.n1606 vdd.n1605 9.3005
R21705 vdd.n1607 vdd.n1518 9.3005
R21706 vdd.n1609 vdd.n1608 9.3005
R21707 vdd.n1610 vdd.n1511 9.3005
R21708 vdd.n1612 vdd.n1611 9.3005
R21709 vdd.n1613 vdd.n1510 9.3005
R21710 vdd.n1615 vdd.n1614 9.3005
R21711 vdd.n1616 vdd.n1503 9.3005
R21712 vdd.n1618 vdd.n1617 9.3005
R21713 vdd.n1619 vdd.n1502 9.3005
R21714 vdd.n1621 vdd.n1620 9.3005
R21715 vdd.n1622 vdd.n1495 9.3005
R21716 vdd.n1624 vdd.n1623 9.3005
R21717 vdd.n1625 vdd.n1494 9.3005
R21718 vdd.n1627 vdd.n1626 9.3005
R21719 vdd.n1628 vdd.n1487 9.3005
R21720 vdd.n1630 vdd.n1629 9.3005
R21721 vdd.n1631 vdd.n1486 9.3005
R21722 vdd.n1633 vdd.n1632 9.3005
R21723 vdd.n1634 vdd.n1479 9.3005
R21724 vdd.n1636 vdd.n1635 9.3005
R21725 vdd.n1637 vdd.n1478 9.3005
R21726 vdd.n1639 vdd.n1638 9.3005
R21727 vdd.n1640 vdd.n1469 9.3005
R21728 vdd.n1642 vdd.n1641 9.3005
R21729 vdd.n1643 vdd.n1468 9.3005
R21730 vdd.n1645 vdd.n1644 9.3005
R21731 vdd.n1646 vdd.n1461 9.3005
R21732 vdd.n1648 vdd.n1647 9.3005
R21733 vdd.n1649 vdd.n1460 9.3005
R21734 vdd.n1651 vdd.n1650 9.3005
R21735 vdd.n1652 vdd.n1453 9.3005
R21736 vdd.n1654 vdd.n1653 9.3005
R21737 vdd.n1655 vdd.n1452 9.3005
R21738 vdd.n1657 vdd.n1656 9.3005
R21739 vdd.n1658 vdd.n1445 9.3005
R21740 vdd.n1660 vdd.n1659 9.3005
R21741 vdd.n1661 vdd.n1444 9.3005
R21742 vdd.n1663 vdd.n1662 9.3005
R21743 vdd.n1664 vdd.n1440 9.3005
R21744 vdd.n1666 vdd.n1665 9.3005
R21745 vdd.n1564 vdd.n1435 9.3005
R21746 vdd.n1431 vdd.n1430 9.3005
R21747 vdd.n1681 vdd.n1680 9.3005
R21748 vdd.n1682 vdd.n1429 9.3005
R21749 vdd.n1684 vdd.n1683 9.3005
R21750 vdd.n1419 vdd.n1418 9.3005
R21751 vdd.n1697 vdd.n1696 9.3005
R21752 vdd.n1698 vdd.n1417 9.3005
R21753 vdd.n1700 vdd.n1699 9.3005
R21754 vdd.n1407 vdd.n1406 9.3005
R21755 vdd.n1714 vdd.n1713 9.3005
R21756 vdd.n1715 vdd.n1405 9.3005
R21757 vdd.n1717 vdd.n1716 9.3005
R21758 vdd.n1396 vdd.n1395 9.3005
R21759 vdd.n1668 vdd.n1667 9.3005
R21760 vdd.n2012 vdd.n1729 9.3005
R21761 vdd.n1933 vdd.n1932 9.3005
R21762 vdd.n1928 vdd.n1927 9.3005
R21763 vdd.n1939 vdd.n1938 9.3005
R21764 vdd.n1941 vdd.n1940 9.3005
R21765 vdd.n1924 vdd.n1923 9.3005
R21766 vdd.n1947 vdd.n1946 9.3005
R21767 vdd.n1949 vdd.n1948 9.3005
R21768 vdd.n1921 vdd.n1918 9.3005
R21769 vdd.n1956 vdd.n1955 9.3005
R21770 vdd.n1984 vdd.n1983 9.3005
R21771 vdd.n1979 vdd.n1978 9.3005
R21772 vdd.n1990 vdd.n1989 9.3005
R21773 vdd.n1992 vdd.n1991 9.3005
R21774 vdd.n1975 vdd.n1974 9.3005
R21775 vdd.n1998 vdd.n1997 9.3005
R21776 vdd.n2000 vdd.n1999 9.3005
R21777 vdd.n1972 vdd.n1969 9.3005
R21778 vdd.n2007 vdd.n2006 9.3005
R21779 vdd.n1839 vdd.n1838 9.3005
R21780 vdd.n1834 vdd.n1833 9.3005
R21781 vdd.n1845 vdd.n1844 9.3005
R21782 vdd.n1847 vdd.n1846 9.3005
R21783 vdd.n1830 vdd.n1829 9.3005
R21784 vdd.n1853 vdd.n1852 9.3005
R21785 vdd.n1855 vdd.n1854 9.3005
R21786 vdd.n1827 vdd.n1824 9.3005
R21787 vdd.n1862 vdd.n1861 9.3005
R21788 vdd.n1890 vdd.n1889 9.3005
R21789 vdd.n1885 vdd.n1884 9.3005
R21790 vdd.n1896 vdd.n1895 9.3005
R21791 vdd.n1898 vdd.n1897 9.3005
R21792 vdd.n1881 vdd.n1880 9.3005
R21793 vdd.n1904 vdd.n1903 9.3005
R21794 vdd.n1906 vdd.n1905 9.3005
R21795 vdd.n1878 vdd.n1875 9.3005
R21796 vdd.n1913 vdd.n1912 9.3005
R21797 vdd.n1746 vdd.n1745 9.3005
R21798 vdd.n1741 vdd.n1740 9.3005
R21799 vdd.n1752 vdd.n1751 9.3005
R21800 vdd.n1754 vdd.n1753 9.3005
R21801 vdd.n1737 vdd.n1736 9.3005
R21802 vdd.n1760 vdd.n1759 9.3005
R21803 vdd.n1762 vdd.n1761 9.3005
R21804 vdd.n1734 vdd.n1731 9.3005
R21805 vdd.n1769 vdd.n1768 9.3005
R21806 vdd.n1797 vdd.n1796 9.3005
R21807 vdd.n1792 vdd.n1791 9.3005
R21808 vdd.n1803 vdd.n1802 9.3005
R21809 vdd.n1805 vdd.n1804 9.3005
R21810 vdd.n1788 vdd.n1787 9.3005
R21811 vdd.n1811 vdd.n1810 9.3005
R21812 vdd.n1813 vdd.n1812 9.3005
R21813 vdd.n1785 vdd.n1782 9.3005
R21814 vdd.n1820 vdd.n1819 9.3005
R21815 vdd.n288 vdd.n287 8.92171
R21816 vdd.n237 vdd.n236 8.92171
R21817 vdd.n194 vdd.n193 8.92171
R21818 vdd.n143 vdd.n142 8.92171
R21819 vdd.n101 vdd.n100 8.92171
R21820 vdd.n50 vdd.n49 8.92171
R21821 vdd.n1938 vdd.n1937 8.92171
R21822 vdd.n1989 vdd.n1988 8.92171
R21823 vdd.n1844 vdd.n1843 8.92171
R21824 vdd.n1895 vdd.n1894 8.92171
R21825 vdd.n1751 vdd.n1750 8.92171
R21826 vdd.n1802 vdd.n1801 8.92171
R21827 vdd.n215 vdd.n121 8.81535
R21828 vdd.n1916 vdd.n1822 8.81535
R21829 vdd.n2051 vdd.t14 8.72962
R21830 vdd.n3228 vdd.t2 8.72962
R21831 vdd.t135 vdd.n2025 8.50289
R21832 vdd.n493 vdd.t103 8.50289
R21833 vdd.n28 vdd.n14 8.42249
R21834 vdd.n1727 vdd.t6 8.27616
R21835 vdd.n3436 vdd.t106 8.27616
R21836 vdd.n3440 vdd.n3439 8.16225
R21837 vdd.n2012 vdd.n2011 8.16225
R21838 vdd.n284 vdd.n278 8.14595
R21839 vdd.n233 vdd.n227 8.14595
R21840 vdd.n190 vdd.n184 8.14595
R21841 vdd.n139 vdd.n133 8.14595
R21842 vdd.n97 vdd.n91 8.14595
R21843 vdd.n46 vdd.n40 8.14595
R21844 vdd.n1934 vdd.n1928 8.14595
R21845 vdd.n1985 vdd.n1979 8.14595
R21846 vdd.n1840 vdd.n1834 8.14595
R21847 vdd.n1891 vdd.n1885 8.14595
R21848 vdd.n1747 vdd.n1741 8.14595
R21849 vdd.n1798 vdd.n1792 8.14595
R21850 vdd.t114 vdd.n1415 8.04943
R21851 vdd.n3427 vdd.t12 8.04943
R21852 vdd.n2225 vdd.n962 7.70933
R21853 vdd.n2225 vdd.n965 7.70933
R21854 vdd.n2231 vdd.n951 7.70933
R21855 vdd.n2237 vdd.n951 7.70933
R21856 vdd.n2237 vdd.n944 7.70933
R21857 vdd.n2243 vdd.n944 7.70933
R21858 vdd.n2243 vdd.n947 7.70933
R21859 vdd.n2249 vdd.n940 7.70933
R21860 vdd.n2255 vdd.n934 7.70933
R21861 vdd.n2261 vdd.n921 7.70933
R21862 vdd.n2267 vdd.n921 7.70933
R21863 vdd.n2273 vdd.n915 7.70933
R21864 vdd.n2279 vdd.n908 7.70933
R21865 vdd.n2279 vdd.n911 7.70933
R21866 vdd.n2285 vdd.n904 7.70933
R21867 vdd.n2292 vdd.n890 7.70933
R21868 vdd.n2298 vdd.n890 7.70933
R21869 vdd.n2304 vdd.n884 7.70933
R21870 vdd.n2310 vdd.n880 7.70933
R21871 vdd.n2316 vdd.n874 7.70933
R21872 vdd.n2334 vdd.n856 7.70933
R21873 vdd.n2334 vdd.n849 7.70933
R21874 vdd.n2342 vdd.n849 7.70933
R21875 vdd.n2424 vdd.n833 7.70933
R21876 vdd.n2807 vdd.n785 7.70933
R21877 vdd.n2819 vdd.n774 7.70933
R21878 vdd.n2819 vdd.n768 7.70933
R21879 vdd.n2825 vdd.n768 7.70933
R21880 vdd.n2837 vdd.n759 7.70933
R21881 vdd.n2843 vdd.n753 7.70933
R21882 vdd.n2855 vdd.n740 7.70933
R21883 vdd.n2862 vdd.n733 7.70933
R21884 vdd.n2862 vdd.n736 7.70933
R21885 vdd.n2868 vdd.n729 7.70933
R21886 vdd.n2874 vdd.n715 7.70933
R21887 vdd.n2880 vdd.n715 7.70933
R21888 vdd.n2886 vdd.n709 7.70933
R21889 vdd.n2892 vdd.n702 7.70933
R21890 vdd.n2892 vdd.n705 7.70933
R21891 vdd.n2898 vdd.n698 7.70933
R21892 vdd.n2904 vdd.n692 7.70933
R21893 vdd.n2910 vdd.n679 7.70933
R21894 vdd.n2916 vdd.n679 7.70933
R21895 vdd.n2916 vdd.n671 7.70933
R21896 vdd.n2967 vdd.n671 7.70933
R21897 vdd.n2967 vdd.n674 7.70933
R21898 vdd.n2973 vdd.n631 7.70933
R21899 vdd.n3043 vdd.n631 7.70933
R21900 vdd.n283 vdd.n280 7.3702
R21901 vdd.n232 vdd.n229 7.3702
R21902 vdd.n189 vdd.n186 7.3702
R21903 vdd.n138 vdd.n135 7.3702
R21904 vdd.n96 vdd.n93 7.3702
R21905 vdd.n45 vdd.n42 7.3702
R21906 vdd.n1933 vdd.n1930 7.3702
R21907 vdd.n1984 vdd.n1981 7.3702
R21908 vdd.n1839 vdd.n1836 7.3702
R21909 vdd.n1890 vdd.n1887 7.3702
R21910 vdd.n1746 vdd.n1743 7.3702
R21911 vdd.n1797 vdd.n1794 7.3702
R21912 vdd.n934 vdd.t213 7.36923
R21913 vdd.n2898 vdd.t190 7.36923
R21914 vdd.n1694 vdd.t8 7.1425
R21915 vdd.n2249 vdd.t167 7.1425
R21916 vdd.n1253 vdd.t161 7.1425
R21917 vdd.n2831 vdd.t166 7.1425
R21918 vdd.n692 vdd.t176 7.1425
R21919 vdd.n3420 vdd.t122 7.1425
R21920 vdd.n1605 vdd.n1604 6.98232
R21921 vdd.n2113 vdd.n2112 6.98232
R21922 vdd.n3335 vdd.n3334 6.98232
R21923 vdd.n3127 vdd.n3126 6.98232
R21924 vdd.n1710 vdd.t137 6.91577
R21925 vdd.n325 vdd.t139 6.91577
R21926 vdd.n1253 vdd.t162 6.80241
R21927 vdd.n2831 vdd.t206 6.80241
R21928 vdd.n2017 vdd.t10 6.68904
R21929 vdd.n3261 vdd.t110 6.68904
R21930 vdd.n1380 vdd.t20 6.46231
R21931 vdd.n2273 vdd.t174 6.46231
R21932 vdd.t177 vdd.n884 6.46231
R21933 vdd.n2855 vdd.t182 6.46231
R21934 vdd.t198 vdd.n709 6.46231
R21935 vdd.t0 vdd.n492 6.46231
R21936 vdd.n2349 vdd.t210 6.34895
R21937 vdd.n2728 vdd.t195 6.34895
R21938 vdd.n3440 vdd.n309 6.27748
R21939 vdd.n2011 vdd.n2010 6.27748
R21940 vdd.n2870 vdd.n725 6.2444
R21941 vdd.n2289 vdd.n2288 6.2444
R21942 vdd.n2310 vdd.t203 5.89549
R21943 vdd.n753 vdd.t178 5.89549
R21944 vdd.n284 vdd.n283 5.81868
R21945 vdd.n233 vdd.n232 5.81868
R21946 vdd.n190 vdd.n189 5.81868
R21947 vdd.n139 vdd.n138 5.81868
R21948 vdd.n97 vdd.n96 5.81868
R21949 vdd.n46 vdd.n45 5.81868
R21950 vdd.n1934 vdd.n1933 5.81868
R21951 vdd.n1985 vdd.n1984 5.81868
R21952 vdd.n1840 vdd.n1839 5.81868
R21953 vdd.n1891 vdd.n1890 5.81868
R21954 vdd.n1747 vdd.n1746 5.81868
R21955 vdd.n1798 vdd.n1797 5.81868
R21956 vdd.n2432 vdd.n2431 5.77611
R21957 vdd.n1177 vdd.n1176 5.77611
R21958 vdd.n2740 vdd.n2739 5.77611
R21959 vdd.n2982 vdd.n663 5.77611
R21960 vdd.n3048 vdd.n627 5.77611
R21961 vdd.n2603 vdd.n2537 5.77611
R21962 vdd.n2357 vdd.n840 5.77611
R21963 vdd.n1313 vdd.n1145 5.77611
R21964 vdd.n1567 vdd.n1564 5.62474
R21965 vdd.n2076 vdd.n2073 5.62474
R21966 vdd.n3295 vdd.n3292 5.62474
R21967 vdd.n3082 vdd.n3079 5.62474
R21968 vdd.n2285 vdd.t192 5.55539
R21969 vdd.n729 vdd.t170 5.55539
R21970 vdd.n287 vdd.n278 5.04292
R21971 vdd.n236 vdd.n227 5.04292
R21972 vdd.n193 vdd.n184 5.04292
R21973 vdd.n142 vdd.n133 5.04292
R21974 vdd.n100 vdd.n91 5.04292
R21975 vdd.n49 vdd.n40 5.04292
R21976 vdd.n1937 vdd.n1928 5.04292
R21977 vdd.n1988 vdd.n1979 5.04292
R21978 vdd.n1843 vdd.n1834 5.04292
R21979 vdd.n1894 vdd.n1885 5.04292
R21980 vdd.n1750 vdd.n1741 5.04292
R21981 vdd.n1801 vdd.n1792 5.04292
R21982 vdd.n2043 vdd.t20 4.8752
R21983 vdd.t173 vdd.t183 4.8752
R21984 vdd.t214 vdd.t160 4.8752
R21985 vdd.n3236 vdd.t0 4.8752
R21986 vdd.n2433 vdd.n2432 4.83952
R21987 vdd.n1176 vdd.n1175 4.83952
R21988 vdd.n2741 vdd.n2740 4.83952
R21989 vdd.n663 vdd.n658 4.83952
R21990 vdd.n627 vdd.n622 4.83952
R21991 vdd.n2600 vdd.n2537 4.83952
R21992 vdd.n2360 vdd.n840 4.83952
R21993 vdd.n1316 vdd.n1145 4.83952
R21994 vdd.n1227 vdd.t180 4.76184
R21995 vdd.n2813 vdd.t168 4.76184
R21996 vdd.n2081 vdd.n2080 4.74817
R21997 vdd.n1349 vdd.n1344 4.74817
R21998 vdd.n1011 vdd.n1008 4.74817
R21999 vdd.n2174 vdd.n1007 4.74817
R22000 vdd.n2179 vdd.n1008 4.74817
R22001 vdd.n2178 vdd.n1007 4.74817
R22002 vdd.n521 vdd.n519 4.74817
R22003 vdd.n3197 vdd.n522 4.74817
R22004 vdd.n3200 vdd.n522 4.74817
R22005 vdd.n3201 vdd.n521 4.74817
R22006 vdd.n3089 vdd.n606 4.74817
R22007 vdd.n3085 vdd.n608 4.74817
R22008 vdd.n3088 vdd.n608 4.74817
R22009 vdd.n3093 vdd.n606 4.74817
R22010 vdd.n2080 vdd.n1107 4.74817
R22011 vdd.n1346 vdd.n1344 4.74817
R22012 vdd.n309 vdd.n308 4.7074
R22013 vdd.n215 vdd.n214 4.7074
R22014 vdd.n2010 vdd.n2009 4.7074
R22015 vdd.n1916 vdd.n1915 4.7074
R22016 vdd.t10 vdd.n1386 4.64847
R22017 vdd.t175 vdd.n915 4.64847
R22018 vdd.n2304 vdd.t212 4.64847
R22019 vdd.t201 vdd.n740 4.64847
R22020 vdd.n2886 vdd.t197 4.64847
R22021 vdd.n3252 vdd.t110 4.64847
R22022 vdd.n904 vdd.t88 4.53511
R22023 vdd.n2868 vdd.t51 4.53511
R22024 vdd.n1719 vdd.t137 4.42174
R22025 vdd.n2231 vdd.t29 4.42174
R22026 vdd.n1227 vdd.t74 4.42174
R22027 vdd.n2813 vdd.t81 4.42174
R22028 vdd.n674 vdd.t25 4.42174
R22029 vdd.n3434 vdd.t139 4.42174
R22030 vdd.n2859 vdd.n725 4.37123
R22031 vdd.n2290 vdd.n2289 4.37123
R22032 vdd.n2328 vdd.t199 4.30838
R22033 vdd.n2716 vdd.t186 4.30838
R22034 vdd.n288 vdd.n276 4.26717
R22035 vdd.n237 vdd.n225 4.26717
R22036 vdd.n194 vdd.n182 4.26717
R22037 vdd.n143 vdd.n131 4.26717
R22038 vdd.n101 vdd.n89 4.26717
R22039 vdd.n50 vdd.n38 4.26717
R22040 vdd.n1938 vdd.n1926 4.26717
R22041 vdd.n1989 vdd.n1977 4.26717
R22042 vdd.n1844 vdd.n1832 4.26717
R22043 vdd.n1895 vdd.n1883 4.26717
R22044 vdd.n1751 vdd.n1739 4.26717
R22045 vdd.n1802 vdd.n1790 4.26717
R22046 vdd.t8 vdd.n1414 4.19501
R22047 vdd.t122 vdd.n329 4.19501
R22048 vdd.n309 vdd.n215 4.10845
R22049 vdd.n2010 vdd.n1916 4.10845
R22050 vdd.n265 vdd.t130 4.06363
R22051 vdd.n265 vdd.t158 4.06363
R22052 vdd.n263 vdd.t148 4.06363
R22053 vdd.n263 vdd.t225 4.06363
R22054 vdd.n261 vdd.t238 4.06363
R22055 vdd.n261 vdd.t119 4.06363
R22056 vdd.n259 vdd.t112 4.06363
R22057 vdd.n259 vdd.t151 4.06363
R22058 vdd.n257 vdd.t1 4.06363
R22059 vdd.n257 vdd.t101 4.06363
R22060 vdd.n171 vdd.t13 4.06363
R22061 vdd.n171 vdd.t123 4.06363
R22062 vdd.n169 vdd.t233 4.06363
R22063 vdd.n169 vdd.t150 4.06363
R22064 vdd.n167 vdd.t134 4.06363
R22065 vdd.n167 vdd.t107 4.06363
R22066 vdd.n165 vdd.t104 4.06363
R22067 vdd.n165 vdd.t111 4.06363
R22068 vdd.n163 vdd.t218 4.06363
R22069 vdd.n163 vdd.t143 4.06363
R22070 vdd.n78 vdd.t17 4.06363
R22071 vdd.n78 vdd.t232 4.06363
R22072 vdd.n76 vdd.t140 4.06363
R22073 vdd.n76 vdd.t129 4.06363
R22074 vdd.n74 vdd.t239 4.06363
R22075 vdd.n74 vdd.t149 4.06363
R22076 vdd.n72 vdd.t236 4.06363
R22077 vdd.n72 vdd.t223 4.06363
R22078 vdd.n70 vdd.t241 4.06363
R22079 vdd.n70 vdd.t217 4.06363
R22080 vdd.n1958 vdd.t156 4.06363
R22081 vdd.n1958 vdd.t157 4.06363
R22082 vdd.n1960 vdd.t11 4.06363
R22083 vdd.n1960 vdd.t145 4.06363
R22084 vdd.n1962 vdd.t226 4.06363
R22085 vdd.n1962 vdd.t118 4.06363
R22086 vdd.n1964 vdd.t109 4.06363
R22087 vdd.n1964 vdd.t146 4.06363
R22088 vdd.n1966 vdd.t237 4.06363
R22089 vdd.n1966 vdd.t159 4.06363
R22090 vdd.n1864 vdd.t243 4.06363
R22091 vdd.n1864 vdd.t113 4.06363
R22092 vdd.n1866 vdd.t229 4.06363
R22093 vdd.n1866 vdd.t136 4.06363
R22094 vdd.n1868 vdd.t7 4.06363
R22095 vdd.n1868 vdd.t19 4.06363
R22096 vdd.n1870 vdd.t221 4.06363
R22097 vdd.n1870 vdd.t224 4.06363
R22098 vdd.n1872 vdd.t9 4.06363
R22099 vdd.n1872 vdd.t124 4.06363
R22100 vdd.n1771 vdd.t216 4.06363
R22101 vdd.n1771 vdd.t21 4.06363
R22102 vdd.n1773 vdd.t222 4.06363
R22103 vdd.n1773 vdd.t227 4.06363
R22104 vdd.n1775 vdd.t242 4.06363
R22105 vdd.n1775 vdd.t228 4.06363
R22106 vdd.n1777 vdd.t127 4.06363
R22107 vdd.n1777 vdd.t138 4.06363
R22108 vdd.n1779 vdd.t105 4.06363
R22109 vdd.n1779 vdd.t115 4.06363
R22110 vdd.n940 vdd.t205 3.96828
R22111 vdd.n2322 vdd.t185 3.96828
R22112 vdd.n2710 vdd.t202 3.96828
R22113 vdd.n2904 vdd.t191 3.96828
R22114 vdd.n26 vdd.t152 3.9605
R22115 vdd.n26 vdd.t121 3.9605
R22116 vdd.n23 vdd.t125 3.9605
R22117 vdd.n23 vdd.t116 3.9605
R22118 vdd.n21 vdd.t120 3.9605
R22119 vdd.n21 vdd.t231 3.9605
R22120 vdd.n20 vdd.t117 3.9605
R22121 vdd.n20 vdd.t5 3.9605
R22122 vdd.n15 vdd.t126 3.9605
R22123 vdd.n15 vdd.t141 3.9605
R22124 vdd.n16 vdd.t235 3.9605
R22125 vdd.n16 vdd.t4 3.9605
R22126 vdd.n18 vdd.t234 3.9605
R22127 vdd.n18 vdd.t142 3.9605
R22128 vdd.n25 vdd.t147 3.9605
R22129 vdd.n25 vdd.t230 3.9605
R22130 vdd.n2255 vdd.t205 3.74155
R22131 vdd.n874 vdd.t185 3.74155
R22132 vdd.n2837 vdd.t202 3.74155
R22133 vdd.n698 vdd.t191 3.74155
R22134 vdd.n7 vdd.t215 3.61217
R22135 vdd.n7 vdd.t179 3.61217
R22136 vdd.n8 vdd.t187 3.61217
R22137 vdd.n8 vdd.t207 3.61217
R22138 vdd.n10 vdd.t196 3.61217
R22139 vdd.n10 vdd.t169 3.61217
R22140 vdd.n12 vdd.t165 3.61217
R22141 vdd.n12 vdd.t194 3.61217
R22142 vdd.n5 vdd.t209 3.61217
R22143 vdd.n5 vdd.t189 3.61217
R22144 vdd.n3 vdd.t181 3.61217
R22145 vdd.n3 vdd.t211 3.61217
R22146 vdd.n1 vdd.t163 3.61217
R22147 vdd.n1 vdd.t200 3.61217
R22148 vdd.n0 vdd.t204 3.61217
R22149 vdd.n0 vdd.t184 3.61217
R22150 vdd.n292 vdd.n291 3.49141
R22151 vdd.n241 vdd.n240 3.49141
R22152 vdd.n198 vdd.n197 3.49141
R22153 vdd.n147 vdd.n146 3.49141
R22154 vdd.n105 vdd.n104 3.49141
R22155 vdd.n54 vdd.n53 3.49141
R22156 vdd.n1942 vdd.n1941 3.49141
R22157 vdd.n1993 vdd.n1992 3.49141
R22158 vdd.n1848 vdd.n1847 3.49141
R22159 vdd.n1899 vdd.n1898 3.49141
R22160 vdd.n1755 vdd.n1754 3.49141
R22161 vdd.n1806 vdd.n1805 3.49141
R22162 vdd.t199 vdd.n856 3.40145
R22163 vdd.n2496 vdd.t208 3.40145
R22164 vdd.n2800 vdd.t193 3.40145
R22165 vdd.n2825 vdd.t186 3.40145
R22166 vdd.n1702 vdd.t114 3.28809
R22167 vdd.n965 vdd.t29 3.28809
R22168 vdd.n2349 vdd.t74 3.28809
R22169 vdd.n2728 vdd.t81 3.28809
R22170 vdd.n2973 vdd.t25 3.28809
R22171 vdd.t12 vdd.n3426 3.28809
R22172 vdd.n1403 vdd.t6 3.06136
R22173 vdd.n2267 vdd.t175 3.06136
R22174 vdd.n1265 vdd.t212 3.06136
R22175 vdd.n2849 vdd.t201 3.06136
R22176 vdd.t197 vdd.n702 3.06136
R22177 vdd.t106 vdd.n3435 3.06136
R22178 vdd.n2342 vdd.t180 2.94799
R22179 vdd.t168 vdd.n774 2.94799
R22180 vdd.n2026 vdd.t135 2.83463
R22181 vdd.n3253 vdd.t103 2.83463
R22182 vdd.n295 vdd.n274 2.71565
R22183 vdd.n244 vdd.n223 2.71565
R22184 vdd.n201 vdd.n180 2.71565
R22185 vdd.n150 vdd.n129 2.71565
R22186 vdd.n108 vdd.n87 2.71565
R22187 vdd.n57 vdd.n36 2.71565
R22188 vdd.n1945 vdd.n1924 2.71565
R22189 vdd.n1996 vdd.n1975 2.71565
R22190 vdd.n1851 vdd.n1830 2.71565
R22191 vdd.n1902 vdd.n1881 2.71565
R22192 vdd.n1758 vdd.n1737 2.71565
R22193 vdd.n1809 vdd.n1788 2.71565
R22194 vdd.n2042 vdd.t14 2.6079
R22195 vdd.t2 vdd.n499 2.6079
R22196 vdd.n2316 vdd.t183 2.49453
R22197 vdd.n759 vdd.t214 2.49453
R22198 vdd.n282 vdd.n281 2.4129
R22199 vdd.n231 vdd.n230 2.4129
R22200 vdd.n188 vdd.n187 2.4129
R22201 vdd.n137 vdd.n136 2.4129
R22202 vdd.n95 vdd.n94 2.4129
R22203 vdd.n44 vdd.n43 2.4129
R22204 vdd.n1932 vdd.n1931 2.4129
R22205 vdd.n1983 vdd.n1982 2.4129
R22206 vdd.n1838 vdd.n1837 2.4129
R22207 vdd.n1889 vdd.n1888 2.4129
R22208 vdd.n1745 vdd.n1744 2.4129
R22209 vdd.n1796 vdd.n1795 2.4129
R22210 vdd.n2186 vdd.n1008 2.27742
R22211 vdd.n2186 vdd.n1007 2.27742
R22212 vdd.n3009 vdd.n522 2.27742
R22213 vdd.n3009 vdd.n521 2.27742
R22214 vdd.n3077 vdd.n608 2.27742
R22215 vdd.n3077 vdd.n606 2.27742
R22216 vdd.n2080 vdd.n2079 2.27742
R22217 vdd.n2079 vdd.n1344 2.27742
R22218 vdd.n911 vdd.t192 2.15444
R22219 vdd.n2292 vdd.t172 2.15444
R22220 vdd.n736 vdd.t171 2.15444
R22221 vdd.n2874 vdd.t170 2.15444
R22222 vdd.n296 vdd.n272 1.93989
R22223 vdd.n245 vdd.n221 1.93989
R22224 vdd.n202 vdd.n178 1.93989
R22225 vdd.n151 vdd.n127 1.93989
R22226 vdd.n109 vdd.n85 1.93989
R22227 vdd.n58 vdd.n34 1.93989
R22228 vdd.n1946 vdd.n1922 1.93989
R22229 vdd.n1997 vdd.n1973 1.93989
R22230 vdd.n1852 vdd.n1828 1.93989
R22231 vdd.n1903 vdd.n1879 1.93989
R22232 vdd.n1759 vdd.n1735 1.93989
R22233 vdd.n1810 vdd.n1786 1.93989
R22234 vdd.n1265 vdd.t203 1.81434
R22235 vdd.n2849 vdd.t178 1.81434
R22236 vdd.n1438 vdd.t61 1.47425
R22237 vdd.t47 vdd.n3411 1.47425
R22238 vdd.t210 vdd.n833 1.36088
R22239 vdd.n2807 vdd.t195 1.36088
R22240 vdd.t174 vdd.n908 1.24752
R22241 vdd.n2298 vdd.t177 1.24752
R22242 vdd.t182 vdd.n733 1.24752
R22243 vdd.n2880 vdd.t198 1.24752
R22244 vdd.n307 vdd.n267 1.16414
R22245 vdd.n300 vdd.n299 1.16414
R22246 vdd.n256 vdd.n216 1.16414
R22247 vdd.n249 vdd.n248 1.16414
R22248 vdd.n213 vdd.n173 1.16414
R22249 vdd.n206 vdd.n205 1.16414
R22250 vdd.n162 vdd.n122 1.16414
R22251 vdd.n155 vdd.n154 1.16414
R22252 vdd.n120 vdd.n80 1.16414
R22253 vdd.n113 vdd.n112 1.16414
R22254 vdd.n69 vdd.n29 1.16414
R22255 vdd.n62 vdd.n61 1.16414
R22256 vdd.n1957 vdd.n1917 1.16414
R22257 vdd.n1950 vdd.n1949 1.16414
R22258 vdd.n2008 vdd.n1968 1.16414
R22259 vdd.n2001 vdd.n2000 1.16414
R22260 vdd.n1863 vdd.n1823 1.16414
R22261 vdd.n1856 vdd.n1855 1.16414
R22262 vdd.n1914 vdd.n1874 1.16414
R22263 vdd.n1907 vdd.n1906 1.16414
R22264 vdd.n1770 vdd.n1730 1.16414
R22265 vdd.n1763 vdd.n1762 1.16414
R22266 vdd.n1821 vdd.n1781 1.16414
R22267 vdd.n1814 vdd.n1813 1.16414
R22268 vdd.n2011 vdd.n28 1.11236
R22269 vdd vdd.n3440 1.10453
R22270 vdd.n2034 vdd.t155 1.02079
R22271 vdd.t88 vdd.t172 1.02079
R22272 vdd.t171 vdd.t51 1.02079
R22273 vdd.n3244 vdd.t100 1.02079
R22274 vdd.n1568 vdd.n1567 0.970197
R22275 vdd.n2077 vdd.n2076 0.970197
R22276 vdd.n3296 vdd.n3295 0.970197
R22277 vdd.n3084 vdd.n3082 0.970197
R22278 vdd.n2322 vdd.t162 0.907421
R22279 vdd.n2710 vdd.t206 0.907421
R22280 vdd.t18 vdd.n1392 0.794056
R22281 vdd.n2061 vdd.t33 0.794056
R22282 vdd.t43 vdd.n511 0.794056
R22283 vdd.n481 vdd.t133 0.794056
R22284 vdd.n1711 vdd.t108 0.567326
R22285 vdd.n947 vdd.t167 0.567326
R22286 vdd.n2328 vdd.t161 0.567326
R22287 vdd.n2716 vdd.t166 0.567326
R22288 vdd.n2910 vdd.t176 0.567326
R22289 vdd.n3428 vdd.t128 0.567326
R22290 vdd.n2067 vdd.n1009 0.509646
R22291 vdd.n3209 vdd.n3208 0.509646
R22292 vdd.n3407 vdd.n3406 0.509646
R22293 vdd.n3289 vdd.n3288 0.509646
R22294 vdd.n3215 vdd.n514 0.509646
R22295 vdd.n2056 vdd.n1345 0.509646
R22296 vdd.n1673 vdd.n1435 0.509646
R22297 vdd.n1667 vdd.n1666 0.509646
R22298 vdd.n4 vdd.n2 0.459552
R22299 vdd.n11 vdd.n9 0.459552
R22300 vdd.n305 vdd.n304 0.388379
R22301 vdd.n271 vdd.n269 0.388379
R22302 vdd.n254 vdd.n253 0.388379
R22303 vdd.n220 vdd.n218 0.388379
R22304 vdd.n211 vdd.n210 0.388379
R22305 vdd.n177 vdd.n175 0.388379
R22306 vdd.n160 vdd.n159 0.388379
R22307 vdd.n126 vdd.n124 0.388379
R22308 vdd.n118 vdd.n117 0.388379
R22309 vdd.n84 vdd.n82 0.388379
R22310 vdd.n67 vdd.n66 0.388379
R22311 vdd.n33 vdd.n31 0.388379
R22312 vdd.n1955 vdd.n1954 0.388379
R22313 vdd.n1921 vdd.n1919 0.388379
R22314 vdd.n2006 vdd.n2005 0.388379
R22315 vdd.n1972 vdd.n1970 0.388379
R22316 vdd.n1861 vdd.n1860 0.388379
R22317 vdd.n1827 vdd.n1825 0.388379
R22318 vdd.n1912 vdd.n1911 0.388379
R22319 vdd.n1878 vdd.n1876 0.388379
R22320 vdd.n1768 vdd.n1767 0.388379
R22321 vdd.n1734 vdd.n1732 0.388379
R22322 vdd.n1819 vdd.n1818 0.388379
R22323 vdd.n1785 vdd.n1783 0.388379
R22324 vdd.n19 vdd.n17 0.387128
R22325 vdd.n24 vdd.n22 0.387128
R22326 vdd.n6 vdd.n4 0.358259
R22327 vdd.n13 vdd.n11 0.358259
R22328 vdd.n260 vdd.n258 0.358259
R22329 vdd.n262 vdd.n260 0.358259
R22330 vdd.n264 vdd.n262 0.358259
R22331 vdd.n266 vdd.n264 0.358259
R22332 vdd.n308 vdd.n266 0.358259
R22333 vdd.n166 vdd.n164 0.358259
R22334 vdd.n168 vdd.n166 0.358259
R22335 vdd.n170 vdd.n168 0.358259
R22336 vdd.n172 vdd.n170 0.358259
R22337 vdd.n214 vdd.n172 0.358259
R22338 vdd.n73 vdd.n71 0.358259
R22339 vdd.n75 vdd.n73 0.358259
R22340 vdd.n77 vdd.n75 0.358259
R22341 vdd.n79 vdd.n77 0.358259
R22342 vdd.n121 vdd.n79 0.358259
R22343 vdd.n2009 vdd.n1967 0.358259
R22344 vdd.n1967 vdd.n1965 0.358259
R22345 vdd.n1965 vdd.n1963 0.358259
R22346 vdd.n1963 vdd.n1961 0.358259
R22347 vdd.n1961 vdd.n1959 0.358259
R22348 vdd.n1915 vdd.n1873 0.358259
R22349 vdd.n1873 vdd.n1871 0.358259
R22350 vdd.n1871 vdd.n1869 0.358259
R22351 vdd.n1869 vdd.n1867 0.358259
R22352 vdd.n1867 vdd.n1865 0.358259
R22353 vdd.n1822 vdd.n1780 0.358259
R22354 vdd.n1780 vdd.n1778 0.358259
R22355 vdd.n1778 vdd.n1776 0.358259
R22356 vdd.n1776 vdd.n1774 0.358259
R22357 vdd.n1774 vdd.n1772 0.358259
R22358 vdd.t131 vdd.n1421 0.340595
R22359 vdd.n2261 vdd.t213 0.340595
R22360 vdd.n880 vdd.t173 0.340595
R22361 vdd.n2843 vdd.t160 0.340595
R22362 vdd.n705 vdd.t190 0.340595
R22363 vdd.n3419 vdd.t22 0.340595
R22364 vdd.n14 vdd.n6 0.334552
R22365 vdd.n14 vdd.n13 0.334552
R22366 vdd.n27 vdd.n19 0.21707
R22367 vdd.n27 vdd.n24 0.21707
R22368 vdd.n306 vdd.n268 0.155672
R22369 vdd.n298 vdd.n268 0.155672
R22370 vdd.n298 vdd.n297 0.155672
R22371 vdd.n297 vdd.n273 0.155672
R22372 vdd.n290 vdd.n273 0.155672
R22373 vdd.n290 vdd.n289 0.155672
R22374 vdd.n289 vdd.n277 0.155672
R22375 vdd.n282 vdd.n277 0.155672
R22376 vdd.n255 vdd.n217 0.155672
R22377 vdd.n247 vdd.n217 0.155672
R22378 vdd.n247 vdd.n246 0.155672
R22379 vdd.n246 vdd.n222 0.155672
R22380 vdd.n239 vdd.n222 0.155672
R22381 vdd.n239 vdd.n238 0.155672
R22382 vdd.n238 vdd.n226 0.155672
R22383 vdd.n231 vdd.n226 0.155672
R22384 vdd.n212 vdd.n174 0.155672
R22385 vdd.n204 vdd.n174 0.155672
R22386 vdd.n204 vdd.n203 0.155672
R22387 vdd.n203 vdd.n179 0.155672
R22388 vdd.n196 vdd.n179 0.155672
R22389 vdd.n196 vdd.n195 0.155672
R22390 vdd.n195 vdd.n183 0.155672
R22391 vdd.n188 vdd.n183 0.155672
R22392 vdd.n161 vdd.n123 0.155672
R22393 vdd.n153 vdd.n123 0.155672
R22394 vdd.n153 vdd.n152 0.155672
R22395 vdd.n152 vdd.n128 0.155672
R22396 vdd.n145 vdd.n128 0.155672
R22397 vdd.n145 vdd.n144 0.155672
R22398 vdd.n144 vdd.n132 0.155672
R22399 vdd.n137 vdd.n132 0.155672
R22400 vdd.n119 vdd.n81 0.155672
R22401 vdd.n111 vdd.n81 0.155672
R22402 vdd.n111 vdd.n110 0.155672
R22403 vdd.n110 vdd.n86 0.155672
R22404 vdd.n103 vdd.n86 0.155672
R22405 vdd.n103 vdd.n102 0.155672
R22406 vdd.n102 vdd.n90 0.155672
R22407 vdd.n95 vdd.n90 0.155672
R22408 vdd.n68 vdd.n30 0.155672
R22409 vdd.n60 vdd.n30 0.155672
R22410 vdd.n60 vdd.n59 0.155672
R22411 vdd.n59 vdd.n35 0.155672
R22412 vdd.n52 vdd.n35 0.155672
R22413 vdd.n52 vdd.n51 0.155672
R22414 vdd.n51 vdd.n39 0.155672
R22415 vdd.n44 vdd.n39 0.155672
R22416 vdd.n1956 vdd.n1918 0.155672
R22417 vdd.n1948 vdd.n1918 0.155672
R22418 vdd.n1948 vdd.n1947 0.155672
R22419 vdd.n1947 vdd.n1923 0.155672
R22420 vdd.n1940 vdd.n1923 0.155672
R22421 vdd.n1940 vdd.n1939 0.155672
R22422 vdd.n1939 vdd.n1927 0.155672
R22423 vdd.n1932 vdd.n1927 0.155672
R22424 vdd.n2007 vdd.n1969 0.155672
R22425 vdd.n1999 vdd.n1969 0.155672
R22426 vdd.n1999 vdd.n1998 0.155672
R22427 vdd.n1998 vdd.n1974 0.155672
R22428 vdd.n1991 vdd.n1974 0.155672
R22429 vdd.n1991 vdd.n1990 0.155672
R22430 vdd.n1990 vdd.n1978 0.155672
R22431 vdd.n1983 vdd.n1978 0.155672
R22432 vdd.n1862 vdd.n1824 0.155672
R22433 vdd.n1854 vdd.n1824 0.155672
R22434 vdd.n1854 vdd.n1853 0.155672
R22435 vdd.n1853 vdd.n1829 0.155672
R22436 vdd.n1846 vdd.n1829 0.155672
R22437 vdd.n1846 vdd.n1845 0.155672
R22438 vdd.n1845 vdd.n1833 0.155672
R22439 vdd.n1838 vdd.n1833 0.155672
R22440 vdd.n1913 vdd.n1875 0.155672
R22441 vdd.n1905 vdd.n1875 0.155672
R22442 vdd.n1905 vdd.n1904 0.155672
R22443 vdd.n1904 vdd.n1880 0.155672
R22444 vdd.n1897 vdd.n1880 0.155672
R22445 vdd.n1897 vdd.n1896 0.155672
R22446 vdd.n1896 vdd.n1884 0.155672
R22447 vdd.n1889 vdd.n1884 0.155672
R22448 vdd.n1769 vdd.n1731 0.155672
R22449 vdd.n1761 vdd.n1731 0.155672
R22450 vdd.n1761 vdd.n1760 0.155672
R22451 vdd.n1760 vdd.n1736 0.155672
R22452 vdd.n1753 vdd.n1736 0.155672
R22453 vdd.n1753 vdd.n1752 0.155672
R22454 vdd.n1752 vdd.n1740 0.155672
R22455 vdd.n1745 vdd.n1740 0.155672
R22456 vdd.n1820 vdd.n1782 0.155672
R22457 vdd.n1812 vdd.n1782 0.155672
R22458 vdd.n1812 vdd.n1811 0.155672
R22459 vdd.n1811 vdd.n1787 0.155672
R22460 vdd.n1804 vdd.n1787 0.155672
R22461 vdd.n1804 vdd.n1803 0.155672
R22462 vdd.n1803 vdd.n1791 0.155672
R22463 vdd.n1796 vdd.n1791 0.155672
R22464 vdd.n1014 vdd.n1006 0.152939
R22465 vdd.n1018 vdd.n1014 0.152939
R22466 vdd.n1019 vdd.n1018 0.152939
R22467 vdd.n1020 vdd.n1019 0.152939
R22468 vdd.n1021 vdd.n1020 0.152939
R22469 vdd.n1025 vdd.n1021 0.152939
R22470 vdd.n1026 vdd.n1025 0.152939
R22471 vdd.n1027 vdd.n1026 0.152939
R22472 vdd.n1028 vdd.n1027 0.152939
R22473 vdd.n1032 vdd.n1028 0.152939
R22474 vdd.n1033 vdd.n1032 0.152939
R22475 vdd.n1034 vdd.n1033 0.152939
R22476 vdd.n2150 vdd.n1034 0.152939
R22477 vdd.n2150 vdd.n2149 0.152939
R22478 vdd.n2149 vdd.n2148 0.152939
R22479 vdd.n2148 vdd.n1040 0.152939
R22480 vdd.n1045 vdd.n1040 0.152939
R22481 vdd.n1046 vdd.n1045 0.152939
R22482 vdd.n1047 vdd.n1046 0.152939
R22483 vdd.n1051 vdd.n1047 0.152939
R22484 vdd.n1052 vdd.n1051 0.152939
R22485 vdd.n1053 vdd.n1052 0.152939
R22486 vdd.n1054 vdd.n1053 0.152939
R22487 vdd.n1058 vdd.n1054 0.152939
R22488 vdd.n1059 vdd.n1058 0.152939
R22489 vdd.n1060 vdd.n1059 0.152939
R22490 vdd.n1061 vdd.n1060 0.152939
R22491 vdd.n1065 vdd.n1061 0.152939
R22492 vdd.n1066 vdd.n1065 0.152939
R22493 vdd.n1067 vdd.n1066 0.152939
R22494 vdd.n1068 vdd.n1067 0.152939
R22495 vdd.n1072 vdd.n1068 0.152939
R22496 vdd.n1073 vdd.n1072 0.152939
R22497 vdd.n1074 vdd.n1073 0.152939
R22498 vdd.n2111 vdd.n1074 0.152939
R22499 vdd.n2111 vdd.n2110 0.152939
R22500 vdd.n2110 vdd.n2109 0.152939
R22501 vdd.n2109 vdd.n1080 0.152939
R22502 vdd.n1085 vdd.n1080 0.152939
R22503 vdd.n1086 vdd.n1085 0.152939
R22504 vdd.n1087 vdd.n1086 0.152939
R22505 vdd.n1091 vdd.n1087 0.152939
R22506 vdd.n1092 vdd.n1091 0.152939
R22507 vdd.n1093 vdd.n1092 0.152939
R22508 vdd.n1094 vdd.n1093 0.152939
R22509 vdd.n1098 vdd.n1094 0.152939
R22510 vdd.n1099 vdd.n1098 0.152939
R22511 vdd.n1100 vdd.n1099 0.152939
R22512 vdd.n1101 vdd.n1100 0.152939
R22513 vdd.n1105 vdd.n1101 0.152939
R22514 vdd.n1106 vdd.n1105 0.152939
R22515 vdd.n2185 vdd.n1009 0.152939
R22516 vdd.n2014 vdd.n2013 0.152939
R22517 vdd.n2014 vdd.n1383 0.152939
R22518 vdd.n2029 vdd.n1383 0.152939
R22519 vdd.n2030 vdd.n2029 0.152939
R22520 vdd.n2031 vdd.n2030 0.152939
R22521 vdd.n2031 vdd.n1372 0.152939
R22522 vdd.n2046 vdd.n1372 0.152939
R22523 vdd.n2047 vdd.n2046 0.152939
R22524 vdd.n2048 vdd.n2047 0.152939
R22525 vdd.n2048 vdd.n1360 0.152939
R22526 vdd.n2065 vdd.n1360 0.152939
R22527 vdd.n2066 vdd.n2065 0.152939
R22528 vdd.n2067 vdd.n2066 0.152939
R22529 vdd.n527 vdd.n524 0.152939
R22530 vdd.n528 vdd.n527 0.152939
R22531 vdd.n529 vdd.n528 0.152939
R22532 vdd.n530 vdd.n529 0.152939
R22533 vdd.n533 vdd.n530 0.152939
R22534 vdd.n534 vdd.n533 0.152939
R22535 vdd.n535 vdd.n534 0.152939
R22536 vdd.n536 vdd.n535 0.152939
R22537 vdd.n539 vdd.n536 0.152939
R22538 vdd.n540 vdd.n539 0.152939
R22539 vdd.n541 vdd.n540 0.152939
R22540 vdd.n542 vdd.n541 0.152939
R22541 vdd.n547 vdd.n542 0.152939
R22542 vdd.n548 vdd.n547 0.152939
R22543 vdd.n549 vdd.n548 0.152939
R22544 vdd.n550 vdd.n549 0.152939
R22545 vdd.n553 vdd.n550 0.152939
R22546 vdd.n554 vdd.n553 0.152939
R22547 vdd.n555 vdd.n554 0.152939
R22548 vdd.n556 vdd.n555 0.152939
R22549 vdd.n559 vdd.n556 0.152939
R22550 vdd.n560 vdd.n559 0.152939
R22551 vdd.n561 vdd.n560 0.152939
R22552 vdd.n562 vdd.n561 0.152939
R22553 vdd.n565 vdd.n562 0.152939
R22554 vdd.n566 vdd.n565 0.152939
R22555 vdd.n567 vdd.n566 0.152939
R22556 vdd.n568 vdd.n567 0.152939
R22557 vdd.n571 vdd.n568 0.152939
R22558 vdd.n572 vdd.n571 0.152939
R22559 vdd.n573 vdd.n572 0.152939
R22560 vdd.n574 vdd.n573 0.152939
R22561 vdd.n577 vdd.n574 0.152939
R22562 vdd.n578 vdd.n577 0.152939
R22563 vdd.n3125 vdd.n578 0.152939
R22564 vdd.n3125 vdd.n3124 0.152939
R22565 vdd.n3124 vdd.n3123 0.152939
R22566 vdd.n3123 vdd.n582 0.152939
R22567 vdd.n587 vdd.n582 0.152939
R22568 vdd.n588 vdd.n587 0.152939
R22569 vdd.n591 vdd.n588 0.152939
R22570 vdd.n592 vdd.n591 0.152939
R22571 vdd.n593 vdd.n592 0.152939
R22572 vdd.n594 vdd.n593 0.152939
R22573 vdd.n597 vdd.n594 0.152939
R22574 vdd.n598 vdd.n597 0.152939
R22575 vdd.n599 vdd.n598 0.152939
R22576 vdd.n600 vdd.n599 0.152939
R22577 vdd.n603 vdd.n600 0.152939
R22578 vdd.n604 vdd.n603 0.152939
R22579 vdd.n605 vdd.n604 0.152939
R22580 vdd.n3208 vdd.n518 0.152939
R22581 vdd.n3209 vdd.n508 0.152939
R22582 vdd.n3223 vdd.n508 0.152939
R22583 vdd.n3224 vdd.n3223 0.152939
R22584 vdd.n3225 vdd.n3224 0.152939
R22585 vdd.n3225 vdd.n496 0.152939
R22586 vdd.n3239 vdd.n496 0.152939
R22587 vdd.n3240 vdd.n3239 0.152939
R22588 vdd.n3241 vdd.n3240 0.152939
R22589 vdd.n3241 vdd.n484 0.152939
R22590 vdd.n3256 vdd.n484 0.152939
R22591 vdd.n3257 vdd.n3256 0.152939
R22592 vdd.n3258 vdd.n3257 0.152939
R22593 vdd.n3258 vdd.n310 0.152939
R22594 vdd.n320 vdd.n311 0.152939
R22595 vdd.n321 vdd.n320 0.152939
R22596 vdd.n322 vdd.n321 0.152939
R22597 vdd.n331 vdd.n322 0.152939
R22598 vdd.n332 vdd.n331 0.152939
R22599 vdd.n333 vdd.n332 0.152939
R22600 vdd.n334 vdd.n333 0.152939
R22601 vdd.n342 vdd.n334 0.152939
R22602 vdd.n343 vdd.n342 0.152939
R22603 vdd.n344 vdd.n343 0.152939
R22604 vdd.n345 vdd.n344 0.152939
R22605 vdd.n353 vdd.n345 0.152939
R22606 vdd.n3407 vdd.n353 0.152939
R22607 vdd.n3406 vdd.n354 0.152939
R22608 vdd.n357 vdd.n354 0.152939
R22609 vdd.n361 vdd.n357 0.152939
R22610 vdd.n362 vdd.n361 0.152939
R22611 vdd.n363 vdd.n362 0.152939
R22612 vdd.n364 vdd.n363 0.152939
R22613 vdd.n365 vdd.n364 0.152939
R22614 vdd.n369 vdd.n365 0.152939
R22615 vdd.n370 vdd.n369 0.152939
R22616 vdd.n371 vdd.n370 0.152939
R22617 vdd.n372 vdd.n371 0.152939
R22618 vdd.n376 vdd.n372 0.152939
R22619 vdd.n377 vdd.n376 0.152939
R22620 vdd.n378 vdd.n377 0.152939
R22621 vdd.n379 vdd.n378 0.152939
R22622 vdd.n383 vdd.n379 0.152939
R22623 vdd.n384 vdd.n383 0.152939
R22624 vdd.n385 vdd.n384 0.152939
R22625 vdd.n3372 vdd.n385 0.152939
R22626 vdd.n3372 vdd.n3371 0.152939
R22627 vdd.n3371 vdd.n3370 0.152939
R22628 vdd.n3370 vdd.n391 0.152939
R22629 vdd.n396 vdd.n391 0.152939
R22630 vdd.n397 vdd.n396 0.152939
R22631 vdd.n398 vdd.n397 0.152939
R22632 vdd.n402 vdd.n398 0.152939
R22633 vdd.n403 vdd.n402 0.152939
R22634 vdd.n404 vdd.n403 0.152939
R22635 vdd.n405 vdd.n404 0.152939
R22636 vdd.n409 vdd.n405 0.152939
R22637 vdd.n410 vdd.n409 0.152939
R22638 vdd.n411 vdd.n410 0.152939
R22639 vdd.n412 vdd.n411 0.152939
R22640 vdd.n416 vdd.n412 0.152939
R22641 vdd.n417 vdd.n416 0.152939
R22642 vdd.n418 vdd.n417 0.152939
R22643 vdd.n419 vdd.n418 0.152939
R22644 vdd.n423 vdd.n419 0.152939
R22645 vdd.n424 vdd.n423 0.152939
R22646 vdd.n425 vdd.n424 0.152939
R22647 vdd.n3333 vdd.n425 0.152939
R22648 vdd.n3333 vdd.n3332 0.152939
R22649 vdd.n3332 vdd.n3331 0.152939
R22650 vdd.n3331 vdd.n431 0.152939
R22651 vdd.n436 vdd.n431 0.152939
R22652 vdd.n437 vdd.n436 0.152939
R22653 vdd.n438 vdd.n437 0.152939
R22654 vdd.n442 vdd.n438 0.152939
R22655 vdd.n443 vdd.n442 0.152939
R22656 vdd.n444 vdd.n443 0.152939
R22657 vdd.n445 vdd.n444 0.152939
R22658 vdd.n449 vdd.n445 0.152939
R22659 vdd.n450 vdd.n449 0.152939
R22660 vdd.n451 vdd.n450 0.152939
R22661 vdd.n452 vdd.n451 0.152939
R22662 vdd.n456 vdd.n452 0.152939
R22663 vdd.n457 vdd.n456 0.152939
R22664 vdd.n458 vdd.n457 0.152939
R22665 vdd.n459 vdd.n458 0.152939
R22666 vdd.n463 vdd.n459 0.152939
R22667 vdd.n464 vdd.n463 0.152939
R22668 vdd.n465 vdd.n464 0.152939
R22669 vdd.n3289 vdd.n465 0.152939
R22670 vdd.n3216 vdd.n3215 0.152939
R22671 vdd.n3217 vdd.n3216 0.152939
R22672 vdd.n3217 vdd.n502 0.152939
R22673 vdd.n3231 vdd.n502 0.152939
R22674 vdd.n3232 vdd.n3231 0.152939
R22675 vdd.n3233 vdd.n3232 0.152939
R22676 vdd.n3233 vdd.n489 0.152939
R22677 vdd.n3247 vdd.n489 0.152939
R22678 vdd.n3248 vdd.n3247 0.152939
R22679 vdd.n3249 vdd.n3248 0.152939
R22680 vdd.n3249 vdd.n477 0.152939
R22681 vdd.n3264 vdd.n477 0.152939
R22682 vdd.n3265 vdd.n3264 0.152939
R22683 vdd.n3266 vdd.n3265 0.152939
R22684 vdd.n3266 vdd.n475 0.152939
R22685 vdd.n3270 vdd.n475 0.152939
R22686 vdd.n3271 vdd.n3270 0.152939
R22687 vdd.n3272 vdd.n3271 0.152939
R22688 vdd.n3272 vdd.n472 0.152939
R22689 vdd.n3276 vdd.n472 0.152939
R22690 vdd.n3277 vdd.n3276 0.152939
R22691 vdd.n3278 vdd.n3277 0.152939
R22692 vdd.n3278 vdd.n469 0.152939
R22693 vdd.n3282 vdd.n469 0.152939
R22694 vdd.n3283 vdd.n3282 0.152939
R22695 vdd.n3284 vdd.n3283 0.152939
R22696 vdd.n3284 vdd.n466 0.152939
R22697 vdd.n3288 vdd.n466 0.152939
R22698 vdd.n3078 vdd.n514 0.152939
R22699 vdd.n2078 vdd.n1345 0.152939
R22700 vdd.n1674 vdd.n1673 0.152939
R22701 vdd.n1675 vdd.n1674 0.152939
R22702 vdd.n1675 vdd.n1424 0.152939
R22703 vdd.n1689 vdd.n1424 0.152939
R22704 vdd.n1690 vdd.n1689 0.152939
R22705 vdd.n1691 vdd.n1690 0.152939
R22706 vdd.n1691 vdd.n1411 0.152939
R22707 vdd.n1705 vdd.n1411 0.152939
R22708 vdd.n1706 vdd.n1705 0.152939
R22709 vdd.n1707 vdd.n1706 0.152939
R22710 vdd.n1707 vdd.n1400 0.152939
R22711 vdd.n1722 vdd.n1400 0.152939
R22712 vdd.n1723 vdd.n1722 0.152939
R22713 vdd.n1724 vdd.n1723 0.152939
R22714 vdd.n1724 vdd.n1389 0.152939
R22715 vdd.n2020 vdd.n1389 0.152939
R22716 vdd.n2021 vdd.n2020 0.152939
R22717 vdd.n2022 vdd.n2021 0.152939
R22718 vdd.n2022 vdd.n1377 0.152939
R22719 vdd.n2037 vdd.n1377 0.152939
R22720 vdd.n2038 vdd.n2037 0.152939
R22721 vdd.n2039 vdd.n2038 0.152939
R22722 vdd.n2039 vdd.n1367 0.152939
R22723 vdd.n2054 vdd.n1367 0.152939
R22724 vdd.n2055 vdd.n2054 0.152939
R22725 vdd.n2058 vdd.n2055 0.152939
R22726 vdd.n2058 vdd.n2057 0.152939
R22727 vdd.n2057 vdd.n2056 0.152939
R22728 vdd.n1666 vdd.n1440 0.152939
R22729 vdd.n1662 vdd.n1440 0.152939
R22730 vdd.n1662 vdd.n1661 0.152939
R22731 vdd.n1661 vdd.n1660 0.152939
R22732 vdd.n1660 vdd.n1445 0.152939
R22733 vdd.n1656 vdd.n1445 0.152939
R22734 vdd.n1656 vdd.n1655 0.152939
R22735 vdd.n1655 vdd.n1654 0.152939
R22736 vdd.n1654 vdd.n1453 0.152939
R22737 vdd.n1650 vdd.n1453 0.152939
R22738 vdd.n1650 vdd.n1649 0.152939
R22739 vdd.n1649 vdd.n1648 0.152939
R22740 vdd.n1648 vdd.n1461 0.152939
R22741 vdd.n1644 vdd.n1461 0.152939
R22742 vdd.n1644 vdd.n1643 0.152939
R22743 vdd.n1643 vdd.n1642 0.152939
R22744 vdd.n1642 vdd.n1469 0.152939
R22745 vdd.n1638 vdd.n1469 0.152939
R22746 vdd.n1638 vdd.n1637 0.152939
R22747 vdd.n1637 vdd.n1636 0.152939
R22748 vdd.n1636 vdd.n1479 0.152939
R22749 vdd.n1632 vdd.n1479 0.152939
R22750 vdd.n1632 vdd.n1631 0.152939
R22751 vdd.n1631 vdd.n1630 0.152939
R22752 vdd.n1630 vdd.n1487 0.152939
R22753 vdd.n1626 vdd.n1487 0.152939
R22754 vdd.n1626 vdd.n1625 0.152939
R22755 vdd.n1625 vdd.n1624 0.152939
R22756 vdd.n1624 vdd.n1495 0.152939
R22757 vdd.n1620 vdd.n1495 0.152939
R22758 vdd.n1620 vdd.n1619 0.152939
R22759 vdd.n1619 vdd.n1618 0.152939
R22760 vdd.n1618 vdd.n1503 0.152939
R22761 vdd.n1614 vdd.n1503 0.152939
R22762 vdd.n1614 vdd.n1613 0.152939
R22763 vdd.n1613 vdd.n1612 0.152939
R22764 vdd.n1612 vdd.n1511 0.152939
R22765 vdd.n1608 vdd.n1511 0.152939
R22766 vdd.n1608 vdd.n1607 0.152939
R22767 vdd.n1607 vdd.n1606 0.152939
R22768 vdd.n1606 vdd.n1519 0.152939
R22769 vdd.n1526 vdd.n1519 0.152939
R22770 vdd.n1596 vdd.n1526 0.152939
R22771 vdd.n1596 vdd.n1595 0.152939
R22772 vdd.n1595 vdd.n1594 0.152939
R22773 vdd.n1594 vdd.n1527 0.152939
R22774 vdd.n1590 vdd.n1527 0.152939
R22775 vdd.n1590 vdd.n1589 0.152939
R22776 vdd.n1589 vdd.n1588 0.152939
R22777 vdd.n1588 vdd.n1534 0.152939
R22778 vdd.n1584 vdd.n1534 0.152939
R22779 vdd.n1584 vdd.n1583 0.152939
R22780 vdd.n1583 vdd.n1582 0.152939
R22781 vdd.n1582 vdd.n1542 0.152939
R22782 vdd.n1578 vdd.n1542 0.152939
R22783 vdd.n1578 vdd.n1577 0.152939
R22784 vdd.n1577 vdd.n1576 0.152939
R22785 vdd.n1576 vdd.n1550 0.152939
R22786 vdd.n1572 vdd.n1550 0.152939
R22787 vdd.n1572 vdd.n1571 0.152939
R22788 vdd.n1571 vdd.n1570 0.152939
R22789 vdd.n1570 vdd.n1558 0.152939
R22790 vdd.n1558 vdd.n1435 0.152939
R22791 vdd.n1667 vdd.n1430 0.152939
R22792 vdd.n1681 vdd.n1430 0.152939
R22793 vdd.n1682 vdd.n1681 0.152939
R22794 vdd.n1683 vdd.n1682 0.152939
R22795 vdd.n1683 vdd.n1418 0.152939
R22796 vdd.n1697 vdd.n1418 0.152939
R22797 vdd.n1698 vdd.n1697 0.152939
R22798 vdd.n1699 vdd.n1698 0.152939
R22799 vdd.n1699 vdd.n1406 0.152939
R22800 vdd.n1714 vdd.n1406 0.152939
R22801 vdd.n1715 vdd.n1714 0.152939
R22802 vdd.n1716 vdd.n1715 0.152939
R22803 vdd.n1716 vdd.n1395 0.152939
R22804 vdd.n2013 vdd.n2012 0.145814
R22805 vdd.n3439 vdd.n310 0.145814
R22806 vdd.n3439 vdd.n311 0.145814
R22807 vdd.n2012 vdd.n1395 0.145814
R22808 vdd.n2186 vdd.n2185 0.110256
R22809 vdd.n3009 vdd.n518 0.110256
R22810 vdd.n3078 vdd.n3077 0.110256
R22811 vdd.n2079 vdd.n2078 0.110256
R22812 vdd.n2186 vdd.n1006 0.0431829
R22813 vdd.n2079 vdd.n1106 0.0431829
R22814 vdd.n3009 vdd.n524 0.0431829
R22815 vdd.n3077 vdd.n605 0.0431829
R22816 vdd vdd.n28 0.00833333
R22817 CSoutput.n19 CSoutput.t209 184.661
R22818 CSoutput.n78 CSoutput.n77 165.8
R22819 CSoutput.n76 CSoutput.n0 165.8
R22820 CSoutput.n75 CSoutput.n74 165.8
R22821 CSoutput.n73 CSoutput.n72 165.8
R22822 CSoutput.n71 CSoutput.n2 165.8
R22823 CSoutput.n69 CSoutput.n68 165.8
R22824 CSoutput.n67 CSoutput.n3 165.8
R22825 CSoutput.n66 CSoutput.n65 165.8
R22826 CSoutput.n63 CSoutput.n4 165.8
R22827 CSoutput.n61 CSoutput.n60 165.8
R22828 CSoutput.n59 CSoutput.n5 165.8
R22829 CSoutput.n58 CSoutput.n57 165.8
R22830 CSoutput.n55 CSoutput.n6 165.8
R22831 CSoutput.n54 CSoutput.n53 165.8
R22832 CSoutput.n52 CSoutput.n51 165.8
R22833 CSoutput.n50 CSoutput.n8 165.8
R22834 CSoutput.n48 CSoutput.n47 165.8
R22835 CSoutput.n46 CSoutput.n9 165.8
R22836 CSoutput.n45 CSoutput.n44 165.8
R22837 CSoutput.n42 CSoutput.n10 165.8
R22838 CSoutput.n41 CSoutput.n40 165.8
R22839 CSoutput.n39 CSoutput.n38 165.8
R22840 CSoutput.n37 CSoutput.n12 165.8
R22841 CSoutput.n35 CSoutput.n34 165.8
R22842 CSoutput.n33 CSoutput.n13 165.8
R22843 CSoutput.n32 CSoutput.n31 165.8
R22844 CSoutput.n29 CSoutput.n14 165.8
R22845 CSoutput.n28 CSoutput.n27 165.8
R22846 CSoutput.n26 CSoutput.n25 165.8
R22847 CSoutput.n24 CSoutput.n16 165.8
R22848 CSoutput.n22 CSoutput.n21 165.8
R22849 CSoutput.n20 CSoutput.n17 165.8
R22850 CSoutput.n77 CSoutput.t212 162.194
R22851 CSoutput.n18 CSoutput.t205 120.501
R22852 CSoutput.n23 CSoutput.t198 120.501
R22853 CSoutput.n15 CSoutput.t193 120.501
R22854 CSoutput.n30 CSoutput.t207 120.501
R22855 CSoutput.n36 CSoutput.t208 120.501
R22856 CSoutput.n11 CSoutput.t195 120.501
R22857 CSoutput.n43 CSoutput.t192 120.501
R22858 CSoutput.n49 CSoutput.t211 120.501
R22859 CSoutput.n7 CSoutput.t199 120.501
R22860 CSoutput.n56 CSoutput.t202 120.501
R22861 CSoutput.n62 CSoutput.t213 120.501
R22862 CSoutput.n64 CSoutput.t203 120.501
R22863 CSoutput.n70 CSoutput.t204 120.501
R22864 CSoutput.n1 CSoutput.t197 120.501
R22865 CSoutput.n290 CSoutput.n288 103.469
R22866 CSoutput.n278 CSoutput.n276 103.469
R22867 CSoutput.n267 CSoutput.n265 103.469
R22868 CSoutput.n104 CSoutput.n102 103.469
R22869 CSoutput.n92 CSoutput.n90 103.469
R22870 CSoutput.n81 CSoutput.n79 103.469
R22871 CSoutput.n296 CSoutput.n295 103.111
R22872 CSoutput.n294 CSoutput.n293 103.111
R22873 CSoutput.n292 CSoutput.n291 103.111
R22874 CSoutput.n290 CSoutput.n289 103.111
R22875 CSoutput.n286 CSoutput.n285 103.111
R22876 CSoutput.n284 CSoutput.n283 103.111
R22877 CSoutput.n282 CSoutput.n281 103.111
R22878 CSoutput.n280 CSoutput.n279 103.111
R22879 CSoutput.n278 CSoutput.n277 103.111
R22880 CSoutput.n275 CSoutput.n274 103.111
R22881 CSoutput.n273 CSoutput.n272 103.111
R22882 CSoutput.n271 CSoutput.n270 103.111
R22883 CSoutput.n269 CSoutput.n268 103.111
R22884 CSoutput.n267 CSoutput.n266 103.111
R22885 CSoutput.n104 CSoutput.n103 103.111
R22886 CSoutput.n106 CSoutput.n105 103.111
R22887 CSoutput.n108 CSoutput.n107 103.111
R22888 CSoutput.n110 CSoutput.n109 103.111
R22889 CSoutput.n112 CSoutput.n111 103.111
R22890 CSoutput.n92 CSoutput.n91 103.111
R22891 CSoutput.n94 CSoutput.n93 103.111
R22892 CSoutput.n96 CSoutput.n95 103.111
R22893 CSoutput.n98 CSoutput.n97 103.111
R22894 CSoutput.n100 CSoutput.n99 103.111
R22895 CSoutput.n81 CSoutput.n80 103.111
R22896 CSoutput.n83 CSoutput.n82 103.111
R22897 CSoutput.n85 CSoutput.n84 103.111
R22898 CSoutput.n87 CSoutput.n86 103.111
R22899 CSoutput.n89 CSoutput.n88 103.111
R22900 CSoutput.n298 CSoutput.n297 103.111
R22901 CSoutput.n342 CSoutput.n340 81.5057
R22902 CSoutput.n322 CSoutput.n320 81.5057
R22903 CSoutput.n303 CSoutput.n301 81.5057
R22904 CSoutput.n402 CSoutput.n400 81.5057
R22905 CSoutput.n382 CSoutput.n380 81.5057
R22906 CSoutput.n363 CSoutput.n361 81.5057
R22907 CSoutput.n358 CSoutput.n357 80.9324
R22908 CSoutput.n356 CSoutput.n355 80.9324
R22909 CSoutput.n354 CSoutput.n353 80.9324
R22910 CSoutput.n352 CSoutput.n351 80.9324
R22911 CSoutput.n350 CSoutput.n349 80.9324
R22912 CSoutput.n348 CSoutput.n347 80.9324
R22913 CSoutput.n346 CSoutput.n345 80.9324
R22914 CSoutput.n344 CSoutput.n343 80.9324
R22915 CSoutput.n342 CSoutput.n341 80.9324
R22916 CSoutput.n338 CSoutput.n337 80.9324
R22917 CSoutput.n336 CSoutput.n335 80.9324
R22918 CSoutput.n334 CSoutput.n333 80.9324
R22919 CSoutput.n332 CSoutput.n331 80.9324
R22920 CSoutput.n330 CSoutput.n329 80.9324
R22921 CSoutput.n328 CSoutput.n327 80.9324
R22922 CSoutput.n326 CSoutput.n325 80.9324
R22923 CSoutput.n324 CSoutput.n323 80.9324
R22924 CSoutput.n322 CSoutput.n321 80.9324
R22925 CSoutput.n319 CSoutput.n318 80.9324
R22926 CSoutput.n317 CSoutput.n316 80.9324
R22927 CSoutput.n315 CSoutput.n314 80.9324
R22928 CSoutput.n313 CSoutput.n312 80.9324
R22929 CSoutput.n311 CSoutput.n310 80.9324
R22930 CSoutput.n309 CSoutput.n308 80.9324
R22931 CSoutput.n307 CSoutput.n306 80.9324
R22932 CSoutput.n305 CSoutput.n304 80.9324
R22933 CSoutput.n303 CSoutput.n302 80.9324
R22934 CSoutput.n402 CSoutput.n401 80.9324
R22935 CSoutput.n404 CSoutput.n403 80.9324
R22936 CSoutput.n406 CSoutput.n405 80.9324
R22937 CSoutput.n408 CSoutput.n407 80.9324
R22938 CSoutput.n410 CSoutput.n409 80.9324
R22939 CSoutput.n412 CSoutput.n411 80.9324
R22940 CSoutput.n414 CSoutput.n413 80.9324
R22941 CSoutput.n416 CSoutput.n415 80.9324
R22942 CSoutput.n418 CSoutput.n417 80.9324
R22943 CSoutput.n382 CSoutput.n381 80.9324
R22944 CSoutput.n384 CSoutput.n383 80.9324
R22945 CSoutput.n386 CSoutput.n385 80.9324
R22946 CSoutput.n388 CSoutput.n387 80.9324
R22947 CSoutput.n390 CSoutput.n389 80.9324
R22948 CSoutput.n392 CSoutput.n391 80.9324
R22949 CSoutput.n394 CSoutput.n393 80.9324
R22950 CSoutput.n396 CSoutput.n395 80.9324
R22951 CSoutput.n398 CSoutput.n397 80.9324
R22952 CSoutput.n363 CSoutput.n362 80.9324
R22953 CSoutput.n365 CSoutput.n364 80.9324
R22954 CSoutput.n367 CSoutput.n366 80.9324
R22955 CSoutput.n369 CSoutput.n368 80.9324
R22956 CSoutput.n371 CSoutput.n370 80.9324
R22957 CSoutput.n373 CSoutput.n372 80.9324
R22958 CSoutput.n375 CSoutput.n374 80.9324
R22959 CSoutput.n377 CSoutput.n376 80.9324
R22960 CSoutput.n379 CSoutput.n378 80.9324
R22961 CSoutput.n25 CSoutput.n24 48.1486
R22962 CSoutput.n69 CSoutput.n3 48.1486
R22963 CSoutput.n38 CSoutput.n37 48.1486
R22964 CSoutput.n42 CSoutput.n41 48.1486
R22965 CSoutput.n51 CSoutput.n50 48.1486
R22966 CSoutput.n55 CSoutput.n54 48.1486
R22967 CSoutput.n22 CSoutput.n17 46.462
R22968 CSoutput.n72 CSoutput.n71 46.462
R22969 CSoutput.n20 CSoutput.n19 44.9055
R22970 CSoutput.n29 CSoutput.n28 43.7635
R22971 CSoutput.n65 CSoutput.n63 43.7635
R22972 CSoutput.n35 CSoutput.n13 41.7396
R22973 CSoutput.n57 CSoutput.n5 41.7396
R22974 CSoutput.n44 CSoutput.n9 37.0171
R22975 CSoutput.n48 CSoutput.n9 37.0171
R22976 CSoutput.n76 CSoutput.n75 34.9932
R22977 CSoutput.n31 CSoutput.n13 32.2947
R22978 CSoutput.n61 CSoutput.n5 32.2947
R22979 CSoutput.n30 CSoutput.n29 29.6014
R22980 CSoutput.n63 CSoutput.n62 29.6014
R22981 CSoutput.n19 CSoutput.n18 28.4085
R22982 CSoutput.n18 CSoutput.n17 25.1176
R22983 CSoutput.n72 CSoutput.n1 25.1176
R22984 CSoutput.n43 CSoutput.n42 22.0922
R22985 CSoutput.n50 CSoutput.n49 22.0922
R22986 CSoutput.n77 CSoutput.n76 21.8586
R22987 CSoutput.n37 CSoutput.n36 18.9681
R22988 CSoutput.n56 CSoutput.n55 18.9681
R22989 CSoutput.n25 CSoutput.n15 17.6292
R22990 CSoutput.n64 CSoutput.n3 17.6292
R22991 CSoutput.n24 CSoutput.n23 15.844
R22992 CSoutput.n70 CSoutput.n69 15.844
R22993 CSoutput.n38 CSoutput.n11 14.5051
R22994 CSoutput.n54 CSoutput.n7 14.5051
R22995 CSoutput.n421 CSoutput.n78 11.4982
R22996 CSoutput.n41 CSoutput.n11 11.3811
R22997 CSoutput.n51 CSoutput.n7 11.3811
R22998 CSoutput.n23 CSoutput.n22 10.0422
R22999 CSoutput.n71 CSoutput.n70 10.0422
R23000 CSoutput.n287 CSoutput.n275 9.25285
R23001 CSoutput.n101 CSoutput.n89 9.25285
R23002 CSoutput.n360 CSoutput.n300 8.99065
R23003 CSoutput.n339 CSoutput.n319 8.98182
R23004 CSoutput.n399 CSoutput.n379 8.98182
R23005 CSoutput.n28 CSoutput.n15 8.25698
R23006 CSoutput.n65 CSoutput.n64 8.25698
R23007 CSoutput.n300 CSoutput.n299 7.12641
R23008 CSoutput.n114 CSoutput.n113 7.12641
R23009 CSoutput.n36 CSoutput.n35 6.91809
R23010 CSoutput.n57 CSoutput.n56 6.91809
R23011 CSoutput.n360 CSoutput.n359 6.02792
R23012 CSoutput.n420 CSoutput.n419 6.02792
R23013 CSoutput.n421 CSoutput.n114 5.39821
R23014 CSoutput.n359 CSoutput.n358 5.25266
R23015 CSoutput.n339 CSoutput.n338 5.25266
R23016 CSoutput.n419 CSoutput.n418 5.25266
R23017 CSoutput.n399 CSoutput.n398 5.25266
R23018 CSoutput.n299 CSoutput.n298 5.1449
R23019 CSoutput.n287 CSoutput.n286 5.1449
R23020 CSoutput.n113 CSoutput.n112 5.1449
R23021 CSoutput.n101 CSoutput.n100 5.1449
R23022 CSoutput.n205 CSoutput.n158 4.5005
R23023 CSoutput.n174 CSoutput.n158 4.5005
R23024 CSoutput.n169 CSoutput.n153 4.5005
R23025 CSoutput.n169 CSoutput.n155 4.5005
R23026 CSoutput.n169 CSoutput.n152 4.5005
R23027 CSoutput.n169 CSoutput.n156 4.5005
R23028 CSoutput.n169 CSoutput.n151 4.5005
R23029 CSoutput.n169 CSoutput.t196 4.5005
R23030 CSoutput.n169 CSoutput.n150 4.5005
R23031 CSoutput.n169 CSoutput.n157 4.5005
R23032 CSoutput.n169 CSoutput.n158 4.5005
R23033 CSoutput.n167 CSoutput.n153 4.5005
R23034 CSoutput.n167 CSoutput.n155 4.5005
R23035 CSoutput.n167 CSoutput.n152 4.5005
R23036 CSoutput.n167 CSoutput.n156 4.5005
R23037 CSoutput.n167 CSoutput.n151 4.5005
R23038 CSoutput.n167 CSoutput.t196 4.5005
R23039 CSoutput.n167 CSoutput.n150 4.5005
R23040 CSoutput.n167 CSoutput.n157 4.5005
R23041 CSoutput.n167 CSoutput.n158 4.5005
R23042 CSoutput.n166 CSoutput.n153 4.5005
R23043 CSoutput.n166 CSoutput.n155 4.5005
R23044 CSoutput.n166 CSoutput.n152 4.5005
R23045 CSoutput.n166 CSoutput.n156 4.5005
R23046 CSoutput.n166 CSoutput.n151 4.5005
R23047 CSoutput.n166 CSoutput.t196 4.5005
R23048 CSoutput.n166 CSoutput.n150 4.5005
R23049 CSoutput.n166 CSoutput.n157 4.5005
R23050 CSoutput.n166 CSoutput.n158 4.5005
R23051 CSoutput.n251 CSoutput.n153 4.5005
R23052 CSoutput.n251 CSoutput.n155 4.5005
R23053 CSoutput.n251 CSoutput.n152 4.5005
R23054 CSoutput.n251 CSoutput.n156 4.5005
R23055 CSoutput.n251 CSoutput.n151 4.5005
R23056 CSoutput.n251 CSoutput.t196 4.5005
R23057 CSoutput.n251 CSoutput.n150 4.5005
R23058 CSoutput.n251 CSoutput.n157 4.5005
R23059 CSoutput.n251 CSoutput.n158 4.5005
R23060 CSoutput.n249 CSoutput.n153 4.5005
R23061 CSoutput.n249 CSoutput.n155 4.5005
R23062 CSoutput.n249 CSoutput.n152 4.5005
R23063 CSoutput.n249 CSoutput.n156 4.5005
R23064 CSoutput.n249 CSoutput.n151 4.5005
R23065 CSoutput.n249 CSoutput.t196 4.5005
R23066 CSoutput.n249 CSoutput.n150 4.5005
R23067 CSoutput.n249 CSoutput.n157 4.5005
R23068 CSoutput.n247 CSoutput.n153 4.5005
R23069 CSoutput.n247 CSoutput.n155 4.5005
R23070 CSoutput.n247 CSoutput.n152 4.5005
R23071 CSoutput.n247 CSoutput.n156 4.5005
R23072 CSoutput.n247 CSoutput.n151 4.5005
R23073 CSoutput.n247 CSoutput.t196 4.5005
R23074 CSoutput.n247 CSoutput.n150 4.5005
R23075 CSoutput.n247 CSoutput.n157 4.5005
R23076 CSoutput.n177 CSoutput.n153 4.5005
R23077 CSoutput.n177 CSoutput.n155 4.5005
R23078 CSoutput.n177 CSoutput.n152 4.5005
R23079 CSoutput.n177 CSoutput.n156 4.5005
R23080 CSoutput.n177 CSoutput.n151 4.5005
R23081 CSoutput.n177 CSoutput.t196 4.5005
R23082 CSoutput.n177 CSoutput.n150 4.5005
R23083 CSoutput.n177 CSoutput.n157 4.5005
R23084 CSoutput.n177 CSoutput.n158 4.5005
R23085 CSoutput.n176 CSoutput.n153 4.5005
R23086 CSoutput.n176 CSoutput.n155 4.5005
R23087 CSoutput.n176 CSoutput.n152 4.5005
R23088 CSoutput.n176 CSoutput.n156 4.5005
R23089 CSoutput.n176 CSoutput.n151 4.5005
R23090 CSoutput.n176 CSoutput.t196 4.5005
R23091 CSoutput.n176 CSoutput.n150 4.5005
R23092 CSoutput.n176 CSoutput.n157 4.5005
R23093 CSoutput.n176 CSoutput.n158 4.5005
R23094 CSoutput.n180 CSoutput.n153 4.5005
R23095 CSoutput.n180 CSoutput.n155 4.5005
R23096 CSoutput.n180 CSoutput.n152 4.5005
R23097 CSoutput.n180 CSoutput.n156 4.5005
R23098 CSoutput.n180 CSoutput.n151 4.5005
R23099 CSoutput.n180 CSoutput.t196 4.5005
R23100 CSoutput.n180 CSoutput.n150 4.5005
R23101 CSoutput.n180 CSoutput.n157 4.5005
R23102 CSoutput.n180 CSoutput.n158 4.5005
R23103 CSoutput.n179 CSoutput.n153 4.5005
R23104 CSoutput.n179 CSoutput.n155 4.5005
R23105 CSoutput.n179 CSoutput.n152 4.5005
R23106 CSoutput.n179 CSoutput.n156 4.5005
R23107 CSoutput.n179 CSoutput.n151 4.5005
R23108 CSoutput.n179 CSoutput.t196 4.5005
R23109 CSoutput.n179 CSoutput.n150 4.5005
R23110 CSoutput.n179 CSoutput.n157 4.5005
R23111 CSoutput.n179 CSoutput.n158 4.5005
R23112 CSoutput.n162 CSoutput.n153 4.5005
R23113 CSoutput.n162 CSoutput.n155 4.5005
R23114 CSoutput.n162 CSoutput.n152 4.5005
R23115 CSoutput.n162 CSoutput.n156 4.5005
R23116 CSoutput.n162 CSoutput.n151 4.5005
R23117 CSoutput.n162 CSoutput.t196 4.5005
R23118 CSoutput.n162 CSoutput.n150 4.5005
R23119 CSoutput.n162 CSoutput.n157 4.5005
R23120 CSoutput.n162 CSoutput.n158 4.5005
R23121 CSoutput.n254 CSoutput.n153 4.5005
R23122 CSoutput.n254 CSoutput.n155 4.5005
R23123 CSoutput.n254 CSoutput.n152 4.5005
R23124 CSoutput.n254 CSoutput.n156 4.5005
R23125 CSoutput.n254 CSoutput.n151 4.5005
R23126 CSoutput.n254 CSoutput.t196 4.5005
R23127 CSoutput.n254 CSoutput.n150 4.5005
R23128 CSoutput.n254 CSoutput.n157 4.5005
R23129 CSoutput.n254 CSoutput.n158 4.5005
R23130 CSoutput.n241 CSoutput.n212 4.5005
R23131 CSoutput.n241 CSoutput.n218 4.5005
R23132 CSoutput.n199 CSoutput.n188 4.5005
R23133 CSoutput.n199 CSoutput.n190 4.5005
R23134 CSoutput.n199 CSoutput.n187 4.5005
R23135 CSoutput.n199 CSoutput.n191 4.5005
R23136 CSoutput.n199 CSoutput.n186 4.5005
R23137 CSoutput.n199 CSoutput.t200 4.5005
R23138 CSoutput.n199 CSoutput.n185 4.5005
R23139 CSoutput.n199 CSoutput.n192 4.5005
R23140 CSoutput.n241 CSoutput.n199 4.5005
R23141 CSoutput.n220 CSoutput.n188 4.5005
R23142 CSoutput.n220 CSoutput.n190 4.5005
R23143 CSoutput.n220 CSoutput.n187 4.5005
R23144 CSoutput.n220 CSoutput.n191 4.5005
R23145 CSoutput.n220 CSoutput.n186 4.5005
R23146 CSoutput.n220 CSoutput.t200 4.5005
R23147 CSoutput.n220 CSoutput.n185 4.5005
R23148 CSoutput.n220 CSoutput.n192 4.5005
R23149 CSoutput.n241 CSoutput.n220 4.5005
R23150 CSoutput.n198 CSoutput.n188 4.5005
R23151 CSoutput.n198 CSoutput.n190 4.5005
R23152 CSoutput.n198 CSoutput.n187 4.5005
R23153 CSoutput.n198 CSoutput.n191 4.5005
R23154 CSoutput.n198 CSoutput.n186 4.5005
R23155 CSoutput.n198 CSoutput.t200 4.5005
R23156 CSoutput.n198 CSoutput.n185 4.5005
R23157 CSoutput.n198 CSoutput.n192 4.5005
R23158 CSoutput.n241 CSoutput.n198 4.5005
R23159 CSoutput.n222 CSoutput.n188 4.5005
R23160 CSoutput.n222 CSoutput.n190 4.5005
R23161 CSoutput.n222 CSoutput.n187 4.5005
R23162 CSoutput.n222 CSoutput.n191 4.5005
R23163 CSoutput.n222 CSoutput.n186 4.5005
R23164 CSoutput.n222 CSoutput.t200 4.5005
R23165 CSoutput.n222 CSoutput.n185 4.5005
R23166 CSoutput.n222 CSoutput.n192 4.5005
R23167 CSoutput.n241 CSoutput.n222 4.5005
R23168 CSoutput.n188 CSoutput.n183 4.5005
R23169 CSoutput.n190 CSoutput.n183 4.5005
R23170 CSoutput.n187 CSoutput.n183 4.5005
R23171 CSoutput.n191 CSoutput.n183 4.5005
R23172 CSoutput.n186 CSoutput.n183 4.5005
R23173 CSoutput.t200 CSoutput.n183 4.5005
R23174 CSoutput.n185 CSoutput.n183 4.5005
R23175 CSoutput.n192 CSoutput.n183 4.5005
R23176 CSoutput.n244 CSoutput.n188 4.5005
R23177 CSoutput.n244 CSoutput.n190 4.5005
R23178 CSoutput.n244 CSoutput.n187 4.5005
R23179 CSoutput.n244 CSoutput.n191 4.5005
R23180 CSoutput.n244 CSoutput.n186 4.5005
R23181 CSoutput.n244 CSoutput.t200 4.5005
R23182 CSoutput.n244 CSoutput.n185 4.5005
R23183 CSoutput.n244 CSoutput.n192 4.5005
R23184 CSoutput.n242 CSoutput.n188 4.5005
R23185 CSoutput.n242 CSoutput.n190 4.5005
R23186 CSoutput.n242 CSoutput.n187 4.5005
R23187 CSoutput.n242 CSoutput.n191 4.5005
R23188 CSoutput.n242 CSoutput.n186 4.5005
R23189 CSoutput.n242 CSoutput.t200 4.5005
R23190 CSoutput.n242 CSoutput.n185 4.5005
R23191 CSoutput.n242 CSoutput.n192 4.5005
R23192 CSoutput.n242 CSoutput.n241 4.5005
R23193 CSoutput.n224 CSoutput.n188 4.5005
R23194 CSoutput.n224 CSoutput.n190 4.5005
R23195 CSoutput.n224 CSoutput.n187 4.5005
R23196 CSoutput.n224 CSoutput.n191 4.5005
R23197 CSoutput.n224 CSoutput.n186 4.5005
R23198 CSoutput.n224 CSoutput.t200 4.5005
R23199 CSoutput.n224 CSoutput.n185 4.5005
R23200 CSoutput.n224 CSoutput.n192 4.5005
R23201 CSoutput.n241 CSoutput.n224 4.5005
R23202 CSoutput.n196 CSoutput.n188 4.5005
R23203 CSoutput.n196 CSoutput.n190 4.5005
R23204 CSoutput.n196 CSoutput.n187 4.5005
R23205 CSoutput.n196 CSoutput.n191 4.5005
R23206 CSoutput.n196 CSoutput.n186 4.5005
R23207 CSoutput.n196 CSoutput.t200 4.5005
R23208 CSoutput.n196 CSoutput.n185 4.5005
R23209 CSoutput.n196 CSoutput.n192 4.5005
R23210 CSoutput.n241 CSoutput.n196 4.5005
R23211 CSoutput.n226 CSoutput.n188 4.5005
R23212 CSoutput.n226 CSoutput.n190 4.5005
R23213 CSoutput.n226 CSoutput.n187 4.5005
R23214 CSoutput.n226 CSoutput.n191 4.5005
R23215 CSoutput.n226 CSoutput.n186 4.5005
R23216 CSoutput.n226 CSoutput.t200 4.5005
R23217 CSoutput.n226 CSoutput.n185 4.5005
R23218 CSoutput.n226 CSoutput.n192 4.5005
R23219 CSoutput.n241 CSoutput.n226 4.5005
R23220 CSoutput.n195 CSoutput.n188 4.5005
R23221 CSoutput.n195 CSoutput.n190 4.5005
R23222 CSoutput.n195 CSoutput.n187 4.5005
R23223 CSoutput.n195 CSoutput.n191 4.5005
R23224 CSoutput.n195 CSoutput.n186 4.5005
R23225 CSoutput.n195 CSoutput.t200 4.5005
R23226 CSoutput.n195 CSoutput.n185 4.5005
R23227 CSoutput.n195 CSoutput.n192 4.5005
R23228 CSoutput.n241 CSoutput.n195 4.5005
R23229 CSoutput.n240 CSoutput.n188 4.5005
R23230 CSoutput.n240 CSoutput.n190 4.5005
R23231 CSoutput.n240 CSoutput.n187 4.5005
R23232 CSoutput.n240 CSoutput.n191 4.5005
R23233 CSoutput.n240 CSoutput.n186 4.5005
R23234 CSoutput.n240 CSoutput.t200 4.5005
R23235 CSoutput.n240 CSoutput.n185 4.5005
R23236 CSoutput.n240 CSoutput.n192 4.5005
R23237 CSoutput.n241 CSoutput.n240 4.5005
R23238 CSoutput.n239 CSoutput.n124 4.5005
R23239 CSoutput.n140 CSoutput.n124 4.5005
R23240 CSoutput.n135 CSoutput.n119 4.5005
R23241 CSoutput.n135 CSoutput.n121 4.5005
R23242 CSoutput.n135 CSoutput.n118 4.5005
R23243 CSoutput.n135 CSoutput.n122 4.5005
R23244 CSoutput.n135 CSoutput.n117 4.5005
R23245 CSoutput.n135 CSoutput.t201 4.5005
R23246 CSoutput.n135 CSoutput.n116 4.5005
R23247 CSoutput.n135 CSoutput.n123 4.5005
R23248 CSoutput.n135 CSoutput.n124 4.5005
R23249 CSoutput.n133 CSoutput.n119 4.5005
R23250 CSoutput.n133 CSoutput.n121 4.5005
R23251 CSoutput.n133 CSoutput.n118 4.5005
R23252 CSoutput.n133 CSoutput.n122 4.5005
R23253 CSoutput.n133 CSoutput.n117 4.5005
R23254 CSoutput.n133 CSoutput.t201 4.5005
R23255 CSoutput.n133 CSoutput.n116 4.5005
R23256 CSoutput.n133 CSoutput.n123 4.5005
R23257 CSoutput.n133 CSoutput.n124 4.5005
R23258 CSoutput.n132 CSoutput.n119 4.5005
R23259 CSoutput.n132 CSoutput.n121 4.5005
R23260 CSoutput.n132 CSoutput.n118 4.5005
R23261 CSoutput.n132 CSoutput.n122 4.5005
R23262 CSoutput.n132 CSoutput.n117 4.5005
R23263 CSoutput.n132 CSoutput.t201 4.5005
R23264 CSoutput.n132 CSoutput.n116 4.5005
R23265 CSoutput.n132 CSoutput.n123 4.5005
R23266 CSoutput.n132 CSoutput.n124 4.5005
R23267 CSoutput.n261 CSoutput.n119 4.5005
R23268 CSoutput.n261 CSoutput.n121 4.5005
R23269 CSoutput.n261 CSoutput.n118 4.5005
R23270 CSoutput.n261 CSoutput.n122 4.5005
R23271 CSoutput.n261 CSoutput.n117 4.5005
R23272 CSoutput.n261 CSoutput.t201 4.5005
R23273 CSoutput.n261 CSoutput.n116 4.5005
R23274 CSoutput.n261 CSoutput.n123 4.5005
R23275 CSoutput.n261 CSoutput.n124 4.5005
R23276 CSoutput.n259 CSoutput.n119 4.5005
R23277 CSoutput.n259 CSoutput.n121 4.5005
R23278 CSoutput.n259 CSoutput.n118 4.5005
R23279 CSoutput.n259 CSoutput.n122 4.5005
R23280 CSoutput.n259 CSoutput.n117 4.5005
R23281 CSoutput.n259 CSoutput.t201 4.5005
R23282 CSoutput.n259 CSoutput.n116 4.5005
R23283 CSoutput.n259 CSoutput.n123 4.5005
R23284 CSoutput.n257 CSoutput.n119 4.5005
R23285 CSoutput.n257 CSoutput.n121 4.5005
R23286 CSoutput.n257 CSoutput.n118 4.5005
R23287 CSoutput.n257 CSoutput.n122 4.5005
R23288 CSoutput.n257 CSoutput.n117 4.5005
R23289 CSoutput.n257 CSoutput.t201 4.5005
R23290 CSoutput.n257 CSoutput.n116 4.5005
R23291 CSoutput.n257 CSoutput.n123 4.5005
R23292 CSoutput.n143 CSoutput.n119 4.5005
R23293 CSoutput.n143 CSoutput.n121 4.5005
R23294 CSoutput.n143 CSoutput.n118 4.5005
R23295 CSoutput.n143 CSoutput.n122 4.5005
R23296 CSoutput.n143 CSoutput.n117 4.5005
R23297 CSoutput.n143 CSoutput.t201 4.5005
R23298 CSoutput.n143 CSoutput.n116 4.5005
R23299 CSoutput.n143 CSoutput.n123 4.5005
R23300 CSoutput.n143 CSoutput.n124 4.5005
R23301 CSoutput.n142 CSoutput.n119 4.5005
R23302 CSoutput.n142 CSoutput.n121 4.5005
R23303 CSoutput.n142 CSoutput.n118 4.5005
R23304 CSoutput.n142 CSoutput.n122 4.5005
R23305 CSoutput.n142 CSoutput.n117 4.5005
R23306 CSoutput.n142 CSoutput.t201 4.5005
R23307 CSoutput.n142 CSoutput.n116 4.5005
R23308 CSoutput.n142 CSoutput.n123 4.5005
R23309 CSoutput.n142 CSoutput.n124 4.5005
R23310 CSoutput.n146 CSoutput.n119 4.5005
R23311 CSoutput.n146 CSoutput.n121 4.5005
R23312 CSoutput.n146 CSoutput.n118 4.5005
R23313 CSoutput.n146 CSoutput.n122 4.5005
R23314 CSoutput.n146 CSoutput.n117 4.5005
R23315 CSoutput.n146 CSoutput.t201 4.5005
R23316 CSoutput.n146 CSoutput.n116 4.5005
R23317 CSoutput.n146 CSoutput.n123 4.5005
R23318 CSoutput.n146 CSoutput.n124 4.5005
R23319 CSoutput.n145 CSoutput.n119 4.5005
R23320 CSoutput.n145 CSoutput.n121 4.5005
R23321 CSoutput.n145 CSoutput.n118 4.5005
R23322 CSoutput.n145 CSoutput.n122 4.5005
R23323 CSoutput.n145 CSoutput.n117 4.5005
R23324 CSoutput.n145 CSoutput.t201 4.5005
R23325 CSoutput.n145 CSoutput.n116 4.5005
R23326 CSoutput.n145 CSoutput.n123 4.5005
R23327 CSoutput.n145 CSoutput.n124 4.5005
R23328 CSoutput.n128 CSoutput.n119 4.5005
R23329 CSoutput.n128 CSoutput.n121 4.5005
R23330 CSoutput.n128 CSoutput.n118 4.5005
R23331 CSoutput.n128 CSoutput.n122 4.5005
R23332 CSoutput.n128 CSoutput.n117 4.5005
R23333 CSoutput.n128 CSoutput.t201 4.5005
R23334 CSoutput.n128 CSoutput.n116 4.5005
R23335 CSoutput.n128 CSoutput.n123 4.5005
R23336 CSoutput.n128 CSoutput.n124 4.5005
R23337 CSoutput.n264 CSoutput.n119 4.5005
R23338 CSoutput.n264 CSoutput.n121 4.5005
R23339 CSoutput.n264 CSoutput.n118 4.5005
R23340 CSoutput.n264 CSoutput.n122 4.5005
R23341 CSoutput.n264 CSoutput.n117 4.5005
R23342 CSoutput.n264 CSoutput.t201 4.5005
R23343 CSoutput.n264 CSoutput.n116 4.5005
R23344 CSoutput.n264 CSoutput.n123 4.5005
R23345 CSoutput.n264 CSoutput.n124 4.5005
R23346 CSoutput.n299 CSoutput.n287 4.10845
R23347 CSoutput.n113 CSoutput.n101 4.10845
R23348 CSoutput.n297 CSoutput.t46 4.06363
R23349 CSoutput.n297 CSoutput.t35 4.06363
R23350 CSoutput.n295 CSoutput.t177 4.06363
R23351 CSoutput.n295 CSoutput.t28 4.06363
R23352 CSoutput.n293 CSoutput.t23 4.06363
R23353 CSoutput.n293 CSoutput.t38 4.06363
R23354 CSoutput.n291 CSoutput.t41 4.06363
R23355 CSoutput.n291 CSoutput.t186 4.06363
R23356 CSoutput.n289 CSoutput.t12 4.06363
R23357 CSoutput.n289 CSoutput.t19 4.06363
R23358 CSoutput.n288 CSoutput.t1 4.06363
R23359 CSoutput.n288 CSoutput.t0 4.06363
R23360 CSoutput.n285 CSoutput.t24 4.06363
R23361 CSoutput.n285 CSoutput.t11 4.06363
R23362 CSoutput.n283 CSoutput.t40 4.06363
R23363 CSoutput.n283 CSoutput.t5 4.06363
R23364 CSoutput.n281 CSoutput.t16 4.06363
R23365 CSoutput.n281 CSoutput.t183 4.06363
R23366 CSoutput.n279 CSoutput.t18 4.06363
R23367 CSoutput.n279 CSoutput.t30 4.06363
R23368 CSoutput.n277 CSoutput.t34 4.06363
R23369 CSoutput.n277 CSoutput.t14 4.06363
R23370 CSoutput.n276 CSoutput.t171 4.06363
R23371 CSoutput.n276 CSoutput.t170 4.06363
R23372 CSoutput.n274 CSoutput.t182 4.06363
R23373 CSoutput.n274 CSoutput.t43 4.06363
R23374 CSoutput.n272 CSoutput.t27 4.06363
R23375 CSoutput.n272 CSoutput.t8 4.06363
R23376 CSoutput.n270 CSoutput.t39 4.06363
R23377 CSoutput.n270 CSoutput.t33 4.06363
R23378 CSoutput.n268 CSoutput.t175 4.06363
R23379 CSoutput.n268 CSoutput.t187 4.06363
R23380 CSoutput.n266 CSoutput.t169 4.06363
R23381 CSoutput.n266 CSoutput.t184 4.06363
R23382 CSoutput.n265 CSoutput.t7 4.06363
R23383 CSoutput.n265 CSoutput.t189 4.06363
R23384 CSoutput.n102 CSoutput.t45 4.06363
R23385 CSoutput.n102 CSoutput.t172 4.06363
R23386 CSoutput.n103 CSoutput.t36 4.06363
R23387 CSoutput.n103 CSoutput.t44 4.06363
R23388 CSoutput.n105 CSoutput.t22 4.06363
R23389 CSoutput.n105 CSoutput.t4 4.06363
R23390 CSoutput.n107 CSoutput.t37 4.06363
R23391 CSoutput.n107 CSoutput.t178 4.06363
R23392 CSoutput.n109 CSoutput.t47 4.06363
R23393 CSoutput.n109 CSoutput.t17 4.06363
R23394 CSoutput.n111 CSoutput.t29 4.06363
R23395 CSoutput.n111 CSoutput.t185 4.06363
R23396 CSoutput.n90 CSoutput.t20 4.06363
R23397 CSoutput.n90 CSoutput.t13 4.06363
R23398 CSoutput.n91 CSoutput.t31 4.06363
R23399 CSoutput.n91 CSoutput.t191 4.06363
R23400 CSoutput.n93 CSoutput.t9 4.06363
R23401 CSoutput.n93 CSoutput.t181 4.06363
R23402 CSoutput.n95 CSoutput.t176 4.06363
R23403 CSoutput.n95 CSoutput.t2 4.06363
R23404 CSoutput.n97 CSoutput.t25 4.06363
R23405 CSoutput.n97 CSoutput.t173 4.06363
R23406 CSoutput.n99 CSoutput.t42 4.06363
R23407 CSoutput.n99 CSoutput.t3 4.06363
R23408 CSoutput.n79 CSoutput.t10 4.06363
R23409 CSoutput.n79 CSoutput.t6 4.06363
R23410 CSoutput.n80 CSoutput.t179 4.06363
R23411 CSoutput.n80 CSoutput.t168 4.06363
R23412 CSoutput.n82 CSoutput.t180 4.06363
R23413 CSoutput.n82 CSoutput.t174 4.06363
R23414 CSoutput.n84 CSoutput.t32 4.06363
R23415 CSoutput.n84 CSoutput.t190 4.06363
R23416 CSoutput.n86 CSoutput.t21 4.06363
R23417 CSoutput.n86 CSoutput.t26 4.06363
R23418 CSoutput.n88 CSoutput.t188 4.06363
R23419 CSoutput.n88 CSoutput.t15 4.06363
R23420 CSoutput.n44 CSoutput.n43 3.79402
R23421 CSoutput.n49 CSoutput.n48 3.79402
R23422 CSoutput.n359 CSoutput.n339 3.72967
R23423 CSoutput.n419 CSoutput.n399 3.72967
R23424 CSoutput.n420 CSoutput.n360 3.71319
R23425 CSoutput.n421 CSoutput.n420 3.57343
R23426 CSoutput.n357 CSoutput.t96 2.82907
R23427 CSoutput.n357 CSoutput.t63 2.82907
R23428 CSoutput.n355 CSoutput.t166 2.82907
R23429 CSoutput.n355 CSoutput.t148 2.82907
R23430 CSoutput.n353 CSoutput.t70 2.82907
R23431 CSoutput.n353 CSoutput.t77 2.82907
R23432 CSoutput.n351 CSoutput.t61 2.82907
R23433 CSoutput.n351 CSoutput.t155 2.82907
R23434 CSoutput.n349 CSoutput.t117 2.82907
R23435 CSoutput.n349 CSoutput.t49 2.82907
R23436 CSoutput.n347 CSoutput.t159 2.82907
R23437 CSoutput.n347 CSoutput.t139 2.82907
R23438 CSoutput.n345 CSoutput.t97 2.82907
R23439 CSoutput.n345 CSoutput.t106 2.82907
R23440 CSoutput.n343 CSoutput.t48 2.82907
R23441 CSoutput.n343 CSoutput.t149 2.82907
R23442 CSoutput.n341 CSoutput.t140 2.82907
R23443 CSoutput.n341 CSoutput.t79 2.82907
R23444 CSoutput.n340 CSoutput.t64 2.82907
R23445 CSoutput.n340 CSoutput.t158 2.82907
R23446 CSoutput.n337 CSoutput.t167 2.82907
R23447 CSoutput.n337 CSoutput.t153 2.82907
R23448 CSoutput.n335 CSoutput.t152 2.82907
R23449 CSoutput.n335 CSoutput.t157 2.82907
R23450 CSoutput.n333 CSoutput.t78 2.82907
R23451 CSoutput.n333 CSoutput.t165 2.82907
R23452 CSoutput.n331 CSoutput.t57 2.82907
R23453 CSoutput.n331 CSoutput.t156 2.82907
R23454 CSoutput.n329 CSoutput.t72 2.82907
R23455 CSoutput.n329 CSoutput.t90 2.82907
R23456 CSoutput.n327 CSoutput.t88 2.82907
R23457 CSoutput.n327 CSoutput.t62 2.82907
R23458 CSoutput.n325 CSoutput.t103 2.82907
R23459 CSoutput.n325 CSoutput.t73 2.82907
R23460 CSoutput.n323 CSoutput.t74 2.82907
R23461 CSoutput.n323 CSoutput.t89 2.82907
R23462 CSoutput.n321 CSoutput.t87 2.82907
R23463 CSoutput.n321 CSoutput.t101 2.82907
R23464 CSoutput.n320 CSoutput.t102 2.82907
R23465 CSoutput.n320 CSoutput.t75 2.82907
R23466 CSoutput.n318 CSoutput.t116 2.82907
R23467 CSoutput.n318 CSoutput.t147 2.82907
R23468 CSoutput.n316 CSoutput.t124 2.82907
R23469 CSoutput.n316 CSoutput.t163 2.82907
R23470 CSoutput.n314 CSoutput.t65 2.82907
R23471 CSoutput.n314 CSoutput.t81 2.82907
R23472 CSoutput.n312 CSoutput.t107 2.82907
R23473 CSoutput.n312 CSoutput.t138 2.82907
R23474 CSoutput.n310 CSoutput.t128 2.82907
R23475 CSoutput.n310 CSoutput.t92 2.82907
R23476 CSoutput.n308 CSoutput.t54 2.82907
R23477 CSoutput.n308 CSoutput.t111 2.82907
R23478 CSoutput.n306 CSoutput.t91 2.82907
R23479 CSoutput.n306 CSoutput.t104 2.82907
R23480 CSoutput.n304 CSoutput.t105 2.82907
R23481 CSoutput.n304 CSoutput.t146 2.82907
R23482 CSoutput.n302 CSoutput.t123 2.82907
R23483 CSoutput.n302 CSoutput.t50 2.82907
R23484 CSoutput.n301 CSoutput.t143 2.82907
R23485 CSoutput.n301 CSoutput.t66 2.82907
R23486 CSoutput.n400 CSoutput.t134 2.82907
R23487 CSoutput.n400 CSoutput.t154 2.82907
R23488 CSoutput.n401 CSoutput.t162 2.82907
R23489 CSoutput.n401 CSoutput.t122 2.82907
R23490 CSoutput.n403 CSoutput.t127 2.82907
R23491 CSoutput.n403 CSoutput.t144 2.82907
R23492 CSoutput.n405 CSoutput.t68 2.82907
R23493 CSoutput.n405 CSoutput.t114 2.82907
R23494 CSoutput.n407 CSoutput.t121 2.82907
R23495 CSoutput.n407 CSoutput.t135 2.82907
R23496 CSoutput.n409 CSoutput.t145 2.82907
R23497 CSoutput.n409 CSoutput.t126 2.82907
R23498 CSoutput.n411 CSoutput.t131 2.82907
R23499 CSoutput.n411 CSoutput.t151 2.82907
R23500 CSoutput.n413 CSoutput.t69 2.82907
R23501 CSoutput.n413 CSoutput.t80 2.82907
R23502 CSoutput.n415 CSoutput.t141 2.82907
R23503 CSoutput.n415 CSoutput.t160 2.82907
R23504 CSoutput.n417 CSoutput.t51 2.82907
R23505 CSoutput.n417 CSoutput.t82 2.82907
R23506 CSoutput.n380 CSoutput.t99 2.82907
R23507 CSoutput.n380 CSoutput.t118 2.82907
R23508 CSoutput.n381 CSoutput.t119 2.82907
R23509 CSoutput.n381 CSoutput.t108 2.82907
R23510 CSoutput.n383 CSoutput.t109 2.82907
R23511 CSoutput.n383 CSoutput.t100 2.82907
R23512 CSoutput.n385 CSoutput.t93 2.82907
R23513 CSoutput.n385 CSoutput.t85 2.82907
R23514 CSoutput.n387 CSoutput.t86 2.82907
R23515 CSoutput.n387 CSoutput.t110 2.82907
R23516 CSoutput.n389 CSoutput.t112 2.82907
R23517 CSoutput.n389 CSoutput.t52 2.82907
R23518 CSoutput.n391 CSoutput.t53 2.82907
R23519 CSoutput.n391 CSoutput.t76 2.82907
R23520 CSoutput.n393 CSoutput.t83 2.82907
R23521 CSoutput.n393 CSoutput.t71 2.82907
R23522 CSoutput.n395 CSoutput.t67 2.82907
R23523 CSoutput.n395 CSoutput.t58 2.82907
R23524 CSoutput.n397 CSoutput.t59 2.82907
R23525 CSoutput.n397 CSoutput.t84 2.82907
R23526 CSoutput.n361 CSoutput.t113 2.82907
R23527 CSoutput.n361 CSoutput.t56 2.82907
R23528 CSoutput.n362 CSoutput.t95 2.82907
R23529 CSoutput.n362 CSoutput.t150 2.82907
R23530 CSoutput.n364 CSoutput.t60 2.82907
R23531 CSoutput.n364 CSoutput.t130 2.82907
R23532 CSoutput.n366 CSoutput.t129 2.82907
R23533 CSoutput.n366 CSoutput.t115 2.82907
R23534 CSoutput.n368 CSoutput.t133 2.82907
R23535 CSoutput.n368 CSoutput.t98 2.82907
R23536 CSoutput.n370 CSoutput.t125 2.82907
R23537 CSoutput.n370 CSoutput.t142 2.82907
R23538 CSoutput.n372 CSoutput.t164 2.82907
R23539 CSoutput.n372 CSoutput.t132 2.82907
R23540 CSoutput.n374 CSoutput.t137 2.82907
R23541 CSoutput.n374 CSoutput.t136 2.82907
R23542 CSoutput.n376 CSoutput.t120 2.82907
R23543 CSoutput.n376 CSoutput.t55 2.82907
R23544 CSoutput.n378 CSoutput.t94 2.82907
R23545 CSoutput.n378 CSoutput.t161 2.82907
R23546 CSoutput.n300 CSoutput.n114 2.78353
R23547 CSoutput.n75 CSoutput.n1 2.45513
R23548 CSoutput.n205 CSoutput.n203 2.251
R23549 CSoutput.n205 CSoutput.n202 2.251
R23550 CSoutput.n205 CSoutput.n201 2.251
R23551 CSoutput.n205 CSoutput.n200 2.251
R23552 CSoutput.n174 CSoutput.n173 2.251
R23553 CSoutput.n174 CSoutput.n172 2.251
R23554 CSoutput.n174 CSoutput.n171 2.251
R23555 CSoutput.n174 CSoutput.n170 2.251
R23556 CSoutput.n247 CSoutput.n246 2.251
R23557 CSoutput.n212 CSoutput.n210 2.251
R23558 CSoutput.n212 CSoutput.n209 2.251
R23559 CSoutput.n212 CSoutput.n208 2.251
R23560 CSoutput.n230 CSoutput.n212 2.251
R23561 CSoutput.n218 CSoutput.n217 2.251
R23562 CSoutput.n218 CSoutput.n216 2.251
R23563 CSoutput.n218 CSoutput.n215 2.251
R23564 CSoutput.n218 CSoutput.n214 2.251
R23565 CSoutput.n244 CSoutput.n184 2.251
R23566 CSoutput.n239 CSoutput.n237 2.251
R23567 CSoutput.n239 CSoutput.n236 2.251
R23568 CSoutput.n239 CSoutput.n235 2.251
R23569 CSoutput.n239 CSoutput.n234 2.251
R23570 CSoutput.n140 CSoutput.n139 2.251
R23571 CSoutput.n140 CSoutput.n138 2.251
R23572 CSoutput.n140 CSoutput.n137 2.251
R23573 CSoutput.n140 CSoutput.n136 2.251
R23574 CSoutput.n257 CSoutput.n256 2.251
R23575 CSoutput.n174 CSoutput.n154 2.2505
R23576 CSoutput.n169 CSoutput.n154 2.2505
R23577 CSoutput.n167 CSoutput.n154 2.2505
R23578 CSoutput.n166 CSoutput.n154 2.2505
R23579 CSoutput.n251 CSoutput.n154 2.2505
R23580 CSoutput.n249 CSoutput.n154 2.2505
R23581 CSoutput.n247 CSoutput.n154 2.2505
R23582 CSoutput.n177 CSoutput.n154 2.2505
R23583 CSoutput.n176 CSoutput.n154 2.2505
R23584 CSoutput.n180 CSoutput.n154 2.2505
R23585 CSoutput.n179 CSoutput.n154 2.2505
R23586 CSoutput.n162 CSoutput.n154 2.2505
R23587 CSoutput.n254 CSoutput.n154 2.2505
R23588 CSoutput.n254 CSoutput.n253 2.2505
R23589 CSoutput.n218 CSoutput.n189 2.2505
R23590 CSoutput.n199 CSoutput.n189 2.2505
R23591 CSoutput.n220 CSoutput.n189 2.2505
R23592 CSoutput.n198 CSoutput.n189 2.2505
R23593 CSoutput.n222 CSoutput.n189 2.2505
R23594 CSoutput.n189 CSoutput.n183 2.2505
R23595 CSoutput.n244 CSoutput.n189 2.2505
R23596 CSoutput.n242 CSoutput.n189 2.2505
R23597 CSoutput.n224 CSoutput.n189 2.2505
R23598 CSoutput.n196 CSoutput.n189 2.2505
R23599 CSoutput.n226 CSoutput.n189 2.2505
R23600 CSoutput.n195 CSoutput.n189 2.2505
R23601 CSoutput.n240 CSoutput.n189 2.2505
R23602 CSoutput.n240 CSoutput.n193 2.2505
R23603 CSoutput.n140 CSoutput.n120 2.2505
R23604 CSoutput.n135 CSoutput.n120 2.2505
R23605 CSoutput.n133 CSoutput.n120 2.2505
R23606 CSoutput.n132 CSoutput.n120 2.2505
R23607 CSoutput.n261 CSoutput.n120 2.2505
R23608 CSoutput.n259 CSoutput.n120 2.2505
R23609 CSoutput.n257 CSoutput.n120 2.2505
R23610 CSoutput.n143 CSoutput.n120 2.2505
R23611 CSoutput.n142 CSoutput.n120 2.2505
R23612 CSoutput.n146 CSoutput.n120 2.2505
R23613 CSoutput.n145 CSoutput.n120 2.2505
R23614 CSoutput.n128 CSoutput.n120 2.2505
R23615 CSoutput.n264 CSoutput.n120 2.2505
R23616 CSoutput.n264 CSoutput.n263 2.2505
R23617 CSoutput.n182 CSoutput.n175 2.25024
R23618 CSoutput.n182 CSoutput.n168 2.25024
R23619 CSoutput.n250 CSoutput.n182 2.25024
R23620 CSoutput.n182 CSoutput.n178 2.25024
R23621 CSoutput.n182 CSoutput.n181 2.25024
R23622 CSoutput.n182 CSoutput.n149 2.25024
R23623 CSoutput.n232 CSoutput.n229 2.25024
R23624 CSoutput.n232 CSoutput.n228 2.25024
R23625 CSoutput.n232 CSoutput.n227 2.25024
R23626 CSoutput.n232 CSoutput.n194 2.25024
R23627 CSoutput.n232 CSoutput.n231 2.25024
R23628 CSoutput.n233 CSoutput.n232 2.25024
R23629 CSoutput.n148 CSoutput.n141 2.25024
R23630 CSoutput.n148 CSoutput.n134 2.25024
R23631 CSoutput.n260 CSoutput.n148 2.25024
R23632 CSoutput.n148 CSoutput.n144 2.25024
R23633 CSoutput.n148 CSoutput.n147 2.25024
R23634 CSoutput.n148 CSoutput.n115 2.25024
R23635 CSoutput.n249 CSoutput.n159 1.50111
R23636 CSoutput.n197 CSoutput.n183 1.50111
R23637 CSoutput.n259 CSoutput.n125 1.50111
R23638 CSoutput.n205 CSoutput.n204 1.501
R23639 CSoutput.n212 CSoutput.n211 1.501
R23640 CSoutput.n239 CSoutput.n238 1.501
R23641 CSoutput.n253 CSoutput.n164 1.12536
R23642 CSoutput.n253 CSoutput.n165 1.12536
R23643 CSoutput.n253 CSoutput.n252 1.12536
R23644 CSoutput.n213 CSoutput.n193 1.12536
R23645 CSoutput.n219 CSoutput.n193 1.12536
R23646 CSoutput.n221 CSoutput.n193 1.12536
R23647 CSoutput.n263 CSoutput.n130 1.12536
R23648 CSoutput.n263 CSoutput.n131 1.12536
R23649 CSoutput.n263 CSoutput.n262 1.12536
R23650 CSoutput.n253 CSoutput.n160 1.12536
R23651 CSoutput.n253 CSoutput.n161 1.12536
R23652 CSoutput.n253 CSoutput.n163 1.12536
R23653 CSoutput.n243 CSoutput.n193 1.12536
R23654 CSoutput.n223 CSoutput.n193 1.12536
R23655 CSoutput.n225 CSoutput.n193 1.12536
R23656 CSoutput.n263 CSoutput.n126 1.12536
R23657 CSoutput.n263 CSoutput.n127 1.12536
R23658 CSoutput.n263 CSoutput.n129 1.12536
R23659 CSoutput.n31 CSoutput.n30 0.669944
R23660 CSoutput.n62 CSoutput.n61 0.669944
R23661 CSoutput.n344 CSoutput.n342 0.573776
R23662 CSoutput.n346 CSoutput.n344 0.573776
R23663 CSoutput.n348 CSoutput.n346 0.573776
R23664 CSoutput.n350 CSoutput.n348 0.573776
R23665 CSoutput.n352 CSoutput.n350 0.573776
R23666 CSoutput.n354 CSoutput.n352 0.573776
R23667 CSoutput.n356 CSoutput.n354 0.573776
R23668 CSoutput.n358 CSoutput.n356 0.573776
R23669 CSoutput.n324 CSoutput.n322 0.573776
R23670 CSoutput.n326 CSoutput.n324 0.573776
R23671 CSoutput.n328 CSoutput.n326 0.573776
R23672 CSoutput.n330 CSoutput.n328 0.573776
R23673 CSoutput.n332 CSoutput.n330 0.573776
R23674 CSoutput.n334 CSoutput.n332 0.573776
R23675 CSoutput.n336 CSoutput.n334 0.573776
R23676 CSoutput.n338 CSoutput.n336 0.573776
R23677 CSoutput.n305 CSoutput.n303 0.573776
R23678 CSoutput.n307 CSoutput.n305 0.573776
R23679 CSoutput.n309 CSoutput.n307 0.573776
R23680 CSoutput.n311 CSoutput.n309 0.573776
R23681 CSoutput.n313 CSoutput.n311 0.573776
R23682 CSoutput.n315 CSoutput.n313 0.573776
R23683 CSoutput.n317 CSoutput.n315 0.573776
R23684 CSoutput.n319 CSoutput.n317 0.573776
R23685 CSoutput.n418 CSoutput.n416 0.573776
R23686 CSoutput.n416 CSoutput.n414 0.573776
R23687 CSoutput.n414 CSoutput.n412 0.573776
R23688 CSoutput.n412 CSoutput.n410 0.573776
R23689 CSoutput.n410 CSoutput.n408 0.573776
R23690 CSoutput.n408 CSoutput.n406 0.573776
R23691 CSoutput.n406 CSoutput.n404 0.573776
R23692 CSoutput.n404 CSoutput.n402 0.573776
R23693 CSoutput.n398 CSoutput.n396 0.573776
R23694 CSoutput.n396 CSoutput.n394 0.573776
R23695 CSoutput.n394 CSoutput.n392 0.573776
R23696 CSoutput.n392 CSoutput.n390 0.573776
R23697 CSoutput.n390 CSoutput.n388 0.573776
R23698 CSoutput.n388 CSoutput.n386 0.573776
R23699 CSoutput.n386 CSoutput.n384 0.573776
R23700 CSoutput.n384 CSoutput.n382 0.573776
R23701 CSoutput.n379 CSoutput.n377 0.573776
R23702 CSoutput.n377 CSoutput.n375 0.573776
R23703 CSoutput.n375 CSoutput.n373 0.573776
R23704 CSoutput.n373 CSoutput.n371 0.573776
R23705 CSoutput.n371 CSoutput.n369 0.573776
R23706 CSoutput.n369 CSoutput.n367 0.573776
R23707 CSoutput.n367 CSoutput.n365 0.573776
R23708 CSoutput.n365 CSoutput.n363 0.573776
R23709 CSoutput.n421 CSoutput.n264 0.53442
R23710 CSoutput.n292 CSoutput.n290 0.358259
R23711 CSoutput.n294 CSoutput.n292 0.358259
R23712 CSoutput.n296 CSoutput.n294 0.358259
R23713 CSoutput.n298 CSoutput.n296 0.358259
R23714 CSoutput.n280 CSoutput.n278 0.358259
R23715 CSoutput.n282 CSoutput.n280 0.358259
R23716 CSoutput.n284 CSoutput.n282 0.358259
R23717 CSoutput.n286 CSoutput.n284 0.358259
R23718 CSoutput.n269 CSoutput.n267 0.358259
R23719 CSoutput.n271 CSoutput.n269 0.358259
R23720 CSoutput.n273 CSoutput.n271 0.358259
R23721 CSoutput.n275 CSoutput.n273 0.358259
R23722 CSoutput.n112 CSoutput.n110 0.358259
R23723 CSoutput.n110 CSoutput.n108 0.358259
R23724 CSoutput.n108 CSoutput.n106 0.358259
R23725 CSoutput.n106 CSoutput.n104 0.358259
R23726 CSoutput.n100 CSoutput.n98 0.358259
R23727 CSoutput.n98 CSoutput.n96 0.358259
R23728 CSoutput.n96 CSoutput.n94 0.358259
R23729 CSoutput.n94 CSoutput.n92 0.358259
R23730 CSoutput.n89 CSoutput.n87 0.358259
R23731 CSoutput.n87 CSoutput.n85 0.358259
R23732 CSoutput.n85 CSoutput.n83 0.358259
R23733 CSoutput.n83 CSoutput.n81 0.358259
R23734 CSoutput.n21 CSoutput.n20 0.169105
R23735 CSoutput.n21 CSoutput.n16 0.169105
R23736 CSoutput.n26 CSoutput.n16 0.169105
R23737 CSoutput.n27 CSoutput.n26 0.169105
R23738 CSoutput.n27 CSoutput.n14 0.169105
R23739 CSoutput.n32 CSoutput.n14 0.169105
R23740 CSoutput.n33 CSoutput.n32 0.169105
R23741 CSoutput.n34 CSoutput.n33 0.169105
R23742 CSoutput.n34 CSoutput.n12 0.169105
R23743 CSoutput.n39 CSoutput.n12 0.169105
R23744 CSoutput.n40 CSoutput.n39 0.169105
R23745 CSoutput.n40 CSoutput.n10 0.169105
R23746 CSoutput.n45 CSoutput.n10 0.169105
R23747 CSoutput.n46 CSoutput.n45 0.169105
R23748 CSoutput.n47 CSoutput.n46 0.169105
R23749 CSoutput.n47 CSoutput.n8 0.169105
R23750 CSoutput.n52 CSoutput.n8 0.169105
R23751 CSoutput.n53 CSoutput.n52 0.169105
R23752 CSoutput.n53 CSoutput.n6 0.169105
R23753 CSoutput.n58 CSoutput.n6 0.169105
R23754 CSoutput.n59 CSoutput.n58 0.169105
R23755 CSoutput.n60 CSoutput.n59 0.169105
R23756 CSoutput.n60 CSoutput.n4 0.169105
R23757 CSoutput.n66 CSoutput.n4 0.169105
R23758 CSoutput.n67 CSoutput.n66 0.169105
R23759 CSoutput.n68 CSoutput.n67 0.169105
R23760 CSoutput.n68 CSoutput.n2 0.169105
R23761 CSoutput.n73 CSoutput.n2 0.169105
R23762 CSoutput.n74 CSoutput.n73 0.169105
R23763 CSoutput.n74 CSoutput.n0 0.169105
R23764 CSoutput.n78 CSoutput.n0 0.169105
R23765 CSoutput.n207 CSoutput.n206 0.0910737
R23766 CSoutput.n258 CSoutput.n255 0.0723685
R23767 CSoutput.n212 CSoutput.n207 0.0522944
R23768 CSoutput.n255 CSoutput.n254 0.0499135
R23769 CSoutput.n206 CSoutput.n205 0.0499135
R23770 CSoutput.n240 CSoutput.n239 0.0464294
R23771 CSoutput.n248 CSoutput.n245 0.0391444
R23772 CSoutput.n207 CSoutput.t210 0.023435
R23773 CSoutput.n255 CSoutput.t194 0.02262
R23774 CSoutput.n206 CSoutput.t206 0.02262
R23775 CSoutput CSoutput.n421 0.0052
R23776 CSoutput.n177 CSoutput.n160 0.00365111
R23777 CSoutput.n180 CSoutput.n161 0.00365111
R23778 CSoutput.n163 CSoutput.n162 0.00365111
R23779 CSoutput.n205 CSoutput.n164 0.00365111
R23780 CSoutput.n169 CSoutput.n165 0.00365111
R23781 CSoutput.n252 CSoutput.n166 0.00365111
R23782 CSoutput.n243 CSoutput.n242 0.00365111
R23783 CSoutput.n223 CSoutput.n196 0.00365111
R23784 CSoutput.n225 CSoutput.n195 0.00365111
R23785 CSoutput.n213 CSoutput.n212 0.00365111
R23786 CSoutput.n219 CSoutput.n199 0.00365111
R23787 CSoutput.n221 CSoutput.n198 0.00365111
R23788 CSoutput.n143 CSoutput.n126 0.00365111
R23789 CSoutput.n146 CSoutput.n127 0.00365111
R23790 CSoutput.n129 CSoutput.n128 0.00365111
R23791 CSoutput.n239 CSoutput.n130 0.00365111
R23792 CSoutput.n135 CSoutput.n131 0.00365111
R23793 CSoutput.n262 CSoutput.n132 0.00365111
R23794 CSoutput.n174 CSoutput.n164 0.00340054
R23795 CSoutput.n167 CSoutput.n165 0.00340054
R23796 CSoutput.n252 CSoutput.n251 0.00340054
R23797 CSoutput.n247 CSoutput.n160 0.00340054
R23798 CSoutput.n176 CSoutput.n161 0.00340054
R23799 CSoutput.n179 CSoutput.n163 0.00340054
R23800 CSoutput.n218 CSoutput.n213 0.00340054
R23801 CSoutput.n220 CSoutput.n219 0.00340054
R23802 CSoutput.n222 CSoutput.n221 0.00340054
R23803 CSoutput.n244 CSoutput.n243 0.00340054
R23804 CSoutput.n224 CSoutput.n223 0.00340054
R23805 CSoutput.n226 CSoutput.n225 0.00340054
R23806 CSoutput.n140 CSoutput.n130 0.00340054
R23807 CSoutput.n133 CSoutput.n131 0.00340054
R23808 CSoutput.n262 CSoutput.n261 0.00340054
R23809 CSoutput.n257 CSoutput.n126 0.00340054
R23810 CSoutput.n142 CSoutput.n127 0.00340054
R23811 CSoutput.n145 CSoutput.n129 0.00340054
R23812 CSoutput.n175 CSoutput.n169 0.00252698
R23813 CSoutput.n168 CSoutput.n166 0.00252698
R23814 CSoutput.n250 CSoutput.n249 0.00252698
R23815 CSoutput.n178 CSoutput.n176 0.00252698
R23816 CSoutput.n181 CSoutput.n179 0.00252698
R23817 CSoutput.n254 CSoutput.n149 0.00252698
R23818 CSoutput.n175 CSoutput.n174 0.00252698
R23819 CSoutput.n168 CSoutput.n167 0.00252698
R23820 CSoutput.n251 CSoutput.n250 0.00252698
R23821 CSoutput.n178 CSoutput.n177 0.00252698
R23822 CSoutput.n181 CSoutput.n180 0.00252698
R23823 CSoutput.n162 CSoutput.n149 0.00252698
R23824 CSoutput.n229 CSoutput.n199 0.00252698
R23825 CSoutput.n228 CSoutput.n198 0.00252698
R23826 CSoutput.n227 CSoutput.n183 0.00252698
R23827 CSoutput.n224 CSoutput.n194 0.00252698
R23828 CSoutput.n231 CSoutput.n226 0.00252698
R23829 CSoutput.n240 CSoutput.n233 0.00252698
R23830 CSoutput.n229 CSoutput.n218 0.00252698
R23831 CSoutput.n228 CSoutput.n220 0.00252698
R23832 CSoutput.n227 CSoutput.n222 0.00252698
R23833 CSoutput.n242 CSoutput.n194 0.00252698
R23834 CSoutput.n231 CSoutput.n196 0.00252698
R23835 CSoutput.n233 CSoutput.n195 0.00252698
R23836 CSoutput.n141 CSoutput.n135 0.00252698
R23837 CSoutput.n134 CSoutput.n132 0.00252698
R23838 CSoutput.n260 CSoutput.n259 0.00252698
R23839 CSoutput.n144 CSoutput.n142 0.00252698
R23840 CSoutput.n147 CSoutput.n145 0.00252698
R23841 CSoutput.n264 CSoutput.n115 0.00252698
R23842 CSoutput.n141 CSoutput.n140 0.00252698
R23843 CSoutput.n134 CSoutput.n133 0.00252698
R23844 CSoutput.n261 CSoutput.n260 0.00252698
R23845 CSoutput.n144 CSoutput.n143 0.00252698
R23846 CSoutput.n147 CSoutput.n146 0.00252698
R23847 CSoutput.n128 CSoutput.n115 0.00252698
R23848 CSoutput.n249 CSoutput.n248 0.0020275
R23849 CSoutput.n248 CSoutput.n247 0.0020275
R23850 CSoutput.n245 CSoutput.n183 0.0020275
R23851 CSoutput.n245 CSoutput.n244 0.0020275
R23852 CSoutput.n259 CSoutput.n258 0.0020275
R23853 CSoutput.n258 CSoutput.n257 0.0020275
R23854 CSoutput.n159 CSoutput.n158 0.00166668
R23855 CSoutput.n241 CSoutput.n197 0.00166668
R23856 CSoutput.n125 CSoutput.n124 0.00166668
R23857 CSoutput.n263 CSoutput.n125 0.00133328
R23858 CSoutput.n197 CSoutput.n193 0.00133328
R23859 CSoutput.n253 CSoutput.n159 0.00133328
R23860 CSoutput.n256 CSoutput.n148 0.001
R23861 CSoutput.n234 CSoutput.n148 0.001
R23862 CSoutput.n136 CSoutput.n116 0.001
R23863 CSoutput.n235 CSoutput.n116 0.001
R23864 CSoutput.n137 CSoutput.n117 0.001
R23865 CSoutput.n236 CSoutput.n117 0.001
R23866 CSoutput.n138 CSoutput.n118 0.001
R23867 CSoutput.n237 CSoutput.n118 0.001
R23868 CSoutput.n139 CSoutput.n119 0.001
R23869 CSoutput.n238 CSoutput.n119 0.001
R23870 CSoutput.n232 CSoutput.n184 0.001
R23871 CSoutput.n232 CSoutput.n230 0.001
R23872 CSoutput.n214 CSoutput.n185 0.001
R23873 CSoutput.n208 CSoutput.n185 0.001
R23874 CSoutput.n215 CSoutput.n186 0.001
R23875 CSoutput.n209 CSoutput.n186 0.001
R23876 CSoutput.n216 CSoutput.n187 0.001
R23877 CSoutput.n210 CSoutput.n187 0.001
R23878 CSoutput.n217 CSoutput.n188 0.001
R23879 CSoutput.n211 CSoutput.n188 0.001
R23880 CSoutput.n246 CSoutput.n182 0.001
R23881 CSoutput.n200 CSoutput.n182 0.001
R23882 CSoutput.n170 CSoutput.n150 0.001
R23883 CSoutput.n201 CSoutput.n150 0.001
R23884 CSoutput.n171 CSoutput.n151 0.001
R23885 CSoutput.n202 CSoutput.n151 0.001
R23886 CSoutput.n172 CSoutput.n152 0.001
R23887 CSoutput.n203 CSoutput.n152 0.001
R23888 CSoutput.n173 CSoutput.n153 0.001
R23889 CSoutput.n204 CSoutput.n153 0.001
R23890 CSoutput.n204 CSoutput.n154 0.001
R23891 CSoutput.n203 CSoutput.n155 0.001
R23892 CSoutput.n202 CSoutput.n156 0.001
R23893 CSoutput.n201 CSoutput.t196 0.001
R23894 CSoutput.n200 CSoutput.n157 0.001
R23895 CSoutput.n173 CSoutput.n155 0.001
R23896 CSoutput.n172 CSoutput.n156 0.001
R23897 CSoutput.n171 CSoutput.t196 0.001
R23898 CSoutput.n170 CSoutput.n157 0.001
R23899 CSoutput.n246 CSoutput.n158 0.001
R23900 CSoutput.n211 CSoutput.n189 0.001
R23901 CSoutput.n210 CSoutput.n190 0.001
R23902 CSoutput.n209 CSoutput.n191 0.001
R23903 CSoutput.n208 CSoutput.t200 0.001
R23904 CSoutput.n230 CSoutput.n192 0.001
R23905 CSoutput.n217 CSoutput.n190 0.001
R23906 CSoutput.n216 CSoutput.n191 0.001
R23907 CSoutput.n215 CSoutput.t200 0.001
R23908 CSoutput.n214 CSoutput.n192 0.001
R23909 CSoutput.n241 CSoutput.n184 0.001
R23910 CSoutput.n238 CSoutput.n120 0.001
R23911 CSoutput.n237 CSoutput.n121 0.001
R23912 CSoutput.n236 CSoutput.n122 0.001
R23913 CSoutput.n235 CSoutput.t201 0.001
R23914 CSoutput.n234 CSoutput.n123 0.001
R23915 CSoutput.n139 CSoutput.n121 0.001
R23916 CSoutput.n138 CSoutput.n122 0.001
R23917 CSoutput.n137 CSoutput.t201 0.001
R23918 CSoutput.n136 CSoutput.n123 0.001
R23919 CSoutput.n256 CSoutput.n124 0.001
R23920 a_n8300_8799.n142 a_n8300_8799.t109 490.524
R23921 a_n8300_8799.n153 a_n8300_8799.t45 490.524
R23922 a_n8300_8799.n165 a_n8300_8799.t93 490.524
R23923 a_n8300_8799.n108 a_n8300_8799.t85 490.524
R23924 a_n8300_8799.n119 a_n8300_8799.t92 490.524
R23925 a_n8300_8799.n131 a_n8300_8799.t94 490.524
R23926 a_n8300_8799.n33 a_n8300_8799.t47 484.3
R23927 a_n8300_8799.n148 a_n8300_8799.t46 464.166
R23928 a_n8300_8799.n147 a_n8300_8799.t96 464.166
R23929 a_n8300_8799.n138 a_n8300_8799.t57 464.166
R23930 a_n8300_8799.n146 a_n8300_8799.t49 464.166
R23931 a_n8300_8799.n145 a_n8300_8799.t100 464.166
R23932 a_n8300_8799.n139 a_n8300_8799.t73 464.166
R23933 a_n8300_8799.n144 a_n8300_8799.t58 464.166
R23934 a_n8300_8799.n143 a_n8300_8799.t113 464.166
R23935 a_n8300_8799.n140 a_n8300_8799.t84 464.166
R23936 a_n8300_8799.n141 a_n8300_8799.t60 464.166
R23937 a_n8300_8799.n42 a_n8300_8799.t53 484.3
R23938 a_n8300_8799.n159 a_n8300_8799.t52 464.166
R23939 a_n8300_8799.n158 a_n8300_8799.t108 464.166
R23940 a_n8300_8799.n149 a_n8300_8799.t62 464.166
R23941 a_n8300_8799.n157 a_n8300_8799.t56 464.166
R23942 a_n8300_8799.n156 a_n8300_8799.t110 464.166
R23943 a_n8300_8799.n150 a_n8300_8799.t82 464.166
R23944 a_n8300_8799.n155 a_n8300_8799.t65 464.166
R23945 a_n8300_8799.n154 a_n8300_8799.t48 464.166
R23946 a_n8300_8799.n151 a_n8300_8799.t91 464.166
R23947 a_n8300_8799.n152 a_n8300_8799.t66 464.166
R23948 a_n8300_8799.n51 a_n8300_8799.t81 484.3
R23949 a_n8300_8799.n171 a_n8300_8799.t95 464.166
R23950 a_n8300_8799.n170 a_n8300_8799.t55 464.166
R23951 a_n8300_8799.n161 a_n8300_8799.t106 464.166
R23952 a_n8300_8799.n169 a_n8300_8799.t69 464.166
R23953 a_n8300_8799.n168 a_n8300_8799.t101 464.166
R23954 a_n8300_8799.n162 a_n8300_8799.t59 464.166
R23955 a_n8300_8799.n167 a_n8300_8799.t87 464.166
R23956 a_n8300_8799.n166 a_n8300_8799.t51 464.166
R23957 a_n8300_8799.n163 a_n8300_8799.t78 464.166
R23958 a_n8300_8799.n164 a_n8300_8799.t64 464.166
R23959 a_n8300_8799.n107 a_n8300_8799.t107 464.166
R23960 a_n8300_8799.n106 a_n8300_8799.t61 464.166
R23961 a_n8300_8799.n109 a_n8300_8799.t83 464.166
R23962 a_n8300_8799.n105 a_n8300_8799.t103 464.166
R23963 a_n8300_8799.n110 a_n8300_8799.t104 464.166
R23964 a_n8300_8799.n111 a_n8300_8799.t72 464.166
R23965 a_n8300_8799.n104 a_n8300_8799.t90 464.166
R23966 a_n8300_8799.n112 a_n8300_8799.t102 464.166
R23967 a_n8300_8799.n103 a_n8300_8799.t70 464.166
R23968 a_n8300_8799.n113 a_n8300_8799.t71 464.166
R23969 a_n8300_8799.n118 a_n8300_8799.t115 464.166
R23970 a_n8300_8799.n117 a_n8300_8799.t67 464.166
R23971 a_n8300_8799.n120 a_n8300_8799.t89 464.166
R23972 a_n8300_8799.n116 a_n8300_8799.t112 464.166
R23973 a_n8300_8799.n121 a_n8300_8799.t114 464.166
R23974 a_n8300_8799.n122 a_n8300_8799.t79 464.166
R23975 a_n8300_8799.n115 a_n8300_8799.t99 464.166
R23976 a_n8300_8799.n123 a_n8300_8799.t111 464.166
R23977 a_n8300_8799.n114 a_n8300_8799.t75 464.166
R23978 a_n8300_8799.n124 a_n8300_8799.t76 464.166
R23979 a_n8300_8799.n130 a_n8300_8799.t63 464.166
R23980 a_n8300_8799.n129 a_n8300_8799.t77 464.166
R23981 a_n8300_8799.n132 a_n8300_8799.t50 464.166
R23982 a_n8300_8799.n128 a_n8300_8799.t86 464.166
R23983 a_n8300_8799.n133 a_n8300_8799.t74 464.166
R23984 a_n8300_8799.n134 a_n8300_8799.t98 464.166
R23985 a_n8300_8799.n127 a_n8300_8799.t68 464.166
R23986 a_n8300_8799.n135 a_n8300_8799.t105 464.166
R23987 a_n8300_8799.n126 a_n8300_8799.t54 464.166
R23988 a_n8300_8799.n136 a_n8300_8799.t44 464.166
R23989 a_n8300_8799.n41 a_n8300_8799.n40 75.3623
R23990 a_n8300_8799.n39 a_n8300_8799.n24 70.3058
R23991 a_n8300_8799.n24 a_n8300_8799.n38 70.1674
R23992 a_n8300_8799.n38 a_n8300_8799.n139 20.9683
R23993 a_n8300_8799.n37 a_n8300_8799.n25 75.0448
R23994 a_n8300_8799.n145 a_n8300_8799.n37 11.2134
R23995 a_n8300_8799.n36 a_n8300_8799.n25 80.4688
R23996 a_n8300_8799.n27 a_n8300_8799.n35 74.73
R23997 a_n8300_8799.n34 a_n8300_8799.n27 70.1674
R23998 a_n8300_8799.n148 a_n8300_8799.n34 20.9683
R23999 a_n8300_8799.n26 a_n8300_8799.n33 70.5844
R24000 a_n8300_8799.n50 a_n8300_8799.n49 75.3623
R24001 a_n8300_8799.n48 a_n8300_8799.n20 70.3058
R24002 a_n8300_8799.n20 a_n8300_8799.n47 70.1674
R24003 a_n8300_8799.n47 a_n8300_8799.n150 20.9683
R24004 a_n8300_8799.n46 a_n8300_8799.n21 75.0448
R24005 a_n8300_8799.n156 a_n8300_8799.n46 11.2134
R24006 a_n8300_8799.n45 a_n8300_8799.n21 80.4688
R24007 a_n8300_8799.n23 a_n8300_8799.n44 74.73
R24008 a_n8300_8799.n43 a_n8300_8799.n23 70.1674
R24009 a_n8300_8799.n159 a_n8300_8799.n43 20.9683
R24010 a_n8300_8799.n22 a_n8300_8799.n42 70.5844
R24011 a_n8300_8799.n59 a_n8300_8799.n58 75.3623
R24012 a_n8300_8799.n57 a_n8300_8799.n16 70.3058
R24013 a_n8300_8799.n16 a_n8300_8799.n56 70.1674
R24014 a_n8300_8799.n56 a_n8300_8799.n162 20.9683
R24015 a_n8300_8799.n55 a_n8300_8799.n17 75.0448
R24016 a_n8300_8799.n168 a_n8300_8799.n55 11.2134
R24017 a_n8300_8799.n54 a_n8300_8799.n17 80.4688
R24018 a_n8300_8799.n19 a_n8300_8799.n53 74.73
R24019 a_n8300_8799.n52 a_n8300_8799.n19 70.1674
R24020 a_n8300_8799.n171 a_n8300_8799.n52 20.9683
R24021 a_n8300_8799.n18 a_n8300_8799.n51 70.5844
R24022 a_n8300_8799.n12 a_n8300_8799.n68 70.5844
R24023 a_n8300_8799.n67 a_n8300_8799.n13 70.1674
R24024 a_n8300_8799.n67 a_n8300_8799.n103 20.9683
R24025 a_n8300_8799.n13 a_n8300_8799.n66 74.73
R24026 a_n8300_8799.n112 a_n8300_8799.n66 11.843
R24027 a_n8300_8799.n65 a_n8300_8799.n14 80.4688
R24028 a_n8300_8799.n65 a_n8300_8799.n104 0.365327
R24029 a_n8300_8799.n14 a_n8300_8799.n64 75.0448
R24030 a_n8300_8799.n63 a_n8300_8799.n15 70.1674
R24031 a_n8300_8799.n63 a_n8300_8799.n105 20.9683
R24032 a_n8300_8799.n15 a_n8300_8799.n62 70.3058
R24033 a_n8300_8799.n109 a_n8300_8799.n62 20.6913
R24034 a_n8300_8799.n61 a_n8300_8799.n60 75.3623
R24035 a_n8300_8799.n8 a_n8300_8799.n77 70.5844
R24036 a_n8300_8799.n76 a_n8300_8799.n9 70.1674
R24037 a_n8300_8799.n76 a_n8300_8799.n114 20.9683
R24038 a_n8300_8799.n9 a_n8300_8799.n75 74.73
R24039 a_n8300_8799.n123 a_n8300_8799.n75 11.843
R24040 a_n8300_8799.n74 a_n8300_8799.n10 80.4688
R24041 a_n8300_8799.n74 a_n8300_8799.n115 0.365327
R24042 a_n8300_8799.n10 a_n8300_8799.n73 75.0448
R24043 a_n8300_8799.n72 a_n8300_8799.n11 70.1674
R24044 a_n8300_8799.n72 a_n8300_8799.n116 20.9683
R24045 a_n8300_8799.n11 a_n8300_8799.n71 70.3058
R24046 a_n8300_8799.n120 a_n8300_8799.n71 20.6913
R24047 a_n8300_8799.n70 a_n8300_8799.n69 75.3623
R24048 a_n8300_8799.n4 a_n8300_8799.n86 70.5844
R24049 a_n8300_8799.n85 a_n8300_8799.n5 70.1674
R24050 a_n8300_8799.n85 a_n8300_8799.n126 20.9683
R24051 a_n8300_8799.n5 a_n8300_8799.n84 74.73
R24052 a_n8300_8799.n135 a_n8300_8799.n84 11.843
R24053 a_n8300_8799.n83 a_n8300_8799.n6 80.4688
R24054 a_n8300_8799.n83 a_n8300_8799.n127 0.365327
R24055 a_n8300_8799.n6 a_n8300_8799.n82 75.0448
R24056 a_n8300_8799.n81 a_n8300_8799.n7 70.1674
R24057 a_n8300_8799.n81 a_n8300_8799.n128 20.9683
R24058 a_n8300_8799.n7 a_n8300_8799.n80 70.3058
R24059 a_n8300_8799.n132 a_n8300_8799.n80 20.6913
R24060 a_n8300_8799.n79 a_n8300_8799.n78 75.3623
R24061 a_n8300_8799.n28 a_n8300_8799.n87 98.9633
R24062 a_n8300_8799.n31 a_n8300_8799.n176 98.9631
R24063 a_n8300_8799.n31 a_n8300_8799.n177 98.6055
R24064 a_n8300_8799.n31 a_n8300_8799.n178 98.6055
R24065 a_n8300_8799.n32 a_n8300_8799.n179 98.6055
R24066 a_n8300_8799.n32 a_n8300_8799.n180 98.6055
R24067 a_n8300_8799.n30 a_n8300_8799.n92 98.6055
R24068 a_n8300_8799.n30 a_n8300_8799.n91 98.6055
R24069 a_n8300_8799.n29 a_n8300_8799.n90 98.6055
R24070 a_n8300_8799.n29 a_n8300_8799.n89 98.6055
R24071 a_n8300_8799.n28 a_n8300_8799.n88 98.6055
R24072 a_n8300_8799.n182 a_n8300_8799.n181 98.6054
R24073 a_n8300_8799.n3 a_n8300_8799.n93 81.4626
R24074 a_n8300_8799.n1 a_n8300_8799.n99 81.4626
R24075 a_n8300_8799.n0 a_n8300_8799.n96 81.4626
R24076 a_n8300_8799.n2 a_n8300_8799.n101 80.9324
R24077 a_n8300_8799.n2 a_n8300_8799.n102 80.9324
R24078 a_n8300_8799.n3 a_n8300_8799.n95 80.9324
R24079 a_n8300_8799.n3 a_n8300_8799.n94 80.9324
R24080 a_n8300_8799.n1 a_n8300_8799.n100 80.9324
R24081 a_n8300_8799.n1 a_n8300_8799.n98 80.9324
R24082 a_n8300_8799.n0 a_n8300_8799.n97 80.9324
R24083 a_n8300_8799.n34 a_n8300_8799.n147 20.9683
R24084 a_n8300_8799.n146 a_n8300_8799.n145 48.2005
R24085 a_n8300_8799.n144 a_n8300_8799.n38 20.9683
R24086 a_n8300_8799.n141 a_n8300_8799.n140 48.2005
R24087 a_n8300_8799.n43 a_n8300_8799.n158 20.9683
R24088 a_n8300_8799.n157 a_n8300_8799.n156 48.2005
R24089 a_n8300_8799.n155 a_n8300_8799.n47 20.9683
R24090 a_n8300_8799.n152 a_n8300_8799.n151 48.2005
R24091 a_n8300_8799.n52 a_n8300_8799.n170 20.9683
R24092 a_n8300_8799.n169 a_n8300_8799.n168 48.2005
R24093 a_n8300_8799.n167 a_n8300_8799.n56 20.9683
R24094 a_n8300_8799.n164 a_n8300_8799.n163 48.2005
R24095 a_n8300_8799.n107 a_n8300_8799.n106 48.2005
R24096 a_n8300_8799.n110 a_n8300_8799.n63 20.9683
R24097 a_n8300_8799.n111 a_n8300_8799.n104 48.2005
R24098 a_n8300_8799.n113 a_n8300_8799.n67 20.9683
R24099 a_n8300_8799.n118 a_n8300_8799.n117 48.2005
R24100 a_n8300_8799.n121 a_n8300_8799.n72 20.9683
R24101 a_n8300_8799.n122 a_n8300_8799.n115 48.2005
R24102 a_n8300_8799.n124 a_n8300_8799.n76 20.9683
R24103 a_n8300_8799.n130 a_n8300_8799.n129 48.2005
R24104 a_n8300_8799.n133 a_n8300_8799.n81 20.9683
R24105 a_n8300_8799.n134 a_n8300_8799.n127 48.2005
R24106 a_n8300_8799.n136 a_n8300_8799.n85 20.9683
R24107 a_n8300_8799.n36 a_n8300_8799.n138 47.835
R24108 a_n8300_8799.n39 a_n8300_8799.n143 20.6913
R24109 a_n8300_8799.n45 a_n8300_8799.n149 47.835
R24110 a_n8300_8799.n48 a_n8300_8799.n154 20.6913
R24111 a_n8300_8799.n54 a_n8300_8799.n161 47.835
R24112 a_n8300_8799.n57 a_n8300_8799.n166 20.6913
R24113 a_n8300_8799.n105 a_n8300_8799.n62 21.4216
R24114 a_n8300_8799.n116 a_n8300_8799.n71 21.4216
R24115 a_n8300_8799.n128 a_n8300_8799.n80 21.4216
R24116 a_n8300_8799.t88 a_n8300_8799.n68 484.3
R24117 a_n8300_8799.t97 a_n8300_8799.n77 484.3
R24118 a_n8300_8799.t80 a_n8300_8799.n86 484.3
R24119 a_n8300_8799.n61 a_n8300_8799.n108 45.0871
R24120 a_n8300_8799.n70 a_n8300_8799.n119 45.0871
R24121 a_n8300_8799.n79 a_n8300_8799.n131 45.0871
R24122 a_n8300_8799.n41 a_n8300_8799.n142 45.0871
R24123 a_n8300_8799.n50 a_n8300_8799.n153 45.0871
R24124 a_n8300_8799.n59 a_n8300_8799.n165 45.0871
R24125 a_n8300_8799.n181 a_n8300_8799.n175 34.1489
R24126 a_n8300_8799.n2 a_n8300_8799.n1 33.5285
R24127 a_n8300_8799.n35 a_n8300_8799.n138 11.843
R24128 a_n8300_8799.n143 a_n8300_8799.n40 36.139
R24129 a_n8300_8799.n44 a_n8300_8799.n149 11.843
R24130 a_n8300_8799.n154 a_n8300_8799.n49 36.139
R24131 a_n8300_8799.n53 a_n8300_8799.n161 11.843
R24132 a_n8300_8799.n166 a_n8300_8799.n58 36.139
R24133 a_n8300_8799.n109 a_n8300_8799.n60 36.139
R24134 a_n8300_8799.n103 a_n8300_8799.n66 34.4824
R24135 a_n8300_8799.n120 a_n8300_8799.n69 36.139
R24136 a_n8300_8799.n114 a_n8300_8799.n75 34.4824
R24137 a_n8300_8799.n132 a_n8300_8799.n78 36.139
R24138 a_n8300_8799.n126 a_n8300_8799.n84 34.4824
R24139 a_n8300_8799.n37 a_n8300_8799.n139 35.3134
R24140 a_n8300_8799.n46 a_n8300_8799.n150 35.3134
R24141 a_n8300_8799.n55 a_n8300_8799.n162 35.3134
R24142 a_n8300_8799.n64 a_n8300_8799.n110 35.3134
R24143 a_n8300_8799.n111 a_n8300_8799.n64 11.2134
R24144 a_n8300_8799.n73 a_n8300_8799.n121 35.3134
R24145 a_n8300_8799.n122 a_n8300_8799.n73 11.2134
R24146 a_n8300_8799.n82 a_n8300_8799.n133 35.3134
R24147 a_n8300_8799.n134 a_n8300_8799.n82 11.2134
R24148 a_n8300_8799.n147 a_n8300_8799.n35 34.4824
R24149 a_n8300_8799.n40 a_n8300_8799.n140 10.5784
R24150 a_n8300_8799.n158 a_n8300_8799.n44 34.4824
R24151 a_n8300_8799.n49 a_n8300_8799.n151 10.5784
R24152 a_n8300_8799.n170 a_n8300_8799.n53 34.4824
R24153 a_n8300_8799.n58 a_n8300_8799.n163 10.5784
R24154 a_n8300_8799.n60 a_n8300_8799.n106 10.5784
R24155 a_n8300_8799.n69 a_n8300_8799.n117 10.5784
R24156 a_n8300_8799.n78 a_n8300_8799.n129 10.5784
R24157 a_n8300_8799.n175 a_n8300_8799.n30 20.7404
R24158 a_n8300_8799.n142 a_n8300_8799.n141 14.1472
R24159 a_n8300_8799.n153 a_n8300_8799.n152 14.1472
R24160 a_n8300_8799.n165 a_n8300_8799.n164 14.1472
R24161 a_n8300_8799.n108 a_n8300_8799.n107 14.1472
R24162 a_n8300_8799.n119 a_n8300_8799.n118 14.1472
R24163 a_n8300_8799.n131 a_n8300_8799.n130 14.1472
R24164 a_n8300_8799.n174 a_n8300_8799.n3 12.3339
R24165 a_n8300_8799.n175 a_n8300_8799.n174 11.4887
R24166 a_n8300_8799.n160 a_n8300_8799.n26 9.01755
R24167 a_n8300_8799.n125 a_n8300_8799.n12 9.01755
R24168 a_n8300_8799.n173 a_n8300_8799.n137 7.21326
R24169 a_n8300_8799.n173 a_n8300_8799.n172 6.79371
R24170 a_n8300_8799.n160 a_n8300_8799.n22 4.90959
R24171 a_n8300_8799.n172 a_n8300_8799.n18 4.90959
R24172 a_n8300_8799.n125 a_n8300_8799.n8 4.90959
R24173 a_n8300_8799.n137 a_n8300_8799.n4 4.90959
R24174 a_n8300_8799.n172 a_n8300_8799.n160 4.10845
R24175 a_n8300_8799.n137 a_n8300_8799.n125 4.10845
R24176 a_n8300_8799.n176 a_n8300_8799.t34 3.61217
R24177 a_n8300_8799.n176 a_n8300_8799.t29 3.61217
R24178 a_n8300_8799.n177 a_n8300_8799.t25 3.61217
R24179 a_n8300_8799.n177 a_n8300_8799.t18 3.61217
R24180 a_n8300_8799.n178 a_n8300_8799.t36 3.61217
R24181 a_n8300_8799.n178 a_n8300_8799.t14 3.61217
R24182 a_n8300_8799.n179 a_n8300_8799.t30 3.61217
R24183 a_n8300_8799.n179 a_n8300_8799.t24 3.61217
R24184 a_n8300_8799.n180 a_n8300_8799.t20 3.61217
R24185 a_n8300_8799.n180 a_n8300_8799.t31 3.61217
R24186 a_n8300_8799.n92 a_n8300_8799.t33 3.61217
R24187 a_n8300_8799.n92 a_n8300_8799.t16 3.61217
R24188 a_n8300_8799.n91 a_n8300_8799.t32 3.61217
R24189 a_n8300_8799.n91 a_n8300_8799.t22 3.61217
R24190 a_n8300_8799.n90 a_n8300_8799.t23 3.61217
R24191 a_n8300_8799.n90 a_n8300_8799.t15 3.61217
R24192 a_n8300_8799.n89 a_n8300_8799.t19 3.61217
R24193 a_n8300_8799.n89 a_n8300_8799.t17 3.61217
R24194 a_n8300_8799.n88 a_n8300_8799.t35 3.61217
R24195 a_n8300_8799.n88 a_n8300_8799.t27 3.61217
R24196 a_n8300_8799.n87 a_n8300_8799.t28 3.61217
R24197 a_n8300_8799.n87 a_n8300_8799.t21 3.61217
R24198 a_n8300_8799.t13 a_n8300_8799.n182 3.61217
R24199 a_n8300_8799.n182 a_n8300_8799.t26 3.61217
R24200 a_n8300_8799.n174 a_n8300_8799.n173 3.4105
R24201 a_n8300_8799.n101 a_n8300_8799.t11 2.82907
R24202 a_n8300_8799.n101 a_n8300_8799.t42 2.82907
R24203 a_n8300_8799.n102 a_n8300_8799.t6 2.82907
R24204 a_n8300_8799.n102 a_n8300_8799.t3 2.82907
R24205 a_n8300_8799.n95 a_n8300_8799.t10 2.82907
R24206 a_n8300_8799.n95 a_n8300_8799.t43 2.82907
R24207 a_n8300_8799.n94 a_n8300_8799.t38 2.82907
R24208 a_n8300_8799.n94 a_n8300_8799.t37 2.82907
R24209 a_n8300_8799.n93 a_n8300_8799.t8 2.82907
R24210 a_n8300_8799.n93 a_n8300_8799.t1 2.82907
R24211 a_n8300_8799.n99 a_n8300_8799.t39 2.82907
R24212 a_n8300_8799.n99 a_n8300_8799.t40 2.82907
R24213 a_n8300_8799.n100 a_n8300_8799.t12 2.82907
R24214 a_n8300_8799.n100 a_n8300_8799.t2 2.82907
R24215 a_n8300_8799.n98 a_n8300_8799.t41 2.82907
R24216 a_n8300_8799.n98 a_n8300_8799.t7 2.82907
R24217 a_n8300_8799.n97 a_n8300_8799.t0 2.82907
R24218 a_n8300_8799.n97 a_n8300_8799.t4 2.82907
R24219 a_n8300_8799.n96 a_n8300_8799.t5 2.82907
R24220 a_n8300_8799.n96 a_n8300_8799.t9 2.82907
R24221 a_n8300_8799.n33 a_n8300_8799.n148 22.3251
R24222 a_n8300_8799.n42 a_n8300_8799.n159 22.3251
R24223 a_n8300_8799.n51 a_n8300_8799.n171 22.3251
R24224 a_n8300_8799.n68 a_n8300_8799.n113 22.3251
R24225 a_n8300_8799.n77 a_n8300_8799.n124 22.3251
R24226 a_n8300_8799.n86 a_n8300_8799.n136 22.3251
R24227 a_n8300_8799.n36 a_n8300_8799.n146 0.365327
R24228 a_n8300_8799.n144 a_n8300_8799.n39 21.4216
R24229 a_n8300_8799.n45 a_n8300_8799.n157 0.365327
R24230 a_n8300_8799.n155 a_n8300_8799.n48 21.4216
R24231 a_n8300_8799.n54 a_n8300_8799.n169 0.365327
R24232 a_n8300_8799.n167 a_n8300_8799.n57 21.4216
R24233 a_n8300_8799.n112 a_n8300_8799.n65 47.835
R24234 a_n8300_8799.n123 a_n8300_8799.n74 47.835
R24235 a_n8300_8799.n135 a_n8300_8799.n83 47.835
R24236 a_n8300_8799.n3 a_n8300_8799.n2 1.59102
R24237 a_n8300_8799.n1 a_n8300_8799.n0 1.06084
R24238 a_n8300_8799.n27 a_n8300_8799.n25 0.758076
R24239 a_n8300_8799.n25 a_n8300_8799.n24 0.758076
R24240 a_n8300_8799.n41 a_n8300_8799.n24 0.758076
R24241 a_n8300_8799.n23 a_n8300_8799.n21 0.758076
R24242 a_n8300_8799.n21 a_n8300_8799.n20 0.758076
R24243 a_n8300_8799.n50 a_n8300_8799.n20 0.758076
R24244 a_n8300_8799.n19 a_n8300_8799.n17 0.758076
R24245 a_n8300_8799.n17 a_n8300_8799.n16 0.758076
R24246 a_n8300_8799.n59 a_n8300_8799.n16 0.758076
R24247 a_n8300_8799.n15 a_n8300_8799.n14 0.758076
R24248 a_n8300_8799.n14 a_n8300_8799.n13 0.758076
R24249 a_n8300_8799.n13 a_n8300_8799.n12 0.758076
R24250 a_n8300_8799.n11 a_n8300_8799.n10 0.758076
R24251 a_n8300_8799.n10 a_n8300_8799.n9 0.758076
R24252 a_n8300_8799.n9 a_n8300_8799.n8 0.758076
R24253 a_n8300_8799.n7 a_n8300_8799.n6 0.758076
R24254 a_n8300_8799.n6 a_n8300_8799.n5 0.758076
R24255 a_n8300_8799.n5 a_n8300_8799.n4 0.758076
R24256 a_n8300_8799.n32 a_n8300_8799.n31 0.716017
R24257 a_n8300_8799.n181 a_n8300_8799.n32 0.716017
R24258 a_n8300_8799.n30 a_n8300_8799.n29 0.716017
R24259 a_n8300_8799.n29 a_n8300_8799.n28 0.716017
R24260 a_n8300_8799.n79 a_n8300_8799.n7 0.568682
R24261 a_n8300_8799.n70 a_n8300_8799.n11 0.568682
R24262 a_n8300_8799.n61 a_n8300_8799.n15 0.568682
R24263 a_n8300_8799.n19 a_n8300_8799.n18 0.568682
R24264 a_n8300_8799.n23 a_n8300_8799.n22 0.568682
R24265 a_n8300_8799.n27 a_n8300_8799.n26 0.568682
R24266 plus.n61 plus.t11 251.488
R24267 plus.n12 plus.t14 251.488
R24268 plus.n100 plus.t1 243.97
R24269 plus.n96 plus.t23 231.093
R24270 plus.n47 plus.t6 231.093
R24271 plus.n100 plus.n99 223.454
R24272 plus.n102 plus.n101 223.454
R24273 plus.n60 plus.t5 187.445
R24274 plus.n65 plus.t21 187.445
R24275 plus.n71 plus.t20 187.445
R24276 plus.n56 plus.t16 187.445
R24277 plus.n54 plus.t17 187.445
R24278 plus.n83 plus.t13 187.445
R24279 plus.n89 plus.t15 187.445
R24280 plus.n50 plus.t10 187.445
R24281 plus.n1 plus.t12 187.445
R24282 plus.n40 plus.t8 187.445
R24283 plus.n34 plus.t7 187.445
R24284 plus.n5 plus.t19 187.445
R24285 plus.n7 plus.t18 187.445
R24286 plus.n22 plus.t24 187.445
R24287 plus.n16 plus.t22 187.445
R24288 plus.n11 plus.t9 187.445
R24289 plus.n97 plus.n96 161.3
R24290 plus.n95 plus.n49 161.3
R24291 plus.n94 plus.n93 161.3
R24292 plus.n92 plus.n91 161.3
R24293 plus.n90 plus.n51 161.3
R24294 plus.n88 plus.n87 161.3
R24295 plus.n86 plus.n52 161.3
R24296 plus.n85 plus.n84 161.3
R24297 plus.n82 plus.n53 161.3
R24298 plus.n81 plus.n80 161.3
R24299 plus.n79 plus.n78 161.3
R24300 plus.n77 plus.n55 161.3
R24301 plus.n76 plus.n75 161.3
R24302 plus.n74 plus.n73 161.3
R24303 plus.n72 plus.n57 161.3
R24304 plus.n70 plus.n69 161.3
R24305 plus.n68 plus.n58 161.3
R24306 plus.n67 plus.n66 161.3
R24307 plus.n64 plus.n59 161.3
R24308 plus.n63 plus.n62 161.3
R24309 plus.n14 plus.n13 161.3
R24310 plus.n15 plus.n10 161.3
R24311 plus.n18 plus.n17 161.3
R24312 plus.n19 plus.n9 161.3
R24313 plus.n21 plus.n20 161.3
R24314 plus.n23 plus.n8 161.3
R24315 plus.n25 plus.n24 161.3
R24316 plus.n27 plus.n26 161.3
R24317 plus.n28 plus.n6 161.3
R24318 plus.n30 plus.n29 161.3
R24319 plus.n32 plus.n31 161.3
R24320 plus.n33 plus.n4 161.3
R24321 plus.n36 plus.n35 161.3
R24322 plus.n37 plus.n3 161.3
R24323 plus.n39 plus.n38 161.3
R24324 plus.n41 plus.n2 161.3
R24325 plus.n43 plus.n42 161.3
R24326 plus.n45 plus.n44 161.3
R24327 plus.n46 plus.n0 161.3
R24328 plus.n48 plus.n47 161.3
R24329 plus.n64 plus.n63 56.5617
R24330 plus.n91 plus.n90 56.5617
R24331 plus.n42 plus.n41 56.5617
R24332 plus.n15 plus.n14 56.5617
R24333 plus.n73 plus.n72 56.5617
R24334 plus.n82 plus.n81 56.5617
R24335 plus.n33 plus.n32 56.5617
R24336 plus.n24 plus.n23 56.5617
R24337 plus.n95 plus.n94 48.3272
R24338 plus.n46 plus.n45 48.3272
R24339 plus.n70 plus.n58 44.4521
R24340 plus.n84 plus.n52 44.4521
R24341 plus.n35 plus.n3 44.4521
R24342 plus.n21 plus.n9 44.4521
R24343 plus.n62 plus.n61 43.0014
R24344 plus.n13 plus.n12 43.0014
R24345 plus.n77 plus.n76 40.577
R24346 plus.n78 plus.n77 40.577
R24347 plus.n29 plus.n28 40.577
R24348 plus.n28 plus.n27 40.577
R24349 plus.n61 plus.n60 39.4345
R24350 plus.n12 plus.n11 39.4345
R24351 plus.n66 plus.n58 36.702
R24352 plus.n88 plus.n52 36.702
R24353 plus.n39 plus.n3 36.702
R24354 plus.n17 plus.n9 36.702
R24355 plus.n98 plus.n97 33.3471
R24356 plus.n65 plus.n64 20.9036
R24357 plus.n90 plus.n89 20.9036
R24358 plus.n41 plus.n40 20.9036
R24359 plus.n16 plus.n15 20.9036
R24360 plus.n99 plus.t2 19.8005
R24361 plus.n99 plus.t4 19.8005
R24362 plus.n101 plus.t0 19.8005
R24363 plus.n101 plus.t3 19.8005
R24364 plus.n73 plus.n56 18.9362
R24365 plus.n81 plus.n54 18.9362
R24366 plus.n32 plus.n5 18.9362
R24367 plus.n24 plus.n7 18.9362
R24368 plus.n72 plus.n71 16.9689
R24369 plus.n83 plus.n82 16.9689
R24370 plus.n34 plus.n33 16.9689
R24371 plus.n23 plus.n22 16.9689
R24372 plus plus.n103 15.204
R24373 plus.n63 plus.n60 15.0015
R24374 plus.n91 plus.n50 15.0015
R24375 plus.n42 plus.n1 15.0015
R24376 plus.n14 plus.n11 15.0015
R24377 plus.n96 plus.n95 12.4157
R24378 plus.n47 plus.n46 12.4157
R24379 plus.n98 plus.n48 11.9418
R24380 plus.n94 plus.n50 9.59132
R24381 plus.n45 plus.n1 9.59132
R24382 plus.n71 plus.n70 7.62397
R24383 plus.n84 plus.n83 7.62397
R24384 plus.n35 plus.n34 7.62397
R24385 plus.n22 plus.n21 7.62397
R24386 plus.n76 plus.n56 5.65662
R24387 plus.n78 plus.n54 5.65662
R24388 plus.n29 plus.n5 5.65662
R24389 plus.n27 plus.n7 5.65662
R24390 plus.n103 plus.n102 5.40567
R24391 plus.n66 plus.n65 3.68928
R24392 plus.n89 plus.n88 3.68928
R24393 plus.n40 plus.n39 3.68928
R24394 plus.n17 plus.n16 3.68928
R24395 plus.n103 plus.n98 1.188
R24396 plus.n102 plus.n100 0.716017
R24397 plus.n62 plus.n59 0.189894
R24398 plus.n67 plus.n59 0.189894
R24399 plus.n68 plus.n67 0.189894
R24400 plus.n69 plus.n68 0.189894
R24401 plus.n69 plus.n57 0.189894
R24402 plus.n74 plus.n57 0.189894
R24403 plus.n75 plus.n74 0.189894
R24404 plus.n75 plus.n55 0.189894
R24405 plus.n79 plus.n55 0.189894
R24406 plus.n80 plus.n79 0.189894
R24407 plus.n80 plus.n53 0.189894
R24408 plus.n85 plus.n53 0.189894
R24409 plus.n86 plus.n85 0.189894
R24410 plus.n87 plus.n86 0.189894
R24411 plus.n87 plus.n51 0.189894
R24412 plus.n92 plus.n51 0.189894
R24413 plus.n93 plus.n92 0.189894
R24414 plus.n93 plus.n49 0.189894
R24415 plus.n97 plus.n49 0.189894
R24416 plus.n48 plus.n0 0.189894
R24417 plus.n44 plus.n0 0.189894
R24418 plus.n44 plus.n43 0.189894
R24419 plus.n43 plus.n2 0.189894
R24420 plus.n38 plus.n2 0.189894
R24421 plus.n38 plus.n37 0.189894
R24422 plus.n37 plus.n36 0.189894
R24423 plus.n36 plus.n4 0.189894
R24424 plus.n31 plus.n4 0.189894
R24425 plus.n31 plus.n30 0.189894
R24426 plus.n30 plus.n6 0.189894
R24427 plus.n26 plus.n6 0.189894
R24428 plus.n26 plus.n25 0.189894
R24429 plus.n25 plus.n8 0.189894
R24430 plus.n20 plus.n8 0.189894
R24431 plus.n20 plus.n19 0.189894
R24432 plus.n19 plus.n18 0.189894
R24433 plus.n18 plus.n10 0.189894
R24434 plus.n13 plus.n10 0.189894
R24435 a_n3827_n3924.n12 a_n3827_n3924.t38 214.994
R24436 a_n3827_n3924.n1 a_n3827_n3924.t45 214.766
R24437 a_n3827_n3924.n13 a_n3827_n3924.t31 214.321
R24438 a_n3827_n3924.n14 a_n3827_n3924.t37 214.321
R24439 a_n3827_n3924.n15 a_n3827_n3924.t35 214.321
R24440 a_n3827_n3924.n16 a_n3827_n3924.t0 214.321
R24441 a_n3827_n3924.n17 a_n3827_n3924.t29 214.321
R24442 a_n3827_n3924.n18 a_n3827_n3924.t3 214.321
R24443 a_n3827_n3924.n19 a_n3827_n3924.t28 214.321
R24444 a_n3827_n3924.n12 a_n3827_n3924.t39 214.321
R24445 a_n3827_n3924.n0 a_n3827_n3924.t19 55.8337
R24446 a_n3827_n3924.n2 a_n3827_n3924.t26 55.8337
R24447 a_n3827_n3924.n11 a_n3827_n3924.t30 55.8337
R24448 a_n3827_n3924.n43 a_n3827_n3924.t7 55.8335
R24449 a_n3827_n3924.n41 a_n3827_n3924.t47 55.8335
R24450 a_n3827_n3924.n32 a_n3827_n3924.t42 55.8335
R24451 a_n3827_n3924.n31 a_n3827_n3924.t16 55.8335
R24452 a_n3827_n3924.n22 a_n3827_n3924.t24 55.8335
R24453 a_n3827_n3924.n45 a_n3827_n3924.n44 53.0052
R24454 a_n3827_n3924.n47 a_n3827_n3924.n46 53.0052
R24455 a_n3827_n3924.n49 a_n3827_n3924.n48 53.0052
R24456 a_n3827_n3924.n4 a_n3827_n3924.n3 53.0052
R24457 a_n3827_n3924.n6 a_n3827_n3924.n5 53.0052
R24458 a_n3827_n3924.n8 a_n3827_n3924.n7 53.0052
R24459 a_n3827_n3924.n10 a_n3827_n3924.n9 53.0052
R24460 a_n3827_n3924.n40 a_n3827_n3924.n39 53.0051
R24461 a_n3827_n3924.n38 a_n3827_n3924.n37 53.0051
R24462 a_n3827_n3924.n36 a_n3827_n3924.n35 53.0051
R24463 a_n3827_n3924.n34 a_n3827_n3924.n33 53.0051
R24464 a_n3827_n3924.n30 a_n3827_n3924.n29 53.0051
R24465 a_n3827_n3924.n28 a_n3827_n3924.n27 53.0051
R24466 a_n3827_n3924.n26 a_n3827_n3924.n25 53.0051
R24467 a_n3827_n3924.n24 a_n3827_n3924.n23 53.0051
R24468 a_n3827_n3924.n51 a_n3827_n3924.n50 53.0051
R24469 a_n3827_n3924.n21 a_n3827_n3924.n11 12.2417
R24470 a_n3827_n3924.n43 a_n3827_n3924.n42 12.2417
R24471 a_n3827_n3924.n22 a_n3827_n3924.n21 5.16214
R24472 a_n3827_n3924.n42 a_n3827_n3924.n41 5.16214
R24473 a_n3827_n3924.n44 a_n3827_n3924.t15 2.82907
R24474 a_n3827_n3924.n44 a_n3827_n3924.t20 2.82907
R24475 a_n3827_n3924.n46 a_n3827_n3924.t13 2.82907
R24476 a_n3827_n3924.n46 a_n3827_n3924.t17 2.82907
R24477 a_n3827_n3924.n48 a_n3827_n3924.t10 2.82907
R24478 a_n3827_n3924.n48 a_n3827_n3924.t14 2.82907
R24479 a_n3827_n3924.n3 a_n3827_n3924.t27 2.82907
R24480 a_n3827_n3924.n3 a_n3827_n3924.t41 2.82907
R24481 a_n3827_n3924.n5 a_n3827_n3924.t36 2.82907
R24482 a_n3827_n3924.n5 a_n3827_n3924.t32 2.82907
R24483 a_n3827_n3924.n7 a_n3827_n3924.t34 2.82907
R24484 a_n3827_n3924.n7 a_n3827_n3924.t33 2.82907
R24485 a_n3827_n3924.n9 a_n3827_n3924.t1 2.82907
R24486 a_n3827_n3924.n9 a_n3827_n3924.t48 2.82907
R24487 a_n3827_n3924.n39 a_n3827_n3924.t40 2.82907
R24488 a_n3827_n3924.n39 a_n3827_n3924.t43 2.82907
R24489 a_n3827_n3924.n37 a_n3827_n3924.t5 2.82907
R24490 a_n3827_n3924.n37 a_n3827_n3924.t46 2.82907
R24491 a_n3827_n3924.n35 a_n3827_n3924.t4 2.82907
R24492 a_n3827_n3924.n35 a_n3827_n3924.t2 2.82907
R24493 a_n3827_n3924.n33 a_n3827_n3924.t49 2.82907
R24494 a_n3827_n3924.n33 a_n3827_n3924.t44 2.82907
R24495 a_n3827_n3924.n29 a_n3827_n3924.t8 2.82907
R24496 a_n3827_n3924.n29 a_n3827_n3924.t21 2.82907
R24497 a_n3827_n3924.n27 a_n3827_n3924.t12 2.82907
R24498 a_n3827_n3924.n27 a_n3827_n3924.t6 2.82907
R24499 a_n3827_n3924.n25 a_n3827_n3924.t23 2.82907
R24500 a_n3827_n3924.n25 a_n3827_n3924.t11 2.82907
R24501 a_n3827_n3924.n23 a_n3827_n3924.t18 2.82907
R24502 a_n3827_n3924.n23 a_n3827_n3924.t22 2.82907
R24503 a_n3827_n3924.t25 a_n3827_n3924.n51 2.82907
R24504 a_n3827_n3924.n51 a_n3827_n3924.t9 2.82907
R24505 a_n3827_n3924.n42 a_n3827_n3924.n1 1.95694
R24506 a_n3827_n3924.n21 a_n3827_n3924.n20 1.95694
R24507 a_n3827_n3924.n19 a_n3827_n3924.n18 0.672012
R24508 a_n3827_n3924.n18 a_n3827_n3924.n17 0.672012
R24509 a_n3827_n3924.n17 a_n3827_n3924.n16 0.672012
R24510 a_n3827_n3924.n16 a_n3827_n3924.n15 0.672012
R24511 a_n3827_n3924.n15 a_n3827_n3924.n14 0.672012
R24512 a_n3827_n3924.n14 a_n3827_n3924.n13 0.672012
R24513 a_n3827_n3924.n24 a_n3827_n3924.n22 0.530672
R24514 a_n3827_n3924.n26 a_n3827_n3924.n24 0.530672
R24515 a_n3827_n3924.n28 a_n3827_n3924.n26 0.530672
R24516 a_n3827_n3924.n30 a_n3827_n3924.n28 0.530672
R24517 a_n3827_n3924.n31 a_n3827_n3924.n30 0.530672
R24518 a_n3827_n3924.n34 a_n3827_n3924.n32 0.530672
R24519 a_n3827_n3924.n36 a_n3827_n3924.n34 0.530672
R24520 a_n3827_n3924.n38 a_n3827_n3924.n36 0.530672
R24521 a_n3827_n3924.n40 a_n3827_n3924.n38 0.530672
R24522 a_n3827_n3924.n41 a_n3827_n3924.n40 0.530672
R24523 a_n3827_n3924.n11 a_n3827_n3924.n10 0.530672
R24524 a_n3827_n3924.n10 a_n3827_n3924.n8 0.530672
R24525 a_n3827_n3924.n8 a_n3827_n3924.n6 0.530672
R24526 a_n3827_n3924.n6 a_n3827_n3924.n4 0.530672
R24527 a_n3827_n3924.n4 a_n3827_n3924.n2 0.530672
R24528 a_n3827_n3924.n50 a_n3827_n3924.n0 0.530672
R24529 a_n3827_n3924.n50 a_n3827_n3924.n49 0.530672
R24530 a_n3827_n3924.n49 a_n3827_n3924.n47 0.530672
R24531 a_n3827_n3924.n47 a_n3827_n3924.n45 0.530672
R24532 a_n3827_n3924.n45 a_n3827_n3924.n43 0.530672
R24533 a_n3827_n3924.n20 a_n3827_n3924.n19 0.370413
R24534 a_n3827_n3924.n20 a_n3827_n3924.n12 0.302099
R24535 a_n3827_n3924.n32 a_n3827_n3924.n31 0.235414
R24536 a_n3827_n3924.n2 a_n3827_n3924.n0 0.235414
R24537 a_n3827_n3924.n13 a_n3827_n3924.n1 0.227971
R24538 diffpairibias.n0 diffpairibias.t27 436.822
R24539 diffpairibias.n27 diffpairibias.t24 435.479
R24540 diffpairibias.n26 diffpairibias.t21 435.479
R24541 diffpairibias.n25 diffpairibias.t22 435.479
R24542 diffpairibias.n24 diffpairibias.t26 435.479
R24543 diffpairibias.n23 diffpairibias.t20 435.479
R24544 diffpairibias.n0 diffpairibias.t23 435.479
R24545 diffpairibias.n1 diffpairibias.t28 435.479
R24546 diffpairibias.n2 diffpairibias.t25 435.479
R24547 diffpairibias.n3 diffpairibias.t29 435.479
R24548 diffpairibias.n13 diffpairibias.t14 377.536
R24549 diffpairibias.n13 diffpairibias.t0 376.193
R24550 diffpairibias.n14 diffpairibias.t10 376.193
R24551 diffpairibias.n15 diffpairibias.t12 376.193
R24552 diffpairibias.n16 diffpairibias.t6 376.193
R24553 diffpairibias.n17 diffpairibias.t2 376.193
R24554 diffpairibias.n18 diffpairibias.t16 376.193
R24555 diffpairibias.n19 diffpairibias.t4 376.193
R24556 diffpairibias.n20 diffpairibias.t18 376.193
R24557 diffpairibias.n21 diffpairibias.t8 376.193
R24558 diffpairibias.n4 diffpairibias.t15 113.368
R24559 diffpairibias.n4 diffpairibias.t1 112.698
R24560 diffpairibias.n5 diffpairibias.t11 112.698
R24561 diffpairibias.n6 diffpairibias.t13 112.698
R24562 diffpairibias.n7 diffpairibias.t7 112.698
R24563 diffpairibias.n8 diffpairibias.t3 112.698
R24564 diffpairibias.n9 diffpairibias.t17 112.698
R24565 diffpairibias.n10 diffpairibias.t5 112.698
R24566 diffpairibias.n11 diffpairibias.t19 112.698
R24567 diffpairibias.n12 diffpairibias.t9 112.698
R24568 diffpairibias.n22 diffpairibias.n21 4.77242
R24569 diffpairibias.n22 diffpairibias.n12 4.30807
R24570 diffpairibias.n23 diffpairibias.n22 4.13945
R24571 diffpairibias.n21 diffpairibias.n20 1.34352
R24572 diffpairibias.n20 diffpairibias.n19 1.34352
R24573 diffpairibias.n19 diffpairibias.n18 1.34352
R24574 diffpairibias.n18 diffpairibias.n17 1.34352
R24575 diffpairibias.n17 diffpairibias.n16 1.34352
R24576 diffpairibias.n16 diffpairibias.n15 1.34352
R24577 diffpairibias.n15 diffpairibias.n14 1.34352
R24578 diffpairibias.n14 diffpairibias.n13 1.34352
R24579 diffpairibias.n3 diffpairibias.n2 1.34352
R24580 diffpairibias.n2 diffpairibias.n1 1.34352
R24581 diffpairibias.n1 diffpairibias.n0 1.34352
R24582 diffpairibias.n24 diffpairibias.n23 1.34352
R24583 diffpairibias.n25 diffpairibias.n24 1.34352
R24584 diffpairibias.n26 diffpairibias.n25 1.34352
R24585 diffpairibias.n27 diffpairibias.n26 1.34352
R24586 diffpairibias.n28 diffpairibias.n27 0.862419
R24587 diffpairibias diffpairibias.n28 0.684875
R24588 diffpairibias.n12 diffpairibias.n11 0.672012
R24589 diffpairibias.n11 diffpairibias.n10 0.672012
R24590 diffpairibias.n10 diffpairibias.n9 0.672012
R24591 diffpairibias.n9 diffpairibias.n8 0.672012
R24592 diffpairibias.n8 diffpairibias.n7 0.672012
R24593 diffpairibias.n7 diffpairibias.n6 0.672012
R24594 diffpairibias.n6 diffpairibias.n5 0.672012
R24595 diffpairibias.n5 diffpairibias.n4 0.672012
R24596 diffpairibias.n28 diffpairibias.n3 0.190907
R24597 a_n2982_8322.n28 a_n2982_8322.t20 74.6477
R24598 a_n2982_8322.n13 a_n2982_8322.t9 74.6477
R24599 a_n2982_8322.n1 a_n2982_8322.t35 74.6474
R24600 a_n2982_8322.n20 a_n2982_8322.t14 74.2899
R24601 a_n2982_8322.n10 a_n2982_8322.t15 74.2899
R24602 a_n2982_8322.n14 a_n2982_8322.t7 74.2899
R24603 a_n2982_8322.n15 a_n2982_8322.t10 74.2899
R24604 a_n2982_8322.n18 a_n2982_8322.t11 74.2899
R24605 a_n2982_8322.n28 a_n2982_8322.n27 70.6783
R24606 a_n2982_8322.n26 a_n2982_8322.n25 70.6783
R24607 a_n2982_8322.n24 a_n2982_8322.n23 70.6783
R24608 a_n2982_8322.n22 a_n2982_8322.n21 70.6783
R24609 a_n2982_8322.n1 a_n2982_8322.n0 70.6783
R24610 a_n2982_8322.n3 a_n2982_8322.n2 70.6783
R24611 a_n2982_8322.n5 a_n2982_8322.n4 70.6783
R24612 a_n2982_8322.n7 a_n2982_8322.n6 70.6783
R24613 a_n2982_8322.n9 a_n2982_8322.n8 70.6783
R24614 a_n2982_8322.n13 a_n2982_8322.n12 70.6783
R24615 a_n2982_8322.n17 a_n2982_8322.n16 70.6783
R24616 a_n2982_8322.n30 a_n2982_8322.n29 70.6782
R24617 a_n2982_8322.n20 a_n2982_8322.n19 24.9022
R24618 a_n2982_8322.n11 a_n2982_8322.t0 9.96358
R24619 a_n2982_8322.n19 a_n2982_8322.n18 8.38735
R24620 a_n2982_8322.n11 a_n2982_8322.n10 6.90998
R24621 a_n2982_8322.n19 a_n2982_8322.n11 5.3452
R24622 a_n2982_8322.n27 a_n2982_8322.t33 3.61217
R24623 a_n2982_8322.n27 a_n2982_8322.t29 3.61217
R24624 a_n2982_8322.n25 a_n2982_8322.t17 3.61217
R24625 a_n2982_8322.n25 a_n2982_8322.t16 3.61217
R24626 a_n2982_8322.n23 a_n2982_8322.t30 3.61217
R24627 a_n2982_8322.n23 a_n2982_8322.t23 3.61217
R24628 a_n2982_8322.n21 a_n2982_8322.t27 3.61217
R24629 a_n2982_8322.n21 a_n2982_8322.t25 3.61217
R24630 a_n2982_8322.n0 a_n2982_8322.t28 3.61217
R24631 a_n2982_8322.n0 a_n2982_8322.t24 3.61217
R24632 a_n2982_8322.n2 a_n2982_8322.t21 3.61217
R24633 a_n2982_8322.n2 a_n2982_8322.t37 3.61217
R24634 a_n2982_8322.n4 a_n2982_8322.t34 3.61217
R24635 a_n2982_8322.n4 a_n2982_8322.t22 3.61217
R24636 a_n2982_8322.n6 a_n2982_8322.t19 3.61217
R24637 a_n2982_8322.n6 a_n2982_8322.t18 3.61217
R24638 a_n2982_8322.n8 a_n2982_8322.t32 3.61217
R24639 a_n2982_8322.n8 a_n2982_8322.t31 3.61217
R24640 a_n2982_8322.n12 a_n2982_8322.t13 3.61217
R24641 a_n2982_8322.n12 a_n2982_8322.t12 3.61217
R24642 a_n2982_8322.n16 a_n2982_8322.t8 3.61217
R24643 a_n2982_8322.n16 a_n2982_8322.t6 3.61217
R24644 a_n2982_8322.t36 a_n2982_8322.n30 3.61217
R24645 a_n2982_8322.n30 a_n2982_8322.t26 3.61217
R24646 a_n2982_8322.n10 a_n2982_8322.n9 0.358259
R24647 a_n2982_8322.n9 a_n2982_8322.n7 0.358259
R24648 a_n2982_8322.n7 a_n2982_8322.n5 0.358259
R24649 a_n2982_8322.n5 a_n2982_8322.n3 0.358259
R24650 a_n2982_8322.n3 a_n2982_8322.n1 0.358259
R24651 a_n2982_8322.n18 a_n2982_8322.n17 0.358259
R24652 a_n2982_8322.n17 a_n2982_8322.n15 0.358259
R24653 a_n2982_8322.n14 a_n2982_8322.n13 0.358259
R24654 a_n2982_8322.n22 a_n2982_8322.n20 0.358259
R24655 a_n2982_8322.n24 a_n2982_8322.n22 0.358259
R24656 a_n2982_8322.n26 a_n2982_8322.n24 0.358259
R24657 a_n2982_8322.n29 a_n2982_8322.n26 0.358259
R24658 a_n2982_8322.n29 a_n2982_8322.n28 0.358259
R24659 a_n2982_8322.n15 a_n2982_8322.n14 0.101793
R24660 a_n2982_8322.t5 a_n2982_8322.t2 0.0788333
R24661 a_n2982_8322.t4 a_n2982_8322.t3 0.0788333
R24662 a_n2982_8322.t0 a_n2982_8322.t1 0.0788333
R24663 a_n2982_8322.t4 a_n2982_8322.t5 0.0318333
R24664 a_n2982_8322.t0 a_n2982_8322.t3 0.0318333
R24665 a_n2982_8322.t2 a_n2982_8322.t3 0.0318333
R24666 a_n2982_8322.t1 a_n2982_8322.t4 0.0318333
R24667 minus.n61 minus.t24 251.488
R24668 minus.n12 minus.t16 251.488
R24669 minus.n102 minus.t4 243.255
R24670 minus.n96 minus.t14 231.093
R24671 minus.n47 minus.t9 231.093
R24672 minus.n101 minus.n99 224.169
R24673 minus.n101 minus.n100 223.454
R24674 minus.n50 minus.t21 187.445
R24675 minus.n89 minus.t18 187.445
R24676 minus.n83 minus.t15 187.445
R24677 minus.n54 minus.t7 187.445
R24678 minus.n56 minus.t6 187.445
R24679 minus.n71 minus.t12 187.445
R24680 minus.n65 minus.t11 187.445
R24681 minus.n60 minus.t19 187.445
R24682 minus.n11 minus.t10 187.445
R24683 minus.n16 minus.t8 187.445
R24684 minus.n22 minus.t5 187.445
R24685 minus.n7 minus.t22 187.445
R24686 minus.n5 minus.t23 187.445
R24687 minus.n34 minus.t17 187.445
R24688 minus.n40 minus.t20 187.445
R24689 minus.n1 minus.t13 187.445
R24690 minus.n63 minus.n62 161.3
R24691 minus.n64 minus.n59 161.3
R24692 minus.n67 minus.n66 161.3
R24693 minus.n68 minus.n58 161.3
R24694 minus.n70 minus.n69 161.3
R24695 minus.n72 minus.n57 161.3
R24696 minus.n74 minus.n73 161.3
R24697 minus.n76 minus.n75 161.3
R24698 minus.n77 minus.n55 161.3
R24699 minus.n79 minus.n78 161.3
R24700 minus.n81 minus.n80 161.3
R24701 minus.n82 minus.n53 161.3
R24702 minus.n85 minus.n84 161.3
R24703 minus.n86 minus.n52 161.3
R24704 minus.n88 minus.n87 161.3
R24705 minus.n90 minus.n51 161.3
R24706 minus.n92 minus.n91 161.3
R24707 minus.n94 minus.n93 161.3
R24708 minus.n95 minus.n49 161.3
R24709 minus.n97 minus.n96 161.3
R24710 minus.n48 minus.n47 161.3
R24711 minus.n46 minus.n0 161.3
R24712 minus.n45 minus.n44 161.3
R24713 minus.n43 minus.n42 161.3
R24714 minus.n41 minus.n2 161.3
R24715 minus.n39 minus.n38 161.3
R24716 minus.n37 minus.n3 161.3
R24717 minus.n36 minus.n35 161.3
R24718 minus.n33 minus.n4 161.3
R24719 minus.n32 minus.n31 161.3
R24720 minus.n30 minus.n29 161.3
R24721 minus.n28 minus.n6 161.3
R24722 minus.n27 minus.n26 161.3
R24723 minus.n25 minus.n24 161.3
R24724 minus.n23 minus.n8 161.3
R24725 minus.n21 minus.n20 161.3
R24726 minus.n19 minus.n9 161.3
R24727 minus.n18 minus.n17 161.3
R24728 minus.n15 minus.n10 161.3
R24729 minus.n14 minus.n13 161.3
R24730 minus.n91 minus.n90 56.5617
R24731 minus.n64 minus.n63 56.5617
R24732 minus.n15 minus.n14 56.5617
R24733 minus.n42 minus.n41 56.5617
R24734 minus.n82 minus.n81 56.5617
R24735 minus.n73 minus.n72 56.5617
R24736 minus.n24 minus.n23 56.5617
R24737 minus.n33 minus.n32 56.5617
R24738 minus.n95 minus.n94 48.3272
R24739 minus.n46 minus.n45 48.3272
R24740 minus.n84 minus.n52 44.4521
R24741 minus.n70 minus.n58 44.4521
R24742 minus.n21 minus.n9 44.4521
R24743 minus.n35 minus.n3 44.4521
R24744 minus.n13 minus.n12 43.0014
R24745 minus.n62 minus.n61 43.0014
R24746 minus.n78 minus.n77 40.577
R24747 minus.n77 minus.n76 40.577
R24748 minus.n28 minus.n27 40.577
R24749 minus.n29 minus.n28 40.577
R24750 minus.n61 minus.n60 39.4345
R24751 minus.n12 minus.n11 39.4345
R24752 minus.n88 minus.n52 36.702
R24753 minus.n66 minus.n58 36.702
R24754 minus.n17 minus.n9 36.702
R24755 minus.n39 minus.n3 36.702
R24756 minus.n98 minus.n97 33.563
R24757 minus.n90 minus.n89 20.9036
R24758 minus.n65 minus.n64 20.9036
R24759 minus.n16 minus.n15 20.9036
R24760 minus.n41 minus.n40 20.9036
R24761 minus.n100 minus.t3 19.8005
R24762 minus.n100 minus.t0 19.8005
R24763 minus.n99 minus.t2 19.8005
R24764 minus.n99 minus.t1 19.8005
R24765 minus.n81 minus.n54 18.9362
R24766 minus.n73 minus.n56 18.9362
R24767 minus.n24 minus.n7 18.9362
R24768 minus.n32 minus.n5 18.9362
R24769 minus.n83 minus.n82 16.9689
R24770 minus.n72 minus.n71 16.9689
R24771 minus.n23 minus.n22 16.9689
R24772 minus.n34 minus.n33 16.9689
R24773 minus.n91 minus.n50 15.0015
R24774 minus.n63 minus.n60 15.0015
R24775 minus.n14 minus.n11 15.0015
R24776 minus.n42 minus.n1 15.0015
R24777 minus.n96 minus.n95 12.4157
R24778 minus.n47 minus.n46 12.4157
R24779 minus.n98 minus.n48 12.1577
R24780 minus minus.n103 12.0243
R24781 minus.n94 minus.n50 9.59132
R24782 minus.n45 minus.n1 9.59132
R24783 minus.n84 minus.n83 7.62397
R24784 minus.n71 minus.n70 7.62397
R24785 minus.n22 minus.n21 7.62397
R24786 minus.n35 minus.n34 7.62397
R24787 minus.n78 minus.n54 5.65662
R24788 minus.n76 minus.n56 5.65662
R24789 minus.n27 minus.n7 5.65662
R24790 minus.n29 minus.n5 5.65662
R24791 minus.n103 minus.n102 4.80222
R24792 minus.n89 minus.n88 3.68928
R24793 minus.n66 minus.n65 3.68928
R24794 minus.n17 minus.n16 3.68928
R24795 minus.n40 minus.n39 3.68928
R24796 minus.n103 minus.n98 0.972091
R24797 minus.n102 minus.n101 0.716017
R24798 minus.n97 minus.n49 0.189894
R24799 minus.n93 minus.n49 0.189894
R24800 minus.n93 minus.n92 0.189894
R24801 minus.n92 minus.n51 0.189894
R24802 minus.n87 minus.n51 0.189894
R24803 minus.n87 minus.n86 0.189894
R24804 minus.n86 minus.n85 0.189894
R24805 minus.n85 minus.n53 0.189894
R24806 minus.n80 minus.n53 0.189894
R24807 minus.n80 minus.n79 0.189894
R24808 minus.n79 minus.n55 0.189894
R24809 minus.n75 minus.n55 0.189894
R24810 minus.n75 minus.n74 0.189894
R24811 minus.n74 minus.n57 0.189894
R24812 minus.n69 minus.n57 0.189894
R24813 minus.n69 minus.n68 0.189894
R24814 minus.n68 minus.n67 0.189894
R24815 minus.n67 minus.n59 0.189894
R24816 minus.n62 minus.n59 0.189894
R24817 minus.n13 minus.n10 0.189894
R24818 minus.n18 minus.n10 0.189894
R24819 minus.n19 minus.n18 0.189894
R24820 minus.n20 minus.n19 0.189894
R24821 minus.n20 minus.n8 0.189894
R24822 minus.n25 minus.n8 0.189894
R24823 minus.n26 minus.n25 0.189894
R24824 minus.n26 minus.n6 0.189894
R24825 minus.n30 minus.n6 0.189894
R24826 minus.n31 minus.n30 0.189894
R24827 minus.n31 minus.n4 0.189894
R24828 minus.n36 minus.n4 0.189894
R24829 minus.n37 minus.n36 0.189894
R24830 minus.n38 minus.n37 0.189894
R24831 minus.n38 minus.n2 0.189894
R24832 minus.n43 minus.n2 0.189894
R24833 minus.n44 minus.n43 0.189894
R24834 minus.n44 minus.n0 0.189894
R24835 minus.n48 minus.n0 0.189894
R24836 outputibias.n27 outputibias.n1 289.615
R24837 outputibias.n58 outputibias.n32 289.615
R24838 outputibias.n90 outputibias.n64 289.615
R24839 outputibias.n122 outputibias.n96 289.615
R24840 outputibias.n28 outputibias.n27 185
R24841 outputibias.n26 outputibias.n25 185
R24842 outputibias.n5 outputibias.n4 185
R24843 outputibias.n20 outputibias.n19 185
R24844 outputibias.n18 outputibias.n17 185
R24845 outputibias.n9 outputibias.n8 185
R24846 outputibias.n12 outputibias.n11 185
R24847 outputibias.n59 outputibias.n58 185
R24848 outputibias.n57 outputibias.n56 185
R24849 outputibias.n36 outputibias.n35 185
R24850 outputibias.n51 outputibias.n50 185
R24851 outputibias.n49 outputibias.n48 185
R24852 outputibias.n40 outputibias.n39 185
R24853 outputibias.n43 outputibias.n42 185
R24854 outputibias.n91 outputibias.n90 185
R24855 outputibias.n89 outputibias.n88 185
R24856 outputibias.n68 outputibias.n67 185
R24857 outputibias.n83 outputibias.n82 185
R24858 outputibias.n81 outputibias.n80 185
R24859 outputibias.n72 outputibias.n71 185
R24860 outputibias.n75 outputibias.n74 185
R24861 outputibias.n123 outputibias.n122 185
R24862 outputibias.n121 outputibias.n120 185
R24863 outputibias.n100 outputibias.n99 185
R24864 outputibias.n115 outputibias.n114 185
R24865 outputibias.n113 outputibias.n112 185
R24866 outputibias.n104 outputibias.n103 185
R24867 outputibias.n107 outputibias.n106 185
R24868 outputibias.n0 outputibias.t11 178.945
R24869 outputibias.n133 outputibias.t8 177.018
R24870 outputibias.n132 outputibias.t10 177.018
R24871 outputibias.n0 outputibias.t9 177.018
R24872 outputibias.t5 outputibias.n10 147.661
R24873 outputibias.t7 outputibias.n41 147.661
R24874 outputibias.t3 outputibias.n73 147.661
R24875 outputibias.t1 outputibias.n105 147.661
R24876 outputibias.n128 outputibias.t4 132.363
R24877 outputibias.n128 outputibias.t6 130.436
R24878 outputibias.n129 outputibias.t2 130.436
R24879 outputibias.n130 outputibias.t0 130.436
R24880 outputibias.n27 outputibias.n26 104.615
R24881 outputibias.n26 outputibias.n4 104.615
R24882 outputibias.n19 outputibias.n4 104.615
R24883 outputibias.n19 outputibias.n18 104.615
R24884 outputibias.n18 outputibias.n8 104.615
R24885 outputibias.n11 outputibias.n8 104.615
R24886 outputibias.n58 outputibias.n57 104.615
R24887 outputibias.n57 outputibias.n35 104.615
R24888 outputibias.n50 outputibias.n35 104.615
R24889 outputibias.n50 outputibias.n49 104.615
R24890 outputibias.n49 outputibias.n39 104.615
R24891 outputibias.n42 outputibias.n39 104.615
R24892 outputibias.n90 outputibias.n89 104.615
R24893 outputibias.n89 outputibias.n67 104.615
R24894 outputibias.n82 outputibias.n67 104.615
R24895 outputibias.n82 outputibias.n81 104.615
R24896 outputibias.n81 outputibias.n71 104.615
R24897 outputibias.n74 outputibias.n71 104.615
R24898 outputibias.n122 outputibias.n121 104.615
R24899 outputibias.n121 outputibias.n99 104.615
R24900 outputibias.n114 outputibias.n99 104.615
R24901 outputibias.n114 outputibias.n113 104.615
R24902 outputibias.n113 outputibias.n103 104.615
R24903 outputibias.n106 outputibias.n103 104.615
R24904 outputibias.n63 outputibias.n31 95.6354
R24905 outputibias.n63 outputibias.n62 94.6732
R24906 outputibias.n95 outputibias.n94 94.6732
R24907 outputibias.n127 outputibias.n126 94.6732
R24908 outputibias.n11 outputibias.t5 52.3082
R24909 outputibias.n42 outputibias.t7 52.3082
R24910 outputibias.n74 outputibias.t3 52.3082
R24911 outputibias.n106 outputibias.t1 52.3082
R24912 outputibias.n12 outputibias.n10 15.6674
R24913 outputibias.n43 outputibias.n41 15.6674
R24914 outputibias.n75 outputibias.n73 15.6674
R24915 outputibias.n107 outputibias.n105 15.6674
R24916 outputibias.n13 outputibias.n9 12.8005
R24917 outputibias.n44 outputibias.n40 12.8005
R24918 outputibias.n76 outputibias.n72 12.8005
R24919 outputibias.n108 outputibias.n104 12.8005
R24920 outputibias.n17 outputibias.n16 12.0247
R24921 outputibias.n48 outputibias.n47 12.0247
R24922 outputibias.n80 outputibias.n79 12.0247
R24923 outputibias.n112 outputibias.n111 12.0247
R24924 outputibias.n20 outputibias.n7 11.249
R24925 outputibias.n51 outputibias.n38 11.249
R24926 outputibias.n83 outputibias.n70 11.249
R24927 outputibias.n115 outputibias.n102 11.249
R24928 outputibias.n21 outputibias.n5 10.4732
R24929 outputibias.n52 outputibias.n36 10.4732
R24930 outputibias.n84 outputibias.n68 10.4732
R24931 outputibias.n116 outputibias.n100 10.4732
R24932 outputibias.n25 outputibias.n24 9.69747
R24933 outputibias.n56 outputibias.n55 9.69747
R24934 outputibias.n88 outputibias.n87 9.69747
R24935 outputibias.n120 outputibias.n119 9.69747
R24936 outputibias.n31 outputibias.n30 9.45567
R24937 outputibias.n62 outputibias.n61 9.45567
R24938 outputibias.n94 outputibias.n93 9.45567
R24939 outputibias.n126 outputibias.n125 9.45567
R24940 outputibias.n30 outputibias.n29 9.3005
R24941 outputibias.n3 outputibias.n2 9.3005
R24942 outputibias.n24 outputibias.n23 9.3005
R24943 outputibias.n22 outputibias.n21 9.3005
R24944 outputibias.n7 outputibias.n6 9.3005
R24945 outputibias.n16 outputibias.n15 9.3005
R24946 outputibias.n14 outputibias.n13 9.3005
R24947 outputibias.n61 outputibias.n60 9.3005
R24948 outputibias.n34 outputibias.n33 9.3005
R24949 outputibias.n55 outputibias.n54 9.3005
R24950 outputibias.n53 outputibias.n52 9.3005
R24951 outputibias.n38 outputibias.n37 9.3005
R24952 outputibias.n47 outputibias.n46 9.3005
R24953 outputibias.n45 outputibias.n44 9.3005
R24954 outputibias.n93 outputibias.n92 9.3005
R24955 outputibias.n66 outputibias.n65 9.3005
R24956 outputibias.n87 outputibias.n86 9.3005
R24957 outputibias.n85 outputibias.n84 9.3005
R24958 outputibias.n70 outputibias.n69 9.3005
R24959 outputibias.n79 outputibias.n78 9.3005
R24960 outputibias.n77 outputibias.n76 9.3005
R24961 outputibias.n125 outputibias.n124 9.3005
R24962 outputibias.n98 outputibias.n97 9.3005
R24963 outputibias.n119 outputibias.n118 9.3005
R24964 outputibias.n117 outputibias.n116 9.3005
R24965 outputibias.n102 outputibias.n101 9.3005
R24966 outputibias.n111 outputibias.n110 9.3005
R24967 outputibias.n109 outputibias.n108 9.3005
R24968 outputibias.n28 outputibias.n3 8.92171
R24969 outputibias.n59 outputibias.n34 8.92171
R24970 outputibias.n91 outputibias.n66 8.92171
R24971 outputibias.n123 outputibias.n98 8.92171
R24972 outputibias.n29 outputibias.n1 8.14595
R24973 outputibias.n60 outputibias.n32 8.14595
R24974 outputibias.n92 outputibias.n64 8.14595
R24975 outputibias.n124 outputibias.n96 8.14595
R24976 outputibias.n31 outputibias.n1 5.81868
R24977 outputibias.n62 outputibias.n32 5.81868
R24978 outputibias.n94 outputibias.n64 5.81868
R24979 outputibias.n126 outputibias.n96 5.81868
R24980 outputibias.n131 outputibias.n130 5.20947
R24981 outputibias.n29 outputibias.n28 5.04292
R24982 outputibias.n60 outputibias.n59 5.04292
R24983 outputibias.n92 outputibias.n91 5.04292
R24984 outputibias.n124 outputibias.n123 5.04292
R24985 outputibias.n131 outputibias.n127 4.42209
R24986 outputibias.n14 outputibias.n10 4.38594
R24987 outputibias.n45 outputibias.n41 4.38594
R24988 outputibias.n77 outputibias.n73 4.38594
R24989 outputibias.n109 outputibias.n105 4.38594
R24990 outputibias.n132 outputibias.n131 4.28454
R24991 outputibias.n25 outputibias.n3 4.26717
R24992 outputibias.n56 outputibias.n34 4.26717
R24993 outputibias.n88 outputibias.n66 4.26717
R24994 outputibias.n120 outputibias.n98 4.26717
R24995 outputibias.n24 outputibias.n5 3.49141
R24996 outputibias.n55 outputibias.n36 3.49141
R24997 outputibias.n87 outputibias.n68 3.49141
R24998 outputibias.n119 outputibias.n100 3.49141
R24999 outputibias.n21 outputibias.n20 2.71565
R25000 outputibias.n52 outputibias.n51 2.71565
R25001 outputibias.n84 outputibias.n83 2.71565
R25002 outputibias.n116 outputibias.n115 2.71565
R25003 outputibias.n17 outputibias.n7 1.93989
R25004 outputibias.n48 outputibias.n38 1.93989
R25005 outputibias.n80 outputibias.n70 1.93989
R25006 outputibias.n112 outputibias.n102 1.93989
R25007 outputibias.n130 outputibias.n129 1.9266
R25008 outputibias.n129 outputibias.n128 1.9266
R25009 outputibias.n133 outputibias.n132 1.92658
R25010 outputibias.n134 outputibias.n133 1.29913
R25011 outputibias.n16 outputibias.n9 1.16414
R25012 outputibias.n47 outputibias.n40 1.16414
R25013 outputibias.n79 outputibias.n72 1.16414
R25014 outputibias.n111 outputibias.n104 1.16414
R25015 outputibias.n127 outputibias.n95 0.962709
R25016 outputibias.n95 outputibias.n63 0.962709
R25017 outputibias.n13 outputibias.n12 0.388379
R25018 outputibias.n44 outputibias.n43 0.388379
R25019 outputibias.n76 outputibias.n75 0.388379
R25020 outputibias.n108 outputibias.n107 0.388379
R25021 outputibias.n134 outputibias.n0 0.337251
R25022 outputibias outputibias.n134 0.302375
R25023 outputibias.n30 outputibias.n2 0.155672
R25024 outputibias.n23 outputibias.n2 0.155672
R25025 outputibias.n23 outputibias.n22 0.155672
R25026 outputibias.n22 outputibias.n6 0.155672
R25027 outputibias.n15 outputibias.n6 0.155672
R25028 outputibias.n15 outputibias.n14 0.155672
R25029 outputibias.n61 outputibias.n33 0.155672
R25030 outputibias.n54 outputibias.n33 0.155672
R25031 outputibias.n54 outputibias.n53 0.155672
R25032 outputibias.n53 outputibias.n37 0.155672
R25033 outputibias.n46 outputibias.n37 0.155672
R25034 outputibias.n46 outputibias.n45 0.155672
R25035 outputibias.n93 outputibias.n65 0.155672
R25036 outputibias.n86 outputibias.n65 0.155672
R25037 outputibias.n86 outputibias.n85 0.155672
R25038 outputibias.n85 outputibias.n69 0.155672
R25039 outputibias.n78 outputibias.n69 0.155672
R25040 outputibias.n78 outputibias.n77 0.155672
R25041 outputibias.n125 outputibias.n97 0.155672
R25042 outputibias.n118 outputibias.n97 0.155672
R25043 outputibias.n118 outputibias.n117 0.155672
R25044 outputibias.n117 outputibias.n101 0.155672
R25045 outputibias.n110 outputibias.n101 0.155672
R25046 outputibias.n110 outputibias.n109 0.155672
R25047 output.n41 output.n15 289.615
R25048 output.n72 output.n46 289.615
R25049 output.n104 output.n78 289.615
R25050 output.n136 output.n110 289.615
R25051 output.n77 output.n45 197.26
R25052 output.n77 output.n76 196.298
R25053 output.n109 output.n108 196.298
R25054 output.n141 output.n140 196.298
R25055 output.n42 output.n41 185
R25056 output.n40 output.n39 185
R25057 output.n19 output.n18 185
R25058 output.n34 output.n33 185
R25059 output.n32 output.n31 185
R25060 output.n23 output.n22 185
R25061 output.n26 output.n25 185
R25062 output.n73 output.n72 185
R25063 output.n71 output.n70 185
R25064 output.n50 output.n49 185
R25065 output.n65 output.n64 185
R25066 output.n63 output.n62 185
R25067 output.n54 output.n53 185
R25068 output.n57 output.n56 185
R25069 output.n105 output.n104 185
R25070 output.n103 output.n102 185
R25071 output.n82 output.n81 185
R25072 output.n97 output.n96 185
R25073 output.n95 output.n94 185
R25074 output.n86 output.n85 185
R25075 output.n89 output.n88 185
R25076 output.n137 output.n136 185
R25077 output.n135 output.n134 185
R25078 output.n114 output.n113 185
R25079 output.n129 output.n128 185
R25080 output.n127 output.n126 185
R25081 output.n118 output.n117 185
R25082 output.n121 output.n120 185
R25083 output.t0 output.n24 147.661
R25084 output.t2 output.n55 147.661
R25085 output.t3 output.n87 147.661
R25086 output.t1 output.n119 147.661
R25087 output.n41 output.n40 104.615
R25088 output.n40 output.n18 104.615
R25089 output.n33 output.n18 104.615
R25090 output.n33 output.n32 104.615
R25091 output.n32 output.n22 104.615
R25092 output.n25 output.n22 104.615
R25093 output.n72 output.n71 104.615
R25094 output.n71 output.n49 104.615
R25095 output.n64 output.n49 104.615
R25096 output.n64 output.n63 104.615
R25097 output.n63 output.n53 104.615
R25098 output.n56 output.n53 104.615
R25099 output.n104 output.n103 104.615
R25100 output.n103 output.n81 104.615
R25101 output.n96 output.n81 104.615
R25102 output.n96 output.n95 104.615
R25103 output.n95 output.n85 104.615
R25104 output.n88 output.n85 104.615
R25105 output.n136 output.n135 104.615
R25106 output.n135 output.n113 104.615
R25107 output.n128 output.n113 104.615
R25108 output.n128 output.n127 104.615
R25109 output.n127 output.n117 104.615
R25110 output.n120 output.n117 104.615
R25111 output.n1 output.t5 77.056
R25112 output.n14 output.t7 76.6694
R25113 output.n1 output.n0 72.7095
R25114 output.n3 output.n2 72.7095
R25115 output.n5 output.n4 72.7095
R25116 output.n7 output.n6 72.7095
R25117 output.n9 output.n8 72.7095
R25118 output.n11 output.n10 72.7095
R25119 output.n13 output.n12 72.7095
R25120 output.n25 output.t0 52.3082
R25121 output.n56 output.t2 52.3082
R25122 output.n88 output.t3 52.3082
R25123 output.n120 output.t1 52.3082
R25124 output.n26 output.n24 15.6674
R25125 output.n57 output.n55 15.6674
R25126 output.n89 output.n87 15.6674
R25127 output.n121 output.n119 15.6674
R25128 output.n27 output.n23 12.8005
R25129 output.n58 output.n54 12.8005
R25130 output.n90 output.n86 12.8005
R25131 output.n122 output.n118 12.8005
R25132 output.n31 output.n30 12.0247
R25133 output.n62 output.n61 12.0247
R25134 output.n94 output.n93 12.0247
R25135 output.n126 output.n125 12.0247
R25136 output.n34 output.n21 11.249
R25137 output.n65 output.n52 11.249
R25138 output.n97 output.n84 11.249
R25139 output.n129 output.n116 11.249
R25140 output.n35 output.n19 10.4732
R25141 output.n66 output.n50 10.4732
R25142 output.n98 output.n82 10.4732
R25143 output.n130 output.n114 10.4732
R25144 output.n39 output.n38 9.69747
R25145 output.n70 output.n69 9.69747
R25146 output.n102 output.n101 9.69747
R25147 output.n134 output.n133 9.69747
R25148 output.n45 output.n44 9.45567
R25149 output.n76 output.n75 9.45567
R25150 output.n108 output.n107 9.45567
R25151 output.n140 output.n139 9.45567
R25152 output.n44 output.n43 9.3005
R25153 output.n17 output.n16 9.3005
R25154 output.n38 output.n37 9.3005
R25155 output.n36 output.n35 9.3005
R25156 output.n21 output.n20 9.3005
R25157 output.n30 output.n29 9.3005
R25158 output.n28 output.n27 9.3005
R25159 output.n75 output.n74 9.3005
R25160 output.n48 output.n47 9.3005
R25161 output.n69 output.n68 9.3005
R25162 output.n67 output.n66 9.3005
R25163 output.n52 output.n51 9.3005
R25164 output.n61 output.n60 9.3005
R25165 output.n59 output.n58 9.3005
R25166 output.n107 output.n106 9.3005
R25167 output.n80 output.n79 9.3005
R25168 output.n101 output.n100 9.3005
R25169 output.n99 output.n98 9.3005
R25170 output.n84 output.n83 9.3005
R25171 output.n93 output.n92 9.3005
R25172 output.n91 output.n90 9.3005
R25173 output.n139 output.n138 9.3005
R25174 output.n112 output.n111 9.3005
R25175 output.n133 output.n132 9.3005
R25176 output.n131 output.n130 9.3005
R25177 output.n116 output.n115 9.3005
R25178 output.n125 output.n124 9.3005
R25179 output.n123 output.n122 9.3005
R25180 output.n42 output.n17 8.92171
R25181 output.n73 output.n48 8.92171
R25182 output.n105 output.n80 8.92171
R25183 output.n137 output.n112 8.92171
R25184 output output.n141 8.15037
R25185 output.n43 output.n15 8.14595
R25186 output.n74 output.n46 8.14595
R25187 output.n106 output.n78 8.14595
R25188 output.n138 output.n110 8.14595
R25189 output.n45 output.n15 5.81868
R25190 output.n76 output.n46 5.81868
R25191 output.n108 output.n78 5.81868
R25192 output.n140 output.n110 5.81868
R25193 output.n43 output.n42 5.04292
R25194 output.n74 output.n73 5.04292
R25195 output.n106 output.n105 5.04292
R25196 output.n138 output.n137 5.04292
R25197 output.n28 output.n24 4.38594
R25198 output.n59 output.n55 4.38594
R25199 output.n91 output.n87 4.38594
R25200 output.n123 output.n119 4.38594
R25201 output.n39 output.n17 4.26717
R25202 output.n70 output.n48 4.26717
R25203 output.n102 output.n80 4.26717
R25204 output.n134 output.n112 4.26717
R25205 output.n0 output.t11 3.9605
R25206 output.n0 output.t16 3.9605
R25207 output.n2 output.t4 3.9605
R25208 output.n2 output.t12 3.9605
R25209 output.n4 output.t14 3.9605
R25210 output.n4 output.t13 3.9605
R25211 output.n6 output.t19 3.9605
R25212 output.n6 output.t6 3.9605
R25213 output.n8 output.t8 3.9605
R25214 output.n8 output.t17 3.9605
R25215 output.n10 output.t18 3.9605
R25216 output.n10 output.t9 3.9605
R25217 output.n12 output.t10 3.9605
R25218 output.n12 output.t15 3.9605
R25219 output.n38 output.n19 3.49141
R25220 output.n69 output.n50 3.49141
R25221 output.n101 output.n82 3.49141
R25222 output.n133 output.n114 3.49141
R25223 output.n35 output.n34 2.71565
R25224 output.n66 output.n65 2.71565
R25225 output.n98 output.n97 2.71565
R25226 output.n130 output.n129 2.71565
R25227 output.n31 output.n21 1.93989
R25228 output.n62 output.n52 1.93989
R25229 output.n94 output.n84 1.93989
R25230 output.n126 output.n116 1.93989
R25231 output.n30 output.n23 1.16414
R25232 output.n61 output.n54 1.16414
R25233 output.n93 output.n86 1.16414
R25234 output.n125 output.n118 1.16414
R25235 output.n141 output.n109 0.962709
R25236 output.n109 output.n77 0.962709
R25237 output.n27 output.n26 0.388379
R25238 output.n58 output.n57 0.388379
R25239 output.n90 output.n89 0.388379
R25240 output.n122 output.n121 0.388379
R25241 output.n14 output.n13 0.387128
R25242 output.n13 output.n11 0.387128
R25243 output.n11 output.n9 0.387128
R25244 output.n9 output.n7 0.387128
R25245 output.n7 output.n5 0.387128
R25246 output.n5 output.n3 0.387128
R25247 output.n3 output.n1 0.387128
R25248 output.n44 output.n16 0.155672
R25249 output.n37 output.n16 0.155672
R25250 output.n37 output.n36 0.155672
R25251 output.n36 output.n20 0.155672
R25252 output.n29 output.n20 0.155672
R25253 output.n29 output.n28 0.155672
R25254 output.n75 output.n47 0.155672
R25255 output.n68 output.n47 0.155672
R25256 output.n68 output.n67 0.155672
R25257 output.n67 output.n51 0.155672
R25258 output.n60 output.n51 0.155672
R25259 output.n60 output.n59 0.155672
R25260 output.n107 output.n79 0.155672
R25261 output.n100 output.n79 0.155672
R25262 output.n100 output.n99 0.155672
R25263 output.n99 output.n83 0.155672
R25264 output.n92 output.n83 0.155672
R25265 output.n92 output.n91 0.155672
R25266 output.n139 output.n111 0.155672
R25267 output.n132 output.n111 0.155672
R25268 output.n132 output.n131 0.155672
R25269 output.n131 output.n115 0.155672
R25270 output.n124 output.n115 0.155672
R25271 output.n124 output.n123 0.155672
R25272 output output.n14 0.126227
C0 output outputibias 2.34152f
C1 vdd output 7.23429f
C2 CSoutput output 6.13881f
C3 CSoutput outputibias 0.032386f
C4 vdd CSoutput 92.9043f
C5 minus diffpairibias 5.12e-19
C6 commonsourceibias output 0.006808f
C7 vdd plus 0.087969f
C8 CSoutput minus 3.16311f
C9 plus diffpairibias 4.13e-19
C10 commonsourceibias outputibias 0.003832f
C11 vdd commonsourceibias 0.004218f
C12 CSoutput plus 0.913039f
C13 commonsourceibias diffpairibias 0.064336f
C14 minus plus 10.3236f
C15 CSoutput commonsourceibias 66.8263f
C16 minus commonsourceibias 0.337885f
C17 plus commonsourceibias 0.284038f
C18 diffpairibias gnd 60.00283f
C19 outputibias gnd 32.465668f
C20 output gnd 15.47879f
C21 commonsourceibias gnd 0.223204p
C22 plus gnd 37.3376f
C23 minus gnd 30.87907f
C24 CSoutput gnd 0.14452p
C25 vdd gnd 0.480516p
C26 output.t5 gnd 0.464308f
C27 output.t11 gnd 0.044422f
C28 output.t16 gnd 0.044422f
C29 output.n0 gnd 0.364624f
C30 output.n1 gnd 0.614102f
C31 output.t4 gnd 0.044422f
C32 output.t12 gnd 0.044422f
C33 output.n2 gnd 0.364624f
C34 output.n3 gnd 0.350265f
C35 output.t14 gnd 0.044422f
C36 output.t13 gnd 0.044422f
C37 output.n4 gnd 0.364624f
C38 output.n5 gnd 0.350265f
C39 output.t19 gnd 0.044422f
C40 output.t6 gnd 0.044422f
C41 output.n6 gnd 0.364624f
C42 output.n7 gnd 0.350265f
C43 output.t8 gnd 0.044422f
C44 output.t17 gnd 0.044422f
C45 output.n8 gnd 0.364624f
C46 output.n9 gnd 0.350265f
C47 output.t18 gnd 0.044422f
C48 output.t9 gnd 0.044422f
C49 output.n10 gnd 0.364624f
C50 output.n11 gnd 0.350265f
C51 output.t10 gnd 0.044422f
C52 output.t15 gnd 0.044422f
C53 output.n12 gnd 0.364624f
C54 output.n13 gnd 0.350265f
C55 output.t7 gnd 0.462979f
C56 output.n14 gnd 0.28994f
C57 output.n15 gnd 0.015803f
C58 output.n16 gnd 0.011243f
C59 output.n17 gnd 0.006041f
C60 output.n18 gnd 0.01428f
C61 output.n19 gnd 0.006397f
C62 output.n20 gnd 0.011243f
C63 output.n21 gnd 0.006041f
C64 output.n22 gnd 0.01428f
C65 output.n23 gnd 0.006397f
C66 output.n24 gnd 0.048111f
C67 output.t0 gnd 0.023274f
C68 output.n25 gnd 0.01071f
C69 output.n26 gnd 0.008435f
C70 output.n27 gnd 0.006041f
C71 output.n28 gnd 0.267512f
C72 output.n29 gnd 0.011243f
C73 output.n30 gnd 0.006041f
C74 output.n31 gnd 0.006397f
C75 output.n32 gnd 0.01428f
C76 output.n33 gnd 0.01428f
C77 output.n34 gnd 0.006397f
C78 output.n35 gnd 0.006041f
C79 output.n36 gnd 0.011243f
C80 output.n37 gnd 0.011243f
C81 output.n38 gnd 0.006041f
C82 output.n39 gnd 0.006397f
C83 output.n40 gnd 0.01428f
C84 output.n41 gnd 0.030913f
C85 output.n42 gnd 0.006397f
C86 output.n43 gnd 0.006041f
C87 output.n44 gnd 0.025987f
C88 output.n45 gnd 0.097665f
C89 output.n46 gnd 0.015803f
C90 output.n47 gnd 0.011243f
C91 output.n48 gnd 0.006041f
C92 output.n49 gnd 0.01428f
C93 output.n50 gnd 0.006397f
C94 output.n51 gnd 0.011243f
C95 output.n52 gnd 0.006041f
C96 output.n53 gnd 0.01428f
C97 output.n54 gnd 0.006397f
C98 output.n55 gnd 0.048111f
C99 output.t2 gnd 0.023274f
C100 output.n56 gnd 0.01071f
C101 output.n57 gnd 0.008435f
C102 output.n58 gnd 0.006041f
C103 output.n59 gnd 0.267512f
C104 output.n60 gnd 0.011243f
C105 output.n61 gnd 0.006041f
C106 output.n62 gnd 0.006397f
C107 output.n63 gnd 0.01428f
C108 output.n64 gnd 0.01428f
C109 output.n65 gnd 0.006397f
C110 output.n66 gnd 0.006041f
C111 output.n67 gnd 0.011243f
C112 output.n68 gnd 0.011243f
C113 output.n69 gnd 0.006041f
C114 output.n70 gnd 0.006397f
C115 output.n71 gnd 0.01428f
C116 output.n72 gnd 0.030913f
C117 output.n73 gnd 0.006397f
C118 output.n74 gnd 0.006041f
C119 output.n75 gnd 0.025987f
C120 output.n76 gnd 0.09306f
C121 output.n77 gnd 1.65264f
C122 output.n78 gnd 0.015803f
C123 output.n79 gnd 0.011243f
C124 output.n80 gnd 0.006041f
C125 output.n81 gnd 0.01428f
C126 output.n82 gnd 0.006397f
C127 output.n83 gnd 0.011243f
C128 output.n84 gnd 0.006041f
C129 output.n85 gnd 0.01428f
C130 output.n86 gnd 0.006397f
C131 output.n87 gnd 0.048111f
C132 output.t3 gnd 0.023274f
C133 output.n88 gnd 0.01071f
C134 output.n89 gnd 0.008435f
C135 output.n90 gnd 0.006041f
C136 output.n91 gnd 0.267512f
C137 output.n92 gnd 0.011243f
C138 output.n93 gnd 0.006041f
C139 output.n94 gnd 0.006397f
C140 output.n95 gnd 0.01428f
C141 output.n96 gnd 0.01428f
C142 output.n97 gnd 0.006397f
C143 output.n98 gnd 0.006041f
C144 output.n99 gnd 0.011243f
C145 output.n100 gnd 0.011243f
C146 output.n101 gnd 0.006041f
C147 output.n102 gnd 0.006397f
C148 output.n103 gnd 0.01428f
C149 output.n104 gnd 0.030913f
C150 output.n105 gnd 0.006397f
C151 output.n106 gnd 0.006041f
C152 output.n107 gnd 0.025987f
C153 output.n108 gnd 0.09306f
C154 output.n109 gnd 0.713089f
C155 output.n110 gnd 0.015803f
C156 output.n111 gnd 0.011243f
C157 output.n112 gnd 0.006041f
C158 output.n113 gnd 0.01428f
C159 output.n114 gnd 0.006397f
C160 output.n115 gnd 0.011243f
C161 output.n116 gnd 0.006041f
C162 output.n117 gnd 0.01428f
C163 output.n118 gnd 0.006397f
C164 output.n119 gnd 0.048111f
C165 output.t1 gnd 0.023274f
C166 output.n120 gnd 0.01071f
C167 output.n121 gnd 0.008435f
C168 output.n122 gnd 0.006041f
C169 output.n123 gnd 0.267512f
C170 output.n124 gnd 0.011243f
C171 output.n125 gnd 0.006041f
C172 output.n126 gnd 0.006397f
C173 output.n127 gnd 0.01428f
C174 output.n128 gnd 0.01428f
C175 output.n129 gnd 0.006397f
C176 output.n130 gnd 0.006041f
C177 output.n131 gnd 0.011243f
C178 output.n132 gnd 0.011243f
C179 output.n133 gnd 0.006041f
C180 output.n134 gnd 0.006397f
C181 output.n135 gnd 0.01428f
C182 output.n136 gnd 0.030913f
C183 output.n137 gnd 0.006397f
C184 output.n138 gnd 0.006041f
C185 output.n139 gnd 0.025987f
C186 output.n140 gnd 0.09306f
C187 output.n141 gnd 1.67353f
C188 outputibias.t9 gnd 0.11477f
C189 outputibias.t11 gnd 0.115567f
C190 outputibias.n0 gnd 0.130108f
C191 outputibias.n1 gnd 0.001372f
C192 outputibias.n2 gnd 9.76e-19
C193 outputibias.n3 gnd 5.24e-19
C194 outputibias.n4 gnd 0.001239f
C195 outputibias.n5 gnd 5.55e-19
C196 outputibias.n6 gnd 9.76e-19
C197 outputibias.n7 gnd 5.24e-19
C198 outputibias.n8 gnd 0.001239f
C199 outputibias.n9 gnd 5.55e-19
C200 outputibias.n10 gnd 0.004176f
C201 outputibias.t5 gnd 0.00202f
C202 outputibias.n11 gnd 9.3e-19
C203 outputibias.n12 gnd 7.32e-19
C204 outputibias.n13 gnd 5.24e-19
C205 outputibias.n14 gnd 0.02322f
C206 outputibias.n15 gnd 9.76e-19
C207 outputibias.n16 gnd 5.24e-19
C208 outputibias.n17 gnd 5.55e-19
C209 outputibias.n18 gnd 0.001239f
C210 outputibias.n19 gnd 0.001239f
C211 outputibias.n20 gnd 5.55e-19
C212 outputibias.n21 gnd 5.24e-19
C213 outputibias.n22 gnd 9.76e-19
C214 outputibias.n23 gnd 9.76e-19
C215 outputibias.n24 gnd 5.24e-19
C216 outputibias.n25 gnd 5.55e-19
C217 outputibias.n26 gnd 0.001239f
C218 outputibias.n27 gnd 0.002683f
C219 outputibias.n28 gnd 5.55e-19
C220 outputibias.n29 gnd 5.24e-19
C221 outputibias.n30 gnd 0.002256f
C222 outputibias.n31 gnd 0.005781f
C223 outputibias.n32 gnd 0.001372f
C224 outputibias.n33 gnd 9.76e-19
C225 outputibias.n34 gnd 5.24e-19
C226 outputibias.n35 gnd 0.001239f
C227 outputibias.n36 gnd 5.55e-19
C228 outputibias.n37 gnd 9.76e-19
C229 outputibias.n38 gnd 5.24e-19
C230 outputibias.n39 gnd 0.001239f
C231 outputibias.n40 gnd 5.55e-19
C232 outputibias.n41 gnd 0.004176f
C233 outputibias.t7 gnd 0.00202f
C234 outputibias.n42 gnd 9.3e-19
C235 outputibias.n43 gnd 7.32e-19
C236 outputibias.n44 gnd 5.24e-19
C237 outputibias.n45 gnd 0.02322f
C238 outputibias.n46 gnd 9.76e-19
C239 outputibias.n47 gnd 5.24e-19
C240 outputibias.n48 gnd 5.55e-19
C241 outputibias.n49 gnd 0.001239f
C242 outputibias.n50 gnd 0.001239f
C243 outputibias.n51 gnd 5.55e-19
C244 outputibias.n52 gnd 5.24e-19
C245 outputibias.n53 gnd 9.76e-19
C246 outputibias.n54 gnd 9.76e-19
C247 outputibias.n55 gnd 5.24e-19
C248 outputibias.n56 gnd 5.55e-19
C249 outputibias.n57 gnd 0.001239f
C250 outputibias.n58 gnd 0.002683f
C251 outputibias.n59 gnd 5.55e-19
C252 outputibias.n60 gnd 5.24e-19
C253 outputibias.n61 gnd 0.002256f
C254 outputibias.n62 gnd 0.005197f
C255 outputibias.n63 gnd 0.121892f
C256 outputibias.n64 gnd 0.001372f
C257 outputibias.n65 gnd 9.76e-19
C258 outputibias.n66 gnd 5.24e-19
C259 outputibias.n67 gnd 0.001239f
C260 outputibias.n68 gnd 5.55e-19
C261 outputibias.n69 gnd 9.76e-19
C262 outputibias.n70 gnd 5.24e-19
C263 outputibias.n71 gnd 0.001239f
C264 outputibias.n72 gnd 5.55e-19
C265 outputibias.n73 gnd 0.004176f
C266 outputibias.t3 gnd 0.00202f
C267 outputibias.n74 gnd 9.3e-19
C268 outputibias.n75 gnd 7.32e-19
C269 outputibias.n76 gnd 5.24e-19
C270 outputibias.n77 gnd 0.02322f
C271 outputibias.n78 gnd 9.76e-19
C272 outputibias.n79 gnd 5.24e-19
C273 outputibias.n80 gnd 5.55e-19
C274 outputibias.n81 gnd 0.001239f
C275 outputibias.n82 gnd 0.001239f
C276 outputibias.n83 gnd 5.55e-19
C277 outputibias.n84 gnd 5.24e-19
C278 outputibias.n85 gnd 9.76e-19
C279 outputibias.n86 gnd 9.76e-19
C280 outputibias.n87 gnd 5.24e-19
C281 outputibias.n88 gnd 5.55e-19
C282 outputibias.n89 gnd 0.001239f
C283 outputibias.n90 gnd 0.002683f
C284 outputibias.n91 gnd 5.55e-19
C285 outputibias.n92 gnd 5.24e-19
C286 outputibias.n93 gnd 0.002256f
C287 outputibias.n94 gnd 0.005197f
C288 outputibias.n95 gnd 0.064513f
C289 outputibias.n96 gnd 0.001372f
C290 outputibias.n97 gnd 9.76e-19
C291 outputibias.n98 gnd 5.24e-19
C292 outputibias.n99 gnd 0.001239f
C293 outputibias.n100 gnd 5.55e-19
C294 outputibias.n101 gnd 9.76e-19
C295 outputibias.n102 gnd 5.24e-19
C296 outputibias.n103 gnd 0.001239f
C297 outputibias.n104 gnd 5.55e-19
C298 outputibias.n105 gnd 0.004176f
C299 outputibias.t1 gnd 0.00202f
C300 outputibias.n106 gnd 9.3e-19
C301 outputibias.n107 gnd 7.32e-19
C302 outputibias.n108 gnd 5.24e-19
C303 outputibias.n109 gnd 0.02322f
C304 outputibias.n110 gnd 9.76e-19
C305 outputibias.n111 gnd 5.24e-19
C306 outputibias.n112 gnd 5.55e-19
C307 outputibias.n113 gnd 0.001239f
C308 outputibias.n114 gnd 0.001239f
C309 outputibias.n115 gnd 5.55e-19
C310 outputibias.n116 gnd 5.24e-19
C311 outputibias.n117 gnd 9.76e-19
C312 outputibias.n118 gnd 9.76e-19
C313 outputibias.n119 gnd 5.24e-19
C314 outputibias.n120 gnd 5.55e-19
C315 outputibias.n121 gnd 0.001239f
C316 outputibias.n122 gnd 0.002683f
C317 outputibias.n123 gnd 5.55e-19
C318 outputibias.n124 gnd 5.24e-19
C319 outputibias.n125 gnd 0.002256f
C320 outputibias.n126 gnd 0.005197f
C321 outputibias.n127 gnd 0.084814f
C322 outputibias.t0 gnd 0.108319f
C323 outputibias.t2 gnd 0.108319f
C324 outputibias.t6 gnd 0.108319f
C325 outputibias.t4 gnd 0.109238f
C326 outputibias.n128 gnd 0.134674f
C327 outputibias.n129 gnd 0.07244f
C328 outputibias.n130 gnd 0.079818f
C329 outputibias.n131 gnd 0.164901f
C330 outputibias.t10 gnd 0.11477f
C331 outputibias.n132 gnd 0.067481f
C332 outputibias.t8 gnd 0.11477f
C333 outputibias.n133 gnd 0.065115f
C334 outputibias.n134 gnd 0.029159f
C335 minus.n0 gnd 0.029643f
C336 minus.t13 gnd 0.498449f
C337 minus.n1 gnd 0.201595f
C338 minus.n2 gnd 0.029643f
C339 minus.t20 gnd 0.498449f
C340 minus.n3 gnd 0.024552f
C341 minus.n4 gnd 0.029643f
C342 minus.t17 gnd 0.498449f
C343 minus.t23 gnd 0.498449f
C344 minus.n5 gnd 0.201595f
C345 minus.n6 gnd 0.029643f
C346 minus.t22 gnd 0.498449f
C347 minus.n7 gnd 0.201595f
C348 minus.n8 gnd 0.029643f
C349 minus.t5 gnd 0.498449f
C350 minus.n9 gnd 0.024552f
C351 minus.n10 gnd 0.029643f
C352 minus.t8 gnd 0.498449f
C353 minus.t10 gnd 0.498449f
C354 minus.n11 gnd 0.231826f
C355 minus.t16 gnd 0.55863f
C356 minus.n12 gnd 0.234793f
C357 minus.n13 gnd 0.126525f
C358 minus.n14 gnd 0.037428f
C359 minus.n15 gnd 0.0341f
C360 minus.n16 gnd 0.201595f
C361 minus.n17 gnd 0.036381f
C362 minus.n18 gnd 0.029643f
C363 minus.n19 gnd 0.029643f
C364 minus.n20 gnd 0.029643f
C365 minus.n21 gnd 0.038428f
C366 minus.n22 gnd 0.201595f
C367 minus.n23 gnd 0.036319f
C368 minus.n24 gnd 0.035209f
C369 minus.n25 gnd 0.029643f
C370 minus.n26 gnd 0.029643f
C371 minus.n27 gnd 0.03771f
C372 minus.n28 gnd 0.023942f
C373 minus.n29 gnd 0.03771f
C374 minus.n30 gnd 0.029643f
C375 minus.n31 gnd 0.029643f
C376 minus.n32 gnd 0.035209f
C377 minus.n33 gnd 0.036319f
C378 minus.n34 gnd 0.201595f
C379 minus.n35 gnd 0.038428f
C380 minus.n36 gnd 0.029643f
C381 minus.n37 gnd 0.029643f
C382 minus.n38 gnd 0.029643f
C383 minus.n39 gnd 0.036381f
C384 minus.n40 gnd 0.201595f
C385 minus.n41 gnd 0.0341f
C386 minus.n42 gnd 0.037428f
C387 minus.n43 gnd 0.029643f
C388 minus.n44 gnd 0.029643f
C389 minus.n45 gnd 0.038684f
C390 minus.n46 gnd 0.011481f
C391 minus.t9 gnd 0.539073f
C392 minus.n47 gnd 0.233779f
C393 minus.n48 gnd 0.347788f
C394 minus.n49 gnd 0.029643f
C395 minus.t14 gnd 0.539073f
C396 minus.t21 gnd 0.498449f
C397 minus.n50 gnd 0.201595f
C398 minus.n51 gnd 0.029643f
C399 minus.t18 gnd 0.498449f
C400 minus.n52 gnd 0.024552f
C401 minus.n53 gnd 0.029643f
C402 minus.t15 gnd 0.498449f
C403 minus.t7 gnd 0.498449f
C404 minus.n54 gnd 0.201595f
C405 minus.n55 gnd 0.029643f
C406 minus.t6 gnd 0.498449f
C407 minus.n56 gnd 0.201595f
C408 minus.n57 gnd 0.029643f
C409 minus.t12 gnd 0.498449f
C410 minus.n58 gnd 0.024552f
C411 minus.n59 gnd 0.029643f
C412 minus.t11 gnd 0.498449f
C413 minus.t19 gnd 0.498449f
C414 minus.n60 gnd 0.231826f
C415 minus.t24 gnd 0.55863f
C416 minus.n61 gnd 0.234793f
C417 minus.n62 gnd 0.126525f
C418 minus.n63 gnd 0.037428f
C419 minus.n64 gnd 0.0341f
C420 minus.n65 gnd 0.201595f
C421 minus.n66 gnd 0.036381f
C422 minus.n67 gnd 0.029643f
C423 minus.n68 gnd 0.029643f
C424 minus.n69 gnd 0.029643f
C425 minus.n70 gnd 0.038428f
C426 minus.n71 gnd 0.201595f
C427 minus.n72 gnd 0.036319f
C428 minus.n73 gnd 0.035209f
C429 minus.n74 gnd 0.029643f
C430 minus.n75 gnd 0.029643f
C431 minus.n76 gnd 0.03771f
C432 minus.n77 gnd 0.023942f
C433 minus.n78 gnd 0.03771f
C434 minus.n79 gnd 0.029643f
C435 minus.n80 gnd 0.029643f
C436 minus.n81 gnd 0.035209f
C437 minus.n82 gnd 0.036319f
C438 minus.n83 gnd 0.201595f
C439 minus.n84 gnd 0.038428f
C440 minus.n85 gnd 0.029643f
C441 minus.n86 gnd 0.029643f
C442 minus.n87 gnd 0.029643f
C443 minus.n88 gnd 0.036381f
C444 minus.n89 gnd 0.201595f
C445 minus.n90 gnd 0.0341f
C446 minus.n91 gnd 0.037428f
C447 minus.n92 gnd 0.029643f
C448 minus.n93 gnd 0.029643f
C449 minus.n94 gnd 0.038684f
C450 minus.n95 gnd 0.011481f
C451 minus.n96 gnd 0.233779f
C452 minus.n97 gnd 1.00193f
C453 minus.n98 gnd 1.489f
C454 minus.t2 gnd 0.009138f
C455 minus.t1 gnd 0.009138f
C456 minus.n99 gnd 0.030049f
C457 minus.t3 gnd 0.009138f
C458 minus.t0 gnd 0.009138f
C459 minus.n100 gnd 0.029637f
C460 minus.n101 gnd 0.252936f
C461 minus.t4 gnd 0.050862f
C462 minus.n102 gnd 0.138025f
C463 minus.n103 gnd 2.19148f
C464 a_n2982_8322.t26 gnd 0.100069f
C465 a_n2982_8322.t3 gnd 20.7601f
C466 a_n2982_8322.t2 gnd 20.6146f
C467 a_n2982_8322.t5 gnd 20.6146f
C468 a_n2982_8322.t4 gnd 20.7601f
C469 a_n2982_8322.t1 gnd 20.6146f
C470 a_n2982_8322.t0 gnd 30.2036f
C471 a_n2982_8322.t35 gnd 0.936988f
C472 a_n2982_8322.t28 gnd 0.100069f
C473 a_n2982_8322.t24 gnd 0.100069f
C474 a_n2982_8322.n0 gnd 0.704883f
C475 a_n2982_8322.n1 gnd 0.787605f
C476 a_n2982_8322.t21 gnd 0.100069f
C477 a_n2982_8322.t37 gnd 0.100069f
C478 a_n2982_8322.n2 gnd 0.704883f
C479 a_n2982_8322.n3 gnd 0.400171f
C480 a_n2982_8322.t34 gnd 0.100069f
C481 a_n2982_8322.t22 gnd 0.100069f
C482 a_n2982_8322.n4 gnd 0.704883f
C483 a_n2982_8322.n5 gnd 0.400171f
C484 a_n2982_8322.t19 gnd 0.100069f
C485 a_n2982_8322.t18 gnd 0.100069f
C486 a_n2982_8322.n6 gnd 0.704883f
C487 a_n2982_8322.n7 gnd 0.400171f
C488 a_n2982_8322.t32 gnd 0.100069f
C489 a_n2982_8322.t31 gnd 0.100069f
C490 a_n2982_8322.n8 gnd 0.704883f
C491 a_n2982_8322.n9 gnd 0.400171f
C492 a_n2982_8322.t15 gnd 0.935125f
C493 a_n2982_8322.n10 gnd 1.11045f
C494 a_n2982_8322.n11 gnd 3.82915f
C495 a_n2982_8322.t9 gnd 0.936991f
C496 a_n2982_8322.t13 gnd 0.100069f
C497 a_n2982_8322.t12 gnd 0.100069f
C498 a_n2982_8322.n12 gnd 0.704883f
C499 a_n2982_8322.n13 gnd 0.787602f
C500 a_n2982_8322.t7 gnd 0.935125f
C501 a_n2982_8322.n14 gnd 0.396333f
C502 a_n2982_8322.t10 gnd 0.935125f
C503 a_n2982_8322.n15 gnd 0.396333f
C504 a_n2982_8322.t8 gnd 0.100069f
C505 a_n2982_8322.t6 gnd 0.100069f
C506 a_n2982_8322.n16 gnd 0.704883f
C507 a_n2982_8322.n17 gnd 0.400171f
C508 a_n2982_8322.t11 gnd 0.935125f
C509 a_n2982_8322.n18 gnd 1.47007f
C510 a_n2982_8322.n19 gnd 2.34921f
C511 a_n2982_8322.t14 gnd 0.935125f
C512 a_n2982_8322.n20 gnd 1.86969f
C513 a_n2982_8322.t27 gnd 0.100069f
C514 a_n2982_8322.t25 gnd 0.100069f
C515 a_n2982_8322.n21 gnd 0.704883f
C516 a_n2982_8322.n22 gnd 0.400171f
C517 a_n2982_8322.t30 gnd 0.100069f
C518 a_n2982_8322.t23 gnd 0.100069f
C519 a_n2982_8322.n23 gnd 0.704883f
C520 a_n2982_8322.n24 gnd 0.400171f
C521 a_n2982_8322.t17 gnd 0.100069f
C522 a_n2982_8322.t16 gnd 0.100069f
C523 a_n2982_8322.n25 gnd 0.704883f
C524 a_n2982_8322.n26 gnd 0.400171f
C525 a_n2982_8322.t20 gnd 0.936991f
C526 a_n2982_8322.t33 gnd 0.100069f
C527 a_n2982_8322.t29 gnd 0.100069f
C528 a_n2982_8322.n27 gnd 0.704883f
C529 a_n2982_8322.n28 gnd 0.787602f
C530 a_n2982_8322.n29 gnd 0.400169f
C531 a_n2982_8322.n30 gnd 0.704885f
C532 a_n2982_8322.t36 gnd 0.100069f
C533 diffpairibias.t27 gnd 0.090128f
C534 diffpairibias.t23 gnd 0.08996f
C535 diffpairibias.n0 gnd 0.105991f
C536 diffpairibias.t28 gnd 0.08996f
C537 diffpairibias.n1 gnd 0.051736f
C538 diffpairibias.t25 gnd 0.08996f
C539 diffpairibias.n2 gnd 0.051736f
C540 diffpairibias.t29 gnd 0.08996f
C541 diffpairibias.n3 gnd 0.041084f
C542 diffpairibias.t15 gnd 0.086371f
C543 diffpairibias.t1 gnd 0.085993f
C544 diffpairibias.n4 gnd 0.13579f
C545 diffpairibias.t11 gnd 0.085993f
C546 diffpairibias.n5 gnd 0.072463f
C547 diffpairibias.t13 gnd 0.085993f
C548 diffpairibias.n6 gnd 0.072463f
C549 diffpairibias.t7 gnd 0.085993f
C550 diffpairibias.n7 gnd 0.072463f
C551 diffpairibias.t3 gnd 0.085993f
C552 diffpairibias.n8 gnd 0.072463f
C553 diffpairibias.t17 gnd 0.085993f
C554 diffpairibias.n9 gnd 0.072463f
C555 diffpairibias.t5 gnd 0.085993f
C556 diffpairibias.n10 gnd 0.072463f
C557 diffpairibias.t19 gnd 0.085993f
C558 diffpairibias.n11 gnd 0.072463f
C559 diffpairibias.t9 gnd 0.085993f
C560 diffpairibias.n12 gnd 0.102883f
C561 diffpairibias.t14 gnd 0.086899f
C562 diffpairibias.t0 gnd 0.086748f
C563 diffpairibias.n13 gnd 0.094648f
C564 diffpairibias.t10 gnd 0.086748f
C565 diffpairibias.n14 gnd 0.052262f
C566 diffpairibias.t12 gnd 0.086748f
C567 diffpairibias.n15 gnd 0.052262f
C568 diffpairibias.t6 gnd 0.086748f
C569 diffpairibias.n16 gnd 0.052262f
C570 diffpairibias.t2 gnd 0.086748f
C571 diffpairibias.n17 gnd 0.052262f
C572 diffpairibias.t16 gnd 0.086748f
C573 diffpairibias.n18 gnd 0.052262f
C574 diffpairibias.t4 gnd 0.086748f
C575 diffpairibias.n19 gnd 0.052262f
C576 diffpairibias.t18 gnd 0.086748f
C577 diffpairibias.n20 gnd 0.052262f
C578 diffpairibias.t8 gnd 0.086748f
C579 diffpairibias.n21 gnd 0.061849f
C580 diffpairibias.n22 gnd 0.233513f
C581 diffpairibias.t20 gnd 0.08996f
C582 diffpairibias.n23 gnd 0.051747f
C583 diffpairibias.t26 gnd 0.08996f
C584 diffpairibias.n24 gnd 0.051736f
C585 diffpairibias.t22 gnd 0.08996f
C586 diffpairibias.n25 gnd 0.051736f
C587 diffpairibias.t21 gnd 0.08996f
C588 diffpairibias.n26 gnd 0.051736f
C589 diffpairibias.t24 gnd 0.08996f
C590 diffpairibias.n27 gnd 0.04729f
C591 diffpairibias.n28 gnd 0.047711f
C592 a_n3827_n3924.t9 gnd 0.089565f
C593 a_n3827_n3924.t19 gnd 0.930867f
C594 a_n3827_n3924.n0 gnd 0.351909f
C595 a_n3827_n3924.t45 gnd 1.15846f
C596 a_n3827_n3924.n1 gnd 1.34803f
C597 a_n3827_n3924.t26 gnd 0.930867f
C598 a_n3827_n3924.n2 gnd 0.351909f
C599 a_n3827_n3924.t27 gnd 0.089565f
C600 a_n3827_n3924.t41 gnd 0.089565f
C601 a_n3827_n3924.n3 gnd 0.731494f
C602 a_n3827_n3924.n4 gnd 0.368632f
C603 a_n3827_n3924.t36 gnd 0.089565f
C604 a_n3827_n3924.t32 gnd 0.089565f
C605 a_n3827_n3924.n5 gnd 0.731494f
C606 a_n3827_n3924.n6 gnd 0.368632f
C607 a_n3827_n3924.t34 gnd 0.089565f
C608 a_n3827_n3924.t33 gnd 0.089565f
C609 a_n3827_n3924.n7 gnd 0.731494f
C610 a_n3827_n3924.n8 gnd 0.368632f
C611 a_n3827_n3924.t1 gnd 0.089565f
C612 a_n3827_n3924.t48 gnd 0.089565f
C613 a_n3827_n3924.n9 gnd 0.731494f
C614 a_n3827_n3924.n10 gnd 0.368632f
C615 a_n3827_n3924.t30 gnd 0.930867f
C616 a_n3827_n3924.n11 gnd 0.871363f
C617 a_n3827_n3924.t38 gnd 1.15823f
C618 a_n3827_n3924.t39 gnd 1.15658f
C619 a_n3827_n3924.n12 gnd 1.17173f
C620 a_n3827_n3924.t31 gnd 1.15658f
C621 a_n3827_n3924.n13 gnd 0.610864f
C622 a_n3827_n3924.t37 gnd 1.15658f
C623 a_n3827_n3924.n14 gnd 0.8146f
C624 a_n3827_n3924.t35 gnd 1.15658f
C625 a_n3827_n3924.n15 gnd 0.8146f
C626 a_n3827_n3924.t0 gnd 1.15658f
C627 a_n3827_n3924.n16 gnd 0.8146f
C628 a_n3827_n3924.t29 gnd 1.15658f
C629 a_n3827_n3924.n17 gnd 0.8146f
C630 a_n3827_n3924.t3 gnd 1.15658f
C631 a_n3827_n3924.n18 gnd 0.8146f
C632 a_n3827_n3924.t28 gnd 1.15658f
C633 a_n3827_n3924.n19 gnd 0.676219f
C634 a_n3827_n3924.n20 gnd 0.440277f
C635 a_n3827_n3924.n21 gnd 0.844371f
C636 a_n3827_n3924.t24 gnd 0.930864f
C637 a_n3827_n3924.n22 gnd 0.578206f
C638 a_n3827_n3924.t18 gnd 0.089565f
C639 a_n3827_n3924.t22 gnd 0.089565f
C640 a_n3827_n3924.n23 gnd 0.731493f
C641 a_n3827_n3924.n24 gnd 0.368633f
C642 a_n3827_n3924.t23 gnd 0.089565f
C643 a_n3827_n3924.t11 gnd 0.089565f
C644 a_n3827_n3924.n25 gnd 0.731493f
C645 a_n3827_n3924.n26 gnd 0.368633f
C646 a_n3827_n3924.t12 gnd 0.089565f
C647 a_n3827_n3924.t6 gnd 0.089565f
C648 a_n3827_n3924.n27 gnd 0.731493f
C649 a_n3827_n3924.n28 gnd 0.368633f
C650 a_n3827_n3924.t8 gnd 0.089565f
C651 a_n3827_n3924.t21 gnd 0.089565f
C652 a_n3827_n3924.n29 gnd 0.731493f
C653 a_n3827_n3924.n30 gnd 0.368633f
C654 a_n3827_n3924.t16 gnd 0.930864f
C655 a_n3827_n3924.n31 gnd 0.351913f
C656 a_n3827_n3924.t42 gnd 0.930864f
C657 a_n3827_n3924.n32 gnd 0.351913f
C658 a_n3827_n3924.t49 gnd 0.089565f
C659 a_n3827_n3924.t44 gnd 0.089565f
C660 a_n3827_n3924.n33 gnd 0.731493f
C661 a_n3827_n3924.n34 gnd 0.368633f
C662 a_n3827_n3924.t4 gnd 0.089565f
C663 a_n3827_n3924.t2 gnd 0.089565f
C664 a_n3827_n3924.n35 gnd 0.731493f
C665 a_n3827_n3924.n36 gnd 0.368633f
C666 a_n3827_n3924.t5 gnd 0.089565f
C667 a_n3827_n3924.t46 gnd 0.089565f
C668 a_n3827_n3924.n37 gnd 0.731493f
C669 a_n3827_n3924.n38 gnd 0.368633f
C670 a_n3827_n3924.t40 gnd 0.089565f
C671 a_n3827_n3924.t43 gnd 0.089565f
C672 a_n3827_n3924.n39 gnd 0.731493f
C673 a_n3827_n3924.n40 gnd 0.368633f
C674 a_n3827_n3924.t47 gnd 0.930864f
C675 a_n3827_n3924.n41 gnd 0.578206f
C676 a_n3827_n3924.n42 gnd 0.844371f
C677 a_n3827_n3924.t7 gnd 0.930864f
C678 a_n3827_n3924.n43 gnd 0.871367f
C679 a_n3827_n3924.t15 gnd 0.089565f
C680 a_n3827_n3924.t20 gnd 0.089565f
C681 a_n3827_n3924.n44 gnd 0.731494f
C682 a_n3827_n3924.n45 gnd 0.368632f
C683 a_n3827_n3924.t13 gnd 0.089565f
C684 a_n3827_n3924.t17 gnd 0.089565f
C685 a_n3827_n3924.n46 gnd 0.731494f
C686 a_n3827_n3924.n47 gnd 0.368632f
C687 a_n3827_n3924.t10 gnd 0.089565f
C688 a_n3827_n3924.t14 gnd 0.089565f
C689 a_n3827_n3924.n48 gnd 0.731494f
C690 a_n3827_n3924.n49 gnd 0.368632f
C691 a_n3827_n3924.n50 gnd 0.368631f
C692 a_n3827_n3924.n51 gnd 0.731495f
C693 a_n3827_n3924.t25 gnd 0.089565f
C694 plus.n0 gnd 0.021953f
C695 plus.t6 gnd 0.399228f
C696 plus.t12 gnd 0.369143f
C697 plus.n1 gnd 0.149298f
C698 plus.n2 gnd 0.021953f
C699 plus.t8 gnd 0.369143f
C700 plus.n3 gnd 0.018183f
C701 plus.n4 gnd 0.021953f
C702 plus.t7 gnd 0.369143f
C703 plus.t19 gnd 0.369143f
C704 plus.n5 gnd 0.149298f
C705 plus.n6 gnd 0.021953f
C706 plus.t18 gnd 0.369143f
C707 plus.n7 gnd 0.149298f
C708 plus.n8 gnd 0.021953f
C709 plus.t24 gnd 0.369143f
C710 plus.n9 gnd 0.018183f
C711 plus.n10 gnd 0.021953f
C712 plus.t22 gnd 0.369143f
C713 plus.t9 gnd 0.369143f
C714 plus.n11 gnd 0.171686f
C715 plus.t14 gnd 0.413712f
C716 plus.n12 gnd 0.173884f
C717 plus.n13 gnd 0.093702f
C718 plus.n14 gnd 0.027719f
C719 plus.n15 gnd 0.025254f
C720 plus.n16 gnd 0.149298f
C721 plus.n17 gnd 0.026943f
C722 plus.n18 gnd 0.021953f
C723 plus.n19 gnd 0.021953f
C724 plus.n20 gnd 0.021953f
C725 plus.n21 gnd 0.028459f
C726 plus.n22 gnd 0.149298f
C727 plus.n23 gnd 0.026897f
C728 plus.n24 gnd 0.026075f
C729 plus.n25 gnd 0.021953f
C730 plus.n26 gnd 0.021953f
C731 plus.n27 gnd 0.027927f
C732 plus.n28 gnd 0.017731f
C733 plus.n29 gnd 0.027927f
C734 plus.n30 gnd 0.021953f
C735 plus.n31 gnd 0.021953f
C736 plus.n32 gnd 0.026075f
C737 plus.n33 gnd 0.026897f
C738 plus.n34 gnd 0.149298f
C739 plus.n35 gnd 0.028459f
C740 plus.n36 gnd 0.021953f
C741 plus.n37 gnd 0.021953f
C742 plus.n38 gnd 0.021953f
C743 plus.n39 gnd 0.026943f
C744 plus.n40 gnd 0.149298f
C745 plus.n41 gnd 0.025254f
C746 plus.n42 gnd 0.027719f
C747 plus.n43 gnd 0.021953f
C748 plus.n44 gnd 0.021953f
C749 plus.n45 gnd 0.028648f
C750 plus.n46 gnd 0.008502f
C751 plus.n47 gnd 0.173132f
C752 plus.n48 gnd 0.251919f
C753 plus.n49 gnd 0.021953f
C754 plus.t10 gnd 0.369143f
C755 plus.n50 gnd 0.149298f
C756 plus.n51 gnd 0.021953f
C757 plus.t15 gnd 0.369143f
C758 plus.n52 gnd 0.018183f
C759 plus.n53 gnd 0.021953f
C760 plus.t13 gnd 0.369143f
C761 plus.t17 gnd 0.369143f
C762 plus.n54 gnd 0.149298f
C763 plus.n55 gnd 0.021953f
C764 plus.t16 gnd 0.369143f
C765 plus.n56 gnd 0.149298f
C766 plus.n57 gnd 0.021953f
C767 plus.t20 gnd 0.369143f
C768 plus.n58 gnd 0.018183f
C769 plus.n59 gnd 0.021953f
C770 plus.t21 gnd 0.369143f
C771 plus.t5 gnd 0.369143f
C772 plus.n60 gnd 0.171686f
C773 plus.t11 gnd 0.413712f
C774 plus.n61 gnd 0.173884f
C775 plus.n62 gnd 0.093702f
C776 plus.n63 gnd 0.027719f
C777 plus.n64 gnd 0.025254f
C778 plus.n65 gnd 0.149298f
C779 plus.n66 gnd 0.026943f
C780 plus.n67 gnd 0.021953f
C781 plus.n68 gnd 0.021953f
C782 plus.n69 gnd 0.021953f
C783 plus.n70 gnd 0.028459f
C784 plus.n71 gnd 0.149298f
C785 plus.n72 gnd 0.026897f
C786 plus.n73 gnd 0.026075f
C787 plus.n74 gnd 0.021953f
C788 plus.n75 gnd 0.021953f
C789 plus.n76 gnd 0.027927f
C790 plus.n77 gnd 0.017731f
C791 plus.n78 gnd 0.027927f
C792 plus.n79 gnd 0.021953f
C793 plus.n80 gnd 0.021953f
C794 plus.n81 gnd 0.026075f
C795 plus.n82 gnd 0.026897f
C796 plus.n83 gnd 0.149298f
C797 plus.n84 gnd 0.028459f
C798 plus.n85 gnd 0.021953f
C799 plus.n86 gnd 0.021953f
C800 plus.n87 gnd 0.021953f
C801 plus.n88 gnd 0.026943f
C802 plus.n89 gnd 0.149298f
C803 plus.n90 gnd 0.025254f
C804 plus.n91 gnd 0.027719f
C805 plus.n92 gnd 0.021953f
C806 plus.n93 gnd 0.021953f
C807 plus.n94 gnd 0.028648f
C808 plus.n95 gnd 0.008502f
C809 plus.t23 gnd 0.399228f
C810 plus.n96 gnd 0.173132f
C811 plus.n97 gnd 0.733225f
C812 plus.n98 gnd 1.09402f
C813 plus.t1 gnd 0.037898f
C814 plus.t2 gnd 0.006768f
C815 plus.t4 gnd 0.006768f
C816 plus.n99 gnd 0.021948f
C817 plus.n100 gnd 0.170388f
C818 plus.t0 gnd 0.006768f
C819 plus.t3 gnd 0.006768f
C820 plus.n101 gnd 0.021948f
C821 plus.n102 gnd 0.127897f
C822 plus.n103 gnd 3.01173f
C823 a_n8300_8799.n0 gnd 0.884806f
C824 a_n8300_8799.n1 gnd 3.63607f
C825 a_n8300_8799.n2 gnd 3.37542f
C826 a_n8300_8799.n3 gnd 1.67746f
C827 a_n8300_8799.n4 gnd 0.17874f
C828 a_n8300_8799.n5 gnd 0.209316f
C829 a_n8300_8799.n6 gnd 0.209316f
C830 a_n8300_8799.n7 gnd 0.209316f
C831 a_n8300_8799.n8 gnd 0.17874f
C832 a_n8300_8799.n9 gnd 0.209316f
C833 a_n8300_8799.n10 gnd 0.209316f
C834 a_n8300_8799.n11 gnd 0.209316f
C835 a_n8300_8799.n12 gnd 0.345263f
C836 a_n8300_8799.n13 gnd 0.209316f
C837 a_n8300_8799.n14 gnd 0.209316f
C838 a_n8300_8799.n15 gnd 0.209316f
C839 a_n8300_8799.n16 gnd 0.209316f
C840 a_n8300_8799.n17 gnd 0.209316f
C841 a_n8300_8799.n18 gnd 0.17874f
C842 a_n8300_8799.n19 gnd 0.209316f
C843 a_n8300_8799.n20 gnd 0.209316f
C844 a_n8300_8799.n21 gnd 0.209316f
C845 a_n8300_8799.n22 gnd 0.17874f
C846 a_n8300_8799.n23 gnd 0.209316f
C847 a_n8300_8799.n24 gnd 0.209316f
C848 a_n8300_8799.n25 gnd 0.209316f
C849 a_n8300_8799.n26 gnd 0.345263f
C850 a_n8300_8799.n27 gnd 0.209316f
C851 a_n8300_8799.n28 gnd 1.0276f
C852 a_n8300_8799.n29 gnd 1.01304f
C853 a_n8300_8799.n30 gnd 3.00728f
C854 a_n8300_8799.n31 gnd 1.53412f
C855 a_n8300_8799.n32 gnd 1.01304f
C856 a_n8300_8799.n33 gnd 0.253132f
C857 a_n8300_8799.n35 gnd 0.007796f
C858 a_n8300_8799.n36 gnd 0.011784f
C859 a_n8300_8799.n37 gnd 0.008104f
C860 a_n8300_8799.n39 gnd 4.05e-19
C861 a_n8300_8799.n40 gnd 0.008399f
C862 a_n8300_8799.n41 gnd 0.264806f
C863 a_n8300_8799.n42 gnd 0.253132f
C864 a_n8300_8799.n44 gnd 0.007796f
C865 a_n8300_8799.n45 gnd 0.011784f
C866 a_n8300_8799.n46 gnd 0.008104f
C867 a_n8300_8799.n48 gnd 4.05e-19
C868 a_n8300_8799.n49 gnd 0.008399f
C869 a_n8300_8799.n50 gnd 0.264806f
C870 a_n8300_8799.n51 gnd 0.253132f
C871 a_n8300_8799.n53 gnd 0.007796f
C872 a_n8300_8799.n54 gnd 0.011784f
C873 a_n8300_8799.n55 gnd 0.008104f
C874 a_n8300_8799.n57 gnd 4.05e-19
C875 a_n8300_8799.n58 gnd 0.008399f
C876 a_n8300_8799.n59 gnd 0.264806f
C877 a_n8300_8799.n60 gnd 0.008399f
C878 a_n8300_8799.n61 gnd 0.264806f
C879 a_n8300_8799.n62 gnd 4.05e-19
C880 a_n8300_8799.n64 gnd 0.008104f
C881 a_n8300_8799.n65 gnd 0.011784f
C882 a_n8300_8799.n66 gnd 0.007796f
C883 a_n8300_8799.n68 gnd 0.253132f
C884 a_n8300_8799.n69 gnd 0.008399f
C885 a_n8300_8799.n70 gnd 0.264806f
C886 a_n8300_8799.n71 gnd 4.05e-19
C887 a_n8300_8799.n73 gnd 0.008104f
C888 a_n8300_8799.n74 gnd 0.011784f
C889 a_n8300_8799.n75 gnd 0.007796f
C890 a_n8300_8799.n77 gnd 0.253132f
C891 a_n8300_8799.n78 gnd 0.008399f
C892 a_n8300_8799.n79 gnd 0.264806f
C893 a_n8300_8799.n80 gnd 4.05e-19
C894 a_n8300_8799.n82 gnd 0.008104f
C895 a_n8300_8799.n83 gnd 0.011784f
C896 a_n8300_8799.n84 gnd 0.007796f
C897 a_n8300_8799.n86 gnd 0.253132f
C898 a_n8300_8799.t26 gnd 0.145184f
C899 a_n8300_8799.t28 gnd 0.145184f
C900 a_n8300_8799.t21 gnd 0.145184f
C901 a_n8300_8799.n87 gnd 1.14509f
C902 a_n8300_8799.t35 gnd 0.145184f
C903 a_n8300_8799.t27 gnd 0.145184f
C904 a_n8300_8799.n88 gnd 1.1432f
C905 a_n8300_8799.t19 gnd 0.145184f
C906 a_n8300_8799.t17 gnd 0.145184f
C907 a_n8300_8799.n89 gnd 1.1432f
C908 a_n8300_8799.t23 gnd 0.145184f
C909 a_n8300_8799.t15 gnd 0.145184f
C910 a_n8300_8799.n90 gnd 1.1432f
C911 a_n8300_8799.t32 gnd 0.145184f
C912 a_n8300_8799.t22 gnd 0.145184f
C913 a_n8300_8799.n91 gnd 1.1432f
C914 a_n8300_8799.t33 gnd 0.145184f
C915 a_n8300_8799.t16 gnd 0.145184f
C916 a_n8300_8799.n92 gnd 1.1432f
C917 a_n8300_8799.t8 gnd 0.112921f
C918 a_n8300_8799.t1 gnd 0.112921f
C919 a_n8300_8799.n93 gnd 1.00075f
C920 a_n8300_8799.t38 gnd 0.112921f
C921 a_n8300_8799.t37 gnd 0.112921f
C922 a_n8300_8799.n94 gnd 0.997808f
C923 a_n8300_8799.t10 gnd 0.112921f
C924 a_n8300_8799.t43 gnd 0.112921f
C925 a_n8300_8799.n95 gnd 0.997808f
C926 a_n8300_8799.t5 gnd 0.112921f
C927 a_n8300_8799.t9 gnd 0.112921f
C928 a_n8300_8799.n96 gnd 1.00075f
C929 a_n8300_8799.t0 gnd 0.112921f
C930 a_n8300_8799.t4 gnd 0.112921f
C931 a_n8300_8799.n97 gnd 0.997807f
C932 a_n8300_8799.t41 gnd 0.112921f
C933 a_n8300_8799.t7 gnd 0.112921f
C934 a_n8300_8799.n98 gnd 0.997807f
C935 a_n8300_8799.t39 gnd 0.112921f
C936 a_n8300_8799.t40 gnd 0.112921f
C937 a_n8300_8799.n99 gnd 1.00075f
C938 a_n8300_8799.t12 gnd 0.112921f
C939 a_n8300_8799.t2 gnd 0.112921f
C940 a_n8300_8799.n100 gnd 0.997807f
C941 a_n8300_8799.t11 gnd 0.112921f
C942 a_n8300_8799.t42 gnd 0.112921f
C943 a_n8300_8799.n101 gnd 0.997808f
C944 a_n8300_8799.t6 gnd 0.112921f
C945 a_n8300_8799.t3 gnd 0.112921f
C946 a_n8300_8799.n102 gnd 0.997808f
C947 a_n8300_8799.t70 gnd 0.602f
C948 a_n8300_8799.n103 gnd 0.272459f
C949 a_n8300_8799.t71 gnd 0.602f
C950 a_n8300_8799.t90 gnd 0.602f
C951 a_n8300_8799.n104 gnd 0.263541f
C952 a_n8300_8799.t103 gnd 0.602f
C953 a_n8300_8799.n105 gnd 0.275011f
C954 a_n8300_8799.t104 gnd 0.602f
C955 a_n8300_8799.t61 gnd 0.602f
C956 a_n8300_8799.n106 gnd 0.268381f
C957 a_n8300_8799.t85 gnd 0.616149f
C958 a_n8300_8799.t107 gnd 0.602f
C959 a_n8300_8799.n107 gnd 0.274573f
C960 a_n8300_8799.n108 gnd 0.250946f
C961 a_n8300_8799.t83 gnd 0.602f
C962 a_n8300_8799.n109 gnd 0.27234f
C963 a_n8300_8799.n110 gnd 0.272474f
C964 a_n8300_8799.t72 gnd 0.602f
C965 a_n8300_8799.n111 gnd 0.268703f
C966 a_n8300_8799.t102 gnd 0.602f
C967 a_n8300_8799.n112 gnd 0.268955f
C968 a_n8300_8799.n113 gnd 0.274573f
C969 a_n8300_8799.t88 gnd 0.612929f
C970 a_n8300_8799.t75 gnd 0.602f
C971 a_n8300_8799.n114 gnd 0.272459f
C972 a_n8300_8799.t76 gnd 0.602f
C973 a_n8300_8799.t99 gnd 0.602f
C974 a_n8300_8799.n115 gnd 0.263541f
C975 a_n8300_8799.t112 gnd 0.602f
C976 a_n8300_8799.n116 gnd 0.275011f
C977 a_n8300_8799.t114 gnd 0.602f
C978 a_n8300_8799.t67 gnd 0.602f
C979 a_n8300_8799.n117 gnd 0.268381f
C980 a_n8300_8799.t92 gnd 0.616149f
C981 a_n8300_8799.t115 gnd 0.602f
C982 a_n8300_8799.n118 gnd 0.274573f
C983 a_n8300_8799.n119 gnd 0.250946f
C984 a_n8300_8799.t89 gnd 0.602f
C985 a_n8300_8799.n120 gnd 0.27234f
C986 a_n8300_8799.n121 gnd 0.272474f
C987 a_n8300_8799.t79 gnd 0.602f
C988 a_n8300_8799.n122 gnd 0.268703f
C989 a_n8300_8799.t111 gnd 0.602f
C990 a_n8300_8799.n123 gnd 0.268955f
C991 a_n8300_8799.n124 gnd 0.274573f
C992 a_n8300_8799.t97 gnd 0.612929f
C993 a_n8300_8799.n125 gnd 0.903767f
C994 a_n8300_8799.t54 gnd 0.602f
C995 a_n8300_8799.n126 gnd 0.272459f
C996 a_n8300_8799.t44 gnd 0.602f
C997 a_n8300_8799.t68 gnd 0.602f
C998 a_n8300_8799.n127 gnd 0.263541f
C999 a_n8300_8799.t86 gnd 0.602f
C1000 a_n8300_8799.n128 gnd 0.275011f
C1001 a_n8300_8799.t74 gnd 0.602f
C1002 a_n8300_8799.t77 gnd 0.602f
C1003 a_n8300_8799.n129 gnd 0.268381f
C1004 a_n8300_8799.t94 gnd 0.616149f
C1005 a_n8300_8799.t63 gnd 0.602f
C1006 a_n8300_8799.n130 gnd 0.274573f
C1007 a_n8300_8799.n131 gnd 0.250946f
C1008 a_n8300_8799.t50 gnd 0.602f
C1009 a_n8300_8799.n132 gnd 0.27234f
C1010 a_n8300_8799.n133 gnd 0.272474f
C1011 a_n8300_8799.t98 gnd 0.602f
C1012 a_n8300_8799.n134 gnd 0.268703f
C1013 a_n8300_8799.t105 gnd 0.602f
C1014 a_n8300_8799.n135 gnd 0.268955f
C1015 a_n8300_8799.n136 gnd 0.274573f
C1016 a_n8300_8799.t80 gnd 0.612929f
C1017 a_n8300_8799.n137 gnd 1.91075f
C1018 a_n8300_8799.t47 gnd 0.612929f
C1019 a_n8300_8799.t46 gnd 0.602f
C1020 a_n8300_8799.t96 gnd 0.602f
C1021 a_n8300_8799.t57 gnd 0.602f
C1022 a_n8300_8799.n138 gnd 0.268955f
C1023 a_n8300_8799.t49 gnd 0.602f
C1024 a_n8300_8799.t100 gnd 0.602f
C1025 a_n8300_8799.t73 gnd 0.602f
C1026 a_n8300_8799.n139 gnd 0.272474f
C1027 a_n8300_8799.t58 gnd 0.602f
C1028 a_n8300_8799.t113 gnd 0.602f
C1029 a_n8300_8799.t84 gnd 0.602f
C1030 a_n8300_8799.n140 gnd 0.268381f
C1031 a_n8300_8799.t109 gnd 0.616149f
C1032 a_n8300_8799.t60 gnd 0.602f
C1033 a_n8300_8799.n141 gnd 0.274573f
C1034 a_n8300_8799.n142 gnd 0.250946f
C1035 a_n8300_8799.n143 gnd 0.27234f
C1036 a_n8300_8799.n144 gnd 0.275011f
C1037 a_n8300_8799.n145 gnd 0.268703f
C1038 a_n8300_8799.n146 gnd 0.263541f
C1039 a_n8300_8799.n147 gnd 0.272459f
C1040 a_n8300_8799.n148 gnd 0.274573f
C1041 a_n8300_8799.t53 gnd 0.612929f
C1042 a_n8300_8799.t52 gnd 0.602f
C1043 a_n8300_8799.t108 gnd 0.602f
C1044 a_n8300_8799.t62 gnd 0.602f
C1045 a_n8300_8799.n149 gnd 0.268955f
C1046 a_n8300_8799.t56 gnd 0.602f
C1047 a_n8300_8799.t110 gnd 0.602f
C1048 a_n8300_8799.t82 gnd 0.602f
C1049 a_n8300_8799.n150 gnd 0.272474f
C1050 a_n8300_8799.t65 gnd 0.602f
C1051 a_n8300_8799.t48 gnd 0.602f
C1052 a_n8300_8799.t91 gnd 0.602f
C1053 a_n8300_8799.n151 gnd 0.268381f
C1054 a_n8300_8799.t45 gnd 0.616149f
C1055 a_n8300_8799.t66 gnd 0.602f
C1056 a_n8300_8799.n152 gnd 0.274573f
C1057 a_n8300_8799.n153 gnd 0.250946f
C1058 a_n8300_8799.n154 gnd 0.27234f
C1059 a_n8300_8799.n155 gnd 0.275011f
C1060 a_n8300_8799.n156 gnd 0.268703f
C1061 a_n8300_8799.n157 gnd 0.263541f
C1062 a_n8300_8799.n158 gnd 0.272459f
C1063 a_n8300_8799.n159 gnd 0.274573f
C1064 a_n8300_8799.n160 gnd 0.903767f
C1065 a_n8300_8799.t81 gnd 0.612929f
C1066 a_n8300_8799.t95 gnd 0.602f
C1067 a_n8300_8799.t55 gnd 0.602f
C1068 a_n8300_8799.t106 gnd 0.602f
C1069 a_n8300_8799.n161 gnd 0.268955f
C1070 a_n8300_8799.t69 gnd 0.602f
C1071 a_n8300_8799.t101 gnd 0.602f
C1072 a_n8300_8799.t59 gnd 0.602f
C1073 a_n8300_8799.n162 gnd 0.272474f
C1074 a_n8300_8799.t87 gnd 0.602f
C1075 a_n8300_8799.t51 gnd 0.602f
C1076 a_n8300_8799.t78 gnd 0.602f
C1077 a_n8300_8799.n163 gnd 0.268381f
C1078 a_n8300_8799.t93 gnd 0.616149f
C1079 a_n8300_8799.t64 gnd 0.602f
C1080 a_n8300_8799.n164 gnd 0.274573f
C1081 a_n8300_8799.n165 gnd 0.250946f
C1082 a_n8300_8799.n166 gnd 0.27234f
C1083 a_n8300_8799.n167 gnd 0.275011f
C1084 a_n8300_8799.n168 gnd 0.268703f
C1085 a_n8300_8799.n169 gnd 0.263541f
C1086 a_n8300_8799.n170 gnd 0.272459f
C1087 a_n8300_8799.n171 gnd 0.274573f
C1088 a_n8300_8799.n172 gnd 1.38704f
C1089 a_n8300_8799.n173 gnd 17.483099f
C1090 a_n8300_8799.n174 gnd 4.40577f
C1091 a_n8300_8799.n175 gnd 7.68044f
C1092 a_n8300_8799.t34 gnd 0.145184f
C1093 a_n8300_8799.t29 gnd 0.145184f
C1094 a_n8300_8799.n176 gnd 1.14508f
C1095 a_n8300_8799.t25 gnd 0.145184f
C1096 a_n8300_8799.t18 gnd 0.145184f
C1097 a_n8300_8799.n177 gnd 1.1432f
C1098 a_n8300_8799.t36 gnd 0.145184f
C1099 a_n8300_8799.t14 gnd 0.145184f
C1100 a_n8300_8799.n178 gnd 1.1432f
C1101 a_n8300_8799.t30 gnd 0.145184f
C1102 a_n8300_8799.t24 gnd 0.145184f
C1103 a_n8300_8799.n179 gnd 1.1432f
C1104 a_n8300_8799.t20 gnd 0.145184f
C1105 a_n8300_8799.t31 gnd 0.145184f
C1106 a_n8300_8799.n180 gnd 1.1432f
C1107 a_n8300_8799.n181 gnd 3.73873f
C1108 a_n8300_8799.n182 gnd 1.1432f
C1109 a_n8300_8799.t13 gnd 0.145184f
C1110 CSoutput.n0 gnd 0.042073f
C1111 CSoutput.t197 gnd 0.278303f
C1112 CSoutput.n1 gnd 0.125668f
C1113 CSoutput.n2 gnd 0.042073f
C1114 CSoutput.t204 gnd 0.278303f
C1115 CSoutput.n3 gnd 0.033346f
C1116 CSoutput.n4 gnd 0.042073f
C1117 CSoutput.t213 gnd 0.278303f
C1118 CSoutput.n5 gnd 0.028755f
C1119 CSoutput.n6 gnd 0.042073f
C1120 CSoutput.t202 gnd 0.278303f
C1121 CSoutput.t199 gnd 0.278303f
C1122 CSoutput.n7 gnd 0.124298f
C1123 CSoutput.n8 gnd 0.042073f
C1124 CSoutput.t211 gnd 0.278303f
C1125 CSoutput.n9 gnd 0.027416f
C1126 CSoutput.n10 gnd 0.042073f
C1127 CSoutput.t192 gnd 0.278303f
C1128 CSoutput.t195 gnd 0.278303f
C1129 CSoutput.n11 gnd 0.124298f
C1130 CSoutput.n12 gnd 0.042073f
C1131 CSoutput.t208 gnd 0.278303f
C1132 CSoutput.n13 gnd 0.028755f
C1133 CSoutput.n14 gnd 0.042073f
C1134 CSoutput.t207 gnd 0.278303f
C1135 CSoutput.t193 gnd 0.278303f
C1136 CSoutput.n15 gnd 0.124298f
C1137 CSoutput.n16 gnd 0.042073f
C1138 CSoutput.t198 gnd 0.278303f
C1139 CSoutput.n17 gnd 0.030711f
C1140 CSoutput.t209 gnd 0.33258f
C1141 CSoutput.t205 gnd 0.278303f
C1142 CSoutput.n18 gnd 0.15868f
C1143 CSoutput.n19 gnd 0.153975f
C1144 CSoutput.n20 gnd 0.178629f
C1145 CSoutput.n21 gnd 0.042073f
C1146 CSoutput.n22 gnd 0.035114f
C1147 CSoutput.n23 gnd 0.124298f
C1148 CSoutput.n24 gnd 0.033849f
C1149 CSoutput.n25 gnd 0.033346f
C1150 CSoutput.n26 gnd 0.042073f
C1151 CSoutput.n27 gnd 0.042073f
C1152 CSoutput.n28 gnd 0.034844f
C1153 CSoutput.n29 gnd 0.029584f
C1154 CSoutput.n30 gnd 0.127065f
C1155 CSoutput.n31 gnd 0.029991f
C1156 CSoutput.n32 gnd 0.042073f
C1157 CSoutput.n33 gnd 0.042073f
C1158 CSoutput.n34 gnd 0.042073f
C1159 CSoutput.n35 gnd 0.034473f
C1160 CSoutput.n36 gnd 0.124298f
C1161 CSoutput.n37 gnd 0.032969f
C1162 CSoutput.n38 gnd 0.034227f
C1163 CSoutput.n39 gnd 0.042073f
C1164 CSoutput.n40 gnd 0.042073f
C1165 CSoutput.n41 gnd 0.035107f
C1166 CSoutput.n42 gnd 0.032088f
C1167 CSoutput.n43 gnd 0.124298f
C1168 CSoutput.n44 gnd 0.032902f
C1169 CSoutput.n45 gnd 0.042073f
C1170 CSoutput.n46 gnd 0.042073f
C1171 CSoutput.n47 gnd 0.042073f
C1172 CSoutput.n48 gnd 0.032902f
C1173 CSoutput.n49 gnd 0.124298f
C1174 CSoutput.n50 gnd 0.032088f
C1175 CSoutput.n51 gnd 0.035107f
C1176 CSoutput.n52 gnd 0.042073f
C1177 CSoutput.n53 gnd 0.042073f
C1178 CSoutput.n54 gnd 0.034227f
C1179 CSoutput.n55 gnd 0.032969f
C1180 CSoutput.n56 gnd 0.124298f
C1181 CSoutput.n57 gnd 0.034473f
C1182 CSoutput.n58 gnd 0.042073f
C1183 CSoutput.n59 gnd 0.042073f
C1184 CSoutput.n60 gnd 0.042073f
C1185 CSoutput.n61 gnd 0.029991f
C1186 CSoutput.n62 gnd 0.127065f
C1187 CSoutput.n63 gnd 0.029584f
C1188 CSoutput.t203 gnd 0.278303f
C1189 CSoutput.n64 gnd 0.124298f
C1190 CSoutput.n65 gnd 0.034844f
C1191 CSoutput.n66 gnd 0.042073f
C1192 CSoutput.n67 gnd 0.042073f
C1193 CSoutput.n68 gnd 0.042073f
C1194 CSoutput.n69 gnd 0.033849f
C1195 CSoutput.n70 gnd 0.124298f
C1196 CSoutput.n71 gnd 0.035114f
C1197 CSoutput.n72 gnd 0.030711f
C1198 CSoutput.n73 gnd 0.042073f
C1199 CSoutput.n74 gnd 0.042073f
C1200 CSoutput.n75 gnd 0.03185f
C1201 CSoutput.n76 gnd 0.018916f
C1202 CSoutput.t212 gnd 0.312693f
C1203 CSoutput.n77 gnd 0.155333f
C1204 CSoutput.n78 gnd 0.635462f
C1205 CSoutput.t10 gnd 0.05248f
C1206 CSoutput.t6 gnd 0.05248f
C1207 CSoutput.n79 gnd 0.406318f
C1208 CSoutput.t179 gnd 0.05248f
C1209 CSoutput.t168 gnd 0.05248f
C1210 CSoutput.n80 gnd 0.405593f
C1211 CSoutput.n81 gnd 0.411677f
C1212 CSoutput.t180 gnd 0.05248f
C1213 CSoutput.t174 gnd 0.05248f
C1214 CSoutput.n82 gnd 0.405593f
C1215 CSoutput.n83 gnd 0.202857f
C1216 CSoutput.t32 gnd 0.05248f
C1217 CSoutput.t190 gnd 0.05248f
C1218 CSoutput.n84 gnd 0.405593f
C1219 CSoutput.n85 gnd 0.202857f
C1220 CSoutput.t21 gnd 0.05248f
C1221 CSoutput.t26 gnd 0.05248f
C1222 CSoutput.n86 gnd 0.405593f
C1223 CSoutput.n87 gnd 0.202857f
C1224 CSoutput.t188 gnd 0.05248f
C1225 CSoutput.t15 gnd 0.05248f
C1226 CSoutput.n88 gnd 0.405593f
C1227 CSoutput.n89 gnd 0.371993f
C1228 CSoutput.t20 gnd 0.05248f
C1229 CSoutput.t13 gnd 0.05248f
C1230 CSoutput.n90 gnd 0.406318f
C1231 CSoutput.t31 gnd 0.05248f
C1232 CSoutput.t191 gnd 0.05248f
C1233 CSoutput.n91 gnd 0.405593f
C1234 CSoutput.n92 gnd 0.411677f
C1235 CSoutput.t9 gnd 0.05248f
C1236 CSoutput.t181 gnd 0.05248f
C1237 CSoutput.n93 gnd 0.405593f
C1238 CSoutput.n94 gnd 0.202857f
C1239 CSoutput.t176 gnd 0.05248f
C1240 CSoutput.t2 gnd 0.05248f
C1241 CSoutput.n95 gnd 0.405593f
C1242 CSoutput.n96 gnd 0.202857f
C1243 CSoutput.t25 gnd 0.05248f
C1244 CSoutput.t173 gnd 0.05248f
C1245 CSoutput.n97 gnd 0.405593f
C1246 CSoutput.n98 gnd 0.202857f
C1247 CSoutput.t42 gnd 0.05248f
C1248 CSoutput.t3 gnd 0.05248f
C1249 CSoutput.n99 gnd 0.405593f
C1250 CSoutput.n100 gnd 0.302511f
C1251 CSoutput.n101 gnd 0.381464f
C1252 CSoutput.t45 gnd 0.05248f
C1253 CSoutput.t172 gnd 0.05248f
C1254 CSoutput.n102 gnd 0.406318f
C1255 CSoutput.t36 gnd 0.05248f
C1256 CSoutput.t44 gnd 0.05248f
C1257 CSoutput.n103 gnd 0.405593f
C1258 CSoutput.n104 gnd 0.411677f
C1259 CSoutput.t22 gnd 0.05248f
C1260 CSoutput.t4 gnd 0.05248f
C1261 CSoutput.n105 gnd 0.405593f
C1262 CSoutput.n106 gnd 0.202857f
C1263 CSoutput.t37 gnd 0.05248f
C1264 CSoutput.t178 gnd 0.05248f
C1265 CSoutput.n107 gnd 0.405593f
C1266 CSoutput.n108 gnd 0.202857f
C1267 CSoutput.t47 gnd 0.05248f
C1268 CSoutput.t17 gnd 0.05248f
C1269 CSoutput.n109 gnd 0.405593f
C1270 CSoutput.n110 gnd 0.202857f
C1271 CSoutput.t29 gnd 0.05248f
C1272 CSoutput.t185 gnd 0.05248f
C1273 CSoutput.n111 gnd 0.405593f
C1274 CSoutput.n112 gnd 0.302511f
C1275 CSoutput.n113 gnd 0.426379f
C1276 CSoutput.n114 gnd 8.95057f
C1277 CSoutput.n116 gnd 0.744262f
C1278 CSoutput.n117 gnd 0.558197f
C1279 CSoutput.n118 gnd 0.744262f
C1280 CSoutput.n119 gnd 0.744262f
C1281 CSoutput.n120 gnd 2.00378f
C1282 CSoutput.n121 gnd 0.744262f
C1283 CSoutput.n122 gnd 0.744262f
C1284 CSoutput.t201 gnd 0.930328f
C1285 CSoutput.n123 gnd 0.744262f
C1286 CSoutput.n124 gnd 0.744262f
C1287 CSoutput.n128 gnd 0.744262f
C1288 CSoutput.n132 gnd 0.744262f
C1289 CSoutput.n133 gnd 0.744262f
C1290 CSoutput.n135 gnd 0.744262f
C1291 CSoutput.n140 gnd 0.744262f
C1292 CSoutput.n142 gnd 0.744262f
C1293 CSoutput.n143 gnd 0.744262f
C1294 CSoutput.n145 gnd 0.744262f
C1295 CSoutput.n146 gnd 0.744262f
C1296 CSoutput.n148 gnd 0.744262f
C1297 CSoutput.t194 gnd 12.436501f
C1298 CSoutput.n150 gnd 0.744262f
C1299 CSoutput.n151 gnd 0.558197f
C1300 CSoutput.n152 gnd 0.744262f
C1301 CSoutput.n153 gnd 0.744262f
C1302 CSoutput.n154 gnd 2.00378f
C1303 CSoutput.n155 gnd 0.744262f
C1304 CSoutput.n156 gnd 0.744262f
C1305 CSoutput.t196 gnd 0.930328f
C1306 CSoutput.n157 gnd 0.744262f
C1307 CSoutput.n158 gnd 0.744262f
C1308 CSoutput.n162 gnd 0.744262f
C1309 CSoutput.n166 gnd 0.744262f
C1310 CSoutput.n167 gnd 0.744262f
C1311 CSoutput.n169 gnd 0.744262f
C1312 CSoutput.n174 gnd 0.744262f
C1313 CSoutput.n176 gnd 0.744262f
C1314 CSoutput.n177 gnd 0.744262f
C1315 CSoutput.n179 gnd 0.744262f
C1316 CSoutput.n180 gnd 0.744262f
C1317 CSoutput.n182 gnd 0.744262f
C1318 CSoutput.n183 gnd 0.558197f
C1319 CSoutput.n185 gnd 0.744262f
C1320 CSoutput.n186 gnd 0.558197f
C1321 CSoutput.n187 gnd 0.744262f
C1322 CSoutput.n188 gnd 0.744262f
C1323 CSoutput.n189 gnd 2.00378f
C1324 CSoutput.n190 gnd 0.744262f
C1325 CSoutput.n191 gnd 0.744262f
C1326 CSoutput.t200 gnd 0.930328f
C1327 CSoutput.n192 gnd 0.744262f
C1328 CSoutput.n193 gnd 2.00378f
C1329 CSoutput.n195 gnd 0.744262f
C1330 CSoutput.n196 gnd 0.744262f
C1331 CSoutput.n198 gnd 0.744262f
C1332 CSoutput.n199 gnd 0.744262f
C1333 CSoutput.t210 gnd 12.2339f
C1334 CSoutput.t206 gnd 12.436501f
C1335 CSoutput.n205 gnd 2.33486f
C1336 CSoutput.n206 gnd 9.511371f
C1337 CSoutput.n207 gnd 9.909361f
C1338 CSoutput.n212 gnd 2.52928f
C1339 CSoutput.n218 gnd 0.744262f
C1340 CSoutput.n220 gnd 0.744262f
C1341 CSoutput.n222 gnd 0.744262f
C1342 CSoutput.n224 gnd 0.744262f
C1343 CSoutput.n226 gnd 0.744262f
C1344 CSoutput.n232 gnd 0.744262f
C1345 CSoutput.n239 gnd 1.36543f
C1346 CSoutput.n240 gnd 1.36543f
C1347 CSoutput.n241 gnd 0.744262f
C1348 CSoutput.n242 gnd 0.744262f
C1349 CSoutput.n244 gnd 0.558197f
C1350 CSoutput.n245 gnd 0.478045f
C1351 CSoutput.n247 gnd 0.558197f
C1352 CSoutput.n248 gnd 0.478045f
C1353 CSoutput.n249 gnd 0.558197f
C1354 CSoutput.n251 gnd 0.744262f
C1355 CSoutput.n253 gnd 2.00378f
C1356 CSoutput.n254 gnd 2.33486f
C1357 CSoutput.n255 gnd 8.74801f
C1358 CSoutput.n257 gnd 0.558197f
C1359 CSoutput.n258 gnd 1.43627f
C1360 CSoutput.n259 gnd 0.558197f
C1361 CSoutput.n261 gnd 0.744262f
C1362 CSoutput.n263 gnd 2.00378f
C1363 CSoutput.n264 gnd 4.36456f
C1364 CSoutput.t7 gnd 0.05248f
C1365 CSoutput.t189 gnd 0.05248f
C1366 CSoutput.n265 gnd 0.406318f
C1367 CSoutput.t169 gnd 0.05248f
C1368 CSoutput.t184 gnd 0.05248f
C1369 CSoutput.n266 gnd 0.405593f
C1370 CSoutput.n267 gnd 0.411677f
C1371 CSoutput.t175 gnd 0.05248f
C1372 CSoutput.t187 gnd 0.05248f
C1373 CSoutput.n268 gnd 0.405593f
C1374 CSoutput.n269 gnd 0.202857f
C1375 CSoutput.t39 gnd 0.05248f
C1376 CSoutput.t33 gnd 0.05248f
C1377 CSoutput.n270 gnd 0.405593f
C1378 CSoutput.n271 gnd 0.202857f
C1379 CSoutput.t27 gnd 0.05248f
C1380 CSoutput.t8 gnd 0.05248f
C1381 CSoutput.n272 gnd 0.405593f
C1382 CSoutput.n273 gnd 0.202857f
C1383 CSoutput.t182 gnd 0.05248f
C1384 CSoutput.t43 gnd 0.05248f
C1385 CSoutput.n274 gnd 0.405593f
C1386 CSoutput.n275 gnd 0.371993f
C1387 CSoutput.t171 gnd 0.05248f
C1388 CSoutput.t170 gnd 0.05248f
C1389 CSoutput.n276 gnd 0.406318f
C1390 CSoutput.t34 gnd 0.05248f
C1391 CSoutput.t14 gnd 0.05248f
C1392 CSoutput.n277 gnd 0.405593f
C1393 CSoutput.n278 gnd 0.411677f
C1394 CSoutput.t18 gnd 0.05248f
C1395 CSoutput.t30 gnd 0.05248f
C1396 CSoutput.n279 gnd 0.405593f
C1397 CSoutput.n280 gnd 0.202857f
C1398 CSoutput.t16 gnd 0.05248f
C1399 CSoutput.t183 gnd 0.05248f
C1400 CSoutput.n281 gnd 0.405593f
C1401 CSoutput.n282 gnd 0.202857f
C1402 CSoutput.t40 gnd 0.05248f
C1403 CSoutput.t5 gnd 0.05248f
C1404 CSoutput.n283 gnd 0.405593f
C1405 CSoutput.n284 gnd 0.202857f
C1406 CSoutput.t24 gnd 0.05248f
C1407 CSoutput.t11 gnd 0.05248f
C1408 CSoutput.n285 gnd 0.405593f
C1409 CSoutput.n286 gnd 0.302511f
C1410 CSoutput.n287 gnd 0.381464f
C1411 CSoutput.t1 gnd 0.05248f
C1412 CSoutput.t0 gnd 0.05248f
C1413 CSoutput.n288 gnd 0.406318f
C1414 CSoutput.t12 gnd 0.05248f
C1415 CSoutput.t19 gnd 0.05248f
C1416 CSoutput.n289 gnd 0.405593f
C1417 CSoutput.n290 gnd 0.411677f
C1418 CSoutput.t41 gnd 0.05248f
C1419 CSoutput.t186 gnd 0.05248f
C1420 CSoutput.n291 gnd 0.405593f
C1421 CSoutput.n292 gnd 0.202857f
C1422 CSoutput.t23 gnd 0.05248f
C1423 CSoutput.t38 gnd 0.05248f
C1424 CSoutput.n293 gnd 0.405593f
C1425 CSoutput.n294 gnd 0.202857f
C1426 CSoutput.t177 gnd 0.05248f
C1427 CSoutput.t28 gnd 0.05248f
C1428 CSoutput.n295 gnd 0.405593f
C1429 CSoutput.n296 gnd 0.202857f
C1430 CSoutput.t46 gnd 0.05248f
C1431 CSoutput.t35 gnd 0.05248f
C1432 CSoutput.n297 gnd 0.405592f
C1433 CSoutput.n298 gnd 0.302512f
C1434 CSoutput.n299 gnd 0.426379f
C1435 CSoutput.n300 gnd 12.3032f
C1436 CSoutput.t143 gnd 0.04592f
C1437 CSoutput.t66 gnd 0.04592f
C1438 CSoutput.n301 gnd 0.407123f
C1439 CSoutput.t123 gnd 0.04592f
C1440 CSoutput.t50 gnd 0.04592f
C1441 CSoutput.n302 gnd 0.405765f
C1442 CSoutput.n303 gnd 0.378098f
C1443 CSoutput.t105 gnd 0.04592f
C1444 CSoutput.t146 gnd 0.04592f
C1445 CSoutput.n304 gnd 0.405765f
C1446 CSoutput.n305 gnd 0.186384f
C1447 CSoutput.t91 gnd 0.04592f
C1448 CSoutput.t104 gnd 0.04592f
C1449 CSoutput.n306 gnd 0.405765f
C1450 CSoutput.n307 gnd 0.186384f
C1451 CSoutput.t54 gnd 0.04592f
C1452 CSoutput.t111 gnd 0.04592f
C1453 CSoutput.n308 gnd 0.405765f
C1454 CSoutput.n309 gnd 0.186384f
C1455 CSoutput.t128 gnd 0.04592f
C1456 CSoutput.t92 gnd 0.04592f
C1457 CSoutput.n310 gnd 0.405765f
C1458 CSoutput.n311 gnd 0.186384f
C1459 CSoutput.t107 gnd 0.04592f
C1460 CSoutput.t138 gnd 0.04592f
C1461 CSoutput.n312 gnd 0.405765f
C1462 CSoutput.n313 gnd 0.186384f
C1463 CSoutput.t65 gnd 0.04592f
C1464 CSoutput.t81 gnd 0.04592f
C1465 CSoutput.n314 gnd 0.405765f
C1466 CSoutput.n315 gnd 0.186384f
C1467 CSoutput.t124 gnd 0.04592f
C1468 CSoutput.t163 gnd 0.04592f
C1469 CSoutput.n316 gnd 0.405765f
C1470 CSoutput.n317 gnd 0.186384f
C1471 CSoutput.t116 gnd 0.04592f
C1472 CSoutput.t147 gnd 0.04592f
C1473 CSoutput.n318 gnd 0.405765f
C1474 CSoutput.n319 gnd 0.343776f
C1475 CSoutput.t102 gnd 0.04592f
C1476 CSoutput.t75 gnd 0.04592f
C1477 CSoutput.n320 gnd 0.407123f
C1478 CSoutput.t87 gnd 0.04592f
C1479 CSoutput.t101 gnd 0.04592f
C1480 CSoutput.n321 gnd 0.405765f
C1481 CSoutput.n322 gnd 0.378098f
C1482 CSoutput.t74 gnd 0.04592f
C1483 CSoutput.t89 gnd 0.04592f
C1484 CSoutput.n323 gnd 0.405765f
C1485 CSoutput.n324 gnd 0.186384f
C1486 CSoutput.t103 gnd 0.04592f
C1487 CSoutput.t73 gnd 0.04592f
C1488 CSoutput.n325 gnd 0.405765f
C1489 CSoutput.n326 gnd 0.186384f
C1490 CSoutput.t88 gnd 0.04592f
C1491 CSoutput.t62 gnd 0.04592f
C1492 CSoutput.n327 gnd 0.405765f
C1493 CSoutput.n328 gnd 0.186384f
C1494 CSoutput.t72 gnd 0.04592f
C1495 CSoutput.t90 gnd 0.04592f
C1496 CSoutput.n329 gnd 0.405765f
C1497 CSoutput.n330 gnd 0.186384f
C1498 CSoutput.t57 gnd 0.04592f
C1499 CSoutput.t156 gnd 0.04592f
C1500 CSoutput.n331 gnd 0.405765f
C1501 CSoutput.n332 gnd 0.186384f
C1502 CSoutput.t78 gnd 0.04592f
C1503 CSoutput.t165 gnd 0.04592f
C1504 CSoutput.n333 gnd 0.405765f
C1505 CSoutput.n334 gnd 0.186384f
C1506 CSoutput.t152 gnd 0.04592f
C1507 CSoutput.t157 gnd 0.04592f
C1508 CSoutput.n335 gnd 0.405765f
C1509 CSoutput.n336 gnd 0.186384f
C1510 CSoutput.t167 gnd 0.04592f
C1511 CSoutput.t153 gnd 0.04592f
C1512 CSoutput.n337 gnd 0.405765f
C1513 CSoutput.n338 gnd 0.282971f
C1514 CSoutput.n339 gnd 0.356915f
C1515 CSoutput.t64 gnd 0.04592f
C1516 CSoutput.t158 gnd 0.04592f
C1517 CSoutput.n340 gnd 0.407123f
C1518 CSoutput.t140 gnd 0.04592f
C1519 CSoutput.t79 gnd 0.04592f
C1520 CSoutput.n341 gnd 0.405765f
C1521 CSoutput.n342 gnd 0.378098f
C1522 CSoutput.t48 gnd 0.04592f
C1523 CSoutput.t149 gnd 0.04592f
C1524 CSoutput.n343 gnd 0.405765f
C1525 CSoutput.n344 gnd 0.186384f
C1526 CSoutput.t97 gnd 0.04592f
C1527 CSoutput.t106 gnd 0.04592f
C1528 CSoutput.n345 gnd 0.405765f
C1529 CSoutput.n346 gnd 0.186384f
C1530 CSoutput.t159 gnd 0.04592f
C1531 CSoutput.t139 gnd 0.04592f
C1532 CSoutput.n347 gnd 0.405765f
C1533 CSoutput.n348 gnd 0.186384f
C1534 CSoutput.t117 gnd 0.04592f
C1535 CSoutput.t49 gnd 0.04592f
C1536 CSoutput.n349 gnd 0.405765f
C1537 CSoutput.n350 gnd 0.186384f
C1538 CSoutput.t61 gnd 0.04592f
C1539 CSoutput.t155 gnd 0.04592f
C1540 CSoutput.n351 gnd 0.405765f
C1541 CSoutput.n352 gnd 0.186384f
C1542 CSoutput.t70 gnd 0.04592f
C1543 CSoutput.t77 gnd 0.04592f
C1544 CSoutput.n353 gnd 0.405765f
C1545 CSoutput.n354 gnd 0.186384f
C1546 CSoutput.t166 gnd 0.04592f
C1547 CSoutput.t148 gnd 0.04592f
C1548 CSoutput.n355 gnd 0.405765f
C1549 CSoutput.n356 gnd 0.186384f
C1550 CSoutput.t96 gnd 0.04592f
C1551 CSoutput.t63 gnd 0.04592f
C1552 CSoutput.n357 gnd 0.405765f
C1553 CSoutput.n358 gnd 0.282971f
C1554 CSoutput.n359 gnd 0.38327f
C1555 CSoutput.n360 gnd 12.9105f
C1556 CSoutput.t113 gnd 0.04592f
C1557 CSoutput.t56 gnd 0.04592f
C1558 CSoutput.n361 gnd 0.407123f
C1559 CSoutput.t95 gnd 0.04592f
C1560 CSoutput.t150 gnd 0.04592f
C1561 CSoutput.n362 gnd 0.405765f
C1562 CSoutput.n363 gnd 0.378098f
C1563 CSoutput.t60 gnd 0.04592f
C1564 CSoutput.t130 gnd 0.04592f
C1565 CSoutput.n364 gnd 0.405765f
C1566 CSoutput.n365 gnd 0.186384f
C1567 CSoutput.t129 gnd 0.04592f
C1568 CSoutput.t115 gnd 0.04592f
C1569 CSoutput.n366 gnd 0.405765f
C1570 CSoutput.n367 gnd 0.186384f
C1571 CSoutput.t133 gnd 0.04592f
C1572 CSoutput.t98 gnd 0.04592f
C1573 CSoutput.n368 gnd 0.405765f
C1574 CSoutput.n369 gnd 0.186384f
C1575 CSoutput.t125 gnd 0.04592f
C1576 CSoutput.t142 gnd 0.04592f
C1577 CSoutput.n370 gnd 0.405765f
C1578 CSoutput.n371 gnd 0.186384f
C1579 CSoutput.t164 gnd 0.04592f
C1580 CSoutput.t132 gnd 0.04592f
C1581 CSoutput.n372 gnd 0.405765f
C1582 CSoutput.n373 gnd 0.186384f
C1583 CSoutput.t137 gnd 0.04592f
C1584 CSoutput.t136 gnd 0.04592f
C1585 CSoutput.n374 gnd 0.405765f
C1586 CSoutput.n375 gnd 0.186384f
C1587 CSoutput.t120 gnd 0.04592f
C1588 CSoutput.t55 gnd 0.04592f
C1589 CSoutput.n376 gnd 0.405765f
C1590 CSoutput.n377 gnd 0.186384f
C1591 CSoutput.t94 gnd 0.04592f
C1592 CSoutput.t161 gnd 0.04592f
C1593 CSoutput.n378 gnd 0.405765f
C1594 CSoutput.n379 gnd 0.343776f
C1595 CSoutput.t99 gnd 0.04592f
C1596 CSoutput.t118 gnd 0.04592f
C1597 CSoutput.n380 gnd 0.407123f
C1598 CSoutput.t119 gnd 0.04592f
C1599 CSoutput.t108 gnd 0.04592f
C1600 CSoutput.n381 gnd 0.405765f
C1601 CSoutput.n382 gnd 0.378098f
C1602 CSoutput.t109 gnd 0.04592f
C1603 CSoutput.t100 gnd 0.04592f
C1604 CSoutput.n383 gnd 0.405765f
C1605 CSoutput.n384 gnd 0.186384f
C1606 CSoutput.t93 gnd 0.04592f
C1607 CSoutput.t85 gnd 0.04592f
C1608 CSoutput.n385 gnd 0.405765f
C1609 CSoutput.n386 gnd 0.186384f
C1610 CSoutput.t86 gnd 0.04592f
C1611 CSoutput.t110 gnd 0.04592f
C1612 CSoutput.n387 gnd 0.405765f
C1613 CSoutput.n388 gnd 0.186384f
C1614 CSoutput.t112 gnd 0.04592f
C1615 CSoutput.t52 gnd 0.04592f
C1616 CSoutput.n389 gnd 0.405765f
C1617 CSoutput.n390 gnd 0.186384f
C1618 CSoutput.t53 gnd 0.04592f
C1619 CSoutput.t76 gnd 0.04592f
C1620 CSoutput.n391 gnd 0.405765f
C1621 CSoutput.n392 gnd 0.186384f
C1622 CSoutput.t83 gnd 0.04592f
C1623 CSoutput.t71 gnd 0.04592f
C1624 CSoutput.n393 gnd 0.405765f
C1625 CSoutput.n394 gnd 0.186384f
C1626 CSoutput.t67 gnd 0.04592f
C1627 CSoutput.t58 gnd 0.04592f
C1628 CSoutput.n395 gnd 0.405765f
C1629 CSoutput.n396 gnd 0.186384f
C1630 CSoutput.t59 gnd 0.04592f
C1631 CSoutput.t84 gnd 0.04592f
C1632 CSoutput.n397 gnd 0.405765f
C1633 CSoutput.n398 gnd 0.282971f
C1634 CSoutput.n399 gnd 0.356915f
C1635 CSoutput.t134 gnd 0.04592f
C1636 CSoutput.t154 gnd 0.04592f
C1637 CSoutput.n400 gnd 0.407123f
C1638 CSoutput.t162 gnd 0.04592f
C1639 CSoutput.t122 gnd 0.04592f
C1640 CSoutput.n401 gnd 0.405765f
C1641 CSoutput.n402 gnd 0.378098f
C1642 CSoutput.t127 gnd 0.04592f
C1643 CSoutput.t144 gnd 0.04592f
C1644 CSoutput.n403 gnd 0.405765f
C1645 CSoutput.n404 gnd 0.186384f
C1646 CSoutput.t68 gnd 0.04592f
C1647 CSoutput.t114 gnd 0.04592f
C1648 CSoutput.n405 gnd 0.405765f
C1649 CSoutput.n406 gnd 0.186384f
C1650 CSoutput.t121 gnd 0.04592f
C1651 CSoutput.t135 gnd 0.04592f
C1652 CSoutput.n407 gnd 0.405765f
C1653 CSoutput.n408 gnd 0.186384f
C1654 CSoutput.t145 gnd 0.04592f
C1655 CSoutput.t126 gnd 0.04592f
C1656 CSoutput.n409 gnd 0.405765f
C1657 CSoutput.n410 gnd 0.186384f
C1658 CSoutput.t131 gnd 0.04592f
C1659 CSoutput.t151 gnd 0.04592f
C1660 CSoutput.n411 gnd 0.405765f
C1661 CSoutput.n412 gnd 0.186384f
C1662 CSoutput.t69 gnd 0.04592f
C1663 CSoutput.t80 gnd 0.04592f
C1664 CSoutput.n413 gnd 0.405765f
C1665 CSoutput.n414 gnd 0.186384f
C1666 CSoutput.t141 gnd 0.04592f
C1667 CSoutput.t160 gnd 0.04592f
C1668 CSoutput.n415 gnd 0.405765f
C1669 CSoutput.n416 gnd 0.186384f
C1670 CSoutput.t51 gnd 0.04592f
C1671 CSoutput.t82 gnd 0.04592f
C1672 CSoutput.n417 gnd 0.405765f
C1673 CSoutput.n418 gnd 0.282971f
C1674 CSoutput.n419 gnd 0.38327f
C1675 CSoutput.n420 gnd 7.872509f
C1676 CSoutput.n421 gnd 12.8911f
C1677 vdd.t204 gnd 0.032436f
C1678 vdd.t184 gnd 0.032436f
C1679 vdd.n0 gnd 0.255824f
C1680 vdd.t163 gnd 0.032436f
C1681 vdd.t200 gnd 0.032436f
C1682 vdd.n1 gnd 0.255401f
C1683 vdd.n2 gnd 0.235529f
C1684 vdd.t181 gnd 0.032436f
C1685 vdd.t211 gnd 0.032436f
C1686 vdd.n3 gnd 0.255401f
C1687 vdd.n4 gnd 0.119116f
C1688 vdd.t209 gnd 0.032436f
C1689 vdd.t189 gnd 0.032436f
C1690 vdd.n5 gnd 0.255401f
C1691 vdd.n6 gnd 0.111768f
C1692 vdd.t215 gnd 0.032436f
C1693 vdd.t179 gnd 0.032436f
C1694 vdd.n7 gnd 0.255824f
C1695 vdd.t187 gnd 0.032436f
C1696 vdd.t207 gnd 0.032436f
C1697 vdd.n8 gnd 0.255401f
C1698 vdd.n9 gnd 0.235529f
C1699 vdd.t196 gnd 0.032436f
C1700 vdd.t169 gnd 0.032436f
C1701 vdd.n10 gnd 0.255401f
C1702 vdd.n11 gnd 0.119116f
C1703 vdd.t165 gnd 0.032436f
C1704 vdd.t194 gnd 0.032436f
C1705 vdd.n12 gnd 0.255401f
C1706 vdd.n13 gnd 0.111768f
C1707 vdd.n14 gnd 0.079018f
C1708 vdd.t126 gnd 0.01802f
C1709 vdd.t141 gnd 0.01802f
C1710 vdd.n15 gnd 0.165864f
C1711 vdd.t235 gnd 0.01802f
C1712 vdd.t4 gnd 0.01802f
C1713 vdd.n16 gnd 0.165378f
C1714 vdd.n17 gnd 0.28781f
C1715 vdd.t234 gnd 0.01802f
C1716 vdd.t142 gnd 0.01802f
C1717 vdd.n18 gnd 0.165378f
C1718 vdd.n19 gnd 0.119071f
C1719 vdd.t117 gnd 0.01802f
C1720 vdd.t5 gnd 0.01802f
C1721 vdd.n20 gnd 0.165864f
C1722 vdd.t120 gnd 0.01802f
C1723 vdd.t231 gnd 0.01802f
C1724 vdd.n21 gnd 0.165378f
C1725 vdd.n22 gnd 0.28781f
C1726 vdd.t125 gnd 0.01802f
C1727 vdd.t116 gnd 0.01802f
C1728 vdd.n23 gnd 0.165378f
C1729 vdd.n24 gnd 0.119071f
C1730 vdd.t147 gnd 0.01802f
C1731 vdd.t230 gnd 0.01802f
C1732 vdd.n25 gnd 0.165378f
C1733 vdd.t152 gnd 0.01802f
C1734 vdd.t121 gnd 0.01802f
C1735 vdd.n26 gnd 0.165378f
C1736 vdd.n27 gnd 18.5015f
C1737 vdd.n28 gnd 7.436759f
C1738 vdd.n29 gnd 0.004915f
C1739 vdd.n30 gnd 0.004561f
C1740 vdd.n31 gnd 0.002523f
C1741 vdd.n32 gnd 0.005793f
C1742 vdd.n33 gnd 0.002451f
C1743 vdd.n34 gnd 0.002595f
C1744 vdd.n35 gnd 0.004561f
C1745 vdd.n36 gnd 0.002451f
C1746 vdd.n37 gnd 0.005793f
C1747 vdd.n38 gnd 0.002595f
C1748 vdd.n39 gnd 0.004561f
C1749 vdd.n40 gnd 0.002451f
C1750 vdd.n41 gnd 0.004344f
C1751 vdd.n42 gnd 0.004357f
C1752 vdd.t16 gnd 0.012445f
C1753 vdd.n43 gnd 0.027689f
C1754 vdd.n44 gnd 0.144102f
C1755 vdd.n45 gnd 0.002451f
C1756 vdd.n46 gnd 0.002595f
C1757 vdd.n47 gnd 0.005793f
C1758 vdd.n48 gnd 0.005793f
C1759 vdd.n49 gnd 0.002595f
C1760 vdd.n50 gnd 0.002451f
C1761 vdd.n51 gnd 0.004561f
C1762 vdd.n52 gnd 0.004561f
C1763 vdd.n53 gnd 0.002451f
C1764 vdd.n54 gnd 0.002595f
C1765 vdd.n55 gnd 0.005793f
C1766 vdd.n56 gnd 0.005793f
C1767 vdd.n57 gnd 0.002595f
C1768 vdd.n58 gnd 0.002451f
C1769 vdd.n59 gnd 0.004561f
C1770 vdd.n60 gnd 0.004561f
C1771 vdd.n61 gnd 0.002451f
C1772 vdd.n62 gnd 0.002595f
C1773 vdd.n63 gnd 0.005793f
C1774 vdd.n64 gnd 0.005793f
C1775 vdd.n65 gnd 0.013695f
C1776 vdd.n66 gnd 0.002523f
C1777 vdd.n67 gnd 0.002451f
C1778 vdd.n68 gnd 0.011788f
C1779 vdd.n69 gnd 0.00823f
C1780 vdd.t241 gnd 0.028831f
C1781 vdd.t217 gnd 0.028831f
C1782 vdd.n70 gnd 0.19815f
C1783 vdd.n71 gnd 0.155815f
C1784 vdd.t236 gnd 0.028831f
C1785 vdd.t223 gnd 0.028831f
C1786 vdd.n72 gnd 0.19815f
C1787 vdd.n73 gnd 0.125742f
C1788 vdd.t239 gnd 0.028831f
C1789 vdd.t149 gnd 0.028831f
C1790 vdd.n74 gnd 0.19815f
C1791 vdd.n75 gnd 0.125742f
C1792 vdd.t140 gnd 0.028831f
C1793 vdd.t129 gnd 0.028831f
C1794 vdd.n76 gnd 0.19815f
C1795 vdd.n77 gnd 0.125742f
C1796 vdd.t17 gnd 0.028831f
C1797 vdd.t232 gnd 0.028831f
C1798 vdd.n78 gnd 0.19815f
C1799 vdd.n79 gnd 0.125742f
C1800 vdd.n80 gnd 0.004915f
C1801 vdd.n81 gnd 0.004561f
C1802 vdd.n82 gnd 0.002523f
C1803 vdd.n83 gnd 0.005793f
C1804 vdd.n84 gnd 0.002451f
C1805 vdd.n85 gnd 0.002595f
C1806 vdd.n86 gnd 0.004561f
C1807 vdd.n87 gnd 0.002451f
C1808 vdd.n88 gnd 0.005793f
C1809 vdd.n89 gnd 0.002595f
C1810 vdd.n90 gnd 0.004561f
C1811 vdd.n91 gnd 0.002451f
C1812 vdd.n92 gnd 0.004344f
C1813 vdd.n93 gnd 0.004357f
C1814 vdd.t154 gnd 0.012445f
C1815 vdd.n94 gnd 0.027689f
C1816 vdd.n95 gnd 0.144102f
C1817 vdd.n96 gnd 0.002451f
C1818 vdd.n97 gnd 0.002595f
C1819 vdd.n98 gnd 0.005793f
C1820 vdd.n99 gnd 0.005793f
C1821 vdd.n100 gnd 0.002595f
C1822 vdd.n101 gnd 0.002451f
C1823 vdd.n102 gnd 0.004561f
C1824 vdd.n103 gnd 0.004561f
C1825 vdd.n104 gnd 0.002451f
C1826 vdd.n105 gnd 0.002595f
C1827 vdd.n106 gnd 0.005793f
C1828 vdd.n107 gnd 0.005793f
C1829 vdd.n108 gnd 0.002595f
C1830 vdd.n109 gnd 0.002451f
C1831 vdd.n110 gnd 0.004561f
C1832 vdd.n111 gnd 0.004561f
C1833 vdd.n112 gnd 0.002451f
C1834 vdd.n113 gnd 0.002595f
C1835 vdd.n114 gnd 0.005793f
C1836 vdd.n115 gnd 0.005793f
C1837 vdd.n116 gnd 0.013695f
C1838 vdd.n117 gnd 0.002523f
C1839 vdd.n118 gnd 0.002451f
C1840 vdd.n119 gnd 0.011788f
C1841 vdd.n120 gnd 0.007971f
C1842 vdd.n121 gnd 0.093552f
C1843 vdd.n122 gnd 0.004915f
C1844 vdd.n123 gnd 0.004561f
C1845 vdd.n124 gnd 0.002523f
C1846 vdd.n125 gnd 0.005793f
C1847 vdd.n126 gnd 0.002451f
C1848 vdd.n127 gnd 0.002595f
C1849 vdd.n128 gnd 0.004561f
C1850 vdd.n129 gnd 0.002451f
C1851 vdd.n130 gnd 0.005793f
C1852 vdd.n131 gnd 0.002595f
C1853 vdd.n132 gnd 0.004561f
C1854 vdd.n133 gnd 0.002451f
C1855 vdd.n134 gnd 0.004344f
C1856 vdd.n135 gnd 0.004357f
C1857 vdd.t219 gnd 0.012445f
C1858 vdd.n136 gnd 0.027689f
C1859 vdd.n137 gnd 0.144102f
C1860 vdd.n138 gnd 0.002451f
C1861 vdd.n139 gnd 0.002595f
C1862 vdd.n140 gnd 0.005793f
C1863 vdd.n141 gnd 0.005793f
C1864 vdd.n142 gnd 0.002595f
C1865 vdd.n143 gnd 0.002451f
C1866 vdd.n144 gnd 0.004561f
C1867 vdd.n145 gnd 0.004561f
C1868 vdd.n146 gnd 0.002451f
C1869 vdd.n147 gnd 0.002595f
C1870 vdd.n148 gnd 0.005793f
C1871 vdd.n149 gnd 0.005793f
C1872 vdd.n150 gnd 0.002595f
C1873 vdd.n151 gnd 0.002451f
C1874 vdd.n152 gnd 0.004561f
C1875 vdd.n153 gnd 0.004561f
C1876 vdd.n154 gnd 0.002451f
C1877 vdd.n155 gnd 0.002595f
C1878 vdd.n156 gnd 0.005793f
C1879 vdd.n157 gnd 0.005793f
C1880 vdd.n158 gnd 0.013695f
C1881 vdd.n159 gnd 0.002523f
C1882 vdd.n160 gnd 0.002451f
C1883 vdd.n161 gnd 0.011788f
C1884 vdd.n162 gnd 0.00823f
C1885 vdd.t218 gnd 0.028831f
C1886 vdd.t143 gnd 0.028831f
C1887 vdd.n163 gnd 0.19815f
C1888 vdd.n164 gnd 0.155815f
C1889 vdd.t104 gnd 0.028831f
C1890 vdd.t111 gnd 0.028831f
C1891 vdd.n165 gnd 0.19815f
C1892 vdd.n166 gnd 0.125742f
C1893 vdd.t134 gnd 0.028831f
C1894 vdd.t107 gnd 0.028831f
C1895 vdd.n167 gnd 0.19815f
C1896 vdd.n168 gnd 0.125742f
C1897 vdd.t233 gnd 0.028831f
C1898 vdd.t150 gnd 0.028831f
C1899 vdd.n169 gnd 0.19815f
C1900 vdd.n170 gnd 0.125742f
C1901 vdd.t13 gnd 0.028831f
C1902 vdd.t123 gnd 0.028831f
C1903 vdd.n171 gnd 0.19815f
C1904 vdd.n172 gnd 0.125742f
C1905 vdd.n173 gnd 0.004915f
C1906 vdd.n174 gnd 0.004561f
C1907 vdd.n175 gnd 0.002523f
C1908 vdd.n176 gnd 0.005793f
C1909 vdd.n177 gnd 0.002451f
C1910 vdd.n178 gnd 0.002595f
C1911 vdd.n179 gnd 0.004561f
C1912 vdd.n180 gnd 0.002451f
C1913 vdd.n181 gnd 0.005793f
C1914 vdd.n182 gnd 0.002595f
C1915 vdd.n183 gnd 0.004561f
C1916 vdd.n184 gnd 0.002451f
C1917 vdd.n185 gnd 0.004344f
C1918 vdd.n186 gnd 0.004357f
C1919 vdd.t23 gnd 0.012445f
C1920 vdd.n187 gnd 0.027689f
C1921 vdd.n188 gnd 0.144102f
C1922 vdd.n189 gnd 0.002451f
C1923 vdd.n190 gnd 0.002595f
C1924 vdd.n191 gnd 0.005793f
C1925 vdd.n192 gnd 0.005793f
C1926 vdd.n193 gnd 0.002595f
C1927 vdd.n194 gnd 0.002451f
C1928 vdd.n195 gnd 0.004561f
C1929 vdd.n196 gnd 0.004561f
C1930 vdd.n197 gnd 0.002451f
C1931 vdd.n198 gnd 0.002595f
C1932 vdd.n199 gnd 0.005793f
C1933 vdd.n200 gnd 0.005793f
C1934 vdd.n201 gnd 0.002595f
C1935 vdd.n202 gnd 0.002451f
C1936 vdd.n203 gnd 0.004561f
C1937 vdd.n204 gnd 0.004561f
C1938 vdd.n205 gnd 0.002451f
C1939 vdd.n206 gnd 0.002595f
C1940 vdd.n207 gnd 0.005793f
C1941 vdd.n208 gnd 0.005793f
C1942 vdd.n209 gnd 0.013695f
C1943 vdd.n210 gnd 0.002523f
C1944 vdd.n211 gnd 0.002451f
C1945 vdd.n212 gnd 0.011788f
C1946 vdd.n213 gnd 0.007971f
C1947 vdd.n214 gnd 0.055654f
C1948 vdd.n215 gnd 0.200537f
C1949 vdd.n216 gnd 0.004915f
C1950 vdd.n217 gnd 0.004561f
C1951 vdd.n218 gnd 0.002523f
C1952 vdd.n219 gnd 0.005793f
C1953 vdd.n220 gnd 0.002451f
C1954 vdd.n221 gnd 0.002595f
C1955 vdd.n222 gnd 0.004561f
C1956 vdd.n223 gnd 0.002451f
C1957 vdd.n224 gnd 0.005793f
C1958 vdd.n225 gnd 0.002595f
C1959 vdd.n226 gnd 0.004561f
C1960 vdd.n227 gnd 0.002451f
C1961 vdd.n228 gnd 0.004344f
C1962 vdd.n229 gnd 0.004357f
C1963 vdd.t3 gnd 0.012445f
C1964 vdd.n230 gnd 0.027689f
C1965 vdd.n231 gnd 0.144102f
C1966 vdd.n232 gnd 0.002451f
C1967 vdd.n233 gnd 0.002595f
C1968 vdd.n234 gnd 0.005793f
C1969 vdd.n235 gnd 0.005793f
C1970 vdd.n236 gnd 0.002595f
C1971 vdd.n237 gnd 0.002451f
C1972 vdd.n238 gnd 0.004561f
C1973 vdd.n239 gnd 0.004561f
C1974 vdd.n240 gnd 0.002451f
C1975 vdd.n241 gnd 0.002595f
C1976 vdd.n242 gnd 0.005793f
C1977 vdd.n243 gnd 0.005793f
C1978 vdd.n244 gnd 0.002595f
C1979 vdd.n245 gnd 0.002451f
C1980 vdd.n246 gnd 0.004561f
C1981 vdd.n247 gnd 0.004561f
C1982 vdd.n248 gnd 0.002451f
C1983 vdd.n249 gnd 0.002595f
C1984 vdd.n250 gnd 0.005793f
C1985 vdd.n251 gnd 0.005793f
C1986 vdd.n252 gnd 0.013695f
C1987 vdd.n253 gnd 0.002523f
C1988 vdd.n254 gnd 0.002451f
C1989 vdd.n255 gnd 0.011788f
C1990 vdd.n256 gnd 0.00823f
C1991 vdd.t1 gnd 0.028831f
C1992 vdd.t101 gnd 0.028831f
C1993 vdd.n257 gnd 0.19815f
C1994 vdd.n258 gnd 0.155815f
C1995 vdd.t112 gnd 0.028831f
C1996 vdd.t151 gnd 0.028831f
C1997 vdd.n259 gnd 0.19815f
C1998 vdd.n260 gnd 0.125742f
C1999 vdd.t238 gnd 0.028831f
C2000 vdd.t119 gnd 0.028831f
C2001 vdd.n261 gnd 0.19815f
C2002 vdd.n262 gnd 0.125742f
C2003 vdd.t148 gnd 0.028831f
C2004 vdd.t225 gnd 0.028831f
C2005 vdd.n263 gnd 0.19815f
C2006 vdd.n264 gnd 0.125742f
C2007 vdd.t130 gnd 0.028831f
C2008 vdd.t158 gnd 0.028831f
C2009 vdd.n265 gnd 0.19815f
C2010 vdd.n266 gnd 0.125742f
C2011 vdd.n267 gnd 0.004915f
C2012 vdd.n268 gnd 0.004561f
C2013 vdd.n269 gnd 0.002523f
C2014 vdd.n270 gnd 0.005793f
C2015 vdd.n271 gnd 0.002451f
C2016 vdd.n272 gnd 0.002595f
C2017 vdd.n273 gnd 0.004561f
C2018 vdd.n274 gnd 0.002451f
C2019 vdd.n275 gnd 0.005793f
C2020 vdd.n276 gnd 0.002595f
C2021 vdd.n277 gnd 0.004561f
C2022 vdd.n278 gnd 0.002451f
C2023 vdd.n279 gnd 0.004344f
C2024 vdd.n280 gnd 0.004357f
C2025 vdd.t144 gnd 0.012445f
C2026 vdd.n281 gnd 0.027689f
C2027 vdd.n282 gnd 0.144102f
C2028 vdd.n283 gnd 0.002451f
C2029 vdd.n284 gnd 0.002595f
C2030 vdd.n285 gnd 0.005793f
C2031 vdd.n286 gnd 0.005793f
C2032 vdd.n287 gnd 0.002595f
C2033 vdd.n288 gnd 0.002451f
C2034 vdd.n289 gnd 0.004561f
C2035 vdd.n290 gnd 0.004561f
C2036 vdd.n291 gnd 0.002451f
C2037 vdd.n292 gnd 0.002595f
C2038 vdd.n293 gnd 0.005793f
C2039 vdd.n294 gnd 0.005793f
C2040 vdd.n295 gnd 0.002595f
C2041 vdd.n296 gnd 0.002451f
C2042 vdd.n297 gnd 0.004561f
C2043 vdd.n298 gnd 0.004561f
C2044 vdd.n299 gnd 0.002451f
C2045 vdd.n300 gnd 0.002595f
C2046 vdd.n301 gnd 0.005793f
C2047 vdd.n302 gnd 0.005793f
C2048 vdd.n303 gnd 0.013695f
C2049 vdd.n304 gnd 0.002523f
C2050 vdd.n305 gnd 0.002451f
C2051 vdd.n306 gnd 0.011788f
C2052 vdd.n307 gnd 0.007971f
C2053 vdd.n308 gnd 0.055654f
C2054 vdd.n309 gnd 0.220396f
C2055 vdd.n310 gnd 0.008925f
C2056 vdd.n311 gnd 0.008925f
C2057 vdd.n312 gnd 0.007208f
C2058 vdd.n313 gnd 0.007208f
C2059 vdd.n314 gnd 0.008955f
C2060 vdd.n315 gnd 0.008955f
C2061 vdd.t133 gnd 0.457591f
C2062 vdd.n316 gnd 0.008955f
C2063 vdd.n317 gnd 0.008955f
C2064 vdd.n318 gnd 0.008955f
C2065 vdd.t139 gnd 0.457591f
C2066 vdd.n319 gnd 0.008955f
C2067 vdd.n320 gnd 0.008955f
C2068 vdd.n321 gnd 0.008955f
C2069 vdd.n322 gnd 0.008955f
C2070 vdd.n323 gnd 0.007208f
C2071 vdd.n324 gnd 0.008955f
C2072 vdd.n325 gnd 0.736722f
C2073 vdd.n326 gnd 0.008955f
C2074 vdd.n327 gnd 0.008955f
C2075 vdd.n328 gnd 0.008955f
C2076 vdd.n329 gnd 0.6269f
C2077 vdd.n330 gnd 0.008955f
C2078 vdd.n331 gnd 0.008955f
C2079 vdd.n332 gnd 0.008955f
C2080 vdd.n333 gnd 0.008955f
C2081 vdd.n334 gnd 0.008955f
C2082 vdd.n335 gnd 0.007208f
C2083 vdd.n336 gnd 0.008955f
C2084 vdd.t122 gnd 0.457591f
C2085 vdd.n337 gnd 0.008955f
C2086 vdd.n338 gnd 0.008955f
C2087 vdd.n339 gnd 0.008955f
C2088 vdd.n340 gnd 0.915183f
C2089 vdd.n341 gnd 0.008955f
C2090 vdd.n342 gnd 0.008955f
C2091 vdd.n343 gnd 0.008955f
C2092 vdd.n344 gnd 0.008955f
C2093 vdd.n345 gnd 0.008955f
C2094 vdd.n346 gnd 0.007208f
C2095 vdd.n347 gnd 0.008955f
C2096 vdd.n348 gnd 0.008955f
C2097 vdd.n349 gnd 0.008955f
C2098 vdd.n350 gnd 0.021104f
C2099 vdd.n351 gnd 2.10492f
C2100 vdd.n352 gnd 0.021434f
C2101 vdd.n353 gnd 0.008955f
C2102 vdd.n354 gnd 0.008955f
C2103 vdd.n356 gnd 0.008955f
C2104 vdd.n357 gnd 0.008955f
C2105 vdd.n358 gnd 0.007208f
C2106 vdd.n359 gnd 0.007208f
C2107 vdd.n360 gnd 0.008955f
C2108 vdd.n361 gnd 0.008955f
C2109 vdd.n362 gnd 0.008955f
C2110 vdd.n363 gnd 0.008955f
C2111 vdd.n364 gnd 0.008955f
C2112 vdd.n365 gnd 0.008955f
C2113 vdd.n366 gnd 0.007208f
C2114 vdd.n368 gnd 0.008955f
C2115 vdd.n369 gnd 0.008955f
C2116 vdd.n370 gnd 0.008955f
C2117 vdd.n371 gnd 0.008955f
C2118 vdd.n372 gnd 0.008955f
C2119 vdd.n373 gnd 0.007208f
C2120 vdd.n375 gnd 0.008955f
C2121 vdd.n376 gnd 0.008955f
C2122 vdd.n377 gnd 0.008955f
C2123 vdd.n378 gnd 0.008955f
C2124 vdd.n379 gnd 0.008955f
C2125 vdd.n380 gnd 0.007208f
C2126 vdd.n382 gnd 0.008955f
C2127 vdd.n383 gnd 0.008955f
C2128 vdd.n384 gnd 0.008955f
C2129 vdd.n385 gnd 0.008955f
C2130 vdd.n386 gnd 0.006019f
C2131 vdd.t66 gnd 0.110173f
C2132 vdd.t65 gnd 0.117745f
C2133 vdd.t64 gnd 0.143884f
C2134 vdd.n387 gnd 0.184439f
C2135 vdd.n388 gnd 0.155683f
C2136 vdd.n390 gnd 0.008955f
C2137 vdd.n391 gnd 0.008955f
C2138 vdd.n392 gnd 0.007208f
C2139 vdd.n393 gnd 0.008955f
C2140 vdd.n395 gnd 0.008955f
C2141 vdd.n396 gnd 0.008955f
C2142 vdd.n397 gnd 0.008955f
C2143 vdd.n398 gnd 0.008955f
C2144 vdd.n399 gnd 0.007208f
C2145 vdd.n401 gnd 0.008955f
C2146 vdd.n402 gnd 0.008955f
C2147 vdd.n403 gnd 0.008955f
C2148 vdd.n404 gnd 0.008955f
C2149 vdd.n405 gnd 0.008955f
C2150 vdd.n406 gnd 0.007208f
C2151 vdd.n408 gnd 0.008955f
C2152 vdd.n409 gnd 0.008955f
C2153 vdd.n410 gnd 0.008955f
C2154 vdd.n411 gnd 0.008955f
C2155 vdd.n412 gnd 0.008955f
C2156 vdd.n413 gnd 0.007208f
C2157 vdd.n415 gnd 0.008955f
C2158 vdd.n416 gnd 0.008955f
C2159 vdd.n417 gnd 0.008955f
C2160 vdd.n418 gnd 0.008955f
C2161 vdd.n419 gnd 0.008955f
C2162 vdd.n420 gnd 0.007208f
C2163 vdd.n422 gnd 0.008955f
C2164 vdd.n423 gnd 0.008955f
C2165 vdd.n424 gnd 0.008955f
C2166 vdd.n425 gnd 0.008955f
C2167 vdd.n426 gnd 0.007136f
C2168 vdd.t49 gnd 0.110173f
C2169 vdd.t48 gnd 0.117745f
C2170 vdd.t46 gnd 0.143884f
C2171 vdd.n427 gnd 0.184439f
C2172 vdd.n428 gnd 0.155683f
C2173 vdd.n430 gnd 0.008955f
C2174 vdd.n431 gnd 0.008955f
C2175 vdd.n432 gnd 0.007208f
C2176 vdd.n433 gnd 0.008955f
C2177 vdd.n435 gnd 0.008955f
C2178 vdd.n436 gnd 0.008955f
C2179 vdd.n437 gnd 0.008955f
C2180 vdd.n438 gnd 0.008955f
C2181 vdd.n439 gnd 0.007208f
C2182 vdd.n441 gnd 0.008955f
C2183 vdd.n442 gnd 0.008955f
C2184 vdd.n443 gnd 0.008955f
C2185 vdd.n444 gnd 0.008955f
C2186 vdd.n445 gnd 0.008955f
C2187 vdd.n446 gnd 0.007208f
C2188 vdd.n448 gnd 0.008955f
C2189 vdd.n449 gnd 0.008955f
C2190 vdd.n450 gnd 0.008955f
C2191 vdd.n451 gnd 0.008955f
C2192 vdd.n452 gnd 0.008955f
C2193 vdd.n453 gnd 0.007208f
C2194 vdd.n455 gnd 0.008955f
C2195 vdd.n456 gnd 0.008955f
C2196 vdd.n457 gnd 0.008955f
C2197 vdd.n458 gnd 0.008955f
C2198 vdd.n459 gnd 0.008955f
C2199 vdd.n460 gnd 0.007208f
C2200 vdd.n462 gnd 0.008955f
C2201 vdd.n463 gnd 0.008955f
C2202 vdd.n464 gnd 0.008955f
C2203 vdd.n465 gnd 0.008955f
C2204 vdd.n466 gnd 0.008955f
C2205 vdd.n467 gnd 0.008955f
C2206 vdd.n468 gnd 0.007208f
C2207 vdd.n469 gnd 0.008955f
C2208 vdd.n470 gnd 0.008955f
C2209 vdd.n471 gnd 0.007208f
C2210 vdd.n472 gnd 0.008955f
C2211 vdd.n473 gnd 0.008955f
C2212 vdd.n474 gnd 0.007208f
C2213 vdd.n475 gnd 0.008955f
C2214 vdd.n476 gnd 0.007208f
C2215 vdd.n477 gnd 0.008955f
C2216 vdd.n478 gnd 0.007208f
C2217 vdd.n479 gnd 0.008955f
C2218 vdd.n480 gnd 0.008955f
C2219 vdd.t110 gnd 0.457591f
C2220 vdd.n481 gnd 0.489623f
C2221 vdd.n482 gnd 0.008955f
C2222 vdd.n483 gnd 0.007208f
C2223 vdd.n484 gnd 0.008955f
C2224 vdd.n485 gnd 0.007208f
C2225 vdd.n486 gnd 0.008955f
C2226 vdd.t103 gnd 0.457591f
C2227 vdd.n487 gnd 0.008955f
C2228 vdd.n488 gnd 0.007208f
C2229 vdd.n489 gnd 0.008955f
C2230 vdd.n490 gnd 0.007208f
C2231 vdd.n491 gnd 0.008955f
C2232 vdd.n492 gnd 0.718418f
C2233 vdd.n493 gnd 0.759602f
C2234 vdd.t100 gnd 0.457591f
C2235 vdd.n494 gnd 0.008955f
C2236 vdd.n495 gnd 0.007208f
C2237 vdd.n496 gnd 0.008955f
C2238 vdd.n497 gnd 0.007208f
C2239 vdd.n498 gnd 0.008955f
C2240 vdd.n499 gnd 0.562837f
C2241 vdd.n500 gnd 0.008955f
C2242 vdd.n501 gnd 0.007208f
C2243 vdd.n502 gnd 0.008955f
C2244 vdd.n503 gnd 0.007208f
C2245 vdd.n504 gnd 0.008955f
C2246 vdd.n505 gnd 0.915183f
C2247 vdd.t2 gnd 0.457591f
C2248 vdd.n506 gnd 0.008955f
C2249 vdd.n507 gnd 0.007208f
C2250 vdd.n508 gnd 0.008955f
C2251 vdd.n509 gnd 0.007208f
C2252 vdd.n510 gnd 0.008955f
C2253 vdd.n511 gnd 0.489623f
C2254 vdd.n512 gnd 0.008955f
C2255 vdd.n513 gnd 0.007208f
C2256 vdd.n514 gnd 0.021434f
C2257 vdd.n515 gnd 0.021434f
C2258 vdd.n516 gnd 11.1103f
C2259 vdd.t43 gnd 0.457591f
C2260 vdd.n517 gnd 0.021434f
C2261 vdd.n518 gnd 0.007702f
C2262 vdd.n519 gnd 0.007208f
C2263 vdd.n524 gnd 0.005731f
C2264 vdd.n525 gnd 0.007208f
C2265 vdd.n526 gnd 0.008955f
C2266 vdd.n527 gnd 0.008955f
C2267 vdd.n528 gnd 0.008955f
C2268 vdd.n529 gnd 0.008955f
C2269 vdd.n530 gnd 0.008955f
C2270 vdd.n531 gnd 0.007208f
C2271 vdd.n532 gnd 0.008955f
C2272 vdd.n533 gnd 0.008955f
C2273 vdd.n534 gnd 0.008955f
C2274 vdd.n535 gnd 0.008955f
C2275 vdd.n536 gnd 0.008955f
C2276 vdd.n537 gnd 0.007208f
C2277 vdd.n538 gnd 0.008955f
C2278 vdd.n539 gnd 0.008955f
C2279 vdd.n540 gnd 0.008955f
C2280 vdd.n541 gnd 0.008955f
C2281 vdd.n542 gnd 0.008955f
C2282 vdd.t78 gnd 0.110173f
C2283 vdd.t79 gnd 0.117745f
C2284 vdd.t77 gnd 0.143884f
C2285 vdd.n543 gnd 0.184439f
C2286 vdd.n544 gnd 0.154963f
C2287 vdd.n545 gnd 0.014704f
C2288 vdd.n546 gnd 0.008955f
C2289 vdd.n547 gnd 0.008955f
C2290 vdd.n548 gnd 0.008955f
C2291 vdd.n549 gnd 0.008955f
C2292 vdd.n550 gnd 0.008955f
C2293 vdd.n551 gnd 0.007208f
C2294 vdd.n552 gnd 0.008955f
C2295 vdd.n553 gnd 0.008955f
C2296 vdd.n554 gnd 0.008955f
C2297 vdd.n555 gnd 0.008955f
C2298 vdd.n556 gnd 0.008955f
C2299 vdd.n557 gnd 0.007208f
C2300 vdd.n558 gnd 0.008955f
C2301 vdd.n559 gnd 0.008955f
C2302 vdd.n560 gnd 0.008955f
C2303 vdd.n561 gnd 0.008955f
C2304 vdd.n562 gnd 0.008955f
C2305 vdd.n563 gnd 0.007208f
C2306 vdd.n564 gnd 0.008955f
C2307 vdd.n565 gnd 0.008955f
C2308 vdd.n566 gnd 0.008955f
C2309 vdd.n567 gnd 0.008955f
C2310 vdd.n568 gnd 0.008955f
C2311 vdd.n569 gnd 0.007208f
C2312 vdd.n570 gnd 0.008955f
C2313 vdd.n571 gnd 0.008955f
C2314 vdd.n572 gnd 0.008955f
C2315 vdd.n573 gnd 0.008955f
C2316 vdd.n574 gnd 0.008955f
C2317 vdd.n575 gnd 0.007208f
C2318 vdd.n576 gnd 0.008955f
C2319 vdd.n577 gnd 0.008955f
C2320 vdd.n578 gnd 0.008955f
C2321 vdd.n579 gnd 0.007136f
C2322 vdd.t68 gnd 0.110173f
C2323 vdd.t69 gnd 0.117745f
C2324 vdd.t67 gnd 0.143884f
C2325 vdd.n580 gnd 0.184439f
C2326 vdd.n581 gnd 0.154963f
C2327 vdd.n582 gnd 0.008955f
C2328 vdd.n583 gnd 0.007208f
C2329 vdd.n585 gnd 0.008955f
C2330 vdd.n587 gnd 0.008955f
C2331 vdd.n588 gnd 0.008955f
C2332 vdd.n589 gnd 0.007208f
C2333 vdd.n590 gnd 0.008955f
C2334 vdd.n591 gnd 0.008955f
C2335 vdd.n592 gnd 0.008955f
C2336 vdd.n593 gnd 0.008955f
C2337 vdd.n594 gnd 0.008955f
C2338 vdd.n595 gnd 0.007208f
C2339 vdd.n596 gnd 0.008955f
C2340 vdd.n597 gnd 0.008955f
C2341 vdd.n598 gnd 0.008955f
C2342 vdd.n599 gnd 0.008955f
C2343 vdd.n600 gnd 0.008955f
C2344 vdd.n601 gnd 0.007208f
C2345 vdd.n602 gnd 0.008955f
C2346 vdd.n603 gnd 0.008955f
C2347 vdd.n604 gnd 0.008955f
C2348 vdd.n605 gnd 0.005731f
C2349 vdd.n610 gnd 0.00609f
C2350 vdd.n611 gnd 0.00609f
C2351 vdd.n612 gnd 0.00609f
C2352 vdd.n613 gnd 10.8083f
C2353 vdd.n614 gnd 0.00609f
C2354 vdd.n615 gnd 0.00609f
C2355 vdd.n616 gnd 0.00609f
C2356 vdd.n618 gnd 0.00609f
C2357 vdd.n619 gnd 0.00609f
C2358 vdd.n621 gnd 0.00609f
C2359 vdd.n622 gnd 0.004433f
C2360 vdd.n624 gnd 0.00609f
C2361 vdd.t27 gnd 0.246078f
C2362 vdd.t26 gnd 0.251892f
C2363 vdd.t24 gnd 0.160649f
C2364 vdd.n625 gnd 0.086822f
C2365 vdd.n626 gnd 0.049248f
C2366 vdd.n627 gnd 0.008703f
C2367 vdd.n628 gnd 0.013827f
C2368 vdd.n630 gnd 0.00609f
C2369 vdd.n631 gnd 0.622324f
C2370 vdd.n632 gnd 0.013039f
C2371 vdd.n633 gnd 0.013039f
C2372 vdd.n634 gnd 0.00609f
C2373 vdd.n635 gnd 0.013827f
C2374 vdd.n636 gnd 0.00609f
C2375 vdd.n637 gnd 0.00609f
C2376 vdd.n638 gnd 0.00609f
C2377 vdd.n639 gnd 0.00609f
C2378 vdd.n640 gnd 0.00609f
C2379 vdd.n642 gnd 0.00609f
C2380 vdd.n643 gnd 0.00609f
C2381 vdd.n645 gnd 0.00609f
C2382 vdd.n646 gnd 0.00609f
C2383 vdd.n648 gnd 0.00609f
C2384 vdd.n649 gnd 0.00609f
C2385 vdd.n651 gnd 0.00609f
C2386 vdd.n652 gnd 0.00609f
C2387 vdd.n654 gnd 0.00609f
C2388 vdd.n655 gnd 0.00609f
C2389 vdd.n657 gnd 0.00609f
C2390 vdd.n658 gnd 0.004433f
C2391 vdd.n660 gnd 0.00609f
C2392 vdd.t41 gnd 0.246078f
C2393 vdd.t40 gnd 0.251892f
C2394 vdd.t39 gnd 0.160649f
C2395 vdd.n661 gnd 0.086822f
C2396 vdd.n662 gnd 0.049248f
C2397 vdd.n663 gnd 0.008703f
C2398 vdd.n664 gnd 0.00609f
C2399 vdd.n665 gnd 0.00609f
C2400 vdd.t25 gnd 0.311162f
C2401 vdd.n666 gnd 0.00609f
C2402 vdd.n667 gnd 0.00609f
C2403 vdd.n668 gnd 0.00609f
C2404 vdd.n669 gnd 0.00609f
C2405 vdd.n670 gnd 0.00609f
C2406 vdd.n671 gnd 0.622324f
C2407 vdd.n672 gnd 0.00609f
C2408 vdd.n673 gnd 0.00609f
C2409 vdd.n674 gnd 0.489623f
C2410 vdd.n675 gnd 0.00609f
C2411 vdd.n676 gnd 0.00609f
C2412 vdd.n677 gnd 0.00609f
C2413 vdd.n678 gnd 0.00609f
C2414 vdd.n679 gnd 0.622324f
C2415 vdd.n680 gnd 0.00609f
C2416 vdd.n681 gnd 0.00609f
C2417 vdd.n682 gnd 0.00609f
C2418 vdd.n683 gnd 0.00609f
C2419 vdd.n684 gnd 0.00609f
C2420 vdd.t176 gnd 0.311162f
C2421 vdd.n685 gnd 0.00609f
C2422 vdd.n686 gnd 0.00609f
C2423 vdd.n687 gnd 0.00609f
C2424 vdd.n688 gnd 0.00609f
C2425 vdd.n689 gnd 0.00609f
C2426 vdd.t191 gnd 0.311162f
C2427 vdd.n690 gnd 0.00609f
C2428 vdd.n691 gnd 0.00609f
C2429 vdd.n692 gnd 0.599445f
C2430 vdd.n693 gnd 0.00609f
C2431 vdd.n694 gnd 0.00609f
C2432 vdd.n695 gnd 0.00609f
C2433 vdd.t190 gnd 0.311162f
C2434 vdd.n696 gnd 0.00609f
C2435 vdd.n697 gnd 0.00609f
C2436 vdd.n698 gnd 0.462167f
C2437 vdd.n699 gnd 0.00609f
C2438 vdd.n700 gnd 0.00609f
C2439 vdd.n701 gnd 0.00609f
C2440 vdd.n702 gnd 0.434712f
C2441 vdd.n703 gnd 0.00609f
C2442 vdd.n704 gnd 0.00609f
C2443 vdd.n705 gnd 0.32489f
C2444 vdd.n706 gnd 0.00609f
C2445 vdd.n707 gnd 0.00609f
C2446 vdd.n708 gnd 0.00609f
C2447 vdd.n709 gnd 0.571989f
C2448 vdd.n710 gnd 0.00609f
C2449 vdd.n711 gnd 0.00609f
C2450 vdd.t197 gnd 0.311162f
C2451 vdd.n712 gnd 0.00609f
C2452 vdd.n713 gnd 0.00609f
C2453 vdd.n714 gnd 0.00609f
C2454 vdd.n715 gnd 0.622324f
C2455 vdd.n716 gnd 0.00609f
C2456 vdd.n717 gnd 0.00609f
C2457 vdd.t198 gnd 0.311162f
C2458 vdd.n718 gnd 0.00609f
C2459 vdd.n719 gnd 0.00609f
C2460 vdd.n720 gnd 0.00609f
C2461 vdd.t170 gnd 0.311162f
C2462 vdd.n721 gnd 0.00609f
C2463 vdd.n722 gnd 0.00609f
C2464 vdd.n723 gnd 0.00609f
C2465 vdd.t52 gnd 0.251892f
C2466 vdd.t50 gnd 0.160649f
C2467 vdd.t53 gnd 0.251892f
C2468 vdd.n724 gnd 0.141573f
C2469 vdd.n725 gnd 0.017641f
C2470 vdd.n726 gnd 0.00609f
C2471 vdd.t51 gnd 0.22422f
C2472 vdd.n727 gnd 0.00609f
C2473 vdd.n728 gnd 0.00609f
C2474 vdd.n729 gnd 0.535382f
C2475 vdd.n730 gnd 0.00609f
C2476 vdd.n731 gnd 0.00609f
C2477 vdd.n732 gnd 0.00609f
C2478 vdd.n733 gnd 0.361497f
C2479 vdd.n734 gnd 0.00609f
C2480 vdd.n735 gnd 0.00609f
C2481 vdd.t171 gnd 0.128126f
C2482 vdd.n736 gnd 0.398104f
C2483 vdd.n737 gnd 0.00609f
C2484 vdd.n738 gnd 0.00609f
C2485 vdd.n739 gnd 0.00609f
C2486 vdd.n740 gnd 0.498775f
C2487 vdd.n741 gnd 0.00609f
C2488 vdd.n742 gnd 0.00609f
C2489 vdd.t182 gnd 0.311162f
C2490 vdd.n743 gnd 0.00609f
C2491 vdd.n744 gnd 0.00609f
C2492 vdd.n745 gnd 0.00609f
C2493 vdd.t178 gnd 0.311162f
C2494 vdd.n746 gnd 0.00609f
C2495 vdd.n747 gnd 0.00609f
C2496 vdd.t201 gnd 0.311162f
C2497 vdd.n748 gnd 0.00609f
C2498 vdd.n749 gnd 0.00609f
C2499 vdd.n750 gnd 0.00609f
C2500 vdd.t160 gnd 0.210492f
C2501 vdd.n751 gnd 0.00609f
C2502 vdd.n752 gnd 0.00609f
C2503 vdd.n753 gnd 0.54911f
C2504 vdd.n754 gnd 0.00609f
C2505 vdd.n755 gnd 0.00609f
C2506 vdd.n756 gnd 0.00609f
C2507 vdd.t202 gnd 0.311162f
C2508 vdd.n757 gnd 0.00609f
C2509 vdd.n758 gnd 0.00609f
C2510 vdd.t214 gnd 0.297434f
C2511 vdd.n759 gnd 0.411832f
C2512 vdd.n760 gnd 0.00609f
C2513 vdd.n761 gnd 0.00609f
C2514 vdd.n762 gnd 0.00609f
C2515 vdd.t166 gnd 0.311162f
C2516 vdd.n763 gnd 0.00609f
C2517 vdd.n764 gnd 0.00609f
C2518 vdd.t206 gnd 0.311162f
C2519 vdd.n765 gnd 0.00609f
C2520 vdd.n766 gnd 0.00609f
C2521 vdd.n767 gnd 0.00609f
C2522 vdd.n768 gnd 0.622324f
C2523 vdd.n769 gnd 0.00609f
C2524 vdd.n770 gnd 0.00609f
C2525 vdd.t186 gnd 0.311162f
C2526 vdd.n771 gnd 0.00609f
C2527 vdd.n772 gnd 0.00609f
C2528 vdd.n773 gnd 0.00609f
C2529 vdd.n774 gnd 0.430136f
C2530 vdd.n775 gnd 0.00609f
C2531 vdd.n776 gnd 0.00609f
C2532 vdd.n777 gnd 0.00609f
C2533 vdd.n778 gnd 0.00609f
C2534 vdd.n779 gnd 0.00609f
C2535 vdd.t81 gnd 0.311162f
C2536 vdd.n780 gnd 0.00609f
C2537 vdd.n781 gnd 0.00609f
C2538 vdd.t168 gnd 0.311162f
C2539 vdd.n782 gnd 0.00609f
C2540 vdd.n783 gnd 0.013039f
C2541 vdd.n784 gnd 0.013039f
C2542 vdd.n785 gnd 0.704691f
C2543 vdd.n786 gnd 0.00609f
C2544 vdd.n787 gnd 0.00609f
C2545 vdd.t195 gnd 0.311162f
C2546 vdd.n788 gnd 0.013039f
C2547 vdd.n789 gnd 0.00609f
C2548 vdd.n790 gnd 0.00609f
C2549 vdd.t208 gnd 0.530806f
C2550 vdd.n808 gnd 0.013827f
C2551 vdd.n826 gnd 0.013039f
C2552 vdd.n827 gnd 0.00609f
C2553 vdd.n828 gnd 0.013039f
C2554 vdd.t99 gnd 0.246078f
C2555 vdd.t98 gnd 0.251892f
C2556 vdd.t97 gnd 0.160649f
C2557 vdd.n829 gnd 0.086822f
C2558 vdd.n830 gnd 0.049248f
C2559 vdd.n831 gnd 0.013827f
C2560 vdd.n832 gnd 0.00609f
C2561 vdd.n833 gnd 0.366073f
C2562 vdd.n834 gnd 0.013039f
C2563 vdd.n835 gnd 0.00609f
C2564 vdd.n836 gnd 0.013827f
C2565 vdd.n837 gnd 0.00609f
C2566 vdd.t76 gnd 0.246078f
C2567 vdd.t75 gnd 0.251892f
C2568 vdd.t73 gnd 0.160649f
C2569 vdd.n838 gnd 0.086822f
C2570 vdd.n839 gnd 0.049248f
C2571 vdd.n840 gnd 0.008703f
C2572 vdd.n841 gnd 0.00609f
C2573 vdd.n842 gnd 0.00609f
C2574 vdd.t74 gnd 0.311162f
C2575 vdd.n843 gnd 0.00609f
C2576 vdd.t210 gnd 0.311162f
C2577 vdd.n844 gnd 0.00609f
C2578 vdd.n845 gnd 0.00609f
C2579 vdd.n846 gnd 0.00609f
C2580 vdd.n847 gnd 0.00609f
C2581 vdd.n848 gnd 0.00609f
C2582 vdd.n849 gnd 0.622324f
C2583 vdd.n850 gnd 0.00609f
C2584 vdd.n851 gnd 0.00609f
C2585 vdd.t180 gnd 0.311162f
C2586 vdd.n852 gnd 0.00609f
C2587 vdd.n853 gnd 0.00609f
C2588 vdd.n854 gnd 0.00609f
C2589 vdd.n855 gnd 0.00609f
C2590 vdd.n856 gnd 0.448439f
C2591 vdd.n857 gnd 0.00609f
C2592 vdd.n858 gnd 0.00609f
C2593 vdd.n859 gnd 0.00609f
C2594 vdd.n860 gnd 0.00609f
C2595 vdd.n861 gnd 0.00609f
C2596 vdd.t161 gnd 0.311162f
C2597 vdd.n862 gnd 0.00609f
C2598 vdd.n863 gnd 0.00609f
C2599 vdd.t199 gnd 0.311162f
C2600 vdd.n864 gnd 0.00609f
C2601 vdd.n865 gnd 0.00609f
C2602 vdd.n866 gnd 0.00609f
C2603 vdd.t185 gnd 0.311162f
C2604 vdd.n867 gnd 0.00609f
C2605 vdd.n868 gnd 0.00609f
C2606 vdd.t162 gnd 0.311162f
C2607 vdd.n869 gnd 0.00609f
C2608 vdd.n870 gnd 0.00609f
C2609 vdd.n871 gnd 0.00609f
C2610 vdd.t183 gnd 0.297434f
C2611 vdd.n872 gnd 0.00609f
C2612 vdd.n873 gnd 0.00609f
C2613 vdd.n874 gnd 0.462167f
C2614 vdd.n875 gnd 0.00609f
C2615 vdd.n876 gnd 0.00609f
C2616 vdd.n877 gnd 0.00609f
C2617 vdd.t203 gnd 0.311162f
C2618 vdd.n878 gnd 0.00609f
C2619 vdd.n879 gnd 0.00609f
C2620 vdd.t173 gnd 0.210492f
C2621 vdd.n880 gnd 0.32489f
C2622 vdd.n881 gnd 0.00609f
C2623 vdd.n882 gnd 0.00609f
C2624 vdd.n883 gnd 0.00609f
C2625 vdd.n884 gnd 0.571989f
C2626 vdd.n885 gnd 0.00609f
C2627 vdd.n886 gnd 0.00609f
C2628 vdd.t212 gnd 0.311162f
C2629 vdd.n887 gnd 0.00609f
C2630 vdd.n888 gnd 0.00609f
C2631 vdd.n889 gnd 0.00609f
C2632 vdd.n890 gnd 0.622324f
C2633 vdd.n891 gnd 0.00609f
C2634 vdd.n892 gnd 0.00609f
C2635 vdd.t177 gnd 0.311162f
C2636 vdd.n893 gnd 0.00609f
C2637 vdd.n894 gnd 0.00609f
C2638 vdd.n895 gnd 0.00609f
C2639 vdd.t172 gnd 0.128126f
C2640 vdd.n896 gnd 0.00609f
C2641 vdd.n897 gnd 0.00609f
C2642 vdd.n898 gnd 0.00609f
C2643 vdd.t89 gnd 0.251892f
C2644 vdd.t87 gnd 0.160649f
C2645 vdd.t90 gnd 0.251892f
C2646 vdd.n899 gnd 0.141573f
C2647 vdd.n900 gnd 0.00609f
C2648 vdd.n901 gnd 0.00609f
C2649 vdd.t192 gnd 0.311162f
C2650 vdd.n902 gnd 0.00609f
C2651 vdd.n903 gnd 0.00609f
C2652 vdd.t88 gnd 0.22422f
C2653 vdd.n904 gnd 0.494199f
C2654 vdd.n905 gnd 0.00609f
C2655 vdd.n906 gnd 0.00609f
C2656 vdd.n907 gnd 0.00609f
C2657 vdd.n908 gnd 0.361497f
C2658 vdd.n909 gnd 0.00609f
C2659 vdd.n910 gnd 0.00609f
C2660 vdd.n911 gnd 0.398104f
C2661 vdd.n912 gnd 0.00609f
C2662 vdd.n913 gnd 0.00609f
C2663 vdd.n914 gnd 0.00609f
C2664 vdd.n915 gnd 0.498775f
C2665 vdd.n916 gnd 0.00609f
C2666 vdd.n917 gnd 0.00609f
C2667 vdd.t174 gnd 0.311162f
C2668 vdd.n918 gnd 0.00609f
C2669 vdd.n919 gnd 0.00609f
C2670 vdd.n920 gnd 0.00609f
C2671 vdd.n921 gnd 0.622324f
C2672 vdd.n922 gnd 0.00609f
C2673 vdd.n923 gnd 0.00609f
C2674 vdd.t175 gnd 0.311162f
C2675 vdd.n924 gnd 0.00609f
C2676 vdd.n925 gnd 0.00609f
C2677 vdd.n926 gnd 0.00609f
C2678 vdd.t213 gnd 0.311162f
C2679 vdd.n927 gnd 0.00609f
C2680 vdd.n928 gnd 0.00609f
C2681 vdd.n929 gnd 0.00609f
C2682 vdd.n930 gnd 0.00609f
C2683 vdd.n931 gnd 0.00609f
C2684 vdd.t205 gnd 0.311162f
C2685 vdd.n932 gnd 0.00609f
C2686 vdd.n933 gnd 0.00609f
C2687 vdd.n934 gnd 0.608596f
C2688 vdd.n935 gnd 0.00609f
C2689 vdd.n936 gnd 0.00609f
C2690 vdd.n937 gnd 0.00609f
C2691 vdd.t167 gnd 0.311162f
C2692 vdd.n938 gnd 0.00609f
C2693 vdd.n939 gnd 0.00609f
C2694 vdd.n940 gnd 0.471319f
C2695 vdd.n941 gnd 0.00609f
C2696 vdd.n942 gnd 0.00609f
C2697 vdd.n943 gnd 0.00609f
C2698 vdd.n944 gnd 0.622324f
C2699 vdd.n945 gnd 0.00609f
C2700 vdd.n946 gnd 0.00609f
C2701 vdd.n947 gnd 0.334042f
C2702 vdd.n948 gnd 0.00609f
C2703 vdd.n949 gnd 0.00609f
C2704 vdd.n950 gnd 0.00609f
C2705 vdd.n951 gnd 0.622324f
C2706 vdd.n952 gnd 0.00609f
C2707 vdd.n953 gnd 0.00609f
C2708 vdd.n954 gnd 0.00609f
C2709 vdd.n955 gnd 0.00609f
C2710 vdd.n956 gnd 0.00609f
C2711 vdd.t29 gnd 0.311162f
C2712 vdd.n957 gnd 0.00609f
C2713 vdd.n958 gnd 0.00609f
C2714 vdd.n959 gnd 0.00609f
C2715 vdd.n960 gnd 0.013039f
C2716 vdd.n961 gnd 0.013039f
C2717 vdd.n962 gnd 0.841968f
C2718 vdd.n963 gnd 0.00609f
C2719 vdd.n964 gnd 0.00609f
C2720 vdd.n965 gnd 0.443864f
C2721 vdd.n966 gnd 0.013039f
C2722 vdd.n967 gnd 0.00609f
C2723 vdd.n968 gnd 0.00609f
C2724 vdd.n969 gnd 11.1103f
C2725 vdd.n1003 gnd 0.013827f
C2726 vdd.n1004 gnd 0.00609f
C2727 vdd.n1005 gnd 0.00609f
C2728 vdd.n1006 gnd 0.005731f
C2729 vdd.n1009 gnd 0.021434f
C2730 vdd.n1010 gnd 0.005983f
C2731 vdd.n1011 gnd 0.007208f
C2732 vdd.n1013 gnd 0.008955f
C2733 vdd.n1014 gnd 0.008955f
C2734 vdd.n1015 gnd 0.007208f
C2735 vdd.n1017 gnd 0.008955f
C2736 vdd.n1018 gnd 0.008955f
C2737 vdd.n1019 gnd 0.008955f
C2738 vdd.n1020 gnd 0.008955f
C2739 vdd.n1021 gnd 0.008955f
C2740 vdd.n1022 gnd 0.007208f
C2741 vdd.n1024 gnd 0.008955f
C2742 vdd.n1025 gnd 0.008955f
C2743 vdd.n1026 gnd 0.008955f
C2744 vdd.n1027 gnd 0.008955f
C2745 vdd.n1028 gnd 0.008955f
C2746 vdd.n1029 gnd 0.007208f
C2747 vdd.n1031 gnd 0.008955f
C2748 vdd.n1032 gnd 0.008955f
C2749 vdd.n1033 gnd 0.008955f
C2750 vdd.n1034 gnd 0.008955f
C2751 vdd.n1035 gnd 0.006019f
C2752 vdd.t38 gnd 0.110173f
C2753 vdd.t37 gnd 0.117745f
C2754 vdd.t36 gnd 0.143884f
C2755 vdd.n1036 gnd 0.184439f
C2756 vdd.n1037 gnd 0.154963f
C2757 vdd.n1039 gnd 0.008955f
C2758 vdd.n1040 gnd 0.008955f
C2759 vdd.n1041 gnd 0.007208f
C2760 vdd.n1042 gnd 0.008955f
C2761 vdd.n1044 gnd 0.008955f
C2762 vdd.n1045 gnd 0.008955f
C2763 vdd.n1046 gnd 0.008955f
C2764 vdd.n1047 gnd 0.008955f
C2765 vdd.n1048 gnd 0.007208f
C2766 vdd.n1050 gnd 0.008955f
C2767 vdd.n1051 gnd 0.008955f
C2768 vdd.n1052 gnd 0.008955f
C2769 vdd.n1053 gnd 0.008955f
C2770 vdd.n1054 gnd 0.008955f
C2771 vdd.n1055 gnd 0.007208f
C2772 vdd.n1057 gnd 0.008955f
C2773 vdd.n1058 gnd 0.008955f
C2774 vdd.n1059 gnd 0.008955f
C2775 vdd.n1060 gnd 0.008955f
C2776 vdd.n1061 gnd 0.008955f
C2777 vdd.n1062 gnd 0.007208f
C2778 vdd.n1064 gnd 0.008955f
C2779 vdd.n1065 gnd 0.008955f
C2780 vdd.n1066 gnd 0.008955f
C2781 vdd.n1067 gnd 0.008955f
C2782 vdd.n1068 gnd 0.008955f
C2783 vdd.n1069 gnd 0.007208f
C2784 vdd.n1071 gnd 0.008955f
C2785 vdd.n1072 gnd 0.008955f
C2786 vdd.n1073 gnd 0.008955f
C2787 vdd.n1074 gnd 0.008955f
C2788 vdd.n1075 gnd 0.007136f
C2789 vdd.t35 gnd 0.110173f
C2790 vdd.t34 gnd 0.117745f
C2791 vdd.t32 gnd 0.143884f
C2792 vdd.n1076 gnd 0.184439f
C2793 vdd.n1077 gnd 0.154963f
C2794 vdd.n1079 gnd 0.008955f
C2795 vdd.n1080 gnd 0.008955f
C2796 vdd.n1081 gnd 0.007208f
C2797 vdd.n1082 gnd 0.008955f
C2798 vdd.n1084 gnd 0.008955f
C2799 vdd.n1085 gnd 0.008955f
C2800 vdd.n1086 gnd 0.008955f
C2801 vdd.n1087 gnd 0.008955f
C2802 vdd.n1088 gnd 0.007208f
C2803 vdd.n1090 gnd 0.008955f
C2804 vdd.n1091 gnd 0.008955f
C2805 vdd.n1092 gnd 0.008955f
C2806 vdd.n1093 gnd 0.008955f
C2807 vdd.n1094 gnd 0.008955f
C2808 vdd.n1095 gnd 0.007208f
C2809 vdd.n1097 gnd 0.008955f
C2810 vdd.n1098 gnd 0.008955f
C2811 vdd.n1099 gnd 0.008955f
C2812 vdd.n1100 gnd 0.008955f
C2813 vdd.n1101 gnd 0.008955f
C2814 vdd.n1102 gnd 0.007208f
C2815 vdd.n1104 gnd 0.008955f
C2816 vdd.n1105 gnd 0.008955f
C2817 vdd.n1106 gnd 0.005731f
C2818 vdd.n1107 gnd 0.007208f
C2819 vdd.n1108 gnd 0.013827f
C2820 vdd.n1109 gnd 0.013827f
C2821 vdd.n1110 gnd 0.00609f
C2822 vdd.n1111 gnd 0.00609f
C2823 vdd.n1112 gnd 0.00609f
C2824 vdd.n1113 gnd 0.00609f
C2825 vdd.n1114 gnd 0.00609f
C2826 vdd.n1115 gnd 0.00609f
C2827 vdd.n1116 gnd 0.00609f
C2828 vdd.n1117 gnd 0.00609f
C2829 vdd.n1118 gnd 0.00609f
C2830 vdd.n1119 gnd 0.00609f
C2831 vdd.n1120 gnd 0.00609f
C2832 vdd.n1121 gnd 0.00609f
C2833 vdd.n1122 gnd 0.00609f
C2834 vdd.n1123 gnd 0.00609f
C2835 vdd.n1124 gnd 0.00609f
C2836 vdd.n1125 gnd 0.00609f
C2837 vdd.n1126 gnd 0.00609f
C2838 vdd.n1127 gnd 0.00609f
C2839 vdd.n1128 gnd 0.00609f
C2840 vdd.n1129 gnd 0.00609f
C2841 vdd.n1130 gnd 0.00609f
C2842 vdd.n1131 gnd 0.00609f
C2843 vdd.n1132 gnd 0.00609f
C2844 vdd.n1133 gnd 0.00609f
C2845 vdd.n1134 gnd 0.00609f
C2846 vdd.n1135 gnd 0.00609f
C2847 vdd.n1136 gnd 0.00609f
C2848 vdd.n1137 gnd 0.00609f
C2849 vdd.n1138 gnd 0.00609f
C2850 vdd.n1139 gnd 0.00609f
C2851 vdd.n1140 gnd 0.00609f
C2852 vdd.n1141 gnd 0.00609f
C2853 vdd.n1142 gnd 0.00609f
C2854 vdd.t30 gnd 0.246078f
C2855 vdd.t31 gnd 0.251892f
C2856 vdd.t28 gnd 0.160649f
C2857 vdd.n1143 gnd 0.086822f
C2858 vdd.n1144 gnd 0.049248f
C2859 vdd.n1145 gnd 0.008703f
C2860 vdd.n1146 gnd 0.00609f
C2861 vdd.t71 gnd 0.246078f
C2862 vdd.t72 gnd 0.251892f
C2863 vdd.t70 gnd 0.160649f
C2864 vdd.n1147 gnd 0.086822f
C2865 vdd.n1148 gnd 0.049248f
C2866 vdd.n1149 gnd 0.00609f
C2867 vdd.n1150 gnd 0.00609f
C2868 vdd.n1151 gnd 0.00609f
C2869 vdd.n1152 gnd 0.00609f
C2870 vdd.n1153 gnd 0.00609f
C2871 vdd.n1154 gnd 0.00609f
C2872 vdd.n1155 gnd 0.00609f
C2873 vdd.n1156 gnd 0.00609f
C2874 vdd.n1157 gnd 0.00609f
C2875 vdd.n1158 gnd 0.00609f
C2876 vdd.n1159 gnd 0.00609f
C2877 vdd.n1160 gnd 0.00609f
C2878 vdd.n1161 gnd 0.00609f
C2879 vdd.n1162 gnd 0.00609f
C2880 vdd.n1163 gnd 0.00609f
C2881 vdd.n1164 gnd 0.00609f
C2882 vdd.n1165 gnd 0.00609f
C2883 vdd.n1166 gnd 0.00609f
C2884 vdd.n1167 gnd 0.00609f
C2885 vdd.n1168 gnd 0.00609f
C2886 vdd.n1169 gnd 0.00609f
C2887 vdd.n1170 gnd 0.00609f
C2888 vdd.n1171 gnd 0.00609f
C2889 vdd.n1172 gnd 0.00609f
C2890 vdd.n1173 gnd 0.00609f
C2891 vdd.n1174 gnd 0.00609f
C2892 vdd.n1175 gnd 0.004433f
C2893 vdd.n1176 gnd 0.008703f
C2894 vdd.n1177 gnd 0.004701f
C2895 vdd.n1178 gnd 0.00609f
C2896 vdd.n1179 gnd 0.00609f
C2897 vdd.n1180 gnd 0.00609f
C2898 vdd.n1181 gnd 0.013827f
C2899 vdd.n1182 gnd 0.013827f
C2900 vdd.n1183 gnd 0.013039f
C2901 vdd.n1184 gnd 0.013039f
C2902 vdd.n1185 gnd 0.00609f
C2903 vdd.n1186 gnd 0.00609f
C2904 vdd.n1187 gnd 0.00609f
C2905 vdd.n1188 gnd 0.00609f
C2906 vdd.n1189 gnd 0.00609f
C2907 vdd.n1190 gnd 0.00609f
C2908 vdd.n1191 gnd 0.00609f
C2909 vdd.n1192 gnd 0.00609f
C2910 vdd.n1193 gnd 0.00609f
C2911 vdd.n1194 gnd 0.00609f
C2912 vdd.n1195 gnd 0.00609f
C2913 vdd.n1196 gnd 0.00609f
C2914 vdd.n1197 gnd 0.00609f
C2915 vdd.n1198 gnd 0.00609f
C2916 vdd.n1199 gnd 0.00609f
C2917 vdd.n1200 gnd 0.00609f
C2918 vdd.n1201 gnd 0.00609f
C2919 vdd.n1202 gnd 0.00609f
C2920 vdd.n1203 gnd 0.00609f
C2921 vdd.n1204 gnd 0.00609f
C2922 vdd.n1205 gnd 0.00609f
C2923 vdd.n1206 gnd 0.00609f
C2924 vdd.n1207 gnd 0.00609f
C2925 vdd.n1208 gnd 0.00609f
C2926 vdd.n1209 gnd 0.00609f
C2927 vdd.n1210 gnd 0.00609f
C2928 vdd.n1211 gnd 0.00609f
C2929 vdd.n1212 gnd 0.00609f
C2930 vdd.n1213 gnd 0.00609f
C2931 vdd.n1214 gnd 0.00609f
C2932 vdd.n1215 gnd 0.00609f
C2933 vdd.n1216 gnd 0.00609f
C2934 vdd.n1217 gnd 0.00609f
C2935 vdd.n1218 gnd 0.00609f
C2936 vdd.n1219 gnd 0.00609f
C2937 vdd.n1220 gnd 0.00609f
C2938 vdd.n1221 gnd 0.00609f
C2939 vdd.n1222 gnd 0.00609f
C2940 vdd.n1223 gnd 0.00609f
C2941 vdd.n1224 gnd 0.00609f
C2942 vdd.n1225 gnd 0.00609f
C2943 vdd.n1226 gnd 0.00609f
C2944 vdd.n1227 gnd 0.370649f
C2945 vdd.n1228 gnd 0.00609f
C2946 vdd.n1229 gnd 0.00609f
C2947 vdd.n1230 gnd 0.00609f
C2948 vdd.n1231 gnd 0.00609f
C2949 vdd.n1232 gnd 0.00609f
C2950 vdd.n1233 gnd 0.00609f
C2951 vdd.n1234 gnd 0.00609f
C2952 vdd.n1235 gnd 0.00609f
C2953 vdd.n1236 gnd 0.00609f
C2954 vdd.n1237 gnd 0.00609f
C2955 vdd.n1238 gnd 0.00609f
C2956 vdd.n1239 gnd 0.00609f
C2957 vdd.n1240 gnd 0.00609f
C2958 vdd.n1241 gnd 0.00609f
C2959 vdd.n1242 gnd 0.00609f
C2960 vdd.n1243 gnd 0.00609f
C2961 vdd.n1244 gnd 0.00609f
C2962 vdd.n1245 gnd 0.00609f
C2963 vdd.n1246 gnd 0.00609f
C2964 vdd.n1247 gnd 0.00609f
C2965 vdd.n1248 gnd 0.00609f
C2966 vdd.n1249 gnd 0.00609f
C2967 vdd.n1250 gnd 0.00609f
C2968 vdd.n1251 gnd 0.00609f
C2969 vdd.n1252 gnd 0.00609f
C2970 vdd.n1253 gnd 0.562837f
C2971 vdd.n1254 gnd 0.00609f
C2972 vdd.n1255 gnd 0.00609f
C2973 vdd.n1256 gnd 0.00609f
C2974 vdd.n1257 gnd 0.00609f
C2975 vdd.n1258 gnd 0.00609f
C2976 vdd.n1259 gnd 0.00609f
C2977 vdd.n1260 gnd 0.00609f
C2978 vdd.n1261 gnd 0.00609f
C2979 vdd.n1262 gnd 0.00609f
C2980 vdd.n1263 gnd 0.00609f
C2981 vdd.n1264 gnd 0.00609f
C2982 vdd.n1265 gnd 0.196764f
C2983 vdd.n1266 gnd 0.00609f
C2984 vdd.n1267 gnd 0.00609f
C2985 vdd.n1268 gnd 0.00609f
C2986 vdd.n1269 gnd 0.00609f
C2987 vdd.n1270 gnd 0.00609f
C2988 vdd.n1271 gnd 0.00609f
C2989 vdd.n1272 gnd 0.00609f
C2990 vdd.n1273 gnd 0.00609f
C2991 vdd.n1274 gnd 0.00609f
C2992 vdd.n1275 gnd 0.00609f
C2993 vdd.n1276 gnd 0.00609f
C2994 vdd.n1277 gnd 0.00609f
C2995 vdd.n1278 gnd 0.00609f
C2996 vdd.n1279 gnd 0.00609f
C2997 vdd.n1280 gnd 0.00609f
C2998 vdd.n1281 gnd 0.00609f
C2999 vdd.n1282 gnd 0.00609f
C3000 vdd.n1283 gnd 0.00609f
C3001 vdd.n1284 gnd 0.00609f
C3002 vdd.n1285 gnd 0.00609f
C3003 vdd.n1286 gnd 0.00609f
C3004 vdd.n1287 gnd 0.00609f
C3005 vdd.n1288 gnd 0.00609f
C3006 vdd.n1289 gnd 0.00609f
C3007 vdd.n1290 gnd 0.00609f
C3008 vdd.n1291 gnd 0.00609f
C3009 vdd.n1292 gnd 0.00609f
C3010 vdd.n1293 gnd 0.00609f
C3011 vdd.n1294 gnd 0.00609f
C3012 vdd.n1295 gnd 0.00609f
C3013 vdd.n1296 gnd 0.00609f
C3014 vdd.n1297 gnd 0.00609f
C3015 vdd.n1298 gnd 0.00609f
C3016 vdd.n1299 gnd 0.00609f
C3017 vdd.n1300 gnd 0.00609f
C3018 vdd.n1301 gnd 0.00609f
C3019 vdd.n1302 gnd 0.00609f
C3020 vdd.n1303 gnd 0.00609f
C3021 vdd.n1304 gnd 0.00609f
C3022 vdd.n1305 gnd 0.00609f
C3023 vdd.n1306 gnd 0.00609f
C3024 vdd.n1307 gnd 0.00609f
C3025 vdd.n1308 gnd 0.013039f
C3026 vdd.n1309 gnd 0.013039f
C3027 vdd.n1310 gnd 0.013827f
C3028 vdd.n1311 gnd 0.00609f
C3029 vdd.n1312 gnd 0.00609f
C3030 vdd.n1313 gnd 0.004701f
C3031 vdd.n1314 gnd 0.00609f
C3032 vdd.n1315 gnd 0.00609f
C3033 vdd.n1316 gnd 0.004433f
C3034 vdd.n1317 gnd 0.00609f
C3035 vdd.n1318 gnd 0.00609f
C3036 vdd.n1319 gnd 0.00609f
C3037 vdd.n1320 gnd 0.00609f
C3038 vdd.n1321 gnd 0.00609f
C3039 vdd.n1322 gnd 0.00609f
C3040 vdd.n1323 gnd 0.00609f
C3041 vdd.n1324 gnd 0.00609f
C3042 vdd.n1325 gnd 0.00609f
C3043 vdd.n1326 gnd 0.00609f
C3044 vdd.n1327 gnd 0.00609f
C3045 vdd.n1328 gnd 0.00609f
C3046 vdd.n1329 gnd 0.00609f
C3047 vdd.n1330 gnd 0.00609f
C3048 vdd.n1331 gnd 0.00609f
C3049 vdd.n1332 gnd 0.00609f
C3050 vdd.n1333 gnd 0.00609f
C3051 vdd.n1334 gnd 0.00609f
C3052 vdd.n1335 gnd 0.00609f
C3053 vdd.n1336 gnd 0.00609f
C3054 vdd.n1337 gnd 0.00609f
C3055 vdd.n1338 gnd 0.00609f
C3056 vdd.n1339 gnd 0.00609f
C3057 vdd.n1340 gnd 0.00609f
C3058 vdd.n1341 gnd 0.00609f
C3059 vdd.n1342 gnd 0.00609f
C3060 vdd.n1343 gnd 0.041023f
C3061 vdd.n1345 gnd 0.021434f
C3062 vdd.n1346 gnd 0.007208f
C3063 vdd.n1348 gnd 0.008955f
C3064 vdd.n1349 gnd 0.007208f
C3065 vdd.n1350 gnd 0.008955f
C3066 vdd.n1352 gnd 0.008955f
C3067 vdd.n1353 gnd 0.008955f
C3068 vdd.n1355 gnd 0.008955f
C3069 vdd.n1356 gnd 0.005983f
C3070 vdd.t33 gnd 0.457591f
C3071 vdd.n1357 gnd 0.008955f
C3072 vdd.n1358 gnd 0.021434f
C3073 vdd.n1359 gnd 0.007208f
C3074 vdd.n1360 gnd 0.008955f
C3075 vdd.n1361 gnd 0.007208f
C3076 vdd.n1362 gnd 0.008955f
C3077 vdd.n1363 gnd 0.915183f
C3078 vdd.n1364 gnd 0.008955f
C3079 vdd.n1365 gnd 0.007208f
C3080 vdd.n1366 gnd 0.007208f
C3081 vdd.n1367 gnd 0.008955f
C3082 vdd.n1368 gnd 0.007208f
C3083 vdd.n1369 gnd 0.008955f
C3084 vdd.t14 gnd 0.457591f
C3085 vdd.n1370 gnd 0.008955f
C3086 vdd.n1371 gnd 0.007208f
C3087 vdd.n1372 gnd 0.008955f
C3088 vdd.n1373 gnd 0.007208f
C3089 vdd.n1374 gnd 0.008955f
C3090 vdd.t20 gnd 0.457591f
C3091 vdd.n1375 gnd 0.008955f
C3092 vdd.n1376 gnd 0.007208f
C3093 vdd.n1377 gnd 0.008955f
C3094 vdd.n1378 gnd 0.007208f
C3095 vdd.n1379 gnd 0.008955f
C3096 vdd.t155 gnd 0.457591f
C3097 vdd.n1380 gnd 0.718418f
C3098 vdd.n1381 gnd 0.008955f
C3099 vdd.n1382 gnd 0.007208f
C3100 vdd.n1383 gnd 0.008955f
C3101 vdd.n1384 gnd 0.007208f
C3102 vdd.n1385 gnd 0.008955f
C3103 vdd.n1386 gnd 0.645204f
C3104 vdd.n1387 gnd 0.008955f
C3105 vdd.n1388 gnd 0.007208f
C3106 vdd.n1389 gnd 0.008955f
C3107 vdd.n1390 gnd 0.007208f
C3108 vdd.n1391 gnd 0.008955f
C3109 vdd.n1392 gnd 0.489623f
C3110 vdd.t10 gnd 0.457591f
C3111 vdd.n1393 gnd 0.008955f
C3112 vdd.n1394 gnd 0.007208f
C3113 vdd.n1395 gnd 0.008925f
C3114 vdd.n1396 gnd 0.007208f
C3115 vdd.n1397 gnd 0.008955f
C3116 vdd.t6 gnd 0.457591f
C3117 vdd.n1398 gnd 0.008955f
C3118 vdd.n1399 gnd 0.007208f
C3119 vdd.n1400 gnd 0.008955f
C3120 vdd.n1401 gnd 0.007208f
C3121 vdd.n1402 gnd 0.008955f
C3122 vdd.t137 gnd 0.457591f
C3123 vdd.n1403 gnd 0.581141f
C3124 vdd.n1404 gnd 0.008955f
C3125 vdd.n1405 gnd 0.007208f
C3126 vdd.n1406 gnd 0.008955f
C3127 vdd.n1407 gnd 0.007208f
C3128 vdd.n1408 gnd 0.008955f
C3129 vdd.t108 gnd 0.457591f
C3130 vdd.n1409 gnd 0.008955f
C3131 vdd.n1410 gnd 0.007208f
C3132 vdd.n1411 gnd 0.008955f
C3133 vdd.n1412 gnd 0.007208f
C3134 vdd.n1413 gnd 0.008955f
C3135 vdd.n1414 gnd 0.6269f
C3136 vdd.n1415 gnd 0.759602f
C3137 vdd.t114 gnd 0.457591f
C3138 vdd.n1416 gnd 0.008955f
C3139 vdd.n1417 gnd 0.007208f
C3140 vdd.n1418 gnd 0.008955f
C3141 vdd.n1419 gnd 0.007208f
C3142 vdd.n1420 gnd 0.008955f
C3143 vdd.n1421 gnd 0.471319f
C3144 vdd.n1422 gnd 0.008955f
C3145 vdd.n1423 gnd 0.007208f
C3146 vdd.n1424 gnd 0.008955f
C3147 vdd.n1425 gnd 0.007208f
C3148 vdd.n1426 gnd 0.008955f
C3149 vdd.n1427 gnd 0.915183f
C3150 vdd.t131 gnd 0.457591f
C3151 vdd.n1428 gnd 0.008955f
C3152 vdd.n1429 gnd 0.007208f
C3153 vdd.n1430 gnd 0.008955f
C3154 vdd.n1431 gnd 0.007208f
C3155 vdd.n1432 gnd 0.008955f
C3156 vdd.t61 gnd 0.457591f
C3157 vdd.n1433 gnd 0.008955f
C3158 vdd.n1434 gnd 0.007208f
C3159 vdd.n1435 gnd 0.021434f
C3160 vdd.n1436 gnd 0.021434f
C3161 vdd.n1437 gnd 2.10492f
C3162 vdd.n1438 gnd 0.517078f
C3163 vdd.n1439 gnd 0.021434f
C3164 vdd.n1440 gnd 0.008955f
C3165 vdd.n1442 gnd 0.008955f
C3166 vdd.n1443 gnd 0.008955f
C3167 vdd.n1444 gnd 0.007208f
C3168 vdd.n1445 gnd 0.008955f
C3169 vdd.n1446 gnd 0.008955f
C3170 vdd.n1448 gnd 0.008955f
C3171 vdd.n1449 gnd 0.008955f
C3172 vdd.n1451 gnd 0.008955f
C3173 vdd.n1452 gnd 0.007208f
C3174 vdd.n1453 gnd 0.008955f
C3175 vdd.n1454 gnd 0.008955f
C3176 vdd.n1456 gnd 0.008955f
C3177 vdd.n1457 gnd 0.008955f
C3178 vdd.n1459 gnd 0.008955f
C3179 vdd.n1460 gnd 0.007208f
C3180 vdd.n1461 gnd 0.008955f
C3181 vdd.n1462 gnd 0.008955f
C3182 vdd.n1464 gnd 0.008955f
C3183 vdd.n1465 gnd 0.008955f
C3184 vdd.n1467 gnd 0.008955f
C3185 vdd.n1468 gnd 0.007208f
C3186 vdd.n1469 gnd 0.008955f
C3187 vdd.n1470 gnd 0.008955f
C3188 vdd.n1472 gnd 0.008955f
C3189 vdd.n1473 gnd 0.008955f
C3190 vdd.n1475 gnd 0.008955f
C3191 vdd.t95 gnd 0.110173f
C3192 vdd.t96 gnd 0.117745f
C3193 vdd.t94 gnd 0.143884f
C3194 vdd.n1476 gnd 0.184439f
C3195 vdd.n1477 gnd 0.155683f
C3196 vdd.n1478 gnd 0.015425f
C3197 vdd.n1479 gnd 0.008955f
C3198 vdd.n1480 gnd 0.008955f
C3199 vdd.n1482 gnd 0.008955f
C3200 vdd.n1483 gnd 0.008955f
C3201 vdd.n1485 gnd 0.008955f
C3202 vdd.n1486 gnd 0.007208f
C3203 vdd.n1487 gnd 0.008955f
C3204 vdd.n1488 gnd 0.008955f
C3205 vdd.n1490 gnd 0.008955f
C3206 vdd.n1491 gnd 0.008955f
C3207 vdd.n1493 gnd 0.008955f
C3208 vdd.n1494 gnd 0.007208f
C3209 vdd.n1495 gnd 0.008955f
C3210 vdd.n1496 gnd 0.008955f
C3211 vdd.n1498 gnd 0.008955f
C3212 vdd.n1499 gnd 0.008955f
C3213 vdd.n1501 gnd 0.008955f
C3214 vdd.n1502 gnd 0.007208f
C3215 vdd.n1503 gnd 0.008955f
C3216 vdd.n1504 gnd 0.008955f
C3217 vdd.n1506 gnd 0.008955f
C3218 vdd.n1507 gnd 0.008955f
C3219 vdd.n1509 gnd 0.008955f
C3220 vdd.n1510 gnd 0.007208f
C3221 vdd.n1511 gnd 0.008955f
C3222 vdd.n1512 gnd 0.008955f
C3223 vdd.n1514 gnd 0.008955f
C3224 vdd.n1515 gnd 0.008955f
C3225 vdd.n1517 gnd 0.008955f
C3226 vdd.n1518 gnd 0.007208f
C3227 vdd.n1519 gnd 0.008955f
C3228 vdd.n1520 gnd 0.008955f
C3229 vdd.n1522 gnd 0.008955f
C3230 vdd.n1523 gnd 0.007136f
C3231 vdd.n1525 gnd 0.007208f
C3232 vdd.n1526 gnd 0.008955f
C3233 vdd.n1527 gnd 0.008955f
C3234 vdd.n1528 gnd 0.008955f
C3235 vdd.n1529 gnd 0.008955f
C3236 vdd.n1531 gnd 0.008955f
C3237 vdd.n1532 gnd 0.008955f
C3238 vdd.n1533 gnd 0.007208f
C3239 vdd.n1534 gnd 0.008955f
C3240 vdd.n1536 gnd 0.008955f
C3241 vdd.n1537 gnd 0.008955f
C3242 vdd.n1539 gnd 0.008955f
C3243 vdd.n1540 gnd 0.008955f
C3244 vdd.n1541 gnd 0.007208f
C3245 vdd.n1542 gnd 0.008955f
C3246 vdd.n1544 gnd 0.008955f
C3247 vdd.n1545 gnd 0.008955f
C3248 vdd.n1547 gnd 0.008955f
C3249 vdd.n1548 gnd 0.008955f
C3250 vdd.n1549 gnd 0.007208f
C3251 vdd.n1550 gnd 0.008955f
C3252 vdd.n1552 gnd 0.008955f
C3253 vdd.n1553 gnd 0.008955f
C3254 vdd.n1555 gnd 0.008955f
C3255 vdd.n1556 gnd 0.008955f
C3256 vdd.n1557 gnd 0.007208f
C3257 vdd.n1558 gnd 0.008955f
C3258 vdd.n1560 gnd 0.008955f
C3259 vdd.n1561 gnd 0.008955f
C3260 vdd.n1563 gnd 0.008955f
C3261 vdd.n1564 gnd 0.003424f
C3262 vdd.t62 gnd 0.110173f
C3263 vdd.t63 gnd 0.117745f
C3264 vdd.t60 gnd 0.143884f
C3265 vdd.n1565 gnd 0.184439f
C3266 vdd.n1566 gnd 0.155683f
C3267 vdd.n1567 gnd 0.011821f
C3268 vdd.n1568 gnd 0.003784f
C3269 vdd.n1569 gnd 0.007208f
C3270 vdd.n1570 gnd 0.008955f
C3271 vdd.n1571 gnd 0.008955f
C3272 vdd.n1572 gnd 0.008955f
C3273 vdd.n1573 gnd 0.007208f
C3274 vdd.n1574 gnd 0.007208f
C3275 vdd.n1575 gnd 0.007208f
C3276 vdd.n1576 gnd 0.008955f
C3277 vdd.n1577 gnd 0.008955f
C3278 vdd.n1578 gnd 0.008955f
C3279 vdd.n1579 gnd 0.007208f
C3280 vdd.n1580 gnd 0.007208f
C3281 vdd.n1581 gnd 0.007208f
C3282 vdd.n1582 gnd 0.008955f
C3283 vdd.n1583 gnd 0.008955f
C3284 vdd.n1584 gnd 0.008955f
C3285 vdd.n1585 gnd 0.007208f
C3286 vdd.n1586 gnd 0.007208f
C3287 vdd.n1587 gnd 0.007208f
C3288 vdd.n1588 gnd 0.008955f
C3289 vdd.n1589 gnd 0.008955f
C3290 vdd.n1590 gnd 0.008955f
C3291 vdd.n1591 gnd 0.007208f
C3292 vdd.n1592 gnd 0.007208f
C3293 vdd.n1593 gnd 0.007208f
C3294 vdd.n1594 gnd 0.008955f
C3295 vdd.n1595 gnd 0.008955f
C3296 vdd.n1596 gnd 0.008955f
C3297 vdd.n1597 gnd 0.007208f
C3298 vdd.n1598 gnd 0.008955f
C3299 vdd.n1599 gnd 0.008955f
C3300 vdd.n1601 gnd 0.008955f
C3301 vdd.t85 gnd 0.110173f
C3302 vdd.t86 gnd 0.117745f
C3303 vdd.t84 gnd 0.143884f
C3304 vdd.n1602 gnd 0.184439f
C3305 vdd.n1603 gnd 0.155683f
C3306 vdd.n1604 gnd 0.015425f
C3307 vdd.n1605 gnd 0.004901f
C3308 vdd.n1606 gnd 0.008955f
C3309 vdd.n1607 gnd 0.008955f
C3310 vdd.n1608 gnd 0.008955f
C3311 vdd.n1609 gnd 0.007208f
C3312 vdd.n1610 gnd 0.007208f
C3313 vdd.n1611 gnd 0.007208f
C3314 vdd.n1612 gnd 0.008955f
C3315 vdd.n1613 gnd 0.008955f
C3316 vdd.n1614 gnd 0.008955f
C3317 vdd.n1615 gnd 0.007208f
C3318 vdd.n1616 gnd 0.007208f
C3319 vdd.n1617 gnd 0.007208f
C3320 vdd.n1618 gnd 0.008955f
C3321 vdd.n1619 gnd 0.008955f
C3322 vdd.n1620 gnd 0.008955f
C3323 vdd.n1621 gnd 0.007208f
C3324 vdd.n1622 gnd 0.007208f
C3325 vdd.n1623 gnd 0.007208f
C3326 vdd.n1624 gnd 0.008955f
C3327 vdd.n1625 gnd 0.008955f
C3328 vdd.n1626 gnd 0.008955f
C3329 vdd.n1627 gnd 0.007208f
C3330 vdd.n1628 gnd 0.007208f
C3331 vdd.n1629 gnd 0.007208f
C3332 vdd.n1630 gnd 0.008955f
C3333 vdd.n1631 gnd 0.008955f
C3334 vdd.n1632 gnd 0.008955f
C3335 vdd.n1633 gnd 0.007208f
C3336 vdd.n1634 gnd 0.007208f
C3337 vdd.n1635 gnd 0.006019f
C3338 vdd.n1636 gnd 0.008955f
C3339 vdd.n1637 gnd 0.008955f
C3340 vdd.n1638 gnd 0.008955f
C3341 vdd.n1639 gnd 0.006019f
C3342 vdd.n1640 gnd 0.007208f
C3343 vdd.n1641 gnd 0.007208f
C3344 vdd.n1642 gnd 0.008955f
C3345 vdd.n1643 gnd 0.008955f
C3346 vdd.n1644 gnd 0.008955f
C3347 vdd.n1645 gnd 0.007208f
C3348 vdd.n1646 gnd 0.007208f
C3349 vdd.n1647 gnd 0.007208f
C3350 vdd.n1648 gnd 0.008955f
C3351 vdd.n1649 gnd 0.008955f
C3352 vdd.n1650 gnd 0.008955f
C3353 vdd.n1651 gnd 0.007208f
C3354 vdd.n1652 gnd 0.007208f
C3355 vdd.n1653 gnd 0.007208f
C3356 vdd.n1654 gnd 0.008955f
C3357 vdd.n1655 gnd 0.008955f
C3358 vdd.n1656 gnd 0.008955f
C3359 vdd.n1657 gnd 0.007208f
C3360 vdd.n1658 gnd 0.007208f
C3361 vdd.n1659 gnd 0.007208f
C3362 vdd.n1660 gnd 0.008955f
C3363 vdd.n1661 gnd 0.008955f
C3364 vdd.n1662 gnd 0.008955f
C3365 vdd.n1663 gnd 0.007208f
C3366 vdd.n1664 gnd 0.007208f
C3367 vdd.n1665 gnd 0.005983f
C3368 vdd.n1666 gnd 0.021434f
C3369 vdd.n1667 gnd 0.021104f
C3370 vdd.n1668 gnd 0.005983f
C3371 vdd.n1669 gnd 0.021104f
C3372 vdd.n1670 gnd 1.29041f
C3373 vdd.n1671 gnd 0.021104f
C3374 vdd.n1672 gnd 0.005983f
C3375 vdd.n1673 gnd 0.021104f
C3376 vdd.n1674 gnd 0.008955f
C3377 vdd.n1675 gnd 0.008955f
C3378 vdd.n1676 gnd 0.007208f
C3379 vdd.n1677 gnd 0.008955f
C3380 vdd.n1678 gnd 0.855696f
C3381 vdd.n1679 gnd 0.008955f
C3382 vdd.n1680 gnd 0.007208f
C3383 vdd.n1681 gnd 0.008955f
C3384 vdd.n1682 gnd 0.008955f
C3385 vdd.n1683 gnd 0.008955f
C3386 vdd.n1684 gnd 0.007208f
C3387 vdd.n1685 gnd 0.008955f
C3388 vdd.n1686 gnd 0.901455f
C3389 vdd.n1687 gnd 0.008955f
C3390 vdd.n1688 gnd 0.007208f
C3391 vdd.n1689 gnd 0.008955f
C3392 vdd.n1690 gnd 0.008955f
C3393 vdd.n1691 gnd 0.008955f
C3394 vdd.n1692 gnd 0.007208f
C3395 vdd.n1693 gnd 0.008955f
C3396 vdd.t8 gnd 0.457591f
C3397 vdd.n1694 gnd 0.745874f
C3398 vdd.n1695 gnd 0.008955f
C3399 vdd.n1696 gnd 0.007208f
C3400 vdd.n1697 gnd 0.008955f
C3401 vdd.n1698 gnd 0.008955f
C3402 vdd.n1699 gnd 0.008955f
C3403 vdd.n1700 gnd 0.007208f
C3404 vdd.n1701 gnd 0.008955f
C3405 vdd.n1702 gnd 0.590293f
C3406 vdd.n1703 gnd 0.008955f
C3407 vdd.n1704 gnd 0.007208f
C3408 vdd.n1705 gnd 0.008955f
C3409 vdd.n1706 gnd 0.008955f
C3410 vdd.n1707 gnd 0.008955f
C3411 vdd.n1708 gnd 0.007208f
C3412 vdd.n1709 gnd 0.008955f
C3413 vdd.n1710 gnd 0.736722f
C3414 vdd.n1711 gnd 0.480471f
C3415 vdd.n1712 gnd 0.008955f
C3416 vdd.n1713 gnd 0.007208f
C3417 vdd.n1714 gnd 0.008955f
C3418 vdd.n1715 gnd 0.008955f
C3419 vdd.n1716 gnd 0.008955f
C3420 vdd.n1717 gnd 0.007208f
C3421 vdd.n1718 gnd 0.008955f
C3422 vdd.n1719 gnd 0.636052f
C3423 vdd.n1720 gnd 0.008955f
C3424 vdd.n1721 gnd 0.007208f
C3425 vdd.n1722 gnd 0.008955f
C3426 vdd.n1723 gnd 0.008955f
C3427 vdd.n1724 gnd 0.008955f
C3428 vdd.n1725 gnd 0.007208f
C3429 vdd.n1726 gnd 0.008955f
C3430 vdd.t18 gnd 0.457591f
C3431 vdd.n1727 gnd 0.759602f
C3432 vdd.n1728 gnd 0.008955f
C3433 vdd.n1729 gnd 0.007208f
C3434 vdd.n1730 gnd 0.004915f
C3435 vdd.n1731 gnd 0.004561f
C3436 vdd.n1732 gnd 0.002523f
C3437 vdd.n1733 gnd 0.005793f
C3438 vdd.n1734 gnd 0.002451f
C3439 vdd.n1735 gnd 0.002595f
C3440 vdd.n1736 gnd 0.004561f
C3441 vdd.n1737 gnd 0.002451f
C3442 vdd.n1738 gnd 0.005793f
C3443 vdd.n1739 gnd 0.002595f
C3444 vdd.n1740 gnd 0.004561f
C3445 vdd.n1741 gnd 0.002451f
C3446 vdd.n1742 gnd 0.004344f
C3447 vdd.n1743 gnd 0.004357f
C3448 vdd.t15 gnd 0.012445f
C3449 vdd.n1744 gnd 0.027689f
C3450 vdd.n1745 gnd 0.144102f
C3451 vdd.n1746 gnd 0.002451f
C3452 vdd.n1747 gnd 0.002595f
C3453 vdd.n1748 gnd 0.005793f
C3454 vdd.n1749 gnd 0.005793f
C3455 vdd.n1750 gnd 0.002595f
C3456 vdd.n1751 gnd 0.002451f
C3457 vdd.n1752 gnd 0.004561f
C3458 vdd.n1753 gnd 0.004561f
C3459 vdd.n1754 gnd 0.002451f
C3460 vdd.n1755 gnd 0.002595f
C3461 vdd.n1756 gnd 0.005793f
C3462 vdd.n1757 gnd 0.005793f
C3463 vdd.n1758 gnd 0.002595f
C3464 vdd.n1759 gnd 0.002451f
C3465 vdd.n1760 gnd 0.004561f
C3466 vdd.n1761 gnd 0.004561f
C3467 vdd.n1762 gnd 0.002451f
C3468 vdd.n1763 gnd 0.002595f
C3469 vdd.n1764 gnd 0.005793f
C3470 vdd.n1765 gnd 0.005793f
C3471 vdd.n1766 gnd 0.013695f
C3472 vdd.n1767 gnd 0.002523f
C3473 vdd.n1768 gnd 0.002451f
C3474 vdd.n1769 gnd 0.011788f
C3475 vdd.n1770 gnd 0.00823f
C3476 vdd.t216 gnd 0.028831f
C3477 vdd.t21 gnd 0.028831f
C3478 vdd.n1771 gnd 0.19815f
C3479 vdd.n1772 gnd 0.155815f
C3480 vdd.t222 gnd 0.028831f
C3481 vdd.t227 gnd 0.028831f
C3482 vdd.n1773 gnd 0.19815f
C3483 vdd.n1774 gnd 0.125742f
C3484 vdd.t242 gnd 0.028831f
C3485 vdd.t228 gnd 0.028831f
C3486 vdd.n1775 gnd 0.19815f
C3487 vdd.n1776 gnd 0.125742f
C3488 vdd.t127 gnd 0.028831f
C3489 vdd.t138 gnd 0.028831f
C3490 vdd.n1777 gnd 0.19815f
C3491 vdd.n1778 gnd 0.125742f
C3492 vdd.t105 gnd 0.028831f
C3493 vdd.t115 gnd 0.028831f
C3494 vdd.n1779 gnd 0.19815f
C3495 vdd.n1780 gnd 0.125742f
C3496 vdd.n1781 gnd 0.004915f
C3497 vdd.n1782 gnd 0.004561f
C3498 vdd.n1783 gnd 0.002523f
C3499 vdd.n1784 gnd 0.005793f
C3500 vdd.n1785 gnd 0.002451f
C3501 vdd.n1786 gnd 0.002595f
C3502 vdd.n1787 gnd 0.004561f
C3503 vdd.n1788 gnd 0.002451f
C3504 vdd.n1789 gnd 0.005793f
C3505 vdd.n1790 gnd 0.002595f
C3506 vdd.n1791 gnd 0.004561f
C3507 vdd.n1792 gnd 0.002451f
C3508 vdd.n1793 gnd 0.004344f
C3509 vdd.n1794 gnd 0.004357f
C3510 vdd.t240 gnd 0.012445f
C3511 vdd.n1795 gnd 0.027689f
C3512 vdd.n1796 gnd 0.144102f
C3513 vdd.n1797 gnd 0.002451f
C3514 vdd.n1798 gnd 0.002595f
C3515 vdd.n1799 gnd 0.005793f
C3516 vdd.n1800 gnd 0.005793f
C3517 vdd.n1801 gnd 0.002595f
C3518 vdd.n1802 gnd 0.002451f
C3519 vdd.n1803 gnd 0.004561f
C3520 vdd.n1804 gnd 0.004561f
C3521 vdd.n1805 gnd 0.002451f
C3522 vdd.n1806 gnd 0.002595f
C3523 vdd.n1807 gnd 0.005793f
C3524 vdd.n1808 gnd 0.005793f
C3525 vdd.n1809 gnd 0.002595f
C3526 vdd.n1810 gnd 0.002451f
C3527 vdd.n1811 gnd 0.004561f
C3528 vdd.n1812 gnd 0.004561f
C3529 vdd.n1813 gnd 0.002451f
C3530 vdd.n1814 gnd 0.002595f
C3531 vdd.n1815 gnd 0.005793f
C3532 vdd.n1816 gnd 0.005793f
C3533 vdd.n1817 gnd 0.013695f
C3534 vdd.n1818 gnd 0.002523f
C3535 vdd.n1819 gnd 0.002451f
C3536 vdd.n1820 gnd 0.011788f
C3537 vdd.n1821 gnd 0.007971f
C3538 vdd.n1822 gnd 0.093552f
C3539 vdd.n1823 gnd 0.004915f
C3540 vdd.n1824 gnd 0.004561f
C3541 vdd.n1825 gnd 0.002523f
C3542 vdd.n1826 gnd 0.005793f
C3543 vdd.n1827 gnd 0.002451f
C3544 vdd.n1828 gnd 0.002595f
C3545 vdd.n1829 gnd 0.004561f
C3546 vdd.n1830 gnd 0.002451f
C3547 vdd.n1831 gnd 0.005793f
C3548 vdd.n1832 gnd 0.002595f
C3549 vdd.n1833 gnd 0.004561f
C3550 vdd.n1834 gnd 0.002451f
C3551 vdd.n1835 gnd 0.004344f
C3552 vdd.n1836 gnd 0.004357f
C3553 vdd.t102 gnd 0.012445f
C3554 vdd.n1837 gnd 0.027689f
C3555 vdd.n1838 gnd 0.144102f
C3556 vdd.n1839 gnd 0.002451f
C3557 vdd.n1840 gnd 0.002595f
C3558 vdd.n1841 gnd 0.005793f
C3559 vdd.n1842 gnd 0.005793f
C3560 vdd.n1843 gnd 0.002595f
C3561 vdd.n1844 gnd 0.002451f
C3562 vdd.n1845 gnd 0.004561f
C3563 vdd.n1846 gnd 0.004561f
C3564 vdd.n1847 gnd 0.002451f
C3565 vdd.n1848 gnd 0.002595f
C3566 vdd.n1849 gnd 0.005793f
C3567 vdd.n1850 gnd 0.005793f
C3568 vdd.n1851 gnd 0.002595f
C3569 vdd.n1852 gnd 0.002451f
C3570 vdd.n1853 gnd 0.004561f
C3571 vdd.n1854 gnd 0.004561f
C3572 vdd.n1855 gnd 0.002451f
C3573 vdd.n1856 gnd 0.002595f
C3574 vdd.n1857 gnd 0.005793f
C3575 vdd.n1858 gnd 0.005793f
C3576 vdd.n1859 gnd 0.013695f
C3577 vdd.n1860 gnd 0.002523f
C3578 vdd.n1861 gnd 0.002451f
C3579 vdd.n1862 gnd 0.011788f
C3580 vdd.n1863 gnd 0.00823f
C3581 vdd.t243 gnd 0.028831f
C3582 vdd.t113 gnd 0.028831f
C3583 vdd.n1864 gnd 0.19815f
C3584 vdd.n1865 gnd 0.155815f
C3585 vdd.t229 gnd 0.028831f
C3586 vdd.t136 gnd 0.028831f
C3587 vdd.n1866 gnd 0.19815f
C3588 vdd.n1867 gnd 0.125742f
C3589 vdd.t7 gnd 0.028831f
C3590 vdd.t19 gnd 0.028831f
C3591 vdd.n1868 gnd 0.19815f
C3592 vdd.n1869 gnd 0.125742f
C3593 vdd.t221 gnd 0.028831f
C3594 vdd.t224 gnd 0.028831f
C3595 vdd.n1870 gnd 0.19815f
C3596 vdd.n1871 gnd 0.125742f
C3597 vdd.t9 gnd 0.028831f
C3598 vdd.t124 gnd 0.028831f
C3599 vdd.n1872 gnd 0.19815f
C3600 vdd.n1873 gnd 0.125742f
C3601 vdd.n1874 gnd 0.004915f
C3602 vdd.n1875 gnd 0.004561f
C3603 vdd.n1876 gnd 0.002523f
C3604 vdd.n1877 gnd 0.005793f
C3605 vdd.n1878 gnd 0.002451f
C3606 vdd.n1879 gnd 0.002595f
C3607 vdd.n1880 gnd 0.004561f
C3608 vdd.n1881 gnd 0.002451f
C3609 vdd.n1882 gnd 0.005793f
C3610 vdd.n1883 gnd 0.002595f
C3611 vdd.n1884 gnd 0.004561f
C3612 vdd.n1885 gnd 0.002451f
C3613 vdd.n1886 gnd 0.004344f
C3614 vdd.n1887 gnd 0.004357f
C3615 vdd.t153 gnd 0.012445f
C3616 vdd.n1888 gnd 0.027689f
C3617 vdd.n1889 gnd 0.144102f
C3618 vdd.n1890 gnd 0.002451f
C3619 vdd.n1891 gnd 0.002595f
C3620 vdd.n1892 gnd 0.005793f
C3621 vdd.n1893 gnd 0.005793f
C3622 vdd.n1894 gnd 0.002595f
C3623 vdd.n1895 gnd 0.002451f
C3624 vdd.n1896 gnd 0.004561f
C3625 vdd.n1897 gnd 0.004561f
C3626 vdd.n1898 gnd 0.002451f
C3627 vdd.n1899 gnd 0.002595f
C3628 vdd.n1900 gnd 0.005793f
C3629 vdd.n1901 gnd 0.005793f
C3630 vdd.n1902 gnd 0.002595f
C3631 vdd.n1903 gnd 0.002451f
C3632 vdd.n1904 gnd 0.004561f
C3633 vdd.n1905 gnd 0.004561f
C3634 vdd.n1906 gnd 0.002451f
C3635 vdd.n1907 gnd 0.002595f
C3636 vdd.n1908 gnd 0.005793f
C3637 vdd.n1909 gnd 0.005793f
C3638 vdd.n1910 gnd 0.013695f
C3639 vdd.n1911 gnd 0.002523f
C3640 vdd.n1912 gnd 0.002451f
C3641 vdd.n1913 gnd 0.011788f
C3642 vdd.n1914 gnd 0.007971f
C3643 vdd.n1915 gnd 0.055654f
C3644 vdd.n1916 gnd 0.200537f
C3645 vdd.n1917 gnd 0.004915f
C3646 vdd.n1918 gnd 0.004561f
C3647 vdd.n1919 gnd 0.002523f
C3648 vdd.n1920 gnd 0.005793f
C3649 vdd.n1921 gnd 0.002451f
C3650 vdd.n1922 gnd 0.002595f
C3651 vdd.n1923 gnd 0.004561f
C3652 vdd.n1924 gnd 0.002451f
C3653 vdd.n1925 gnd 0.005793f
C3654 vdd.n1926 gnd 0.002595f
C3655 vdd.n1927 gnd 0.004561f
C3656 vdd.n1928 gnd 0.002451f
C3657 vdd.n1929 gnd 0.004344f
C3658 vdd.n1930 gnd 0.004357f
C3659 vdd.t220 gnd 0.012445f
C3660 vdd.n1931 gnd 0.027689f
C3661 vdd.n1932 gnd 0.144102f
C3662 vdd.n1933 gnd 0.002451f
C3663 vdd.n1934 gnd 0.002595f
C3664 vdd.n1935 gnd 0.005793f
C3665 vdd.n1936 gnd 0.005793f
C3666 vdd.n1937 gnd 0.002595f
C3667 vdd.n1938 gnd 0.002451f
C3668 vdd.n1939 gnd 0.004561f
C3669 vdd.n1940 gnd 0.004561f
C3670 vdd.n1941 gnd 0.002451f
C3671 vdd.n1942 gnd 0.002595f
C3672 vdd.n1943 gnd 0.005793f
C3673 vdd.n1944 gnd 0.005793f
C3674 vdd.n1945 gnd 0.002595f
C3675 vdd.n1946 gnd 0.002451f
C3676 vdd.n1947 gnd 0.004561f
C3677 vdd.n1948 gnd 0.004561f
C3678 vdd.n1949 gnd 0.002451f
C3679 vdd.n1950 gnd 0.002595f
C3680 vdd.n1951 gnd 0.005793f
C3681 vdd.n1952 gnd 0.005793f
C3682 vdd.n1953 gnd 0.013695f
C3683 vdd.n1954 gnd 0.002523f
C3684 vdd.n1955 gnd 0.002451f
C3685 vdd.n1956 gnd 0.011788f
C3686 vdd.n1957 gnd 0.00823f
C3687 vdd.t156 gnd 0.028831f
C3688 vdd.t157 gnd 0.028831f
C3689 vdd.n1958 gnd 0.19815f
C3690 vdd.n1959 gnd 0.155815f
C3691 vdd.t11 gnd 0.028831f
C3692 vdd.t145 gnd 0.028831f
C3693 vdd.n1960 gnd 0.19815f
C3694 vdd.n1961 gnd 0.125742f
C3695 vdd.t226 gnd 0.028831f
C3696 vdd.t118 gnd 0.028831f
C3697 vdd.n1962 gnd 0.19815f
C3698 vdd.n1963 gnd 0.125742f
C3699 vdd.t109 gnd 0.028831f
C3700 vdd.t146 gnd 0.028831f
C3701 vdd.n1964 gnd 0.19815f
C3702 vdd.n1965 gnd 0.125742f
C3703 vdd.t237 gnd 0.028831f
C3704 vdd.t159 gnd 0.028831f
C3705 vdd.n1966 gnd 0.19815f
C3706 vdd.n1967 gnd 0.125742f
C3707 vdd.n1968 gnd 0.004915f
C3708 vdd.n1969 gnd 0.004561f
C3709 vdd.n1970 gnd 0.002523f
C3710 vdd.n1971 gnd 0.005793f
C3711 vdd.n1972 gnd 0.002451f
C3712 vdd.n1973 gnd 0.002595f
C3713 vdd.n1974 gnd 0.004561f
C3714 vdd.n1975 gnd 0.002451f
C3715 vdd.n1976 gnd 0.005793f
C3716 vdd.n1977 gnd 0.002595f
C3717 vdd.n1978 gnd 0.004561f
C3718 vdd.n1979 gnd 0.002451f
C3719 vdd.n1980 gnd 0.004344f
C3720 vdd.n1981 gnd 0.004357f
C3721 vdd.t132 gnd 0.012445f
C3722 vdd.n1982 gnd 0.027689f
C3723 vdd.n1983 gnd 0.144102f
C3724 vdd.n1984 gnd 0.002451f
C3725 vdd.n1985 gnd 0.002595f
C3726 vdd.n1986 gnd 0.005793f
C3727 vdd.n1987 gnd 0.005793f
C3728 vdd.n1988 gnd 0.002595f
C3729 vdd.n1989 gnd 0.002451f
C3730 vdd.n1990 gnd 0.004561f
C3731 vdd.n1991 gnd 0.004561f
C3732 vdd.n1992 gnd 0.002451f
C3733 vdd.n1993 gnd 0.002595f
C3734 vdd.n1994 gnd 0.005793f
C3735 vdd.n1995 gnd 0.005793f
C3736 vdd.n1996 gnd 0.002595f
C3737 vdd.n1997 gnd 0.002451f
C3738 vdd.n1998 gnd 0.004561f
C3739 vdd.n1999 gnd 0.004561f
C3740 vdd.n2000 gnd 0.002451f
C3741 vdd.n2001 gnd 0.002595f
C3742 vdd.n2002 gnd 0.005793f
C3743 vdd.n2003 gnd 0.005793f
C3744 vdd.n2004 gnd 0.013695f
C3745 vdd.n2005 gnd 0.002523f
C3746 vdd.n2006 gnd 0.002451f
C3747 vdd.n2007 gnd 0.011788f
C3748 vdd.n2008 gnd 0.007971f
C3749 vdd.n2009 gnd 0.055654f
C3750 vdd.n2010 gnd 0.220396f
C3751 vdd.n2011 gnd 2.30824f
C3752 vdd.n2012 gnd 0.533085f
C3753 vdd.n2013 gnd 0.008925f
C3754 vdd.n2014 gnd 0.008955f
C3755 vdd.n2015 gnd 0.007208f
C3756 vdd.n2016 gnd 0.008955f
C3757 vdd.n2017 gnd 0.72757f
C3758 vdd.n2018 gnd 0.008955f
C3759 vdd.n2019 gnd 0.007208f
C3760 vdd.n2020 gnd 0.008955f
C3761 vdd.n2021 gnd 0.008955f
C3762 vdd.n2022 gnd 0.008955f
C3763 vdd.n2023 gnd 0.007208f
C3764 vdd.n2024 gnd 0.008955f
C3765 vdd.n2025 gnd 0.759602f
C3766 vdd.t135 gnd 0.457591f
C3767 vdd.n2026 gnd 0.571989f
C3768 vdd.n2027 gnd 0.008955f
C3769 vdd.n2028 gnd 0.007208f
C3770 vdd.n2029 gnd 0.008955f
C3771 vdd.n2030 gnd 0.008955f
C3772 vdd.n2031 gnd 0.008955f
C3773 vdd.n2032 gnd 0.007208f
C3774 vdd.n2033 gnd 0.008955f
C3775 vdd.n2034 gnd 0.498775f
C3776 vdd.n2035 gnd 0.008955f
C3777 vdd.n2036 gnd 0.007208f
C3778 vdd.n2037 gnd 0.008955f
C3779 vdd.n2038 gnd 0.008955f
C3780 vdd.n2039 gnd 0.008955f
C3781 vdd.n2040 gnd 0.007208f
C3782 vdd.n2041 gnd 0.008955f
C3783 vdd.n2042 gnd 0.562837f
C3784 vdd.n2043 gnd 0.654356f
C3785 vdd.n2044 gnd 0.008955f
C3786 vdd.n2045 gnd 0.007208f
C3787 vdd.n2046 gnd 0.008955f
C3788 vdd.n2047 gnd 0.008955f
C3789 vdd.n2048 gnd 0.008955f
C3790 vdd.n2049 gnd 0.007208f
C3791 vdd.n2050 gnd 0.008955f
C3792 vdd.n2051 gnd 0.809937f
C3793 vdd.n2052 gnd 0.008955f
C3794 vdd.n2053 gnd 0.007208f
C3795 vdd.n2054 gnd 0.008955f
C3796 vdd.n2055 gnd 0.008955f
C3797 vdd.n2056 gnd 0.021104f
C3798 vdd.n2057 gnd 0.008955f
C3799 vdd.n2058 gnd 0.008955f
C3800 vdd.n2059 gnd 0.007208f
C3801 vdd.n2060 gnd 0.008955f
C3802 vdd.n2061 gnd 0.489623f
C3803 vdd.n2062 gnd 0.915183f
C3804 vdd.n2063 gnd 0.008955f
C3805 vdd.n2064 gnd 0.007208f
C3806 vdd.n2065 gnd 0.008955f
C3807 vdd.n2066 gnd 0.008955f
C3808 vdd.n2067 gnd 0.021104f
C3809 vdd.n2068 gnd 0.005983f
C3810 vdd.n2069 gnd 0.021104f
C3811 vdd.n2070 gnd 1.25838f
C3812 vdd.n2071 gnd 0.021104f
C3813 vdd.n2072 gnd 0.021434f
C3814 vdd.n2073 gnd 0.003424f
C3815 vdd.t56 gnd 0.110173f
C3816 vdd.t55 gnd 0.117745f
C3817 vdd.t54 gnd 0.143884f
C3818 vdd.n2074 gnd 0.184439f
C3819 vdd.n2075 gnd 0.154963f
C3820 vdd.n2076 gnd 0.0111f
C3821 vdd.n2077 gnd 0.003784f
C3822 vdd.n2078 gnd 0.007702f
C3823 vdd.n2079 gnd 0.95069f
C3824 vdd.n2081 gnd 0.007208f
C3825 vdd.n2082 gnd 0.007208f
C3826 vdd.n2083 gnd 0.008955f
C3827 vdd.n2085 gnd 0.008955f
C3828 vdd.n2086 gnd 0.008955f
C3829 vdd.n2087 gnd 0.007208f
C3830 vdd.n2088 gnd 0.007208f
C3831 vdd.n2089 gnd 0.007208f
C3832 vdd.n2090 gnd 0.008955f
C3833 vdd.n2092 gnd 0.008955f
C3834 vdd.n2093 gnd 0.008955f
C3835 vdd.n2094 gnd 0.007208f
C3836 vdd.n2095 gnd 0.007208f
C3837 vdd.n2096 gnd 0.007208f
C3838 vdd.n2097 gnd 0.008955f
C3839 vdd.n2099 gnd 0.008955f
C3840 vdd.n2100 gnd 0.008955f
C3841 vdd.n2101 gnd 0.007208f
C3842 vdd.n2102 gnd 0.007208f
C3843 vdd.n2103 gnd 0.007208f
C3844 vdd.n2104 gnd 0.008955f
C3845 vdd.n2106 gnd 0.008955f
C3846 vdd.n2107 gnd 0.008955f
C3847 vdd.n2108 gnd 0.007208f
C3848 vdd.n2109 gnd 0.008955f
C3849 vdd.n2110 gnd 0.008955f
C3850 vdd.n2111 gnd 0.008955f
C3851 vdd.n2112 gnd 0.014704f
C3852 vdd.n2113 gnd 0.004901f
C3853 vdd.n2114 gnd 0.007208f
C3854 vdd.n2115 gnd 0.008955f
C3855 vdd.n2117 gnd 0.008955f
C3856 vdd.n2118 gnd 0.008955f
C3857 vdd.n2119 gnd 0.007208f
C3858 vdd.n2120 gnd 0.007208f
C3859 vdd.n2121 gnd 0.007208f
C3860 vdd.n2122 gnd 0.008955f
C3861 vdd.n2124 gnd 0.008955f
C3862 vdd.n2125 gnd 0.008955f
C3863 vdd.n2126 gnd 0.007208f
C3864 vdd.n2127 gnd 0.007208f
C3865 vdd.n2128 gnd 0.007208f
C3866 vdd.n2129 gnd 0.008955f
C3867 vdd.n2131 gnd 0.008955f
C3868 vdd.n2132 gnd 0.008955f
C3869 vdd.n2133 gnd 0.007208f
C3870 vdd.n2134 gnd 0.007208f
C3871 vdd.n2135 gnd 0.007208f
C3872 vdd.n2136 gnd 0.008955f
C3873 vdd.n2138 gnd 0.008955f
C3874 vdd.n2139 gnd 0.008955f
C3875 vdd.n2140 gnd 0.007208f
C3876 vdd.n2141 gnd 0.007208f
C3877 vdd.n2142 gnd 0.007208f
C3878 vdd.n2143 gnd 0.008955f
C3879 vdd.n2145 gnd 0.008955f
C3880 vdd.n2146 gnd 0.008955f
C3881 vdd.n2147 gnd 0.007208f
C3882 vdd.n2148 gnd 0.008955f
C3883 vdd.n2149 gnd 0.008955f
C3884 vdd.n2150 gnd 0.008955f
C3885 vdd.n2151 gnd 0.014704f
C3886 vdd.n2152 gnd 0.006019f
C3887 vdd.n2153 gnd 0.007208f
C3888 vdd.n2154 gnd 0.008955f
C3889 vdd.n2156 gnd 0.008955f
C3890 vdd.n2157 gnd 0.008955f
C3891 vdd.n2158 gnd 0.007208f
C3892 vdd.n2159 gnd 0.007208f
C3893 vdd.n2160 gnd 0.007208f
C3894 vdd.n2161 gnd 0.008955f
C3895 vdd.n2163 gnd 0.008955f
C3896 vdd.n2164 gnd 0.008955f
C3897 vdd.n2165 gnd 0.007208f
C3898 vdd.n2166 gnd 0.007208f
C3899 vdd.n2167 gnd 0.007208f
C3900 vdd.n2168 gnd 0.008955f
C3901 vdd.n2170 gnd 0.008955f
C3902 vdd.n2171 gnd 0.008955f
C3903 vdd.n2172 gnd 0.007208f
C3904 vdd.n2173 gnd 0.007208f
C3905 vdd.n2174 gnd 0.007208f
C3906 vdd.n2175 gnd 0.008955f
C3907 vdd.n2177 gnd 0.008955f
C3908 vdd.n2178 gnd 0.007208f
C3909 vdd.n2179 gnd 0.007208f
C3910 vdd.n2180 gnd 0.008955f
C3911 vdd.n2182 gnd 0.008955f
C3912 vdd.n2183 gnd 0.008955f
C3913 vdd.n2184 gnd 0.007208f
C3914 vdd.n2185 gnd 0.007702f
C3915 vdd.n2186 gnd 0.95069f
C3916 vdd.n2187 gnd 0.041023f
C3917 vdd.n2188 gnd 0.00609f
C3918 vdd.n2189 gnd 0.00609f
C3919 vdd.n2190 gnd 0.00609f
C3920 vdd.n2191 gnd 0.00609f
C3921 vdd.n2192 gnd 0.00609f
C3922 vdd.n2193 gnd 0.00609f
C3923 vdd.n2194 gnd 0.00609f
C3924 vdd.n2195 gnd 0.00609f
C3925 vdd.n2196 gnd 0.00609f
C3926 vdd.n2197 gnd 0.00609f
C3927 vdd.n2198 gnd 0.00609f
C3928 vdd.n2199 gnd 0.00609f
C3929 vdd.n2200 gnd 0.00609f
C3930 vdd.n2201 gnd 0.00609f
C3931 vdd.n2202 gnd 0.00609f
C3932 vdd.n2203 gnd 0.00609f
C3933 vdd.n2204 gnd 0.00609f
C3934 vdd.n2205 gnd 0.00609f
C3935 vdd.n2206 gnd 0.00609f
C3936 vdd.n2207 gnd 0.00609f
C3937 vdd.n2208 gnd 0.00609f
C3938 vdd.n2209 gnd 0.00609f
C3939 vdd.n2210 gnd 0.00609f
C3940 vdd.n2211 gnd 0.00609f
C3941 vdd.n2212 gnd 0.00609f
C3942 vdd.n2213 gnd 0.00609f
C3943 vdd.n2214 gnd 0.00609f
C3944 vdd.n2215 gnd 0.00609f
C3945 vdd.n2216 gnd 0.00609f
C3946 vdd.n2217 gnd 0.00609f
C3947 vdd.n2218 gnd 10.8083f
C3948 vdd.n2220 gnd 0.013827f
C3949 vdd.n2221 gnd 0.013827f
C3950 vdd.n2222 gnd 0.013039f
C3951 vdd.n2223 gnd 0.00609f
C3952 vdd.n2224 gnd 0.00609f
C3953 vdd.n2225 gnd 0.622324f
C3954 vdd.n2226 gnd 0.00609f
C3955 vdd.n2227 gnd 0.00609f
C3956 vdd.n2228 gnd 0.00609f
C3957 vdd.n2229 gnd 0.00609f
C3958 vdd.n2230 gnd 0.00609f
C3959 vdd.n2231 gnd 0.489623f
C3960 vdd.n2232 gnd 0.00609f
C3961 vdd.n2233 gnd 0.00609f
C3962 vdd.n2234 gnd 0.00609f
C3963 vdd.n2235 gnd 0.00609f
C3964 vdd.n2236 gnd 0.00609f
C3965 vdd.n2237 gnd 0.622324f
C3966 vdd.n2238 gnd 0.00609f
C3967 vdd.n2239 gnd 0.00609f
C3968 vdd.n2240 gnd 0.00609f
C3969 vdd.n2241 gnd 0.00609f
C3970 vdd.n2242 gnd 0.00609f
C3971 vdd.n2243 gnd 0.622324f
C3972 vdd.n2244 gnd 0.00609f
C3973 vdd.n2245 gnd 0.00609f
C3974 vdd.n2246 gnd 0.00609f
C3975 vdd.n2247 gnd 0.00609f
C3976 vdd.n2248 gnd 0.00609f
C3977 vdd.n2249 gnd 0.599445f
C3978 vdd.n2250 gnd 0.00609f
C3979 vdd.n2251 gnd 0.00609f
C3980 vdd.n2252 gnd 0.00609f
C3981 vdd.n2253 gnd 0.00609f
C3982 vdd.n2254 gnd 0.00609f
C3983 vdd.n2255 gnd 0.462167f
C3984 vdd.n2256 gnd 0.00609f
C3985 vdd.n2257 gnd 0.00609f
C3986 vdd.n2258 gnd 0.00609f
C3987 vdd.n2259 gnd 0.00609f
C3988 vdd.n2260 gnd 0.00609f
C3989 vdd.n2261 gnd 0.32489f
C3990 vdd.n2262 gnd 0.00609f
C3991 vdd.n2263 gnd 0.00609f
C3992 vdd.n2264 gnd 0.00609f
C3993 vdd.n2265 gnd 0.00609f
C3994 vdd.n2266 gnd 0.00609f
C3995 vdd.n2267 gnd 0.434712f
C3996 vdd.n2268 gnd 0.00609f
C3997 vdd.n2269 gnd 0.00609f
C3998 vdd.n2270 gnd 0.00609f
C3999 vdd.n2271 gnd 0.00609f
C4000 vdd.n2272 gnd 0.00609f
C4001 vdd.n2273 gnd 0.571989f
C4002 vdd.n2274 gnd 0.00609f
C4003 vdd.n2275 gnd 0.00609f
C4004 vdd.n2276 gnd 0.00609f
C4005 vdd.n2277 gnd 0.00609f
C4006 vdd.n2278 gnd 0.00609f
C4007 vdd.n2279 gnd 0.622324f
C4008 vdd.n2280 gnd 0.00609f
C4009 vdd.n2281 gnd 0.00609f
C4010 vdd.n2282 gnd 0.00609f
C4011 vdd.n2283 gnd 0.00609f
C4012 vdd.n2284 gnd 0.00609f
C4013 vdd.n2285 gnd 0.535382f
C4014 vdd.n2286 gnd 0.00609f
C4015 vdd.n2287 gnd 0.00609f
C4016 vdd.n2288 gnd 0.004836f
C4017 vdd.n2289 gnd 0.017641f
C4018 vdd.n2290 gnd 0.004299f
C4019 vdd.n2291 gnd 0.00609f
C4020 vdd.n2292 gnd 0.398104f
C4021 vdd.n2293 gnd 0.00609f
C4022 vdd.n2294 gnd 0.00609f
C4023 vdd.n2295 gnd 0.00609f
C4024 vdd.n2296 gnd 0.00609f
C4025 vdd.n2297 gnd 0.00609f
C4026 vdd.n2298 gnd 0.361497f
C4027 vdd.n2299 gnd 0.00609f
C4028 vdd.n2300 gnd 0.00609f
C4029 vdd.n2301 gnd 0.00609f
C4030 vdd.n2302 gnd 0.00609f
C4031 vdd.n2303 gnd 0.00609f
C4032 vdd.n2304 gnd 0.498775f
C4033 vdd.n2305 gnd 0.00609f
C4034 vdd.n2306 gnd 0.00609f
C4035 vdd.n2307 gnd 0.00609f
C4036 vdd.n2308 gnd 0.00609f
C4037 vdd.n2309 gnd 0.00609f
C4038 vdd.n2310 gnd 0.54911f
C4039 vdd.n2311 gnd 0.00609f
C4040 vdd.n2312 gnd 0.00609f
C4041 vdd.n2313 gnd 0.00609f
C4042 vdd.n2314 gnd 0.00609f
C4043 vdd.n2315 gnd 0.00609f
C4044 vdd.n2316 gnd 0.411832f
C4045 vdd.n2317 gnd 0.00609f
C4046 vdd.n2318 gnd 0.00609f
C4047 vdd.n2319 gnd 0.00609f
C4048 vdd.n2320 gnd 0.00609f
C4049 vdd.n2321 gnd 0.00609f
C4050 vdd.n2322 gnd 0.196764f
C4051 vdd.n2323 gnd 0.00609f
C4052 vdd.n2324 gnd 0.00609f
C4053 vdd.n2325 gnd 0.00609f
C4054 vdd.n2326 gnd 0.00609f
C4055 vdd.n2327 gnd 0.00609f
C4056 vdd.n2328 gnd 0.196764f
C4057 vdd.n2329 gnd 0.00609f
C4058 vdd.n2330 gnd 0.00609f
C4059 vdd.n2331 gnd 0.00609f
C4060 vdd.n2332 gnd 0.00609f
C4061 vdd.n2333 gnd 0.00609f
C4062 vdd.n2334 gnd 0.622324f
C4063 vdd.n2335 gnd 0.00609f
C4064 vdd.n2336 gnd 0.00609f
C4065 vdd.n2337 gnd 0.00609f
C4066 vdd.n2338 gnd 0.00609f
C4067 vdd.n2339 gnd 0.00609f
C4068 vdd.n2340 gnd 0.00609f
C4069 vdd.n2341 gnd 0.00609f
C4070 vdd.n2342 gnd 0.430136f
C4071 vdd.n2343 gnd 0.00609f
C4072 vdd.n2344 gnd 0.00609f
C4073 vdd.n2345 gnd 0.00609f
C4074 vdd.n2346 gnd 0.00609f
C4075 vdd.n2347 gnd 0.00609f
C4076 vdd.n2348 gnd 0.00609f
C4077 vdd.n2349 gnd 0.388953f
C4078 vdd.n2350 gnd 0.00609f
C4079 vdd.n2351 gnd 0.00609f
C4080 vdd.n2352 gnd 0.00609f
C4081 vdd.n2353 gnd 0.013827f
C4082 vdd.n2354 gnd 0.013039f
C4083 vdd.n2355 gnd 0.00609f
C4084 vdd.n2356 gnd 0.00609f
C4085 vdd.n2357 gnd 0.004701f
C4086 vdd.n2358 gnd 0.00609f
C4087 vdd.n2359 gnd 0.00609f
C4088 vdd.n2360 gnd 0.004433f
C4089 vdd.n2361 gnd 0.00609f
C4090 vdd.n2362 gnd 0.00609f
C4091 vdd.n2363 gnd 0.00609f
C4092 vdd.n2364 gnd 0.00609f
C4093 vdd.n2365 gnd 0.00609f
C4094 vdd.n2366 gnd 0.00609f
C4095 vdd.n2367 gnd 0.00609f
C4096 vdd.n2368 gnd 0.00609f
C4097 vdd.n2369 gnd 0.00609f
C4098 vdd.n2370 gnd 0.00609f
C4099 vdd.n2371 gnd 0.00609f
C4100 vdd.n2372 gnd 0.00609f
C4101 vdd.n2373 gnd 0.00609f
C4102 vdd.n2374 gnd 0.00609f
C4103 vdd.n2375 gnd 0.00609f
C4104 vdd.n2376 gnd 0.00609f
C4105 vdd.n2377 gnd 0.00609f
C4106 vdd.n2378 gnd 0.00609f
C4107 vdd.n2379 gnd 0.00609f
C4108 vdd.n2380 gnd 0.00609f
C4109 vdd.n2381 gnd 0.00609f
C4110 vdd.n2382 gnd 0.00609f
C4111 vdd.n2383 gnd 0.00609f
C4112 vdd.n2384 gnd 0.00609f
C4113 vdd.n2385 gnd 0.00609f
C4114 vdd.n2386 gnd 0.00609f
C4115 vdd.n2387 gnd 0.00609f
C4116 vdd.n2388 gnd 0.00609f
C4117 vdd.n2389 gnd 0.00609f
C4118 vdd.n2390 gnd 0.00609f
C4119 vdd.n2391 gnd 0.00609f
C4120 vdd.n2392 gnd 0.00609f
C4121 vdd.n2393 gnd 0.00609f
C4122 vdd.n2394 gnd 0.00609f
C4123 vdd.n2395 gnd 0.00609f
C4124 vdd.n2396 gnd 0.00609f
C4125 vdd.n2397 gnd 0.00609f
C4126 vdd.n2398 gnd 0.00609f
C4127 vdd.n2399 gnd 0.00609f
C4128 vdd.n2400 gnd 0.00609f
C4129 vdd.n2401 gnd 0.00609f
C4130 vdd.n2402 gnd 0.00609f
C4131 vdd.n2403 gnd 0.00609f
C4132 vdd.n2404 gnd 0.00609f
C4133 vdd.n2405 gnd 0.00609f
C4134 vdd.n2406 gnd 0.00609f
C4135 vdd.n2407 gnd 0.00609f
C4136 vdd.n2408 gnd 0.00609f
C4137 vdd.n2409 gnd 0.00609f
C4138 vdd.n2410 gnd 0.00609f
C4139 vdd.n2411 gnd 0.00609f
C4140 vdd.n2412 gnd 0.00609f
C4141 vdd.n2413 gnd 0.00609f
C4142 vdd.n2414 gnd 0.00609f
C4143 vdd.n2415 gnd 0.00609f
C4144 vdd.n2416 gnd 0.00609f
C4145 vdd.n2417 gnd 0.00609f
C4146 vdd.n2418 gnd 0.00609f
C4147 vdd.n2419 gnd 0.00609f
C4148 vdd.n2420 gnd 0.00609f
C4149 vdd.n2421 gnd 0.013827f
C4150 vdd.n2422 gnd 0.013039f
C4151 vdd.n2423 gnd 0.013039f
C4152 vdd.n2424 gnd 0.704691f
C4153 vdd.n2425 gnd 0.013039f
C4154 vdd.n2426 gnd 0.013827f
C4155 vdd.n2427 gnd 0.013039f
C4156 vdd.n2428 gnd 0.00609f
C4157 vdd.n2429 gnd 0.00609f
C4158 vdd.n2430 gnd 0.00609f
C4159 vdd.n2431 gnd 0.004701f
C4160 vdd.n2432 gnd 0.008703f
C4161 vdd.n2433 gnd 0.004433f
C4162 vdd.n2434 gnd 0.00609f
C4163 vdd.n2435 gnd 0.00609f
C4164 vdd.n2436 gnd 0.00609f
C4165 vdd.n2437 gnd 0.00609f
C4166 vdd.n2438 gnd 0.00609f
C4167 vdd.n2439 gnd 0.00609f
C4168 vdd.n2440 gnd 0.00609f
C4169 vdd.n2441 gnd 0.00609f
C4170 vdd.n2442 gnd 0.00609f
C4171 vdd.n2443 gnd 0.00609f
C4172 vdd.n2444 gnd 0.00609f
C4173 vdd.n2445 gnd 0.00609f
C4174 vdd.n2446 gnd 0.00609f
C4175 vdd.n2447 gnd 0.00609f
C4176 vdd.n2448 gnd 0.00609f
C4177 vdd.n2449 gnd 0.00609f
C4178 vdd.n2450 gnd 0.00609f
C4179 vdd.n2451 gnd 0.00609f
C4180 vdd.n2452 gnd 0.00609f
C4181 vdd.n2453 gnd 0.00609f
C4182 vdd.n2454 gnd 0.00609f
C4183 vdd.n2455 gnd 0.00609f
C4184 vdd.n2456 gnd 0.00609f
C4185 vdd.n2457 gnd 0.00609f
C4186 vdd.n2458 gnd 0.00609f
C4187 vdd.n2459 gnd 0.00609f
C4188 vdd.n2460 gnd 0.00609f
C4189 vdd.n2461 gnd 0.00609f
C4190 vdd.n2462 gnd 0.00609f
C4191 vdd.n2463 gnd 0.00609f
C4192 vdd.n2464 gnd 0.00609f
C4193 vdd.n2465 gnd 0.00609f
C4194 vdd.n2466 gnd 0.00609f
C4195 vdd.n2467 gnd 0.00609f
C4196 vdd.n2468 gnd 0.00609f
C4197 vdd.n2469 gnd 0.00609f
C4198 vdd.n2470 gnd 0.00609f
C4199 vdd.n2471 gnd 0.00609f
C4200 vdd.n2472 gnd 0.00609f
C4201 vdd.n2473 gnd 0.00609f
C4202 vdd.n2474 gnd 0.00609f
C4203 vdd.n2475 gnd 0.00609f
C4204 vdd.n2476 gnd 0.00609f
C4205 vdd.n2477 gnd 0.00609f
C4206 vdd.n2478 gnd 0.00609f
C4207 vdd.n2479 gnd 0.00609f
C4208 vdd.n2480 gnd 0.00609f
C4209 vdd.n2481 gnd 0.00609f
C4210 vdd.n2482 gnd 0.00609f
C4211 vdd.n2483 gnd 0.00609f
C4212 vdd.n2484 gnd 0.00609f
C4213 vdd.n2485 gnd 0.00609f
C4214 vdd.n2486 gnd 0.00609f
C4215 vdd.n2487 gnd 0.00609f
C4216 vdd.n2488 gnd 0.00609f
C4217 vdd.n2489 gnd 0.00609f
C4218 vdd.n2490 gnd 0.00609f
C4219 vdd.n2491 gnd 0.00609f
C4220 vdd.n2492 gnd 0.00609f
C4221 vdd.n2493 gnd 0.00609f
C4222 vdd.n2494 gnd 0.013827f
C4223 vdd.n2495 gnd 0.013827f
C4224 vdd.n2496 gnd 0.759602f
C4225 vdd.t188 gnd 2.69979f
C4226 vdd.t164 gnd 2.69979f
C4227 vdd.n2530 gnd 0.013827f
C4228 vdd.t193 gnd 0.530806f
C4229 vdd.n2531 gnd 0.00609f
C4230 vdd.t82 gnd 0.246078f
C4231 vdd.t83 gnd 0.251892f
C4232 vdd.t80 gnd 0.160649f
C4233 vdd.n2532 gnd 0.086822f
C4234 vdd.n2533 gnd 0.049248f
C4235 vdd.n2534 gnd 0.00609f
C4236 vdd.t92 gnd 0.246078f
C4237 vdd.t93 gnd 0.251892f
C4238 vdd.t91 gnd 0.160649f
C4239 vdd.n2535 gnd 0.086822f
C4240 vdd.n2536 gnd 0.049248f
C4241 vdd.n2537 gnd 0.008703f
C4242 vdd.n2538 gnd 0.013827f
C4243 vdd.n2539 gnd 0.013827f
C4244 vdd.n2540 gnd 0.00609f
C4245 vdd.n2541 gnd 0.00609f
C4246 vdd.n2542 gnd 0.00609f
C4247 vdd.n2543 gnd 0.00609f
C4248 vdd.n2544 gnd 0.00609f
C4249 vdd.n2545 gnd 0.00609f
C4250 vdd.n2546 gnd 0.00609f
C4251 vdd.n2547 gnd 0.00609f
C4252 vdd.n2548 gnd 0.00609f
C4253 vdd.n2549 gnd 0.00609f
C4254 vdd.n2550 gnd 0.00609f
C4255 vdd.n2551 gnd 0.00609f
C4256 vdd.n2552 gnd 0.00609f
C4257 vdd.n2553 gnd 0.00609f
C4258 vdd.n2554 gnd 0.00609f
C4259 vdd.n2555 gnd 0.00609f
C4260 vdd.n2556 gnd 0.00609f
C4261 vdd.n2557 gnd 0.00609f
C4262 vdd.n2558 gnd 0.00609f
C4263 vdd.n2559 gnd 0.00609f
C4264 vdd.n2560 gnd 0.00609f
C4265 vdd.n2561 gnd 0.00609f
C4266 vdd.n2562 gnd 0.00609f
C4267 vdd.n2563 gnd 0.00609f
C4268 vdd.n2564 gnd 0.00609f
C4269 vdd.n2565 gnd 0.00609f
C4270 vdd.n2566 gnd 0.00609f
C4271 vdd.n2567 gnd 0.00609f
C4272 vdd.n2568 gnd 0.00609f
C4273 vdd.n2569 gnd 0.00609f
C4274 vdd.n2570 gnd 0.00609f
C4275 vdd.n2571 gnd 0.00609f
C4276 vdd.n2572 gnd 0.00609f
C4277 vdd.n2573 gnd 0.00609f
C4278 vdd.n2574 gnd 0.00609f
C4279 vdd.n2575 gnd 0.00609f
C4280 vdd.n2576 gnd 0.00609f
C4281 vdd.n2577 gnd 0.00609f
C4282 vdd.n2578 gnd 0.00609f
C4283 vdd.n2579 gnd 0.00609f
C4284 vdd.n2580 gnd 0.00609f
C4285 vdd.n2581 gnd 0.00609f
C4286 vdd.n2582 gnd 0.00609f
C4287 vdd.n2583 gnd 0.00609f
C4288 vdd.n2584 gnd 0.00609f
C4289 vdd.n2585 gnd 0.00609f
C4290 vdd.n2586 gnd 0.00609f
C4291 vdd.n2587 gnd 0.00609f
C4292 vdd.n2588 gnd 0.00609f
C4293 vdd.n2589 gnd 0.00609f
C4294 vdd.n2590 gnd 0.00609f
C4295 vdd.n2591 gnd 0.00609f
C4296 vdd.n2592 gnd 0.00609f
C4297 vdd.n2593 gnd 0.00609f
C4298 vdd.n2594 gnd 0.00609f
C4299 vdd.n2595 gnd 0.00609f
C4300 vdd.n2596 gnd 0.00609f
C4301 vdd.n2597 gnd 0.00609f
C4302 vdd.n2598 gnd 0.00609f
C4303 vdd.n2599 gnd 0.00609f
C4304 vdd.n2600 gnd 0.004433f
C4305 vdd.n2601 gnd 0.00609f
C4306 vdd.n2602 gnd 0.00609f
C4307 vdd.n2603 gnd 0.004701f
C4308 vdd.n2604 gnd 0.00609f
C4309 vdd.n2605 gnd 0.00609f
C4310 vdd.n2606 gnd 0.013827f
C4311 vdd.n2607 gnd 0.013039f
C4312 vdd.n2608 gnd 0.013039f
C4313 vdd.n2609 gnd 0.00609f
C4314 vdd.n2610 gnd 0.00609f
C4315 vdd.n2611 gnd 0.00609f
C4316 vdd.n2612 gnd 0.00609f
C4317 vdd.n2613 gnd 0.00609f
C4318 vdd.n2614 gnd 0.00609f
C4319 vdd.n2615 gnd 0.00609f
C4320 vdd.n2616 gnd 0.00609f
C4321 vdd.n2617 gnd 0.00609f
C4322 vdd.n2618 gnd 0.00609f
C4323 vdd.n2619 gnd 0.00609f
C4324 vdd.n2620 gnd 0.00609f
C4325 vdd.n2621 gnd 0.00609f
C4326 vdd.n2622 gnd 0.00609f
C4327 vdd.n2623 gnd 0.00609f
C4328 vdd.n2624 gnd 0.00609f
C4329 vdd.n2625 gnd 0.00609f
C4330 vdd.n2626 gnd 0.00609f
C4331 vdd.n2627 gnd 0.00609f
C4332 vdd.n2628 gnd 0.00609f
C4333 vdd.n2629 gnd 0.00609f
C4334 vdd.n2630 gnd 0.00609f
C4335 vdd.n2631 gnd 0.00609f
C4336 vdd.n2632 gnd 0.00609f
C4337 vdd.n2633 gnd 0.00609f
C4338 vdd.n2634 gnd 0.00609f
C4339 vdd.n2635 gnd 0.00609f
C4340 vdd.n2636 gnd 0.00609f
C4341 vdd.n2637 gnd 0.00609f
C4342 vdd.n2638 gnd 0.00609f
C4343 vdd.n2639 gnd 0.00609f
C4344 vdd.n2640 gnd 0.00609f
C4345 vdd.n2641 gnd 0.00609f
C4346 vdd.n2642 gnd 0.00609f
C4347 vdd.n2643 gnd 0.00609f
C4348 vdd.n2644 gnd 0.00609f
C4349 vdd.n2645 gnd 0.00609f
C4350 vdd.n2646 gnd 0.00609f
C4351 vdd.n2647 gnd 0.00609f
C4352 vdd.n2648 gnd 0.00609f
C4353 vdd.n2649 gnd 0.00609f
C4354 vdd.n2650 gnd 0.00609f
C4355 vdd.n2651 gnd 0.00609f
C4356 vdd.n2652 gnd 0.00609f
C4357 vdd.n2653 gnd 0.00609f
C4358 vdd.n2654 gnd 0.00609f
C4359 vdd.n2655 gnd 0.00609f
C4360 vdd.n2656 gnd 0.00609f
C4361 vdd.n2657 gnd 0.00609f
C4362 vdd.n2658 gnd 0.00609f
C4363 vdd.n2659 gnd 0.00609f
C4364 vdd.n2660 gnd 0.00609f
C4365 vdd.n2661 gnd 0.00609f
C4366 vdd.n2662 gnd 0.00609f
C4367 vdd.n2663 gnd 0.00609f
C4368 vdd.n2664 gnd 0.00609f
C4369 vdd.n2665 gnd 0.00609f
C4370 vdd.n2666 gnd 0.00609f
C4371 vdd.n2667 gnd 0.00609f
C4372 vdd.n2668 gnd 0.00609f
C4373 vdd.n2669 gnd 0.00609f
C4374 vdd.n2670 gnd 0.00609f
C4375 vdd.n2671 gnd 0.00609f
C4376 vdd.n2672 gnd 0.00609f
C4377 vdd.n2673 gnd 0.00609f
C4378 vdd.n2674 gnd 0.00609f
C4379 vdd.n2675 gnd 0.00609f
C4380 vdd.n2676 gnd 0.00609f
C4381 vdd.n2677 gnd 0.00609f
C4382 vdd.n2678 gnd 0.00609f
C4383 vdd.n2679 gnd 0.00609f
C4384 vdd.n2680 gnd 0.00609f
C4385 vdd.n2681 gnd 0.00609f
C4386 vdd.n2682 gnd 0.00609f
C4387 vdd.n2683 gnd 0.00609f
C4388 vdd.n2684 gnd 0.00609f
C4389 vdd.n2685 gnd 0.00609f
C4390 vdd.n2686 gnd 0.00609f
C4391 vdd.n2687 gnd 0.00609f
C4392 vdd.n2688 gnd 0.00609f
C4393 vdd.n2689 gnd 0.00609f
C4394 vdd.n2690 gnd 0.00609f
C4395 vdd.n2691 gnd 0.00609f
C4396 vdd.n2692 gnd 0.00609f
C4397 vdd.n2693 gnd 0.00609f
C4398 vdd.n2694 gnd 0.00609f
C4399 vdd.n2695 gnd 0.00609f
C4400 vdd.n2696 gnd 0.00609f
C4401 vdd.n2697 gnd 0.00609f
C4402 vdd.n2698 gnd 0.00609f
C4403 vdd.n2699 gnd 0.00609f
C4404 vdd.n2700 gnd 0.00609f
C4405 vdd.n2701 gnd 0.00609f
C4406 vdd.n2702 gnd 0.00609f
C4407 vdd.n2703 gnd 0.00609f
C4408 vdd.n2704 gnd 0.00609f
C4409 vdd.n2705 gnd 0.00609f
C4410 vdd.n2706 gnd 0.00609f
C4411 vdd.n2707 gnd 0.00609f
C4412 vdd.n2708 gnd 0.00609f
C4413 vdd.n2709 gnd 0.00609f
C4414 vdd.n2710 gnd 0.196764f
C4415 vdd.n2711 gnd 0.00609f
C4416 vdd.n2712 gnd 0.00609f
C4417 vdd.n2713 gnd 0.00609f
C4418 vdd.n2714 gnd 0.00609f
C4419 vdd.n2715 gnd 0.00609f
C4420 vdd.n2716 gnd 0.196764f
C4421 vdd.n2717 gnd 0.00609f
C4422 vdd.n2718 gnd 0.00609f
C4423 vdd.n2719 gnd 0.00609f
C4424 vdd.n2720 gnd 0.00609f
C4425 vdd.n2721 gnd 0.00609f
C4426 vdd.n2722 gnd 0.00609f
C4427 vdd.n2723 gnd 0.00609f
C4428 vdd.n2724 gnd 0.00609f
C4429 vdd.n2725 gnd 0.00609f
C4430 vdd.n2726 gnd 0.00609f
C4431 vdd.n2727 gnd 0.00609f
C4432 vdd.n2728 gnd 0.388953f
C4433 vdd.n2729 gnd 0.00609f
C4434 vdd.n2730 gnd 0.00609f
C4435 vdd.n2731 gnd 0.00609f
C4436 vdd.n2732 gnd 0.013039f
C4437 vdd.n2733 gnd 0.013039f
C4438 vdd.n2734 gnd 0.013827f
C4439 vdd.n2735 gnd 0.013827f
C4440 vdd.n2736 gnd 0.00609f
C4441 vdd.n2737 gnd 0.00609f
C4442 vdd.n2738 gnd 0.00609f
C4443 vdd.n2739 gnd 0.004701f
C4444 vdd.n2740 gnd 0.008703f
C4445 vdd.n2741 gnd 0.004433f
C4446 vdd.n2742 gnd 0.00609f
C4447 vdd.n2743 gnd 0.00609f
C4448 vdd.n2744 gnd 0.00609f
C4449 vdd.n2745 gnd 0.00609f
C4450 vdd.n2746 gnd 0.00609f
C4451 vdd.n2747 gnd 0.00609f
C4452 vdd.n2748 gnd 0.00609f
C4453 vdd.n2749 gnd 0.00609f
C4454 vdd.n2750 gnd 0.00609f
C4455 vdd.n2751 gnd 0.00609f
C4456 vdd.n2752 gnd 0.00609f
C4457 vdd.n2753 gnd 0.00609f
C4458 vdd.n2754 gnd 0.00609f
C4459 vdd.n2755 gnd 0.00609f
C4460 vdd.n2756 gnd 0.00609f
C4461 vdd.n2757 gnd 0.00609f
C4462 vdd.n2758 gnd 0.00609f
C4463 vdd.n2759 gnd 0.00609f
C4464 vdd.n2760 gnd 0.00609f
C4465 vdd.n2761 gnd 0.00609f
C4466 vdd.n2762 gnd 0.00609f
C4467 vdd.n2763 gnd 0.00609f
C4468 vdd.n2764 gnd 0.00609f
C4469 vdd.n2765 gnd 0.00609f
C4470 vdd.n2766 gnd 0.00609f
C4471 vdd.n2767 gnd 0.00609f
C4472 vdd.n2768 gnd 0.00609f
C4473 vdd.n2769 gnd 0.00609f
C4474 vdd.n2770 gnd 0.00609f
C4475 vdd.n2771 gnd 0.00609f
C4476 vdd.n2772 gnd 0.00609f
C4477 vdd.n2773 gnd 0.00609f
C4478 vdd.n2774 gnd 0.00609f
C4479 vdd.n2775 gnd 0.00609f
C4480 vdd.n2776 gnd 0.00609f
C4481 vdd.n2777 gnd 0.00609f
C4482 vdd.n2778 gnd 0.00609f
C4483 vdd.n2779 gnd 0.00609f
C4484 vdd.n2780 gnd 0.00609f
C4485 vdd.n2781 gnd 0.00609f
C4486 vdd.n2782 gnd 0.00609f
C4487 vdd.n2783 gnd 0.00609f
C4488 vdd.n2784 gnd 0.00609f
C4489 vdd.n2785 gnd 0.00609f
C4490 vdd.n2786 gnd 0.00609f
C4491 vdd.n2787 gnd 0.00609f
C4492 vdd.n2788 gnd 0.00609f
C4493 vdd.n2789 gnd 0.00609f
C4494 vdd.n2790 gnd 0.00609f
C4495 vdd.n2791 gnd 0.00609f
C4496 vdd.n2792 gnd 0.00609f
C4497 vdd.n2793 gnd 0.00609f
C4498 vdd.n2794 gnd 0.00609f
C4499 vdd.n2795 gnd 0.00609f
C4500 vdd.n2796 gnd 0.00609f
C4501 vdd.n2797 gnd 0.00609f
C4502 vdd.n2798 gnd 0.00609f
C4503 vdd.n2799 gnd 0.00609f
C4504 vdd.n2800 gnd 0.759602f
C4505 vdd.n2802 gnd 0.013827f
C4506 vdd.n2803 gnd 0.013827f
C4507 vdd.n2804 gnd 0.013039f
C4508 vdd.n2805 gnd 0.00609f
C4509 vdd.n2806 gnd 0.00609f
C4510 vdd.n2807 gnd 0.366073f
C4511 vdd.n2808 gnd 0.00609f
C4512 vdd.n2809 gnd 0.00609f
C4513 vdd.n2810 gnd 0.00609f
C4514 vdd.n2811 gnd 0.00609f
C4515 vdd.n2812 gnd 0.00609f
C4516 vdd.n2813 gnd 0.370649f
C4517 vdd.n2814 gnd 0.00609f
C4518 vdd.n2815 gnd 0.00609f
C4519 vdd.n2816 gnd 0.00609f
C4520 vdd.n2817 gnd 0.00609f
C4521 vdd.n2818 gnd 0.00609f
C4522 vdd.n2819 gnd 0.622324f
C4523 vdd.n2820 gnd 0.00609f
C4524 vdd.n2821 gnd 0.00609f
C4525 vdd.n2822 gnd 0.00609f
C4526 vdd.n2823 gnd 0.00609f
C4527 vdd.n2824 gnd 0.00609f
C4528 vdd.n2825 gnd 0.448439f
C4529 vdd.n2826 gnd 0.00609f
C4530 vdd.n2827 gnd 0.00609f
C4531 vdd.n2828 gnd 0.00609f
C4532 vdd.n2829 gnd 0.00609f
C4533 vdd.n2830 gnd 0.00609f
C4534 vdd.n2831 gnd 0.562837f
C4535 vdd.n2832 gnd 0.00609f
C4536 vdd.n2833 gnd 0.00609f
C4537 vdd.n2834 gnd 0.00609f
C4538 vdd.n2835 gnd 0.00609f
C4539 vdd.n2836 gnd 0.00609f
C4540 vdd.n2837 gnd 0.462167f
C4541 vdd.n2838 gnd 0.00609f
C4542 vdd.n2839 gnd 0.00609f
C4543 vdd.n2840 gnd 0.00609f
C4544 vdd.n2841 gnd 0.00609f
C4545 vdd.n2842 gnd 0.00609f
C4546 vdd.n2843 gnd 0.32489f
C4547 vdd.n2844 gnd 0.00609f
C4548 vdd.n2845 gnd 0.00609f
C4549 vdd.n2846 gnd 0.00609f
C4550 vdd.n2847 gnd 0.00609f
C4551 vdd.n2848 gnd 0.00609f
C4552 vdd.n2849 gnd 0.196764f
C4553 vdd.n2850 gnd 0.00609f
C4554 vdd.n2851 gnd 0.00609f
C4555 vdd.n2852 gnd 0.00609f
C4556 vdd.n2853 gnd 0.00609f
C4557 vdd.n2854 gnd 0.00609f
C4558 vdd.n2855 gnd 0.571989f
C4559 vdd.n2856 gnd 0.00609f
C4560 vdd.n2857 gnd 0.00609f
C4561 vdd.n2858 gnd 0.00609f
C4562 vdd.n2859 gnd 0.004299f
C4563 vdd.n2860 gnd 0.00609f
C4564 vdd.n2861 gnd 0.00609f
C4565 vdd.n2862 gnd 0.622324f
C4566 vdd.n2863 gnd 0.00609f
C4567 vdd.n2864 gnd 0.00609f
C4568 vdd.n2865 gnd 0.00609f
C4569 vdd.n2866 gnd 0.00609f
C4570 vdd.n2867 gnd 0.00609f
C4571 vdd.n2868 gnd 0.494199f
C4572 vdd.n2869 gnd 0.00609f
C4573 vdd.n2870 gnd 0.004836f
C4574 vdd.n2871 gnd 0.00609f
C4575 vdd.n2872 gnd 0.00609f
C4576 vdd.n2873 gnd 0.00609f
C4577 vdd.n2874 gnd 0.398104f
C4578 vdd.n2875 gnd 0.00609f
C4579 vdd.n2876 gnd 0.00609f
C4580 vdd.n2877 gnd 0.00609f
C4581 vdd.n2878 gnd 0.00609f
C4582 vdd.n2879 gnd 0.00609f
C4583 vdd.n2880 gnd 0.361497f
C4584 vdd.n2881 gnd 0.00609f
C4585 vdd.n2882 gnd 0.00609f
C4586 vdd.n2883 gnd 0.00609f
C4587 vdd.n2884 gnd 0.00609f
C4588 vdd.n2885 gnd 0.00609f
C4589 vdd.n2886 gnd 0.498775f
C4590 vdd.n2887 gnd 0.00609f
C4591 vdd.n2888 gnd 0.00609f
C4592 vdd.n2889 gnd 0.00609f
C4593 vdd.n2890 gnd 0.00609f
C4594 vdd.n2891 gnd 0.00609f
C4595 vdd.n2892 gnd 0.622324f
C4596 vdd.n2893 gnd 0.00609f
C4597 vdd.n2894 gnd 0.00609f
C4598 vdd.n2895 gnd 0.00609f
C4599 vdd.n2896 gnd 0.00609f
C4600 vdd.n2897 gnd 0.00609f
C4601 vdd.n2898 gnd 0.608596f
C4602 vdd.n2899 gnd 0.00609f
C4603 vdd.n2900 gnd 0.00609f
C4604 vdd.n2901 gnd 0.00609f
C4605 vdd.n2902 gnd 0.00609f
C4606 vdd.n2903 gnd 0.00609f
C4607 vdd.n2904 gnd 0.471319f
C4608 vdd.n2905 gnd 0.00609f
C4609 vdd.n2906 gnd 0.00609f
C4610 vdd.n2907 gnd 0.00609f
C4611 vdd.n2908 gnd 0.00609f
C4612 vdd.n2909 gnd 0.00609f
C4613 vdd.n2910 gnd 0.334042f
C4614 vdd.n2911 gnd 0.00609f
C4615 vdd.n2912 gnd 0.00609f
C4616 vdd.n2913 gnd 0.00609f
C4617 vdd.n2914 gnd 0.00609f
C4618 vdd.n2915 gnd 0.00609f
C4619 vdd.n2916 gnd 0.622324f
C4620 vdd.n2917 gnd 0.00609f
C4621 vdd.n2918 gnd 0.00609f
C4622 vdd.n2919 gnd 0.00609f
C4623 vdd.n2920 gnd 0.00609f
C4624 vdd.n2921 gnd 0.00609f
C4625 vdd.n2922 gnd 0.00609f
C4626 vdd.n2924 gnd 0.00609f
C4627 vdd.n2925 gnd 0.00609f
C4628 vdd.n2927 gnd 0.00609f
C4629 vdd.n2928 gnd 0.00609f
C4630 vdd.n2931 gnd 0.00609f
C4631 vdd.n2932 gnd 0.00609f
C4632 vdd.n2933 gnd 0.00609f
C4633 vdd.n2934 gnd 0.00609f
C4634 vdd.n2936 gnd 0.00609f
C4635 vdd.n2937 gnd 0.00609f
C4636 vdd.n2938 gnd 0.00609f
C4637 vdd.n2939 gnd 0.00609f
C4638 vdd.n2940 gnd 0.00609f
C4639 vdd.n2941 gnd 0.00609f
C4640 vdd.n2943 gnd 0.00609f
C4641 vdd.n2944 gnd 0.00609f
C4642 vdd.n2945 gnd 0.00609f
C4643 vdd.n2946 gnd 0.00609f
C4644 vdd.n2947 gnd 0.00609f
C4645 vdd.n2948 gnd 0.00609f
C4646 vdd.n2950 gnd 0.00609f
C4647 vdd.n2951 gnd 0.00609f
C4648 vdd.n2952 gnd 0.00609f
C4649 vdd.n2953 gnd 0.00609f
C4650 vdd.n2954 gnd 0.00609f
C4651 vdd.n2955 gnd 0.00609f
C4652 vdd.n2957 gnd 0.00609f
C4653 vdd.n2958 gnd 0.013827f
C4654 vdd.n2959 gnd 0.013827f
C4655 vdd.n2960 gnd 0.013039f
C4656 vdd.n2961 gnd 0.00609f
C4657 vdd.n2962 gnd 0.00609f
C4658 vdd.n2963 gnd 0.00609f
C4659 vdd.n2964 gnd 0.00609f
C4660 vdd.n2965 gnd 0.00609f
C4661 vdd.n2966 gnd 0.00609f
C4662 vdd.n2967 gnd 0.622324f
C4663 vdd.n2968 gnd 0.00609f
C4664 vdd.n2969 gnd 0.00609f
C4665 vdd.n2970 gnd 0.00609f
C4666 vdd.n2971 gnd 0.00609f
C4667 vdd.n2972 gnd 0.00609f
C4668 vdd.n2973 gnd 0.443864f
C4669 vdd.n2974 gnd 0.00609f
C4670 vdd.n2975 gnd 0.00609f
C4671 vdd.n2976 gnd 0.00609f
C4672 vdd.n2977 gnd 0.013827f
C4673 vdd.n2979 gnd 0.013827f
C4674 vdd.n2980 gnd 0.013039f
C4675 vdd.n2981 gnd 0.00609f
C4676 vdd.n2982 gnd 0.004701f
C4677 vdd.n2983 gnd 0.00609f
C4678 vdd.n2985 gnd 0.00609f
C4679 vdd.n2986 gnd 0.00609f
C4680 vdd.n2987 gnd 0.00609f
C4681 vdd.n2988 gnd 0.00609f
C4682 vdd.n2989 gnd 0.00609f
C4683 vdd.n2990 gnd 0.00609f
C4684 vdd.n2992 gnd 0.00609f
C4685 vdd.n2993 gnd 0.00609f
C4686 vdd.n2994 gnd 0.00609f
C4687 vdd.n2995 gnd 0.00609f
C4688 vdd.n2996 gnd 0.00609f
C4689 vdd.n2997 gnd 0.00609f
C4690 vdd.n2999 gnd 0.00609f
C4691 vdd.n3000 gnd 0.00609f
C4692 vdd.n3001 gnd 0.00609f
C4693 vdd.n3002 gnd 0.00609f
C4694 vdd.n3003 gnd 0.00609f
C4695 vdd.n3004 gnd 0.00609f
C4696 vdd.n3006 gnd 0.00609f
C4697 vdd.n3007 gnd 0.00609f
C4698 vdd.n3008 gnd 0.00609f
C4699 vdd.n3009 gnd 0.954111f
C4700 vdd.n3010 gnd 0.037602f
C4701 vdd.n3011 gnd 0.00609f
C4702 vdd.n3012 gnd 0.00609f
C4703 vdd.n3014 gnd 0.00609f
C4704 vdd.n3015 gnd 0.00609f
C4705 vdd.n3016 gnd 0.00609f
C4706 vdd.n3017 gnd 0.00609f
C4707 vdd.n3018 gnd 0.00609f
C4708 vdd.n3019 gnd 0.00609f
C4709 vdd.n3021 gnd 0.00609f
C4710 vdd.n3022 gnd 0.00609f
C4711 vdd.n3023 gnd 0.00609f
C4712 vdd.n3024 gnd 0.00609f
C4713 vdd.n3025 gnd 0.00609f
C4714 vdd.n3026 gnd 0.00609f
C4715 vdd.n3028 gnd 0.00609f
C4716 vdd.n3029 gnd 0.00609f
C4717 vdd.n3030 gnd 0.00609f
C4718 vdd.n3031 gnd 0.00609f
C4719 vdd.n3032 gnd 0.00609f
C4720 vdd.n3033 gnd 0.00609f
C4721 vdd.n3035 gnd 0.00609f
C4722 vdd.n3036 gnd 0.00609f
C4723 vdd.n3038 gnd 0.00609f
C4724 vdd.n3039 gnd 0.00609f
C4725 vdd.n3040 gnd 0.013827f
C4726 vdd.n3041 gnd 0.013039f
C4727 vdd.n3042 gnd 0.013039f
C4728 vdd.n3043 gnd 0.841968f
C4729 vdd.n3044 gnd 0.013039f
C4730 vdd.n3045 gnd 0.013827f
C4731 vdd.n3046 gnd 0.013039f
C4732 vdd.n3047 gnd 0.00609f
C4733 vdd.n3048 gnd 0.004701f
C4734 vdd.n3049 gnd 0.00609f
C4735 vdd.n3051 gnd 0.00609f
C4736 vdd.n3052 gnd 0.00609f
C4737 vdd.n3053 gnd 0.00609f
C4738 vdd.n3054 gnd 0.00609f
C4739 vdd.n3055 gnd 0.00609f
C4740 vdd.n3056 gnd 0.00609f
C4741 vdd.n3058 gnd 0.00609f
C4742 vdd.n3059 gnd 0.00609f
C4743 vdd.n3060 gnd 0.00609f
C4744 vdd.n3061 gnd 0.00609f
C4745 vdd.n3062 gnd 0.00609f
C4746 vdd.n3063 gnd 0.00609f
C4747 vdd.n3065 gnd 0.00609f
C4748 vdd.n3066 gnd 0.00609f
C4749 vdd.n3067 gnd 0.00609f
C4750 vdd.n3068 gnd 0.00609f
C4751 vdd.n3069 gnd 0.00609f
C4752 vdd.n3070 gnd 0.00609f
C4753 vdd.n3072 gnd 0.00609f
C4754 vdd.n3073 gnd 0.00609f
C4755 vdd.n3075 gnd 0.00609f
C4756 vdd.n3076 gnd 0.037602f
C4757 vdd.n3077 gnd 0.954111f
C4758 vdd.n3078 gnd 0.007702f
C4759 vdd.n3079 gnd 0.003424f
C4760 vdd.t44 gnd 0.110173f
C4761 vdd.t45 gnd 0.117745f
C4762 vdd.t42 gnd 0.143884f
C4763 vdd.n3080 gnd 0.184439f
C4764 vdd.n3081 gnd 0.154963f
C4765 vdd.n3082 gnd 0.0111f
C4766 vdd.n3083 gnd 0.008955f
C4767 vdd.n3084 gnd 0.003784f
C4768 vdd.n3085 gnd 0.007208f
C4769 vdd.n3086 gnd 0.008955f
C4770 vdd.n3087 gnd 0.008955f
C4771 vdd.n3088 gnd 0.007208f
C4772 vdd.n3089 gnd 0.007208f
C4773 vdd.n3090 gnd 0.008955f
C4774 vdd.n3092 gnd 0.008955f
C4775 vdd.n3093 gnd 0.007208f
C4776 vdd.n3094 gnd 0.007208f
C4777 vdd.n3095 gnd 0.007208f
C4778 vdd.n3096 gnd 0.008955f
C4779 vdd.n3098 gnd 0.008955f
C4780 vdd.n3100 gnd 0.008955f
C4781 vdd.n3101 gnd 0.007208f
C4782 vdd.n3102 gnd 0.007208f
C4783 vdd.n3103 gnd 0.007208f
C4784 vdd.n3104 gnd 0.008955f
C4785 vdd.n3106 gnd 0.008955f
C4786 vdd.n3108 gnd 0.008955f
C4787 vdd.n3109 gnd 0.007208f
C4788 vdd.n3110 gnd 0.007208f
C4789 vdd.n3111 gnd 0.007208f
C4790 vdd.n3112 gnd 0.008955f
C4791 vdd.n3114 gnd 0.008955f
C4792 vdd.n3115 gnd 0.008955f
C4793 vdd.n3116 gnd 0.007208f
C4794 vdd.n3117 gnd 0.007208f
C4795 vdd.n3118 gnd 0.008955f
C4796 vdd.n3119 gnd 0.008955f
C4797 vdd.n3121 gnd 0.008955f
C4798 vdd.n3122 gnd 0.007208f
C4799 vdd.n3123 gnd 0.008955f
C4800 vdd.n3124 gnd 0.008955f
C4801 vdd.n3125 gnd 0.008955f
C4802 vdd.n3126 gnd 0.014704f
C4803 vdd.n3127 gnd 0.004901f
C4804 vdd.n3128 gnd 0.008955f
C4805 vdd.n3130 gnd 0.008955f
C4806 vdd.n3132 gnd 0.008955f
C4807 vdd.n3133 gnd 0.007208f
C4808 vdd.n3134 gnd 0.007208f
C4809 vdd.n3135 gnd 0.007208f
C4810 vdd.n3136 gnd 0.008955f
C4811 vdd.n3138 gnd 0.008955f
C4812 vdd.n3140 gnd 0.008955f
C4813 vdd.n3141 gnd 0.007208f
C4814 vdd.n3142 gnd 0.007208f
C4815 vdd.n3143 gnd 0.007208f
C4816 vdd.n3144 gnd 0.008955f
C4817 vdd.n3146 gnd 0.008955f
C4818 vdd.n3148 gnd 0.008955f
C4819 vdd.n3149 gnd 0.007208f
C4820 vdd.n3150 gnd 0.007208f
C4821 vdd.n3151 gnd 0.007208f
C4822 vdd.n3152 gnd 0.008955f
C4823 vdd.n3154 gnd 0.008955f
C4824 vdd.n3156 gnd 0.008955f
C4825 vdd.n3157 gnd 0.007208f
C4826 vdd.n3158 gnd 0.007208f
C4827 vdd.n3159 gnd 0.007208f
C4828 vdd.n3160 gnd 0.008955f
C4829 vdd.n3162 gnd 0.008955f
C4830 vdd.n3164 gnd 0.008955f
C4831 vdd.n3165 gnd 0.007208f
C4832 vdd.n3166 gnd 0.007208f
C4833 vdd.n3167 gnd 0.006019f
C4834 vdd.n3168 gnd 0.008955f
C4835 vdd.n3170 gnd 0.008955f
C4836 vdd.n3172 gnd 0.008955f
C4837 vdd.n3173 gnd 0.006019f
C4838 vdd.n3174 gnd 0.007208f
C4839 vdd.n3175 gnd 0.007208f
C4840 vdd.n3176 gnd 0.008955f
C4841 vdd.n3178 gnd 0.008955f
C4842 vdd.n3180 gnd 0.008955f
C4843 vdd.n3181 gnd 0.007208f
C4844 vdd.n3182 gnd 0.007208f
C4845 vdd.n3183 gnd 0.007208f
C4846 vdd.n3184 gnd 0.008955f
C4847 vdd.n3186 gnd 0.008955f
C4848 vdd.n3188 gnd 0.008955f
C4849 vdd.n3189 gnd 0.007208f
C4850 vdd.n3190 gnd 0.007208f
C4851 vdd.n3191 gnd 0.007208f
C4852 vdd.n3192 gnd 0.008955f
C4853 vdd.n3194 gnd 0.008955f
C4854 vdd.n3195 gnd 0.008955f
C4855 vdd.n3196 gnd 0.007208f
C4856 vdd.n3197 gnd 0.007208f
C4857 vdd.n3198 gnd 0.008955f
C4858 vdd.n3199 gnd 0.008955f
C4859 vdd.n3200 gnd 0.007208f
C4860 vdd.n3201 gnd 0.007208f
C4861 vdd.n3202 gnd 0.008955f
C4862 vdd.n3203 gnd 0.008955f
C4863 vdd.n3205 gnd 0.008955f
C4864 vdd.n3206 gnd 0.007208f
C4865 vdd.n3207 gnd 0.005983f
C4866 vdd.n3208 gnd 0.021434f
C4867 vdd.n3209 gnd 0.021104f
C4868 vdd.n3210 gnd 0.005983f
C4869 vdd.n3211 gnd 0.021104f
C4870 vdd.n3212 gnd 1.25838f
C4871 vdd.n3213 gnd 0.021104f
C4872 vdd.n3214 gnd 0.005983f
C4873 vdd.n3215 gnd 0.021104f
C4874 vdd.n3216 gnd 0.008955f
C4875 vdd.n3217 gnd 0.008955f
C4876 vdd.n3218 gnd 0.007208f
C4877 vdd.n3219 gnd 0.008955f
C4878 vdd.n3220 gnd 0.915183f
C4879 vdd.n3221 gnd 0.008955f
C4880 vdd.n3222 gnd 0.007208f
C4881 vdd.n3223 gnd 0.008955f
C4882 vdd.n3224 gnd 0.008955f
C4883 vdd.n3225 gnd 0.008955f
C4884 vdd.n3226 gnd 0.007208f
C4885 vdd.n3227 gnd 0.008955f
C4886 vdd.n3228 gnd 0.809937f
C4887 vdd.n3229 gnd 0.008955f
C4888 vdd.n3230 gnd 0.007208f
C4889 vdd.n3231 gnd 0.008955f
C4890 vdd.n3232 gnd 0.008955f
C4891 vdd.n3233 gnd 0.008955f
C4892 vdd.n3234 gnd 0.007208f
C4893 vdd.n3235 gnd 0.008955f
C4894 vdd.t0 gnd 0.457591f
C4895 vdd.n3236 gnd 0.654356f
C4896 vdd.n3237 gnd 0.008955f
C4897 vdd.n3238 gnd 0.007208f
C4898 vdd.n3239 gnd 0.008955f
C4899 vdd.n3240 gnd 0.008955f
C4900 vdd.n3241 gnd 0.008955f
C4901 vdd.n3242 gnd 0.007208f
C4902 vdd.n3243 gnd 0.008955f
C4903 vdd.n3244 gnd 0.498775f
C4904 vdd.n3245 gnd 0.008955f
C4905 vdd.n3246 gnd 0.007208f
C4906 vdd.n3247 gnd 0.008955f
C4907 vdd.n3248 gnd 0.008955f
C4908 vdd.n3249 gnd 0.008955f
C4909 vdd.n3250 gnd 0.007208f
C4910 vdd.n3251 gnd 0.008955f
C4911 vdd.n3252 gnd 0.645204f
C4912 vdd.n3253 gnd 0.571989f
C4913 vdd.n3254 gnd 0.008955f
C4914 vdd.n3255 gnd 0.007208f
C4915 vdd.n3256 gnd 0.008955f
C4916 vdd.n3257 gnd 0.008955f
C4917 vdd.n3258 gnd 0.008955f
C4918 vdd.n3259 gnd 0.007208f
C4919 vdd.n3260 gnd 0.008955f
C4920 vdd.n3261 gnd 0.72757f
C4921 vdd.n3262 gnd 0.008955f
C4922 vdd.n3263 gnd 0.007208f
C4923 vdd.n3264 gnd 0.008955f
C4924 vdd.n3265 gnd 0.008955f
C4925 vdd.n3266 gnd 0.008955f
C4926 vdd.n3267 gnd 0.007208f
C4927 vdd.n3268 gnd 0.007208f
C4928 vdd.n3269 gnd 0.007208f
C4929 vdd.n3270 gnd 0.008955f
C4930 vdd.n3271 gnd 0.008955f
C4931 vdd.n3272 gnd 0.008955f
C4932 vdd.n3273 gnd 0.007208f
C4933 vdd.n3274 gnd 0.007208f
C4934 vdd.n3275 gnd 0.007208f
C4935 vdd.n3276 gnd 0.008955f
C4936 vdd.n3277 gnd 0.008955f
C4937 vdd.n3278 gnd 0.008955f
C4938 vdd.n3279 gnd 0.007208f
C4939 vdd.n3280 gnd 0.007208f
C4940 vdd.n3281 gnd 0.007208f
C4941 vdd.n3282 gnd 0.008955f
C4942 vdd.n3283 gnd 0.008955f
C4943 vdd.n3284 gnd 0.008955f
C4944 vdd.n3285 gnd 0.007208f
C4945 vdd.n3286 gnd 0.007208f
C4946 vdd.n3287 gnd 0.005983f
C4947 vdd.n3288 gnd 0.021104f
C4948 vdd.n3289 gnd 0.021434f
C4949 vdd.n3291 gnd 0.021434f
C4950 vdd.n3292 gnd 0.003424f
C4951 vdd.t59 gnd 0.110173f
C4952 vdd.t58 gnd 0.117745f
C4953 vdd.t57 gnd 0.143884f
C4954 vdd.n3293 gnd 0.184439f
C4955 vdd.n3294 gnd 0.155683f
C4956 vdd.n3295 gnd 0.011821f
C4957 vdd.n3296 gnd 0.003784f
C4958 vdd.n3297 gnd 0.007208f
C4959 vdd.n3298 gnd 0.008955f
C4960 vdd.n3300 gnd 0.008955f
C4961 vdd.n3301 gnd 0.008955f
C4962 vdd.n3302 gnd 0.007208f
C4963 vdd.n3303 gnd 0.007208f
C4964 vdd.n3304 gnd 0.007208f
C4965 vdd.n3305 gnd 0.008955f
C4966 vdd.n3307 gnd 0.008955f
C4967 vdd.n3308 gnd 0.008955f
C4968 vdd.n3309 gnd 0.007208f
C4969 vdd.n3310 gnd 0.007208f
C4970 vdd.n3311 gnd 0.007208f
C4971 vdd.n3312 gnd 0.008955f
C4972 vdd.n3314 gnd 0.008955f
C4973 vdd.n3315 gnd 0.008955f
C4974 vdd.n3316 gnd 0.007208f
C4975 vdd.n3317 gnd 0.007208f
C4976 vdd.n3318 gnd 0.007208f
C4977 vdd.n3319 gnd 0.008955f
C4978 vdd.n3321 gnd 0.008955f
C4979 vdd.n3322 gnd 0.008955f
C4980 vdd.n3323 gnd 0.007208f
C4981 vdd.n3324 gnd 0.007208f
C4982 vdd.n3325 gnd 0.007208f
C4983 vdd.n3326 gnd 0.008955f
C4984 vdd.n3328 gnd 0.008955f
C4985 vdd.n3329 gnd 0.008955f
C4986 vdd.n3330 gnd 0.007208f
C4987 vdd.n3331 gnd 0.008955f
C4988 vdd.n3332 gnd 0.008955f
C4989 vdd.n3333 gnd 0.008955f
C4990 vdd.n3334 gnd 0.015425f
C4991 vdd.n3335 gnd 0.004901f
C4992 vdd.n3336 gnd 0.007208f
C4993 vdd.n3337 gnd 0.008955f
C4994 vdd.n3339 gnd 0.008955f
C4995 vdd.n3340 gnd 0.008955f
C4996 vdd.n3341 gnd 0.007208f
C4997 vdd.n3342 gnd 0.007208f
C4998 vdd.n3343 gnd 0.007208f
C4999 vdd.n3344 gnd 0.008955f
C5000 vdd.n3346 gnd 0.008955f
C5001 vdd.n3347 gnd 0.008955f
C5002 vdd.n3348 gnd 0.007208f
C5003 vdd.n3349 gnd 0.007208f
C5004 vdd.n3350 gnd 0.007208f
C5005 vdd.n3351 gnd 0.008955f
C5006 vdd.n3353 gnd 0.008955f
C5007 vdd.n3354 gnd 0.008955f
C5008 vdd.n3355 gnd 0.007208f
C5009 vdd.n3356 gnd 0.007208f
C5010 vdd.n3357 gnd 0.007208f
C5011 vdd.n3358 gnd 0.008955f
C5012 vdd.n3360 gnd 0.008955f
C5013 vdd.n3361 gnd 0.008955f
C5014 vdd.n3362 gnd 0.007208f
C5015 vdd.n3363 gnd 0.007208f
C5016 vdd.n3364 gnd 0.007208f
C5017 vdd.n3365 gnd 0.008955f
C5018 vdd.n3367 gnd 0.008955f
C5019 vdd.n3368 gnd 0.008955f
C5020 vdd.n3369 gnd 0.007208f
C5021 vdd.n3370 gnd 0.008955f
C5022 vdd.n3371 gnd 0.008955f
C5023 vdd.n3372 gnd 0.008955f
C5024 vdd.n3373 gnd 0.015425f
C5025 vdd.n3374 gnd 0.006019f
C5026 vdd.n3375 gnd 0.007208f
C5027 vdd.n3376 gnd 0.008955f
C5028 vdd.n3378 gnd 0.008955f
C5029 vdd.n3379 gnd 0.008955f
C5030 vdd.n3380 gnd 0.007208f
C5031 vdd.n3381 gnd 0.007208f
C5032 vdd.n3382 gnd 0.007208f
C5033 vdd.n3383 gnd 0.008955f
C5034 vdd.n3385 gnd 0.008955f
C5035 vdd.n3386 gnd 0.008955f
C5036 vdd.n3387 gnd 0.007208f
C5037 vdd.n3388 gnd 0.007208f
C5038 vdd.n3389 gnd 0.007208f
C5039 vdd.n3390 gnd 0.008955f
C5040 vdd.n3392 gnd 0.008955f
C5041 vdd.n3393 gnd 0.008955f
C5042 vdd.n3394 gnd 0.007208f
C5043 vdd.n3395 gnd 0.007208f
C5044 vdd.n3396 gnd 0.007208f
C5045 vdd.n3397 gnd 0.008955f
C5046 vdd.n3399 gnd 0.008955f
C5047 vdd.n3400 gnd 0.008955f
C5048 vdd.n3402 gnd 0.008955f
C5049 vdd.n3403 gnd 0.007208f
C5050 vdd.n3404 gnd 0.007208f
C5051 vdd.n3405 gnd 0.005983f
C5052 vdd.n3406 gnd 0.021434f
C5053 vdd.n3407 gnd 0.021104f
C5054 vdd.n3408 gnd 0.005983f
C5055 vdd.n3409 gnd 0.021104f
C5056 vdd.n3410 gnd 1.29041f
C5057 vdd.n3411 gnd 0.517078f
C5058 vdd.t47 gnd 0.457591f
C5059 vdd.n3412 gnd 0.855696f
C5060 vdd.n3413 gnd 0.008955f
C5061 vdd.n3414 gnd 0.007208f
C5062 vdd.n3415 gnd 0.007208f
C5063 vdd.n3416 gnd 0.007208f
C5064 vdd.n3417 gnd 0.008955f
C5065 vdd.n3418 gnd 0.901455f
C5066 vdd.t22 gnd 0.457591f
C5067 vdd.n3419 gnd 0.471319f
C5068 vdd.n3420 gnd 0.745874f
C5069 vdd.n3421 gnd 0.008955f
C5070 vdd.n3422 gnd 0.007208f
C5071 vdd.n3423 gnd 0.007208f
C5072 vdd.n3424 gnd 0.007208f
C5073 vdd.n3425 gnd 0.008955f
C5074 vdd.n3426 gnd 0.590293f
C5075 vdd.t12 gnd 0.457591f
C5076 vdd.n3427 gnd 0.759602f
C5077 vdd.t128 gnd 0.457591f
C5078 vdd.n3428 gnd 0.480471f
C5079 vdd.n3429 gnd 0.008955f
C5080 vdd.n3430 gnd 0.007208f
C5081 vdd.n3431 gnd 0.007208f
C5082 vdd.n3432 gnd 0.007208f
C5083 vdd.n3433 gnd 0.008955f
C5084 vdd.n3434 gnd 0.636052f
C5085 vdd.n3435 gnd 0.581141f
C5086 vdd.t106 gnd 0.457591f
C5087 vdd.n3436 gnd 0.759602f
C5088 vdd.n3437 gnd 0.008955f
C5089 vdd.n3438 gnd 0.007208f
C5090 vdd.n3439 gnd 0.533085f
C5091 vdd.n3440 gnd 2.29851f
C5092 a_n2804_13878.t23 gnd 0.194556f
C5093 a_n2804_13878.t10 gnd 0.194556f
C5094 a_n2804_13878.t20 gnd 0.194556f
C5095 a_n2804_13878.n0 gnd 1.53358f
C5096 a_n2804_13878.t25 gnd 0.194556f
C5097 a_n2804_13878.t15 gnd 0.194556f
C5098 a_n2804_13878.n1 gnd 1.53196f
C5099 a_n2804_13878.n2 gnd 2.14061f
C5100 a_n2804_13878.t21 gnd 0.194556f
C5101 a_n2804_13878.t14 gnd 0.194556f
C5102 a_n2804_13878.n3 gnd 1.53196f
C5103 a_n2804_13878.n4 gnd 1.04414f
C5104 a_n2804_13878.t8 gnd 0.194556f
C5105 a_n2804_13878.t11 gnd 0.194556f
C5106 a_n2804_13878.n5 gnd 1.53196f
C5107 a_n2804_13878.n6 gnd 1.04414f
C5108 a_n2804_13878.t24 gnd 0.194556f
C5109 a_n2804_13878.t9 gnd 0.194556f
C5110 a_n2804_13878.n7 gnd 1.53196f
C5111 a_n2804_13878.n8 gnd 1.04414f
C5112 a_n2804_13878.t19 gnd 0.194556f
C5113 a_n2804_13878.t7 gnd 0.194556f
C5114 a_n2804_13878.n9 gnd 1.53196f
C5115 a_n2804_13878.n10 gnd 4.90178f
C5116 a_n2804_13878.t2 gnd 1.82172f
C5117 a_n2804_13878.t30 gnd 0.194556f
C5118 a_n2804_13878.t1 gnd 0.194556f
C5119 a_n2804_13878.n11 gnd 1.37045f
C5120 a_n2804_13878.n12 gnd 1.53128f
C5121 a_n2804_13878.t5 gnd 1.81809f
C5122 a_n2804_13878.n13 gnd 0.770559f
C5123 a_n2804_13878.t4 gnd 1.81809f
C5124 a_n2804_13878.n14 gnd 0.770559f
C5125 a_n2804_13878.t0 gnd 0.194556f
C5126 a_n2804_13878.t3 gnd 0.194556f
C5127 a_n2804_13878.n15 gnd 1.37045f
C5128 a_n2804_13878.n16 gnd 0.778022f
C5129 a_n2804_13878.t31 gnd 1.81809f
C5130 a_n2804_13878.n17 gnd 2.85814f
C5131 a_n2804_13878.n18 gnd 3.74876f
C5132 a_n2804_13878.t13 gnd 0.194556f
C5133 a_n2804_13878.t22 gnd 0.194556f
C5134 a_n2804_13878.n19 gnd 1.53195f
C5135 a_n2804_13878.n20 gnd 2.50239f
C5136 a_n2804_13878.t26 gnd 0.194556f
C5137 a_n2804_13878.t12 gnd 0.194556f
C5138 a_n2804_13878.n21 gnd 1.53196f
C5139 a_n2804_13878.n22 gnd 0.678771f
C5140 a_n2804_13878.t16 gnd 0.194556f
C5141 a_n2804_13878.t17 gnd 0.194556f
C5142 a_n2804_13878.n23 gnd 1.53196f
C5143 a_n2804_13878.n24 gnd 0.678771f
C5144 a_n2804_13878.t27 gnd 0.194556f
C5145 a_n2804_13878.t28 gnd 0.194556f
C5146 a_n2804_13878.n25 gnd 1.53196f
C5147 a_n2804_13878.n26 gnd 0.678771f
C5148 a_n2804_13878.t6 gnd 0.194556f
C5149 a_n2804_13878.t18 gnd 0.194556f
C5150 a_n2804_13878.n27 gnd 1.53196f
C5151 a_n2804_13878.n28 gnd 1.37704f
C5152 a_n2804_13878.n29 gnd 1.5345f
C5153 a_n2804_13878.t29 gnd 0.194556f
C5154 a_n2982_13878.n0 gnd 0.883913f
C5155 a_n2982_13878.n1 gnd 3.58469f
C5156 a_n2982_13878.n2 gnd 3.31432f
C5157 a_n2982_13878.n3 gnd 3.91444f
C5158 a_n2982_13878.n4 gnd 0.902552f
C5159 a_n2982_13878.n5 gnd 0.198406f
C5160 a_n2982_13878.n6 gnd 0.14613f
C5161 a_n2982_13878.n7 gnd 0.22967f
C5162 a_n2982_13878.n8 gnd 0.177393f
C5163 a_n2982_13878.n9 gnd 0.198406f
C5164 a_n2982_13878.n10 gnd 0.14613f
C5165 a_n2982_13878.n11 gnd 0.954828f
C5166 a_n2982_13878.n12 gnd 0.209105f
C5167 a_n2982_13878.n13 gnd 0.735977f
C5168 a_n2982_13878.n14 gnd 0.209105f
C5169 a_n2982_13878.n15 gnd 0.209105f
C5170 a_n2982_13878.n16 gnd 0.476233f
C5171 a_n2982_13878.n17 gnd 0.274168f
C5172 a_n2982_13878.n18 gnd 0.209105f
C5173 a_n2982_13878.n19 gnd 0.528509f
C5174 a_n2982_13878.n20 gnd 0.209105f
C5175 a_n2982_13878.n21 gnd 0.209105f
C5176 a_n2982_13878.n22 gnd 0.930364f
C5177 a_n2982_13878.n23 gnd 0.274168f
C5178 a_n2982_13878.n24 gnd 0.104552f
C5179 a_n2982_13878.n25 gnd 0.209105f
C5180 a_n2982_13878.n26 gnd 0.842549f
C5181 a_n2982_13878.n27 gnd 0.209105f
C5182 a_n2982_13878.n28 gnd 0.274168f
C5183 a_n2982_13878.n29 gnd 0.970217f
C5184 a_n2982_13878.n30 gnd 0.209105f
C5185 a_n2982_13878.n31 gnd 0.209105f
C5186 a_n2982_13878.n32 gnd 0.476233f
C5187 a_n2982_13878.n33 gnd 0.209105f
C5188 a_n2982_13878.n34 gnd 0.274168f
C5189 a_n2982_13878.n35 gnd 3.21642f
C5190 a_n2982_13878.n36 gnd 1.16f
C5191 a_n2982_13878.n37 gnd 2.11818f
C5192 a_n2982_13878.n38 gnd 1.72153f
C5193 a_n2982_13878.n39 gnd 1.16f
C5194 a_n2982_13878.n40 gnd 1.72153f
C5195 a_n2982_13878.n41 gnd 2.31679f
C5196 a_n2982_13878.n42 gnd 0.277359f
C5197 a_n2982_13878.n43 gnd 0.00839f
C5198 a_n2982_13878.n44 gnd 4.04e-19
C5199 a_n2982_13878.n46 gnd 0.008096f
C5200 a_n2982_13878.n47 gnd 0.011772f
C5201 a_n2982_13878.n48 gnd 0.007788f
C5202 a_n2982_13878.n50 gnd 1.64303f
C5203 a_n2982_13878.n51 gnd 0.277359f
C5204 a_n2982_13878.n52 gnd 0.00839f
C5205 a_n2982_13878.n53 gnd 4.04e-19
C5206 a_n2982_13878.n55 gnd 0.008096f
C5207 a_n2982_13878.n56 gnd 0.011772f
C5208 a_n2982_13878.n57 gnd 0.007788f
C5209 a_n2982_13878.n58 gnd 0.00839f
C5210 a_n2982_13878.n59 gnd 4.04e-19
C5211 a_n2982_13878.n61 gnd 0.008096f
C5212 a_n2982_13878.n62 gnd 0.011772f
C5213 a_n2982_13878.n63 gnd 0.007788f
C5214 a_n2982_13878.n65 gnd 0.277359f
C5215 a_n2982_13878.n66 gnd 0.00839f
C5216 a_n2982_13878.n67 gnd 4.04e-19
C5217 a_n2982_13878.n69 gnd 0.008096f
C5218 a_n2982_13878.n70 gnd 0.011772f
C5219 a_n2982_13878.n71 gnd 0.007788f
C5220 a_n2982_13878.n73 gnd 0.277359f
C5221 a_n2982_13878.n74 gnd 0.008096f
C5222 a_n2982_13878.n75 gnd 0.276227f
C5223 a_n2982_13878.n76 gnd 0.008096f
C5224 a_n2982_13878.n77 gnd 0.276227f
C5225 a_n2982_13878.n78 gnd 0.008096f
C5226 a_n2982_13878.n79 gnd 0.276227f
C5227 a_n2982_13878.n80 gnd 0.008096f
C5228 a_n2982_13878.n81 gnd 0.276227f
C5229 a_n2982_13878.n83 gnd 0.296601f
C5230 a_n2982_13878.t58 gnd 0.145037f
C5231 a_n2982_13878.t28 gnd 1.35806f
C5232 a_n2982_13878.t54 gnd 0.145037f
C5233 a_n2982_13878.t34 gnd 0.145037f
C5234 a_n2982_13878.n84 gnd 1.02164f
C5235 a_n2982_13878.t13 gnd 0.674643f
C5236 a_n2982_13878.n85 gnd 0.296601f
C5237 a_n2982_13878.t17 gnd 0.674643f
C5238 a_n2982_13878.t29 gnd 0.674643f
C5239 a_n2982_13878.n86 gnd 0.287692f
C5240 a_n2982_13878.t11 gnd 0.674643f
C5241 a_n2982_13878.n87 gnd 0.29915f
C5242 a_n2982_13878.t39 gnd 0.674643f
C5243 a_n2982_13878.t33 gnd 0.674643f
C5244 a_n2982_13878.n88 gnd 0.292527f
C5245 a_n2982_13878.t27 gnd 0.688688f
C5246 a_n2982_13878.t82 gnd 0.674643f
C5247 a_n2982_13878.n89 gnd 0.296601f
C5248 a_n2982_13878.t91 gnd 0.674643f
C5249 a_n2982_13878.t97 gnd 0.674643f
C5250 a_n2982_13878.n90 gnd 0.287692f
C5251 a_n2982_13878.t101 gnd 0.674643f
C5252 a_n2982_13878.n91 gnd 0.29915f
C5253 a_n2982_13878.t72 gnd 0.674643f
C5254 a_n2982_13878.t75 gnd 0.674643f
C5255 a_n2982_13878.n92 gnd 0.292527f
C5256 a_n2982_13878.t105 gnd 0.688688f
C5257 a_n2982_13878.t49 gnd 0.688688f
C5258 a_n2982_13878.t19 gnd 0.674643f
C5259 a_n2982_13878.t15 gnd 0.674643f
C5260 a_n2982_13878.t55 gnd 0.674643f
C5261 a_n2982_13878.n93 gnd 0.296483f
C5262 a_n2982_13878.t51 gnd 0.674643f
C5263 a_n2982_13878.t37 gnd 0.674643f
C5264 a_n2982_13878.t45 gnd 0.674643f
C5265 a_n2982_13878.n94 gnd 0.292849f
C5266 a_n2982_13878.t35 gnd 0.674643f
C5267 a_n2982_13878.t23 gnd 0.674643f
C5268 a_n2982_13878.t47 gnd 0.674643f
C5269 a_n2982_13878.t25 gnd 0.674643f
C5270 a_n2982_13878.t43 gnd 0.685497f
C5271 a_n2982_13878.t106 gnd 0.688688f
C5272 a_n2982_13878.t83 gnd 0.674643f
C5273 a_n2982_13878.t88 gnd 0.674643f
C5274 a_n2982_13878.t76 gnd 0.674643f
C5275 a_n2982_13878.n95 gnd 0.296483f
C5276 a_n2982_13878.t93 gnd 0.674643f
C5277 a_n2982_13878.t102 gnd 0.674643f
C5278 a_n2982_13878.t103 gnd 0.674643f
C5279 a_n2982_13878.n96 gnd 0.292849f
C5280 a_n2982_13878.t70 gnd 0.674643f
C5281 a_n2982_13878.t85 gnd 0.674643f
C5282 a_n2982_13878.t73 gnd 0.674643f
C5283 a_n2982_13878.n97 gnd 0.296601f
C5284 a_n2982_13878.t80 gnd 0.674643f
C5285 a_n2982_13878.t99 gnd 0.685497f
C5286 a_n2982_13878.n98 gnd 0.298713f
C5287 a_n2982_13878.n99 gnd 0.293101f
C5288 a_n2982_13878.n100 gnd 0.287692f
C5289 a_n2982_13878.n101 gnd 0.296616f
C5290 a_n2982_13878.n102 gnd 0.29915f
C5291 a_n2982_13878.n103 gnd 0.292527f
C5292 a_n2982_13878.n104 gnd 0.298713f
C5293 a_n2982_13878.n105 gnd 0.298713f
C5294 a_n2982_13878.t61 gnd 0.112807f
C5295 a_n2982_13878.t67 gnd 0.112807f
C5296 a_n2982_13878.n106 gnd 0.999739f
C5297 a_n2982_13878.t63 gnd 0.112807f
C5298 a_n2982_13878.t2 gnd 0.112807f
C5299 a_n2982_13878.n107 gnd 0.9968f
C5300 a_n2982_13878.t1 gnd 0.112807f
C5301 a_n2982_13878.t3 gnd 0.112807f
C5302 a_n2982_13878.n108 gnd 0.9968f
C5303 a_n2982_13878.t62 gnd 0.112807f
C5304 a_n2982_13878.t65 gnd 0.112807f
C5305 a_n2982_13878.n109 gnd 0.999739f
C5306 a_n2982_13878.t64 gnd 0.112807f
C5307 a_n2982_13878.t59 gnd 0.112807f
C5308 a_n2982_13878.n110 gnd 0.9968f
C5309 a_n2982_13878.t6 gnd 0.112807f
C5310 a_n2982_13878.t0 gnd 0.112807f
C5311 a_n2982_13878.n111 gnd 0.996801f
C5312 a_n2982_13878.t66 gnd 0.112807f
C5313 a_n2982_13878.t9 gnd 0.112807f
C5314 a_n2982_13878.n112 gnd 0.996801f
C5315 a_n2982_13878.t8 gnd 0.112807f
C5316 a_n2982_13878.t10 gnd 0.112807f
C5317 a_n2982_13878.n113 gnd 0.996801f
C5318 a_n2982_13878.t60 gnd 0.112807f
C5319 a_n2982_13878.t4 gnd 0.112807f
C5320 a_n2982_13878.n114 gnd 0.99974f
C5321 a_n2982_13878.t7 gnd 0.112807f
C5322 a_n2982_13878.t5 gnd 0.112807f
C5323 a_n2982_13878.n115 gnd 0.996801f
C5324 a_n2982_13878.n116 gnd 0.293101f
C5325 a_n2982_13878.n117 gnd 0.287692f
C5326 a_n2982_13878.n118 gnd 0.296616f
C5327 a_n2982_13878.n119 gnd 0.29915f
C5328 a_n2982_13878.n120 gnd 0.292527f
C5329 a_n2982_13878.n121 gnd 0.298713f
C5330 a_n2982_13878.t44 gnd 1.35806f
C5331 a_n2982_13878.t48 gnd 0.145037f
C5332 a_n2982_13878.t26 gnd 0.145037f
C5333 a_n2982_13878.n122 gnd 1.02164f
C5334 a_n2982_13878.t36 gnd 0.145037f
C5335 a_n2982_13878.t24 gnd 0.145037f
C5336 a_n2982_13878.n123 gnd 1.02164f
C5337 a_n2982_13878.t38 gnd 0.145037f
C5338 a_n2982_13878.t46 gnd 0.145037f
C5339 a_n2982_13878.n124 gnd 1.02164f
C5340 a_n2982_13878.t56 gnd 0.145037f
C5341 a_n2982_13878.t52 gnd 0.145037f
C5342 a_n2982_13878.n125 gnd 1.02164f
C5343 a_n2982_13878.t20 gnd 0.145037f
C5344 a_n2982_13878.t16 gnd 0.145037f
C5345 a_n2982_13878.n126 gnd 1.02164f
C5346 a_n2982_13878.t50 gnd 1.35535f
C5347 a_n2982_13878.n127 gnd 0.993167f
C5348 a_n2982_13878.t81 gnd 0.674643f
C5349 a_n2982_13878.t92 gnd 0.674643f
C5350 a_n2982_13878.t107 gnd 0.674643f
C5351 a_n2982_13878.n128 gnd 0.296616f
C5352 a_n2982_13878.t94 gnd 0.674643f
C5353 a_n2982_13878.t77 gnd 0.674643f
C5354 a_n2982_13878.t78 gnd 0.674643f
C5355 a_n2982_13878.n129 gnd 0.296616f
C5356 a_n2982_13878.t98 gnd 0.674643f
C5357 a_n2982_13878.t87 gnd 0.674643f
C5358 a_n2982_13878.t86 gnd 0.674643f
C5359 a_n2982_13878.n130 gnd 0.296616f
C5360 a_n2982_13878.t90 gnd 0.674643f
C5361 a_n2982_13878.t79 gnd 0.674643f
C5362 a_n2982_13878.t68 gnd 0.674643f
C5363 a_n2982_13878.n131 gnd 0.296616f
C5364 a_n2982_13878.t95 gnd 0.685948f
C5365 a_n2982_13878.n132 gnd 0.292849f
C5366 a_n2982_13878.n133 gnd 0.287531f
C5367 a_n2982_13878.t104 gnd 0.685948f
C5368 a_n2982_13878.n134 gnd 0.292849f
C5369 a_n2982_13878.n135 gnd 0.287531f
C5370 a_n2982_13878.t89 gnd 0.685948f
C5371 a_n2982_13878.n136 gnd 0.292849f
C5372 a_n2982_13878.n137 gnd 0.287531f
C5373 a_n2982_13878.t84 gnd 0.685948f
C5374 a_n2982_13878.n138 gnd 0.292849f
C5375 a_n2982_13878.n139 gnd 0.287531f
C5376 a_n2982_13878.n140 gnd 1.32168f
C5377 a_n2982_13878.t74 gnd 0.674643f
C5378 a_n2982_13878.n141 gnd 0.298713f
C5379 a_n2982_13878.t100 gnd 0.674643f
C5380 a_n2982_13878.n142 gnd 0.296483f
C5381 a_n2982_13878.n143 gnd 0.296616f
C5382 a_n2982_13878.t96 gnd 0.674643f
C5383 a_n2982_13878.n144 gnd 0.292849f
C5384 a_n2982_13878.t69 gnd 0.674643f
C5385 a_n2982_13878.n145 gnd 0.293101f
C5386 a_n2982_13878.n146 gnd 0.298713f
C5387 a_n2982_13878.t71 gnd 0.685497f
C5388 a_n2982_13878.t53 gnd 0.674643f
C5389 a_n2982_13878.n147 gnd 0.298713f
C5390 a_n2982_13878.t57 gnd 0.674643f
C5391 a_n2982_13878.n148 gnd 0.296483f
C5392 a_n2982_13878.n149 gnd 0.296616f
C5393 a_n2982_13878.t41 gnd 0.674643f
C5394 a_n2982_13878.n150 gnd 0.292849f
C5395 a_n2982_13878.t31 gnd 0.674643f
C5396 a_n2982_13878.n151 gnd 0.293101f
C5397 a_n2982_13878.n152 gnd 0.298713f
C5398 a_n2982_13878.t21 gnd 0.685497f
C5399 a_n2982_13878.n153 gnd 1.30619f
C5400 a_n2982_13878.t22 gnd 1.35535f
C5401 a_n2982_13878.t14 gnd 0.145037f
C5402 a_n2982_13878.t18 gnd 0.145037f
C5403 a_n2982_13878.n154 gnd 1.02164f
C5404 a_n2982_13878.t30 gnd 0.145037f
C5405 a_n2982_13878.t32 gnd 0.145037f
C5406 a_n2982_13878.n155 gnd 1.02164f
C5407 a_n2982_13878.t40 gnd 0.145037f
C5408 a_n2982_13878.t42 gnd 0.145037f
C5409 a_n2982_13878.n156 gnd 1.02164f
C5410 a_n2982_13878.n157 gnd 1.02165f
C5411 a_n2982_13878.t12 gnd 0.145037f
C5412 commonsourceibias.n0 gnd 0.012818f
C5413 commonsourceibias.t104 gnd 0.19409f
C5414 commonsourceibias.t181 gnd 0.179464f
C5415 commonsourceibias.n1 gnd 0.00935f
C5416 commonsourceibias.n2 gnd 0.009606f
C5417 commonsourceibias.t124 gnd 0.179464f
C5418 commonsourceibias.n3 gnd 0.012358f
C5419 commonsourceibias.n4 gnd 0.009606f
C5420 commonsourceibias.t197 gnd 0.179464f
C5421 commonsourceibias.n5 gnd 0.071606f
C5422 commonsourceibias.t142 gnd 0.179464f
C5423 commonsourceibias.n6 gnd 0.009057f
C5424 commonsourceibias.n7 gnd 0.009606f
C5425 commonsourceibias.t101 gnd 0.179464f
C5426 commonsourceibias.n8 gnd 0.012175f
C5427 commonsourceibias.n9 gnd 0.009606f
C5428 commonsourceibias.t156 gnd 0.179464f
C5429 commonsourceibias.n10 gnd 0.071606f
C5430 commonsourceibias.t143 gnd 0.179464f
C5431 commonsourceibias.n11 gnd 0.008798f
C5432 commonsourceibias.n12 gnd 0.009606f
C5433 commonsourceibias.t193 gnd 0.179464f
C5434 commonsourceibias.n13 gnd 0.01197f
C5435 commonsourceibias.n14 gnd 0.012818f
C5436 commonsourceibias.t72 gnd 0.19409f
C5437 commonsourceibias.t42 gnd 0.179464f
C5438 commonsourceibias.n15 gnd 0.00935f
C5439 commonsourceibias.n16 gnd 0.009606f
C5440 commonsourceibias.t44 gnd 0.179464f
C5441 commonsourceibias.n17 gnd 0.012358f
C5442 commonsourceibias.n18 gnd 0.009606f
C5443 commonsourceibias.t6 gnd 0.179464f
C5444 commonsourceibias.n19 gnd 0.071606f
C5445 commonsourceibias.t52 gnd 0.179464f
C5446 commonsourceibias.n20 gnd 0.009057f
C5447 commonsourceibias.n21 gnd 0.009606f
C5448 commonsourceibias.t74 gnd 0.179464f
C5449 commonsourceibias.n22 gnd 0.012175f
C5450 commonsourceibias.n23 gnd 0.009606f
C5451 commonsourceibias.t16 gnd 0.179464f
C5452 commonsourceibias.n24 gnd 0.071606f
C5453 commonsourceibias.t50 gnd 0.179464f
C5454 commonsourceibias.n25 gnd 0.008798f
C5455 commonsourceibias.n26 gnd 0.009606f
C5456 commonsourceibias.t32 gnd 0.179464f
C5457 commonsourceibias.n27 gnd 0.01197f
C5458 commonsourceibias.n28 gnd 0.009606f
C5459 commonsourceibias.t56 gnd 0.179464f
C5460 commonsourceibias.n29 gnd 0.071606f
C5461 commonsourceibias.t26 gnd 0.179464f
C5462 commonsourceibias.n30 gnd 0.008572f
C5463 commonsourceibias.n31 gnd 0.009606f
C5464 commonsourceibias.t20 gnd 0.179464f
C5465 commonsourceibias.n32 gnd 0.011742f
C5466 commonsourceibias.n33 gnd 0.009606f
C5467 commonsourceibias.t54 gnd 0.179464f
C5468 commonsourceibias.n34 gnd 0.071606f
C5469 commonsourceibias.t68 gnd 0.179464f
C5470 commonsourceibias.n35 gnd 0.008375f
C5471 commonsourceibias.n36 gnd 0.009606f
C5472 commonsourceibias.t38 gnd 0.179464f
C5473 commonsourceibias.n37 gnd 0.011489f
C5474 commonsourceibias.n38 gnd 0.009606f
C5475 commonsourceibias.t14 gnd 0.179464f
C5476 commonsourceibias.n39 gnd 0.071606f
C5477 commonsourceibias.t46 gnd 0.179464f
C5478 commonsourceibias.n40 gnd 0.008208f
C5479 commonsourceibias.n41 gnd 0.009606f
C5480 commonsourceibias.t2 gnd 0.179464f
C5481 commonsourceibias.n42 gnd 0.011208f
C5482 commonsourceibias.t76 gnd 0.199531f
C5483 commonsourceibias.t10 gnd 0.179464f
C5484 commonsourceibias.n43 gnd 0.078223f
C5485 commonsourceibias.n44 gnd 0.08584f
C5486 commonsourceibias.n45 gnd 0.039831f
C5487 commonsourceibias.n46 gnd 0.009606f
C5488 commonsourceibias.n47 gnd 0.00935f
C5489 commonsourceibias.n48 gnd 0.013398f
C5490 commonsourceibias.n49 gnd 0.071606f
C5491 commonsourceibias.n50 gnd 0.013389f
C5492 commonsourceibias.n51 gnd 0.009606f
C5493 commonsourceibias.n52 gnd 0.009606f
C5494 commonsourceibias.n53 gnd 0.009606f
C5495 commonsourceibias.n54 gnd 0.012358f
C5496 commonsourceibias.n55 gnd 0.071606f
C5497 commonsourceibias.n56 gnd 0.012648f
C5498 commonsourceibias.n57 gnd 0.012289f
C5499 commonsourceibias.n58 gnd 0.009606f
C5500 commonsourceibias.n59 gnd 0.009606f
C5501 commonsourceibias.n60 gnd 0.009606f
C5502 commonsourceibias.n61 gnd 0.009057f
C5503 commonsourceibias.n62 gnd 0.01341f
C5504 commonsourceibias.n63 gnd 0.071606f
C5505 commonsourceibias.n64 gnd 0.013406f
C5506 commonsourceibias.n65 gnd 0.009606f
C5507 commonsourceibias.n66 gnd 0.009606f
C5508 commonsourceibias.n67 gnd 0.009606f
C5509 commonsourceibias.n68 gnd 0.012175f
C5510 commonsourceibias.n69 gnd 0.071606f
C5511 commonsourceibias.n70 gnd 0.012558f
C5512 commonsourceibias.n71 gnd 0.012378f
C5513 commonsourceibias.n72 gnd 0.009606f
C5514 commonsourceibias.n73 gnd 0.009606f
C5515 commonsourceibias.n74 gnd 0.009606f
C5516 commonsourceibias.n75 gnd 0.008798f
C5517 commonsourceibias.n76 gnd 0.013416f
C5518 commonsourceibias.n77 gnd 0.071606f
C5519 commonsourceibias.n78 gnd 0.013414f
C5520 commonsourceibias.n79 gnd 0.009606f
C5521 commonsourceibias.n80 gnd 0.009606f
C5522 commonsourceibias.n81 gnd 0.009606f
C5523 commonsourceibias.n82 gnd 0.01197f
C5524 commonsourceibias.n83 gnd 0.071606f
C5525 commonsourceibias.n84 gnd 0.012468f
C5526 commonsourceibias.n85 gnd 0.012468f
C5527 commonsourceibias.n86 gnd 0.009606f
C5528 commonsourceibias.n87 gnd 0.009606f
C5529 commonsourceibias.n88 gnd 0.009606f
C5530 commonsourceibias.n89 gnd 0.008572f
C5531 commonsourceibias.n90 gnd 0.013414f
C5532 commonsourceibias.n91 gnd 0.071606f
C5533 commonsourceibias.n92 gnd 0.013416f
C5534 commonsourceibias.n93 gnd 0.009606f
C5535 commonsourceibias.n94 gnd 0.009606f
C5536 commonsourceibias.n95 gnd 0.009606f
C5537 commonsourceibias.n96 gnd 0.011742f
C5538 commonsourceibias.n97 gnd 0.071606f
C5539 commonsourceibias.n98 gnd 0.012378f
C5540 commonsourceibias.n99 gnd 0.012558f
C5541 commonsourceibias.n100 gnd 0.009606f
C5542 commonsourceibias.n101 gnd 0.009606f
C5543 commonsourceibias.n102 gnd 0.009606f
C5544 commonsourceibias.n103 gnd 0.008375f
C5545 commonsourceibias.n104 gnd 0.013406f
C5546 commonsourceibias.n105 gnd 0.071606f
C5547 commonsourceibias.n106 gnd 0.01341f
C5548 commonsourceibias.n107 gnd 0.009606f
C5549 commonsourceibias.n108 gnd 0.009606f
C5550 commonsourceibias.n109 gnd 0.009606f
C5551 commonsourceibias.n110 gnd 0.011489f
C5552 commonsourceibias.n111 gnd 0.071606f
C5553 commonsourceibias.n112 gnd 0.012289f
C5554 commonsourceibias.n113 gnd 0.012648f
C5555 commonsourceibias.n114 gnd 0.009606f
C5556 commonsourceibias.n115 gnd 0.009606f
C5557 commonsourceibias.n116 gnd 0.009606f
C5558 commonsourceibias.n117 gnd 0.008208f
C5559 commonsourceibias.n118 gnd 0.013389f
C5560 commonsourceibias.n119 gnd 0.071606f
C5561 commonsourceibias.n120 gnd 0.013398f
C5562 commonsourceibias.n121 gnd 0.009606f
C5563 commonsourceibias.n122 gnd 0.009606f
C5564 commonsourceibias.n123 gnd 0.009606f
C5565 commonsourceibias.n124 gnd 0.011208f
C5566 commonsourceibias.n125 gnd 0.071606f
C5567 commonsourceibias.n126 gnd 0.011785f
C5568 commonsourceibias.n127 gnd 0.085921f
C5569 commonsourceibias.n128 gnd 0.095704f
C5570 commonsourceibias.t73 gnd 0.020728f
C5571 commonsourceibias.t43 gnd 0.020728f
C5572 commonsourceibias.n129 gnd 0.183161f
C5573 commonsourceibias.n130 gnd 0.158435f
C5574 commonsourceibias.t45 gnd 0.020728f
C5575 commonsourceibias.t7 gnd 0.020728f
C5576 commonsourceibias.n131 gnd 0.183161f
C5577 commonsourceibias.n132 gnd 0.084133f
C5578 commonsourceibias.t53 gnd 0.020728f
C5579 commonsourceibias.t75 gnd 0.020728f
C5580 commonsourceibias.n133 gnd 0.183161f
C5581 commonsourceibias.n134 gnd 0.084133f
C5582 commonsourceibias.t17 gnd 0.020728f
C5583 commonsourceibias.t51 gnd 0.020728f
C5584 commonsourceibias.n135 gnd 0.183161f
C5585 commonsourceibias.n136 gnd 0.084133f
C5586 commonsourceibias.t33 gnd 0.020728f
C5587 commonsourceibias.t57 gnd 0.020728f
C5588 commonsourceibias.n137 gnd 0.183161f
C5589 commonsourceibias.n138 gnd 0.070289f
C5590 commonsourceibias.t11 gnd 0.020728f
C5591 commonsourceibias.t77 gnd 0.020728f
C5592 commonsourceibias.n139 gnd 0.183774f
C5593 commonsourceibias.t47 gnd 0.020728f
C5594 commonsourceibias.t3 gnd 0.020728f
C5595 commonsourceibias.n140 gnd 0.183161f
C5596 commonsourceibias.n141 gnd 0.170671f
C5597 commonsourceibias.t39 gnd 0.020728f
C5598 commonsourceibias.t15 gnd 0.020728f
C5599 commonsourceibias.n142 gnd 0.183161f
C5600 commonsourceibias.n143 gnd 0.084133f
C5601 commonsourceibias.t55 gnd 0.020728f
C5602 commonsourceibias.t69 gnd 0.020728f
C5603 commonsourceibias.n144 gnd 0.183161f
C5604 commonsourceibias.n145 gnd 0.084133f
C5605 commonsourceibias.t27 gnd 0.020728f
C5606 commonsourceibias.t21 gnd 0.020728f
C5607 commonsourceibias.n146 gnd 0.183161f
C5608 commonsourceibias.n147 gnd 0.070289f
C5609 commonsourceibias.n148 gnd 0.085113f
C5610 commonsourceibias.n149 gnd 0.062168f
C5611 commonsourceibias.t136 gnd 0.179464f
C5612 commonsourceibias.n150 gnd 0.071606f
C5613 commonsourceibias.t119 gnd 0.179464f
C5614 commonsourceibias.n151 gnd 0.071606f
C5615 commonsourceibias.n152 gnd 0.009606f
C5616 commonsourceibias.t155 gnd 0.179464f
C5617 commonsourceibias.n153 gnd 0.071606f
C5618 commonsourceibias.n154 gnd 0.009606f
C5619 commonsourceibias.t140 gnd 0.179464f
C5620 commonsourceibias.n155 gnd 0.071606f
C5621 commonsourceibias.n156 gnd 0.009606f
C5622 commonsourceibias.t109 gnd 0.179464f
C5623 commonsourceibias.n157 gnd 0.008375f
C5624 commonsourceibias.n158 gnd 0.009606f
C5625 commonsourceibias.t182 gnd 0.179464f
C5626 commonsourceibias.n159 gnd 0.011489f
C5627 commonsourceibias.n160 gnd 0.009606f
C5628 commonsourceibias.t166 gnd 0.179464f
C5629 commonsourceibias.n161 gnd 0.071606f
C5630 commonsourceibias.t123 gnd 0.179464f
C5631 commonsourceibias.n162 gnd 0.008208f
C5632 commonsourceibias.n163 gnd 0.009606f
C5633 commonsourceibias.t84 gnd 0.179464f
C5634 commonsourceibias.n164 gnd 0.011208f
C5635 commonsourceibias.t100 gnd 0.199531f
C5636 commonsourceibias.t131 gnd 0.179464f
C5637 commonsourceibias.n165 gnd 0.078223f
C5638 commonsourceibias.n166 gnd 0.08584f
C5639 commonsourceibias.n167 gnd 0.039831f
C5640 commonsourceibias.n168 gnd 0.009606f
C5641 commonsourceibias.n169 gnd 0.00935f
C5642 commonsourceibias.n170 gnd 0.013398f
C5643 commonsourceibias.n171 gnd 0.071606f
C5644 commonsourceibias.n172 gnd 0.013389f
C5645 commonsourceibias.n173 gnd 0.009606f
C5646 commonsourceibias.n174 gnd 0.009606f
C5647 commonsourceibias.n175 gnd 0.009606f
C5648 commonsourceibias.n176 gnd 0.012358f
C5649 commonsourceibias.n177 gnd 0.071606f
C5650 commonsourceibias.n178 gnd 0.012648f
C5651 commonsourceibias.n179 gnd 0.012289f
C5652 commonsourceibias.n180 gnd 0.009606f
C5653 commonsourceibias.n181 gnd 0.009606f
C5654 commonsourceibias.n182 gnd 0.009606f
C5655 commonsourceibias.n183 gnd 0.009057f
C5656 commonsourceibias.n184 gnd 0.01341f
C5657 commonsourceibias.n185 gnd 0.071606f
C5658 commonsourceibias.n186 gnd 0.013406f
C5659 commonsourceibias.n187 gnd 0.009606f
C5660 commonsourceibias.n188 gnd 0.009606f
C5661 commonsourceibias.n189 gnd 0.009606f
C5662 commonsourceibias.n190 gnd 0.012175f
C5663 commonsourceibias.n191 gnd 0.071606f
C5664 commonsourceibias.n192 gnd 0.012558f
C5665 commonsourceibias.n193 gnd 0.012378f
C5666 commonsourceibias.n194 gnd 0.009606f
C5667 commonsourceibias.n195 gnd 0.009606f
C5668 commonsourceibias.n196 gnd 0.011742f
C5669 commonsourceibias.n197 gnd 0.008798f
C5670 commonsourceibias.n198 gnd 0.013416f
C5671 commonsourceibias.n199 gnd 0.009606f
C5672 commonsourceibias.n200 gnd 0.009606f
C5673 commonsourceibias.n201 gnd 0.013414f
C5674 commonsourceibias.n202 gnd 0.008572f
C5675 commonsourceibias.n203 gnd 0.01197f
C5676 commonsourceibias.n204 gnd 0.009606f
C5677 commonsourceibias.n205 gnd 0.008392f
C5678 commonsourceibias.n206 gnd 0.012468f
C5679 commonsourceibias.n207 gnd 0.012468f
C5680 commonsourceibias.n208 gnd 0.008392f
C5681 commonsourceibias.n209 gnd 0.009606f
C5682 commonsourceibias.n210 gnd 0.009606f
C5683 commonsourceibias.n211 gnd 0.008572f
C5684 commonsourceibias.n212 gnd 0.013414f
C5685 commonsourceibias.n213 gnd 0.071606f
C5686 commonsourceibias.n214 gnd 0.013416f
C5687 commonsourceibias.n215 gnd 0.009606f
C5688 commonsourceibias.n216 gnd 0.009606f
C5689 commonsourceibias.n217 gnd 0.009606f
C5690 commonsourceibias.n218 gnd 0.011742f
C5691 commonsourceibias.n219 gnd 0.071606f
C5692 commonsourceibias.n220 gnd 0.012378f
C5693 commonsourceibias.n221 gnd 0.012558f
C5694 commonsourceibias.n222 gnd 0.009606f
C5695 commonsourceibias.n223 gnd 0.009606f
C5696 commonsourceibias.n224 gnd 0.009606f
C5697 commonsourceibias.n225 gnd 0.008375f
C5698 commonsourceibias.n226 gnd 0.013406f
C5699 commonsourceibias.n227 gnd 0.071606f
C5700 commonsourceibias.n228 gnd 0.01341f
C5701 commonsourceibias.n229 gnd 0.009606f
C5702 commonsourceibias.n230 gnd 0.009606f
C5703 commonsourceibias.n231 gnd 0.009606f
C5704 commonsourceibias.n232 gnd 0.011489f
C5705 commonsourceibias.n233 gnd 0.071606f
C5706 commonsourceibias.n234 gnd 0.012289f
C5707 commonsourceibias.n235 gnd 0.012648f
C5708 commonsourceibias.n236 gnd 0.009606f
C5709 commonsourceibias.n237 gnd 0.009606f
C5710 commonsourceibias.n238 gnd 0.009606f
C5711 commonsourceibias.n239 gnd 0.008208f
C5712 commonsourceibias.n240 gnd 0.013389f
C5713 commonsourceibias.n241 gnd 0.071606f
C5714 commonsourceibias.n242 gnd 0.013398f
C5715 commonsourceibias.n243 gnd 0.009606f
C5716 commonsourceibias.n244 gnd 0.009606f
C5717 commonsourceibias.n245 gnd 0.009606f
C5718 commonsourceibias.n246 gnd 0.011208f
C5719 commonsourceibias.n247 gnd 0.071606f
C5720 commonsourceibias.n248 gnd 0.011785f
C5721 commonsourceibias.n249 gnd 0.085921f
C5722 commonsourceibias.n250 gnd 0.056157f
C5723 commonsourceibias.n251 gnd 0.012818f
C5724 commonsourceibias.t145 gnd 0.19409f
C5725 commonsourceibias.t172 gnd 0.179464f
C5726 commonsourceibias.n252 gnd 0.00935f
C5727 commonsourceibias.n253 gnd 0.009606f
C5728 commonsourceibias.t160 gnd 0.179464f
C5729 commonsourceibias.n254 gnd 0.012358f
C5730 commonsourceibias.n255 gnd 0.009606f
C5731 commonsourceibias.t146 gnd 0.179464f
C5732 commonsourceibias.n256 gnd 0.071606f
C5733 commonsourceibias.t173 gnd 0.179464f
C5734 commonsourceibias.n257 gnd 0.009057f
C5735 commonsourceibias.n258 gnd 0.009606f
C5736 commonsourceibias.t158 gnd 0.179464f
C5737 commonsourceibias.n259 gnd 0.012175f
C5738 commonsourceibias.n260 gnd 0.009606f
C5739 commonsourceibias.t144 gnd 0.179464f
C5740 commonsourceibias.n261 gnd 0.071606f
C5741 commonsourceibias.t174 gnd 0.179464f
C5742 commonsourceibias.n262 gnd 0.008798f
C5743 commonsourceibias.n263 gnd 0.009606f
C5744 commonsourceibias.t159 gnd 0.179464f
C5745 commonsourceibias.n264 gnd 0.01197f
C5746 commonsourceibias.n265 gnd 0.009606f
C5747 commonsourceibias.t185 gnd 0.179464f
C5748 commonsourceibias.n266 gnd 0.071606f
C5749 commonsourceibias.t175 gnd 0.179464f
C5750 commonsourceibias.n267 gnd 0.008572f
C5751 commonsourceibias.n268 gnd 0.009606f
C5752 commonsourceibias.t157 gnd 0.179464f
C5753 commonsourceibias.n269 gnd 0.011742f
C5754 commonsourceibias.n270 gnd 0.009606f
C5755 commonsourceibias.t190 gnd 0.179464f
C5756 commonsourceibias.n271 gnd 0.071606f
C5757 commonsourceibias.t91 gnd 0.179464f
C5758 commonsourceibias.n272 gnd 0.008375f
C5759 commonsourceibias.n273 gnd 0.009606f
C5760 commonsourceibias.t169 gnd 0.179464f
C5761 commonsourceibias.n274 gnd 0.011489f
C5762 commonsourceibias.n275 gnd 0.009606f
C5763 commonsourceibias.t82 gnd 0.179464f
C5764 commonsourceibias.n276 gnd 0.071606f
C5765 commonsourceibias.t95 gnd 0.179464f
C5766 commonsourceibias.n277 gnd 0.008208f
C5767 commonsourceibias.n278 gnd 0.009606f
C5768 commonsourceibias.t90 gnd 0.179464f
C5769 commonsourceibias.n279 gnd 0.011208f
C5770 commonsourceibias.t94 gnd 0.199531f
C5771 commonsourceibias.t80 gnd 0.179464f
C5772 commonsourceibias.n280 gnd 0.078223f
C5773 commonsourceibias.n281 gnd 0.08584f
C5774 commonsourceibias.n282 gnd 0.039831f
C5775 commonsourceibias.n283 gnd 0.009606f
C5776 commonsourceibias.n284 gnd 0.00935f
C5777 commonsourceibias.n285 gnd 0.013398f
C5778 commonsourceibias.n286 gnd 0.071606f
C5779 commonsourceibias.n287 gnd 0.013389f
C5780 commonsourceibias.n288 gnd 0.009606f
C5781 commonsourceibias.n289 gnd 0.009606f
C5782 commonsourceibias.n290 gnd 0.009606f
C5783 commonsourceibias.n291 gnd 0.012358f
C5784 commonsourceibias.n292 gnd 0.071606f
C5785 commonsourceibias.n293 gnd 0.012648f
C5786 commonsourceibias.n294 gnd 0.012289f
C5787 commonsourceibias.n295 gnd 0.009606f
C5788 commonsourceibias.n296 gnd 0.009606f
C5789 commonsourceibias.n297 gnd 0.009606f
C5790 commonsourceibias.n298 gnd 0.009057f
C5791 commonsourceibias.n299 gnd 0.01341f
C5792 commonsourceibias.n300 gnd 0.071606f
C5793 commonsourceibias.n301 gnd 0.013406f
C5794 commonsourceibias.n302 gnd 0.009606f
C5795 commonsourceibias.n303 gnd 0.009606f
C5796 commonsourceibias.n304 gnd 0.009606f
C5797 commonsourceibias.n305 gnd 0.012175f
C5798 commonsourceibias.n306 gnd 0.071606f
C5799 commonsourceibias.n307 gnd 0.012558f
C5800 commonsourceibias.n308 gnd 0.012378f
C5801 commonsourceibias.n309 gnd 0.009606f
C5802 commonsourceibias.n310 gnd 0.009606f
C5803 commonsourceibias.n311 gnd 0.009606f
C5804 commonsourceibias.n312 gnd 0.008798f
C5805 commonsourceibias.n313 gnd 0.013416f
C5806 commonsourceibias.n314 gnd 0.071606f
C5807 commonsourceibias.n315 gnd 0.013414f
C5808 commonsourceibias.n316 gnd 0.009606f
C5809 commonsourceibias.n317 gnd 0.009606f
C5810 commonsourceibias.n318 gnd 0.009606f
C5811 commonsourceibias.n319 gnd 0.01197f
C5812 commonsourceibias.n320 gnd 0.071606f
C5813 commonsourceibias.n321 gnd 0.012468f
C5814 commonsourceibias.n322 gnd 0.012468f
C5815 commonsourceibias.n323 gnd 0.009606f
C5816 commonsourceibias.n324 gnd 0.009606f
C5817 commonsourceibias.n325 gnd 0.009606f
C5818 commonsourceibias.n326 gnd 0.008572f
C5819 commonsourceibias.n327 gnd 0.013414f
C5820 commonsourceibias.n328 gnd 0.071606f
C5821 commonsourceibias.n329 gnd 0.013416f
C5822 commonsourceibias.n330 gnd 0.009606f
C5823 commonsourceibias.n331 gnd 0.009606f
C5824 commonsourceibias.n332 gnd 0.009606f
C5825 commonsourceibias.n333 gnd 0.011742f
C5826 commonsourceibias.n334 gnd 0.071606f
C5827 commonsourceibias.n335 gnd 0.012378f
C5828 commonsourceibias.n336 gnd 0.012558f
C5829 commonsourceibias.n337 gnd 0.009606f
C5830 commonsourceibias.n338 gnd 0.009606f
C5831 commonsourceibias.n339 gnd 0.009606f
C5832 commonsourceibias.n340 gnd 0.008375f
C5833 commonsourceibias.n341 gnd 0.013406f
C5834 commonsourceibias.n342 gnd 0.071606f
C5835 commonsourceibias.n343 gnd 0.01341f
C5836 commonsourceibias.n344 gnd 0.009606f
C5837 commonsourceibias.n345 gnd 0.009606f
C5838 commonsourceibias.n346 gnd 0.009606f
C5839 commonsourceibias.n347 gnd 0.011489f
C5840 commonsourceibias.n348 gnd 0.071606f
C5841 commonsourceibias.n349 gnd 0.012289f
C5842 commonsourceibias.n350 gnd 0.012648f
C5843 commonsourceibias.n351 gnd 0.009606f
C5844 commonsourceibias.n352 gnd 0.009606f
C5845 commonsourceibias.n353 gnd 0.009606f
C5846 commonsourceibias.n354 gnd 0.008208f
C5847 commonsourceibias.n355 gnd 0.013389f
C5848 commonsourceibias.n356 gnd 0.071606f
C5849 commonsourceibias.n357 gnd 0.013398f
C5850 commonsourceibias.n358 gnd 0.009606f
C5851 commonsourceibias.n359 gnd 0.009606f
C5852 commonsourceibias.n360 gnd 0.009606f
C5853 commonsourceibias.n361 gnd 0.011208f
C5854 commonsourceibias.n362 gnd 0.071606f
C5855 commonsourceibias.n363 gnd 0.011785f
C5856 commonsourceibias.n364 gnd 0.085921f
C5857 commonsourceibias.n365 gnd 0.029883f
C5858 commonsourceibias.n366 gnd 0.153513f
C5859 commonsourceibias.n367 gnd 0.012818f
C5860 commonsourceibias.t89 gnd 0.179464f
C5861 commonsourceibias.n368 gnd 0.00935f
C5862 commonsourceibias.n369 gnd 0.009606f
C5863 commonsourceibias.t107 gnd 0.179464f
C5864 commonsourceibias.n370 gnd 0.012358f
C5865 commonsourceibias.n371 gnd 0.009606f
C5866 commonsourceibias.t168 gnd 0.179464f
C5867 commonsourceibias.n372 gnd 0.071606f
C5868 commonsourceibias.t199 gnd 0.179464f
C5869 commonsourceibias.n373 gnd 0.009057f
C5870 commonsourceibias.n374 gnd 0.009606f
C5871 commonsourceibias.t98 gnd 0.179464f
C5872 commonsourceibias.n375 gnd 0.012175f
C5873 commonsourceibias.n376 gnd 0.009606f
C5874 commonsourceibias.t150 gnd 0.179464f
C5875 commonsourceibias.n377 gnd 0.071606f
C5876 commonsourceibias.t141 gnd 0.179464f
C5877 commonsourceibias.n378 gnd 0.008798f
C5878 commonsourceibias.n379 gnd 0.009606f
C5879 commonsourceibias.t88 gnd 0.179464f
C5880 commonsourceibias.n380 gnd 0.01197f
C5881 commonsourceibias.n381 gnd 0.009606f
C5882 commonsourceibias.t108 gnd 0.179464f
C5883 commonsourceibias.n382 gnd 0.071606f
C5884 commonsourceibias.t130 gnd 0.179464f
C5885 commonsourceibias.n383 gnd 0.008572f
C5886 commonsourceibias.n384 gnd 0.009606f
C5887 commonsourceibias.t198 gnd 0.179464f
C5888 commonsourceibias.n385 gnd 0.011742f
C5889 commonsourceibias.n386 gnd 0.009606f
C5890 commonsourceibias.t186 gnd 0.179464f
C5891 commonsourceibias.n387 gnd 0.071606f
C5892 commonsourceibias.t92 gnd 0.179464f
C5893 commonsourceibias.n388 gnd 0.008375f
C5894 commonsourceibias.n389 gnd 0.009606f
C5895 commonsourceibias.t177 gnd 0.179464f
C5896 commonsourceibias.n390 gnd 0.011489f
C5897 commonsourceibias.n391 gnd 0.009606f
C5898 commonsourceibias.t170 gnd 0.179464f
C5899 commonsourceibias.n392 gnd 0.071606f
C5900 commonsourceibias.t81 gnd 0.179464f
C5901 commonsourceibias.n393 gnd 0.008208f
C5902 commonsourceibias.n394 gnd 0.009606f
C5903 commonsourceibias.t99 gnd 0.179464f
C5904 commonsourceibias.n395 gnd 0.011208f
C5905 commonsourceibias.t184 gnd 0.199531f
C5906 commonsourceibias.t151 gnd 0.179464f
C5907 commonsourceibias.n396 gnd 0.078223f
C5908 commonsourceibias.n397 gnd 0.08584f
C5909 commonsourceibias.n398 gnd 0.039831f
C5910 commonsourceibias.n399 gnd 0.009606f
C5911 commonsourceibias.n400 gnd 0.00935f
C5912 commonsourceibias.n401 gnd 0.013398f
C5913 commonsourceibias.n402 gnd 0.071606f
C5914 commonsourceibias.n403 gnd 0.013389f
C5915 commonsourceibias.n404 gnd 0.009606f
C5916 commonsourceibias.n405 gnd 0.009606f
C5917 commonsourceibias.n406 gnd 0.009606f
C5918 commonsourceibias.n407 gnd 0.012358f
C5919 commonsourceibias.n408 gnd 0.071606f
C5920 commonsourceibias.n409 gnd 0.012648f
C5921 commonsourceibias.n410 gnd 0.012289f
C5922 commonsourceibias.n411 gnd 0.009606f
C5923 commonsourceibias.n412 gnd 0.009606f
C5924 commonsourceibias.n413 gnd 0.009606f
C5925 commonsourceibias.n414 gnd 0.009057f
C5926 commonsourceibias.n415 gnd 0.01341f
C5927 commonsourceibias.n416 gnd 0.071606f
C5928 commonsourceibias.n417 gnd 0.013406f
C5929 commonsourceibias.n418 gnd 0.009606f
C5930 commonsourceibias.n419 gnd 0.009606f
C5931 commonsourceibias.n420 gnd 0.009606f
C5932 commonsourceibias.n421 gnd 0.012175f
C5933 commonsourceibias.n422 gnd 0.071606f
C5934 commonsourceibias.n423 gnd 0.012558f
C5935 commonsourceibias.n424 gnd 0.012378f
C5936 commonsourceibias.n425 gnd 0.009606f
C5937 commonsourceibias.n426 gnd 0.009606f
C5938 commonsourceibias.n427 gnd 0.009606f
C5939 commonsourceibias.n428 gnd 0.008798f
C5940 commonsourceibias.n429 gnd 0.013416f
C5941 commonsourceibias.n430 gnd 0.071606f
C5942 commonsourceibias.n431 gnd 0.013414f
C5943 commonsourceibias.n432 gnd 0.009606f
C5944 commonsourceibias.n433 gnd 0.009606f
C5945 commonsourceibias.n434 gnd 0.009606f
C5946 commonsourceibias.n435 gnd 0.01197f
C5947 commonsourceibias.n436 gnd 0.071606f
C5948 commonsourceibias.n437 gnd 0.012468f
C5949 commonsourceibias.n438 gnd 0.012468f
C5950 commonsourceibias.n439 gnd 0.009606f
C5951 commonsourceibias.n440 gnd 0.009606f
C5952 commonsourceibias.n441 gnd 0.009606f
C5953 commonsourceibias.n442 gnd 0.008572f
C5954 commonsourceibias.n443 gnd 0.013414f
C5955 commonsourceibias.n444 gnd 0.071606f
C5956 commonsourceibias.n445 gnd 0.013416f
C5957 commonsourceibias.n446 gnd 0.009606f
C5958 commonsourceibias.n447 gnd 0.009606f
C5959 commonsourceibias.n448 gnd 0.009606f
C5960 commonsourceibias.n449 gnd 0.011742f
C5961 commonsourceibias.n450 gnd 0.071606f
C5962 commonsourceibias.n451 gnd 0.012378f
C5963 commonsourceibias.n452 gnd 0.012558f
C5964 commonsourceibias.n453 gnd 0.009606f
C5965 commonsourceibias.n454 gnd 0.009606f
C5966 commonsourceibias.n455 gnd 0.009606f
C5967 commonsourceibias.n456 gnd 0.008375f
C5968 commonsourceibias.n457 gnd 0.013406f
C5969 commonsourceibias.n458 gnd 0.071606f
C5970 commonsourceibias.n459 gnd 0.01341f
C5971 commonsourceibias.n460 gnd 0.009606f
C5972 commonsourceibias.n461 gnd 0.009606f
C5973 commonsourceibias.n462 gnd 0.009606f
C5974 commonsourceibias.n463 gnd 0.011489f
C5975 commonsourceibias.n464 gnd 0.071606f
C5976 commonsourceibias.n465 gnd 0.012289f
C5977 commonsourceibias.n466 gnd 0.012648f
C5978 commonsourceibias.n467 gnd 0.009606f
C5979 commonsourceibias.n468 gnd 0.009606f
C5980 commonsourceibias.n469 gnd 0.009606f
C5981 commonsourceibias.n470 gnd 0.008208f
C5982 commonsourceibias.n471 gnd 0.013389f
C5983 commonsourceibias.n472 gnd 0.071606f
C5984 commonsourceibias.n473 gnd 0.013398f
C5985 commonsourceibias.n474 gnd 0.009606f
C5986 commonsourceibias.n475 gnd 0.009606f
C5987 commonsourceibias.n476 gnd 0.009606f
C5988 commonsourceibias.n477 gnd 0.011208f
C5989 commonsourceibias.n478 gnd 0.071606f
C5990 commonsourceibias.n479 gnd 0.011785f
C5991 commonsourceibias.t183 gnd 0.19409f
C5992 commonsourceibias.n480 gnd 0.085921f
C5993 commonsourceibias.n481 gnd 0.029883f
C5994 commonsourceibias.n482 gnd 0.5392f
C5995 commonsourceibias.n483 gnd 0.012818f
C5996 commonsourceibias.t191 gnd 0.19409f
C5997 commonsourceibias.t134 gnd 0.179464f
C5998 commonsourceibias.n484 gnd 0.00935f
C5999 commonsourceibias.n485 gnd 0.009606f
C6000 commonsourceibias.t97 gnd 0.179464f
C6001 commonsourceibias.n486 gnd 0.012358f
C6002 commonsourceibias.n487 gnd 0.009606f
C6003 commonsourceibias.t117 gnd 0.179464f
C6004 commonsourceibias.n488 gnd 0.009057f
C6005 commonsourceibias.n489 gnd 0.009606f
C6006 commonsourceibias.t187 gnd 0.179464f
C6007 commonsourceibias.n490 gnd 0.012175f
C6008 commonsourceibias.n491 gnd 0.009606f
C6009 commonsourceibias.t118 gnd 0.179464f
C6010 commonsourceibias.n492 gnd 0.008798f
C6011 commonsourceibias.n493 gnd 0.009606f
C6012 commonsourceibias.t149 gnd 0.179464f
C6013 commonsourceibias.n494 gnd 0.01197f
C6014 commonsourceibias.t23 gnd 0.020728f
C6015 commonsourceibias.t1 gnd 0.020728f
C6016 commonsourceibias.n495 gnd 0.183774f
C6017 commonsourceibias.t13 gnd 0.020728f
C6018 commonsourceibias.t35 gnd 0.020728f
C6019 commonsourceibias.n496 gnd 0.183161f
C6020 commonsourceibias.n497 gnd 0.170671f
C6021 commonsourceibias.t67 gnd 0.020728f
C6022 commonsourceibias.t65 gnd 0.020728f
C6023 commonsourceibias.n498 gnd 0.183161f
C6024 commonsourceibias.n499 gnd 0.084133f
C6025 commonsourceibias.t5 gnd 0.020728f
C6026 commonsourceibias.t61 gnd 0.020728f
C6027 commonsourceibias.n500 gnd 0.183161f
C6028 commonsourceibias.n501 gnd 0.084133f
C6029 commonsourceibias.t49 gnd 0.020728f
C6030 commonsourceibias.t71 gnd 0.020728f
C6031 commonsourceibias.n502 gnd 0.183161f
C6032 commonsourceibias.n503 gnd 0.070289f
C6033 commonsourceibias.n504 gnd 0.012818f
C6034 commonsourceibias.t58 gnd 0.179464f
C6035 commonsourceibias.n505 gnd 0.00935f
C6036 commonsourceibias.n506 gnd 0.009606f
C6037 commonsourceibias.t78 gnd 0.179464f
C6038 commonsourceibias.n507 gnd 0.012358f
C6039 commonsourceibias.n508 gnd 0.009606f
C6040 commonsourceibias.t30 gnd 0.179464f
C6041 commonsourceibias.n509 gnd 0.009057f
C6042 commonsourceibias.n510 gnd 0.009606f
C6043 commonsourceibias.t40 gnd 0.179464f
C6044 commonsourceibias.n511 gnd 0.012175f
C6045 commonsourceibias.n512 gnd 0.009606f
C6046 commonsourceibias.t28 gnd 0.179464f
C6047 commonsourceibias.n513 gnd 0.008798f
C6048 commonsourceibias.n514 gnd 0.009606f
C6049 commonsourceibias.t24 gnd 0.179464f
C6050 commonsourceibias.n515 gnd 0.01197f
C6051 commonsourceibias.n516 gnd 0.009606f
C6052 commonsourceibias.t70 gnd 0.179464f
C6053 commonsourceibias.n517 gnd 0.008572f
C6054 commonsourceibias.n518 gnd 0.009606f
C6055 commonsourceibias.t48 gnd 0.179464f
C6056 commonsourceibias.n519 gnd 0.011742f
C6057 commonsourceibias.n520 gnd 0.009606f
C6058 commonsourceibias.t4 gnd 0.179464f
C6059 commonsourceibias.n521 gnd 0.008375f
C6060 commonsourceibias.n522 gnd 0.009606f
C6061 commonsourceibias.t64 gnd 0.179464f
C6062 commonsourceibias.n523 gnd 0.011489f
C6063 commonsourceibias.n524 gnd 0.009606f
C6064 commonsourceibias.t34 gnd 0.179464f
C6065 commonsourceibias.n525 gnd 0.008208f
C6066 commonsourceibias.n526 gnd 0.009606f
C6067 commonsourceibias.t12 gnd 0.179464f
C6068 commonsourceibias.n527 gnd 0.011208f
C6069 commonsourceibias.t22 gnd 0.199531f
C6070 commonsourceibias.t0 gnd 0.179464f
C6071 commonsourceibias.n528 gnd 0.078223f
C6072 commonsourceibias.n529 gnd 0.08584f
C6073 commonsourceibias.n530 gnd 0.039831f
C6074 commonsourceibias.n531 gnd 0.009606f
C6075 commonsourceibias.n532 gnd 0.00935f
C6076 commonsourceibias.n533 gnd 0.013398f
C6077 commonsourceibias.n534 gnd 0.071606f
C6078 commonsourceibias.n535 gnd 0.013389f
C6079 commonsourceibias.n536 gnd 0.009606f
C6080 commonsourceibias.n537 gnd 0.009606f
C6081 commonsourceibias.n538 gnd 0.009606f
C6082 commonsourceibias.n539 gnd 0.012358f
C6083 commonsourceibias.n540 gnd 0.071606f
C6084 commonsourceibias.n541 gnd 0.012648f
C6085 commonsourceibias.t66 gnd 0.179464f
C6086 commonsourceibias.n542 gnd 0.071606f
C6087 commonsourceibias.n543 gnd 0.012289f
C6088 commonsourceibias.n544 gnd 0.009606f
C6089 commonsourceibias.n545 gnd 0.009606f
C6090 commonsourceibias.n546 gnd 0.009606f
C6091 commonsourceibias.n547 gnd 0.009057f
C6092 commonsourceibias.n548 gnd 0.01341f
C6093 commonsourceibias.n549 gnd 0.071606f
C6094 commonsourceibias.n550 gnd 0.013406f
C6095 commonsourceibias.n551 gnd 0.009606f
C6096 commonsourceibias.n552 gnd 0.009606f
C6097 commonsourceibias.n553 gnd 0.009606f
C6098 commonsourceibias.n554 gnd 0.012175f
C6099 commonsourceibias.n555 gnd 0.071606f
C6100 commonsourceibias.n556 gnd 0.012558f
C6101 commonsourceibias.t60 gnd 0.179464f
C6102 commonsourceibias.n557 gnd 0.071606f
C6103 commonsourceibias.n558 gnd 0.012378f
C6104 commonsourceibias.n559 gnd 0.009606f
C6105 commonsourceibias.n560 gnd 0.009606f
C6106 commonsourceibias.n561 gnd 0.009606f
C6107 commonsourceibias.n562 gnd 0.008798f
C6108 commonsourceibias.n563 gnd 0.013416f
C6109 commonsourceibias.n564 gnd 0.071606f
C6110 commonsourceibias.n565 gnd 0.013414f
C6111 commonsourceibias.n566 gnd 0.009606f
C6112 commonsourceibias.n567 gnd 0.009606f
C6113 commonsourceibias.n568 gnd 0.009606f
C6114 commonsourceibias.n569 gnd 0.01197f
C6115 commonsourceibias.n570 gnd 0.071606f
C6116 commonsourceibias.n571 gnd 0.012468f
C6117 commonsourceibias.t62 gnd 0.179464f
C6118 commonsourceibias.n572 gnd 0.071606f
C6119 commonsourceibias.n573 gnd 0.012468f
C6120 commonsourceibias.n574 gnd 0.009606f
C6121 commonsourceibias.n575 gnd 0.009606f
C6122 commonsourceibias.n576 gnd 0.009606f
C6123 commonsourceibias.n577 gnd 0.008572f
C6124 commonsourceibias.n578 gnd 0.013414f
C6125 commonsourceibias.n579 gnd 0.071606f
C6126 commonsourceibias.n580 gnd 0.013416f
C6127 commonsourceibias.n581 gnd 0.009606f
C6128 commonsourceibias.n582 gnd 0.009606f
C6129 commonsourceibias.n583 gnd 0.009606f
C6130 commonsourceibias.n584 gnd 0.011742f
C6131 commonsourceibias.n585 gnd 0.071606f
C6132 commonsourceibias.n586 gnd 0.012378f
C6133 commonsourceibias.t8 gnd 0.179464f
C6134 commonsourceibias.n587 gnd 0.071606f
C6135 commonsourceibias.n588 gnd 0.012558f
C6136 commonsourceibias.n589 gnd 0.009606f
C6137 commonsourceibias.n590 gnd 0.009606f
C6138 commonsourceibias.n591 gnd 0.009606f
C6139 commonsourceibias.n592 gnd 0.008375f
C6140 commonsourceibias.n593 gnd 0.013406f
C6141 commonsourceibias.n594 gnd 0.071606f
C6142 commonsourceibias.n595 gnd 0.01341f
C6143 commonsourceibias.n596 gnd 0.009606f
C6144 commonsourceibias.n597 gnd 0.009606f
C6145 commonsourceibias.n598 gnd 0.009606f
C6146 commonsourceibias.n599 gnd 0.011489f
C6147 commonsourceibias.n600 gnd 0.071606f
C6148 commonsourceibias.n601 gnd 0.012289f
C6149 commonsourceibias.t18 gnd 0.179464f
C6150 commonsourceibias.n602 gnd 0.071606f
C6151 commonsourceibias.n603 gnd 0.012648f
C6152 commonsourceibias.n604 gnd 0.009606f
C6153 commonsourceibias.n605 gnd 0.009606f
C6154 commonsourceibias.n606 gnd 0.009606f
C6155 commonsourceibias.n607 gnd 0.008208f
C6156 commonsourceibias.n608 gnd 0.013389f
C6157 commonsourceibias.n609 gnd 0.071606f
C6158 commonsourceibias.n610 gnd 0.013398f
C6159 commonsourceibias.n611 gnd 0.009606f
C6160 commonsourceibias.n612 gnd 0.009606f
C6161 commonsourceibias.n613 gnd 0.009606f
C6162 commonsourceibias.n614 gnd 0.011208f
C6163 commonsourceibias.n615 gnd 0.071606f
C6164 commonsourceibias.n616 gnd 0.011785f
C6165 commonsourceibias.t36 gnd 0.19409f
C6166 commonsourceibias.n617 gnd 0.085921f
C6167 commonsourceibias.n618 gnd 0.095704f
C6168 commonsourceibias.t59 gnd 0.020728f
C6169 commonsourceibias.t37 gnd 0.020728f
C6170 commonsourceibias.n619 gnd 0.183161f
C6171 commonsourceibias.n620 gnd 0.158435f
C6172 commonsourceibias.t19 gnd 0.020728f
C6173 commonsourceibias.t79 gnd 0.020728f
C6174 commonsourceibias.n621 gnd 0.183161f
C6175 commonsourceibias.n622 gnd 0.084133f
C6176 commonsourceibias.t41 gnd 0.020728f
C6177 commonsourceibias.t31 gnd 0.020728f
C6178 commonsourceibias.n623 gnd 0.183161f
C6179 commonsourceibias.n624 gnd 0.084133f
C6180 commonsourceibias.t29 gnd 0.020728f
C6181 commonsourceibias.t9 gnd 0.020728f
C6182 commonsourceibias.n625 gnd 0.183161f
C6183 commonsourceibias.n626 gnd 0.084133f
C6184 commonsourceibias.t63 gnd 0.020728f
C6185 commonsourceibias.t25 gnd 0.020728f
C6186 commonsourceibias.n627 gnd 0.183161f
C6187 commonsourceibias.n628 gnd 0.070289f
C6188 commonsourceibias.n629 gnd 0.085113f
C6189 commonsourceibias.n630 gnd 0.062168f
C6190 commonsourceibias.t105 gnd 0.179464f
C6191 commonsourceibias.n631 gnd 0.071606f
C6192 commonsourceibias.n632 gnd 0.009606f
C6193 commonsourceibias.t122 gnd 0.179464f
C6194 commonsourceibias.n633 gnd 0.071606f
C6195 commonsourceibias.n634 gnd 0.009606f
C6196 commonsourceibias.t115 gnd 0.179464f
C6197 commonsourceibias.n635 gnd 0.071606f
C6198 commonsourceibias.n636 gnd 0.009606f
C6199 commonsourceibias.t83 gnd 0.179464f
C6200 commonsourceibias.n637 gnd 0.008375f
C6201 commonsourceibias.n638 gnd 0.009606f
C6202 commonsourceibias.t111 gnd 0.179464f
C6203 commonsourceibias.n639 gnd 0.011489f
C6204 commonsourceibias.n640 gnd 0.009606f
C6205 commonsourceibias.t192 gnd 0.179464f
C6206 commonsourceibias.n641 gnd 0.008208f
C6207 commonsourceibias.n642 gnd 0.009606f
C6208 commonsourceibias.t127 gnd 0.179464f
C6209 commonsourceibias.n643 gnd 0.011208f
C6210 commonsourceibias.t153 gnd 0.199531f
C6211 commonsourceibias.t86 gnd 0.179464f
C6212 commonsourceibias.n644 gnd 0.078223f
C6213 commonsourceibias.n645 gnd 0.08584f
C6214 commonsourceibias.n646 gnd 0.039831f
C6215 commonsourceibias.n647 gnd 0.009606f
C6216 commonsourceibias.n648 gnd 0.00935f
C6217 commonsourceibias.n649 gnd 0.013398f
C6218 commonsourceibias.n650 gnd 0.071606f
C6219 commonsourceibias.n651 gnd 0.013389f
C6220 commonsourceibias.n652 gnd 0.009606f
C6221 commonsourceibias.n653 gnd 0.009606f
C6222 commonsourceibias.n654 gnd 0.009606f
C6223 commonsourceibias.n655 gnd 0.012358f
C6224 commonsourceibias.n656 gnd 0.071606f
C6225 commonsourceibias.n657 gnd 0.012648f
C6226 commonsourceibias.t110 gnd 0.179464f
C6227 commonsourceibias.n658 gnd 0.071606f
C6228 commonsourceibias.n659 gnd 0.012289f
C6229 commonsourceibias.n660 gnd 0.009606f
C6230 commonsourceibias.n661 gnd 0.009606f
C6231 commonsourceibias.n662 gnd 0.009606f
C6232 commonsourceibias.n663 gnd 0.009057f
C6233 commonsourceibias.n664 gnd 0.01341f
C6234 commonsourceibias.n665 gnd 0.071606f
C6235 commonsourceibias.n666 gnd 0.013406f
C6236 commonsourceibias.n667 gnd 0.009606f
C6237 commonsourceibias.n668 gnd 0.009606f
C6238 commonsourceibias.n669 gnd 0.009606f
C6239 commonsourceibias.n670 gnd 0.012175f
C6240 commonsourceibias.n671 gnd 0.071606f
C6241 commonsourceibias.n672 gnd 0.012558f
C6242 commonsourceibias.n673 gnd 0.012378f
C6243 commonsourceibias.n674 gnd 0.009606f
C6244 commonsourceibias.n675 gnd 0.009606f
C6245 commonsourceibias.n676 gnd 0.011742f
C6246 commonsourceibias.n677 gnd 0.008798f
C6247 commonsourceibias.n678 gnd 0.013416f
C6248 commonsourceibias.n679 gnd 0.009606f
C6249 commonsourceibias.n680 gnd 0.009606f
C6250 commonsourceibias.n681 gnd 0.013414f
C6251 commonsourceibias.n682 gnd 0.008572f
C6252 commonsourceibias.n683 gnd 0.01197f
C6253 commonsourceibias.n684 gnd 0.009606f
C6254 commonsourceibias.n685 gnd 0.008392f
C6255 commonsourceibias.n686 gnd 0.012468f
C6256 commonsourceibias.t114 gnd 0.179464f
C6257 commonsourceibias.n687 gnd 0.071606f
C6258 commonsourceibias.n688 gnd 0.012468f
C6259 commonsourceibias.n689 gnd 0.008392f
C6260 commonsourceibias.n690 gnd 0.009606f
C6261 commonsourceibias.n691 gnd 0.009606f
C6262 commonsourceibias.n692 gnd 0.008572f
C6263 commonsourceibias.n693 gnd 0.013414f
C6264 commonsourceibias.n694 gnd 0.071606f
C6265 commonsourceibias.n695 gnd 0.013416f
C6266 commonsourceibias.n696 gnd 0.009606f
C6267 commonsourceibias.n697 gnd 0.009606f
C6268 commonsourceibias.n698 gnd 0.009606f
C6269 commonsourceibias.n699 gnd 0.011742f
C6270 commonsourceibias.n700 gnd 0.071606f
C6271 commonsourceibias.n701 gnd 0.012378f
C6272 commonsourceibias.t132 gnd 0.179464f
C6273 commonsourceibias.n702 gnd 0.071606f
C6274 commonsourceibias.n703 gnd 0.012558f
C6275 commonsourceibias.n704 gnd 0.009606f
C6276 commonsourceibias.n705 gnd 0.009606f
C6277 commonsourceibias.n706 gnd 0.009606f
C6278 commonsourceibias.n707 gnd 0.008375f
C6279 commonsourceibias.n708 gnd 0.013406f
C6280 commonsourceibias.n709 gnd 0.071606f
C6281 commonsourceibias.n710 gnd 0.01341f
C6282 commonsourceibias.n711 gnd 0.009606f
C6283 commonsourceibias.n712 gnd 0.009606f
C6284 commonsourceibias.n713 gnd 0.009606f
C6285 commonsourceibias.n714 gnd 0.011489f
C6286 commonsourceibias.n715 gnd 0.071606f
C6287 commonsourceibias.n716 gnd 0.012289f
C6288 commonsourceibias.t152 gnd 0.179464f
C6289 commonsourceibias.n717 gnd 0.071606f
C6290 commonsourceibias.n718 gnd 0.012648f
C6291 commonsourceibias.n719 gnd 0.009606f
C6292 commonsourceibias.n720 gnd 0.009606f
C6293 commonsourceibias.n721 gnd 0.009606f
C6294 commonsourceibias.n722 gnd 0.008208f
C6295 commonsourceibias.n723 gnd 0.013389f
C6296 commonsourceibias.n724 gnd 0.071606f
C6297 commonsourceibias.n725 gnd 0.013398f
C6298 commonsourceibias.n726 gnd 0.009606f
C6299 commonsourceibias.n727 gnd 0.009606f
C6300 commonsourceibias.n728 gnd 0.009606f
C6301 commonsourceibias.n729 gnd 0.011208f
C6302 commonsourceibias.n730 gnd 0.071606f
C6303 commonsourceibias.n731 gnd 0.011785f
C6304 commonsourceibias.n732 gnd 0.085921f
C6305 commonsourceibias.n733 gnd 0.056157f
C6306 commonsourceibias.n734 gnd 0.012818f
C6307 commonsourceibias.t148 gnd 0.179464f
C6308 commonsourceibias.n735 gnd 0.00935f
C6309 commonsourceibias.n736 gnd 0.009606f
C6310 commonsourceibias.t139 gnd 0.179464f
C6311 commonsourceibias.n737 gnd 0.012358f
C6312 commonsourceibias.n738 gnd 0.009606f
C6313 commonsourceibias.t147 gnd 0.179464f
C6314 commonsourceibias.n739 gnd 0.009057f
C6315 commonsourceibias.n740 gnd 0.009606f
C6316 commonsourceibias.t138 gnd 0.179464f
C6317 commonsourceibias.n741 gnd 0.012175f
C6318 commonsourceibias.n742 gnd 0.009606f
C6319 commonsourceibias.t154 gnd 0.179464f
C6320 commonsourceibias.n743 gnd 0.008798f
C6321 commonsourceibias.n744 gnd 0.009606f
C6322 commonsourceibias.t137 gnd 0.179464f
C6323 commonsourceibias.n745 gnd 0.01197f
C6324 commonsourceibias.n746 gnd 0.009606f
C6325 commonsourceibias.t195 gnd 0.179464f
C6326 commonsourceibias.n747 gnd 0.008572f
C6327 commonsourceibias.n748 gnd 0.009606f
C6328 commonsourceibias.t135 gnd 0.179464f
C6329 commonsourceibias.n749 gnd 0.011742f
C6330 commonsourceibias.n750 gnd 0.009606f
C6331 commonsourceibias.t194 gnd 0.179464f
C6332 commonsourceibias.n751 gnd 0.008375f
C6333 commonsourceibias.n752 gnd 0.009606f
C6334 commonsourceibias.t176 gnd 0.179464f
C6335 commonsourceibias.n753 gnd 0.011489f
C6336 commonsourceibias.n754 gnd 0.009606f
C6337 commonsourceibias.t189 gnd 0.179464f
C6338 commonsourceibias.n755 gnd 0.008208f
C6339 commonsourceibias.n756 gnd 0.009606f
C6340 commonsourceibias.t180 gnd 0.179464f
C6341 commonsourceibias.n757 gnd 0.011208f
C6342 commonsourceibias.t188 gnd 0.199531f
C6343 commonsourceibias.t163 gnd 0.179464f
C6344 commonsourceibias.n758 gnd 0.078223f
C6345 commonsourceibias.n759 gnd 0.08584f
C6346 commonsourceibias.n760 gnd 0.039831f
C6347 commonsourceibias.n761 gnd 0.009606f
C6348 commonsourceibias.n762 gnd 0.00935f
C6349 commonsourceibias.n763 gnd 0.013398f
C6350 commonsourceibias.n764 gnd 0.071606f
C6351 commonsourceibias.n765 gnd 0.013389f
C6352 commonsourceibias.n766 gnd 0.009606f
C6353 commonsourceibias.n767 gnd 0.009606f
C6354 commonsourceibias.n768 gnd 0.009606f
C6355 commonsourceibias.n769 gnd 0.012358f
C6356 commonsourceibias.n770 gnd 0.071606f
C6357 commonsourceibias.n771 gnd 0.012648f
C6358 commonsourceibias.t164 gnd 0.179464f
C6359 commonsourceibias.n772 gnd 0.071606f
C6360 commonsourceibias.n773 gnd 0.012289f
C6361 commonsourceibias.n774 gnd 0.009606f
C6362 commonsourceibias.n775 gnd 0.009606f
C6363 commonsourceibias.n776 gnd 0.009606f
C6364 commonsourceibias.n777 gnd 0.009057f
C6365 commonsourceibias.n778 gnd 0.01341f
C6366 commonsourceibias.n779 gnd 0.071606f
C6367 commonsourceibias.n780 gnd 0.013406f
C6368 commonsourceibias.n781 gnd 0.009606f
C6369 commonsourceibias.n782 gnd 0.009606f
C6370 commonsourceibias.n783 gnd 0.009606f
C6371 commonsourceibias.n784 gnd 0.012175f
C6372 commonsourceibias.n785 gnd 0.071606f
C6373 commonsourceibias.n786 gnd 0.012558f
C6374 commonsourceibias.t171 gnd 0.179464f
C6375 commonsourceibias.n787 gnd 0.071606f
C6376 commonsourceibias.n788 gnd 0.012378f
C6377 commonsourceibias.n789 gnd 0.009606f
C6378 commonsourceibias.n790 gnd 0.009606f
C6379 commonsourceibias.n791 gnd 0.009606f
C6380 commonsourceibias.n792 gnd 0.008798f
C6381 commonsourceibias.n793 gnd 0.013416f
C6382 commonsourceibias.n794 gnd 0.071606f
C6383 commonsourceibias.n795 gnd 0.013414f
C6384 commonsourceibias.n796 gnd 0.009606f
C6385 commonsourceibias.n797 gnd 0.009606f
C6386 commonsourceibias.n798 gnd 0.009606f
C6387 commonsourceibias.n799 gnd 0.01197f
C6388 commonsourceibias.n800 gnd 0.071606f
C6389 commonsourceibias.n801 gnd 0.012468f
C6390 commonsourceibias.t161 gnd 0.179464f
C6391 commonsourceibias.n802 gnd 0.071606f
C6392 commonsourceibias.n803 gnd 0.012468f
C6393 commonsourceibias.n804 gnd 0.009606f
C6394 commonsourceibias.n805 gnd 0.009606f
C6395 commonsourceibias.n806 gnd 0.009606f
C6396 commonsourceibias.n807 gnd 0.008572f
C6397 commonsourceibias.n808 gnd 0.013414f
C6398 commonsourceibias.n809 gnd 0.071606f
C6399 commonsourceibias.n810 gnd 0.013416f
C6400 commonsourceibias.n811 gnd 0.009606f
C6401 commonsourceibias.n812 gnd 0.009606f
C6402 commonsourceibias.n813 gnd 0.009606f
C6403 commonsourceibias.n814 gnd 0.011742f
C6404 commonsourceibias.n815 gnd 0.071606f
C6405 commonsourceibias.n816 gnd 0.012378f
C6406 commonsourceibias.t162 gnd 0.179464f
C6407 commonsourceibias.n817 gnd 0.071606f
C6408 commonsourceibias.n818 gnd 0.012558f
C6409 commonsourceibias.n819 gnd 0.009606f
C6410 commonsourceibias.n820 gnd 0.009606f
C6411 commonsourceibias.n821 gnd 0.009606f
C6412 commonsourceibias.n822 gnd 0.008375f
C6413 commonsourceibias.n823 gnd 0.013406f
C6414 commonsourceibias.n824 gnd 0.071606f
C6415 commonsourceibias.n825 gnd 0.01341f
C6416 commonsourceibias.n826 gnd 0.009606f
C6417 commonsourceibias.n827 gnd 0.009606f
C6418 commonsourceibias.n828 gnd 0.009606f
C6419 commonsourceibias.n829 gnd 0.011489f
C6420 commonsourceibias.n830 gnd 0.071606f
C6421 commonsourceibias.n831 gnd 0.012289f
C6422 commonsourceibias.t128 gnd 0.179464f
C6423 commonsourceibias.n832 gnd 0.071606f
C6424 commonsourceibias.n833 gnd 0.012648f
C6425 commonsourceibias.n834 gnd 0.009606f
C6426 commonsourceibias.n835 gnd 0.009606f
C6427 commonsourceibias.n836 gnd 0.009606f
C6428 commonsourceibias.n837 gnd 0.008208f
C6429 commonsourceibias.n838 gnd 0.013389f
C6430 commonsourceibias.n839 gnd 0.071606f
C6431 commonsourceibias.n840 gnd 0.013398f
C6432 commonsourceibias.n841 gnd 0.009606f
C6433 commonsourceibias.n842 gnd 0.009606f
C6434 commonsourceibias.n843 gnd 0.009606f
C6435 commonsourceibias.n844 gnd 0.011208f
C6436 commonsourceibias.n845 gnd 0.071606f
C6437 commonsourceibias.n846 gnd 0.011785f
C6438 commonsourceibias.t129 gnd 0.19409f
C6439 commonsourceibias.n847 gnd 0.085921f
C6440 commonsourceibias.n848 gnd 0.029883f
C6441 commonsourceibias.n849 gnd 0.153513f
C6442 commonsourceibias.n850 gnd 0.012818f
C6443 commonsourceibias.t113 gnd 0.179464f
C6444 commonsourceibias.n851 gnd 0.00935f
C6445 commonsourceibias.n852 gnd 0.009606f
C6446 commonsourceibias.t125 gnd 0.179464f
C6447 commonsourceibias.n853 gnd 0.012358f
C6448 commonsourceibias.n854 gnd 0.009606f
C6449 commonsourceibias.t103 gnd 0.179464f
C6450 commonsourceibias.n855 gnd 0.009057f
C6451 commonsourceibias.n856 gnd 0.009606f
C6452 commonsourceibias.t120 gnd 0.179464f
C6453 commonsourceibias.n857 gnd 0.012175f
C6454 commonsourceibias.n858 gnd 0.009606f
C6455 commonsourceibias.t179 gnd 0.179464f
C6456 commonsourceibias.n859 gnd 0.008798f
C6457 commonsourceibias.n860 gnd 0.009606f
C6458 commonsourceibias.t112 gnd 0.179464f
C6459 commonsourceibias.n861 gnd 0.01197f
C6460 commonsourceibias.n862 gnd 0.009606f
C6461 commonsourceibias.t121 gnd 0.179464f
C6462 commonsourceibias.n863 gnd 0.008572f
C6463 commonsourceibias.n864 gnd 0.009606f
C6464 commonsourceibias.t102 gnd 0.179464f
C6465 commonsourceibias.n865 gnd 0.011742f
C6466 commonsourceibias.n866 gnd 0.009606f
C6467 commonsourceibias.t116 gnd 0.179464f
C6468 commonsourceibias.n867 gnd 0.008375f
C6469 commonsourceibias.n868 gnd 0.009606f
C6470 commonsourceibias.t167 gnd 0.179464f
C6471 commonsourceibias.n869 gnd 0.011489f
C6472 commonsourceibias.n870 gnd 0.009606f
C6473 commonsourceibias.t87 gnd 0.179464f
C6474 commonsourceibias.n871 gnd 0.008208f
C6475 commonsourceibias.n872 gnd 0.009606f
C6476 commonsourceibias.t106 gnd 0.179464f
C6477 commonsourceibias.n873 gnd 0.011208f
C6478 commonsourceibias.t196 gnd 0.199531f
C6479 commonsourceibias.t165 gnd 0.179464f
C6480 commonsourceibias.n874 gnd 0.078223f
C6481 commonsourceibias.n875 gnd 0.08584f
C6482 commonsourceibias.n876 gnd 0.039831f
C6483 commonsourceibias.n877 gnd 0.009606f
C6484 commonsourceibias.n878 gnd 0.00935f
C6485 commonsourceibias.n879 gnd 0.013398f
C6486 commonsourceibias.n880 gnd 0.071606f
C6487 commonsourceibias.n881 gnd 0.013389f
C6488 commonsourceibias.n882 gnd 0.009606f
C6489 commonsourceibias.n883 gnd 0.009606f
C6490 commonsourceibias.n884 gnd 0.009606f
C6491 commonsourceibias.n885 gnd 0.012358f
C6492 commonsourceibias.n886 gnd 0.071606f
C6493 commonsourceibias.n887 gnd 0.012648f
C6494 commonsourceibias.t178 gnd 0.179464f
C6495 commonsourceibias.n888 gnd 0.071606f
C6496 commonsourceibias.n889 gnd 0.012289f
C6497 commonsourceibias.n890 gnd 0.009606f
C6498 commonsourceibias.n891 gnd 0.009606f
C6499 commonsourceibias.n892 gnd 0.009606f
C6500 commonsourceibias.n893 gnd 0.009057f
C6501 commonsourceibias.n894 gnd 0.01341f
C6502 commonsourceibias.n895 gnd 0.071606f
C6503 commonsourceibias.n896 gnd 0.013406f
C6504 commonsourceibias.n897 gnd 0.009606f
C6505 commonsourceibias.n898 gnd 0.009606f
C6506 commonsourceibias.n899 gnd 0.009606f
C6507 commonsourceibias.n900 gnd 0.012175f
C6508 commonsourceibias.n901 gnd 0.071606f
C6509 commonsourceibias.n902 gnd 0.012558f
C6510 commonsourceibias.t96 gnd 0.179464f
C6511 commonsourceibias.n903 gnd 0.071606f
C6512 commonsourceibias.n904 gnd 0.012378f
C6513 commonsourceibias.n905 gnd 0.009606f
C6514 commonsourceibias.n906 gnd 0.009606f
C6515 commonsourceibias.n907 gnd 0.009606f
C6516 commonsourceibias.n908 gnd 0.008798f
C6517 commonsourceibias.n909 gnd 0.013416f
C6518 commonsourceibias.n910 gnd 0.071606f
C6519 commonsourceibias.n911 gnd 0.013414f
C6520 commonsourceibias.n912 gnd 0.009606f
C6521 commonsourceibias.n913 gnd 0.009606f
C6522 commonsourceibias.n914 gnd 0.009606f
C6523 commonsourceibias.n915 gnd 0.01197f
C6524 commonsourceibias.n916 gnd 0.071606f
C6525 commonsourceibias.n917 gnd 0.012468f
C6526 commonsourceibias.t126 gnd 0.179464f
C6527 commonsourceibias.n918 gnd 0.071606f
C6528 commonsourceibias.n919 gnd 0.012468f
C6529 commonsourceibias.n920 gnd 0.009606f
C6530 commonsourceibias.n921 gnd 0.009606f
C6531 commonsourceibias.n922 gnd 0.009606f
C6532 commonsourceibias.n923 gnd 0.008572f
C6533 commonsourceibias.n924 gnd 0.013414f
C6534 commonsourceibias.n925 gnd 0.071606f
C6535 commonsourceibias.n926 gnd 0.013416f
C6536 commonsourceibias.n927 gnd 0.009606f
C6537 commonsourceibias.n928 gnd 0.009606f
C6538 commonsourceibias.n929 gnd 0.009606f
C6539 commonsourceibias.n930 gnd 0.011742f
C6540 commonsourceibias.n931 gnd 0.071606f
C6541 commonsourceibias.n932 gnd 0.012378f
C6542 commonsourceibias.t133 gnd 0.179464f
C6543 commonsourceibias.n933 gnd 0.071606f
C6544 commonsourceibias.n934 gnd 0.012558f
C6545 commonsourceibias.n935 gnd 0.009606f
C6546 commonsourceibias.n936 gnd 0.009606f
C6547 commonsourceibias.n937 gnd 0.009606f
C6548 commonsourceibias.n938 gnd 0.008375f
C6549 commonsourceibias.n939 gnd 0.013406f
C6550 commonsourceibias.n940 gnd 0.071606f
C6551 commonsourceibias.n941 gnd 0.01341f
C6552 commonsourceibias.n942 gnd 0.009606f
C6553 commonsourceibias.n943 gnd 0.009606f
C6554 commonsourceibias.n944 gnd 0.009606f
C6555 commonsourceibias.n945 gnd 0.011489f
C6556 commonsourceibias.n946 gnd 0.071606f
C6557 commonsourceibias.n947 gnd 0.012289f
C6558 commonsourceibias.t85 gnd 0.179464f
C6559 commonsourceibias.n948 gnd 0.071606f
C6560 commonsourceibias.n949 gnd 0.012648f
C6561 commonsourceibias.n950 gnd 0.009606f
C6562 commonsourceibias.n951 gnd 0.009606f
C6563 commonsourceibias.n952 gnd 0.009606f
C6564 commonsourceibias.n953 gnd 0.008208f
C6565 commonsourceibias.n954 gnd 0.013389f
C6566 commonsourceibias.n955 gnd 0.071606f
C6567 commonsourceibias.n956 gnd 0.013398f
C6568 commonsourceibias.n957 gnd 0.009606f
C6569 commonsourceibias.n958 gnd 0.009606f
C6570 commonsourceibias.n959 gnd 0.009606f
C6571 commonsourceibias.n960 gnd 0.011208f
C6572 commonsourceibias.n961 gnd 0.071606f
C6573 commonsourceibias.n962 gnd 0.011785f
C6574 commonsourceibias.t93 gnd 0.19409f
C6575 commonsourceibias.n963 gnd 0.085921f
C6576 commonsourceibias.n964 gnd 0.029883f
C6577 commonsourceibias.n965 gnd 0.202576f
C6578 commonsourceibias.n966 gnd 5.69738f
.ends

