* NGSPICE file created from opamp136.ext - technology: sky130A

.subckt opamp136 gnd CSoutput output vdd plus minus commonsourceibias outputibias
+ diffpairibias
X0 gnd.t350 commonsourceibias.t2 commonsourceibias.t3 gnd.t274 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X1 CSoutput.t95 a_n6972_8799.t36 vdd.t171 vdd.t123 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X2 a_n1808_13878.t11 a_n2848_n452.t17 a_n2848_n452.t18 vdd.t22 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X3 a_n1808_13878.t19 a_n2848_n452.t48 vdd.t263 vdd.t262 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X4 CSoutput.t191 commonsourceibias.t64 gnd.t349 gnd.t243 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=2.73 ps=14.78 w=7 l=1
X5 vdd.t170 a_n6972_8799.t37 CSoutput.t94 vdd.t116 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X6 CSoutput.t93 a_n6972_8799.t38 vdd.t169 vdd.t52 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X7 vdd.t247 vdd.t245 vdd.t246 vdd.t181 sky130_fd_pr__pfet_01v8 ad=3.12 pd=16.78 as=0 ps=0 w=8 l=0.5
X8 commonsourceibias.t1 commonsourceibias.t0 gnd.t348 gnd.t215 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X9 gnd.t347 commonsourceibias.t65 CSoutput.t190 gnd.t203 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X10 a_n6972_8799.t22 plus.t5 a_n3827_n3924.t57 gnd.t64 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.9
X11 gnd.t346 commonsourceibias.t36 commonsourceibias.t37 gnd.t211 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X12 a_n3827_n3924.t13 diffpairibias.t20 gnd.t48 gnd.t47 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=2.73 ps=14.78 w=7 l=1
X13 a_n3827_n3924.t56 plus.t6 a_n6972_8799.t0 gnd.t9 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.9
X14 CSoutput.t92 a_n6972_8799.t39 vdd.t166 vdd.t54 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X15 gnd.t345 commonsourceibias.t34 commonsourceibias.t35 gnd.t191 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X16 a_n1986_8322.t11 a_n2848_n452.t49 a_n6972_8799.t35 vdd.t39 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X17 commonsourceibias.t33 commonsourceibias.t32 gnd.t344 gnd.t233 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X18 gnd.t343 commonsourceibias.t66 CSoutput.t189 gnd.t267 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X19 CSoutput.t91 a_n6972_8799.t40 vdd.t168 vdd.t87 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X20 vdd.t167 a_n6972_8799.t41 CSoutput.t90 vdd.t110 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X21 gnd.t190 gnd.t188 gnd.t189 gnd.t121 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=0 ps=0 w=7 l=1
X22 a_n2848_n452.t32 minus.t5 a_n3827_n3924.t14 gnd.t11 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.9
X23 gnd.t187 gnd.t184 gnd.t186 gnd.t185 sky130_fd_pr__nfet_01v8 ad=2.34 pd=12.78 as=0 ps=0 w=6 l=2
X24 a_n6972_8799.t26 plus.t7 a_n3827_n3924.t55 gnd.t13 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.9
X25 a_n2848_n452.t42 minus.t6 a_n3827_n3924.t27 gnd.t67 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.9
X26 plus.t4 gnd.t181 gnd.t183 gnd.t182 sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.5
X27 vdd.t165 a_n6972_8799.t42 CSoutput.t89 vdd.t132 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X28 CSoutput.t88 a_n6972_8799.t43 vdd.t164 vdd.t89 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X29 commonsourceibias.t31 commonsourceibias.t30 gnd.t342 gnd.t272 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X30 vdd.t162 a_n6972_8799.t44 CSoutput.t87 vdd.t151 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X31 a_n6972_8799.t11 a_n2848_n452.t50 a_n1986_8322.t10 vdd.t12 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=3.51 ps=18.78 w=9 l=0.5
X32 CSoutput.t86 a_n6972_8799.t45 vdd.t163 vdd.t50 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=3.12 ps=16.78 w=8 l=0.5
X33 gnd.t341 commonsourceibias.t67 CSoutput.t188 gnd.t207 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X34 CSoutput.t187 commonsourceibias.t68 gnd.t340 gnd.t222 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X35 gnd.t339 commonsourceibias.t28 commonsourceibias.t29 gnd.t267 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X36 CSoutput.t192 a_n1986_8322.t20 sky130_fd_pr__cap_mim_m3_1 l=12 w=12
X37 CSoutput.t186 commonsourceibias.t69 gnd.t338 gnd.t277 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X38 CSoutput.t85 a_n6972_8799.t46 vdd.t161 vdd.t123 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X39 a_n3827_n3924.t54 plus.t8 a_n6972_8799.t14 gnd.t38 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.9
X40 vdd.t244 vdd.t242 vdd.t243 vdd.t177 sky130_fd_pr__pfet_01v8 ad=3.12 pd=16.78 as=0 ps=0 w=8 l=0.5
X41 a_n3827_n3924.t22 diffpairibias.t21 gnd.t63 gnd.t62 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=2.73 ps=14.78 w=7 l=1
X42 CSoutput.t84 a_n6972_8799.t47 vdd.t160 vdd.t81 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X43 commonsourceibias.t27 commonsourceibias.t26 gnd.t337 gnd.t197 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X44 a_n3827_n3924.t9 minus.t7 a_n2848_n452.t28 gnd.t28 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.9
X45 vdd.t241 vdd.t239 vdd.t240 vdd.t181 sky130_fd_pr__pfet_01v8 ad=3.12 pd=16.78 as=0 ps=0 w=8 l=0.5
X46 CSoutput.t185 commonsourceibias.t70 gnd.t336 gnd.t277 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X47 CSoutput.t83 a_n6972_8799.t48 vdd.t159 vdd.t54 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X48 gnd.t335 commonsourceibias.t24 commonsourceibias.t25 gnd.t261 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X49 CSoutput.t184 commonsourceibias.t71 gnd.t334 gnd.t209 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=2.73 ps=14.78 w=7 l=1
X50 a_n1808_13878.t10 a_n2848_n452.t21 a_n2848_n452.t22 vdd.t0 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=3.51 ps=18.78 w=9 l=0.5
X51 vdd.t158 a_n6972_8799.t49 CSoutput.t82 vdd.t151 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X52 CSoutput.t81 a_n6972_8799.t50 vdd.t157 vdd.t114 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X53 a_n2848_n452.t8 a_n2848_n452.t7 a_n1808_13878.t9 vdd.t13 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X54 output.t3 outputibias.t8 gnd.t366 gnd.t365 sky130_fd_pr__nfet_01v8 ad=2.34 pd=12.78 as=2.34 ps=12.78 w=6 l=2
X55 CSoutput.t193 a_n1986_8322.t21 sky130_fd_pr__cap_mim_m3_1 l=12 w=12
X56 gnd.t180 gnd.t178 gnd.t179 gnd.t107 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=0 ps=0 w=7 l=0.9
X57 CSoutput.t80 a_n6972_8799.t51 vdd.t156 vdd.t87 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X58 vdd.t238 vdd.t236 vdd.t237 vdd.t212 sky130_fd_pr__pfet_01v8 ad=3.51 pd=18.78 as=0 ps=0 w=9 l=0.5
X59 a_n3827_n3924.t53 plus.t9 a_n6972_8799.t7 gnd.t24 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.9
X60 vdd.t155 a_n6972_8799.t52 CSoutput.t79 vdd.t110 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X61 vdd.t30 CSoutput.t194 output.t19 gnd.t41 sky130_fd_pr__nfet_01v8 ad=0.825 pd=5.33 as=0.825 ps=5.33 w=5 l=1
X62 diffpairibias.t19 diffpairibias.t18 gnd.t1 gnd.t0 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=2.73 ps=14.78 w=7 l=1
X63 CSoutput.t183 commonsourceibias.t72 gnd.t333 gnd.t241 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X64 a_n3827_n3924.t52 plus.t10 a_n6972_8799.t15 gnd.t31 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.9
X65 a_n3827_n3924.t11 minus.t8 a_n2848_n452.t30 gnd.t36 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=1.155 ps=7.33 w=7 l=0.9
X66 CSoutput.t182 commonsourceibias.t73 gnd.t332 gnd.t195 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X67 CSoutput.t181 commonsourceibias.t74 gnd.t331 gnd.t259 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X68 CSoutput.t78 a_n6972_8799.t53 vdd.t154 vdd.t118 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X69 commonsourceibias.t53 commonsourceibias.t52 gnd.t330 gnd.t243 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=2.73 ps=14.78 w=7 l=1
X70 gnd.t177 gnd.t175 gnd.t176 gnd.t78 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=0 ps=0 w=7 l=1
X71 vdd.t153 a_n6972_8799.t54 CSoutput.t77 vdd.t62 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X72 vdd.t152 a_n6972_8799.t55 CSoutput.t76 vdd.t151 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X73 vdd.t150 a_n6972_8799.t56 CSoutput.t75 vdd.t107 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X74 diffpairibias.t17 diffpairibias.t16 gnd.t46 gnd.t45 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=2.73 ps=14.78 w=7 l=1
X75 CSoutput.t74 a_n6972_8799.t57 vdd.t149 vdd.t50 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=3.12 ps=16.78 w=8 l=0.5
X76 CSoutput.t73 a_n6972_8799.t58 vdd.t148 vdd.t69 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=3.12 ps=16.78 w=8 l=0.5
X77 gnd.t174 gnd.t172 gnd.t173 gnd.t78 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=0 ps=0 w=7 l=1
X78 vdd.t147 a_n6972_8799.t59 CSoutput.t72 vdd.t48 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X79 CSoutput.t180 commonsourceibias.t75 gnd.t329 gnd.t259 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X80 CSoutput.t71 a_n6972_8799.t60 vdd.t146 vdd.t121 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X81 CSoutput.t70 a_n6972_8799.t61 vdd.t145 vdd.t81 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X82 CSoutput.t69 a_n6972_8799.t62 vdd.t122 vdd.t121 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X83 a_n3827_n3924.t21 minus.t9 a_n2848_n452.t38 gnd.t51 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.9
X84 a_n3827_n3924.t51 plus.t11 a_n6972_8799.t20 gnd.t27 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=1.155 ps=7.33 w=7 l=0.9
X85 vdd.t144 a_n6972_8799.t63 CSoutput.t68 vdd.t134 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X86 gnd.t328 commonsourceibias.t76 CSoutput.t179 gnd.t239 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X87 gnd.t171 gnd.t168 gnd.t170 gnd.t169 sky130_fd_pr__nfet_01v8 ad=2.34 pd=12.78 as=0 ps=0 w=6 l=2
X88 CSoutput.t178 commonsourceibias.t77 gnd.t327 gnd.t255 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X89 a_n6972_8799.t1 plus.t12 a_n3827_n3924.t50 gnd.t10 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.9
X90 gnd.t326 commonsourceibias.t78 CSoutput.t177 gnd.t218 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=1.155 ps=7.33 w=7 l=1
X91 gnd.t167 gnd.t165 gnd.t166 gnd.t121 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=0 ps=0 w=7 l=1
X92 a_n3827_n3924.t0 diffpairibias.t22 gnd.t3 gnd.t2 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=2.73 ps=14.78 w=7 l=1
X93 CSoutput.t176 commonsourceibias.t79 gnd.t325 gnd.t201 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X94 a_n2848_n452.t12 a_n2848_n452.t11 a_n1808_13878.t8 vdd.t39 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X95 vdd.t143 a_n6972_8799.t64 CSoutput.t67 vdd.t91 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X96 a_n3827_n3924.t49 plus.t13 a_n6972_8799.t30 gnd.t54 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.9
X97 a_n6972_8799.t12 a_n2848_n452.t51 a_n1986_8322.t9 vdd.t25 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X98 vdd.t142 a_n6972_8799.t65 CSoutput.t66 vdd.t132 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X99 a_n2848_n452.t10 a_n2848_n452.t9 a_n1808_13878.t7 vdd.t23 sky130_fd_pr__pfet_01v8 ad=3.51 pd=18.78 as=1.485 ps=9.33 w=9 l=0.5
X100 vdd.t138 a_n6972_8799.t66 CSoutput.t65 vdd.t134 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X101 outputibias.t7 outputibias.t6 gnd.t44 gnd.t43 sky130_fd_pr__nfet_01v8 ad=2.34 pd=12.78 as=2.34 ps=12.78 w=6 l=2
X102 commonsourceibias.t51 commonsourceibias.t50 gnd.t324 gnd.t222 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X103 gnd.t323 commonsourceibias.t80 CSoutput.t175 gnd.t236 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X104 gnd.t164 gnd.t162 gnd.t163 gnd.t85 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=0 ps=0 w=7 l=1
X105 CSoutput.t174 commonsourceibias.t81 gnd.t322 gnd.t215 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X106 gnd.t321 commonsourceibias.t48 commonsourceibias.t49 gnd.t220 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X107 vdd.t141 a_n6972_8799.t67 CSoutput.t64 vdd.t66 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X108 CSoutput.t173 commonsourceibias.t82 gnd.t320 gnd.t277 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X109 CSoutput.t63 a_n6972_8799.t68 vdd.t140 vdd.t94 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X110 a_n2848_n452.t33 minus.t10 a_n3827_n3924.t15 gnd.t37 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=2.73 ps=14.78 w=7 l=0.9
X111 diffpairibias.t15 diffpairibias.t14 gnd.t356 gnd.t355 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=2.73 ps=14.78 w=7 l=1
X112 vdd.t235 vdd.t233 vdd.t234 vdd.t220 sky130_fd_pr__pfet_01v8 ad=3.51 pd=18.78 as=0 ps=0 w=9 l=0.5
X113 vdd.t139 a_n6972_8799.t69 CSoutput.t62 vdd.t107 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X114 CSoutput.t61 a_n6972_8799.t70 vdd.t137 vdd.t69 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=3.12 ps=16.78 w=8 l=0.5
X115 vdd.t232 vdd.t229 vdd.t231 vdd.t230 sky130_fd_pr__pfet_01v8 ad=3.51 pd=18.78 as=0 ps=0 w=9 l=0.5
X116 gnd.t319 commonsourceibias.t83 CSoutput.t172 gnd.t226 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=1.155 ps=7.33 w=7 l=1
X117 vdd.t228 vdd.t226 vdd.t227 vdd.t173 sky130_fd_pr__pfet_01v8 ad=3.51 pd=18.78 as=0 ps=0 w=9 l=0.5
X118 vdd.t225 vdd.t223 vdd.t224 vdd.t216 sky130_fd_pr__pfet_01v8 ad=3.51 pd=18.78 as=0 ps=0 w=9 l=0.5
X119 vdd.t9 a_n2848_n452.t52 a_n1986_8322.t19 vdd.t8 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X120 gnd.t318 commonsourceibias.t46 commonsourceibias.t47 gnd.t213 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X121 CSoutput.t171 commonsourceibias.t84 gnd.t317 gnd.t229 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X122 output.t18 CSoutput.t195 vdd.t252 gnd.t359 sky130_fd_pr__nfet_01v8 ad=0.825 pd=5.33 as=0.825 ps=5.33 w=5 l=1
X123 CSoutput.t170 commonsourceibias.t85 gnd.t316 gnd.t272 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X124 a_n1986_8322.t18 a_n2848_n452.t53 vdd.t11 vdd.t10 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X125 a_n3827_n3924.t23 diffpairibias.t23 gnd.t66 gnd.t65 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=2.73 ps=14.78 w=7 l=1
X126 CSoutput.t60 a_n6972_8799.t71 vdd.t136 vdd.t121 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X127 gnd.t315 commonsourceibias.t86 CSoutput.t169 gnd.t274 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X128 gnd.t161 gnd.t159 gnd.t160 gnd.t103 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=0 ps=0 w=7 l=0.9
X129 gnd.t158 gnd.t156 minus.t4 gnd.t157 sky130_fd_pr__nfet_01v8 ad=0.39 pd=2.78 as=0.165 ps=1.33 w=1 l=0.5
X130 vdd.t135 a_n6972_8799.t72 CSoutput.t59 vdd.t134 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X131 commonsourceibias.t45 commonsourceibias.t44 gnd.t314 gnd.t209 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=2.73 ps=14.78 w=7 l=1
X132 vdd.t5 a_n2848_n452.t54 a_n1808_13878.t18 vdd.t4 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X133 gnd.t311 commonsourceibias.t87 CSoutput.t168 gnd.t193 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X134 vdd.t222 vdd.t219 vdd.t221 vdd.t220 sky130_fd_pr__pfet_01v8 ad=3.51 pd=18.78 as=0 ps=0 w=9 l=0.5
X135 gnd.t313 commonsourceibias.t42 commonsourceibias.t43 gnd.t207 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X136 output.t17 CSoutput.t196 vdd.t253 gnd.t360 sky130_fd_pr__nfet_01v8 ad=0.825 pd=5.33 as=0.825 ps=5.33 w=5 l=1
X137 CSoutput.t167 commonsourceibias.t88 gnd.t312 gnd.t241 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X138 gnd.t310 commonsourceibias.t89 CSoutput.t166 gnd.t203 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X139 vdd.t218 vdd.t215 vdd.t217 vdd.t216 sky130_fd_pr__pfet_01v8 ad=3.51 pd=18.78 as=0 ps=0 w=9 l=0.5
X140 vdd.t133 a_n6972_8799.t73 CSoutput.t58 vdd.t132 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X141 gnd.t155 gnd.t153 plus.t3 gnd.t154 sky130_fd_pr__nfet_01v8 ad=0.39 pd=2.78 as=0.165 ps=1.33 w=1 l=0.5
X142 CSoutput.t165 commonsourceibias.t90 gnd.t309 gnd.t255 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X143 a_n6972_8799.t8 plus.t14 a_n3827_n3924.t48 gnd.t25 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=2.73 ps=14.78 w=7 l=0.9
X144 commonsourceibias.t41 commonsourceibias.t40 gnd.t308 gnd.t199 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X145 a_n2848_n452.t37 minus.t11 a_n3827_n3924.t19 gnd.t56 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.9
X146 vdd.t214 vdd.t211 vdd.t213 vdd.t212 sky130_fd_pr__pfet_01v8 ad=3.51 pd=18.78 as=0 ps=0 w=9 l=0.5
X147 a_n1986_8322.t17 a_n2848_n452.t55 vdd.t7 vdd.t6 sky130_fd_pr__pfet_01v8 ad=3.51 pd=18.78 as=1.485 ps=9.33 w=9 l=0.5
X148 a_n6972_8799.t5 a_n2848_n452.t56 a_n1986_8322.t8 vdd.t21 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X149 gnd.t307 commonsourceibias.t91 CSoutput.t164 gnd.t224 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X150 a_n6972_8799.t31 plus.t15 a_n3827_n3924.t47 gnd.t55 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.9
X151 gnd.t152 gnd.t150 gnd.t151 gnd.t96 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=0 ps=0 w=7 l=1
X152 diffpairibias.t13 diffpairibias.t12 gnd.t15 gnd.t14 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=2.73 ps=14.78 w=7 l=1
X153 a_n2848_n452.t47 minus.t12 a_n3827_n3924.t33 gnd.t369 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.9
X154 a_n2848_n452.t6 a_n2848_n452.t5 a_n1808_13878.t6 vdd.t1 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X155 vdd.t131 a_n6972_8799.t74 CSoutput.t57 vdd.t66 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X156 a_n6972_8799.t6 a_n2848_n452.t57 a_n1986_8322.t7 vdd.t22 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X157 CSoutput.t56 a_n6972_8799.t75 vdd.t130 vdd.t94 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X158 gnd.t306 commonsourceibias.t38 commonsourceibias.t39 gnd.t203 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X159 a_n1808_13878.t5 a_n2848_n452.t15 a_n2848_n452.t16 vdd.t25 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X160 gnd.t305 commonsourceibias.t92 CSoutput.t163 gnd.t231 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X161 output.t16 CSoutput.t197 vdd.t28 gnd.t39 sky130_fd_pr__nfet_01v8 ad=0.825 pd=5.33 as=0.825 ps=5.33 w=5 l=1
X162 gnd.t304 commonsourceibias.t93 CSoutput.t162 gnd.t213 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X163 a_n3827_n3924.t29 minus.t13 a_n2848_n452.t43 gnd.t29 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.9
X164 CSoutput.t55 a_n6972_8799.t76 vdd.t129 vdd.t118 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X165 vdd.t33 a_n2848_n452.t58 a_n1986_8322.t16 vdd.t32 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=3.51 ps=18.78 w=9 l=0.5
X166 gnd.t149 gnd.t147 gnd.t148 gnd.t96 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=0 ps=0 w=7 l=1
X167 vdd.t128 a_n6972_8799.t77 CSoutput.t54 vdd.t116 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X168 output.t2 outputibias.t9 gnd.t371 gnd.t370 sky130_fd_pr__nfet_01v8 ad=2.34 pd=12.78 as=2.34 ps=12.78 w=6 l=2
X169 a_n2848_n452.t44 minus.t14 a_n3827_n3924.t30 gnd.t64 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.9
X170 a_n3827_n3924.t46 plus.t16 a_n6972_8799.t18 gnd.t6 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.9
X171 gnd.t146 gnd.t143 gnd.t145 gnd.t144 sky130_fd_pr__nfet_01v8 ad=1.95 pd=10.78 as=0 ps=0 w=5 l=1
X172 gnd.t142 gnd.t140 gnd.t141 gnd.t121 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=0 ps=0 w=7 l=1
X173 CSoutput.t53 a_n6972_8799.t78 vdd.t127 vdd.t114 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X174 outputibias.t5 outputibias.t4 gnd.t373 gnd.t372 sky130_fd_pr__nfet_01v8 ad=2.34 pd=12.78 as=2.34 ps=12.78 w=6 l=2
X175 vdd.t29 CSoutput.t198 output.t15 gnd.t40 sky130_fd_pr__nfet_01v8 ad=0.825 pd=5.33 as=0.825 ps=5.33 w=5 l=1
X176 vdd.t125 a_n6972_8799.t79 CSoutput.t52 vdd.t46 sky130_fd_pr__pfet_01v8 ad=3.12 pd=16.78 as=1.32 ps=8.33 w=8 l=0.5
X177 CSoutput.t161 commonsourceibias.t94 gnd.t303 gnd.t201 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X178 gnd.t302 commonsourceibias.t95 CSoutput.t160 gnd.t239 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X179 gnd.t301 commonsourceibias.t96 CSoutput.t159 gnd.t236 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X180 a_n3827_n3924.t1 diffpairibias.t24 gnd.t5 gnd.t4 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=2.73 ps=14.78 w=7 l=1
X181 a_n3827_n3924.t6 diffpairibias.t25 gnd.t17 gnd.t16 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=2.73 ps=14.78 w=7 l=1
X182 outputibias.t3 outputibias.t2 gnd.t34 gnd.t33 sky130_fd_pr__nfet_01v8 ad=2.34 pd=12.78 as=2.34 ps=12.78 w=6 l=2
X183 a_n6972_8799.t23 plus.t17 a_n3827_n3924.t45 gnd.t12 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.9
X184 vdd.t126 a_n6972_8799.t80 CSoutput.t51 vdd.t79 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X185 gnd.t139 gnd.t137 gnd.t138 gnd.t85 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=0 ps=0 w=7 l=1
X186 a_n6972_8799.t24 plus.t18 a_n3827_n3924.t44 gnd.t67 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.9
X187 gnd.t136 gnd.t134 gnd.t135 gnd.t85 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=0 ps=0 w=7 l=1
X188 CSoutput.t50 a_n6972_8799.t81 vdd.t124 vdd.t123 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X189 vdd.t14 CSoutput.t199 output.t14 gnd.t20 sky130_fd_pr__nfet_01v8 ad=0.825 pd=5.33 as=0.825 ps=5.33 w=5 l=1
X190 minus.t3 gnd.t131 gnd.t133 gnd.t132 sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.5
X191 CSoutput.t49 a_n6972_8799.t82 vdd.t120 vdd.t102 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X192 CSoutput.t158 commonsourceibias.t97 gnd.t300 gnd.t195 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X193 output.t13 CSoutput.t200 vdd.t15 gnd.t21 sky130_fd_pr__nfet_01v8 ad=0.825 pd=5.33 as=0.825 ps=5.33 w=5 l=1
X194 gnd.t130 gnd.t128 gnd.t129 gnd.t78 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=0 ps=0 w=7 l=1
X195 gnd.t194 commonsourceibias.t98 CSoutput.t157 gnd.t193 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X196 diffpairibias.t11 diffpairibias.t10 gnd.t53 gnd.t52 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=2.73 ps=14.78 w=7 l=1
X197 a_n1808_13878.t17 a_n2848_n452.t59 vdd.t35 vdd.t34 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X198 vdd.t210 vdd.t208 vdd.t209 vdd.t192 sky130_fd_pr__pfet_01v8 ad=3.12 pd=16.78 as=0 ps=0 w=8 l=0.5
X199 a_n2848_n452.t46 minus.t15 a_n3827_n3924.t32 gnd.t42 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.9
X200 vdd.t37 a_n2848_n452.t60 a_n1808_13878.t16 vdd.t36 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X201 CSoutput.t48 a_n6972_8799.t83 vdd.t119 vdd.t118 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X202 gnd.t299 commonsourceibias.t99 CSoutput.t156 gnd.t267 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X203 CSoutput.t155 commonsourceibias.t100 gnd.t298 gnd.t209 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=2.73 ps=14.78 w=7 l=1
X204 a_n3827_n3924.t43 plus.t19 a_n6972_8799.t25 gnd.t28 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.9
X205 vdd.t117 a_n6972_8799.t84 CSoutput.t47 vdd.t116 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X206 output.t12 CSoutput.t201 vdd.t40 gnd.t59 sky130_fd_pr__nfet_01v8 ad=0.825 pd=5.33 as=0.825 ps=5.33 w=5 l=1
X207 diffpairibias.t9 diffpairibias.t8 gnd.t58 gnd.t57 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=2.73 ps=14.78 w=7 l=1
X208 gnd.t297 commonsourceibias.t101 CSoutput.t154 gnd.t231 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X209 CSoutput.t46 a_n6972_8799.t85 vdd.t115 vdd.t114 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X210 vdd.t113 a_n6972_8799.t86 CSoutput.t45 vdd.t46 sky130_fd_pr__pfet_01v8 ad=3.12 pd=16.78 as=1.32 ps=8.33 w=8 l=0.5
X211 commonsourceibias.t15 commonsourceibias.t14 gnd.t196 gnd.t195 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X212 a_n3827_n3924.t12 minus.t16 a_n2848_n452.t31 gnd.t26 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.9
X213 a_n1986_8322.t6 a_n2848_n452.t61 a_n6972_8799.t17 vdd.t38 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X214 CSoutput.t44 a_n6972_8799.t87 vdd.t112 vdd.t76 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X215 outputibias.t1 outputibias.t0 gnd.t352 gnd.t351 sky130_fd_pr__nfet_01v8 ad=2.34 pd=12.78 as=2.34 ps=12.78 w=6 l=2
X216 diffpairibias.t7 diffpairibias.t6 gnd.t368 gnd.t367 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=2.73 ps=14.78 w=7 l=1
X217 vdd.t111 a_n6972_8799.t88 CSoutput.t43 vdd.t110 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X218 CSoutput.t42 a_n6972_8799.t89 vdd.t109 vdd.t60 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X219 vdd.t108 a_n6972_8799.t90 CSoutput.t41 vdd.t107 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X220 vdd.t249 a_n2848_n452.t62 a_n1986_8322.t15 vdd.t248 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=3.51 ps=18.78 w=9 l=0.5
X221 vdd.t101 a_n6972_8799.t91 CSoutput.t40 vdd.t79 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X222 output.t1 outputibias.t10 gnd.t50 gnd.t49 sky130_fd_pr__nfet_01v8 ad=2.34 pd=12.78 as=2.34 ps=12.78 w=6 l=2
X223 a_n3827_n3924.t10 minus.t17 a_n2848_n452.t29 gnd.t31 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.9
X224 CSoutput.t153 commonsourceibias.t102 gnd.t296 gnd.t205 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X225 CSoutput.t202 a_n1986_8322.t20 sky130_fd_pr__cap_mim_m3_1 l=12 w=12
X226 a_n3827_n3924.t42 plus.t20 a_n6972_8799.t27 gnd.t36 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=1.155 ps=7.33 w=7 l=0.9
X227 commonsourceibias.t23 commonsourceibias.t22 gnd.t295 gnd.t259 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X228 a_n3827_n3924.t25 minus.t18 a_n2848_n452.t40 gnd.t9 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.9
X229 gnd.t127 gnd.t124 gnd.t126 gnd.t125 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=0 ps=0 w=7 l=1
X230 a_n1808_13878.t15 a_n2848_n452.t63 vdd.t251 vdd.t250 sky130_fd_pr__pfet_01v8 ad=3.51 pd=18.78 as=1.485 ps=9.33 w=9 l=0.5
X231 vdd.t27 CSoutput.t203 output.t11 gnd.t35 sky130_fd_pr__nfet_01v8 ad=0.825 pd=5.33 as=0.825 ps=5.33 w=5 l=1
X232 CSoutput.t152 commonsourceibias.t103 gnd.t294 gnd.t205 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X233 vdd.t106 a_n6972_8799.t92 CSoutput.t39 vdd.t91 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X234 gnd.t293 commonsourceibias.t104 CSoutput.t151 gnd.t274 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X235 CSoutput.t204 a_n1986_8322.t21 sky130_fd_pr__cap_mim_m3_1 l=12 w=12
X236 CSoutput.t38 a_n6972_8799.t93 vdd.t105 vdd.t102 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X237 CSoutput.t37 a_n6972_8799.t94 vdd.t104 vdd.t89 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X238 gnd.t292 commonsourceibias.t20 commonsourceibias.t21 gnd.t218 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=1.155 ps=7.33 w=7 l=1
X239 gnd.t291 commonsourceibias.t105 CSoutput.t150 gnd.t239 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X240 CSoutput.t149 commonsourceibias.t106 gnd.t290 gnd.t215 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X241 gnd.t123 gnd.t120 gnd.t122 gnd.t121 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=0 ps=0 w=7 l=1
X242 CSoutput.t148 commonsourceibias.t107 gnd.t289 gnd.t272 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X243 gnd.t288 commonsourceibias.t108 CSoutput.t147 gnd.t213 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X244 CSoutput.t146 commonsourceibias.t109 gnd.t287 gnd.t195 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X245 vdd.t207 vdd.t205 vdd.t206 vdd.t192 sky130_fd_pr__pfet_01v8 ad=3.12 pd=16.78 as=0 ps=0 w=8 l=0.5
X246 a_n3827_n3924.t20 diffpairibias.t26 gnd.t61 gnd.t60 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=2.73 ps=14.78 w=7 l=1
X247 gnd.t286 commonsourceibias.t110 CSoutput.t145 gnd.t211 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X248 minus.t2 gnd.t117 gnd.t119 gnd.t118 sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.5
X249 a_n1986_8322.t5 a_n2848_n452.t64 a_n6972_8799.t3 vdd.t1 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X250 commonsourceibias.t19 commonsourceibias.t18 gnd.t285 gnd.t201 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X251 vdd.t3 a_n2848_n452.t65 a_n1986_8322.t14 vdd.t2 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X252 CSoutput.t36 a_n6972_8799.t95 vdd.t103 vdd.t102 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X253 a_n6972_8799.t2 plus.t21 a_n3827_n3924.t41 gnd.t11 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.9
X254 vdd.t100 a_n6972_8799.t96 CSoutput.t35 vdd.t44 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X255 vdd.t204 vdd.t202 vdd.t203 vdd.t185 sky130_fd_pr__pfet_01v8 ad=3.12 pd=16.78 as=0 ps=0 w=8 l=0.5
X256 a_n2848_n452.t2 minus.t19 a_n3827_n3924.t5 gnd.t13 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.9
X257 CSoutput.t144 commonsourceibias.t111 gnd.t284 gnd.t233 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X258 CSoutput.t34 a_n6972_8799.t97 vdd.t99 vdd.t64 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X259 gnd.t283 commonsourceibias.t112 CSoutput.t143 gnd.t191 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X260 a_n3827_n3924.t8 minus.t20 a_n2848_n452.t27 gnd.t27 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=1.155 ps=7.33 w=7 l=0.9
X261 vdd.t98 a_n6972_8799.t98 CSoutput.t33 vdd.t84 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X262 vdd.t97 a_n6972_8799.t99 CSoutput.t32 vdd.t58 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X263 CSoutput.t142 commonsourceibias.t113 gnd.t282 gnd.t233 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X264 gnd.t281 commonsourceibias.t114 CSoutput.t141 gnd.t261 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X265 gnd.t280 commonsourceibias.t115 CSoutput.t140 gnd.t218 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=1.155 ps=7.33 w=7 l=1
X266 CSoutput.t139 commonsourceibias.t116 gnd.t279 gnd.t199 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X267 commonsourceibias.t63 commonsourceibias.t62 gnd.t278 gnd.t277 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X268 vdd.t201 vdd.t198 vdd.t200 vdd.t199 sky130_fd_pr__pfet_01v8 ad=3.51 pd=18.78 as=0 ps=0 w=9 l=0.5
X269 a_n3827_n3924.t17 minus.t21 a_n2848_n452.t35 gnd.t54 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.9
X270 a_n3827_n3924.t16 minus.t22 a_n2848_n452.t34 gnd.t38 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.9
X271 a_n1808_13878.t4 a_n2848_n452.t23 a_n2848_n452.t24 vdd.t18 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X272 CSoutput.t31 a_n6972_8799.t100 vdd.t96 vdd.t76 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X273 CSoutput.t138 commonsourceibias.t117 gnd.t276 gnd.t255 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X274 gnd.t116 gnd.t113 gnd.t115 gnd.t114 sky130_fd_pr__nfet_01v8 ad=1.95 pd=10.78 as=0 ps=0 w=5 l=1
X275 a_n1986_8322.t4 a_n2848_n452.t66 a_n6972_8799.t21 vdd.t13 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X276 diffpairibias.t5 diffpairibias.t4 gnd.t354 gnd.t353 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=2.73 ps=14.78 w=7 l=1
X277 gnd.t275 commonsourceibias.t118 CSoutput.t137 gnd.t274 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X278 CSoutput.t136 commonsourceibias.t119 gnd.t273 gnd.t272 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X279 gnd.t271 commonsourceibias.t60 commonsourceibias.t61 gnd.t226 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=1.155 ps=7.33 w=7 l=1
X280 gnd.t112 gnd.t110 gnd.t111 gnd.t96 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=0 ps=0 w=7 l=1
X281 output.t10 CSoutput.t205 vdd.t16 gnd.t22 sky130_fd_pr__nfet_01v8 ad=0.825 pd=5.33 as=0.825 ps=5.33 w=5 l=1
X282 commonsourceibias.t59 commonsourceibias.t58 gnd.t270 gnd.t229 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X283 CSoutput.t30 a_n6972_8799.t101 vdd.t95 vdd.t94 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X284 gnd.t269 commonsourceibias.t120 CSoutput.t135 gnd.t261 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X285 a_n3827_n3924.t7 diffpairibias.t27 gnd.t19 gnd.t18 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=2.73 ps=14.78 w=7 l=1
X286 vdd.t93 a_n6972_8799.t102 CSoutput.t29 vdd.t84 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X287 gnd.t268 commonsourceibias.t121 CSoutput.t134 gnd.t267 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X288 vdd.t92 a_n6972_8799.t103 CSoutput.t28 vdd.t91 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X289 gnd.t109 gnd.t106 gnd.t108 gnd.t107 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=0 ps=0 w=7 l=0.9
X290 a_n1986_8322.t13 a_n2848_n452.t67 vdd.t42 vdd.t41 sky130_fd_pr__pfet_01v8 ad=3.51 pd=18.78 as=1.485 ps=9.33 w=9 l=0.5
X291 gnd.t266 commonsourceibias.t122 CSoutput.t133 gnd.t224 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X292 CSoutput.t132 commonsourceibias.t123 gnd.t265 gnd.t197 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X293 CSoutput.t27 a_n6972_8799.t104 vdd.t90 vdd.t89 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X294 output.t9 CSoutput.t206 vdd.t17 gnd.t23 sky130_fd_pr__nfet_01v8 ad=1.95 pd=10.78 as=0.825 ps=5.33 w=5 l=1
X295 gnd.t264 commonsourceibias.t56 commonsourceibias.t57 gnd.t193 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X296 a_n3827_n3924.t24 minus.t23 a_n2848_n452.t39 gnd.t24 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.9
X297 commonsourceibias.t55 commonsourceibias.t54 gnd.t263 gnd.t241 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X298 vdd.t261 a_n2848_n452.t68 a_n1808_13878.t14 vdd.t260 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=3.51 ps=18.78 w=9 l=0.5
X299 CSoutput.t26 a_n6972_8799.t105 vdd.t88 vdd.t87 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X300 vdd.t197 vdd.t195 vdd.t196 vdd.t185 sky130_fd_pr__pfet_01v8 ad=3.12 pd=16.78 as=0 ps=0 w=8 l=0.5
X301 gnd.t262 commonsourceibias.t124 CSoutput.t131 gnd.t261 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X302 CSoutput.t130 commonsourceibias.t125 gnd.t258 gnd.t197 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X303 CSoutput.t25 a_n6972_8799.t106 vdd.t86 vdd.t64 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X304 CSoutput.t129 commonsourceibias.t126 gnd.t260 gnd.t259 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X305 gnd.t257 commonsourceibias.t127 CSoutput.t128 gnd.t207 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X306 commonsourceibias.t13 commonsourceibias.t12 gnd.t256 gnd.t255 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X307 gnd.t105 gnd.t102 gnd.t104 gnd.t103 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=0 ps=0 w=7 l=0.9
X308 gnd.t254 commonsourceibias.t128 CSoutput.t127 gnd.t236 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X309 gnd.t101 gnd.t99 plus.t2 gnd.t100 sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.5
X310 vdd.t85 a_n6972_8799.t107 CSoutput.t24 vdd.t84 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X311 vdd.t83 a_n6972_8799.t108 CSoutput.t23 vdd.t58 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X312 vdd.t194 vdd.t191 vdd.t193 vdd.t192 sky130_fd_pr__pfet_01v8 ad=3.12 pd=16.78 as=0 ps=0 w=8 l=0.5
X313 gnd.t253 commonsourceibias.t10 commonsourceibias.t11 gnd.t224 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X314 gnd.t98 gnd.t95 gnd.t97 gnd.t96 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=0 ps=0 w=7 l=1
X315 a_n1986_8322.t3 a_n2848_n452.t69 a_n6972_8799.t34 vdd.t31 sky130_fd_pr__pfet_01v8 ad=3.51 pd=18.78 as=1.485 ps=9.33 w=9 l=0.5
X316 vdd.t190 vdd.t188 vdd.t189 vdd.t177 sky130_fd_pr__pfet_01v8 ad=3.12 pd=16.78 as=0 ps=0 w=8 l=0.5
X317 CSoutput.t22 a_n6972_8799.t109 vdd.t82 vdd.t81 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X318 a_n6972_8799.t4 a_n2848_n452.t70 a_n1986_8322.t2 vdd.t18 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X319 gnd.t252 commonsourceibias.t129 CSoutput.t126 gnd.t193 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X320 vdd.t80 a_n6972_8799.t110 CSoutput.t21 vdd.t79 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X321 a_n1808_13878.t13 a_n2848_n452.t71 vdd.t20 vdd.t19 sky130_fd_pr__pfet_01v8 ad=3.51 pd=18.78 as=1.485 ps=9.33 w=9 l=0.5
X322 CSoutput.t125 commonsourceibias.t130 gnd.t251 gnd.t205 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X323 vdd.t78 a_n6972_8799.t111 CSoutput.t20 vdd.t62 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X324 gnd.t250 commonsourceibias.t131 CSoutput.t124 gnd.t226 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=1.155 ps=7.33 w=7 l=1
X325 CSoutput.t19 a_n6972_8799.t112 vdd.t77 vdd.t76 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X326 vdd.t254 CSoutput.t207 output.t8 gnd.t363 sky130_fd_pr__nfet_01v8 ad=0.825 pd=5.33 as=1.95 ps=10.78 w=5 l=1
X327 vdd.t255 CSoutput.t208 output.t7 gnd.t364 sky130_fd_pr__nfet_01v8 ad=0.825 pd=5.33 as=0.825 ps=5.33 w=5 l=1
X328 gnd.t249 commonsourceibias.t8 commonsourceibias.t9 gnd.t231 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X329 CSoutput.t123 commonsourceibias.t132 gnd.t248 gnd.t243 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=2.73 ps=14.78 w=7 l=1
X330 CSoutput.t122 commonsourceibias.t133 gnd.t247 gnd.t229 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X331 a_n3827_n3924.t40 plus.t22 a_n6972_8799.t19 gnd.t51 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.9
X332 a_n2848_n452.t36 minus.t24 a_n3827_n3924.t18 gnd.t55 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.9
X333 CSoutput.t121 commonsourceibias.t134 gnd.t246 gnd.t199 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X334 a_n6972_8799.t32 plus.t23 a_n3827_n3924.t39 gnd.t369 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.9
X335 gnd.t245 commonsourceibias.t135 CSoutput.t120 gnd.t220 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X336 gnd.t94 gnd.t92 minus.t1 gnd.t93 sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.39 ps=2.78 w=1 l=0.5
X337 vdd.t187 vdd.t184 vdd.t186 vdd.t185 sky130_fd_pr__pfet_01v8 ad=3.12 pd=16.78 as=0 ps=0 w=8 l=0.5
X338 CSoutput.t119 commonsourceibias.t136 gnd.t244 gnd.t243 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=2.73 ps=14.78 w=7 l=1
X339 CSoutput.t209 a_n1986_8322.t21 sky130_fd_pr__cap_mim_m3_1 l=12 w=12
X340 vdd.t183 vdd.t180 vdd.t182 vdd.t181 sky130_fd_pr__pfet_01v8 ad=3.12 pd=16.78 as=0 ps=0 w=8 l=0.5
X341 a_n2848_n452.t41 minus.t25 a_n3827_n3924.t26 gnd.t10 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.9
X342 CSoutput.t118 commonsourceibias.t137 gnd.t242 gnd.t241 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X343 CSoutput.t117 commonsourceibias.t138 gnd.t235 gnd.t222 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X344 gnd.t238 commonsourceibias.t139 CSoutput.t116 gnd.t191 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X345 a_n1808_13878.t3 a_n2848_n452.t3 a_n2848_n452.t4 vdd.t21 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X346 CSoutput.t18 a_n6972_8799.t113 vdd.t71 vdd.t60 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X347 vdd.t73 a_n6972_8799.t114 CSoutput.t17 vdd.t56 sky130_fd_pr__pfet_01v8 ad=3.12 pd=16.78 as=1.32 ps=8.33 w=8 l=0.5
X348 gnd.t240 commonsourceibias.t6 commonsourceibias.t7 gnd.t239 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X349 gnd.t237 commonsourceibias.t4 commonsourceibias.t5 gnd.t236 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X350 CSoutput.t16 a_n6972_8799.t115 vdd.t75 vdd.t52 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X351 a_n3827_n3924.t2 minus.t26 a_n2848_n452.t0 gnd.t6 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.9
X352 a_n3827_n3924.t3 diffpairibias.t28 gnd.t8 gnd.t7 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=2.73 ps=14.78 w=7 l=1
X353 vdd.t74 a_n6972_8799.t116 CSoutput.t15 vdd.t48 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X354 CSoutput.t115 commonsourceibias.t140 gnd.t234 gnd.t233 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X355 gnd.t232 commonsourceibias.t141 CSoutput.t114 gnd.t231 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X356 a_n2848_n452.t26 a_n2848_n452.t25 a_n1808_13878.t2 vdd.t31 sky130_fd_pr__pfet_01v8 ad=3.51 pd=18.78 as=1.485 ps=9.33 w=9 l=0.5
X357 a_n6972_8799.t29 a_n2848_n452.t72 a_n1986_8322.t1 vdd.t0 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=3.51 ps=18.78 w=9 l=0.5
X358 a_n6972_8799.t13 plus.t24 a_n3827_n3924.t38 gnd.t37 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=2.73 ps=14.78 w=7 l=0.9
X359 vdd.t72 a_n6972_8799.t117 CSoutput.t14 vdd.t56 sky130_fd_pr__pfet_01v8 ad=3.12 pd=16.78 as=1.32 ps=8.33 w=8 l=0.5
X360 CSoutput.t13 a_n6972_8799.t118 vdd.t70 vdd.t69 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=3.12 ps=16.78 w=8 l=0.5
X361 CSoutput.t113 commonsourceibias.t142 gnd.t230 gnd.t229 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X362 vdd.t68 a_n6972_8799.t119 CSoutput.t12 vdd.t44 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X363 gnd.t91 gnd.t88 gnd.t90 gnd.t89 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=0 ps=0 w=7 l=1
X364 gnd.t228 commonsourceibias.t143 CSoutput.t112 gnd.t220 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X365 gnd.t227 commonsourceibias.t144 CSoutput.t111 gnd.t226 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=1.155 ps=7.33 w=7 l=1
X366 gnd.t225 commonsourceibias.t145 CSoutput.t110 gnd.t224 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X367 diffpairibias.t3 diffpairibias.t2 gnd.t69 gnd.t68 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=2.73 ps=14.78 w=7 l=1
X368 vdd.t67 a_n6972_8799.t120 CSoutput.t11 vdd.t66 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X369 vdd.t179 vdd.t176 vdd.t178 vdd.t177 sky130_fd_pr__pfet_01v8 ad=3.12 pd=16.78 as=0 ps=0 w=8 l=0.5
X370 CSoutput.t109 commonsourceibias.t146 gnd.t223 gnd.t222 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X371 CSoutput.t10 a_n6972_8799.t121 vdd.t65 vdd.t64 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X372 output.t6 CSoutput.t210 vdd.t26 gnd.t32 sky130_fd_pr__nfet_01v8 ad=0.825 pd=5.33 as=0.825 ps=5.33 w=5 l=1
X373 gnd.t87 gnd.t84 gnd.t86 gnd.t85 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=0 ps=0 w=7 l=1
X374 vdd.t43 CSoutput.t211 output.t5 gnd.t70 sky130_fd_pr__nfet_01v8 ad=0.825 pd=5.33 as=0.825 ps=5.33 w=5 l=1
X375 a_n2848_n452.t1 minus.t27 a_n3827_n3924.t4 gnd.t12 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.9
X376 gnd.t221 commonsourceibias.t147 CSoutput.t108 gnd.t220 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X377 gnd.t83 gnd.t81 plus.t1 gnd.t82 sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.39 ps=2.78 w=1 l=0.5
X378 gnd.t219 commonsourceibias.t148 CSoutput.t107 gnd.t218 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=1.155 ps=7.33 w=7 l=1
X379 vdd.t63 a_n6972_8799.t122 CSoutput.t9 vdd.t62 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X380 gnd.t80 gnd.t77 gnd.t79 gnd.t78 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=0 ps=0 w=7 l=1
X381 diffpairibias.t1 diffpairibias.t0 gnd.t375 gnd.t374 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=2.73 ps=14.78 w=7 l=1
X382 CSoutput.t106 commonsourceibias.t149 gnd.t216 gnd.t215 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X383 CSoutput.t212 a_n1986_8322.t20 sky130_fd_pr__cap_mim_m3_1 l=12 w=12
X384 gnd.t217 commonsourceibias.t150 CSoutput.t105 gnd.t211 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X385 vdd.t257 a_n2848_n452.t73 a_n1808_13878.t12 vdd.t256 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=3.51 ps=18.78 w=9 l=0.5
X386 CSoutput.t8 a_n6972_8799.t123 vdd.t61 vdd.t60 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X387 plus.t0 gnd.t74 gnd.t76 gnd.t75 sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.5
X388 vdd.t59 a_n6972_8799.t124 CSoutput.t7 vdd.t58 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X389 gnd.t214 commonsourceibias.t151 CSoutput.t104 gnd.t213 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X390 vdd.t57 a_n6972_8799.t125 CSoutput.t6 vdd.t56 sky130_fd_pr__pfet_01v8 ad=3.12 pd=16.78 as=1.32 ps=8.33 w=8 l=0.5
X391 CSoutput.t5 a_n6972_8799.t126 vdd.t55 vdd.t54 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X392 a_n6972_8799.t16 plus.t25 a_n3827_n3924.t37 gnd.t42 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.9
X393 gnd.t73 gnd.t71 minus.t0 gnd.t72 sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.5
X394 gnd.t212 commonsourceibias.t152 CSoutput.t103 gnd.t211 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X395 a_n2848_n452.t45 minus.t28 a_n3827_n3924.t31 gnd.t25 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=2.73 ps=14.78 w=7 l=0.9
X396 CSoutput.t4 a_n6972_8799.t127 vdd.t53 vdd.t52 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X397 a_n6972_8799.t28 plus.t26 a_n3827_n3924.t36 gnd.t56 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.9
X398 a_n1986_8322.t0 a_n2848_n452.t74 a_n6972_8799.t33 vdd.t23 sky130_fd_pr__pfet_01v8 ad=3.51 pd=18.78 as=1.485 ps=9.33 w=9 l=0.5
X399 CSoutput.t102 commonsourceibias.t153 gnd.t210 gnd.t209 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=2.73 ps=14.78 w=7 l=1
X400 vdd.t49 a_n6972_8799.t128 CSoutput.t3 vdd.t48 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X401 output.t0 outputibias.t11 gnd.t362 gnd.t361 sky130_fd_pr__nfet_01v8 ad=2.34 pd=12.78 as=2.34 ps=12.78 w=6 l=2
X402 CSoutput.t2 a_n6972_8799.t129 vdd.t51 vdd.t50 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=3.12 ps=16.78 w=8 l=0.5
X403 vdd.t47 a_n6972_8799.t130 CSoutput.t1 vdd.t46 sky130_fd_pr__pfet_01v8 ad=3.12 pd=16.78 as=1.32 ps=8.33 w=8 l=0.5
X404 gnd.t208 commonsourceibias.t154 CSoutput.t101 gnd.t207 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X405 commonsourceibias.t17 commonsourceibias.t16 gnd.t206 gnd.t205 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X406 gnd.t204 commonsourceibias.t155 CSoutput.t100 gnd.t203 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X407 CSoutput.t99 commonsourceibias.t156 gnd.t202 gnd.t201 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X408 a_n1986_8322.t12 a_n2848_n452.t75 vdd.t259 vdd.t258 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X409 a_n1808_13878.t1 a_n2848_n452.t19 a_n2848_n452.t20 vdd.t12 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=3.51 ps=18.78 w=9 l=0.5
X410 vdd.t24 CSoutput.t213 output.t4 gnd.t30 sky130_fd_pr__nfet_01v8 ad=0.825 pd=5.33 as=0.825 ps=5.33 w=5 l=1
X411 vdd.t45 a_n6972_8799.t131 CSoutput.t0 vdd.t44 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X412 a_n3827_n3924.t35 plus.t27 a_n6972_8799.t9 gnd.t26 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.9
X413 a_n3827_n3924.t28 diffpairibias.t29 gnd.t358 gnd.t357 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=2.73 ps=14.78 w=7 l=1
X414 CSoutput.t98 commonsourceibias.t157 gnd.t200 gnd.t199 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X415 CSoutput.t97 commonsourceibias.t158 gnd.t198 gnd.t197 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X416 a_n2848_n452.t14 a_n2848_n452.t13 a_n1808_13878.t0 vdd.t38 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X417 gnd.t192 commonsourceibias.t159 CSoutput.t96 gnd.t191 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X418 vdd.t175 vdd.t172 vdd.t174 vdd.t173 sky130_fd_pr__pfet_01v8 ad=3.51 pd=18.78 as=0 ps=0 w=9 l=0.5
X419 a_n3827_n3924.t34 plus.t28 a_n6972_8799.t10 gnd.t29 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.9
R0 commonsourceibias.n35 commonsourceibias.t52 223.028
R1 commonsourceibias.n128 commonsourceibias.t132 223.028
R2 commonsourceibias.n307 commonsourceibias.t136 223.028
R3 commonsourceibias.n217 commonsourceibias.t64 223.028
R4 commonsourceibias.n454 commonsourceibias.t60 223.028
R5 commonsourceibias.n395 commonsourceibias.t83 223.028
R6 commonsourceibias.n679 commonsourceibias.t144 223.028
R7 commonsourceibias.n589 commonsourceibias.t131 223.028
R8 commonsourceibias.n99 commonsourceibias.t20 207.983
R9 commonsourceibias.n192 commonsourceibias.t78 207.983
R10 commonsourceibias.n371 commonsourceibias.t148 207.983
R11 commonsourceibias.n281 commonsourceibias.t115 207.983
R12 commonsourceibias.n520 commonsourceibias.t44 207.983
R13 commonsourceibias.n566 commonsourceibias.t153 207.983
R14 commonsourceibias.n745 commonsourceibias.t71 207.983
R15 commonsourceibias.n655 commonsourceibias.t100 207.983
R16 commonsourceibias.n97 commonsourceibias.t50 168.701
R17 commonsourceibias.n91 commonsourceibias.t4 168.701
R18 commonsourceibias.n17 commonsourceibias.t40 168.701
R19 commonsourceibias.n83 commonsourceibias.t34 168.701
R20 commonsourceibias.n77 commonsourceibias.t22 168.701
R21 commonsourceibias.n22 commonsourceibias.t24 168.701
R22 commonsourceibias.n69 commonsourceibias.t32 168.701
R23 commonsourceibias.n63 commonsourceibias.t42 168.701
R24 commonsourceibias.n25 commonsourceibias.t0 168.701
R25 commonsourceibias.n27 commonsourceibias.t8 168.701
R26 commonsourceibias.n29 commonsourceibias.t26 168.701
R27 commonsourceibias.n46 commonsourceibias.t36 168.701
R28 commonsourceibias.n40 commonsourceibias.t62 168.701
R29 commonsourceibias.n34 commonsourceibias.t48 168.701
R30 commonsourceibias.n190 commonsourceibias.t146 168.701
R31 commonsourceibias.n184 commonsourceibias.t96 168.701
R32 commonsourceibias.n5 commonsourceibias.t157 168.701
R33 commonsourceibias.n176 commonsourceibias.t112 168.701
R34 commonsourceibias.n170 commonsourceibias.t75 168.701
R35 commonsourceibias.n10 commonsourceibias.t124 168.701
R36 commonsourceibias.n162 commonsourceibias.t113 168.701
R37 commonsourceibias.n156 commonsourceibias.t154 168.701
R38 commonsourceibias.n118 commonsourceibias.t106 168.701
R39 commonsourceibias.n120 commonsourceibias.t92 168.701
R40 commonsourceibias.n122 commonsourceibias.t123 168.701
R41 commonsourceibias.n139 commonsourceibias.t110 168.701
R42 commonsourceibias.n133 commonsourceibias.t82 168.701
R43 commonsourceibias.n127 commonsourceibias.t147 168.701
R44 commonsourceibias.n306 commonsourceibias.t143 168.701
R45 commonsourceibias.n312 commonsourceibias.t70 168.701
R46 commonsourceibias.n318 commonsourceibias.t150 168.701
R47 commonsourceibias.n301 commonsourceibias.t158 168.701
R48 commonsourceibias.n299 commonsourceibias.t101 168.701
R49 commonsourceibias.n297 commonsourceibias.t81 168.701
R50 commonsourceibias.n335 commonsourceibias.t67 168.701
R51 commonsourceibias.n341 commonsourceibias.t111 168.701
R52 commonsourceibias.n294 commonsourceibias.t120 168.701
R53 commonsourceibias.n349 commonsourceibias.t74 168.701
R54 commonsourceibias.n355 commonsourceibias.t159 168.701
R55 commonsourceibias.n289 commonsourceibias.t134 168.701
R56 commonsourceibias.n363 commonsourceibias.t80 168.701
R57 commonsourceibias.n369 commonsourceibias.t68 168.701
R58 commonsourceibias.n279 commonsourceibias.t138 168.701
R59 commonsourceibias.n273 commonsourceibias.t128 168.701
R60 commonsourceibias.n199 commonsourceibias.t116 168.701
R61 commonsourceibias.n265 commonsourceibias.t139 168.701
R62 commonsourceibias.n259 commonsourceibias.t126 168.701
R63 commonsourceibias.n204 commonsourceibias.t114 168.701
R64 commonsourceibias.n251 commonsourceibias.t140 168.701
R65 commonsourceibias.n245 commonsourceibias.t127 168.701
R66 commonsourceibias.n207 commonsourceibias.t149 168.701
R67 commonsourceibias.n209 commonsourceibias.t141 168.701
R68 commonsourceibias.n211 commonsourceibias.t125 168.701
R69 commonsourceibias.n228 commonsourceibias.t152 168.701
R70 commonsourceibias.n222 commonsourceibias.t69 168.701
R71 commonsourceibias.n216 commonsourceibias.t135 168.701
R72 commonsourceibias.n453 commonsourceibias.t58 168.701
R73 commonsourceibias.n459 commonsourceibias.t38 168.701
R74 commonsourceibias.n465 commonsourceibias.t54 168.701
R75 commonsourceibias.n448 commonsourceibias.t6 168.701
R76 commonsourceibias.n446 commonsourceibias.t18 168.701
R77 commonsourceibias.n444 commonsourceibias.t56 168.701
R78 commonsourceibias.n482 commonsourceibias.t30 168.701
R79 commonsourceibias.n488 commonsourceibias.t10 168.701
R80 commonsourceibias.n490 commonsourceibias.t16 168.701
R81 commonsourceibias.n497 commonsourceibias.t46 168.701
R82 commonsourceibias.n503 commonsourceibias.t12 168.701
R83 commonsourceibias.n505 commonsourceibias.t28 168.701
R84 commonsourceibias.n512 commonsourceibias.t14 168.701
R85 commonsourceibias.n518 commonsourceibias.t2 168.701
R86 commonsourceibias.n564 commonsourceibias.t104 168.701
R87 commonsourceibias.n558 commonsourceibias.t73 168.701
R88 commonsourceibias.n551 commonsourceibias.t121 168.701
R89 commonsourceibias.n549 commonsourceibias.t90 168.701
R90 commonsourceibias.n543 commonsourceibias.t151 168.701
R91 commonsourceibias.n536 commonsourceibias.t102 168.701
R92 commonsourceibias.n534 commonsourceibias.t91 168.701
R93 commonsourceibias.n394 commonsourceibias.t84 168.701
R94 commonsourceibias.n400 commonsourceibias.t65 168.701
R95 commonsourceibias.n406 commonsourceibias.t88 168.701
R96 commonsourceibias.n389 commonsourceibias.t95 168.701
R97 commonsourceibias.n387 commonsourceibias.t79 168.701
R98 commonsourceibias.n385 commonsourceibias.t87 168.701
R99 commonsourceibias.n423 commonsourceibias.t119 168.701
R100 commonsourceibias.n678 commonsourceibias.t133 168.701
R101 commonsourceibias.n684 commonsourceibias.t89 168.701
R102 commonsourceibias.n690 commonsourceibias.t72 168.701
R103 commonsourceibias.n673 commonsourceibias.t76 168.701
R104 commonsourceibias.n671 commonsourceibias.t94 168.701
R105 commonsourceibias.n669 commonsourceibias.t98 168.701
R106 commonsourceibias.n707 commonsourceibias.t85 168.701
R107 commonsourceibias.n713 commonsourceibias.t145 168.701
R108 commonsourceibias.n715 commonsourceibias.t103 168.701
R109 commonsourceibias.n722 commonsourceibias.t93 168.701
R110 commonsourceibias.n728 commonsourceibias.t77 168.701
R111 commonsourceibias.n730 commonsourceibias.t66 168.701
R112 commonsourceibias.n737 commonsourceibias.t97 168.701
R113 commonsourceibias.n743 commonsourceibias.t86 168.701
R114 commonsourceibias.n588 commonsourceibias.t142 168.701
R115 commonsourceibias.n594 commonsourceibias.t155 168.701
R116 commonsourceibias.n600 commonsourceibias.t137 168.701
R117 commonsourceibias.n583 commonsourceibias.t105 168.701
R118 commonsourceibias.n581 commonsourceibias.t156 168.701
R119 commonsourceibias.n579 commonsourceibias.t129 168.701
R120 commonsourceibias.n617 commonsourceibias.t107 168.701
R121 commonsourceibias.n623 commonsourceibias.t122 168.701
R122 commonsourceibias.n625 commonsourceibias.t130 168.701
R123 commonsourceibias.n632 commonsourceibias.t108 168.701
R124 commonsourceibias.n638 commonsourceibias.t117 168.701
R125 commonsourceibias.n640 commonsourceibias.t99 168.701
R126 commonsourceibias.n647 commonsourceibias.t109 168.701
R127 commonsourceibias.n653 commonsourceibias.t118 168.701
R128 commonsourceibias.n36 commonsourceibias.n33 161.3
R129 commonsourceibias.n38 commonsourceibias.n37 161.3
R130 commonsourceibias.n39 commonsourceibias.n32 161.3
R131 commonsourceibias.n42 commonsourceibias.n41 161.3
R132 commonsourceibias.n43 commonsourceibias.n31 161.3
R133 commonsourceibias.n45 commonsourceibias.n44 161.3
R134 commonsourceibias.n47 commonsourceibias.n30 161.3
R135 commonsourceibias.n49 commonsourceibias.n48 161.3
R136 commonsourceibias.n51 commonsourceibias.n50 161.3
R137 commonsourceibias.n52 commonsourceibias.n28 161.3
R138 commonsourceibias.n54 commonsourceibias.n53 161.3
R139 commonsourceibias.n56 commonsourceibias.n55 161.3
R140 commonsourceibias.n57 commonsourceibias.n26 161.3
R141 commonsourceibias.n59 commonsourceibias.n58 161.3
R142 commonsourceibias.n61 commonsourceibias.n60 161.3
R143 commonsourceibias.n62 commonsourceibias.n24 161.3
R144 commonsourceibias.n65 commonsourceibias.n64 161.3
R145 commonsourceibias.n66 commonsourceibias.n23 161.3
R146 commonsourceibias.n68 commonsourceibias.n67 161.3
R147 commonsourceibias.n70 commonsourceibias.n21 161.3
R148 commonsourceibias.n72 commonsourceibias.n71 161.3
R149 commonsourceibias.n73 commonsourceibias.n20 161.3
R150 commonsourceibias.n75 commonsourceibias.n74 161.3
R151 commonsourceibias.n76 commonsourceibias.n19 161.3
R152 commonsourceibias.n79 commonsourceibias.n78 161.3
R153 commonsourceibias.n80 commonsourceibias.n18 161.3
R154 commonsourceibias.n82 commonsourceibias.n81 161.3
R155 commonsourceibias.n84 commonsourceibias.n16 161.3
R156 commonsourceibias.n86 commonsourceibias.n85 161.3
R157 commonsourceibias.n87 commonsourceibias.n15 161.3
R158 commonsourceibias.n89 commonsourceibias.n88 161.3
R159 commonsourceibias.n90 commonsourceibias.n14 161.3
R160 commonsourceibias.n93 commonsourceibias.n92 161.3
R161 commonsourceibias.n94 commonsourceibias.n13 161.3
R162 commonsourceibias.n96 commonsourceibias.n95 161.3
R163 commonsourceibias.n98 commonsourceibias.n12 161.3
R164 commonsourceibias.n129 commonsourceibias.n126 161.3
R165 commonsourceibias.n131 commonsourceibias.n130 161.3
R166 commonsourceibias.n132 commonsourceibias.n125 161.3
R167 commonsourceibias.n135 commonsourceibias.n134 161.3
R168 commonsourceibias.n136 commonsourceibias.n124 161.3
R169 commonsourceibias.n138 commonsourceibias.n137 161.3
R170 commonsourceibias.n140 commonsourceibias.n123 161.3
R171 commonsourceibias.n142 commonsourceibias.n141 161.3
R172 commonsourceibias.n144 commonsourceibias.n143 161.3
R173 commonsourceibias.n145 commonsourceibias.n121 161.3
R174 commonsourceibias.n147 commonsourceibias.n146 161.3
R175 commonsourceibias.n149 commonsourceibias.n148 161.3
R176 commonsourceibias.n150 commonsourceibias.n119 161.3
R177 commonsourceibias.n152 commonsourceibias.n151 161.3
R178 commonsourceibias.n154 commonsourceibias.n153 161.3
R179 commonsourceibias.n155 commonsourceibias.n117 161.3
R180 commonsourceibias.n158 commonsourceibias.n157 161.3
R181 commonsourceibias.n159 commonsourceibias.n11 161.3
R182 commonsourceibias.n161 commonsourceibias.n160 161.3
R183 commonsourceibias.n163 commonsourceibias.n9 161.3
R184 commonsourceibias.n165 commonsourceibias.n164 161.3
R185 commonsourceibias.n166 commonsourceibias.n8 161.3
R186 commonsourceibias.n168 commonsourceibias.n167 161.3
R187 commonsourceibias.n169 commonsourceibias.n7 161.3
R188 commonsourceibias.n172 commonsourceibias.n171 161.3
R189 commonsourceibias.n173 commonsourceibias.n6 161.3
R190 commonsourceibias.n175 commonsourceibias.n174 161.3
R191 commonsourceibias.n177 commonsourceibias.n4 161.3
R192 commonsourceibias.n179 commonsourceibias.n178 161.3
R193 commonsourceibias.n180 commonsourceibias.n3 161.3
R194 commonsourceibias.n182 commonsourceibias.n181 161.3
R195 commonsourceibias.n183 commonsourceibias.n2 161.3
R196 commonsourceibias.n186 commonsourceibias.n185 161.3
R197 commonsourceibias.n187 commonsourceibias.n1 161.3
R198 commonsourceibias.n189 commonsourceibias.n188 161.3
R199 commonsourceibias.n191 commonsourceibias.n0 161.3
R200 commonsourceibias.n370 commonsourceibias.n284 161.3
R201 commonsourceibias.n368 commonsourceibias.n367 161.3
R202 commonsourceibias.n366 commonsourceibias.n285 161.3
R203 commonsourceibias.n365 commonsourceibias.n364 161.3
R204 commonsourceibias.n362 commonsourceibias.n286 161.3
R205 commonsourceibias.n361 commonsourceibias.n360 161.3
R206 commonsourceibias.n359 commonsourceibias.n287 161.3
R207 commonsourceibias.n358 commonsourceibias.n357 161.3
R208 commonsourceibias.n356 commonsourceibias.n288 161.3
R209 commonsourceibias.n354 commonsourceibias.n353 161.3
R210 commonsourceibias.n352 commonsourceibias.n290 161.3
R211 commonsourceibias.n351 commonsourceibias.n350 161.3
R212 commonsourceibias.n348 commonsourceibias.n291 161.3
R213 commonsourceibias.n347 commonsourceibias.n346 161.3
R214 commonsourceibias.n345 commonsourceibias.n292 161.3
R215 commonsourceibias.n344 commonsourceibias.n343 161.3
R216 commonsourceibias.n342 commonsourceibias.n293 161.3
R217 commonsourceibias.n340 commonsourceibias.n339 161.3
R218 commonsourceibias.n338 commonsourceibias.n295 161.3
R219 commonsourceibias.n337 commonsourceibias.n336 161.3
R220 commonsourceibias.n334 commonsourceibias.n296 161.3
R221 commonsourceibias.n333 commonsourceibias.n332 161.3
R222 commonsourceibias.n331 commonsourceibias.n330 161.3
R223 commonsourceibias.n329 commonsourceibias.n298 161.3
R224 commonsourceibias.n328 commonsourceibias.n327 161.3
R225 commonsourceibias.n326 commonsourceibias.n325 161.3
R226 commonsourceibias.n324 commonsourceibias.n300 161.3
R227 commonsourceibias.n323 commonsourceibias.n322 161.3
R228 commonsourceibias.n321 commonsourceibias.n320 161.3
R229 commonsourceibias.n319 commonsourceibias.n302 161.3
R230 commonsourceibias.n317 commonsourceibias.n316 161.3
R231 commonsourceibias.n315 commonsourceibias.n303 161.3
R232 commonsourceibias.n314 commonsourceibias.n313 161.3
R233 commonsourceibias.n311 commonsourceibias.n304 161.3
R234 commonsourceibias.n310 commonsourceibias.n309 161.3
R235 commonsourceibias.n308 commonsourceibias.n305 161.3
R236 commonsourceibias.n218 commonsourceibias.n215 161.3
R237 commonsourceibias.n220 commonsourceibias.n219 161.3
R238 commonsourceibias.n221 commonsourceibias.n214 161.3
R239 commonsourceibias.n224 commonsourceibias.n223 161.3
R240 commonsourceibias.n225 commonsourceibias.n213 161.3
R241 commonsourceibias.n227 commonsourceibias.n226 161.3
R242 commonsourceibias.n229 commonsourceibias.n212 161.3
R243 commonsourceibias.n231 commonsourceibias.n230 161.3
R244 commonsourceibias.n233 commonsourceibias.n232 161.3
R245 commonsourceibias.n234 commonsourceibias.n210 161.3
R246 commonsourceibias.n236 commonsourceibias.n235 161.3
R247 commonsourceibias.n238 commonsourceibias.n237 161.3
R248 commonsourceibias.n239 commonsourceibias.n208 161.3
R249 commonsourceibias.n241 commonsourceibias.n240 161.3
R250 commonsourceibias.n243 commonsourceibias.n242 161.3
R251 commonsourceibias.n244 commonsourceibias.n206 161.3
R252 commonsourceibias.n247 commonsourceibias.n246 161.3
R253 commonsourceibias.n248 commonsourceibias.n205 161.3
R254 commonsourceibias.n250 commonsourceibias.n249 161.3
R255 commonsourceibias.n252 commonsourceibias.n203 161.3
R256 commonsourceibias.n254 commonsourceibias.n253 161.3
R257 commonsourceibias.n255 commonsourceibias.n202 161.3
R258 commonsourceibias.n257 commonsourceibias.n256 161.3
R259 commonsourceibias.n258 commonsourceibias.n201 161.3
R260 commonsourceibias.n261 commonsourceibias.n260 161.3
R261 commonsourceibias.n262 commonsourceibias.n200 161.3
R262 commonsourceibias.n264 commonsourceibias.n263 161.3
R263 commonsourceibias.n266 commonsourceibias.n198 161.3
R264 commonsourceibias.n268 commonsourceibias.n267 161.3
R265 commonsourceibias.n269 commonsourceibias.n197 161.3
R266 commonsourceibias.n271 commonsourceibias.n270 161.3
R267 commonsourceibias.n272 commonsourceibias.n196 161.3
R268 commonsourceibias.n275 commonsourceibias.n274 161.3
R269 commonsourceibias.n276 commonsourceibias.n195 161.3
R270 commonsourceibias.n278 commonsourceibias.n277 161.3
R271 commonsourceibias.n280 commonsourceibias.n194 161.3
R272 commonsourceibias.n519 commonsourceibias.n433 161.3
R273 commonsourceibias.n517 commonsourceibias.n516 161.3
R274 commonsourceibias.n515 commonsourceibias.n434 161.3
R275 commonsourceibias.n514 commonsourceibias.n513 161.3
R276 commonsourceibias.n511 commonsourceibias.n435 161.3
R277 commonsourceibias.n510 commonsourceibias.n509 161.3
R278 commonsourceibias.n508 commonsourceibias.n436 161.3
R279 commonsourceibias.n507 commonsourceibias.n506 161.3
R280 commonsourceibias.n504 commonsourceibias.n437 161.3
R281 commonsourceibias.n502 commonsourceibias.n501 161.3
R282 commonsourceibias.n500 commonsourceibias.n438 161.3
R283 commonsourceibias.n499 commonsourceibias.n498 161.3
R284 commonsourceibias.n496 commonsourceibias.n439 161.3
R285 commonsourceibias.n495 commonsourceibias.n494 161.3
R286 commonsourceibias.n493 commonsourceibias.n440 161.3
R287 commonsourceibias.n492 commonsourceibias.n491 161.3
R288 commonsourceibias.n489 commonsourceibias.n441 161.3
R289 commonsourceibias.n487 commonsourceibias.n486 161.3
R290 commonsourceibias.n485 commonsourceibias.n442 161.3
R291 commonsourceibias.n484 commonsourceibias.n483 161.3
R292 commonsourceibias.n481 commonsourceibias.n443 161.3
R293 commonsourceibias.n480 commonsourceibias.n479 161.3
R294 commonsourceibias.n478 commonsourceibias.n477 161.3
R295 commonsourceibias.n476 commonsourceibias.n445 161.3
R296 commonsourceibias.n475 commonsourceibias.n474 161.3
R297 commonsourceibias.n473 commonsourceibias.n472 161.3
R298 commonsourceibias.n471 commonsourceibias.n447 161.3
R299 commonsourceibias.n470 commonsourceibias.n469 161.3
R300 commonsourceibias.n468 commonsourceibias.n467 161.3
R301 commonsourceibias.n466 commonsourceibias.n449 161.3
R302 commonsourceibias.n464 commonsourceibias.n463 161.3
R303 commonsourceibias.n462 commonsourceibias.n450 161.3
R304 commonsourceibias.n461 commonsourceibias.n460 161.3
R305 commonsourceibias.n458 commonsourceibias.n451 161.3
R306 commonsourceibias.n457 commonsourceibias.n456 161.3
R307 commonsourceibias.n455 commonsourceibias.n452 161.3
R308 commonsourceibias.n425 commonsourceibias.n424 161.3
R309 commonsourceibias.n422 commonsourceibias.n384 161.3
R310 commonsourceibias.n421 commonsourceibias.n420 161.3
R311 commonsourceibias.n419 commonsourceibias.n418 161.3
R312 commonsourceibias.n417 commonsourceibias.n386 161.3
R313 commonsourceibias.n416 commonsourceibias.n415 161.3
R314 commonsourceibias.n414 commonsourceibias.n413 161.3
R315 commonsourceibias.n412 commonsourceibias.n388 161.3
R316 commonsourceibias.n411 commonsourceibias.n410 161.3
R317 commonsourceibias.n409 commonsourceibias.n408 161.3
R318 commonsourceibias.n407 commonsourceibias.n390 161.3
R319 commonsourceibias.n405 commonsourceibias.n404 161.3
R320 commonsourceibias.n403 commonsourceibias.n391 161.3
R321 commonsourceibias.n402 commonsourceibias.n401 161.3
R322 commonsourceibias.n399 commonsourceibias.n392 161.3
R323 commonsourceibias.n398 commonsourceibias.n397 161.3
R324 commonsourceibias.n396 commonsourceibias.n393 161.3
R325 commonsourceibias.n531 commonsourceibias.n383 161.3
R326 commonsourceibias.n565 commonsourceibias.n374 161.3
R327 commonsourceibias.n563 commonsourceibias.n562 161.3
R328 commonsourceibias.n561 commonsourceibias.n375 161.3
R329 commonsourceibias.n560 commonsourceibias.n559 161.3
R330 commonsourceibias.n557 commonsourceibias.n376 161.3
R331 commonsourceibias.n556 commonsourceibias.n555 161.3
R332 commonsourceibias.n554 commonsourceibias.n377 161.3
R333 commonsourceibias.n553 commonsourceibias.n552 161.3
R334 commonsourceibias.n550 commonsourceibias.n378 161.3
R335 commonsourceibias.n548 commonsourceibias.n547 161.3
R336 commonsourceibias.n546 commonsourceibias.n379 161.3
R337 commonsourceibias.n545 commonsourceibias.n544 161.3
R338 commonsourceibias.n542 commonsourceibias.n380 161.3
R339 commonsourceibias.n541 commonsourceibias.n540 161.3
R340 commonsourceibias.n539 commonsourceibias.n381 161.3
R341 commonsourceibias.n538 commonsourceibias.n537 161.3
R342 commonsourceibias.n535 commonsourceibias.n382 161.3
R343 commonsourceibias.n533 commonsourceibias.n532 161.3
R344 commonsourceibias.n744 commonsourceibias.n658 161.3
R345 commonsourceibias.n742 commonsourceibias.n741 161.3
R346 commonsourceibias.n740 commonsourceibias.n659 161.3
R347 commonsourceibias.n739 commonsourceibias.n738 161.3
R348 commonsourceibias.n736 commonsourceibias.n660 161.3
R349 commonsourceibias.n735 commonsourceibias.n734 161.3
R350 commonsourceibias.n733 commonsourceibias.n661 161.3
R351 commonsourceibias.n732 commonsourceibias.n731 161.3
R352 commonsourceibias.n729 commonsourceibias.n662 161.3
R353 commonsourceibias.n727 commonsourceibias.n726 161.3
R354 commonsourceibias.n725 commonsourceibias.n663 161.3
R355 commonsourceibias.n724 commonsourceibias.n723 161.3
R356 commonsourceibias.n721 commonsourceibias.n664 161.3
R357 commonsourceibias.n720 commonsourceibias.n719 161.3
R358 commonsourceibias.n718 commonsourceibias.n665 161.3
R359 commonsourceibias.n717 commonsourceibias.n716 161.3
R360 commonsourceibias.n714 commonsourceibias.n666 161.3
R361 commonsourceibias.n712 commonsourceibias.n711 161.3
R362 commonsourceibias.n710 commonsourceibias.n667 161.3
R363 commonsourceibias.n709 commonsourceibias.n708 161.3
R364 commonsourceibias.n706 commonsourceibias.n668 161.3
R365 commonsourceibias.n705 commonsourceibias.n704 161.3
R366 commonsourceibias.n703 commonsourceibias.n702 161.3
R367 commonsourceibias.n701 commonsourceibias.n670 161.3
R368 commonsourceibias.n700 commonsourceibias.n699 161.3
R369 commonsourceibias.n698 commonsourceibias.n697 161.3
R370 commonsourceibias.n696 commonsourceibias.n672 161.3
R371 commonsourceibias.n695 commonsourceibias.n694 161.3
R372 commonsourceibias.n693 commonsourceibias.n692 161.3
R373 commonsourceibias.n691 commonsourceibias.n674 161.3
R374 commonsourceibias.n689 commonsourceibias.n688 161.3
R375 commonsourceibias.n687 commonsourceibias.n675 161.3
R376 commonsourceibias.n686 commonsourceibias.n685 161.3
R377 commonsourceibias.n683 commonsourceibias.n676 161.3
R378 commonsourceibias.n682 commonsourceibias.n681 161.3
R379 commonsourceibias.n680 commonsourceibias.n677 161.3
R380 commonsourceibias.n654 commonsourceibias.n568 161.3
R381 commonsourceibias.n652 commonsourceibias.n651 161.3
R382 commonsourceibias.n650 commonsourceibias.n569 161.3
R383 commonsourceibias.n649 commonsourceibias.n648 161.3
R384 commonsourceibias.n646 commonsourceibias.n570 161.3
R385 commonsourceibias.n645 commonsourceibias.n644 161.3
R386 commonsourceibias.n643 commonsourceibias.n571 161.3
R387 commonsourceibias.n642 commonsourceibias.n641 161.3
R388 commonsourceibias.n639 commonsourceibias.n572 161.3
R389 commonsourceibias.n637 commonsourceibias.n636 161.3
R390 commonsourceibias.n635 commonsourceibias.n573 161.3
R391 commonsourceibias.n634 commonsourceibias.n633 161.3
R392 commonsourceibias.n631 commonsourceibias.n574 161.3
R393 commonsourceibias.n630 commonsourceibias.n629 161.3
R394 commonsourceibias.n628 commonsourceibias.n575 161.3
R395 commonsourceibias.n627 commonsourceibias.n626 161.3
R396 commonsourceibias.n624 commonsourceibias.n576 161.3
R397 commonsourceibias.n622 commonsourceibias.n621 161.3
R398 commonsourceibias.n620 commonsourceibias.n577 161.3
R399 commonsourceibias.n619 commonsourceibias.n618 161.3
R400 commonsourceibias.n616 commonsourceibias.n578 161.3
R401 commonsourceibias.n615 commonsourceibias.n614 161.3
R402 commonsourceibias.n613 commonsourceibias.n612 161.3
R403 commonsourceibias.n611 commonsourceibias.n580 161.3
R404 commonsourceibias.n610 commonsourceibias.n609 161.3
R405 commonsourceibias.n608 commonsourceibias.n607 161.3
R406 commonsourceibias.n606 commonsourceibias.n582 161.3
R407 commonsourceibias.n605 commonsourceibias.n604 161.3
R408 commonsourceibias.n603 commonsourceibias.n602 161.3
R409 commonsourceibias.n601 commonsourceibias.n584 161.3
R410 commonsourceibias.n599 commonsourceibias.n598 161.3
R411 commonsourceibias.n597 commonsourceibias.n585 161.3
R412 commonsourceibias.n596 commonsourceibias.n595 161.3
R413 commonsourceibias.n593 commonsourceibias.n586 161.3
R414 commonsourceibias.n592 commonsourceibias.n591 161.3
R415 commonsourceibias.n590 commonsourceibias.n587 161.3
R416 commonsourceibias.n111 commonsourceibias.n109 81.5057
R417 commonsourceibias.n428 commonsourceibias.n426 81.5057
R418 commonsourceibias.n111 commonsourceibias.n110 80.9324
R419 commonsourceibias.n113 commonsourceibias.n112 80.9324
R420 commonsourceibias.n115 commonsourceibias.n114 80.9324
R421 commonsourceibias.n108 commonsourceibias.n107 80.9324
R422 commonsourceibias.n106 commonsourceibias.n105 80.9324
R423 commonsourceibias.n104 commonsourceibias.n103 80.9324
R424 commonsourceibias.n102 commonsourceibias.n101 80.9324
R425 commonsourceibias.n523 commonsourceibias.n522 80.9324
R426 commonsourceibias.n525 commonsourceibias.n524 80.9324
R427 commonsourceibias.n527 commonsourceibias.n526 80.9324
R428 commonsourceibias.n529 commonsourceibias.n528 80.9324
R429 commonsourceibias.n432 commonsourceibias.n431 80.9324
R430 commonsourceibias.n430 commonsourceibias.n429 80.9324
R431 commonsourceibias.n428 commonsourceibias.n427 80.9324
R432 commonsourceibias.n100 commonsourceibias.n99 80.6037
R433 commonsourceibias.n193 commonsourceibias.n192 80.6037
R434 commonsourceibias.n372 commonsourceibias.n371 80.6037
R435 commonsourceibias.n282 commonsourceibias.n281 80.6037
R436 commonsourceibias.n521 commonsourceibias.n520 80.6037
R437 commonsourceibias.n567 commonsourceibias.n566 80.6037
R438 commonsourceibias.n746 commonsourceibias.n745 80.6037
R439 commonsourceibias.n656 commonsourceibias.n655 80.6037
R440 commonsourceibias.n85 commonsourceibias.n84 56.5617
R441 commonsourceibias.n71 commonsourceibias.n70 56.5617
R442 commonsourceibias.n62 commonsourceibias.n61 56.5617
R443 commonsourceibias.n48 commonsourceibias.n47 56.5617
R444 commonsourceibias.n178 commonsourceibias.n177 56.5617
R445 commonsourceibias.n164 commonsourceibias.n163 56.5617
R446 commonsourceibias.n155 commonsourceibias.n154 56.5617
R447 commonsourceibias.n141 commonsourceibias.n140 56.5617
R448 commonsourceibias.n320 commonsourceibias.n319 56.5617
R449 commonsourceibias.n334 commonsourceibias.n333 56.5617
R450 commonsourceibias.n343 commonsourceibias.n342 56.5617
R451 commonsourceibias.n357 commonsourceibias.n356 56.5617
R452 commonsourceibias.n267 commonsourceibias.n266 56.5617
R453 commonsourceibias.n253 commonsourceibias.n252 56.5617
R454 commonsourceibias.n244 commonsourceibias.n243 56.5617
R455 commonsourceibias.n230 commonsourceibias.n229 56.5617
R456 commonsourceibias.n467 commonsourceibias.n466 56.5617
R457 commonsourceibias.n481 commonsourceibias.n480 56.5617
R458 commonsourceibias.n491 commonsourceibias.n489 56.5617
R459 commonsourceibias.n506 commonsourceibias.n504 56.5617
R460 commonsourceibias.n552 commonsourceibias.n550 56.5617
R461 commonsourceibias.n537 commonsourceibias.n535 56.5617
R462 commonsourceibias.n408 commonsourceibias.n407 56.5617
R463 commonsourceibias.n422 commonsourceibias.n421 56.5617
R464 commonsourceibias.n692 commonsourceibias.n691 56.5617
R465 commonsourceibias.n706 commonsourceibias.n705 56.5617
R466 commonsourceibias.n716 commonsourceibias.n714 56.5617
R467 commonsourceibias.n731 commonsourceibias.n729 56.5617
R468 commonsourceibias.n602 commonsourceibias.n601 56.5617
R469 commonsourceibias.n616 commonsourceibias.n615 56.5617
R470 commonsourceibias.n626 commonsourceibias.n624 56.5617
R471 commonsourceibias.n641 commonsourceibias.n639 56.5617
R472 commonsourceibias.n76 commonsourceibias.n75 56.0773
R473 commonsourceibias.n57 commonsourceibias.n56 56.0773
R474 commonsourceibias.n169 commonsourceibias.n168 56.0773
R475 commonsourceibias.n150 commonsourceibias.n149 56.0773
R476 commonsourceibias.n329 commonsourceibias.n328 56.0773
R477 commonsourceibias.n348 commonsourceibias.n347 56.0773
R478 commonsourceibias.n258 commonsourceibias.n257 56.0773
R479 commonsourceibias.n239 commonsourceibias.n238 56.0773
R480 commonsourceibias.n476 commonsourceibias.n475 56.0773
R481 commonsourceibias.n496 commonsourceibias.n495 56.0773
R482 commonsourceibias.n542 commonsourceibias.n541 56.0773
R483 commonsourceibias.n417 commonsourceibias.n416 56.0773
R484 commonsourceibias.n701 commonsourceibias.n700 56.0773
R485 commonsourceibias.n721 commonsourceibias.n720 56.0773
R486 commonsourceibias.n611 commonsourceibias.n610 56.0773
R487 commonsourceibias.n631 commonsourceibias.n630 56.0773
R488 commonsourceibias.n99 commonsourceibias.n98 55.3321
R489 commonsourceibias.n192 commonsourceibias.n191 55.3321
R490 commonsourceibias.n371 commonsourceibias.n370 55.3321
R491 commonsourceibias.n281 commonsourceibias.n280 55.3321
R492 commonsourceibias.n520 commonsourceibias.n519 55.3321
R493 commonsourceibias.n566 commonsourceibias.n565 55.3321
R494 commonsourceibias.n745 commonsourceibias.n744 55.3321
R495 commonsourceibias.n655 commonsourceibias.n654 55.3321
R496 commonsourceibias.n90 commonsourceibias.n89 55.1086
R497 commonsourceibias.n41 commonsourceibias.n31 55.1086
R498 commonsourceibias.n183 commonsourceibias.n182 55.1086
R499 commonsourceibias.n134 commonsourceibias.n124 55.1086
R500 commonsourceibias.n313 commonsourceibias.n303 55.1086
R501 commonsourceibias.n362 commonsourceibias.n361 55.1086
R502 commonsourceibias.n272 commonsourceibias.n271 55.1086
R503 commonsourceibias.n223 commonsourceibias.n213 55.1086
R504 commonsourceibias.n460 commonsourceibias.n450 55.1086
R505 commonsourceibias.n511 commonsourceibias.n510 55.1086
R506 commonsourceibias.n557 commonsourceibias.n556 55.1086
R507 commonsourceibias.n401 commonsourceibias.n391 55.1086
R508 commonsourceibias.n685 commonsourceibias.n675 55.1086
R509 commonsourceibias.n736 commonsourceibias.n735 55.1086
R510 commonsourceibias.n595 commonsourceibias.n585 55.1086
R511 commonsourceibias.n646 commonsourceibias.n645 55.1086
R512 commonsourceibias.n35 commonsourceibias.n34 47.4592
R513 commonsourceibias.n128 commonsourceibias.n127 47.4592
R514 commonsourceibias.n307 commonsourceibias.n306 47.4592
R515 commonsourceibias.n217 commonsourceibias.n216 47.4592
R516 commonsourceibias.n454 commonsourceibias.n453 47.4592
R517 commonsourceibias.n395 commonsourceibias.n394 47.4592
R518 commonsourceibias.n679 commonsourceibias.n678 47.4592
R519 commonsourceibias.n589 commonsourceibias.n588 47.4592
R520 commonsourceibias.n308 commonsourceibias.n307 44.0436
R521 commonsourceibias.n455 commonsourceibias.n454 44.0436
R522 commonsourceibias.n396 commonsourceibias.n395 44.0436
R523 commonsourceibias.n680 commonsourceibias.n679 44.0436
R524 commonsourceibias.n590 commonsourceibias.n589 44.0436
R525 commonsourceibias.n36 commonsourceibias.n35 44.0436
R526 commonsourceibias.n129 commonsourceibias.n128 44.0436
R527 commonsourceibias.n218 commonsourceibias.n217 44.0436
R528 commonsourceibias.n92 commonsourceibias.n13 42.5146
R529 commonsourceibias.n39 commonsourceibias.n38 42.5146
R530 commonsourceibias.n185 commonsourceibias.n1 42.5146
R531 commonsourceibias.n132 commonsourceibias.n131 42.5146
R532 commonsourceibias.n311 commonsourceibias.n310 42.5146
R533 commonsourceibias.n364 commonsourceibias.n285 42.5146
R534 commonsourceibias.n274 commonsourceibias.n195 42.5146
R535 commonsourceibias.n221 commonsourceibias.n220 42.5146
R536 commonsourceibias.n458 commonsourceibias.n457 42.5146
R537 commonsourceibias.n513 commonsourceibias.n434 42.5146
R538 commonsourceibias.n559 commonsourceibias.n375 42.5146
R539 commonsourceibias.n399 commonsourceibias.n398 42.5146
R540 commonsourceibias.n683 commonsourceibias.n682 42.5146
R541 commonsourceibias.n738 commonsourceibias.n659 42.5146
R542 commonsourceibias.n593 commonsourceibias.n592 42.5146
R543 commonsourceibias.n648 commonsourceibias.n569 42.5146
R544 commonsourceibias.n78 commonsourceibias.n18 41.5458
R545 commonsourceibias.n53 commonsourceibias.n52 41.5458
R546 commonsourceibias.n171 commonsourceibias.n6 41.5458
R547 commonsourceibias.n146 commonsourceibias.n145 41.5458
R548 commonsourceibias.n325 commonsourceibias.n324 41.5458
R549 commonsourceibias.n350 commonsourceibias.n290 41.5458
R550 commonsourceibias.n260 commonsourceibias.n200 41.5458
R551 commonsourceibias.n235 commonsourceibias.n234 41.5458
R552 commonsourceibias.n472 commonsourceibias.n471 41.5458
R553 commonsourceibias.n498 commonsourceibias.n438 41.5458
R554 commonsourceibias.n544 commonsourceibias.n379 41.5458
R555 commonsourceibias.n413 commonsourceibias.n412 41.5458
R556 commonsourceibias.n697 commonsourceibias.n696 41.5458
R557 commonsourceibias.n723 commonsourceibias.n663 41.5458
R558 commonsourceibias.n607 commonsourceibias.n606 41.5458
R559 commonsourceibias.n633 commonsourceibias.n573 41.5458
R560 commonsourceibias.n68 commonsourceibias.n23 40.577
R561 commonsourceibias.n64 commonsourceibias.n23 40.577
R562 commonsourceibias.n161 commonsourceibias.n11 40.577
R563 commonsourceibias.n157 commonsourceibias.n11 40.577
R564 commonsourceibias.n336 commonsourceibias.n295 40.577
R565 commonsourceibias.n340 commonsourceibias.n295 40.577
R566 commonsourceibias.n250 commonsourceibias.n205 40.577
R567 commonsourceibias.n246 commonsourceibias.n205 40.577
R568 commonsourceibias.n483 commonsourceibias.n442 40.577
R569 commonsourceibias.n487 commonsourceibias.n442 40.577
R570 commonsourceibias.n533 commonsourceibias.n383 40.577
R571 commonsourceibias.n424 commonsourceibias.n383 40.577
R572 commonsourceibias.n708 commonsourceibias.n667 40.577
R573 commonsourceibias.n712 commonsourceibias.n667 40.577
R574 commonsourceibias.n618 commonsourceibias.n577 40.577
R575 commonsourceibias.n622 commonsourceibias.n577 40.577
R576 commonsourceibias.n82 commonsourceibias.n18 39.6083
R577 commonsourceibias.n52 commonsourceibias.n51 39.6083
R578 commonsourceibias.n175 commonsourceibias.n6 39.6083
R579 commonsourceibias.n145 commonsourceibias.n144 39.6083
R580 commonsourceibias.n324 commonsourceibias.n323 39.6083
R581 commonsourceibias.n354 commonsourceibias.n290 39.6083
R582 commonsourceibias.n264 commonsourceibias.n200 39.6083
R583 commonsourceibias.n234 commonsourceibias.n233 39.6083
R584 commonsourceibias.n471 commonsourceibias.n470 39.6083
R585 commonsourceibias.n502 commonsourceibias.n438 39.6083
R586 commonsourceibias.n548 commonsourceibias.n379 39.6083
R587 commonsourceibias.n412 commonsourceibias.n411 39.6083
R588 commonsourceibias.n696 commonsourceibias.n695 39.6083
R589 commonsourceibias.n727 commonsourceibias.n663 39.6083
R590 commonsourceibias.n606 commonsourceibias.n605 39.6083
R591 commonsourceibias.n637 commonsourceibias.n573 39.6083
R592 commonsourceibias.n96 commonsourceibias.n13 38.6395
R593 commonsourceibias.n38 commonsourceibias.n33 38.6395
R594 commonsourceibias.n189 commonsourceibias.n1 38.6395
R595 commonsourceibias.n131 commonsourceibias.n126 38.6395
R596 commonsourceibias.n310 commonsourceibias.n305 38.6395
R597 commonsourceibias.n368 commonsourceibias.n285 38.6395
R598 commonsourceibias.n278 commonsourceibias.n195 38.6395
R599 commonsourceibias.n220 commonsourceibias.n215 38.6395
R600 commonsourceibias.n457 commonsourceibias.n452 38.6395
R601 commonsourceibias.n517 commonsourceibias.n434 38.6395
R602 commonsourceibias.n563 commonsourceibias.n375 38.6395
R603 commonsourceibias.n398 commonsourceibias.n393 38.6395
R604 commonsourceibias.n682 commonsourceibias.n677 38.6395
R605 commonsourceibias.n742 commonsourceibias.n659 38.6395
R606 commonsourceibias.n592 commonsourceibias.n587 38.6395
R607 commonsourceibias.n652 commonsourceibias.n569 38.6395
R608 commonsourceibias.n89 commonsourceibias.n15 26.0455
R609 commonsourceibias.n45 commonsourceibias.n31 26.0455
R610 commonsourceibias.n182 commonsourceibias.n3 26.0455
R611 commonsourceibias.n138 commonsourceibias.n124 26.0455
R612 commonsourceibias.n317 commonsourceibias.n303 26.0455
R613 commonsourceibias.n361 commonsourceibias.n287 26.0455
R614 commonsourceibias.n271 commonsourceibias.n197 26.0455
R615 commonsourceibias.n227 commonsourceibias.n213 26.0455
R616 commonsourceibias.n464 commonsourceibias.n450 26.0455
R617 commonsourceibias.n510 commonsourceibias.n436 26.0455
R618 commonsourceibias.n556 commonsourceibias.n377 26.0455
R619 commonsourceibias.n405 commonsourceibias.n391 26.0455
R620 commonsourceibias.n689 commonsourceibias.n675 26.0455
R621 commonsourceibias.n735 commonsourceibias.n661 26.0455
R622 commonsourceibias.n599 commonsourceibias.n585 26.0455
R623 commonsourceibias.n645 commonsourceibias.n571 26.0455
R624 commonsourceibias.n75 commonsourceibias.n20 25.0767
R625 commonsourceibias.n58 commonsourceibias.n57 25.0767
R626 commonsourceibias.n168 commonsourceibias.n8 25.0767
R627 commonsourceibias.n151 commonsourceibias.n150 25.0767
R628 commonsourceibias.n330 commonsourceibias.n329 25.0767
R629 commonsourceibias.n347 commonsourceibias.n292 25.0767
R630 commonsourceibias.n257 commonsourceibias.n202 25.0767
R631 commonsourceibias.n240 commonsourceibias.n239 25.0767
R632 commonsourceibias.n477 commonsourceibias.n476 25.0767
R633 commonsourceibias.n495 commonsourceibias.n440 25.0767
R634 commonsourceibias.n541 commonsourceibias.n381 25.0767
R635 commonsourceibias.n418 commonsourceibias.n417 25.0767
R636 commonsourceibias.n702 commonsourceibias.n701 25.0767
R637 commonsourceibias.n720 commonsourceibias.n665 25.0767
R638 commonsourceibias.n612 commonsourceibias.n611 25.0767
R639 commonsourceibias.n630 commonsourceibias.n575 25.0767
R640 commonsourceibias.n71 commonsourceibias.n22 24.3464
R641 commonsourceibias.n61 commonsourceibias.n25 24.3464
R642 commonsourceibias.n164 commonsourceibias.n10 24.3464
R643 commonsourceibias.n154 commonsourceibias.n118 24.3464
R644 commonsourceibias.n333 commonsourceibias.n297 24.3464
R645 commonsourceibias.n343 commonsourceibias.n294 24.3464
R646 commonsourceibias.n253 commonsourceibias.n204 24.3464
R647 commonsourceibias.n243 commonsourceibias.n207 24.3464
R648 commonsourceibias.n480 commonsourceibias.n444 24.3464
R649 commonsourceibias.n491 commonsourceibias.n490 24.3464
R650 commonsourceibias.n537 commonsourceibias.n536 24.3464
R651 commonsourceibias.n421 commonsourceibias.n385 24.3464
R652 commonsourceibias.n705 commonsourceibias.n669 24.3464
R653 commonsourceibias.n716 commonsourceibias.n715 24.3464
R654 commonsourceibias.n615 commonsourceibias.n579 24.3464
R655 commonsourceibias.n626 commonsourceibias.n625 24.3464
R656 commonsourceibias.n85 commonsourceibias.n17 23.8546
R657 commonsourceibias.n47 commonsourceibias.n46 23.8546
R658 commonsourceibias.n178 commonsourceibias.n5 23.8546
R659 commonsourceibias.n140 commonsourceibias.n139 23.8546
R660 commonsourceibias.n319 commonsourceibias.n318 23.8546
R661 commonsourceibias.n357 commonsourceibias.n289 23.8546
R662 commonsourceibias.n267 commonsourceibias.n199 23.8546
R663 commonsourceibias.n229 commonsourceibias.n228 23.8546
R664 commonsourceibias.n466 commonsourceibias.n465 23.8546
R665 commonsourceibias.n506 commonsourceibias.n505 23.8546
R666 commonsourceibias.n552 commonsourceibias.n551 23.8546
R667 commonsourceibias.n407 commonsourceibias.n406 23.8546
R668 commonsourceibias.n691 commonsourceibias.n690 23.8546
R669 commonsourceibias.n731 commonsourceibias.n730 23.8546
R670 commonsourceibias.n601 commonsourceibias.n600 23.8546
R671 commonsourceibias.n641 commonsourceibias.n640 23.8546
R672 commonsourceibias.n98 commonsourceibias.n97 17.4607
R673 commonsourceibias.n191 commonsourceibias.n190 17.4607
R674 commonsourceibias.n370 commonsourceibias.n369 17.4607
R675 commonsourceibias.n280 commonsourceibias.n279 17.4607
R676 commonsourceibias.n519 commonsourceibias.n518 17.4607
R677 commonsourceibias.n565 commonsourceibias.n564 17.4607
R678 commonsourceibias.n744 commonsourceibias.n743 17.4607
R679 commonsourceibias.n654 commonsourceibias.n653 17.4607
R680 commonsourceibias.n84 commonsourceibias.n83 16.9689
R681 commonsourceibias.n48 commonsourceibias.n29 16.9689
R682 commonsourceibias.n177 commonsourceibias.n176 16.9689
R683 commonsourceibias.n141 commonsourceibias.n122 16.9689
R684 commonsourceibias.n320 commonsourceibias.n301 16.9689
R685 commonsourceibias.n356 commonsourceibias.n355 16.9689
R686 commonsourceibias.n266 commonsourceibias.n265 16.9689
R687 commonsourceibias.n230 commonsourceibias.n211 16.9689
R688 commonsourceibias.n467 commonsourceibias.n448 16.9689
R689 commonsourceibias.n504 commonsourceibias.n503 16.9689
R690 commonsourceibias.n550 commonsourceibias.n549 16.9689
R691 commonsourceibias.n408 commonsourceibias.n389 16.9689
R692 commonsourceibias.n692 commonsourceibias.n673 16.9689
R693 commonsourceibias.n729 commonsourceibias.n728 16.9689
R694 commonsourceibias.n602 commonsourceibias.n583 16.9689
R695 commonsourceibias.n639 commonsourceibias.n638 16.9689
R696 commonsourceibias.n70 commonsourceibias.n69 16.477
R697 commonsourceibias.n63 commonsourceibias.n62 16.477
R698 commonsourceibias.n163 commonsourceibias.n162 16.477
R699 commonsourceibias.n156 commonsourceibias.n155 16.477
R700 commonsourceibias.n335 commonsourceibias.n334 16.477
R701 commonsourceibias.n342 commonsourceibias.n341 16.477
R702 commonsourceibias.n252 commonsourceibias.n251 16.477
R703 commonsourceibias.n245 commonsourceibias.n244 16.477
R704 commonsourceibias.n482 commonsourceibias.n481 16.477
R705 commonsourceibias.n489 commonsourceibias.n488 16.477
R706 commonsourceibias.n535 commonsourceibias.n534 16.477
R707 commonsourceibias.n423 commonsourceibias.n422 16.477
R708 commonsourceibias.n707 commonsourceibias.n706 16.477
R709 commonsourceibias.n714 commonsourceibias.n713 16.477
R710 commonsourceibias.n617 commonsourceibias.n616 16.477
R711 commonsourceibias.n624 commonsourceibias.n623 16.477
R712 commonsourceibias.n77 commonsourceibias.n76 15.9852
R713 commonsourceibias.n56 commonsourceibias.n27 15.9852
R714 commonsourceibias.n170 commonsourceibias.n169 15.9852
R715 commonsourceibias.n149 commonsourceibias.n120 15.9852
R716 commonsourceibias.n328 commonsourceibias.n299 15.9852
R717 commonsourceibias.n349 commonsourceibias.n348 15.9852
R718 commonsourceibias.n259 commonsourceibias.n258 15.9852
R719 commonsourceibias.n238 commonsourceibias.n209 15.9852
R720 commonsourceibias.n475 commonsourceibias.n446 15.9852
R721 commonsourceibias.n497 commonsourceibias.n496 15.9852
R722 commonsourceibias.n543 commonsourceibias.n542 15.9852
R723 commonsourceibias.n416 commonsourceibias.n387 15.9852
R724 commonsourceibias.n700 commonsourceibias.n671 15.9852
R725 commonsourceibias.n722 commonsourceibias.n721 15.9852
R726 commonsourceibias.n610 commonsourceibias.n581 15.9852
R727 commonsourceibias.n632 commonsourceibias.n631 15.9852
R728 commonsourceibias.n91 commonsourceibias.n90 15.4934
R729 commonsourceibias.n41 commonsourceibias.n40 15.4934
R730 commonsourceibias.n184 commonsourceibias.n183 15.4934
R731 commonsourceibias.n134 commonsourceibias.n133 15.4934
R732 commonsourceibias.n313 commonsourceibias.n312 15.4934
R733 commonsourceibias.n363 commonsourceibias.n362 15.4934
R734 commonsourceibias.n273 commonsourceibias.n272 15.4934
R735 commonsourceibias.n223 commonsourceibias.n222 15.4934
R736 commonsourceibias.n460 commonsourceibias.n459 15.4934
R737 commonsourceibias.n512 commonsourceibias.n511 15.4934
R738 commonsourceibias.n558 commonsourceibias.n557 15.4934
R739 commonsourceibias.n401 commonsourceibias.n400 15.4934
R740 commonsourceibias.n685 commonsourceibias.n684 15.4934
R741 commonsourceibias.n737 commonsourceibias.n736 15.4934
R742 commonsourceibias.n595 commonsourceibias.n594 15.4934
R743 commonsourceibias.n647 commonsourceibias.n646 15.4934
R744 commonsourceibias.n102 commonsourceibias.n100 13.2663
R745 commonsourceibias.n523 commonsourceibias.n521 13.2663
R746 commonsourceibias.n748 commonsourceibias.n373 10.4122
R747 commonsourceibias.n159 commonsourceibias.n116 9.50363
R748 commonsourceibias.n531 commonsourceibias.n530 9.50363
R749 commonsourceibias.n92 commonsourceibias.n91 9.09948
R750 commonsourceibias.n40 commonsourceibias.n39 9.09948
R751 commonsourceibias.n185 commonsourceibias.n184 9.09948
R752 commonsourceibias.n133 commonsourceibias.n132 9.09948
R753 commonsourceibias.n312 commonsourceibias.n311 9.09948
R754 commonsourceibias.n364 commonsourceibias.n363 9.09948
R755 commonsourceibias.n274 commonsourceibias.n273 9.09948
R756 commonsourceibias.n222 commonsourceibias.n221 9.09948
R757 commonsourceibias.n459 commonsourceibias.n458 9.09948
R758 commonsourceibias.n513 commonsourceibias.n512 9.09948
R759 commonsourceibias.n559 commonsourceibias.n558 9.09948
R760 commonsourceibias.n400 commonsourceibias.n399 9.09948
R761 commonsourceibias.n684 commonsourceibias.n683 9.09948
R762 commonsourceibias.n738 commonsourceibias.n737 9.09948
R763 commonsourceibias.n594 commonsourceibias.n593 9.09948
R764 commonsourceibias.n648 commonsourceibias.n647 9.09948
R765 commonsourceibias.n283 commonsourceibias.n193 8.79451
R766 commonsourceibias.n657 commonsourceibias.n567 8.79451
R767 commonsourceibias.n78 commonsourceibias.n77 8.60764
R768 commonsourceibias.n53 commonsourceibias.n27 8.60764
R769 commonsourceibias.n171 commonsourceibias.n170 8.60764
R770 commonsourceibias.n146 commonsourceibias.n120 8.60764
R771 commonsourceibias.n325 commonsourceibias.n299 8.60764
R772 commonsourceibias.n350 commonsourceibias.n349 8.60764
R773 commonsourceibias.n260 commonsourceibias.n259 8.60764
R774 commonsourceibias.n235 commonsourceibias.n209 8.60764
R775 commonsourceibias.n472 commonsourceibias.n446 8.60764
R776 commonsourceibias.n498 commonsourceibias.n497 8.60764
R777 commonsourceibias.n544 commonsourceibias.n543 8.60764
R778 commonsourceibias.n413 commonsourceibias.n387 8.60764
R779 commonsourceibias.n697 commonsourceibias.n671 8.60764
R780 commonsourceibias.n723 commonsourceibias.n722 8.60764
R781 commonsourceibias.n607 commonsourceibias.n581 8.60764
R782 commonsourceibias.n633 commonsourceibias.n632 8.60764
R783 commonsourceibias.n748 commonsourceibias.n747 8.46921
R784 commonsourceibias.n69 commonsourceibias.n68 8.11581
R785 commonsourceibias.n64 commonsourceibias.n63 8.11581
R786 commonsourceibias.n162 commonsourceibias.n161 8.11581
R787 commonsourceibias.n157 commonsourceibias.n156 8.11581
R788 commonsourceibias.n336 commonsourceibias.n335 8.11581
R789 commonsourceibias.n341 commonsourceibias.n340 8.11581
R790 commonsourceibias.n251 commonsourceibias.n250 8.11581
R791 commonsourceibias.n246 commonsourceibias.n245 8.11581
R792 commonsourceibias.n483 commonsourceibias.n482 8.11581
R793 commonsourceibias.n488 commonsourceibias.n487 8.11581
R794 commonsourceibias.n534 commonsourceibias.n533 8.11581
R795 commonsourceibias.n424 commonsourceibias.n423 8.11581
R796 commonsourceibias.n708 commonsourceibias.n707 8.11581
R797 commonsourceibias.n713 commonsourceibias.n712 8.11581
R798 commonsourceibias.n618 commonsourceibias.n617 8.11581
R799 commonsourceibias.n623 commonsourceibias.n622 8.11581
R800 commonsourceibias.n83 commonsourceibias.n82 7.62397
R801 commonsourceibias.n51 commonsourceibias.n29 7.62397
R802 commonsourceibias.n176 commonsourceibias.n175 7.62397
R803 commonsourceibias.n144 commonsourceibias.n122 7.62397
R804 commonsourceibias.n323 commonsourceibias.n301 7.62397
R805 commonsourceibias.n355 commonsourceibias.n354 7.62397
R806 commonsourceibias.n265 commonsourceibias.n264 7.62397
R807 commonsourceibias.n233 commonsourceibias.n211 7.62397
R808 commonsourceibias.n470 commonsourceibias.n448 7.62397
R809 commonsourceibias.n503 commonsourceibias.n502 7.62397
R810 commonsourceibias.n549 commonsourceibias.n548 7.62397
R811 commonsourceibias.n411 commonsourceibias.n389 7.62397
R812 commonsourceibias.n695 commonsourceibias.n673 7.62397
R813 commonsourceibias.n728 commonsourceibias.n727 7.62397
R814 commonsourceibias.n605 commonsourceibias.n583 7.62397
R815 commonsourceibias.n638 commonsourceibias.n637 7.62397
R816 commonsourceibias.n97 commonsourceibias.n96 7.13213
R817 commonsourceibias.n34 commonsourceibias.n33 7.13213
R818 commonsourceibias.n190 commonsourceibias.n189 7.13213
R819 commonsourceibias.n127 commonsourceibias.n126 7.13213
R820 commonsourceibias.n306 commonsourceibias.n305 7.13213
R821 commonsourceibias.n369 commonsourceibias.n368 7.13213
R822 commonsourceibias.n279 commonsourceibias.n278 7.13213
R823 commonsourceibias.n216 commonsourceibias.n215 7.13213
R824 commonsourceibias.n453 commonsourceibias.n452 7.13213
R825 commonsourceibias.n518 commonsourceibias.n517 7.13213
R826 commonsourceibias.n564 commonsourceibias.n563 7.13213
R827 commonsourceibias.n394 commonsourceibias.n393 7.13213
R828 commonsourceibias.n678 commonsourceibias.n677 7.13213
R829 commonsourceibias.n743 commonsourceibias.n742 7.13213
R830 commonsourceibias.n588 commonsourceibias.n587 7.13213
R831 commonsourceibias.n653 commonsourceibias.n652 7.13213
R832 commonsourceibias.n373 commonsourceibias.n372 5.06534
R833 commonsourceibias.n283 commonsourceibias.n282 5.06534
R834 commonsourceibias.n747 commonsourceibias.n746 5.06534
R835 commonsourceibias.n657 commonsourceibias.n656 5.06534
R836 commonsourceibias commonsourceibias.n748 4.04308
R837 commonsourceibias.n373 commonsourceibias.n283 3.72967
R838 commonsourceibias.n747 commonsourceibias.n657 3.72967
R839 commonsourceibias.n109 commonsourceibias.t49 2.82907
R840 commonsourceibias.n109 commonsourceibias.t53 2.82907
R841 commonsourceibias.n110 commonsourceibias.t37 2.82907
R842 commonsourceibias.n110 commonsourceibias.t63 2.82907
R843 commonsourceibias.n112 commonsourceibias.t9 2.82907
R844 commonsourceibias.n112 commonsourceibias.t27 2.82907
R845 commonsourceibias.n114 commonsourceibias.t43 2.82907
R846 commonsourceibias.n114 commonsourceibias.t1 2.82907
R847 commonsourceibias.n107 commonsourceibias.t25 2.82907
R848 commonsourceibias.n107 commonsourceibias.t33 2.82907
R849 commonsourceibias.n105 commonsourceibias.t35 2.82907
R850 commonsourceibias.n105 commonsourceibias.t23 2.82907
R851 commonsourceibias.n103 commonsourceibias.t5 2.82907
R852 commonsourceibias.n103 commonsourceibias.t41 2.82907
R853 commonsourceibias.n101 commonsourceibias.t21 2.82907
R854 commonsourceibias.n101 commonsourceibias.t51 2.82907
R855 commonsourceibias.n522 commonsourceibias.t3 2.82907
R856 commonsourceibias.n522 commonsourceibias.t45 2.82907
R857 commonsourceibias.n524 commonsourceibias.t29 2.82907
R858 commonsourceibias.n524 commonsourceibias.t15 2.82907
R859 commonsourceibias.n526 commonsourceibias.t47 2.82907
R860 commonsourceibias.n526 commonsourceibias.t13 2.82907
R861 commonsourceibias.n528 commonsourceibias.t11 2.82907
R862 commonsourceibias.n528 commonsourceibias.t17 2.82907
R863 commonsourceibias.n431 commonsourceibias.t57 2.82907
R864 commonsourceibias.n431 commonsourceibias.t31 2.82907
R865 commonsourceibias.n429 commonsourceibias.t7 2.82907
R866 commonsourceibias.n429 commonsourceibias.t19 2.82907
R867 commonsourceibias.n427 commonsourceibias.t39 2.82907
R868 commonsourceibias.n427 commonsourceibias.t55 2.82907
R869 commonsourceibias.n426 commonsourceibias.t61 2.82907
R870 commonsourceibias.n426 commonsourceibias.t59 2.82907
R871 commonsourceibias.n17 commonsourceibias.n15 0.738255
R872 commonsourceibias.n46 commonsourceibias.n45 0.738255
R873 commonsourceibias.n5 commonsourceibias.n3 0.738255
R874 commonsourceibias.n139 commonsourceibias.n138 0.738255
R875 commonsourceibias.n318 commonsourceibias.n317 0.738255
R876 commonsourceibias.n289 commonsourceibias.n287 0.738255
R877 commonsourceibias.n199 commonsourceibias.n197 0.738255
R878 commonsourceibias.n228 commonsourceibias.n227 0.738255
R879 commonsourceibias.n465 commonsourceibias.n464 0.738255
R880 commonsourceibias.n505 commonsourceibias.n436 0.738255
R881 commonsourceibias.n551 commonsourceibias.n377 0.738255
R882 commonsourceibias.n406 commonsourceibias.n405 0.738255
R883 commonsourceibias.n690 commonsourceibias.n689 0.738255
R884 commonsourceibias.n730 commonsourceibias.n661 0.738255
R885 commonsourceibias.n600 commonsourceibias.n599 0.738255
R886 commonsourceibias.n640 commonsourceibias.n571 0.738255
R887 commonsourceibias.n104 commonsourceibias.n102 0.573776
R888 commonsourceibias.n106 commonsourceibias.n104 0.573776
R889 commonsourceibias.n108 commonsourceibias.n106 0.573776
R890 commonsourceibias.n115 commonsourceibias.n113 0.573776
R891 commonsourceibias.n113 commonsourceibias.n111 0.573776
R892 commonsourceibias.n430 commonsourceibias.n428 0.573776
R893 commonsourceibias.n432 commonsourceibias.n430 0.573776
R894 commonsourceibias.n529 commonsourceibias.n527 0.573776
R895 commonsourceibias.n527 commonsourceibias.n525 0.573776
R896 commonsourceibias.n525 commonsourceibias.n523 0.573776
R897 commonsourceibias.n116 commonsourceibias.n108 0.287138
R898 commonsourceibias.n116 commonsourceibias.n115 0.287138
R899 commonsourceibias.n530 commonsourceibias.n432 0.287138
R900 commonsourceibias.n530 commonsourceibias.n529 0.287138
R901 commonsourceibias.n100 commonsourceibias.n12 0.285035
R902 commonsourceibias.n193 commonsourceibias.n0 0.285035
R903 commonsourceibias.n372 commonsourceibias.n284 0.285035
R904 commonsourceibias.n282 commonsourceibias.n194 0.285035
R905 commonsourceibias.n521 commonsourceibias.n433 0.285035
R906 commonsourceibias.n567 commonsourceibias.n374 0.285035
R907 commonsourceibias.n746 commonsourceibias.n658 0.285035
R908 commonsourceibias.n656 commonsourceibias.n568 0.285035
R909 commonsourceibias.n22 commonsourceibias.n20 0.246418
R910 commonsourceibias.n58 commonsourceibias.n25 0.246418
R911 commonsourceibias.n10 commonsourceibias.n8 0.246418
R912 commonsourceibias.n151 commonsourceibias.n118 0.246418
R913 commonsourceibias.n330 commonsourceibias.n297 0.246418
R914 commonsourceibias.n294 commonsourceibias.n292 0.246418
R915 commonsourceibias.n204 commonsourceibias.n202 0.246418
R916 commonsourceibias.n240 commonsourceibias.n207 0.246418
R917 commonsourceibias.n477 commonsourceibias.n444 0.246418
R918 commonsourceibias.n490 commonsourceibias.n440 0.246418
R919 commonsourceibias.n536 commonsourceibias.n381 0.246418
R920 commonsourceibias.n418 commonsourceibias.n385 0.246418
R921 commonsourceibias.n702 commonsourceibias.n669 0.246418
R922 commonsourceibias.n715 commonsourceibias.n665 0.246418
R923 commonsourceibias.n612 commonsourceibias.n579 0.246418
R924 commonsourceibias.n625 commonsourceibias.n575 0.246418
R925 commonsourceibias.n95 commonsourceibias.n12 0.189894
R926 commonsourceibias.n95 commonsourceibias.n94 0.189894
R927 commonsourceibias.n94 commonsourceibias.n93 0.189894
R928 commonsourceibias.n93 commonsourceibias.n14 0.189894
R929 commonsourceibias.n88 commonsourceibias.n14 0.189894
R930 commonsourceibias.n88 commonsourceibias.n87 0.189894
R931 commonsourceibias.n87 commonsourceibias.n86 0.189894
R932 commonsourceibias.n86 commonsourceibias.n16 0.189894
R933 commonsourceibias.n81 commonsourceibias.n16 0.189894
R934 commonsourceibias.n81 commonsourceibias.n80 0.189894
R935 commonsourceibias.n80 commonsourceibias.n79 0.189894
R936 commonsourceibias.n79 commonsourceibias.n19 0.189894
R937 commonsourceibias.n74 commonsourceibias.n19 0.189894
R938 commonsourceibias.n74 commonsourceibias.n73 0.189894
R939 commonsourceibias.n73 commonsourceibias.n72 0.189894
R940 commonsourceibias.n72 commonsourceibias.n21 0.189894
R941 commonsourceibias.n67 commonsourceibias.n21 0.189894
R942 commonsourceibias.n67 commonsourceibias.n66 0.189894
R943 commonsourceibias.n66 commonsourceibias.n65 0.189894
R944 commonsourceibias.n65 commonsourceibias.n24 0.189894
R945 commonsourceibias.n60 commonsourceibias.n24 0.189894
R946 commonsourceibias.n60 commonsourceibias.n59 0.189894
R947 commonsourceibias.n59 commonsourceibias.n26 0.189894
R948 commonsourceibias.n55 commonsourceibias.n26 0.189894
R949 commonsourceibias.n55 commonsourceibias.n54 0.189894
R950 commonsourceibias.n54 commonsourceibias.n28 0.189894
R951 commonsourceibias.n50 commonsourceibias.n28 0.189894
R952 commonsourceibias.n50 commonsourceibias.n49 0.189894
R953 commonsourceibias.n49 commonsourceibias.n30 0.189894
R954 commonsourceibias.n44 commonsourceibias.n30 0.189894
R955 commonsourceibias.n44 commonsourceibias.n43 0.189894
R956 commonsourceibias.n43 commonsourceibias.n42 0.189894
R957 commonsourceibias.n42 commonsourceibias.n32 0.189894
R958 commonsourceibias.n37 commonsourceibias.n32 0.189894
R959 commonsourceibias.n37 commonsourceibias.n36 0.189894
R960 commonsourceibias.n158 commonsourceibias.n117 0.189894
R961 commonsourceibias.n153 commonsourceibias.n117 0.189894
R962 commonsourceibias.n153 commonsourceibias.n152 0.189894
R963 commonsourceibias.n152 commonsourceibias.n119 0.189894
R964 commonsourceibias.n148 commonsourceibias.n119 0.189894
R965 commonsourceibias.n148 commonsourceibias.n147 0.189894
R966 commonsourceibias.n147 commonsourceibias.n121 0.189894
R967 commonsourceibias.n143 commonsourceibias.n121 0.189894
R968 commonsourceibias.n143 commonsourceibias.n142 0.189894
R969 commonsourceibias.n142 commonsourceibias.n123 0.189894
R970 commonsourceibias.n137 commonsourceibias.n123 0.189894
R971 commonsourceibias.n137 commonsourceibias.n136 0.189894
R972 commonsourceibias.n136 commonsourceibias.n135 0.189894
R973 commonsourceibias.n135 commonsourceibias.n125 0.189894
R974 commonsourceibias.n130 commonsourceibias.n125 0.189894
R975 commonsourceibias.n130 commonsourceibias.n129 0.189894
R976 commonsourceibias.n188 commonsourceibias.n0 0.189894
R977 commonsourceibias.n188 commonsourceibias.n187 0.189894
R978 commonsourceibias.n187 commonsourceibias.n186 0.189894
R979 commonsourceibias.n186 commonsourceibias.n2 0.189894
R980 commonsourceibias.n181 commonsourceibias.n2 0.189894
R981 commonsourceibias.n181 commonsourceibias.n180 0.189894
R982 commonsourceibias.n180 commonsourceibias.n179 0.189894
R983 commonsourceibias.n179 commonsourceibias.n4 0.189894
R984 commonsourceibias.n174 commonsourceibias.n4 0.189894
R985 commonsourceibias.n174 commonsourceibias.n173 0.189894
R986 commonsourceibias.n173 commonsourceibias.n172 0.189894
R987 commonsourceibias.n172 commonsourceibias.n7 0.189894
R988 commonsourceibias.n167 commonsourceibias.n7 0.189894
R989 commonsourceibias.n167 commonsourceibias.n166 0.189894
R990 commonsourceibias.n166 commonsourceibias.n165 0.189894
R991 commonsourceibias.n165 commonsourceibias.n9 0.189894
R992 commonsourceibias.n160 commonsourceibias.n9 0.189894
R993 commonsourceibias.n367 commonsourceibias.n284 0.189894
R994 commonsourceibias.n367 commonsourceibias.n366 0.189894
R995 commonsourceibias.n366 commonsourceibias.n365 0.189894
R996 commonsourceibias.n365 commonsourceibias.n286 0.189894
R997 commonsourceibias.n360 commonsourceibias.n286 0.189894
R998 commonsourceibias.n360 commonsourceibias.n359 0.189894
R999 commonsourceibias.n359 commonsourceibias.n358 0.189894
R1000 commonsourceibias.n358 commonsourceibias.n288 0.189894
R1001 commonsourceibias.n353 commonsourceibias.n288 0.189894
R1002 commonsourceibias.n353 commonsourceibias.n352 0.189894
R1003 commonsourceibias.n352 commonsourceibias.n351 0.189894
R1004 commonsourceibias.n351 commonsourceibias.n291 0.189894
R1005 commonsourceibias.n346 commonsourceibias.n291 0.189894
R1006 commonsourceibias.n346 commonsourceibias.n345 0.189894
R1007 commonsourceibias.n345 commonsourceibias.n344 0.189894
R1008 commonsourceibias.n344 commonsourceibias.n293 0.189894
R1009 commonsourceibias.n339 commonsourceibias.n293 0.189894
R1010 commonsourceibias.n339 commonsourceibias.n338 0.189894
R1011 commonsourceibias.n338 commonsourceibias.n337 0.189894
R1012 commonsourceibias.n337 commonsourceibias.n296 0.189894
R1013 commonsourceibias.n332 commonsourceibias.n296 0.189894
R1014 commonsourceibias.n332 commonsourceibias.n331 0.189894
R1015 commonsourceibias.n331 commonsourceibias.n298 0.189894
R1016 commonsourceibias.n327 commonsourceibias.n298 0.189894
R1017 commonsourceibias.n327 commonsourceibias.n326 0.189894
R1018 commonsourceibias.n326 commonsourceibias.n300 0.189894
R1019 commonsourceibias.n322 commonsourceibias.n300 0.189894
R1020 commonsourceibias.n322 commonsourceibias.n321 0.189894
R1021 commonsourceibias.n321 commonsourceibias.n302 0.189894
R1022 commonsourceibias.n316 commonsourceibias.n302 0.189894
R1023 commonsourceibias.n316 commonsourceibias.n315 0.189894
R1024 commonsourceibias.n315 commonsourceibias.n314 0.189894
R1025 commonsourceibias.n314 commonsourceibias.n304 0.189894
R1026 commonsourceibias.n309 commonsourceibias.n304 0.189894
R1027 commonsourceibias.n309 commonsourceibias.n308 0.189894
R1028 commonsourceibias.n277 commonsourceibias.n194 0.189894
R1029 commonsourceibias.n277 commonsourceibias.n276 0.189894
R1030 commonsourceibias.n276 commonsourceibias.n275 0.189894
R1031 commonsourceibias.n275 commonsourceibias.n196 0.189894
R1032 commonsourceibias.n270 commonsourceibias.n196 0.189894
R1033 commonsourceibias.n270 commonsourceibias.n269 0.189894
R1034 commonsourceibias.n269 commonsourceibias.n268 0.189894
R1035 commonsourceibias.n268 commonsourceibias.n198 0.189894
R1036 commonsourceibias.n263 commonsourceibias.n198 0.189894
R1037 commonsourceibias.n263 commonsourceibias.n262 0.189894
R1038 commonsourceibias.n262 commonsourceibias.n261 0.189894
R1039 commonsourceibias.n261 commonsourceibias.n201 0.189894
R1040 commonsourceibias.n256 commonsourceibias.n201 0.189894
R1041 commonsourceibias.n256 commonsourceibias.n255 0.189894
R1042 commonsourceibias.n255 commonsourceibias.n254 0.189894
R1043 commonsourceibias.n254 commonsourceibias.n203 0.189894
R1044 commonsourceibias.n249 commonsourceibias.n203 0.189894
R1045 commonsourceibias.n249 commonsourceibias.n248 0.189894
R1046 commonsourceibias.n248 commonsourceibias.n247 0.189894
R1047 commonsourceibias.n247 commonsourceibias.n206 0.189894
R1048 commonsourceibias.n242 commonsourceibias.n206 0.189894
R1049 commonsourceibias.n242 commonsourceibias.n241 0.189894
R1050 commonsourceibias.n241 commonsourceibias.n208 0.189894
R1051 commonsourceibias.n237 commonsourceibias.n208 0.189894
R1052 commonsourceibias.n237 commonsourceibias.n236 0.189894
R1053 commonsourceibias.n236 commonsourceibias.n210 0.189894
R1054 commonsourceibias.n232 commonsourceibias.n210 0.189894
R1055 commonsourceibias.n232 commonsourceibias.n231 0.189894
R1056 commonsourceibias.n231 commonsourceibias.n212 0.189894
R1057 commonsourceibias.n226 commonsourceibias.n212 0.189894
R1058 commonsourceibias.n226 commonsourceibias.n225 0.189894
R1059 commonsourceibias.n225 commonsourceibias.n224 0.189894
R1060 commonsourceibias.n224 commonsourceibias.n214 0.189894
R1061 commonsourceibias.n219 commonsourceibias.n214 0.189894
R1062 commonsourceibias.n219 commonsourceibias.n218 0.189894
R1063 commonsourceibias.n456 commonsourceibias.n455 0.189894
R1064 commonsourceibias.n456 commonsourceibias.n451 0.189894
R1065 commonsourceibias.n461 commonsourceibias.n451 0.189894
R1066 commonsourceibias.n462 commonsourceibias.n461 0.189894
R1067 commonsourceibias.n463 commonsourceibias.n462 0.189894
R1068 commonsourceibias.n463 commonsourceibias.n449 0.189894
R1069 commonsourceibias.n468 commonsourceibias.n449 0.189894
R1070 commonsourceibias.n469 commonsourceibias.n468 0.189894
R1071 commonsourceibias.n469 commonsourceibias.n447 0.189894
R1072 commonsourceibias.n473 commonsourceibias.n447 0.189894
R1073 commonsourceibias.n474 commonsourceibias.n473 0.189894
R1074 commonsourceibias.n474 commonsourceibias.n445 0.189894
R1075 commonsourceibias.n478 commonsourceibias.n445 0.189894
R1076 commonsourceibias.n479 commonsourceibias.n478 0.189894
R1077 commonsourceibias.n479 commonsourceibias.n443 0.189894
R1078 commonsourceibias.n484 commonsourceibias.n443 0.189894
R1079 commonsourceibias.n485 commonsourceibias.n484 0.189894
R1080 commonsourceibias.n486 commonsourceibias.n485 0.189894
R1081 commonsourceibias.n486 commonsourceibias.n441 0.189894
R1082 commonsourceibias.n492 commonsourceibias.n441 0.189894
R1083 commonsourceibias.n493 commonsourceibias.n492 0.189894
R1084 commonsourceibias.n494 commonsourceibias.n493 0.189894
R1085 commonsourceibias.n494 commonsourceibias.n439 0.189894
R1086 commonsourceibias.n499 commonsourceibias.n439 0.189894
R1087 commonsourceibias.n500 commonsourceibias.n499 0.189894
R1088 commonsourceibias.n501 commonsourceibias.n500 0.189894
R1089 commonsourceibias.n501 commonsourceibias.n437 0.189894
R1090 commonsourceibias.n507 commonsourceibias.n437 0.189894
R1091 commonsourceibias.n508 commonsourceibias.n507 0.189894
R1092 commonsourceibias.n509 commonsourceibias.n508 0.189894
R1093 commonsourceibias.n509 commonsourceibias.n435 0.189894
R1094 commonsourceibias.n514 commonsourceibias.n435 0.189894
R1095 commonsourceibias.n515 commonsourceibias.n514 0.189894
R1096 commonsourceibias.n516 commonsourceibias.n515 0.189894
R1097 commonsourceibias.n516 commonsourceibias.n433 0.189894
R1098 commonsourceibias.n397 commonsourceibias.n396 0.189894
R1099 commonsourceibias.n397 commonsourceibias.n392 0.189894
R1100 commonsourceibias.n402 commonsourceibias.n392 0.189894
R1101 commonsourceibias.n403 commonsourceibias.n402 0.189894
R1102 commonsourceibias.n404 commonsourceibias.n403 0.189894
R1103 commonsourceibias.n404 commonsourceibias.n390 0.189894
R1104 commonsourceibias.n409 commonsourceibias.n390 0.189894
R1105 commonsourceibias.n410 commonsourceibias.n409 0.189894
R1106 commonsourceibias.n410 commonsourceibias.n388 0.189894
R1107 commonsourceibias.n414 commonsourceibias.n388 0.189894
R1108 commonsourceibias.n415 commonsourceibias.n414 0.189894
R1109 commonsourceibias.n415 commonsourceibias.n386 0.189894
R1110 commonsourceibias.n419 commonsourceibias.n386 0.189894
R1111 commonsourceibias.n420 commonsourceibias.n419 0.189894
R1112 commonsourceibias.n420 commonsourceibias.n384 0.189894
R1113 commonsourceibias.n425 commonsourceibias.n384 0.189894
R1114 commonsourceibias.n532 commonsourceibias.n382 0.189894
R1115 commonsourceibias.n538 commonsourceibias.n382 0.189894
R1116 commonsourceibias.n539 commonsourceibias.n538 0.189894
R1117 commonsourceibias.n540 commonsourceibias.n539 0.189894
R1118 commonsourceibias.n540 commonsourceibias.n380 0.189894
R1119 commonsourceibias.n545 commonsourceibias.n380 0.189894
R1120 commonsourceibias.n546 commonsourceibias.n545 0.189894
R1121 commonsourceibias.n547 commonsourceibias.n546 0.189894
R1122 commonsourceibias.n547 commonsourceibias.n378 0.189894
R1123 commonsourceibias.n553 commonsourceibias.n378 0.189894
R1124 commonsourceibias.n554 commonsourceibias.n553 0.189894
R1125 commonsourceibias.n555 commonsourceibias.n554 0.189894
R1126 commonsourceibias.n555 commonsourceibias.n376 0.189894
R1127 commonsourceibias.n560 commonsourceibias.n376 0.189894
R1128 commonsourceibias.n561 commonsourceibias.n560 0.189894
R1129 commonsourceibias.n562 commonsourceibias.n561 0.189894
R1130 commonsourceibias.n562 commonsourceibias.n374 0.189894
R1131 commonsourceibias.n681 commonsourceibias.n680 0.189894
R1132 commonsourceibias.n681 commonsourceibias.n676 0.189894
R1133 commonsourceibias.n686 commonsourceibias.n676 0.189894
R1134 commonsourceibias.n687 commonsourceibias.n686 0.189894
R1135 commonsourceibias.n688 commonsourceibias.n687 0.189894
R1136 commonsourceibias.n688 commonsourceibias.n674 0.189894
R1137 commonsourceibias.n693 commonsourceibias.n674 0.189894
R1138 commonsourceibias.n694 commonsourceibias.n693 0.189894
R1139 commonsourceibias.n694 commonsourceibias.n672 0.189894
R1140 commonsourceibias.n698 commonsourceibias.n672 0.189894
R1141 commonsourceibias.n699 commonsourceibias.n698 0.189894
R1142 commonsourceibias.n699 commonsourceibias.n670 0.189894
R1143 commonsourceibias.n703 commonsourceibias.n670 0.189894
R1144 commonsourceibias.n704 commonsourceibias.n703 0.189894
R1145 commonsourceibias.n704 commonsourceibias.n668 0.189894
R1146 commonsourceibias.n709 commonsourceibias.n668 0.189894
R1147 commonsourceibias.n710 commonsourceibias.n709 0.189894
R1148 commonsourceibias.n711 commonsourceibias.n710 0.189894
R1149 commonsourceibias.n711 commonsourceibias.n666 0.189894
R1150 commonsourceibias.n717 commonsourceibias.n666 0.189894
R1151 commonsourceibias.n718 commonsourceibias.n717 0.189894
R1152 commonsourceibias.n719 commonsourceibias.n718 0.189894
R1153 commonsourceibias.n719 commonsourceibias.n664 0.189894
R1154 commonsourceibias.n724 commonsourceibias.n664 0.189894
R1155 commonsourceibias.n725 commonsourceibias.n724 0.189894
R1156 commonsourceibias.n726 commonsourceibias.n725 0.189894
R1157 commonsourceibias.n726 commonsourceibias.n662 0.189894
R1158 commonsourceibias.n732 commonsourceibias.n662 0.189894
R1159 commonsourceibias.n733 commonsourceibias.n732 0.189894
R1160 commonsourceibias.n734 commonsourceibias.n733 0.189894
R1161 commonsourceibias.n734 commonsourceibias.n660 0.189894
R1162 commonsourceibias.n739 commonsourceibias.n660 0.189894
R1163 commonsourceibias.n740 commonsourceibias.n739 0.189894
R1164 commonsourceibias.n741 commonsourceibias.n740 0.189894
R1165 commonsourceibias.n741 commonsourceibias.n658 0.189894
R1166 commonsourceibias.n591 commonsourceibias.n590 0.189894
R1167 commonsourceibias.n591 commonsourceibias.n586 0.189894
R1168 commonsourceibias.n596 commonsourceibias.n586 0.189894
R1169 commonsourceibias.n597 commonsourceibias.n596 0.189894
R1170 commonsourceibias.n598 commonsourceibias.n597 0.189894
R1171 commonsourceibias.n598 commonsourceibias.n584 0.189894
R1172 commonsourceibias.n603 commonsourceibias.n584 0.189894
R1173 commonsourceibias.n604 commonsourceibias.n603 0.189894
R1174 commonsourceibias.n604 commonsourceibias.n582 0.189894
R1175 commonsourceibias.n608 commonsourceibias.n582 0.189894
R1176 commonsourceibias.n609 commonsourceibias.n608 0.189894
R1177 commonsourceibias.n609 commonsourceibias.n580 0.189894
R1178 commonsourceibias.n613 commonsourceibias.n580 0.189894
R1179 commonsourceibias.n614 commonsourceibias.n613 0.189894
R1180 commonsourceibias.n614 commonsourceibias.n578 0.189894
R1181 commonsourceibias.n619 commonsourceibias.n578 0.189894
R1182 commonsourceibias.n620 commonsourceibias.n619 0.189894
R1183 commonsourceibias.n621 commonsourceibias.n620 0.189894
R1184 commonsourceibias.n621 commonsourceibias.n576 0.189894
R1185 commonsourceibias.n627 commonsourceibias.n576 0.189894
R1186 commonsourceibias.n628 commonsourceibias.n627 0.189894
R1187 commonsourceibias.n629 commonsourceibias.n628 0.189894
R1188 commonsourceibias.n629 commonsourceibias.n574 0.189894
R1189 commonsourceibias.n634 commonsourceibias.n574 0.189894
R1190 commonsourceibias.n635 commonsourceibias.n634 0.189894
R1191 commonsourceibias.n636 commonsourceibias.n635 0.189894
R1192 commonsourceibias.n636 commonsourceibias.n572 0.189894
R1193 commonsourceibias.n642 commonsourceibias.n572 0.189894
R1194 commonsourceibias.n643 commonsourceibias.n642 0.189894
R1195 commonsourceibias.n644 commonsourceibias.n643 0.189894
R1196 commonsourceibias.n644 commonsourceibias.n570 0.189894
R1197 commonsourceibias.n649 commonsourceibias.n570 0.189894
R1198 commonsourceibias.n650 commonsourceibias.n649 0.189894
R1199 commonsourceibias.n651 commonsourceibias.n650 0.189894
R1200 commonsourceibias.n651 commonsourceibias.n568 0.189894
R1201 commonsourceibias.n159 commonsourceibias.n158 0.170955
R1202 commonsourceibias.n160 commonsourceibias.n159 0.170955
R1203 commonsourceibias.n531 commonsourceibias.n425 0.170955
R1204 commonsourceibias.n532 commonsourceibias.n531 0.170955
R1205 gnd.n2853 gnd.n2852 1004.37
R1206 gnd.n5088 gnd.n4774 939.716
R1207 gnd.n7680 gnd.n207 795.207
R1208 gnd.n347 gnd.n210 795.207
R1209 gnd.n7215 gnd.n519 795.207
R1210 gnd.n605 gnd.n523 795.207
R1211 gnd.n5598 gnd.n5597 795.207
R1212 gnd.n5664 gnd.n1682 795.207
R1213 gnd.n4928 gnd.n4811 795.207
R1214 gnd.n4967 gnd.n1982 795.207
R1215 gnd.n4682 gnd.n1993 766.379
R1216 gnd.n4685 gnd.n4684 766.379
R1217 gnd.n3924 gnd.n3827 766.379
R1218 gnd.n3920 gnd.n3825 766.379
R1219 gnd.n4773 gnd.n2015 756.769
R1220 gnd.n4676 gnd.n4675 756.769
R1221 gnd.n4017 gnd.n3734 756.769
R1222 gnd.n4015 gnd.n3737 756.769
R1223 gnd.n7678 gnd.n212 739.952
R1224 gnd.n7569 gnd.n209 739.952
R1225 gnd.n893 gnd.n521 739.952
R1226 gnd.n7213 gnd.n524 739.952
R1227 gnd.n5857 gnd.n1659 739.952
R1228 gnd.n5872 gnd.n1647 739.952
R1229 gnd.n5091 gnd.n5090 739.952
R1230 gnd.n5086 gnd.n1978 739.952
R1231 gnd.n3164 gnd.n2206 723.135
R1232 gnd.n2854 gnd.n2514 723.135
R1233 gnd.n2682 gnd.n409 723.135
R1234 gnd.n2082 gnd.n2081 723.135
R1235 gnd.n5734 gnd.n1705 711.122
R1236 gnd.n7184 gnd.n587 711.122
R1237 gnd.n5738 gnd.n1687 711.122
R1238 gnd.n7186 gnd.n580 711.122
R1239 gnd.n2206 gnd.n2205 585
R1240 gnd.n3166 gnd.n2206 585
R1241 gnd.n3169 gnd.n3168 585
R1242 gnd.n3168 gnd.n3167 585
R1243 gnd.n2203 gnd.n2202 585
R1244 gnd.n2202 gnd.n2201 585
R1245 gnd.n3174 gnd.n3173 585
R1246 gnd.n3175 gnd.n3174 585
R1247 gnd.n2200 gnd.n2199 585
R1248 gnd.n3176 gnd.n2200 585
R1249 gnd.n3179 gnd.n3178 585
R1250 gnd.n3178 gnd.n3177 585
R1251 gnd.n2197 gnd.n2196 585
R1252 gnd.n2196 gnd.n2195 585
R1253 gnd.n3184 gnd.n3183 585
R1254 gnd.n3185 gnd.n3184 585
R1255 gnd.n2194 gnd.n2193 585
R1256 gnd.n3186 gnd.n2194 585
R1257 gnd.n3189 gnd.n3188 585
R1258 gnd.n3188 gnd.n3187 585
R1259 gnd.n2191 gnd.n2190 585
R1260 gnd.n2190 gnd.n2189 585
R1261 gnd.n3194 gnd.n3193 585
R1262 gnd.n3195 gnd.n3194 585
R1263 gnd.n2188 gnd.n2187 585
R1264 gnd.n3196 gnd.n2188 585
R1265 gnd.n3199 gnd.n3198 585
R1266 gnd.n3198 gnd.n3197 585
R1267 gnd.n2185 gnd.n2184 585
R1268 gnd.n2184 gnd.n2183 585
R1269 gnd.n3204 gnd.n3203 585
R1270 gnd.n3205 gnd.n3204 585
R1271 gnd.n2182 gnd.n2181 585
R1272 gnd.n3206 gnd.n2182 585
R1273 gnd.n3209 gnd.n3208 585
R1274 gnd.n3208 gnd.n3207 585
R1275 gnd.n2179 gnd.n2178 585
R1276 gnd.n2178 gnd.n2177 585
R1277 gnd.n3214 gnd.n3213 585
R1278 gnd.n3215 gnd.n3214 585
R1279 gnd.n2176 gnd.n2175 585
R1280 gnd.n3216 gnd.n2176 585
R1281 gnd.n3219 gnd.n3218 585
R1282 gnd.n3218 gnd.n3217 585
R1283 gnd.n2173 gnd.n2172 585
R1284 gnd.n2172 gnd.n2171 585
R1285 gnd.n3224 gnd.n3223 585
R1286 gnd.n3225 gnd.n3224 585
R1287 gnd.n2170 gnd.n2169 585
R1288 gnd.n3226 gnd.n2170 585
R1289 gnd.n3229 gnd.n3228 585
R1290 gnd.n3228 gnd.n3227 585
R1291 gnd.n2167 gnd.n2166 585
R1292 gnd.n2166 gnd.n2165 585
R1293 gnd.n3234 gnd.n3233 585
R1294 gnd.n3235 gnd.n3234 585
R1295 gnd.n2164 gnd.n2163 585
R1296 gnd.n3236 gnd.n2164 585
R1297 gnd.n3239 gnd.n3238 585
R1298 gnd.n3238 gnd.n3237 585
R1299 gnd.n2161 gnd.n2160 585
R1300 gnd.n2160 gnd.n2159 585
R1301 gnd.n3244 gnd.n3243 585
R1302 gnd.n3245 gnd.n3244 585
R1303 gnd.n2158 gnd.n2157 585
R1304 gnd.n3246 gnd.n2158 585
R1305 gnd.n3249 gnd.n3248 585
R1306 gnd.n3248 gnd.n3247 585
R1307 gnd.n2155 gnd.n2154 585
R1308 gnd.n2154 gnd.n2153 585
R1309 gnd.n3254 gnd.n3253 585
R1310 gnd.n3255 gnd.n3254 585
R1311 gnd.n2152 gnd.n2151 585
R1312 gnd.n3256 gnd.n2152 585
R1313 gnd.n3259 gnd.n3258 585
R1314 gnd.n3258 gnd.n3257 585
R1315 gnd.n2149 gnd.n2148 585
R1316 gnd.n2148 gnd.n2147 585
R1317 gnd.n3264 gnd.n3263 585
R1318 gnd.n3265 gnd.n3264 585
R1319 gnd.n2146 gnd.n2145 585
R1320 gnd.n3266 gnd.n2146 585
R1321 gnd.n3269 gnd.n3268 585
R1322 gnd.n3268 gnd.n3267 585
R1323 gnd.n2143 gnd.n2142 585
R1324 gnd.n2142 gnd.n2141 585
R1325 gnd.n3274 gnd.n3273 585
R1326 gnd.n3275 gnd.n3274 585
R1327 gnd.n2140 gnd.n2139 585
R1328 gnd.n3276 gnd.n2140 585
R1329 gnd.n3279 gnd.n3278 585
R1330 gnd.n3278 gnd.n3277 585
R1331 gnd.n2137 gnd.n2136 585
R1332 gnd.n2136 gnd.n2135 585
R1333 gnd.n3284 gnd.n3283 585
R1334 gnd.n3285 gnd.n3284 585
R1335 gnd.n2134 gnd.n2133 585
R1336 gnd.n3286 gnd.n2134 585
R1337 gnd.n3289 gnd.n3288 585
R1338 gnd.n3288 gnd.n3287 585
R1339 gnd.n2131 gnd.n2130 585
R1340 gnd.n2130 gnd.n2129 585
R1341 gnd.n3294 gnd.n3293 585
R1342 gnd.n3295 gnd.n3294 585
R1343 gnd.n2128 gnd.n2127 585
R1344 gnd.n3296 gnd.n2128 585
R1345 gnd.n3299 gnd.n3298 585
R1346 gnd.n3298 gnd.n3297 585
R1347 gnd.n2125 gnd.n2124 585
R1348 gnd.n2124 gnd.n2123 585
R1349 gnd.n3304 gnd.n3303 585
R1350 gnd.n3305 gnd.n3304 585
R1351 gnd.n2122 gnd.n2121 585
R1352 gnd.n3306 gnd.n2122 585
R1353 gnd.n3309 gnd.n3308 585
R1354 gnd.n3308 gnd.n3307 585
R1355 gnd.n2119 gnd.n2118 585
R1356 gnd.n2118 gnd.n2117 585
R1357 gnd.n3314 gnd.n3313 585
R1358 gnd.n3315 gnd.n3314 585
R1359 gnd.n2116 gnd.n2115 585
R1360 gnd.n3316 gnd.n2116 585
R1361 gnd.n3319 gnd.n3318 585
R1362 gnd.n3318 gnd.n3317 585
R1363 gnd.n2113 gnd.n2112 585
R1364 gnd.n2112 gnd.n2111 585
R1365 gnd.n3324 gnd.n3323 585
R1366 gnd.n3325 gnd.n3324 585
R1367 gnd.n2110 gnd.n2109 585
R1368 gnd.n3326 gnd.n2110 585
R1369 gnd.n3329 gnd.n3328 585
R1370 gnd.n3328 gnd.n3327 585
R1371 gnd.n2107 gnd.n2106 585
R1372 gnd.n2106 gnd.n2105 585
R1373 gnd.n3334 gnd.n3333 585
R1374 gnd.n3335 gnd.n3334 585
R1375 gnd.n2104 gnd.n2103 585
R1376 gnd.n3336 gnd.n2104 585
R1377 gnd.n3339 gnd.n3338 585
R1378 gnd.n3338 gnd.n3337 585
R1379 gnd.n2101 gnd.n2100 585
R1380 gnd.n2100 gnd.n2099 585
R1381 gnd.n3344 gnd.n3343 585
R1382 gnd.n3345 gnd.n3344 585
R1383 gnd.n2098 gnd.n2097 585
R1384 gnd.n3346 gnd.n2098 585
R1385 gnd.n3349 gnd.n3348 585
R1386 gnd.n3348 gnd.n3347 585
R1387 gnd.n2095 gnd.n2094 585
R1388 gnd.n2094 gnd.n2093 585
R1389 gnd.n3354 gnd.n3353 585
R1390 gnd.n3355 gnd.n3354 585
R1391 gnd.n2092 gnd.n2091 585
R1392 gnd.n3356 gnd.n2092 585
R1393 gnd.n3359 gnd.n3358 585
R1394 gnd.n3358 gnd.n3357 585
R1395 gnd.n2089 gnd.n2088 585
R1396 gnd.n2088 gnd.n2087 585
R1397 gnd.n3364 gnd.n3363 585
R1398 gnd.n3365 gnd.n3364 585
R1399 gnd.n2086 gnd.n2085 585
R1400 gnd.n3366 gnd.n2086 585
R1401 gnd.n3369 gnd.n3368 585
R1402 gnd.n3368 gnd.n3367 585
R1403 gnd.n2083 gnd.n2075 585
R1404 gnd.n2075 gnd.n2074 585
R1405 gnd.n3376 gnd.n3375 585
R1406 gnd.n3377 gnd.n3376 585
R1407 gnd.n3164 gnd.n3163 585
R1408 gnd.n3165 gnd.n3164 585
R1409 gnd.n2209 gnd.n2208 585
R1410 gnd.n2208 gnd.n2207 585
R1411 gnd.n3159 gnd.n3158 585
R1412 gnd.n3158 gnd.n3157 585
R1413 gnd.n2212 gnd.n2211 585
R1414 gnd.n3156 gnd.n2212 585
R1415 gnd.n3154 gnd.n3153 585
R1416 gnd.n3155 gnd.n3154 585
R1417 gnd.n3152 gnd.n2214 585
R1418 gnd.n2214 gnd.n2213 585
R1419 gnd.n3151 gnd.n3150 585
R1420 gnd.n3150 gnd.n3149 585
R1421 gnd.n2219 gnd.n2218 585
R1422 gnd.n3148 gnd.n2219 585
R1423 gnd.n3146 gnd.n3145 585
R1424 gnd.n3147 gnd.n3146 585
R1425 gnd.n3144 gnd.n2221 585
R1426 gnd.n2221 gnd.n2220 585
R1427 gnd.n3143 gnd.n3142 585
R1428 gnd.n3142 gnd.n3141 585
R1429 gnd.n2227 gnd.n2226 585
R1430 gnd.n3140 gnd.n2227 585
R1431 gnd.n3138 gnd.n3137 585
R1432 gnd.n3139 gnd.n3138 585
R1433 gnd.n3136 gnd.n2229 585
R1434 gnd.n2229 gnd.n2228 585
R1435 gnd.n3135 gnd.n3134 585
R1436 gnd.n3134 gnd.n3133 585
R1437 gnd.n2235 gnd.n2234 585
R1438 gnd.n3132 gnd.n2235 585
R1439 gnd.n3130 gnd.n3129 585
R1440 gnd.n3131 gnd.n3130 585
R1441 gnd.n3128 gnd.n2237 585
R1442 gnd.n2237 gnd.n2236 585
R1443 gnd.n3127 gnd.n3126 585
R1444 gnd.n3126 gnd.n3125 585
R1445 gnd.n2243 gnd.n2242 585
R1446 gnd.n3124 gnd.n2243 585
R1447 gnd.n3122 gnd.n3121 585
R1448 gnd.n3123 gnd.n3122 585
R1449 gnd.n3120 gnd.n2245 585
R1450 gnd.n2245 gnd.n2244 585
R1451 gnd.n3119 gnd.n3118 585
R1452 gnd.n3118 gnd.n3117 585
R1453 gnd.n2251 gnd.n2250 585
R1454 gnd.n3116 gnd.n2251 585
R1455 gnd.n3114 gnd.n3113 585
R1456 gnd.n3115 gnd.n3114 585
R1457 gnd.n3112 gnd.n2253 585
R1458 gnd.n2253 gnd.n2252 585
R1459 gnd.n3111 gnd.n3110 585
R1460 gnd.n3110 gnd.n3109 585
R1461 gnd.n2259 gnd.n2258 585
R1462 gnd.n3108 gnd.n2259 585
R1463 gnd.n3106 gnd.n3105 585
R1464 gnd.n3107 gnd.n3106 585
R1465 gnd.n3104 gnd.n2261 585
R1466 gnd.n2261 gnd.n2260 585
R1467 gnd.n3103 gnd.n3102 585
R1468 gnd.n3102 gnd.n3101 585
R1469 gnd.n2267 gnd.n2266 585
R1470 gnd.n3100 gnd.n2267 585
R1471 gnd.n3098 gnd.n3097 585
R1472 gnd.n3099 gnd.n3098 585
R1473 gnd.n3096 gnd.n2269 585
R1474 gnd.n2269 gnd.n2268 585
R1475 gnd.n3095 gnd.n3094 585
R1476 gnd.n3094 gnd.n3093 585
R1477 gnd.n2275 gnd.n2274 585
R1478 gnd.n3092 gnd.n2275 585
R1479 gnd.n3090 gnd.n3089 585
R1480 gnd.n3091 gnd.n3090 585
R1481 gnd.n3088 gnd.n2277 585
R1482 gnd.n2277 gnd.n2276 585
R1483 gnd.n3087 gnd.n3086 585
R1484 gnd.n3086 gnd.n3085 585
R1485 gnd.n2283 gnd.n2282 585
R1486 gnd.n3084 gnd.n2283 585
R1487 gnd.n3082 gnd.n3081 585
R1488 gnd.n3083 gnd.n3082 585
R1489 gnd.n3080 gnd.n2285 585
R1490 gnd.n2285 gnd.n2284 585
R1491 gnd.n3079 gnd.n3078 585
R1492 gnd.n3078 gnd.n3077 585
R1493 gnd.n2291 gnd.n2290 585
R1494 gnd.n3076 gnd.n2291 585
R1495 gnd.n3074 gnd.n3073 585
R1496 gnd.n3075 gnd.n3074 585
R1497 gnd.n3072 gnd.n2293 585
R1498 gnd.n2293 gnd.n2292 585
R1499 gnd.n3071 gnd.n3070 585
R1500 gnd.n3070 gnd.n3069 585
R1501 gnd.n2299 gnd.n2298 585
R1502 gnd.n3068 gnd.n2299 585
R1503 gnd.n3066 gnd.n3065 585
R1504 gnd.n3067 gnd.n3066 585
R1505 gnd.n3064 gnd.n2301 585
R1506 gnd.n2301 gnd.n2300 585
R1507 gnd.n3063 gnd.n3062 585
R1508 gnd.n3062 gnd.n3061 585
R1509 gnd.n2307 gnd.n2306 585
R1510 gnd.n3060 gnd.n2307 585
R1511 gnd.n3058 gnd.n3057 585
R1512 gnd.n3059 gnd.n3058 585
R1513 gnd.n3056 gnd.n2309 585
R1514 gnd.n2309 gnd.n2308 585
R1515 gnd.n3055 gnd.n3054 585
R1516 gnd.n3054 gnd.n3053 585
R1517 gnd.n2315 gnd.n2314 585
R1518 gnd.n3052 gnd.n2315 585
R1519 gnd.n3050 gnd.n3049 585
R1520 gnd.n3051 gnd.n3050 585
R1521 gnd.n3048 gnd.n2317 585
R1522 gnd.n2317 gnd.n2316 585
R1523 gnd.n3047 gnd.n3046 585
R1524 gnd.n3046 gnd.n3045 585
R1525 gnd.n2323 gnd.n2322 585
R1526 gnd.n3044 gnd.n2323 585
R1527 gnd.n3042 gnd.n3041 585
R1528 gnd.n3043 gnd.n3042 585
R1529 gnd.n3040 gnd.n2325 585
R1530 gnd.n2325 gnd.n2324 585
R1531 gnd.n3039 gnd.n3038 585
R1532 gnd.n3038 gnd.n3037 585
R1533 gnd.n2331 gnd.n2330 585
R1534 gnd.n3036 gnd.n2331 585
R1535 gnd.n3034 gnd.n3033 585
R1536 gnd.n3035 gnd.n3034 585
R1537 gnd.n3032 gnd.n2333 585
R1538 gnd.n2333 gnd.n2332 585
R1539 gnd.n3031 gnd.n3030 585
R1540 gnd.n3030 gnd.n3029 585
R1541 gnd.n2339 gnd.n2338 585
R1542 gnd.n3028 gnd.n2339 585
R1543 gnd.n3026 gnd.n3025 585
R1544 gnd.n3027 gnd.n3026 585
R1545 gnd.n3024 gnd.n2341 585
R1546 gnd.n2341 gnd.n2340 585
R1547 gnd.n3023 gnd.n3022 585
R1548 gnd.n3022 gnd.n3021 585
R1549 gnd.n2347 gnd.n2346 585
R1550 gnd.n3020 gnd.n2347 585
R1551 gnd.n3018 gnd.n3017 585
R1552 gnd.n3019 gnd.n3018 585
R1553 gnd.n3016 gnd.n2349 585
R1554 gnd.n2349 gnd.n2348 585
R1555 gnd.n3015 gnd.n3014 585
R1556 gnd.n3014 gnd.n3013 585
R1557 gnd.n2355 gnd.n2354 585
R1558 gnd.n3012 gnd.n2355 585
R1559 gnd.n3010 gnd.n3009 585
R1560 gnd.n3011 gnd.n3010 585
R1561 gnd.n3008 gnd.n2357 585
R1562 gnd.n2357 gnd.n2356 585
R1563 gnd.n3007 gnd.n3006 585
R1564 gnd.n3006 gnd.n3005 585
R1565 gnd.n2363 gnd.n2362 585
R1566 gnd.n3004 gnd.n2363 585
R1567 gnd.n3002 gnd.n3001 585
R1568 gnd.n3003 gnd.n3002 585
R1569 gnd.n3000 gnd.n2365 585
R1570 gnd.n2365 gnd.n2364 585
R1571 gnd.n2999 gnd.n2998 585
R1572 gnd.n2998 gnd.n2997 585
R1573 gnd.n2371 gnd.n2370 585
R1574 gnd.n2996 gnd.n2371 585
R1575 gnd.n2994 gnd.n2993 585
R1576 gnd.n2995 gnd.n2994 585
R1577 gnd.n2992 gnd.n2373 585
R1578 gnd.n2373 gnd.n2372 585
R1579 gnd.n2991 gnd.n2990 585
R1580 gnd.n2990 gnd.n2989 585
R1581 gnd.n2379 gnd.n2378 585
R1582 gnd.n2988 gnd.n2379 585
R1583 gnd.n2986 gnd.n2985 585
R1584 gnd.n2987 gnd.n2986 585
R1585 gnd.n2984 gnd.n2381 585
R1586 gnd.n2381 gnd.n2380 585
R1587 gnd.n2983 gnd.n2982 585
R1588 gnd.n2982 gnd.n2981 585
R1589 gnd.n2387 gnd.n2386 585
R1590 gnd.n2980 gnd.n2387 585
R1591 gnd.n2978 gnd.n2977 585
R1592 gnd.n2979 gnd.n2978 585
R1593 gnd.n2976 gnd.n2389 585
R1594 gnd.n2389 gnd.n2388 585
R1595 gnd.n2975 gnd.n2974 585
R1596 gnd.n2974 gnd.n2973 585
R1597 gnd.n2395 gnd.n2394 585
R1598 gnd.n2972 gnd.n2395 585
R1599 gnd.n2970 gnd.n2969 585
R1600 gnd.n2971 gnd.n2970 585
R1601 gnd.n2968 gnd.n2397 585
R1602 gnd.n2397 gnd.n2396 585
R1603 gnd.n2967 gnd.n2966 585
R1604 gnd.n2966 gnd.n2965 585
R1605 gnd.n2403 gnd.n2402 585
R1606 gnd.n2964 gnd.n2403 585
R1607 gnd.n2962 gnd.n2961 585
R1608 gnd.n2963 gnd.n2962 585
R1609 gnd.n2960 gnd.n2405 585
R1610 gnd.n2405 gnd.n2404 585
R1611 gnd.n2959 gnd.n2958 585
R1612 gnd.n2958 gnd.n2957 585
R1613 gnd.n2411 gnd.n2410 585
R1614 gnd.n2956 gnd.n2411 585
R1615 gnd.n2954 gnd.n2953 585
R1616 gnd.n2955 gnd.n2954 585
R1617 gnd.n2952 gnd.n2413 585
R1618 gnd.n2413 gnd.n2412 585
R1619 gnd.n2951 gnd.n2950 585
R1620 gnd.n2950 gnd.n2949 585
R1621 gnd.n2419 gnd.n2418 585
R1622 gnd.n2948 gnd.n2419 585
R1623 gnd.n2946 gnd.n2945 585
R1624 gnd.n2947 gnd.n2946 585
R1625 gnd.n2944 gnd.n2421 585
R1626 gnd.n2421 gnd.n2420 585
R1627 gnd.n2943 gnd.n2942 585
R1628 gnd.n2942 gnd.n2941 585
R1629 gnd.n2427 gnd.n2426 585
R1630 gnd.n2940 gnd.n2427 585
R1631 gnd.n2938 gnd.n2937 585
R1632 gnd.n2939 gnd.n2938 585
R1633 gnd.n2936 gnd.n2429 585
R1634 gnd.n2429 gnd.n2428 585
R1635 gnd.n2935 gnd.n2934 585
R1636 gnd.n2934 gnd.n2933 585
R1637 gnd.n2435 gnd.n2434 585
R1638 gnd.n2932 gnd.n2435 585
R1639 gnd.n2930 gnd.n2929 585
R1640 gnd.n2931 gnd.n2930 585
R1641 gnd.n2928 gnd.n2437 585
R1642 gnd.n2437 gnd.n2436 585
R1643 gnd.n2927 gnd.n2926 585
R1644 gnd.n2926 gnd.n2925 585
R1645 gnd.n2443 gnd.n2442 585
R1646 gnd.n2924 gnd.n2443 585
R1647 gnd.n2922 gnd.n2921 585
R1648 gnd.n2923 gnd.n2922 585
R1649 gnd.n2920 gnd.n2445 585
R1650 gnd.n2445 gnd.n2444 585
R1651 gnd.n2919 gnd.n2918 585
R1652 gnd.n2918 gnd.n2917 585
R1653 gnd.n2451 gnd.n2450 585
R1654 gnd.n2916 gnd.n2451 585
R1655 gnd.n2914 gnd.n2913 585
R1656 gnd.n2915 gnd.n2914 585
R1657 gnd.n2912 gnd.n2453 585
R1658 gnd.n2453 gnd.n2452 585
R1659 gnd.n2911 gnd.n2910 585
R1660 gnd.n2910 gnd.n2909 585
R1661 gnd.n2459 gnd.n2458 585
R1662 gnd.n2908 gnd.n2459 585
R1663 gnd.n2906 gnd.n2905 585
R1664 gnd.n2907 gnd.n2906 585
R1665 gnd.n2904 gnd.n2461 585
R1666 gnd.n2461 gnd.n2460 585
R1667 gnd.n2903 gnd.n2902 585
R1668 gnd.n2902 gnd.n2901 585
R1669 gnd.n2467 gnd.n2466 585
R1670 gnd.n2900 gnd.n2467 585
R1671 gnd.n2898 gnd.n2897 585
R1672 gnd.n2899 gnd.n2898 585
R1673 gnd.n2896 gnd.n2469 585
R1674 gnd.n2469 gnd.n2468 585
R1675 gnd.n2895 gnd.n2894 585
R1676 gnd.n2894 gnd.n2893 585
R1677 gnd.n2475 gnd.n2474 585
R1678 gnd.n2892 gnd.n2475 585
R1679 gnd.n2890 gnd.n2889 585
R1680 gnd.n2891 gnd.n2890 585
R1681 gnd.n2888 gnd.n2477 585
R1682 gnd.n2477 gnd.n2476 585
R1683 gnd.n2887 gnd.n2886 585
R1684 gnd.n2886 gnd.n2885 585
R1685 gnd.n2483 gnd.n2482 585
R1686 gnd.n2884 gnd.n2483 585
R1687 gnd.n2882 gnd.n2881 585
R1688 gnd.n2883 gnd.n2882 585
R1689 gnd.n2880 gnd.n2485 585
R1690 gnd.n2485 gnd.n2484 585
R1691 gnd.n2879 gnd.n2878 585
R1692 gnd.n2878 gnd.n2877 585
R1693 gnd.n2491 gnd.n2490 585
R1694 gnd.n2876 gnd.n2491 585
R1695 gnd.n2874 gnd.n2873 585
R1696 gnd.n2875 gnd.n2874 585
R1697 gnd.n2872 gnd.n2493 585
R1698 gnd.n2493 gnd.n2492 585
R1699 gnd.n2871 gnd.n2870 585
R1700 gnd.n2870 gnd.n2869 585
R1701 gnd.n2499 gnd.n2498 585
R1702 gnd.n2868 gnd.n2499 585
R1703 gnd.n2866 gnd.n2865 585
R1704 gnd.n2867 gnd.n2866 585
R1705 gnd.n2864 gnd.n2501 585
R1706 gnd.n2501 gnd.n2500 585
R1707 gnd.n2863 gnd.n2862 585
R1708 gnd.n2862 gnd.n2861 585
R1709 gnd.n2507 gnd.n2506 585
R1710 gnd.n2860 gnd.n2507 585
R1711 gnd.n2858 gnd.n2857 585
R1712 gnd.n2859 gnd.n2858 585
R1713 gnd.n2856 gnd.n2509 585
R1714 gnd.n2509 gnd.n2508 585
R1715 gnd.n2855 gnd.n2854 585
R1716 gnd.n2854 gnd.n2853 585
R1717 gnd.n2685 gnd.n2684 585
R1718 gnd.n2684 gnd.n2683 585
R1719 gnd.n2686 gnd.n2675 585
R1720 gnd.n2675 gnd.n2674 585
R1721 gnd.n2688 gnd.n2687 585
R1722 gnd.n2689 gnd.n2688 585
R1723 gnd.n2673 gnd.n2672 585
R1724 gnd.n2690 gnd.n2673 585
R1725 gnd.n2693 gnd.n2692 585
R1726 gnd.n2692 gnd.n2691 585
R1727 gnd.n2694 gnd.n2667 585
R1728 gnd.n2667 gnd.n2666 585
R1729 gnd.n2696 gnd.n2695 585
R1730 gnd.n2697 gnd.n2696 585
R1731 gnd.n2665 gnd.n2664 585
R1732 gnd.n2698 gnd.n2665 585
R1733 gnd.n2701 gnd.n2700 585
R1734 gnd.n2700 gnd.n2699 585
R1735 gnd.n2702 gnd.n2659 585
R1736 gnd.n2659 gnd.n2658 585
R1737 gnd.n2704 gnd.n2703 585
R1738 gnd.n2705 gnd.n2704 585
R1739 gnd.n2657 gnd.n2656 585
R1740 gnd.n2706 gnd.n2657 585
R1741 gnd.n2709 gnd.n2708 585
R1742 gnd.n2708 gnd.n2707 585
R1743 gnd.n2710 gnd.n2651 585
R1744 gnd.n2651 gnd.n2650 585
R1745 gnd.n2712 gnd.n2711 585
R1746 gnd.n2713 gnd.n2712 585
R1747 gnd.n2649 gnd.n2648 585
R1748 gnd.n2714 gnd.n2649 585
R1749 gnd.n2717 gnd.n2716 585
R1750 gnd.n2716 gnd.n2715 585
R1751 gnd.n2718 gnd.n2643 585
R1752 gnd.n2643 gnd.n2642 585
R1753 gnd.n2720 gnd.n2719 585
R1754 gnd.n2721 gnd.n2720 585
R1755 gnd.n2641 gnd.n2640 585
R1756 gnd.n2722 gnd.n2641 585
R1757 gnd.n2725 gnd.n2724 585
R1758 gnd.n2724 gnd.n2723 585
R1759 gnd.n2726 gnd.n2635 585
R1760 gnd.n2635 gnd.n2634 585
R1761 gnd.n2728 gnd.n2727 585
R1762 gnd.n2729 gnd.n2728 585
R1763 gnd.n2633 gnd.n2632 585
R1764 gnd.n2730 gnd.n2633 585
R1765 gnd.n2733 gnd.n2732 585
R1766 gnd.n2732 gnd.n2731 585
R1767 gnd.n2734 gnd.n2627 585
R1768 gnd.n2627 gnd.n2626 585
R1769 gnd.n2736 gnd.n2735 585
R1770 gnd.n2737 gnd.n2736 585
R1771 gnd.n2625 gnd.n2624 585
R1772 gnd.n2738 gnd.n2625 585
R1773 gnd.n2741 gnd.n2740 585
R1774 gnd.n2740 gnd.n2739 585
R1775 gnd.n2742 gnd.n2619 585
R1776 gnd.n2619 gnd.n2618 585
R1777 gnd.n2744 gnd.n2743 585
R1778 gnd.n2745 gnd.n2744 585
R1779 gnd.n2617 gnd.n2616 585
R1780 gnd.n2746 gnd.n2617 585
R1781 gnd.n2749 gnd.n2748 585
R1782 gnd.n2748 gnd.n2747 585
R1783 gnd.n2750 gnd.n2611 585
R1784 gnd.n2611 gnd.n2610 585
R1785 gnd.n2752 gnd.n2751 585
R1786 gnd.n2753 gnd.n2752 585
R1787 gnd.n2609 gnd.n2608 585
R1788 gnd.n2754 gnd.n2609 585
R1789 gnd.n2757 gnd.n2756 585
R1790 gnd.n2756 gnd.n2755 585
R1791 gnd.n2758 gnd.n2603 585
R1792 gnd.n2603 gnd.n2602 585
R1793 gnd.n2760 gnd.n2759 585
R1794 gnd.n2761 gnd.n2760 585
R1795 gnd.n2601 gnd.n2600 585
R1796 gnd.n2762 gnd.n2601 585
R1797 gnd.n2765 gnd.n2764 585
R1798 gnd.n2764 gnd.n2763 585
R1799 gnd.n2766 gnd.n2595 585
R1800 gnd.n2595 gnd.n2594 585
R1801 gnd.n2768 gnd.n2767 585
R1802 gnd.n2769 gnd.n2768 585
R1803 gnd.n2593 gnd.n2592 585
R1804 gnd.n2770 gnd.n2593 585
R1805 gnd.n2773 gnd.n2772 585
R1806 gnd.n2772 gnd.n2771 585
R1807 gnd.n2774 gnd.n2587 585
R1808 gnd.n2587 gnd.n2586 585
R1809 gnd.n2776 gnd.n2775 585
R1810 gnd.n2777 gnd.n2776 585
R1811 gnd.n2585 gnd.n2584 585
R1812 gnd.n2778 gnd.n2585 585
R1813 gnd.n2781 gnd.n2780 585
R1814 gnd.n2780 gnd.n2779 585
R1815 gnd.n2782 gnd.n2579 585
R1816 gnd.n2579 gnd.n2578 585
R1817 gnd.n2784 gnd.n2783 585
R1818 gnd.n2785 gnd.n2784 585
R1819 gnd.n2577 gnd.n2576 585
R1820 gnd.n2786 gnd.n2577 585
R1821 gnd.n2789 gnd.n2788 585
R1822 gnd.n2788 gnd.n2787 585
R1823 gnd.n2790 gnd.n2571 585
R1824 gnd.n2571 gnd.n2570 585
R1825 gnd.n2792 gnd.n2791 585
R1826 gnd.n2793 gnd.n2792 585
R1827 gnd.n2569 gnd.n2568 585
R1828 gnd.n2794 gnd.n2569 585
R1829 gnd.n2797 gnd.n2796 585
R1830 gnd.n2796 gnd.n2795 585
R1831 gnd.n2798 gnd.n2563 585
R1832 gnd.n2563 gnd.n2562 585
R1833 gnd.n2800 gnd.n2799 585
R1834 gnd.n2801 gnd.n2800 585
R1835 gnd.n2561 gnd.n2560 585
R1836 gnd.n2802 gnd.n2561 585
R1837 gnd.n2805 gnd.n2804 585
R1838 gnd.n2804 gnd.n2803 585
R1839 gnd.n2806 gnd.n2555 585
R1840 gnd.n2555 gnd.n2554 585
R1841 gnd.n2808 gnd.n2807 585
R1842 gnd.n2809 gnd.n2808 585
R1843 gnd.n2553 gnd.n2552 585
R1844 gnd.n2810 gnd.n2553 585
R1845 gnd.n2813 gnd.n2812 585
R1846 gnd.n2812 gnd.n2811 585
R1847 gnd.n2814 gnd.n2547 585
R1848 gnd.n2547 gnd.n2546 585
R1849 gnd.n2816 gnd.n2815 585
R1850 gnd.n2817 gnd.n2816 585
R1851 gnd.n2545 gnd.n2544 585
R1852 gnd.n2818 gnd.n2545 585
R1853 gnd.n2821 gnd.n2820 585
R1854 gnd.n2820 gnd.n2819 585
R1855 gnd.n2822 gnd.n2539 585
R1856 gnd.n2539 gnd.n2538 585
R1857 gnd.n2824 gnd.n2823 585
R1858 gnd.n2825 gnd.n2824 585
R1859 gnd.n2537 gnd.n2536 585
R1860 gnd.n2826 gnd.n2537 585
R1861 gnd.n2829 gnd.n2828 585
R1862 gnd.n2828 gnd.n2827 585
R1863 gnd.n2830 gnd.n2531 585
R1864 gnd.n2531 gnd.n2530 585
R1865 gnd.n2832 gnd.n2831 585
R1866 gnd.n2833 gnd.n2832 585
R1867 gnd.n2529 gnd.n2528 585
R1868 gnd.n2834 gnd.n2529 585
R1869 gnd.n2837 gnd.n2836 585
R1870 gnd.n2836 gnd.n2835 585
R1871 gnd.n2838 gnd.n2524 585
R1872 gnd.n2524 gnd.n2523 585
R1873 gnd.n2840 gnd.n2839 585
R1874 gnd.n2841 gnd.n2840 585
R1875 gnd.n2522 gnd.n2521 585
R1876 gnd.n2842 gnd.n2522 585
R1877 gnd.n2845 gnd.n2844 585
R1878 gnd.n2844 gnd.n2843 585
R1879 gnd.n2518 gnd.n2516 585
R1880 gnd.n2516 gnd.n2515 585
R1881 gnd.n2850 gnd.n2849 585
R1882 gnd.n2851 gnd.n2850 585
R1883 gnd.n2517 gnd.n2514 585
R1884 gnd.n2852 gnd.n2514 585
R1885 gnd.n5597 gnd.n1651 585
R1886 gnd.n5597 gnd.n5596 585
R1887 gnd.n5758 gnd.n1657 585
R1888 gnd.n5864 gnd.n1657 585
R1889 gnd.n5759 gnd.n1669 585
R1890 gnd.n1680 gnd.n1669 585
R1891 gnd.n5761 gnd.n5760 585
R1892 gnd.n5762 gnd.n5761 585
R1893 gnd.n1670 gnd.n1668 585
R1894 gnd.n5752 gnd.n1668 585
R1895 gnd.n5411 gnd.n1727 585
R1896 gnd.n5423 gnd.n1727 585
R1897 gnd.n5412 gnd.n1738 585
R1898 gnd.n1738 gnd.n1726 585
R1899 gnd.n5414 gnd.n5413 585
R1900 gnd.n5415 gnd.n5414 585
R1901 gnd.n1739 gnd.n1737 585
R1902 gnd.n5403 gnd.n1737 585
R1903 gnd.n5376 gnd.n5375 585
R1904 gnd.n5375 gnd.n5374 585
R1905 gnd.n5377 gnd.n1753 585
R1906 gnd.n5391 gnd.n1753 585
R1907 gnd.n5378 gnd.n1764 585
R1908 gnd.n5359 gnd.n1764 585
R1909 gnd.n5380 gnd.n5379 585
R1910 gnd.n5381 gnd.n5380 585
R1911 gnd.n1765 gnd.n1763 585
R1912 gnd.n5352 gnd.n1763 585
R1913 gnd.n5328 gnd.n5327 585
R1914 gnd.n5327 gnd.n5326 585
R1915 gnd.n5329 gnd.n1788 585
R1916 gnd.n5343 gnd.n1788 585
R1917 gnd.n5330 gnd.n1800 585
R1918 gnd.n5279 gnd.n1800 585
R1919 gnd.n5332 gnd.n5331 585
R1920 gnd.n5333 gnd.n5332 585
R1921 gnd.n1801 gnd.n1799 585
R1922 gnd.n5312 gnd.n1799 585
R1923 gnd.n5288 gnd.n5287 585
R1924 gnd.n5287 gnd.n1813 585
R1925 gnd.n5289 gnd.n1824 585
R1926 gnd.n5303 gnd.n1824 585
R1927 gnd.n5290 gnd.n1841 585
R1928 gnd.n5274 gnd.n1841 585
R1929 gnd.n5292 gnd.n5291 585
R1930 gnd.n5293 gnd.n5292 585
R1931 gnd.n1842 gnd.n1840 585
R1932 gnd.n5270 gnd.n1840 585
R1933 gnd.n5251 gnd.n5250 585
R1934 gnd.n5250 gnd.n1850 585
R1935 gnd.n5252 gnd.n1858 585
R1936 gnd.n5261 gnd.n1858 585
R1937 gnd.n5254 gnd.n5253 585
R1938 gnd.n5255 gnd.n5254 585
R1939 gnd.n1865 gnd.n1864 585
R1940 gnd.n1864 gnd.n1862 585
R1941 gnd.n5233 gnd.n1872 585
R1942 gnd.n5242 gnd.n1872 585
R1943 gnd.n5234 gnd.n1878 585
R1944 gnd.n1878 gnd.n1870 585
R1945 gnd.n5236 gnd.n5235 585
R1946 gnd.n5237 gnd.n5236 585
R1947 gnd.n1879 gnd.n1877 585
R1948 gnd.n5226 gnd.n1877 585
R1949 gnd.n5192 gnd.n5191 585
R1950 gnd.n5191 gnd.n1884 585
R1951 gnd.n5193 gnd.n1891 585
R1952 gnd.n5207 gnd.n1891 585
R1953 gnd.n5194 gnd.n1902 585
R1954 gnd.n1902 gnd.n1900 585
R1955 gnd.n5196 gnd.n5195 585
R1956 gnd.n5197 gnd.n5196 585
R1957 gnd.n1903 gnd.n1901 585
R1958 gnd.n5182 gnd.n1901 585
R1959 gnd.n5157 gnd.n5156 585
R1960 gnd.n5156 gnd.n1909 585
R1961 gnd.n5158 gnd.n1916 585
R1962 gnd.n5172 gnd.n1916 585
R1963 gnd.n5159 gnd.n1928 585
R1964 gnd.n1928 gnd.n1926 585
R1965 gnd.n5161 gnd.n5160 585
R1966 gnd.n5162 gnd.n5161 585
R1967 gnd.n1929 gnd.n1927 585
R1968 gnd.n1927 gnd.n1923 585
R1969 gnd.n5134 gnd.n1937 585
R1970 gnd.n5146 gnd.n1937 585
R1971 gnd.n5135 gnd.n1947 585
R1972 gnd.n1947 gnd.n1935 585
R1973 gnd.n5137 gnd.n5136 585
R1974 gnd.n5138 gnd.n5137 585
R1975 gnd.n1948 gnd.n1946 585
R1976 gnd.n1946 gnd.n1943 585
R1977 gnd.n5114 gnd.n1954 585
R1978 gnd.n5126 gnd.n1954 585
R1979 gnd.n5115 gnd.n1965 585
R1980 gnd.n1965 gnd.n1963 585
R1981 gnd.n5117 gnd.n5116 585
R1982 gnd.n5118 gnd.n5117 585
R1983 gnd.n1966 gnd.n1964 585
R1984 gnd.n1964 gnd.n1960 585
R1985 gnd.n1987 gnd.n1973 585
R1986 gnd.n5106 gnd.n1973 585
R1987 gnd.n1985 gnd.n1983 585
R1988 gnd.n1983 gnd.n1971 585
R1989 gnd.n5097 gnd.n5096 585
R1990 gnd.n5098 gnd.n5097 585
R1991 gnd.n1984 gnd.n1982 585
R1992 gnd.n1982 gnd.n1979 585
R1993 gnd.n4968 gnd.n4967 585
R1994 gnd.n4966 gnd.n4965 585
R1995 gnd.n4964 gnd.n4963 585
R1996 gnd.n4962 gnd.n4961 585
R1997 gnd.n4960 gnd.n4959 585
R1998 gnd.n4958 gnd.n4957 585
R1999 gnd.n4956 gnd.n4955 585
R2000 gnd.n4954 gnd.n4953 585
R2001 gnd.n4952 gnd.n4951 585
R2002 gnd.n4950 gnd.n4949 585
R2003 gnd.n4948 gnd.n4947 585
R2004 gnd.n4946 gnd.n4945 585
R2005 gnd.n4944 gnd.n4943 585
R2006 gnd.n4942 gnd.n4941 585
R2007 gnd.n4940 gnd.n4939 585
R2008 gnd.n4938 gnd.n4937 585
R2009 gnd.n4936 gnd.n4935 585
R2010 gnd.n4895 gnd.n4892 585
R2011 gnd.n4931 gnd.n4811 585
R2012 gnd.n5088 gnd.n4811 585
R2013 gnd.n5665 gnd.n5664 585
R2014 gnd.n5666 gnd.n5662 585
R2015 gnd.n5677 gnd.n5659 585
R2016 gnd.n5678 gnd.n5657 585
R2017 gnd.n5656 gnd.n5649 585
R2018 gnd.n5685 gnd.n5648 585
R2019 gnd.n5686 gnd.n5647 585
R2020 gnd.n5645 gnd.n5637 585
R2021 gnd.n5693 gnd.n5636 585
R2022 gnd.n5694 gnd.n5634 585
R2023 gnd.n5633 gnd.n5626 585
R2024 gnd.n5701 gnd.n5625 585
R2025 gnd.n5702 gnd.n5624 585
R2026 gnd.n5622 gnd.n5614 585
R2027 gnd.n5709 gnd.n5613 585
R2028 gnd.n5710 gnd.n5611 585
R2029 gnd.n5610 gnd.n5600 585
R2030 gnd.n5717 gnd.n5599 585
R2031 gnd.n5718 gnd.n5598 585
R2032 gnd.n5598 gnd.n1597 585
R2033 gnd.n5744 gnd.n1682 585
R2034 gnd.n5596 gnd.n1682 585
R2035 gnd.n5745 gnd.n1655 585
R2036 gnd.n5864 gnd.n1655 585
R2037 gnd.n5746 gnd.n1681 585
R2038 gnd.n1681 gnd.n1680 585
R2039 gnd.n1677 gnd.n1666 585
R2040 gnd.n5762 gnd.n1666 585
R2041 gnd.n5751 gnd.n5750 585
R2042 gnd.n5752 gnd.n5751 585
R2043 gnd.n1676 gnd.n1675 585
R2044 gnd.n5423 gnd.n1675 585
R2045 gnd.n5397 gnd.n5396 585
R2046 gnd.n5396 gnd.n1726 585
R2047 gnd.n1747 gnd.n1735 585
R2048 gnd.n5415 gnd.n1735 585
R2049 gnd.n5402 gnd.n5401 585
R2050 gnd.n5403 gnd.n5402 585
R2051 gnd.n1746 gnd.n1745 585
R2052 gnd.n5374 gnd.n1745 585
R2053 gnd.n5393 gnd.n5392 585
R2054 gnd.n5392 gnd.n5391 585
R2055 gnd.n1750 gnd.n1749 585
R2056 gnd.n5359 gnd.n1750 585
R2057 gnd.n1782 gnd.n1762 585
R2058 gnd.n5381 gnd.n1762 585
R2059 gnd.n5351 gnd.n5350 585
R2060 gnd.n5352 gnd.n5351 585
R2061 gnd.n1781 gnd.n1780 585
R2062 gnd.n5326 gnd.n1780 585
R2063 gnd.n5345 gnd.n5344 585
R2064 gnd.n5344 gnd.n5343 585
R2065 gnd.n1785 gnd.n1784 585
R2066 gnd.n5279 gnd.n1785 585
R2067 gnd.n1817 gnd.n1797 585
R2068 gnd.n5333 gnd.n1797 585
R2069 gnd.n5311 gnd.n5310 585
R2070 gnd.n5312 gnd.n5311 585
R2071 gnd.n1816 gnd.n1815 585
R2072 gnd.n1815 gnd.n1813 585
R2073 gnd.n5305 gnd.n5304 585
R2074 gnd.n5304 gnd.n5303 585
R2075 gnd.n1820 gnd.n1819 585
R2076 gnd.n5274 gnd.n1820 585
R2077 gnd.n1853 gnd.n1838 585
R2078 gnd.n5293 gnd.n1838 585
R2079 gnd.n5269 gnd.n5268 585
R2080 gnd.n5270 gnd.n5269 585
R2081 gnd.n1852 gnd.n1851 585
R2082 gnd.n1851 gnd.n1850 585
R2083 gnd.n5263 gnd.n5262 585
R2084 gnd.n5262 gnd.n5261 585
R2085 gnd.n1856 gnd.n1855 585
R2086 gnd.n5255 gnd.n1856 585
R2087 gnd.n5219 gnd.n5218 585
R2088 gnd.n5218 gnd.n1862 585
R2089 gnd.n5220 gnd.n1871 585
R2090 gnd.n5242 gnd.n1871 585
R2091 gnd.n5222 gnd.n5221 585
R2092 gnd.n5221 gnd.n1870 585
R2093 gnd.n5223 gnd.n1876 585
R2094 gnd.n5237 gnd.n1876 585
R2095 gnd.n5225 gnd.n5224 585
R2096 gnd.n5226 gnd.n5225 585
R2097 gnd.n1886 gnd.n1885 585
R2098 gnd.n1885 gnd.n1884 585
R2099 gnd.n5209 gnd.n5208 585
R2100 gnd.n5208 gnd.n5207 585
R2101 gnd.n1889 gnd.n1888 585
R2102 gnd.n1900 gnd.n1889 585
R2103 gnd.n5179 gnd.n1899 585
R2104 gnd.n5197 gnd.n1899 585
R2105 gnd.n5181 gnd.n5180 585
R2106 gnd.n5182 gnd.n5181 585
R2107 gnd.n1911 gnd.n1910 585
R2108 gnd.n1910 gnd.n1909 585
R2109 gnd.n5174 gnd.n5173 585
R2110 gnd.n5173 gnd.n5172 585
R2111 gnd.n1914 gnd.n1913 585
R2112 gnd.n1926 gnd.n1914 585
R2113 gnd.n4909 gnd.n1925 585
R2114 gnd.n5162 gnd.n1925 585
R2115 gnd.n4911 gnd.n4910 585
R2116 gnd.n4910 gnd.n1923 585
R2117 gnd.n4912 gnd.n1936 585
R2118 gnd.n5146 gnd.n1936 585
R2119 gnd.n4914 gnd.n4913 585
R2120 gnd.n4913 gnd.n1935 585
R2121 gnd.n4915 gnd.n1945 585
R2122 gnd.n5138 gnd.n1945 585
R2123 gnd.n4917 gnd.n4916 585
R2124 gnd.n4916 gnd.n1943 585
R2125 gnd.n4918 gnd.n1953 585
R2126 gnd.n5126 gnd.n1953 585
R2127 gnd.n4920 gnd.n4919 585
R2128 gnd.n4919 gnd.n1963 585
R2129 gnd.n4921 gnd.n1962 585
R2130 gnd.n5118 gnd.n1962 585
R2131 gnd.n4923 gnd.n4922 585
R2132 gnd.n4922 gnd.n1960 585
R2133 gnd.n4924 gnd.n1972 585
R2134 gnd.n5106 gnd.n1972 585
R2135 gnd.n4926 gnd.n4925 585
R2136 gnd.n4925 gnd.n1971 585
R2137 gnd.n4927 gnd.n1981 585
R2138 gnd.n5098 gnd.n1981 585
R2139 gnd.n4929 gnd.n4928 585
R2140 gnd.n4928 gnd.n1979 585
R2141 gnd.n4682 gnd.n4681 585
R2142 gnd.n4683 gnd.n4682 585
R2143 gnd.n2068 gnd.n2067 585
R2144 gnd.n3379 gnd.n2067 585
R2145 gnd.n4657 gnd.n3391 585
R2146 gnd.n3391 gnd.n2073 585
R2147 gnd.n4659 gnd.n4658 585
R2148 gnd.n4660 gnd.n4659 585
R2149 gnd.n3392 gnd.n3390 585
R2150 gnd.n3390 gnd.n3386 585
R2151 gnd.n4391 gnd.n4390 585
R2152 gnd.n4390 gnd.n4389 585
R2153 gnd.n3397 gnd.n3396 585
R2154 gnd.n4360 gnd.n3397 585
R2155 gnd.n4380 gnd.n4379 585
R2156 gnd.n4379 gnd.n4378 585
R2157 gnd.n3404 gnd.n3403 585
R2158 gnd.n4366 gnd.n3404 585
R2159 gnd.n4336 gnd.n3424 585
R2160 gnd.n3424 gnd.n3423 585
R2161 gnd.n4338 gnd.n4337 585
R2162 gnd.n4339 gnd.n4338 585
R2163 gnd.n3425 gnd.n3422 585
R2164 gnd.n3433 gnd.n3422 585
R2165 gnd.n4314 gnd.n3445 585
R2166 gnd.n3445 gnd.n3432 585
R2167 gnd.n4316 gnd.n4315 585
R2168 gnd.n4317 gnd.n4316 585
R2169 gnd.n3446 gnd.n3444 585
R2170 gnd.n3444 gnd.n3440 585
R2171 gnd.n4302 gnd.n4301 585
R2172 gnd.n4301 gnd.n4300 585
R2173 gnd.n3451 gnd.n3450 585
R2174 gnd.n3461 gnd.n3451 585
R2175 gnd.n4291 gnd.n4290 585
R2176 gnd.n4290 gnd.n4289 585
R2177 gnd.n3458 gnd.n3457 585
R2178 gnd.n4277 gnd.n3458 585
R2179 gnd.n4251 gnd.n3479 585
R2180 gnd.n3479 gnd.n3468 585
R2181 gnd.n4253 gnd.n4252 585
R2182 gnd.n4254 gnd.n4253 585
R2183 gnd.n3480 gnd.n3478 585
R2184 gnd.n3488 gnd.n3478 585
R2185 gnd.n4229 gnd.n3500 585
R2186 gnd.n3500 gnd.n3487 585
R2187 gnd.n4231 gnd.n4230 585
R2188 gnd.n4232 gnd.n4231 585
R2189 gnd.n3501 gnd.n3499 585
R2190 gnd.n3499 gnd.n3495 585
R2191 gnd.n4217 gnd.n4216 585
R2192 gnd.n4216 gnd.n4215 585
R2193 gnd.n3506 gnd.n3505 585
R2194 gnd.n3515 gnd.n3506 585
R2195 gnd.n4206 gnd.n4205 585
R2196 gnd.n4205 gnd.n4204 585
R2197 gnd.n3513 gnd.n3512 585
R2198 gnd.n4192 gnd.n3513 585
R2199 gnd.n3630 gnd.n3629 585
R2200 gnd.n3630 gnd.n3522 585
R2201 gnd.n4149 gnd.n4148 585
R2202 gnd.n4148 gnd.n4147 585
R2203 gnd.n4150 gnd.n3624 585
R2204 gnd.n3635 gnd.n3624 585
R2205 gnd.n4152 gnd.n4151 585
R2206 gnd.n4153 gnd.n4152 585
R2207 gnd.n3625 gnd.n3623 585
R2208 gnd.n3648 gnd.n3623 585
R2209 gnd.n3608 gnd.n3607 585
R2210 gnd.n3611 gnd.n3608 585
R2211 gnd.n4163 gnd.n4162 585
R2212 gnd.n4162 gnd.n4161 585
R2213 gnd.n4164 gnd.n3602 585
R2214 gnd.n4123 gnd.n3602 585
R2215 gnd.n4166 gnd.n4165 585
R2216 gnd.n4167 gnd.n4166 585
R2217 gnd.n3603 gnd.n3601 585
R2218 gnd.n3662 gnd.n3601 585
R2219 gnd.n4115 gnd.n4114 585
R2220 gnd.n4114 gnd.n4113 585
R2221 gnd.n3659 gnd.n3658 585
R2222 gnd.n4097 gnd.n3659 585
R2223 gnd.n4084 gnd.n3678 585
R2224 gnd.n3678 gnd.n3677 585
R2225 gnd.n4086 gnd.n4085 585
R2226 gnd.n4087 gnd.n4086 585
R2227 gnd.n3679 gnd.n3676 585
R2228 gnd.n3685 gnd.n3676 585
R2229 gnd.n4065 gnd.n4064 585
R2230 gnd.n4066 gnd.n4065 585
R2231 gnd.n3696 gnd.n3695 585
R2232 gnd.n3695 gnd.n3691 585
R2233 gnd.n4055 gnd.n4054 585
R2234 gnd.n4056 gnd.n4055 585
R2235 gnd.n3706 gnd.n3705 585
R2236 gnd.n3711 gnd.n3705 585
R2237 gnd.n4033 gnd.n3724 585
R2238 gnd.n3724 gnd.n3710 585
R2239 gnd.n4035 gnd.n4034 585
R2240 gnd.n4036 gnd.n4035 585
R2241 gnd.n3725 gnd.n3723 585
R2242 gnd.n3723 gnd.n3719 585
R2243 gnd.n4024 gnd.n4023 585
R2244 gnd.n4025 gnd.n4024 585
R2245 gnd.n3732 gnd.n3731 585
R2246 gnd.n3736 gnd.n3731 585
R2247 gnd.n4001 gnd.n3753 585
R2248 gnd.n3753 gnd.n3735 585
R2249 gnd.n4003 gnd.n4002 585
R2250 gnd.n4004 gnd.n4003 585
R2251 gnd.n3754 gnd.n3752 585
R2252 gnd.n3752 gnd.n3743 585
R2253 gnd.n3996 gnd.n3995 585
R2254 gnd.n3995 gnd.n3994 585
R2255 gnd.n3801 gnd.n3800 585
R2256 gnd.n3802 gnd.n3801 585
R2257 gnd.n3955 gnd.n3954 585
R2258 gnd.n3956 gnd.n3955 585
R2259 gnd.n3811 gnd.n3810 585
R2260 gnd.n3810 gnd.n3809 585
R2261 gnd.n3950 gnd.n3949 585
R2262 gnd.n3949 gnd.n3948 585
R2263 gnd.n3814 gnd.n3813 585
R2264 gnd.n3815 gnd.n3814 585
R2265 gnd.n3939 gnd.n3938 585
R2266 gnd.n3940 gnd.n3939 585
R2267 gnd.n3822 gnd.n3821 585
R2268 gnd.n3931 gnd.n3821 585
R2269 gnd.n3934 gnd.n3933 585
R2270 gnd.n3933 gnd.n3932 585
R2271 gnd.n3825 gnd.n3824 585
R2272 gnd.n3826 gnd.n3825 585
R2273 gnd.n3920 gnd.n3919 585
R2274 gnd.n3918 gnd.n3844 585
R2275 gnd.n3917 gnd.n3843 585
R2276 gnd.n3922 gnd.n3843 585
R2277 gnd.n3916 gnd.n3915 585
R2278 gnd.n3914 gnd.n3913 585
R2279 gnd.n3912 gnd.n3911 585
R2280 gnd.n3910 gnd.n3909 585
R2281 gnd.n3908 gnd.n3907 585
R2282 gnd.n3906 gnd.n3905 585
R2283 gnd.n3904 gnd.n3903 585
R2284 gnd.n3902 gnd.n3901 585
R2285 gnd.n3900 gnd.n3899 585
R2286 gnd.n3898 gnd.n3897 585
R2287 gnd.n3896 gnd.n3895 585
R2288 gnd.n3894 gnd.n3893 585
R2289 gnd.n3892 gnd.n3891 585
R2290 gnd.n3890 gnd.n3889 585
R2291 gnd.n3888 gnd.n3887 585
R2292 gnd.n3886 gnd.n3885 585
R2293 gnd.n3884 gnd.n3883 585
R2294 gnd.n3882 gnd.n3881 585
R2295 gnd.n3880 gnd.n3879 585
R2296 gnd.n3878 gnd.n3877 585
R2297 gnd.n3876 gnd.n3875 585
R2298 gnd.n3874 gnd.n3873 585
R2299 gnd.n3831 gnd.n3830 585
R2300 gnd.n3925 gnd.n3924 585
R2301 gnd.n4686 gnd.n4685 585
R2302 gnd.n4688 gnd.n4687 585
R2303 gnd.n4690 gnd.n4689 585
R2304 gnd.n4692 gnd.n4691 585
R2305 gnd.n4694 gnd.n4693 585
R2306 gnd.n4696 gnd.n4695 585
R2307 gnd.n4698 gnd.n4697 585
R2308 gnd.n4700 gnd.n4699 585
R2309 gnd.n4702 gnd.n4701 585
R2310 gnd.n4704 gnd.n4703 585
R2311 gnd.n4706 gnd.n4705 585
R2312 gnd.n4708 gnd.n4707 585
R2313 gnd.n4710 gnd.n4709 585
R2314 gnd.n4712 gnd.n4711 585
R2315 gnd.n4714 gnd.n4713 585
R2316 gnd.n4716 gnd.n4715 585
R2317 gnd.n4718 gnd.n4717 585
R2318 gnd.n4720 gnd.n4719 585
R2319 gnd.n4722 gnd.n4721 585
R2320 gnd.n4724 gnd.n4723 585
R2321 gnd.n4726 gnd.n4725 585
R2322 gnd.n4728 gnd.n4727 585
R2323 gnd.n4730 gnd.n4729 585
R2324 gnd.n4732 gnd.n4731 585
R2325 gnd.n4734 gnd.n4733 585
R2326 gnd.n4735 gnd.n2035 585
R2327 gnd.n4736 gnd.n1993 585
R2328 gnd.n4774 gnd.n1993 585
R2329 gnd.n4684 gnd.n2065 585
R2330 gnd.n4684 gnd.n4683 585
R2331 gnd.n4353 gnd.n2064 585
R2332 gnd.n3379 gnd.n2064 585
R2333 gnd.n4355 gnd.n4354 585
R2334 gnd.n4354 gnd.n2073 585
R2335 gnd.n4356 gnd.n3388 585
R2336 gnd.n4660 gnd.n3388 585
R2337 gnd.n4358 gnd.n4357 585
R2338 gnd.n4357 gnd.n3386 585
R2339 gnd.n4359 gnd.n3399 585
R2340 gnd.n4389 gnd.n3399 585
R2341 gnd.n4362 gnd.n4361 585
R2342 gnd.n4361 gnd.n4360 585
R2343 gnd.n4363 gnd.n3406 585
R2344 gnd.n4378 gnd.n3406 585
R2345 gnd.n4365 gnd.n4364 585
R2346 gnd.n4366 gnd.n4365 585
R2347 gnd.n3416 gnd.n3415 585
R2348 gnd.n3423 gnd.n3415 585
R2349 gnd.n4341 gnd.n4340 585
R2350 gnd.n4340 gnd.n4339 585
R2351 gnd.n3419 gnd.n3418 585
R2352 gnd.n3433 gnd.n3419 585
R2353 gnd.n4267 gnd.n4266 585
R2354 gnd.n4266 gnd.n3432 585
R2355 gnd.n4268 gnd.n3442 585
R2356 gnd.n4317 gnd.n3442 585
R2357 gnd.n4270 gnd.n4269 585
R2358 gnd.n4269 gnd.n3440 585
R2359 gnd.n4271 gnd.n3453 585
R2360 gnd.n4300 gnd.n3453 585
R2361 gnd.n4273 gnd.n4272 585
R2362 gnd.n4272 gnd.n3461 585
R2363 gnd.n4274 gnd.n3460 585
R2364 gnd.n4289 gnd.n3460 585
R2365 gnd.n4276 gnd.n4275 585
R2366 gnd.n4277 gnd.n4276 585
R2367 gnd.n3472 gnd.n3471 585
R2368 gnd.n3471 gnd.n3468 585
R2369 gnd.n4256 gnd.n4255 585
R2370 gnd.n4255 gnd.n4254 585
R2371 gnd.n3475 gnd.n3474 585
R2372 gnd.n3488 gnd.n3475 585
R2373 gnd.n4180 gnd.n4179 585
R2374 gnd.n4179 gnd.n3487 585
R2375 gnd.n4181 gnd.n3497 585
R2376 gnd.n4232 gnd.n3497 585
R2377 gnd.n4183 gnd.n4182 585
R2378 gnd.n4182 gnd.n3495 585
R2379 gnd.n4184 gnd.n3508 585
R2380 gnd.n4215 gnd.n3508 585
R2381 gnd.n4186 gnd.n4185 585
R2382 gnd.n4185 gnd.n3515 585
R2383 gnd.n4187 gnd.n3514 585
R2384 gnd.n4204 gnd.n3514 585
R2385 gnd.n4189 gnd.n4188 585
R2386 gnd.n4192 gnd.n4189 585
R2387 gnd.n3525 gnd.n3524 585
R2388 gnd.n3524 gnd.n3522 585
R2389 gnd.n3632 gnd.n3631 585
R2390 gnd.n4147 gnd.n3631 585
R2391 gnd.n3634 gnd.n3633 585
R2392 gnd.n3635 gnd.n3634 585
R2393 gnd.n3645 gnd.n3621 585
R2394 gnd.n4153 gnd.n3621 585
R2395 gnd.n3647 gnd.n3646 585
R2396 gnd.n3648 gnd.n3647 585
R2397 gnd.n3644 gnd.n3643 585
R2398 gnd.n3644 gnd.n3611 585
R2399 gnd.n3642 gnd.n3609 585
R2400 gnd.n4161 gnd.n3609 585
R2401 gnd.n3598 gnd.n3596 585
R2402 gnd.n4123 gnd.n3598 585
R2403 gnd.n4169 gnd.n4168 585
R2404 gnd.n4168 gnd.n4167 585
R2405 gnd.n3597 gnd.n3595 585
R2406 gnd.n3662 gnd.n3597 585
R2407 gnd.n4094 gnd.n3661 585
R2408 gnd.n4113 gnd.n3661 585
R2409 gnd.n4096 gnd.n4095 585
R2410 gnd.n4097 gnd.n4096 585
R2411 gnd.n3671 gnd.n3670 585
R2412 gnd.n3677 gnd.n3670 585
R2413 gnd.n4089 gnd.n4088 585
R2414 gnd.n4088 gnd.n4087 585
R2415 gnd.n3674 gnd.n3673 585
R2416 gnd.n3685 gnd.n3674 585
R2417 gnd.n3974 gnd.n3693 585
R2418 gnd.n4066 gnd.n3693 585
R2419 gnd.n3976 gnd.n3975 585
R2420 gnd.n3975 gnd.n3691 585
R2421 gnd.n3977 gnd.n3704 585
R2422 gnd.n4056 gnd.n3704 585
R2423 gnd.n3979 gnd.n3978 585
R2424 gnd.n3979 gnd.n3711 585
R2425 gnd.n3981 gnd.n3980 585
R2426 gnd.n3980 gnd.n3710 585
R2427 gnd.n3982 gnd.n3721 585
R2428 gnd.n4036 gnd.n3721 585
R2429 gnd.n3984 gnd.n3983 585
R2430 gnd.n3983 gnd.n3719 585
R2431 gnd.n3985 gnd.n3730 585
R2432 gnd.n4025 gnd.n3730 585
R2433 gnd.n3987 gnd.n3986 585
R2434 gnd.n3987 gnd.n3736 585
R2435 gnd.n3989 gnd.n3988 585
R2436 gnd.n3988 gnd.n3735 585
R2437 gnd.n3990 gnd.n3751 585
R2438 gnd.n4004 gnd.n3751 585
R2439 gnd.n3991 gnd.n3804 585
R2440 gnd.n3804 gnd.n3743 585
R2441 gnd.n3993 gnd.n3992 585
R2442 gnd.n3994 gnd.n3993 585
R2443 gnd.n3805 gnd.n3803 585
R2444 gnd.n3803 gnd.n3802 585
R2445 gnd.n3958 gnd.n3957 585
R2446 gnd.n3957 gnd.n3956 585
R2447 gnd.n3808 gnd.n3807 585
R2448 gnd.n3809 gnd.n3808 585
R2449 gnd.n3947 gnd.n3946 585
R2450 gnd.n3948 gnd.n3947 585
R2451 gnd.n3817 gnd.n3816 585
R2452 gnd.n3816 gnd.n3815 585
R2453 gnd.n3942 gnd.n3941 585
R2454 gnd.n3941 gnd.n3940 585
R2455 gnd.n3820 gnd.n3819 585
R2456 gnd.n3931 gnd.n3820 585
R2457 gnd.n3930 gnd.n3929 585
R2458 gnd.n3932 gnd.n3930 585
R2459 gnd.n3828 gnd.n3827 585
R2460 gnd.n3827 gnd.n3826 585
R2461 gnd.n7681 gnd.n7680 585
R2462 gnd.n7680 gnd.n7679 585
R2463 gnd.n7682 gnd.n203 585
R2464 gnd.n208 gnd.n203 585
R2465 gnd.n7684 gnd.n7683 585
R2466 gnd.n7685 gnd.n7684 585
R2467 gnd.n190 gnd.n189 585
R2468 gnd.n193 gnd.n190 585
R2469 gnd.n7693 gnd.n7692 585
R2470 gnd.n7692 gnd.n7691 585
R2471 gnd.n7694 gnd.n185 585
R2472 gnd.n185 gnd.n184 585
R2473 gnd.n7696 gnd.n7695 585
R2474 gnd.n7697 gnd.n7696 585
R2475 gnd.n170 gnd.n169 585
R2476 gnd.n174 gnd.n170 585
R2477 gnd.n7705 gnd.n7704 585
R2478 gnd.n7704 gnd.n7703 585
R2479 gnd.n7706 gnd.n165 585
R2480 gnd.n7514 gnd.n165 585
R2481 gnd.n7708 gnd.n7707 585
R2482 gnd.n7709 gnd.n7708 585
R2483 gnd.n152 gnd.n151 585
R2484 gnd.n162 gnd.n152 585
R2485 gnd.n7717 gnd.n7716 585
R2486 gnd.n7716 gnd.n7715 585
R2487 gnd.n7718 gnd.n147 585
R2488 gnd.n147 gnd.n146 585
R2489 gnd.n7720 gnd.n7719 585
R2490 gnd.n7721 gnd.n7720 585
R2491 gnd.n132 gnd.n131 585
R2492 gnd.n136 gnd.n132 585
R2493 gnd.n7729 gnd.n7728 585
R2494 gnd.n7728 gnd.n7727 585
R2495 gnd.n7730 gnd.n127 585
R2496 gnd.n133 gnd.n127 585
R2497 gnd.n7732 gnd.n7731 585
R2498 gnd.n7733 gnd.n7732 585
R2499 gnd.n115 gnd.n114 585
R2500 gnd.n124 gnd.n115 585
R2501 gnd.n7741 gnd.n7740 585
R2502 gnd.n7740 gnd.n7739 585
R2503 gnd.n7742 gnd.n109 585
R2504 gnd.n109 gnd.n107 585
R2505 gnd.n7744 gnd.n7743 585
R2506 gnd.n7745 gnd.n7744 585
R2507 gnd.n110 gnd.n108 585
R2508 gnd.n7472 gnd.n108 585
R2509 gnd.n7433 gnd.n7432 585
R2510 gnd.n7432 gnd.n90 585
R2511 gnd.n7431 gnd.n91 585
R2512 gnd.n7753 gnd.n91 585
R2513 gnd.n7430 gnd.n7429 585
R2514 gnd.n7429 gnd.n7428 585
R2515 gnd.n363 gnd.n361 585
R2516 gnd.n364 gnd.n363 585
R2517 gnd.n7421 gnd.n7420 585
R2518 gnd.n7420 gnd.n7419 585
R2519 gnd.n369 gnd.n368 585
R2520 gnd.n370 gnd.n369 585
R2521 gnd.n7410 gnd.n7409 585
R2522 gnd.n7411 gnd.n7410 585
R2523 gnd.n379 gnd.n378 585
R2524 gnd.n7402 gnd.n378 585
R2525 gnd.n7373 gnd.n7372 585
R2526 gnd.n7372 gnd.n7371 585
R2527 gnd.n7374 gnd.n392 585
R2528 gnd.n7388 gnd.n392 585
R2529 gnd.n7375 gnd.n403 585
R2530 gnd.n7365 gnd.n403 585
R2531 gnd.n7377 gnd.n7376 585
R2532 gnd.n7378 gnd.n7377 585
R2533 gnd.n404 gnd.n402 585
R2534 gnd.n7353 gnd.n402 585
R2535 gnd.n7329 gnd.n7328 585
R2536 gnd.n7328 gnd.n7327 585
R2537 gnd.n7330 gnd.n424 585
R2538 gnd.n7344 gnd.n424 585
R2539 gnd.n7331 gnd.n436 585
R2540 gnd.n7319 gnd.n436 585
R2541 gnd.n7333 gnd.n7332 585
R2542 gnd.n7334 gnd.n7333 585
R2543 gnd.n437 gnd.n435 585
R2544 gnd.n7306 gnd.n435 585
R2545 gnd.n7282 gnd.n7281 585
R2546 gnd.n7281 gnd.n449 585
R2547 gnd.n7283 gnd.n459 585
R2548 gnd.n7297 gnd.n459 585
R2549 gnd.n7284 gnd.n471 585
R2550 gnd.n7273 gnd.n471 585
R2551 gnd.n7286 gnd.n7285 585
R2552 gnd.n7287 gnd.n7286 585
R2553 gnd.n472 gnd.n470 585
R2554 gnd.n7260 gnd.n470 585
R2555 gnd.n7236 gnd.n7235 585
R2556 gnd.n7235 gnd.n483 585
R2557 gnd.n7237 gnd.n494 585
R2558 gnd.n7251 gnd.n494 585
R2559 gnd.n7238 gnd.n506 585
R2560 gnd.n7227 gnd.n506 585
R2561 gnd.n7240 gnd.n7239 585
R2562 gnd.n7241 gnd.n7240 585
R2563 gnd.n507 gnd.n505 585
R2564 gnd.n7223 gnd.n505 585
R2565 gnd.n7096 gnd.n7095 585
R2566 gnd.n7097 gnd.n7096 585
R2567 gnd.n7091 gnd.n523 585
R2568 gnd.n7214 gnd.n523 585
R2569 gnd.n606 gnd.n605 585
R2570 gnd.n7163 gnd.n607 585
R2571 gnd.n7162 gnd.n608 585
R2572 gnd.n615 gnd.n609 585
R2573 gnd.n7155 gnd.n616 585
R2574 gnd.n7154 gnd.n617 585
R2575 gnd.n619 gnd.n618 585
R2576 gnd.n7147 gnd.n625 585
R2577 gnd.n7146 gnd.n626 585
R2578 gnd.n633 gnd.n627 585
R2579 gnd.n7139 gnd.n634 585
R2580 gnd.n7138 gnd.n635 585
R2581 gnd.n637 gnd.n636 585
R2582 gnd.n7131 gnd.n643 585
R2583 gnd.n7130 gnd.n644 585
R2584 gnd.n568 gnd.n567 585
R2585 gnd.n7201 gnd.n7200 585
R2586 gnd.n571 gnd.n566 585
R2587 gnd.n7193 gnd.n519 585
R2588 gnd.n7203 gnd.n519 585
R2589 gnd.n348 gnd.n347 585
R2590 gnd.n7535 gnd.n343 585
R2591 gnd.n7537 gnd.n7536 585
R2592 gnd.n7539 gnd.n341 585
R2593 gnd.n7541 gnd.n7540 585
R2594 gnd.n7542 gnd.n336 585
R2595 gnd.n7544 gnd.n7543 585
R2596 gnd.n7546 gnd.n334 585
R2597 gnd.n7548 gnd.n7547 585
R2598 gnd.n7549 gnd.n329 585
R2599 gnd.n7551 gnd.n7550 585
R2600 gnd.n7553 gnd.n327 585
R2601 gnd.n7555 gnd.n7554 585
R2602 gnd.n7556 gnd.n322 585
R2603 gnd.n7558 gnd.n7557 585
R2604 gnd.n7560 gnd.n320 585
R2605 gnd.n7562 gnd.n7561 585
R2606 gnd.n7563 gnd.n318 585
R2607 gnd.n7564 gnd.n207 585
R2608 gnd.n211 gnd.n207 585
R2609 gnd.n7531 gnd.n210 585
R2610 gnd.n7679 gnd.n210 585
R2611 gnd.n7530 gnd.n7529 585
R2612 gnd.n7529 gnd.n208 585
R2613 gnd.n7528 gnd.n202 585
R2614 gnd.n7685 gnd.n202 585
R2615 gnd.n353 gnd.n352 585
R2616 gnd.n352 gnd.n193 585
R2617 gnd.n7524 gnd.n192 585
R2618 gnd.n7691 gnd.n192 585
R2619 gnd.n7523 gnd.n7522 585
R2620 gnd.n7522 gnd.n184 585
R2621 gnd.n7521 gnd.n183 585
R2622 gnd.n7697 gnd.n183 585
R2623 gnd.n356 gnd.n355 585
R2624 gnd.n355 gnd.n174 585
R2625 gnd.n7517 gnd.n173 585
R2626 gnd.n7703 gnd.n173 585
R2627 gnd.n7516 gnd.n7515 585
R2628 gnd.n7515 gnd.n7514 585
R2629 gnd.n358 gnd.n164 585
R2630 gnd.n7709 gnd.n164 585
R2631 gnd.n7453 gnd.n7452 585
R2632 gnd.n7452 gnd.n162 585
R2633 gnd.n7454 gnd.n154 585
R2634 gnd.n7715 gnd.n154 585
R2635 gnd.n7456 gnd.n7455 585
R2636 gnd.n7455 gnd.n146 585
R2637 gnd.n7457 gnd.n145 585
R2638 gnd.n7721 gnd.n145 585
R2639 gnd.n7459 gnd.n7458 585
R2640 gnd.n7458 gnd.n136 585
R2641 gnd.n7460 gnd.n135 585
R2642 gnd.n7727 gnd.n135 585
R2643 gnd.n7462 gnd.n7461 585
R2644 gnd.n7461 gnd.n133 585
R2645 gnd.n7463 gnd.n126 585
R2646 gnd.n7733 gnd.n126 585
R2647 gnd.n7465 gnd.n7464 585
R2648 gnd.n7464 gnd.n124 585
R2649 gnd.n7466 gnd.n117 585
R2650 gnd.n7739 gnd.n117 585
R2651 gnd.n7468 gnd.n7467 585
R2652 gnd.n7467 gnd.n107 585
R2653 gnd.n7469 gnd.n106 585
R2654 gnd.n7745 gnd.n106 585
R2655 gnd.n7471 gnd.n7470 585
R2656 gnd.n7472 gnd.n7471 585
R2657 gnd.n88 gnd.n87 585
R2658 gnd.n90 gnd.n88 585
R2659 gnd.n7755 gnd.n7754 585
R2660 gnd.n7754 gnd.n7753 585
R2661 gnd.n7756 gnd.n86 585
R2662 gnd.n7428 gnd.n86 585
R2663 gnd.n372 gnd.n85 585
R2664 gnd.n372 gnd.n364 585
R2665 gnd.n7395 gnd.n373 585
R2666 gnd.n7419 gnd.n373 585
R2667 gnd.n7396 gnd.n7394 585
R2668 gnd.n7394 gnd.n370 585
R2669 gnd.n386 gnd.n377 585
R2670 gnd.n7411 gnd.n377 585
R2671 gnd.n7401 gnd.n7400 585
R2672 gnd.n7402 gnd.n7401 585
R2673 gnd.n385 gnd.n384 585
R2674 gnd.n7371 gnd.n384 585
R2675 gnd.n7390 gnd.n7389 585
R2676 gnd.n7389 gnd.n7388 585
R2677 gnd.n389 gnd.n388 585
R2678 gnd.n7365 gnd.n389 585
R2679 gnd.n418 gnd.n400 585
R2680 gnd.n7378 gnd.n400 585
R2681 gnd.n7352 gnd.n7351 585
R2682 gnd.n7353 gnd.n7352 585
R2683 gnd.n417 gnd.n416 585
R2684 gnd.n7327 gnd.n416 585
R2685 gnd.n7346 gnd.n7345 585
R2686 gnd.n7345 gnd.n7344 585
R2687 gnd.n421 gnd.n420 585
R2688 gnd.n7319 gnd.n421 585
R2689 gnd.n453 gnd.n433 585
R2690 gnd.n7334 gnd.n433 585
R2691 gnd.n7305 gnd.n7304 585
R2692 gnd.n7306 gnd.n7305 585
R2693 gnd.n452 gnd.n451 585
R2694 gnd.n451 gnd.n449 585
R2695 gnd.n7299 gnd.n7298 585
R2696 gnd.n7298 gnd.n7297 585
R2697 gnd.n456 gnd.n455 585
R2698 gnd.n7273 gnd.n456 585
R2699 gnd.n487 gnd.n468 585
R2700 gnd.n7287 gnd.n468 585
R2701 gnd.n7259 gnd.n7258 585
R2702 gnd.n7260 gnd.n7259 585
R2703 gnd.n486 gnd.n485 585
R2704 gnd.n485 gnd.n483 585
R2705 gnd.n7253 gnd.n7252 585
R2706 gnd.n7252 gnd.n7251 585
R2707 gnd.n490 gnd.n489 585
R2708 gnd.n7227 gnd.n490 585
R2709 gnd.n517 gnd.n503 585
R2710 gnd.n7241 gnd.n503 585
R2711 gnd.n7222 gnd.n7221 585
R2712 gnd.n7223 gnd.n7222 585
R2713 gnd.n516 gnd.n515 585
R2714 gnd.n7097 gnd.n515 585
R2715 gnd.n7216 gnd.n7215 585
R2716 gnd.n7215 gnd.n7214 585
R2717 gnd.n4669 gnd.n2015 585
R2718 gnd.n2015 gnd.n1992 585
R2719 gnd.n4670 gnd.n3381 585
R2720 gnd.n3381 gnd.n2066 585
R2721 gnd.n4672 gnd.n4671 585
R2722 gnd.n4673 gnd.n4672 585
R2723 gnd.n3382 gnd.n3380 585
R2724 gnd.n3389 gnd.n3380 585
R2725 gnd.n4663 gnd.n4662 585
R2726 gnd.n4662 gnd.n4661 585
R2727 gnd.n3385 gnd.n3384 585
R2728 gnd.n4388 gnd.n3385 585
R2729 gnd.n4374 gnd.n3408 585
R2730 gnd.n3408 gnd.n3398 585
R2731 gnd.n4376 gnd.n4375 585
R2732 gnd.n4377 gnd.n4376 585
R2733 gnd.n3409 gnd.n3407 585
R2734 gnd.n3407 gnd.n3405 585
R2735 gnd.n4369 gnd.n4368 585
R2736 gnd.n4368 gnd.n4367 585
R2737 gnd.n3412 gnd.n3411 585
R2738 gnd.n3421 gnd.n3412 585
R2739 gnd.n4325 gnd.n3435 585
R2740 gnd.n3435 gnd.n3420 585
R2741 gnd.n4327 gnd.n4326 585
R2742 gnd.n4328 gnd.n4327 585
R2743 gnd.n3436 gnd.n3434 585
R2744 gnd.n3443 gnd.n3434 585
R2745 gnd.n4320 gnd.n4319 585
R2746 gnd.n4319 gnd.n4318 585
R2747 gnd.n3439 gnd.n3438 585
R2748 gnd.n4299 gnd.n3439 585
R2749 gnd.n4285 gnd.n3463 585
R2750 gnd.n3463 gnd.n3452 585
R2751 gnd.n4287 gnd.n4286 585
R2752 gnd.n4288 gnd.n4287 585
R2753 gnd.n3464 gnd.n3462 585
R2754 gnd.n3462 gnd.n3459 585
R2755 gnd.n4280 gnd.n4279 585
R2756 gnd.n4279 gnd.n4278 585
R2757 gnd.n3467 gnd.n3466 585
R2758 gnd.n3477 gnd.n3467 585
R2759 gnd.n4240 gnd.n3490 585
R2760 gnd.n3490 gnd.n3476 585
R2761 gnd.n4242 gnd.n4241 585
R2762 gnd.n4243 gnd.n4242 585
R2763 gnd.n3491 gnd.n3489 585
R2764 gnd.n3498 gnd.n3489 585
R2765 gnd.n4235 gnd.n4234 585
R2766 gnd.n4234 gnd.n4233 585
R2767 gnd.n3494 gnd.n3493 585
R2768 gnd.n4214 gnd.n3494 585
R2769 gnd.n4200 gnd.n3517 585
R2770 gnd.n3517 gnd.n3507 585
R2771 gnd.n4202 gnd.n4201 585
R2772 gnd.n4203 gnd.n4202 585
R2773 gnd.n3518 gnd.n3516 585
R2774 gnd.n4191 gnd.n3516 585
R2775 gnd.n4195 gnd.n4194 585
R2776 gnd.n4194 gnd.n4193 585
R2777 gnd.n3521 gnd.n3520 585
R2778 gnd.n4146 gnd.n3521 585
R2779 gnd.n3639 gnd.n3638 585
R2780 gnd.n3640 gnd.n3639 585
R2781 gnd.n3619 gnd.n3618 585
R2782 gnd.n3622 gnd.n3619 585
R2783 gnd.n4156 gnd.n4155 585
R2784 gnd.n4155 gnd.n4154 585
R2785 gnd.n4157 gnd.n3613 585
R2786 gnd.n3649 gnd.n3613 585
R2787 gnd.n4159 gnd.n4158 585
R2788 gnd.n4160 gnd.n4159 585
R2789 gnd.n3614 gnd.n3612 585
R2790 gnd.n4124 gnd.n3612 585
R2791 gnd.n4108 gnd.n4107 585
R2792 gnd.n4107 gnd.n3600 585
R2793 gnd.n4109 gnd.n3664 585
R2794 gnd.n3664 gnd.n3599 585
R2795 gnd.n4111 gnd.n4110 585
R2796 gnd.n4112 gnd.n4111 585
R2797 gnd.n3665 gnd.n3663 585
R2798 gnd.n3663 gnd.n3660 585
R2799 gnd.n4100 gnd.n4099 585
R2800 gnd.n4099 gnd.n4098 585
R2801 gnd.n3668 gnd.n3667 585
R2802 gnd.n3675 gnd.n3668 585
R2803 gnd.n4074 gnd.n4073 585
R2804 gnd.n4075 gnd.n4074 585
R2805 gnd.n3687 gnd.n3686 585
R2806 gnd.n3694 gnd.n3686 585
R2807 gnd.n4069 gnd.n4068 585
R2808 gnd.n4068 gnd.n4067 585
R2809 gnd.n3690 gnd.n3689 585
R2810 gnd.n4057 gnd.n3690 585
R2811 gnd.n4044 gnd.n3714 585
R2812 gnd.n3714 gnd.n3713 585
R2813 gnd.n4046 gnd.n4045 585
R2814 gnd.n4047 gnd.n4046 585
R2815 gnd.n3715 gnd.n3712 585
R2816 gnd.n3722 gnd.n3712 585
R2817 gnd.n4039 gnd.n4038 585
R2818 gnd.n4038 gnd.n4037 585
R2819 gnd.n3718 gnd.n3717 585
R2820 gnd.n4026 gnd.n3718 585
R2821 gnd.n4013 gnd.n3739 585
R2822 gnd.n3739 gnd.n3738 585
R2823 gnd.n4015 gnd.n4014 585
R2824 gnd.n4016 gnd.n4015 585
R2825 gnd.n4009 gnd.n3737 585
R2826 gnd.n4008 gnd.n4007 585
R2827 gnd.n3742 gnd.n3741 585
R2828 gnd.n4005 gnd.n3742 585
R2829 gnd.n3764 gnd.n3763 585
R2830 gnd.n3767 gnd.n3766 585
R2831 gnd.n3765 gnd.n3760 585
R2832 gnd.n3772 gnd.n3771 585
R2833 gnd.n3774 gnd.n3773 585
R2834 gnd.n3777 gnd.n3776 585
R2835 gnd.n3775 gnd.n3758 585
R2836 gnd.n3782 gnd.n3781 585
R2837 gnd.n3784 gnd.n3783 585
R2838 gnd.n3787 gnd.n3786 585
R2839 gnd.n3785 gnd.n3756 585
R2840 gnd.n3792 gnd.n3791 585
R2841 gnd.n3796 gnd.n3793 585
R2842 gnd.n3797 gnd.n3734 585
R2843 gnd.n4675 gnd.n2030 585
R2844 gnd.n4742 gnd.n4741 585
R2845 gnd.n4744 gnd.n4743 585
R2846 gnd.n4746 gnd.n4745 585
R2847 gnd.n4748 gnd.n4747 585
R2848 gnd.n4750 gnd.n4749 585
R2849 gnd.n4752 gnd.n4751 585
R2850 gnd.n4754 gnd.n4753 585
R2851 gnd.n4756 gnd.n4755 585
R2852 gnd.n4758 gnd.n4757 585
R2853 gnd.n4760 gnd.n4759 585
R2854 gnd.n4762 gnd.n4761 585
R2855 gnd.n4764 gnd.n4763 585
R2856 gnd.n4767 gnd.n4766 585
R2857 gnd.n4765 gnd.n2018 585
R2858 gnd.n4771 gnd.n2016 585
R2859 gnd.n4773 gnd.n4772 585
R2860 gnd.n4774 gnd.n4773 585
R2861 gnd.n4676 gnd.n2071 585
R2862 gnd.n4676 gnd.n1992 585
R2863 gnd.n4678 gnd.n4677 585
R2864 gnd.n4677 gnd.n2066 585
R2865 gnd.n4674 gnd.n2070 585
R2866 gnd.n4674 gnd.n4673 585
R2867 gnd.n4653 gnd.n2072 585
R2868 gnd.n3389 gnd.n2072 585
R2869 gnd.n4652 gnd.n3387 585
R2870 gnd.n4661 gnd.n3387 585
R2871 gnd.n4387 gnd.n3394 585
R2872 gnd.n4388 gnd.n4387 585
R2873 gnd.n4386 gnd.n4385 585
R2874 gnd.n4386 gnd.n3398 585
R2875 gnd.n4384 gnd.n3400 585
R2876 gnd.n4377 gnd.n3400 585
R2877 gnd.n3413 gnd.n3401 585
R2878 gnd.n3413 gnd.n3405 585
R2879 gnd.n4333 gnd.n3414 585
R2880 gnd.n4367 gnd.n3414 585
R2881 gnd.n4332 gnd.n4331 585
R2882 gnd.n4331 gnd.n3421 585
R2883 gnd.n4330 gnd.n3429 585
R2884 gnd.n4330 gnd.n3420 585
R2885 gnd.n4329 gnd.n3431 585
R2886 gnd.n4329 gnd.n4328 585
R2887 gnd.n4308 gnd.n3430 585
R2888 gnd.n3443 gnd.n3430 585
R2889 gnd.n4307 gnd.n3441 585
R2890 gnd.n4318 gnd.n3441 585
R2891 gnd.n4298 gnd.n3448 585
R2892 gnd.n4299 gnd.n4298 585
R2893 gnd.n4297 gnd.n4296 585
R2894 gnd.n4297 gnd.n3452 585
R2895 gnd.n4295 gnd.n3454 585
R2896 gnd.n4288 gnd.n3454 585
R2897 gnd.n3469 gnd.n3455 585
R2898 gnd.n3469 gnd.n3459 585
R2899 gnd.n4248 gnd.n3470 585
R2900 gnd.n4278 gnd.n3470 585
R2901 gnd.n4247 gnd.n4246 585
R2902 gnd.n4246 gnd.n3477 585
R2903 gnd.n4245 gnd.n3484 585
R2904 gnd.n4245 gnd.n3476 585
R2905 gnd.n4244 gnd.n3486 585
R2906 gnd.n4244 gnd.n4243 585
R2907 gnd.n4223 gnd.n3485 585
R2908 gnd.n3498 gnd.n3485 585
R2909 gnd.n4222 gnd.n3496 585
R2910 gnd.n4233 gnd.n3496 585
R2911 gnd.n4213 gnd.n3503 585
R2912 gnd.n4214 gnd.n4213 585
R2913 gnd.n4212 gnd.n4211 585
R2914 gnd.n4212 gnd.n3507 585
R2915 gnd.n4210 gnd.n3509 585
R2916 gnd.n4203 gnd.n3509 585
R2917 gnd.n4190 gnd.n3510 585
R2918 gnd.n4191 gnd.n4190 585
R2919 gnd.n4143 gnd.n3523 585
R2920 gnd.n4193 gnd.n3523 585
R2921 gnd.n4145 gnd.n4144 585
R2922 gnd.n4146 gnd.n4145 585
R2923 gnd.n4138 gnd.n3641 585
R2924 gnd.n3641 gnd.n3640 585
R2925 gnd.n4136 gnd.n4135 585
R2926 gnd.n4135 gnd.n3622 585
R2927 gnd.n4133 gnd.n3620 585
R2928 gnd.n4154 gnd.n3620 585
R2929 gnd.n3651 gnd.n3650 585
R2930 gnd.n3650 gnd.n3649 585
R2931 gnd.n4127 gnd.n3610 585
R2932 gnd.n4160 gnd.n3610 585
R2933 gnd.n4126 gnd.n4125 585
R2934 gnd.n4125 gnd.n4124 585
R2935 gnd.n4122 gnd.n3653 585
R2936 gnd.n4122 gnd.n3600 585
R2937 gnd.n4121 gnd.n4120 585
R2938 gnd.n4121 gnd.n3599 585
R2939 gnd.n3656 gnd.n3655 585
R2940 gnd.n4112 gnd.n3655 585
R2941 gnd.n4080 gnd.n4079 585
R2942 gnd.n4079 gnd.n3660 585
R2943 gnd.n4081 gnd.n3669 585
R2944 gnd.n4098 gnd.n3669 585
R2945 gnd.n4078 gnd.n4077 585
R2946 gnd.n4077 gnd.n3675 585
R2947 gnd.n4076 gnd.n3683 585
R2948 gnd.n4076 gnd.n4075 585
R2949 gnd.n4061 gnd.n3684 585
R2950 gnd.n3694 gnd.n3684 585
R2951 gnd.n4060 gnd.n3692 585
R2952 gnd.n4067 gnd.n3692 585
R2953 gnd.n4059 gnd.n4058 585
R2954 gnd.n4058 gnd.n4057 585
R2955 gnd.n3703 gnd.n3700 585
R2956 gnd.n3713 gnd.n3703 585
R2957 gnd.n4049 gnd.n4048 585
R2958 gnd.n4048 gnd.n4047 585
R2959 gnd.n3709 gnd.n3708 585
R2960 gnd.n3722 gnd.n3709 585
R2961 gnd.n4029 gnd.n3720 585
R2962 gnd.n4037 gnd.n3720 585
R2963 gnd.n4028 gnd.n4027 585
R2964 gnd.n4027 gnd.n4026 585
R2965 gnd.n3729 gnd.n3727 585
R2966 gnd.n3738 gnd.n3729 585
R2967 gnd.n4018 gnd.n4017 585
R2968 gnd.n4017 gnd.n4016 585
R2969 gnd.n7000 gnd.n739 585
R2970 gnd.n6879 gnd.n739 585
R2971 gnd.n7002 gnd.n7001 585
R2972 gnd.n7003 gnd.n7002 585
R2973 gnd.n740 gnd.n738 585
R2974 gnd.n738 gnd.n734 585
R2975 gnd.n6870 gnd.n6869 585
R2976 gnd.n6871 gnd.n6870 585
R2977 gnd.n6868 gnd.n989 585
R2978 gnd.n6835 gnd.n989 585
R2979 gnd.n6867 gnd.n6866 585
R2980 gnd.n6866 gnd.n6865 585
R2981 gnd.n991 gnd.n990 585
R2982 gnd.n6786 gnd.n991 585
R2983 gnd.n6818 gnd.n6817 585
R2984 gnd.n6817 gnd.n1001 585
R2985 gnd.n6819 gnd.n1017 585
R2986 gnd.n1017 gnd.n999 585
R2987 gnd.n6821 gnd.n6820 585
R2988 gnd.n6822 gnd.n6821 585
R2989 gnd.n6816 gnd.n1016 585
R2990 gnd.n6794 gnd.n1016 585
R2991 gnd.n6815 gnd.n6814 585
R2992 gnd.n6814 gnd.n6813 585
R2993 gnd.n1019 gnd.n1018 585
R2994 gnd.n6776 gnd.n1019 585
R2995 gnd.n6762 gnd.n6761 585
R2996 gnd.n6762 gnd.n1029 585
R2997 gnd.n6764 gnd.n6763 585
R2998 gnd.n6763 gnd.n1027 585
R2999 gnd.n6765 gnd.n1041 585
R3000 gnd.n6656 gnd.n1041 585
R3001 gnd.n6767 gnd.n6766 585
R3002 gnd.n6768 gnd.n6767 585
R3003 gnd.n6760 gnd.n1040 585
R3004 gnd.n1047 gnd.n1040 585
R3005 gnd.n6759 gnd.n6758 585
R3006 gnd.n6758 gnd.n6757 585
R3007 gnd.n1043 gnd.n1042 585
R3008 gnd.n6673 gnd.n1043 585
R3009 gnd.n6745 gnd.n6744 585
R3010 gnd.n6746 gnd.n6745 585
R3011 gnd.n6743 gnd.n1059 585
R3012 gnd.n1059 gnd.n1055 585
R3013 gnd.n6742 gnd.n6741 585
R3014 gnd.n6741 gnd.n6740 585
R3015 gnd.n1061 gnd.n1060 585
R3016 gnd.n6680 gnd.n1061 585
R3017 gnd.n6719 gnd.n6718 585
R3018 gnd.n6720 gnd.n6719 585
R3019 gnd.n6717 gnd.n1072 585
R3020 gnd.n6712 gnd.n1072 585
R3021 gnd.n6716 gnd.n6715 585
R3022 gnd.n6715 gnd.n6714 585
R3023 gnd.n1074 gnd.n1073 585
R3024 gnd.n1087 gnd.n1074 585
R3025 gnd.n6636 gnd.n1109 585
R3026 gnd.n1109 gnd.n1085 585
R3027 gnd.n6638 gnd.n6637 585
R3028 gnd.n6639 gnd.n6638 585
R3029 gnd.n6635 gnd.n1094 585
R3030 gnd.n6693 gnd.n1094 585
R3031 gnd.n6634 gnd.n6633 585
R3032 gnd.n6633 gnd.n6632 585
R3033 gnd.n1111 gnd.n1110 585
R3034 gnd.n6630 gnd.n1111 585
R3035 gnd.n6621 gnd.n1119 585
R3036 gnd.n6609 gnd.n1119 585
R3037 gnd.n6623 gnd.n6622 585
R3038 gnd.n6624 gnd.n6623 585
R3039 gnd.n6620 gnd.n1118 585
R3040 gnd.n1124 gnd.n1118 585
R3041 gnd.n6619 gnd.n6618 585
R3042 gnd.n6618 gnd.n6617 585
R3043 gnd.n1121 gnd.n1120 585
R3044 gnd.n6569 gnd.n1121 585
R3045 gnd.n6572 gnd.n1147 585
R3046 gnd.n6572 gnd.n6571 585
R3047 gnd.n6574 gnd.n6573 585
R3048 gnd.n6573 gnd.n1132 585
R3049 gnd.n6575 gnd.n1145 585
R3050 gnd.n6561 gnd.n1145 585
R3051 gnd.n6577 gnd.n6576 585
R3052 gnd.n6578 gnd.n6577 585
R3053 gnd.n1146 gnd.n1144 585
R3054 gnd.n6537 gnd.n1144 585
R3055 gnd.n6527 gnd.n1162 585
R3056 gnd.n1162 gnd.n1156 585
R3057 gnd.n6529 gnd.n6528 585
R3058 gnd.n6530 gnd.n6529 585
R3059 gnd.n6526 gnd.n1161 585
R3060 gnd.n1168 gnd.n1161 585
R3061 gnd.n6525 gnd.n6524 585
R3062 gnd.n6524 gnd.n6523 585
R3063 gnd.n1164 gnd.n1163 585
R3064 gnd.n6322 gnd.n1164 585
R3065 gnd.n6511 gnd.n6510 585
R3066 gnd.n6512 gnd.n6511 585
R3067 gnd.n6509 gnd.n1179 585
R3068 gnd.n1179 gnd.n1176 585
R3069 gnd.n6508 gnd.n6507 585
R3070 gnd.n6507 gnd.n6506 585
R3071 gnd.n1181 gnd.n1180 585
R3072 gnd.n6465 gnd.n1181 585
R3073 gnd.n6478 gnd.n6477 585
R3074 gnd.n6479 gnd.n6478 585
R3075 gnd.n6476 gnd.n1193 585
R3076 gnd.n6471 gnd.n1193 585
R3077 gnd.n6475 gnd.n6474 585
R3078 gnd.n6474 gnd.n6473 585
R3079 gnd.n1195 gnd.n1194 585
R3080 gnd.n6454 gnd.n1195 585
R3081 gnd.n6441 gnd.n1219 585
R3082 gnd.n1219 gnd.n1206 585
R3083 gnd.n6443 gnd.n6442 585
R3084 gnd.n6444 gnd.n6443 585
R3085 gnd.n6440 gnd.n1218 585
R3086 gnd.n1218 gnd.n1214 585
R3087 gnd.n6439 gnd.n6438 585
R3088 gnd.n6438 gnd.n6437 585
R3089 gnd.n1221 gnd.n1220 585
R3090 gnd.n6345 gnd.n1221 585
R3091 gnd.n6425 gnd.n6424 585
R3092 gnd.n6426 gnd.n6425 585
R3093 gnd.n6423 gnd.n1235 585
R3094 gnd.n1235 gnd.n1231 585
R3095 gnd.n6422 gnd.n6421 585
R3096 gnd.n6421 gnd.n6420 585
R3097 gnd.n1237 gnd.n1236 585
R3098 gnd.n6353 gnd.n1237 585
R3099 gnd.n6407 gnd.n6406 585
R3100 gnd.n6408 gnd.n6407 585
R3101 gnd.n6405 gnd.n1248 585
R3102 gnd.n1254 gnd.n1248 585
R3103 gnd.n6404 gnd.n6403 585
R3104 gnd.n6403 gnd.n6402 585
R3105 gnd.n1250 gnd.n1249 585
R3106 gnd.n1264 gnd.n1250 585
R3107 gnd.n6377 gnd.n6376 585
R3108 gnd.n6376 gnd.n1262 585
R3109 gnd.n6378 gnd.n1274 585
R3110 gnd.n6364 gnd.n1274 585
R3111 gnd.n6380 gnd.n6379 585
R3112 gnd.n6381 gnd.n6380 585
R3113 gnd.n6375 gnd.n1273 585
R3114 gnd.n6370 gnd.n1273 585
R3115 gnd.n6374 gnd.n6373 585
R3116 gnd.n6373 gnd.n6372 585
R3117 gnd.n1276 gnd.n1275 585
R3118 gnd.n1323 gnd.n1276 585
R3119 gnd.n6258 gnd.n6257 585
R3120 gnd.n6259 gnd.n6258 585
R3121 gnd.n1315 gnd.n1314 585
R3122 gnd.n1315 gnd.n1300 585
R3123 gnd.n6267 gnd.n6266 585
R3124 gnd.n6266 gnd.n6265 585
R3125 gnd.n6268 gnd.n1312 585
R3126 gnd.n6245 gnd.n1312 585
R3127 gnd.n6270 gnd.n6269 585
R3128 gnd.n6271 gnd.n6270 585
R3129 gnd.n1313 gnd.n1311 585
R3130 gnd.n1311 gnd.n1308 585
R3131 gnd.n6219 gnd.n1348 585
R3132 gnd.n6219 gnd.n6218 585
R3133 gnd.n6220 gnd.n1347 585
R3134 gnd.n6220 gnd.n1335 585
R3135 gnd.n6222 gnd.n6221 585
R3136 gnd.n6221 gnd.n1333 585
R3137 gnd.n6223 gnd.n1345 585
R3138 gnd.n6207 gnd.n1345 585
R3139 gnd.n6225 gnd.n6224 585
R3140 gnd.n6226 gnd.n6225 585
R3141 gnd.n1346 gnd.n1344 585
R3142 gnd.n6194 gnd.n1344 585
R3143 gnd.n6168 gnd.n6166 585
R3144 gnd.n6168 gnd.n6167 585
R3145 gnd.n6169 gnd.n6165 585
R3146 gnd.n6169 gnd.n1366 585
R3147 gnd.n6171 gnd.n6170 585
R3148 gnd.n6170 gnd.n1364 585
R3149 gnd.n6172 gnd.n1376 585
R3150 gnd.n6153 gnd.n1376 585
R3151 gnd.n6174 gnd.n6173 585
R3152 gnd.n6175 gnd.n6174 585
R3153 gnd.n6164 gnd.n1375 585
R3154 gnd.n6159 gnd.n1375 585
R3155 gnd.n6163 gnd.n6162 585
R3156 gnd.n6162 gnd.n6161 585
R3157 gnd.n1378 gnd.n1377 585
R3158 gnd.n1393 gnd.n1378 585
R3159 gnd.n6106 gnd.n1414 585
R3160 gnd.n6106 gnd.n6105 585
R3161 gnd.n6107 gnd.n1413 585
R3162 gnd.n6107 gnd.n1401 585
R3163 gnd.n6109 gnd.n6108 585
R3164 gnd.n6108 gnd.n1399 585
R3165 gnd.n6110 gnd.n1411 585
R3166 gnd.n6096 gnd.n1411 585
R3167 gnd.n6112 gnd.n6111 585
R3168 gnd.n6113 gnd.n6112 585
R3169 gnd.n1412 gnd.n1410 585
R3170 gnd.n6090 gnd.n1410 585
R3171 gnd.n6049 gnd.n6048 585
R3172 gnd.n6048 gnd.n6047 585
R3173 gnd.n6051 gnd.n6050 585
R3174 gnd.n6051 gnd.n1429 585
R3175 gnd.n6052 gnd.n1446 585
R3176 gnd.n6052 gnd.n1427 585
R3177 gnd.n6056 gnd.n6055 585
R3178 gnd.n6055 gnd.n6054 585
R3179 gnd.n6057 gnd.n1435 585
R3180 gnd.n6072 gnd.n1435 585
R3181 gnd.n6058 gnd.n1444 585
R3182 gnd.n1452 gnd.n1444 585
R3183 gnd.n6060 gnd.n6059 585
R3184 gnd.n6061 gnd.n6060 585
R3185 gnd.n1445 gnd.n1443 585
R3186 gnd.n6021 gnd.n1443 585
R3187 gnd.n6007 gnd.n1470 585
R3188 gnd.n1470 gnd.n1458 585
R3189 gnd.n6009 gnd.n6008 585
R3190 gnd.n6010 gnd.n6009 585
R3191 gnd.n6005 gnd.n1469 585
R3192 gnd.n6004 gnd.n6003 585
R3193 gnd.n1492 gnd.n1491 585
R3194 gnd.n6001 gnd.n1492 585
R3195 gnd.n1532 gnd.n1531 585
R3196 gnd.n1534 gnd.n1533 585
R3197 gnd.n1536 gnd.n1535 585
R3198 gnd.n1538 gnd.n1537 585
R3199 gnd.n1540 gnd.n1539 585
R3200 gnd.n1542 gnd.n1541 585
R3201 gnd.n1544 gnd.n1543 585
R3202 gnd.n1546 gnd.n1545 585
R3203 gnd.n1548 gnd.n1547 585
R3204 gnd.n1550 gnd.n1549 585
R3205 gnd.n1552 gnd.n1551 585
R3206 gnd.n1554 gnd.n1553 585
R3207 gnd.n1556 gnd.n1555 585
R3208 gnd.n1558 gnd.n1557 585
R3209 gnd.n1560 gnd.n1559 585
R3210 gnd.n1562 gnd.n1561 585
R3211 gnd.n1564 gnd.n1563 585
R3212 gnd.n1566 gnd.n1565 585
R3213 gnd.n1568 gnd.n1567 585
R3214 gnd.n1570 gnd.n1569 585
R3215 gnd.n1572 gnd.n1571 585
R3216 gnd.n1574 gnd.n1573 585
R3217 gnd.n1576 gnd.n1575 585
R3218 gnd.n1578 gnd.n1577 585
R3219 gnd.n1580 gnd.n1579 585
R3220 gnd.n1582 gnd.n1581 585
R3221 gnd.n1584 gnd.n1583 585
R3222 gnd.n1586 gnd.n1585 585
R3223 gnd.n1588 gnd.n1587 585
R3224 gnd.n5932 gnd.n5931 585
R3225 gnd.n5934 gnd.n5933 585
R3226 gnd.n5936 gnd.n5935 585
R3227 gnd.n5938 gnd.n5937 585
R3228 gnd.n5941 gnd.n5940 585
R3229 gnd.n5943 gnd.n5942 585
R3230 gnd.n5945 gnd.n5944 585
R3231 gnd.n5947 gnd.n5946 585
R3232 gnd.n5949 gnd.n5948 585
R3233 gnd.n5951 gnd.n5950 585
R3234 gnd.n5953 gnd.n5952 585
R3235 gnd.n5955 gnd.n5954 585
R3236 gnd.n5957 gnd.n5956 585
R3237 gnd.n5959 gnd.n5958 585
R3238 gnd.n5961 gnd.n5960 585
R3239 gnd.n5963 gnd.n5962 585
R3240 gnd.n5965 gnd.n5964 585
R3241 gnd.n5967 gnd.n5966 585
R3242 gnd.n5969 gnd.n5968 585
R3243 gnd.n5971 gnd.n5970 585
R3244 gnd.n5973 gnd.n5972 585
R3245 gnd.n5975 gnd.n5974 585
R3246 gnd.n5977 gnd.n5976 585
R3247 gnd.n5979 gnd.n5978 585
R3248 gnd.n5981 gnd.n5980 585
R3249 gnd.n5983 gnd.n5982 585
R3250 gnd.n5985 gnd.n5984 585
R3251 gnd.n5987 gnd.n5986 585
R3252 gnd.n5989 gnd.n5988 585
R3253 gnd.n5991 gnd.n5990 585
R3254 gnd.n5993 gnd.n5992 585
R3255 gnd.n5994 gnd.n1525 585
R3256 gnd.n5999 gnd.n5998 585
R3257 gnd.n6882 gnd.n6881 585
R3258 gnd.n6883 gnd.n984 585
R3259 gnd.n6885 gnd.n6884 585
R3260 gnd.n6887 gnd.n982 585
R3261 gnd.n6889 gnd.n6888 585
R3262 gnd.n6890 gnd.n981 585
R3263 gnd.n6892 gnd.n6891 585
R3264 gnd.n6894 gnd.n979 585
R3265 gnd.n6896 gnd.n6895 585
R3266 gnd.n6897 gnd.n978 585
R3267 gnd.n6899 gnd.n6898 585
R3268 gnd.n6901 gnd.n976 585
R3269 gnd.n6903 gnd.n6902 585
R3270 gnd.n6904 gnd.n975 585
R3271 gnd.n6906 gnd.n6905 585
R3272 gnd.n6908 gnd.n973 585
R3273 gnd.n6910 gnd.n6909 585
R3274 gnd.n6911 gnd.n972 585
R3275 gnd.n6913 gnd.n6912 585
R3276 gnd.n6915 gnd.n970 585
R3277 gnd.n6917 gnd.n6916 585
R3278 gnd.n6918 gnd.n969 585
R3279 gnd.n6920 gnd.n6919 585
R3280 gnd.n6922 gnd.n967 585
R3281 gnd.n6924 gnd.n6923 585
R3282 gnd.n6925 gnd.n966 585
R3283 gnd.n6927 gnd.n6926 585
R3284 gnd.n6929 gnd.n964 585
R3285 gnd.n6931 gnd.n6930 585
R3286 gnd.n6933 gnd.n961 585
R3287 gnd.n6935 gnd.n6934 585
R3288 gnd.n6937 gnd.n786 585
R3289 gnd.n6938 gnd.n726 585
R3290 gnd.n6940 gnd.n785 585
R3291 gnd.n6942 gnd.n6941 585
R3292 gnd.n6944 gnd.n783 585
R3293 gnd.n6946 gnd.n6945 585
R3294 gnd.n6948 gnd.n780 585
R3295 gnd.n6950 gnd.n6949 585
R3296 gnd.n6952 gnd.n778 585
R3297 gnd.n6954 gnd.n6953 585
R3298 gnd.n6955 gnd.n777 585
R3299 gnd.n6957 gnd.n6956 585
R3300 gnd.n6959 gnd.n775 585
R3301 gnd.n6961 gnd.n6960 585
R3302 gnd.n6962 gnd.n774 585
R3303 gnd.n6964 gnd.n6963 585
R3304 gnd.n6966 gnd.n772 585
R3305 gnd.n6968 gnd.n6967 585
R3306 gnd.n6969 gnd.n771 585
R3307 gnd.n6971 gnd.n6970 585
R3308 gnd.n6973 gnd.n769 585
R3309 gnd.n6975 gnd.n6974 585
R3310 gnd.n6976 gnd.n768 585
R3311 gnd.n6978 gnd.n6977 585
R3312 gnd.n6980 gnd.n766 585
R3313 gnd.n6982 gnd.n6981 585
R3314 gnd.n6983 gnd.n765 585
R3315 gnd.n6985 gnd.n6984 585
R3316 gnd.n6987 gnd.n763 585
R3317 gnd.n6989 gnd.n6988 585
R3318 gnd.n6990 gnd.n762 585
R3319 gnd.n6992 gnd.n6991 585
R3320 gnd.n6994 gnd.n761 585
R3321 gnd.n6995 gnd.n760 585
R3322 gnd.n6998 gnd.n6997 585
R3323 gnd.n6880 gnd.n6876 585
R3324 gnd.n6880 gnd.n6879 585
R3325 gnd.n6875 gnd.n736 585
R3326 gnd.n7003 gnd.n736 585
R3327 gnd.n6874 gnd.n6873 585
R3328 gnd.n6873 gnd.n734 585
R3329 gnd.n6872 gnd.n985 585
R3330 gnd.n6872 gnd.n6871 585
R3331 gnd.n6781 gnd.n986 585
R3332 gnd.n6835 gnd.n986 585
R3333 gnd.n6782 gnd.n992 585
R3334 gnd.n6865 gnd.n992 585
R3335 gnd.n6787 gnd.n6783 585
R3336 gnd.n6787 gnd.n6786 585
R3337 gnd.n6788 gnd.n6780 585
R3338 gnd.n6788 gnd.n1001 585
R3339 gnd.n6790 gnd.n6789 585
R3340 gnd.n6789 gnd.n999 585
R3341 gnd.n6791 gnd.n1015 585
R3342 gnd.n6822 gnd.n1015 585
R3343 gnd.n6793 gnd.n6792 585
R3344 gnd.n6794 gnd.n6793 585
R3345 gnd.n6779 gnd.n1021 585
R3346 gnd.n6813 gnd.n1021 585
R3347 gnd.n6778 gnd.n6777 585
R3348 gnd.n6777 gnd.n6776 585
R3349 gnd.n6774 gnd.n1035 585
R3350 gnd.n6774 gnd.n1029 585
R3351 gnd.n6773 gnd.n6772 585
R3352 gnd.n6773 gnd.n1027 585
R3353 gnd.n6771 gnd.n1036 585
R3354 gnd.n6656 gnd.n1036 585
R3355 gnd.n6770 gnd.n6769 585
R3356 gnd.n6769 gnd.n6768 585
R3357 gnd.n1038 gnd.n1037 585
R3358 gnd.n1047 gnd.n1038 585
R3359 gnd.n1098 gnd.n1045 585
R3360 gnd.n6757 gnd.n1045 585
R3361 gnd.n6675 gnd.n6674 585
R3362 gnd.n6674 gnd.n6673 585
R3363 gnd.n6676 gnd.n1057 585
R3364 gnd.n6746 gnd.n1057 585
R3365 gnd.n6678 gnd.n6677 585
R3366 gnd.n6677 gnd.n1055 585
R3367 gnd.n6679 gnd.n1062 585
R3368 gnd.n6740 gnd.n1062 585
R3369 gnd.n6682 gnd.n6681 585
R3370 gnd.n6681 gnd.n6680 585
R3371 gnd.n6683 gnd.n1070 585
R3372 gnd.n6720 gnd.n1070 585
R3373 gnd.n6684 gnd.n1076 585
R3374 gnd.n6712 gnd.n1076 585
R3375 gnd.n6685 gnd.n1075 585
R3376 gnd.n6714 gnd.n1075 585
R3377 gnd.n6687 gnd.n6686 585
R3378 gnd.n6687 gnd.n1087 585
R3379 gnd.n6689 gnd.n6688 585
R3380 gnd.n6688 gnd.n1085 585
R3381 gnd.n6690 gnd.n1096 585
R3382 gnd.n6639 gnd.n1096 585
R3383 gnd.n6692 gnd.n6691 585
R3384 gnd.n6693 gnd.n6692 585
R3385 gnd.n1097 gnd.n1095 585
R3386 gnd.n6632 gnd.n1095 585
R3387 gnd.n6629 gnd.n6628 585
R3388 gnd.n6630 gnd.n6629 585
R3389 gnd.n6627 gnd.n1113 585
R3390 gnd.n6609 gnd.n1113 585
R3391 gnd.n6626 gnd.n6625 585
R3392 gnd.n6625 gnd.n6624 585
R3393 gnd.n1115 gnd.n1114 585
R3394 gnd.n1124 gnd.n1115 585
R3395 gnd.n6566 gnd.n1123 585
R3396 gnd.n6617 gnd.n1123 585
R3397 gnd.n6568 gnd.n6567 585
R3398 gnd.n6569 gnd.n6568 585
R3399 gnd.n6565 gnd.n1148 585
R3400 gnd.n6571 gnd.n1148 585
R3401 gnd.n6564 gnd.n6563 585
R3402 gnd.n6563 gnd.n1132 585
R3403 gnd.n6562 gnd.n1149 585
R3404 gnd.n6562 gnd.n6561 585
R3405 gnd.n6534 gnd.n1143 585
R3406 gnd.n6578 gnd.n1143 585
R3407 gnd.n6536 gnd.n6535 585
R3408 gnd.n6537 gnd.n6536 585
R3409 gnd.n6533 gnd.n1157 585
R3410 gnd.n1157 gnd.n1156 585
R3411 gnd.n6532 gnd.n6531 585
R3412 gnd.n6531 gnd.n6530 585
R3413 gnd.n1159 gnd.n1158 585
R3414 gnd.n1168 gnd.n1159 585
R3415 gnd.n6319 gnd.n1166 585
R3416 gnd.n6523 gnd.n1166 585
R3417 gnd.n6321 gnd.n6320 585
R3418 gnd.n6322 gnd.n6321 585
R3419 gnd.n6318 gnd.n1178 585
R3420 gnd.n6512 gnd.n1178 585
R3421 gnd.n6317 gnd.n6316 585
R3422 gnd.n6316 gnd.n1176 585
R3423 gnd.n1199 gnd.n1183 585
R3424 gnd.n6506 gnd.n1183 585
R3425 gnd.n6467 gnd.n6466 585
R3426 gnd.n6466 gnd.n6465 585
R3427 gnd.n6468 gnd.n1192 585
R3428 gnd.n6479 gnd.n1192 585
R3429 gnd.n6470 gnd.n6469 585
R3430 gnd.n6471 gnd.n6470 585
R3431 gnd.n1198 gnd.n1197 585
R3432 gnd.n6473 gnd.n1197 585
R3433 gnd.n1281 gnd.n1208 585
R3434 gnd.n6454 gnd.n1208 585
R3435 gnd.n1283 gnd.n1282 585
R3436 gnd.n1282 gnd.n1206 585
R3437 gnd.n1284 gnd.n1216 585
R3438 gnd.n6444 gnd.n1216 585
R3439 gnd.n1286 gnd.n1285 585
R3440 gnd.n1285 gnd.n1214 585
R3441 gnd.n1287 gnd.n1223 585
R3442 gnd.n6437 gnd.n1223 585
R3443 gnd.n6347 gnd.n6346 585
R3444 gnd.n6346 gnd.n6345 585
R3445 gnd.n6348 gnd.n1233 585
R3446 gnd.n6426 gnd.n1233 585
R3447 gnd.n6350 gnd.n6349 585
R3448 gnd.n6349 gnd.n1231 585
R3449 gnd.n6351 gnd.n1239 585
R3450 gnd.n6420 gnd.n1239 585
R3451 gnd.n6355 gnd.n6354 585
R3452 gnd.n6354 gnd.n6353 585
R3453 gnd.n6356 gnd.n1246 585
R3454 gnd.n6408 gnd.n1246 585
R3455 gnd.n6358 gnd.n6357 585
R3456 gnd.n6357 gnd.n1254 585
R3457 gnd.n6359 gnd.n1252 585
R3458 gnd.n6402 gnd.n1252 585
R3459 gnd.n6361 gnd.n6360 585
R3460 gnd.n6361 gnd.n1264 585
R3461 gnd.n6362 gnd.n1280 585
R3462 gnd.n6362 gnd.n1262 585
R3463 gnd.n6366 gnd.n6365 585
R3464 gnd.n6365 gnd.n6364 585
R3465 gnd.n6367 gnd.n1271 585
R3466 gnd.n6381 gnd.n1271 585
R3467 gnd.n6369 gnd.n6368 585
R3468 gnd.n6370 gnd.n6369 585
R3469 gnd.n1279 gnd.n1278 585
R3470 gnd.n6372 gnd.n1278 585
R3471 gnd.n1321 gnd.n1320 585
R3472 gnd.n1323 gnd.n1321 585
R3473 gnd.n6261 gnd.n6260 585
R3474 gnd.n6260 gnd.n6259 585
R3475 gnd.n6262 gnd.n1318 585
R3476 gnd.n1318 gnd.n1300 585
R3477 gnd.n6264 gnd.n6263 585
R3478 gnd.n6265 gnd.n6264 585
R3479 gnd.n1319 gnd.n1317 585
R3480 gnd.n6245 gnd.n1317 585
R3481 gnd.n6198 gnd.n1310 585
R3482 gnd.n6271 gnd.n1310 585
R3483 gnd.n6200 gnd.n6199 585
R3484 gnd.n6199 gnd.n1308 585
R3485 gnd.n6201 gnd.n1350 585
R3486 gnd.n6218 gnd.n1350 585
R3487 gnd.n6203 gnd.n6202 585
R3488 gnd.n6202 gnd.n1335 585
R3489 gnd.n6204 gnd.n1355 585
R3490 gnd.n1355 gnd.n1333 585
R3491 gnd.n6206 gnd.n6205 585
R3492 gnd.n6207 gnd.n6206 585
R3493 gnd.n6197 gnd.n1342 585
R3494 gnd.n6226 gnd.n1342 585
R3495 gnd.n6196 gnd.n6195 585
R3496 gnd.n6195 gnd.n6194 585
R3497 gnd.n1357 gnd.n1356 585
R3498 gnd.n6167 gnd.n1357 585
R3499 gnd.n1385 gnd.n1384 585
R3500 gnd.n1385 gnd.n1366 585
R3501 gnd.n1386 gnd.n1383 585
R3502 gnd.n1386 gnd.n1364 585
R3503 gnd.n6155 gnd.n6154 585
R3504 gnd.n6154 gnd.n6153 585
R3505 gnd.n6156 gnd.n1374 585
R3506 gnd.n6175 gnd.n1374 585
R3507 gnd.n6158 gnd.n6157 585
R3508 gnd.n6159 gnd.n6158 585
R3509 gnd.n1382 gnd.n1380 585
R3510 gnd.n6161 gnd.n1380 585
R3511 gnd.n6101 gnd.n1417 585
R3512 gnd.n1417 gnd.n1393 585
R3513 gnd.n6103 gnd.n6102 585
R3514 gnd.n6105 gnd.n6103 585
R3515 gnd.n6100 gnd.n1416 585
R3516 gnd.n1416 gnd.n1401 585
R3517 gnd.n6099 gnd.n6098 585
R3518 gnd.n6098 gnd.n1399 585
R3519 gnd.n6097 gnd.n6094 585
R3520 gnd.n6097 gnd.n6096 585
R3521 gnd.n6093 gnd.n1408 585
R3522 gnd.n6113 gnd.n1408 585
R3523 gnd.n6092 gnd.n6091 585
R3524 gnd.n6091 gnd.n6090 585
R3525 gnd.n1419 gnd.n1418 585
R3526 gnd.n6047 gnd.n1419 585
R3527 gnd.n6066 gnd.n6065 585
R3528 gnd.n6066 gnd.n1429 585
R3529 gnd.n6068 gnd.n6067 585
R3530 gnd.n6067 gnd.n1427 585
R3531 gnd.n6069 gnd.n1438 585
R3532 gnd.n6054 gnd.n1438 585
R3533 gnd.n6071 gnd.n6070 585
R3534 gnd.n6072 gnd.n6071 585
R3535 gnd.n6064 gnd.n1437 585
R3536 gnd.n1452 gnd.n1437 585
R3537 gnd.n6063 gnd.n6062 585
R3538 gnd.n6062 gnd.n6061 585
R3539 gnd.n1440 gnd.n1439 585
R3540 gnd.n6021 gnd.n1440 585
R3541 gnd.n5996 gnd.n5995 585
R3542 gnd.n5995 gnd.n1458 585
R3543 gnd.n5997 gnd.n1467 585
R3544 gnd.n6010 gnd.n1467 585
R3545 gnd.n5861 gnd.n1659 585
R3546 gnd.n5596 gnd.n1659 585
R3547 gnd.n5863 gnd.n5862 585
R3548 gnd.n5864 gnd.n5863 585
R3549 gnd.n1660 gnd.n1658 585
R3550 gnd.n1680 gnd.n1658 585
R3551 gnd.n5764 gnd.n5763 585
R3552 gnd.n5763 gnd.n5762 585
R3553 gnd.n1663 gnd.n1662 585
R3554 gnd.n5752 gnd.n1663 585
R3555 gnd.n5422 gnd.n5421 585
R3556 gnd.n5423 gnd.n5422 585
R3557 gnd.n1729 gnd.n1728 585
R3558 gnd.n1728 gnd.n1726 585
R3559 gnd.n5417 gnd.n5416 585
R3560 gnd.n5416 gnd.n5415 585
R3561 gnd.n1732 gnd.n1731 585
R3562 gnd.n5403 gnd.n1732 585
R3563 gnd.n5388 gnd.n1755 585
R3564 gnd.n5374 gnd.n1755 585
R3565 gnd.n5390 gnd.n5389 585
R3566 gnd.n5391 gnd.n5390 585
R3567 gnd.n1756 gnd.n1754 585
R3568 gnd.n5359 gnd.n1754 585
R3569 gnd.n5383 gnd.n5382 585
R3570 gnd.n5382 gnd.n5381 585
R3571 gnd.n1759 gnd.n1758 585
R3572 gnd.n5352 gnd.n1759 585
R3573 gnd.n5340 gnd.n1790 585
R3574 gnd.n5326 gnd.n1790 585
R3575 gnd.n5342 gnd.n5341 585
R3576 gnd.n5343 gnd.n5342 585
R3577 gnd.n1791 gnd.n1789 585
R3578 gnd.n5279 gnd.n1789 585
R3579 gnd.n5335 gnd.n5334 585
R3580 gnd.n5334 gnd.n5333 585
R3581 gnd.n1794 gnd.n1793 585
R3582 gnd.n5312 gnd.n1794 585
R3583 gnd.n5300 gnd.n1826 585
R3584 gnd.n1826 gnd.n1813 585
R3585 gnd.n5302 gnd.n5301 585
R3586 gnd.n5303 gnd.n5302 585
R3587 gnd.n1827 gnd.n1825 585
R3588 gnd.n5274 gnd.n1825 585
R3589 gnd.n5295 gnd.n5294 585
R3590 gnd.n5294 gnd.n5293 585
R3591 gnd.n1836 gnd.n1835 585
R3592 gnd.n5270 gnd.n1836 585
R3593 gnd.n5258 gnd.n5257 585
R3594 gnd.n5257 gnd.n1850 585
R3595 gnd.n5260 gnd.n5259 585
R3596 gnd.n5261 gnd.n5260 585
R3597 gnd.n5256 gnd.n1861 585
R3598 gnd.n5256 gnd.n5255 585
R3599 gnd.n1860 gnd.n1859 585
R3600 gnd.n1862 gnd.n1859 585
R3601 gnd.n5241 gnd.n5240 585
R3602 gnd.n5242 gnd.n5241 585
R3603 gnd.n5239 gnd.n1833 585
R3604 gnd.n5239 gnd.n1870 585
R3605 gnd.n5238 gnd.n1874 585
R3606 gnd.n5238 gnd.n5237 585
R3607 gnd.n5203 gnd.n1873 585
R3608 gnd.n5226 gnd.n1873 585
R3609 gnd.n5204 gnd.n1893 585
R3610 gnd.n1893 gnd.n1884 585
R3611 gnd.n5206 gnd.n5205 585
R3612 gnd.n5207 gnd.n5206 585
R3613 gnd.n1894 gnd.n1892 585
R3614 gnd.n1900 gnd.n1892 585
R3615 gnd.n5199 gnd.n5198 585
R3616 gnd.n5198 gnd.n5197 585
R3617 gnd.n1897 gnd.n1896 585
R3618 gnd.n5182 gnd.n1897 585
R3619 gnd.n5169 gnd.n1918 585
R3620 gnd.n1918 gnd.n1909 585
R3621 gnd.n5171 gnd.n5170 585
R3622 gnd.n5172 gnd.n5171 585
R3623 gnd.n1919 gnd.n1917 585
R3624 gnd.n1926 gnd.n1917 585
R3625 gnd.n5164 gnd.n5163 585
R3626 gnd.n5163 gnd.n5162 585
R3627 gnd.n1922 gnd.n1921 585
R3628 gnd.n1923 gnd.n1922 585
R3629 gnd.n5145 gnd.n5144 585
R3630 gnd.n5146 gnd.n5145 585
R3631 gnd.n1939 gnd.n1938 585
R3632 gnd.n1938 gnd.n1935 585
R3633 gnd.n5140 gnd.n5139 585
R3634 gnd.n5139 gnd.n5138 585
R3635 gnd.n1942 gnd.n1941 585
R3636 gnd.n1943 gnd.n1942 585
R3637 gnd.n5125 gnd.n5124 585
R3638 gnd.n5126 gnd.n5125 585
R3639 gnd.n1956 gnd.n1955 585
R3640 gnd.n1963 gnd.n1955 585
R3641 gnd.n5120 gnd.n5119 585
R3642 gnd.n5119 gnd.n5118 585
R3643 gnd.n1959 gnd.n1958 585
R3644 gnd.n1960 gnd.n1959 585
R3645 gnd.n5105 gnd.n5104 585
R3646 gnd.n5106 gnd.n5105 585
R3647 gnd.n1975 gnd.n1974 585
R3648 gnd.n1974 gnd.n1971 585
R3649 gnd.n5100 gnd.n5099 585
R3650 gnd.n5099 gnd.n5098 585
R3651 gnd.n1978 gnd.n1977 585
R3652 gnd.n1979 gnd.n1978 585
R3653 gnd.n5086 gnd.n5085 585
R3654 gnd.n5084 gnd.n4813 585
R3655 gnd.n5083 gnd.n4812 585
R3656 gnd.n5088 gnd.n4812 585
R3657 gnd.n5082 gnd.n5081 585
R3658 gnd.n5080 gnd.n5079 585
R3659 gnd.n5078 gnd.n5077 585
R3660 gnd.n5076 gnd.n5075 585
R3661 gnd.n5074 gnd.n5073 585
R3662 gnd.n5072 gnd.n5071 585
R3663 gnd.n5070 gnd.n5069 585
R3664 gnd.n5068 gnd.n5067 585
R3665 gnd.n5066 gnd.n5065 585
R3666 gnd.n5064 gnd.n5063 585
R3667 gnd.n5062 gnd.n5061 585
R3668 gnd.n5060 gnd.n5059 585
R3669 gnd.n5058 gnd.n5057 585
R3670 gnd.n5056 gnd.n5055 585
R3671 gnd.n5054 gnd.n5053 585
R3672 gnd.n5051 gnd.n5050 585
R3673 gnd.n5049 gnd.n5048 585
R3674 gnd.n5047 gnd.n5046 585
R3675 gnd.n5045 gnd.n5044 585
R3676 gnd.n5043 gnd.n5042 585
R3677 gnd.n5041 gnd.n5040 585
R3678 gnd.n5039 gnd.n5038 585
R3679 gnd.n5037 gnd.n5036 585
R3680 gnd.n5035 gnd.n5034 585
R3681 gnd.n5033 gnd.n5032 585
R3682 gnd.n5031 gnd.n5030 585
R3683 gnd.n5029 gnd.n5028 585
R3684 gnd.n5027 gnd.n5026 585
R3685 gnd.n5025 gnd.n5024 585
R3686 gnd.n5023 gnd.n5022 585
R3687 gnd.n5021 gnd.n5020 585
R3688 gnd.n5019 gnd.n5018 585
R3689 gnd.n5017 gnd.n5016 585
R3690 gnd.n5015 gnd.n5014 585
R3691 gnd.n5013 gnd.n5012 585
R3692 gnd.n5011 gnd.n5010 585
R3693 gnd.n5009 gnd.n5008 585
R3694 gnd.n5007 gnd.n5006 585
R3695 gnd.n5005 gnd.n5004 585
R3696 gnd.n5003 gnd.n5002 585
R3697 gnd.n5001 gnd.n5000 585
R3698 gnd.n4999 gnd.n4998 585
R3699 gnd.n4997 gnd.n4996 585
R3700 gnd.n4995 gnd.n4994 585
R3701 gnd.n4993 gnd.n4992 585
R3702 gnd.n4991 gnd.n4990 585
R3703 gnd.n4989 gnd.n4988 585
R3704 gnd.n4987 gnd.n4986 585
R3705 gnd.n4985 gnd.n4984 585
R3706 gnd.n4983 gnd.n4982 585
R3707 gnd.n4981 gnd.n4980 585
R3708 gnd.n4979 gnd.n4978 585
R3709 gnd.n4977 gnd.n4976 585
R3710 gnd.n4975 gnd.n4974 585
R3711 gnd.n4973 gnd.n1991 585
R3712 gnd.n5090 gnd.n1990 585
R3713 gnd.n5872 gnd.n5871 585
R3714 gnd.n5874 gnd.n1645 585
R3715 gnd.n5876 gnd.n5875 585
R3716 gnd.n5877 gnd.n1638 585
R3717 gnd.n5879 gnd.n5878 585
R3718 gnd.n5881 gnd.n1636 585
R3719 gnd.n5883 gnd.n5882 585
R3720 gnd.n5884 gnd.n1631 585
R3721 gnd.n5886 gnd.n5885 585
R3722 gnd.n5888 gnd.n1629 585
R3723 gnd.n5890 gnd.n5889 585
R3724 gnd.n5891 gnd.n1624 585
R3725 gnd.n5893 gnd.n5892 585
R3726 gnd.n5895 gnd.n1622 585
R3727 gnd.n5897 gnd.n5896 585
R3728 gnd.n5898 gnd.n1617 585
R3729 gnd.n5900 gnd.n5899 585
R3730 gnd.n5902 gnd.n1616 585
R3731 gnd.n5903 gnd.n1613 585
R3732 gnd.n5906 gnd.n5905 585
R3733 gnd.n1615 gnd.n1609 585
R3734 gnd.n5910 gnd.n1606 585
R3735 gnd.n5912 gnd.n5911 585
R3736 gnd.n5914 gnd.n1604 585
R3737 gnd.n5916 gnd.n5915 585
R3738 gnd.n5917 gnd.n1599 585
R3739 gnd.n5919 gnd.n5918 585
R3740 gnd.n5921 gnd.n1598 585
R3741 gnd.n5922 gnd.n1594 585
R3742 gnd.n5925 gnd.n5924 585
R3743 gnd.n1595 gnd.n1589 585
R3744 gnd.n5814 gnd.n1590 585
R3745 gnd.n5816 gnd.n5815 585
R3746 gnd.n5817 gnd.n5807 585
R3747 gnd.n5819 gnd.n5818 585
R3748 gnd.n5821 gnd.n5805 585
R3749 gnd.n5823 gnd.n5822 585
R3750 gnd.n5824 gnd.n5797 585
R3751 gnd.n5826 gnd.n5825 585
R3752 gnd.n5828 gnd.n5795 585
R3753 gnd.n5830 gnd.n5829 585
R3754 gnd.n5831 gnd.n5790 585
R3755 gnd.n5833 gnd.n5832 585
R3756 gnd.n5835 gnd.n5788 585
R3757 gnd.n5837 gnd.n5836 585
R3758 gnd.n5838 gnd.n5783 585
R3759 gnd.n5840 gnd.n5839 585
R3760 gnd.n5842 gnd.n5781 585
R3761 gnd.n5844 gnd.n5843 585
R3762 gnd.n5845 gnd.n5776 585
R3763 gnd.n5847 gnd.n5846 585
R3764 gnd.n5849 gnd.n5774 585
R3765 gnd.n5851 gnd.n5850 585
R3766 gnd.n5852 gnd.n5770 585
R3767 gnd.n5854 gnd.n5853 585
R3768 gnd.n5856 gnd.n5769 585
R3769 gnd.n5858 gnd.n5857 585
R3770 gnd.n5857 gnd.n1597 585
R3771 gnd.n5867 gnd.n1647 585
R3772 gnd.n5596 gnd.n1647 585
R3773 gnd.n5866 gnd.n5865 585
R3774 gnd.n5865 gnd.n5864 585
R3775 gnd.n1653 gnd.n1652 585
R3776 gnd.n1680 gnd.n1653 585
R3777 gnd.n5755 gnd.n1665 585
R3778 gnd.n5762 gnd.n1665 585
R3779 gnd.n5754 gnd.n5753 585
R3780 gnd.n5753 gnd.n5752 585
R3781 gnd.n1673 gnd.n1672 585
R3782 gnd.n5423 gnd.n1673 585
R3783 gnd.n5408 gnd.n5407 585
R3784 gnd.n5407 gnd.n1726 585
R3785 gnd.n5406 gnd.n1734 585
R3786 gnd.n5415 gnd.n1734 585
R3787 gnd.n5405 gnd.n5404 585
R3788 gnd.n5404 gnd.n5403 585
R3789 gnd.n1743 gnd.n1741 585
R3790 gnd.n5374 gnd.n1743 585
R3791 gnd.n5356 gnd.n1752 585
R3792 gnd.n5391 gnd.n1752 585
R3793 gnd.n5358 gnd.n5357 585
R3794 gnd.n5359 gnd.n5358 585
R3795 gnd.n5355 gnd.n1761 585
R3796 gnd.n5381 gnd.n1761 585
R3797 gnd.n5354 gnd.n5353 585
R3798 gnd.n5353 gnd.n5352 585
R3799 gnd.n1778 gnd.n1776 585
R3800 gnd.n5326 gnd.n1778 585
R3801 gnd.n5278 gnd.n1787 585
R3802 gnd.n5343 gnd.n1787 585
R3803 gnd.n5281 gnd.n5280 585
R3804 gnd.n5280 gnd.n5279 585
R3805 gnd.n5282 gnd.n1796 585
R3806 gnd.n5333 gnd.n1796 585
R3807 gnd.n5283 gnd.n1814 585
R3808 gnd.n5312 gnd.n1814 585
R3809 gnd.n5285 gnd.n5284 585
R3810 gnd.n5284 gnd.n1813 585
R3811 gnd.n5277 gnd.n1822 585
R3812 gnd.n5303 gnd.n1822 585
R3813 gnd.n5276 gnd.n5275 585
R3814 gnd.n5275 gnd.n5274 585
R3815 gnd.n5273 gnd.n1837 585
R3816 gnd.n5293 gnd.n1837 585
R3817 gnd.n5272 gnd.n5271 585
R3818 gnd.n5271 gnd.n5270 585
R3819 gnd.n1849 gnd.n1847 585
R3820 gnd.n1850 gnd.n1849 585
R3821 gnd.n5247 gnd.n1857 585
R3822 gnd.n5261 gnd.n1857 585
R3823 gnd.n5246 gnd.n1863 585
R3824 gnd.n5255 gnd.n1863 585
R3825 gnd.n5245 gnd.n5244 585
R3826 gnd.n5244 gnd.n1862 585
R3827 gnd.n5243 gnd.n1867 585
R3828 gnd.n5243 gnd.n5242 585
R3829 gnd.n5230 gnd.n1869 585
R3830 gnd.n1870 gnd.n1869 585
R3831 gnd.n5229 gnd.n1875 585
R3832 gnd.n5237 gnd.n1875 585
R3833 gnd.n5228 gnd.n5227 585
R3834 gnd.n5227 gnd.n5226 585
R3835 gnd.n1883 gnd.n1881 585
R3836 gnd.n1884 gnd.n1883 585
R3837 gnd.n5188 gnd.n1890 585
R3838 gnd.n5207 gnd.n1890 585
R3839 gnd.n5187 gnd.n5186 585
R3840 gnd.n5186 gnd.n1900 585
R3841 gnd.n5185 gnd.n1898 585
R3842 gnd.n5197 gnd.n1898 585
R3843 gnd.n5184 gnd.n5183 585
R3844 gnd.n5183 gnd.n5182 585
R3845 gnd.n1908 gnd.n1906 585
R3846 gnd.n1909 gnd.n1908 585
R3847 gnd.n5153 gnd.n1915 585
R3848 gnd.n5172 gnd.n1915 585
R3849 gnd.n5152 gnd.n5151 585
R3850 gnd.n5151 gnd.n1926 585
R3851 gnd.n5150 gnd.n1924 585
R3852 gnd.n5162 gnd.n1924 585
R3853 gnd.n5149 gnd.n5148 585
R3854 gnd.n5148 gnd.n1923 585
R3855 gnd.n5147 gnd.n1932 585
R3856 gnd.n5147 gnd.n5146 585
R3857 gnd.n5131 gnd.n1934 585
R3858 gnd.n1935 gnd.n1934 585
R3859 gnd.n5130 gnd.n1944 585
R3860 gnd.n5138 gnd.n1944 585
R3861 gnd.n5129 gnd.n5128 585
R3862 gnd.n5128 gnd.n1943 585
R3863 gnd.n5127 gnd.n1950 585
R3864 gnd.n5127 gnd.n5126 585
R3865 gnd.n5111 gnd.n1952 585
R3866 gnd.n1963 gnd.n1952 585
R3867 gnd.n5110 gnd.n1961 585
R3868 gnd.n5118 gnd.n1961 585
R3869 gnd.n5109 gnd.n5108 585
R3870 gnd.n5108 gnd.n1960 585
R3871 gnd.n5107 gnd.n1968 585
R3872 gnd.n5107 gnd.n5106 585
R3873 gnd.n5093 gnd.n1970 585
R3874 gnd.n1971 gnd.n1970 585
R3875 gnd.n5094 gnd.n1980 585
R3876 gnd.n5098 gnd.n1980 585
R3877 gnd.n5092 gnd.n5091 585
R3878 gnd.n5091 gnd.n1979 585
R3879 gnd.n7678 gnd.n7677 585
R3880 gnd.n7679 gnd.n7678 585
R3881 gnd.n200 gnd.n199 585
R3882 gnd.n208 gnd.n200 585
R3883 gnd.n7687 gnd.n7686 585
R3884 gnd.n7686 gnd.n7685 585
R3885 gnd.n7688 gnd.n194 585
R3886 gnd.n194 gnd.n193 585
R3887 gnd.n7690 gnd.n7689 585
R3888 gnd.n7691 gnd.n7690 585
R3889 gnd.n181 gnd.n180 585
R3890 gnd.n184 gnd.n181 585
R3891 gnd.n7699 gnd.n7698 585
R3892 gnd.n7698 gnd.n7697 585
R3893 gnd.n7700 gnd.n175 585
R3894 gnd.n175 gnd.n174 585
R3895 gnd.n7702 gnd.n7701 585
R3896 gnd.n7703 gnd.n7702 585
R3897 gnd.n161 gnd.n160 585
R3898 gnd.n7514 gnd.n161 585
R3899 gnd.n7711 gnd.n7710 585
R3900 gnd.n7710 gnd.n7709 585
R3901 gnd.n7712 gnd.n155 585
R3902 gnd.n162 gnd.n155 585
R3903 gnd.n7714 gnd.n7713 585
R3904 gnd.n7715 gnd.n7714 585
R3905 gnd.n143 gnd.n142 585
R3906 gnd.n146 gnd.n143 585
R3907 gnd.n7723 gnd.n7722 585
R3908 gnd.n7722 gnd.n7721 585
R3909 gnd.n7724 gnd.n137 585
R3910 gnd.n137 gnd.n136 585
R3911 gnd.n7726 gnd.n7725 585
R3912 gnd.n7727 gnd.n7726 585
R3913 gnd.n123 gnd.n122 585
R3914 gnd.n133 gnd.n123 585
R3915 gnd.n7735 gnd.n7734 585
R3916 gnd.n7734 gnd.n7733 585
R3917 gnd.n7736 gnd.n118 585
R3918 gnd.n124 gnd.n118 585
R3919 gnd.n7738 gnd.n7737 585
R3920 gnd.n7739 gnd.n7738 585
R3921 gnd.n104 gnd.n102 585
R3922 gnd.n107 gnd.n104 585
R3923 gnd.n7747 gnd.n7746 585
R3924 gnd.n7746 gnd.n7745 585
R3925 gnd.n103 gnd.n95 585
R3926 gnd.n7472 gnd.n103 585
R3927 gnd.n7750 gnd.n93 585
R3928 gnd.n93 gnd.n90 585
R3929 gnd.n7752 gnd.n7751 585
R3930 gnd.n7753 gnd.n7752 585
R3931 gnd.n7414 gnd.n92 585
R3932 gnd.n7428 gnd.n92 585
R3933 gnd.n7416 gnd.n7415 585
R3934 gnd.n7416 gnd.n364 585
R3935 gnd.n7418 gnd.n7417 585
R3936 gnd.n7419 gnd.n7418 585
R3937 gnd.n7413 gnd.n100 585
R3938 gnd.n7413 gnd.n370 585
R3939 gnd.n7412 gnd.n375 585
R3940 gnd.n7412 gnd.n7411 585
R3941 gnd.n7384 gnd.n374 585
R3942 gnd.n7402 gnd.n374 585
R3943 gnd.n7385 gnd.n394 585
R3944 gnd.n7371 gnd.n394 585
R3945 gnd.n7387 gnd.n7386 585
R3946 gnd.n7388 gnd.n7387 585
R3947 gnd.n395 gnd.n393 585
R3948 gnd.n7365 gnd.n393 585
R3949 gnd.n7380 gnd.n7379 585
R3950 gnd.n7379 gnd.n7378 585
R3951 gnd.n398 gnd.n397 585
R3952 gnd.n7353 gnd.n398 585
R3953 gnd.n7341 gnd.n426 585
R3954 gnd.n7327 gnd.n426 585
R3955 gnd.n7343 gnd.n7342 585
R3956 gnd.n7344 gnd.n7343 585
R3957 gnd.n427 gnd.n425 585
R3958 gnd.n7319 gnd.n425 585
R3959 gnd.n7336 gnd.n7335 585
R3960 gnd.n7335 gnd.n7334 585
R3961 gnd.n430 gnd.n429 585
R3962 gnd.n7306 gnd.n430 585
R3963 gnd.n7294 gnd.n461 585
R3964 gnd.n461 gnd.n449 585
R3965 gnd.n7296 gnd.n7295 585
R3966 gnd.n7297 gnd.n7296 585
R3967 gnd.n462 gnd.n460 585
R3968 gnd.n7273 gnd.n460 585
R3969 gnd.n7289 gnd.n7288 585
R3970 gnd.n7288 gnd.n7287 585
R3971 gnd.n465 gnd.n464 585
R3972 gnd.n7260 gnd.n465 585
R3973 gnd.n7248 gnd.n496 585
R3974 gnd.n496 gnd.n483 585
R3975 gnd.n7250 gnd.n7249 585
R3976 gnd.n7251 gnd.n7250 585
R3977 gnd.n497 gnd.n495 585
R3978 gnd.n7227 gnd.n495 585
R3979 gnd.n7243 gnd.n7242 585
R3980 gnd.n7242 gnd.n7241 585
R3981 gnd.n500 gnd.n499 585
R3982 gnd.n7223 gnd.n500 585
R3983 gnd.n7211 gnd.n525 585
R3984 gnd.n7097 gnd.n525 585
R3985 gnd.n7213 gnd.n7212 585
R3986 gnd.n7214 gnd.n7213 585
R3987 gnd.n7207 gnd.n524 585
R3988 gnd.n7206 gnd.n7205 585
R3989 gnd.n528 gnd.n527 585
R3990 gnd.n7203 gnd.n528 585
R3991 gnd.n805 gnd.n804 585
R3992 gnd.n807 gnd.n806 585
R3993 gnd.n809 gnd.n808 585
R3994 gnd.n813 gnd.n800 585
R3995 gnd.n815 gnd.n814 585
R3996 gnd.n817 gnd.n816 585
R3997 gnd.n819 gnd.n818 585
R3998 gnd.n823 gnd.n798 585
R3999 gnd.n825 gnd.n824 585
R4000 gnd.n827 gnd.n826 585
R4001 gnd.n829 gnd.n828 585
R4002 gnd.n833 gnd.n796 585
R4003 gnd.n835 gnd.n834 585
R4004 gnd.n837 gnd.n836 585
R4005 gnd.n839 gnd.n838 585
R4006 gnd.n843 gnd.n842 585
R4007 gnd.n845 gnd.n844 585
R4008 gnd.n848 gnd.n847 585
R4009 gnd.n846 gnd.n790 585
R4010 gnd.n853 gnd.n852 585
R4011 gnd.n855 gnd.n854 585
R4012 gnd.n858 gnd.n857 585
R4013 gnd.n856 gnd.n787 585
R4014 gnd.n958 gnd.n957 585
R4015 gnd.n956 gnd.n955 585
R4016 gnd.n954 gnd.n953 585
R4017 gnd.n952 gnd.n951 585
R4018 gnd.n950 gnd.n949 585
R4019 gnd.n948 gnd.n947 585
R4020 gnd.n946 gnd.n945 585
R4021 gnd.n944 gnd.n943 585
R4022 gnd.n942 gnd.n941 585
R4023 gnd.n940 gnd.n939 585
R4024 gnd.n938 gnd.n937 585
R4025 gnd.n936 gnd.n935 585
R4026 gnd.n934 gnd.n933 585
R4027 gnd.n932 gnd.n931 585
R4028 gnd.n930 gnd.n929 585
R4029 gnd.n928 gnd.n927 585
R4030 gnd.n926 gnd.n925 585
R4031 gnd.n924 gnd.n923 585
R4032 gnd.n922 gnd.n921 585
R4033 gnd.n920 gnd.n919 585
R4034 gnd.n918 gnd.n917 585
R4035 gnd.n916 gnd.n915 585
R4036 gnd.n914 gnd.n913 585
R4037 gnd.n912 gnd.n911 585
R4038 gnd.n910 gnd.n909 585
R4039 gnd.n908 gnd.n907 585
R4040 gnd.n906 gnd.n905 585
R4041 gnd.n904 gnd.n903 585
R4042 gnd.n902 gnd.n901 585
R4043 gnd.n900 gnd.n899 585
R4044 gnd.n894 gnd.n893 585
R4045 gnd.n7569 gnd.n7568 585
R4046 gnd.n7571 gnd.n314 585
R4047 gnd.n7573 gnd.n7572 585
R4048 gnd.n7574 gnd.n307 585
R4049 gnd.n7576 gnd.n7575 585
R4050 gnd.n7578 gnd.n305 585
R4051 gnd.n7580 gnd.n7579 585
R4052 gnd.n7581 gnd.n300 585
R4053 gnd.n7583 gnd.n7582 585
R4054 gnd.n7585 gnd.n298 585
R4055 gnd.n7587 gnd.n7586 585
R4056 gnd.n7588 gnd.n293 585
R4057 gnd.n7590 gnd.n7589 585
R4058 gnd.n7592 gnd.n291 585
R4059 gnd.n7594 gnd.n7593 585
R4060 gnd.n7595 gnd.n286 585
R4061 gnd.n7597 gnd.n7596 585
R4062 gnd.n7599 gnd.n285 585
R4063 gnd.n7600 gnd.n282 585
R4064 gnd.n7603 gnd.n7602 585
R4065 gnd.n284 gnd.n278 585
R4066 gnd.n7607 gnd.n275 585
R4067 gnd.n7609 gnd.n7608 585
R4068 gnd.n7611 gnd.n273 585
R4069 gnd.n7613 gnd.n7612 585
R4070 gnd.n7614 gnd.n268 585
R4071 gnd.n7616 gnd.n7615 585
R4072 gnd.n7618 gnd.n266 585
R4073 gnd.n7620 gnd.n7619 585
R4074 gnd.n7621 gnd.n261 585
R4075 gnd.n7623 gnd.n7622 585
R4076 gnd.n7625 gnd.n259 585
R4077 gnd.n7627 gnd.n7626 585
R4078 gnd.n7628 gnd.n254 585
R4079 gnd.n7630 gnd.n7629 585
R4080 gnd.n7632 gnd.n252 585
R4081 gnd.n7634 gnd.n7633 585
R4082 gnd.n7635 gnd.n247 585
R4083 gnd.n7637 gnd.n7636 585
R4084 gnd.n7639 gnd.n245 585
R4085 gnd.n7641 gnd.n7640 585
R4086 gnd.n7645 gnd.n240 585
R4087 gnd.n7647 gnd.n7646 585
R4088 gnd.n7649 gnd.n238 585
R4089 gnd.n7651 gnd.n7650 585
R4090 gnd.n7652 gnd.n233 585
R4091 gnd.n7654 gnd.n7653 585
R4092 gnd.n7656 gnd.n231 585
R4093 gnd.n7658 gnd.n7657 585
R4094 gnd.n7659 gnd.n226 585
R4095 gnd.n7661 gnd.n7660 585
R4096 gnd.n7663 gnd.n224 585
R4097 gnd.n7665 gnd.n7664 585
R4098 gnd.n7666 gnd.n219 585
R4099 gnd.n7668 gnd.n7667 585
R4100 gnd.n7670 gnd.n217 585
R4101 gnd.n7672 gnd.n7671 585
R4102 gnd.n7673 gnd.n215 585
R4103 gnd.n7674 gnd.n212 585
R4104 gnd.n212 gnd.n211 585
R4105 gnd.n7499 gnd.n209 585
R4106 gnd.n7679 gnd.n209 585
R4107 gnd.n7501 gnd.n7500 585
R4108 gnd.n7500 gnd.n208 585
R4109 gnd.n7502 gnd.n201 585
R4110 gnd.n7685 gnd.n201 585
R4111 gnd.n7504 gnd.n7503 585
R4112 gnd.n7503 gnd.n193 585
R4113 gnd.n7505 gnd.n191 585
R4114 gnd.n7691 gnd.n191 585
R4115 gnd.n7507 gnd.n7506 585
R4116 gnd.n7506 gnd.n184 585
R4117 gnd.n7508 gnd.n182 585
R4118 gnd.n7697 gnd.n182 585
R4119 gnd.n7510 gnd.n7509 585
R4120 gnd.n7509 gnd.n174 585
R4121 gnd.n7511 gnd.n172 585
R4122 gnd.n7703 gnd.n172 585
R4123 gnd.n7513 gnd.n7512 585
R4124 gnd.n7514 gnd.n7513 585
R4125 gnd.n7496 gnd.n163 585
R4126 gnd.n7709 gnd.n163 585
R4127 gnd.n7495 gnd.n7494 585
R4128 gnd.n7494 gnd.n162 585
R4129 gnd.n7492 gnd.n153 585
R4130 gnd.n7715 gnd.n153 585
R4131 gnd.n7491 gnd.n7490 585
R4132 gnd.n7490 gnd.n146 585
R4133 gnd.n7489 gnd.n144 585
R4134 gnd.n7721 gnd.n144 585
R4135 gnd.n7488 gnd.n7487 585
R4136 gnd.n7487 gnd.n136 585
R4137 gnd.n7485 gnd.n134 585
R4138 gnd.n7727 gnd.n134 585
R4139 gnd.n7484 gnd.n7483 585
R4140 gnd.n7483 gnd.n133 585
R4141 gnd.n7482 gnd.n125 585
R4142 gnd.n7733 gnd.n125 585
R4143 gnd.n7481 gnd.n7480 585
R4144 gnd.n7480 gnd.n124 585
R4145 gnd.n7478 gnd.n116 585
R4146 gnd.n7739 gnd.n116 585
R4147 gnd.n7477 gnd.n7476 585
R4148 gnd.n7476 gnd.n107 585
R4149 gnd.n7475 gnd.n105 585
R4150 gnd.n7745 gnd.n105 585
R4151 gnd.n7474 gnd.n7473 585
R4152 gnd.n7473 gnd.n7472 585
R4153 gnd.n7436 gnd.n359 585
R4154 gnd.n7436 gnd.n90 585
R4155 gnd.n7425 gnd.n89 585
R4156 gnd.n7753 gnd.n89 585
R4157 gnd.n7427 gnd.n7426 585
R4158 gnd.n7428 gnd.n7427 585
R4159 gnd.n7424 gnd.n365 585
R4160 gnd.n365 gnd.n364 585
R4161 gnd.n371 gnd.n366 585
R4162 gnd.n7419 gnd.n371 585
R4163 gnd.n7406 gnd.n7405 585
R4164 gnd.n7405 gnd.n370 585
R4165 gnd.n7407 gnd.n376 585
R4166 gnd.n7411 gnd.n376 585
R4167 gnd.n7404 gnd.n7403 585
R4168 gnd.n7403 gnd.n7402 585
R4169 gnd.n382 gnd.n381 585
R4170 gnd.n7371 gnd.n382 585
R4171 gnd.n7368 gnd.n390 585
R4172 gnd.n7388 gnd.n390 585
R4173 gnd.n7367 gnd.n7366 585
R4174 gnd.n7366 gnd.n7365 585
R4175 gnd.n407 gnd.n399 585
R4176 gnd.n7378 gnd.n399 585
R4177 gnd.n7324 gnd.n415 585
R4178 gnd.n7353 gnd.n415 585
R4179 gnd.n7326 gnd.n7325 585
R4180 gnd.n7327 gnd.n7326 585
R4181 gnd.n7322 gnd.n422 585
R4182 gnd.n7344 gnd.n422 585
R4183 gnd.n7321 gnd.n7320 585
R4184 gnd.n7320 gnd.n7319 585
R4185 gnd.n442 gnd.n432 585
R4186 gnd.n7334 gnd.n432 585
R4187 gnd.n7277 gnd.n450 585
R4188 gnd.n7306 gnd.n450 585
R4189 gnd.n7279 gnd.n7278 585
R4190 gnd.n7278 gnd.n449 585
R4191 gnd.n7276 gnd.n457 585
R4192 gnd.n7297 gnd.n457 585
R4193 gnd.n7275 gnd.n7274 585
R4194 gnd.n7274 gnd.n7273 585
R4195 gnd.n477 gnd.n467 585
R4196 gnd.n7287 gnd.n467 585
R4197 gnd.n7231 gnd.n484 585
R4198 gnd.n7260 gnd.n484 585
R4199 gnd.n7233 gnd.n7232 585
R4200 gnd.n7232 gnd.n483 585
R4201 gnd.n7230 gnd.n492 585
R4202 gnd.n7251 gnd.n492 585
R4203 gnd.n7229 gnd.n7228 585
R4204 gnd.n7228 gnd.n7227 585
R4205 gnd.n7226 gnd.n502 585
R4206 gnd.n7241 gnd.n502 585
R4207 gnd.n7225 gnd.n7224 585
R4208 gnd.n7224 gnd.n7223 585
R4209 gnd.n514 gnd.n512 585
R4210 gnd.n7097 gnd.n514 585
R4211 gnd.n7092 gnd.n521 585
R4212 gnd.n7214 gnd.n521 585
R4213 gnd.n3374 gnd.n2082 585
R4214 gnd.n2082 gnd.n1839 585
R4215 gnd.n2682 gnd.n2681 585
R4216 gnd.n2682 gnd.n383 585
R4217 gnd.n7361 gnd.n409 585
R4218 gnd.n409 gnd.n391 585
R4219 gnd.n7363 gnd.n7362 585
R4220 gnd.n7364 gnd.n7363 585
R4221 gnd.n410 gnd.n408 585
R4222 gnd.n408 gnd.n401 585
R4223 gnd.n7356 gnd.n7355 585
R4224 gnd.n7355 gnd.n7354 585
R4225 gnd.n413 gnd.n412 585
R4226 gnd.n414 gnd.n413 585
R4227 gnd.n7315 gnd.n444 585
R4228 gnd.n444 gnd.n423 585
R4229 gnd.n7317 gnd.n7316 585
R4230 gnd.n7318 gnd.n7317 585
R4231 gnd.n445 gnd.n443 585
R4232 gnd.n443 gnd.n434 585
R4233 gnd.n7310 gnd.n7309 585
R4234 gnd.n7309 gnd.n431 585
R4235 gnd.n7308 gnd.n447 585
R4236 gnd.n7308 gnd.n7307 585
R4237 gnd.n7269 gnd.n448 585
R4238 gnd.n458 gnd.n448 585
R4239 gnd.n7271 gnd.n7270 585
R4240 gnd.n7272 gnd.n7271 585
R4241 gnd.n479 gnd.n478 585
R4242 gnd.n478 gnd.n469 585
R4243 gnd.n7264 gnd.n7263 585
R4244 gnd.n7263 gnd.n466 585
R4245 gnd.n7262 gnd.n481 585
R4246 gnd.n7262 gnd.n7261 585
R4247 gnd.n7108 gnd.n482 585
R4248 gnd.n493 gnd.n482 585
R4249 gnd.n7110 gnd.n7109 585
R4250 gnd.n7110 gnd.n491 585
R4251 gnd.n7111 gnd.n7104 585
R4252 gnd.n7111 gnd.n504 585
R4253 gnd.n7113 gnd.n7112 585
R4254 gnd.n7112 gnd.n501 585
R4255 gnd.n7114 gnd.n7099 585
R4256 gnd.n7099 gnd.n7098 585
R4257 gnd.n7116 gnd.n7115 585
R4258 gnd.n7116 gnd.n522 585
R4259 gnd.n7117 gnd.n7090 585
R4260 gnd.n7117 gnd.n520 585
R4261 gnd.n7119 gnd.n7118 585
R4262 gnd.n7118 gnd.n529 585
R4263 gnd.n7120 gnd.n671 585
R4264 gnd.n671 gnd.n669 585
R4265 gnd.n7122 gnd.n7121 585
R4266 gnd.n7123 gnd.n7122 585
R4267 gnd.n672 gnd.n670 585
R4268 gnd.n670 gnd.n647 585
R4269 gnd.n7084 gnd.n7083 585
R4270 gnd.n7083 gnd.n585 585
R4271 gnd.n7082 gnd.n674 585
R4272 gnd.n7082 gnd.n584 585
R4273 gnd.n7081 gnd.n676 585
R4274 gnd.n7081 gnd.n7080 585
R4275 gnd.n7066 gnd.n675 585
R4276 gnd.n677 gnd.n675 585
R4277 gnd.n7068 gnd.n7067 585
R4278 gnd.n7069 gnd.n7068 585
R4279 gnd.n688 gnd.n687 585
R4280 gnd.n687 gnd.n684 585
R4281 gnd.n7060 gnd.n7059 585
R4282 gnd.n7059 gnd.n7058 585
R4283 gnd.n691 gnd.n690 585
R4284 gnd.n700 gnd.n691 585
R4285 gnd.n7030 gnd.n712 585
R4286 gnd.n712 gnd.n699 585
R4287 gnd.n7032 gnd.n7031 585
R4288 gnd.n7033 gnd.n7032 585
R4289 gnd.n713 gnd.n711 585
R4290 gnd.n711 gnd.n708 585
R4291 gnd.n7025 gnd.n7024 585
R4292 gnd.n7024 gnd.n7023 585
R4293 gnd.n716 gnd.n715 585
R4294 gnd.n725 gnd.n716 585
R4295 gnd.n6857 gnd.n6856 585
R4296 gnd.n6857 gnd.n724 585
R4297 gnd.n6858 gnd.n6853 585
R4298 gnd.n6858 gnd.n737 585
R4299 gnd.n6861 gnd.n6860 585
R4300 gnd.n6860 gnd.n6859 585
R4301 gnd.n6862 gnd.n994 585
R4302 gnd.n994 gnd.n987 585
R4303 gnd.n6864 gnd.n6863 585
R4304 gnd.n6865 gnd.n6864 585
R4305 gnd.n995 gnd.n993 585
R4306 gnd.n6784 gnd.n993 585
R4307 gnd.n6847 gnd.n6846 585
R4308 gnd.n6846 gnd.n6845 585
R4309 gnd.n998 gnd.n997 585
R4310 gnd.n1014 gnd.n998 585
R4311 gnd.n6811 gnd.n6810 585
R4312 gnd.n6812 gnd.n6811 585
R4313 gnd.n1023 gnd.n1022 585
R4314 gnd.n6775 gnd.n1022 585
R4315 gnd.n6806 gnd.n6805 585
R4316 gnd.n6805 gnd.n6804 585
R4317 gnd.n1026 gnd.n1025 585
R4318 gnd.n6655 gnd.n1026 585
R4319 gnd.n6732 gnd.n6730 585
R4320 gnd.n6732 gnd.n6731 585
R4321 gnd.n6734 gnd.n6733 585
R4322 gnd.n6733 gnd.n1044 585
R4323 gnd.n6735 gnd.n1065 585
R4324 gnd.n1065 gnd.n1058 585
R4325 gnd.n6737 gnd.n6736 585
R4326 gnd.n6738 gnd.n6737 585
R4327 gnd.n1066 gnd.n1064 585
R4328 gnd.n1064 gnd.t31 585
R4329 gnd.n6723 gnd.n6722 585
R4330 gnd.n6722 gnd.n6721 585
R4331 gnd.n1069 gnd.n1068 585
R4332 gnd.n6713 gnd.n1069 585
R4333 gnd.n6700 gnd.n6699 585
R4334 gnd.n6701 gnd.n6700 585
R4335 gnd.n1089 gnd.n1088 585
R4336 gnd.n1108 gnd.n1088 585
R4337 gnd.n6695 gnd.n6694 585
R4338 gnd.n6694 gnd.n6693 585
R4339 gnd.n1092 gnd.n1091 585
R4340 gnd.n6631 gnd.n1092 585
R4341 gnd.n6612 gnd.n6611 585
R4342 gnd.n6611 gnd.n6610 585
R4343 gnd.n6613 gnd.n1127 585
R4344 gnd.n1127 gnd.n1116 585
R4345 gnd.n6615 gnd.n6614 585
R4346 gnd.n6616 gnd.n6615 585
R4347 gnd.n1128 gnd.n1126 585
R4348 gnd.n6570 gnd.n1126 585
R4349 gnd.n6603 gnd.n6602 585
R4350 gnd.n6602 gnd.n6601 585
R4351 gnd.n1131 gnd.n1130 585
R4352 gnd.n1150 gnd.n1131 585
R4353 gnd.n6493 gnd.n6489 585
R4354 gnd.n6489 gnd.n1141 585
R4355 gnd.n6496 gnd.n6494 585
R4356 gnd.n6496 gnd.n6495 585
R4357 gnd.n6498 gnd.n6488 585
R4358 gnd.n6498 gnd.n6497 585
R4359 gnd.n6500 gnd.n6499 585
R4360 gnd.n6499 gnd.n1165 585
R4361 gnd.n6501 gnd.n1186 585
R4362 gnd.n6315 gnd.n1186 585
R4363 gnd.n6503 gnd.n6502 585
R4364 gnd.n6504 gnd.n6503 585
R4365 gnd.n1187 gnd.n1185 585
R4366 gnd.n1185 gnd.n1182 585
R4367 gnd.n6482 gnd.n6481 585
R4368 gnd.n6481 gnd.n6480 585
R4369 gnd.n1190 gnd.n1189 585
R4370 gnd.n6472 gnd.n1190 585
R4371 gnd.n6453 gnd.n6452 585
R4372 gnd.n6454 gnd.n6453 585
R4373 gnd.n1210 gnd.n1209 585
R4374 gnd.n1217 gnd.n1209 585
R4375 gnd.n6448 gnd.n6447 585
R4376 gnd.n6447 gnd.n6446 585
R4377 gnd.n1213 gnd.n1212 585
R4378 gnd.n1222 gnd.n1213 585
R4379 gnd.n6416 gnd.n1241 585
R4380 gnd.n1241 gnd.n1234 585
R4381 gnd.n6418 gnd.n6417 585
R4382 gnd.n6419 gnd.n6418 585
R4383 gnd.n1242 gnd.n1240 585
R4384 gnd.n6352 gnd.n1240 585
R4385 gnd.n6411 gnd.n6410 585
R4386 gnd.n6410 gnd.n6409 585
R4387 gnd.n1245 gnd.n1244 585
R4388 gnd.n6401 gnd.n1245 585
R4389 gnd.n6389 gnd.n6388 585
R4390 gnd.n6390 gnd.n6389 585
R4391 gnd.n1266 gnd.n1265 585
R4392 gnd.n6363 gnd.n1265 585
R4393 gnd.n6384 gnd.n6383 585
R4394 gnd.n6383 gnd.n6382 585
R4395 gnd.n1269 gnd.n1268 585
R4396 gnd.n6371 gnd.n1269 585
R4397 gnd.n6254 gnd.n6253 585
R4398 gnd.n6255 gnd.n6254 585
R4399 gnd.n1325 gnd.n1324 585
R4400 gnd.n1324 gnd.n1322 585
R4401 gnd.n6249 gnd.n6248 585
R4402 gnd.n6248 gnd.n1316 585
R4403 gnd.n6247 gnd.n1327 585
R4404 gnd.n6247 gnd.n6246 585
R4405 gnd.n6243 gnd.n6242 585
R4406 gnd.n6243 gnd.n1308 585
R4407 gnd.n1329 gnd.n1328 585
R4408 gnd.n1349 gnd.n1328 585
R4409 gnd.n6238 gnd.n6237 585
R4410 gnd.n6237 gnd.n6236 585
R4411 gnd.n1332 gnd.n1331 585
R4412 gnd.n1343 gnd.n1332 585
R4413 gnd.n6192 gnd.n6191 585
R4414 gnd.n6193 gnd.n6192 585
R4415 gnd.n1360 gnd.n1359 585
R4416 gnd.t10 gnd.n1359 585
R4417 gnd.n6187 gnd.n6186 585
R4418 gnd.n6186 gnd.n6185 585
R4419 gnd.n1363 gnd.n1362 585
R4420 gnd.n1387 gnd.n1363 585
R4421 gnd.n6124 gnd.n6123 585
R4422 gnd.n6124 gnd.n1372 585
R4423 gnd.n6126 gnd.n6125 585
R4424 gnd.n6125 gnd.n1379 585
R4425 gnd.n6127 gnd.n1403 585
R4426 gnd.n6104 gnd.n1403 585
R4427 gnd.n6129 gnd.n6128 585
R4428 gnd.n6130 gnd.n6129 585
R4429 gnd.n1404 gnd.n1402 585
R4430 gnd.n6095 gnd.n1402 585
R4431 gnd.n6116 gnd.n6115 585
R4432 gnd.n6115 gnd.n6114 585
R4433 gnd.n1407 gnd.n1406 585
R4434 gnd.n1420 gnd.n1407 585
R4435 gnd.n6079 gnd.n6078 585
R4436 gnd.n6080 gnd.n6079 585
R4437 gnd.n1431 gnd.n1430 585
R4438 gnd.n6053 gnd.n1430 585
R4439 gnd.n6074 gnd.n6073 585
R4440 gnd.n6073 gnd.n6072 585
R4441 gnd.n1434 gnd.n1433 585
R4442 gnd.n1442 gnd.n1434 585
R4443 gnd.n6019 gnd.n6018 585
R4444 gnd.n6020 gnd.n6019 585
R4445 gnd.n1461 gnd.n1460 585
R4446 gnd.n1468 gnd.n1460 585
R4447 gnd.n6014 gnd.n6013 585
R4448 gnd.n6013 gnd.n6012 585
R4449 gnd.n1464 gnd.n1463 585
R4450 gnd.n1493 gnd.n1464 585
R4451 gnd.n5539 gnd.n5479 585
R4452 gnd.n5479 gnd.n5468 585
R4453 gnd.n5541 gnd.n5540 585
R4454 gnd.n5542 gnd.n5541 585
R4455 gnd.n5480 gnd.n5478 585
R4456 gnd.n5478 gnd.n5476 585
R4457 gnd.n5534 gnd.n5533 585
R4458 gnd.n5533 gnd.n5532 585
R4459 gnd.n5483 gnd.n5482 585
R4460 gnd.n5490 gnd.n5483 585
R4461 gnd.n5520 gnd.n5519 585
R4462 gnd.n5521 gnd.n5520 585
R4463 gnd.n5494 gnd.n5493 585
R4464 gnd.n5493 gnd.n5489 585
R4465 gnd.n5515 gnd.n5514 585
R4466 gnd.n5514 gnd.n5513 585
R4467 gnd.n5498 gnd.n5497 585
R4468 gnd.n5499 gnd.n5498 585
R4469 gnd.n5447 gnd.n5446 585
R4470 gnd.n5451 gnd.n5447 585
R4471 gnd.n5583 gnd.n5582 585
R4472 gnd.n5582 gnd.n5581 585
R4473 gnd.n5584 gnd.n5441 585
R4474 gnd.n5448 gnd.n5441 585
R4475 gnd.n5586 gnd.n5585 585
R4476 gnd.n5586 gnd.n1702 585
R4477 gnd.n5587 gnd.n5440 585
R4478 gnd.n5587 gnd.n1688 585
R4479 gnd.n5591 gnd.n5590 585
R4480 gnd.n5590 gnd.n5589 585
R4481 gnd.n5592 gnd.n1717 585
R4482 gnd.n5588 gnd.n1717 585
R4483 gnd.n5594 gnd.n5593 585
R4484 gnd.n5595 gnd.n5594 585
R4485 gnd.n1718 gnd.n1716 585
R4486 gnd.n1716 gnd.n1656 585
R4487 gnd.n5434 gnd.n5433 585
R4488 gnd.n5433 gnd.n1654 585
R4489 gnd.n5432 gnd.n1720 585
R4490 gnd.n5432 gnd.n1667 585
R4491 gnd.n5431 gnd.n5430 585
R4492 gnd.n5431 gnd.n1664 585
R4493 gnd.n1722 gnd.n1721 585
R4494 gnd.n1721 gnd.n1674 585
R4495 gnd.n5426 gnd.n5425 585
R4496 gnd.n5425 gnd.n5424 585
R4497 gnd.n1725 gnd.n1724 585
R4498 gnd.n1736 gnd.n1725 585
R4499 gnd.n5369 gnd.n5368 585
R4500 gnd.n5368 gnd.n1733 585
R4501 gnd.n5370 gnd.n1771 585
R4502 gnd.n1771 gnd.n1744 585
R4503 gnd.n5372 gnd.n5371 585
R4504 gnd.n5373 gnd.n5372 585
R4505 gnd.n1772 gnd.n1770 585
R4506 gnd.n1770 gnd.n1751 585
R4507 gnd.n5362 gnd.n5361 585
R4508 gnd.n5361 gnd.n5360 585
R4509 gnd.n1775 gnd.n1774 585
R4510 gnd.n1775 gnd.n1760 585
R4511 gnd.n5322 gnd.n1807 585
R4512 gnd.n1807 gnd.n1779 585
R4513 gnd.n5324 gnd.n5323 585
R4514 gnd.n5325 gnd.n5324 585
R4515 gnd.n1808 gnd.n1806 585
R4516 gnd.n1806 gnd.n1786 585
R4517 gnd.n5317 gnd.n5316 585
R4518 gnd.n5316 gnd.n1798 585
R4519 gnd.n5315 gnd.n1810 585
R4520 gnd.n5315 gnd.n1795 585
R4521 gnd.n5314 gnd.n1812 585
R4522 gnd.n5314 gnd.n5313 585
R4523 gnd.n2079 gnd.n1811 585
R4524 gnd.n1823 gnd.n1811 585
R4525 gnd.n2081 gnd.n2080 585
R4526 gnd.n2081 gnd.n1821 585
R4527 gnd.n7184 gnd.n7183 585
R4528 gnd.n7185 gnd.n7184 585
R4529 gnd.n588 gnd.n586 585
R4530 gnd.n7079 gnd.n586 585
R4531 gnd.n7077 gnd.n7076 585
R4532 gnd.n7078 gnd.n7077 585
R4533 gnd.n680 gnd.n679 585
R4534 gnd.n686 gnd.n679 585
R4535 gnd.n7072 gnd.n7071 585
R4536 gnd.n7071 gnd.n7070 585
R4537 gnd.n683 gnd.n682 585
R4538 gnd.n7057 gnd.n683 585
R4539 gnd.n704 gnd.n702 585
R4540 gnd.n702 gnd.n692 585
R4541 gnd.n7042 gnd.n7041 585
R4542 gnd.n7043 gnd.n7042 585
R4543 gnd.n703 gnd.n701 585
R4544 gnd.n710 gnd.n701 585
R4545 gnd.n7036 gnd.n7035 585
R4546 gnd.n7035 gnd.n7034 585
R4547 gnd.n707 gnd.n706 585
R4548 gnd.n7022 gnd.n707 585
R4549 gnd.n730 gnd.n728 585
R4550 gnd.n728 gnd.n717 585
R4551 gnd.n7012 gnd.n7011 585
R4552 gnd.n7013 gnd.n7012 585
R4553 gnd.n729 gnd.n727 585
R4554 gnd.n6878 gnd.n727 585
R4555 gnd.n7006 gnd.n7005 585
R4556 gnd.n7005 gnd.n7004 585
R4557 gnd.n733 gnd.n732 585
R4558 gnd.n988 gnd.n733 585
R4559 gnd.n6838 gnd.n6837 585
R4560 gnd.n6837 gnd.n6836 585
R4561 gnd.n1005 gnd.n1003 585
R4562 gnd.n6785 gnd.n1003 585
R4563 gnd.n6843 gnd.n6842 585
R4564 gnd.n6844 gnd.n6843 585
R4565 gnd.n1004 gnd.n1002 585
R4566 gnd.n6823 gnd.n1002 585
R4567 gnd.n6797 gnd.n6796 585
R4568 gnd.n6796 gnd.n6795 585
R4569 gnd.n1033 gnd.n1031 585
R4570 gnd.n1031 gnd.n1020 585
R4571 gnd.n6802 gnd.n6801 585
R4572 gnd.n6803 gnd.n6802 585
R4573 gnd.n1032 gnd.n1030 585
R4574 gnd.n6657 gnd.n1030 585
R4575 gnd.n1051 gnd.n1049 585
R4576 gnd.n1049 gnd.n1039 585
R4577 gnd.n6755 gnd.n6754 585
R4578 gnd.n6756 gnd.n6755 585
R4579 gnd.n1050 gnd.n1048 585
R4580 gnd.n6672 gnd.n1048 585
R4581 gnd.n6749 gnd.n6748 585
R4582 gnd.n6748 gnd.n6747 585
R4583 gnd.n1054 gnd.n1053 585
R4584 gnd.n6739 gnd.n1054 585
R4585 gnd.n1081 gnd.n1079 585
R4586 gnd.n1079 gnd.n1071 585
R4587 gnd.n6710 gnd.n6709 585
R4588 gnd.n6711 gnd.n6710 585
R4589 gnd.n1080 gnd.n1078 585
R4590 gnd.n1102 gnd.n1078 585
R4591 gnd.n6704 gnd.n6703 585
R4592 gnd.n6703 gnd.n6702 585
R4593 gnd.n1084 gnd.n1083 585
R4594 gnd.n6640 gnd.n1084 585
R4595 gnd.n6589 gnd.n6588 585
R4596 gnd.n6588 gnd.n1093 585
R4597 gnd.n6592 gnd.n6587 585
R4598 gnd.n6587 gnd.n1112 585
R4599 gnd.n6593 gnd.n6586 585
R4600 gnd.n6586 gnd.n1117 585
R4601 gnd.n6594 gnd.n6585 585
R4602 gnd.n6585 gnd.n1125 585
R4603 gnd.n1137 gnd.n1135 585
R4604 gnd.n1135 gnd.n1122 585
R4605 gnd.n6599 gnd.n6598 585
R4606 gnd.n6600 gnd.n6599 585
R4607 gnd.n1136 gnd.n1134 585
R4608 gnd.n6560 gnd.n1134 585
R4609 gnd.n6581 gnd.n6580 585
R4610 gnd.n6580 gnd.n6579 585
R4611 gnd.n1140 gnd.n1139 585
R4612 gnd.n6538 gnd.n1140 585
R4613 gnd.n1172 gnd.n1170 585
R4614 gnd.n1170 gnd.n1160 585
R4615 gnd.n6521 gnd.n6520 585
R4616 gnd.n6522 gnd.n6521 585
R4617 gnd.n1171 gnd.n1169 585
R4618 gnd.n6323 gnd.n1169 585
R4619 gnd.n6515 gnd.n6514 585
R4620 gnd.n6514 gnd.n6513 585
R4621 gnd.n1175 gnd.n1174 585
R4622 gnd.n6505 gnd.n1175 585
R4623 gnd.n6463 gnd.n6462 585
R4624 gnd.n6464 gnd.n6463 585
R4625 gnd.n1202 gnd.n1201 585
R4626 gnd.n1201 gnd.n1191 585
R4627 gnd.n6458 gnd.n6457 585
R4628 gnd.n6457 gnd.n1196 585
R4629 gnd.n6456 gnd.n1204 585
R4630 gnd.n6456 gnd.n6455 585
R4631 gnd.n1227 gnd.n1205 585
R4632 gnd.n6445 gnd.n1205 585
R4633 gnd.n6435 gnd.n6434 585
R4634 gnd.n6436 gnd.n6435 585
R4635 gnd.n1226 gnd.n1225 585
R4636 gnd.n6344 gnd.n1225 585
R4637 gnd.n6429 gnd.n6428 585
R4638 gnd.n6428 gnd.n6427 585
R4639 gnd.n1230 gnd.n1229 585
R4640 gnd.n1238 gnd.n1230 585
R4641 gnd.n1258 gnd.n1256 585
R4642 gnd.n1256 gnd.n1247 585
R4643 gnd.n6399 gnd.n6398 585
R4644 gnd.n6400 gnd.n6399 585
R4645 gnd.n1257 gnd.n1255 585
R4646 gnd.n1255 gnd.n1251 585
R4647 gnd.n6393 gnd.n6392 585
R4648 gnd.n6392 gnd.n6391 585
R4649 gnd.n1261 gnd.n1260 585
R4650 gnd.n1272 gnd.n1261 585
R4651 gnd.n6280 gnd.n6279 585
R4652 gnd.n6279 gnd.n1270 585
R4653 gnd.n6281 gnd.n6278 585
R4654 gnd.n6278 gnd.n1277 585
R4655 gnd.n1304 gnd.n1302 585
R4656 gnd.n6256 gnd.n1302 585
R4657 gnd.n6286 gnd.n6285 585
R4658 gnd.n6287 gnd.n6286 585
R4659 gnd.n1303 gnd.n1301 585
R4660 gnd.n6244 gnd.n1301 585
R4661 gnd.n6274 gnd.n6273 585
R4662 gnd.n6273 gnd.n6272 585
R4663 gnd.n1307 gnd.n1306 585
R4664 gnd.n6217 gnd.n1307 585
R4665 gnd.n6234 gnd.n6233 585
R4666 gnd.n6235 gnd.n6234 585
R4667 gnd.n1337 gnd.n1336 585
R4668 gnd.n6208 gnd.n1336 585
R4669 gnd.n6229 gnd.n6228 585
R4670 gnd.n6228 gnd.n6227 585
R4671 gnd.n1340 gnd.n1339 585
R4672 gnd.n1358 gnd.n1340 585
R4673 gnd.n6183 gnd.n6182 585
R4674 gnd.n6184 gnd.n6183 585
R4675 gnd.n1368 gnd.n1367 585
R4676 gnd.n6152 gnd.n1367 585
R4677 gnd.n6178 gnd.n6177 585
R4678 gnd.n6177 gnd.n6176 585
R4679 gnd.n1371 gnd.n1370 585
R4680 gnd.n6160 gnd.n1371 585
R4681 gnd.n6138 gnd.n6137 585
R4682 gnd.n6139 gnd.n6138 585
R4683 gnd.n1395 gnd.n1394 585
R4684 gnd.n1415 gnd.n1394 585
R4685 gnd.n6133 gnd.n6132 585
R4686 gnd.n6132 gnd.n6131 585
R4687 gnd.n1398 gnd.n1397 585
R4688 gnd.n1409 gnd.n1398 585
R4689 gnd.n6088 gnd.n6087 585
R4690 gnd.n6089 gnd.n6088 585
R4691 gnd.n1423 gnd.n1422 585
R4692 gnd.n6046 gnd.n1422 585
R4693 gnd.n6083 gnd.n6082 585
R4694 gnd.n6082 gnd.n6081 585
R4695 gnd.n1426 gnd.n1425 585
R4696 gnd.n1436 gnd.n1426 585
R4697 gnd.n6029 gnd.n6028 585
R4698 gnd.n6030 gnd.n6029 585
R4699 gnd.n1454 gnd.n1453 585
R4700 gnd.n1453 gnd.n1441 585
R4701 gnd.n6024 gnd.n6023 585
R4702 gnd.n6023 gnd.n6022 585
R4703 gnd.n1457 gnd.n1456 585
R4704 gnd.n6011 gnd.n1457 585
R4705 gnd.n5561 gnd.n5560 585
R4706 gnd.n5560 gnd.n1465 585
R4707 gnd.n5562 gnd.n5559 585
R4708 gnd.n5559 gnd.n5558 585
R4709 gnd.n5467 gnd.n5465 585
R4710 gnd.n5477 gnd.n5467 585
R4711 gnd.n5566 gnd.n5464 585
R4712 gnd.n5543 gnd.n5464 585
R4713 gnd.n5567 gnd.n5463 585
R4714 gnd.n5531 gnd.n5463 585
R4715 gnd.n5568 gnd.n5462 585
R4716 gnd.n5530 gnd.n5462 585
R4717 gnd.n5491 gnd.n5460 585
R4718 gnd.n5492 gnd.n5491 585
R4719 gnd.n5572 gnd.n5459 585
R4720 gnd.n5522 gnd.n5459 585
R4721 gnd.n5573 gnd.n5458 585
R4722 gnd.n5512 gnd.n5458 585
R4723 gnd.n5574 gnd.n5457 585
R4724 gnd.n5511 gnd.n5457 585
R4725 gnd.n5454 gnd.n5452 585
R4726 gnd.n5500 gnd.n5452 585
R4727 gnd.n5579 gnd.n5578 585
R4728 gnd.n5580 gnd.n5579 585
R4729 gnd.n5453 gnd.n1705 585
R4730 gnd.n5449 gnd.n1705 585
R4731 gnd.n5734 gnd.n5733 585
R4732 gnd.n5732 gnd.n1704 585
R4733 gnd.n1707 gnd.n1703 585
R4734 gnd.n5736 gnd.n1703 585
R4735 gnd.n5728 gnd.n1709 585
R4736 gnd.n5727 gnd.n1710 585
R4737 gnd.n5726 gnd.n1711 585
R4738 gnd.n5723 gnd.n1712 585
R4739 gnd.n5722 gnd.n1713 585
R4740 gnd.n5602 gnd.n1714 585
R4741 gnd.n5604 gnd.n5603 585
R4742 gnd.n5714 gnd.n5605 585
R4743 gnd.n5713 gnd.n5606 585
R4744 gnd.n5616 gnd.n5607 585
R4745 gnd.n5706 gnd.n5617 585
R4746 gnd.n5705 gnd.n5618 585
R4747 gnd.n5620 gnd.n5619 585
R4748 gnd.n5698 gnd.n5628 585
R4749 gnd.n5697 gnd.n5629 585
R4750 gnd.n5639 gnd.n5630 585
R4751 gnd.n5690 gnd.n5640 585
R4752 gnd.n5689 gnd.n5641 585
R4753 gnd.n5643 gnd.n5642 585
R4754 gnd.n5682 gnd.n5651 585
R4755 gnd.n5681 gnd.n5652 585
R4756 gnd.n5672 gnd.n5653 585
R4757 gnd.n5674 gnd.n5673 585
R4758 gnd.n1700 gnd.n1685 585
R4759 gnd.n5740 gnd.n1686 585
R4760 gnd.n5739 gnd.n5738 585
R4761 gnd.n7187 gnd.n7186 585
R4762 gnd.n7186 gnd.n7185 585
R4763 gnd.n583 gnd.n582 585
R4764 gnd.n7079 gnd.n583 585
R4765 gnd.n7050 gnd.n678 585
R4766 gnd.n7078 gnd.n678 585
R4767 gnd.n7051 gnd.n7049 585
R4768 gnd.n7049 gnd.n686 585
R4769 gnd.n695 gnd.n685 585
R4770 gnd.n7070 gnd.n685 585
R4771 gnd.n7056 gnd.n7055 585
R4772 gnd.n7057 gnd.n7056 585
R4773 gnd.n694 gnd.n693 585
R4774 gnd.n693 gnd.n692 585
R4775 gnd.n7045 gnd.n7044 585
R4776 gnd.n7044 gnd.n7043 585
R4777 gnd.n698 gnd.n697 585
R4778 gnd.n710 gnd.n698 585
R4779 gnd.n720 gnd.n709 585
R4780 gnd.n7034 gnd.n709 585
R4781 gnd.n7021 gnd.n7020 585
R4782 gnd.n7022 gnd.n7021 585
R4783 gnd.n719 gnd.n718 585
R4784 gnd.n718 gnd.n717 585
R4785 gnd.n7015 gnd.n7014 585
R4786 gnd.n7014 gnd.n7013 585
R4787 gnd.n723 gnd.n722 585
R4788 gnd.n6878 gnd.n723 585
R4789 gnd.n6829 gnd.n735 585
R4790 gnd.n7004 gnd.n735 585
R4791 gnd.n1010 gnd.n1008 585
R4792 gnd.n1008 gnd.n988 585
R4793 gnd.n6834 gnd.n6833 585
R4794 gnd.n6836 gnd.n6834 585
R4795 gnd.n1009 gnd.n1007 585
R4796 gnd.n6785 gnd.n1007 585
R4797 gnd.n6826 gnd.n1000 585
R4798 gnd.n6844 gnd.n1000 585
R4799 gnd.n6825 gnd.n6824 585
R4800 gnd.n6824 gnd.n6823 585
R4801 gnd.n1013 gnd.n1012 585
R4802 gnd.n6795 gnd.n1013 585
R4803 gnd.n6660 gnd.n6659 585
R4804 gnd.n6659 gnd.n1020 585
R4805 gnd.n6664 gnd.n1028 585
R4806 gnd.n6803 gnd.n1028 585
R4807 gnd.n6665 gnd.n6658 585
R4808 gnd.n6658 gnd.n6657 585
R4809 gnd.n6666 gnd.n6654 585
R4810 gnd.n6654 gnd.n1039 585
R4811 gnd.n1100 gnd.n1046 585
R4812 gnd.n6756 gnd.n1046 585
R4813 gnd.n6671 gnd.n6670 585
R4814 gnd.n6672 gnd.n6671 585
R4815 gnd.n1099 gnd.n1056 585
R4816 gnd.n6747 gnd.n1056 585
R4817 gnd.n6650 gnd.n1063 585
R4818 gnd.n6739 gnd.n1063 585
R4819 gnd.n6649 gnd.n6648 585
R4820 gnd.n6648 gnd.n1071 585
R4821 gnd.n6647 gnd.n1077 585
R4822 gnd.n6711 gnd.n1077 585
R4823 gnd.n1104 gnd.n1103 585
R4824 gnd.n1103 gnd.n1102 585
R4825 gnd.n6643 gnd.n1086 585
R4826 gnd.n6702 gnd.n1086 585
R4827 gnd.n6642 gnd.n6641 585
R4828 gnd.n6641 gnd.n6640 585
R4829 gnd.n1107 gnd.n1106 585
R4830 gnd.n1107 gnd.n1093 585
R4831 gnd.n6548 gnd.n6547 585
R4832 gnd.n6547 gnd.n1112 585
R4833 gnd.n6552 gnd.n6546 585
R4834 gnd.n6546 gnd.n1117 585
R4835 gnd.n6553 gnd.n6545 585
R4836 gnd.n6545 gnd.n1125 585
R4837 gnd.n6554 gnd.n6544 585
R4838 gnd.n6544 gnd.n1122 585
R4839 gnd.n1152 gnd.n1133 585
R4840 gnd.n6600 gnd.n1133 585
R4841 gnd.n6559 gnd.n6558 585
R4842 gnd.n6560 gnd.n6559 585
R4843 gnd.n1151 gnd.n1142 585
R4844 gnd.n6579 gnd.n1142 585
R4845 gnd.n6540 gnd.n6539 585
R4846 gnd.n6539 gnd.n6538 585
R4847 gnd.n1155 gnd.n1154 585
R4848 gnd.n1160 gnd.n1155 585
R4849 gnd.n6326 gnd.n1167 585
R4850 gnd.n6522 gnd.n1167 585
R4851 gnd.n6325 gnd.n6324 585
R4852 gnd.n6324 gnd.n6323 585
R4853 gnd.n6330 gnd.n1177 585
R4854 gnd.n6513 gnd.n1177 585
R4855 gnd.n6331 gnd.n1184 585
R4856 gnd.n6505 gnd.n1184 585
R4857 gnd.n6332 gnd.n1200 585
R4858 gnd.n6464 gnd.n1200 585
R4859 gnd.n6313 gnd.n6312 585
R4860 gnd.n6312 gnd.n1191 585
R4861 gnd.n6336 gnd.n6311 585
R4862 gnd.n6311 gnd.n1196 585
R4863 gnd.n6337 gnd.n1207 585
R4864 gnd.n6455 gnd.n1207 585
R4865 gnd.n6338 gnd.n1215 585
R4866 gnd.n6445 gnd.n1215 585
R4867 gnd.n1289 gnd.n1224 585
R4868 gnd.n6436 gnd.n1224 585
R4869 gnd.n6343 gnd.n6342 585
R4870 gnd.n6344 gnd.n6343 585
R4871 gnd.n1288 gnd.n1232 585
R4872 gnd.n6427 gnd.n1232 585
R4873 gnd.n6307 gnd.n6306 585
R4874 gnd.n6306 gnd.n1238 585
R4875 gnd.n6305 gnd.n6304 585
R4876 gnd.n6305 gnd.n1247 585
R4877 gnd.n6303 gnd.n1253 585
R4878 gnd.n6400 gnd.n1253 585
R4879 gnd.n1292 gnd.n1291 585
R4880 gnd.n1291 gnd.n1251 585
R4881 gnd.n6299 gnd.n1263 585
R4882 gnd.n6391 gnd.n1263 585
R4883 gnd.n6298 gnd.n6297 585
R4884 gnd.n6297 gnd.n1272 585
R4885 gnd.n6296 gnd.n1294 585
R4886 gnd.n6296 gnd.n1270 585
R4887 gnd.n6295 gnd.n6294 585
R4888 gnd.n6295 gnd.n1277 585
R4889 gnd.n1296 gnd.n1295 585
R4890 gnd.n6256 gnd.n1295 585
R4891 gnd.n6289 gnd.n6288 585
R4892 gnd.n6288 gnd.n6287 585
R4893 gnd.n1299 gnd.n1298 585
R4894 gnd.n6244 gnd.n1299 585
R4895 gnd.n1352 gnd.n1309 585
R4896 gnd.n6272 gnd.n1309 585
R4897 gnd.n6216 gnd.n6215 585
R4898 gnd.n6217 gnd.n6216 585
R4899 gnd.n1351 gnd.n1334 585
R4900 gnd.n6235 gnd.n1334 585
R4901 gnd.n6210 gnd.n6209 585
R4902 gnd.n6209 gnd.n6208 585
R4903 gnd.n1354 gnd.n1341 585
R4904 gnd.n6227 gnd.n1341 585
R4905 gnd.n6146 gnd.n6145 585
R4906 gnd.n6145 gnd.n1358 585
R4907 gnd.n1389 gnd.n1365 585
R4908 gnd.n6184 gnd.n1365 585
R4909 gnd.n6151 gnd.n6150 585
R4910 gnd.n6152 gnd.n6151 585
R4911 gnd.n1388 gnd.n1373 585
R4912 gnd.n6176 gnd.n1373 585
R4913 gnd.n6142 gnd.n1381 585
R4914 gnd.n6160 gnd.n1381 585
R4915 gnd.n6141 gnd.n6140 585
R4916 gnd.n6140 gnd.n6139 585
R4917 gnd.n1392 gnd.n1391 585
R4918 gnd.n1415 gnd.n1392 585
R4919 gnd.n6039 gnd.n1400 585
R4920 gnd.n6131 gnd.n1400 585
R4921 gnd.n6040 gnd.n6038 585
R4922 gnd.n6038 gnd.n1409 585
R4923 gnd.n1448 gnd.n1421 585
R4924 gnd.n6089 gnd.n1421 585
R4925 gnd.n6045 gnd.n6044 585
R4926 gnd.n6046 gnd.n6045 585
R4927 gnd.n1447 gnd.n1428 585
R4928 gnd.n6081 gnd.n1428 585
R4929 gnd.n6033 gnd.n6032 585
R4930 gnd.n6032 gnd.n1436 585
R4931 gnd.n6031 gnd.n1450 585
R4932 gnd.n6031 gnd.n6030 585
R4933 gnd.n5550 gnd.n1451 585
R4934 gnd.n1451 gnd.n1441 585
R4935 gnd.n5551 gnd.n1459 585
R4936 gnd.n6022 gnd.n1459 585
R4937 gnd.n5552 gnd.n1466 585
R4938 gnd.n6011 gnd.n1466 585
R4939 gnd.n5472 gnd.n5470 585
R4940 gnd.n5470 gnd.n1465 585
R4941 gnd.n5557 gnd.n5556 585
R4942 gnd.n5558 gnd.n5557 585
R4943 gnd.n5471 gnd.n5469 585
R4944 gnd.n5477 gnd.n5469 585
R4945 gnd.n5545 gnd.n5544 585
R4946 gnd.n5544 gnd.n5543 585
R4947 gnd.n5475 gnd.n5474 585
R4948 gnd.n5531 gnd.n5475 585
R4949 gnd.n5529 gnd.n5528 585
R4950 gnd.n5530 gnd.n5529 585
R4951 gnd.n5485 gnd.n5484 585
R4952 gnd.n5492 gnd.n5484 585
R4953 gnd.n5524 gnd.n5523 585
R4954 gnd.n5523 gnd.n5522 585
R4955 gnd.n5488 gnd.n5487 585
R4956 gnd.n5512 gnd.n5488 585
R4957 gnd.n5510 gnd.n5509 585
R4958 gnd.n5511 gnd.n5510 585
R4959 gnd.n5502 gnd.n5501 585
R4960 gnd.n5501 gnd.n5500 585
R4961 gnd.n5505 gnd.n5450 585
R4962 gnd.n5580 gnd.n5450 585
R4963 gnd.n5504 gnd.n1687 585
R4964 gnd.n5449 gnd.n1687 585
R4965 gnd.n7126 gnd.n7125 585
R4966 gnd.n7125 gnd.n7124 585
R4967 gnd.n7127 gnd.n646 585
R4968 gnd.n665 gnd.n641 585
R4969 gnd.n7134 gnd.n640 585
R4970 gnd.n7135 gnd.n639 585
R4971 gnd.n662 gnd.n631 585
R4972 gnd.n7142 gnd.n630 585
R4973 gnd.n7143 gnd.n629 585
R4974 gnd.n660 gnd.n623 585
R4975 gnd.n7150 gnd.n622 585
R4976 gnd.n7151 gnd.n621 585
R4977 gnd.n657 gnd.n613 585
R4978 gnd.n7158 gnd.n612 585
R4979 gnd.n7159 gnd.n611 585
R4980 gnd.n655 gnd.n603 585
R4981 gnd.n7166 gnd.n602 585
R4982 gnd.n7167 gnd.n601 585
R4983 gnd.n652 gnd.n598 585
R4984 gnd.n7172 gnd.n597 585
R4985 gnd.n7173 gnd.n596 585
R4986 gnd.n7174 gnd.n595 585
R4987 gnd.n649 gnd.n593 585
R4988 gnd.n7178 gnd.n592 585
R4989 gnd.n7179 gnd.n591 585
R4990 gnd.n7180 gnd.n587 585
R4991 gnd.n7190 gnd.n580 585
R4992 gnd.n7191 gnd.n579 585
R4993 gnd.n7196 gnd.n578 585
R4994 gnd.n7197 gnd.n577 585
R4995 gnd.n6997 gnd.n739 506.916
R4996 gnd.n6881 gnd.n6880 506.916
R4997 gnd.n5999 gnd.n1467 506.916
R4998 gnd.n6009 gnd.n1469 506.916
R4999 gnd.n3166 gnd.n3165 417.911
R5000 gnd.n1526 gnd.t178 389.64
R5001 gnd.n962 gnd.t102 389.64
R5002 gnd.n1528 gnd.t106 389.64
R5003 gnd.n781 gnd.t159 389.64
R5004 gnd.n5669 gnd.t124 371.625
R5005 gnd.n569 gnd.t77 371.625
R5006 gnd.n5660 gnd.t120 371.625
R5007 gnd.n792 gnd.t172 371.625
R5008 gnd.n872 gnd.t175 371.625
R5009 gnd.n895 gnd.t128 371.625
R5010 gnd.n312 gnd.t150 371.625
R5011 gnd.n279 gnd.t110 371.625
R5012 gnd.n7642 gnd.t147 371.625
R5013 gnd.n349 gnd.t95 371.625
R5014 gnd.n4832 gnd.t134 371.625
R5015 gnd.n4854 gnd.t137 371.625
R5016 gnd.n4875 gnd.t84 371.625
R5017 gnd.n4893 gnd.t162 371.625
R5018 gnd.n5798 gnd.t140 371.625
R5019 gnd.n1643 gnd.t165 371.625
R5020 gnd.n1610 gnd.t188 371.625
R5021 gnd.n574 gnd.t88 371.625
R5022 gnd.n3794 gnd.t113 323.425
R5023 gnd.n2031 gnd.t143 323.425
R5024 gnd.n4642 gnd.n4616 289.615
R5025 gnd.n4610 gnd.n4584 289.615
R5026 gnd.n4578 gnd.n4552 289.615
R5027 gnd.n4547 gnd.n4521 289.615
R5028 gnd.n4515 gnd.n4489 289.615
R5029 gnd.n4483 gnd.n4457 289.615
R5030 gnd.n4451 gnd.n4425 289.615
R5031 gnd.n4420 gnd.n4394 289.615
R5032 gnd.n3868 gnd.t184 279.217
R5033 gnd.n2057 gnd.t168 279.217
R5034 gnd.n1477 gnd.t155 260.649
R5035 gnd.n752 gnd.t158 260.649
R5036 gnd.n6002 gnd.n6001 256.663
R5037 gnd.n6001 gnd.n1494 256.663
R5038 gnd.n6001 gnd.n1495 256.663
R5039 gnd.n6001 gnd.n1496 256.663
R5040 gnd.n6001 gnd.n1497 256.663
R5041 gnd.n6001 gnd.n1498 256.663
R5042 gnd.n6001 gnd.n1499 256.663
R5043 gnd.n6001 gnd.n1500 256.663
R5044 gnd.n6001 gnd.n1501 256.663
R5045 gnd.n6001 gnd.n1502 256.663
R5046 gnd.n6001 gnd.n1503 256.663
R5047 gnd.n6001 gnd.n1504 256.663
R5048 gnd.n6001 gnd.n1505 256.663
R5049 gnd.n6001 gnd.n1506 256.663
R5050 gnd.n6001 gnd.n1507 256.663
R5051 gnd.n6001 gnd.n1508 256.663
R5052 gnd.n5931 gnd.n5930 256.663
R5053 gnd.n6001 gnd.n1509 256.663
R5054 gnd.n6001 gnd.n1510 256.663
R5055 gnd.n6001 gnd.n1511 256.663
R5056 gnd.n6001 gnd.n1512 256.663
R5057 gnd.n6001 gnd.n1513 256.663
R5058 gnd.n6001 gnd.n1514 256.663
R5059 gnd.n6001 gnd.n1515 256.663
R5060 gnd.n6001 gnd.n1516 256.663
R5061 gnd.n6001 gnd.n1517 256.663
R5062 gnd.n6001 gnd.n1518 256.663
R5063 gnd.n6001 gnd.n1519 256.663
R5064 gnd.n6001 gnd.n1520 256.663
R5065 gnd.n6001 gnd.n1521 256.663
R5066 gnd.n6001 gnd.n1522 256.663
R5067 gnd.n6001 gnd.n1523 256.663
R5068 gnd.n6001 gnd.n1524 256.663
R5069 gnd.n6001 gnd.n6000 256.663
R5070 gnd.n6877 gnd.n726 256.663
R5071 gnd.n6886 gnd.n726 256.663
R5072 gnd.n983 gnd.n726 256.663
R5073 gnd.n6893 gnd.n726 256.663
R5074 gnd.n980 gnd.n726 256.663
R5075 gnd.n6900 gnd.n726 256.663
R5076 gnd.n977 gnd.n726 256.663
R5077 gnd.n6907 gnd.n726 256.663
R5078 gnd.n974 gnd.n726 256.663
R5079 gnd.n6914 gnd.n726 256.663
R5080 gnd.n971 gnd.n726 256.663
R5081 gnd.n6921 gnd.n726 256.663
R5082 gnd.n968 gnd.n726 256.663
R5083 gnd.n6928 gnd.n726 256.663
R5084 gnd.n965 gnd.n726 256.663
R5085 gnd.n6936 gnd.n726 256.663
R5086 gnd.n6940 gnd.n6939 256.663
R5087 gnd.n960 gnd.n726 256.663
R5088 gnd.n6943 gnd.n726 256.663
R5089 gnd.n784 gnd.n726 256.663
R5090 gnd.n6951 gnd.n726 256.663
R5091 gnd.n779 gnd.n726 256.663
R5092 gnd.n6958 gnd.n726 256.663
R5093 gnd.n776 gnd.n726 256.663
R5094 gnd.n6965 gnd.n726 256.663
R5095 gnd.n773 gnd.n726 256.663
R5096 gnd.n6972 gnd.n726 256.663
R5097 gnd.n770 gnd.n726 256.663
R5098 gnd.n6979 gnd.n726 256.663
R5099 gnd.n767 gnd.n726 256.663
R5100 gnd.n6986 gnd.n726 256.663
R5101 gnd.n764 gnd.n726 256.663
R5102 gnd.n6993 gnd.n726 256.663
R5103 gnd.n6996 gnd.n726 256.663
R5104 gnd.n5088 gnd.n4802 242.672
R5105 gnd.n5088 gnd.n4803 242.672
R5106 gnd.n5088 gnd.n4804 242.672
R5107 gnd.n5088 gnd.n4805 242.672
R5108 gnd.n5088 gnd.n4806 242.672
R5109 gnd.n5088 gnd.n4807 242.672
R5110 gnd.n5088 gnd.n4808 242.672
R5111 gnd.n5088 gnd.n4809 242.672
R5112 gnd.n5088 gnd.n4810 242.672
R5113 gnd.n5663 gnd.n1597 242.672
R5114 gnd.n5658 gnd.n1597 242.672
R5115 gnd.n5655 gnd.n1597 242.672
R5116 gnd.n5646 gnd.n1597 242.672
R5117 gnd.n5635 gnd.n1597 242.672
R5118 gnd.n5632 gnd.n1597 242.672
R5119 gnd.n5623 gnd.n1597 242.672
R5120 gnd.n5612 gnd.n1597 242.672
R5121 gnd.n5609 gnd.n1597 242.672
R5122 gnd.n3922 gnd.n3921 242.672
R5123 gnd.n3922 gnd.n3832 242.672
R5124 gnd.n3922 gnd.n3833 242.672
R5125 gnd.n3922 gnd.n3834 242.672
R5126 gnd.n3922 gnd.n3835 242.672
R5127 gnd.n3922 gnd.n3836 242.672
R5128 gnd.n3922 gnd.n3837 242.672
R5129 gnd.n3922 gnd.n3838 242.672
R5130 gnd.n3922 gnd.n3839 242.672
R5131 gnd.n3922 gnd.n3840 242.672
R5132 gnd.n3922 gnd.n3841 242.672
R5133 gnd.n3922 gnd.n3842 242.672
R5134 gnd.n3923 gnd.n3922 242.672
R5135 gnd.n4774 gnd.n2006 242.672
R5136 gnd.n4774 gnd.n2005 242.672
R5137 gnd.n4774 gnd.n2004 242.672
R5138 gnd.n4774 gnd.n2003 242.672
R5139 gnd.n4774 gnd.n2002 242.672
R5140 gnd.n4774 gnd.n2001 242.672
R5141 gnd.n4774 gnd.n2000 242.672
R5142 gnd.n4774 gnd.n1999 242.672
R5143 gnd.n4774 gnd.n1998 242.672
R5144 gnd.n4774 gnd.n1997 242.672
R5145 gnd.n4774 gnd.n1996 242.672
R5146 gnd.n4774 gnd.n1995 242.672
R5147 gnd.n4774 gnd.n1994 242.672
R5148 gnd.n7203 gnd.n558 242.672
R5149 gnd.n7203 gnd.n559 242.672
R5150 gnd.n7203 gnd.n560 242.672
R5151 gnd.n7203 gnd.n561 242.672
R5152 gnd.n7203 gnd.n562 242.672
R5153 gnd.n7203 gnd.n563 242.672
R5154 gnd.n7203 gnd.n564 242.672
R5155 gnd.n7203 gnd.n565 242.672
R5156 gnd.n7203 gnd.n7202 242.672
R5157 gnd.n346 gnd.n211 242.672
R5158 gnd.n7538 gnd.n211 242.672
R5159 gnd.n342 gnd.n211 242.672
R5160 gnd.n7545 gnd.n211 242.672
R5161 gnd.n335 gnd.n211 242.672
R5162 gnd.n7552 gnd.n211 242.672
R5163 gnd.n328 gnd.n211 242.672
R5164 gnd.n7559 gnd.n211 242.672
R5165 gnd.n321 gnd.n211 242.672
R5166 gnd.n4006 gnd.n4005 242.672
R5167 gnd.n4005 gnd.n3744 242.672
R5168 gnd.n4005 gnd.n3745 242.672
R5169 gnd.n4005 gnd.n3746 242.672
R5170 gnd.n4005 gnd.n3747 242.672
R5171 gnd.n4005 gnd.n3748 242.672
R5172 gnd.n4005 gnd.n3749 242.672
R5173 gnd.n4005 gnd.n3750 242.672
R5174 gnd.n4774 gnd.n2007 242.672
R5175 gnd.n4774 gnd.n2008 242.672
R5176 gnd.n4774 gnd.n2009 242.672
R5177 gnd.n4774 gnd.n2010 242.672
R5178 gnd.n4774 gnd.n2011 242.672
R5179 gnd.n4774 gnd.n2012 242.672
R5180 gnd.n4774 gnd.n2013 242.672
R5181 gnd.n4774 gnd.n2014 242.672
R5182 gnd.n5088 gnd.n5087 242.672
R5183 gnd.n5088 gnd.n4775 242.672
R5184 gnd.n5088 gnd.n4776 242.672
R5185 gnd.n5088 gnd.n4777 242.672
R5186 gnd.n5088 gnd.n4778 242.672
R5187 gnd.n5088 gnd.n4779 242.672
R5188 gnd.n5088 gnd.n4780 242.672
R5189 gnd.n5088 gnd.n4781 242.672
R5190 gnd.n5088 gnd.n4782 242.672
R5191 gnd.n5088 gnd.n4783 242.672
R5192 gnd.n5088 gnd.n4784 242.672
R5193 gnd.n5088 gnd.n4785 242.672
R5194 gnd.n5088 gnd.n4786 242.672
R5195 gnd.n5088 gnd.n4787 242.672
R5196 gnd.n5088 gnd.n4788 242.672
R5197 gnd.n5088 gnd.n4789 242.672
R5198 gnd.n5088 gnd.n4790 242.672
R5199 gnd.n5088 gnd.n4791 242.672
R5200 gnd.n5088 gnd.n4792 242.672
R5201 gnd.n5088 gnd.n4793 242.672
R5202 gnd.n5088 gnd.n4794 242.672
R5203 gnd.n5088 gnd.n4795 242.672
R5204 gnd.n5088 gnd.n4796 242.672
R5205 gnd.n5088 gnd.n4797 242.672
R5206 gnd.n5088 gnd.n4798 242.672
R5207 gnd.n5088 gnd.n4799 242.672
R5208 gnd.n5088 gnd.n4800 242.672
R5209 gnd.n5088 gnd.n4801 242.672
R5210 gnd.n5089 gnd.n5088 242.672
R5211 gnd.n5873 gnd.n1597 242.672
R5212 gnd.n1646 gnd.n1597 242.672
R5213 gnd.n5880 gnd.n1597 242.672
R5214 gnd.n1637 gnd.n1597 242.672
R5215 gnd.n5887 gnd.n1597 242.672
R5216 gnd.n1630 gnd.n1597 242.672
R5217 gnd.n5894 gnd.n1597 242.672
R5218 gnd.n1623 gnd.n1597 242.672
R5219 gnd.n5901 gnd.n1597 242.672
R5220 gnd.n5904 gnd.n1597 242.672
R5221 gnd.n1614 gnd.n1597 242.672
R5222 gnd.n5913 gnd.n1597 242.672
R5223 gnd.n1605 gnd.n1597 242.672
R5224 gnd.n5920 gnd.n1597 242.672
R5225 gnd.n5923 gnd.n1597 242.672
R5226 gnd.n1597 gnd.n1596 242.672
R5227 gnd.n5929 gnd.n1591 242.672
R5228 gnd.n5813 gnd.n1597 242.672
R5229 gnd.n5812 gnd.n1597 242.672
R5230 gnd.n5820 gnd.n1597 242.672
R5231 gnd.n5806 gnd.n1597 242.672
R5232 gnd.n5827 gnd.n1597 242.672
R5233 gnd.n5796 gnd.n1597 242.672
R5234 gnd.n5834 gnd.n1597 242.672
R5235 gnd.n5789 gnd.n1597 242.672
R5236 gnd.n5841 gnd.n1597 242.672
R5237 gnd.n5782 gnd.n1597 242.672
R5238 gnd.n5848 gnd.n1597 242.672
R5239 gnd.n5775 gnd.n1597 242.672
R5240 gnd.n5855 gnd.n1597 242.672
R5241 gnd.n7204 gnd.n7203 242.672
R5242 gnd.n7203 gnd.n530 242.672
R5243 gnd.n7203 gnd.n531 242.672
R5244 gnd.n7203 gnd.n532 242.672
R5245 gnd.n7203 gnd.n533 242.672
R5246 gnd.n7203 gnd.n534 242.672
R5247 gnd.n7203 gnd.n535 242.672
R5248 gnd.n7203 gnd.n536 242.672
R5249 gnd.n7203 gnd.n537 242.672
R5250 gnd.n7203 gnd.n538 242.672
R5251 gnd.n7203 gnd.n539 242.672
R5252 gnd.n7203 gnd.n540 242.672
R5253 gnd.n7203 gnd.n541 242.672
R5254 gnd.n959 gnd.n788 242.672
R5255 gnd.n7203 gnd.n542 242.672
R5256 gnd.n7203 gnd.n543 242.672
R5257 gnd.n7203 gnd.n544 242.672
R5258 gnd.n7203 gnd.n545 242.672
R5259 gnd.n7203 gnd.n546 242.672
R5260 gnd.n7203 gnd.n547 242.672
R5261 gnd.n7203 gnd.n548 242.672
R5262 gnd.n7203 gnd.n549 242.672
R5263 gnd.n7203 gnd.n550 242.672
R5264 gnd.n7203 gnd.n551 242.672
R5265 gnd.n7203 gnd.n552 242.672
R5266 gnd.n7203 gnd.n553 242.672
R5267 gnd.n7203 gnd.n554 242.672
R5268 gnd.n7203 gnd.n555 242.672
R5269 gnd.n7203 gnd.n556 242.672
R5270 gnd.n7203 gnd.n557 242.672
R5271 gnd.n7570 gnd.n211 242.672
R5272 gnd.n315 gnd.n211 242.672
R5273 gnd.n7577 gnd.n211 242.672
R5274 gnd.n306 gnd.n211 242.672
R5275 gnd.n7584 gnd.n211 242.672
R5276 gnd.n299 gnd.n211 242.672
R5277 gnd.n7591 gnd.n211 242.672
R5278 gnd.n292 gnd.n211 242.672
R5279 gnd.n7598 gnd.n211 242.672
R5280 gnd.n7601 gnd.n211 242.672
R5281 gnd.n283 gnd.n211 242.672
R5282 gnd.n7610 gnd.n211 242.672
R5283 gnd.n274 gnd.n211 242.672
R5284 gnd.n7617 gnd.n211 242.672
R5285 gnd.n267 gnd.n211 242.672
R5286 gnd.n7624 gnd.n211 242.672
R5287 gnd.n260 gnd.n211 242.672
R5288 gnd.n7631 gnd.n211 242.672
R5289 gnd.n253 gnd.n211 242.672
R5290 gnd.n7638 gnd.n211 242.672
R5291 gnd.n246 gnd.n211 242.672
R5292 gnd.n7648 gnd.n211 242.672
R5293 gnd.n239 gnd.n211 242.672
R5294 gnd.n7655 gnd.n211 242.672
R5295 gnd.n232 gnd.n211 242.672
R5296 gnd.n7662 gnd.n211 242.672
R5297 gnd.n225 gnd.n211 242.672
R5298 gnd.n7669 gnd.n211 242.672
R5299 gnd.n218 gnd.n211 242.672
R5300 gnd.n5736 gnd.n5735 242.672
R5301 gnd.n5736 gnd.n1689 242.672
R5302 gnd.n5736 gnd.n1690 242.672
R5303 gnd.n5736 gnd.n1691 242.672
R5304 gnd.n5736 gnd.n1692 242.672
R5305 gnd.n5736 gnd.n1693 242.672
R5306 gnd.n5736 gnd.n1694 242.672
R5307 gnd.n5736 gnd.n1695 242.672
R5308 gnd.n5736 gnd.n1696 242.672
R5309 gnd.n5736 gnd.n1697 242.672
R5310 gnd.n5736 gnd.n1698 242.672
R5311 gnd.n5736 gnd.n1699 242.672
R5312 gnd.n5736 gnd.n1701 242.672
R5313 gnd.n5737 gnd.n5736 242.672
R5314 gnd.n7124 gnd.n666 242.672
R5315 gnd.n7124 gnd.n664 242.672
R5316 gnd.n7124 gnd.n663 242.672
R5317 gnd.n7124 gnd.n661 242.672
R5318 gnd.n7124 gnd.n659 242.672
R5319 gnd.n7124 gnd.n658 242.672
R5320 gnd.n7124 gnd.n656 242.672
R5321 gnd.n7124 gnd.n654 242.672
R5322 gnd.n7124 gnd.n653 242.672
R5323 gnd.n7124 gnd.n651 242.672
R5324 gnd.n7124 gnd.n650 242.672
R5325 gnd.n7124 gnd.n648 242.672
R5326 gnd.n7124 gnd.n668 242.672
R5327 gnd.n7124 gnd.n667 242.672
R5328 gnd.n215 gnd.n212 240.244
R5329 gnd.n7671 gnd.n7670 240.244
R5330 gnd.n7668 gnd.n219 240.244
R5331 gnd.n7664 gnd.n7663 240.244
R5332 gnd.n7661 gnd.n226 240.244
R5333 gnd.n7657 gnd.n7656 240.244
R5334 gnd.n7654 gnd.n233 240.244
R5335 gnd.n7650 gnd.n7649 240.244
R5336 gnd.n7647 gnd.n240 240.244
R5337 gnd.n7640 gnd.n7639 240.244
R5338 gnd.n7637 gnd.n247 240.244
R5339 gnd.n7633 gnd.n7632 240.244
R5340 gnd.n7630 gnd.n254 240.244
R5341 gnd.n7626 gnd.n7625 240.244
R5342 gnd.n7623 gnd.n261 240.244
R5343 gnd.n7619 gnd.n7618 240.244
R5344 gnd.n7616 gnd.n268 240.244
R5345 gnd.n7612 gnd.n7611 240.244
R5346 gnd.n7609 gnd.n275 240.244
R5347 gnd.n7602 gnd.n284 240.244
R5348 gnd.n7600 gnd.n7599 240.244
R5349 gnd.n7597 gnd.n286 240.244
R5350 gnd.n7593 gnd.n7592 240.244
R5351 gnd.n7590 gnd.n293 240.244
R5352 gnd.n7586 gnd.n7585 240.244
R5353 gnd.n7583 gnd.n300 240.244
R5354 gnd.n7579 gnd.n7578 240.244
R5355 gnd.n7576 gnd.n307 240.244
R5356 gnd.n7572 gnd.n7571 240.244
R5357 gnd.n521 gnd.n514 240.244
R5358 gnd.n7224 gnd.n514 240.244
R5359 gnd.n7224 gnd.n502 240.244
R5360 gnd.n7228 gnd.n502 240.244
R5361 gnd.n7228 gnd.n492 240.244
R5362 gnd.n7232 gnd.n492 240.244
R5363 gnd.n7232 gnd.n484 240.244
R5364 gnd.n484 gnd.n467 240.244
R5365 gnd.n7274 gnd.n467 240.244
R5366 gnd.n7274 gnd.n457 240.244
R5367 gnd.n7278 gnd.n457 240.244
R5368 gnd.n7278 gnd.n450 240.244
R5369 gnd.n450 gnd.n432 240.244
R5370 gnd.n7320 gnd.n432 240.244
R5371 gnd.n7320 gnd.n422 240.244
R5372 gnd.n7326 gnd.n422 240.244
R5373 gnd.n7326 gnd.n415 240.244
R5374 gnd.n415 gnd.n399 240.244
R5375 gnd.n7366 gnd.n399 240.244
R5376 gnd.n7366 gnd.n390 240.244
R5377 gnd.n390 gnd.n382 240.244
R5378 gnd.n7403 gnd.n382 240.244
R5379 gnd.n7403 gnd.n376 240.244
R5380 gnd.n7405 gnd.n376 240.244
R5381 gnd.n7405 gnd.n371 240.244
R5382 gnd.n371 gnd.n365 240.244
R5383 gnd.n7427 gnd.n365 240.244
R5384 gnd.n7427 gnd.n89 240.244
R5385 gnd.n7436 gnd.n89 240.244
R5386 gnd.n7473 gnd.n7436 240.244
R5387 gnd.n7473 gnd.n105 240.244
R5388 gnd.n7476 gnd.n105 240.244
R5389 gnd.n7476 gnd.n116 240.244
R5390 gnd.n7480 gnd.n116 240.244
R5391 gnd.n7480 gnd.n125 240.244
R5392 gnd.n7483 gnd.n125 240.244
R5393 gnd.n7483 gnd.n134 240.244
R5394 gnd.n7487 gnd.n134 240.244
R5395 gnd.n7487 gnd.n144 240.244
R5396 gnd.n7490 gnd.n144 240.244
R5397 gnd.n7490 gnd.n153 240.244
R5398 gnd.n7494 gnd.n153 240.244
R5399 gnd.n7494 gnd.n163 240.244
R5400 gnd.n7513 gnd.n163 240.244
R5401 gnd.n7513 gnd.n172 240.244
R5402 gnd.n7509 gnd.n172 240.244
R5403 gnd.n7509 gnd.n182 240.244
R5404 gnd.n7506 gnd.n182 240.244
R5405 gnd.n7506 gnd.n191 240.244
R5406 gnd.n7503 gnd.n191 240.244
R5407 gnd.n7503 gnd.n201 240.244
R5408 gnd.n7500 gnd.n201 240.244
R5409 gnd.n7500 gnd.n209 240.244
R5410 gnd.n7205 gnd.n528 240.244
R5411 gnd.n804 gnd.n528 240.244
R5412 gnd.n808 gnd.n807 240.244
R5413 gnd.n814 gnd.n813 240.244
R5414 gnd.n818 gnd.n817 240.244
R5415 gnd.n824 gnd.n823 240.244
R5416 gnd.n828 gnd.n827 240.244
R5417 gnd.n834 gnd.n833 240.244
R5418 gnd.n838 gnd.n837 240.244
R5419 gnd.n844 gnd.n843 240.244
R5420 gnd.n847 gnd.n846 240.244
R5421 gnd.n854 gnd.n853 240.244
R5422 gnd.n857 gnd.n856 240.244
R5423 gnd.n957 gnd.n956 240.244
R5424 gnd.n953 gnd.n952 240.244
R5425 gnd.n949 gnd.n948 240.244
R5426 gnd.n945 gnd.n944 240.244
R5427 gnd.n941 gnd.n940 240.244
R5428 gnd.n937 gnd.n936 240.244
R5429 gnd.n933 gnd.n932 240.244
R5430 gnd.n929 gnd.n928 240.244
R5431 gnd.n925 gnd.n924 240.244
R5432 gnd.n921 gnd.n920 240.244
R5433 gnd.n917 gnd.n916 240.244
R5434 gnd.n913 gnd.n912 240.244
R5435 gnd.n909 gnd.n908 240.244
R5436 gnd.n905 gnd.n904 240.244
R5437 gnd.n901 gnd.n900 240.244
R5438 gnd.n7213 gnd.n525 240.244
R5439 gnd.n525 gnd.n500 240.244
R5440 gnd.n7242 gnd.n500 240.244
R5441 gnd.n7242 gnd.n495 240.244
R5442 gnd.n7250 gnd.n495 240.244
R5443 gnd.n7250 gnd.n496 240.244
R5444 gnd.n496 gnd.n465 240.244
R5445 gnd.n7288 gnd.n465 240.244
R5446 gnd.n7288 gnd.n460 240.244
R5447 gnd.n7296 gnd.n460 240.244
R5448 gnd.n7296 gnd.n461 240.244
R5449 gnd.n461 gnd.n430 240.244
R5450 gnd.n7335 gnd.n430 240.244
R5451 gnd.n7335 gnd.n425 240.244
R5452 gnd.n7343 gnd.n425 240.244
R5453 gnd.n7343 gnd.n426 240.244
R5454 gnd.n426 gnd.n398 240.244
R5455 gnd.n7379 gnd.n398 240.244
R5456 gnd.n7379 gnd.n393 240.244
R5457 gnd.n7387 gnd.n393 240.244
R5458 gnd.n7387 gnd.n394 240.244
R5459 gnd.n394 gnd.n374 240.244
R5460 gnd.n7412 gnd.n374 240.244
R5461 gnd.n7413 gnd.n7412 240.244
R5462 gnd.n7418 gnd.n7413 240.244
R5463 gnd.n7418 gnd.n7416 240.244
R5464 gnd.n7416 gnd.n92 240.244
R5465 gnd.n7752 gnd.n92 240.244
R5466 gnd.n7752 gnd.n93 240.244
R5467 gnd.n103 gnd.n93 240.244
R5468 gnd.n7746 gnd.n103 240.244
R5469 gnd.n7746 gnd.n104 240.244
R5470 gnd.n7738 gnd.n104 240.244
R5471 gnd.n7738 gnd.n118 240.244
R5472 gnd.n7734 gnd.n118 240.244
R5473 gnd.n7734 gnd.n123 240.244
R5474 gnd.n7726 gnd.n123 240.244
R5475 gnd.n7726 gnd.n137 240.244
R5476 gnd.n7722 gnd.n137 240.244
R5477 gnd.n7722 gnd.n143 240.244
R5478 gnd.n7714 gnd.n143 240.244
R5479 gnd.n7714 gnd.n155 240.244
R5480 gnd.n7710 gnd.n155 240.244
R5481 gnd.n7710 gnd.n161 240.244
R5482 gnd.n7702 gnd.n161 240.244
R5483 gnd.n7702 gnd.n175 240.244
R5484 gnd.n7698 gnd.n175 240.244
R5485 gnd.n7698 gnd.n181 240.244
R5486 gnd.n7690 gnd.n181 240.244
R5487 gnd.n7690 gnd.n194 240.244
R5488 gnd.n7686 gnd.n194 240.244
R5489 gnd.n7686 gnd.n200 240.244
R5490 gnd.n7678 gnd.n200 240.244
R5491 gnd.n5857 gnd.n5856 240.244
R5492 gnd.n5854 gnd.n5770 240.244
R5493 gnd.n5850 gnd.n5849 240.244
R5494 gnd.n5847 gnd.n5776 240.244
R5495 gnd.n5843 gnd.n5842 240.244
R5496 gnd.n5840 gnd.n5783 240.244
R5497 gnd.n5836 gnd.n5835 240.244
R5498 gnd.n5833 gnd.n5790 240.244
R5499 gnd.n5829 gnd.n5828 240.244
R5500 gnd.n5826 gnd.n5797 240.244
R5501 gnd.n5822 gnd.n5821 240.244
R5502 gnd.n5819 gnd.n5807 240.244
R5503 gnd.n5815 gnd.n5814 240.244
R5504 gnd.n5924 gnd.n1595 240.244
R5505 gnd.n5922 gnd.n5921 240.244
R5506 gnd.n5919 gnd.n1599 240.244
R5507 gnd.n5915 gnd.n5914 240.244
R5508 gnd.n5912 gnd.n1606 240.244
R5509 gnd.n5905 gnd.n1615 240.244
R5510 gnd.n5903 gnd.n5902 240.244
R5511 gnd.n5900 gnd.n1617 240.244
R5512 gnd.n5896 gnd.n5895 240.244
R5513 gnd.n5893 gnd.n1624 240.244
R5514 gnd.n5889 gnd.n5888 240.244
R5515 gnd.n5886 gnd.n1631 240.244
R5516 gnd.n5882 gnd.n5881 240.244
R5517 gnd.n5879 gnd.n1638 240.244
R5518 gnd.n5875 gnd.n5874 240.244
R5519 gnd.n5091 gnd.n1980 240.244
R5520 gnd.n1980 gnd.n1970 240.244
R5521 gnd.n5107 gnd.n1970 240.244
R5522 gnd.n5108 gnd.n5107 240.244
R5523 gnd.n5108 gnd.n1961 240.244
R5524 gnd.n1961 gnd.n1952 240.244
R5525 gnd.n5127 gnd.n1952 240.244
R5526 gnd.n5128 gnd.n5127 240.244
R5527 gnd.n5128 gnd.n1944 240.244
R5528 gnd.n1944 gnd.n1934 240.244
R5529 gnd.n5147 gnd.n1934 240.244
R5530 gnd.n5148 gnd.n5147 240.244
R5531 gnd.n5148 gnd.n1924 240.244
R5532 gnd.n5151 gnd.n1924 240.244
R5533 gnd.n5151 gnd.n1915 240.244
R5534 gnd.n1915 gnd.n1908 240.244
R5535 gnd.n5183 gnd.n1908 240.244
R5536 gnd.n5183 gnd.n1898 240.244
R5537 gnd.n5186 gnd.n1898 240.244
R5538 gnd.n5186 gnd.n1890 240.244
R5539 gnd.n1890 gnd.n1883 240.244
R5540 gnd.n5227 gnd.n1883 240.244
R5541 gnd.n5227 gnd.n1875 240.244
R5542 gnd.n1875 gnd.n1869 240.244
R5543 gnd.n5243 gnd.n1869 240.244
R5544 gnd.n5244 gnd.n5243 240.244
R5545 gnd.n5244 gnd.n1863 240.244
R5546 gnd.n1863 gnd.n1857 240.244
R5547 gnd.n1857 gnd.n1849 240.244
R5548 gnd.n5271 gnd.n1849 240.244
R5549 gnd.n5271 gnd.n1837 240.244
R5550 gnd.n5275 gnd.n1837 240.244
R5551 gnd.n5275 gnd.n1822 240.244
R5552 gnd.n5284 gnd.n1822 240.244
R5553 gnd.n5284 gnd.n1814 240.244
R5554 gnd.n1814 gnd.n1796 240.244
R5555 gnd.n5280 gnd.n1796 240.244
R5556 gnd.n5280 gnd.n1787 240.244
R5557 gnd.n1787 gnd.n1778 240.244
R5558 gnd.n5353 gnd.n1778 240.244
R5559 gnd.n5353 gnd.n1761 240.244
R5560 gnd.n5358 gnd.n1761 240.244
R5561 gnd.n5358 gnd.n1752 240.244
R5562 gnd.n1752 gnd.n1743 240.244
R5563 gnd.n5404 gnd.n1743 240.244
R5564 gnd.n5404 gnd.n1734 240.244
R5565 gnd.n5407 gnd.n1734 240.244
R5566 gnd.n5407 gnd.n1673 240.244
R5567 gnd.n5753 gnd.n1673 240.244
R5568 gnd.n5753 gnd.n1665 240.244
R5569 gnd.n1665 gnd.n1653 240.244
R5570 gnd.n5865 gnd.n1653 240.244
R5571 gnd.n5865 gnd.n1647 240.244
R5572 gnd.n4813 gnd.n4812 240.244
R5573 gnd.n5081 gnd.n4812 240.244
R5574 gnd.n5079 gnd.n5078 240.244
R5575 gnd.n5075 gnd.n5074 240.244
R5576 gnd.n5071 gnd.n5070 240.244
R5577 gnd.n5067 gnd.n5066 240.244
R5578 gnd.n5063 gnd.n5062 240.244
R5579 gnd.n5059 gnd.n5058 240.244
R5580 gnd.n5055 gnd.n5054 240.244
R5581 gnd.n5050 gnd.n5049 240.244
R5582 gnd.n5046 gnd.n5045 240.244
R5583 gnd.n5042 gnd.n5041 240.244
R5584 gnd.n5038 gnd.n5037 240.244
R5585 gnd.n5034 gnd.n5033 240.244
R5586 gnd.n5030 gnd.n5029 240.244
R5587 gnd.n5026 gnd.n5025 240.244
R5588 gnd.n5022 gnd.n5021 240.244
R5589 gnd.n5018 gnd.n5017 240.244
R5590 gnd.n5014 gnd.n5013 240.244
R5591 gnd.n5010 gnd.n5009 240.244
R5592 gnd.n5006 gnd.n5005 240.244
R5593 gnd.n5002 gnd.n5001 240.244
R5594 gnd.n4998 gnd.n4997 240.244
R5595 gnd.n4994 gnd.n4993 240.244
R5596 gnd.n4990 gnd.n4989 240.244
R5597 gnd.n4986 gnd.n4985 240.244
R5598 gnd.n4982 gnd.n4981 240.244
R5599 gnd.n4978 gnd.n4977 240.244
R5600 gnd.n4974 gnd.n1991 240.244
R5601 gnd.n5099 gnd.n1978 240.244
R5602 gnd.n5099 gnd.n1974 240.244
R5603 gnd.n5105 gnd.n1974 240.244
R5604 gnd.n5105 gnd.n1959 240.244
R5605 gnd.n5119 gnd.n1959 240.244
R5606 gnd.n5119 gnd.n1955 240.244
R5607 gnd.n5125 gnd.n1955 240.244
R5608 gnd.n5125 gnd.n1942 240.244
R5609 gnd.n5139 gnd.n1942 240.244
R5610 gnd.n5139 gnd.n1938 240.244
R5611 gnd.n5145 gnd.n1938 240.244
R5612 gnd.n5145 gnd.n1922 240.244
R5613 gnd.n5163 gnd.n1922 240.244
R5614 gnd.n5163 gnd.n1917 240.244
R5615 gnd.n5171 gnd.n1917 240.244
R5616 gnd.n5171 gnd.n1918 240.244
R5617 gnd.n1918 gnd.n1897 240.244
R5618 gnd.n5198 gnd.n1897 240.244
R5619 gnd.n5198 gnd.n1892 240.244
R5620 gnd.n5206 gnd.n1892 240.244
R5621 gnd.n5206 gnd.n1893 240.244
R5622 gnd.n1893 gnd.n1873 240.244
R5623 gnd.n5238 gnd.n1873 240.244
R5624 gnd.n5239 gnd.n5238 240.244
R5625 gnd.n5241 gnd.n5239 240.244
R5626 gnd.n5241 gnd.n1859 240.244
R5627 gnd.n5256 gnd.n1859 240.244
R5628 gnd.n5260 gnd.n5256 240.244
R5629 gnd.n5260 gnd.n5257 240.244
R5630 gnd.n5257 gnd.n1836 240.244
R5631 gnd.n5294 gnd.n1836 240.244
R5632 gnd.n5294 gnd.n1825 240.244
R5633 gnd.n5302 gnd.n1825 240.244
R5634 gnd.n5302 gnd.n1826 240.244
R5635 gnd.n1826 gnd.n1794 240.244
R5636 gnd.n5334 gnd.n1794 240.244
R5637 gnd.n5334 gnd.n1789 240.244
R5638 gnd.n5342 gnd.n1789 240.244
R5639 gnd.n5342 gnd.n1790 240.244
R5640 gnd.n1790 gnd.n1759 240.244
R5641 gnd.n5382 gnd.n1759 240.244
R5642 gnd.n5382 gnd.n1754 240.244
R5643 gnd.n5390 gnd.n1754 240.244
R5644 gnd.n5390 gnd.n1755 240.244
R5645 gnd.n1755 gnd.n1732 240.244
R5646 gnd.n5416 gnd.n1732 240.244
R5647 gnd.n5416 gnd.n1728 240.244
R5648 gnd.n5422 gnd.n1728 240.244
R5649 gnd.n5422 gnd.n1663 240.244
R5650 gnd.n5763 gnd.n1663 240.244
R5651 gnd.n5763 gnd.n1658 240.244
R5652 gnd.n5863 gnd.n1658 240.244
R5653 gnd.n5863 gnd.n1659 240.244
R5654 gnd.n4773 gnd.n2016 240.244
R5655 gnd.n4766 gnd.n4765 240.244
R5656 gnd.n4763 gnd.n4762 240.244
R5657 gnd.n4759 gnd.n4758 240.244
R5658 gnd.n4755 gnd.n4754 240.244
R5659 gnd.n4751 gnd.n4750 240.244
R5660 gnd.n4747 gnd.n4746 240.244
R5661 gnd.n4743 gnd.n4742 240.244
R5662 gnd.n4017 gnd.n3729 240.244
R5663 gnd.n4027 gnd.n3729 240.244
R5664 gnd.n4027 gnd.n3720 240.244
R5665 gnd.n3720 gnd.n3709 240.244
R5666 gnd.n4048 gnd.n3709 240.244
R5667 gnd.n4048 gnd.n3703 240.244
R5668 gnd.n4058 gnd.n3703 240.244
R5669 gnd.n4058 gnd.n3692 240.244
R5670 gnd.n3692 gnd.n3684 240.244
R5671 gnd.n4076 gnd.n3684 240.244
R5672 gnd.n4077 gnd.n4076 240.244
R5673 gnd.n4077 gnd.n3669 240.244
R5674 gnd.n4079 gnd.n3669 240.244
R5675 gnd.n4079 gnd.n3655 240.244
R5676 gnd.n4121 gnd.n3655 240.244
R5677 gnd.n4122 gnd.n4121 240.244
R5678 gnd.n4125 gnd.n4122 240.244
R5679 gnd.n4125 gnd.n3610 240.244
R5680 gnd.n3650 gnd.n3610 240.244
R5681 gnd.n3650 gnd.n3620 240.244
R5682 gnd.n4135 gnd.n3620 240.244
R5683 gnd.n4135 gnd.n3641 240.244
R5684 gnd.n4145 gnd.n3641 240.244
R5685 gnd.n4145 gnd.n3523 240.244
R5686 gnd.n4190 gnd.n3523 240.244
R5687 gnd.n4190 gnd.n3509 240.244
R5688 gnd.n4212 gnd.n3509 240.244
R5689 gnd.n4213 gnd.n4212 240.244
R5690 gnd.n4213 gnd.n3496 240.244
R5691 gnd.n3496 gnd.n3485 240.244
R5692 gnd.n4244 gnd.n3485 240.244
R5693 gnd.n4245 gnd.n4244 240.244
R5694 gnd.n4246 gnd.n4245 240.244
R5695 gnd.n4246 gnd.n3470 240.244
R5696 gnd.n3470 gnd.n3469 240.244
R5697 gnd.n3469 gnd.n3454 240.244
R5698 gnd.n4297 gnd.n3454 240.244
R5699 gnd.n4298 gnd.n4297 240.244
R5700 gnd.n4298 gnd.n3441 240.244
R5701 gnd.n3441 gnd.n3430 240.244
R5702 gnd.n4329 gnd.n3430 240.244
R5703 gnd.n4330 gnd.n4329 240.244
R5704 gnd.n4331 gnd.n4330 240.244
R5705 gnd.n4331 gnd.n3414 240.244
R5706 gnd.n3414 gnd.n3413 240.244
R5707 gnd.n3413 gnd.n3400 240.244
R5708 gnd.n4386 gnd.n3400 240.244
R5709 gnd.n4387 gnd.n4386 240.244
R5710 gnd.n4387 gnd.n3387 240.244
R5711 gnd.n3387 gnd.n2072 240.244
R5712 gnd.n4674 gnd.n2072 240.244
R5713 gnd.n4677 gnd.n4674 240.244
R5714 gnd.n4677 gnd.n4676 240.244
R5715 gnd.n4007 gnd.n3742 240.244
R5716 gnd.n3763 gnd.n3742 240.244
R5717 gnd.n3766 gnd.n3765 240.244
R5718 gnd.n3773 gnd.n3772 240.244
R5719 gnd.n3776 gnd.n3775 240.244
R5720 gnd.n3783 gnd.n3782 240.244
R5721 gnd.n3786 gnd.n3785 240.244
R5722 gnd.n3793 gnd.n3792 240.244
R5723 gnd.n4015 gnd.n3739 240.244
R5724 gnd.n3739 gnd.n3718 240.244
R5725 gnd.n4038 gnd.n3718 240.244
R5726 gnd.n4038 gnd.n3712 240.244
R5727 gnd.n4046 gnd.n3712 240.244
R5728 gnd.n4046 gnd.n3714 240.244
R5729 gnd.n3714 gnd.n3690 240.244
R5730 gnd.n4068 gnd.n3690 240.244
R5731 gnd.n4068 gnd.n3686 240.244
R5732 gnd.n4074 gnd.n3686 240.244
R5733 gnd.n4074 gnd.n3668 240.244
R5734 gnd.n4099 gnd.n3668 240.244
R5735 gnd.n4099 gnd.n3663 240.244
R5736 gnd.n4111 gnd.n3663 240.244
R5737 gnd.n4111 gnd.n3664 240.244
R5738 gnd.n4107 gnd.n3664 240.244
R5739 gnd.n4107 gnd.n3612 240.244
R5740 gnd.n4159 gnd.n3612 240.244
R5741 gnd.n4159 gnd.n3613 240.244
R5742 gnd.n4155 gnd.n3613 240.244
R5743 gnd.n4155 gnd.n3619 240.244
R5744 gnd.n3639 gnd.n3619 240.244
R5745 gnd.n3639 gnd.n3521 240.244
R5746 gnd.n4194 gnd.n3521 240.244
R5747 gnd.n4194 gnd.n3516 240.244
R5748 gnd.n4202 gnd.n3516 240.244
R5749 gnd.n4202 gnd.n3517 240.244
R5750 gnd.n3517 gnd.n3494 240.244
R5751 gnd.n4234 gnd.n3494 240.244
R5752 gnd.n4234 gnd.n3489 240.244
R5753 gnd.n4242 gnd.n3489 240.244
R5754 gnd.n4242 gnd.n3490 240.244
R5755 gnd.n3490 gnd.n3467 240.244
R5756 gnd.n4279 gnd.n3467 240.244
R5757 gnd.n4279 gnd.n3462 240.244
R5758 gnd.n4287 gnd.n3462 240.244
R5759 gnd.n4287 gnd.n3463 240.244
R5760 gnd.n3463 gnd.n3439 240.244
R5761 gnd.n4319 gnd.n3439 240.244
R5762 gnd.n4319 gnd.n3434 240.244
R5763 gnd.n4327 gnd.n3434 240.244
R5764 gnd.n4327 gnd.n3435 240.244
R5765 gnd.n3435 gnd.n3412 240.244
R5766 gnd.n4368 gnd.n3412 240.244
R5767 gnd.n4368 gnd.n3407 240.244
R5768 gnd.n4376 gnd.n3407 240.244
R5769 gnd.n4376 gnd.n3408 240.244
R5770 gnd.n3408 gnd.n3385 240.244
R5771 gnd.n4662 gnd.n3385 240.244
R5772 gnd.n4662 gnd.n3380 240.244
R5773 gnd.n4672 gnd.n3380 240.244
R5774 gnd.n4672 gnd.n3381 240.244
R5775 gnd.n3381 gnd.n2015 240.244
R5776 gnd.n318 gnd.n207 240.244
R5777 gnd.n7561 gnd.n7560 240.244
R5778 gnd.n7558 gnd.n322 240.244
R5779 gnd.n7554 gnd.n7553 240.244
R5780 gnd.n7551 gnd.n329 240.244
R5781 gnd.n7547 gnd.n7546 240.244
R5782 gnd.n7544 gnd.n336 240.244
R5783 gnd.n7540 gnd.n7539 240.244
R5784 gnd.n7537 gnd.n343 240.244
R5785 gnd.n7215 gnd.n515 240.244
R5786 gnd.n7222 gnd.n515 240.244
R5787 gnd.n7222 gnd.n503 240.244
R5788 gnd.n503 gnd.n490 240.244
R5789 gnd.n7252 gnd.n490 240.244
R5790 gnd.n7252 gnd.n485 240.244
R5791 gnd.n7259 gnd.n485 240.244
R5792 gnd.n7259 gnd.n468 240.244
R5793 gnd.n468 gnd.n456 240.244
R5794 gnd.n7298 gnd.n456 240.244
R5795 gnd.n7298 gnd.n451 240.244
R5796 gnd.n7305 gnd.n451 240.244
R5797 gnd.n7305 gnd.n433 240.244
R5798 gnd.n433 gnd.n421 240.244
R5799 gnd.n7345 gnd.n421 240.244
R5800 gnd.n7345 gnd.n416 240.244
R5801 gnd.n7352 gnd.n416 240.244
R5802 gnd.n7352 gnd.n400 240.244
R5803 gnd.n400 gnd.n389 240.244
R5804 gnd.n7389 gnd.n389 240.244
R5805 gnd.n7389 gnd.n384 240.244
R5806 gnd.n7401 gnd.n384 240.244
R5807 gnd.n7401 gnd.n377 240.244
R5808 gnd.n7394 gnd.n377 240.244
R5809 gnd.n7394 gnd.n373 240.244
R5810 gnd.n373 gnd.n372 240.244
R5811 gnd.n372 gnd.n86 240.244
R5812 gnd.n7754 gnd.n86 240.244
R5813 gnd.n7754 gnd.n88 240.244
R5814 gnd.n7471 gnd.n88 240.244
R5815 gnd.n7471 gnd.n106 240.244
R5816 gnd.n7467 gnd.n106 240.244
R5817 gnd.n7467 gnd.n117 240.244
R5818 gnd.n7464 gnd.n117 240.244
R5819 gnd.n7464 gnd.n126 240.244
R5820 gnd.n7461 gnd.n126 240.244
R5821 gnd.n7461 gnd.n135 240.244
R5822 gnd.n7458 gnd.n135 240.244
R5823 gnd.n7458 gnd.n145 240.244
R5824 gnd.n7455 gnd.n145 240.244
R5825 gnd.n7455 gnd.n154 240.244
R5826 gnd.n7452 gnd.n154 240.244
R5827 gnd.n7452 gnd.n164 240.244
R5828 gnd.n7515 gnd.n164 240.244
R5829 gnd.n7515 gnd.n173 240.244
R5830 gnd.n355 gnd.n173 240.244
R5831 gnd.n355 gnd.n183 240.244
R5832 gnd.n7522 gnd.n183 240.244
R5833 gnd.n7522 gnd.n192 240.244
R5834 gnd.n352 gnd.n192 240.244
R5835 gnd.n352 gnd.n202 240.244
R5836 gnd.n7529 gnd.n202 240.244
R5837 gnd.n7529 gnd.n210 240.244
R5838 gnd.n608 gnd.n607 240.244
R5839 gnd.n616 gnd.n615 240.244
R5840 gnd.n618 gnd.n617 240.244
R5841 gnd.n626 gnd.n625 240.244
R5842 gnd.n634 gnd.n633 240.244
R5843 gnd.n636 gnd.n635 240.244
R5844 gnd.n644 gnd.n643 240.244
R5845 gnd.n7201 gnd.n567 240.244
R5846 gnd.n566 gnd.n519 240.244
R5847 gnd.n7096 gnd.n523 240.244
R5848 gnd.n7096 gnd.n505 240.244
R5849 gnd.n7240 gnd.n505 240.244
R5850 gnd.n7240 gnd.n506 240.244
R5851 gnd.n506 gnd.n494 240.244
R5852 gnd.n7235 gnd.n494 240.244
R5853 gnd.n7235 gnd.n470 240.244
R5854 gnd.n7286 gnd.n470 240.244
R5855 gnd.n7286 gnd.n471 240.244
R5856 gnd.n471 gnd.n459 240.244
R5857 gnd.n7281 gnd.n459 240.244
R5858 gnd.n7281 gnd.n435 240.244
R5859 gnd.n7333 gnd.n435 240.244
R5860 gnd.n7333 gnd.n436 240.244
R5861 gnd.n436 gnd.n424 240.244
R5862 gnd.n7328 gnd.n424 240.244
R5863 gnd.n7328 gnd.n402 240.244
R5864 gnd.n7377 gnd.n402 240.244
R5865 gnd.n7377 gnd.n403 240.244
R5866 gnd.n403 gnd.n392 240.244
R5867 gnd.n7372 gnd.n392 240.244
R5868 gnd.n7372 gnd.n378 240.244
R5869 gnd.n7410 gnd.n378 240.244
R5870 gnd.n7410 gnd.n369 240.244
R5871 gnd.n7420 gnd.n369 240.244
R5872 gnd.n7420 gnd.n363 240.244
R5873 gnd.n7429 gnd.n363 240.244
R5874 gnd.n7429 gnd.n91 240.244
R5875 gnd.n7432 gnd.n91 240.244
R5876 gnd.n7432 gnd.n108 240.244
R5877 gnd.n7744 gnd.n108 240.244
R5878 gnd.n7744 gnd.n109 240.244
R5879 gnd.n7740 gnd.n109 240.244
R5880 gnd.n7740 gnd.n115 240.244
R5881 gnd.n7732 gnd.n115 240.244
R5882 gnd.n7732 gnd.n127 240.244
R5883 gnd.n7728 gnd.n127 240.244
R5884 gnd.n7728 gnd.n132 240.244
R5885 gnd.n7720 gnd.n132 240.244
R5886 gnd.n7720 gnd.n147 240.244
R5887 gnd.n7716 gnd.n147 240.244
R5888 gnd.n7716 gnd.n152 240.244
R5889 gnd.n7708 gnd.n152 240.244
R5890 gnd.n7708 gnd.n165 240.244
R5891 gnd.n7704 gnd.n165 240.244
R5892 gnd.n7704 gnd.n170 240.244
R5893 gnd.n7696 gnd.n170 240.244
R5894 gnd.n7696 gnd.n185 240.244
R5895 gnd.n7692 gnd.n185 240.244
R5896 gnd.n7692 gnd.n190 240.244
R5897 gnd.n7684 gnd.n190 240.244
R5898 gnd.n7684 gnd.n203 240.244
R5899 gnd.n7680 gnd.n203 240.244
R5900 gnd.n2035 gnd.n1993 240.244
R5901 gnd.n4733 gnd.n4732 240.244
R5902 gnd.n4729 gnd.n4728 240.244
R5903 gnd.n4725 gnd.n4724 240.244
R5904 gnd.n4721 gnd.n4720 240.244
R5905 gnd.n4717 gnd.n4716 240.244
R5906 gnd.n4713 gnd.n4712 240.244
R5907 gnd.n4709 gnd.n4708 240.244
R5908 gnd.n4705 gnd.n4704 240.244
R5909 gnd.n4701 gnd.n4700 240.244
R5910 gnd.n4697 gnd.n4696 240.244
R5911 gnd.n4693 gnd.n4692 240.244
R5912 gnd.n4689 gnd.n4688 240.244
R5913 gnd.n3930 gnd.n3827 240.244
R5914 gnd.n3930 gnd.n3820 240.244
R5915 gnd.n3941 gnd.n3820 240.244
R5916 gnd.n3941 gnd.n3816 240.244
R5917 gnd.n3947 gnd.n3816 240.244
R5918 gnd.n3947 gnd.n3808 240.244
R5919 gnd.n3957 gnd.n3808 240.244
R5920 gnd.n3957 gnd.n3803 240.244
R5921 gnd.n3993 gnd.n3803 240.244
R5922 gnd.n3993 gnd.n3804 240.244
R5923 gnd.n3804 gnd.n3751 240.244
R5924 gnd.n3988 gnd.n3751 240.244
R5925 gnd.n3988 gnd.n3987 240.244
R5926 gnd.n3987 gnd.n3730 240.244
R5927 gnd.n3983 gnd.n3730 240.244
R5928 gnd.n3983 gnd.n3721 240.244
R5929 gnd.n3980 gnd.n3721 240.244
R5930 gnd.n3980 gnd.n3979 240.244
R5931 gnd.n3979 gnd.n3704 240.244
R5932 gnd.n3975 gnd.n3704 240.244
R5933 gnd.n3975 gnd.n3693 240.244
R5934 gnd.n3693 gnd.n3674 240.244
R5935 gnd.n4088 gnd.n3674 240.244
R5936 gnd.n4088 gnd.n3670 240.244
R5937 gnd.n4096 gnd.n3670 240.244
R5938 gnd.n4096 gnd.n3661 240.244
R5939 gnd.n3661 gnd.n3597 240.244
R5940 gnd.n4168 gnd.n3597 240.244
R5941 gnd.n4168 gnd.n3598 240.244
R5942 gnd.n3609 gnd.n3598 240.244
R5943 gnd.n3644 gnd.n3609 240.244
R5944 gnd.n3647 gnd.n3644 240.244
R5945 gnd.n3647 gnd.n3621 240.244
R5946 gnd.n3634 gnd.n3621 240.244
R5947 gnd.n3634 gnd.n3631 240.244
R5948 gnd.n3631 gnd.n3524 240.244
R5949 gnd.n4189 gnd.n3524 240.244
R5950 gnd.n4189 gnd.n3514 240.244
R5951 gnd.n4185 gnd.n3514 240.244
R5952 gnd.n4185 gnd.n3508 240.244
R5953 gnd.n4182 gnd.n3508 240.244
R5954 gnd.n4182 gnd.n3497 240.244
R5955 gnd.n4179 gnd.n3497 240.244
R5956 gnd.n4179 gnd.n3475 240.244
R5957 gnd.n4255 gnd.n3475 240.244
R5958 gnd.n4255 gnd.n3471 240.244
R5959 gnd.n4276 gnd.n3471 240.244
R5960 gnd.n4276 gnd.n3460 240.244
R5961 gnd.n4272 gnd.n3460 240.244
R5962 gnd.n4272 gnd.n3453 240.244
R5963 gnd.n4269 gnd.n3453 240.244
R5964 gnd.n4269 gnd.n3442 240.244
R5965 gnd.n4266 gnd.n3442 240.244
R5966 gnd.n4266 gnd.n3419 240.244
R5967 gnd.n4340 gnd.n3419 240.244
R5968 gnd.n4340 gnd.n3415 240.244
R5969 gnd.n4365 gnd.n3415 240.244
R5970 gnd.n4365 gnd.n3406 240.244
R5971 gnd.n4361 gnd.n3406 240.244
R5972 gnd.n4361 gnd.n3399 240.244
R5973 gnd.n4357 gnd.n3399 240.244
R5974 gnd.n4357 gnd.n3388 240.244
R5975 gnd.n4354 gnd.n3388 240.244
R5976 gnd.n4354 gnd.n2064 240.244
R5977 gnd.n4684 gnd.n2064 240.244
R5978 gnd.n3844 gnd.n3843 240.244
R5979 gnd.n3915 gnd.n3843 240.244
R5980 gnd.n3913 gnd.n3912 240.244
R5981 gnd.n3909 gnd.n3908 240.244
R5982 gnd.n3905 gnd.n3904 240.244
R5983 gnd.n3901 gnd.n3900 240.244
R5984 gnd.n3897 gnd.n3896 240.244
R5985 gnd.n3893 gnd.n3892 240.244
R5986 gnd.n3889 gnd.n3888 240.244
R5987 gnd.n3885 gnd.n3884 240.244
R5988 gnd.n3881 gnd.n3880 240.244
R5989 gnd.n3877 gnd.n3876 240.244
R5990 gnd.n3873 gnd.n3831 240.244
R5991 gnd.n3933 gnd.n3825 240.244
R5992 gnd.n3933 gnd.n3821 240.244
R5993 gnd.n3939 gnd.n3821 240.244
R5994 gnd.n3939 gnd.n3814 240.244
R5995 gnd.n3949 gnd.n3814 240.244
R5996 gnd.n3949 gnd.n3810 240.244
R5997 gnd.n3955 gnd.n3810 240.244
R5998 gnd.n3955 gnd.n3801 240.244
R5999 gnd.n3995 gnd.n3801 240.244
R6000 gnd.n3995 gnd.n3752 240.244
R6001 gnd.n4003 gnd.n3752 240.244
R6002 gnd.n4003 gnd.n3753 240.244
R6003 gnd.n3753 gnd.n3731 240.244
R6004 gnd.n4024 gnd.n3731 240.244
R6005 gnd.n4024 gnd.n3723 240.244
R6006 gnd.n4035 gnd.n3723 240.244
R6007 gnd.n4035 gnd.n3724 240.244
R6008 gnd.n3724 gnd.n3705 240.244
R6009 gnd.n4055 gnd.n3705 240.244
R6010 gnd.n4055 gnd.n3695 240.244
R6011 gnd.n4065 gnd.n3695 240.244
R6012 gnd.n4065 gnd.n3676 240.244
R6013 gnd.n4086 gnd.n3676 240.244
R6014 gnd.n4086 gnd.n3678 240.244
R6015 gnd.n3678 gnd.n3659 240.244
R6016 gnd.n4114 gnd.n3659 240.244
R6017 gnd.n4114 gnd.n3601 240.244
R6018 gnd.n4166 gnd.n3601 240.244
R6019 gnd.n4166 gnd.n3602 240.244
R6020 gnd.n4162 gnd.n3602 240.244
R6021 gnd.n4162 gnd.n3608 240.244
R6022 gnd.n3623 gnd.n3608 240.244
R6023 gnd.n4152 gnd.n3623 240.244
R6024 gnd.n4152 gnd.n3624 240.244
R6025 gnd.n4148 gnd.n3624 240.244
R6026 gnd.n4148 gnd.n3630 240.244
R6027 gnd.n3630 gnd.n3513 240.244
R6028 gnd.n4205 gnd.n3513 240.244
R6029 gnd.n4205 gnd.n3506 240.244
R6030 gnd.n4216 gnd.n3506 240.244
R6031 gnd.n4216 gnd.n3499 240.244
R6032 gnd.n4231 gnd.n3499 240.244
R6033 gnd.n4231 gnd.n3500 240.244
R6034 gnd.n3500 gnd.n3478 240.244
R6035 gnd.n4253 gnd.n3478 240.244
R6036 gnd.n4253 gnd.n3479 240.244
R6037 gnd.n3479 gnd.n3458 240.244
R6038 gnd.n4290 gnd.n3458 240.244
R6039 gnd.n4290 gnd.n3451 240.244
R6040 gnd.n4301 gnd.n3451 240.244
R6041 gnd.n4301 gnd.n3444 240.244
R6042 gnd.n4316 gnd.n3444 240.244
R6043 gnd.n4316 gnd.n3445 240.244
R6044 gnd.n3445 gnd.n3422 240.244
R6045 gnd.n4338 gnd.n3422 240.244
R6046 gnd.n4338 gnd.n3424 240.244
R6047 gnd.n3424 gnd.n3404 240.244
R6048 gnd.n4379 gnd.n3404 240.244
R6049 gnd.n4379 gnd.n3397 240.244
R6050 gnd.n4390 gnd.n3397 240.244
R6051 gnd.n4390 gnd.n3390 240.244
R6052 gnd.n4659 gnd.n3390 240.244
R6053 gnd.n4659 gnd.n3391 240.244
R6054 gnd.n3391 gnd.n2067 240.244
R6055 gnd.n4682 gnd.n2067 240.244
R6056 gnd.n5599 gnd.n5598 240.244
R6057 gnd.n5611 gnd.n5610 240.244
R6058 gnd.n5622 gnd.n5613 240.244
R6059 gnd.n5625 gnd.n5624 240.244
R6060 gnd.n5634 gnd.n5633 240.244
R6061 gnd.n5645 gnd.n5636 240.244
R6062 gnd.n5648 gnd.n5647 240.244
R6063 gnd.n5657 gnd.n5656 240.244
R6064 gnd.n5662 gnd.n5659 240.244
R6065 gnd.n4928 gnd.n1981 240.244
R6066 gnd.n4925 gnd.n1981 240.244
R6067 gnd.n4925 gnd.n1972 240.244
R6068 gnd.n4922 gnd.n1972 240.244
R6069 gnd.n4922 gnd.n1962 240.244
R6070 gnd.n4919 gnd.n1962 240.244
R6071 gnd.n4919 gnd.n1953 240.244
R6072 gnd.n4916 gnd.n1953 240.244
R6073 gnd.n4916 gnd.n1945 240.244
R6074 gnd.n4913 gnd.n1945 240.244
R6075 gnd.n4913 gnd.n1936 240.244
R6076 gnd.n4910 gnd.n1936 240.244
R6077 gnd.n4910 gnd.n1925 240.244
R6078 gnd.n1925 gnd.n1914 240.244
R6079 gnd.n5173 gnd.n1914 240.244
R6080 gnd.n5173 gnd.n1910 240.244
R6081 gnd.n5181 gnd.n1910 240.244
R6082 gnd.n5181 gnd.n1899 240.244
R6083 gnd.n1899 gnd.n1889 240.244
R6084 gnd.n5208 gnd.n1889 240.244
R6085 gnd.n5208 gnd.n1885 240.244
R6086 gnd.n5225 gnd.n1885 240.244
R6087 gnd.n5225 gnd.n1876 240.244
R6088 gnd.n5221 gnd.n1876 240.244
R6089 gnd.n5221 gnd.n1871 240.244
R6090 gnd.n5218 gnd.n1871 240.244
R6091 gnd.n5218 gnd.n1856 240.244
R6092 gnd.n5262 gnd.n1856 240.244
R6093 gnd.n5262 gnd.n1851 240.244
R6094 gnd.n5269 gnd.n1851 240.244
R6095 gnd.n5269 gnd.n1838 240.244
R6096 gnd.n1838 gnd.n1820 240.244
R6097 gnd.n5304 gnd.n1820 240.244
R6098 gnd.n5304 gnd.n1815 240.244
R6099 gnd.n5311 gnd.n1815 240.244
R6100 gnd.n5311 gnd.n1797 240.244
R6101 gnd.n1797 gnd.n1785 240.244
R6102 gnd.n5344 gnd.n1785 240.244
R6103 gnd.n5344 gnd.n1780 240.244
R6104 gnd.n5351 gnd.n1780 240.244
R6105 gnd.n5351 gnd.n1762 240.244
R6106 gnd.n1762 gnd.n1750 240.244
R6107 gnd.n5392 gnd.n1750 240.244
R6108 gnd.n5392 gnd.n1745 240.244
R6109 gnd.n5402 gnd.n1745 240.244
R6110 gnd.n5402 gnd.n1735 240.244
R6111 gnd.n5396 gnd.n1735 240.244
R6112 gnd.n5396 gnd.n1675 240.244
R6113 gnd.n5751 gnd.n1675 240.244
R6114 gnd.n5751 gnd.n1666 240.244
R6115 gnd.n1681 gnd.n1666 240.244
R6116 gnd.n1681 gnd.n1655 240.244
R6117 gnd.n1682 gnd.n1655 240.244
R6118 gnd.n4965 gnd.n4964 240.244
R6119 gnd.n4961 gnd.n4960 240.244
R6120 gnd.n4957 gnd.n4956 240.244
R6121 gnd.n4953 gnd.n4952 240.244
R6122 gnd.n4949 gnd.n4948 240.244
R6123 gnd.n4945 gnd.n4944 240.244
R6124 gnd.n4941 gnd.n4940 240.244
R6125 gnd.n4937 gnd.n4936 240.244
R6126 gnd.n4892 gnd.n4811 240.244
R6127 gnd.n5097 gnd.n1982 240.244
R6128 gnd.n5097 gnd.n1983 240.244
R6129 gnd.n1983 gnd.n1973 240.244
R6130 gnd.n1973 gnd.n1964 240.244
R6131 gnd.n5117 gnd.n1964 240.244
R6132 gnd.n5117 gnd.n1965 240.244
R6133 gnd.n1965 gnd.n1954 240.244
R6134 gnd.n1954 gnd.n1946 240.244
R6135 gnd.n5137 gnd.n1946 240.244
R6136 gnd.n5137 gnd.n1947 240.244
R6137 gnd.n1947 gnd.n1937 240.244
R6138 gnd.n1937 gnd.n1927 240.244
R6139 gnd.n5161 gnd.n1927 240.244
R6140 gnd.n5161 gnd.n1928 240.244
R6141 gnd.n1928 gnd.n1916 240.244
R6142 gnd.n5156 gnd.n1916 240.244
R6143 gnd.n5156 gnd.n1901 240.244
R6144 gnd.n5196 gnd.n1901 240.244
R6145 gnd.n5196 gnd.n1902 240.244
R6146 gnd.n1902 gnd.n1891 240.244
R6147 gnd.n5191 gnd.n1891 240.244
R6148 gnd.n5191 gnd.n1877 240.244
R6149 gnd.n5236 gnd.n1877 240.244
R6150 gnd.n5236 gnd.n1878 240.244
R6151 gnd.n1878 gnd.n1872 240.244
R6152 gnd.n1872 gnd.n1864 240.244
R6153 gnd.n5254 gnd.n1864 240.244
R6154 gnd.n5254 gnd.n1858 240.244
R6155 gnd.n5250 gnd.n1858 240.244
R6156 gnd.n5250 gnd.n1840 240.244
R6157 gnd.n5292 gnd.n1840 240.244
R6158 gnd.n5292 gnd.n1841 240.244
R6159 gnd.n1841 gnd.n1824 240.244
R6160 gnd.n5287 gnd.n1824 240.244
R6161 gnd.n5287 gnd.n1799 240.244
R6162 gnd.n5332 gnd.n1799 240.244
R6163 gnd.n5332 gnd.n1800 240.244
R6164 gnd.n1800 gnd.n1788 240.244
R6165 gnd.n5327 gnd.n1788 240.244
R6166 gnd.n5327 gnd.n1763 240.244
R6167 gnd.n5380 gnd.n1763 240.244
R6168 gnd.n5380 gnd.n1764 240.244
R6169 gnd.n1764 gnd.n1753 240.244
R6170 gnd.n5375 gnd.n1753 240.244
R6171 gnd.n5375 gnd.n1737 240.244
R6172 gnd.n5414 gnd.n1737 240.244
R6173 gnd.n5414 gnd.n1738 240.244
R6174 gnd.n1738 gnd.n1727 240.244
R6175 gnd.n1727 gnd.n1668 240.244
R6176 gnd.n5761 gnd.n1668 240.244
R6177 gnd.n5761 gnd.n1669 240.244
R6178 gnd.n1669 gnd.n1657 240.244
R6179 gnd.n5597 gnd.n1657 240.244
R6180 gnd.n3164 gnd.n2208 240.244
R6181 gnd.n3158 gnd.n2208 240.244
R6182 gnd.n3158 gnd.n2212 240.244
R6183 gnd.n3154 gnd.n2212 240.244
R6184 gnd.n3154 gnd.n2214 240.244
R6185 gnd.n3150 gnd.n2214 240.244
R6186 gnd.n3150 gnd.n2219 240.244
R6187 gnd.n3146 gnd.n2219 240.244
R6188 gnd.n3146 gnd.n2221 240.244
R6189 gnd.n3142 gnd.n2221 240.244
R6190 gnd.n3142 gnd.n2227 240.244
R6191 gnd.n3138 gnd.n2227 240.244
R6192 gnd.n3138 gnd.n2229 240.244
R6193 gnd.n3134 gnd.n2229 240.244
R6194 gnd.n3134 gnd.n2235 240.244
R6195 gnd.n3130 gnd.n2235 240.244
R6196 gnd.n3130 gnd.n2237 240.244
R6197 gnd.n3126 gnd.n2237 240.244
R6198 gnd.n3126 gnd.n2243 240.244
R6199 gnd.n3122 gnd.n2243 240.244
R6200 gnd.n3122 gnd.n2245 240.244
R6201 gnd.n3118 gnd.n2245 240.244
R6202 gnd.n3118 gnd.n2251 240.244
R6203 gnd.n3114 gnd.n2251 240.244
R6204 gnd.n3114 gnd.n2253 240.244
R6205 gnd.n3110 gnd.n2253 240.244
R6206 gnd.n3110 gnd.n2259 240.244
R6207 gnd.n3106 gnd.n2259 240.244
R6208 gnd.n3106 gnd.n2261 240.244
R6209 gnd.n3102 gnd.n2261 240.244
R6210 gnd.n3102 gnd.n2267 240.244
R6211 gnd.n3098 gnd.n2267 240.244
R6212 gnd.n3098 gnd.n2269 240.244
R6213 gnd.n3094 gnd.n2269 240.244
R6214 gnd.n3094 gnd.n2275 240.244
R6215 gnd.n3090 gnd.n2275 240.244
R6216 gnd.n3090 gnd.n2277 240.244
R6217 gnd.n3086 gnd.n2277 240.244
R6218 gnd.n3086 gnd.n2283 240.244
R6219 gnd.n3082 gnd.n2283 240.244
R6220 gnd.n3082 gnd.n2285 240.244
R6221 gnd.n3078 gnd.n2285 240.244
R6222 gnd.n3078 gnd.n2291 240.244
R6223 gnd.n3074 gnd.n2291 240.244
R6224 gnd.n3074 gnd.n2293 240.244
R6225 gnd.n3070 gnd.n2293 240.244
R6226 gnd.n3070 gnd.n2299 240.244
R6227 gnd.n3066 gnd.n2299 240.244
R6228 gnd.n3066 gnd.n2301 240.244
R6229 gnd.n3062 gnd.n2301 240.244
R6230 gnd.n3062 gnd.n2307 240.244
R6231 gnd.n3058 gnd.n2307 240.244
R6232 gnd.n3058 gnd.n2309 240.244
R6233 gnd.n3054 gnd.n2309 240.244
R6234 gnd.n3054 gnd.n2315 240.244
R6235 gnd.n3050 gnd.n2315 240.244
R6236 gnd.n3050 gnd.n2317 240.244
R6237 gnd.n3046 gnd.n2317 240.244
R6238 gnd.n3046 gnd.n2323 240.244
R6239 gnd.n3042 gnd.n2323 240.244
R6240 gnd.n3042 gnd.n2325 240.244
R6241 gnd.n3038 gnd.n2325 240.244
R6242 gnd.n3038 gnd.n2331 240.244
R6243 gnd.n3034 gnd.n2331 240.244
R6244 gnd.n3034 gnd.n2333 240.244
R6245 gnd.n3030 gnd.n2333 240.244
R6246 gnd.n3030 gnd.n2339 240.244
R6247 gnd.n3026 gnd.n2339 240.244
R6248 gnd.n3026 gnd.n2341 240.244
R6249 gnd.n3022 gnd.n2341 240.244
R6250 gnd.n3022 gnd.n2347 240.244
R6251 gnd.n3018 gnd.n2347 240.244
R6252 gnd.n3018 gnd.n2349 240.244
R6253 gnd.n3014 gnd.n2349 240.244
R6254 gnd.n3014 gnd.n2355 240.244
R6255 gnd.n3010 gnd.n2355 240.244
R6256 gnd.n3010 gnd.n2357 240.244
R6257 gnd.n3006 gnd.n2357 240.244
R6258 gnd.n3006 gnd.n2363 240.244
R6259 gnd.n3002 gnd.n2363 240.244
R6260 gnd.n3002 gnd.n2365 240.244
R6261 gnd.n2998 gnd.n2365 240.244
R6262 gnd.n2998 gnd.n2371 240.244
R6263 gnd.n2994 gnd.n2371 240.244
R6264 gnd.n2994 gnd.n2373 240.244
R6265 gnd.n2990 gnd.n2373 240.244
R6266 gnd.n2990 gnd.n2379 240.244
R6267 gnd.n2986 gnd.n2379 240.244
R6268 gnd.n2986 gnd.n2381 240.244
R6269 gnd.n2982 gnd.n2381 240.244
R6270 gnd.n2982 gnd.n2387 240.244
R6271 gnd.n2978 gnd.n2387 240.244
R6272 gnd.n2978 gnd.n2389 240.244
R6273 gnd.n2974 gnd.n2389 240.244
R6274 gnd.n2974 gnd.n2395 240.244
R6275 gnd.n2970 gnd.n2395 240.244
R6276 gnd.n2970 gnd.n2397 240.244
R6277 gnd.n2966 gnd.n2397 240.244
R6278 gnd.n2966 gnd.n2403 240.244
R6279 gnd.n2962 gnd.n2403 240.244
R6280 gnd.n2962 gnd.n2405 240.244
R6281 gnd.n2958 gnd.n2405 240.244
R6282 gnd.n2958 gnd.n2411 240.244
R6283 gnd.n2954 gnd.n2411 240.244
R6284 gnd.n2954 gnd.n2413 240.244
R6285 gnd.n2950 gnd.n2413 240.244
R6286 gnd.n2950 gnd.n2419 240.244
R6287 gnd.n2946 gnd.n2419 240.244
R6288 gnd.n2946 gnd.n2421 240.244
R6289 gnd.n2942 gnd.n2421 240.244
R6290 gnd.n2942 gnd.n2427 240.244
R6291 gnd.n2938 gnd.n2427 240.244
R6292 gnd.n2938 gnd.n2429 240.244
R6293 gnd.n2934 gnd.n2429 240.244
R6294 gnd.n2934 gnd.n2435 240.244
R6295 gnd.n2930 gnd.n2435 240.244
R6296 gnd.n2930 gnd.n2437 240.244
R6297 gnd.n2926 gnd.n2437 240.244
R6298 gnd.n2926 gnd.n2443 240.244
R6299 gnd.n2922 gnd.n2443 240.244
R6300 gnd.n2922 gnd.n2445 240.244
R6301 gnd.n2918 gnd.n2445 240.244
R6302 gnd.n2918 gnd.n2451 240.244
R6303 gnd.n2914 gnd.n2451 240.244
R6304 gnd.n2914 gnd.n2453 240.244
R6305 gnd.n2910 gnd.n2453 240.244
R6306 gnd.n2910 gnd.n2459 240.244
R6307 gnd.n2906 gnd.n2459 240.244
R6308 gnd.n2906 gnd.n2461 240.244
R6309 gnd.n2902 gnd.n2461 240.244
R6310 gnd.n2902 gnd.n2467 240.244
R6311 gnd.n2898 gnd.n2467 240.244
R6312 gnd.n2898 gnd.n2469 240.244
R6313 gnd.n2894 gnd.n2469 240.244
R6314 gnd.n2894 gnd.n2475 240.244
R6315 gnd.n2890 gnd.n2475 240.244
R6316 gnd.n2890 gnd.n2477 240.244
R6317 gnd.n2886 gnd.n2477 240.244
R6318 gnd.n2886 gnd.n2483 240.244
R6319 gnd.n2882 gnd.n2483 240.244
R6320 gnd.n2882 gnd.n2485 240.244
R6321 gnd.n2878 gnd.n2485 240.244
R6322 gnd.n2878 gnd.n2491 240.244
R6323 gnd.n2874 gnd.n2491 240.244
R6324 gnd.n2874 gnd.n2493 240.244
R6325 gnd.n2870 gnd.n2493 240.244
R6326 gnd.n2870 gnd.n2499 240.244
R6327 gnd.n2866 gnd.n2499 240.244
R6328 gnd.n2866 gnd.n2501 240.244
R6329 gnd.n2862 gnd.n2501 240.244
R6330 gnd.n2862 gnd.n2507 240.244
R6331 gnd.n2858 gnd.n2507 240.244
R6332 gnd.n2858 gnd.n2509 240.244
R6333 gnd.n2854 gnd.n2509 240.244
R6334 gnd.n2850 gnd.n2514 240.244
R6335 gnd.n2850 gnd.n2516 240.244
R6336 gnd.n2844 gnd.n2516 240.244
R6337 gnd.n2844 gnd.n2522 240.244
R6338 gnd.n2840 gnd.n2522 240.244
R6339 gnd.n2840 gnd.n2524 240.244
R6340 gnd.n2836 gnd.n2524 240.244
R6341 gnd.n2836 gnd.n2529 240.244
R6342 gnd.n2832 gnd.n2529 240.244
R6343 gnd.n2832 gnd.n2531 240.244
R6344 gnd.n2828 gnd.n2531 240.244
R6345 gnd.n2828 gnd.n2537 240.244
R6346 gnd.n2824 gnd.n2537 240.244
R6347 gnd.n2824 gnd.n2539 240.244
R6348 gnd.n2820 gnd.n2539 240.244
R6349 gnd.n2820 gnd.n2545 240.244
R6350 gnd.n2816 gnd.n2545 240.244
R6351 gnd.n2816 gnd.n2547 240.244
R6352 gnd.n2812 gnd.n2547 240.244
R6353 gnd.n2812 gnd.n2553 240.244
R6354 gnd.n2808 gnd.n2553 240.244
R6355 gnd.n2808 gnd.n2555 240.244
R6356 gnd.n2804 gnd.n2555 240.244
R6357 gnd.n2804 gnd.n2561 240.244
R6358 gnd.n2800 gnd.n2561 240.244
R6359 gnd.n2800 gnd.n2563 240.244
R6360 gnd.n2796 gnd.n2563 240.244
R6361 gnd.n2796 gnd.n2569 240.244
R6362 gnd.n2792 gnd.n2569 240.244
R6363 gnd.n2792 gnd.n2571 240.244
R6364 gnd.n2788 gnd.n2571 240.244
R6365 gnd.n2788 gnd.n2577 240.244
R6366 gnd.n2784 gnd.n2577 240.244
R6367 gnd.n2784 gnd.n2579 240.244
R6368 gnd.n2780 gnd.n2579 240.244
R6369 gnd.n2780 gnd.n2585 240.244
R6370 gnd.n2776 gnd.n2585 240.244
R6371 gnd.n2776 gnd.n2587 240.244
R6372 gnd.n2772 gnd.n2587 240.244
R6373 gnd.n2772 gnd.n2593 240.244
R6374 gnd.n2768 gnd.n2593 240.244
R6375 gnd.n2768 gnd.n2595 240.244
R6376 gnd.n2764 gnd.n2595 240.244
R6377 gnd.n2764 gnd.n2601 240.244
R6378 gnd.n2760 gnd.n2601 240.244
R6379 gnd.n2760 gnd.n2603 240.244
R6380 gnd.n2756 gnd.n2603 240.244
R6381 gnd.n2756 gnd.n2609 240.244
R6382 gnd.n2752 gnd.n2609 240.244
R6383 gnd.n2752 gnd.n2611 240.244
R6384 gnd.n2748 gnd.n2611 240.244
R6385 gnd.n2748 gnd.n2617 240.244
R6386 gnd.n2744 gnd.n2617 240.244
R6387 gnd.n2744 gnd.n2619 240.244
R6388 gnd.n2740 gnd.n2619 240.244
R6389 gnd.n2740 gnd.n2625 240.244
R6390 gnd.n2736 gnd.n2625 240.244
R6391 gnd.n2736 gnd.n2627 240.244
R6392 gnd.n2732 gnd.n2627 240.244
R6393 gnd.n2732 gnd.n2633 240.244
R6394 gnd.n2728 gnd.n2633 240.244
R6395 gnd.n2728 gnd.n2635 240.244
R6396 gnd.n2724 gnd.n2635 240.244
R6397 gnd.n2724 gnd.n2641 240.244
R6398 gnd.n2720 gnd.n2641 240.244
R6399 gnd.n2720 gnd.n2643 240.244
R6400 gnd.n2716 gnd.n2643 240.244
R6401 gnd.n2716 gnd.n2649 240.244
R6402 gnd.n2712 gnd.n2649 240.244
R6403 gnd.n2712 gnd.n2651 240.244
R6404 gnd.n2708 gnd.n2651 240.244
R6405 gnd.n2708 gnd.n2657 240.244
R6406 gnd.n2704 gnd.n2657 240.244
R6407 gnd.n2704 gnd.n2659 240.244
R6408 gnd.n2700 gnd.n2659 240.244
R6409 gnd.n2700 gnd.n2665 240.244
R6410 gnd.n2696 gnd.n2665 240.244
R6411 gnd.n2696 gnd.n2667 240.244
R6412 gnd.n2692 gnd.n2667 240.244
R6413 gnd.n2692 gnd.n2673 240.244
R6414 gnd.n2688 gnd.n2673 240.244
R6415 gnd.n2688 gnd.n2675 240.244
R6416 gnd.n2684 gnd.n2675 240.244
R6417 gnd.n2684 gnd.n2682 240.244
R6418 gnd.n2081 gnd.n1811 240.244
R6419 gnd.n5314 gnd.n1811 240.244
R6420 gnd.n5315 gnd.n5314 240.244
R6421 gnd.n5316 gnd.n5315 240.244
R6422 gnd.n5316 gnd.n1806 240.244
R6423 gnd.n5324 gnd.n1806 240.244
R6424 gnd.n5324 gnd.n1807 240.244
R6425 gnd.n1807 gnd.n1775 240.244
R6426 gnd.n5361 gnd.n1775 240.244
R6427 gnd.n5361 gnd.n1770 240.244
R6428 gnd.n5372 gnd.n1770 240.244
R6429 gnd.n5372 gnd.n1771 240.244
R6430 gnd.n5368 gnd.n1771 240.244
R6431 gnd.n5368 gnd.n1725 240.244
R6432 gnd.n5425 gnd.n1725 240.244
R6433 gnd.n5425 gnd.n1721 240.244
R6434 gnd.n5431 gnd.n1721 240.244
R6435 gnd.n5432 gnd.n5431 240.244
R6436 gnd.n5433 gnd.n5432 240.244
R6437 gnd.n5433 gnd.n1716 240.244
R6438 gnd.n5594 gnd.n1716 240.244
R6439 gnd.n5594 gnd.n1717 240.244
R6440 gnd.n5590 gnd.n1717 240.244
R6441 gnd.n5590 gnd.n5587 240.244
R6442 gnd.n5587 gnd.n5586 240.244
R6443 gnd.n5586 gnd.n5441 240.244
R6444 gnd.n5582 gnd.n5441 240.244
R6445 gnd.n5582 gnd.n5447 240.244
R6446 gnd.n5498 gnd.n5447 240.244
R6447 gnd.n5514 gnd.n5498 240.244
R6448 gnd.n5514 gnd.n5493 240.244
R6449 gnd.n5520 gnd.n5493 240.244
R6450 gnd.n5520 gnd.n5483 240.244
R6451 gnd.n5533 gnd.n5483 240.244
R6452 gnd.n5533 gnd.n5478 240.244
R6453 gnd.n5541 gnd.n5478 240.244
R6454 gnd.n5541 gnd.n5479 240.244
R6455 gnd.n5479 gnd.n1464 240.244
R6456 gnd.n6013 gnd.n1464 240.244
R6457 gnd.n6013 gnd.n1460 240.244
R6458 gnd.n6019 gnd.n1460 240.244
R6459 gnd.n6019 gnd.n1434 240.244
R6460 gnd.n6073 gnd.n1434 240.244
R6461 gnd.n6073 gnd.n1430 240.244
R6462 gnd.n6079 gnd.n1430 240.244
R6463 gnd.n6079 gnd.n1407 240.244
R6464 gnd.n6115 gnd.n1407 240.244
R6465 gnd.n6115 gnd.n1402 240.244
R6466 gnd.n6129 gnd.n1402 240.244
R6467 gnd.n6129 gnd.n1403 240.244
R6468 gnd.n6125 gnd.n1403 240.244
R6469 gnd.n6125 gnd.n6124 240.244
R6470 gnd.n6124 gnd.n1363 240.244
R6471 gnd.n6186 gnd.n1363 240.244
R6472 gnd.n6186 gnd.n1359 240.244
R6473 gnd.n6192 gnd.n1359 240.244
R6474 gnd.n6192 gnd.n1332 240.244
R6475 gnd.n6237 gnd.n1332 240.244
R6476 gnd.n6237 gnd.n1328 240.244
R6477 gnd.n6243 gnd.n1328 240.244
R6478 gnd.n6247 gnd.n6243 240.244
R6479 gnd.n6248 gnd.n6247 240.244
R6480 gnd.n6248 gnd.n1324 240.244
R6481 gnd.n6254 gnd.n1324 240.244
R6482 gnd.n6254 gnd.n1269 240.244
R6483 gnd.n6383 gnd.n1269 240.244
R6484 gnd.n6383 gnd.n1265 240.244
R6485 gnd.n6389 gnd.n1265 240.244
R6486 gnd.n6389 gnd.n1245 240.244
R6487 gnd.n6410 gnd.n1245 240.244
R6488 gnd.n6410 gnd.n1240 240.244
R6489 gnd.n6418 gnd.n1240 240.244
R6490 gnd.n6418 gnd.n1241 240.244
R6491 gnd.n1241 gnd.n1213 240.244
R6492 gnd.n6447 gnd.n1213 240.244
R6493 gnd.n6447 gnd.n1209 240.244
R6494 gnd.n6453 gnd.n1209 240.244
R6495 gnd.n6453 gnd.n1190 240.244
R6496 gnd.n6481 gnd.n1190 240.244
R6497 gnd.n6481 gnd.n1185 240.244
R6498 gnd.n6503 gnd.n1185 240.244
R6499 gnd.n6503 gnd.n1186 240.244
R6500 gnd.n6499 gnd.n1186 240.244
R6501 gnd.n6499 gnd.n6498 240.244
R6502 gnd.n6498 gnd.n6496 240.244
R6503 gnd.n6496 gnd.n6489 240.244
R6504 gnd.n6489 gnd.n1131 240.244
R6505 gnd.n6602 gnd.n1131 240.244
R6506 gnd.n6602 gnd.n1126 240.244
R6507 gnd.n6615 gnd.n1126 240.244
R6508 gnd.n6615 gnd.n1127 240.244
R6509 gnd.n6611 gnd.n1127 240.244
R6510 gnd.n6611 gnd.n1092 240.244
R6511 gnd.n6694 gnd.n1092 240.244
R6512 gnd.n6694 gnd.n1088 240.244
R6513 gnd.n6700 gnd.n1088 240.244
R6514 gnd.n6700 gnd.n1069 240.244
R6515 gnd.n6722 gnd.n1069 240.244
R6516 gnd.n6722 gnd.n1064 240.244
R6517 gnd.n6737 gnd.n1064 240.244
R6518 gnd.n6737 gnd.n1065 240.244
R6519 gnd.n6733 gnd.n1065 240.244
R6520 gnd.n6733 gnd.n6732 240.244
R6521 gnd.n6732 gnd.n1026 240.244
R6522 gnd.n6805 gnd.n1026 240.244
R6523 gnd.n6805 gnd.n1022 240.244
R6524 gnd.n6811 gnd.n1022 240.244
R6525 gnd.n6811 gnd.n998 240.244
R6526 gnd.n6846 gnd.n998 240.244
R6527 gnd.n6846 gnd.n993 240.244
R6528 gnd.n6864 gnd.n993 240.244
R6529 gnd.n6864 gnd.n994 240.244
R6530 gnd.n6860 gnd.n994 240.244
R6531 gnd.n6860 gnd.n6858 240.244
R6532 gnd.n6858 gnd.n6857 240.244
R6533 gnd.n6857 gnd.n716 240.244
R6534 gnd.n7024 gnd.n716 240.244
R6535 gnd.n7024 gnd.n711 240.244
R6536 gnd.n7032 gnd.n711 240.244
R6537 gnd.n7032 gnd.n712 240.244
R6538 gnd.n712 gnd.n691 240.244
R6539 gnd.n7059 gnd.n691 240.244
R6540 gnd.n7059 gnd.n687 240.244
R6541 gnd.n7068 gnd.n687 240.244
R6542 gnd.n7068 gnd.n675 240.244
R6543 gnd.n7081 gnd.n675 240.244
R6544 gnd.n7082 gnd.n7081 240.244
R6545 gnd.n7083 gnd.n7082 240.244
R6546 gnd.n7083 gnd.n670 240.244
R6547 gnd.n7122 gnd.n670 240.244
R6548 gnd.n7122 gnd.n671 240.244
R6549 gnd.n7118 gnd.n671 240.244
R6550 gnd.n7118 gnd.n7117 240.244
R6551 gnd.n7117 gnd.n7116 240.244
R6552 gnd.n7116 gnd.n7099 240.244
R6553 gnd.n7112 gnd.n7099 240.244
R6554 gnd.n7112 gnd.n7111 240.244
R6555 gnd.n7111 gnd.n7110 240.244
R6556 gnd.n7110 gnd.n482 240.244
R6557 gnd.n7262 gnd.n482 240.244
R6558 gnd.n7263 gnd.n7262 240.244
R6559 gnd.n7263 gnd.n478 240.244
R6560 gnd.n7271 gnd.n478 240.244
R6561 gnd.n7271 gnd.n448 240.244
R6562 gnd.n7308 gnd.n448 240.244
R6563 gnd.n7309 gnd.n7308 240.244
R6564 gnd.n7309 gnd.n443 240.244
R6565 gnd.n7317 gnd.n443 240.244
R6566 gnd.n7317 gnd.n444 240.244
R6567 gnd.n444 gnd.n413 240.244
R6568 gnd.n7355 gnd.n413 240.244
R6569 gnd.n7355 gnd.n408 240.244
R6570 gnd.n7363 gnd.n408 240.244
R6571 gnd.n7363 gnd.n409 240.244
R6572 gnd.n3168 gnd.n2206 240.244
R6573 gnd.n3168 gnd.n2202 240.244
R6574 gnd.n3174 gnd.n2202 240.244
R6575 gnd.n3174 gnd.n2200 240.244
R6576 gnd.n3178 gnd.n2200 240.244
R6577 gnd.n3178 gnd.n2196 240.244
R6578 gnd.n3184 gnd.n2196 240.244
R6579 gnd.n3184 gnd.n2194 240.244
R6580 gnd.n3188 gnd.n2194 240.244
R6581 gnd.n3188 gnd.n2190 240.244
R6582 gnd.n3194 gnd.n2190 240.244
R6583 gnd.n3194 gnd.n2188 240.244
R6584 gnd.n3198 gnd.n2188 240.244
R6585 gnd.n3198 gnd.n2184 240.244
R6586 gnd.n3204 gnd.n2184 240.244
R6587 gnd.n3204 gnd.n2182 240.244
R6588 gnd.n3208 gnd.n2182 240.244
R6589 gnd.n3208 gnd.n2178 240.244
R6590 gnd.n3214 gnd.n2178 240.244
R6591 gnd.n3214 gnd.n2176 240.244
R6592 gnd.n3218 gnd.n2176 240.244
R6593 gnd.n3218 gnd.n2172 240.244
R6594 gnd.n3224 gnd.n2172 240.244
R6595 gnd.n3224 gnd.n2170 240.244
R6596 gnd.n3228 gnd.n2170 240.244
R6597 gnd.n3228 gnd.n2166 240.244
R6598 gnd.n3234 gnd.n2166 240.244
R6599 gnd.n3234 gnd.n2164 240.244
R6600 gnd.n3238 gnd.n2164 240.244
R6601 gnd.n3238 gnd.n2160 240.244
R6602 gnd.n3244 gnd.n2160 240.244
R6603 gnd.n3244 gnd.n2158 240.244
R6604 gnd.n3248 gnd.n2158 240.244
R6605 gnd.n3248 gnd.n2154 240.244
R6606 gnd.n3254 gnd.n2154 240.244
R6607 gnd.n3254 gnd.n2152 240.244
R6608 gnd.n3258 gnd.n2152 240.244
R6609 gnd.n3258 gnd.n2148 240.244
R6610 gnd.n3264 gnd.n2148 240.244
R6611 gnd.n3264 gnd.n2146 240.244
R6612 gnd.n3268 gnd.n2146 240.244
R6613 gnd.n3268 gnd.n2142 240.244
R6614 gnd.n3274 gnd.n2142 240.244
R6615 gnd.n3274 gnd.n2140 240.244
R6616 gnd.n3278 gnd.n2140 240.244
R6617 gnd.n3278 gnd.n2136 240.244
R6618 gnd.n3284 gnd.n2136 240.244
R6619 gnd.n3284 gnd.n2134 240.244
R6620 gnd.n3288 gnd.n2134 240.244
R6621 gnd.n3288 gnd.n2130 240.244
R6622 gnd.n3294 gnd.n2130 240.244
R6623 gnd.n3294 gnd.n2128 240.244
R6624 gnd.n3298 gnd.n2128 240.244
R6625 gnd.n3298 gnd.n2124 240.244
R6626 gnd.n3304 gnd.n2124 240.244
R6627 gnd.n3304 gnd.n2122 240.244
R6628 gnd.n3308 gnd.n2122 240.244
R6629 gnd.n3308 gnd.n2118 240.244
R6630 gnd.n3314 gnd.n2118 240.244
R6631 gnd.n3314 gnd.n2116 240.244
R6632 gnd.n3318 gnd.n2116 240.244
R6633 gnd.n3318 gnd.n2112 240.244
R6634 gnd.n3324 gnd.n2112 240.244
R6635 gnd.n3324 gnd.n2110 240.244
R6636 gnd.n3328 gnd.n2110 240.244
R6637 gnd.n3328 gnd.n2106 240.244
R6638 gnd.n3334 gnd.n2106 240.244
R6639 gnd.n3334 gnd.n2104 240.244
R6640 gnd.n3338 gnd.n2104 240.244
R6641 gnd.n3338 gnd.n2100 240.244
R6642 gnd.n3344 gnd.n2100 240.244
R6643 gnd.n3344 gnd.n2098 240.244
R6644 gnd.n3348 gnd.n2098 240.244
R6645 gnd.n3348 gnd.n2094 240.244
R6646 gnd.n3354 gnd.n2094 240.244
R6647 gnd.n3354 gnd.n2092 240.244
R6648 gnd.n3358 gnd.n2092 240.244
R6649 gnd.n3358 gnd.n2088 240.244
R6650 gnd.n3364 gnd.n2088 240.244
R6651 gnd.n3364 gnd.n2086 240.244
R6652 gnd.n3368 gnd.n2086 240.244
R6653 gnd.n3368 gnd.n2075 240.244
R6654 gnd.n3376 gnd.n2075 240.244
R6655 gnd.n3376 gnd.n2082 240.244
R6656 gnd.n5579 gnd.n1705 240.244
R6657 gnd.n5579 gnd.n5452 240.244
R6658 gnd.n5457 gnd.n5452 240.244
R6659 gnd.n5458 gnd.n5457 240.244
R6660 gnd.n5459 gnd.n5458 240.244
R6661 gnd.n5491 gnd.n5459 240.244
R6662 gnd.n5491 gnd.n5462 240.244
R6663 gnd.n5463 gnd.n5462 240.244
R6664 gnd.n5464 gnd.n5463 240.244
R6665 gnd.n5467 gnd.n5464 240.244
R6666 gnd.n5559 gnd.n5467 240.244
R6667 gnd.n5560 gnd.n5559 240.244
R6668 gnd.n5560 gnd.n1457 240.244
R6669 gnd.n6023 gnd.n1457 240.244
R6670 gnd.n6023 gnd.n1453 240.244
R6671 gnd.n6029 gnd.n1453 240.244
R6672 gnd.n6029 gnd.n1426 240.244
R6673 gnd.n6082 gnd.n1426 240.244
R6674 gnd.n6082 gnd.n1422 240.244
R6675 gnd.n6088 gnd.n1422 240.244
R6676 gnd.n6088 gnd.n1398 240.244
R6677 gnd.n6132 gnd.n1398 240.244
R6678 gnd.n6132 gnd.n1394 240.244
R6679 gnd.n6138 gnd.n1394 240.244
R6680 gnd.n6138 gnd.n1371 240.244
R6681 gnd.n6177 gnd.n1371 240.244
R6682 gnd.n6177 gnd.n1367 240.244
R6683 gnd.n6183 gnd.n1367 240.244
R6684 gnd.n6183 gnd.n1340 240.244
R6685 gnd.n6228 gnd.n1340 240.244
R6686 gnd.n6228 gnd.n1336 240.244
R6687 gnd.n6234 gnd.n1336 240.244
R6688 gnd.n6234 gnd.n1307 240.244
R6689 gnd.n6273 gnd.n1307 240.244
R6690 gnd.n6273 gnd.n1301 240.244
R6691 gnd.n6286 gnd.n1301 240.244
R6692 gnd.n6286 gnd.n1302 240.244
R6693 gnd.n6278 gnd.n1302 240.244
R6694 gnd.n6279 gnd.n6278 240.244
R6695 gnd.n6279 gnd.n1261 240.244
R6696 gnd.n6392 gnd.n1261 240.244
R6697 gnd.n6392 gnd.n1255 240.244
R6698 gnd.n6399 gnd.n1255 240.244
R6699 gnd.n6399 gnd.n1256 240.244
R6700 gnd.n1256 gnd.n1230 240.244
R6701 gnd.n6428 gnd.n1230 240.244
R6702 gnd.n6428 gnd.n1225 240.244
R6703 gnd.n6435 gnd.n1225 240.244
R6704 gnd.n6435 gnd.n1205 240.244
R6705 gnd.n6456 gnd.n1205 240.244
R6706 gnd.n6457 gnd.n6456 240.244
R6707 gnd.n6457 gnd.n1201 240.244
R6708 gnd.n6463 gnd.n1201 240.244
R6709 gnd.n6463 gnd.n1175 240.244
R6710 gnd.n6514 gnd.n1175 240.244
R6711 gnd.n6514 gnd.n1169 240.244
R6712 gnd.n6521 gnd.n1169 240.244
R6713 gnd.n6521 gnd.n1170 240.244
R6714 gnd.n1170 gnd.n1140 240.244
R6715 gnd.n6580 gnd.n1140 240.244
R6716 gnd.n6580 gnd.n1134 240.244
R6717 gnd.n6599 gnd.n1134 240.244
R6718 gnd.n6599 gnd.n1135 240.244
R6719 gnd.n6585 gnd.n1135 240.244
R6720 gnd.n6586 gnd.n6585 240.244
R6721 gnd.n6587 gnd.n6586 240.244
R6722 gnd.n6588 gnd.n6587 240.244
R6723 gnd.n6588 gnd.n1084 240.244
R6724 gnd.n6703 gnd.n1084 240.244
R6725 gnd.n6703 gnd.n1078 240.244
R6726 gnd.n6710 gnd.n1078 240.244
R6727 gnd.n6710 gnd.n1079 240.244
R6728 gnd.n1079 gnd.n1054 240.244
R6729 gnd.n6748 gnd.n1054 240.244
R6730 gnd.n6748 gnd.n1048 240.244
R6731 gnd.n6755 gnd.n1048 240.244
R6732 gnd.n6755 gnd.n1049 240.244
R6733 gnd.n1049 gnd.n1030 240.244
R6734 gnd.n6802 gnd.n1030 240.244
R6735 gnd.n6802 gnd.n1031 240.244
R6736 gnd.n6796 gnd.n1031 240.244
R6737 gnd.n6796 gnd.n1002 240.244
R6738 gnd.n6843 gnd.n1002 240.244
R6739 gnd.n6843 gnd.n1003 240.244
R6740 gnd.n6837 gnd.n1003 240.244
R6741 gnd.n6837 gnd.n733 240.244
R6742 gnd.n7005 gnd.n733 240.244
R6743 gnd.n7005 gnd.n727 240.244
R6744 gnd.n7012 gnd.n727 240.244
R6745 gnd.n7012 gnd.n728 240.244
R6746 gnd.n728 gnd.n707 240.244
R6747 gnd.n7035 gnd.n707 240.244
R6748 gnd.n7035 gnd.n701 240.244
R6749 gnd.n7042 gnd.n701 240.244
R6750 gnd.n7042 gnd.n702 240.244
R6751 gnd.n702 gnd.n683 240.244
R6752 gnd.n7071 gnd.n683 240.244
R6753 gnd.n7071 gnd.n679 240.244
R6754 gnd.n7077 gnd.n679 240.244
R6755 gnd.n7077 gnd.n586 240.244
R6756 gnd.n7184 gnd.n586 240.244
R6757 gnd.n1704 gnd.n1703 240.244
R6758 gnd.n1709 gnd.n1703 240.244
R6759 gnd.n1711 gnd.n1710 240.244
R6760 gnd.n1713 gnd.n1712 240.244
R6761 gnd.n5603 gnd.n5602 240.244
R6762 gnd.n5606 gnd.n5605 240.244
R6763 gnd.n5617 gnd.n5616 240.244
R6764 gnd.n5619 gnd.n5618 240.244
R6765 gnd.n5629 gnd.n5628 240.244
R6766 gnd.n5640 gnd.n5639 240.244
R6767 gnd.n5642 gnd.n5641 240.244
R6768 gnd.n5652 gnd.n5651 240.244
R6769 gnd.n5673 gnd.n5672 240.244
R6770 gnd.n1700 gnd.n1686 240.244
R6771 gnd.n5450 gnd.n1687 240.244
R6772 gnd.n5501 gnd.n5450 240.244
R6773 gnd.n5510 gnd.n5501 240.244
R6774 gnd.n5510 gnd.n5488 240.244
R6775 gnd.n5523 gnd.n5488 240.244
R6776 gnd.n5523 gnd.n5484 240.244
R6777 gnd.n5529 gnd.n5484 240.244
R6778 gnd.n5529 gnd.n5475 240.244
R6779 gnd.n5544 gnd.n5475 240.244
R6780 gnd.n5544 gnd.n5469 240.244
R6781 gnd.n5557 gnd.n5469 240.244
R6782 gnd.n5557 gnd.n5470 240.244
R6783 gnd.n5470 gnd.n1466 240.244
R6784 gnd.n1466 gnd.n1459 240.244
R6785 gnd.n1459 gnd.n1451 240.244
R6786 gnd.n6031 gnd.n1451 240.244
R6787 gnd.n6032 gnd.n6031 240.244
R6788 gnd.n6032 gnd.n1428 240.244
R6789 gnd.n6045 gnd.n1428 240.244
R6790 gnd.n6045 gnd.n1421 240.244
R6791 gnd.n6038 gnd.n1421 240.244
R6792 gnd.n6038 gnd.n1400 240.244
R6793 gnd.n1400 gnd.n1392 240.244
R6794 gnd.n6140 gnd.n1392 240.244
R6795 gnd.n6140 gnd.n1381 240.244
R6796 gnd.n1381 gnd.n1373 240.244
R6797 gnd.n6151 gnd.n1373 240.244
R6798 gnd.n6151 gnd.n1365 240.244
R6799 gnd.n6145 gnd.n1365 240.244
R6800 gnd.n6145 gnd.n1341 240.244
R6801 gnd.n6209 gnd.n1341 240.244
R6802 gnd.n6209 gnd.n1334 240.244
R6803 gnd.n6216 gnd.n1334 240.244
R6804 gnd.n6216 gnd.n1309 240.244
R6805 gnd.n1309 gnd.n1299 240.244
R6806 gnd.n6288 gnd.n1299 240.244
R6807 gnd.n6288 gnd.n1295 240.244
R6808 gnd.n6295 gnd.n1295 240.244
R6809 gnd.n6296 gnd.n6295 240.244
R6810 gnd.n6297 gnd.n6296 240.244
R6811 gnd.n6297 gnd.n1263 240.244
R6812 gnd.n1291 gnd.n1263 240.244
R6813 gnd.n1291 gnd.n1253 240.244
R6814 gnd.n6305 gnd.n1253 240.244
R6815 gnd.n6306 gnd.n6305 240.244
R6816 gnd.n6306 gnd.n1232 240.244
R6817 gnd.n6343 gnd.n1232 240.244
R6818 gnd.n6343 gnd.n1224 240.244
R6819 gnd.n1224 gnd.n1215 240.244
R6820 gnd.n1215 gnd.n1207 240.244
R6821 gnd.n6311 gnd.n1207 240.244
R6822 gnd.n6312 gnd.n6311 240.244
R6823 gnd.n6312 gnd.n1200 240.244
R6824 gnd.n1200 gnd.n1184 240.244
R6825 gnd.n1184 gnd.n1177 240.244
R6826 gnd.n6324 gnd.n1177 240.244
R6827 gnd.n6324 gnd.n1167 240.244
R6828 gnd.n1167 gnd.n1155 240.244
R6829 gnd.n6539 gnd.n1155 240.244
R6830 gnd.n6539 gnd.n1142 240.244
R6831 gnd.n6559 gnd.n1142 240.244
R6832 gnd.n6559 gnd.n1133 240.244
R6833 gnd.n6544 gnd.n1133 240.244
R6834 gnd.n6545 gnd.n6544 240.244
R6835 gnd.n6546 gnd.n6545 240.244
R6836 gnd.n6547 gnd.n6546 240.244
R6837 gnd.n6547 gnd.n1107 240.244
R6838 gnd.n6641 gnd.n1107 240.244
R6839 gnd.n6641 gnd.n1086 240.244
R6840 gnd.n1103 gnd.n1086 240.244
R6841 gnd.n1103 gnd.n1077 240.244
R6842 gnd.n6648 gnd.n1077 240.244
R6843 gnd.n6648 gnd.n1063 240.244
R6844 gnd.n1063 gnd.n1056 240.244
R6845 gnd.n6671 gnd.n1056 240.244
R6846 gnd.n6671 gnd.n1046 240.244
R6847 gnd.n6654 gnd.n1046 240.244
R6848 gnd.n6658 gnd.n6654 240.244
R6849 gnd.n6658 gnd.n1028 240.244
R6850 gnd.n6659 gnd.n1028 240.244
R6851 gnd.n6659 gnd.n1013 240.244
R6852 gnd.n6824 gnd.n1013 240.244
R6853 gnd.n6824 gnd.n1000 240.244
R6854 gnd.n1007 gnd.n1000 240.244
R6855 gnd.n6834 gnd.n1007 240.244
R6856 gnd.n6834 gnd.n1008 240.244
R6857 gnd.n1008 gnd.n735 240.244
R6858 gnd.n735 gnd.n723 240.244
R6859 gnd.n7014 gnd.n723 240.244
R6860 gnd.n7014 gnd.n718 240.244
R6861 gnd.n7021 gnd.n718 240.244
R6862 gnd.n7021 gnd.n709 240.244
R6863 gnd.n709 gnd.n698 240.244
R6864 gnd.n7044 gnd.n698 240.244
R6865 gnd.n7044 gnd.n693 240.244
R6866 gnd.n7056 gnd.n693 240.244
R6867 gnd.n7056 gnd.n685 240.244
R6868 gnd.n7049 gnd.n685 240.244
R6869 gnd.n7049 gnd.n678 240.244
R6870 gnd.n678 gnd.n583 240.244
R6871 gnd.n7186 gnd.n583 240.244
R6872 gnd.n592 gnd.n591 240.244
R6873 gnd.n649 gnd.n595 240.244
R6874 gnd.n597 gnd.n596 240.244
R6875 gnd.n652 gnd.n601 240.244
R6876 gnd.n655 gnd.n602 240.244
R6877 gnd.n612 gnd.n611 240.244
R6878 gnd.n657 gnd.n621 240.244
R6879 gnd.n660 gnd.n622 240.244
R6880 gnd.n630 gnd.n629 240.244
R6881 gnd.n662 gnd.n639 240.244
R6882 gnd.n665 gnd.n640 240.244
R6883 gnd.n7125 gnd.n646 240.244
R6884 gnd.n7125 gnd.n577 240.244
R6885 gnd.n579 gnd.n578 240.244
R6886 gnd.n1477 gnd.n1476 240.132
R6887 gnd.n752 gnd.n751 240.132
R6888 gnd.n3165 gnd.n2207 225.874
R6889 gnd.n3157 gnd.n2207 225.874
R6890 gnd.n3157 gnd.n3156 225.874
R6891 gnd.n3156 gnd.n3155 225.874
R6892 gnd.n3155 gnd.n2213 225.874
R6893 gnd.n3149 gnd.n2213 225.874
R6894 gnd.n3149 gnd.n3148 225.874
R6895 gnd.n3148 gnd.n3147 225.874
R6896 gnd.n3147 gnd.n2220 225.874
R6897 gnd.n3141 gnd.n2220 225.874
R6898 gnd.n3141 gnd.n3140 225.874
R6899 gnd.n3140 gnd.n3139 225.874
R6900 gnd.n3139 gnd.n2228 225.874
R6901 gnd.n3133 gnd.n2228 225.874
R6902 gnd.n3133 gnd.n3132 225.874
R6903 gnd.n3132 gnd.n3131 225.874
R6904 gnd.n3131 gnd.n2236 225.874
R6905 gnd.n3125 gnd.n2236 225.874
R6906 gnd.n3125 gnd.n3124 225.874
R6907 gnd.n3124 gnd.n3123 225.874
R6908 gnd.n3123 gnd.n2244 225.874
R6909 gnd.n3117 gnd.n2244 225.874
R6910 gnd.n3117 gnd.n3116 225.874
R6911 gnd.n3116 gnd.n3115 225.874
R6912 gnd.n3115 gnd.n2252 225.874
R6913 gnd.n3109 gnd.n2252 225.874
R6914 gnd.n3109 gnd.n3108 225.874
R6915 gnd.n3108 gnd.n3107 225.874
R6916 gnd.n3107 gnd.n2260 225.874
R6917 gnd.n3101 gnd.n2260 225.874
R6918 gnd.n3101 gnd.n3100 225.874
R6919 gnd.n3100 gnd.n3099 225.874
R6920 gnd.n3099 gnd.n2268 225.874
R6921 gnd.n3093 gnd.n2268 225.874
R6922 gnd.n3093 gnd.n3092 225.874
R6923 gnd.n3092 gnd.n3091 225.874
R6924 gnd.n3091 gnd.n2276 225.874
R6925 gnd.n3085 gnd.n2276 225.874
R6926 gnd.n3085 gnd.n3084 225.874
R6927 gnd.n3084 gnd.n3083 225.874
R6928 gnd.n3083 gnd.n2284 225.874
R6929 gnd.n3077 gnd.n2284 225.874
R6930 gnd.n3077 gnd.n3076 225.874
R6931 gnd.n3076 gnd.n3075 225.874
R6932 gnd.n3075 gnd.n2292 225.874
R6933 gnd.n3069 gnd.n2292 225.874
R6934 gnd.n3069 gnd.n3068 225.874
R6935 gnd.n3068 gnd.n3067 225.874
R6936 gnd.n3067 gnd.n2300 225.874
R6937 gnd.n3061 gnd.n2300 225.874
R6938 gnd.n3061 gnd.n3060 225.874
R6939 gnd.n3060 gnd.n3059 225.874
R6940 gnd.n3059 gnd.n2308 225.874
R6941 gnd.n3053 gnd.n2308 225.874
R6942 gnd.n3053 gnd.n3052 225.874
R6943 gnd.n3052 gnd.n3051 225.874
R6944 gnd.n3051 gnd.n2316 225.874
R6945 gnd.n3045 gnd.n2316 225.874
R6946 gnd.n3045 gnd.n3044 225.874
R6947 gnd.n3044 gnd.n3043 225.874
R6948 gnd.n3043 gnd.n2324 225.874
R6949 gnd.n3037 gnd.n2324 225.874
R6950 gnd.n3037 gnd.n3036 225.874
R6951 gnd.n3036 gnd.n3035 225.874
R6952 gnd.n3035 gnd.n2332 225.874
R6953 gnd.n3029 gnd.n2332 225.874
R6954 gnd.n3029 gnd.n3028 225.874
R6955 gnd.n3028 gnd.n3027 225.874
R6956 gnd.n3027 gnd.n2340 225.874
R6957 gnd.n3021 gnd.n2340 225.874
R6958 gnd.n3021 gnd.n3020 225.874
R6959 gnd.n3020 gnd.n3019 225.874
R6960 gnd.n3019 gnd.n2348 225.874
R6961 gnd.n3013 gnd.n2348 225.874
R6962 gnd.n3013 gnd.n3012 225.874
R6963 gnd.n3012 gnd.n3011 225.874
R6964 gnd.n3011 gnd.n2356 225.874
R6965 gnd.n3005 gnd.n2356 225.874
R6966 gnd.n3005 gnd.n3004 225.874
R6967 gnd.n3004 gnd.n3003 225.874
R6968 gnd.n3003 gnd.n2364 225.874
R6969 gnd.n2997 gnd.n2364 225.874
R6970 gnd.n2997 gnd.n2996 225.874
R6971 gnd.n2996 gnd.n2995 225.874
R6972 gnd.n2995 gnd.n2372 225.874
R6973 gnd.n2989 gnd.n2372 225.874
R6974 gnd.n2989 gnd.n2988 225.874
R6975 gnd.n2988 gnd.n2987 225.874
R6976 gnd.n2987 gnd.n2380 225.874
R6977 gnd.n2981 gnd.n2380 225.874
R6978 gnd.n2981 gnd.n2980 225.874
R6979 gnd.n2980 gnd.n2979 225.874
R6980 gnd.n2979 gnd.n2388 225.874
R6981 gnd.n2973 gnd.n2388 225.874
R6982 gnd.n2973 gnd.n2972 225.874
R6983 gnd.n2972 gnd.n2971 225.874
R6984 gnd.n2971 gnd.n2396 225.874
R6985 gnd.n2965 gnd.n2396 225.874
R6986 gnd.n2965 gnd.n2964 225.874
R6987 gnd.n2964 gnd.n2963 225.874
R6988 gnd.n2963 gnd.n2404 225.874
R6989 gnd.n2957 gnd.n2404 225.874
R6990 gnd.n2957 gnd.n2956 225.874
R6991 gnd.n2956 gnd.n2955 225.874
R6992 gnd.n2955 gnd.n2412 225.874
R6993 gnd.n2949 gnd.n2412 225.874
R6994 gnd.n2949 gnd.n2948 225.874
R6995 gnd.n2948 gnd.n2947 225.874
R6996 gnd.n2947 gnd.n2420 225.874
R6997 gnd.n2941 gnd.n2420 225.874
R6998 gnd.n2941 gnd.n2940 225.874
R6999 gnd.n2940 gnd.n2939 225.874
R7000 gnd.n2939 gnd.n2428 225.874
R7001 gnd.n2933 gnd.n2428 225.874
R7002 gnd.n2933 gnd.n2932 225.874
R7003 gnd.n2932 gnd.n2931 225.874
R7004 gnd.n2931 gnd.n2436 225.874
R7005 gnd.n2925 gnd.n2436 225.874
R7006 gnd.n2925 gnd.n2924 225.874
R7007 gnd.n2924 gnd.n2923 225.874
R7008 gnd.n2923 gnd.n2444 225.874
R7009 gnd.n2917 gnd.n2444 225.874
R7010 gnd.n2917 gnd.n2916 225.874
R7011 gnd.n2916 gnd.n2915 225.874
R7012 gnd.n2915 gnd.n2452 225.874
R7013 gnd.n2909 gnd.n2452 225.874
R7014 gnd.n2909 gnd.n2908 225.874
R7015 gnd.n2908 gnd.n2907 225.874
R7016 gnd.n2907 gnd.n2460 225.874
R7017 gnd.n2901 gnd.n2460 225.874
R7018 gnd.n2901 gnd.n2900 225.874
R7019 gnd.n2900 gnd.n2899 225.874
R7020 gnd.n2899 gnd.n2468 225.874
R7021 gnd.n2893 gnd.n2468 225.874
R7022 gnd.n2893 gnd.n2892 225.874
R7023 gnd.n2892 gnd.n2891 225.874
R7024 gnd.n2891 gnd.n2476 225.874
R7025 gnd.n2885 gnd.n2476 225.874
R7026 gnd.n2885 gnd.n2884 225.874
R7027 gnd.n2884 gnd.n2883 225.874
R7028 gnd.n2883 gnd.n2484 225.874
R7029 gnd.n2877 gnd.n2484 225.874
R7030 gnd.n2877 gnd.n2876 225.874
R7031 gnd.n2876 gnd.n2875 225.874
R7032 gnd.n2875 gnd.n2492 225.874
R7033 gnd.n2869 gnd.n2492 225.874
R7034 gnd.n2869 gnd.n2868 225.874
R7035 gnd.n2868 gnd.n2867 225.874
R7036 gnd.n2867 gnd.n2500 225.874
R7037 gnd.n2861 gnd.n2500 225.874
R7038 gnd.n2861 gnd.n2860 225.874
R7039 gnd.n2860 gnd.n2859 225.874
R7040 gnd.n2859 gnd.n2508 225.874
R7041 gnd.n2853 gnd.n2508 225.874
R7042 gnd.n3868 gnd.t187 224.174
R7043 gnd.n2057 gnd.t170 224.174
R7044 gnd.n788 gnd.n541 199.319
R7045 gnd.n788 gnd.n542 199.319
R7046 gnd.n5813 gnd.n1591 199.319
R7047 gnd.n1596 gnd.n1591 199.319
R7048 gnd.n1478 gnd.n1475 186.49
R7049 gnd.n753 gnd.n750 186.49
R7050 gnd.n4643 gnd.n4642 185
R7051 gnd.n4641 gnd.n4640 185
R7052 gnd.n4620 gnd.n4619 185
R7053 gnd.n4635 gnd.n4634 185
R7054 gnd.n4633 gnd.n4632 185
R7055 gnd.n4624 gnd.n4623 185
R7056 gnd.n4627 gnd.n4626 185
R7057 gnd.n4611 gnd.n4610 185
R7058 gnd.n4609 gnd.n4608 185
R7059 gnd.n4588 gnd.n4587 185
R7060 gnd.n4603 gnd.n4602 185
R7061 gnd.n4601 gnd.n4600 185
R7062 gnd.n4592 gnd.n4591 185
R7063 gnd.n4595 gnd.n4594 185
R7064 gnd.n4579 gnd.n4578 185
R7065 gnd.n4577 gnd.n4576 185
R7066 gnd.n4556 gnd.n4555 185
R7067 gnd.n4571 gnd.n4570 185
R7068 gnd.n4569 gnd.n4568 185
R7069 gnd.n4560 gnd.n4559 185
R7070 gnd.n4563 gnd.n4562 185
R7071 gnd.n4548 gnd.n4547 185
R7072 gnd.n4546 gnd.n4545 185
R7073 gnd.n4525 gnd.n4524 185
R7074 gnd.n4540 gnd.n4539 185
R7075 gnd.n4538 gnd.n4537 185
R7076 gnd.n4529 gnd.n4528 185
R7077 gnd.n4532 gnd.n4531 185
R7078 gnd.n4516 gnd.n4515 185
R7079 gnd.n4514 gnd.n4513 185
R7080 gnd.n4493 gnd.n4492 185
R7081 gnd.n4508 gnd.n4507 185
R7082 gnd.n4506 gnd.n4505 185
R7083 gnd.n4497 gnd.n4496 185
R7084 gnd.n4500 gnd.n4499 185
R7085 gnd.n4484 gnd.n4483 185
R7086 gnd.n4482 gnd.n4481 185
R7087 gnd.n4461 gnd.n4460 185
R7088 gnd.n4476 gnd.n4475 185
R7089 gnd.n4474 gnd.n4473 185
R7090 gnd.n4465 gnd.n4464 185
R7091 gnd.n4468 gnd.n4467 185
R7092 gnd.n4452 gnd.n4451 185
R7093 gnd.n4450 gnd.n4449 185
R7094 gnd.n4429 gnd.n4428 185
R7095 gnd.n4444 gnd.n4443 185
R7096 gnd.n4442 gnd.n4441 185
R7097 gnd.n4433 gnd.n4432 185
R7098 gnd.n4436 gnd.n4435 185
R7099 gnd.n4421 gnd.n4420 185
R7100 gnd.n4419 gnd.n4418 185
R7101 gnd.n4398 gnd.n4397 185
R7102 gnd.n4413 gnd.n4412 185
R7103 gnd.n4411 gnd.n4410 185
R7104 gnd.n4402 gnd.n4401 185
R7105 gnd.n4405 gnd.n4404 185
R7106 gnd.n3869 gnd.t186 178.987
R7107 gnd.n2058 gnd.t171 178.987
R7108 gnd.n1 gnd.t48 170.774
R7109 gnd.n9 gnd.t19 170.103
R7110 gnd.n8 gnd.t66 170.103
R7111 gnd.n7 gnd.t8 170.103
R7112 gnd.n6 gnd.t17 170.103
R7113 gnd.n5 gnd.t358 170.103
R7114 gnd.n4 gnd.t5 170.103
R7115 gnd.n3 gnd.t63 170.103
R7116 gnd.n2 gnd.t3 170.103
R7117 gnd.n1 gnd.t61 170.103
R7118 gnd.n6995 gnd.n6994 163.367
R7119 gnd.n6992 gnd.n762 163.367
R7120 gnd.n6988 gnd.n6987 163.367
R7121 gnd.n6985 gnd.n765 163.367
R7122 gnd.n6981 gnd.n6980 163.367
R7123 gnd.n6978 gnd.n768 163.367
R7124 gnd.n6974 gnd.n6973 163.367
R7125 gnd.n6971 gnd.n771 163.367
R7126 gnd.n6967 gnd.n6966 163.367
R7127 gnd.n6964 gnd.n774 163.367
R7128 gnd.n6960 gnd.n6959 163.367
R7129 gnd.n6957 gnd.n777 163.367
R7130 gnd.n6953 gnd.n6952 163.367
R7131 gnd.n6950 gnd.n780 163.367
R7132 gnd.n6945 gnd.n6944 163.367
R7133 gnd.n6942 gnd.n785 163.367
R7134 gnd.n6938 gnd.n6937 163.367
R7135 gnd.n6935 gnd.n961 163.367
R7136 gnd.n6930 gnd.n6929 163.367
R7137 gnd.n6927 gnd.n966 163.367
R7138 gnd.n6923 gnd.n6922 163.367
R7139 gnd.n6920 gnd.n969 163.367
R7140 gnd.n6916 gnd.n6915 163.367
R7141 gnd.n6913 gnd.n972 163.367
R7142 gnd.n6909 gnd.n6908 163.367
R7143 gnd.n6906 gnd.n975 163.367
R7144 gnd.n6902 gnd.n6901 163.367
R7145 gnd.n6899 gnd.n978 163.367
R7146 gnd.n6895 gnd.n6894 163.367
R7147 gnd.n6892 gnd.n981 163.367
R7148 gnd.n6888 gnd.n6887 163.367
R7149 gnd.n6885 gnd.n984 163.367
R7150 gnd.n5995 gnd.n1467 163.367
R7151 gnd.n5995 gnd.n1440 163.367
R7152 gnd.n6062 gnd.n1440 163.367
R7153 gnd.n6062 gnd.n1437 163.367
R7154 gnd.n6071 gnd.n1437 163.367
R7155 gnd.n6071 gnd.n1438 163.367
R7156 gnd.n6067 gnd.n1438 163.367
R7157 gnd.n6067 gnd.n6066 163.367
R7158 gnd.n6066 gnd.n1419 163.367
R7159 gnd.n6091 gnd.n1419 163.367
R7160 gnd.n6091 gnd.n1408 163.367
R7161 gnd.n6097 gnd.n1408 163.367
R7162 gnd.n6098 gnd.n6097 163.367
R7163 gnd.n6098 gnd.n1416 163.367
R7164 gnd.n6103 gnd.n1416 163.367
R7165 gnd.n6103 gnd.n1417 163.367
R7166 gnd.n1417 gnd.n1380 163.367
R7167 gnd.n6158 gnd.n1380 163.367
R7168 gnd.n6158 gnd.n1374 163.367
R7169 gnd.n6154 gnd.n1374 163.367
R7170 gnd.n6154 gnd.n1386 163.367
R7171 gnd.n1386 gnd.n1385 163.367
R7172 gnd.n1385 gnd.n1357 163.367
R7173 gnd.n6195 gnd.n1357 163.367
R7174 gnd.n6195 gnd.n1342 163.367
R7175 gnd.n6206 gnd.n1342 163.367
R7176 gnd.n6206 gnd.n1355 163.367
R7177 gnd.n6202 gnd.n1355 163.367
R7178 gnd.n6202 gnd.n1350 163.367
R7179 gnd.n6199 gnd.n1350 163.367
R7180 gnd.n6199 gnd.n1310 163.367
R7181 gnd.n1317 gnd.n1310 163.367
R7182 gnd.n6264 gnd.n1317 163.367
R7183 gnd.n6264 gnd.n1318 163.367
R7184 gnd.n6260 gnd.n1318 163.367
R7185 gnd.n6260 gnd.n1321 163.367
R7186 gnd.n1321 gnd.n1278 163.367
R7187 gnd.n6369 gnd.n1278 163.367
R7188 gnd.n6369 gnd.n1271 163.367
R7189 gnd.n6365 gnd.n1271 163.367
R7190 gnd.n6365 gnd.n6362 163.367
R7191 gnd.n6362 gnd.n6361 163.367
R7192 gnd.n6361 gnd.n1252 163.367
R7193 gnd.n6357 gnd.n1252 163.367
R7194 gnd.n6357 gnd.n1246 163.367
R7195 gnd.n6354 gnd.n1246 163.367
R7196 gnd.n6354 gnd.n1239 163.367
R7197 gnd.n6349 gnd.n1239 163.367
R7198 gnd.n6349 gnd.n1233 163.367
R7199 gnd.n6346 gnd.n1233 163.367
R7200 gnd.n6346 gnd.n1223 163.367
R7201 gnd.n1285 gnd.n1223 163.367
R7202 gnd.n1285 gnd.n1216 163.367
R7203 gnd.n1282 gnd.n1216 163.367
R7204 gnd.n1282 gnd.n1208 163.367
R7205 gnd.n1208 gnd.n1197 163.367
R7206 gnd.n6470 gnd.n1197 163.367
R7207 gnd.n6470 gnd.n1192 163.367
R7208 gnd.n6466 gnd.n1192 163.367
R7209 gnd.n6466 gnd.n1183 163.367
R7210 gnd.n6316 gnd.n1183 163.367
R7211 gnd.n6316 gnd.n1178 163.367
R7212 gnd.n6321 gnd.n1178 163.367
R7213 gnd.n6321 gnd.n1166 163.367
R7214 gnd.n1166 gnd.n1159 163.367
R7215 gnd.n6531 gnd.n1159 163.367
R7216 gnd.n6531 gnd.n1157 163.367
R7217 gnd.n6536 gnd.n1157 163.367
R7218 gnd.n6536 gnd.n1143 163.367
R7219 gnd.n6562 gnd.n1143 163.367
R7220 gnd.n6563 gnd.n6562 163.367
R7221 gnd.n6563 gnd.n1148 163.367
R7222 gnd.n6568 gnd.n1148 163.367
R7223 gnd.n6568 gnd.n1123 163.367
R7224 gnd.n1123 gnd.n1115 163.367
R7225 gnd.n6625 gnd.n1115 163.367
R7226 gnd.n6625 gnd.n1113 163.367
R7227 gnd.n6629 gnd.n1113 163.367
R7228 gnd.n6629 gnd.n1095 163.367
R7229 gnd.n6692 gnd.n1095 163.367
R7230 gnd.n6692 gnd.n1096 163.367
R7231 gnd.n6688 gnd.n1096 163.367
R7232 gnd.n6688 gnd.n6687 163.367
R7233 gnd.n6687 gnd.n1075 163.367
R7234 gnd.n1076 gnd.n1075 163.367
R7235 gnd.n1076 gnd.n1070 163.367
R7236 gnd.n6681 gnd.n1070 163.367
R7237 gnd.n6681 gnd.n1062 163.367
R7238 gnd.n6677 gnd.n1062 163.367
R7239 gnd.n6677 gnd.n1057 163.367
R7240 gnd.n6674 gnd.n1057 163.367
R7241 gnd.n6674 gnd.n1045 163.367
R7242 gnd.n1045 gnd.n1038 163.367
R7243 gnd.n6769 gnd.n1038 163.367
R7244 gnd.n6769 gnd.n1036 163.367
R7245 gnd.n6773 gnd.n1036 163.367
R7246 gnd.n6774 gnd.n6773 163.367
R7247 gnd.n6777 gnd.n6774 163.367
R7248 gnd.n6777 gnd.n1021 163.367
R7249 gnd.n6793 gnd.n1021 163.367
R7250 gnd.n6793 gnd.n1015 163.367
R7251 gnd.n6789 gnd.n1015 163.367
R7252 gnd.n6789 gnd.n6788 163.367
R7253 gnd.n6788 gnd.n6787 163.367
R7254 gnd.n6787 gnd.n992 163.367
R7255 gnd.n992 gnd.n986 163.367
R7256 gnd.n6872 gnd.n986 163.367
R7257 gnd.n6873 gnd.n6872 163.367
R7258 gnd.n6873 gnd.n736 163.367
R7259 gnd.n6880 gnd.n736 163.367
R7260 gnd.n6003 gnd.n1492 163.367
R7261 gnd.n1531 gnd.n1492 163.367
R7262 gnd.n1535 gnd.n1534 163.367
R7263 gnd.n1539 gnd.n1538 163.367
R7264 gnd.n1543 gnd.n1542 163.367
R7265 gnd.n1547 gnd.n1546 163.367
R7266 gnd.n1551 gnd.n1550 163.367
R7267 gnd.n1555 gnd.n1554 163.367
R7268 gnd.n1559 gnd.n1558 163.367
R7269 gnd.n1563 gnd.n1562 163.367
R7270 gnd.n1567 gnd.n1566 163.367
R7271 gnd.n1571 gnd.n1570 163.367
R7272 gnd.n1575 gnd.n1574 163.367
R7273 gnd.n1579 gnd.n1578 163.367
R7274 gnd.n1583 gnd.n1582 163.367
R7275 gnd.n1587 gnd.n1586 163.367
R7276 gnd.n5933 gnd.n5932 163.367
R7277 gnd.n5937 gnd.n5936 163.367
R7278 gnd.n5942 gnd.n5941 163.367
R7279 gnd.n5946 gnd.n5945 163.367
R7280 gnd.n5950 gnd.n5949 163.367
R7281 gnd.n5954 gnd.n5953 163.367
R7282 gnd.n5958 gnd.n5957 163.367
R7283 gnd.n5962 gnd.n5961 163.367
R7284 gnd.n5966 gnd.n5965 163.367
R7285 gnd.n5970 gnd.n5969 163.367
R7286 gnd.n5974 gnd.n5973 163.367
R7287 gnd.n5978 gnd.n5977 163.367
R7288 gnd.n5982 gnd.n5981 163.367
R7289 gnd.n5986 gnd.n5985 163.367
R7290 gnd.n5990 gnd.n5989 163.367
R7291 gnd.n5992 gnd.n1525 163.367
R7292 gnd.n6009 gnd.n1470 163.367
R7293 gnd.n1470 gnd.n1443 163.367
R7294 gnd.n6060 gnd.n1443 163.367
R7295 gnd.n6060 gnd.n1444 163.367
R7296 gnd.n1444 gnd.n1435 163.367
R7297 gnd.n6055 gnd.n1435 163.367
R7298 gnd.n6055 gnd.n6052 163.367
R7299 gnd.n6052 gnd.n6051 163.367
R7300 gnd.n6051 gnd.n6048 163.367
R7301 gnd.n6048 gnd.n1410 163.367
R7302 gnd.n6112 gnd.n1410 163.367
R7303 gnd.n6112 gnd.n1411 163.367
R7304 gnd.n6108 gnd.n1411 163.367
R7305 gnd.n6108 gnd.n6107 163.367
R7306 gnd.n6107 gnd.n6106 163.367
R7307 gnd.n6106 gnd.n1378 163.367
R7308 gnd.n6162 gnd.n1378 163.367
R7309 gnd.n6162 gnd.n1375 163.367
R7310 gnd.n6174 gnd.n1375 163.367
R7311 gnd.n6174 gnd.n1376 163.367
R7312 gnd.n6170 gnd.n1376 163.367
R7313 gnd.n6170 gnd.n6169 163.367
R7314 gnd.n6169 gnd.n6168 163.367
R7315 gnd.n6168 gnd.n1344 163.367
R7316 gnd.n6225 gnd.n1344 163.367
R7317 gnd.n6225 gnd.n1345 163.367
R7318 gnd.n6221 gnd.n1345 163.367
R7319 gnd.n6221 gnd.n6220 163.367
R7320 gnd.n6220 gnd.n6219 163.367
R7321 gnd.n6219 gnd.n1311 163.367
R7322 gnd.n6270 gnd.n1311 163.367
R7323 gnd.n6270 gnd.n1312 163.367
R7324 gnd.n6266 gnd.n1312 163.367
R7325 gnd.n6266 gnd.n1315 163.367
R7326 gnd.n6258 gnd.n1315 163.367
R7327 gnd.n6258 gnd.n1276 163.367
R7328 gnd.n6373 gnd.n1276 163.367
R7329 gnd.n6373 gnd.n1273 163.367
R7330 gnd.n6380 gnd.n1273 163.367
R7331 gnd.n6380 gnd.n1274 163.367
R7332 gnd.n6376 gnd.n1274 163.367
R7333 gnd.n6376 gnd.n1250 163.367
R7334 gnd.n6403 gnd.n1250 163.367
R7335 gnd.n6403 gnd.n1248 163.367
R7336 gnd.n6407 gnd.n1248 163.367
R7337 gnd.n6407 gnd.n1237 163.367
R7338 gnd.n6421 gnd.n1237 163.367
R7339 gnd.n6421 gnd.n1235 163.367
R7340 gnd.n6425 gnd.n1235 163.367
R7341 gnd.n6425 gnd.n1221 163.367
R7342 gnd.n6438 gnd.n1221 163.367
R7343 gnd.n6438 gnd.n1218 163.367
R7344 gnd.n6443 gnd.n1218 163.367
R7345 gnd.n6443 gnd.n1219 163.367
R7346 gnd.n1219 gnd.n1195 163.367
R7347 gnd.n6474 gnd.n1195 163.367
R7348 gnd.n6474 gnd.n1193 163.367
R7349 gnd.n6478 gnd.n1193 163.367
R7350 gnd.n6478 gnd.n1181 163.367
R7351 gnd.n6507 gnd.n1181 163.367
R7352 gnd.n6507 gnd.n1179 163.367
R7353 gnd.n6511 gnd.n1179 163.367
R7354 gnd.n6511 gnd.n1164 163.367
R7355 gnd.n6524 gnd.n1164 163.367
R7356 gnd.n6524 gnd.n1161 163.367
R7357 gnd.n6529 gnd.n1161 163.367
R7358 gnd.n6529 gnd.n1162 163.367
R7359 gnd.n1162 gnd.n1144 163.367
R7360 gnd.n6577 gnd.n1144 163.367
R7361 gnd.n6577 gnd.n1145 163.367
R7362 gnd.n6573 gnd.n1145 163.367
R7363 gnd.n6573 gnd.n6572 163.367
R7364 gnd.n6572 gnd.n1121 163.367
R7365 gnd.n6618 gnd.n1121 163.367
R7366 gnd.n6618 gnd.n1118 163.367
R7367 gnd.n6623 gnd.n1118 163.367
R7368 gnd.n6623 gnd.n1119 163.367
R7369 gnd.n1119 gnd.n1111 163.367
R7370 gnd.n6633 gnd.n1111 163.367
R7371 gnd.n6633 gnd.n1094 163.367
R7372 gnd.n6638 gnd.n1094 163.367
R7373 gnd.n6638 gnd.n1109 163.367
R7374 gnd.n1109 gnd.n1074 163.367
R7375 gnd.n6715 gnd.n1074 163.367
R7376 gnd.n6715 gnd.n1072 163.367
R7377 gnd.n6719 gnd.n1072 163.367
R7378 gnd.n6719 gnd.n1061 163.367
R7379 gnd.n6741 gnd.n1061 163.367
R7380 gnd.n6741 gnd.n1059 163.367
R7381 gnd.n6745 gnd.n1059 163.367
R7382 gnd.n6745 gnd.n1043 163.367
R7383 gnd.n6758 gnd.n1043 163.367
R7384 gnd.n6758 gnd.n1040 163.367
R7385 gnd.n6767 gnd.n1040 163.367
R7386 gnd.n6767 gnd.n1041 163.367
R7387 gnd.n6763 gnd.n1041 163.367
R7388 gnd.n6763 gnd.n6762 163.367
R7389 gnd.n6762 gnd.n1019 163.367
R7390 gnd.n6814 gnd.n1019 163.367
R7391 gnd.n6814 gnd.n1016 163.367
R7392 gnd.n6821 gnd.n1016 163.367
R7393 gnd.n6821 gnd.n1017 163.367
R7394 gnd.n6817 gnd.n1017 163.367
R7395 gnd.n6817 gnd.n991 163.367
R7396 gnd.n6866 gnd.n991 163.367
R7397 gnd.n6866 gnd.n989 163.367
R7398 gnd.n6870 gnd.n989 163.367
R7399 gnd.n6870 gnd.n738 163.367
R7400 gnd.n7002 gnd.n738 163.367
R7401 gnd.n7002 gnd.n739 163.367
R7402 gnd.n759 gnd.n758 156.462
R7403 gnd.n4583 gnd.n4551 153.042
R7404 gnd.n4647 gnd.n4646 152.079
R7405 gnd.n4615 gnd.n4614 152.079
R7406 gnd.n4583 gnd.n4582 152.079
R7407 gnd.n1483 gnd.n1482 152
R7408 gnd.n1484 gnd.n1473 152
R7409 gnd.n1486 gnd.n1485 152
R7410 gnd.n1488 gnd.n1471 152
R7411 gnd.n1490 gnd.n1489 152
R7412 gnd.n757 gnd.n741 152
R7413 gnd.n749 gnd.n742 152
R7414 gnd.n748 gnd.n747 152
R7415 gnd.n746 gnd.n743 152
R7416 gnd.n744 gnd.t156 150.546
R7417 gnd.t371 gnd.n4625 147.661
R7418 gnd.t50 gnd.n4593 147.661
R7419 gnd.t366 gnd.n4561 147.661
R7420 gnd.t362 gnd.n4530 147.661
R7421 gnd.t373 gnd.n4498 147.661
R7422 gnd.t44 gnd.n4466 147.661
R7423 gnd.t352 gnd.n4434 147.661
R7424 gnd.t34 gnd.n4403 147.661
R7425 gnd.n6939 gnd.n960 143.351
R7426 gnd.n5930 gnd.n1508 143.351
R7427 gnd.n5930 gnd.n1509 143.351
R7428 gnd.n1480 gnd.t81 130.484
R7429 gnd.n1489 gnd.t153 126.766
R7430 gnd.n1487 gnd.t74 126.766
R7431 gnd.n1473 gnd.t99 126.766
R7432 gnd.n1481 gnd.t181 126.766
R7433 gnd.n745 gnd.t131 126.766
R7434 gnd.n747 gnd.t71 126.766
R7435 gnd.n756 gnd.t117 126.766
R7436 gnd.n758 gnd.t92 126.766
R7437 gnd.n6940 gnd.n959 104.897
R7438 gnd.n5931 gnd.n5929 104.897
R7439 gnd.n4642 gnd.n4641 104.615
R7440 gnd.n4641 gnd.n4619 104.615
R7441 gnd.n4634 gnd.n4619 104.615
R7442 gnd.n4634 gnd.n4633 104.615
R7443 gnd.n4633 gnd.n4623 104.615
R7444 gnd.n4626 gnd.n4623 104.615
R7445 gnd.n4610 gnd.n4609 104.615
R7446 gnd.n4609 gnd.n4587 104.615
R7447 gnd.n4602 gnd.n4587 104.615
R7448 gnd.n4602 gnd.n4601 104.615
R7449 gnd.n4601 gnd.n4591 104.615
R7450 gnd.n4594 gnd.n4591 104.615
R7451 gnd.n4578 gnd.n4577 104.615
R7452 gnd.n4577 gnd.n4555 104.615
R7453 gnd.n4570 gnd.n4555 104.615
R7454 gnd.n4570 gnd.n4569 104.615
R7455 gnd.n4569 gnd.n4559 104.615
R7456 gnd.n4562 gnd.n4559 104.615
R7457 gnd.n4547 gnd.n4546 104.615
R7458 gnd.n4546 gnd.n4524 104.615
R7459 gnd.n4539 gnd.n4524 104.615
R7460 gnd.n4539 gnd.n4538 104.615
R7461 gnd.n4538 gnd.n4528 104.615
R7462 gnd.n4531 gnd.n4528 104.615
R7463 gnd.n4515 gnd.n4514 104.615
R7464 gnd.n4514 gnd.n4492 104.615
R7465 gnd.n4507 gnd.n4492 104.615
R7466 gnd.n4507 gnd.n4506 104.615
R7467 gnd.n4506 gnd.n4496 104.615
R7468 gnd.n4499 gnd.n4496 104.615
R7469 gnd.n4483 gnd.n4482 104.615
R7470 gnd.n4482 gnd.n4460 104.615
R7471 gnd.n4475 gnd.n4460 104.615
R7472 gnd.n4475 gnd.n4474 104.615
R7473 gnd.n4474 gnd.n4464 104.615
R7474 gnd.n4467 gnd.n4464 104.615
R7475 gnd.n4451 gnd.n4450 104.615
R7476 gnd.n4450 gnd.n4428 104.615
R7477 gnd.n4443 gnd.n4428 104.615
R7478 gnd.n4443 gnd.n4442 104.615
R7479 gnd.n4442 gnd.n4432 104.615
R7480 gnd.n4435 gnd.n4432 104.615
R7481 gnd.n4420 gnd.n4419 104.615
R7482 gnd.n4419 gnd.n4397 104.615
R7483 gnd.n4412 gnd.n4397 104.615
R7484 gnd.n4412 gnd.n4411 104.615
R7485 gnd.n4411 gnd.n4401 104.615
R7486 gnd.n4404 gnd.n4401 104.615
R7487 gnd.n3794 gnd.t116 100.632
R7488 gnd.n2031 gnd.t145 100.632
R7489 gnd.n7671 gnd.n218 99.6594
R7490 gnd.n7669 gnd.n7668 99.6594
R7491 gnd.n7664 gnd.n225 99.6594
R7492 gnd.n7662 gnd.n7661 99.6594
R7493 gnd.n7657 gnd.n232 99.6594
R7494 gnd.n7655 gnd.n7654 99.6594
R7495 gnd.n7650 gnd.n239 99.6594
R7496 gnd.n7648 gnd.n7647 99.6594
R7497 gnd.n7640 gnd.n246 99.6594
R7498 gnd.n7638 gnd.n7637 99.6594
R7499 gnd.n7633 gnd.n253 99.6594
R7500 gnd.n7631 gnd.n7630 99.6594
R7501 gnd.n7626 gnd.n260 99.6594
R7502 gnd.n7624 gnd.n7623 99.6594
R7503 gnd.n7619 gnd.n267 99.6594
R7504 gnd.n7617 gnd.n7616 99.6594
R7505 gnd.n7612 gnd.n274 99.6594
R7506 gnd.n7610 gnd.n7609 99.6594
R7507 gnd.n284 gnd.n283 99.6594
R7508 gnd.n7601 gnd.n7600 99.6594
R7509 gnd.n7598 gnd.n7597 99.6594
R7510 gnd.n7593 gnd.n292 99.6594
R7511 gnd.n7591 gnd.n7590 99.6594
R7512 gnd.n7586 gnd.n299 99.6594
R7513 gnd.n7584 gnd.n7583 99.6594
R7514 gnd.n7579 gnd.n306 99.6594
R7515 gnd.n7577 gnd.n7576 99.6594
R7516 gnd.n7572 gnd.n315 99.6594
R7517 gnd.n7570 gnd.n7569 99.6594
R7518 gnd.n7204 gnd.n524 99.6594
R7519 gnd.n804 gnd.n530 99.6594
R7520 gnd.n808 gnd.n531 99.6594
R7521 gnd.n814 gnd.n532 99.6594
R7522 gnd.n818 gnd.n533 99.6594
R7523 gnd.n824 gnd.n534 99.6594
R7524 gnd.n828 gnd.n535 99.6594
R7525 gnd.n834 gnd.n536 99.6594
R7526 gnd.n838 gnd.n537 99.6594
R7527 gnd.n844 gnd.n538 99.6594
R7528 gnd.n846 gnd.n539 99.6594
R7529 gnd.n854 gnd.n540 99.6594
R7530 gnd.n856 gnd.n541 99.6594
R7531 gnd.n956 gnd.n543 99.6594
R7532 gnd.n952 gnd.n544 99.6594
R7533 gnd.n948 gnd.n545 99.6594
R7534 gnd.n944 gnd.n546 99.6594
R7535 gnd.n940 gnd.n547 99.6594
R7536 gnd.n936 gnd.n548 99.6594
R7537 gnd.n932 gnd.n549 99.6594
R7538 gnd.n928 gnd.n550 99.6594
R7539 gnd.n924 gnd.n551 99.6594
R7540 gnd.n920 gnd.n552 99.6594
R7541 gnd.n916 gnd.n553 99.6594
R7542 gnd.n912 gnd.n554 99.6594
R7543 gnd.n908 gnd.n555 99.6594
R7544 gnd.n904 gnd.n556 99.6594
R7545 gnd.n900 gnd.n557 99.6594
R7546 gnd.n5855 gnd.n5854 99.6594
R7547 gnd.n5850 gnd.n5775 99.6594
R7548 gnd.n5848 gnd.n5847 99.6594
R7549 gnd.n5843 gnd.n5782 99.6594
R7550 gnd.n5841 gnd.n5840 99.6594
R7551 gnd.n5836 gnd.n5789 99.6594
R7552 gnd.n5834 gnd.n5833 99.6594
R7553 gnd.n5829 gnd.n5796 99.6594
R7554 gnd.n5827 gnd.n5826 99.6594
R7555 gnd.n5822 gnd.n5806 99.6594
R7556 gnd.n5820 gnd.n5819 99.6594
R7557 gnd.n5815 gnd.n5812 99.6594
R7558 gnd.n1596 gnd.n1595 99.6594
R7559 gnd.n5923 gnd.n5922 99.6594
R7560 gnd.n5920 gnd.n5919 99.6594
R7561 gnd.n5915 gnd.n1605 99.6594
R7562 gnd.n5913 gnd.n5912 99.6594
R7563 gnd.n1615 gnd.n1614 99.6594
R7564 gnd.n5904 gnd.n5903 99.6594
R7565 gnd.n5901 gnd.n5900 99.6594
R7566 gnd.n5896 gnd.n1623 99.6594
R7567 gnd.n5894 gnd.n5893 99.6594
R7568 gnd.n5889 gnd.n1630 99.6594
R7569 gnd.n5887 gnd.n5886 99.6594
R7570 gnd.n5882 gnd.n1637 99.6594
R7571 gnd.n5880 gnd.n5879 99.6594
R7572 gnd.n5875 gnd.n1646 99.6594
R7573 gnd.n5873 gnd.n5872 99.6594
R7574 gnd.n5087 gnd.n5086 99.6594
R7575 gnd.n5081 gnd.n4775 99.6594
R7576 gnd.n5078 gnd.n4776 99.6594
R7577 gnd.n5074 gnd.n4777 99.6594
R7578 gnd.n5070 gnd.n4778 99.6594
R7579 gnd.n5066 gnd.n4779 99.6594
R7580 gnd.n5062 gnd.n4780 99.6594
R7581 gnd.n5058 gnd.n4781 99.6594
R7582 gnd.n5054 gnd.n4782 99.6594
R7583 gnd.n5049 gnd.n4783 99.6594
R7584 gnd.n5045 gnd.n4784 99.6594
R7585 gnd.n5041 gnd.n4785 99.6594
R7586 gnd.n5037 gnd.n4786 99.6594
R7587 gnd.n5033 gnd.n4787 99.6594
R7588 gnd.n5029 gnd.n4788 99.6594
R7589 gnd.n5025 gnd.n4789 99.6594
R7590 gnd.n5021 gnd.n4790 99.6594
R7591 gnd.n5017 gnd.n4791 99.6594
R7592 gnd.n5013 gnd.n4792 99.6594
R7593 gnd.n5009 gnd.n4793 99.6594
R7594 gnd.n5005 gnd.n4794 99.6594
R7595 gnd.n5001 gnd.n4795 99.6594
R7596 gnd.n4997 gnd.n4796 99.6594
R7597 gnd.n4993 gnd.n4797 99.6594
R7598 gnd.n4989 gnd.n4798 99.6594
R7599 gnd.n4985 gnd.n4799 99.6594
R7600 gnd.n4981 gnd.n4800 99.6594
R7601 gnd.n4977 gnd.n4801 99.6594
R7602 gnd.n5089 gnd.n1991 99.6594
R7603 gnd.n4765 gnd.n2014 99.6594
R7604 gnd.n4763 gnd.n2013 99.6594
R7605 gnd.n4759 gnd.n2012 99.6594
R7606 gnd.n4755 gnd.n2011 99.6594
R7607 gnd.n4751 gnd.n2010 99.6594
R7608 gnd.n4747 gnd.n2009 99.6594
R7609 gnd.n4743 gnd.n2008 99.6594
R7610 gnd.n4675 gnd.n2007 99.6594
R7611 gnd.n4006 gnd.n3737 99.6594
R7612 gnd.n3763 gnd.n3744 99.6594
R7613 gnd.n3765 gnd.n3745 99.6594
R7614 gnd.n3773 gnd.n3746 99.6594
R7615 gnd.n3775 gnd.n3747 99.6594
R7616 gnd.n3783 gnd.n3748 99.6594
R7617 gnd.n3785 gnd.n3749 99.6594
R7618 gnd.n3793 gnd.n3750 99.6594
R7619 gnd.n7561 gnd.n321 99.6594
R7620 gnd.n7559 gnd.n7558 99.6594
R7621 gnd.n7554 gnd.n328 99.6594
R7622 gnd.n7552 gnd.n7551 99.6594
R7623 gnd.n7547 gnd.n335 99.6594
R7624 gnd.n7545 gnd.n7544 99.6594
R7625 gnd.n7540 gnd.n342 99.6594
R7626 gnd.n7538 gnd.n7537 99.6594
R7627 gnd.n347 gnd.n346 99.6594
R7628 gnd.n605 gnd.n558 99.6594
R7629 gnd.n608 gnd.n559 99.6594
R7630 gnd.n616 gnd.n560 99.6594
R7631 gnd.n618 gnd.n561 99.6594
R7632 gnd.n626 gnd.n562 99.6594
R7633 gnd.n634 gnd.n563 99.6594
R7634 gnd.n636 gnd.n564 99.6594
R7635 gnd.n644 gnd.n565 99.6594
R7636 gnd.n7202 gnd.n7201 99.6594
R7637 gnd.n4733 gnd.n1994 99.6594
R7638 gnd.n4729 gnd.n1995 99.6594
R7639 gnd.n4725 gnd.n1996 99.6594
R7640 gnd.n4721 gnd.n1997 99.6594
R7641 gnd.n4717 gnd.n1998 99.6594
R7642 gnd.n4713 gnd.n1999 99.6594
R7643 gnd.n4709 gnd.n2000 99.6594
R7644 gnd.n4705 gnd.n2001 99.6594
R7645 gnd.n4701 gnd.n2002 99.6594
R7646 gnd.n4697 gnd.n2003 99.6594
R7647 gnd.n4693 gnd.n2004 99.6594
R7648 gnd.n4689 gnd.n2005 99.6594
R7649 gnd.n4685 gnd.n2006 99.6594
R7650 gnd.n3921 gnd.n3920 99.6594
R7651 gnd.n3915 gnd.n3832 99.6594
R7652 gnd.n3912 gnd.n3833 99.6594
R7653 gnd.n3908 gnd.n3834 99.6594
R7654 gnd.n3904 gnd.n3835 99.6594
R7655 gnd.n3900 gnd.n3836 99.6594
R7656 gnd.n3896 gnd.n3837 99.6594
R7657 gnd.n3892 gnd.n3838 99.6594
R7658 gnd.n3888 gnd.n3839 99.6594
R7659 gnd.n3884 gnd.n3840 99.6594
R7660 gnd.n3880 gnd.n3841 99.6594
R7661 gnd.n3876 gnd.n3842 99.6594
R7662 gnd.n3923 gnd.n3831 99.6594
R7663 gnd.n5610 gnd.n5609 99.6594
R7664 gnd.n5613 gnd.n5612 99.6594
R7665 gnd.n5624 gnd.n5623 99.6594
R7666 gnd.n5633 gnd.n5632 99.6594
R7667 gnd.n5636 gnd.n5635 99.6594
R7668 gnd.n5647 gnd.n5646 99.6594
R7669 gnd.n5656 gnd.n5655 99.6594
R7670 gnd.n5659 gnd.n5658 99.6594
R7671 gnd.n5664 gnd.n5663 99.6594
R7672 gnd.n4967 gnd.n4802 99.6594
R7673 gnd.n4964 gnd.n4803 99.6594
R7674 gnd.n4960 gnd.n4804 99.6594
R7675 gnd.n4956 gnd.n4805 99.6594
R7676 gnd.n4952 gnd.n4806 99.6594
R7677 gnd.n4948 gnd.n4807 99.6594
R7678 gnd.n4944 gnd.n4808 99.6594
R7679 gnd.n4940 gnd.n4809 99.6594
R7680 gnd.n4936 gnd.n4810 99.6594
R7681 gnd.n4965 gnd.n4802 99.6594
R7682 gnd.n4961 gnd.n4803 99.6594
R7683 gnd.n4957 gnd.n4804 99.6594
R7684 gnd.n4953 gnd.n4805 99.6594
R7685 gnd.n4949 gnd.n4806 99.6594
R7686 gnd.n4945 gnd.n4807 99.6594
R7687 gnd.n4941 gnd.n4808 99.6594
R7688 gnd.n4937 gnd.n4809 99.6594
R7689 gnd.n4892 gnd.n4810 99.6594
R7690 gnd.n5663 gnd.n5662 99.6594
R7691 gnd.n5658 gnd.n5657 99.6594
R7692 gnd.n5655 gnd.n5648 99.6594
R7693 gnd.n5646 gnd.n5645 99.6594
R7694 gnd.n5635 gnd.n5634 99.6594
R7695 gnd.n5632 gnd.n5625 99.6594
R7696 gnd.n5623 gnd.n5622 99.6594
R7697 gnd.n5612 gnd.n5611 99.6594
R7698 gnd.n5609 gnd.n5599 99.6594
R7699 gnd.n3921 gnd.n3844 99.6594
R7700 gnd.n3913 gnd.n3832 99.6594
R7701 gnd.n3909 gnd.n3833 99.6594
R7702 gnd.n3905 gnd.n3834 99.6594
R7703 gnd.n3901 gnd.n3835 99.6594
R7704 gnd.n3897 gnd.n3836 99.6594
R7705 gnd.n3893 gnd.n3837 99.6594
R7706 gnd.n3889 gnd.n3838 99.6594
R7707 gnd.n3885 gnd.n3839 99.6594
R7708 gnd.n3881 gnd.n3840 99.6594
R7709 gnd.n3877 gnd.n3841 99.6594
R7710 gnd.n3873 gnd.n3842 99.6594
R7711 gnd.n3924 gnd.n3923 99.6594
R7712 gnd.n4688 gnd.n2006 99.6594
R7713 gnd.n4692 gnd.n2005 99.6594
R7714 gnd.n4696 gnd.n2004 99.6594
R7715 gnd.n4700 gnd.n2003 99.6594
R7716 gnd.n4704 gnd.n2002 99.6594
R7717 gnd.n4708 gnd.n2001 99.6594
R7718 gnd.n4712 gnd.n2000 99.6594
R7719 gnd.n4716 gnd.n1999 99.6594
R7720 gnd.n4720 gnd.n1998 99.6594
R7721 gnd.n4724 gnd.n1997 99.6594
R7722 gnd.n4728 gnd.n1996 99.6594
R7723 gnd.n4732 gnd.n1995 99.6594
R7724 gnd.n2035 gnd.n1994 99.6594
R7725 gnd.n607 gnd.n558 99.6594
R7726 gnd.n615 gnd.n559 99.6594
R7727 gnd.n617 gnd.n560 99.6594
R7728 gnd.n625 gnd.n561 99.6594
R7729 gnd.n633 gnd.n562 99.6594
R7730 gnd.n635 gnd.n563 99.6594
R7731 gnd.n643 gnd.n564 99.6594
R7732 gnd.n567 gnd.n565 99.6594
R7733 gnd.n7202 gnd.n566 99.6594
R7734 gnd.n346 gnd.n343 99.6594
R7735 gnd.n7539 gnd.n7538 99.6594
R7736 gnd.n342 gnd.n336 99.6594
R7737 gnd.n7546 gnd.n7545 99.6594
R7738 gnd.n335 gnd.n329 99.6594
R7739 gnd.n7553 gnd.n7552 99.6594
R7740 gnd.n328 gnd.n322 99.6594
R7741 gnd.n7560 gnd.n7559 99.6594
R7742 gnd.n321 gnd.n318 99.6594
R7743 gnd.n4007 gnd.n4006 99.6594
R7744 gnd.n3766 gnd.n3744 99.6594
R7745 gnd.n3772 gnd.n3745 99.6594
R7746 gnd.n3776 gnd.n3746 99.6594
R7747 gnd.n3782 gnd.n3747 99.6594
R7748 gnd.n3786 gnd.n3748 99.6594
R7749 gnd.n3792 gnd.n3749 99.6594
R7750 gnd.n3750 gnd.n3734 99.6594
R7751 gnd.n4742 gnd.n2007 99.6594
R7752 gnd.n4746 gnd.n2008 99.6594
R7753 gnd.n4750 gnd.n2009 99.6594
R7754 gnd.n4754 gnd.n2010 99.6594
R7755 gnd.n4758 gnd.n2011 99.6594
R7756 gnd.n4762 gnd.n2012 99.6594
R7757 gnd.n4766 gnd.n2013 99.6594
R7758 gnd.n2016 gnd.n2014 99.6594
R7759 gnd.n5087 gnd.n4813 99.6594
R7760 gnd.n5079 gnd.n4775 99.6594
R7761 gnd.n5075 gnd.n4776 99.6594
R7762 gnd.n5071 gnd.n4777 99.6594
R7763 gnd.n5067 gnd.n4778 99.6594
R7764 gnd.n5063 gnd.n4779 99.6594
R7765 gnd.n5059 gnd.n4780 99.6594
R7766 gnd.n5055 gnd.n4781 99.6594
R7767 gnd.n5050 gnd.n4782 99.6594
R7768 gnd.n5046 gnd.n4783 99.6594
R7769 gnd.n5042 gnd.n4784 99.6594
R7770 gnd.n5038 gnd.n4785 99.6594
R7771 gnd.n5034 gnd.n4786 99.6594
R7772 gnd.n5030 gnd.n4787 99.6594
R7773 gnd.n5026 gnd.n4788 99.6594
R7774 gnd.n5022 gnd.n4789 99.6594
R7775 gnd.n5018 gnd.n4790 99.6594
R7776 gnd.n5014 gnd.n4791 99.6594
R7777 gnd.n5010 gnd.n4792 99.6594
R7778 gnd.n5006 gnd.n4793 99.6594
R7779 gnd.n5002 gnd.n4794 99.6594
R7780 gnd.n4998 gnd.n4795 99.6594
R7781 gnd.n4994 gnd.n4796 99.6594
R7782 gnd.n4990 gnd.n4797 99.6594
R7783 gnd.n4986 gnd.n4798 99.6594
R7784 gnd.n4982 gnd.n4799 99.6594
R7785 gnd.n4978 gnd.n4800 99.6594
R7786 gnd.n4974 gnd.n4801 99.6594
R7787 gnd.n5090 gnd.n5089 99.6594
R7788 gnd.n5874 gnd.n5873 99.6594
R7789 gnd.n1646 gnd.n1638 99.6594
R7790 gnd.n5881 gnd.n5880 99.6594
R7791 gnd.n1637 gnd.n1631 99.6594
R7792 gnd.n5888 gnd.n5887 99.6594
R7793 gnd.n1630 gnd.n1624 99.6594
R7794 gnd.n5895 gnd.n5894 99.6594
R7795 gnd.n1623 gnd.n1617 99.6594
R7796 gnd.n5902 gnd.n5901 99.6594
R7797 gnd.n5905 gnd.n5904 99.6594
R7798 gnd.n1614 gnd.n1606 99.6594
R7799 gnd.n5914 gnd.n5913 99.6594
R7800 gnd.n1605 gnd.n1599 99.6594
R7801 gnd.n5921 gnd.n5920 99.6594
R7802 gnd.n5924 gnd.n5923 99.6594
R7803 gnd.n5814 gnd.n5813 99.6594
R7804 gnd.n5812 gnd.n5807 99.6594
R7805 gnd.n5821 gnd.n5820 99.6594
R7806 gnd.n5806 gnd.n5797 99.6594
R7807 gnd.n5828 gnd.n5827 99.6594
R7808 gnd.n5796 gnd.n5790 99.6594
R7809 gnd.n5835 gnd.n5834 99.6594
R7810 gnd.n5789 gnd.n5783 99.6594
R7811 gnd.n5842 gnd.n5841 99.6594
R7812 gnd.n5782 gnd.n5776 99.6594
R7813 gnd.n5849 gnd.n5848 99.6594
R7814 gnd.n5775 gnd.n5770 99.6594
R7815 gnd.n5856 gnd.n5855 99.6594
R7816 gnd.n7205 gnd.n7204 99.6594
R7817 gnd.n807 gnd.n530 99.6594
R7818 gnd.n813 gnd.n531 99.6594
R7819 gnd.n817 gnd.n532 99.6594
R7820 gnd.n823 gnd.n533 99.6594
R7821 gnd.n827 gnd.n534 99.6594
R7822 gnd.n833 gnd.n535 99.6594
R7823 gnd.n837 gnd.n536 99.6594
R7824 gnd.n843 gnd.n537 99.6594
R7825 gnd.n847 gnd.n538 99.6594
R7826 gnd.n853 gnd.n539 99.6594
R7827 gnd.n857 gnd.n540 99.6594
R7828 gnd.n957 gnd.n542 99.6594
R7829 gnd.n953 gnd.n543 99.6594
R7830 gnd.n949 gnd.n544 99.6594
R7831 gnd.n945 gnd.n545 99.6594
R7832 gnd.n941 gnd.n546 99.6594
R7833 gnd.n937 gnd.n547 99.6594
R7834 gnd.n933 gnd.n548 99.6594
R7835 gnd.n929 gnd.n549 99.6594
R7836 gnd.n925 gnd.n550 99.6594
R7837 gnd.n921 gnd.n551 99.6594
R7838 gnd.n917 gnd.n552 99.6594
R7839 gnd.n913 gnd.n553 99.6594
R7840 gnd.n909 gnd.n554 99.6594
R7841 gnd.n905 gnd.n555 99.6594
R7842 gnd.n901 gnd.n556 99.6594
R7843 gnd.n893 gnd.n557 99.6594
R7844 gnd.n7571 gnd.n7570 99.6594
R7845 gnd.n315 gnd.n307 99.6594
R7846 gnd.n7578 gnd.n7577 99.6594
R7847 gnd.n306 gnd.n300 99.6594
R7848 gnd.n7585 gnd.n7584 99.6594
R7849 gnd.n299 gnd.n293 99.6594
R7850 gnd.n7592 gnd.n7591 99.6594
R7851 gnd.n292 gnd.n286 99.6594
R7852 gnd.n7599 gnd.n7598 99.6594
R7853 gnd.n7602 gnd.n7601 99.6594
R7854 gnd.n283 gnd.n275 99.6594
R7855 gnd.n7611 gnd.n7610 99.6594
R7856 gnd.n274 gnd.n268 99.6594
R7857 gnd.n7618 gnd.n7617 99.6594
R7858 gnd.n267 gnd.n261 99.6594
R7859 gnd.n7625 gnd.n7624 99.6594
R7860 gnd.n260 gnd.n254 99.6594
R7861 gnd.n7632 gnd.n7631 99.6594
R7862 gnd.n253 gnd.n247 99.6594
R7863 gnd.n7639 gnd.n7638 99.6594
R7864 gnd.n246 gnd.n240 99.6594
R7865 gnd.n7649 gnd.n7648 99.6594
R7866 gnd.n239 gnd.n233 99.6594
R7867 gnd.n7656 gnd.n7655 99.6594
R7868 gnd.n232 gnd.n226 99.6594
R7869 gnd.n7663 gnd.n7662 99.6594
R7870 gnd.n225 gnd.n219 99.6594
R7871 gnd.n7670 gnd.n7669 99.6594
R7872 gnd.n218 gnd.n215 99.6594
R7873 gnd.n5735 gnd.n5734 99.6594
R7874 gnd.n1709 gnd.n1689 99.6594
R7875 gnd.n1711 gnd.n1690 99.6594
R7876 gnd.n1713 gnd.n1691 99.6594
R7877 gnd.n5603 gnd.n1692 99.6594
R7878 gnd.n5606 gnd.n1693 99.6594
R7879 gnd.n5617 gnd.n1694 99.6594
R7880 gnd.n5619 gnd.n1695 99.6594
R7881 gnd.n5629 gnd.n1696 99.6594
R7882 gnd.n5640 gnd.n1697 99.6594
R7883 gnd.n5642 gnd.n1698 99.6594
R7884 gnd.n5652 gnd.n1699 99.6594
R7885 gnd.n5673 gnd.n1701 99.6594
R7886 gnd.n5737 gnd.n1686 99.6594
R7887 gnd.n5735 gnd.n1704 99.6594
R7888 gnd.n1710 gnd.n1689 99.6594
R7889 gnd.n1712 gnd.n1690 99.6594
R7890 gnd.n5602 gnd.n1691 99.6594
R7891 gnd.n5605 gnd.n1692 99.6594
R7892 gnd.n5616 gnd.n1693 99.6594
R7893 gnd.n5618 gnd.n1694 99.6594
R7894 gnd.n5628 gnd.n1695 99.6594
R7895 gnd.n5639 gnd.n1696 99.6594
R7896 gnd.n5641 gnd.n1697 99.6594
R7897 gnd.n5651 gnd.n1698 99.6594
R7898 gnd.n5672 gnd.n1699 99.6594
R7899 gnd.n1701 gnd.n1700 99.6594
R7900 gnd.n5738 gnd.n5737 99.6594
R7901 gnd.n648 gnd.n591 99.6594
R7902 gnd.n650 gnd.n649 99.6594
R7903 gnd.n651 gnd.n596 99.6594
R7904 gnd.n653 gnd.n652 99.6594
R7905 gnd.n654 gnd.n602 99.6594
R7906 gnd.n656 gnd.n611 99.6594
R7907 gnd.n658 gnd.n657 99.6594
R7908 gnd.n659 gnd.n622 99.6594
R7909 gnd.n661 gnd.n629 99.6594
R7910 gnd.n663 gnd.n662 99.6594
R7911 gnd.n664 gnd.n640 99.6594
R7912 gnd.n666 gnd.n646 99.6594
R7913 gnd.n667 gnd.n577 99.6594
R7914 gnd.n668 gnd.n579 99.6594
R7915 gnd.n666 gnd.n665 99.6594
R7916 gnd.n664 gnd.n639 99.6594
R7917 gnd.n663 gnd.n630 99.6594
R7918 gnd.n661 gnd.n660 99.6594
R7919 gnd.n659 gnd.n621 99.6594
R7920 gnd.n658 gnd.n612 99.6594
R7921 gnd.n656 gnd.n655 99.6594
R7922 gnd.n654 gnd.n601 99.6594
R7923 gnd.n653 gnd.n597 99.6594
R7924 gnd.n651 gnd.n595 99.6594
R7925 gnd.n650 gnd.n592 99.6594
R7926 gnd.n648 gnd.n587 99.6594
R7927 gnd.n668 gnd.n580 99.6594
R7928 gnd.n667 gnd.n578 99.6594
R7929 gnd.n5669 gnd.t127 98.63
R7930 gnd.n569 gnd.t80 98.63
R7931 gnd.n5660 gnd.t122 98.63
R7932 gnd.n792 gnd.t174 98.63
R7933 gnd.n872 gnd.t177 98.63
R7934 gnd.n895 gnd.t130 98.63
R7935 gnd.n312 gnd.t151 98.63
R7936 gnd.n279 gnd.t111 98.63
R7937 gnd.n7642 gnd.t148 98.63
R7938 gnd.n349 gnd.t97 98.63
R7939 gnd.n4832 gnd.t136 98.63
R7940 gnd.n4854 gnd.t139 98.63
R7941 gnd.n4875 gnd.t87 98.63
R7942 gnd.n4893 gnd.t164 98.63
R7943 gnd.n5798 gnd.t141 98.63
R7944 gnd.n1643 gnd.t166 98.63
R7945 gnd.n1610 gnd.t189 98.63
R7946 gnd.n574 gnd.t90 98.63
R7947 gnd.n1526 gnd.t180 96.6984
R7948 gnd.n962 gnd.t104 96.6984
R7949 gnd.n1528 gnd.t109 96.6906
R7950 gnd.n781 gnd.t160 96.6906
R7951 gnd.n2852 gnd.n2851 91.9545
R7952 gnd.n2851 gnd.n2515 91.9545
R7953 gnd.n2843 gnd.n2515 91.9545
R7954 gnd.n2843 gnd.n2842 91.9545
R7955 gnd.n2842 gnd.n2841 91.9545
R7956 gnd.n2841 gnd.n2523 91.9545
R7957 gnd.n2835 gnd.n2523 91.9545
R7958 gnd.n2835 gnd.n2834 91.9545
R7959 gnd.n2834 gnd.n2833 91.9545
R7960 gnd.n2833 gnd.n2530 91.9545
R7961 gnd.n2827 gnd.n2530 91.9545
R7962 gnd.n2827 gnd.n2826 91.9545
R7963 gnd.n2826 gnd.n2825 91.9545
R7964 gnd.n2825 gnd.n2538 91.9545
R7965 gnd.n2819 gnd.n2538 91.9545
R7966 gnd.n2819 gnd.n2818 91.9545
R7967 gnd.n2818 gnd.n2817 91.9545
R7968 gnd.n2817 gnd.n2546 91.9545
R7969 gnd.n2811 gnd.n2546 91.9545
R7970 gnd.n2811 gnd.n2810 91.9545
R7971 gnd.n2810 gnd.n2809 91.9545
R7972 gnd.n2809 gnd.n2554 91.9545
R7973 gnd.n2803 gnd.n2554 91.9545
R7974 gnd.n2803 gnd.n2802 91.9545
R7975 gnd.n2802 gnd.n2801 91.9545
R7976 gnd.n2801 gnd.n2562 91.9545
R7977 gnd.n2795 gnd.n2562 91.9545
R7978 gnd.n2795 gnd.n2794 91.9545
R7979 gnd.n2794 gnd.n2793 91.9545
R7980 gnd.n2793 gnd.n2570 91.9545
R7981 gnd.n2787 gnd.n2570 91.9545
R7982 gnd.n2787 gnd.n2786 91.9545
R7983 gnd.n2786 gnd.n2785 91.9545
R7984 gnd.n2785 gnd.n2578 91.9545
R7985 gnd.n2779 gnd.n2578 91.9545
R7986 gnd.n2779 gnd.n2778 91.9545
R7987 gnd.n2778 gnd.n2777 91.9545
R7988 gnd.n2777 gnd.n2586 91.9545
R7989 gnd.n2771 gnd.n2586 91.9545
R7990 gnd.n2771 gnd.n2770 91.9545
R7991 gnd.n2770 gnd.n2769 91.9545
R7992 gnd.n2769 gnd.n2594 91.9545
R7993 gnd.n2763 gnd.n2594 91.9545
R7994 gnd.n2763 gnd.n2762 91.9545
R7995 gnd.n2762 gnd.n2761 91.9545
R7996 gnd.n2761 gnd.n2602 91.9545
R7997 gnd.n2755 gnd.n2602 91.9545
R7998 gnd.n2755 gnd.n2754 91.9545
R7999 gnd.n2754 gnd.n2753 91.9545
R8000 gnd.n2753 gnd.n2610 91.9545
R8001 gnd.n2747 gnd.n2610 91.9545
R8002 gnd.n2747 gnd.n2746 91.9545
R8003 gnd.n2746 gnd.n2745 91.9545
R8004 gnd.n2745 gnd.n2618 91.9545
R8005 gnd.n2739 gnd.n2618 91.9545
R8006 gnd.n2739 gnd.n2738 91.9545
R8007 gnd.n2738 gnd.n2737 91.9545
R8008 gnd.n2737 gnd.n2626 91.9545
R8009 gnd.n2731 gnd.n2626 91.9545
R8010 gnd.n2731 gnd.n2730 91.9545
R8011 gnd.n2730 gnd.n2729 91.9545
R8012 gnd.n2729 gnd.n2634 91.9545
R8013 gnd.n2723 gnd.n2634 91.9545
R8014 gnd.n2723 gnd.n2722 91.9545
R8015 gnd.n2722 gnd.n2721 91.9545
R8016 gnd.n2721 gnd.n2642 91.9545
R8017 gnd.n2715 gnd.n2642 91.9545
R8018 gnd.n2715 gnd.n2714 91.9545
R8019 gnd.n2714 gnd.n2713 91.9545
R8020 gnd.n2713 gnd.n2650 91.9545
R8021 gnd.n2707 gnd.n2650 91.9545
R8022 gnd.n2707 gnd.n2706 91.9545
R8023 gnd.n2706 gnd.n2705 91.9545
R8024 gnd.n2705 gnd.n2658 91.9545
R8025 gnd.n2699 gnd.n2658 91.9545
R8026 gnd.n2699 gnd.n2698 91.9545
R8027 gnd.n2698 gnd.n2697 91.9545
R8028 gnd.n2697 gnd.n2666 91.9545
R8029 gnd.n2691 gnd.n2666 91.9545
R8030 gnd.n2691 gnd.n2690 91.9545
R8031 gnd.n2690 gnd.n2689 91.9545
R8032 gnd.n2689 gnd.n2674 91.9545
R8033 gnd.n2683 gnd.n2674 91.9545
R8034 gnd.n1480 gnd.n1479 81.8399
R8035 gnd.n3795 gnd.t115 74.8376
R8036 gnd.n2032 gnd.t146 74.8376
R8037 gnd.n1527 gnd.t179 72.8438
R8038 gnd.n963 gnd.t105 72.8438
R8039 gnd.n1481 gnd.n1474 72.8411
R8040 gnd.n1487 gnd.n1472 72.8411
R8041 gnd.n756 gnd.n755 72.8411
R8042 gnd.n5670 gnd.t126 72.836
R8043 gnd.n1529 gnd.t108 72.836
R8044 gnd.n782 gnd.t161 72.836
R8045 gnd.n570 gnd.t79 72.836
R8046 gnd.n5661 gnd.t123 72.836
R8047 gnd.n793 gnd.t173 72.836
R8048 gnd.n873 gnd.t176 72.836
R8049 gnd.n896 gnd.t129 72.836
R8050 gnd.n313 gnd.t152 72.836
R8051 gnd.n280 gnd.t112 72.836
R8052 gnd.n7643 gnd.t149 72.836
R8053 gnd.n350 gnd.t98 72.836
R8054 gnd.n4833 gnd.t135 72.836
R8055 gnd.n4855 gnd.t138 72.836
R8056 gnd.n4876 gnd.t86 72.836
R8057 gnd.n4894 gnd.t163 72.836
R8058 gnd.n5799 gnd.t142 72.836
R8059 gnd.n1644 gnd.t167 72.836
R8060 gnd.n1611 gnd.t190 72.836
R8061 gnd.n575 gnd.t91 72.836
R8062 gnd.n6996 gnd.n6995 71.676
R8063 gnd.n6993 gnd.n6992 71.676
R8064 gnd.n6988 gnd.n764 71.676
R8065 gnd.n6986 gnd.n6985 71.676
R8066 gnd.n6981 gnd.n767 71.676
R8067 gnd.n6979 gnd.n6978 71.676
R8068 gnd.n6974 gnd.n770 71.676
R8069 gnd.n6972 gnd.n6971 71.676
R8070 gnd.n6967 gnd.n773 71.676
R8071 gnd.n6965 gnd.n6964 71.676
R8072 gnd.n6960 gnd.n776 71.676
R8073 gnd.n6958 gnd.n6957 71.676
R8074 gnd.n6953 gnd.n779 71.676
R8075 gnd.n6951 gnd.n6950 71.676
R8076 gnd.n6945 gnd.n784 71.676
R8077 gnd.n6943 gnd.n6942 71.676
R8078 gnd.n6939 gnd.n6938 71.676
R8079 gnd.n6936 gnd.n6935 71.676
R8080 gnd.n6930 gnd.n965 71.676
R8081 gnd.n6928 gnd.n6927 71.676
R8082 gnd.n6923 gnd.n968 71.676
R8083 gnd.n6921 gnd.n6920 71.676
R8084 gnd.n6916 gnd.n971 71.676
R8085 gnd.n6914 gnd.n6913 71.676
R8086 gnd.n6909 gnd.n974 71.676
R8087 gnd.n6907 gnd.n6906 71.676
R8088 gnd.n6902 gnd.n977 71.676
R8089 gnd.n6900 gnd.n6899 71.676
R8090 gnd.n6895 gnd.n980 71.676
R8091 gnd.n6893 gnd.n6892 71.676
R8092 gnd.n6888 gnd.n983 71.676
R8093 gnd.n6886 gnd.n6885 71.676
R8094 gnd.n6881 gnd.n6877 71.676
R8095 gnd.n6002 gnd.n1469 71.676
R8096 gnd.n1531 gnd.n1494 71.676
R8097 gnd.n1535 gnd.n1495 71.676
R8098 gnd.n1539 gnd.n1496 71.676
R8099 gnd.n1543 gnd.n1497 71.676
R8100 gnd.n1547 gnd.n1498 71.676
R8101 gnd.n1551 gnd.n1499 71.676
R8102 gnd.n1555 gnd.n1500 71.676
R8103 gnd.n1559 gnd.n1501 71.676
R8104 gnd.n1563 gnd.n1502 71.676
R8105 gnd.n1567 gnd.n1503 71.676
R8106 gnd.n1571 gnd.n1504 71.676
R8107 gnd.n1575 gnd.n1505 71.676
R8108 gnd.n1579 gnd.n1506 71.676
R8109 gnd.n1583 gnd.n1507 71.676
R8110 gnd.n1587 gnd.n1508 71.676
R8111 gnd.n5933 gnd.n1510 71.676
R8112 gnd.n5937 gnd.n1511 71.676
R8113 gnd.n5942 gnd.n1512 71.676
R8114 gnd.n5946 gnd.n1513 71.676
R8115 gnd.n5950 gnd.n1514 71.676
R8116 gnd.n5954 gnd.n1515 71.676
R8117 gnd.n5958 gnd.n1516 71.676
R8118 gnd.n5962 gnd.n1517 71.676
R8119 gnd.n5966 gnd.n1518 71.676
R8120 gnd.n5970 gnd.n1519 71.676
R8121 gnd.n5974 gnd.n1520 71.676
R8122 gnd.n5978 gnd.n1521 71.676
R8123 gnd.n5982 gnd.n1522 71.676
R8124 gnd.n5986 gnd.n1523 71.676
R8125 gnd.n5990 gnd.n1524 71.676
R8126 gnd.n6000 gnd.n1525 71.676
R8127 gnd.n6003 gnd.n6002 71.676
R8128 gnd.n1534 gnd.n1494 71.676
R8129 gnd.n1538 gnd.n1495 71.676
R8130 gnd.n1542 gnd.n1496 71.676
R8131 gnd.n1546 gnd.n1497 71.676
R8132 gnd.n1550 gnd.n1498 71.676
R8133 gnd.n1554 gnd.n1499 71.676
R8134 gnd.n1558 gnd.n1500 71.676
R8135 gnd.n1562 gnd.n1501 71.676
R8136 gnd.n1566 gnd.n1502 71.676
R8137 gnd.n1570 gnd.n1503 71.676
R8138 gnd.n1574 gnd.n1504 71.676
R8139 gnd.n1578 gnd.n1505 71.676
R8140 gnd.n1582 gnd.n1506 71.676
R8141 gnd.n1586 gnd.n1507 71.676
R8142 gnd.n5932 gnd.n1509 71.676
R8143 gnd.n5936 gnd.n1510 71.676
R8144 gnd.n5941 gnd.n1511 71.676
R8145 gnd.n5945 gnd.n1512 71.676
R8146 gnd.n5949 gnd.n1513 71.676
R8147 gnd.n5953 gnd.n1514 71.676
R8148 gnd.n5957 gnd.n1515 71.676
R8149 gnd.n5961 gnd.n1516 71.676
R8150 gnd.n5965 gnd.n1517 71.676
R8151 gnd.n5969 gnd.n1518 71.676
R8152 gnd.n5973 gnd.n1519 71.676
R8153 gnd.n5977 gnd.n1520 71.676
R8154 gnd.n5981 gnd.n1521 71.676
R8155 gnd.n5985 gnd.n1522 71.676
R8156 gnd.n5989 gnd.n1523 71.676
R8157 gnd.n5992 gnd.n1524 71.676
R8158 gnd.n6000 gnd.n5999 71.676
R8159 gnd.n6877 gnd.n984 71.676
R8160 gnd.n6887 gnd.n6886 71.676
R8161 gnd.n983 gnd.n981 71.676
R8162 gnd.n6894 gnd.n6893 71.676
R8163 gnd.n980 gnd.n978 71.676
R8164 gnd.n6901 gnd.n6900 71.676
R8165 gnd.n977 gnd.n975 71.676
R8166 gnd.n6908 gnd.n6907 71.676
R8167 gnd.n974 gnd.n972 71.676
R8168 gnd.n6915 gnd.n6914 71.676
R8169 gnd.n971 gnd.n969 71.676
R8170 gnd.n6922 gnd.n6921 71.676
R8171 gnd.n968 gnd.n966 71.676
R8172 gnd.n6929 gnd.n6928 71.676
R8173 gnd.n965 gnd.n961 71.676
R8174 gnd.n6937 gnd.n6936 71.676
R8175 gnd.n960 gnd.n785 71.676
R8176 gnd.n6944 gnd.n6943 71.676
R8177 gnd.n784 gnd.n780 71.676
R8178 gnd.n6952 gnd.n6951 71.676
R8179 gnd.n779 gnd.n777 71.676
R8180 gnd.n6959 gnd.n6958 71.676
R8181 gnd.n776 gnd.n774 71.676
R8182 gnd.n6966 gnd.n6965 71.676
R8183 gnd.n773 gnd.n771 71.676
R8184 gnd.n6973 gnd.n6972 71.676
R8185 gnd.n770 gnd.n768 71.676
R8186 gnd.n6980 gnd.n6979 71.676
R8187 gnd.n767 gnd.n765 71.676
R8188 gnd.n6987 gnd.n6986 71.676
R8189 gnd.n764 gnd.n762 71.676
R8190 gnd.n6994 gnd.n6993 71.676
R8191 gnd.n6997 gnd.n6996 71.676
R8192 gnd.n10 gnd.t58 69.1507
R8193 gnd.n18 gnd.t356 68.4792
R8194 gnd.n17 gnd.t375 68.4792
R8195 gnd.n16 gnd.t53 68.4792
R8196 gnd.n15 gnd.t15 68.4792
R8197 gnd.n14 gnd.t368 68.4792
R8198 gnd.n13 gnd.t69 68.4792
R8199 gnd.n12 gnd.t46 68.4792
R8200 gnd.n11 gnd.t354 68.4792
R8201 gnd.n10 gnd.t1 68.4792
R8202 gnd.n3922 gnd.n3826 64.369
R8203 gnd.n5939 gnd.n1527 59.5399
R8204 gnd.n6932 gnd.n963 59.5399
R8205 gnd.n1530 gnd.n1529 59.5399
R8206 gnd.n6947 gnd.n782 59.5399
R8207 gnd.n6006 gnd.n1490 59.1804
R8208 gnd.n4774 gnd.n1992 57.3586
R8209 gnd.n5088 gnd.n1979 57.3586
R8210 gnd.n7679 gnd.n211 57.3586
R8211 gnd.n3577 gnd.t314 56.407
R8212 gnd.n3530 gnd.t334 56.407
R8213 gnd.n3545 gnd.t298 56.407
R8214 gnd.n3561 gnd.t210 56.407
R8215 gnd.n68 gnd.t292 56.407
R8216 gnd.n21 gnd.t219 56.407
R8217 gnd.n36 gnd.t280 56.407
R8218 gnd.n52 gnd.t326 56.407
R8219 gnd.n3590 gnd.t271 55.8337
R8220 gnd.n3543 gnd.t227 55.8337
R8221 gnd.n3558 gnd.t250 55.8337
R8222 gnd.n3574 gnd.t319 55.8337
R8223 gnd.n81 gnd.t330 55.8337
R8224 gnd.n34 gnd.t244 55.8337
R8225 gnd.n49 gnd.t349 55.8337
R8226 gnd.n65 gnd.t248 55.8337
R8227 gnd.n2683 gnd.n171 55.1729
R8228 gnd.n1478 gnd.n1477 54.358
R8229 gnd.n753 gnd.n752 54.358
R8230 gnd.n3577 gnd.n3576 53.0052
R8231 gnd.n3579 gnd.n3578 53.0052
R8232 gnd.n3581 gnd.n3580 53.0052
R8233 gnd.n3583 gnd.n3582 53.0052
R8234 gnd.n3585 gnd.n3584 53.0052
R8235 gnd.n3587 gnd.n3586 53.0052
R8236 gnd.n3589 gnd.n3588 53.0052
R8237 gnd.n3530 gnd.n3529 53.0052
R8238 gnd.n3532 gnd.n3531 53.0052
R8239 gnd.n3534 gnd.n3533 53.0052
R8240 gnd.n3536 gnd.n3535 53.0052
R8241 gnd.n3538 gnd.n3537 53.0052
R8242 gnd.n3540 gnd.n3539 53.0052
R8243 gnd.n3542 gnd.n3541 53.0052
R8244 gnd.n3545 gnd.n3544 53.0052
R8245 gnd.n3547 gnd.n3546 53.0052
R8246 gnd.n3549 gnd.n3548 53.0052
R8247 gnd.n3551 gnd.n3550 53.0052
R8248 gnd.n3553 gnd.n3552 53.0052
R8249 gnd.n3555 gnd.n3554 53.0052
R8250 gnd.n3557 gnd.n3556 53.0052
R8251 gnd.n3561 gnd.n3560 53.0052
R8252 gnd.n3563 gnd.n3562 53.0052
R8253 gnd.n3565 gnd.n3564 53.0052
R8254 gnd.n3567 gnd.n3566 53.0052
R8255 gnd.n3569 gnd.n3568 53.0052
R8256 gnd.n3571 gnd.n3570 53.0052
R8257 gnd.n3573 gnd.n3572 53.0052
R8258 gnd.n80 gnd.n79 53.0052
R8259 gnd.n78 gnd.n77 53.0052
R8260 gnd.n76 gnd.n75 53.0052
R8261 gnd.n74 gnd.n73 53.0052
R8262 gnd.n72 gnd.n71 53.0052
R8263 gnd.n70 gnd.n69 53.0052
R8264 gnd.n68 gnd.n67 53.0052
R8265 gnd.n33 gnd.n32 53.0052
R8266 gnd.n31 gnd.n30 53.0052
R8267 gnd.n29 gnd.n28 53.0052
R8268 gnd.n27 gnd.n26 53.0052
R8269 gnd.n25 gnd.n24 53.0052
R8270 gnd.n23 gnd.n22 53.0052
R8271 gnd.n21 gnd.n20 53.0052
R8272 gnd.n48 gnd.n47 53.0052
R8273 gnd.n46 gnd.n45 53.0052
R8274 gnd.n44 gnd.n43 53.0052
R8275 gnd.n42 gnd.n41 53.0052
R8276 gnd.n40 gnd.n39 53.0052
R8277 gnd.n38 gnd.n37 53.0052
R8278 gnd.n36 gnd.n35 53.0052
R8279 gnd.n64 gnd.n63 53.0052
R8280 gnd.n62 gnd.n61 53.0052
R8281 gnd.n60 gnd.n59 53.0052
R8282 gnd.n58 gnd.n57 53.0052
R8283 gnd.n56 gnd.n55 53.0052
R8284 gnd.n54 gnd.n53 53.0052
R8285 gnd.n52 gnd.n51 53.0052
R8286 gnd.n744 gnd.n743 52.4801
R8287 gnd.n4626 gnd.t371 52.3082
R8288 gnd.n4594 gnd.t50 52.3082
R8289 gnd.n4562 gnd.t366 52.3082
R8290 gnd.n4531 gnd.t362 52.3082
R8291 gnd.n4499 gnd.t373 52.3082
R8292 gnd.n4467 gnd.t44 52.3082
R8293 gnd.n4435 gnd.t352 52.3082
R8294 gnd.n4404 gnd.t34 52.3082
R8295 gnd.n4456 gnd.n4424 51.4173
R8296 gnd.n4520 gnd.n4519 50.455
R8297 gnd.n4488 gnd.n4487 50.455
R8298 gnd.n4456 gnd.n4455 50.455
R8299 gnd.n3869 gnd.n3868 45.1884
R8300 gnd.n2058 gnd.n2057 45.1884
R8301 gnd.n6999 gnd.n759 44.3322
R8302 gnd.n1481 gnd.n1480 44.3189
R8303 gnd.n5671 gnd.n5670 42.4732
R8304 gnd.n576 gnd.n575 42.4732
R8305 gnd.n571 gnd.n570 42.2793
R8306 gnd.n3870 gnd.n3869 42.2793
R8307 gnd.n2059 gnd.n2058 42.2793
R8308 gnd.n3796 gnd.n3795 42.2793
R8309 gnd.n4741 gnd.n2032 42.2793
R8310 gnd.n5666 gnd.n5661 42.2793
R8311 gnd.n794 gnd.n793 42.2793
R8312 gnd.n939 gnd.n873 42.2793
R8313 gnd.n899 gnd.n896 42.2793
R8314 gnd.n314 gnd.n313 42.2793
R8315 gnd.n7607 gnd.n280 42.2793
R8316 gnd.n7644 gnd.n7643 42.2793
R8317 gnd.n7535 gnd.n350 42.2793
R8318 gnd.n5052 gnd.n4833 42.2793
R8319 gnd.n5012 gnd.n4855 42.2793
R8320 gnd.n4973 gnd.n4876 42.2793
R8321 gnd.n4895 gnd.n4894 42.2793
R8322 gnd.n5800 gnd.n5799 42.2793
R8323 gnd.n1645 gnd.n1644 42.2793
R8324 gnd.n5910 gnd.n1611 42.2793
R8325 gnd.n1479 gnd.n1478 41.6274
R8326 gnd.n754 gnd.n753 41.6274
R8327 gnd.n1488 gnd.n1487 40.8975
R8328 gnd.n757 gnd.n756 40.8975
R8329 gnd.n1487 gnd.n1486 35.055
R8330 gnd.n1482 gnd.n1481 35.055
R8331 gnd.n746 gnd.n745 35.055
R8332 gnd.n756 gnd.n742 35.055
R8333 gnd.n3167 gnd.n3166 32.9544
R8334 gnd.n3167 gnd.n2201 32.9544
R8335 gnd.n3175 gnd.n2201 32.9544
R8336 gnd.n3176 gnd.n3175 32.9544
R8337 gnd.n3177 gnd.n3176 32.9544
R8338 gnd.n3177 gnd.n2195 32.9544
R8339 gnd.n3185 gnd.n2195 32.9544
R8340 gnd.n3186 gnd.n3185 32.9544
R8341 gnd.n3187 gnd.n3186 32.9544
R8342 gnd.n3187 gnd.n2189 32.9544
R8343 gnd.n3195 gnd.n2189 32.9544
R8344 gnd.n3196 gnd.n3195 32.9544
R8345 gnd.n3197 gnd.n3196 32.9544
R8346 gnd.n3197 gnd.n2183 32.9544
R8347 gnd.n3205 gnd.n2183 32.9544
R8348 gnd.n3206 gnd.n3205 32.9544
R8349 gnd.n3207 gnd.n3206 32.9544
R8350 gnd.n3207 gnd.n2177 32.9544
R8351 gnd.n3215 gnd.n2177 32.9544
R8352 gnd.n3216 gnd.n3215 32.9544
R8353 gnd.n3217 gnd.n3216 32.9544
R8354 gnd.n3217 gnd.n2171 32.9544
R8355 gnd.n3225 gnd.n2171 32.9544
R8356 gnd.n3226 gnd.n3225 32.9544
R8357 gnd.n3227 gnd.n3226 32.9544
R8358 gnd.n3227 gnd.n2165 32.9544
R8359 gnd.n3235 gnd.n2165 32.9544
R8360 gnd.n3236 gnd.n3235 32.9544
R8361 gnd.n3237 gnd.n3236 32.9544
R8362 gnd.n3237 gnd.n2159 32.9544
R8363 gnd.n3245 gnd.n2159 32.9544
R8364 gnd.n3246 gnd.n3245 32.9544
R8365 gnd.n3247 gnd.n3246 32.9544
R8366 gnd.n3247 gnd.n2153 32.9544
R8367 gnd.n3255 gnd.n2153 32.9544
R8368 gnd.n3256 gnd.n3255 32.9544
R8369 gnd.n3257 gnd.n3256 32.9544
R8370 gnd.n3257 gnd.n2147 32.9544
R8371 gnd.n3265 gnd.n2147 32.9544
R8372 gnd.n3266 gnd.n3265 32.9544
R8373 gnd.n3267 gnd.n3266 32.9544
R8374 gnd.n3267 gnd.n2141 32.9544
R8375 gnd.n3275 gnd.n2141 32.9544
R8376 gnd.n3276 gnd.n3275 32.9544
R8377 gnd.n3277 gnd.n3276 32.9544
R8378 gnd.n3277 gnd.n2135 32.9544
R8379 gnd.n3285 gnd.n2135 32.9544
R8380 gnd.n3286 gnd.n3285 32.9544
R8381 gnd.n3287 gnd.n3286 32.9544
R8382 gnd.n3287 gnd.n2129 32.9544
R8383 gnd.n3295 gnd.n2129 32.9544
R8384 gnd.n3296 gnd.n3295 32.9544
R8385 gnd.n3297 gnd.n3296 32.9544
R8386 gnd.n3297 gnd.n2123 32.9544
R8387 gnd.n3305 gnd.n2123 32.9544
R8388 gnd.n3306 gnd.n3305 32.9544
R8389 gnd.n3307 gnd.n3306 32.9544
R8390 gnd.n3307 gnd.n2117 32.9544
R8391 gnd.n3315 gnd.n2117 32.9544
R8392 gnd.n3316 gnd.n3315 32.9544
R8393 gnd.n3317 gnd.n3316 32.9544
R8394 gnd.n3317 gnd.n2111 32.9544
R8395 gnd.n3325 gnd.n2111 32.9544
R8396 gnd.n3326 gnd.n3325 32.9544
R8397 gnd.n3327 gnd.n3326 32.9544
R8398 gnd.n3327 gnd.n2105 32.9544
R8399 gnd.n3335 gnd.n2105 32.9544
R8400 gnd.n3336 gnd.n3335 32.9544
R8401 gnd.n3337 gnd.n3336 32.9544
R8402 gnd.n3337 gnd.n2099 32.9544
R8403 gnd.n3345 gnd.n2099 32.9544
R8404 gnd.n3346 gnd.n3345 32.9544
R8405 gnd.n3347 gnd.n3346 32.9544
R8406 gnd.n3347 gnd.n2093 32.9544
R8407 gnd.n3355 gnd.n2093 32.9544
R8408 gnd.n3356 gnd.n3355 32.9544
R8409 gnd.n3357 gnd.n3356 32.9544
R8410 gnd.n3357 gnd.n2087 32.9544
R8411 gnd.n3365 gnd.n2087 32.9544
R8412 gnd.n3366 gnd.n3365 32.9544
R8413 gnd.n3367 gnd.n3366 32.9544
R8414 gnd.n3367 gnd.n2074 32.9544
R8415 gnd.n3377 gnd.n2074 32.9544
R8416 gnd.n6882 gnd.n6876 32.9371
R8417 gnd.n5998 gnd.n5997 32.9371
R8418 gnd.n3932 gnd.n3826 31.8661
R8419 gnd.n3932 gnd.n3931 31.8661
R8420 gnd.n3940 gnd.n3815 31.8661
R8421 gnd.n3948 gnd.n3815 31.8661
R8422 gnd.n3948 gnd.n3809 31.8661
R8423 gnd.n3956 gnd.n3809 31.8661
R8424 gnd.n3956 gnd.n3802 31.8661
R8425 gnd.n3994 gnd.n3802 31.8661
R8426 gnd.n4004 gnd.n3735 31.8661
R8427 gnd.n5098 gnd.n1979 31.8661
R8428 gnd.n5106 gnd.n1971 31.8661
R8429 gnd.n5106 gnd.n1960 31.8661
R8430 gnd.n5118 gnd.n1960 31.8661
R8431 gnd.n5118 gnd.n1963 31.8661
R8432 gnd.n5126 gnd.n1943 31.8661
R8433 gnd.n5138 gnd.n1943 31.8661
R8434 gnd.n5146 gnd.n1935 31.8661
R8435 gnd.n5162 gnd.n1923 31.8661
R8436 gnd.n5162 gnd.n1926 31.8661
R8437 gnd.n5172 gnd.n1909 31.8661
R8438 gnd.n5182 gnd.n1909 31.8661
R8439 gnd.n5197 gnd.n1900 31.8661
R8440 gnd.n5207 gnd.n1884 31.8661
R8441 gnd.n5226 gnd.n1884 31.8661
R8442 gnd.n5237 gnd.n1870 31.8661
R8443 gnd.n5242 gnd.n1870 31.8661
R8444 gnd.n5255 gnd.n1862 31.8661
R8445 gnd.n5261 gnd.n1850 31.8661
R8446 gnd.n5270 gnd.n1850 31.8661
R8447 gnd.n5589 gnd.n5588 31.8661
R8448 gnd.n5589 gnd.n1688 31.8661
R8449 gnd.n5448 gnd.n1702 31.8661
R8450 gnd.n647 gnd.n585 31.8661
R8451 gnd.n7123 gnd.n669 31.8661
R8452 gnd.n669 gnd.n529 31.8661
R8453 gnd.n7411 gnd.n370 31.8661
R8454 gnd.n7419 gnd.n370 31.8661
R8455 gnd.n7428 gnd.n364 31.8661
R8456 gnd.n7753 gnd.n90 31.8661
R8457 gnd.n7472 gnd.n90 31.8661
R8458 gnd.n7745 gnd.n107 31.8661
R8459 gnd.n7739 gnd.n107 31.8661
R8460 gnd.n7733 gnd.n124 31.8661
R8461 gnd.n7727 gnd.n133 31.8661
R8462 gnd.n7727 gnd.n136 31.8661
R8463 gnd.n7721 gnd.n146 31.8661
R8464 gnd.n7715 gnd.n146 31.8661
R8465 gnd.n7709 gnd.n162 31.8661
R8466 gnd.n7703 gnd.n174 31.8661
R8467 gnd.n7697 gnd.n184 31.8661
R8468 gnd.n7691 gnd.n184 31.8661
R8469 gnd.n7691 gnd.n193 31.8661
R8470 gnd.n7685 gnd.n193 31.8661
R8471 gnd.n7679 gnd.n208 31.8661
R8472 gnd.n5274 gnd.n1821 29.3168
R8473 gnd.n5313 gnd.n1813 29.3168
R8474 gnd.n5333 gnd.n1798 29.3168
R8475 gnd.n5279 gnd.n1786 29.3168
R8476 gnd.n5326 gnd.n1779 29.3168
R8477 gnd.n5352 gnd.n1760 29.3168
R8478 gnd.n5359 gnd.n1751 29.3168
R8479 gnd.n5374 gnd.n1744 29.3168
R8480 gnd.n5403 gnd.n1733 29.3168
R8481 gnd.n5424 gnd.n1726 29.3168
R8482 gnd.n5423 gnd.n1674 29.3168
R8483 gnd.n5752 gnd.n1664 29.3168
R8484 gnd.n5762 gnd.n1667 29.3168
R8485 gnd.n5864 gnd.n1656 29.3168
R8486 gnd.n5596 gnd.n5595 29.3168
R8487 gnd.n7214 gnd.n520 29.3168
R8488 gnd.n7097 gnd.n522 29.3168
R8489 gnd.n7241 gnd.n501 29.3168
R8490 gnd.n7227 gnd.n504 29.3168
R8491 gnd.n7251 gnd.n491 29.3168
R8492 gnd.n493 gnd.n483 29.3168
R8493 gnd.n7287 gnd.n466 29.3168
R8494 gnd.n7273 gnd.n469 29.3168
R8495 gnd.n458 gnd.n449 29.3168
R8496 gnd.n7334 gnd.n431 29.3168
R8497 gnd.n7319 gnd.n434 29.3168
R8498 gnd.n7327 gnd.n423 29.3168
R8499 gnd.n7353 gnd.n414 29.3168
R8500 gnd.n7365 gnd.n401 29.3168
R8501 gnd.n7371 gnd.n391 29.3168
R8502 gnd.n5274 gnd.n1839 28.3609
R8503 gnd.n7371 gnd.n383 28.3609
R8504 gnd.n5595 gnd.n1597 28.0422
R8505 gnd.n7203 gnd.n520 28.0422
R8506 gnd.n5146 gnd.t203 27.7236
R8507 gnd.n162 gnd.t277 27.7236
R8508 gnd.n1900 gnd.t201 27.0862
R8509 gnd.n124 gnd.t231 27.0862
R8510 gnd.t272 gnd.n1862 26.4489
R8511 gnd.n5255 gnd.t224 26.4489
R8512 gnd.t233 gnd.n364 26.4489
R8513 gnd.n7428 gnd.t207 26.4489
R8514 gnd.n5197 gnd.t239 25.8116
R8515 gnd.n5312 gnd.t255 25.8116
R8516 gnd.n7378 gnd.t191 25.8116
R8517 gnd.n7733 gnd.t197 25.8116
R8518 gnd.n5670 gnd.n5669 25.7944
R8519 gnd.n570 gnd.n569 25.7944
R8520 gnd.n3795 gnd.n3794 25.7944
R8521 gnd.n2032 gnd.n2031 25.7944
R8522 gnd.n5661 gnd.n5660 25.7944
R8523 gnd.n793 gnd.n792 25.7944
R8524 gnd.n873 gnd.n872 25.7944
R8525 gnd.n896 gnd.n895 25.7944
R8526 gnd.n313 gnd.n312 25.7944
R8527 gnd.n280 gnd.n279 25.7944
R8528 gnd.n7643 gnd.n7642 25.7944
R8529 gnd.n350 gnd.n349 25.7944
R8530 gnd.n4833 gnd.n4832 25.7944
R8531 gnd.n4855 gnd.n4854 25.7944
R8532 gnd.n4876 gnd.n4875 25.7944
R8533 gnd.n4894 gnd.n4893 25.7944
R8534 gnd.n5799 gnd.n5798 25.7944
R8535 gnd.n1644 gnd.n1643 25.7944
R8536 gnd.n1611 gnd.n1610 25.7944
R8537 gnd.n575 gnd.n574 25.7944
R8538 gnd.t229 gnd.n1935 25.1743
R8539 gnd.n5360 gnd.t195 25.1743
R8540 gnd.n5391 gnd.t274 25.1743
R8541 gnd.n7297 gnd.t222 25.1743
R8542 gnd.n7307 gnd.t236 25.1743
R8543 gnd.n7709 gnd.t220 25.1743
R8544 gnd.n4016 gnd.n3736 24.8557
R8545 gnd.n4026 gnd.n3719 24.8557
R8546 gnd.n3722 gnd.n3710 24.8557
R8547 gnd.n4047 gnd.n3711 24.8557
R8548 gnd.n4057 gnd.n3691 24.8557
R8549 gnd.n4067 gnd.n4066 24.8557
R8550 gnd.n3677 gnd.n3675 24.8557
R8551 gnd.n4098 gnd.n4097 24.8557
R8552 gnd.n4113 gnd.n3660 24.8557
R8553 gnd.n4167 gnd.n3599 24.8557
R8554 gnd.n4123 gnd.n3600 24.8557
R8555 gnd.n4160 gnd.n3611 24.8557
R8556 gnd.n3649 gnd.n3648 24.8557
R8557 gnd.n4154 gnd.n4153 24.8557
R8558 gnd.n3635 gnd.n3622 24.8557
R8559 gnd.n4193 gnd.n4192 24.8557
R8560 gnd.n4203 gnd.n3515 24.8557
R8561 gnd.n4215 gnd.n3507 24.8557
R8562 gnd.n4214 gnd.n3495 24.8557
R8563 gnd.n4233 gnd.n4232 24.8557
R8564 gnd.n4243 gnd.n3488 24.8557
R8565 gnd.n4254 gnd.n3476 24.8557
R8566 gnd.n4278 gnd.n4277 24.8557
R8567 gnd.n4289 gnd.n3459 24.8557
R8568 gnd.n4288 gnd.n3461 24.8557
R8569 gnd.n4300 gnd.n3452 24.8557
R8570 gnd.n4318 gnd.n4317 24.8557
R8571 gnd.n3443 gnd.n3432 24.8557
R8572 gnd.n4339 gnd.n3420 24.8557
R8573 gnd.n4367 gnd.n4366 24.8557
R8574 gnd.n4378 gnd.n3405 24.8557
R8575 gnd.n4389 gnd.n3398 24.8557
R8576 gnd.n4388 gnd.n3386 24.8557
R8577 gnd.n4661 gnd.n4660 24.8557
R8578 gnd.n4683 gnd.n2066 24.8557
R8579 gnd.t213 gnd.n1823 24.537
R8580 gnd.n7364 gnd.t259 24.537
R8581 gnd.n5736 gnd.n1688 23.8997
R8582 gnd.n7124 gnd.n7123 23.8997
R8583 gnd.n1527 gnd.n1526 23.855
R8584 gnd.n963 gnd.n962 23.855
R8585 gnd.n1529 gnd.n1528 23.855
R8586 gnd.n782 gnd.n781 23.855
R8587 gnd.n4037 gnd.t33 23.2624
R8588 gnd.n3738 gnd.t114 22.6251
R8589 gnd.n5098 gnd.t85 22.6251
R8590 gnd.n208 gnd.t96 22.6251
R8591 gnd.t361 gnd.n3743 21.3504
R8592 gnd.n6008 gnd.n6006 20.7615
R8593 gnd.n7000 gnd.n6999 20.7615
R8594 gnd.t20 gnd.n3433 20.7131
R8595 gnd.t39 gnd.n3468 20.0758
R8596 gnd.t121 gnd.n1654 20.0758
R8597 gnd.n7098 gnd.t78 20.0758
R8598 gnd.n1476 gnd.t76 19.8005
R8599 gnd.n1476 gnd.t101 19.8005
R8600 gnd.n1475 gnd.t183 19.8005
R8601 gnd.n1475 gnd.t83 19.8005
R8602 gnd.n751 gnd.t133 19.8005
R8603 gnd.n751 gnd.t73 19.8005
R8604 gnd.n750 gnd.t119 19.8005
R8605 gnd.n750 gnd.t94 19.8005
R8606 gnd.n3378 gnd.n3377 19.7728
R8607 gnd.n1472 gnd.n1471 19.5087
R8608 gnd.n1485 gnd.n1472 19.5087
R8609 gnd.n1483 gnd.n1474 19.5087
R8610 gnd.n755 gnd.n749 19.5087
R8611 gnd.n4204 gnd.t30 19.4385
R8612 gnd.n5505 gnd.n5504 19.3944
R8613 gnd.n5505 gnd.n5502 19.3944
R8614 gnd.n5509 gnd.n5502 19.3944
R8615 gnd.n5509 gnd.n5487 19.3944
R8616 gnd.n5524 gnd.n5487 19.3944
R8617 gnd.n5524 gnd.n5485 19.3944
R8618 gnd.n5528 gnd.n5485 19.3944
R8619 gnd.n5528 gnd.n5474 19.3944
R8620 gnd.n5545 gnd.n5474 19.3944
R8621 gnd.n5545 gnd.n5471 19.3944
R8622 gnd.n5556 gnd.n5471 19.3944
R8623 gnd.n5556 gnd.n5472 19.3944
R8624 gnd.n5552 gnd.n5472 19.3944
R8625 gnd.n5552 gnd.n5551 19.3944
R8626 gnd.n5551 gnd.n5550 19.3944
R8627 gnd.n5550 gnd.n1450 19.3944
R8628 gnd.n6033 gnd.n1450 19.3944
R8629 gnd.n6033 gnd.n1447 19.3944
R8630 gnd.n6044 gnd.n1447 19.3944
R8631 gnd.n6044 gnd.n1448 19.3944
R8632 gnd.n6040 gnd.n1448 19.3944
R8633 gnd.n6040 gnd.n6039 19.3944
R8634 gnd.n6039 gnd.n1391 19.3944
R8635 gnd.n6141 gnd.n1391 19.3944
R8636 gnd.n6142 gnd.n6141 19.3944
R8637 gnd.n6142 gnd.n1388 19.3944
R8638 gnd.n6150 gnd.n1388 19.3944
R8639 gnd.n6150 gnd.n1389 19.3944
R8640 gnd.n6146 gnd.n1389 19.3944
R8641 gnd.n6146 gnd.n1354 19.3944
R8642 gnd.n6210 gnd.n1354 19.3944
R8643 gnd.n6210 gnd.n1351 19.3944
R8644 gnd.n6215 gnd.n1351 19.3944
R8645 gnd.n6215 gnd.n1352 19.3944
R8646 gnd.n1352 gnd.n1298 19.3944
R8647 gnd.n6289 gnd.n1298 19.3944
R8648 gnd.n6289 gnd.n1296 19.3944
R8649 gnd.n6294 gnd.n1296 19.3944
R8650 gnd.n6294 gnd.n1294 19.3944
R8651 gnd.n6298 gnd.n1294 19.3944
R8652 gnd.n6299 gnd.n6298 19.3944
R8653 gnd.n6299 gnd.n1292 19.3944
R8654 gnd.n6303 gnd.n1292 19.3944
R8655 gnd.n6304 gnd.n6303 19.3944
R8656 gnd.n6307 gnd.n6304 19.3944
R8657 gnd.n6307 gnd.n1288 19.3944
R8658 gnd.n6342 gnd.n1288 19.3944
R8659 gnd.n6342 gnd.n1289 19.3944
R8660 gnd.n6338 gnd.n1289 19.3944
R8661 gnd.n6338 gnd.n6337 19.3944
R8662 gnd.n6337 gnd.n6336 19.3944
R8663 gnd.n6336 gnd.n6313 19.3944
R8664 gnd.n6332 gnd.n6313 19.3944
R8665 gnd.n6332 gnd.n6331 19.3944
R8666 gnd.n6331 gnd.n6330 19.3944
R8667 gnd.n6330 gnd.n6325 19.3944
R8668 gnd.n6326 gnd.n6325 19.3944
R8669 gnd.n6326 gnd.n1154 19.3944
R8670 gnd.n6540 gnd.n1154 19.3944
R8671 gnd.n6540 gnd.n1151 19.3944
R8672 gnd.n6558 gnd.n1151 19.3944
R8673 gnd.n6558 gnd.n1152 19.3944
R8674 gnd.n6554 gnd.n1152 19.3944
R8675 gnd.n6554 gnd.n6553 19.3944
R8676 gnd.n6553 gnd.n6552 19.3944
R8677 gnd.n6552 gnd.n6548 19.3944
R8678 gnd.n6548 gnd.n1106 19.3944
R8679 gnd.n6642 gnd.n1106 19.3944
R8680 gnd.n6643 gnd.n6642 19.3944
R8681 gnd.n6643 gnd.n1104 19.3944
R8682 gnd.n6647 gnd.n1104 19.3944
R8683 gnd.n6649 gnd.n6647 19.3944
R8684 gnd.n6650 gnd.n6649 19.3944
R8685 gnd.n6650 gnd.n1099 19.3944
R8686 gnd.n6670 gnd.n1099 19.3944
R8687 gnd.n6670 gnd.n1100 19.3944
R8688 gnd.n6666 gnd.n1100 19.3944
R8689 gnd.n6666 gnd.n6665 19.3944
R8690 gnd.n6665 gnd.n6664 19.3944
R8691 gnd.n6664 gnd.n6660 19.3944
R8692 gnd.n6660 gnd.n1012 19.3944
R8693 gnd.n6825 gnd.n1012 19.3944
R8694 gnd.n6826 gnd.n6825 19.3944
R8695 gnd.n6826 gnd.n1009 19.3944
R8696 gnd.n6833 gnd.n1009 19.3944
R8697 gnd.n6833 gnd.n1010 19.3944
R8698 gnd.n6829 gnd.n1010 19.3944
R8699 gnd.n6829 gnd.n722 19.3944
R8700 gnd.n7015 gnd.n722 19.3944
R8701 gnd.n7015 gnd.n719 19.3944
R8702 gnd.n7020 gnd.n719 19.3944
R8703 gnd.n7020 gnd.n720 19.3944
R8704 gnd.n720 gnd.n697 19.3944
R8705 gnd.n7045 gnd.n697 19.3944
R8706 gnd.n7045 gnd.n694 19.3944
R8707 gnd.n7055 gnd.n694 19.3944
R8708 gnd.n7055 gnd.n695 19.3944
R8709 gnd.n7051 gnd.n695 19.3944
R8710 gnd.n7051 gnd.n7050 19.3944
R8711 gnd.n7050 gnd.n582 19.3944
R8712 gnd.n7187 gnd.n582 19.3944
R8713 gnd.n5674 gnd.n1685 19.3944
R8714 gnd.n5740 gnd.n1685 19.3944
R8715 gnd.n5740 gnd.n5739 19.3944
R8716 gnd.n5733 gnd.n5732 19.3944
R8717 gnd.n5732 gnd.n1707 19.3944
R8718 gnd.n5728 gnd.n1707 19.3944
R8719 gnd.n5728 gnd.n5727 19.3944
R8720 gnd.n5727 gnd.n5726 19.3944
R8721 gnd.n5726 gnd.n5723 19.3944
R8722 gnd.n5723 gnd.n5722 19.3944
R8723 gnd.n5722 gnd.n1714 19.3944
R8724 gnd.n5604 gnd.n1714 19.3944
R8725 gnd.n5714 gnd.n5604 19.3944
R8726 gnd.n5714 gnd.n5713 19.3944
R8727 gnd.n5713 gnd.n5607 19.3944
R8728 gnd.n5706 gnd.n5607 19.3944
R8729 gnd.n5706 gnd.n5705 19.3944
R8730 gnd.n5705 gnd.n5620 19.3944
R8731 gnd.n5698 gnd.n5620 19.3944
R8732 gnd.n5698 gnd.n5697 19.3944
R8733 gnd.n5697 gnd.n5630 19.3944
R8734 gnd.n5690 gnd.n5630 19.3944
R8735 gnd.n5690 gnd.n5689 19.3944
R8736 gnd.n5689 gnd.n5643 19.3944
R8737 gnd.n5682 gnd.n5643 19.3944
R8738 gnd.n5682 gnd.n5681 19.3944
R8739 gnd.n5681 gnd.n5653 19.3944
R8740 gnd.n7163 gnd.n606 19.3944
R8741 gnd.n7163 gnd.n7162 19.3944
R8742 gnd.n7162 gnd.n609 19.3944
R8743 gnd.n7155 gnd.n609 19.3944
R8744 gnd.n7155 gnd.n7154 19.3944
R8745 gnd.n7154 gnd.n619 19.3944
R8746 gnd.n7147 gnd.n619 19.3944
R8747 gnd.n7147 gnd.n7146 19.3944
R8748 gnd.n7146 gnd.n627 19.3944
R8749 gnd.n7139 gnd.n627 19.3944
R8750 gnd.n7139 gnd.n7138 19.3944
R8751 gnd.n7138 gnd.n637 19.3944
R8752 gnd.n7131 gnd.n637 19.3944
R8753 gnd.n7131 gnd.n7130 19.3944
R8754 gnd.n7130 gnd.n568 19.3944
R8755 gnd.n7200 gnd.n568 19.3944
R8756 gnd.n3919 gnd.n3918 19.3944
R8757 gnd.n3918 gnd.n3917 19.3944
R8758 gnd.n3917 gnd.n3916 19.3944
R8759 gnd.n3916 gnd.n3914 19.3944
R8760 gnd.n3914 gnd.n3911 19.3944
R8761 gnd.n3911 gnd.n3910 19.3944
R8762 gnd.n3910 gnd.n3907 19.3944
R8763 gnd.n3907 gnd.n3906 19.3944
R8764 gnd.n3906 gnd.n3903 19.3944
R8765 gnd.n3903 gnd.n3902 19.3944
R8766 gnd.n3902 gnd.n3899 19.3944
R8767 gnd.n3899 gnd.n3898 19.3944
R8768 gnd.n3898 gnd.n3895 19.3944
R8769 gnd.n3895 gnd.n3894 19.3944
R8770 gnd.n3894 gnd.n3891 19.3944
R8771 gnd.n3891 gnd.n3890 19.3944
R8772 gnd.n3890 gnd.n3887 19.3944
R8773 gnd.n3887 gnd.n3886 19.3944
R8774 gnd.n3886 gnd.n3883 19.3944
R8775 gnd.n3883 gnd.n3882 19.3944
R8776 gnd.n3882 gnd.n3879 19.3944
R8777 gnd.n3879 gnd.n3878 19.3944
R8778 gnd.n3875 gnd.n3874 19.3944
R8779 gnd.n3874 gnd.n3830 19.3944
R8780 gnd.n3925 gnd.n3830 19.3944
R8781 gnd.n4691 gnd.n4690 19.3944
R8782 gnd.n4690 gnd.n4687 19.3944
R8783 gnd.n4687 gnd.n4686 19.3944
R8784 gnd.n4736 gnd.n4735 19.3944
R8785 gnd.n4735 gnd.n4734 19.3944
R8786 gnd.n4734 gnd.n4731 19.3944
R8787 gnd.n4731 gnd.n4730 19.3944
R8788 gnd.n4730 gnd.n4727 19.3944
R8789 gnd.n4727 gnd.n4726 19.3944
R8790 gnd.n4726 gnd.n4723 19.3944
R8791 gnd.n4723 gnd.n4722 19.3944
R8792 gnd.n4722 gnd.n4719 19.3944
R8793 gnd.n4719 gnd.n4718 19.3944
R8794 gnd.n4718 gnd.n4715 19.3944
R8795 gnd.n4715 gnd.n4714 19.3944
R8796 gnd.n4714 gnd.n4711 19.3944
R8797 gnd.n4711 gnd.n4710 19.3944
R8798 gnd.n4710 gnd.n4707 19.3944
R8799 gnd.n4707 gnd.n4706 19.3944
R8800 gnd.n4706 gnd.n4703 19.3944
R8801 gnd.n4703 gnd.n4702 19.3944
R8802 gnd.n4702 gnd.n4699 19.3944
R8803 gnd.n4699 gnd.n4698 19.3944
R8804 gnd.n4698 gnd.n4695 19.3944
R8805 gnd.n4695 gnd.n4694 19.3944
R8806 gnd.n4018 gnd.n3727 19.3944
R8807 gnd.n4028 gnd.n3727 19.3944
R8808 gnd.n4029 gnd.n4028 19.3944
R8809 gnd.n4029 gnd.n3708 19.3944
R8810 gnd.n4049 gnd.n3708 19.3944
R8811 gnd.n4049 gnd.n3700 19.3944
R8812 gnd.n4059 gnd.n3700 19.3944
R8813 gnd.n4060 gnd.n4059 19.3944
R8814 gnd.n4061 gnd.n4060 19.3944
R8815 gnd.n4061 gnd.n3683 19.3944
R8816 gnd.n4078 gnd.n3683 19.3944
R8817 gnd.n4081 gnd.n4078 19.3944
R8818 gnd.n4081 gnd.n4080 19.3944
R8819 gnd.n4080 gnd.n3656 19.3944
R8820 gnd.n4120 gnd.n3656 19.3944
R8821 gnd.n4120 gnd.n3653 19.3944
R8822 gnd.n4126 gnd.n3653 19.3944
R8823 gnd.n4127 gnd.n4126 19.3944
R8824 gnd.n4127 gnd.n3651 19.3944
R8825 gnd.n4133 gnd.n3651 19.3944
R8826 gnd.n4136 gnd.n4133 19.3944
R8827 gnd.n4138 gnd.n4136 19.3944
R8828 gnd.n4144 gnd.n4138 19.3944
R8829 gnd.n4144 gnd.n4143 19.3944
R8830 gnd.n4143 gnd.n3510 19.3944
R8831 gnd.n4210 gnd.n3510 19.3944
R8832 gnd.n4211 gnd.n4210 19.3944
R8833 gnd.n4211 gnd.n3503 19.3944
R8834 gnd.n4222 gnd.n3503 19.3944
R8835 gnd.n4223 gnd.n4222 19.3944
R8836 gnd.n4223 gnd.n3486 19.3944
R8837 gnd.n3486 gnd.n3484 19.3944
R8838 gnd.n4247 gnd.n3484 19.3944
R8839 gnd.n4248 gnd.n4247 19.3944
R8840 gnd.n4248 gnd.n3455 19.3944
R8841 gnd.n4295 gnd.n3455 19.3944
R8842 gnd.n4296 gnd.n4295 19.3944
R8843 gnd.n4296 gnd.n3448 19.3944
R8844 gnd.n4307 gnd.n3448 19.3944
R8845 gnd.n4308 gnd.n4307 19.3944
R8846 gnd.n4308 gnd.n3431 19.3944
R8847 gnd.n3431 gnd.n3429 19.3944
R8848 gnd.n4332 gnd.n3429 19.3944
R8849 gnd.n4333 gnd.n4332 19.3944
R8850 gnd.n4333 gnd.n3401 19.3944
R8851 gnd.n4384 gnd.n3401 19.3944
R8852 gnd.n4385 gnd.n4384 19.3944
R8853 gnd.n4385 gnd.n3394 19.3944
R8854 gnd.n4652 gnd.n3394 19.3944
R8855 gnd.n4653 gnd.n4652 19.3944
R8856 gnd.n4653 gnd.n2070 19.3944
R8857 gnd.n4678 gnd.n2070 19.3944
R8858 gnd.n4678 gnd.n2071 19.3944
R8859 gnd.n4009 gnd.n4008 19.3944
R8860 gnd.n4008 gnd.n3741 19.3944
R8861 gnd.n3764 gnd.n3741 19.3944
R8862 gnd.n3767 gnd.n3764 19.3944
R8863 gnd.n3767 gnd.n3760 19.3944
R8864 gnd.n3771 gnd.n3760 19.3944
R8865 gnd.n3774 gnd.n3771 19.3944
R8866 gnd.n3777 gnd.n3774 19.3944
R8867 gnd.n3777 gnd.n3758 19.3944
R8868 gnd.n3781 gnd.n3758 19.3944
R8869 gnd.n3784 gnd.n3781 19.3944
R8870 gnd.n3787 gnd.n3784 19.3944
R8871 gnd.n3787 gnd.n3756 19.3944
R8872 gnd.n3791 gnd.n3756 19.3944
R8873 gnd.n4014 gnd.n4013 19.3944
R8874 gnd.n4013 gnd.n3717 19.3944
R8875 gnd.n4039 gnd.n3717 19.3944
R8876 gnd.n4039 gnd.n3715 19.3944
R8877 gnd.n4045 gnd.n3715 19.3944
R8878 gnd.n4045 gnd.n4044 19.3944
R8879 gnd.n4044 gnd.n3689 19.3944
R8880 gnd.n4069 gnd.n3689 19.3944
R8881 gnd.n4069 gnd.n3687 19.3944
R8882 gnd.n4073 gnd.n3687 19.3944
R8883 gnd.n4073 gnd.n3667 19.3944
R8884 gnd.n4100 gnd.n3667 19.3944
R8885 gnd.n4100 gnd.n3665 19.3944
R8886 gnd.n4110 gnd.n3665 19.3944
R8887 gnd.n4110 gnd.n4109 19.3944
R8888 gnd.n4109 gnd.n4108 19.3944
R8889 gnd.n4108 gnd.n3614 19.3944
R8890 gnd.n4158 gnd.n3614 19.3944
R8891 gnd.n4158 gnd.n4157 19.3944
R8892 gnd.n4157 gnd.n4156 19.3944
R8893 gnd.n4156 gnd.n3618 19.3944
R8894 gnd.n3638 gnd.n3618 19.3944
R8895 gnd.n3638 gnd.n3520 19.3944
R8896 gnd.n4195 gnd.n3520 19.3944
R8897 gnd.n4195 gnd.n3518 19.3944
R8898 gnd.n4201 gnd.n3518 19.3944
R8899 gnd.n4201 gnd.n4200 19.3944
R8900 gnd.n4200 gnd.n3493 19.3944
R8901 gnd.n4235 gnd.n3493 19.3944
R8902 gnd.n4235 gnd.n3491 19.3944
R8903 gnd.n4241 gnd.n3491 19.3944
R8904 gnd.n4241 gnd.n4240 19.3944
R8905 gnd.n4240 gnd.n3466 19.3944
R8906 gnd.n4280 gnd.n3466 19.3944
R8907 gnd.n4280 gnd.n3464 19.3944
R8908 gnd.n4286 gnd.n3464 19.3944
R8909 gnd.n4286 gnd.n4285 19.3944
R8910 gnd.n4285 gnd.n3438 19.3944
R8911 gnd.n4320 gnd.n3438 19.3944
R8912 gnd.n4320 gnd.n3436 19.3944
R8913 gnd.n4326 gnd.n3436 19.3944
R8914 gnd.n4326 gnd.n4325 19.3944
R8915 gnd.n4325 gnd.n3411 19.3944
R8916 gnd.n4369 gnd.n3411 19.3944
R8917 gnd.n4369 gnd.n3409 19.3944
R8918 gnd.n4375 gnd.n3409 19.3944
R8919 gnd.n4375 gnd.n4374 19.3944
R8920 gnd.n4374 gnd.n3384 19.3944
R8921 gnd.n4663 gnd.n3384 19.3944
R8922 gnd.n4663 gnd.n3382 19.3944
R8923 gnd.n4671 gnd.n3382 19.3944
R8924 gnd.n4671 gnd.n4670 19.3944
R8925 gnd.n4670 gnd.n4669 19.3944
R8926 gnd.n4772 gnd.n4771 19.3944
R8927 gnd.n4771 gnd.n2018 19.3944
R8928 gnd.n4767 gnd.n2018 19.3944
R8929 gnd.n4767 gnd.n4764 19.3944
R8930 gnd.n4764 gnd.n4761 19.3944
R8931 gnd.n4761 gnd.n4760 19.3944
R8932 gnd.n4760 gnd.n4757 19.3944
R8933 gnd.n4757 gnd.n4756 19.3944
R8934 gnd.n4756 gnd.n4753 19.3944
R8935 gnd.n4753 gnd.n4752 19.3944
R8936 gnd.n4752 gnd.n4749 19.3944
R8937 gnd.n4749 gnd.n4748 19.3944
R8938 gnd.n4748 gnd.n4745 19.3944
R8939 gnd.n4745 gnd.n4744 19.3944
R8940 gnd.n3929 gnd.n3828 19.3944
R8941 gnd.n3929 gnd.n3819 19.3944
R8942 gnd.n3942 gnd.n3819 19.3944
R8943 gnd.n3942 gnd.n3817 19.3944
R8944 gnd.n3946 gnd.n3817 19.3944
R8945 gnd.n3946 gnd.n3807 19.3944
R8946 gnd.n3958 gnd.n3807 19.3944
R8947 gnd.n3958 gnd.n3805 19.3944
R8948 gnd.n3992 gnd.n3805 19.3944
R8949 gnd.n3992 gnd.n3991 19.3944
R8950 gnd.n3991 gnd.n3990 19.3944
R8951 gnd.n3990 gnd.n3989 19.3944
R8952 gnd.n3989 gnd.n3986 19.3944
R8953 gnd.n3986 gnd.n3985 19.3944
R8954 gnd.n3985 gnd.n3984 19.3944
R8955 gnd.n3984 gnd.n3982 19.3944
R8956 gnd.n3982 gnd.n3981 19.3944
R8957 gnd.n3981 gnd.n3978 19.3944
R8958 gnd.n3978 gnd.n3977 19.3944
R8959 gnd.n3977 gnd.n3976 19.3944
R8960 gnd.n3976 gnd.n3974 19.3944
R8961 gnd.n3974 gnd.n3673 19.3944
R8962 gnd.n4089 gnd.n3673 19.3944
R8963 gnd.n4089 gnd.n3671 19.3944
R8964 gnd.n4095 gnd.n3671 19.3944
R8965 gnd.n4095 gnd.n4094 19.3944
R8966 gnd.n4094 gnd.n3595 19.3944
R8967 gnd.n4169 gnd.n3595 19.3944
R8968 gnd.n4169 gnd.n3596 19.3944
R8969 gnd.n3643 gnd.n3642 19.3944
R8970 gnd.n3646 gnd.n3645 19.3944
R8971 gnd.n3633 gnd.n3632 19.3944
R8972 gnd.n4188 gnd.n3525 19.3944
R8973 gnd.n4188 gnd.n4187 19.3944
R8974 gnd.n4187 gnd.n4186 19.3944
R8975 gnd.n4186 gnd.n4184 19.3944
R8976 gnd.n4184 gnd.n4183 19.3944
R8977 gnd.n4183 gnd.n4181 19.3944
R8978 gnd.n4181 gnd.n4180 19.3944
R8979 gnd.n4180 gnd.n3474 19.3944
R8980 gnd.n4256 gnd.n3474 19.3944
R8981 gnd.n4256 gnd.n3472 19.3944
R8982 gnd.n4275 gnd.n3472 19.3944
R8983 gnd.n4275 gnd.n4274 19.3944
R8984 gnd.n4274 gnd.n4273 19.3944
R8985 gnd.n4273 gnd.n4271 19.3944
R8986 gnd.n4271 gnd.n4270 19.3944
R8987 gnd.n4270 gnd.n4268 19.3944
R8988 gnd.n4268 gnd.n4267 19.3944
R8989 gnd.n4267 gnd.n3418 19.3944
R8990 gnd.n4341 gnd.n3418 19.3944
R8991 gnd.n4341 gnd.n3416 19.3944
R8992 gnd.n4364 gnd.n3416 19.3944
R8993 gnd.n4364 gnd.n4363 19.3944
R8994 gnd.n4363 gnd.n4362 19.3944
R8995 gnd.n4362 gnd.n4359 19.3944
R8996 gnd.n4359 gnd.n4358 19.3944
R8997 gnd.n4358 gnd.n4356 19.3944
R8998 gnd.n4356 gnd.n4355 19.3944
R8999 gnd.n4355 gnd.n4353 19.3944
R9000 gnd.n4353 gnd.n2065 19.3944
R9001 gnd.n3934 gnd.n3824 19.3944
R9002 gnd.n3934 gnd.n3822 19.3944
R9003 gnd.n3938 gnd.n3822 19.3944
R9004 gnd.n3938 gnd.n3813 19.3944
R9005 gnd.n3950 gnd.n3813 19.3944
R9006 gnd.n3950 gnd.n3811 19.3944
R9007 gnd.n3954 gnd.n3811 19.3944
R9008 gnd.n3954 gnd.n3800 19.3944
R9009 gnd.n3996 gnd.n3800 19.3944
R9010 gnd.n3996 gnd.n3754 19.3944
R9011 gnd.n4002 gnd.n3754 19.3944
R9012 gnd.n4002 gnd.n4001 19.3944
R9013 gnd.n4001 gnd.n3732 19.3944
R9014 gnd.n4023 gnd.n3732 19.3944
R9015 gnd.n4023 gnd.n3725 19.3944
R9016 gnd.n4034 gnd.n3725 19.3944
R9017 gnd.n4034 gnd.n4033 19.3944
R9018 gnd.n4033 gnd.n3706 19.3944
R9019 gnd.n4054 gnd.n3706 19.3944
R9020 gnd.n4054 gnd.n3696 19.3944
R9021 gnd.n4064 gnd.n3696 19.3944
R9022 gnd.n4064 gnd.n3679 19.3944
R9023 gnd.n4085 gnd.n3679 19.3944
R9024 gnd.n4085 gnd.n4084 19.3944
R9025 gnd.n4084 gnd.n3658 19.3944
R9026 gnd.n4115 gnd.n3658 19.3944
R9027 gnd.n4115 gnd.n3603 19.3944
R9028 gnd.n4165 gnd.n3603 19.3944
R9029 gnd.n4165 gnd.n4164 19.3944
R9030 gnd.n4164 gnd.n4163 19.3944
R9031 gnd.n4163 gnd.n3607 19.3944
R9032 gnd.n3625 gnd.n3607 19.3944
R9033 gnd.n4151 gnd.n3625 19.3944
R9034 gnd.n4151 gnd.n4150 19.3944
R9035 gnd.n4150 gnd.n4149 19.3944
R9036 gnd.n4149 gnd.n3629 19.3944
R9037 gnd.n3629 gnd.n3512 19.3944
R9038 gnd.n4206 gnd.n3512 19.3944
R9039 gnd.n4206 gnd.n3505 19.3944
R9040 gnd.n4217 gnd.n3505 19.3944
R9041 gnd.n4217 gnd.n3501 19.3944
R9042 gnd.n4230 gnd.n3501 19.3944
R9043 gnd.n4230 gnd.n4229 19.3944
R9044 gnd.n4229 gnd.n3480 19.3944
R9045 gnd.n4252 gnd.n3480 19.3944
R9046 gnd.n4252 gnd.n4251 19.3944
R9047 gnd.n4251 gnd.n3457 19.3944
R9048 gnd.n4291 gnd.n3457 19.3944
R9049 gnd.n4291 gnd.n3450 19.3944
R9050 gnd.n4302 gnd.n3450 19.3944
R9051 gnd.n4302 gnd.n3446 19.3944
R9052 gnd.n4315 gnd.n3446 19.3944
R9053 gnd.n4315 gnd.n4314 19.3944
R9054 gnd.n4314 gnd.n3425 19.3944
R9055 gnd.n4337 gnd.n3425 19.3944
R9056 gnd.n4337 gnd.n4336 19.3944
R9057 gnd.n4336 gnd.n3403 19.3944
R9058 gnd.n4380 gnd.n3403 19.3944
R9059 gnd.n4380 gnd.n3396 19.3944
R9060 gnd.n4391 gnd.n3396 19.3944
R9061 gnd.n4391 gnd.n3392 19.3944
R9062 gnd.n4658 gnd.n3392 19.3944
R9063 gnd.n4658 gnd.n4657 19.3944
R9064 gnd.n4657 gnd.n2068 19.3944
R9065 gnd.n4681 gnd.n2068 19.3944
R9066 gnd.n5718 gnd.n5717 19.3944
R9067 gnd.n5717 gnd.n5600 19.3944
R9068 gnd.n5710 gnd.n5600 19.3944
R9069 gnd.n5710 gnd.n5709 19.3944
R9070 gnd.n5709 gnd.n5614 19.3944
R9071 gnd.n5702 gnd.n5614 19.3944
R9072 gnd.n5702 gnd.n5701 19.3944
R9073 gnd.n5701 gnd.n5626 19.3944
R9074 gnd.n5694 gnd.n5626 19.3944
R9075 gnd.n5694 gnd.n5693 19.3944
R9076 gnd.n5693 gnd.n5637 19.3944
R9077 gnd.n5686 gnd.n5637 19.3944
R9078 gnd.n5686 gnd.n5685 19.3944
R9079 gnd.n5685 gnd.n5649 19.3944
R9080 gnd.n5678 gnd.n5649 19.3944
R9081 gnd.n5678 gnd.n5677 19.3944
R9082 gnd.n2080 gnd.n2079 19.3944
R9083 gnd.n2079 gnd.n1812 19.3944
R9084 gnd.n1812 gnd.n1810 19.3944
R9085 gnd.n5317 gnd.n1810 19.3944
R9086 gnd.n5317 gnd.n1808 19.3944
R9087 gnd.n5323 gnd.n1808 19.3944
R9088 gnd.n5323 gnd.n5322 19.3944
R9089 gnd.n5322 gnd.n1774 19.3944
R9090 gnd.n5362 gnd.n1774 19.3944
R9091 gnd.n5362 gnd.n1772 19.3944
R9092 gnd.n5371 gnd.n1772 19.3944
R9093 gnd.n5371 gnd.n5370 19.3944
R9094 gnd.n5370 gnd.n5369 19.3944
R9095 gnd.n5369 gnd.n1724 19.3944
R9096 gnd.n5426 gnd.n1724 19.3944
R9097 gnd.n5426 gnd.n1722 19.3944
R9098 gnd.n5430 gnd.n1722 19.3944
R9099 gnd.n5430 gnd.n1720 19.3944
R9100 gnd.n5434 gnd.n1720 19.3944
R9101 gnd.n5434 gnd.n1718 19.3944
R9102 gnd.n5593 gnd.n1718 19.3944
R9103 gnd.n5593 gnd.n5592 19.3944
R9104 gnd.n5592 gnd.n5591 19.3944
R9105 gnd.n5591 gnd.n5440 19.3944
R9106 gnd.n5585 gnd.n5440 19.3944
R9107 gnd.n5585 gnd.n5584 19.3944
R9108 gnd.n5584 gnd.n5583 19.3944
R9109 gnd.n5583 gnd.n5446 19.3944
R9110 gnd.n5497 gnd.n5446 19.3944
R9111 gnd.n5515 gnd.n5497 19.3944
R9112 gnd.n5515 gnd.n5494 19.3944
R9113 gnd.n5519 gnd.n5494 19.3944
R9114 gnd.n5519 gnd.n5482 19.3944
R9115 gnd.n5534 gnd.n5482 19.3944
R9116 gnd.n5534 gnd.n5480 19.3944
R9117 gnd.n5540 gnd.n5480 19.3944
R9118 gnd.n5540 gnd.n5539 19.3944
R9119 gnd.n5539 gnd.n1463 19.3944
R9120 gnd.n6014 gnd.n1463 19.3944
R9121 gnd.n6014 gnd.n1461 19.3944
R9122 gnd.n6018 gnd.n1461 19.3944
R9123 gnd.n6018 gnd.n1433 19.3944
R9124 gnd.n6074 gnd.n1433 19.3944
R9125 gnd.n6074 gnd.n1431 19.3944
R9126 gnd.n6078 gnd.n1431 19.3944
R9127 gnd.n6078 gnd.n1406 19.3944
R9128 gnd.n6116 gnd.n1406 19.3944
R9129 gnd.n6116 gnd.n1404 19.3944
R9130 gnd.n6128 gnd.n1404 19.3944
R9131 gnd.n6128 gnd.n6127 19.3944
R9132 gnd.n6127 gnd.n6126 19.3944
R9133 gnd.n6126 gnd.n6123 19.3944
R9134 gnd.n6123 gnd.n1362 19.3944
R9135 gnd.n6187 gnd.n1362 19.3944
R9136 gnd.n6187 gnd.n1360 19.3944
R9137 gnd.n6191 gnd.n1360 19.3944
R9138 gnd.n6191 gnd.n1331 19.3944
R9139 gnd.n6238 gnd.n1331 19.3944
R9140 gnd.n6238 gnd.n1329 19.3944
R9141 gnd.n6242 gnd.n1329 19.3944
R9142 gnd.n6242 gnd.n1327 19.3944
R9143 gnd.n6249 gnd.n1327 19.3944
R9144 gnd.n6249 gnd.n1325 19.3944
R9145 gnd.n6253 gnd.n1325 19.3944
R9146 gnd.n6253 gnd.n1268 19.3944
R9147 gnd.n6384 gnd.n1268 19.3944
R9148 gnd.n6384 gnd.n1266 19.3944
R9149 gnd.n6388 gnd.n1266 19.3944
R9150 gnd.n6388 gnd.n1244 19.3944
R9151 gnd.n6411 gnd.n1244 19.3944
R9152 gnd.n6411 gnd.n1242 19.3944
R9153 gnd.n6417 gnd.n1242 19.3944
R9154 gnd.n6417 gnd.n6416 19.3944
R9155 gnd.n6416 gnd.n1212 19.3944
R9156 gnd.n6448 gnd.n1212 19.3944
R9157 gnd.n6448 gnd.n1210 19.3944
R9158 gnd.n6452 gnd.n1210 19.3944
R9159 gnd.n6452 gnd.n1189 19.3944
R9160 gnd.n6482 gnd.n1189 19.3944
R9161 gnd.n6482 gnd.n1187 19.3944
R9162 gnd.n6502 gnd.n1187 19.3944
R9163 gnd.n6502 gnd.n6501 19.3944
R9164 gnd.n6501 gnd.n6500 19.3944
R9165 gnd.n6500 gnd.n6488 19.3944
R9166 gnd.n6494 gnd.n6488 19.3944
R9167 gnd.n6494 gnd.n6493 19.3944
R9168 gnd.n6493 gnd.n1130 19.3944
R9169 gnd.n6603 gnd.n1130 19.3944
R9170 gnd.n6603 gnd.n1128 19.3944
R9171 gnd.n6614 gnd.n1128 19.3944
R9172 gnd.n6614 gnd.n6613 19.3944
R9173 gnd.n6613 gnd.n6612 19.3944
R9174 gnd.n6612 gnd.n1091 19.3944
R9175 gnd.n6695 gnd.n1091 19.3944
R9176 gnd.n6695 gnd.n1089 19.3944
R9177 gnd.n6699 gnd.n1089 19.3944
R9178 gnd.n6699 gnd.n1068 19.3944
R9179 gnd.n6723 gnd.n1068 19.3944
R9180 gnd.n6723 gnd.n1066 19.3944
R9181 gnd.n6736 gnd.n1066 19.3944
R9182 gnd.n6736 gnd.n6735 19.3944
R9183 gnd.n6735 gnd.n6734 19.3944
R9184 gnd.n6734 gnd.n6730 19.3944
R9185 gnd.n6730 gnd.n1025 19.3944
R9186 gnd.n6806 gnd.n1025 19.3944
R9187 gnd.n6806 gnd.n1023 19.3944
R9188 gnd.n6810 gnd.n1023 19.3944
R9189 gnd.n6810 gnd.n997 19.3944
R9190 gnd.n6847 gnd.n997 19.3944
R9191 gnd.n6847 gnd.n995 19.3944
R9192 gnd.n6863 gnd.n995 19.3944
R9193 gnd.n6863 gnd.n6862 19.3944
R9194 gnd.n6862 gnd.n6861 19.3944
R9195 gnd.n6861 gnd.n6853 19.3944
R9196 gnd.n6856 gnd.n6853 19.3944
R9197 gnd.n6856 gnd.n715 19.3944
R9198 gnd.n7025 gnd.n715 19.3944
R9199 gnd.n7025 gnd.n713 19.3944
R9200 gnd.n7031 gnd.n713 19.3944
R9201 gnd.n7031 gnd.n7030 19.3944
R9202 gnd.n7030 gnd.n690 19.3944
R9203 gnd.n7060 gnd.n690 19.3944
R9204 gnd.n7060 gnd.n688 19.3944
R9205 gnd.n7067 gnd.n688 19.3944
R9206 gnd.n7067 gnd.n7066 19.3944
R9207 gnd.n7066 gnd.n676 19.3944
R9208 gnd.n676 gnd.n674 19.3944
R9209 gnd.n7084 gnd.n674 19.3944
R9210 gnd.n7084 gnd.n672 19.3944
R9211 gnd.n7121 gnd.n672 19.3944
R9212 gnd.n7121 gnd.n7120 19.3944
R9213 gnd.n7120 gnd.n7119 19.3944
R9214 gnd.n7119 gnd.n7090 19.3944
R9215 gnd.n7115 gnd.n7090 19.3944
R9216 gnd.n7115 gnd.n7114 19.3944
R9217 gnd.n7114 gnd.n7113 19.3944
R9218 gnd.n7113 gnd.n7104 19.3944
R9219 gnd.n7109 gnd.n7104 19.3944
R9220 gnd.n7109 gnd.n7108 19.3944
R9221 gnd.n7108 gnd.n481 19.3944
R9222 gnd.n7264 gnd.n481 19.3944
R9223 gnd.n7264 gnd.n479 19.3944
R9224 gnd.n7270 gnd.n479 19.3944
R9225 gnd.n7270 gnd.n7269 19.3944
R9226 gnd.n7269 gnd.n447 19.3944
R9227 gnd.n7310 gnd.n447 19.3944
R9228 gnd.n7310 gnd.n445 19.3944
R9229 gnd.n7316 gnd.n445 19.3944
R9230 gnd.n7316 gnd.n7315 19.3944
R9231 gnd.n7315 gnd.n412 19.3944
R9232 gnd.n7356 gnd.n412 19.3944
R9233 gnd.n7356 gnd.n410 19.3944
R9234 gnd.n7362 gnd.n410 19.3944
R9235 gnd.n7362 gnd.n7361 19.3944
R9236 gnd.n2849 gnd.n2517 19.3944
R9237 gnd.n2849 gnd.n2518 19.3944
R9238 gnd.n2845 gnd.n2518 19.3944
R9239 gnd.n2845 gnd.n2521 19.3944
R9240 gnd.n2839 gnd.n2521 19.3944
R9241 gnd.n2839 gnd.n2838 19.3944
R9242 gnd.n2838 gnd.n2837 19.3944
R9243 gnd.n2837 gnd.n2528 19.3944
R9244 gnd.n2831 gnd.n2528 19.3944
R9245 gnd.n2831 gnd.n2830 19.3944
R9246 gnd.n2830 gnd.n2829 19.3944
R9247 gnd.n2829 gnd.n2536 19.3944
R9248 gnd.n2823 gnd.n2536 19.3944
R9249 gnd.n2823 gnd.n2822 19.3944
R9250 gnd.n2822 gnd.n2821 19.3944
R9251 gnd.n2821 gnd.n2544 19.3944
R9252 gnd.n2815 gnd.n2544 19.3944
R9253 gnd.n2815 gnd.n2814 19.3944
R9254 gnd.n2814 gnd.n2813 19.3944
R9255 gnd.n2813 gnd.n2552 19.3944
R9256 gnd.n2807 gnd.n2552 19.3944
R9257 gnd.n2807 gnd.n2806 19.3944
R9258 gnd.n2806 gnd.n2805 19.3944
R9259 gnd.n2805 gnd.n2560 19.3944
R9260 gnd.n2799 gnd.n2560 19.3944
R9261 gnd.n2799 gnd.n2798 19.3944
R9262 gnd.n2798 gnd.n2797 19.3944
R9263 gnd.n2797 gnd.n2568 19.3944
R9264 gnd.n2791 gnd.n2568 19.3944
R9265 gnd.n2791 gnd.n2790 19.3944
R9266 gnd.n2790 gnd.n2789 19.3944
R9267 gnd.n2789 gnd.n2576 19.3944
R9268 gnd.n2783 gnd.n2576 19.3944
R9269 gnd.n2783 gnd.n2782 19.3944
R9270 gnd.n2782 gnd.n2781 19.3944
R9271 gnd.n2781 gnd.n2584 19.3944
R9272 gnd.n2775 gnd.n2584 19.3944
R9273 gnd.n2775 gnd.n2774 19.3944
R9274 gnd.n2774 gnd.n2773 19.3944
R9275 gnd.n2773 gnd.n2592 19.3944
R9276 gnd.n2767 gnd.n2592 19.3944
R9277 gnd.n2767 gnd.n2766 19.3944
R9278 gnd.n2766 gnd.n2765 19.3944
R9279 gnd.n2765 gnd.n2600 19.3944
R9280 gnd.n2759 gnd.n2600 19.3944
R9281 gnd.n2759 gnd.n2758 19.3944
R9282 gnd.n2758 gnd.n2757 19.3944
R9283 gnd.n2757 gnd.n2608 19.3944
R9284 gnd.n2751 gnd.n2608 19.3944
R9285 gnd.n2751 gnd.n2750 19.3944
R9286 gnd.n2750 gnd.n2749 19.3944
R9287 gnd.n2749 gnd.n2616 19.3944
R9288 gnd.n2743 gnd.n2616 19.3944
R9289 gnd.n2743 gnd.n2742 19.3944
R9290 gnd.n2742 gnd.n2741 19.3944
R9291 gnd.n2741 gnd.n2624 19.3944
R9292 gnd.n2735 gnd.n2624 19.3944
R9293 gnd.n2735 gnd.n2734 19.3944
R9294 gnd.n2734 gnd.n2733 19.3944
R9295 gnd.n2733 gnd.n2632 19.3944
R9296 gnd.n2727 gnd.n2632 19.3944
R9297 gnd.n2727 gnd.n2726 19.3944
R9298 gnd.n2726 gnd.n2725 19.3944
R9299 gnd.n2725 gnd.n2640 19.3944
R9300 gnd.n2719 gnd.n2640 19.3944
R9301 gnd.n2719 gnd.n2718 19.3944
R9302 gnd.n2718 gnd.n2717 19.3944
R9303 gnd.n2717 gnd.n2648 19.3944
R9304 gnd.n2711 gnd.n2648 19.3944
R9305 gnd.n2711 gnd.n2710 19.3944
R9306 gnd.n2710 gnd.n2709 19.3944
R9307 gnd.n2709 gnd.n2656 19.3944
R9308 gnd.n2703 gnd.n2656 19.3944
R9309 gnd.n2703 gnd.n2702 19.3944
R9310 gnd.n2702 gnd.n2701 19.3944
R9311 gnd.n2701 gnd.n2664 19.3944
R9312 gnd.n2695 gnd.n2664 19.3944
R9313 gnd.n2695 gnd.n2694 19.3944
R9314 gnd.n2694 gnd.n2693 19.3944
R9315 gnd.n2693 gnd.n2672 19.3944
R9316 gnd.n2687 gnd.n2672 19.3944
R9317 gnd.n2687 gnd.n2686 19.3944
R9318 gnd.n2686 gnd.n2685 19.3944
R9319 gnd.n2685 gnd.n2681 19.3944
R9320 gnd.n3163 gnd.n2209 19.3944
R9321 gnd.n3159 gnd.n2209 19.3944
R9322 gnd.n3159 gnd.n2211 19.3944
R9323 gnd.n3153 gnd.n2211 19.3944
R9324 gnd.n3153 gnd.n3152 19.3944
R9325 gnd.n3152 gnd.n3151 19.3944
R9326 gnd.n3151 gnd.n2218 19.3944
R9327 gnd.n3145 gnd.n2218 19.3944
R9328 gnd.n3145 gnd.n3144 19.3944
R9329 gnd.n3144 gnd.n3143 19.3944
R9330 gnd.n3143 gnd.n2226 19.3944
R9331 gnd.n3137 gnd.n2226 19.3944
R9332 gnd.n3137 gnd.n3136 19.3944
R9333 gnd.n3136 gnd.n3135 19.3944
R9334 gnd.n3135 gnd.n2234 19.3944
R9335 gnd.n3129 gnd.n2234 19.3944
R9336 gnd.n3129 gnd.n3128 19.3944
R9337 gnd.n3128 gnd.n3127 19.3944
R9338 gnd.n3127 gnd.n2242 19.3944
R9339 gnd.n3121 gnd.n2242 19.3944
R9340 gnd.n3121 gnd.n3120 19.3944
R9341 gnd.n3120 gnd.n3119 19.3944
R9342 gnd.n3119 gnd.n2250 19.3944
R9343 gnd.n3113 gnd.n2250 19.3944
R9344 gnd.n3113 gnd.n3112 19.3944
R9345 gnd.n3112 gnd.n3111 19.3944
R9346 gnd.n3111 gnd.n2258 19.3944
R9347 gnd.n3105 gnd.n2258 19.3944
R9348 gnd.n3105 gnd.n3104 19.3944
R9349 gnd.n3104 gnd.n3103 19.3944
R9350 gnd.n3103 gnd.n2266 19.3944
R9351 gnd.n3097 gnd.n2266 19.3944
R9352 gnd.n3097 gnd.n3096 19.3944
R9353 gnd.n3096 gnd.n3095 19.3944
R9354 gnd.n3095 gnd.n2274 19.3944
R9355 gnd.n3089 gnd.n2274 19.3944
R9356 gnd.n3089 gnd.n3088 19.3944
R9357 gnd.n3088 gnd.n3087 19.3944
R9358 gnd.n3087 gnd.n2282 19.3944
R9359 gnd.n3081 gnd.n2282 19.3944
R9360 gnd.n3081 gnd.n3080 19.3944
R9361 gnd.n3080 gnd.n3079 19.3944
R9362 gnd.n3079 gnd.n2290 19.3944
R9363 gnd.n3073 gnd.n2290 19.3944
R9364 gnd.n3073 gnd.n3072 19.3944
R9365 gnd.n3072 gnd.n3071 19.3944
R9366 gnd.n3071 gnd.n2298 19.3944
R9367 gnd.n3065 gnd.n2298 19.3944
R9368 gnd.n3065 gnd.n3064 19.3944
R9369 gnd.n3064 gnd.n3063 19.3944
R9370 gnd.n3063 gnd.n2306 19.3944
R9371 gnd.n3057 gnd.n2306 19.3944
R9372 gnd.n3057 gnd.n3056 19.3944
R9373 gnd.n3056 gnd.n3055 19.3944
R9374 gnd.n3055 gnd.n2314 19.3944
R9375 gnd.n3049 gnd.n2314 19.3944
R9376 gnd.n3049 gnd.n3048 19.3944
R9377 gnd.n3048 gnd.n3047 19.3944
R9378 gnd.n3047 gnd.n2322 19.3944
R9379 gnd.n3041 gnd.n2322 19.3944
R9380 gnd.n3041 gnd.n3040 19.3944
R9381 gnd.n3040 gnd.n3039 19.3944
R9382 gnd.n3039 gnd.n2330 19.3944
R9383 gnd.n3033 gnd.n2330 19.3944
R9384 gnd.n3033 gnd.n3032 19.3944
R9385 gnd.n3032 gnd.n3031 19.3944
R9386 gnd.n3031 gnd.n2338 19.3944
R9387 gnd.n3025 gnd.n2338 19.3944
R9388 gnd.n3025 gnd.n3024 19.3944
R9389 gnd.n3024 gnd.n3023 19.3944
R9390 gnd.n3023 gnd.n2346 19.3944
R9391 gnd.n3017 gnd.n2346 19.3944
R9392 gnd.n3017 gnd.n3016 19.3944
R9393 gnd.n3016 gnd.n3015 19.3944
R9394 gnd.n3015 gnd.n2354 19.3944
R9395 gnd.n3009 gnd.n2354 19.3944
R9396 gnd.n3009 gnd.n3008 19.3944
R9397 gnd.n3008 gnd.n3007 19.3944
R9398 gnd.n3007 gnd.n2362 19.3944
R9399 gnd.n3001 gnd.n2362 19.3944
R9400 gnd.n3001 gnd.n3000 19.3944
R9401 gnd.n3000 gnd.n2999 19.3944
R9402 gnd.n2999 gnd.n2370 19.3944
R9403 gnd.n2993 gnd.n2370 19.3944
R9404 gnd.n2993 gnd.n2992 19.3944
R9405 gnd.n2992 gnd.n2991 19.3944
R9406 gnd.n2991 gnd.n2378 19.3944
R9407 gnd.n2985 gnd.n2378 19.3944
R9408 gnd.n2985 gnd.n2984 19.3944
R9409 gnd.n2984 gnd.n2983 19.3944
R9410 gnd.n2983 gnd.n2386 19.3944
R9411 gnd.n2977 gnd.n2386 19.3944
R9412 gnd.n2977 gnd.n2976 19.3944
R9413 gnd.n2976 gnd.n2975 19.3944
R9414 gnd.n2975 gnd.n2394 19.3944
R9415 gnd.n2969 gnd.n2394 19.3944
R9416 gnd.n2969 gnd.n2968 19.3944
R9417 gnd.n2968 gnd.n2967 19.3944
R9418 gnd.n2967 gnd.n2402 19.3944
R9419 gnd.n2961 gnd.n2402 19.3944
R9420 gnd.n2961 gnd.n2960 19.3944
R9421 gnd.n2960 gnd.n2959 19.3944
R9422 gnd.n2959 gnd.n2410 19.3944
R9423 gnd.n2953 gnd.n2410 19.3944
R9424 gnd.n2953 gnd.n2952 19.3944
R9425 gnd.n2952 gnd.n2951 19.3944
R9426 gnd.n2951 gnd.n2418 19.3944
R9427 gnd.n2945 gnd.n2418 19.3944
R9428 gnd.n2945 gnd.n2944 19.3944
R9429 gnd.n2944 gnd.n2943 19.3944
R9430 gnd.n2943 gnd.n2426 19.3944
R9431 gnd.n2937 gnd.n2426 19.3944
R9432 gnd.n2937 gnd.n2936 19.3944
R9433 gnd.n2936 gnd.n2935 19.3944
R9434 gnd.n2935 gnd.n2434 19.3944
R9435 gnd.n2929 gnd.n2434 19.3944
R9436 gnd.n2929 gnd.n2928 19.3944
R9437 gnd.n2928 gnd.n2927 19.3944
R9438 gnd.n2927 gnd.n2442 19.3944
R9439 gnd.n2921 gnd.n2442 19.3944
R9440 gnd.n2921 gnd.n2920 19.3944
R9441 gnd.n2920 gnd.n2919 19.3944
R9442 gnd.n2919 gnd.n2450 19.3944
R9443 gnd.n2913 gnd.n2450 19.3944
R9444 gnd.n2913 gnd.n2912 19.3944
R9445 gnd.n2912 gnd.n2911 19.3944
R9446 gnd.n2911 gnd.n2458 19.3944
R9447 gnd.n2905 gnd.n2458 19.3944
R9448 gnd.n2905 gnd.n2904 19.3944
R9449 gnd.n2904 gnd.n2903 19.3944
R9450 gnd.n2903 gnd.n2466 19.3944
R9451 gnd.n2897 gnd.n2466 19.3944
R9452 gnd.n2897 gnd.n2896 19.3944
R9453 gnd.n2896 gnd.n2895 19.3944
R9454 gnd.n2895 gnd.n2474 19.3944
R9455 gnd.n2889 gnd.n2474 19.3944
R9456 gnd.n2889 gnd.n2888 19.3944
R9457 gnd.n2888 gnd.n2887 19.3944
R9458 gnd.n2887 gnd.n2482 19.3944
R9459 gnd.n2881 gnd.n2482 19.3944
R9460 gnd.n2881 gnd.n2880 19.3944
R9461 gnd.n2880 gnd.n2879 19.3944
R9462 gnd.n2879 gnd.n2490 19.3944
R9463 gnd.n2873 gnd.n2490 19.3944
R9464 gnd.n2873 gnd.n2872 19.3944
R9465 gnd.n2872 gnd.n2871 19.3944
R9466 gnd.n2871 gnd.n2498 19.3944
R9467 gnd.n2865 gnd.n2498 19.3944
R9468 gnd.n2865 gnd.n2864 19.3944
R9469 gnd.n2864 gnd.n2863 19.3944
R9470 gnd.n2863 gnd.n2506 19.3944
R9471 gnd.n2857 gnd.n2506 19.3944
R9472 gnd.n2857 gnd.n2856 19.3944
R9473 gnd.n2856 gnd.n2855 19.3944
R9474 gnd.n7207 gnd.n7206 19.3944
R9475 gnd.n7206 gnd.n527 19.3944
R9476 gnd.n805 gnd.n527 19.3944
R9477 gnd.n806 gnd.n805 19.3944
R9478 gnd.n809 gnd.n806 19.3944
R9479 gnd.n809 gnd.n800 19.3944
R9480 gnd.n815 gnd.n800 19.3944
R9481 gnd.n816 gnd.n815 19.3944
R9482 gnd.n819 gnd.n816 19.3944
R9483 gnd.n819 gnd.n798 19.3944
R9484 gnd.n825 gnd.n798 19.3944
R9485 gnd.n826 gnd.n825 19.3944
R9486 gnd.n829 gnd.n826 19.3944
R9487 gnd.n829 gnd.n796 19.3944
R9488 gnd.n835 gnd.n796 19.3944
R9489 gnd.n836 gnd.n835 19.3944
R9490 gnd.n839 gnd.n836 19.3944
R9491 gnd.n845 gnd.n842 19.3944
R9492 gnd.n848 gnd.n845 19.3944
R9493 gnd.n848 gnd.n790 19.3944
R9494 gnd.n852 gnd.n790 19.3944
R9495 gnd.n855 gnd.n852 19.3944
R9496 gnd.n858 gnd.n855 19.3944
R9497 gnd.n858 gnd.n787 19.3944
R9498 gnd.n958 gnd.n955 19.3944
R9499 gnd.n955 gnd.n954 19.3944
R9500 gnd.n954 gnd.n951 19.3944
R9501 gnd.n951 gnd.n950 19.3944
R9502 gnd.n950 gnd.n947 19.3944
R9503 gnd.n947 gnd.n946 19.3944
R9504 gnd.n946 gnd.n943 19.3944
R9505 gnd.n943 gnd.n942 19.3944
R9506 gnd.n938 gnd.n935 19.3944
R9507 gnd.n935 gnd.n934 19.3944
R9508 gnd.n934 gnd.n931 19.3944
R9509 gnd.n931 gnd.n930 19.3944
R9510 gnd.n930 gnd.n927 19.3944
R9511 gnd.n927 gnd.n926 19.3944
R9512 gnd.n926 gnd.n923 19.3944
R9513 gnd.n923 gnd.n922 19.3944
R9514 gnd.n922 gnd.n919 19.3944
R9515 gnd.n919 gnd.n918 19.3944
R9516 gnd.n918 gnd.n915 19.3944
R9517 gnd.n915 gnd.n914 19.3944
R9518 gnd.n914 gnd.n911 19.3944
R9519 gnd.n911 gnd.n910 19.3944
R9520 gnd.n910 gnd.n907 19.3944
R9521 gnd.n907 gnd.n906 19.3944
R9522 gnd.n906 gnd.n903 19.3944
R9523 gnd.n903 gnd.n902 19.3944
R9524 gnd.n7092 gnd.n512 19.3944
R9525 gnd.n7225 gnd.n512 19.3944
R9526 gnd.n7226 gnd.n7225 19.3944
R9527 gnd.n7229 gnd.n7226 19.3944
R9528 gnd.n7230 gnd.n7229 19.3944
R9529 gnd.n7233 gnd.n7230 19.3944
R9530 gnd.n7233 gnd.n7231 19.3944
R9531 gnd.n7231 gnd.n477 19.3944
R9532 gnd.n7275 gnd.n477 19.3944
R9533 gnd.n7276 gnd.n7275 19.3944
R9534 gnd.n7279 gnd.n7276 19.3944
R9535 gnd.n7279 gnd.n7277 19.3944
R9536 gnd.n7277 gnd.n442 19.3944
R9537 gnd.n7321 gnd.n442 19.3944
R9538 gnd.n7322 gnd.n7321 19.3944
R9539 gnd.n7325 gnd.n7322 19.3944
R9540 gnd.n7325 gnd.n7324 19.3944
R9541 gnd.n7324 gnd.n407 19.3944
R9542 gnd.n7367 gnd.n407 19.3944
R9543 gnd.n7368 gnd.n7367 19.3944
R9544 gnd.n7368 gnd.n381 19.3944
R9545 gnd.n7404 gnd.n381 19.3944
R9546 gnd.n7407 gnd.n7404 19.3944
R9547 gnd.n7407 gnd.n7406 19.3944
R9548 gnd.n7406 gnd.n366 19.3944
R9549 gnd.n7424 gnd.n366 19.3944
R9550 gnd.n7426 gnd.n7424 19.3944
R9551 gnd.n7426 gnd.n7425 19.3944
R9552 gnd.n7425 gnd.n359 19.3944
R9553 gnd.n7474 gnd.n359 19.3944
R9554 gnd.n7475 gnd.n7474 19.3944
R9555 gnd.n7477 gnd.n7475 19.3944
R9556 gnd.n7478 gnd.n7477 19.3944
R9557 gnd.n7481 gnd.n7478 19.3944
R9558 gnd.n7482 gnd.n7481 19.3944
R9559 gnd.n7484 gnd.n7482 19.3944
R9560 gnd.n7485 gnd.n7484 19.3944
R9561 gnd.n7488 gnd.n7485 19.3944
R9562 gnd.n7489 gnd.n7488 19.3944
R9563 gnd.n7491 gnd.n7489 19.3944
R9564 gnd.n7492 gnd.n7491 19.3944
R9565 gnd.n7495 gnd.n7492 19.3944
R9566 gnd.n7496 gnd.n7495 19.3944
R9567 gnd.n7512 gnd.n7496 19.3944
R9568 gnd.n7512 gnd.n7511 19.3944
R9569 gnd.n7511 gnd.n7510 19.3944
R9570 gnd.n7510 gnd.n7508 19.3944
R9571 gnd.n7508 gnd.n7507 19.3944
R9572 gnd.n7507 gnd.n7505 19.3944
R9573 gnd.n7505 gnd.n7504 19.3944
R9574 gnd.n7504 gnd.n7502 19.3944
R9575 gnd.n7502 gnd.n7501 19.3944
R9576 gnd.n7501 gnd.n7499 19.3944
R9577 gnd.n7095 gnd.n7091 19.3944
R9578 gnd.n7095 gnd.n507 19.3944
R9579 gnd.n7239 gnd.n507 19.3944
R9580 gnd.n7239 gnd.n7238 19.3944
R9581 gnd.n7238 gnd.n7237 19.3944
R9582 gnd.n7237 gnd.n7236 19.3944
R9583 gnd.n7236 gnd.n472 19.3944
R9584 gnd.n7285 gnd.n472 19.3944
R9585 gnd.n7285 gnd.n7284 19.3944
R9586 gnd.n7284 gnd.n7283 19.3944
R9587 gnd.n7283 gnd.n7282 19.3944
R9588 gnd.n7282 gnd.n437 19.3944
R9589 gnd.n7332 gnd.n437 19.3944
R9590 gnd.n7332 gnd.n7331 19.3944
R9591 gnd.n7331 gnd.n7330 19.3944
R9592 gnd.n7330 gnd.n7329 19.3944
R9593 gnd.n7329 gnd.n404 19.3944
R9594 gnd.n7376 gnd.n404 19.3944
R9595 gnd.n7376 gnd.n7375 19.3944
R9596 gnd.n7375 gnd.n7374 19.3944
R9597 gnd.n7374 gnd.n7373 19.3944
R9598 gnd.n7373 gnd.n379 19.3944
R9599 gnd.n7409 gnd.n379 19.3944
R9600 gnd.n7409 gnd.n368 19.3944
R9601 gnd.n7421 gnd.n368 19.3944
R9602 gnd.n7421 gnd.n361 19.3944
R9603 gnd.n7430 gnd.n361 19.3944
R9604 gnd.n7431 gnd.n7430 19.3944
R9605 gnd.n7433 gnd.n7431 19.3944
R9606 gnd.n7433 gnd.n110 19.3944
R9607 gnd.n7743 gnd.n110 19.3944
R9608 gnd.n7743 gnd.n7742 19.3944
R9609 gnd.n7742 gnd.n7741 19.3944
R9610 gnd.n7741 gnd.n114 19.3944
R9611 gnd.n7731 gnd.n114 19.3944
R9612 gnd.n7731 gnd.n7730 19.3944
R9613 gnd.n7730 gnd.n7729 19.3944
R9614 gnd.n7729 gnd.n131 19.3944
R9615 gnd.n7719 gnd.n131 19.3944
R9616 gnd.n7719 gnd.n7718 19.3944
R9617 gnd.n7718 gnd.n7717 19.3944
R9618 gnd.n7717 gnd.n151 19.3944
R9619 gnd.n7707 gnd.n151 19.3944
R9620 gnd.n7707 gnd.n7706 19.3944
R9621 gnd.n7706 gnd.n7705 19.3944
R9622 gnd.n7705 gnd.n169 19.3944
R9623 gnd.n7695 gnd.n169 19.3944
R9624 gnd.n7695 gnd.n7694 19.3944
R9625 gnd.n7694 gnd.n7693 19.3944
R9626 gnd.n7693 gnd.n189 19.3944
R9627 gnd.n7683 gnd.n189 19.3944
R9628 gnd.n7683 gnd.n7682 19.3944
R9629 gnd.n7682 gnd.n7681 19.3944
R9630 gnd.n7603 gnd.n278 19.3944
R9631 gnd.n7603 gnd.n282 19.3944
R9632 gnd.n285 gnd.n282 19.3944
R9633 gnd.n7596 gnd.n285 19.3944
R9634 gnd.n7596 gnd.n7595 19.3944
R9635 gnd.n7595 gnd.n7594 19.3944
R9636 gnd.n7594 gnd.n291 19.3944
R9637 gnd.n7589 gnd.n291 19.3944
R9638 gnd.n7589 gnd.n7588 19.3944
R9639 gnd.n7588 gnd.n7587 19.3944
R9640 gnd.n7587 gnd.n298 19.3944
R9641 gnd.n7582 gnd.n298 19.3944
R9642 gnd.n7582 gnd.n7581 19.3944
R9643 gnd.n7581 gnd.n7580 19.3944
R9644 gnd.n7580 gnd.n305 19.3944
R9645 gnd.n7575 gnd.n305 19.3944
R9646 gnd.n7575 gnd.n7574 19.3944
R9647 gnd.n7574 gnd.n7573 19.3944
R9648 gnd.n7641 gnd.n245 19.3944
R9649 gnd.n7636 gnd.n245 19.3944
R9650 gnd.n7636 gnd.n7635 19.3944
R9651 gnd.n7635 gnd.n7634 19.3944
R9652 gnd.n7634 gnd.n252 19.3944
R9653 gnd.n7629 gnd.n252 19.3944
R9654 gnd.n7629 gnd.n7628 19.3944
R9655 gnd.n7628 gnd.n7627 19.3944
R9656 gnd.n7627 gnd.n259 19.3944
R9657 gnd.n7622 gnd.n259 19.3944
R9658 gnd.n7622 gnd.n7621 19.3944
R9659 gnd.n7621 gnd.n7620 19.3944
R9660 gnd.n7620 gnd.n266 19.3944
R9661 gnd.n7615 gnd.n266 19.3944
R9662 gnd.n7615 gnd.n7614 19.3944
R9663 gnd.n7614 gnd.n7613 19.3944
R9664 gnd.n7613 gnd.n273 19.3944
R9665 gnd.n7608 gnd.n273 19.3944
R9666 gnd.n7674 gnd.n7673 19.3944
R9667 gnd.n7673 gnd.n7672 19.3944
R9668 gnd.n7672 gnd.n217 19.3944
R9669 gnd.n7667 gnd.n217 19.3944
R9670 gnd.n7667 gnd.n7666 19.3944
R9671 gnd.n7666 gnd.n7665 19.3944
R9672 gnd.n7665 gnd.n224 19.3944
R9673 gnd.n7660 gnd.n224 19.3944
R9674 gnd.n7660 gnd.n7659 19.3944
R9675 gnd.n7659 gnd.n7658 19.3944
R9676 gnd.n7658 gnd.n231 19.3944
R9677 gnd.n7653 gnd.n231 19.3944
R9678 gnd.n7653 gnd.n7652 19.3944
R9679 gnd.n7652 gnd.n7651 19.3944
R9680 gnd.n7651 gnd.n238 19.3944
R9681 gnd.n7646 gnd.n238 19.3944
R9682 gnd.n7646 gnd.n7645 19.3944
R9683 gnd.n7564 gnd.n7563 19.3944
R9684 gnd.n7563 gnd.n7562 19.3944
R9685 gnd.n7562 gnd.n320 19.3944
R9686 gnd.n7557 gnd.n320 19.3944
R9687 gnd.n7557 gnd.n7556 19.3944
R9688 gnd.n7556 gnd.n7555 19.3944
R9689 gnd.n7555 gnd.n327 19.3944
R9690 gnd.n7550 gnd.n327 19.3944
R9691 gnd.n7550 gnd.n7549 19.3944
R9692 gnd.n7549 gnd.n7548 19.3944
R9693 gnd.n7548 gnd.n334 19.3944
R9694 gnd.n7543 gnd.n334 19.3944
R9695 gnd.n7543 gnd.n7542 19.3944
R9696 gnd.n7542 gnd.n7541 19.3944
R9697 gnd.n7541 gnd.n341 19.3944
R9698 gnd.n7536 gnd.n341 19.3944
R9699 gnd.n7216 gnd.n516 19.3944
R9700 gnd.n7221 gnd.n516 19.3944
R9701 gnd.n7221 gnd.n517 19.3944
R9702 gnd.n517 gnd.n489 19.3944
R9703 gnd.n7253 gnd.n489 19.3944
R9704 gnd.n7253 gnd.n486 19.3944
R9705 gnd.n7258 gnd.n486 19.3944
R9706 gnd.n7258 gnd.n487 19.3944
R9707 gnd.n487 gnd.n455 19.3944
R9708 gnd.n7299 gnd.n455 19.3944
R9709 gnd.n7299 gnd.n452 19.3944
R9710 gnd.n7304 gnd.n452 19.3944
R9711 gnd.n7304 gnd.n453 19.3944
R9712 gnd.n453 gnd.n420 19.3944
R9713 gnd.n7346 gnd.n420 19.3944
R9714 gnd.n7346 gnd.n417 19.3944
R9715 gnd.n7351 gnd.n417 19.3944
R9716 gnd.n7351 gnd.n418 19.3944
R9717 gnd.n418 gnd.n388 19.3944
R9718 gnd.n7390 gnd.n388 19.3944
R9719 gnd.n7390 gnd.n385 19.3944
R9720 gnd.n7400 gnd.n385 19.3944
R9721 gnd.n7400 gnd.n386 19.3944
R9722 gnd.n7396 gnd.n386 19.3944
R9723 gnd.n7396 gnd.n7395 19.3944
R9724 gnd.n7395 gnd.n85 19.3944
R9725 gnd.n7756 gnd.n85 19.3944
R9726 gnd.n7756 gnd.n7755 19.3944
R9727 gnd.n7755 gnd.n87 19.3944
R9728 gnd.n7470 gnd.n87 19.3944
R9729 gnd.n7470 gnd.n7469 19.3944
R9730 gnd.n7469 gnd.n7468 19.3944
R9731 gnd.n7468 gnd.n7466 19.3944
R9732 gnd.n7466 gnd.n7465 19.3944
R9733 gnd.n7465 gnd.n7463 19.3944
R9734 gnd.n7463 gnd.n7462 19.3944
R9735 gnd.n7462 gnd.n7460 19.3944
R9736 gnd.n7460 gnd.n7459 19.3944
R9737 gnd.n7459 gnd.n7457 19.3944
R9738 gnd.n7457 gnd.n7456 19.3944
R9739 gnd.n7456 gnd.n7454 19.3944
R9740 gnd.n7454 gnd.n7453 19.3944
R9741 gnd.n7453 gnd.n358 19.3944
R9742 gnd.n7516 gnd.n358 19.3944
R9743 gnd.n7517 gnd.n7516 19.3944
R9744 gnd.n7517 gnd.n356 19.3944
R9745 gnd.n7521 gnd.n356 19.3944
R9746 gnd.n7523 gnd.n7521 19.3944
R9747 gnd.n7524 gnd.n7523 19.3944
R9748 gnd.n7524 gnd.n353 19.3944
R9749 gnd.n7528 gnd.n353 19.3944
R9750 gnd.n7530 gnd.n7528 19.3944
R9751 gnd.n7531 gnd.n7530 19.3944
R9752 gnd.n7212 gnd.n7211 19.3944
R9753 gnd.n7211 gnd.n499 19.3944
R9754 gnd.n7243 gnd.n499 19.3944
R9755 gnd.n7243 gnd.n497 19.3944
R9756 gnd.n7249 gnd.n497 19.3944
R9757 gnd.n7249 gnd.n7248 19.3944
R9758 gnd.n7248 gnd.n464 19.3944
R9759 gnd.n7289 gnd.n464 19.3944
R9760 gnd.n7289 gnd.n462 19.3944
R9761 gnd.n7295 gnd.n462 19.3944
R9762 gnd.n7295 gnd.n7294 19.3944
R9763 gnd.n7294 gnd.n429 19.3944
R9764 gnd.n7336 gnd.n429 19.3944
R9765 gnd.n7336 gnd.n427 19.3944
R9766 gnd.n7342 gnd.n427 19.3944
R9767 gnd.n7342 gnd.n7341 19.3944
R9768 gnd.n7341 gnd.n397 19.3944
R9769 gnd.n7380 gnd.n397 19.3944
R9770 gnd.n7380 gnd.n395 19.3944
R9771 gnd.n7386 gnd.n395 19.3944
R9772 gnd.n7386 gnd.n7385 19.3944
R9773 gnd.n7385 gnd.n7384 19.3944
R9774 gnd.n375 gnd.n100 19.3944
R9775 gnd.n7417 gnd.n100 19.3944
R9776 gnd.n7415 gnd.n7414 19.3944
R9777 gnd.n7751 gnd.n7750 19.3944
R9778 gnd.n7747 gnd.n95 19.3944
R9779 gnd.n7747 gnd.n102 19.3944
R9780 gnd.n7737 gnd.n102 19.3944
R9781 gnd.n7737 gnd.n7736 19.3944
R9782 gnd.n7736 gnd.n7735 19.3944
R9783 gnd.n7735 gnd.n122 19.3944
R9784 gnd.n7725 gnd.n122 19.3944
R9785 gnd.n7725 gnd.n7724 19.3944
R9786 gnd.n7724 gnd.n7723 19.3944
R9787 gnd.n7723 gnd.n142 19.3944
R9788 gnd.n7713 gnd.n142 19.3944
R9789 gnd.n7713 gnd.n7712 19.3944
R9790 gnd.n7712 gnd.n7711 19.3944
R9791 gnd.n7711 gnd.n160 19.3944
R9792 gnd.n7701 gnd.n160 19.3944
R9793 gnd.n7701 gnd.n7700 19.3944
R9794 gnd.n7700 gnd.n7699 19.3944
R9795 gnd.n7699 gnd.n180 19.3944
R9796 gnd.n7689 gnd.n180 19.3944
R9797 gnd.n7689 gnd.n7688 19.3944
R9798 gnd.n7688 gnd.n7687 19.3944
R9799 gnd.n7687 gnd.n199 19.3944
R9800 gnd.n7677 gnd.n199 19.3944
R9801 gnd.n5085 gnd.n5084 19.3944
R9802 gnd.n5084 gnd.n5083 19.3944
R9803 gnd.n5083 gnd.n5082 19.3944
R9804 gnd.n5082 gnd.n5080 19.3944
R9805 gnd.n5080 gnd.n5077 19.3944
R9806 gnd.n5077 gnd.n5076 19.3944
R9807 gnd.n5076 gnd.n5073 19.3944
R9808 gnd.n5073 gnd.n5072 19.3944
R9809 gnd.n5072 gnd.n5069 19.3944
R9810 gnd.n5069 gnd.n5068 19.3944
R9811 gnd.n5068 gnd.n5065 19.3944
R9812 gnd.n5065 gnd.n5064 19.3944
R9813 gnd.n5064 gnd.n5061 19.3944
R9814 gnd.n5061 gnd.n5060 19.3944
R9815 gnd.n5060 gnd.n5057 19.3944
R9816 gnd.n5057 gnd.n5056 19.3944
R9817 gnd.n5056 gnd.n5053 19.3944
R9818 gnd.n5051 gnd.n5048 19.3944
R9819 gnd.n5048 gnd.n5047 19.3944
R9820 gnd.n5047 gnd.n5044 19.3944
R9821 gnd.n5044 gnd.n5043 19.3944
R9822 gnd.n5043 gnd.n5040 19.3944
R9823 gnd.n5040 gnd.n5039 19.3944
R9824 gnd.n5039 gnd.n5036 19.3944
R9825 gnd.n5036 gnd.n5035 19.3944
R9826 gnd.n5035 gnd.n5032 19.3944
R9827 gnd.n5032 gnd.n5031 19.3944
R9828 gnd.n5031 gnd.n5028 19.3944
R9829 gnd.n5028 gnd.n5027 19.3944
R9830 gnd.n5027 gnd.n5024 19.3944
R9831 gnd.n5024 gnd.n5023 19.3944
R9832 gnd.n5023 gnd.n5020 19.3944
R9833 gnd.n5020 gnd.n5019 19.3944
R9834 gnd.n5019 gnd.n5016 19.3944
R9835 gnd.n5016 gnd.n5015 19.3944
R9836 gnd.n5011 gnd.n5008 19.3944
R9837 gnd.n5008 gnd.n5007 19.3944
R9838 gnd.n5007 gnd.n5004 19.3944
R9839 gnd.n5004 gnd.n5003 19.3944
R9840 gnd.n5003 gnd.n5000 19.3944
R9841 gnd.n5000 gnd.n4999 19.3944
R9842 gnd.n4999 gnd.n4996 19.3944
R9843 gnd.n4996 gnd.n4995 19.3944
R9844 gnd.n4995 gnd.n4992 19.3944
R9845 gnd.n4992 gnd.n4991 19.3944
R9846 gnd.n4991 gnd.n4988 19.3944
R9847 gnd.n4988 gnd.n4987 19.3944
R9848 gnd.n4987 gnd.n4984 19.3944
R9849 gnd.n4984 gnd.n4983 19.3944
R9850 gnd.n4983 gnd.n4980 19.3944
R9851 gnd.n4980 gnd.n4979 19.3944
R9852 gnd.n4979 gnd.n4976 19.3944
R9853 gnd.n4976 gnd.n4975 19.3944
R9854 gnd.n4968 gnd.n4966 19.3944
R9855 gnd.n4966 gnd.n4963 19.3944
R9856 gnd.n4963 gnd.n4962 19.3944
R9857 gnd.n4962 gnd.n4959 19.3944
R9858 gnd.n4959 gnd.n4958 19.3944
R9859 gnd.n4958 gnd.n4955 19.3944
R9860 gnd.n4955 gnd.n4954 19.3944
R9861 gnd.n4954 gnd.n4951 19.3944
R9862 gnd.n4951 gnd.n4950 19.3944
R9863 gnd.n4950 gnd.n4947 19.3944
R9864 gnd.n4947 gnd.n4946 19.3944
R9865 gnd.n4946 gnd.n4943 19.3944
R9866 gnd.n4943 gnd.n4942 19.3944
R9867 gnd.n4942 gnd.n4939 19.3944
R9868 gnd.n4939 gnd.n4938 19.3944
R9869 gnd.n4938 gnd.n4935 19.3944
R9870 gnd.n4929 gnd.n4927 19.3944
R9871 gnd.n4927 gnd.n4926 19.3944
R9872 gnd.n4926 gnd.n4924 19.3944
R9873 gnd.n4924 gnd.n4923 19.3944
R9874 gnd.n4923 gnd.n4921 19.3944
R9875 gnd.n4921 gnd.n4920 19.3944
R9876 gnd.n4920 gnd.n4918 19.3944
R9877 gnd.n4918 gnd.n4917 19.3944
R9878 gnd.n4917 gnd.n4915 19.3944
R9879 gnd.n4915 gnd.n4914 19.3944
R9880 gnd.n4914 gnd.n4912 19.3944
R9881 gnd.n4912 gnd.n4911 19.3944
R9882 gnd.n4911 gnd.n4909 19.3944
R9883 gnd.n4909 gnd.n1913 19.3944
R9884 gnd.n5174 gnd.n1913 19.3944
R9885 gnd.n5174 gnd.n1911 19.3944
R9886 gnd.n5180 gnd.n1911 19.3944
R9887 gnd.n5180 gnd.n5179 19.3944
R9888 gnd.n5179 gnd.n1888 19.3944
R9889 gnd.n5209 gnd.n1888 19.3944
R9890 gnd.n5209 gnd.n1886 19.3944
R9891 gnd.n5224 gnd.n1886 19.3944
R9892 gnd.n5224 gnd.n5223 19.3944
R9893 gnd.n5223 gnd.n5222 19.3944
R9894 gnd.n5222 gnd.n5220 19.3944
R9895 gnd.n5220 gnd.n5219 19.3944
R9896 gnd.n5219 gnd.n1855 19.3944
R9897 gnd.n5263 gnd.n1855 19.3944
R9898 gnd.n5263 gnd.n1852 19.3944
R9899 gnd.n5268 gnd.n1852 19.3944
R9900 gnd.n5268 gnd.n1853 19.3944
R9901 gnd.n1853 gnd.n1819 19.3944
R9902 gnd.n5305 gnd.n1819 19.3944
R9903 gnd.n5305 gnd.n1816 19.3944
R9904 gnd.n5310 gnd.n1816 19.3944
R9905 gnd.n5310 gnd.n1817 19.3944
R9906 gnd.n1817 gnd.n1784 19.3944
R9907 gnd.n5345 gnd.n1784 19.3944
R9908 gnd.n5345 gnd.n1781 19.3944
R9909 gnd.n5350 gnd.n1781 19.3944
R9910 gnd.n5350 gnd.n1782 19.3944
R9911 gnd.n1782 gnd.n1749 19.3944
R9912 gnd.n5393 gnd.n1749 19.3944
R9913 gnd.n5393 gnd.n1746 19.3944
R9914 gnd.n5401 gnd.n1746 19.3944
R9915 gnd.n5401 gnd.n1747 19.3944
R9916 gnd.n5397 gnd.n1747 19.3944
R9917 gnd.n5397 gnd.n1676 19.3944
R9918 gnd.n5750 gnd.n1676 19.3944
R9919 gnd.n5750 gnd.n1677 19.3944
R9920 gnd.n5746 gnd.n1677 19.3944
R9921 gnd.n5746 gnd.n5745 19.3944
R9922 gnd.n5745 gnd.n5744 19.3944
R9923 gnd.n5094 gnd.n5092 19.3944
R9924 gnd.n5094 gnd.n5093 19.3944
R9925 gnd.n5093 gnd.n1968 19.3944
R9926 gnd.n5109 gnd.n1968 19.3944
R9927 gnd.n5110 gnd.n5109 19.3944
R9928 gnd.n5111 gnd.n5110 19.3944
R9929 gnd.n5111 gnd.n1950 19.3944
R9930 gnd.n5129 gnd.n1950 19.3944
R9931 gnd.n5130 gnd.n5129 19.3944
R9932 gnd.n5131 gnd.n5130 19.3944
R9933 gnd.n5131 gnd.n1932 19.3944
R9934 gnd.n5149 gnd.n1932 19.3944
R9935 gnd.n5150 gnd.n5149 19.3944
R9936 gnd.n5152 gnd.n5150 19.3944
R9937 gnd.n5153 gnd.n5152 19.3944
R9938 gnd.n5153 gnd.n1906 19.3944
R9939 gnd.n5184 gnd.n1906 19.3944
R9940 gnd.n5185 gnd.n5184 19.3944
R9941 gnd.n5187 gnd.n5185 19.3944
R9942 gnd.n5188 gnd.n5187 19.3944
R9943 gnd.n5188 gnd.n1881 19.3944
R9944 gnd.n5228 gnd.n1881 19.3944
R9945 gnd.n5229 gnd.n5228 19.3944
R9946 gnd.n5230 gnd.n5229 19.3944
R9947 gnd.n5230 gnd.n1867 19.3944
R9948 gnd.n5245 gnd.n1867 19.3944
R9949 gnd.n5246 gnd.n5245 19.3944
R9950 gnd.n5247 gnd.n5246 19.3944
R9951 gnd.n5247 gnd.n1847 19.3944
R9952 gnd.n5272 gnd.n1847 19.3944
R9953 gnd.n5273 gnd.n5272 19.3944
R9954 gnd.n5276 gnd.n5273 19.3944
R9955 gnd.n5277 gnd.n5276 19.3944
R9956 gnd.n5285 gnd.n5277 19.3944
R9957 gnd.n5285 gnd.n5283 19.3944
R9958 gnd.n5283 gnd.n5282 19.3944
R9959 gnd.n5282 gnd.n5281 19.3944
R9960 gnd.n5281 gnd.n5278 19.3944
R9961 gnd.n5278 gnd.n1776 19.3944
R9962 gnd.n5354 gnd.n1776 19.3944
R9963 gnd.n5355 gnd.n5354 19.3944
R9964 gnd.n5357 gnd.n5355 19.3944
R9965 gnd.n5357 gnd.n5356 19.3944
R9966 gnd.n5356 gnd.n1741 19.3944
R9967 gnd.n5405 gnd.n1741 19.3944
R9968 gnd.n5406 gnd.n5405 19.3944
R9969 gnd.n5408 gnd.n5406 19.3944
R9970 gnd.n5408 gnd.n1672 19.3944
R9971 gnd.n5754 gnd.n1672 19.3944
R9972 gnd.n5755 gnd.n5754 19.3944
R9973 gnd.n5755 gnd.n1652 19.3944
R9974 gnd.n5866 gnd.n1652 19.3944
R9975 gnd.n5867 gnd.n5866 19.3944
R9976 gnd.n5096 gnd.n1984 19.3944
R9977 gnd.n5096 gnd.n1985 19.3944
R9978 gnd.n1987 gnd.n1985 19.3944
R9979 gnd.n1987 gnd.n1966 19.3944
R9980 gnd.n5116 gnd.n1966 19.3944
R9981 gnd.n5116 gnd.n5115 19.3944
R9982 gnd.n5115 gnd.n5114 19.3944
R9983 gnd.n5114 gnd.n1948 19.3944
R9984 gnd.n5136 gnd.n1948 19.3944
R9985 gnd.n5136 gnd.n5135 19.3944
R9986 gnd.n5135 gnd.n5134 19.3944
R9987 gnd.n5134 gnd.n1929 19.3944
R9988 gnd.n5160 gnd.n1929 19.3944
R9989 gnd.n5160 gnd.n5159 19.3944
R9990 gnd.n5159 gnd.n5158 19.3944
R9991 gnd.n5158 gnd.n5157 19.3944
R9992 gnd.n5157 gnd.n1903 19.3944
R9993 gnd.n5195 gnd.n1903 19.3944
R9994 gnd.n5195 gnd.n5194 19.3944
R9995 gnd.n5194 gnd.n5193 19.3944
R9996 gnd.n5193 gnd.n5192 19.3944
R9997 gnd.n5192 gnd.n1879 19.3944
R9998 gnd.n5235 gnd.n1879 19.3944
R9999 gnd.n5235 gnd.n5234 19.3944
R10000 gnd.n5234 gnd.n5233 19.3944
R10001 gnd.n5233 gnd.n1865 19.3944
R10002 gnd.n5253 gnd.n1865 19.3944
R10003 gnd.n5253 gnd.n5252 19.3944
R10004 gnd.n5252 gnd.n5251 19.3944
R10005 gnd.n5251 gnd.n1842 19.3944
R10006 gnd.n5291 gnd.n1842 19.3944
R10007 gnd.n5291 gnd.n5290 19.3944
R10008 gnd.n5290 gnd.n5289 19.3944
R10009 gnd.n5289 gnd.n5288 19.3944
R10010 gnd.n5288 gnd.n1801 19.3944
R10011 gnd.n5331 gnd.n1801 19.3944
R10012 gnd.n5331 gnd.n5330 19.3944
R10013 gnd.n5330 gnd.n5329 19.3944
R10014 gnd.n5329 gnd.n5328 19.3944
R10015 gnd.n5328 gnd.n1765 19.3944
R10016 gnd.n5379 gnd.n1765 19.3944
R10017 gnd.n5379 gnd.n5378 19.3944
R10018 gnd.n5378 gnd.n5377 19.3944
R10019 gnd.n5377 gnd.n5376 19.3944
R10020 gnd.n5376 gnd.n1739 19.3944
R10021 gnd.n5413 gnd.n1739 19.3944
R10022 gnd.n5413 gnd.n5412 19.3944
R10023 gnd.n5412 gnd.n5411 19.3944
R10024 gnd.n5411 gnd.n1670 19.3944
R10025 gnd.n5760 gnd.n1670 19.3944
R10026 gnd.n5760 gnd.n5759 19.3944
R10027 gnd.n5759 gnd.n5758 19.3944
R10028 gnd.n5758 gnd.n1651 19.3944
R10029 gnd.n5858 gnd.n5769 19.3944
R10030 gnd.n5853 gnd.n5769 19.3944
R10031 gnd.n5853 gnd.n5852 19.3944
R10032 gnd.n5852 gnd.n5851 19.3944
R10033 gnd.n5851 gnd.n5774 19.3944
R10034 gnd.n5846 gnd.n5774 19.3944
R10035 gnd.n5846 gnd.n5845 19.3944
R10036 gnd.n5845 gnd.n5844 19.3944
R10037 gnd.n5844 gnd.n5781 19.3944
R10038 gnd.n5839 gnd.n5781 19.3944
R10039 gnd.n5839 gnd.n5838 19.3944
R10040 gnd.n5838 gnd.n5837 19.3944
R10041 gnd.n5837 gnd.n5788 19.3944
R10042 gnd.n5832 gnd.n5788 19.3944
R10043 gnd.n5832 gnd.n5831 19.3944
R10044 gnd.n5831 gnd.n5830 19.3944
R10045 gnd.n5830 gnd.n5795 19.3944
R10046 gnd.n5906 gnd.n1609 19.3944
R10047 gnd.n5906 gnd.n1613 19.3944
R10048 gnd.n1616 gnd.n1613 19.3944
R10049 gnd.n5899 gnd.n1616 19.3944
R10050 gnd.n5899 gnd.n5898 19.3944
R10051 gnd.n5898 gnd.n5897 19.3944
R10052 gnd.n5897 gnd.n1622 19.3944
R10053 gnd.n5892 gnd.n1622 19.3944
R10054 gnd.n5892 gnd.n5891 19.3944
R10055 gnd.n5891 gnd.n5890 19.3944
R10056 gnd.n5890 gnd.n1629 19.3944
R10057 gnd.n5885 gnd.n1629 19.3944
R10058 gnd.n5885 gnd.n5884 19.3944
R10059 gnd.n5884 gnd.n5883 19.3944
R10060 gnd.n5883 gnd.n1636 19.3944
R10061 gnd.n5878 gnd.n1636 19.3944
R10062 gnd.n5878 gnd.n5877 19.3944
R10063 gnd.n5877 gnd.n5876 19.3944
R10064 gnd.n5925 gnd.n1589 19.3944
R10065 gnd.n5925 gnd.n1594 19.3944
R10066 gnd.n1598 gnd.n1594 19.3944
R10067 gnd.n5918 gnd.n1598 19.3944
R10068 gnd.n5918 gnd.n5917 19.3944
R10069 gnd.n5917 gnd.n5916 19.3944
R10070 gnd.n5916 gnd.n1604 19.3944
R10071 gnd.n5911 gnd.n1604 19.3944
R10072 gnd.n5825 gnd.n5824 19.3944
R10073 gnd.n5824 gnd.n5823 19.3944
R10074 gnd.n5823 gnd.n5805 19.3944
R10075 gnd.n5818 gnd.n5805 19.3944
R10076 gnd.n5818 gnd.n5817 19.3944
R10077 gnd.n5817 gnd.n5816 19.3944
R10078 gnd.n5816 gnd.n1590 19.3944
R10079 gnd.n5100 gnd.n1977 19.3944
R10080 gnd.n5100 gnd.n1975 19.3944
R10081 gnd.n5104 gnd.n1975 19.3944
R10082 gnd.n5104 gnd.n1958 19.3944
R10083 gnd.n5120 gnd.n1958 19.3944
R10084 gnd.n5120 gnd.n1956 19.3944
R10085 gnd.n5124 gnd.n1956 19.3944
R10086 gnd.n5124 gnd.n1941 19.3944
R10087 gnd.n5140 gnd.n1941 19.3944
R10088 gnd.n5140 gnd.n1939 19.3944
R10089 gnd.n5144 gnd.n1939 19.3944
R10090 gnd.n5144 gnd.n1921 19.3944
R10091 gnd.n5164 gnd.n1921 19.3944
R10092 gnd.n5164 gnd.n1919 19.3944
R10093 gnd.n5170 gnd.n1919 19.3944
R10094 gnd.n5170 gnd.n5169 19.3944
R10095 gnd.n5169 gnd.n1896 19.3944
R10096 gnd.n5199 gnd.n1896 19.3944
R10097 gnd.n5199 gnd.n1894 19.3944
R10098 gnd.n5205 gnd.n1894 19.3944
R10099 gnd.n5205 gnd.n5204 19.3944
R10100 gnd.n5204 gnd.n5203 19.3944
R10101 gnd.n1874 gnd.n1833 19.3944
R10102 gnd.n5240 gnd.n1833 19.3944
R10103 gnd.n1861 gnd.n1860 19.3944
R10104 gnd.n5259 gnd.n5258 19.3944
R10105 gnd.n5295 gnd.n1835 19.3944
R10106 gnd.n5295 gnd.n1827 19.3944
R10107 gnd.n5301 gnd.n1827 19.3944
R10108 gnd.n5301 gnd.n5300 19.3944
R10109 gnd.n5300 gnd.n1793 19.3944
R10110 gnd.n5335 gnd.n1793 19.3944
R10111 gnd.n5335 gnd.n1791 19.3944
R10112 gnd.n5341 gnd.n1791 19.3944
R10113 gnd.n5341 gnd.n5340 19.3944
R10114 gnd.n5340 gnd.n1758 19.3944
R10115 gnd.n5383 gnd.n1758 19.3944
R10116 gnd.n5383 gnd.n1756 19.3944
R10117 gnd.n5389 gnd.n1756 19.3944
R10118 gnd.n5389 gnd.n5388 19.3944
R10119 gnd.n5388 gnd.n1731 19.3944
R10120 gnd.n5417 gnd.n1731 19.3944
R10121 gnd.n5417 gnd.n1729 19.3944
R10122 gnd.n5421 gnd.n1729 19.3944
R10123 gnd.n5421 gnd.n1662 19.3944
R10124 gnd.n5764 gnd.n1662 19.3944
R10125 gnd.n5764 gnd.n1660 19.3944
R10126 gnd.n5862 gnd.n1660 19.3944
R10127 gnd.n5862 gnd.n5861 19.3944
R10128 gnd.n3169 gnd.n2205 19.3944
R10129 gnd.n3169 gnd.n2203 19.3944
R10130 gnd.n3173 gnd.n2203 19.3944
R10131 gnd.n3173 gnd.n2199 19.3944
R10132 gnd.n3179 gnd.n2199 19.3944
R10133 gnd.n3179 gnd.n2197 19.3944
R10134 gnd.n3183 gnd.n2197 19.3944
R10135 gnd.n3183 gnd.n2193 19.3944
R10136 gnd.n3189 gnd.n2193 19.3944
R10137 gnd.n3189 gnd.n2191 19.3944
R10138 gnd.n3193 gnd.n2191 19.3944
R10139 gnd.n3193 gnd.n2187 19.3944
R10140 gnd.n3199 gnd.n2187 19.3944
R10141 gnd.n3199 gnd.n2185 19.3944
R10142 gnd.n3203 gnd.n2185 19.3944
R10143 gnd.n3203 gnd.n2181 19.3944
R10144 gnd.n3209 gnd.n2181 19.3944
R10145 gnd.n3209 gnd.n2179 19.3944
R10146 gnd.n3213 gnd.n2179 19.3944
R10147 gnd.n3213 gnd.n2175 19.3944
R10148 gnd.n3219 gnd.n2175 19.3944
R10149 gnd.n3219 gnd.n2173 19.3944
R10150 gnd.n3223 gnd.n2173 19.3944
R10151 gnd.n3223 gnd.n2169 19.3944
R10152 gnd.n3229 gnd.n2169 19.3944
R10153 gnd.n3229 gnd.n2167 19.3944
R10154 gnd.n3233 gnd.n2167 19.3944
R10155 gnd.n3233 gnd.n2163 19.3944
R10156 gnd.n3239 gnd.n2163 19.3944
R10157 gnd.n3239 gnd.n2161 19.3944
R10158 gnd.n3243 gnd.n2161 19.3944
R10159 gnd.n3243 gnd.n2157 19.3944
R10160 gnd.n3249 gnd.n2157 19.3944
R10161 gnd.n3249 gnd.n2155 19.3944
R10162 gnd.n3253 gnd.n2155 19.3944
R10163 gnd.n3253 gnd.n2151 19.3944
R10164 gnd.n3259 gnd.n2151 19.3944
R10165 gnd.n3259 gnd.n2149 19.3944
R10166 gnd.n3263 gnd.n2149 19.3944
R10167 gnd.n3263 gnd.n2145 19.3944
R10168 gnd.n3269 gnd.n2145 19.3944
R10169 gnd.n3269 gnd.n2143 19.3944
R10170 gnd.n3273 gnd.n2143 19.3944
R10171 gnd.n3273 gnd.n2139 19.3944
R10172 gnd.n3279 gnd.n2139 19.3944
R10173 gnd.n3279 gnd.n2137 19.3944
R10174 gnd.n3283 gnd.n2137 19.3944
R10175 gnd.n3283 gnd.n2133 19.3944
R10176 gnd.n3289 gnd.n2133 19.3944
R10177 gnd.n3289 gnd.n2131 19.3944
R10178 gnd.n3293 gnd.n2131 19.3944
R10179 gnd.n3293 gnd.n2127 19.3944
R10180 gnd.n3299 gnd.n2127 19.3944
R10181 gnd.n3299 gnd.n2125 19.3944
R10182 gnd.n3303 gnd.n2125 19.3944
R10183 gnd.n3303 gnd.n2121 19.3944
R10184 gnd.n3309 gnd.n2121 19.3944
R10185 gnd.n3309 gnd.n2119 19.3944
R10186 gnd.n3313 gnd.n2119 19.3944
R10187 gnd.n3313 gnd.n2115 19.3944
R10188 gnd.n3319 gnd.n2115 19.3944
R10189 gnd.n3319 gnd.n2113 19.3944
R10190 gnd.n3323 gnd.n2113 19.3944
R10191 gnd.n3323 gnd.n2109 19.3944
R10192 gnd.n3329 gnd.n2109 19.3944
R10193 gnd.n3329 gnd.n2107 19.3944
R10194 gnd.n3333 gnd.n2107 19.3944
R10195 gnd.n3333 gnd.n2103 19.3944
R10196 gnd.n3339 gnd.n2103 19.3944
R10197 gnd.n3339 gnd.n2101 19.3944
R10198 gnd.n3343 gnd.n2101 19.3944
R10199 gnd.n3343 gnd.n2097 19.3944
R10200 gnd.n3349 gnd.n2097 19.3944
R10201 gnd.n3349 gnd.n2095 19.3944
R10202 gnd.n3353 gnd.n2095 19.3944
R10203 gnd.n3353 gnd.n2091 19.3944
R10204 gnd.n3359 gnd.n2091 19.3944
R10205 gnd.n3359 gnd.n2089 19.3944
R10206 gnd.n3363 gnd.n2089 19.3944
R10207 gnd.n3363 gnd.n2085 19.3944
R10208 gnd.n3369 gnd.n2085 19.3944
R10209 gnd.n3369 gnd.n2083 19.3944
R10210 gnd.n3375 gnd.n2083 19.3944
R10211 gnd.n3375 gnd.n3374 19.3944
R10212 gnd.n5578 gnd.n5453 19.3944
R10213 gnd.n5578 gnd.n5454 19.3944
R10214 gnd.n5574 gnd.n5454 19.3944
R10215 gnd.n5574 gnd.n5573 19.3944
R10216 gnd.n5573 gnd.n5572 19.3944
R10217 gnd.n5572 gnd.n5460 19.3944
R10218 gnd.n5568 gnd.n5460 19.3944
R10219 gnd.n5568 gnd.n5567 19.3944
R10220 gnd.n5567 gnd.n5566 19.3944
R10221 gnd.n5566 gnd.n5465 19.3944
R10222 gnd.n5562 gnd.n5465 19.3944
R10223 gnd.n5562 gnd.n5561 19.3944
R10224 gnd.n5561 gnd.n1456 19.3944
R10225 gnd.n6024 gnd.n1456 19.3944
R10226 gnd.n6024 gnd.n1454 19.3944
R10227 gnd.n6028 gnd.n1454 19.3944
R10228 gnd.n6028 gnd.n1425 19.3944
R10229 gnd.n6083 gnd.n1425 19.3944
R10230 gnd.n6083 gnd.n1423 19.3944
R10231 gnd.n6087 gnd.n1423 19.3944
R10232 gnd.n6087 gnd.n1397 19.3944
R10233 gnd.n6133 gnd.n1397 19.3944
R10234 gnd.n6133 gnd.n1395 19.3944
R10235 gnd.n6137 gnd.n1395 19.3944
R10236 gnd.n6137 gnd.n1370 19.3944
R10237 gnd.n6178 gnd.n1370 19.3944
R10238 gnd.n6178 gnd.n1368 19.3944
R10239 gnd.n6182 gnd.n1368 19.3944
R10240 gnd.n6182 gnd.n1339 19.3944
R10241 gnd.n6229 gnd.n1339 19.3944
R10242 gnd.n6229 gnd.n1337 19.3944
R10243 gnd.n6233 gnd.n1337 19.3944
R10244 gnd.n6233 gnd.n1306 19.3944
R10245 gnd.n6274 gnd.n1306 19.3944
R10246 gnd.n6274 gnd.n1303 19.3944
R10247 gnd.n6285 gnd.n1303 19.3944
R10248 gnd.n6285 gnd.n1304 19.3944
R10249 gnd.n6281 gnd.n1304 19.3944
R10250 gnd.n6281 gnd.n6280 19.3944
R10251 gnd.n6280 gnd.n1260 19.3944
R10252 gnd.n6393 gnd.n1260 19.3944
R10253 gnd.n6393 gnd.n1257 19.3944
R10254 gnd.n6398 gnd.n1257 19.3944
R10255 gnd.n6398 gnd.n1258 19.3944
R10256 gnd.n1258 gnd.n1229 19.3944
R10257 gnd.n6429 gnd.n1229 19.3944
R10258 gnd.n6429 gnd.n1226 19.3944
R10259 gnd.n6434 gnd.n1226 19.3944
R10260 gnd.n6434 gnd.n1227 19.3944
R10261 gnd.n1227 gnd.n1204 19.3944
R10262 gnd.n6458 gnd.n1204 19.3944
R10263 gnd.n6458 gnd.n1202 19.3944
R10264 gnd.n6462 gnd.n1202 19.3944
R10265 gnd.n6462 gnd.n1174 19.3944
R10266 gnd.n6515 gnd.n1174 19.3944
R10267 gnd.n6515 gnd.n1171 19.3944
R10268 gnd.n6520 gnd.n1171 19.3944
R10269 gnd.n6520 gnd.n1172 19.3944
R10270 gnd.n1172 gnd.n1139 19.3944
R10271 gnd.n6581 gnd.n1139 19.3944
R10272 gnd.n6581 gnd.n1136 19.3944
R10273 gnd.n6598 gnd.n1136 19.3944
R10274 gnd.n6598 gnd.n1137 19.3944
R10275 gnd.n6594 gnd.n1137 19.3944
R10276 gnd.n6594 gnd.n6593 19.3944
R10277 gnd.n6593 gnd.n6592 19.3944
R10278 gnd.n6592 gnd.n6589 19.3944
R10279 gnd.n6589 gnd.n1083 19.3944
R10280 gnd.n6704 gnd.n1083 19.3944
R10281 gnd.n6704 gnd.n1080 19.3944
R10282 gnd.n6709 gnd.n1080 19.3944
R10283 gnd.n6709 gnd.n1081 19.3944
R10284 gnd.n1081 gnd.n1053 19.3944
R10285 gnd.n6749 gnd.n1053 19.3944
R10286 gnd.n6749 gnd.n1050 19.3944
R10287 gnd.n6754 gnd.n1050 19.3944
R10288 gnd.n6754 gnd.n1051 19.3944
R10289 gnd.n1051 gnd.n1032 19.3944
R10290 gnd.n6801 gnd.n1032 19.3944
R10291 gnd.n6801 gnd.n1033 19.3944
R10292 gnd.n6797 gnd.n1033 19.3944
R10293 gnd.n6797 gnd.n1004 19.3944
R10294 gnd.n6842 gnd.n1004 19.3944
R10295 gnd.n6842 gnd.n1005 19.3944
R10296 gnd.n6838 gnd.n1005 19.3944
R10297 gnd.n6838 gnd.n732 19.3944
R10298 gnd.n7006 gnd.n732 19.3944
R10299 gnd.n7006 gnd.n729 19.3944
R10300 gnd.n7011 gnd.n729 19.3944
R10301 gnd.n7011 gnd.n730 19.3944
R10302 gnd.n730 gnd.n706 19.3944
R10303 gnd.n7036 gnd.n706 19.3944
R10304 gnd.n7036 gnd.n703 19.3944
R10305 gnd.n7041 gnd.n703 19.3944
R10306 gnd.n7041 gnd.n704 19.3944
R10307 gnd.n704 gnd.n682 19.3944
R10308 gnd.n7072 gnd.n682 19.3944
R10309 gnd.n7072 gnd.n680 19.3944
R10310 gnd.n7076 gnd.n680 19.3944
R10311 gnd.n7076 gnd.n588 19.3944
R10312 gnd.n7183 gnd.n588 19.3944
R10313 gnd.n7180 gnd.n7179 19.3944
R10314 gnd.n7179 gnd.n7178 19.3944
R10315 gnd.n7178 gnd.n593 19.3944
R10316 gnd.n7174 gnd.n593 19.3944
R10317 gnd.n7174 gnd.n7173 19.3944
R10318 gnd.n7173 gnd.n7172 19.3944
R10319 gnd.n7172 gnd.n598 19.3944
R10320 gnd.n7167 gnd.n598 19.3944
R10321 gnd.n7167 gnd.n7166 19.3944
R10322 gnd.n7166 gnd.n603 19.3944
R10323 gnd.n7159 gnd.n603 19.3944
R10324 gnd.n7159 gnd.n7158 19.3944
R10325 gnd.n7158 gnd.n613 19.3944
R10326 gnd.n7151 gnd.n613 19.3944
R10327 gnd.n7151 gnd.n7150 19.3944
R10328 gnd.n7150 gnd.n623 19.3944
R10329 gnd.n7143 gnd.n623 19.3944
R10330 gnd.n7143 gnd.n7142 19.3944
R10331 gnd.n7142 gnd.n631 19.3944
R10332 gnd.n7135 gnd.n631 19.3944
R10333 gnd.n7135 gnd.n7134 19.3944
R10334 gnd.n7134 gnd.n641 19.3944
R10335 gnd.n7127 gnd.n641 19.3944
R10336 gnd.n7127 gnd.n7126 19.3944
R10337 gnd.n7197 gnd.n7196 19.3944
R10338 gnd.n7196 gnd.n7191 19.3944
R10339 gnd.n7191 gnd.n7190 19.3944
R10340 gnd.n4161 gnd.t32 18.8012
R10341 gnd.n4146 gnd.t49 18.8012
R10342 gnd.n7703 gnd.n171 18.8012
R10343 gnd.n4005 gnd.n4004 18.4825
R10344 gnd.n959 gnd.n787 18.4247
R10345 gnd.n5929 gnd.n1590 18.4247
R10346 gnd.n7200 gnd.n571 18.2308
R10347 gnd.n5677 gnd.n5666 18.2308
R10348 gnd.n7536 gnd.n7535 18.2308
R10349 gnd.n4935 gnd.n4895 18.2308
R10350 gnd.t364 gnd.n3685 18.1639
R10351 gnd.n3713 gnd.t23 17.5266
R10352 gnd.n1963 gnd.t226 17.5266
R10353 gnd.n7697 gnd.t243 17.5266
R10354 gnd.n4112 gnd.t41 16.8893
R10355 gnd.n1926 gnd.t241 16.8893
R10356 gnd.n7721 gnd.t211 16.8893
R10357 gnd.n942 gnd.n939 16.6793
R10358 gnd.n7608 gnd.n7607 16.6793
R10359 gnd.n5015 gnd.n5012 16.6793
R10360 gnd.n5911 gnd.n5910 16.6793
R10361 gnd.n3940 gnd.t185 16.2519
R10362 gnd.n3640 gnd.t21 16.2519
R10363 gnd.n5226 gnd.t193 16.2519
R10364 gnd.n5293 gnd.t205 16.2519
R10365 gnd.n7402 gnd.t261 16.2519
R10366 gnd.n7745 gnd.t215 16.2519
R10367 gnd.n5449 gnd.n5448 15.9333
R10368 gnd.n5581 gnd.n5449 15.9333
R10369 gnd.n5581 gnd.n5580 15.9333
R10370 gnd.n5580 gnd.n5451 15.9333
R10371 gnd.n5500 gnd.n5499 15.9333
R10372 gnd.n5511 gnd.n5499 15.9333
R10373 gnd.n5513 gnd.n5511 15.9333
R10374 gnd.n5513 gnd.n5512 15.9333
R10375 gnd.n5512 gnd.n5489 15.9333
R10376 gnd.n5522 gnd.n5489 15.9333
R10377 gnd.n5522 gnd.n5521 15.9333
R10378 gnd.n5521 gnd.n5492 15.9333
R10379 gnd.n5492 gnd.n5490 15.9333
R10380 gnd.n5532 gnd.n5530 15.9333
R10381 gnd.n5532 gnd.n5531 15.9333
R10382 gnd.n5531 gnd.n5476 15.9333
R10383 gnd.n5543 gnd.n5476 15.9333
R10384 gnd.n5543 gnd.n5542 15.9333
R10385 gnd.n5542 gnd.n5477 15.9333
R10386 gnd.n5477 gnd.n5468 15.9333
R10387 gnd.n5558 gnd.n5468 15.9333
R10388 gnd.n6012 gnd.n1465 15.9333
R10389 gnd.n6020 gnd.n1441 15.9333
R10390 gnd.n6072 gnd.n1436 15.9333
R10391 gnd.n6081 gnd.n6080 15.9333
R10392 gnd.n6131 gnd.n6130 15.9333
R10393 gnd.n6139 gnd.n1379 15.9333
R10394 gnd.n6176 gnd.n1372 15.9333
R10395 gnd.n6185 gnd.n6184 15.9333
R10396 gnd.n6236 gnd.n6235 15.9333
R10397 gnd.n6272 gnd.n1308 15.9333
R10398 gnd.n6244 gnd.n1316 15.9333
R10399 gnd.n6256 gnd.n6255 15.9333
R10400 gnd.n6382 gnd.n1270 15.9333
R10401 gnd.n6391 gnd.n6390 15.9333
R10402 gnd.n6401 gnd.n6400 15.9333
R10403 gnd.n6352 gnd.n1238 15.9333
R10404 gnd.n6344 gnd.n1234 15.9333
R10405 gnd.n6446 gnd.n6445 15.9333
R10406 gnd.n6455 gnd.n6454 15.9333
R10407 gnd.n6454 gnd.n1196 15.9333
R10408 gnd.n6480 gnd.n1191 15.9333
R10409 gnd.n6505 gnd.n6504 15.9333
R10410 gnd.n6323 gnd.n1165 15.9333
R10411 gnd.n6495 gnd.n1160 15.9333
R10412 gnd.n6579 gnd.n1141 15.9333
R10413 gnd.n6601 gnd.n6600 15.9333
R10414 gnd.n6616 gnd.n1125 15.9333
R10415 gnd.n6610 gnd.n1112 15.9333
R10416 gnd.n6693 gnd.n1093 15.9333
R10417 gnd.n6702 gnd.n6701 15.9333
R10418 gnd.n6739 gnd.n6738 15.9333
R10419 gnd.n6672 gnd.n1044 15.9333
R10420 gnd.n6731 gnd.n1039 15.9333
R10421 gnd.n6804 gnd.n6803 15.9333
R10422 gnd.n6878 gnd.n724 15.9333
R10423 gnd.n7013 gnd.n724 15.9333
R10424 gnd.n7023 gnd.n717 15.9333
R10425 gnd.n7023 gnd.n7022 15.9333
R10426 gnd.n7022 gnd.n708 15.9333
R10427 gnd.n7034 gnd.n708 15.9333
R10428 gnd.n7034 gnd.n7033 15.9333
R10429 gnd.n7033 gnd.n710 15.9333
R10430 gnd.n710 gnd.n699 15.9333
R10431 gnd.n7043 gnd.n699 15.9333
R10432 gnd.n700 gnd.n692 15.9333
R10433 gnd.n7058 gnd.n692 15.9333
R10434 gnd.n7058 gnd.n7057 15.9333
R10435 gnd.n7057 gnd.n684 15.9333
R10436 gnd.n7070 gnd.n684 15.9333
R10437 gnd.n7070 gnd.n7069 15.9333
R10438 gnd.n7069 gnd.n686 15.9333
R10439 gnd.n686 gnd.n677 15.9333
R10440 gnd.n7078 gnd.n677 15.9333
R10441 gnd.n7080 gnd.n7079 15.9333
R10442 gnd.n7079 gnd.n584 15.9333
R10443 gnd.n7185 gnd.n584 15.9333
R10444 gnd.n7185 gnd.n585 15.9333
R10445 gnd.n4627 gnd.n4625 15.6674
R10446 gnd.n4595 gnd.n4593 15.6674
R10447 gnd.n4563 gnd.n4561 15.6674
R10448 gnd.n4532 gnd.n4530 15.6674
R10449 gnd.n4500 gnd.n4498 15.6674
R10450 gnd.n4468 gnd.n4466 15.6674
R10451 gnd.n4436 gnd.n4434 15.6674
R10452 gnd.n4405 gnd.n4403 15.6674
R10453 gnd.n3931 gnd.t185 15.6146
R10454 gnd.t169 gnd.n2073 15.6146
R10455 gnd.t144 gnd.n3379 15.6146
R10456 gnd.n5237 gnd.t193 15.6146
R10457 gnd.n5270 gnd.t205 15.6146
R10458 gnd.n7411 gnd.t261 15.6146
R10459 gnd.n7472 gnd.t215 15.6146
R10460 gnd.n899 gnd.n894 15.3217
R10461 gnd.n7568 gnd.n314 15.3217
R10462 gnd.n4973 gnd.n1990 15.3217
R10463 gnd.n5871 gnd.n1645 15.3217
R10464 gnd.n6836 gnd.t103 15.296
R10465 gnd.n745 gnd.n744 15.0827
R10466 gnd.n1479 gnd.n1474 15.0481
R10467 gnd.n755 gnd.n754 15.0481
R10468 gnd.n4299 gnd.t22 14.9773
R10469 gnd.n5172 gnd.t241 14.9773
R10470 gnd.n5343 gnd.t267 14.9773
R10471 gnd.t209 gnd.n1736 14.9773
R10472 gnd.n6089 gnd.t0 14.9773
R10473 gnd.n6795 gnd.t65 14.9773
R10474 gnd.n7261 gnd.t218 14.9773
R10475 gnd.n7344 gnd.t199 14.9773
R10476 gnd.t211 gnd.n136 14.9773
R10477 gnd.n6046 gnd.n1429 14.6587
R10478 gnd.n1387 gnd.t9 14.6587
R10479 gnd.n6208 gnd.n1333 14.6587
R10480 gnd.n1102 gnd.n1087 14.6587
R10481 gnd.t56 gnd.n1058 14.6587
R10482 gnd.n6823 gnd.n999 14.6587
R10483 gnd.n7004 gnd.n734 14.6587
R10484 gnd.t372 gnd.n3421 14.34
R10485 gnd.n4377 gnd.t363 14.34
R10486 gnd.n5126 gnd.t226 14.34
R10487 gnd.n5325 gnd.t267 14.34
R10488 gnd.n5415 gnd.t209 14.34
R10489 gnd.t218 gnd.n7260 14.34
R10490 gnd.n7318 gnd.t199 14.34
R10491 gnd.t243 gnd.n174 14.34
R10492 gnd.n6095 gnd.n1399 14.0214
R10493 gnd.t10 gnd.n1366 14.0214
R10494 gnd.n6371 gnd.n6370 14.0214
R10495 gnd.n6420 gnd.n6419 14.0214
R10496 gnd.n6322 gnd.n6315 14.0214
R10497 gnd.n6571 gnd.n6570 14.0214
R10498 gnd.n6740 gnd.t31 14.0214
R10499 gnd.n6775 gnd.n1029 14.0214
R10500 gnd.n6859 gnd.t72 14.0214
R10501 gnd.n4087 gnd.t365 13.7027
R10502 gnd.n3797 gnd.n3796 13.5763
R10503 gnd.n4741 gnd.n2030 13.5763
R10504 gnd.n4005 gnd.n3743 13.384
R10505 gnd.n6022 gnd.t75 13.384
R10506 gnd.n6113 gnd.n1409 13.384
R10507 gnd.n6194 gnd.n1358 13.384
R10508 gnd.n6217 gnd.t13 13.384
R10509 gnd.n1323 gnd.n1277 13.384
R10510 gnd.n6427 gnd.n6426 13.384
R10511 gnd.n6513 gnd.n1176 13.384
R10512 gnd.n6617 gnd.n1122 13.384
R10513 gnd.n6640 gnd.t54 13.384
R10514 gnd.n6720 gnd.n1071 13.384
R10515 gnd.n6813 gnd.n1020 13.384
R10516 gnd.n1490 gnd.n1471 13.1884
R10517 gnd.n1485 gnd.n1484 13.1884
R10518 gnd.n1484 gnd.n1483 13.1884
R10519 gnd.n748 gnd.n743 13.1884
R10520 gnd.n749 gnd.n748 13.1884
R10521 gnd.n1486 gnd.n1473 13.146
R10522 gnd.n1482 gnd.n1473 13.146
R10523 gnd.n747 gnd.n746 13.146
R10524 gnd.n747 gnd.n742 13.146
R10525 gnd.n7514 gnd.n171 13.0654
R10526 gnd.n4628 gnd.n4624 12.8005
R10527 gnd.n4596 gnd.n4592 12.8005
R10528 gnd.n4564 gnd.n4560 12.8005
R10529 gnd.n4533 gnd.n4529 12.8005
R10530 gnd.n4501 gnd.n4497 12.8005
R10531 gnd.n4469 gnd.n4465 12.8005
R10532 gnd.n4437 gnd.n4433 12.8005
R10533 gnd.n4406 gnd.n4402 12.8005
R10534 gnd.n6010 gnd.n1468 12.7467
R10535 gnd.t100 gnd.t107 12.7467
R10536 gnd.n6090 gnd.n1420 12.7467
R10537 gnd.t369 gnd.n1393 12.7467
R10538 gnd.n6226 gnd.n1343 12.7467
R10539 gnd.n6259 gnd.n1322 12.7467
R10540 gnd.n6345 gnd.n1222 12.7467
R10541 gnd.n6506 gnd.n1182 12.7467
R10542 gnd.n1124 gnd.n1116 12.7467
R10543 gnd.n6713 gnd.n6712 12.7467
R10544 gnd.n6768 gnd.t29 12.7467
R10545 gnd.n6794 gnd.n1014 12.7467
R10546 gnd.n6785 gnd.t132 12.7467
R10547 gnd.n5530 gnd.t47 12.4281
R10548 gnd.n7043 gnd.t355 12.4281
R10549 gnd.n3796 gnd.n3791 12.4126
R10550 gnd.n4744 gnd.n4741 12.4126
R10551 gnd.n6006 gnd.n6005 12.1761
R10552 gnd.n6999 gnd.n6998 12.1761
R10553 gnd.n1415 gnd.n1401 12.1094
R10554 gnd.n6152 gnd.n1364 12.1094
R10555 gnd.n6381 gnd.n1272 12.1094
R10556 gnd.n6353 gnd.n1247 12.1094
R10557 gnd.n6523 gnd.n6522 12.1094
R10558 gnd.n6560 gnd.n1132 12.1094
R10559 gnd.n6747 gnd.n1055 12.1094
R10560 gnd.n6657 gnd.n1027 12.1094
R10561 gnd.n4632 gnd.n4631 12.0247
R10562 gnd.n4600 gnd.n4599 12.0247
R10563 gnd.n4568 gnd.n4567 12.0247
R10564 gnd.n4537 gnd.n4536 12.0247
R10565 gnd.n4505 gnd.n4504 12.0247
R10566 gnd.n4473 gnd.n4472 12.0247
R10567 gnd.n4441 gnd.n4440 12.0247
R10568 gnd.n4410 gnd.n4409 12.0247
R10569 gnd.n6061 gnd.n1442 11.4721
R10570 gnd.n1349 gnd.n1335 11.4721
R10571 gnd.n6246 gnd.n6245 11.4721
R10572 gnd.n6444 gnd.n1217 11.4721
R10573 gnd.n6472 gnd.n6471 11.4721
R10574 gnd.n6631 gnd.n6630 11.4721
R10575 gnd.n1108 gnd.n1085 11.4721
R10576 gnd.n6784 gnd.n1001 11.4721
R10577 gnd.n6871 gnd.n987 11.4721
R10578 gnd.n4635 gnd.n4622 11.249
R10579 gnd.n4603 gnd.n4590 11.249
R10580 gnd.n4571 gnd.n4558 11.249
R10581 gnd.n4540 gnd.n4527 11.249
R10582 gnd.n4508 gnd.n4495 11.249
R10583 gnd.n4476 gnd.n4463 11.249
R10584 gnd.n4444 gnd.n4431 11.249
R10585 gnd.n4413 gnd.n4400 11.249
R10586 gnd.n4075 gnd.t365 11.1535
R10587 gnd.n6161 gnd.n6160 10.8348
R10588 gnd.n6265 gnd.t28 10.8348
R10589 gnd.n1264 gnd.n1251 10.8348
R10590 gnd.n6402 gnd.n1251 10.8348
R10591 gnd.n6538 gnd.n1156 10.8348
R10592 gnd.n6538 gnd.n6537 10.8348
R10593 gnd.n6609 gnd.t12 10.8348
R10594 gnd.n6756 gnd.n1047 10.8348
R10595 gnd.n902 gnd.n899 10.6672
R10596 gnd.n7573 gnd.n314 10.6672
R10597 gnd.n4975 gnd.n4973 10.6672
R10598 gnd.n5876 gnd.n1645 10.6672
R10599 gnd.n6934 gnd.n786 10.6151
R10600 gnd.n6934 gnd.n6933 10.6151
R10601 gnd.n6931 gnd.n964 10.6151
R10602 gnd.n6926 gnd.n964 10.6151
R10603 gnd.n6926 gnd.n6925 10.6151
R10604 gnd.n6925 gnd.n6924 10.6151
R10605 gnd.n6924 gnd.n967 10.6151
R10606 gnd.n6919 gnd.n967 10.6151
R10607 gnd.n6919 gnd.n6918 10.6151
R10608 gnd.n6918 gnd.n6917 10.6151
R10609 gnd.n6917 gnd.n970 10.6151
R10610 gnd.n6912 gnd.n970 10.6151
R10611 gnd.n6912 gnd.n6911 10.6151
R10612 gnd.n6911 gnd.n6910 10.6151
R10613 gnd.n6910 gnd.n973 10.6151
R10614 gnd.n6905 gnd.n973 10.6151
R10615 gnd.n6905 gnd.n6904 10.6151
R10616 gnd.n6904 gnd.n6903 10.6151
R10617 gnd.n6903 gnd.n976 10.6151
R10618 gnd.n6898 gnd.n976 10.6151
R10619 gnd.n6898 gnd.n6897 10.6151
R10620 gnd.n6897 gnd.n6896 10.6151
R10621 gnd.n6896 gnd.n979 10.6151
R10622 gnd.n6891 gnd.n979 10.6151
R10623 gnd.n6891 gnd.n6890 10.6151
R10624 gnd.n6890 gnd.n6889 10.6151
R10625 gnd.n6889 gnd.n982 10.6151
R10626 gnd.n6884 gnd.n982 10.6151
R10627 gnd.n6884 gnd.n6883 10.6151
R10628 gnd.n6883 gnd.n6882 10.6151
R10629 gnd.n5997 gnd.n5996 10.6151
R10630 gnd.n5996 gnd.n1439 10.6151
R10631 gnd.n6063 gnd.n1439 10.6151
R10632 gnd.n6064 gnd.n6063 10.6151
R10633 gnd.n6070 gnd.n6064 10.6151
R10634 gnd.n6070 gnd.n6069 10.6151
R10635 gnd.n6069 gnd.n6068 10.6151
R10636 gnd.n6068 gnd.n6065 10.6151
R10637 gnd.n6065 gnd.n1418 10.6151
R10638 gnd.n6092 gnd.n1418 10.6151
R10639 gnd.n6093 gnd.n6092 10.6151
R10640 gnd.n6094 gnd.n6093 10.6151
R10641 gnd.n6099 gnd.n6094 10.6151
R10642 gnd.n6100 gnd.n6099 10.6151
R10643 gnd.n6102 gnd.n6100 10.6151
R10644 gnd.n6102 gnd.n6101 10.6151
R10645 gnd.n6101 gnd.n1382 10.6151
R10646 gnd.n6157 gnd.n1382 10.6151
R10647 gnd.n6157 gnd.n6156 10.6151
R10648 gnd.n6156 gnd.n6155 10.6151
R10649 gnd.n6155 gnd.n1383 10.6151
R10650 gnd.n1384 gnd.n1383 10.6151
R10651 gnd.n1384 gnd.n1356 10.6151
R10652 gnd.n6196 gnd.n1356 10.6151
R10653 gnd.n6197 gnd.n6196 10.6151
R10654 gnd.n6205 gnd.n6197 10.6151
R10655 gnd.n6205 gnd.n6204 10.6151
R10656 gnd.n6204 gnd.n6203 10.6151
R10657 gnd.n6203 gnd.n6201 10.6151
R10658 gnd.n6201 gnd.n6200 10.6151
R10659 gnd.n6200 gnd.n6198 10.6151
R10660 gnd.n6198 gnd.n1319 10.6151
R10661 gnd.n6263 gnd.n1319 10.6151
R10662 gnd.n6263 gnd.n6262 10.6151
R10663 gnd.n6262 gnd.n6261 10.6151
R10664 gnd.n6261 gnd.n1320 10.6151
R10665 gnd.n1320 gnd.n1279 10.6151
R10666 gnd.n6368 gnd.n1279 10.6151
R10667 gnd.n6368 gnd.n6367 10.6151
R10668 gnd.n6367 gnd.n6366 10.6151
R10669 gnd.n6366 gnd.n1280 10.6151
R10670 gnd.n6360 gnd.n1280 10.6151
R10671 gnd.n6360 gnd.n6359 10.6151
R10672 gnd.n6359 gnd.n6358 10.6151
R10673 gnd.n6358 gnd.n6356 10.6151
R10674 gnd.n6356 gnd.n6355 10.6151
R10675 gnd.n6355 gnd.n6351 10.6151
R10676 gnd.n6351 gnd.n6350 10.6151
R10677 gnd.n6350 gnd.n6348 10.6151
R10678 gnd.n6348 gnd.n6347 10.6151
R10679 gnd.n6347 gnd.n1287 10.6151
R10680 gnd.n1287 gnd.n1286 10.6151
R10681 gnd.n1286 gnd.n1284 10.6151
R10682 gnd.n1284 gnd.n1283 10.6151
R10683 gnd.n1283 gnd.n1281 10.6151
R10684 gnd.n1281 gnd.n1198 10.6151
R10685 gnd.n6469 gnd.n1198 10.6151
R10686 gnd.n6469 gnd.n6468 10.6151
R10687 gnd.n6468 gnd.n6467 10.6151
R10688 gnd.n6467 gnd.n1199 10.6151
R10689 gnd.n6317 gnd.n1199 10.6151
R10690 gnd.n6318 gnd.n6317 10.6151
R10691 gnd.n6320 gnd.n6318 10.6151
R10692 gnd.n6320 gnd.n6319 10.6151
R10693 gnd.n6319 gnd.n1158 10.6151
R10694 gnd.n6532 gnd.n1158 10.6151
R10695 gnd.n6533 gnd.n6532 10.6151
R10696 gnd.n6535 gnd.n6533 10.6151
R10697 gnd.n6535 gnd.n6534 10.6151
R10698 gnd.n6534 gnd.n1149 10.6151
R10699 gnd.n6564 gnd.n1149 10.6151
R10700 gnd.n6565 gnd.n6564 10.6151
R10701 gnd.n6567 gnd.n6565 10.6151
R10702 gnd.n6567 gnd.n6566 10.6151
R10703 gnd.n6566 gnd.n1114 10.6151
R10704 gnd.n6626 gnd.n1114 10.6151
R10705 gnd.n6627 gnd.n6626 10.6151
R10706 gnd.n6628 gnd.n6627 10.6151
R10707 gnd.n6628 gnd.n1097 10.6151
R10708 gnd.n6691 gnd.n1097 10.6151
R10709 gnd.n6691 gnd.n6690 10.6151
R10710 gnd.n6690 gnd.n6689 10.6151
R10711 gnd.n6689 gnd.n6686 10.6151
R10712 gnd.n6686 gnd.n6685 10.6151
R10713 gnd.n6685 gnd.n6684 10.6151
R10714 gnd.n6684 gnd.n6683 10.6151
R10715 gnd.n6683 gnd.n6682 10.6151
R10716 gnd.n6682 gnd.n6679 10.6151
R10717 gnd.n6679 gnd.n6678 10.6151
R10718 gnd.n6678 gnd.n6676 10.6151
R10719 gnd.n6676 gnd.n6675 10.6151
R10720 gnd.n6675 gnd.n1098 10.6151
R10721 gnd.n1098 gnd.n1037 10.6151
R10722 gnd.n6770 gnd.n1037 10.6151
R10723 gnd.n6771 gnd.n6770 10.6151
R10724 gnd.n6772 gnd.n6771 10.6151
R10725 gnd.n6772 gnd.n1035 10.6151
R10726 gnd.n6778 gnd.n1035 10.6151
R10727 gnd.n6779 gnd.n6778 10.6151
R10728 gnd.n6792 gnd.n6779 10.6151
R10729 gnd.n6792 gnd.n6791 10.6151
R10730 gnd.n6791 gnd.n6790 10.6151
R10731 gnd.n6790 gnd.n6780 10.6151
R10732 gnd.n6783 gnd.n6780 10.6151
R10733 gnd.n6783 gnd.n6782 10.6151
R10734 gnd.n6782 gnd.n6781 10.6151
R10735 gnd.n6781 gnd.n985 10.6151
R10736 gnd.n6874 gnd.n985 10.6151
R10737 gnd.n6875 gnd.n6874 10.6151
R10738 gnd.n6876 gnd.n6875 10.6151
R10739 gnd.n5935 gnd.n5934 10.6151
R10740 gnd.n5938 gnd.n5935 10.6151
R10741 gnd.n5943 gnd.n5940 10.6151
R10742 gnd.n5944 gnd.n5943 10.6151
R10743 gnd.n5947 gnd.n5944 10.6151
R10744 gnd.n5948 gnd.n5947 10.6151
R10745 gnd.n5951 gnd.n5948 10.6151
R10746 gnd.n5952 gnd.n5951 10.6151
R10747 gnd.n5955 gnd.n5952 10.6151
R10748 gnd.n5956 gnd.n5955 10.6151
R10749 gnd.n5959 gnd.n5956 10.6151
R10750 gnd.n5960 gnd.n5959 10.6151
R10751 gnd.n5963 gnd.n5960 10.6151
R10752 gnd.n5964 gnd.n5963 10.6151
R10753 gnd.n5967 gnd.n5964 10.6151
R10754 gnd.n5968 gnd.n5967 10.6151
R10755 gnd.n5971 gnd.n5968 10.6151
R10756 gnd.n5972 gnd.n5971 10.6151
R10757 gnd.n5975 gnd.n5972 10.6151
R10758 gnd.n5976 gnd.n5975 10.6151
R10759 gnd.n5979 gnd.n5976 10.6151
R10760 gnd.n5980 gnd.n5979 10.6151
R10761 gnd.n5983 gnd.n5980 10.6151
R10762 gnd.n5984 gnd.n5983 10.6151
R10763 gnd.n5987 gnd.n5984 10.6151
R10764 gnd.n5988 gnd.n5987 10.6151
R10765 gnd.n5991 gnd.n5988 10.6151
R10766 gnd.n5993 gnd.n5991 10.6151
R10767 gnd.n5994 gnd.n5993 10.6151
R10768 gnd.n5998 gnd.n5994 10.6151
R10769 gnd.n6005 gnd.n6004 10.6151
R10770 gnd.n6004 gnd.n1491 10.6151
R10771 gnd.n1532 gnd.n1491 10.6151
R10772 gnd.n1533 gnd.n1532 10.6151
R10773 gnd.n1536 gnd.n1533 10.6151
R10774 gnd.n1537 gnd.n1536 10.6151
R10775 gnd.n1540 gnd.n1537 10.6151
R10776 gnd.n1541 gnd.n1540 10.6151
R10777 gnd.n1544 gnd.n1541 10.6151
R10778 gnd.n1545 gnd.n1544 10.6151
R10779 gnd.n1548 gnd.n1545 10.6151
R10780 gnd.n1549 gnd.n1548 10.6151
R10781 gnd.n1552 gnd.n1549 10.6151
R10782 gnd.n1553 gnd.n1552 10.6151
R10783 gnd.n1556 gnd.n1553 10.6151
R10784 gnd.n1557 gnd.n1556 10.6151
R10785 gnd.n1560 gnd.n1557 10.6151
R10786 gnd.n1561 gnd.n1560 10.6151
R10787 gnd.n1564 gnd.n1561 10.6151
R10788 gnd.n1565 gnd.n1564 10.6151
R10789 gnd.n1568 gnd.n1565 10.6151
R10790 gnd.n1569 gnd.n1568 10.6151
R10791 gnd.n1572 gnd.n1569 10.6151
R10792 gnd.n1573 gnd.n1572 10.6151
R10793 gnd.n1576 gnd.n1573 10.6151
R10794 gnd.n1577 gnd.n1576 10.6151
R10795 gnd.n1580 gnd.n1577 10.6151
R10796 gnd.n1581 gnd.n1580 10.6151
R10797 gnd.n1585 gnd.n1584 10.6151
R10798 gnd.n1588 gnd.n1585 10.6151
R10799 gnd.n6998 gnd.n760 10.6151
R10800 gnd.n761 gnd.n760 10.6151
R10801 gnd.n6991 gnd.n761 10.6151
R10802 gnd.n6991 gnd.n6990 10.6151
R10803 gnd.n6990 gnd.n6989 10.6151
R10804 gnd.n6989 gnd.n763 10.6151
R10805 gnd.n6984 gnd.n763 10.6151
R10806 gnd.n6984 gnd.n6983 10.6151
R10807 gnd.n6983 gnd.n6982 10.6151
R10808 gnd.n6982 gnd.n766 10.6151
R10809 gnd.n6977 gnd.n766 10.6151
R10810 gnd.n6977 gnd.n6976 10.6151
R10811 gnd.n6976 gnd.n6975 10.6151
R10812 gnd.n6975 gnd.n769 10.6151
R10813 gnd.n6970 gnd.n769 10.6151
R10814 gnd.n6970 gnd.n6969 10.6151
R10815 gnd.n6969 gnd.n6968 10.6151
R10816 gnd.n6968 gnd.n772 10.6151
R10817 gnd.n6963 gnd.n772 10.6151
R10818 gnd.n6963 gnd.n6962 10.6151
R10819 gnd.n6962 gnd.n6961 10.6151
R10820 gnd.n6961 gnd.n775 10.6151
R10821 gnd.n6956 gnd.n775 10.6151
R10822 gnd.n6956 gnd.n6955 10.6151
R10823 gnd.n6955 gnd.n6954 10.6151
R10824 gnd.n6954 gnd.n778 10.6151
R10825 gnd.n6949 gnd.n778 10.6151
R10826 gnd.n6949 gnd.n6948 10.6151
R10827 gnd.n6946 gnd.n783 10.6151
R10828 gnd.n6941 gnd.n783 10.6151
R10829 gnd.n6008 gnd.n6007 10.6151
R10830 gnd.n6007 gnd.n1445 10.6151
R10831 gnd.n6059 gnd.n1445 10.6151
R10832 gnd.n6059 gnd.n6058 10.6151
R10833 gnd.n6058 gnd.n6057 10.6151
R10834 gnd.n6057 gnd.n6056 10.6151
R10835 gnd.n6056 gnd.n1446 10.6151
R10836 gnd.n6050 gnd.n1446 10.6151
R10837 gnd.n6050 gnd.n6049 10.6151
R10838 gnd.n6049 gnd.n1412 10.6151
R10839 gnd.n6111 gnd.n1412 10.6151
R10840 gnd.n6111 gnd.n6110 10.6151
R10841 gnd.n6110 gnd.n6109 10.6151
R10842 gnd.n6109 gnd.n1413 10.6151
R10843 gnd.n1414 gnd.n1413 10.6151
R10844 gnd.n1414 gnd.n1377 10.6151
R10845 gnd.n6163 gnd.n1377 10.6151
R10846 gnd.n6164 gnd.n6163 10.6151
R10847 gnd.n6173 gnd.n6164 10.6151
R10848 gnd.n6173 gnd.n6172 10.6151
R10849 gnd.n6172 gnd.n6171 10.6151
R10850 gnd.n6171 gnd.n6165 10.6151
R10851 gnd.n6166 gnd.n6165 10.6151
R10852 gnd.n6166 gnd.n1346 10.6151
R10853 gnd.n6224 gnd.n1346 10.6151
R10854 gnd.n6224 gnd.n6223 10.6151
R10855 gnd.n6223 gnd.n6222 10.6151
R10856 gnd.n6222 gnd.n1347 10.6151
R10857 gnd.n1348 gnd.n1347 10.6151
R10858 gnd.n1348 gnd.n1313 10.6151
R10859 gnd.n6269 gnd.n1313 10.6151
R10860 gnd.n6269 gnd.n6268 10.6151
R10861 gnd.n6268 gnd.n6267 10.6151
R10862 gnd.n6267 gnd.n1314 10.6151
R10863 gnd.n6257 gnd.n1314 10.6151
R10864 gnd.n6257 gnd.n1275 10.6151
R10865 gnd.n6374 gnd.n1275 10.6151
R10866 gnd.n6375 gnd.n6374 10.6151
R10867 gnd.n6379 gnd.n6375 10.6151
R10868 gnd.n6379 gnd.n6378 10.6151
R10869 gnd.n6378 gnd.n6377 10.6151
R10870 gnd.n6377 gnd.n1249 10.6151
R10871 gnd.n6404 gnd.n1249 10.6151
R10872 gnd.n6405 gnd.n6404 10.6151
R10873 gnd.n6406 gnd.n6405 10.6151
R10874 gnd.n6406 gnd.n1236 10.6151
R10875 gnd.n6422 gnd.n1236 10.6151
R10876 gnd.n6423 gnd.n6422 10.6151
R10877 gnd.n6424 gnd.n6423 10.6151
R10878 gnd.n6424 gnd.n1220 10.6151
R10879 gnd.n6439 gnd.n1220 10.6151
R10880 gnd.n6440 gnd.n6439 10.6151
R10881 gnd.n6442 gnd.n6440 10.6151
R10882 gnd.n6442 gnd.n6441 10.6151
R10883 gnd.n6441 gnd.n1194 10.6151
R10884 gnd.n6475 gnd.n1194 10.6151
R10885 gnd.n6476 gnd.n6475 10.6151
R10886 gnd.n6477 gnd.n6476 10.6151
R10887 gnd.n6477 gnd.n1180 10.6151
R10888 gnd.n6508 gnd.n1180 10.6151
R10889 gnd.n6509 gnd.n6508 10.6151
R10890 gnd.n6510 gnd.n6509 10.6151
R10891 gnd.n6510 gnd.n1163 10.6151
R10892 gnd.n6525 gnd.n1163 10.6151
R10893 gnd.n6526 gnd.n6525 10.6151
R10894 gnd.n6528 gnd.n6526 10.6151
R10895 gnd.n6528 gnd.n6527 10.6151
R10896 gnd.n6527 gnd.n1146 10.6151
R10897 gnd.n6576 gnd.n1146 10.6151
R10898 gnd.n6576 gnd.n6575 10.6151
R10899 gnd.n6575 gnd.n6574 10.6151
R10900 gnd.n6574 gnd.n1147 10.6151
R10901 gnd.n1147 gnd.n1120 10.6151
R10902 gnd.n6619 gnd.n1120 10.6151
R10903 gnd.n6620 gnd.n6619 10.6151
R10904 gnd.n6622 gnd.n6620 10.6151
R10905 gnd.n6622 gnd.n6621 10.6151
R10906 gnd.n6621 gnd.n1110 10.6151
R10907 gnd.n6634 gnd.n1110 10.6151
R10908 gnd.n6635 gnd.n6634 10.6151
R10909 gnd.n6637 gnd.n6635 10.6151
R10910 gnd.n6637 gnd.n6636 10.6151
R10911 gnd.n6636 gnd.n1073 10.6151
R10912 gnd.n6716 gnd.n1073 10.6151
R10913 gnd.n6717 gnd.n6716 10.6151
R10914 gnd.n6718 gnd.n6717 10.6151
R10915 gnd.n6718 gnd.n1060 10.6151
R10916 gnd.n6742 gnd.n1060 10.6151
R10917 gnd.n6743 gnd.n6742 10.6151
R10918 gnd.n6744 gnd.n6743 10.6151
R10919 gnd.n6744 gnd.n1042 10.6151
R10920 gnd.n6759 gnd.n1042 10.6151
R10921 gnd.n6760 gnd.n6759 10.6151
R10922 gnd.n6766 gnd.n6760 10.6151
R10923 gnd.n6766 gnd.n6765 10.6151
R10924 gnd.n6765 gnd.n6764 10.6151
R10925 gnd.n6764 gnd.n6761 10.6151
R10926 gnd.n6761 gnd.n1018 10.6151
R10927 gnd.n6815 gnd.n1018 10.6151
R10928 gnd.n6816 gnd.n6815 10.6151
R10929 gnd.n6820 gnd.n6816 10.6151
R10930 gnd.n6820 gnd.n6819 10.6151
R10931 gnd.n6819 gnd.n6818 10.6151
R10932 gnd.n6818 gnd.n990 10.6151
R10933 gnd.n6867 gnd.n990 10.6151
R10934 gnd.n6868 gnd.n6867 10.6151
R10935 gnd.n6869 gnd.n6868 10.6151
R10936 gnd.n6869 gnd.n740 10.6151
R10937 gnd.n7001 gnd.n740 10.6151
R10938 gnd.n7001 gnd.n7000 10.6151
R10939 gnd.n3994 gnd.t361 10.5161
R10940 gnd.n3423 gnd.t372 10.5161
R10941 gnd.n4360 gnd.t363 10.5161
R10942 gnd.n4636 gnd.n4620 10.4732
R10943 gnd.n4604 gnd.n4588 10.4732
R10944 gnd.n4572 gnd.n4556 10.4732
R10945 gnd.n4541 gnd.n4525 10.4732
R10946 gnd.n4509 gnd.n4493 10.4732
R10947 gnd.n4477 gnd.n4461 10.4732
R10948 gnd.n4445 gnd.n4429 10.4732
R10949 gnd.n4414 gnd.n4398 10.4732
R10950 gnd.n1452 gnd.n1442 10.1975
R10951 gnd.n6054 gnd.n6053 10.1975
R10952 gnd.n6218 gnd.n1349 10.1975
R10953 gnd.n1217 gnd.n1206 10.1975
R10954 gnd.n6473 gnd.n6472 10.1975
R10955 gnd.n6639 gnd.n1108 10.1975
R10956 gnd.n6786 gnd.n6784 10.1975
R10957 gnd.n6835 gnd.n987 10.1975
R10958 gnd.t22 gnd.n3440 9.87883
R10959 gnd.n4640 gnd.n4639 9.69747
R10960 gnd.n4608 gnd.n4607 9.69747
R10961 gnd.n4576 gnd.n4575 9.69747
R10962 gnd.n4545 gnd.n4544 9.69747
R10963 gnd.n4513 gnd.n4512 9.69747
R10964 gnd.n4481 gnd.n4480 9.69747
R10965 gnd.n4449 gnd.n4448 9.69747
R10966 gnd.n4418 gnd.n4417 9.69747
R10967 gnd.n6105 gnd.n1415 9.56018
R10968 gnd.n6153 gnd.n6152 9.56018
R10969 gnd.n6364 gnd.n1272 9.56018
R10970 gnd.n6363 gnd.t26 9.56018
R10971 gnd.n6408 gnd.n1247 9.56018
R10972 gnd.n6522 gnd.n1168 9.56018
R10973 gnd.n1150 gnd.t11 9.56018
R10974 gnd.n6561 gnd.n6560 9.56018
R10975 gnd.n6747 gnd.n6746 9.56018
R10976 gnd.n6657 gnd.n6656 9.56018
R10977 gnd.n4646 gnd.n4645 9.45567
R10978 gnd.n4614 gnd.n4613 9.45567
R10979 gnd.n4582 gnd.n4581 9.45567
R10980 gnd.n4551 gnd.n4550 9.45567
R10981 gnd.n4519 gnd.n4518 9.45567
R10982 gnd.n4487 gnd.n4486 9.45567
R10983 gnd.n4455 gnd.n4454 9.45567
R10984 gnd.n4424 gnd.n4423 9.45567
R10985 gnd.n939 gnd.n938 9.30959
R10986 gnd.n7607 gnd.n278 9.30959
R10987 gnd.n5012 gnd.n5011 9.30959
R10988 gnd.n5910 gnd.n1609 9.30959
R10989 gnd.n4645 gnd.n4644 9.3005
R10990 gnd.n4618 gnd.n4617 9.3005
R10991 gnd.n4639 gnd.n4638 9.3005
R10992 gnd.n4637 gnd.n4636 9.3005
R10993 gnd.n4622 gnd.n4621 9.3005
R10994 gnd.n4631 gnd.n4630 9.3005
R10995 gnd.n4629 gnd.n4628 9.3005
R10996 gnd.n4613 gnd.n4612 9.3005
R10997 gnd.n4586 gnd.n4585 9.3005
R10998 gnd.n4607 gnd.n4606 9.3005
R10999 gnd.n4605 gnd.n4604 9.3005
R11000 gnd.n4590 gnd.n4589 9.3005
R11001 gnd.n4599 gnd.n4598 9.3005
R11002 gnd.n4597 gnd.n4596 9.3005
R11003 gnd.n4581 gnd.n4580 9.3005
R11004 gnd.n4554 gnd.n4553 9.3005
R11005 gnd.n4575 gnd.n4574 9.3005
R11006 gnd.n4573 gnd.n4572 9.3005
R11007 gnd.n4558 gnd.n4557 9.3005
R11008 gnd.n4567 gnd.n4566 9.3005
R11009 gnd.n4565 gnd.n4564 9.3005
R11010 gnd.n4550 gnd.n4549 9.3005
R11011 gnd.n4523 gnd.n4522 9.3005
R11012 gnd.n4544 gnd.n4543 9.3005
R11013 gnd.n4542 gnd.n4541 9.3005
R11014 gnd.n4527 gnd.n4526 9.3005
R11015 gnd.n4536 gnd.n4535 9.3005
R11016 gnd.n4534 gnd.n4533 9.3005
R11017 gnd.n4518 gnd.n4517 9.3005
R11018 gnd.n4491 gnd.n4490 9.3005
R11019 gnd.n4512 gnd.n4511 9.3005
R11020 gnd.n4510 gnd.n4509 9.3005
R11021 gnd.n4495 gnd.n4494 9.3005
R11022 gnd.n4504 gnd.n4503 9.3005
R11023 gnd.n4502 gnd.n4501 9.3005
R11024 gnd.n4486 gnd.n4485 9.3005
R11025 gnd.n4459 gnd.n4458 9.3005
R11026 gnd.n4480 gnd.n4479 9.3005
R11027 gnd.n4478 gnd.n4477 9.3005
R11028 gnd.n4463 gnd.n4462 9.3005
R11029 gnd.n4472 gnd.n4471 9.3005
R11030 gnd.n4470 gnd.n4469 9.3005
R11031 gnd.n4454 gnd.n4453 9.3005
R11032 gnd.n4427 gnd.n4426 9.3005
R11033 gnd.n4448 gnd.n4447 9.3005
R11034 gnd.n4446 gnd.n4445 9.3005
R11035 gnd.n4431 gnd.n4430 9.3005
R11036 gnd.n4440 gnd.n4439 9.3005
R11037 gnd.n4438 gnd.n4437 9.3005
R11038 gnd.n4423 gnd.n4422 9.3005
R11039 gnd.n4396 gnd.n4395 9.3005
R11040 gnd.n4417 gnd.n4416 9.3005
R11041 gnd.n4415 gnd.n4414 9.3005
R11042 gnd.n4400 gnd.n4399 9.3005
R11043 gnd.n4409 gnd.n4408 9.3005
R11044 gnd.n4407 gnd.n4406 9.3005
R11045 gnd.n4771 gnd.n4770 9.3005
R11046 gnd.n4769 gnd.n2018 9.3005
R11047 gnd.n4768 gnd.n4767 9.3005
R11048 gnd.n4764 gnd.n2019 9.3005
R11049 gnd.n4761 gnd.n2020 9.3005
R11050 gnd.n4760 gnd.n2021 9.3005
R11051 gnd.n4757 gnd.n2022 9.3005
R11052 gnd.n4756 gnd.n2023 9.3005
R11053 gnd.n4753 gnd.n2024 9.3005
R11054 gnd.n4752 gnd.n2025 9.3005
R11055 gnd.n4749 gnd.n2026 9.3005
R11056 gnd.n4748 gnd.n2027 9.3005
R11057 gnd.n4745 gnd.n2028 9.3005
R11058 gnd.n4744 gnd.n2029 9.3005
R11059 gnd.n4741 gnd.n4740 9.3005
R11060 gnd.n4739 gnd.n2030 9.3005
R11061 gnd.n4772 gnd.n2017 9.3005
R11062 gnd.n4013 gnd.n4012 9.3005
R11063 gnd.n3717 gnd.n3716 9.3005
R11064 gnd.n4040 gnd.n4039 9.3005
R11065 gnd.n4041 gnd.n3715 9.3005
R11066 gnd.n4045 gnd.n4042 9.3005
R11067 gnd.n4044 gnd.n4043 9.3005
R11068 gnd.n3689 gnd.n3688 9.3005
R11069 gnd.n4070 gnd.n4069 9.3005
R11070 gnd.n4071 gnd.n3687 9.3005
R11071 gnd.n4073 gnd.n4072 9.3005
R11072 gnd.n3667 gnd.n3666 9.3005
R11073 gnd.n4101 gnd.n4100 9.3005
R11074 gnd.n4102 gnd.n3665 9.3005
R11075 gnd.n4110 gnd.n4103 9.3005
R11076 gnd.n4109 gnd.n4104 9.3005
R11077 gnd.n4108 gnd.n4106 9.3005
R11078 gnd.n4105 gnd.n3614 9.3005
R11079 gnd.n4158 gnd.n3615 9.3005
R11080 gnd.n4157 gnd.n3616 9.3005
R11081 gnd.n4156 gnd.n3617 9.3005
R11082 gnd.n3636 gnd.n3618 9.3005
R11083 gnd.n3638 gnd.n3637 9.3005
R11084 gnd.n3520 gnd.n3519 9.3005
R11085 gnd.n4196 gnd.n4195 9.3005
R11086 gnd.n4197 gnd.n3518 9.3005
R11087 gnd.n4201 gnd.n4198 9.3005
R11088 gnd.n4200 gnd.n4199 9.3005
R11089 gnd.n3493 gnd.n3492 9.3005
R11090 gnd.n4236 gnd.n4235 9.3005
R11091 gnd.n4237 gnd.n3491 9.3005
R11092 gnd.n4241 gnd.n4238 9.3005
R11093 gnd.n4240 gnd.n4239 9.3005
R11094 gnd.n3466 gnd.n3465 9.3005
R11095 gnd.n4281 gnd.n4280 9.3005
R11096 gnd.n4282 gnd.n3464 9.3005
R11097 gnd.n4286 gnd.n4283 9.3005
R11098 gnd.n4285 gnd.n4284 9.3005
R11099 gnd.n3438 gnd.n3437 9.3005
R11100 gnd.n4321 gnd.n4320 9.3005
R11101 gnd.n4322 gnd.n3436 9.3005
R11102 gnd.n4326 gnd.n4323 9.3005
R11103 gnd.n4325 gnd.n4324 9.3005
R11104 gnd.n3411 gnd.n3410 9.3005
R11105 gnd.n4370 gnd.n4369 9.3005
R11106 gnd.n4371 gnd.n3409 9.3005
R11107 gnd.n4375 gnd.n4372 9.3005
R11108 gnd.n4374 gnd.n4373 9.3005
R11109 gnd.n3384 gnd.n3383 9.3005
R11110 gnd.n4664 gnd.n4663 9.3005
R11111 gnd.n4665 gnd.n3382 9.3005
R11112 gnd.n4671 gnd.n4666 9.3005
R11113 gnd.n4670 gnd.n4667 9.3005
R11114 gnd.n4669 gnd.n4668 9.3005
R11115 gnd.n4014 gnd.n4011 9.3005
R11116 gnd.n3796 gnd.n3755 9.3005
R11117 gnd.n3791 gnd.n3790 9.3005
R11118 gnd.n3789 gnd.n3756 9.3005
R11119 gnd.n3788 gnd.n3787 9.3005
R11120 gnd.n3784 gnd.n3757 9.3005
R11121 gnd.n3781 gnd.n3780 9.3005
R11122 gnd.n3779 gnd.n3758 9.3005
R11123 gnd.n3778 gnd.n3777 9.3005
R11124 gnd.n3774 gnd.n3759 9.3005
R11125 gnd.n3771 gnd.n3770 9.3005
R11126 gnd.n3769 gnd.n3760 9.3005
R11127 gnd.n3768 gnd.n3767 9.3005
R11128 gnd.n3764 gnd.n3762 9.3005
R11129 gnd.n3761 gnd.n3741 9.3005
R11130 gnd.n4008 gnd.n3740 9.3005
R11131 gnd.n4010 gnd.n4009 9.3005
R11132 gnd.n3798 gnd.n3797 9.3005
R11133 gnd.n4021 gnd.n3727 9.3005
R11134 gnd.n4028 gnd.n3728 9.3005
R11135 gnd.n4030 gnd.n4029 9.3005
R11136 gnd.n4031 gnd.n3708 9.3005
R11137 gnd.n4050 gnd.n4049 9.3005
R11138 gnd.n4052 gnd.n3700 9.3005
R11139 gnd.n4059 gnd.n3702 9.3005
R11140 gnd.n4060 gnd.n3697 9.3005
R11141 gnd.n4062 gnd.n4061 9.3005
R11142 gnd.n3698 gnd.n3683 9.3005
R11143 gnd.n4078 gnd.n3681 9.3005
R11144 gnd.n4082 gnd.n4081 9.3005
R11145 gnd.n4080 gnd.n3657 9.3005
R11146 gnd.n4117 gnd.n3656 9.3005
R11147 gnd.n4120 gnd.n4119 9.3005
R11148 gnd.n3653 gnd.n3652 9.3005
R11149 gnd.n4126 gnd.n3654 9.3005
R11150 gnd.n4128 gnd.n4127 9.3005
R11151 gnd.n4130 gnd.n3651 9.3005
R11152 gnd.n4133 gnd.n4132 9.3005
R11153 gnd.n4136 gnd.n4134 9.3005
R11154 gnd.n4138 gnd.n4137 9.3005
R11155 gnd.n4144 gnd.n4139 9.3005
R11156 gnd.n4143 gnd.n4142 9.3005
R11157 gnd.n3511 gnd.n3510 9.3005
R11158 gnd.n4210 gnd.n4209 9.3005
R11159 gnd.n4211 gnd.n3504 9.3005
R11160 gnd.n4219 gnd.n3503 9.3005
R11161 gnd.n4222 gnd.n4221 9.3005
R11162 gnd.n4224 gnd.n4223 9.3005
R11163 gnd.n4227 gnd.n3486 9.3005
R11164 gnd.n4225 gnd.n3484 9.3005
R11165 gnd.n4247 gnd.n3482 9.3005
R11166 gnd.n4249 gnd.n4248 9.3005
R11167 gnd.n3456 gnd.n3455 9.3005
R11168 gnd.n4295 gnd.n4294 9.3005
R11169 gnd.n4296 gnd.n3449 9.3005
R11170 gnd.n4304 gnd.n3448 9.3005
R11171 gnd.n4307 gnd.n4306 9.3005
R11172 gnd.n4309 gnd.n4308 9.3005
R11173 gnd.n4312 gnd.n3431 9.3005
R11174 gnd.n4310 gnd.n3429 9.3005
R11175 gnd.n4332 gnd.n3427 9.3005
R11176 gnd.n4334 gnd.n4333 9.3005
R11177 gnd.n3402 gnd.n3401 9.3005
R11178 gnd.n4384 gnd.n4383 9.3005
R11179 gnd.n4385 gnd.n3395 9.3005
R11180 gnd.n4393 gnd.n3394 9.3005
R11181 gnd.n4652 gnd.n4651 9.3005
R11182 gnd.n4654 gnd.n4653 9.3005
R11183 gnd.n4655 gnd.n2070 9.3005
R11184 gnd.n4679 gnd.n4678 9.3005
R11185 gnd.n2071 gnd.n2033 9.3005
R11186 gnd.n4019 gnd.n4018 9.3005
R11187 gnd.n4735 gnd.n2034 9.3005
R11188 gnd.n4734 gnd.n2036 9.3005
R11189 gnd.n4731 gnd.n2037 9.3005
R11190 gnd.n4730 gnd.n2038 9.3005
R11191 gnd.n4727 gnd.n2039 9.3005
R11192 gnd.n4726 gnd.n2040 9.3005
R11193 gnd.n4723 gnd.n2041 9.3005
R11194 gnd.n4722 gnd.n2042 9.3005
R11195 gnd.n4719 gnd.n2043 9.3005
R11196 gnd.n4718 gnd.n2044 9.3005
R11197 gnd.n4715 gnd.n2045 9.3005
R11198 gnd.n4714 gnd.n2046 9.3005
R11199 gnd.n4711 gnd.n2047 9.3005
R11200 gnd.n4710 gnd.n2048 9.3005
R11201 gnd.n4707 gnd.n2049 9.3005
R11202 gnd.n4706 gnd.n2050 9.3005
R11203 gnd.n4703 gnd.n2051 9.3005
R11204 gnd.n4702 gnd.n2052 9.3005
R11205 gnd.n4699 gnd.n2053 9.3005
R11206 gnd.n4698 gnd.n2054 9.3005
R11207 gnd.n4695 gnd.n2055 9.3005
R11208 gnd.n4694 gnd.n2056 9.3005
R11209 gnd.n4691 gnd.n2060 9.3005
R11210 gnd.n4690 gnd.n2061 9.3005
R11211 gnd.n4687 gnd.n2062 9.3005
R11212 gnd.n4686 gnd.n2063 9.3005
R11213 gnd.n4737 gnd.n4736 9.3005
R11214 gnd.n4188 gnd.n4172 9.3005
R11215 gnd.n4187 gnd.n4173 9.3005
R11216 gnd.n4186 gnd.n4174 9.3005
R11217 gnd.n4184 gnd.n4175 9.3005
R11218 gnd.n4183 gnd.n4176 9.3005
R11219 gnd.n4181 gnd.n4177 9.3005
R11220 gnd.n4180 gnd.n4178 9.3005
R11221 gnd.n3474 gnd.n3473 9.3005
R11222 gnd.n4257 gnd.n4256 9.3005
R11223 gnd.n4258 gnd.n3472 9.3005
R11224 gnd.n4275 gnd.n4259 9.3005
R11225 gnd.n4274 gnd.n4260 9.3005
R11226 gnd.n4273 gnd.n4261 9.3005
R11227 gnd.n4271 gnd.n4262 9.3005
R11228 gnd.n4270 gnd.n4263 9.3005
R11229 gnd.n4268 gnd.n4264 9.3005
R11230 gnd.n4267 gnd.n4265 9.3005
R11231 gnd.n3418 gnd.n3417 9.3005
R11232 gnd.n4342 gnd.n4341 9.3005
R11233 gnd.n4343 gnd.n3416 9.3005
R11234 gnd.n4364 gnd.n4344 9.3005
R11235 gnd.n4363 gnd.n4345 9.3005
R11236 gnd.n4362 gnd.n4346 9.3005
R11237 gnd.n4359 gnd.n4347 9.3005
R11238 gnd.n4358 gnd.n4348 9.3005
R11239 gnd.n4356 gnd.n4349 9.3005
R11240 gnd.n4355 gnd.n4350 9.3005
R11241 gnd.n4353 gnd.n4352 9.3005
R11242 gnd.n4351 gnd.n2065 9.3005
R11243 gnd.n3929 gnd.n3928 9.3005
R11244 gnd.n3819 gnd.n3818 9.3005
R11245 gnd.n3943 gnd.n3942 9.3005
R11246 gnd.n3944 gnd.n3817 9.3005
R11247 gnd.n3946 gnd.n3945 9.3005
R11248 gnd.n3807 gnd.n3806 9.3005
R11249 gnd.n3959 gnd.n3958 9.3005
R11250 gnd.n3960 gnd.n3805 9.3005
R11251 gnd.n3992 gnd.n3961 9.3005
R11252 gnd.n3991 gnd.n3962 9.3005
R11253 gnd.n3990 gnd.n3963 9.3005
R11254 gnd.n3989 gnd.n3964 9.3005
R11255 gnd.n3986 gnd.n3965 9.3005
R11256 gnd.n3985 gnd.n3966 9.3005
R11257 gnd.n3984 gnd.n3967 9.3005
R11258 gnd.n3982 gnd.n3968 9.3005
R11259 gnd.n3981 gnd.n3969 9.3005
R11260 gnd.n3978 gnd.n3970 9.3005
R11261 gnd.n3977 gnd.n3971 9.3005
R11262 gnd.n3976 gnd.n3972 9.3005
R11263 gnd.n3974 gnd.n3973 9.3005
R11264 gnd.n3673 gnd.n3672 9.3005
R11265 gnd.n4090 gnd.n4089 9.3005
R11266 gnd.n4091 gnd.n3671 9.3005
R11267 gnd.n4095 gnd.n4092 9.3005
R11268 gnd.n4094 gnd.n4093 9.3005
R11269 gnd.n3595 gnd.n3594 9.3005
R11270 gnd.n4170 gnd.n4169 9.3005
R11271 gnd.n3927 gnd.n3828 9.3005
R11272 gnd.n3830 gnd.n3829 9.3005
R11273 gnd.n3874 gnd.n3872 9.3005
R11274 gnd.n3875 gnd.n3871 9.3005
R11275 gnd.n3878 gnd.n3867 9.3005
R11276 gnd.n3879 gnd.n3866 9.3005
R11277 gnd.n3882 gnd.n3865 9.3005
R11278 gnd.n3883 gnd.n3864 9.3005
R11279 gnd.n3886 gnd.n3863 9.3005
R11280 gnd.n3887 gnd.n3862 9.3005
R11281 gnd.n3890 gnd.n3861 9.3005
R11282 gnd.n3891 gnd.n3860 9.3005
R11283 gnd.n3894 gnd.n3859 9.3005
R11284 gnd.n3895 gnd.n3858 9.3005
R11285 gnd.n3898 gnd.n3857 9.3005
R11286 gnd.n3899 gnd.n3856 9.3005
R11287 gnd.n3902 gnd.n3855 9.3005
R11288 gnd.n3903 gnd.n3854 9.3005
R11289 gnd.n3906 gnd.n3853 9.3005
R11290 gnd.n3907 gnd.n3852 9.3005
R11291 gnd.n3910 gnd.n3851 9.3005
R11292 gnd.n3911 gnd.n3850 9.3005
R11293 gnd.n3914 gnd.n3849 9.3005
R11294 gnd.n3916 gnd.n3848 9.3005
R11295 gnd.n3917 gnd.n3847 9.3005
R11296 gnd.n3918 gnd.n3846 9.3005
R11297 gnd.n3919 gnd.n3845 9.3005
R11298 gnd.n3926 gnd.n3925 9.3005
R11299 gnd.n3935 gnd.n3934 9.3005
R11300 gnd.n3936 gnd.n3822 9.3005
R11301 gnd.n3938 gnd.n3937 9.3005
R11302 gnd.n3813 gnd.n3812 9.3005
R11303 gnd.n3951 gnd.n3950 9.3005
R11304 gnd.n3952 gnd.n3811 9.3005
R11305 gnd.n3954 gnd.n3953 9.3005
R11306 gnd.n3800 gnd.n3799 9.3005
R11307 gnd.n3997 gnd.n3996 9.3005
R11308 gnd.n3998 gnd.n3754 9.3005
R11309 gnd.n4002 gnd.n4000 9.3005
R11310 gnd.n4001 gnd.n3733 9.3005
R11311 gnd.n4020 gnd.n3732 9.3005
R11312 gnd.n4023 gnd.n4022 9.3005
R11313 gnd.n3726 gnd.n3725 9.3005
R11314 gnd.n4034 gnd.n4032 9.3005
R11315 gnd.n4033 gnd.n3707 9.3005
R11316 gnd.n4051 gnd.n3706 9.3005
R11317 gnd.n4054 gnd.n4053 9.3005
R11318 gnd.n3701 gnd.n3696 9.3005
R11319 gnd.n4064 gnd.n4063 9.3005
R11320 gnd.n3699 gnd.n3679 9.3005
R11321 gnd.n4085 gnd.n3680 9.3005
R11322 gnd.n4084 gnd.n4083 9.3005
R11323 gnd.n3682 gnd.n3658 9.3005
R11324 gnd.n4116 gnd.n4115 9.3005
R11325 gnd.n4118 gnd.n3603 9.3005
R11326 gnd.n4165 gnd.n3604 9.3005
R11327 gnd.n4164 gnd.n3605 9.3005
R11328 gnd.n4163 gnd.n3606 9.3005
R11329 gnd.n4129 gnd.n3607 9.3005
R11330 gnd.n4131 gnd.n3625 9.3005
R11331 gnd.n4151 gnd.n3626 9.3005
R11332 gnd.n4150 gnd.n3627 9.3005
R11333 gnd.n4149 gnd.n3628 9.3005
R11334 gnd.n4140 gnd.n3629 9.3005
R11335 gnd.n4141 gnd.n3512 9.3005
R11336 gnd.n4207 gnd.n4206 9.3005
R11337 gnd.n4208 gnd.n3505 9.3005
R11338 gnd.n4218 gnd.n4217 9.3005
R11339 gnd.n4220 gnd.n3501 9.3005
R11340 gnd.n4230 gnd.n3502 9.3005
R11341 gnd.n4229 gnd.n4228 9.3005
R11342 gnd.n4226 gnd.n3480 9.3005
R11343 gnd.n4252 gnd.n3481 9.3005
R11344 gnd.n4251 gnd.n4250 9.3005
R11345 gnd.n3483 gnd.n3457 9.3005
R11346 gnd.n4292 gnd.n4291 9.3005
R11347 gnd.n4293 gnd.n3450 9.3005
R11348 gnd.n4303 gnd.n4302 9.3005
R11349 gnd.n4305 gnd.n3446 9.3005
R11350 gnd.n4315 gnd.n3447 9.3005
R11351 gnd.n4314 gnd.n4313 9.3005
R11352 gnd.n4311 gnd.n3425 9.3005
R11353 gnd.n4337 gnd.n3426 9.3005
R11354 gnd.n4336 gnd.n4335 9.3005
R11355 gnd.n3428 gnd.n3403 9.3005
R11356 gnd.n4381 gnd.n4380 9.3005
R11357 gnd.n4382 gnd.n3396 9.3005
R11358 gnd.n4392 gnd.n4391 9.3005
R11359 gnd.n4650 gnd.n3392 9.3005
R11360 gnd.n4658 gnd.n3393 9.3005
R11361 gnd.n4657 gnd.n4656 9.3005
R11362 gnd.n2069 gnd.n2068 9.3005
R11363 gnd.n4681 gnd.n4680 9.3005
R11364 gnd.n3824 gnd.n3823 9.3005
R11365 gnd.n3163 gnd.n3162 9.3005
R11366 gnd.n3161 gnd.n2209 9.3005
R11367 gnd.n3160 gnd.n3159 9.3005
R11368 gnd.n2211 gnd.n2210 9.3005
R11369 gnd.n3153 gnd.n2215 9.3005
R11370 gnd.n3152 gnd.n2216 9.3005
R11371 gnd.n3151 gnd.n2217 9.3005
R11372 gnd.n2222 gnd.n2218 9.3005
R11373 gnd.n3145 gnd.n2223 9.3005
R11374 gnd.n3144 gnd.n2224 9.3005
R11375 gnd.n3143 gnd.n2225 9.3005
R11376 gnd.n2230 gnd.n2226 9.3005
R11377 gnd.n3137 gnd.n2231 9.3005
R11378 gnd.n3136 gnd.n2232 9.3005
R11379 gnd.n3135 gnd.n2233 9.3005
R11380 gnd.n2238 gnd.n2234 9.3005
R11381 gnd.n3129 gnd.n2239 9.3005
R11382 gnd.n3128 gnd.n2240 9.3005
R11383 gnd.n3127 gnd.n2241 9.3005
R11384 gnd.n2246 gnd.n2242 9.3005
R11385 gnd.n3121 gnd.n2247 9.3005
R11386 gnd.n3120 gnd.n2248 9.3005
R11387 gnd.n3119 gnd.n2249 9.3005
R11388 gnd.n2254 gnd.n2250 9.3005
R11389 gnd.n3113 gnd.n2255 9.3005
R11390 gnd.n3112 gnd.n2256 9.3005
R11391 gnd.n3111 gnd.n2257 9.3005
R11392 gnd.n2262 gnd.n2258 9.3005
R11393 gnd.n3105 gnd.n2263 9.3005
R11394 gnd.n3104 gnd.n2264 9.3005
R11395 gnd.n3103 gnd.n2265 9.3005
R11396 gnd.n2270 gnd.n2266 9.3005
R11397 gnd.n3097 gnd.n2271 9.3005
R11398 gnd.n3096 gnd.n2272 9.3005
R11399 gnd.n3095 gnd.n2273 9.3005
R11400 gnd.n2278 gnd.n2274 9.3005
R11401 gnd.n3089 gnd.n2279 9.3005
R11402 gnd.n3088 gnd.n2280 9.3005
R11403 gnd.n3087 gnd.n2281 9.3005
R11404 gnd.n2286 gnd.n2282 9.3005
R11405 gnd.n3081 gnd.n2287 9.3005
R11406 gnd.n3080 gnd.n2288 9.3005
R11407 gnd.n3079 gnd.n2289 9.3005
R11408 gnd.n2294 gnd.n2290 9.3005
R11409 gnd.n3073 gnd.n2295 9.3005
R11410 gnd.n3072 gnd.n2296 9.3005
R11411 gnd.n3071 gnd.n2297 9.3005
R11412 gnd.n2302 gnd.n2298 9.3005
R11413 gnd.n3065 gnd.n2303 9.3005
R11414 gnd.n3064 gnd.n2304 9.3005
R11415 gnd.n3063 gnd.n2305 9.3005
R11416 gnd.n2310 gnd.n2306 9.3005
R11417 gnd.n3057 gnd.n2311 9.3005
R11418 gnd.n3056 gnd.n2312 9.3005
R11419 gnd.n3055 gnd.n2313 9.3005
R11420 gnd.n2318 gnd.n2314 9.3005
R11421 gnd.n3049 gnd.n2319 9.3005
R11422 gnd.n3048 gnd.n2320 9.3005
R11423 gnd.n3047 gnd.n2321 9.3005
R11424 gnd.n2326 gnd.n2322 9.3005
R11425 gnd.n3041 gnd.n2327 9.3005
R11426 gnd.n3040 gnd.n2328 9.3005
R11427 gnd.n3039 gnd.n2329 9.3005
R11428 gnd.n2334 gnd.n2330 9.3005
R11429 gnd.n3033 gnd.n2335 9.3005
R11430 gnd.n3032 gnd.n2336 9.3005
R11431 gnd.n3031 gnd.n2337 9.3005
R11432 gnd.n2342 gnd.n2338 9.3005
R11433 gnd.n3025 gnd.n2343 9.3005
R11434 gnd.n3024 gnd.n2344 9.3005
R11435 gnd.n3023 gnd.n2345 9.3005
R11436 gnd.n2350 gnd.n2346 9.3005
R11437 gnd.n3017 gnd.n2351 9.3005
R11438 gnd.n3016 gnd.n2352 9.3005
R11439 gnd.n3015 gnd.n2353 9.3005
R11440 gnd.n2358 gnd.n2354 9.3005
R11441 gnd.n3009 gnd.n2359 9.3005
R11442 gnd.n3008 gnd.n2360 9.3005
R11443 gnd.n3007 gnd.n2361 9.3005
R11444 gnd.n2366 gnd.n2362 9.3005
R11445 gnd.n3001 gnd.n2367 9.3005
R11446 gnd.n3000 gnd.n2368 9.3005
R11447 gnd.n2999 gnd.n2369 9.3005
R11448 gnd.n2374 gnd.n2370 9.3005
R11449 gnd.n2993 gnd.n2375 9.3005
R11450 gnd.n2992 gnd.n2376 9.3005
R11451 gnd.n2991 gnd.n2377 9.3005
R11452 gnd.n2382 gnd.n2378 9.3005
R11453 gnd.n2985 gnd.n2383 9.3005
R11454 gnd.n2984 gnd.n2384 9.3005
R11455 gnd.n2983 gnd.n2385 9.3005
R11456 gnd.n2390 gnd.n2386 9.3005
R11457 gnd.n2977 gnd.n2391 9.3005
R11458 gnd.n2976 gnd.n2392 9.3005
R11459 gnd.n2975 gnd.n2393 9.3005
R11460 gnd.n2398 gnd.n2394 9.3005
R11461 gnd.n2969 gnd.n2399 9.3005
R11462 gnd.n2968 gnd.n2400 9.3005
R11463 gnd.n2967 gnd.n2401 9.3005
R11464 gnd.n2406 gnd.n2402 9.3005
R11465 gnd.n2961 gnd.n2407 9.3005
R11466 gnd.n2960 gnd.n2408 9.3005
R11467 gnd.n2959 gnd.n2409 9.3005
R11468 gnd.n2414 gnd.n2410 9.3005
R11469 gnd.n2953 gnd.n2415 9.3005
R11470 gnd.n2952 gnd.n2416 9.3005
R11471 gnd.n2951 gnd.n2417 9.3005
R11472 gnd.n2422 gnd.n2418 9.3005
R11473 gnd.n2945 gnd.n2423 9.3005
R11474 gnd.n2944 gnd.n2424 9.3005
R11475 gnd.n2943 gnd.n2425 9.3005
R11476 gnd.n2430 gnd.n2426 9.3005
R11477 gnd.n2937 gnd.n2431 9.3005
R11478 gnd.n2936 gnd.n2432 9.3005
R11479 gnd.n2935 gnd.n2433 9.3005
R11480 gnd.n2438 gnd.n2434 9.3005
R11481 gnd.n2929 gnd.n2439 9.3005
R11482 gnd.n2928 gnd.n2440 9.3005
R11483 gnd.n2927 gnd.n2441 9.3005
R11484 gnd.n2446 gnd.n2442 9.3005
R11485 gnd.n2921 gnd.n2447 9.3005
R11486 gnd.n2920 gnd.n2448 9.3005
R11487 gnd.n2919 gnd.n2449 9.3005
R11488 gnd.n2454 gnd.n2450 9.3005
R11489 gnd.n2913 gnd.n2455 9.3005
R11490 gnd.n2912 gnd.n2456 9.3005
R11491 gnd.n2911 gnd.n2457 9.3005
R11492 gnd.n2462 gnd.n2458 9.3005
R11493 gnd.n2905 gnd.n2463 9.3005
R11494 gnd.n2904 gnd.n2464 9.3005
R11495 gnd.n2903 gnd.n2465 9.3005
R11496 gnd.n2470 gnd.n2466 9.3005
R11497 gnd.n2897 gnd.n2471 9.3005
R11498 gnd.n2896 gnd.n2472 9.3005
R11499 gnd.n2895 gnd.n2473 9.3005
R11500 gnd.n2478 gnd.n2474 9.3005
R11501 gnd.n2889 gnd.n2479 9.3005
R11502 gnd.n2888 gnd.n2480 9.3005
R11503 gnd.n2887 gnd.n2481 9.3005
R11504 gnd.n2486 gnd.n2482 9.3005
R11505 gnd.n2881 gnd.n2487 9.3005
R11506 gnd.n2880 gnd.n2488 9.3005
R11507 gnd.n2879 gnd.n2489 9.3005
R11508 gnd.n2494 gnd.n2490 9.3005
R11509 gnd.n2873 gnd.n2495 9.3005
R11510 gnd.n2872 gnd.n2496 9.3005
R11511 gnd.n2871 gnd.n2497 9.3005
R11512 gnd.n2502 gnd.n2498 9.3005
R11513 gnd.n2865 gnd.n2503 9.3005
R11514 gnd.n2864 gnd.n2504 9.3005
R11515 gnd.n2863 gnd.n2505 9.3005
R11516 gnd.n2510 gnd.n2506 9.3005
R11517 gnd.n2857 gnd.n2511 9.3005
R11518 gnd.n2856 gnd.n2512 9.3005
R11519 gnd.n2855 gnd.n2513 9.3005
R11520 gnd.n2849 gnd.n2848 9.3005
R11521 gnd.n2847 gnd.n2518 9.3005
R11522 gnd.n2846 gnd.n2845 9.3005
R11523 gnd.n2521 gnd.n2520 9.3005
R11524 gnd.n2839 gnd.n2525 9.3005
R11525 gnd.n2838 gnd.n2526 9.3005
R11526 gnd.n2837 gnd.n2527 9.3005
R11527 gnd.n2532 gnd.n2528 9.3005
R11528 gnd.n2831 gnd.n2533 9.3005
R11529 gnd.n2830 gnd.n2534 9.3005
R11530 gnd.n2829 gnd.n2535 9.3005
R11531 gnd.n2540 gnd.n2536 9.3005
R11532 gnd.n2823 gnd.n2541 9.3005
R11533 gnd.n2822 gnd.n2542 9.3005
R11534 gnd.n2821 gnd.n2543 9.3005
R11535 gnd.n2548 gnd.n2544 9.3005
R11536 gnd.n2815 gnd.n2549 9.3005
R11537 gnd.n2814 gnd.n2550 9.3005
R11538 gnd.n2813 gnd.n2551 9.3005
R11539 gnd.n2556 gnd.n2552 9.3005
R11540 gnd.n2807 gnd.n2557 9.3005
R11541 gnd.n2806 gnd.n2558 9.3005
R11542 gnd.n2805 gnd.n2559 9.3005
R11543 gnd.n2564 gnd.n2560 9.3005
R11544 gnd.n2799 gnd.n2565 9.3005
R11545 gnd.n2798 gnd.n2566 9.3005
R11546 gnd.n2797 gnd.n2567 9.3005
R11547 gnd.n2572 gnd.n2568 9.3005
R11548 gnd.n2791 gnd.n2573 9.3005
R11549 gnd.n2790 gnd.n2574 9.3005
R11550 gnd.n2789 gnd.n2575 9.3005
R11551 gnd.n2580 gnd.n2576 9.3005
R11552 gnd.n2783 gnd.n2581 9.3005
R11553 gnd.n2782 gnd.n2582 9.3005
R11554 gnd.n2781 gnd.n2583 9.3005
R11555 gnd.n2588 gnd.n2584 9.3005
R11556 gnd.n2775 gnd.n2589 9.3005
R11557 gnd.n2774 gnd.n2590 9.3005
R11558 gnd.n2773 gnd.n2591 9.3005
R11559 gnd.n2596 gnd.n2592 9.3005
R11560 gnd.n2767 gnd.n2597 9.3005
R11561 gnd.n2766 gnd.n2598 9.3005
R11562 gnd.n2765 gnd.n2599 9.3005
R11563 gnd.n2604 gnd.n2600 9.3005
R11564 gnd.n2759 gnd.n2605 9.3005
R11565 gnd.n2758 gnd.n2606 9.3005
R11566 gnd.n2757 gnd.n2607 9.3005
R11567 gnd.n2612 gnd.n2608 9.3005
R11568 gnd.n2751 gnd.n2613 9.3005
R11569 gnd.n2750 gnd.n2614 9.3005
R11570 gnd.n2749 gnd.n2615 9.3005
R11571 gnd.n2620 gnd.n2616 9.3005
R11572 gnd.n2743 gnd.n2621 9.3005
R11573 gnd.n2742 gnd.n2622 9.3005
R11574 gnd.n2741 gnd.n2623 9.3005
R11575 gnd.n2628 gnd.n2624 9.3005
R11576 gnd.n2735 gnd.n2629 9.3005
R11577 gnd.n2734 gnd.n2630 9.3005
R11578 gnd.n2733 gnd.n2631 9.3005
R11579 gnd.n2636 gnd.n2632 9.3005
R11580 gnd.n2727 gnd.n2637 9.3005
R11581 gnd.n2726 gnd.n2638 9.3005
R11582 gnd.n2725 gnd.n2639 9.3005
R11583 gnd.n2644 gnd.n2640 9.3005
R11584 gnd.n2719 gnd.n2645 9.3005
R11585 gnd.n2718 gnd.n2646 9.3005
R11586 gnd.n2717 gnd.n2647 9.3005
R11587 gnd.n2652 gnd.n2648 9.3005
R11588 gnd.n2711 gnd.n2653 9.3005
R11589 gnd.n2710 gnd.n2654 9.3005
R11590 gnd.n2709 gnd.n2655 9.3005
R11591 gnd.n2660 gnd.n2656 9.3005
R11592 gnd.n2703 gnd.n2661 9.3005
R11593 gnd.n2702 gnd.n2662 9.3005
R11594 gnd.n2701 gnd.n2663 9.3005
R11595 gnd.n2668 gnd.n2664 9.3005
R11596 gnd.n2695 gnd.n2669 9.3005
R11597 gnd.n2694 gnd.n2670 9.3005
R11598 gnd.n2693 gnd.n2671 9.3005
R11599 gnd.n2676 gnd.n2672 9.3005
R11600 gnd.n2687 gnd.n2677 9.3005
R11601 gnd.n2686 gnd.n2678 9.3005
R11602 gnd.n2685 gnd.n2679 9.3005
R11603 gnd.n2681 gnd.n2680 9.3005
R11604 gnd.n2519 gnd.n2517 9.3005
R11605 gnd.n7757 gnd.n7756 9.3005
R11606 gnd.n7755 gnd.n84 9.3005
R11607 gnd.n7437 gnd.n87 9.3005
R11608 gnd.n7470 gnd.n7438 9.3005
R11609 gnd.n7469 gnd.n7439 9.3005
R11610 gnd.n7468 gnd.n7440 9.3005
R11611 gnd.n7466 gnd.n7441 9.3005
R11612 gnd.n7465 gnd.n7442 9.3005
R11613 gnd.n7463 gnd.n7443 9.3005
R11614 gnd.n7462 gnd.n7444 9.3005
R11615 gnd.n7460 gnd.n7445 9.3005
R11616 gnd.n7459 gnd.n7446 9.3005
R11617 gnd.n7457 gnd.n7447 9.3005
R11618 gnd.n7456 gnd.n7448 9.3005
R11619 gnd.n7454 gnd.n7449 9.3005
R11620 gnd.n7453 gnd.n7451 9.3005
R11621 gnd.n7450 gnd.n358 9.3005
R11622 gnd.n7516 gnd.n357 9.3005
R11623 gnd.n7518 gnd.n7517 9.3005
R11624 gnd.n7519 gnd.n356 9.3005
R11625 gnd.n7521 gnd.n7520 9.3005
R11626 gnd.n7523 gnd.n354 9.3005
R11627 gnd.n7525 gnd.n7524 9.3005
R11628 gnd.n7526 gnd.n353 9.3005
R11629 gnd.n7528 gnd.n7527 9.3005
R11630 gnd.n7530 gnd.n351 9.3005
R11631 gnd.n7532 gnd.n7531 9.3005
R11632 gnd.n7563 gnd.n317 9.3005
R11633 gnd.n7562 gnd.n319 9.3005
R11634 gnd.n323 gnd.n320 9.3005
R11635 gnd.n7557 gnd.n324 9.3005
R11636 gnd.n7556 gnd.n325 9.3005
R11637 gnd.n7555 gnd.n326 9.3005
R11638 gnd.n330 gnd.n327 9.3005
R11639 gnd.n7550 gnd.n331 9.3005
R11640 gnd.n7549 gnd.n332 9.3005
R11641 gnd.n7548 gnd.n333 9.3005
R11642 gnd.n337 gnd.n334 9.3005
R11643 gnd.n7543 gnd.n338 9.3005
R11644 gnd.n7542 gnd.n339 9.3005
R11645 gnd.n7541 gnd.n340 9.3005
R11646 gnd.n344 gnd.n341 9.3005
R11647 gnd.n7536 gnd.n345 9.3005
R11648 gnd.n7535 gnd.n7534 9.3005
R11649 gnd.n7533 gnd.n348 9.3005
R11650 gnd.n7565 gnd.n7564 9.3005
R11651 gnd.n7673 gnd.n214 9.3005
R11652 gnd.n7672 gnd.n216 9.3005
R11653 gnd.n220 gnd.n217 9.3005
R11654 gnd.n7667 gnd.n221 9.3005
R11655 gnd.n7666 gnd.n222 9.3005
R11656 gnd.n7665 gnd.n223 9.3005
R11657 gnd.n227 gnd.n224 9.3005
R11658 gnd.n7660 gnd.n228 9.3005
R11659 gnd.n7659 gnd.n229 9.3005
R11660 gnd.n7658 gnd.n230 9.3005
R11661 gnd.n234 gnd.n231 9.3005
R11662 gnd.n7653 gnd.n235 9.3005
R11663 gnd.n7652 gnd.n236 9.3005
R11664 gnd.n7651 gnd.n237 9.3005
R11665 gnd.n241 gnd.n238 9.3005
R11666 gnd.n7646 gnd.n242 9.3005
R11667 gnd.n7645 gnd.n243 9.3005
R11668 gnd.n7641 gnd.n244 9.3005
R11669 gnd.n248 gnd.n245 9.3005
R11670 gnd.n7636 gnd.n249 9.3005
R11671 gnd.n7635 gnd.n250 9.3005
R11672 gnd.n7634 gnd.n251 9.3005
R11673 gnd.n255 gnd.n252 9.3005
R11674 gnd.n7629 gnd.n256 9.3005
R11675 gnd.n7628 gnd.n257 9.3005
R11676 gnd.n7627 gnd.n258 9.3005
R11677 gnd.n262 gnd.n259 9.3005
R11678 gnd.n7622 gnd.n263 9.3005
R11679 gnd.n7621 gnd.n264 9.3005
R11680 gnd.n7620 gnd.n265 9.3005
R11681 gnd.n269 gnd.n266 9.3005
R11682 gnd.n7615 gnd.n270 9.3005
R11683 gnd.n7614 gnd.n271 9.3005
R11684 gnd.n7613 gnd.n272 9.3005
R11685 gnd.n276 gnd.n273 9.3005
R11686 gnd.n7608 gnd.n277 9.3005
R11687 gnd.n7607 gnd.n7606 9.3005
R11688 gnd.n7605 gnd.n278 9.3005
R11689 gnd.n7604 gnd.n7603 9.3005
R11690 gnd.n282 gnd.n281 9.3005
R11691 gnd.n287 gnd.n285 9.3005
R11692 gnd.n7596 gnd.n288 9.3005
R11693 gnd.n7595 gnd.n289 9.3005
R11694 gnd.n7594 gnd.n290 9.3005
R11695 gnd.n294 gnd.n291 9.3005
R11696 gnd.n7589 gnd.n295 9.3005
R11697 gnd.n7588 gnd.n296 9.3005
R11698 gnd.n7587 gnd.n297 9.3005
R11699 gnd.n301 gnd.n298 9.3005
R11700 gnd.n7582 gnd.n302 9.3005
R11701 gnd.n7581 gnd.n303 9.3005
R11702 gnd.n7580 gnd.n304 9.3005
R11703 gnd.n308 gnd.n305 9.3005
R11704 gnd.n7575 gnd.n309 9.3005
R11705 gnd.n7574 gnd.n310 9.3005
R11706 gnd.n7573 gnd.n311 9.3005
R11707 gnd.n316 gnd.n314 9.3005
R11708 gnd.n7568 gnd.n7567 9.3005
R11709 gnd.n7675 gnd.n7674 9.3005
R11710 gnd.n7095 gnd.n7094 9.3005
R11711 gnd.n513 gnd.n507 9.3005
R11712 gnd.n7239 gnd.n508 9.3005
R11713 gnd.n7238 gnd.n509 9.3005
R11714 gnd.n7237 gnd.n510 9.3005
R11715 gnd.n7236 gnd.n7234 9.3005
R11716 gnd.n511 gnd.n472 9.3005
R11717 gnd.n7285 gnd.n473 9.3005
R11718 gnd.n7284 gnd.n474 9.3005
R11719 gnd.n7283 gnd.n475 9.3005
R11720 gnd.n7282 gnd.n7280 9.3005
R11721 gnd.n476 gnd.n437 9.3005
R11722 gnd.n7332 gnd.n438 9.3005
R11723 gnd.n7331 gnd.n439 9.3005
R11724 gnd.n7330 gnd.n440 9.3005
R11725 gnd.n7329 gnd.n441 9.3005
R11726 gnd.n7323 gnd.n404 9.3005
R11727 gnd.n7376 gnd.n405 9.3005
R11728 gnd.n7375 gnd.n406 9.3005
R11729 gnd.n7374 gnd.n7369 9.3005
R11730 gnd.n7373 gnd.n7370 9.3005
R11731 gnd.n380 gnd.n379 9.3005
R11732 gnd.n7409 gnd.n7408 9.3005
R11733 gnd.n368 gnd.n367 9.3005
R11734 gnd.n7422 gnd.n7421 9.3005
R11735 gnd.n7423 gnd.n361 9.3005
R11736 gnd.n7430 gnd.n362 9.3005
R11737 gnd.n7431 gnd.n360 9.3005
R11738 gnd.n7434 gnd.n7433 9.3005
R11739 gnd.n7435 gnd.n110 9.3005
R11740 gnd.n7743 gnd.n111 9.3005
R11741 gnd.n7742 gnd.n112 9.3005
R11742 gnd.n7741 gnd.n113 9.3005
R11743 gnd.n7479 gnd.n114 9.3005
R11744 gnd.n7731 gnd.n128 9.3005
R11745 gnd.n7730 gnd.n129 9.3005
R11746 gnd.n7729 gnd.n130 9.3005
R11747 gnd.n7486 gnd.n131 9.3005
R11748 gnd.n7719 gnd.n148 9.3005
R11749 gnd.n7718 gnd.n149 9.3005
R11750 gnd.n7717 gnd.n150 9.3005
R11751 gnd.n7493 gnd.n151 9.3005
R11752 gnd.n7707 gnd.n166 9.3005
R11753 gnd.n7706 gnd.n167 9.3005
R11754 gnd.n7705 gnd.n168 9.3005
R11755 gnd.n7497 gnd.n169 9.3005
R11756 gnd.n7695 gnd.n186 9.3005
R11757 gnd.n7694 gnd.n187 9.3005
R11758 gnd.n7693 gnd.n188 9.3005
R11759 gnd.n7498 gnd.n189 9.3005
R11760 gnd.n7683 gnd.n204 9.3005
R11761 gnd.n7682 gnd.n205 9.3005
R11762 gnd.n7681 gnd.n206 9.3005
R11763 gnd.n7093 gnd.n7091 9.3005
R11764 gnd.n7094 gnd.n512 9.3005
R11765 gnd.n7225 gnd.n513 9.3005
R11766 gnd.n7226 gnd.n508 9.3005
R11767 gnd.n7229 gnd.n509 9.3005
R11768 gnd.n7230 gnd.n510 9.3005
R11769 gnd.n7234 gnd.n7233 9.3005
R11770 gnd.n7231 gnd.n511 9.3005
R11771 gnd.n477 gnd.n473 9.3005
R11772 gnd.n7275 gnd.n474 9.3005
R11773 gnd.n7276 gnd.n475 9.3005
R11774 gnd.n7280 gnd.n7279 9.3005
R11775 gnd.n7277 gnd.n476 9.3005
R11776 gnd.n442 gnd.n438 9.3005
R11777 gnd.n7321 gnd.n439 9.3005
R11778 gnd.n7322 gnd.n440 9.3005
R11779 gnd.n7325 gnd.n441 9.3005
R11780 gnd.n7324 gnd.n7323 9.3005
R11781 gnd.n407 gnd.n405 9.3005
R11782 gnd.n7367 gnd.n406 9.3005
R11783 gnd.n7369 gnd.n7368 9.3005
R11784 gnd.n7370 gnd.n381 9.3005
R11785 gnd.n7404 gnd.n380 9.3005
R11786 gnd.n7408 gnd.n7407 9.3005
R11787 gnd.n7406 gnd.n367 9.3005
R11788 gnd.n7422 gnd.n366 9.3005
R11789 gnd.n7424 gnd.n7423 9.3005
R11790 gnd.n7426 gnd.n362 9.3005
R11791 gnd.n7425 gnd.n360 9.3005
R11792 gnd.n7434 gnd.n359 9.3005
R11793 gnd.n7474 gnd.n7435 9.3005
R11794 gnd.n7475 gnd.n111 9.3005
R11795 gnd.n7477 gnd.n112 9.3005
R11796 gnd.n7478 gnd.n113 9.3005
R11797 gnd.n7481 gnd.n7479 9.3005
R11798 gnd.n7482 gnd.n128 9.3005
R11799 gnd.n7484 gnd.n129 9.3005
R11800 gnd.n7485 gnd.n130 9.3005
R11801 gnd.n7488 gnd.n7486 9.3005
R11802 gnd.n7489 gnd.n148 9.3005
R11803 gnd.n7491 gnd.n149 9.3005
R11804 gnd.n7492 gnd.n150 9.3005
R11805 gnd.n7495 gnd.n7493 9.3005
R11806 gnd.n7496 gnd.n166 9.3005
R11807 gnd.n7512 gnd.n167 9.3005
R11808 gnd.n7511 gnd.n168 9.3005
R11809 gnd.n7510 gnd.n7497 9.3005
R11810 gnd.n7508 gnd.n186 9.3005
R11811 gnd.n7507 gnd.n187 9.3005
R11812 gnd.n7505 gnd.n188 9.3005
R11813 gnd.n7504 gnd.n7498 9.3005
R11814 gnd.n7502 gnd.n204 9.3005
R11815 gnd.n7501 gnd.n205 9.3005
R11816 gnd.n7499 gnd.n206 9.3005
R11817 gnd.n7093 gnd.n7092 9.3005
R11818 gnd.n899 gnd.n898 9.3005
R11819 gnd.n902 gnd.n892 9.3005
R11820 gnd.n903 gnd.n891 9.3005
R11821 gnd.n906 gnd.n890 9.3005
R11822 gnd.n907 gnd.n889 9.3005
R11823 gnd.n910 gnd.n888 9.3005
R11824 gnd.n911 gnd.n887 9.3005
R11825 gnd.n914 gnd.n886 9.3005
R11826 gnd.n915 gnd.n885 9.3005
R11827 gnd.n918 gnd.n884 9.3005
R11828 gnd.n919 gnd.n883 9.3005
R11829 gnd.n922 gnd.n882 9.3005
R11830 gnd.n923 gnd.n881 9.3005
R11831 gnd.n926 gnd.n880 9.3005
R11832 gnd.n927 gnd.n879 9.3005
R11833 gnd.n930 gnd.n878 9.3005
R11834 gnd.n931 gnd.n877 9.3005
R11835 gnd.n934 gnd.n876 9.3005
R11836 gnd.n935 gnd.n875 9.3005
R11837 gnd.n938 gnd.n874 9.3005
R11838 gnd.n942 gnd.n870 9.3005
R11839 gnd.n943 gnd.n869 9.3005
R11840 gnd.n946 gnd.n868 9.3005
R11841 gnd.n947 gnd.n867 9.3005
R11842 gnd.n950 gnd.n866 9.3005
R11843 gnd.n951 gnd.n865 9.3005
R11844 gnd.n954 gnd.n864 9.3005
R11845 gnd.n955 gnd.n863 9.3005
R11846 gnd.n958 gnd.n862 9.3005
R11847 gnd.n860 gnd.n787 9.3005
R11848 gnd.n859 gnd.n858 9.3005
R11849 gnd.n855 gnd.n789 9.3005
R11850 gnd.n852 gnd.n851 9.3005
R11851 gnd.n850 gnd.n790 9.3005
R11852 gnd.n849 gnd.n848 9.3005
R11853 gnd.n845 gnd.n791 9.3005
R11854 gnd.n842 gnd.n841 9.3005
R11855 gnd.n840 gnd.n839 9.3005
R11856 gnd.n836 gnd.n795 9.3005
R11857 gnd.n835 gnd.n832 9.3005
R11858 gnd.n831 gnd.n796 9.3005
R11859 gnd.n830 gnd.n829 9.3005
R11860 gnd.n826 gnd.n797 9.3005
R11861 gnd.n825 gnd.n822 9.3005
R11862 gnd.n821 gnd.n798 9.3005
R11863 gnd.n820 gnd.n819 9.3005
R11864 gnd.n816 gnd.n799 9.3005
R11865 gnd.n815 gnd.n812 9.3005
R11866 gnd.n811 gnd.n800 9.3005
R11867 gnd.n810 gnd.n809 9.3005
R11868 gnd.n806 gnd.n801 9.3005
R11869 gnd.n805 gnd.n803 9.3005
R11870 gnd.n802 gnd.n527 9.3005
R11871 gnd.n7206 gnd.n526 9.3005
R11872 gnd.n7208 gnd.n7207 9.3005
R11873 gnd.n939 gnd.n871 9.3005
R11874 gnd.n897 gnd.n894 9.3005
R11875 gnd.n7211 gnd.n7210 9.3005
R11876 gnd.n499 gnd.n498 9.3005
R11877 gnd.n7244 gnd.n7243 9.3005
R11878 gnd.n7245 gnd.n497 9.3005
R11879 gnd.n7249 gnd.n7246 9.3005
R11880 gnd.n7248 gnd.n7247 9.3005
R11881 gnd.n464 gnd.n463 9.3005
R11882 gnd.n7290 gnd.n7289 9.3005
R11883 gnd.n7291 gnd.n462 9.3005
R11884 gnd.n7295 gnd.n7292 9.3005
R11885 gnd.n7294 gnd.n7293 9.3005
R11886 gnd.n429 gnd.n428 9.3005
R11887 gnd.n7337 gnd.n7336 9.3005
R11888 gnd.n7338 gnd.n427 9.3005
R11889 gnd.n7342 gnd.n7339 9.3005
R11890 gnd.n7341 gnd.n7340 9.3005
R11891 gnd.n397 gnd.n396 9.3005
R11892 gnd.n7381 gnd.n7380 9.3005
R11893 gnd.n7382 gnd.n395 9.3005
R11894 gnd.n7386 gnd.n7383 9.3005
R11895 gnd.n7385 gnd.n97 9.3005
R11896 gnd.n102 gnd.n96 9.3005
R11897 gnd.n7737 gnd.n119 9.3005
R11898 gnd.n7736 gnd.n120 9.3005
R11899 gnd.n7735 gnd.n121 9.3005
R11900 gnd.n138 gnd.n122 9.3005
R11901 gnd.n7725 gnd.n139 9.3005
R11902 gnd.n7724 gnd.n140 9.3005
R11903 gnd.n7723 gnd.n141 9.3005
R11904 gnd.n156 gnd.n142 9.3005
R11905 gnd.n7713 gnd.n157 9.3005
R11906 gnd.n7712 gnd.n158 9.3005
R11907 gnd.n7711 gnd.n159 9.3005
R11908 gnd.n176 gnd.n160 9.3005
R11909 gnd.n7701 gnd.n177 9.3005
R11910 gnd.n7700 gnd.n178 9.3005
R11911 gnd.n7699 gnd.n179 9.3005
R11912 gnd.n195 gnd.n180 9.3005
R11913 gnd.n7689 gnd.n196 9.3005
R11914 gnd.n7688 gnd.n197 9.3005
R11915 gnd.n7687 gnd.n198 9.3005
R11916 gnd.n213 gnd.n199 9.3005
R11917 gnd.n7677 gnd.n7676 9.3005
R11918 gnd.n7212 gnd.n7209 9.3005
R11919 gnd.n7748 gnd.n100 9.3005
R11920 gnd.n7748 gnd.n7747 9.3005
R11921 gnd.n4927 gnd.n4896 9.3005
R11922 gnd.n4926 gnd.n4897 9.3005
R11923 gnd.n4924 gnd.n4898 9.3005
R11924 gnd.n4923 gnd.n4899 9.3005
R11925 gnd.n4921 gnd.n4900 9.3005
R11926 gnd.n4920 gnd.n4901 9.3005
R11927 gnd.n4918 gnd.n4902 9.3005
R11928 gnd.n4917 gnd.n4903 9.3005
R11929 gnd.n4915 gnd.n4904 9.3005
R11930 gnd.n4914 gnd.n4905 9.3005
R11931 gnd.n4912 gnd.n4906 9.3005
R11932 gnd.n4911 gnd.n4907 9.3005
R11933 gnd.n4909 gnd.n4908 9.3005
R11934 gnd.n1913 gnd.n1912 9.3005
R11935 gnd.n5175 gnd.n5174 9.3005
R11936 gnd.n5176 gnd.n1911 9.3005
R11937 gnd.n5180 gnd.n5177 9.3005
R11938 gnd.n5179 gnd.n5178 9.3005
R11939 gnd.n1888 gnd.n1887 9.3005
R11940 gnd.n5210 gnd.n5209 9.3005
R11941 gnd.n5211 gnd.n1886 9.3005
R11942 gnd.n5224 gnd.n5212 9.3005
R11943 gnd.n5223 gnd.n5213 9.3005
R11944 gnd.n5222 gnd.n5214 9.3005
R11945 gnd.n5220 gnd.n5215 9.3005
R11946 gnd.n5219 gnd.n5217 9.3005
R11947 gnd.n4930 gnd.n4929 9.3005
R11948 gnd.n4935 gnd.n4934 9.3005
R11949 gnd.n4938 gnd.n4891 9.3005
R11950 gnd.n4939 gnd.n4890 9.3005
R11951 gnd.n4942 gnd.n4889 9.3005
R11952 gnd.n4943 gnd.n4888 9.3005
R11953 gnd.n4946 gnd.n4887 9.3005
R11954 gnd.n4947 gnd.n4886 9.3005
R11955 gnd.n4950 gnd.n4885 9.3005
R11956 gnd.n4951 gnd.n4884 9.3005
R11957 gnd.n4954 gnd.n4883 9.3005
R11958 gnd.n4955 gnd.n4882 9.3005
R11959 gnd.n4958 gnd.n4881 9.3005
R11960 gnd.n4959 gnd.n4880 9.3005
R11961 gnd.n4962 gnd.n4879 9.3005
R11962 gnd.n4963 gnd.n4878 9.3005
R11963 gnd.n4966 gnd.n4877 9.3005
R11964 gnd.n4969 gnd.n4968 9.3005
R11965 gnd.n4933 gnd.n4895 9.3005
R11966 gnd.n4932 gnd.n4931 9.3005
R11967 gnd.n1592 gnd.n1590 9.3005
R11968 gnd.n5816 gnd.n5811 9.3005
R11969 gnd.n5817 gnd.n5810 9.3005
R11970 gnd.n5818 gnd.n5809 9.3005
R11971 gnd.n5808 gnd.n5805 9.3005
R11972 gnd.n5823 gnd.n5804 9.3005
R11973 gnd.n5824 gnd.n5803 9.3005
R11974 gnd.n5825 gnd.n5802 9.3005
R11975 gnd.n5801 gnd.n5795 9.3005
R11976 gnd.n5830 gnd.n5794 9.3005
R11977 gnd.n5831 gnd.n5793 9.3005
R11978 gnd.n5832 gnd.n5792 9.3005
R11979 gnd.n5791 gnd.n5788 9.3005
R11980 gnd.n5837 gnd.n5787 9.3005
R11981 gnd.n5838 gnd.n5786 9.3005
R11982 gnd.n5839 gnd.n5785 9.3005
R11983 gnd.n5784 gnd.n5781 9.3005
R11984 gnd.n5844 gnd.n5780 9.3005
R11985 gnd.n5845 gnd.n5779 9.3005
R11986 gnd.n5846 gnd.n5778 9.3005
R11987 gnd.n5777 gnd.n5774 9.3005
R11988 gnd.n5851 gnd.n5773 9.3005
R11989 gnd.n5852 gnd.n5772 9.3005
R11990 gnd.n5853 gnd.n5771 9.3005
R11991 gnd.n5769 gnd.n5768 9.3005
R11992 gnd.n5859 gnd.n5858 9.3005
R11993 gnd.n5926 gnd.n5925 9.3005
R11994 gnd.n1594 gnd.n1593 9.3005
R11995 gnd.n1600 gnd.n1598 9.3005
R11996 gnd.n5918 gnd.n1601 9.3005
R11997 gnd.n5917 gnd.n1602 9.3005
R11998 gnd.n5916 gnd.n1603 9.3005
R11999 gnd.n1607 gnd.n1604 9.3005
R12000 gnd.n5911 gnd.n1608 9.3005
R12001 gnd.n5910 gnd.n5909 9.3005
R12002 gnd.n5908 gnd.n1609 9.3005
R12003 gnd.n5907 gnd.n5906 9.3005
R12004 gnd.n1613 gnd.n1612 9.3005
R12005 gnd.n1618 gnd.n1616 9.3005
R12006 gnd.n5899 gnd.n1619 9.3005
R12007 gnd.n5898 gnd.n1620 9.3005
R12008 gnd.n5897 gnd.n1621 9.3005
R12009 gnd.n1625 gnd.n1622 9.3005
R12010 gnd.n5892 gnd.n1626 9.3005
R12011 gnd.n5891 gnd.n1627 9.3005
R12012 gnd.n5890 gnd.n1628 9.3005
R12013 gnd.n1632 gnd.n1629 9.3005
R12014 gnd.n5885 gnd.n1633 9.3005
R12015 gnd.n5884 gnd.n1634 9.3005
R12016 gnd.n5883 gnd.n1635 9.3005
R12017 gnd.n1639 gnd.n1636 9.3005
R12018 gnd.n5878 gnd.n1640 9.3005
R12019 gnd.n5877 gnd.n1641 9.3005
R12020 gnd.n5876 gnd.n1642 9.3005
R12021 gnd.n1648 gnd.n1645 9.3005
R12022 gnd.n5871 gnd.n5870 9.3005
R12023 gnd.n5927 gnd.n1589 9.3005
R12024 gnd.n5096 gnd.n5095 9.3005
R12025 gnd.n1989 gnd.n1985 9.3005
R12026 gnd.n1988 gnd.n1987 9.3005
R12027 gnd.n1969 gnd.n1966 9.3005
R12028 gnd.n5116 gnd.n1967 9.3005
R12029 gnd.n5115 gnd.n5112 9.3005
R12030 gnd.n5114 gnd.n5113 9.3005
R12031 gnd.n1951 gnd.n1948 9.3005
R12032 gnd.n5136 gnd.n1949 9.3005
R12033 gnd.n5135 gnd.n5132 9.3005
R12034 gnd.n5134 gnd.n5133 9.3005
R12035 gnd.n1933 gnd.n1929 9.3005
R12036 gnd.n5160 gnd.n1930 9.3005
R12037 gnd.n5159 gnd.n1931 9.3005
R12038 gnd.n5158 gnd.n5154 9.3005
R12039 gnd.n5157 gnd.n5155 9.3005
R12040 gnd.n1907 gnd.n1903 9.3005
R12041 gnd.n5195 gnd.n1904 9.3005
R12042 gnd.n5194 gnd.n1905 9.3005
R12043 gnd.n5193 gnd.n5189 9.3005
R12044 gnd.n5192 gnd.n5190 9.3005
R12045 gnd.n1882 gnd.n1879 9.3005
R12046 gnd.n5235 gnd.n1880 9.3005
R12047 gnd.n5234 gnd.n5231 9.3005
R12048 gnd.n5233 gnd.n5232 9.3005
R12049 gnd.n1868 gnd.n1865 9.3005
R12050 gnd.n5253 gnd.n1866 9.3005
R12051 gnd.n5252 gnd.n5248 9.3005
R12052 gnd.n5251 gnd.n5249 9.3005
R12053 gnd.n1848 gnd.n1842 9.3005
R12054 gnd.n5291 gnd.n1843 9.3005
R12055 gnd.n5290 gnd.n1844 9.3005
R12056 gnd.n5289 gnd.n1845 9.3005
R12057 gnd.n5288 gnd.n5286 9.3005
R12058 gnd.n1846 gnd.n1801 9.3005
R12059 gnd.n5331 gnd.n1802 9.3005
R12060 gnd.n5330 gnd.n1803 9.3005
R12061 gnd.n5329 gnd.n1804 9.3005
R12062 gnd.n5328 gnd.n1805 9.3005
R12063 gnd.n1777 gnd.n1765 9.3005
R12064 gnd.n5379 gnd.n1766 9.3005
R12065 gnd.n5378 gnd.n1767 9.3005
R12066 gnd.n5377 gnd.n1768 9.3005
R12067 gnd.n5376 gnd.n1769 9.3005
R12068 gnd.n1742 gnd.n1739 9.3005
R12069 gnd.n5413 gnd.n1740 9.3005
R12070 gnd.n5412 gnd.n5409 9.3005
R12071 gnd.n5411 gnd.n5410 9.3005
R12072 gnd.n1671 gnd.n1670 9.3005
R12073 gnd.n5760 gnd.n5756 9.3005
R12074 gnd.n5759 gnd.n5757 9.3005
R12075 gnd.n5758 gnd.n1650 9.3005
R12076 gnd.n5868 gnd.n1651 9.3005
R12077 gnd.n1986 gnd.n1984 9.3005
R12078 gnd.n5095 gnd.n5094 9.3005
R12079 gnd.n5093 gnd.n1989 9.3005
R12080 gnd.n1988 gnd.n1968 9.3005
R12081 gnd.n5109 gnd.n1969 9.3005
R12082 gnd.n5110 gnd.n1967 9.3005
R12083 gnd.n5112 gnd.n5111 9.3005
R12084 gnd.n5113 gnd.n1950 9.3005
R12085 gnd.n5129 gnd.n1951 9.3005
R12086 gnd.n5130 gnd.n1949 9.3005
R12087 gnd.n5132 gnd.n5131 9.3005
R12088 gnd.n5133 gnd.n1932 9.3005
R12089 gnd.n5149 gnd.n1933 9.3005
R12090 gnd.n5150 gnd.n1930 9.3005
R12091 gnd.n5152 gnd.n1931 9.3005
R12092 gnd.n5154 gnd.n5153 9.3005
R12093 gnd.n5155 gnd.n1906 9.3005
R12094 gnd.n5184 gnd.n1907 9.3005
R12095 gnd.n5185 gnd.n1904 9.3005
R12096 gnd.n5187 gnd.n1905 9.3005
R12097 gnd.n5189 gnd.n5188 9.3005
R12098 gnd.n5190 gnd.n1881 9.3005
R12099 gnd.n5228 gnd.n1882 9.3005
R12100 gnd.n5229 gnd.n1880 9.3005
R12101 gnd.n5231 gnd.n5230 9.3005
R12102 gnd.n5232 gnd.n1867 9.3005
R12103 gnd.n5245 gnd.n1868 9.3005
R12104 gnd.n5246 gnd.n1866 9.3005
R12105 gnd.n5248 gnd.n5247 9.3005
R12106 gnd.n5249 gnd.n1847 9.3005
R12107 gnd.n5272 gnd.n1848 9.3005
R12108 gnd.n5273 gnd.n1843 9.3005
R12109 gnd.n5276 gnd.n1844 9.3005
R12110 gnd.n5277 gnd.n1845 9.3005
R12111 gnd.n5286 gnd.n5285 9.3005
R12112 gnd.n5283 gnd.n1846 9.3005
R12113 gnd.n5282 gnd.n1802 9.3005
R12114 gnd.n5281 gnd.n1803 9.3005
R12115 gnd.n5278 gnd.n1804 9.3005
R12116 gnd.n1805 gnd.n1776 9.3005
R12117 gnd.n5354 gnd.n1777 9.3005
R12118 gnd.n5355 gnd.n1766 9.3005
R12119 gnd.n5357 gnd.n1767 9.3005
R12120 gnd.n5356 gnd.n1768 9.3005
R12121 gnd.n1769 gnd.n1741 9.3005
R12122 gnd.n5405 gnd.n1742 9.3005
R12123 gnd.n5406 gnd.n1740 9.3005
R12124 gnd.n5409 gnd.n5408 9.3005
R12125 gnd.n5410 gnd.n1672 9.3005
R12126 gnd.n5754 gnd.n1671 9.3005
R12127 gnd.n5756 gnd.n5755 9.3005
R12128 gnd.n5757 gnd.n1652 9.3005
R12129 gnd.n5866 gnd.n1650 9.3005
R12130 gnd.n5868 gnd.n5867 9.3005
R12131 gnd.n5092 gnd.n1986 9.3005
R12132 gnd.n4973 gnd.n4972 9.3005
R12133 gnd.n4975 gnd.n4874 9.3005
R12134 gnd.n4976 gnd.n4873 9.3005
R12135 gnd.n4979 gnd.n4872 9.3005
R12136 gnd.n4980 gnd.n4871 9.3005
R12137 gnd.n4983 gnd.n4870 9.3005
R12138 gnd.n4984 gnd.n4869 9.3005
R12139 gnd.n4987 gnd.n4868 9.3005
R12140 gnd.n4988 gnd.n4867 9.3005
R12141 gnd.n4991 gnd.n4866 9.3005
R12142 gnd.n4992 gnd.n4865 9.3005
R12143 gnd.n4995 gnd.n4864 9.3005
R12144 gnd.n4996 gnd.n4863 9.3005
R12145 gnd.n4999 gnd.n4862 9.3005
R12146 gnd.n5000 gnd.n4861 9.3005
R12147 gnd.n5003 gnd.n4860 9.3005
R12148 gnd.n5004 gnd.n4859 9.3005
R12149 gnd.n5007 gnd.n4858 9.3005
R12150 gnd.n5008 gnd.n4857 9.3005
R12151 gnd.n5011 gnd.n4856 9.3005
R12152 gnd.n5015 gnd.n4852 9.3005
R12153 gnd.n5016 gnd.n4851 9.3005
R12154 gnd.n5019 gnd.n4850 9.3005
R12155 gnd.n5020 gnd.n4849 9.3005
R12156 gnd.n5023 gnd.n4848 9.3005
R12157 gnd.n5024 gnd.n4847 9.3005
R12158 gnd.n5027 gnd.n4846 9.3005
R12159 gnd.n5028 gnd.n4845 9.3005
R12160 gnd.n5031 gnd.n4844 9.3005
R12161 gnd.n5032 gnd.n4843 9.3005
R12162 gnd.n5035 gnd.n4842 9.3005
R12163 gnd.n5036 gnd.n4841 9.3005
R12164 gnd.n5039 gnd.n4840 9.3005
R12165 gnd.n5040 gnd.n4839 9.3005
R12166 gnd.n5043 gnd.n4838 9.3005
R12167 gnd.n5044 gnd.n4837 9.3005
R12168 gnd.n5047 gnd.n4836 9.3005
R12169 gnd.n5048 gnd.n4835 9.3005
R12170 gnd.n5051 gnd.n4834 9.3005
R12171 gnd.n5053 gnd.n4831 9.3005
R12172 gnd.n5056 gnd.n4830 9.3005
R12173 gnd.n5057 gnd.n4829 9.3005
R12174 gnd.n5060 gnd.n4828 9.3005
R12175 gnd.n5061 gnd.n4827 9.3005
R12176 gnd.n5064 gnd.n4826 9.3005
R12177 gnd.n5065 gnd.n4825 9.3005
R12178 gnd.n5068 gnd.n4824 9.3005
R12179 gnd.n5069 gnd.n4823 9.3005
R12180 gnd.n5072 gnd.n4822 9.3005
R12181 gnd.n5073 gnd.n4821 9.3005
R12182 gnd.n5076 gnd.n4820 9.3005
R12183 gnd.n5077 gnd.n4819 9.3005
R12184 gnd.n5080 gnd.n4818 9.3005
R12185 gnd.n5082 gnd.n4817 9.3005
R12186 gnd.n5083 gnd.n4816 9.3005
R12187 gnd.n5084 gnd.n4815 9.3005
R12188 gnd.n5085 gnd.n4814 9.3005
R12189 gnd.n5012 gnd.n4853 9.3005
R12190 gnd.n4971 gnd.n1990 9.3005
R12191 gnd.n5101 gnd.n5100 9.3005
R12192 gnd.n5102 gnd.n1975 9.3005
R12193 gnd.n5104 gnd.n5103 9.3005
R12194 gnd.n1958 gnd.n1957 9.3005
R12195 gnd.n5121 gnd.n5120 9.3005
R12196 gnd.n5122 gnd.n1956 9.3005
R12197 gnd.n5124 gnd.n5123 9.3005
R12198 gnd.n1941 gnd.n1940 9.3005
R12199 gnd.n5141 gnd.n5140 9.3005
R12200 gnd.n5142 gnd.n1939 9.3005
R12201 gnd.n5144 gnd.n5143 9.3005
R12202 gnd.n1921 gnd.n1920 9.3005
R12203 gnd.n5165 gnd.n5164 9.3005
R12204 gnd.n5166 gnd.n1919 9.3005
R12205 gnd.n5170 gnd.n5167 9.3005
R12206 gnd.n5169 gnd.n5168 9.3005
R12207 gnd.n1896 gnd.n1895 9.3005
R12208 gnd.n5200 gnd.n5199 9.3005
R12209 gnd.n5201 gnd.n1894 9.3005
R12210 gnd.n5205 gnd.n5202 9.3005
R12211 gnd.n5204 gnd.n1828 9.3005
R12212 gnd.n5297 gnd.n1827 9.3005
R12213 gnd.n5301 gnd.n5298 9.3005
R12214 gnd.n5300 gnd.n5299 9.3005
R12215 gnd.n1793 gnd.n1792 9.3005
R12216 gnd.n5336 gnd.n5335 9.3005
R12217 gnd.n5337 gnd.n1791 9.3005
R12218 gnd.n5341 gnd.n5338 9.3005
R12219 gnd.n5340 gnd.n5339 9.3005
R12220 gnd.n1758 gnd.n1757 9.3005
R12221 gnd.n5384 gnd.n5383 9.3005
R12222 gnd.n5385 gnd.n1756 9.3005
R12223 gnd.n5389 gnd.n5386 9.3005
R12224 gnd.n5388 gnd.n5387 9.3005
R12225 gnd.n1731 gnd.n1730 9.3005
R12226 gnd.n5418 gnd.n5417 9.3005
R12227 gnd.n5419 gnd.n1729 9.3005
R12228 gnd.n5421 gnd.n5420 9.3005
R12229 gnd.n1662 gnd.n1661 9.3005
R12230 gnd.n5765 gnd.n5764 9.3005
R12231 gnd.n5766 gnd.n1660 9.3005
R12232 gnd.n5862 gnd.n5767 9.3005
R12233 gnd.n5861 gnd.n5860 9.3005
R12234 gnd.n1977 gnd.n1976 9.3005
R12235 gnd.n5296 gnd.n1833 9.3005
R12236 gnd.n5296 gnd.n5295 9.3005
R12237 gnd.n2079 gnd.n2078 9.3005
R12238 gnd.n2077 gnd.n1812 9.3005
R12239 gnd.n1810 gnd.n1809 9.3005
R12240 gnd.n5318 gnd.n5317 9.3005
R12241 gnd.n5319 gnd.n1808 9.3005
R12242 gnd.n5323 gnd.n5320 9.3005
R12243 gnd.n5322 gnd.n5321 9.3005
R12244 gnd.n1774 gnd.n1773 9.3005
R12245 gnd.n5363 gnd.n5362 9.3005
R12246 gnd.n5364 gnd.n1772 9.3005
R12247 gnd.n5371 gnd.n5365 9.3005
R12248 gnd.n5370 gnd.n5366 9.3005
R12249 gnd.n5369 gnd.n5367 9.3005
R12250 gnd.n1724 gnd.n1723 9.3005
R12251 gnd.n5427 gnd.n5426 9.3005
R12252 gnd.n5428 gnd.n1722 9.3005
R12253 gnd.n5430 gnd.n5429 9.3005
R12254 gnd.n1720 gnd.n1719 9.3005
R12255 gnd.n5435 gnd.n5434 9.3005
R12256 gnd.n5436 gnd.n1718 9.3005
R12257 gnd.n5593 gnd.n5437 9.3005
R12258 gnd.n5592 gnd.n5438 9.3005
R12259 gnd.n5591 gnd.n5439 9.3005
R12260 gnd.n5442 gnd.n5440 9.3005
R12261 gnd.n5585 gnd.n5443 9.3005
R12262 gnd.n5584 gnd.n5444 9.3005
R12263 gnd.n5583 gnd.n5445 9.3005
R12264 gnd.n5495 gnd.n5446 9.3005
R12265 gnd.n5497 gnd.n5496 9.3005
R12266 gnd.n5516 gnd.n5515 9.3005
R12267 gnd.n5517 gnd.n5494 9.3005
R12268 gnd.n5519 gnd.n5518 9.3005
R12269 gnd.n5482 gnd.n5481 9.3005
R12270 gnd.n5535 gnd.n5534 9.3005
R12271 gnd.n5536 gnd.n5480 9.3005
R12272 gnd.n5540 gnd.n5537 9.3005
R12273 gnd.n5539 gnd.n5538 9.3005
R12274 gnd.n1463 gnd.n1462 9.3005
R12275 gnd.n6015 gnd.n6014 9.3005
R12276 gnd.n6016 gnd.n1461 9.3005
R12277 gnd.n6018 gnd.n6017 9.3005
R12278 gnd.n1433 gnd.n1432 9.3005
R12279 gnd.n6075 gnd.n6074 9.3005
R12280 gnd.n6076 gnd.n1431 9.3005
R12281 gnd.n6078 gnd.n6077 9.3005
R12282 gnd.n1406 gnd.n1405 9.3005
R12283 gnd.n6117 gnd.n6116 9.3005
R12284 gnd.n6118 gnd.n1404 9.3005
R12285 gnd.n6128 gnd.n6119 9.3005
R12286 gnd.n6127 gnd.n6120 9.3005
R12287 gnd.n6126 gnd.n6121 9.3005
R12288 gnd.n6123 gnd.n6122 9.3005
R12289 gnd.n1362 gnd.n1361 9.3005
R12290 gnd.n6188 gnd.n6187 9.3005
R12291 gnd.n6189 gnd.n1360 9.3005
R12292 gnd.n6191 gnd.n6190 9.3005
R12293 gnd.n1331 gnd.n1330 9.3005
R12294 gnd.n6239 gnd.n6238 9.3005
R12295 gnd.n6240 gnd.n1329 9.3005
R12296 gnd.n6242 gnd.n6241 9.3005
R12297 gnd.n1327 gnd.n1326 9.3005
R12298 gnd.n6250 gnd.n6249 9.3005
R12299 gnd.n6251 gnd.n1325 9.3005
R12300 gnd.n6253 gnd.n6252 9.3005
R12301 gnd.n1268 gnd.n1267 9.3005
R12302 gnd.n6385 gnd.n6384 9.3005
R12303 gnd.n6386 gnd.n1266 9.3005
R12304 gnd.n6388 gnd.n6387 9.3005
R12305 gnd.n1244 gnd.n1243 9.3005
R12306 gnd.n6412 gnd.n6411 9.3005
R12307 gnd.n6413 gnd.n1242 9.3005
R12308 gnd.n6417 gnd.n6414 9.3005
R12309 gnd.n6416 gnd.n6415 9.3005
R12310 gnd.n1212 gnd.n1211 9.3005
R12311 gnd.n6449 gnd.n6448 9.3005
R12312 gnd.n6450 gnd.n1210 9.3005
R12313 gnd.n6452 gnd.n6451 9.3005
R12314 gnd.n1189 gnd.n1188 9.3005
R12315 gnd.n6483 gnd.n6482 9.3005
R12316 gnd.n6484 gnd.n1187 9.3005
R12317 gnd.n6502 gnd.n6485 9.3005
R12318 gnd.n6501 gnd.n6486 9.3005
R12319 gnd.n6500 gnd.n6487 9.3005
R12320 gnd.n6490 gnd.n6488 9.3005
R12321 gnd.n6494 gnd.n6491 9.3005
R12322 gnd.n6493 gnd.n6492 9.3005
R12323 gnd.n1130 gnd.n1129 9.3005
R12324 gnd.n6604 gnd.n6603 9.3005
R12325 gnd.n6605 gnd.n1128 9.3005
R12326 gnd.n6614 gnd.n6606 9.3005
R12327 gnd.n6613 gnd.n6607 9.3005
R12328 gnd.n6612 gnd.n6608 9.3005
R12329 gnd.n1091 gnd.n1090 9.3005
R12330 gnd.n6696 gnd.n6695 9.3005
R12331 gnd.n6697 gnd.n1089 9.3005
R12332 gnd.n6699 gnd.n6698 9.3005
R12333 gnd.n1068 gnd.n1067 9.3005
R12334 gnd.n6724 gnd.n6723 9.3005
R12335 gnd.n6725 gnd.n1066 9.3005
R12336 gnd.n6736 gnd.n6726 9.3005
R12337 gnd.n6735 gnd.n6727 9.3005
R12338 gnd.n6734 gnd.n6728 9.3005
R12339 gnd.n6730 gnd.n6729 9.3005
R12340 gnd.n1025 gnd.n1024 9.3005
R12341 gnd.n6807 gnd.n6806 9.3005
R12342 gnd.n6808 gnd.n1023 9.3005
R12343 gnd.n6810 gnd.n6809 9.3005
R12344 gnd.n997 gnd.n996 9.3005
R12345 gnd.n6848 gnd.n6847 9.3005
R12346 gnd.n6849 gnd.n995 9.3005
R12347 gnd.n6863 gnd.n6850 9.3005
R12348 gnd.n6862 gnd.n6851 9.3005
R12349 gnd.n6861 gnd.n6852 9.3005
R12350 gnd.n6854 gnd.n6853 9.3005
R12351 gnd.n6856 gnd.n6855 9.3005
R12352 gnd.n715 gnd.n714 9.3005
R12353 gnd.n7026 gnd.n7025 9.3005
R12354 gnd.n7027 gnd.n713 9.3005
R12355 gnd.n7031 gnd.n7028 9.3005
R12356 gnd.n7030 gnd.n7029 9.3005
R12357 gnd.n690 gnd.n689 9.3005
R12358 gnd.n7061 gnd.n7060 9.3005
R12359 gnd.n7062 gnd.n688 9.3005
R12360 gnd.n7067 gnd.n7063 9.3005
R12361 gnd.n7066 gnd.n7065 9.3005
R12362 gnd.n7064 gnd.n676 9.3005
R12363 gnd.n674 gnd.n673 9.3005
R12364 gnd.n7085 gnd.n7084 9.3005
R12365 gnd.n7086 gnd.n672 9.3005
R12366 gnd.n7121 gnd.n7087 9.3005
R12367 gnd.n7120 gnd.n7088 9.3005
R12368 gnd.n7119 gnd.n7089 9.3005
R12369 gnd.n7100 gnd.n7090 9.3005
R12370 gnd.n7115 gnd.n7101 9.3005
R12371 gnd.n7114 gnd.n7102 9.3005
R12372 gnd.n7113 gnd.n7103 9.3005
R12373 gnd.n7105 gnd.n7104 9.3005
R12374 gnd.n7109 gnd.n7106 9.3005
R12375 gnd.n7108 gnd.n7107 9.3005
R12376 gnd.n481 gnd.n480 9.3005
R12377 gnd.n7265 gnd.n7264 9.3005
R12378 gnd.n7266 gnd.n479 9.3005
R12379 gnd.n7270 gnd.n7267 9.3005
R12380 gnd.n7269 gnd.n7268 9.3005
R12381 gnd.n447 gnd.n446 9.3005
R12382 gnd.n7311 gnd.n7310 9.3005
R12383 gnd.n7312 gnd.n445 9.3005
R12384 gnd.n7316 gnd.n7313 9.3005
R12385 gnd.n7315 gnd.n7314 9.3005
R12386 gnd.n412 gnd.n411 9.3005
R12387 gnd.n7357 gnd.n7356 9.3005
R12388 gnd.n7358 gnd.n410 9.3005
R12389 gnd.n7362 gnd.n7359 9.3005
R12390 gnd.n7361 gnd.n7360 9.3005
R12391 gnd.n2080 gnd.n2076 9.3005
R12392 gnd.n3375 gnd.n3372 9.3005
R12393 gnd.n3371 gnd.n2083 9.3005
R12394 gnd.n3370 gnd.n3369 9.3005
R12395 gnd.n2085 gnd.n2084 9.3005
R12396 gnd.n3363 gnd.n3362 9.3005
R12397 gnd.n3361 gnd.n2089 9.3005
R12398 gnd.n3360 gnd.n3359 9.3005
R12399 gnd.n2091 gnd.n2090 9.3005
R12400 gnd.n3353 gnd.n3352 9.3005
R12401 gnd.n3351 gnd.n2095 9.3005
R12402 gnd.n3350 gnd.n3349 9.3005
R12403 gnd.n2097 gnd.n2096 9.3005
R12404 gnd.n3343 gnd.n3342 9.3005
R12405 gnd.n3341 gnd.n2101 9.3005
R12406 gnd.n3340 gnd.n3339 9.3005
R12407 gnd.n2103 gnd.n2102 9.3005
R12408 gnd.n3333 gnd.n3332 9.3005
R12409 gnd.n3331 gnd.n2107 9.3005
R12410 gnd.n3330 gnd.n3329 9.3005
R12411 gnd.n2109 gnd.n2108 9.3005
R12412 gnd.n3323 gnd.n3322 9.3005
R12413 gnd.n3321 gnd.n2113 9.3005
R12414 gnd.n3320 gnd.n3319 9.3005
R12415 gnd.n2115 gnd.n2114 9.3005
R12416 gnd.n3313 gnd.n3312 9.3005
R12417 gnd.n3311 gnd.n2119 9.3005
R12418 gnd.n3310 gnd.n3309 9.3005
R12419 gnd.n2121 gnd.n2120 9.3005
R12420 gnd.n3303 gnd.n3302 9.3005
R12421 gnd.n3301 gnd.n2125 9.3005
R12422 gnd.n3300 gnd.n3299 9.3005
R12423 gnd.n2127 gnd.n2126 9.3005
R12424 gnd.n3293 gnd.n3292 9.3005
R12425 gnd.n3291 gnd.n2131 9.3005
R12426 gnd.n3290 gnd.n3289 9.3005
R12427 gnd.n2133 gnd.n2132 9.3005
R12428 gnd.n3283 gnd.n3282 9.3005
R12429 gnd.n3281 gnd.n2137 9.3005
R12430 gnd.n3280 gnd.n3279 9.3005
R12431 gnd.n2139 gnd.n2138 9.3005
R12432 gnd.n3273 gnd.n3272 9.3005
R12433 gnd.n3271 gnd.n2143 9.3005
R12434 gnd.n3270 gnd.n3269 9.3005
R12435 gnd.n2145 gnd.n2144 9.3005
R12436 gnd.n3263 gnd.n3262 9.3005
R12437 gnd.n3261 gnd.n2149 9.3005
R12438 gnd.n3260 gnd.n3259 9.3005
R12439 gnd.n2151 gnd.n2150 9.3005
R12440 gnd.n3253 gnd.n3252 9.3005
R12441 gnd.n3251 gnd.n2155 9.3005
R12442 gnd.n3250 gnd.n3249 9.3005
R12443 gnd.n2157 gnd.n2156 9.3005
R12444 gnd.n3243 gnd.n3242 9.3005
R12445 gnd.n3241 gnd.n2161 9.3005
R12446 gnd.n3240 gnd.n3239 9.3005
R12447 gnd.n2163 gnd.n2162 9.3005
R12448 gnd.n3233 gnd.n3232 9.3005
R12449 gnd.n3231 gnd.n2167 9.3005
R12450 gnd.n3230 gnd.n3229 9.3005
R12451 gnd.n2169 gnd.n2168 9.3005
R12452 gnd.n3223 gnd.n3222 9.3005
R12453 gnd.n3221 gnd.n2173 9.3005
R12454 gnd.n3220 gnd.n3219 9.3005
R12455 gnd.n2175 gnd.n2174 9.3005
R12456 gnd.n3213 gnd.n3212 9.3005
R12457 gnd.n3211 gnd.n2179 9.3005
R12458 gnd.n3210 gnd.n3209 9.3005
R12459 gnd.n2181 gnd.n2180 9.3005
R12460 gnd.n3203 gnd.n3202 9.3005
R12461 gnd.n3201 gnd.n2185 9.3005
R12462 gnd.n3200 gnd.n3199 9.3005
R12463 gnd.n2187 gnd.n2186 9.3005
R12464 gnd.n3193 gnd.n3192 9.3005
R12465 gnd.n3191 gnd.n2191 9.3005
R12466 gnd.n3190 gnd.n3189 9.3005
R12467 gnd.n2193 gnd.n2192 9.3005
R12468 gnd.n3183 gnd.n3182 9.3005
R12469 gnd.n3181 gnd.n2197 9.3005
R12470 gnd.n3180 gnd.n3179 9.3005
R12471 gnd.n2199 gnd.n2198 9.3005
R12472 gnd.n3173 gnd.n3172 9.3005
R12473 gnd.n3171 gnd.n2203 9.3005
R12474 gnd.n3170 gnd.n3169 9.3005
R12475 gnd.n2205 gnd.n2204 9.3005
R12476 gnd.n3374 gnd.n3373 9.3005
R12477 gnd.n7190 gnd.n7189 9.3005
R12478 gnd.n5506 gnd.n5505 9.3005
R12479 gnd.n5507 gnd.n5502 9.3005
R12480 gnd.n5509 gnd.n5508 9.3005
R12481 gnd.n5487 gnd.n5486 9.3005
R12482 gnd.n5525 gnd.n5524 9.3005
R12483 gnd.n5526 gnd.n5485 9.3005
R12484 gnd.n5528 gnd.n5527 9.3005
R12485 gnd.n5474 gnd.n5473 9.3005
R12486 gnd.n5546 gnd.n5545 9.3005
R12487 gnd.n5547 gnd.n5471 9.3005
R12488 gnd.n5556 gnd.n5555 9.3005
R12489 gnd.n5554 gnd.n5472 9.3005
R12490 gnd.n5553 gnd.n5552 9.3005
R12491 gnd.n5551 gnd.n5548 9.3005
R12492 gnd.n5550 gnd.n5549 9.3005
R12493 gnd.n1450 gnd.n1449 9.3005
R12494 gnd.n6034 gnd.n6033 9.3005
R12495 gnd.n6035 gnd.n1447 9.3005
R12496 gnd.n6044 gnd.n6043 9.3005
R12497 gnd.n6042 gnd.n1448 9.3005
R12498 gnd.n6041 gnd.n6040 9.3005
R12499 gnd.n6039 gnd.n6037 9.3005
R12500 gnd.n6036 gnd.n1391 9.3005
R12501 gnd.n6141 gnd.n1390 9.3005
R12502 gnd.n6143 gnd.n6142 9.3005
R12503 gnd.n6144 gnd.n1388 9.3005
R12504 gnd.n6150 gnd.n6149 9.3005
R12505 gnd.n6148 gnd.n1389 9.3005
R12506 gnd.n6147 gnd.n6146 9.3005
R12507 gnd.n1354 gnd.n1353 9.3005
R12508 gnd.n6211 gnd.n6210 9.3005
R12509 gnd.n6212 gnd.n1351 9.3005
R12510 gnd.n6215 gnd.n6214 9.3005
R12511 gnd.n6213 gnd.n1352 9.3005
R12512 gnd.n1298 gnd.n1297 9.3005
R12513 gnd.n6290 gnd.n6289 9.3005
R12514 gnd.n6291 gnd.n1296 9.3005
R12515 gnd.n6294 gnd.n6293 9.3005
R12516 gnd.n6292 gnd.n1294 9.3005
R12517 gnd.n6298 gnd.n1293 9.3005
R12518 gnd.n6300 gnd.n6299 9.3005
R12519 gnd.n6301 gnd.n1292 9.3005
R12520 gnd.n6303 gnd.n6302 9.3005
R12521 gnd.n6304 gnd.n1290 9.3005
R12522 gnd.n6308 gnd.n6307 9.3005
R12523 gnd.n6309 gnd.n1288 9.3005
R12524 gnd.n6342 gnd.n6341 9.3005
R12525 gnd.n6340 gnd.n1289 9.3005
R12526 gnd.n6339 gnd.n6338 9.3005
R12527 gnd.n6337 gnd.n6310 9.3005
R12528 gnd.n6336 gnd.n6335 9.3005
R12529 gnd.n6334 gnd.n6313 9.3005
R12530 gnd.n6333 gnd.n6332 9.3005
R12531 gnd.n6331 gnd.n6314 9.3005
R12532 gnd.n6330 gnd.n6329 9.3005
R12533 gnd.n6328 gnd.n6325 9.3005
R12534 gnd.n6327 gnd.n6326 9.3005
R12535 gnd.n1154 gnd.n1153 9.3005
R12536 gnd.n6541 gnd.n6540 9.3005
R12537 gnd.n6542 gnd.n1151 9.3005
R12538 gnd.n6558 gnd.n6557 9.3005
R12539 gnd.n6556 gnd.n1152 9.3005
R12540 gnd.n6555 gnd.n6554 9.3005
R12541 gnd.n6553 gnd.n6543 9.3005
R12542 gnd.n6552 gnd.n6551 9.3005
R12543 gnd.n6550 gnd.n6548 9.3005
R12544 gnd.n6549 gnd.n1106 9.3005
R12545 gnd.n6642 gnd.n1105 9.3005
R12546 gnd.n6644 gnd.n6643 9.3005
R12547 gnd.n6645 gnd.n1104 9.3005
R12548 gnd.n6647 gnd.n6646 9.3005
R12549 gnd.n6649 gnd.n1101 9.3005
R12550 gnd.n6651 gnd.n6650 9.3005
R12551 gnd.n6652 gnd.n1099 9.3005
R12552 gnd.n6670 gnd.n6669 9.3005
R12553 gnd.n6668 gnd.n1100 9.3005
R12554 gnd.n6667 gnd.n6666 9.3005
R12555 gnd.n6665 gnd.n6653 9.3005
R12556 gnd.n6664 gnd.n6663 9.3005
R12557 gnd.n6662 gnd.n6660 9.3005
R12558 gnd.n6661 gnd.n1012 9.3005
R12559 gnd.n6825 gnd.n1011 9.3005
R12560 gnd.n6827 gnd.n6826 9.3005
R12561 gnd.n6828 gnd.n1009 9.3005
R12562 gnd.n6833 gnd.n6832 9.3005
R12563 gnd.n6831 gnd.n1010 9.3005
R12564 gnd.n6830 gnd.n6829 9.3005
R12565 gnd.n722 gnd.n721 9.3005
R12566 gnd.n7016 gnd.n7015 9.3005
R12567 gnd.n7017 gnd.n719 9.3005
R12568 gnd.n7020 gnd.n7019 9.3005
R12569 gnd.n7018 gnd.n720 9.3005
R12570 gnd.n697 gnd.n696 9.3005
R12571 gnd.n7046 gnd.n7045 9.3005
R12572 gnd.n7047 gnd.n694 9.3005
R12573 gnd.n7055 gnd.n7054 9.3005
R12574 gnd.n7053 gnd.n695 9.3005
R12575 gnd.n7052 gnd.n7051 9.3005
R12576 gnd.n7050 gnd.n7048 9.3005
R12577 gnd.n582 gnd.n581 9.3005
R12578 gnd.n7188 gnd.n7187 9.3005
R12579 gnd.n5504 gnd.n5503 9.3005
R12580 gnd.n5739 gnd.n1683 9.3005
R12581 gnd.n1855 gnd.n1854 9.3005
R12582 gnd.n5264 gnd.n5263 9.3005
R12583 gnd.n5265 gnd.n1852 9.3005
R12584 gnd.n5268 gnd.n5267 9.3005
R12585 gnd.n5266 gnd.n1853 9.3005
R12586 gnd.n1819 gnd.n1818 9.3005
R12587 gnd.n5306 gnd.n5305 9.3005
R12588 gnd.n5307 gnd.n1816 9.3005
R12589 gnd.n5310 gnd.n5309 9.3005
R12590 gnd.n5308 gnd.n1817 9.3005
R12591 gnd.n1784 gnd.n1783 9.3005
R12592 gnd.n5346 gnd.n5345 9.3005
R12593 gnd.n5347 gnd.n1781 9.3005
R12594 gnd.n5350 gnd.n5349 9.3005
R12595 gnd.n5348 gnd.n1782 9.3005
R12596 gnd.n1749 gnd.n1748 9.3005
R12597 gnd.n5394 gnd.n5393 9.3005
R12598 gnd.n5395 gnd.n1746 9.3005
R12599 gnd.n5401 gnd.n5400 9.3005
R12600 gnd.n5399 gnd.n1747 9.3005
R12601 gnd.n5398 gnd.n5397 9.3005
R12602 gnd.n1678 gnd.n1676 9.3005
R12603 gnd.n5750 gnd.n5749 9.3005
R12604 gnd.n5748 gnd.n1677 9.3005
R12605 gnd.n5747 gnd.n5746 9.3005
R12606 gnd.n5745 gnd.n1679 9.3005
R12607 gnd.n5744 gnd.n5743 9.3005
R12608 gnd.n5717 gnd.n5716 9.3005
R12609 gnd.n5601 gnd.n5600 9.3005
R12610 gnd.n5711 gnd.n5710 9.3005
R12611 gnd.n5709 gnd.n5708 9.3005
R12612 gnd.n5615 gnd.n5614 9.3005
R12613 gnd.n5703 gnd.n5702 9.3005
R12614 gnd.n5701 gnd.n5700 9.3005
R12615 gnd.n5627 gnd.n5626 9.3005
R12616 gnd.n5695 gnd.n5694 9.3005
R12617 gnd.n5693 gnd.n5692 9.3005
R12618 gnd.n5638 gnd.n5637 9.3005
R12619 gnd.n5687 gnd.n5686 9.3005
R12620 gnd.n5685 gnd.n5684 9.3005
R12621 gnd.n5650 gnd.n5649 9.3005
R12622 gnd.n5679 gnd.n5678 9.3005
R12623 gnd.n5677 gnd.n5676 9.3005
R12624 gnd.n5668 gnd.n5666 9.3005
R12625 gnd.n5665 gnd.n1684 9.3005
R12626 gnd.n5719 gnd.n5718 9.3005
R12627 gnd.n5741 gnd.n5740 9.3005
R12628 gnd.n5667 gnd.n1685 9.3005
R12629 gnd.n5675 gnd.n5674 9.3005
R12630 gnd.n5654 gnd.n5653 9.3005
R12631 gnd.n5681 gnd.n5680 9.3005
R12632 gnd.n5683 gnd.n5682 9.3005
R12633 gnd.n5644 gnd.n5643 9.3005
R12634 gnd.n5689 gnd.n5688 9.3005
R12635 gnd.n5691 gnd.n5690 9.3005
R12636 gnd.n5631 gnd.n5630 9.3005
R12637 gnd.n5697 gnd.n5696 9.3005
R12638 gnd.n5699 gnd.n5698 9.3005
R12639 gnd.n5621 gnd.n5620 9.3005
R12640 gnd.n5705 gnd.n5704 9.3005
R12641 gnd.n5707 gnd.n5706 9.3005
R12642 gnd.n5608 gnd.n5607 9.3005
R12643 gnd.n5713 gnd.n5712 9.3005
R12644 gnd.n5715 gnd.n5714 9.3005
R12645 gnd.n5604 gnd.n1715 9.3005
R12646 gnd.n5720 gnd.n1714 9.3005
R12647 gnd.n5722 gnd.n5721 9.3005
R12648 gnd.n5724 gnd.n5723 9.3005
R12649 gnd.n5726 gnd.n5725 9.3005
R12650 gnd.n5727 gnd.n1708 9.3005
R12651 gnd.n5729 gnd.n5728 9.3005
R12652 gnd.n5730 gnd.n1707 9.3005
R12653 gnd.n5732 gnd.n5731 9.3005
R12654 gnd.n5733 gnd.n1706 9.3005
R12655 gnd.n5578 gnd.n5577 9.3005
R12656 gnd.n5576 gnd.n5454 9.3005
R12657 gnd.n5575 gnd.n5574 9.3005
R12658 gnd.n5573 gnd.n5456 9.3005
R12659 gnd.n5572 gnd.n5571 9.3005
R12660 gnd.n5570 gnd.n5460 9.3005
R12661 gnd.n5569 gnd.n5568 9.3005
R12662 gnd.n5567 gnd.n5461 9.3005
R12663 gnd.n5566 gnd.n5565 9.3005
R12664 gnd.n5564 gnd.n5465 9.3005
R12665 gnd.n5563 gnd.n5562 9.3005
R12666 gnd.n5561 gnd.n5466 9.3005
R12667 gnd.n1456 gnd.n1455 9.3005
R12668 gnd.n6025 gnd.n6024 9.3005
R12669 gnd.n6026 gnd.n1454 9.3005
R12670 gnd.n6028 gnd.n6027 9.3005
R12671 gnd.n1425 gnd.n1424 9.3005
R12672 gnd.n6084 gnd.n6083 9.3005
R12673 gnd.n6085 gnd.n1423 9.3005
R12674 gnd.n6087 gnd.n6086 9.3005
R12675 gnd.n1397 gnd.n1396 9.3005
R12676 gnd.n6134 gnd.n6133 9.3005
R12677 gnd.n6135 gnd.n1395 9.3005
R12678 gnd.n6137 gnd.n6136 9.3005
R12679 gnd.n1370 gnd.n1369 9.3005
R12680 gnd.n6179 gnd.n6178 9.3005
R12681 gnd.n6180 gnd.n1368 9.3005
R12682 gnd.n6182 gnd.n6181 9.3005
R12683 gnd.n1339 gnd.n1338 9.3005
R12684 gnd.n6230 gnd.n6229 9.3005
R12685 gnd.n6231 gnd.n1337 9.3005
R12686 gnd.n6233 gnd.n6232 9.3005
R12687 gnd.n1306 gnd.n1305 9.3005
R12688 gnd.n6275 gnd.n6274 9.3005
R12689 gnd.n6276 gnd.n1303 9.3005
R12690 gnd.n6285 gnd.n6284 9.3005
R12691 gnd.n6283 gnd.n1304 9.3005
R12692 gnd.n6282 gnd.n6281 9.3005
R12693 gnd.n6280 gnd.n6277 9.3005
R12694 gnd.n1260 gnd.n1259 9.3005
R12695 gnd.n6394 gnd.n6393 9.3005
R12696 gnd.n6395 gnd.n1257 9.3005
R12697 gnd.n6398 gnd.n6397 9.3005
R12698 gnd.n6396 gnd.n1258 9.3005
R12699 gnd.n1229 gnd.n1228 9.3005
R12700 gnd.n6430 gnd.n6429 9.3005
R12701 gnd.n6431 gnd.n1226 9.3005
R12702 gnd.n6434 gnd.n6433 9.3005
R12703 gnd.n6432 gnd.n1227 9.3005
R12704 gnd.n1204 gnd.n1203 9.3005
R12705 gnd.n6459 gnd.n6458 9.3005
R12706 gnd.n6460 gnd.n1202 9.3005
R12707 gnd.n6462 gnd.n6461 9.3005
R12708 gnd.n1174 gnd.n1173 9.3005
R12709 gnd.n6516 gnd.n6515 9.3005
R12710 gnd.n6517 gnd.n1171 9.3005
R12711 gnd.n6520 gnd.n6519 9.3005
R12712 gnd.n6518 gnd.n1172 9.3005
R12713 gnd.n1139 gnd.n1138 9.3005
R12714 gnd.n6582 gnd.n6581 9.3005
R12715 gnd.n6583 gnd.n1136 9.3005
R12716 gnd.n6598 gnd.n6597 9.3005
R12717 gnd.n6596 gnd.n1137 9.3005
R12718 gnd.n6595 gnd.n6594 9.3005
R12719 gnd.n6593 gnd.n6584 9.3005
R12720 gnd.n6592 gnd.n6591 9.3005
R12721 gnd.n6590 gnd.n6589 9.3005
R12722 gnd.n1083 gnd.n1082 9.3005
R12723 gnd.n6705 gnd.n6704 9.3005
R12724 gnd.n6706 gnd.n1080 9.3005
R12725 gnd.n6709 gnd.n6708 9.3005
R12726 gnd.n6707 gnd.n1081 9.3005
R12727 gnd.n1053 gnd.n1052 9.3005
R12728 gnd.n6750 gnd.n6749 9.3005
R12729 gnd.n6751 gnd.n1050 9.3005
R12730 gnd.n6754 gnd.n6753 9.3005
R12731 gnd.n6752 gnd.n1051 9.3005
R12732 gnd.n1034 gnd.n1032 9.3005
R12733 gnd.n6801 gnd.n6800 9.3005
R12734 gnd.n6799 gnd.n1033 9.3005
R12735 gnd.n6798 gnd.n6797 9.3005
R12736 gnd.n1006 gnd.n1004 9.3005
R12737 gnd.n6842 gnd.n6841 9.3005
R12738 gnd.n6840 gnd.n1005 9.3005
R12739 gnd.n6839 gnd.n6838 9.3005
R12740 gnd.n732 gnd.n731 9.3005
R12741 gnd.n7007 gnd.n7006 9.3005
R12742 gnd.n7008 gnd.n729 9.3005
R12743 gnd.n7011 gnd.n7010 9.3005
R12744 gnd.n7009 gnd.n730 9.3005
R12745 gnd.n706 gnd.n705 9.3005
R12746 gnd.n7037 gnd.n7036 9.3005
R12747 gnd.n7038 gnd.n703 9.3005
R12748 gnd.n7041 gnd.n7040 9.3005
R12749 gnd.n7039 gnd.n704 9.3005
R12750 gnd.n682 gnd.n681 9.3005
R12751 gnd.n7073 gnd.n7072 9.3005
R12752 gnd.n7074 gnd.n680 9.3005
R12753 gnd.n7076 gnd.n7075 9.3005
R12754 gnd.n589 gnd.n588 9.3005
R12755 gnd.n7183 gnd.n7182 9.3005
R12756 gnd.n5455 gnd.n5453 9.3005
R12757 gnd.n7179 gnd.n590 9.3005
R12758 gnd.n7178 gnd.n7177 9.3005
R12759 gnd.n7176 gnd.n593 9.3005
R12760 gnd.n7175 gnd.n7174 9.3005
R12761 gnd.n7173 gnd.n594 9.3005
R12762 gnd.n7172 gnd.n7171 9.3005
R12763 gnd.n7181 gnd.n7180 9.3005
R12764 gnd.n7200 gnd.n7199 9.3005
R12765 gnd.n645 gnd.n568 9.3005
R12766 gnd.n7130 gnd.n7129 9.3005
R12767 gnd.n7132 gnd.n7131 9.3005
R12768 gnd.n638 gnd.n637 9.3005
R12769 gnd.n7138 gnd.n7137 9.3005
R12770 gnd.n7140 gnd.n7139 9.3005
R12771 gnd.n628 gnd.n627 9.3005
R12772 gnd.n7146 gnd.n7145 9.3005
R12773 gnd.n7148 gnd.n7147 9.3005
R12774 gnd.n620 gnd.n619 9.3005
R12775 gnd.n7154 gnd.n7153 9.3005
R12776 gnd.n7156 gnd.n7155 9.3005
R12777 gnd.n610 gnd.n609 9.3005
R12778 gnd.n7162 gnd.n7161 9.3005
R12779 gnd.n7164 gnd.n7163 9.3005
R12780 gnd.n606 gnd.n600 9.3005
R12781 gnd.n573 gnd.n571 9.3005
R12782 gnd.n7194 gnd.n7193 9.3005
R12783 gnd.n7169 gnd.n598 9.3005
R12784 gnd.n7168 gnd.n7167 9.3005
R12785 gnd.n7166 gnd.n7165 9.3005
R12786 gnd.n604 gnd.n603 9.3005
R12787 gnd.n7160 gnd.n7159 9.3005
R12788 gnd.n7158 gnd.n7157 9.3005
R12789 gnd.n614 gnd.n613 9.3005
R12790 gnd.n7152 gnd.n7151 9.3005
R12791 gnd.n7150 gnd.n7149 9.3005
R12792 gnd.n624 gnd.n623 9.3005
R12793 gnd.n7144 gnd.n7143 9.3005
R12794 gnd.n7142 gnd.n7141 9.3005
R12795 gnd.n632 gnd.n631 9.3005
R12796 gnd.n7136 gnd.n7135 9.3005
R12797 gnd.n7134 gnd.n7133 9.3005
R12798 gnd.n642 gnd.n641 9.3005
R12799 gnd.n7128 gnd.n7127 9.3005
R12800 gnd.n7126 gnd.n572 9.3005
R12801 gnd.n7198 gnd.n7197 9.3005
R12802 gnd.n7196 gnd.n7195 9.3005
R12803 gnd.n7192 gnd.n7191 9.3005
R12804 gnd.n7218 gnd.n516 9.3005
R12805 gnd.n7221 gnd.n7220 9.3005
R12806 gnd.n7219 gnd.n517 9.3005
R12807 gnd.n489 gnd.n488 9.3005
R12808 gnd.n7254 gnd.n7253 9.3005
R12809 gnd.n7255 gnd.n486 9.3005
R12810 gnd.n7258 gnd.n7257 9.3005
R12811 gnd.n7256 gnd.n487 9.3005
R12812 gnd.n455 gnd.n454 9.3005
R12813 gnd.n7300 gnd.n7299 9.3005
R12814 gnd.n7301 gnd.n452 9.3005
R12815 gnd.n7304 gnd.n7303 9.3005
R12816 gnd.n7302 gnd.n453 9.3005
R12817 gnd.n420 gnd.n419 9.3005
R12818 gnd.n7347 gnd.n7346 9.3005
R12819 gnd.n7348 gnd.n417 9.3005
R12820 gnd.n7351 gnd.n7350 9.3005
R12821 gnd.n7349 gnd.n418 9.3005
R12822 gnd.n388 gnd.n387 9.3005
R12823 gnd.n7391 gnd.n7390 9.3005
R12824 gnd.n7392 gnd.n385 9.3005
R12825 gnd.n7400 gnd.n7399 9.3005
R12826 gnd.n7398 gnd.n386 9.3005
R12827 gnd.n7397 gnd.n7396 9.3005
R12828 gnd.n7395 gnd.n7393 9.3005
R12829 gnd.n85 gnd.n83 9.3005
R12830 gnd.n7217 gnd.n7216 9.3005
R12831 gnd.t35 gnd.n3487 9.24152
R12832 gnd.n3389 gnd.t169 9.24152
R12833 gnd.n4673 gnd.t144 9.24152
R12834 gnd.t85 gnd.n1971 9.24152
R12835 gnd.n1680 gnd.t121 9.24152
R12836 gnd.n6227 gnd.t353 9.24152
R12837 gnd.n6711 gnd.t7 9.24152
R12838 gnd.n7223 gnd.t78 9.24152
R12839 gnd.n7685 gnd.t96 9.24152
R12840 gnd.t43 gnd.t35 8.92286
R12841 gnd.n1468 gnd.n1458 8.92286
R12842 gnd.n6207 gnd.n1343 8.92286
R12843 gnd.n1322 gnd.n1300 8.92286
R12844 gnd.n6437 gnd.n1222 8.92286
R12845 gnd.n6465 gnd.n1182 8.92286
R12846 gnd.n6624 gnd.n1116 8.92286
R12847 gnd.n6714 gnd.n6713 8.92286
R12848 gnd.n6822 gnd.n1014 8.92286
R12849 gnd.n7003 gnd.n737 8.92286
R12850 gnd.n4643 gnd.n4618 8.92171
R12851 gnd.n4611 gnd.n4586 8.92171
R12852 gnd.n4579 gnd.n4554 8.92171
R12853 gnd.n4548 gnd.n4523 8.92171
R12854 gnd.n4516 gnd.n4491 8.92171
R12855 gnd.n4484 gnd.n4459 8.92171
R12856 gnd.n4452 gnd.n4427 8.92171
R12857 gnd.n4421 gnd.n4396 8.92171
R12858 gnd.n759 gnd.n741 8.72777
R12859 gnd.n4147 gnd.t21 8.60421
R12860 gnd.t125 gnd.n5451 8.60421
R12861 gnd.t57 gnd.n1493 8.60421
R12862 gnd.n6001 gnd.n1493 8.60421
R12863 gnd.t68 gnd.n1214 8.60421
R12864 gnd.n6479 gnd.t357 8.60421
R12865 gnd.n725 gnd.t18 8.60421
R12866 gnd.n7080 gnd.t89 8.60421
R12867 gnd.n3559 gnd.n3543 8.43656
R12868 gnd.n50 gnd.n34 8.43656
R12869 gnd.n6012 gnd.t154 8.28555
R12870 gnd.n6167 gnd.n1358 8.28555
R12871 gnd.n6372 gnd.n1277 8.28555
R12872 gnd.n6427 gnd.n1231 8.28555
R12873 gnd.n6513 gnd.n6512 8.28555
R12874 gnd.n6569 gnd.n1122 8.28555
R12875 gnd.n6680 gnd.n1071 8.28555
R12876 gnd.t157 gnd.n6844 8.28555
R12877 gnd.n4644 gnd.n4616 8.14595
R12878 gnd.n4612 gnd.n4584 8.14595
R12879 gnd.n4580 gnd.n4552 8.14595
R12880 gnd.n4549 gnd.n4521 8.14595
R12881 gnd.n4517 gnd.n4489 8.14595
R12882 gnd.n4485 gnd.n4457 8.14595
R12883 gnd.n4453 gnd.n4425 8.14595
R12884 gnd.n4422 gnd.n4394 8.14595
R12885 gnd.n5216 gnd.n0 8.10675
R12886 gnd.n7759 gnd.n7758 8.10675
R12887 gnd.n4649 gnd.n4648 7.97301
R12888 gnd.t41 gnd.n3662 7.9669
R12889 gnd.n5736 gnd.n1702 7.9669
R12890 gnd.t2 gnd.n6159 7.9669
R12891 gnd.n6757 gnd.t52 7.9669
R12892 gnd.n7124 gnd.n647 7.9669
R12893 gnd.n7759 gnd.n82 7.86902
R12894 gnd.n7193 gnd.n571 7.75808
R12895 gnd.n5666 gnd.n5665 7.75808
R12896 gnd.n7535 gnd.n348 7.75808
R12897 gnd.n4931 gnd.n4895 7.75808
R12898 gnd.t154 gnd.n6011 7.64824
R12899 gnd.n6053 gnd.t182 7.64824
R12900 gnd.n6096 gnd.n6095 7.64824
R12901 gnd.n6167 gnd.t10 7.64824
R12902 gnd.n1254 gnd.t42 7.64824
R12903 gnd.n6409 gnd.t42 7.64824
R12904 gnd.n6497 gnd.t51 7.64824
R12905 gnd.n6530 gnd.t51 7.64824
R12906 gnd.n6680 gnd.t31 7.64824
R12907 gnd.n6776 gnd.n6775 7.64824
R12908 gnd.n6845 gnd.t157 7.64824
R12909 gnd.n3592 gnd.n3591 7.53171
R12910 gnd.n4056 gnd.t23 7.32958
R12911 gnd.n5500 gnd.t125 7.32958
R12912 gnd.n5558 gnd.t57 7.32958
R12913 gnd.n6001 gnd.n1465 7.32958
R12914 gnd.n7013 gnd.n726 7.32958
R12915 gnd.t18 gnd.n717 7.32958
R12916 gnd.t89 gnd.n7078 7.32958
R12917 gnd.n1489 gnd.n1488 7.30353
R12918 gnd.n758 gnd.n757 7.30353
R12919 gnd.n4016 gnd.n3735 7.01093
R12920 gnd.n3738 gnd.n3736 7.01093
R12921 gnd.n4026 gnd.n4025 7.01093
R12922 gnd.n4037 gnd.n3719 7.01093
R12923 gnd.n4036 gnd.n3722 7.01093
R12924 gnd.n4047 gnd.n3710 7.01093
R12925 gnd.n3713 gnd.n3711 7.01093
R12926 gnd.n4057 gnd.n4056 7.01093
R12927 gnd.n4067 gnd.n3691 7.01093
R12928 gnd.n4066 gnd.n3694 7.01093
R12929 gnd.n4075 gnd.n3685 7.01093
R12930 gnd.n4087 gnd.n3675 7.01093
R12931 gnd.n4097 gnd.n3660 7.01093
R12932 gnd.n4113 gnd.n4112 7.01093
R12933 gnd.n3662 gnd.n3599 7.01093
R12934 gnd.n4167 gnd.n3600 7.01093
R12935 gnd.n4161 gnd.n4160 7.01093
R12936 gnd.n3649 gnd.n3611 7.01093
R12937 gnd.n4153 gnd.n3622 7.01093
R12938 gnd.n3640 gnd.n3635 7.01093
R12939 gnd.n4147 gnd.n4146 7.01093
R12940 gnd.n4193 gnd.n3522 7.01093
R12941 gnd.n4192 gnd.n4191 7.01093
R12942 gnd.n4204 gnd.n4203 7.01093
R12943 gnd.n3515 gnd.n3507 7.01093
R12944 gnd.n4233 gnd.n3495 7.01093
R12945 gnd.n4232 gnd.n3498 7.01093
R12946 gnd.n4243 gnd.n3487 7.01093
R12947 gnd.n3488 gnd.n3476 7.01093
R12948 gnd.n4254 gnd.n3477 7.01093
R12949 gnd.n4278 gnd.n3468 7.01093
R12950 gnd.n4277 gnd.n3459 7.01093
R12951 gnd.n4300 gnd.n4299 7.01093
R12952 gnd.n4318 gnd.n3440 7.01093
R12953 gnd.n4317 gnd.n3443 7.01093
R12954 gnd.n4328 gnd.n3432 7.01093
R12955 gnd.n3433 gnd.n3420 7.01093
R12956 gnd.n4339 gnd.n3421 7.01093
R12957 gnd.n4366 gnd.n3405 7.01093
R12958 gnd.n4378 gnd.n4377 7.01093
R12959 gnd.n4360 gnd.n3398 7.01093
R12960 gnd.n4389 gnd.n4388 7.01093
R12961 gnd.n4661 gnd.n3386 7.01093
R12962 gnd.n4660 gnd.n3389 7.01093
R12963 gnd.n4673 gnd.n2073 7.01093
R12964 gnd.n4683 gnd.n1992 7.01093
R12965 gnd.n6022 gnd.n1458 7.01093
R12966 gnd.n6047 gnd.n6046 7.01093
R12967 gnd.n6287 gnd.n1300 7.01093
R12968 gnd.n6419 gnd.t24 7.01093
R12969 gnd.n6437 gnd.n6436 7.01093
R12970 gnd.n6465 gnd.n6464 7.01093
R12971 gnd.n6315 gnd.t64 7.01093
R12972 gnd.n6624 gnd.n1117 7.01093
R12973 gnd.n6823 gnd.n6822 7.01093
R12974 gnd.n7004 gnd.n7003 7.01093
R12975 gnd.t118 gnd.n737 7.01093
R12976 gnd.n3694 gnd.t364 6.69227
R12977 gnd.n3498 gnd.t43 6.69227
R12978 gnd.n4367 gnd.t359 6.69227
R12979 gnd.n5138 gnd.t229 6.69227
R12980 gnd.n6193 gnd.t353 6.69227
R12981 gnd.n6721 gnd.t7 6.69227
R12982 gnd.n7514 gnd.t220 6.69227
R12983 gnd.n6933 gnd.n6932 6.5566
R12984 gnd.n5939 gnd.n5938 6.5566
R12985 gnd.n1584 gnd.n1530 6.5566
R12986 gnd.n6947 gnd.n6946 6.5566
R12987 gnd.n6105 gnd.n6104 6.37362
R12988 gnd.n6153 gnd.n1387 6.37362
R12989 gnd.n6364 gnd.n6363 6.37362
R12990 gnd.n6561 gnd.n1150 6.37362
R12991 gnd.n6746 gnd.n1058 6.37362
R12992 gnd.n6656 gnd.n6655 6.37362
R12993 gnd.n5674 gnd.n5671 6.20656
R12994 gnd.n7197 gnd.n576 6.20656
R12995 gnd.t351 gnd.n4123 6.05496
R12996 gnd.n4124 gnd.t32 6.05496
R12997 gnd.t49 gnd.n3522 6.05496
R12998 gnd.t70 gnd.n4288 6.05496
R12999 gnd.n5182 gnd.t239 6.05496
R13000 gnd.n133 gnd.t197 6.05496
R13001 gnd.n4646 gnd.n4616 5.81868
R13002 gnd.n4614 gnd.n4584 5.81868
R13003 gnd.n4582 gnd.n4552 5.81868
R13004 gnd.n4551 gnd.n4521 5.81868
R13005 gnd.n4519 gnd.n4489 5.81868
R13006 gnd.n4487 gnd.n4457 5.81868
R13007 gnd.n4455 gnd.n4425 5.81868
R13008 gnd.n4424 gnd.n4394 5.81868
R13009 gnd.n6054 gnd.n1436 5.73631
R13010 gnd.n6047 gnd.t82 5.73631
R13011 gnd.t38 gnd.n6207 5.73631
R13012 gnd.n6218 gnd.n6217 5.73631
R13013 gnd.n6272 gnd.n6271 5.73631
R13014 gnd.t26 gnd.n1262 5.73631
R13015 gnd.n6436 gnd.t25 5.73631
R13016 gnd.n6455 gnd.n1206 5.73631
R13017 gnd.n6473 gnd.n1196 5.73631
R13018 gnd.n6464 gnd.t27 5.73631
R13019 gnd.n6578 gnd.t11 5.73631
R13020 gnd.n6632 gnd.n1093 5.73631
R13021 gnd.n6640 gnd.n6639 5.73631
R13022 gnd.n6714 gnd.t55 5.73631
R13023 gnd.n6786 gnd.n6785 5.73631
R13024 gnd.n6879 gnd.t118 5.73631
R13025 gnd.n6940 gnd.n786 5.62001
R13026 gnd.n5934 gnd.n5931 5.62001
R13027 gnd.n5931 gnd.n1588 5.62001
R13028 gnd.n6941 gnd.n6940 5.62001
R13029 gnd.n3875 gnd.n3870 5.4308
R13030 gnd.n4691 gnd.n2059 5.4308
R13031 gnd.n4191 gnd.t30 5.41765
R13032 gnd.t59 gnd.n4214 5.41765
R13033 gnd.t370 gnd.n3452 5.41765
R13034 gnd.n5242 gnd.t272 5.41765
R13035 gnd.n5261 gnd.t224 5.41765
R13036 gnd.n6246 gnd.t62 5.41765
R13037 gnd.t14 gnd.n6631 5.41765
R13038 gnd.n7419 gnd.t233 5.41765
R13039 gnd.n7753 gnd.t207 5.41765
R13040 gnd.n6161 gnd.n1379 5.09899
R13041 gnd.n6159 gnd.n1372 5.09899
R13042 gnd.t67 gnd.n6371 5.09899
R13043 gnd.n6390 gnd.n1264 5.09899
R13044 gnd.n6402 gnd.n6401 5.09899
R13045 gnd.n6495 gnd.n1156 5.09899
R13046 gnd.n6537 gnd.n1141 5.09899
R13047 gnd.n6570 gnd.t6 5.09899
R13048 gnd.n6757 gnd.n1044 5.09899
R13049 gnd.n6731 gnd.n1047 5.09899
R13050 gnd.n4644 gnd.n4643 5.04292
R13051 gnd.n4612 gnd.n4611 5.04292
R13052 gnd.n4580 gnd.n4579 5.04292
R13053 gnd.n4549 gnd.n4548 5.04292
R13054 gnd.n4517 gnd.n4516 5.04292
R13055 gnd.n4485 gnd.n4484 5.04292
R13056 gnd.n4453 gnd.n4452 5.04292
R13057 gnd.n4422 gnd.n4421 5.04292
R13058 gnd.n4154 gnd.t40 4.78034
R13059 gnd.n3477 gnd.t39 4.78034
R13060 gnd.n3378 gnd.n2066 4.78034
R13061 gnd.n5207 gnd.t201 4.78034
R13062 gnd.n5303 gnd.t213 4.78034
R13063 gnd.n6030 gnd.t60 4.78034
R13064 gnd.n6271 gnd.t62 4.78034
R13065 gnd.n6632 gnd.t14 4.78034
R13066 gnd.n6836 gnd.t374 4.78034
R13067 gnd.n726 gnd.t93 4.78034
R13068 gnd.n7388 gnd.t259 4.78034
R13069 gnd.n7739 gnd.t231 4.78034
R13070 gnd.n3596 gnd.n3593 4.74817
R13071 gnd.n3646 gnd.n3528 4.74817
R13072 gnd.n3633 gnd.n3527 4.74817
R13073 gnd.n3526 gnd.n3525 4.74817
R13074 gnd.n3642 gnd.n3593 4.74817
R13075 gnd.n3643 gnd.n3528 4.74817
R13076 gnd.n3645 gnd.n3527 4.74817
R13077 gnd.n3632 gnd.n3526 4.74817
R13078 gnd.n7384 gnd.n101 4.74817
R13079 gnd.n7415 gnd.n99 4.74817
R13080 gnd.n7751 gnd.n94 4.74817
R13081 gnd.n7749 gnd.n95 4.74817
R13082 gnd.n375 gnd.n101 4.74817
R13083 gnd.n7417 gnd.n99 4.74817
R13084 gnd.n7414 gnd.n94 4.74817
R13085 gnd.n7750 gnd.n7749 4.74817
R13086 gnd.n5203 gnd.n1834 4.74817
R13087 gnd.n1860 gnd.n1832 4.74817
R13088 gnd.n5259 gnd.n1831 4.74817
R13089 gnd.n1835 gnd.n1830 4.74817
R13090 gnd.n1874 gnd.n1834 4.74817
R13091 gnd.n5240 gnd.n1832 4.74817
R13092 gnd.n1861 gnd.n1831 4.74817
R13093 gnd.n5258 gnd.n1830 4.74817
R13094 gnd.n3591 gnd.n3590 4.74296
R13095 gnd.n82 gnd.n81 4.74296
R13096 gnd.n3559 gnd.n3558 4.7074
R13097 gnd.n3575 gnd.n3574 4.7074
R13098 gnd.n50 gnd.n49 4.7074
R13099 gnd.n66 gnd.n65 4.7074
R13100 gnd.n3591 gnd.n3575 4.65959
R13101 gnd.n82 gnd.n66 4.65959
R13102 gnd.n959 gnd.n861 4.6132
R13103 gnd.n5929 gnd.n5928 4.6132
R13104 gnd.n6061 gnd.n1441 4.46168
R13105 gnd.n6081 gnd.n1427 4.46168
R13106 gnd.n6096 gnd.t36 4.46168
R13107 gnd.n6235 gnd.n1335 4.46168
R13108 gnd.n6245 gnd.n6244 4.46168
R13109 gnd.n6445 gnd.n6444 4.46168
R13110 gnd.n6471 gnd.n1191 4.46168
R13111 gnd.n6630 gnd.n1112 4.46168
R13112 gnd.n6702 gnd.n1085 4.46168
R13113 gnd.n6776 gnd.t37 4.46168
R13114 gnd.n6844 gnd.n1001 4.46168
R13115 gnd.n6871 gnd.n988 4.46168
R13116 gnd.n754 gnd.n741 4.46111
R13117 gnd.n4629 gnd.n4625 4.38594
R13118 gnd.n4597 gnd.n4593 4.38594
R13119 gnd.n4565 gnd.n4561 4.38594
R13120 gnd.n4534 gnd.n4530 4.38594
R13121 gnd.n4502 gnd.n4498 4.38594
R13122 gnd.n4470 gnd.n4466 4.38594
R13123 gnd.n4438 gnd.n4434 4.38594
R13124 gnd.n4407 gnd.n4403 4.38594
R13125 gnd.n4640 gnd.n4618 4.26717
R13126 gnd.n4608 gnd.n4586 4.26717
R13127 gnd.n4576 gnd.n4554 4.26717
R13128 gnd.n4545 gnd.n4523 4.26717
R13129 gnd.n4513 gnd.n4491 4.26717
R13130 gnd.n4481 gnd.n4459 4.26717
R13131 gnd.n4449 gnd.n4427 4.26717
R13132 gnd.n4418 gnd.n4396 4.26717
R13133 gnd.n4098 gnd.t360 4.14303
R13134 gnd.n4328 gnd.t20 4.14303
R13135 gnd.t203 gnd.n1923 4.14303
R13136 gnd.n5381 gnd.t195 4.14303
R13137 gnd.n5373 gnd.t274 4.14303
R13138 gnd.t4 gnd.n6408 4.14303
R13139 gnd.t367 gnd.n1168 4.14303
R13140 gnd.n7272 gnd.t222 4.14303
R13141 gnd.t236 gnd.n7306 4.14303
R13142 gnd.n7715 gnd.t277 4.14303
R13143 gnd.n4648 gnd.n4647 4.08274
R13144 gnd.n6932 gnd.n6931 4.05904
R13145 gnd.n5940 gnd.n5939 4.05904
R13146 gnd.n1581 gnd.n1530 4.05904
R13147 gnd.n6948 gnd.n6947 4.05904
R13148 gnd.n19 gnd.n9 3.99943
R13149 gnd.n5588 gnd.n1597 3.82437
R13150 gnd.t182 gnd.n1427 3.82437
R13151 gnd.t36 gnd.n1409 3.82437
R13152 gnd.n6130 gnd.n1401 3.82437
R13153 gnd.n6185 gnd.n1364 3.82437
R13154 gnd.n6287 gnd.t28 3.82437
R13155 gnd.n6382 gnd.n6381 3.82437
R13156 gnd.n6353 gnd.n6352 3.82437
R13157 gnd.n6523 gnd.n1165 3.82437
R13158 gnd.n6601 gnd.n1132 3.82437
R13159 gnd.t12 gnd.n1117 3.82437
R13160 gnd.n6738 gnd.n1055 3.82437
R13161 gnd.n6804 gnd.n1027 3.82437
R13162 gnd.t37 gnd.n1020 3.82437
R13163 gnd.t93 gnd.n725 3.82437
R13164 gnd.n7203 gnd.n529 3.82437
R13165 gnd.n4171 gnd.n3592 3.81325
R13166 gnd.n3575 gnd.n3559 3.72967
R13167 gnd.n66 gnd.n50 3.72967
R13168 gnd.n4648 gnd.n4520 3.70378
R13169 gnd.n19 gnd.n18 3.60163
R13170 gnd.n5293 gnd.n1839 3.50571
R13171 gnd.t255 gnd.n1795 3.50571
R13172 gnd.n5490 gnd.t47 3.50571
R13173 gnd.t355 gnd.n700 3.50571
R13174 gnd.n7354 gnd.t191 3.50571
R13175 gnd.n7402 gnd.n383 3.50571
R13176 gnd.n4639 gnd.n4620 3.49141
R13177 gnd.n4607 gnd.n4588 3.49141
R13178 gnd.n4575 gnd.n4556 3.49141
R13179 gnd.n4544 gnd.n4525 3.49141
R13180 gnd.n4512 gnd.n4493 3.49141
R13181 gnd.n4480 gnd.n4461 3.49141
R13182 gnd.n4448 gnd.n4429 3.49141
R13183 gnd.n4417 gnd.n4398 3.49141
R13184 gnd.n839 gnd.n794 3.29747
R13185 gnd.n842 gnd.n794 3.29747
R13186 gnd.n7644 gnd.n7641 3.29747
R13187 gnd.n7645 gnd.n7644 3.29747
R13188 gnd.n5053 gnd.n5052 3.29747
R13189 gnd.n5052 gnd.n5051 3.29747
R13190 gnd.n5800 gnd.n5795 3.29747
R13191 gnd.n5825 gnd.n5800 3.29747
R13192 gnd.n6011 gnd.n6010 3.18706
R13193 gnd.t82 gnd.n1420 3.18706
R13194 gnd.n6090 gnd.n6089 3.18706
R13195 gnd.n6227 gnd.n6226 3.18706
R13196 gnd.n6259 gnd.n6256 3.18706
R13197 gnd.n6345 gnd.n6344 3.18706
R13198 gnd.n6506 gnd.n6505 3.18706
R13199 gnd.n1125 gnd.n1124 3.18706
R13200 gnd.n6712 gnd.n6711 3.18706
R13201 gnd.n6795 gnd.n6794 3.18706
R13202 gnd.n6865 gnd.t132 3.18706
R13203 gnd.n6879 gnd.n6878 3.18706
R13204 gnd.n3677 gnd.t360 2.8684
R13205 gnd.n6160 gnd.t2 2.8684
R13206 gnd.t52 gnd.n6756 2.8684
R13207 gnd.n3576 gnd.t196 2.82907
R13208 gnd.n3576 gnd.t350 2.82907
R13209 gnd.n3578 gnd.t256 2.82907
R13210 gnd.n3578 gnd.t339 2.82907
R13211 gnd.n3580 gnd.t206 2.82907
R13212 gnd.n3580 gnd.t318 2.82907
R13213 gnd.n3582 gnd.t342 2.82907
R13214 gnd.n3582 gnd.t253 2.82907
R13215 gnd.n3584 gnd.t285 2.82907
R13216 gnd.n3584 gnd.t264 2.82907
R13217 gnd.n3586 gnd.t263 2.82907
R13218 gnd.n3586 gnd.t240 2.82907
R13219 gnd.n3588 gnd.t270 2.82907
R13220 gnd.n3588 gnd.t306 2.82907
R13221 gnd.n3529 gnd.t300 2.82907
R13222 gnd.n3529 gnd.t315 2.82907
R13223 gnd.n3531 gnd.t327 2.82907
R13224 gnd.n3531 gnd.t343 2.82907
R13225 gnd.n3533 gnd.t294 2.82907
R13226 gnd.n3533 gnd.t304 2.82907
R13227 gnd.n3535 gnd.t316 2.82907
R13228 gnd.n3535 gnd.t225 2.82907
R13229 gnd.n3537 gnd.t303 2.82907
R13230 gnd.n3537 gnd.t194 2.82907
R13231 gnd.n3539 gnd.t333 2.82907
R13232 gnd.n3539 gnd.t328 2.82907
R13233 gnd.n3541 gnd.t247 2.82907
R13234 gnd.n3541 gnd.t310 2.82907
R13235 gnd.n3544 gnd.t287 2.82907
R13236 gnd.n3544 gnd.t275 2.82907
R13237 gnd.n3546 gnd.t276 2.82907
R13238 gnd.n3546 gnd.t299 2.82907
R13239 gnd.n3548 gnd.t251 2.82907
R13240 gnd.n3548 gnd.t288 2.82907
R13241 gnd.n3550 gnd.t289 2.82907
R13242 gnd.n3550 gnd.t266 2.82907
R13243 gnd.n3552 gnd.t202 2.82907
R13244 gnd.n3552 gnd.t252 2.82907
R13245 gnd.n3554 gnd.t242 2.82907
R13246 gnd.n3554 gnd.t291 2.82907
R13247 gnd.n3556 gnd.t230 2.82907
R13248 gnd.n3556 gnd.t204 2.82907
R13249 gnd.n3560 gnd.t332 2.82907
R13250 gnd.n3560 gnd.t293 2.82907
R13251 gnd.n3562 gnd.t309 2.82907
R13252 gnd.n3562 gnd.t268 2.82907
R13253 gnd.n3564 gnd.t296 2.82907
R13254 gnd.n3564 gnd.t214 2.82907
R13255 gnd.n3566 gnd.t273 2.82907
R13256 gnd.n3566 gnd.t307 2.82907
R13257 gnd.n3568 gnd.t325 2.82907
R13258 gnd.n3568 gnd.t311 2.82907
R13259 gnd.n3570 gnd.t312 2.82907
R13260 gnd.n3570 gnd.t302 2.82907
R13261 gnd.n3572 gnd.t317 2.82907
R13262 gnd.n3572 gnd.t347 2.82907
R13263 gnd.n79 gnd.t278 2.82907
R13264 gnd.n79 gnd.t321 2.82907
R13265 gnd.n77 gnd.t337 2.82907
R13266 gnd.n77 gnd.t346 2.82907
R13267 gnd.n75 gnd.t348 2.82907
R13268 gnd.n75 gnd.t249 2.82907
R13269 gnd.n73 gnd.t344 2.82907
R13270 gnd.n73 gnd.t313 2.82907
R13271 gnd.n71 gnd.t295 2.82907
R13272 gnd.n71 gnd.t335 2.82907
R13273 gnd.n69 gnd.t308 2.82907
R13274 gnd.n69 gnd.t345 2.82907
R13275 gnd.n67 gnd.t324 2.82907
R13276 gnd.n67 gnd.t237 2.82907
R13277 gnd.n32 gnd.t336 2.82907
R13278 gnd.n32 gnd.t228 2.82907
R13279 gnd.n30 gnd.t198 2.82907
R13280 gnd.n30 gnd.t217 2.82907
R13281 gnd.n28 gnd.t322 2.82907
R13282 gnd.n28 gnd.t297 2.82907
R13283 gnd.n26 gnd.t284 2.82907
R13284 gnd.n26 gnd.t341 2.82907
R13285 gnd.n24 gnd.t331 2.82907
R13286 gnd.n24 gnd.t269 2.82907
R13287 gnd.n22 gnd.t246 2.82907
R13288 gnd.n22 gnd.t192 2.82907
R13289 gnd.n20 gnd.t340 2.82907
R13290 gnd.n20 gnd.t323 2.82907
R13291 gnd.n47 gnd.t338 2.82907
R13292 gnd.n47 gnd.t245 2.82907
R13293 gnd.n45 gnd.t258 2.82907
R13294 gnd.n45 gnd.t212 2.82907
R13295 gnd.n43 gnd.t216 2.82907
R13296 gnd.n43 gnd.t232 2.82907
R13297 gnd.n41 gnd.t234 2.82907
R13298 gnd.n41 gnd.t257 2.82907
R13299 gnd.n39 gnd.t260 2.82907
R13300 gnd.n39 gnd.t281 2.82907
R13301 gnd.n37 gnd.t279 2.82907
R13302 gnd.n37 gnd.t238 2.82907
R13303 gnd.n35 gnd.t235 2.82907
R13304 gnd.n35 gnd.t254 2.82907
R13305 gnd.n63 gnd.t320 2.82907
R13306 gnd.n63 gnd.t221 2.82907
R13307 gnd.n61 gnd.t265 2.82907
R13308 gnd.n61 gnd.t286 2.82907
R13309 gnd.n59 gnd.t290 2.82907
R13310 gnd.n59 gnd.t305 2.82907
R13311 gnd.n57 gnd.t282 2.82907
R13312 gnd.n57 gnd.t208 2.82907
R13313 gnd.n55 gnd.t329 2.82907
R13314 gnd.n55 gnd.t262 2.82907
R13315 gnd.n53 gnd.t200 2.82907
R13316 gnd.n53 gnd.t283 2.82907
R13317 gnd.n51 gnd.t223 2.82907
R13318 gnd.n51 gnd.t301 2.82907
R13319 gnd.n4636 gnd.n4635 2.71565
R13320 gnd.n4604 gnd.n4603 2.71565
R13321 gnd.n4572 gnd.n4571 2.71565
R13322 gnd.n4541 gnd.n4540 2.71565
R13323 gnd.n4509 gnd.n4508 2.71565
R13324 gnd.n4477 gnd.n4476 2.71565
R13325 gnd.n4445 gnd.n4444 2.71565
R13326 gnd.n4414 gnd.n4413 2.71565
R13327 gnd.n5303 gnd.n1821 2.54975
R13328 gnd.n1823 gnd.n1813 2.54975
R13329 gnd.n5313 gnd.n5312 2.54975
R13330 gnd.n5333 gnd.n1795 2.54975
R13331 gnd.n5279 gnd.n1798 2.54975
R13332 gnd.n5343 gnd.n1786 2.54975
R13333 gnd.n5326 gnd.n5325 2.54975
R13334 gnd.n5352 gnd.n1779 2.54975
R13335 gnd.n5381 gnd.n1760 2.54975
R13336 gnd.n5360 gnd.n5359 2.54975
R13337 gnd.n5391 gnd.n1751 2.54975
R13338 gnd.n5374 gnd.n5373 2.54975
R13339 gnd.n5403 gnd.n1744 2.54975
R13340 gnd.n5415 gnd.n1733 2.54975
R13341 gnd.n1736 gnd.n1726 2.54975
R13342 gnd.n5424 gnd.n5423 2.54975
R13343 gnd.n5752 gnd.n1674 2.54975
R13344 gnd.n5762 gnd.n1664 2.54975
R13345 gnd.n1680 gnd.n1667 2.54975
R13346 gnd.n5864 gnd.n1654 2.54975
R13347 gnd.n5596 gnd.n1656 2.54975
R13348 gnd.n6030 gnd.t100 2.54975
R13349 gnd.n6114 gnd.n6113 2.54975
R13350 gnd.n6104 gnd.t369 2.54975
R13351 gnd.n6194 gnd.n6193 2.54975
R13352 gnd.t13 gnd.n1308 2.54975
R13353 gnd.n6255 gnd.n1323 2.54975
R13354 gnd.n6372 gnd.t67 2.54975
R13355 gnd.n6426 gnd.n1234 2.54975
R13356 gnd.n6504 gnd.n1176 2.54975
R13357 gnd.t6 gnd.n6569 2.54975
R13358 gnd.n6617 gnd.n6616 2.54975
R13359 gnd.n6693 gnd.t54 2.54975
R13360 gnd.n6721 gnd.n6720 2.54975
R13361 gnd.n6655 gnd.t29 2.54975
R13362 gnd.n6813 gnd.n6812 2.54975
R13363 gnd.n7214 gnd.n522 2.54975
R13364 gnd.n7098 gnd.n7097 2.54975
R13365 gnd.n7223 gnd.n501 2.54975
R13366 gnd.n7241 gnd.n504 2.54975
R13367 gnd.n7227 gnd.n491 2.54975
R13368 gnd.n7251 gnd.n493 2.54975
R13369 gnd.n7261 gnd.n483 2.54975
R13370 gnd.n7260 gnd.n466 2.54975
R13371 gnd.n7287 gnd.n469 2.54975
R13372 gnd.n7273 gnd.n7272 2.54975
R13373 gnd.n7297 gnd.n458 2.54975
R13374 gnd.n7307 gnd.n449 2.54975
R13375 gnd.n7306 gnd.n431 2.54975
R13376 gnd.n7334 gnd.n434 2.54975
R13377 gnd.n7319 gnd.n7318 2.54975
R13378 gnd.n7344 gnd.n423 2.54975
R13379 gnd.n7327 gnd.n414 2.54975
R13380 gnd.n7354 gnd.n7353 2.54975
R13381 gnd.n7378 gnd.n401 2.54975
R13382 gnd.n7365 gnd.n7364 2.54975
R13383 gnd.n7388 gnd.n391 2.54975
R13384 gnd.n4171 gnd.n3593 2.27742
R13385 gnd.n4171 gnd.n3528 2.27742
R13386 gnd.n4171 gnd.n3527 2.27742
R13387 gnd.n4171 gnd.n3526 2.27742
R13388 gnd.n7748 gnd.n101 2.27742
R13389 gnd.n7748 gnd.n99 2.27742
R13390 gnd.n7748 gnd.n94 2.27742
R13391 gnd.n7749 gnd.n7748 2.27742
R13392 gnd.n5296 gnd.n1834 2.27742
R13393 gnd.n5296 gnd.n1832 2.27742
R13394 gnd.n5296 gnd.n1831 2.27742
R13395 gnd.n5296 gnd.n1830 2.27742
R13396 gnd.n4025 gnd.t114 2.23109
R13397 gnd.n3648 gnd.t40 2.23109
R13398 gnd.n3379 gnd.n3378 2.23109
R13399 gnd.n6409 gnd.t4 2.23109
R13400 gnd.n6497 gnd.t367 2.23109
R13401 gnd.n4632 gnd.n4622 1.93989
R13402 gnd.n4600 gnd.n4590 1.93989
R13403 gnd.n4568 gnd.n4558 1.93989
R13404 gnd.n4537 gnd.n4527 1.93989
R13405 gnd.n4505 gnd.n4495 1.93989
R13406 gnd.n4473 gnd.n4463 1.93989
R13407 gnd.n4441 gnd.n4431 1.93989
R13408 gnd.n4410 gnd.n4400 1.93989
R13409 gnd.n6131 gnd.n1399 1.91244
R13410 gnd.n6184 gnd.n1366 1.91244
R13411 gnd.n6420 gnd.n1238 1.91244
R13412 gnd.n6323 gnd.n6322 1.91244
R13413 gnd.n6740 gnd.n6739 1.91244
R13414 gnd.n6803 gnd.n1029 1.91244
R13415 gnd.t72 gnd.n988 1.91244
R13416 gnd.t33 gnd.n4036 1.59378
R13417 gnd.n4215 gnd.t59 1.59378
R13418 gnd.n3461 gnd.t370 1.59378
R13419 gnd.t45 gnd.n1270 1.59378
R13420 gnd.n6600 gnd.t16 1.59378
R13421 gnd.t75 gnd.n6021 1.27512
R13422 gnd.n6021 gnd.n6020 1.27512
R13423 gnd.n6080 gnd.n1429 1.27512
R13424 gnd.n6208 gnd.t38 1.27512
R13425 gnd.n6236 gnd.n1333 1.27512
R13426 gnd.n6265 gnd.n1316 1.27512
R13427 gnd.n6446 gnd.n1214 1.27512
R13428 gnd.n6480 gnd.n6479 1.27512
R13429 gnd.n6610 gnd.n6609 1.27512
R13430 gnd.n6701 gnd.n1087 1.27512
R13431 gnd.n1102 gnd.t55 1.27512
R13432 gnd.n6845 gnd.n999 1.27512
R13433 gnd.n6859 gnd.n734 1.27512
R13434 gnd.n3878 gnd.n3870 1.16414
R13435 gnd.n4694 gnd.n2059 1.16414
R13436 gnd.n4631 gnd.n4624 1.16414
R13437 gnd.n4599 gnd.n4592 1.16414
R13438 gnd.n4567 gnd.n4560 1.16414
R13439 gnd.n4536 gnd.n4529 1.16414
R13440 gnd.n4504 gnd.n4497 1.16414
R13441 gnd.n4472 gnd.n4465 1.16414
R13442 gnd.n4440 gnd.n4433 1.16414
R13443 gnd.n4409 gnd.n4402 1.16414
R13444 gnd.n959 gnd.n958 0.970197
R13445 gnd.n5929 gnd.n1589 0.970197
R13446 gnd.n4615 gnd.n4583 0.962709
R13447 gnd.n4647 gnd.n4615 0.962709
R13448 gnd.n4488 gnd.n4456 0.962709
R13449 gnd.n4520 gnd.n4488 0.962709
R13450 gnd.n4124 gnd.t351 0.956468
R13451 gnd.n4289 gnd.t70 0.956468
R13452 gnd.t60 gnd.n1452 0.956468
R13453 gnd.n6114 gnd.t0 0.956468
R13454 gnd.n6812 gnd.t65 0.956468
R13455 gnd.t374 gnd.n6835 0.956468
R13456 gnd.n2 gnd.n1 0.672012
R13457 gnd.n3 gnd.n2 0.672012
R13458 gnd.n4 gnd.n3 0.672012
R13459 gnd.n5 gnd.n4 0.672012
R13460 gnd.n6 gnd.n5 0.672012
R13461 gnd.n7 gnd.n6 0.672012
R13462 gnd.n8 gnd.n7 0.672012
R13463 gnd.n9 gnd.n8 0.672012
R13464 gnd.n11 gnd.n10 0.672012
R13465 gnd.n12 gnd.n11 0.672012
R13466 gnd.n13 gnd.n12 0.672012
R13467 gnd.n14 gnd.n13 0.672012
R13468 gnd.n15 gnd.n14 0.672012
R13469 gnd.n16 gnd.n15 0.672012
R13470 gnd.n17 gnd.n16 0.672012
R13471 gnd.n18 gnd.n17 0.672012
R13472 gnd gnd.n0 0.665707
R13473 gnd.n6072 gnd.t107 0.637812
R13474 gnd.n6139 gnd.n1393 0.637812
R13475 gnd.n6176 gnd.n6175 0.637812
R13476 gnd.n6175 gnd.t9 0.637812
R13477 gnd.n6391 gnd.n1262 0.637812
R13478 gnd.n6400 gnd.n1254 0.637812
R13479 gnd.t24 gnd.n1231 0.637812
R13480 gnd.n6512 gnd.t64 0.637812
R13481 gnd.n6530 gnd.n1160 0.637812
R13482 gnd.n6579 gnd.n6578 0.637812
R13483 gnd.n6673 gnd.t56 0.637812
R13484 gnd.n6673 gnd.n6672 0.637812
R13485 gnd.n6768 gnd.n1039 0.637812
R13486 gnd.n6865 gnd.t103 0.637812
R13487 gnd.n3590 gnd.n3589 0.573776
R13488 gnd.n3589 gnd.n3587 0.573776
R13489 gnd.n3587 gnd.n3585 0.573776
R13490 gnd.n3585 gnd.n3583 0.573776
R13491 gnd.n3583 gnd.n3581 0.573776
R13492 gnd.n3581 gnd.n3579 0.573776
R13493 gnd.n3579 gnd.n3577 0.573776
R13494 gnd.n3543 gnd.n3542 0.573776
R13495 gnd.n3542 gnd.n3540 0.573776
R13496 gnd.n3540 gnd.n3538 0.573776
R13497 gnd.n3538 gnd.n3536 0.573776
R13498 gnd.n3536 gnd.n3534 0.573776
R13499 gnd.n3534 gnd.n3532 0.573776
R13500 gnd.n3532 gnd.n3530 0.573776
R13501 gnd.n3558 gnd.n3557 0.573776
R13502 gnd.n3557 gnd.n3555 0.573776
R13503 gnd.n3555 gnd.n3553 0.573776
R13504 gnd.n3553 gnd.n3551 0.573776
R13505 gnd.n3551 gnd.n3549 0.573776
R13506 gnd.n3549 gnd.n3547 0.573776
R13507 gnd.n3547 gnd.n3545 0.573776
R13508 gnd.n3574 gnd.n3573 0.573776
R13509 gnd.n3573 gnd.n3571 0.573776
R13510 gnd.n3571 gnd.n3569 0.573776
R13511 gnd.n3569 gnd.n3567 0.573776
R13512 gnd.n3567 gnd.n3565 0.573776
R13513 gnd.n3565 gnd.n3563 0.573776
R13514 gnd.n3563 gnd.n3561 0.573776
R13515 gnd.n70 gnd.n68 0.573776
R13516 gnd.n72 gnd.n70 0.573776
R13517 gnd.n74 gnd.n72 0.573776
R13518 gnd.n76 gnd.n74 0.573776
R13519 gnd.n78 gnd.n76 0.573776
R13520 gnd.n80 gnd.n78 0.573776
R13521 gnd.n81 gnd.n80 0.573776
R13522 gnd.n23 gnd.n21 0.573776
R13523 gnd.n25 gnd.n23 0.573776
R13524 gnd.n27 gnd.n25 0.573776
R13525 gnd.n29 gnd.n27 0.573776
R13526 gnd.n31 gnd.n29 0.573776
R13527 gnd.n33 gnd.n31 0.573776
R13528 gnd.n34 gnd.n33 0.573776
R13529 gnd.n38 gnd.n36 0.573776
R13530 gnd.n40 gnd.n38 0.573776
R13531 gnd.n42 gnd.n40 0.573776
R13532 gnd.n44 gnd.n42 0.573776
R13533 gnd.n46 gnd.n44 0.573776
R13534 gnd.n48 gnd.n46 0.573776
R13535 gnd.n49 gnd.n48 0.573776
R13536 gnd.n54 gnd.n52 0.573776
R13537 gnd.n56 gnd.n54 0.573776
R13538 gnd.n58 gnd.n56 0.573776
R13539 gnd.n60 gnd.n58 0.573776
R13540 gnd.n62 gnd.n60 0.573776
R13541 gnd.n64 gnd.n62 0.573776
R13542 gnd.n65 gnd.n64 0.573776
R13543 gnd.n7760 gnd.n7759 0.553847
R13544 gnd.n7533 gnd.n7532 0.505073
R13545 gnd.n4932 gnd.n4930 0.505073
R13546 gnd.n4351 gnd.n2063 0.486781
R13547 gnd.n3927 gnd.n3926 0.48678
R13548 gnd.n4668 gnd.n2017 0.480683
R13549 gnd.n4011 gnd.n4010 0.480683
R13550 gnd.n7676 gnd.n7675 0.470012
R13551 gnd.n7209 gnd.n7208 0.470012
R13552 gnd.n5860 gnd.n5859 0.470012
R13553 gnd.n4814 gnd.n1976 0.470012
R13554 gnd.n3162 gnd.n2204 0.459342
R13555 gnd.n2519 gnd.n2513 0.459342
R13556 gnd.n7189 gnd.n7188 0.451719
R13557 gnd.n5503 gnd.n1683 0.451719
R13558 gnd.n5455 gnd.n1706 0.451719
R13559 gnd.n7182 gnd.n7181 0.451719
R13560 gnd.n7748 gnd.n98 0.421899
R13561 gnd.n5296 gnd.n1829 0.421899
R13562 gnd.n5671 gnd.n5653 0.388379
R13563 gnd.n4628 gnd.n4627 0.388379
R13564 gnd.n4596 gnd.n4595 0.388379
R13565 gnd.n4564 gnd.n4563 0.388379
R13566 gnd.n4533 gnd.n4532 0.388379
R13567 gnd.n4501 gnd.n4500 0.388379
R13568 gnd.n4469 gnd.n4468 0.388379
R13569 gnd.n4437 gnd.n4436 0.388379
R13570 gnd.n4406 gnd.n4405 0.388379
R13571 gnd.n7126 gnd.n576 0.388379
R13572 gnd.n7760 gnd.n19 0.374463
R13573 gnd gnd.n7760 0.367492
R13574 gnd.n3423 gnd.t359 0.319156
R13575 gnd.n6370 gnd.t45 0.319156
R13576 gnd.t25 gnd.t68 0.319156
R13577 gnd.t27 gnd.t357 0.319156
R13578 gnd.n6571 gnd.t16 0.319156
R13579 gnd.n3845 gnd.n3823 0.311721
R13580 gnd.n7566 gnd.n7565 0.293183
R13581 gnd.n4970 gnd.n4969 0.293183
R13582 gnd.n2076 gnd.n1829 0.276415
R13583 gnd.n7360 gnd.n98 0.276415
R13584 gnd.n5743 gnd.n5742 0.27489
R13585 gnd.n7217 gnd.n518 0.27489
R13586 gnd.n4739 gnd.n4738 0.268793
R13587 gnd.n7567 gnd.n7566 0.258122
R13588 gnd.n897 gnd.n599 0.258122
R13589 gnd.n5870 gnd.n5869 0.258122
R13590 gnd.n4971 gnd.n4970 0.258122
R13591 gnd.n4738 gnd.n4737 0.241354
R13592 gnd.n861 gnd.n860 0.229039
R13593 gnd.n862 gnd.n861 0.229039
R13594 gnd.n5928 gnd.n1592 0.229039
R13595 gnd.n5928 gnd.n5927 0.229039
R13596 gnd.n3999 gnd.n3798 0.206293
R13597 gnd.n2680 gnd.n98 0.183427
R13598 gnd.n3373 gnd.n1829 0.183427
R13599 gnd.n3592 gnd.n0 0.169152
R13600 gnd.n4645 gnd.n4617 0.155672
R13601 gnd.n4638 gnd.n4617 0.155672
R13602 gnd.n4638 gnd.n4637 0.155672
R13603 gnd.n4637 gnd.n4621 0.155672
R13604 gnd.n4630 gnd.n4621 0.155672
R13605 gnd.n4630 gnd.n4629 0.155672
R13606 gnd.n4613 gnd.n4585 0.155672
R13607 gnd.n4606 gnd.n4585 0.155672
R13608 gnd.n4606 gnd.n4605 0.155672
R13609 gnd.n4605 gnd.n4589 0.155672
R13610 gnd.n4598 gnd.n4589 0.155672
R13611 gnd.n4598 gnd.n4597 0.155672
R13612 gnd.n4581 gnd.n4553 0.155672
R13613 gnd.n4574 gnd.n4553 0.155672
R13614 gnd.n4574 gnd.n4573 0.155672
R13615 gnd.n4573 gnd.n4557 0.155672
R13616 gnd.n4566 gnd.n4557 0.155672
R13617 gnd.n4566 gnd.n4565 0.155672
R13618 gnd.n4550 gnd.n4522 0.155672
R13619 gnd.n4543 gnd.n4522 0.155672
R13620 gnd.n4543 gnd.n4542 0.155672
R13621 gnd.n4542 gnd.n4526 0.155672
R13622 gnd.n4535 gnd.n4526 0.155672
R13623 gnd.n4535 gnd.n4534 0.155672
R13624 gnd.n4518 gnd.n4490 0.155672
R13625 gnd.n4511 gnd.n4490 0.155672
R13626 gnd.n4511 gnd.n4510 0.155672
R13627 gnd.n4510 gnd.n4494 0.155672
R13628 gnd.n4503 gnd.n4494 0.155672
R13629 gnd.n4503 gnd.n4502 0.155672
R13630 gnd.n4486 gnd.n4458 0.155672
R13631 gnd.n4479 gnd.n4458 0.155672
R13632 gnd.n4479 gnd.n4478 0.155672
R13633 gnd.n4478 gnd.n4462 0.155672
R13634 gnd.n4471 gnd.n4462 0.155672
R13635 gnd.n4471 gnd.n4470 0.155672
R13636 gnd.n4454 gnd.n4426 0.155672
R13637 gnd.n4447 gnd.n4426 0.155672
R13638 gnd.n4447 gnd.n4446 0.155672
R13639 gnd.n4446 gnd.n4430 0.155672
R13640 gnd.n4439 gnd.n4430 0.155672
R13641 gnd.n4439 gnd.n4438 0.155672
R13642 gnd.n4423 gnd.n4395 0.155672
R13643 gnd.n4416 gnd.n4395 0.155672
R13644 gnd.n4416 gnd.n4415 0.155672
R13645 gnd.n4415 gnd.n4399 0.155672
R13646 gnd.n4408 gnd.n4399 0.155672
R13647 gnd.n4408 gnd.n4407 0.155672
R13648 gnd.n4770 gnd.n2017 0.152939
R13649 gnd.n4770 gnd.n4769 0.152939
R13650 gnd.n4769 gnd.n4768 0.152939
R13651 gnd.n4768 gnd.n2019 0.152939
R13652 gnd.n2020 gnd.n2019 0.152939
R13653 gnd.n2021 gnd.n2020 0.152939
R13654 gnd.n2022 gnd.n2021 0.152939
R13655 gnd.n2023 gnd.n2022 0.152939
R13656 gnd.n2024 gnd.n2023 0.152939
R13657 gnd.n2025 gnd.n2024 0.152939
R13658 gnd.n2026 gnd.n2025 0.152939
R13659 gnd.n2027 gnd.n2026 0.152939
R13660 gnd.n2028 gnd.n2027 0.152939
R13661 gnd.n2029 gnd.n2028 0.152939
R13662 gnd.n4740 gnd.n2029 0.152939
R13663 gnd.n4740 gnd.n4739 0.152939
R13664 gnd.n4012 gnd.n4011 0.152939
R13665 gnd.n4012 gnd.n3716 0.152939
R13666 gnd.n4040 gnd.n3716 0.152939
R13667 gnd.n4041 gnd.n4040 0.152939
R13668 gnd.n4042 gnd.n4041 0.152939
R13669 gnd.n4043 gnd.n4042 0.152939
R13670 gnd.n4043 gnd.n3688 0.152939
R13671 gnd.n4070 gnd.n3688 0.152939
R13672 gnd.n4071 gnd.n4070 0.152939
R13673 gnd.n4072 gnd.n4071 0.152939
R13674 gnd.n4072 gnd.n3666 0.152939
R13675 gnd.n4101 gnd.n3666 0.152939
R13676 gnd.n4102 gnd.n4101 0.152939
R13677 gnd.n4103 gnd.n4102 0.152939
R13678 gnd.n4104 gnd.n4103 0.152939
R13679 gnd.n4106 gnd.n4104 0.152939
R13680 gnd.n4106 gnd.n4105 0.152939
R13681 gnd.n4105 gnd.n3615 0.152939
R13682 gnd.n3616 gnd.n3615 0.152939
R13683 gnd.n3617 gnd.n3616 0.152939
R13684 gnd.n3636 gnd.n3617 0.152939
R13685 gnd.n3637 gnd.n3636 0.152939
R13686 gnd.n3637 gnd.n3519 0.152939
R13687 gnd.n4196 gnd.n3519 0.152939
R13688 gnd.n4197 gnd.n4196 0.152939
R13689 gnd.n4198 gnd.n4197 0.152939
R13690 gnd.n4199 gnd.n4198 0.152939
R13691 gnd.n4199 gnd.n3492 0.152939
R13692 gnd.n4236 gnd.n3492 0.152939
R13693 gnd.n4237 gnd.n4236 0.152939
R13694 gnd.n4238 gnd.n4237 0.152939
R13695 gnd.n4239 gnd.n4238 0.152939
R13696 gnd.n4239 gnd.n3465 0.152939
R13697 gnd.n4281 gnd.n3465 0.152939
R13698 gnd.n4282 gnd.n4281 0.152939
R13699 gnd.n4283 gnd.n4282 0.152939
R13700 gnd.n4284 gnd.n4283 0.152939
R13701 gnd.n4284 gnd.n3437 0.152939
R13702 gnd.n4321 gnd.n3437 0.152939
R13703 gnd.n4322 gnd.n4321 0.152939
R13704 gnd.n4323 gnd.n4322 0.152939
R13705 gnd.n4324 gnd.n4323 0.152939
R13706 gnd.n4324 gnd.n3410 0.152939
R13707 gnd.n4370 gnd.n3410 0.152939
R13708 gnd.n4371 gnd.n4370 0.152939
R13709 gnd.n4372 gnd.n4371 0.152939
R13710 gnd.n4373 gnd.n4372 0.152939
R13711 gnd.n4373 gnd.n3383 0.152939
R13712 gnd.n4664 gnd.n3383 0.152939
R13713 gnd.n4665 gnd.n4664 0.152939
R13714 gnd.n4666 gnd.n4665 0.152939
R13715 gnd.n4667 gnd.n4666 0.152939
R13716 gnd.n4668 gnd.n4667 0.152939
R13717 gnd.n4010 gnd.n3740 0.152939
R13718 gnd.n3761 gnd.n3740 0.152939
R13719 gnd.n3762 gnd.n3761 0.152939
R13720 gnd.n3768 gnd.n3762 0.152939
R13721 gnd.n3769 gnd.n3768 0.152939
R13722 gnd.n3770 gnd.n3769 0.152939
R13723 gnd.n3770 gnd.n3759 0.152939
R13724 gnd.n3778 gnd.n3759 0.152939
R13725 gnd.n3779 gnd.n3778 0.152939
R13726 gnd.n3780 gnd.n3779 0.152939
R13727 gnd.n3780 gnd.n3757 0.152939
R13728 gnd.n3788 gnd.n3757 0.152939
R13729 gnd.n3789 gnd.n3788 0.152939
R13730 gnd.n3790 gnd.n3789 0.152939
R13731 gnd.n3790 gnd.n3755 0.152939
R13732 gnd.n3798 gnd.n3755 0.152939
R13733 gnd.n4737 gnd.n2034 0.152939
R13734 gnd.n2036 gnd.n2034 0.152939
R13735 gnd.n2037 gnd.n2036 0.152939
R13736 gnd.n2038 gnd.n2037 0.152939
R13737 gnd.n2039 gnd.n2038 0.152939
R13738 gnd.n2040 gnd.n2039 0.152939
R13739 gnd.n2041 gnd.n2040 0.152939
R13740 gnd.n2042 gnd.n2041 0.152939
R13741 gnd.n2043 gnd.n2042 0.152939
R13742 gnd.n2044 gnd.n2043 0.152939
R13743 gnd.n2045 gnd.n2044 0.152939
R13744 gnd.n2046 gnd.n2045 0.152939
R13745 gnd.n2047 gnd.n2046 0.152939
R13746 gnd.n2048 gnd.n2047 0.152939
R13747 gnd.n2049 gnd.n2048 0.152939
R13748 gnd.n2050 gnd.n2049 0.152939
R13749 gnd.n2051 gnd.n2050 0.152939
R13750 gnd.n2052 gnd.n2051 0.152939
R13751 gnd.n2053 gnd.n2052 0.152939
R13752 gnd.n2054 gnd.n2053 0.152939
R13753 gnd.n2055 gnd.n2054 0.152939
R13754 gnd.n2056 gnd.n2055 0.152939
R13755 gnd.n2060 gnd.n2056 0.152939
R13756 gnd.n2061 gnd.n2060 0.152939
R13757 gnd.n2062 gnd.n2061 0.152939
R13758 gnd.n2063 gnd.n2062 0.152939
R13759 gnd.n4173 gnd.n4172 0.152939
R13760 gnd.n4174 gnd.n4173 0.152939
R13761 gnd.n4175 gnd.n4174 0.152939
R13762 gnd.n4176 gnd.n4175 0.152939
R13763 gnd.n4177 gnd.n4176 0.152939
R13764 gnd.n4178 gnd.n4177 0.152939
R13765 gnd.n4178 gnd.n3473 0.152939
R13766 gnd.n4257 gnd.n3473 0.152939
R13767 gnd.n4258 gnd.n4257 0.152939
R13768 gnd.n4259 gnd.n4258 0.152939
R13769 gnd.n4260 gnd.n4259 0.152939
R13770 gnd.n4261 gnd.n4260 0.152939
R13771 gnd.n4262 gnd.n4261 0.152939
R13772 gnd.n4263 gnd.n4262 0.152939
R13773 gnd.n4264 gnd.n4263 0.152939
R13774 gnd.n4265 gnd.n4264 0.152939
R13775 gnd.n4265 gnd.n3417 0.152939
R13776 gnd.n4342 gnd.n3417 0.152939
R13777 gnd.n4343 gnd.n4342 0.152939
R13778 gnd.n4344 gnd.n4343 0.152939
R13779 gnd.n4345 gnd.n4344 0.152939
R13780 gnd.n4346 gnd.n4345 0.152939
R13781 gnd.n4347 gnd.n4346 0.152939
R13782 gnd.n4348 gnd.n4347 0.152939
R13783 gnd.n4349 gnd.n4348 0.152939
R13784 gnd.n4350 gnd.n4349 0.152939
R13785 gnd.n4352 gnd.n4350 0.152939
R13786 gnd.n4352 gnd.n4351 0.152939
R13787 gnd.n3928 gnd.n3927 0.152939
R13788 gnd.n3928 gnd.n3818 0.152939
R13789 gnd.n3943 gnd.n3818 0.152939
R13790 gnd.n3944 gnd.n3943 0.152939
R13791 gnd.n3945 gnd.n3944 0.152939
R13792 gnd.n3945 gnd.n3806 0.152939
R13793 gnd.n3959 gnd.n3806 0.152939
R13794 gnd.n3960 gnd.n3959 0.152939
R13795 gnd.n3961 gnd.n3960 0.152939
R13796 gnd.n3962 gnd.n3961 0.152939
R13797 gnd.n3963 gnd.n3962 0.152939
R13798 gnd.n3964 gnd.n3963 0.152939
R13799 gnd.n3965 gnd.n3964 0.152939
R13800 gnd.n3966 gnd.n3965 0.152939
R13801 gnd.n3967 gnd.n3966 0.152939
R13802 gnd.n3968 gnd.n3967 0.152939
R13803 gnd.n3969 gnd.n3968 0.152939
R13804 gnd.n3970 gnd.n3969 0.152939
R13805 gnd.n3971 gnd.n3970 0.152939
R13806 gnd.n3972 gnd.n3971 0.152939
R13807 gnd.n3973 gnd.n3972 0.152939
R13808 gnd.n3973 gnd.n3672 0.152939
R13809 gnd.n4090 gnd.n3672 0.152939
R13810 gnd.n4091 gnd.n4090 0.152939
R13811 gnd.n4092 gnd.n4091 0.152939
R13812 gnd.n4093 gnd.n4092 0.152939
R13813 gnd.n4093 gnd.n3594 0.152939
R13814 gnd.n4170 gnd.n3594 0.152939
R13815 gnd.n3846 gnd.n3845 0.152939
R13816 gnd.n3847 gnd.n3846 0.152939
R13817 gnd.n3848 gnd.n3847 0.152939
R13818 gnd.n3849 gnd.n3848 0.152939
R13819 gnd.n3850 gnd.n3849 0.152939
R13820 gnd.n3851 gnd.n3850 0.152939
R13821 gnd.n3852 gnd.n3851 0.152939
R13822 gnd.n3853 gnd.n3852 0.152939
R13823 gnd.n3854 gnd.n3853 0.152939
R13824 gnd.n3855 gnd.n3854 0.152939
R13825 gnd.n3856 gnd.n3855 0.152939
R13826 gnd.n3857 gnd.n3856 0.152939
R13827 gnd.n3858 gnd.n3857 0.152939
R13828 gnd.n3859 gnd.n3858 0.152939
R13829 gnd.n3860 gnd.n3859 0.152939
R13830 gnd.n3861 gnd.n3860 0.152939
R13831 gnd.n3862 gnd.n3861 0.152939
R13832 gnd.n3863 gnd.n3862 0.152939
R13833 gnd.n3864 gnd.n3863 0.152939
R13834 gnd.n3865 gnd.n3864 0.152939
R13835 gnd.n3866 gnd.n3865 0.152939
R13836 gnd.n3867 gnd.n3866 0.152939
R13837 gnd.n3871 gnd.n3867 0.152939
R13838 gnd.n3872 gnd.n3871 0.152939
R13839 gnd.n3872 gnd.n3829 0.152939
R13840 gnd.n3926 gnd.n3829 0.152939
R13841 gnd.n3162 gnd.n3161 0.152939
R13842 gnd.n3161 gnd.n3160 0.152939
R13843 gnd.n3160 gnd.n2210 0.152939
R13844 gnd.n2215 gnd.n2210 0.152939
R13845 gnd.n2216 gnd.n2215 0.152939
R13846 gnd.n2217 gnd.n2216 0.152939
R13847 gnd.n2222 gnd.n2217 0.152939
R13848 gnd.n2223 gnd.n2222 0.152939
R13849 gnd.n2224 gnd.n2223 0.152939
R13850 gnd.n2225 gnd.n2224 0.152939
R13851 gnd.n2230 gnd.n2225 0.152939
R13852 gnd.n2231 gnd.n2230 0.152939
R13853 gnd.n2232 gnd.n2231 0.152939
R13854 gnd.n2233 gnd.n2232 0.152939
R13855 gnd.n2238 gnd.n2233 0.152939
R13856 gnd.n2239 gnd.n2238 0.152939
R13857 gnd.n2240 gnd.n2239 0.152939
R13858 gnd.n2241 gnd.n2240 0.152939
R13859 gnd.n2246 gnd.n2241 0.152939
R13860 gnd.n2247 gnd.n2246 0.152939
R13861 gnd.n2248 gnd.n2247 0.152939
R13862 gnd.n2249 gnd.n2248 0.152939
R13863 gnd.n2254 gnd.n2249 0.152939
R13864 gnd.n2255 gnd.n2254 0.152939
R13865 gnd.n2256 gnd.n2255 0.152939
R13866 gnd.n2257 gnd.n2256 0.152939
R13867 gnd.n2262 gnd.n2257 0.152939
R13868 gnd.n2263 gnd.n2262 0.152939
R13869 gnd.n2264 gnd.n2263 0.152939
R13870 gnd.n2265 gnd.n2264 0.152939
R13871 gnd.n2270 gnd.n2265 0.152939
R13872 gnd.n2271 gnd.n2270 0.152939
R13873 gnd.n2272 gnd.n2271 0.152939
R13874 gnd.n2273 gnd.n2272 0.152939
R13875 gnd.n2278 gnd.n2273 0.152939
R13876 gnd.n2279 gnd.n2278 0.152939
R13877 gnd.n2280 gnd.n2279 0.152939
R13878 gnd.n2281 gnd.n2280 0.152939
R13879 gnd.n2286 gnd.n2281 0.152939
R13880 gnd.n2287 gnd.n2286 0.152939
R13881 gnd.n2288 gnd.n2287 0.152939
R13882 gnd.n2289 gnd.n2288 0.152939
R13883 gnd.n2294 gnd.n2289 0.152939
R13884 gnd.n2295 gnd.n2294 0.152939
R13885 gnd.n2296 gnd.n2295 0.152939
R13886 gnd.n2297 gnd.n2296 0.152939
R13887 gnd.n2302 gnd.n2297 0.152939
R13888 gnd.n2303 gnd.n2302 0.152939
R13889 gnd.n2304 gnd.n2303 0.152939
R13890 gnd.n2305 gnd.n2304 0.152939
R13891 gnd.n2310 gnd.n2305 0.152939
R13892 gnd.n2311 gnd.n2310 0.152939
R13893 gnd.n2312 gnd.n2311 0.152939
R13894 gnd.n2313 gnd.n2312 0.152939
R13895 gnd.n2318 gnd.n2313 0.152939
R13896 gnd.n2319 gnd.n2318 0.152939
R13897 gnd.n2320 gnd.n2319 0.152939
R13898 gnd.n2321 gnd.n2320 0.152939
R13899 gnd.n2326 gnd.n2321 0.152939
R13900 gnd.n2327 gnd.n2326 0.152939
R13901 gnd.n2328 gnd.n2327 0.152939
R13902 gnd.n2329 gnd.n2328 0.152939
R13903 gnd.n2334 gnd.n2329 0.152939
R13904 gnd.n2335 gnd.n2334 0.152939
R13905 gnd.n2336 gnd.n2335 0.152939
R13906 gnd.n2337 gnd.n2336 0.152939
R13907 gnd.n2342 gnd.n2337 0.152939
R13908 gnd.n2343 gnd.n2342 0.152939
R13909 gnd.n2344 gnd.n2343 0.152939
R13910 gnd.n2345 gnd.n2344 0.152939
R13911 gnd.n2350 gnd.n2345 0.152939
R13912 gnd.n2351 gnd.n2350 0.152939
R13913 gnd.n2352 gnd.n2351 0.152939
R13914 gnd.n2353 gnd.n2352 0.152939
R13915 gnd.n2358 gnd.n2353 0.152939
R13916 gnd.n2359 gnd.n2358 0.152939
R13917 gnd.n2360 gnd.n2359 0.152939
R13918 gnd.n2361 gnd.n2360 0.152939
R13919 gnd.n2366 gnd.n2361 0.152939
R13920 gnd.n2367 gnd.n2366 0.152939
R13921 gnd.n2368 gnd.n2367 0.152939
R13922 gnd.n2369 gnd.n2368 0.152939
R13923 gnd.n2374 gnd.n2369 0.152939
R13924 gnd.n2375 gnd.n2374 0.152939
R13925 gnd.n2376 gnd.n2375 0.152939
R13926 gnd.n2377 gnd.n2376 0.152939
R13927 gnd.n2382 gnd.n2377 0.152939
R13928 gnd.n2383 gnd.n2382 0.152939
R13929 gnd.n2384 gnd.n2383 0.152939
R13930 gnd.n2385 gnd.n2384 0.152939
R13931 gnd.n2390 gnd.n2385 0.152939
R13932 gnd.n2391 gnd.n2390 0.152939
R13933 gnd.n2392 gnd.n2391 0.152939
R13934 gnd.n2393 gnd.n2392 0.152939
R13935 gnd.n2398 gnd.n2393 0.152939
R13936 gnd.n2399 gnd.n2398 0.152939
R13937 gnd.n2400 gnd.n2399 0.152939
R13938 gnd.n2401 gnd.n2400 0.152939
R13939 gnd.n2406 gnd.n2401 0.152939
R13940 gnd.n2407 gnd.n2406 0.152939
R13941 gnd.n2408 gnd.n2407 0.152939
R13942 gnd.n2409 gnd.n2408 0.152939
R13943 gnd.n2414 gnd.n2409 0.152939
R13944 gnd.n2415 gnd.n2414 0.152939
R13945 gnd.n2416 gnd.n2415 0.152939
R13946 gnd.n2417 gnd.n2416 0.152939
R13947 gnd.n2422 gnd.n2417 0.152939
R13948 gnd.n2423 gnd.n2422 0.152939
R13949 gnd.n2424 gnd.n2423 0.152939
R13950 gnd.n2425 gnd.n2424 0.152939
R13951 gnd.n2430 gnd.n2425 0.152939
R13952 gnd.n2431 gnd.n2430 0.152939
R13953 gnd.n2432 gnd.n2431 0.152939
R13954 gnd.n2433 gnd.n2432 0.152939
R13955 gnd.n2438 gnd.n2433 0.152939
R13956 gnd.n2439 gnd.n2438 0.152939
R13957 gnd.n2440 gnd.n2439 0.152939
R13958 gnd.n2441 gnd.n2440 0.152939
R13959 gnd.n2446 gnd.n2441 0.152939
R13960 gnd.n2447 gnd.n2446 0.152939
R13961 gnd.n2448 gnd.n2447 0.152939
R13962 gnd.n2449 gnd.n2448 0.152939
R13963 gnd.n2454 gnd.n2449 0.152939
R13964 gnd.n2455 gnd.n2454 0.152939
R13965 gnd.n2456 gnd.n2455 0.152939
R13966 gnd.n2457 gnd.n2456 0.152939
R13967 gnd.n2462 gnd.n2457 0.152939
R13968 gnd.n2463 gnd.n2462 0.152939
R13969 gnd.n2464 gnd.n2463 0.152939
R13970 gnd.n2465 gnd.n2464 0.152939
R13971 gnd.n2470 gnd.n2465 0.152939
R13972 gnd.n2471 gnd.n2470 0.152939
R13973 gnd.n2472 gnd.n2471 0.152939
R13974 gnd.n2473 gnd.n2472 0.152939
R13975 gnd.n2478 gnd.n2473 0.152939
R13976 gnd.n2479 gnd.n2478 0.152939
R13977 gnd.n2480 gnd.n2479 0.152939
R13978 gnd.n2481 gnd.n2480 0.152939
R13979 gnd.n2486 gnd.n2481 0.152939
R13980 gnd.n2487 gnd.n2486 0.152939
R13981 gnd.n2488 gnd.n2487 0.152939
R13982 gnd.n2489 gnd.n2488 0.152939
R13983 gnd.n2494 gnd.n2489 0.152939
R13984 gnd.n2495 gnd.n2494 0.152939
R13985 gnd.n2496 gnd.n2495 0.152939
R13986 gnd.n2497 gnd.n2496 0.152939
R13987 gnd.n2502 gnd.n2497 0.152939
R13988 gnd.n2503 gnd.n2502 0.152939
R13989 gnd.n2504 gnd.n2503 0.152939
R13990 gnd.n2505 gnd.n2504 0.152939
R13991 gnd.n2510 gnd.n2505 0.152939
R13992 gnd.n2511 gnd.n2510 0.152939
R13993 gnd.n2512 gnd.n2511 0.152939
R13994 gnd.n2513 gnd.n2512 0.152939
R13995 gnd.n2848 gnd.n2519 0.152939
R13996 gnd.n2848 gnd.n2847 0.152939
R13997 gnd.n2847 gnd.n2846 0.152939
R13998 gnd.n2846 gnd.n2520 0.152939
R13999 gnd.n2525 gnd.n2520 0.152939
R14000 gnd.n2526 gnd.n2525 0.152939
R14001 gnd.n2527 gnd.n2526 0.152939
R14002 gnd.n2532 gnd.n2527 0.152939
R14003 gnd.n2533 gnd.n2532 0.152939
R14004 gnd.n2534 gnd.n2533 0.152939
R14005 gnd.n2535 gnd.n2534 0.152939
R14006 gnd.n2540 gnd.n2535 0.152939
R14007 gnd.n2541 gnd.n2540 0.152939
R14008 gnd.n2542 gnd.n2541 0.152939
R14009 gnd.n2543 gnd.n2542 0.152939
R14010 gnd.n2548 gnd.n2543 0.152939
R14011 gnd.n2549 gnd.n2548 0.152939
R14012 gnd.n2550 gnd.n2549 0.152939
R14013 gnd.n2551 gnd.n2550 0.152939
R14014 gnd.n2556 gnd.n2551 0.152939
R14015 gnd.n2557 gnd.n2556 0.152939
R14016 gnd.n2558 gnd.n2557 0.152939
R14017 gnd.n2559 gnd.n2558 0.152939
R14018 gnd.n2564 gnd.n2559 0.152939
R14019 gnd.n2565 gnd.n2564 0.152939
R14020 gnd.n2566 gnd.n2565 0.152939
R14021 gnd.n2567 gnd.n2566 0.152939
R14022 gnd.n2572 gnd.n2567 0.152939
R14023 gnd.n2573 gnd.n2572 0.152939
R14024 gnd.n2574 gnd.n2573 0.152939
R14025 gnd.n2575 gnd.n2574 0.152939
R14026 gnd.n2580 gnd.n2575 0.152939
R14027 gnd.n2581 gnd.n2580 0.152939
R14028 gnd.n2582 gnd.n2581 0.152939
R14029 gnd.n2583 gnd.n2582 0.152939
R14030 gnd.n2588 gnd.n2583 0.152939
R14031 gnd.n2589 gnd.n2588 0.152939
R14032 gnd.n2590 gnd.n2589 0.152939
R14033 gnd.n2591 gnd.n2590 0.152939
R14034 gnd.n2596 gnd.n2591 0.152939
R14035 gnd.n2597 gnd.n2596 0.152939
R14036 gnd.n2598 gnd.n2597 0.152939
R14037 gnd.n2599 gnd.n2598 0.152939
R14038 gnd.n2604 gnd.n2599 0.152939
R14039 gnd.n2605 gnd.n2604 0.152939
R14040 gnd.n2606 gnd.n2605 0.152939
R14041 gnd.n2607 gnd.n2606 0.152939
R14042 gnd.n2612 gnd.n2607 0.152939
R14043 gnd.n2613 gnd.n2612 0.152939
R14044 gnd.n2614 gnd.n2613 0.152939
R14045 gnd.n2615 gnd.n2614 0.152939
R14046 gnd.n2620 gnd.n2615 0.152939
R14047 gnd.n2621 gnd.n2620 0.152939
R14048 gnd.n2622 gnd.n2621 0.152939
R14049 gnd.n2623 gnd.n2622 0.152939
R14050 gnd.n2628 gnd.n2623 0.152939
R14051 gnd.n2629 gnd.n2628 0.152939
R14052 gnd.n2630 gnd.n2629 0.152939
R14053 gnd.n2631 gnd.n2630 0.152939
R14054 gnd.n2636 gnd.n2631 0.152939
R14055 gnd.n2637 gnd.n2636 0.152939
R14056 gnd.n2638 gnd.n2637 0.152939
R14057 gnd.n2639 gnd.n2638 0.152939
R14058 gnd.n2644 gnd.n2639 0.152939
R14059 gnd.n2645 gnd.n2644 0.152939
R14060 gnd.n2646 gnd.n2645 0.152939
R14061 gnd.n2647 gnd.n2646 0.152939
R14062 gnd.n2652 gnd.n2647 0.152939
R14063 gnd.n2653 gnd.n2652 0.152939
R14064 gnd.n2654 gnd.n2653 0.152939
R14065 gnd.n2655 gnd.n2654 0.152939
R14066 gnd.n2660 gnd.n2655 0.152939
R14067 gnd.n2661 gnd.n2660 0.152939
R14068 gnd.n2662 gnd.n2661 0.152939
R14069 gnd.n2663 gnd.n2662 0.152939
R14070 gnd.n2668 gnd.n2663 0.152939
R14071 gnd.n2669 gnd.n2668 0.152939
R14072 gnd.n2670 gnd.n2669 0.152939
R14073 gnd.n2671 gnd.n2670 0.152939
R14074 gnd.n2676 gnd.n2671 0.152939
R14075 gnd.n2677 gnd.n2676 0.152939
R14076 gnd.n2678 gnd.n2677 0.152939
R14077 gnd.n2679 gnd.n2678 0.152939
R14078 gnd.n2680 gnd.n2679 0.152939
R14079 gnd.n119 gnd.n96 0.152939
R14080 gnd.n120 gnd.n119 0.152939
R14081 gnd.n121 gnd.n120 0.152939
R14082 gnd.n138 gnd.n121 0.152939
R14083 gnd.n139 gnd.n138 0.152939
R14084 gnd.n140 gnd.n139 0.152939
R14085 gnd.n141 gnd.n140 0.152939
R14086 gnd.n156 gnd.n141 0.152939
R14087 gnd.n157 gnd.n156 0.152939
R14088 gnd.n158 gnd.n157 0.152939
R14089 gnd.n159 gnd.n158 0.152939
R14090 gnd.n176 gnd.n159 0.152939
R14091 gnd.n177 gnd.n176 0.152939
R14092 gnd.n178 gnd.n177 0.152939
R14093 gnd.n179 gnd.n178 0.152939
R14094 gnd.n195 gnd.n179 0.152939
R14095 gnd.n196 gnd.n195 0.152939
R14096 gnd.n197 gnd.n196 0.152939
R14097 gnd.n198 gnd.n197 0.152939
R14098 gnd.n213 gnd.n198 0.152939
R14099 gnd.n7676 gnd.n213 0.152939
R14100 gnd.n7757 gnd.n84 0.152939
R14101 gnd.n7437 gnd.n84 0.152939
R14102 gnd.n7438 gnd.n7437 0.152939
R14103 gnd.n7439 gnd.n7438 0.152939
R14104 gnd.n7440 gnd.n7439 0.152939
R14105 gnd.n7441 gnd.n7440 0.152939
R14106 gnd.n7442 gnd.n7441 0.152939
R14107 gnd.n7443 gnd.n7442 0.152939
R14108 gnd.n7444 gnd.n7443 0.152939
R14109 gnd.n7445 gnd.n7444 0.152939
R14110 gnd.n7446 gnd.n7445 0.152939
R14111 gnd.n7447 gnd.n7446 0.152939
R14112 gnd.n7448 gnd.n7447 0.152939
R14113 gnd.n7449 gnd.n7448 0.152939
R14114 gnd.n7451 gnd.n7449 0.152939
R14115 gnd.n7451 gnd.n7450 0.152939
R14116 gnd.n7450 gnd.n357 0.152939
R14117 gnd.n7518 gnd.n357 0.152939
R14118 gnd.n7519 gnd.n7518 0.152939
R14119 gnd.n7520 gnd.n7519 0.152939
R14120 gnd.n7520 gnd.n354 0.152939
R14121 gnd.n7525 gnd.n354 0.152939
R14122 gnd.n7526 gnd.n7525 0.152939
R14123 gnd.n7527 gnd.n7526 0.152939
R14124 gnd.n7527 gnd.n351 0.152939
R14125 gnd.n7532 gnd.n351 0.152939
R14126 gnd.n7565 gnd.n317 0.152939
R14127 gnd.n319 gnd.n317 0.152939
R14128 gnd.n323 gnd.n319 0.152939
R14129 gnd.n324 gnd.n323 0.152939
R14130 gnd.n325 gnd.n324 0.152939
R14131 gnd.n326 gnd.n325 0.152939
R14132 gnd.n330 gnd.n326 0.152939
R14133 gnd.n331 gnd.n330 0.152939
R14134 gnd.n332 gnd.n331 0.152939
R14135 gnd.n333 gnd.n332 0.152939
R14136 gnd.n337 gnd.n333 0.152939
R14137 gnd.n338 gnd.n337 0.152939
R14138 gnd.n339 gnd.n338 0.152939
R14139 gnd.n340 gnd.n339 0.152939
R14140 gnd.n344 gnd.n340 0.152939
R14141 gnd.n345 gnd.n344 0.152939
R14142 gnd.n7534 gnd.n345 0.152939
R14143 gnd.n7534 gnd.n7533 0.152939
R14144 gnd.n7675 gnd.n214 0.152939
R14145 gnd.n216 gnd.n214 0.152939
R14146 gnd.n220 gnd.n216 0.152939
R14147 gnd.n221 gnd.n220 0.152939
R14148 gnd.n222 gnd.n221 0.152939
R14149 gnd.n223 gnd.n222 0.152939
R14150 gnd.n227 gnd.n223 0.152939
R14151 gnd.n228 gnd.n227 0.152939
R14152 gnd.n229 gnd.n228 0.152939
R14153 gnd.n230 gnd.n229 0.152939
R14154 gnd.n234 gnd.n230 0.152939
R14155 gnd.n235 gnd.n234 0.152939
R14156 gnd.n236 gnd.n235 0.152939
R14157 gnd.n237 gnd.n236 0.152939
R14158 gnd.n241 gnd.n237 0.152939
R14159 gnd.n242 gnd.n241 0.152939
R14160 gnd.n243 gnd.n242 0.152939
R14161 gnd.n244 gnd.n243 0.152939
R14162 gnd.n248 gnd.n244 0.152939
R14163 gnd.n249 gnd.n248 0.152939
R14164 gnd.n250 gnd.n249 0.152939
R14165 gnd.n251 gnd.n250 0.152939
R14166 gnd.n255 gnd.n251 0.152939
R14167 gnd.n256 gnd.n255 0.152939
R14168 gnd.n257 gnd.n256 0.152939
R14169 gnd.n258 gnd.n257 0.152939
R14170 gnd.n262 gnd.n258 0.152939
R14171 gnd.n263 gnd.n262 0.152939
R14172 gnd.n264 gnd.n263 0.152939
R14173 gnd.n265 gnd.n264 0.152939
R14174 gnd.n269 gnd.n265 0.152939
R14175 gnd.n270 gnd.n269 0.152939
R14176 gnd.n271 gnd.n270 0.152939
R14177 gnd.n272 gnd.n271 0.152939
R14178 gnd.n276 gnd.n272 0.152939
R14179 gnd.n277 gnd.n276 0.152939
R14180 gnd.n7606 gnd.n277 0.152939
R14181 gnd.n7606 gnd.n7605 0.152939
R14182 gnd.n7605 gnd.n7604 0.152939
R14183 gnd.n7604 gnd.n281 0.152939
R14184 gnd.n287 gnd.n281 0.152939
R14185 gnd.n288 gnd.n287 0.152939
R14186 gnd.n289 gnd.n288 0.152939
R14187 gnd.n290 gnd.n289 0.152939
R14188 gnd.n294 gnd.n290 0.152939
R14189 gnd.n295 gnd.n294 0.152939
R14190 gnd.n296 gnd.n295 0.152939
R14191 gnd.n297 gnd.n296 0.152939
R14192 gnd.n301 gnd.n297 0.152939
R14193 gnd.n302 gnd.n301 0.152939
R14194 gnd.n303 gnd.n302 0.152939
R14195 gnd.n304 gnd.n303 0.152939
R14196 gnd.n308 gnd.n304 0.152939
R14197 gnd.n309 gnd.n308 0.152939
R14198 gnd.n310 gnd.n309 0.152939
R14199 gnd.n311 gnd.n310 0.152939
R14200 gnd.n316 gnd.n311 0.152939
R14201 gnd.n7567 gnd.n316 0.152939
R14202 gnd.n7208 gnd.n526 0.152939
R14203 gnd.n802 gnd.n526 0.152939
R14204 gnd.n803 gnd.n802 0.152939
R14205 gnd.n803 gnd.n801 0.152939
R14206 gnd.n810 gnd.n801 0.152939
R14207 gnd.n811 gnd.n810 0.152939
R14208 gnd.n812 gnd.n811 0.152939
R14209 gnd.n812 gnd.n799 0.152939
R14210 gnd.n820 gnd.n799 0.152939
R14211 gnd.n821 gnd.n820 0.152939
R14212 gnd.n822 gnd.n821 0.152939
R14213 gnd.n822 gnd.n797 0.152939
R14214 gnd.n830 gnd.n797 0.152939
R14215 gnd.n831 gnd.n830 0.152939
R14216 gnd.n832 gnd.n831 0.152939
R14217 gnd.n832 gnd.n795 0.152939
R14218 gnd.n840 gnd.n795 0.152939
R14219 gnd.n841 gnd.n840 0.152939
R14220 gnd.n841 gnd.n791 0.152939
R14221 gnd.n849 gnd.n791 0.152939
R14222 gnd.n850 gnd.n849 0.152939
R14223 gnd.n851 gnd.n850 0.152939
R14224 gnd.n851 gnd.n789 0.152939
R14225 gnd.n859 gnd.n789 0.152939
R14226 gnd.n860 gnd.n859 0.152939
R14227 gnd.n863 gnd.n862 0.152939
R14228 gnd.n864 gnd.n863 0.152939
R14229 gnd.n865 gnd.n864 0.152939
R14230 gnd.n866 gnd.n865 0.152939
R14231 gnd.n867 gnd.n866 0.152939
R14232 gnd.n868 gnd.n867 0.152939
R14233 gnd.n869 gnd.n868 0.152939
R14234 gnd.n870 gnd.n869 0.152939
R14235 gnd.n871 gnd.n870 0.152939
R14236 gnd.n874 gnd.n871 0.152939
R14237 gnd.n875 gnd.n874 0.152939
R14238 gnd.n876 gnd.n875 0.152939
R14239 gnd.n877 gnd.n876 0.152939
R14240 gnd.n878 gnd.n877 0.152939
R14241 gnd.n879 gnd.n878 0.152939
R14242 gnd.n880 gnd.n879 0.152939
R14243 gnd.n881 gnd.n880 0.152939
R14244 gnd.n882 gnd.n881 0.152939
R14245 gnd.n883 gnd.n882 0.152939
R14246 gnd.n884 gnd.n883 0.152939
R14247 gnd.n885 gnd.n884 0.152939
R14248 gnd.n886 gnd.n885 0.152939
R14249 gnd.n887 gnd.n886 0.152939
R14250 gnd.n888 gnd.n887 0.152939
R14251 gnd.n889 gnd.n888 0.152939
R14252 gnd.n890 gnd.n889 0.152939
R14253 gnd.n891 gnd.n890 0.152939
R14254 gnd.n892 gnd.n891 0.152939
R14255 gnd.n898 gnd.n892 0.152939
R14256 gnd.n898 gnd.n897 0.152939
R14257 gnd.n7210 gnd.n7209 0.152939
R14258 gnd.n7210 gnd.n498 0.152939
R14259 gnd.n7244 gnd.n498 0.152939
R14260 gnd.n7245 gnd.n7244 0.152939
R14261 gnd.n7246 gnd.n7245 0.152939
R14262 gnd.n7247 gnd.n7246 0.152939
R14263 gnd.n7247 gnd.n463 0.152939
R14264 gnd.n7290 gnd.n463 0.152939
R14265 gnd.n7291 gnd.n7290 0.152939
R14266 gnd.n7292 gnd.n7291 0.152939
R14267 gnd.n7293 gnd.n7292 0.152939
R14268 gnd.n7293 gnd.n428 0.152939
R14269 gnd.n7337 gnd.n428 0.152939
R14270 gnd.n7338 gnd.n7337 0.152939
R14271 gnd.n7339 gnd.n7338 0.152939
R14272 gnd.n7340 gnd.n7339 0.152939
R14273 gnd.n7340 gnd.n396 0.152939
R14274 gnd.n7381 gnd.n396 0.152939
R14275 gnd.n7382 gnd.n7381 0.152939
R14276 gnd.n7383 gnd.n7382 0.152939
R14277 gnd.n7383 gnd.n97 0.152939
R14278 gnd.n4930 gnd.n4896 0.152939
R14279 gnd.n4897 gnd.n4896 0.152939
R14280 gnd.n4898 gnd.n4897 0.152939
R14281 gnd.n4899 gnd.n4898 0.152939
R14282 gnd.n4900 gnd.n4899 0.152939
R14283 gnd.n4901 gnd.n4900 0.152939
R14284 gnd.n4902 gnd.n4901 0.152939
R14285 gnd.n4903 gnd.n4902 0.152939
R14286 gnd.n4904 gnd.n4903 0.152939
R14287 gnd.n4905 gnd.n4904 0.152939
R14288 gnd.n4906 gnd.n4905 0.152939
R14289 gnd.n4907 gnd.n4906 0.152939
R14290 gnd.n4908 gnd.n4907 0.152939
R14291 gnd.n4908 gnd.n1912 0.152939
R14292 gnd.n5175 gnd.n1912 0.152939
R14293 gnd.n5176 gnd.n5175 0.152939
R14294 gnd.n5177 gnd.n5176 0.152939
R14295 gnd.n5178 gnd.n5177 0.152939
R14296 gnd.n5178 gnd.n1887 0.152939
R14297 gnd.n5210 gnd.n1887 0.152939
R14298 gnd.n5211 gnd.n5210 0.152939
R14299 gnd.n5212 gnd.n5211 0.152939
R14300 gnd.n5213 gnd.n5212 0.152939
R14301 gnd.n5214 gnd.n5213 0.152939
R14302 gnd.n5215 gnd.n5214 0.152939
R14303 gnd.n5217 gnd.n5215 0.152939
R14304 gnd.n4969 gnd.n4877 0.152939
R14305 gnd.n4878 gnd.n4877 0.152939
R14306 gnd.n4879 gnd.n4878 0.152939
R14307 gnd.n4880 gnd.n4879 0.152939
R14308 gnd.n4881 gnd.n4880 0.152939
R14309 gnd.n4882 gnd.n4881 0.152939
R14310 gnd.n4883 gnd.n4882 0.152939
R14311 gnd.n4884 gnd.n4883 0.152939
R14312 gnd.n4885 gnd.n4884 0.152939
R14313 gnd.n4886 gnd.n4885 0.152939
R14314 gnd.n4887 gnd.n4886 0.152939
R14315 gnd.n4888 gnd.n4887 0.152939
R14316 gnd.n4889 gnd.n4888 0.152939
R14317 gnd.n4890 gnd.n4889 0.152939
R14318 gnd.n4891 gnd.n4890 0.152939
R14319 gnd.n4934 gnd.n4891 0.152939
R14320 gnd.n4934 gnd.n4933 0.152939
R14321 gnd.n4933 gnd.n4932 0.152939
R14322 gnd.n5298 gnd.n5297 0.152939
R14323 gnd.n5299 gnd.n5298 0.152939
R14324 gnd.n5299 gnd.n1792 0.152939
R14325 gnd.n5336 gnd.n1792 0.152939
R14326 gnd.n5337 gnd.n5336 0.152939
R14327 gnd.n5338 gnd.n5337 0.152939
R14328 gnd.n5339 gnd.n5338 0.152939
R14329 gnd.n5339 gnd.n1757 0.152939
R14330 gnd.n5384 gnd.n1757 0.152939
R14331 gnd.n5385 gnd.n5384 0.152939
R14332 gnd.n5386 gnd.n5385 0.152939
R14333 gnd.n5387 gnd.n5386 0.152939
R14334 gnd.n5387 gnd.n1730 0.152939
R14335 gnd.n5418 gnd.n1730 0.152939
R14336 gnd.n5419 gnd.n5418 0.152939
R14337 gnd.n5420 gnd.n5419 0.152939
R14338 gnd.n5420 gnd.n1661 0.152939
R14339 gnd.n5765 gnd.n1661 0.152939
R14340 gnd.n5766 gnd.n5765 0.152939
R14341 gnd.n5767 gnd.n5766 0.152939
R14342 gnd.n5860 gnd.n5767 0.152939
R14343 gnd.n5859 gnd.n5768 0.152939
R14344 gnd.n5771 gnd.n5768 0.152939
R14345 gnd.n5772 gnd.n5771 0.152939
R14346 gnd.n5773 gnd.n5772 0.152939
R14347 gnd.n5777 gnd.n5773 0.152939
R14348 gnd.n5778 gnd.n5777 0.152939
R14349 gnd.n5779 gnd.n5778 0.152939
R14350 gnd.n5780 gnd.n5779 0.152939
R14351 gnd.n5784 gnd.n5780 0.152939
R14352 gnd.n5785 gnd.n5784 0.152939
R14353 gnd.n5786 gnd.n5785 0.152939
R14354 gnd.n5787 gnd.n5786 0.152939
R14355 gnd.n5791 gnd.n5787 0.152939
R14356 gnd.n5792 gnd.n5791 0.152939
R14357 gnd.n5793 gnd.n5792 0.152939
R14358 gnd.n5794 gnd.n5793 0.152939
R14359 gnd.n5801 gnd.n5794 0.152939
R14360 gnd.n5802 gnd.n5801 0.152939
R14361 gnd.n5803 gnd.n5802 0.152939
R14362 gnd.n5804 gnd.n5803 0.152939
R14363 gnd.n5808 gnd.n5804 0.152939
R14364 gnd.n5809 gnd.n5808 0.152939
R14365 gnd.n5810 gnd.n5809 0.152939
R14366 gnd.n5811 gnd.n5810 0.152939
R14367 gnd.n5811 gnd.n1592 0.152939
R14368 gnd.n5927 gnd.n5926 0.152939
R14369 gnd.n5926 gnd.n1593 0.152939
R14370 gnd.n1600 gnd.n1593 0.152939
R14371 gnd.n1601 gnd.n1600 0.152939
R14372 gnd.n1602 gnd.n1601 0.152939
R14373 gnd.n1603 gnd.n1602 0.152939
R14374 gnd.n1607 gnd.n1603 0.152939
R14375 gnd.n1608 gnd.n1607 0.152939
R14376 gnd.n5909 gnd.n1608 0.152939
R14377 gnd.n5909 gnd.n5908 0.152939
R14378 gnd.n5908 gnd.n5907 0.152939
R14379 gnd.n5907 gnd.n1612 0.152939
R14380 gnd.n1618 gnd.n1612 0.152939
R14381 gnd.n1619 gnd.n1618 0.152939
R14382 gnd.n1620 gnd.n1619 0.152939
R14383 gnd.n1621 gnd.n1620 0.152939
R14384 gnd.n1625 gnd.n1621 0.152939
R14385 gnd.n1626 gnd.n1625 0.152939
R14386 gnd.n1627 gnd.n1626 0.152939
R14387 gnd.n1628 gnd.n1627 0.152939
R14388 gnd.n1632 gnd.n1628 0.152939
R14389 gnd.n1633 gnd.n1632 0.152939
R14390 gnd.n1634 gnd.n1633 0.152939
R14391 gnd.n1635 gnd.n1634 0.152939
R14392 gnd.n1639 gnd.n1635 0.152939
R14393 gnd.n1640 gnd.n1639 0.152939
R14394 gnd.n1641 gnd.n1640 0.152939
R14395 gnd.n1642 gnd.n1641 0.152939
R14396 gnd.n1648 gnd.n1642 0.152939
R14397 gnd.n5870 gnd.n1648 0.152939
R14398 gnd.n4815 gnd.n4814 0.152939
R14399 gnd.n4816 gnd.n4815 0.152939
R14400 gnd.n4817 gnd.n4816 0.152939
R14401 gnd.n4818 gnd.n4817 0.152939
R14402 gnd.n4819 gnd.n4818 0.152939
R14403 gnd.n4820 gnd.n4819 0.152939
R14404 gnd.n4821 gnd.n4820 0.152939
R14405 gnd.n4822 gnd.n4821 0.152939
R14406 gnd.n4823 gnd.n4822 0.152939
R14407 gnd.n4824 gnd.n4823 0.152939
R14408 gnd.n4825 gnd.n4824 0.152939
R14409 gnd.n4826 gnd.n4825 0.152939
R14410 gnd.n4827 gnd.n4826 0.152939
R14411 gnd.n4828 gnd.n4827 0.152939
R14412 gnd.n4829 gnd.n4828 0.152939
R14413 gnd.n4830 gnd.n4829 0.152939
R14414 gnd.n4831 gnd.n4830 0.152939
R14415 gnd.n4834 gnd.n4831 0.152939
R14416 gnd.n4835 gnd.n4834 0.152939
R14417 gnd.n4836 gnd.n4835 0.152939
R14418 gnd.n4837 gnd.n4836 0.152939
R14419 gnd.n4838 gnd.n4837 0.152939
R14420 gnd.n4839 gnd.n4838 0.152939
R14421 gnd.n4840 gnd.n4839 0.152939
R14422 gnd.n4841 gnd.n4840 0.152939
R14423 gnd.n4842 gnd.n4841 0.152939
R14424 gnd.n4843 gnd.n4842 0.152939
R14425 gnd.n4844 gnd.n4843 0.152939
R14426 gnd.n4845 gnd.n4844 0.152939
R14427 gnd.n4846 gnd.n4845 0.152939
R14428 gnd.n4847 gnd.n4846 0.152939
R14429 gnd.n4848 gnd.n4847 0.152939
R14430 gnd.n4849 gnd.n4848 0.152939
R14431 gnd.n4850 gnd.n4849 0.152939
R14432 gnd.n4851 gnd.n4850 0.152939
R14433 gnd.n4852 gnd.n4851 0.152939
R14434 gnd.n4853 gnd.n4852 0.152939
R14435 gnd.n4856 gnd.n4853 0.152939
R14436 gnd.n4857 gnd.n4856 0.152939
R14437 gnd.n4858 gnd.n4857 0.152939
R14438 gnd.n4859 gnd.n4858 0.152939
R14439 gnd.n4860 gnd.n4859 0.152939
R14440 gnd.n4861 gnd.n4860 0.152939
R14441 gnd.n4862 gnd.n4861 0.152939
R14442 gnd.n4863 gnd.n4862 0.152939
R14443 gnd.n4864 gnd.n4863 0.152939
R14444 gnd.n4865 gnd.n4864 0.152939
R14445 gnd.n4866 gnd.n4865 0.152939
R14446 gnd.n4867 gnd.n4866 0.152939
R14447 gnd.n4868 gnd.n4867 0.152939
R14448 gnd.n4869 gnd.n4868 0.152939
R14449 gnd.n4870 gnd.n4869 0.152939
R14450 gnd.n4871 gnd.n4870 0.152939
R14451 gnd.n4872 gnd.n4871 0.152939
R14452 gnd.n4873 gnd.n4872 0.152939
R14453 gnd.n4874 gnd.n4873 0.152939
R14454 gnd.n4972 gnd.n4874 0.152939
R14455 gnd.n4972 gnd.n4971 0.152939
R14456 gnd.n5101 gnd.n1976 0.152939
R14457 gnd.n5102 gnd.n5101 0.152939
R14458 gnd.n5103 gnd.n5102 0.152939
R14459 gnd.n5103 gnd.n1957 0.152939
R14460 gnd.n5121 gnd.n1957 0.152939
R14461 gnd.n5122 gnd.n5121 0.152939
R14462 gnd.n5123 gnd.n5122 0.152939
R14463 gnd.n5123 gnd.n1940 0.152939
R14464 gnd.n5141 gnd.n1940 0.152939
R14465 gnd.n5142 gnd.n5141 0.152939
R14466 gnd.n5143 gnd.n5142 0.152939
R14467 gnd.n5143 gnd.n1920 0.152939
R14468 gnd.n5165 gnd.n1920 0.152939
R14469 gnd.n5166 gnd.n5165 0.152939
R14470 gnd.n5167 gnd.n5166 0.152939
R14471 gnd.n5168 gnd.n5167 0.152939
R14472 gnd.n5168 gnd.n1895 0.152939
R14473 gnd.n5200 gnd.n1895 0.152939
R14474 gnd.n5201 gnd.n5200 0.152939
R14475 gnd.n5202 gnd.n5201 0.152939
R14476 gnd.n5202 gnd.n1828 0.152939
R14477 gnd.n2078 gnd.n2076 0.152939
R14478 gnd.n2078 gnd.n2077 0.152939
R14479 gnd.n2077 gnd.n1809 0.152939
R14480 gnd.n5318 gnd.n1809 0.152939
R14481 gnd.n5319 gnd.n5318 0.152939
R14482 gnd.n5320 gnd.n5319 0.152939
R14483 gnd.n5321 gnd.n5320 0.152939
R14484 gnd.n5321 gnd.n1773 0.152939
R14485 gnd.n5363 gnd.n1773 0.152939
R14486 gnd.n5364 gnd.n5363 0.152939
R14487 gnd.n5365 gnd.n5364 0.152939
R14488 gnd.n5366 gnd.n5365 0.152939
R14489 gnd.n5367 gnd.n5366 0.152939
R14490 gnd.n5367 gnd.n1723 0.152939
R14491 gnd.n5427 gnd.n1723 0.152939
R14492 gnd.n5428 gnd.n5427 0.152939
R14493 gnd.n5429 gnd.n5428 0.152939
R14494 gnd.n5429 gnd.n1719 0.152939
R14495 gnd.n5435 gnd.n1719 0.152939
R14496 gnd.n5436 gnd.n5435 0.152939
R14497 gnd.n5437 gnd.n5436 0.152939
R14498 gnd.n5438 gnd.n5437 0.152939
R14499 gnd.n5439 gnd.n5438 0.152939
R14500 gnd.n5442 gnd.n5439 0.152939
R14501 gnd.n5443 gnd.n5442 0.152939
R14502 gnd.n5444 gnd.n5443 0.152939
R14503 gnd.n5445 gnd.n5444 0.152939
R14504 gnd.n5495 gnd.n5445 0.152939
R14505 gnd.n5496 gnd.n5495 0.152939
R14506 gnd.n5516 gnd.n5496 0.152939
R14507 gnd.n5517 gnd.n5516 0.152939
R14508 gnd.n5518 gnd.n5517 0.152939
R14509 gnd.n5518 gnd.n5481 0.152939
R14510 gnd.n5535 gnd.n5481 0.152939
R14511 gnd.n5536 gnd.n5535 0.152939
R14512 gnd.n5537 gnd.n5536 0.152939
R14513 gnd.n5538 gnd.n5537 0.152939
R14514 gnd.n5538 gnd.n1462 0.152939
R14515 gnd.n6015 gnd.n1462 0.152939
R14516 gnd.n6016 gnd.n6015 0.152939
R14517 gnd.n6017 gnd.n6016 0.152939
R14518 gnd.n6017 gnd.n1432 0.152939
R14519 gnd.n6075 gnd.n1432 0.152939
R14520 gnd.n6076 gnd.n6075 0.152939
R14521 gnd.n6077 gnd.n6076 0.152939
R14522 gnd.n6077 gnd.n1405 0.152939
R14523 gnd.n6117 gnd.n1405 0.152939
R14524 gnd.n6118 gnd.n6117 0.152939
R14525 gnd.n6119 gnd.n6118 0.152939
R14526 gnd.n6120 gnd.n6119 0.152939
R14527 gnd.n6121 gnd.n6120 0.152939
R14528 gnd.n6122 gnd.n6121 0.152939
R14529 gnd.n6122 gnd.n1361 0.152939
R14530 gnd.n6188 gnd.n1361 0.152939
R14531 gnd.n6189 gnd.n6188 0.152939
R14532 gnd.n6190 gnd.n6189 0.152939
R14533 gnd.n6190 gnd.n1330 0.152939
R14534 gnd.n6239 gnd.n1330 0.152939
R14535 gnd.n6240 gnd.n6239 0.152939
R14536 gnd.n6241 gnd.n6240 0.152939
R14537 gnd.n6241 gnd.n1326 0.152939
R14538 gnd.n6250 gnd.n1326 0.152939
R14539 gnd.n6251 gnd.n6250 0.152939
R14540 gnd.n6252 gnd.n6251 0.152939
R14541 gnd.n6252 gnd.n1267 0.152939
R14542 gnd.n6385 gnd.n1267 0.152939
R14543 gnd.n6386 gnd.n6385 0.152939
R14544 gnd.n6387 gnd.n6386 0.152939
R14545 gnd.n6387 gnd.n1243 0.152939
R14546 gnd.n6412 gnd.n1243 0.152939
R14547 gnd.n6413 gnd.n6412 0.152939
R14548 gnd.n6414 gnd.n6413 0.152939
R14549 gnd.n6415 gnd.n6414 0.152939
R14550 gnd.n6415 gnd.n1211 0.152939
R14551 gnd.n6449 gnd.n1211 0.152939
R14552 gnd.n6450 gnd.n6449 0.152939
R14553 gnd.n6451 gnd.n6450 0.152939
R14554 gnd.n6451 gnd.n1188 0.152939
R14555 gnd.n6483 gnd.n1188 0.152939
R14556 gnd.n6484 gnd.n6483 0.152939
R14557 gnd.n6485 gnd.n6484 0.152939
R14558 gnd.n6486 gnd.n6485 0.152939
R14559 gnd.n6487 gnd.n6486 0.152939
R14560 gnd.n6490 gnd.n6487 0.152939
R14561 gnd.n6491 gnd.n6490 0.152939
R14562 gnd.n6492 gnd.n6491 0.152939
R14563 gnd.n6492 gnd.n1129 0.152939
R14564 gnd.n6604 gnd.n1129 0.152939
R14565 gnd.n6605 gnd.n6604 0.152939
R14566 gnd.n6606 gnd.n6605 0.152939
R14567 gnd.n6607 gnd.n6606 0.152939
R14568 gnd.n6608 gnd.n6607 0.152939
R14569 gnd.n6608 gnd.n1090 0.152939
R14570 gnd.n6696 gnd.n1090 0.152939
R14571 gnd.n6697 gnd.n6696 0.152939
R14572 gnd.n6698 gnd.n6697 0.152939
R14573 gnd.n6698 gnd.n1067 0.152939
R14574 gnd.n6724 gnd.n1067 0.152939
R14575 gnd.n6725 gnd.n6724 0.152939
R14576 gnd.n6726 gnd.n6725 0.152939
R14577 gnd.n6727 gnd.n6726 0.152939
R14578 gnd.n6728 gnd.n6727 0.152939
R14579 gnd.n6729 gnd.n6728 0.152939
R14580 gnd.n6729 gnd.n1024 0.152939
R14581 gnd.n6807 gnd.n1024 0.152939
R14582 gnd.n6808 gnd.n6807 0.152939
R14583 gnd.n6809 gnd.n6808 0.152939
R14584 gnd.n6809 gnd.n996 0.152939
R14585 gnd.n6848 gnd.n996 0.152939
R14586 gnd.n6849 gnd.n6848 0.152939
R14587 gnd.n6850 gnd.n6849 0.152939
R14588 gnd.n6851 gnd.n6850 0.152939
R14589 gnd.n6852 gnd.n6851 0.152939
R14590 gnd.n6854 gnd.n6852 0.152939
R14591 gnd.n6855 gnd.n6854 0.152939
R14592 gnd.n6855 gnd.n714 0.152939
R14593 gnd.n7026 gnd.n714 0.152939
R14594 gnd.n7027 gnd.n7026 0.152939
R14595 gnd.n7028 gnd.n7027 0.152939
R14596 gnd.n7029 gnd.n7028 0.152939
R14597 gnd.n7029 gnd.n689 0.152939
R14598 gnd.n7061 gnd.n689 0.152939
R14599 gnd.n7062 gnd.n7061 0.152939
R14600 gnd.n7063 gnd.n7062 0.152939
R14601 gnd.n7065 gnd.n7063 0.152939
R14602 gnd.n7065 gnd.n7064 0.152939
R14603 gnd.n7064 gnd.n673 0.152939
R14604 gnd.n7085 gnd.n673 0.152939
R14605 gnd.n7086 gnd.n7085 0.152939
R14606 gnd.n7087 gnd.n7086 0.152939
R14607 gnd.n7088 gnd.n7087 0.152939
R14608 gnd.n7089 gnd.n7088 0.152939
R14609 gnd.n7100 gnd.n7089 0.152939
R14610 gnd.n7101 gnd.n7100 0.152939
R14611 gnd.n7102 gnd.n7101 0.152939
R14612 gnd.n7103 gnd.n7102 0.152939
R14613 gnd.n7105 gnd.n7103 0.152939
R14614 gnd.n7106 gnd.n7105 0.152939
R14615 gnd.n7107 gnd.n7106 0.152939
R14616 gnd.n7107 gnd.n480 0.152939
R14617 gnd.n7265 gnd.n480 0.152939
R14618 gnd.n7266 gnd.n7265 0.152939
R14619 gnd.n7267 gnd.n7266 0.152939
R14620 gnd.n7268 gnd.n7267 0.152939
R14621 gnd.n7268 gnd.n446 0.152939
R14622 gnd.n7311 gnd.n446 0.152939
R14623 gnd.n7312 gnd.n7311 0.152939
R14624 gnd.n7313 gnd.n7312 0.152939
R14625 gnd.n7314 gnd.n7313 0.152939
R14626 gnd.n7314 gnd.n411 0.152939
R14627 gnd.n7357 gnd.n411 0.152939
R14628 gnd.n7358 gnd.n7357 0.152939
R14629 gnd.n7359 gnd.n7358 0.152939
R14630 gnd.n7360 gnd.n7359 0.152939
R14631 gnd.n3170 gnd.n2204 0.152939
R14632 gnd.n3171 gnd.n3170 0.152939
R14633 gnd.n3172 gnd.n3171 0.152939
R14634 gnd.n3172 gnd.n2198 0.152939
R14635 gnd.n3180 gnd.n2198 0.152939
R14636 gnd.n3181 gnd.n3180 0.152939
R14637 gnd.n3182 gnd.n3181 0.152939
R14638 gnd.n3182 gnd.n2192 0.152939
R14639 gnd.n3190 gnd.n2192 0.152939
R14640 gnd.n3191 gnd.n3190 0.152939
R14641 gnd.n3192 gnd.n3191 0.152939
R14642 gnd.n3192 gnd.n2186 0.152939
R14643 gnd.n3200 gnd.n2186 0.152939
R14644 gnd.n3201 gnd.n3200 0.152939
R14645 gnd.n3202 gnd.n3201 0.152939
R14646 gnd.n3202 gnd.n2180 0.152939
R14647 gnd.n3210 gnd.n2180 0.152939
R14648 gnd.n3211 gnd.n3210 0.152939
R14649 gnd.n3212 gnd.n3211 0.152939
R14650 gnd.n3212 gnd.n2174 0.152939
R14651 gnd.n3220 gnd.n2174 0.152939
R14652 gnd.n3221 gnd.n3220 0.152939
R14653 gnd.n3222 gnd.n3221 0.152939
R14654 gnd.n3222 gnd.n2168 0.152939
R14655 gnd.n3230 gnd.n2168 0.152939
R14656 gnd.n3231 gnd.n3230 0.152939
R14657 gnd.n3232 gnd.n3231 0.152939
R14658 gnd.n3232 gnd.n2162 0.152939
R14659 gnd.n3240 gnd.n2162 0.152939
R14660 gnd.n3241 gnd.n3240 0.152939
R14661 gnd.n3242 gnd.n3241 0.152939
R14662 gnd.n3242 gnd.n2156 0.152939
R14663 gnd.n3250 gnd.n2156 0.152939
R14664 gnd.n3251 gnd.n3250 0.152939
R14665 gnd.n3252 gnd.n3251 0.152939
R14666 gnd.n3252 gnd.n2150 0.152939
R14667 gnd.n3260 gnd.n2150 0.152939
R14668 gnd.n3261 gnd.n3260 0.152939
R14669 gnd.n3262 gnd.n3261 0.152939
R14670 gnd.n3262 gnd.n2144 0.152939
R14671 gnd.n3270 gnd.n2144 0.152939
R14672 gnd.n3271 gnd.n3270 0.152939
R14673 gnd.n3272 gnd.n3271 0.152939
R14674 gnd.n3272 gnd.n2138 0.152939
R14675 gnd.n3280 gnd.n2138 0.152939
R14676 gnd.n3281 gnd.n3280 0.152939
R14677 gnd.n3282 gnd.n3281 0.152939
R14678 gnd.n3282 gnd.n2132 0.152939
R14679 gnd.n3290 gnd.n2132 0.152939
R14680 gnd.n3291 gnd.n3290 0.152939
R14681 gnd.n3292 gnd.n3291 0.152939
R14682 gnd.n3292 gnd.n2126 0.152939
R14683 gnd.n3300 gnd.n2126 0.152939
R14684 gnd.n3301 gnd.n3300 0.152939
R14685 gnd.n3302 gnd.n3301 0.152939
R14686 gnd.n3302 gnd.n2120 0.152939
R14687 gnd.n3310 gnd.n2120 0.152939
R14688 gnd.n3311 gnd.n3310 0.152939
R14689 gnd.n3312 gnd.n3311 0.152939
R14690 gnd.n3312 gnd.n2114 0.152939
R14691 gnd.n3320 gnd.n2114 0.152939
R14692 gnd.n3321 gnd.n3320 0.152939
R14693 gnd.n3322 gnd.n3321 0.152939
R14694 gnd.n3322 gnd.n2108 0.152939
R14695 gnd.n3330 gnd.n2108 0.152939
R14696 gnd.n3331 gnd.n3330 0.152939
R14697 gnd.n3332 gnd.n3331 0.152939
R14698 gnd.n3332 gnd.n2102 0.152939
R14699 gnd.n3340 gnd.n2102 0.152939
R14700 gnd.n3341 gnd.n3340 0.152939
R14701 gnd.n3342 gnd.n3341 0.152939
R14702 gnd.n3342 gnd.n2096 0.152939
R14703 gnd.n3350 gnd.n2096 0.152939
R14704 gnd.n3351 gnd.n3350 0.152939
R14705 gnd.n3352 gnd.n3351 0.152939
R14706 gnd.n3352 gnd.n2090 0.152939
R14707 gnd.n3360 gnd.n2090 0.152939
R14708 gnd.n3361 gnd.n3360 0.152939
R14709 gnd.n3362 gnd.n3361 0.152939
R14710 gnd.n3362 gnd.n2084 0.152939
R14711 gnd.n3370 gnd.n2084 0.152939
R14712 gnd.n3371 gnd.n3370 0.152939
R14713 gnd.n3372 gnd.n3371 0.152939
R14714 gnd.n3373 gnd.n3372 0.152939
R14715 gnd.n5506 gnd.n5503 0.152939
R14716 gnd.n5507 gnd.n5506 0.152939
R14717 gnd.n5508 gnd.n5507 0.152939
R14718 gnd.n5508 gnd.n5486 0.152939
R14719 gnd.n5525 gnd.n5486 0.152939
R14720 gnd.n5526 gnd.n5525 0.152939
R14721 gnd.n5527 gnd.n5526 0.152939
R14722 gnd.n5527 gnd.n5473 0.152939
R14723 gnd.n5546 gnd.n5473 0.152939
R14724 gnd.n5547 gnd.n5546 0.152939
R14725 gnd.n5555 gnd.n5547 0.152939
R14726 gnd.n5555 gnd.n5554 0.152939
R14727 gnd.n5554 gnd.n5553 0.152939
R14728 gnd.n5553 gnd.n5548 0.152939
R14729 gnd.n5549 gnd.n5548 0.152939
R14730 gnd.n5549 gnd.n1449 0.152939
R14731 gnd.n6034 gnd.n1449 0.152939
R14732 gnd.n6035 gnd.n6034 0.152939
R14733 gnd.n6043 gnd.n6035 0.152939
R14734 gnd.n6043 gnd.n6042 0.152939
R14735 gnd.n6042 gnd.n6041 0.152939
R14736 gnd.n6041 gnd.n6037 0.152939
R14737 gnd.n6037 gnd.n6036 0.152939
R14738 gnd.n6036 gnd.n1390 0.152939
R14739 gnd.n6143 gnd.n1390 0.152939
R14740 gnd.n6144 gnd.n6143 0.152939
R14741 gnd.n6149 gnd.n6144 0.152939
R14742 gnd.n6149 gnd.n6148 0.152939
R14743 gnd.n6148 gnd.n6147 0.152939
R14744 gnd.n6147 gnd.n1353 0.152939
R14745 gnd.n6211 gnd.n1353 0.152939
R14746 gnd.n6212 gnd.n6211 0.152939
R14747 gnd.n6214 gnd.n6212 0.152939
R14748 gnd.n6214 gnd.n6213 0.152939
R14749 gnd.n6213 gnd.n1297 0.152939
R14750 gnd.n6290 gnd.n1297 0.152939
R14751 gnd.n6291 gnd.n6290 0.152939
R14752 gnd.n6293 gnd.n6291 0.152939
R14753 gnd.n6293 gnd.n6292 0.152939
R14754 gnd.n6292 gnd.n1293 0.152939
R14755 gnd.n6300 gnd.n1293 0.152939
R14756 gnd.n6301 gnd.n6300 0.152939
R14757 gnd.n6302 gnd.n6301 0.152939
R14758 gnd.n6302 gnd.n1290 0.152939
R14759 gnd.n6308 gnd.n1290 0.152939
R14760 gnd.n6309 gnd.n6308 0.152939
R14761 gnd.n6341 gnd.n6309 0.152939
R14762 gnd.n6341 gnd.n6340 0.152939
R14763 gnd.n6340 gnd.n6339 0.152939
R14764 gnd.n6339 gnd.n6310 0.152939
R14765 gnd.n6335 gnd.n6310 0.152939
R14766 gnd.n6335 gnd.n6334 0.152939
R14767 gnd.n6334 gnd.n6333 0.152939
R14768 gnd.n6333 gnd.n6314 0.152939
R14769 gnd.n6329 gnd.n6314 0.152939
R14770 gnd.n6329 gnd.n6328 0.152939
R14771 gnd.n6328 gnd.n6327 0.152939
R14772 gnd.n6327 gnd.n1153 0.152939
R14773 gnd.n6541 gnd.n1153 0.152939
R14774 gnd.n6542 gnd.n6541 0.152939
R14775 gnd.n6557 gnd.n6542 0.152939
R14776 gnd.n6557 gnd.n6556 0.152939
R14777 gnd.n6556 gnd.n6555 0.152939
R14778 gnd.n6555 gnd.n6543 0.152939
R14779 gnd.n6551 gnd.n6543 0.152939
R14780 gnd.n6551 gnd.n6550 0.152939
R14781 gnd.n6550 gnd.n6549 0.152939
R14782 gnd.n6549 gnd.n1105 0.152939
R14783 gnd.n6644 gnd.n1105 0.152939
R14784 gnd.n6645 gnd.n6644 0.152939
R14785 gnd.n6646 gnd.n6645 0.152939
R14786 gnd.n6646 gnd.n1101 0.152939
R14787 gnd.n6651 gnd.n1101 0.152939
R14788 gnd.n6652 gnd.n6651 0.152939
R14789 gnd.n6669 gnd.n6652 0.152939
R14790 gnd.n6669 gnd.n6668 0.152939
R14791 gnd.n6668 gnd.n6667 0.152939
R14792 gnd.n6667 gnd.n6653 0.152939
R14793 gnd.n6663 gnd.n6653 0.152939
R14794 gnd.n6663 gnd.n6662 0.152939
R14795 gnd.n6662 gnd.n6661 0.152939
R14796 gnd.n6661 gnd.n1011 0.152939
R14797 gnd.n6827 gnd.n1011 0.152939
R14798 gnd.n6828 gnd.n6827 0.152939
R14799 gnd.n6832 gnd.n6828 0.152939
R14800 gnd.n6832 gnd.n6831 0.152939
R14801 gnd.n6831 gnd.n6830 0.152939
R14802 gnd.n6830 gnd.n721 0.152939
R14803 gnd.n7016 gnd.n721 0.152939
R14804 gnd.n7017 gnd.n7016 0.152939
R14805 gnd.n7019 gnd.n7017 0.152939
R14806 gnd.n7019 gnd.n7018 0.152939
R14807 gnd.n7018 gnd.n696 0.152939
R14808 gnd.n7046 gnd.n696 0.152939
R14809 gnd.n7047 gnd.n7046 0.152939
R14810 gnd.n7054 gnd.n7047 0.152939
R14811 gnd.n7054 gnd.n7053 0.152939
R14812 gnd.n7053 gnd.n7052 0.152939
R14813 gnd.n7052 gnd.n7048 0.152939
R14814 gnd.n7048 gnd.n581 0.152939
R14815 gnd.n7188 gnd.n581 0.152939
R14816 gnd.n5264 gnd.n1854 0.152939
R14817 gnd.n5265 gnd.n5264 0.152939
R14818 gnd.n5267 gnd.n5265 0.152939
R14819 gnd.n5267 gnd.n5266 0.152939
R14820 gnd.n5266 gnd.n1818 0.152939
R14821 gnd.n5306 gnd.n1818 0.152939
R14822 gnd.n5307 gnd.n5306 0.152939
R14823 gnd.n5309 gnd.n5307 0.152939
R14824 gnd.n5309 gnd.n5308 0.152939
R14825 gnd.n5308 gnd.n1783 0.152939
R14826 gnd.n5346 gnd.n1783 0.152939
R14827 gnd.n5347 gnd.n5346 0.152939
R14828 gnd.n5349 gnd.n5347 0.152939
R14829 gnd.n5349 gnd.n5348 0.152939
R14830 gnd.n5348 gnd.n1748 0.152939
R14831 gnd.n5394 gnd.n1748 0.152939
R14832 gnd.n5395 gnd.n5394 0.152939
R14833 gnd.n5400 gnd.n5395 0.152939
R14834 gnd.n5400 gnd.n5399 0.152939
R14835 gnd.n5399 gnd.n5398 0.152939
R14836 gnd.n5398 gnd.n1678 0.152939
R14837 gnd.n5749 gnd.n1678 0.152939
R14838 gnd.n5749 gnd.n5748 0.152939
R14839 gnd.n5748 gnd.n5747 0.152939
R14840 gnd.n5747 gnd.n1679 0.152939
R14841 gnd.n5743 gnd.n1679 0.152939
R14842 gnd.n5731 gnd.n1706 0.152939
R14843 gnd.n5731 gnd.n5730 0.152939
R14844 gnd.n5730 gnd.n5729 0.152939
R14845 gnd.n5729 gnd.n1708 0.152939
R14846 gnd.n5725 gnd.n1708 0.152939
R14847 gnd.n5725 gnd.n5724 0.152939
R14848 gnd.n5577 gnd.n5455 0.152939
R14849 gnd.n5577 gnd.n5576 0.152939
R14850 gnd.n5576 gnd.n5575 0.152939
R14851 gnd.n5575 gnd.n5456 0.152939
R14852 gnd.n5571 gnd.n5456 0.152939
R14853 gnd.n5571 gnd.n5570 0.152939
R14854 gnd.n5570 gnd.n5569 0.152939
R14855 gnd.n5569 gnd.n5461 0.152939
R14856 gnd.n5565 gnd.n5461 0.152939
R14857 gnd.n5565 gnd.n5564 0.152939
R14858 gnd.n5564 gnd.n5563 0.152939
R14859 gnd.n5563 gnd.n5466 0.152939
R14860 gnd.n5466 gnd.n1455 0.152939
R14861 gnd.n6025 gnd.n1455 0.152939
R14862 gnd.n6026 gnd.n6025 0.152939
R14863 gnd.n6027 gnd.n6026 0.152939
R14864 gnd.n6027 gnd.n1424 0.152939
R14865 gnd.n6084 gnd.n1424 0.152939
R14866 gnd.n6085 gnd.n6084 0.152939
R14867 gnd.n6086 gnd.n6085 0.152939
R14868 gnd.n6086 gnd.n1396 0.152939
R14869 gnd.n6134 gnd.n1396 0.152939
R14870 gnd.n6135 gnd.n6134 0.152939
R14871 gnd.n6136 gnd.n6135 0.152939
R14872 gnd.n6136 gnd.n1369 0.152939
R14873 gnd.n6179 gnd.n1369 0.152939
R14874 gnd.n6180 gnd.n6179 0.152939
R14875 gnd.n6181 gnd.n6180 0.152939
R14876 gnd.n6181 gnd.n1338 0.152939
R14877 gnd.n6230 gnd.n1338 0.152939
R14878 gnd.n6231 gnd.n6230 0.152939
R14879 gnd.n6232 gnd.n6231 0.152939
R14880 gnd.n6232 gnd.n1305 0.152939
R14881 gnd.n6275 gnd.n1305 0.152939
R14882 gnd.n6276 gnd.n6275 0.152939
R14883 gnd.n6284 gnd.n6276 0.152939
R14884 gnd.n6284 gnd.n6283 0.152939
R14885 gnd.n6283 gnd.n6282 0.152939
R14886 gnd.n6282 gnd.n6277 0.152939
R14887 gnd.n6277 gnd.n1259 0.152939
R14888 gnd.n6394 gnd.n1259 0.152939
R14889 gnd.n6395 gnd.n6394 0.152939
R14890 gnd.n6397 gnd.n6395 0.152939
R14891 gnd.n6397 gnd.n6396 0.152939
R14892 gnd.n6396 gnd.n1228 0.152939
R14893 gnd.n6430 gnd.n1228 0.152939
R14894 gnd.n6431 gnd.n6430 0.152939
R14895 gnd.n6433 gnd.n6431 0.152939
R14896 gnd.n6433 gnd.n6432 0.152939
R14897 gnd.n6432 gnd.n1203 0.152939
R14898 gnd.n6459 gnd.n1203 0.152939
R14899 gnd.n6460 gnd.n6459 0.152939
R14900 gnd.n6461 gnd.n6460 0.152939
R14901 gnd.n6461 gnd.n1173 0.152939
R14902 gnd.n6516 gnd.n1173 0.152939
R14903 gnd.n6517 gnd.n6516 0.152939
R14904 gnd.n6519 gnd.n6517 0.152939
R14905 gnd.n6519 gnd.n6518 0.152939
R14906 gnd.n6518 gnd.n1138 0.152939
R14907 gnd.n6582 gnd.n1138 0.152939
R14908 gnd.n6583 gnd.n6582 0.152939
R14909 gnd.n6597 gnd.n6583 0.152939
R14910 gnd.n6597 gnd.n6596 0.152939
R14911 gnd.n6596 gnd.n6595 0.152939
R14912 gnd.n6595 gnd.n6584 0.152939
R14913 gnd.n6591 gnd.n6584 0.152939
R14914 gnd.n6591 gnd.n6590 0.152939
R14915 gnd.n6590 gnd.n1082 0.152939
R14916 gnd.n6705 gnd.n1082 0.152939
R14917 gnd.n6706 gnd.n6705 0.152939
R14918 gnd.n6708 gnd.n6706 0.152939
R14919 gnd.n6708 gnd.n6707 0.152939
R14920 gnd.n6707 gnd.n1052 0.152939
R14921 gnd.n6750 gnd.n1052 0.152939
R14922 gnd.n6751 gnd.n6750 0.152939
R14923 gnd.n6753 gnd.n6751 0.152939
R14924 gnd.n6753 gnd.n6752 0.152939
R14925 gnd.n6752 gnd.n1034 0.152939
R14926 gnd.n6800 gnd.n1034 0.152939
R14927 gnd.n6800 gnd.n6799 0.152939
R14928 gnd.n6799 gnd.n6798 0.152939
R14929 gnd.n6798 gnd.n1006 0.152939
R14930 gnd.n6841 gnd.n1006 0.152939
R14931 gnd.n6841 gnd.n6840 0.152939
R14932 gnd.n6840 gnd.n6839 0.152939
R14933 gnd.n6839 gnd.n731 0.152939
R14934 gnd.n7007 gnd.n731 0.152939
R14935 gnd.n7008 gnd.n7007 0.152939
R14936 gnd.n7010 gnd.n7008 0.152939
R14937 gnd.n7010 gnd.n7009 0.152939
R14938 gnd.n7009 gnd.n705 0.152939
R14939 gnd.n7037 gnd.n705 0.152939
R14940 gnd.n7038 gnd.n7037 0.152939
R14941 gnd.n7040 gnd.n7038 0.152939
R14942 gnd.n7040 gnd.n7039 0.152939
R14943 gnd.n7039 gnd.n681 0.152939
R14944 gnd.n7073 gnd.n681 0.152939
R14945 gnd.n7074 gnd.n7073 0.152939
R14946 gnd.n7075 gnd.n7074 0.152939
R14947 gnd.n7075 gnd.n589 0.152939
R14948 gnd.n7182 gnd.n589 0.152939
R14949 gnd.n7181 gnd.n590 0.152939
R14950 gnd.n7177 gnd.n590 0.152939
R14951 gnd.n7177 gnd.n7176 0.152939
R14952 gnd.n7176 gnd.n7175 0.152939
R14953 gnd.n7175 gnd.n594 0.152939
R14954 gnd.n7171 gnd.n594 0.152939
R14955 gnd.n7218 gnd.n7217 0.152939
R14956 gnd.n7220 gnd.n7218 0.152939
R14957 gnd.n7220 gnd.n7219 0.152939
R14958 gnd.n7219 gnd.n488 0.152939
R14959 gnd.n7254 gnd.n488 0.152939
R14960 gnd.n7255 gnd.n7254 0.152939
R14961 gnd.n7257 gnd.n7255 0.152939
R14962 gnd.n7257 gnd.n7256 0.152939
R14963 gnd.n7256 gnd.n454 0.152939
R14964 gnd.n7300 gnd.n454 0.152939
R14965 gnd.n7301 gnd.n7300 0.152939
R14966 gnd.n7303 gnd.n7301 0.152939
R14967 gnd.n7303 gnd.n7302 0.152939
R14968 gnd.n7302 gnd.n419 0.152939
R14969 gnd.n7347 gnd.n419 0.152939
R14970 gnd.n7348 gnd.n7347 0.152939
R14971 gnd.n7350 gnd.n7348 0.152939
R14972 gnd.n7350 gnd.n7349 0.152939
R14973 gnd.n7349 gnd.n387 0.152939
R14974 gnd.n7391 gnd.n387 0.152939
R14975 gnd.n7392 gnd.n7391 0.152939
R14976 gnd.n7399 gnd.n7392 0.152939
R14977 gnd.n7399 gnd.n7398 0.152939
R14978 gnd.n7398 gnd.n7397 0.152939
R14979 gnd.n7397 gnd.n7393 0.152939
R14980 gnd.n7393 gnd.n83 0.152939
R14981 gnd.n5724 gnd.n1649 0.128549
R14982 gnd.n7171 gnd.n7170 0.128549
R14983 gnd.n4172 gnd.n4171 0.0767195
R14984 gnd.n4171 gnd.n4170 0.0767195
R14985 gnd.n7748 gnd.n96 0.0767195
R14986 gnd.n7748 gnd.n97 0.0767195
R14987 gnd.n5297 gnd.n5296 0.0767195
R14988 gnd.n5296 gnd.n1828 0.0767195
R14989 gnd.n7758 gnd.n7757 0.0695946
R14990 gnd.n5217 gnd.n5216 0.0695946
R14991 gnd.n5216 gnd.n1854 0.0695946
R14992 gnd.n7758 gnd.n83 0.0695946
R14993 gnd.n5869 gnd.n1649 0.063
R14994 gnd.n7170 gnd.n599 0.063
R14995 gnd.n4738 gnd.n2033 0.0477147
R14996 gnd.n7093 gnd.n599 0.0477147
R14997 gnd.n7566 gnd.n206 0.0477147
R14998 gnd.n4970 gnd.n1986 0.0477147
R14999 gnd.n5869 gnd.n5868 0.0477147
R15000 gnd.n3935 gnd.n3823 0.0442063
R15001 gnd.n3936 gnd.n3935 0.0442063
R15002 gnd.n3937 gnd.n3936 0.0442063
R15003 gnd.n3937 gnd.n3812 0.0442063
R15004 gnd.n3951 gnd.n3812 0.0442063
R15005 gnd.n3952 gnd.n3951 0.0442063
R15006 gnd.n3953 gnd.n3952 0.0442063
R15007 gnd.n3953 gnd.n3799 0.0442063
R15008 gnd.n3997 gnd.n3799 0.0442063
R15009 gnd.n3998 gnd.n3997 0.0442063
R15010 gnd.n4000 gnd.n3733 0.0344674
R15011 gnd.n7094 gnd.n7093 0.0344674
R15012 gnd.n7094 gnd.n513 0.0344674
R15013 gnd.n513 gnd.n508 0.0344674
R15014 gnd.n509 gnd.n508 0.0344674
R15015 gnd.n510 gnd.n509 0.0344674
R15016 gnd.n7234 gnd.n510 0.0344674
R15017 gnd.n7234 gnd.n511 0.0344674
R15018 gnd.n511 gnd.n473 0.0344674
R15019 gnd.n474 gnd.n473 0.0344674
R15020 gnd.n475 gnd.n474 0.0344674
R15021 gnd.n7280 gnd.n475 0.0344674
R15022 gnd.n7280 gnd.n476 0.0344674
R15023 gnd.n476 gnd.n438 0.0344674
R15024 gnd.n439 gnd.n438 0.0344674
R15025 gnd.n440 gnd.n439 0.0344674
R15026 gnd.n441 gnd.n440 0.0344674
R15027 gnd.n7323 gnd.n441 0.0344674
R15028 gnd.n7323 gnd.n405 0.0344674
R15029 gnd.n406 gnd.n405 0.0344674
R15030 gnd.n7369 gnd.n406 0.0344674
R15031 gnd.n7370 gnd.n7369 0.0344674
R15032 gnd.n7370 gnd.n380 0.0344674
R15033 gnd.n7408 gnd.n380 0.0344674
R15034 gnd.n7408 gnd.n367 0.0344674
R15035 gnd.n7422 gnd.n367 0.0344674
R15036 gnd.n7423 gnd.n7422 0.0344674
R15037 gnd.n7423 gnd.n362 0.0344674
R15038 gnd.n362 gnd.n360 0.0344674
R15039 gnd.n7434 gnd.n360 0.0344674
R15040 gnd.n7435 gnd.n7434 0.0344674
R15041 gnd.n7435 gnd.n111 0.0344674
R15042 gnd.n112 gnd.n111 0.0344674
R15043 gnd.n113 gnd.n112 0.0344674
R15044 gnd.n7479 gnd.n113 0.0344674
R15045 gnd.n7479 gnd.n128 0.0344674
R15046 gnd.n129 gnd.n128 0.0344674
R15047 gnd.n130 gnd.n129 0.0344674
R15048 gnd.n7486 gnd.n130 0.0344674
R15049 gnd.n7486 gnd.n148 0.0344674
R15050 gnd.n149 gnd.n148 0.0344674
R15051 gnd.n150 gnd.n149 0.0344674
R15052 gnd.n7493 gnd.n150 0.0344674
R15053 gnd.n7493 gnd.n166 0.0344674
R15054 gnd.n167 gnd.n166 0.0344674
R15055 gnd.n168 gnd.n167 0.0344674
R15056 gnd.n7497 gnd.n168 0.0344674
R15057 gnd.n7497 gnd.n186 0.0344674
R15058 gnd.n187 gnd.n186 0.0344674
R15059 gnd.n188 gnd.n187 0.0344674
R15060 gnd.n7498 gnd.n188 0.0344674
R15061 gnd.n7498 gnd.n204 0.0344674
R15062 gnd.n205 gnd.n204 0.0344674
R15063 gnd.n206 gnd.n205 0.0344674
R15064 gnd.n5095 gnd.n1986 0.0344674
R15065 gnd.n5095 gnd.n1989 0.0344674
R15066 gnd.n1989 gnd.n1988 0.0344674
R15067 gnd.n1988 gnd.n1969 0.0344674
R15068 gnd.n1969 gnd.n1967 0.0344674
R15069 gnd.n5112 gnd.n1967 0.0344674
R15070 gnd.n5113 gnd.n5112 0.0344674
R15071 gnd.n5113 gnd.n1951 0.0344674
R15072 gnd.n1951 gnd.n1949 0.0344674
R15073 gnd.n5132 gnd.n1949 0.0344674
R15074 gnd.n5133 gnd.n5132 0.0344674
R15075 gnd.n5133 gnd.n1933 0.0344674
R15076 gnd.n1933 gnd.n1930 0.0344674
R15077 gnd.n1931 gnd.n1930 0.0344674
R15078 gnd.n5154 gnd.n1931 0.0344674
R15079 gnd.n5155 gnd.n5154 0.0344674
R15080 gnd.n5155 gnd.n1907 0.0344674
R15081 gnd.n1907 gnd.n1904 0.0344674
R15082 gnd.n1905 gnd.n1904 0.0344674
R15083 gnd.n5189 gnd.n1905 0.0344674
R15084 gnd.n5190 gnd.n5189 0.0344674
R15085 gnd.n5190 gnd.n1882 0.0344674
R15086 gnd.n1882 gnd.n1880 0.0344674
R15087 gnd.n5231 gnd.n1880 0.0344674
R15088 gnd.n5232 gnd.n5231 0.0344674
R15089 gnd.n5232 gnd.n1868 0.0344674
R15090 gnd.n1868 gnd.n1866 0.0344674
R15091 gnd.n5248 gnd.n1866 0.0344674
R15092 gnd.n5249 gnd.n5248 0.0344674
R15093 gnd.n5249 gnd.n1848 0.0344674
R15094 gnd.n1848 gnd.n1843 0.0344674
R15095 gnd.n1844 gnd.n1843 0.0344674
R15096 gnd.n1845 gnd.n1844 0.0344674
R15097 gnd.n5286 gnd.n1845 0.0344674
R15098 gnd.n5286 gnd.n1846 0.0344674
R15099 gnd.n1846 gnd.n1802 0.0344674
R15100 gnd.n1803 gnd.n1802 0.0344674
R15101 gnd.n1804 gnd.n1803 0.0344674
R15102 gnd.n1805 gnd.n1804 0.0344674
R15103 gnd.n1805 gnd.n1777 0.0344674
R15104 gnd.n1777 gnd.n1766 0.0344674
R15105 gnd.n1767 gnd.n1766 0.0344674
R15106 gnd.n1768 gnd.n1767 0.0344674
R15107 gnd.n1769 gnd.n1768 0.0344674
R15108 gnd.n1769 gnd.n1742 0.0344674
R15109 gnd.n1742 gnd.n1740 0.0344674
R15110 gnd.n5409 gnd.n1740 0.0344674
R15111 gnd.n5410 gnd.n5409 0.0344674
R15112 gnd.n5410 gnd.n1671 0.0344674
R15113 gnd.n5756 gnd.n1671 0.0344674
R15114 gnd.n5757 gnd.n5756 0.0344674
R15115 gnd.n5757 gnd.n1650 0.0344674
R15116 gnd.n5868 gnd.n1650 0.0344674
R15117 gnd.n5721 gnd.n5720 0.0343753
R15118 gnd.n7169 gnd.n7168 0.0343753
R15119 gnd.n5742 gnd.n5741 0.0296328
R15120 gnd.n7192 gnd.n518 0.0296328
R15121 gnd.n4020 gnd.n4019 0.0269946
R15122 gnd.n4022 gnd.n4021 0.0269946
R15123 gnd.n3728 gnd.n3726 0.0269946
R15124 gnd.n4032 gnd.n4030 0.0269946
R15125 gnd.n4031 gnd.n3707 0.0269946
R15126 gnd.n4051 gnd.n4050 0.0269946
R15127 gnd.n4053 gnd.n4052 0.0269946
R15128 gnd.n3702 gnd.n3701 0.0269946
R15129 gnd.n4063 gnd.n3697 0.0269946
R15130 gnd.n4062 gnd.n3699 0.0269946
R15131 gnd.n3698 gnd.n3680 0.0269946
R15132 gnd.n4083 gnd.n3681 0.0269946
R15133 gnd.n4082 gnd.n3682 0.0269946
R15134 gnd.n4116 gnd.n3657 0.0269946
R15135 gnd.n4118 gnd.n4117 0.0269946
R15136 gnd.n4119 gnd.n3604 0.0269946
R15137 gnd.n3652 gnd.n3605 0.0269946
R15138 gnd.n3654 gnd.n3606 0.0269946
R15139 gnd.n4129 gnd.n4128 0.0269946
R15140 gnd.n4131 gnd.n4130 0.0269946
R15141 gnd.n4132 gnd.n3626 0.0269946
R15142 gnd.n4134 gnd.n3627 0.0269946
R15143 gnd.n4137 gnd.n3628 0.0269946
R15144 gnd.n4140 gnd.n4139 0.0269946
R15145 gnd.n4142 gnd.n4141 0.0269946
R15146 gnd.n4207 gnd.n3511 0.0269946
R15147 gnd.n4209 gnd.n4208 0.0269946
R15148 gnd.n4218 gnd.n3504 0.0269946
R15149 gnd.n4220 gnd.n4219 0.0269946
R15150 gnd.n4221 gnd.n3502 0.0269946
R15151 gnd.n4228 gnd.n4224 0.0269946
R15152 gnd.n4227 gnd.n4226 0.0269946
R15153 gnd.n4225 gnd.n3481 0.0269946
R15154 gnd.n4250 gnd.n3482 0.0269946
R15155 gnd.n4249 gnd.n3483 0.0269946
R15156 gnd.n4292 gnd.n3456 0.0269946
R15157 gnd.n4294 gnd.n4293 0.0269946
R15158 gnd.n4303 gnd.n3449 0.0269946
R15159 gnd.n4305 gnd.n4304 0.0269946
R15160 gnd.n4306 gnd.n3447 0.0269946
R15161 gnd.n4313 gnd.n4309 0.0269946
R15162 gnd.n4312 gnd.n4311 0.0269946
R15163 gnd.n4310 gnd.n3426 0.0269946
R15164 gnd.n4335 gnd.n3427 0.0269946
R15165 gnd.n4334 gnd.n3428 0.0269946
R15166 gnd.n4381 gnd.n3402 0.0269946
R15167 gnd.n4383 gnd.n4382 0.0269946
R15168 gnd.n4392 gnd.n3395 0.0269946
R15169 gnd.n4651 gnd.n3393 0.0269946
R15170 gnd.n4656 gnd.n4654 0.0269946
R15171 gnd.n4655 gnd.n2069 0.0269946
R15172 gnd.n4680 gnd.n4679 0.0269946
R15173 gnd.n5719 gnd.n1715 0.022519
R15174 gnd.n5716 gnd.n5715 0.022519
R15175 gnd.n5712 gnd.n5601 0.022519
R15176 gnd.n5711 gnd.n5608 0.022519
R15177 gnd.n5708 gnd.n5707 0.022519
R15178 gnd.n5704 gnd.n5615 0.022519
R15179 gnd.n5703 gnd.n5621 0.022519
R15180 gnd.n5700 gnd.n5699 0.022519
R15181 gnd.n5696 gnd.n5627 0.022519
R15182 gnd.n5695 gnd.n5631 0.022519
R15183 gnd.n5692 gnd.n5691 0.022519
R15184 gnd.n5688 gnd.n5638 0.022519
R15185 gnd.n5687 gnd.n5644 0.022519
R15186 gnd.n5684 gnd.n5683 0.022519
R15187 gnd.n5680 gnd.n5650 0.022519
R15188 gnd.n5679 gnd.n5654 0.022519
R15189 gnd.n5676 gnd.n5675 0.022519
R15190 gnd.n5668 gnd.n5667 0.022519
R15191 gnd.n5741 gnd.n1684 0.022519
R15192 gnd.n7165 gnd.n600 0.022519
R15193 gnd.n7164 gnd.n604 0.022519
R15194 gnd.n7161 gnd.n7160 0.022519
R15195 gnd.n7157 gnd.n610 0.022519
R15196 gnd.n7156 gnd.n614 0.022519
R15197 gnd.n7153 gnd.n7152 0.022519
R15198 gnd.n7149 gnd.n620 0.022519
R15199 gnd.n7148 gnd.n624 0.022519
R15200 gnd.n7145 gnd.n7144 0.022519
R15201 gnd.n7141 gnd.n628 0.022519
R15202 gnd.n7140 gnd.n632 0.022519
R15203 gnd.n7137 gnd.n7136 0.022519
R15204 gnd.n7133 gnd.n638 0.022519
R15205 gnd.n7132 gnd.n642 0.022519
R15206 gnd.n7129 gnd.n7128 0.022519
R15207 gnd.n645 gnd.n572 0.022519
R15208 gnd.n7199 gnd.n7198 0.022519
R15209 gnd.n7195 gnd.n573 0.022519
R15210 gnd.n7194 gnd.n7192 0.022519
R15211 gnd.n7189 gnd.n518 0.0218415
R15212 gnd.n5742 gnd.n1683 0.0218415
R15213 gnd.n4000 gnd.n3999 0.0202011
R15214 gnd.n3999 gnd.n3998 0.0148637
R15215 gnd.n4649 gnd.n4393 0.0144266
R15216 gnd.n4650 gnd.n4649 0.0130679
R15217 gnd.n5720 gnd.n5719 0.0123564
R15218 gnd.n5716 gnd.n1715 0.0123564
R15219 gnd.n5715 gnd.n5601 0.0123564
R15220 gnd.n5712 gnd.n5711 0.0123564
R15221 gnd.n5708 gnd.n5608 0.0123564
R15222 gnd.n5707 gnd.n5615 0.0123564
R15223 gnd.n5704 gnd.n5703 0.0123564
R15224 gnd.n5700 gnd.n5621 0.0123564
R15225 gnd.n5699 gnd.n5627 0.0123564
R15226 gnd.n5696 gnd.n5695 0.0123564
R15227 gnd.n5692 gnd.n5631 0.0123564
R15228 gnd.n5691 gnd.n5638 0.0123564
R15229 gnd.n5688 gnd.n5687 0.0123564
R15230 gnd.n5684 gnd.n5644 0.0123564
R15231 gnd.n5683 gnd.n5650 0.0123564
R15232 gnd.n5680 gnd.n5679 0.0123564
R15233 gnd.n5676 gnd.n5654 0.0123564
R15234 gnd.n5675 gnd.n5668 0.0123564
R15235 gnd.n5667 gnd.n1684 0.0123564
R15236 gnd.n7168 gnd.n600 0.0123564
R15237 gnd.n7165 gnd.n7164 0.0123564
R15238 gnd.n7161 gnd.n604 0.0123564
R15239 gnd.n7160 gnd.n610 0.0123564
R15240 gnd.n7157 gnd.n7156 0.0123564
R15241 gnd.n7153 gnd.n614 0.0123564
R15242 gnd.n7152 gnd.n620 0.0123564
R15243 gnd.n7149 gnd.n7148 0.0123564
R15244 gnd.n7145 gnd.n624 0.0123564
R15245 gnd.n7144 gnd.n628 0.0123564
R15246 gnd.n7141 gnd.n7140 0.0123564
R15247 gnd.n7137 gnd.n632 0.0123564
R15248 gnd.n7136 gnd.n638 0.0123564
R15249 gnd.n7133 gnd.n7132 0.0123564
R15250 gnd.n7129 gnd.n642 0.0123564
R15251 gnd.n7128 gnd.n645 0.0123564
R15252 gnd.n7199 gnd.n572 0.0123564
R15253 gnd.n7198 gnd.n573 0.0123564
R15254 gnd.n7195 gnd.n7194 0.0123564
R15255 gnd.n4019 gnd.n3733 0.00797283
R15256 gnd.n4021 gnd.n4020 0.00797283
R15257 gnd.n4022 gnd.n3728 0.00797283
R15258 gnd.n4030 gnd.n3726 0.00797283
R15259 gnd.n4032 gnd.n4031 0.00797283
R15260 gnd.n4050 gnd.n3707 0.00797283
R15261 gnd.n4052 gnd.n4051 0.00797283
R15262 gnd.n4053 gnd.n3702 0.00797283
R15263 gnd.n3701 gnd.n3697 0.00797283
R15264 gnd.n4063 gnd.n4062 0.00797283
R15265 gnd.n3699 gnd.n3698 0.00797283
R15266 gnd.n3681 gnd.n3680 0.00797283
R15267 gnd.n4083 gnd.n4082 0.00797283
R15268 gnd.n3682 gnd.n3657 0.00797283
R15269 gnd.n4117 gnd.n4116 0.00797283
R15270 gnd.n4119 gnd.n4118 0.00797283
R15271 gnd.n3652 gnd.n3604 0.00797283
R15272 gnd.n3654 gnd.n3605 0.00797283
R15273 gnd.n4128 gnd.n3606 0.00797283
R15274 gnd.n4130 gnd.n4129 0.00797283
R15275 gnd.n4132 gnd.n4131 0.00797283
R15276 gnd.n4134 gnd.n3626 0.00797283
R15277 gnd.n4137 gnd.n3627 0.00797283
R15278 gnd.n4139 gnd.n3628 0.00797283
R15279 gnd.n4142 gnd.n4140 0.00797283
R15280 gnd.n4141 gnd.n3511 0.00797283
R15281 gnd.n4209 gnd.n4207 0.00797283
R15282 gnd.n4208 gnd.n3504 0.00797283
R15283 gnd.n4219 gnd.n4218 0.00797283
R15284 gnd.n4221 gnd.n4220 0.00797283
R15285 gnd.n4224 gnd.n3502 0.00797283
R15286 gnd.n4228 gnd.n4227 0.00797283
R15287 gnd.n4226 gnd.n4225 0.00797283
R15288 gnd.n3482 gnd.n3481 0.00797283
R15289 gnd.n4250 gnd.n4249 0.00797283
R15290 gnd.n3483 gnd.n3456 0.00797283
R15291 gnd.n4294 gnd.n4292 0.00797283
R15292 gnd.n4293 gnd.n3449 0.00797283
R15293 gnd.n4304 gnd.n4303 0.00797283
R15294 gnd.n4306 gnd.n4305 0.00797283
R15295 gnd.n4309 gnd.n3447 0.00797283
R15296 gnd.n4313 gnd.n4312 0.00797283
R15297 gnd.n4311 gnd.n4310 0.00797283
R15298 gnd.n3427 gnd.n3426 0.00797283
R15299 gnd.n4335 gnd.n4334 0.00797283
R15300 gnd.n3428 gnd.n3402 0.00797283
R15301 gnd.n4383 gnd.n4381 0.00797283
R15302 gnd.n4382 gnd.n3395 0.00797283
R15303 gnd.n4393 gnd.n4392 0.00797283
R15304 gnd.n4651 gnd.n4650 0.00797283
R15305 gnd.n4654 gnd.n3393 0.00797283
R15306 gnd.n4656 gnd.n4655 0.00797283
R15307 gnd.n4679 gnd.n2069 0.00797283
R15308 gnd.n4680 gnd.n2033 0.00797283
R15309 gnd.n5721 gnd.n1649 0.00592005
R15310 gnd.n7170 gnd.n7169 0.00592005
R15311 a_n6972_8799.n178 a_n6972_8799.t58 485.149
R15312 a_n6972_8799.n194 a_n6972_8799.t70 485.149
R15313 a_n6972_8799.n211 a_n6972_8799.t118 485.149
R15314 a_n6972_8799.n127 a_n6972_8799.t114 485.149
R15315 a_n6972_8799.n143 a_n6972_8799.t125 485.149
R15316 a_n6972_8799.n160 a_n6972_8799.t117 485.149
R15317 a_n6972_8799.n188 a_n6972_8799.t79 464.166
R15318 a_n6972_8799.n187 a_n6972_8799.t78 464.166
R15319 a_n6972_8799.n173 a_n6972_8799.t56 464.166
R15320 a_n6972_8799.n186 a_n6972_8799.t115 464.166
R15321 a_n6972_8799.n185 a_n6972_8799.t80 464.166
R15322 a_n6972_8799.n174 a_n6972_8799.t62 464.166
R15323 a_n6972_8799.n184 a_n6972_8799.t119 464.166
R15324 a_n6972_8799.n183 a_n6972_8799.t94 464.166
R15325 a_n6972_8799.n175 a_n6972_8799.t92 464.166
R15326 a_n6972_8799.n182 a_n6972_8799.t39 464.166
R15327 a_n6972_8799.n181 a_n6972_8799.t98 464.166
R15328 a_n6972_8799.n176 a_n6972_8799.t97 464.166
R15329 a_n6972_8799.n180 a_n6972_8799.t41 464.166
R15330 a_n6972_8799.n179 a_n6972_8799.t40 464.166
R15331 a_n6972_8799.n177 a_n6972_8799.t111 464.166
R15332 a_n6972_8799.n204 a_n6972_8799.t86 464.166
R15333 a_n6972_8799.n203 a_n6972_8799.t85 464.166
R15334 a_n6972_8799.n189 a_n6972_8799.t69 464.166
R15335 a_n6972_8799.n202 a_n6972_8799.t127 464.166
R15336 a_n6972_8799.n201 a_n6972_8799.t91 464.166
R15337 a_n6972_8799.n190 a_n6972_8799.t71 464.166
R15338 a_n6972_8799.n200 a_n6972_8799.t131 464.166
R15339 a_n6972_8799.n199 a_n6972_8799.t104 464.166
R15340 a_n6972_8799.n191 a_n6972_8799.t103 464.166
R15341 a_n6972_8799.n198 a_n6972_8799.t48 464.166
R15342 a_n6972_8799.n197 a_n6972_8799.t107 464.166
R15343 a_n6972_8799.n192 a_n6972_8799.t106 464.166
R15344 a_n6972_8799.n196 a_n6972_8799.t52 464.166
R15345 a_n6972_8799.n195 a_n6972_8799.t51 464.166
R15346 a_n6972_8799.n193 a_n6972_8799.t122 464.166
R15347 a_n6972_8799.n221 a_n6972_8799.t130 464.166
R15348 a_n6972_8799.n220 a_n6972_8799.t50 464.166
R15349 a_n6972_8799.n206 a_n6972_8799.t90 464.166
R15350 a_n6972_8799.n219 a_n6972_8799.t38 464.166
R15351 a_n6972_8799.n218 a_n6972_8799.t110 464.166
R15352 a_n6972_8799.n207 a_n6972_8799.t60 464.166
R15353 a_n6972_8799.n217 a_n6972_8799.t96 464.166
R15354 a_n6972_8799.n216 a_n6972_8799.t43 464.166
R15355 a_n6972_8799.n208 a_n6972_8799.t64 464.166
R15356 a_n6972_8799.n215 a_n6972_8799.t126 464.166
R15357 a_n6972_8799.n214 a_n6972_8799.t102 464.166
R15358 a_n6972_8799.n209 a_n6972_8799.t121 464.166
R15359 a_n6972_8799.n213 a_n6972_8799.t88 464.166
R15360 a_n6972_8799.n212 a_n6972_8799.t105 464.166
R15361 a_n6972_8799.n210 a_n6972_8799.t54 464.166
R15362 a_n6972_8799.n126 a_n6972_8799.t76 464.166
R15363 a_n6972_8799.n129 a_n6972_8799.t77 464.166
R15364 a_n6972_8799.n125 a_n6972_8799.t100 464.166
R15365 a_n6972_8799.n130 a_n6972_8799.t67 464.166
R15366 a_n6972_8799.n131 a_n6972_8799.t68 464.166
R15367 a_n6972_8799.n132 a_n6972_8799.t99 464.166
R15368 a_n6972_8799.n133 a_n6972_8799.t36 464.166
R15369 a_n6972_8799.n124 a_n6972_8799.t65 464.166
R15370 a_n6972_8799.n134 a_n6972_8799.t82 464.166
R15371 a_n6972_8799.n135 a_n6972_8799.t116 464.166
R15372 a_n6972_8799.n136 a_n6972_8799.t47 464.166
R15373 a_n6972_8799.n137 a_n6972_8799.t63 464.166
R15374 a_n6972_8799.n123 a_n6972_8799.t113 464.166
R15375 a_n6972_8799.n138 a_n6972_8799.t44 464.166
R15376 a_n6972_8799.n142 a_n6972_8799.t83 464.166
R15377 a_n6972_8799.n145 a_n6972_8799.t84 464.166
R15378 a_n6972_8799.n141 a_n6972_8799.t112 464.166
R15379 a_n6972_8799.n146 a_n6972_8799.t74 464.166
R15380 a_n6972_8799.n147 a_n6972_8799.t75 464.166
R15381 a_n6972_8799.n148 a_n6972_8799.t108 464.166
R15382 a_n6972_8799.n149 a_n6972_8799.t46 464.166
R15383 a_n6972_8799.n140 a_n6972_8799.t73 464.166
R15384 a_n6972_8799.n150 a_n6972_8799.t93 464.166
R15385 a_n6972_8799.n151 a_n6972_8799.t128 464.166
R15386 a_n6972_8799.n152 a_n6972_8799.t61 464.166
R15387 a_n6972_8799.n153 a_n6972_8799.t72 464.166
R15388 a_n6972_8799.n139 a_n6972_8799.t123 464.166
R15389 a_n6972_8799.n154 a_n6972_8799.t55 464.166
R15390 a_n6972_8799.n159 a_n6972_8799.t53 464.166
R15391 a_n6972_8799.n162 a_n6972_8799.t37 464.166
R15392 a_n6972_8799.n158 a_n6972_8799.t87 464.166
R15393 a_n6972_8799.n163 a_n6972_8799.t120 464.166
R15394 a_n6972_8799.n164 a_n6972_8799.t101 464.166
R15395 a_n6972_8799.n165 a_n6972_8799.t124 464.166
R15396 a_n6972_8799.n166 a_n6972_8799.t81 464.166
R15397 a_n6972_8799.n157 a_n6972_8799.t42 464.166
R15398 a_n6972_8799.n167 a_n6972_8799.t95 464.166
R15399 a_n6972_8799.n168 a_n6972_8799.t59 464.166
R15400 a_n6972_8799.n169 a_n6972_8799.t109 464.166
R15401 a_n6972_8799.n170 a_n6972_8799.t66 464.166
R15402 a_n6972_8799.n156 a_n6972_8799.t89 464.166
R15403 a_n6972_8799.n171 a_n6972_8799.t49 464.166
R15404 a_n6972_8799.n52 a_n6972_8799.n34 74.4178
R15405 a_n6972_8799.n179 a_n6972_8799.n52 12.4674
R15406 a_n6972_8799.n51 a_n6972_8799.n34 80.107
R15407 a_n6972_8799.n51 a_n6972_8799.n180 1.08907
R15408 a_n6972_8799.n35 a_n6972_8799.n50 75.3623
R15409 a_n6972_8799.n49 a_n6972_8799.n35 70.3058
R15410 a_n6972_8799.n37 a_n6972_8799.n48 70.1674
R15411 a_n6972_8799.n48 a_n6972_8799.n175 20.9683
R15412 a_n6972_8799.n47 a_n6972_8799.n37 75.0448
R15413 a_n6972_8799.n183 a_n6972_8799.n47 11.2134
R15414 a_n6972_8799.n46 a_n6972_8799.n36 80.4688
R15415 a_n6972_8799.n36 a_n6972_8799.n45 74.73
R15416 a_n6972_8799.n44 a_n6972_8799.n38 70.1674
R15417 a_n6972_8799.n186 a_n6972_8799.n44 20.9683
R15418 a_n6972_8799.n38 a_n6972_8799.n43 70.5844
R15419 a_n6972_8799.n43 a_n6972_8799.n173 20.1342
R15420 a_n6972_8799.n42 a_n6972_8799.n39 75.6825
R15421 a_n6972_8799.n187 a_n6972_8799.n42 9.93802
R15422 a_n6972_8799.n39 a_n6972_8799.n188 161.3
R15423 a_n6972_8799.n63 a_n6972_8799.n28 74.4178
R15424 a_n6972_8799.n195 a_n6972_8799.n63 12.4674
R15425 a_n6972_8799.n62 a_n6972_8799.n28 80.107
R15426 a_n6972_8799.n62 a_n6972_8799.n196 1.08907
R15427 a_n6972_8799.n29 a_n6972_8799.n61 75.3623
R15428 a_n6972_8799.n60 a_n6972_8799.n29 70.3058
R15429 a_n6972_8799.n31 a_n6972_8799.n59 70.1674
R15430 a_n6972_8799.n59 a_n6972_8799.n191 20.9683
R15431 a_n6972_8799.n58 a_n6972_8799.n31 75.0448
R15432 a_n6972_8799.n199 a_n6972_8799.n58 11.2134
R15433 a_n6972_8799.n57 a_n6972_8799.n30 80.4688
R15434 a_n6972_8799.n30 a_n6972_8799.n56 74.73
R15435 a_n6972_8799.n55 a_n6972_8799.n32 70.1674
R15436 a_n6972_8799.n202 a_n6972_8799.n55 20.9683
R15437 a_n6972_8799.n32 a_n6972_8799.n54 70.5844
R15438 a_n6972_8799.n54 a_n6972_8799.n189 20.1342
R15439 a_n6972_8799.n53 a_n6972_8799.n33 75.6825
R15440 a_n6972_8799.n203 a_n6972_8799.n53 9.93802
R15441 a_n6972_8799.n33 a_n6972_8799.n204 161.3
R15442 a_n6972_8799.n74 a_n6972_8799.n22 74.4178
R15443 a_n6972_8799.n212 a_n6972_8799.n74 12.4674
R15444 a_n6972_8799.n73 a_n6972_8799.n22 80.107
R15445 a_n6972_8799.n73 a_n6972_8799.n213 1.08907
R15446 a_n6972_8799.n23 a_n6972_8799.n72 75.3623
R15447 a_n6972_8799.n71 a_n6972_8799.n23 70.3058
R15448 a_n6972_8799.n25 a_n6972_8799.n70 70.1674
R15449 a_n6972_8799.n70 a_n6972_8799.n208 20.9683
R15450 a_n6972_8799.n69 a_n6972_8799.n25 75.0448
R15451 a_n6972_8799.n216 a_n6972_8799.n69 11.2134
R15452 a_n6972_8799.n68 a_n6972_8799.n24 80.4688
R15453 a_n6972_8799.n24 a_n6972_8799.n67 74.73
R15454 a_n6972_8799.n66 a_n6972_8799.n26 70.1674
R15455 a_n6972_8799.n219 a_n6972_8799.n66 20.9683
R15456 a_n6972_8799.n26 a_n6972_8799.n65 70.5844
R15457 a_n6972_8799.n65 a_n6972_8799.n206 20.1342
R15458 a_n6972_8799.n64 a_n6972_8799.n27 75.6825
R15459 a_n6972_8799.n220 a_n6972_8799.n64 9.93802
R15460 a_n6972_8799.n27 a_n6972_8799.n221 161.3
R15461 a_n6972_8799.n17 a_n6972_8799.n85 70.1674
R15462 a_n6972_8799.n138 a_n6972_8799.n85 20.9683
R15463 a_n6972_8799.n84 a_n6972_8799.n17 74.4178
R15464 a_n6972_8799.n84 a_n6972_8799.n123 12.4674
R15465 a_n6972_8799.n16 a_n6972_8799.n83 80.107
R15466 a_n6972_8799.n137 a_n6972_8799.n83 1.08907
R15467 a_n6972_8799.n82 a_n6972_8799.n16 75.3623
R15468 a_n6972_8799.n18 a_n6972_8799.n81 70.3058
R15469 a_n6972_8799.n80 a_n6972_8799.n18 70.1674
R15470 a_n6972_8799.n80 a_n6972_8799.n124 20.9683
R15471 a_n6972_8799.n19 a_n6972_8799.n79 75.0448
R15472 a_n6972_8799.n133 a_n6972_8799.n79 11.2134
R15473 a_n6972_8799.n78 a_n6972_8799.n19 80.4688
R15474 a_n6972_8799.n20 a_n6972_8799.n77 74.73
R15475 a_n6972_8799.n76 a_n6972_8799.n20 70.1674
R15476 a_n6972_8799.n76 a_n6972_8799.n125 20.9683
R15477 a_n6972_8799.n21 a_n6972_8799.n75 70.5844
R15478 a_n6972_8799.n129 a_n6972_8799.n75 20.1342
R15479 a_n6972_8799.n128 a_n6972_8799.n21 161.3
R15480 a_n6972_8799.n11 a_n6972_8799.n96 70.1674
R15481 a_n6972_8799.n154 a_n6972_8799.n96 20.9683
R15482 a_n6972_8799.n95 a_n6972_8799.n11 74.4178
R15483 a_n6972_8799.n95 a_n6972_8799.n139 12.4674
R15484 a_n6972_8799.n10 a_n6972_8799.n94 80.107
R15485 a_n6972_8799.n153 a_n6972_8799.n94 1.08907
R15486 a_n6972_8799.n93 a_n6972_8799.n10 75.3623
R15487 a_n6972_8799.n12 a_n6972_8799.n92 70.3058
R15488 a_n6972_8799.n91 a_n6972_8799.n12 70.1674
R15489 a_n6972_8799.n91 a_n6972_8799.n140 20.9683
R15490 a_n6972_8799.n13 a_n6972_8799.n90 75.0448
R15491 a_n6972_8799.n149 a_n6972_8799.n90 11.2134
R15492 a_n6972_8799.n89 a_n6972_8799.n13 80.4688
R15493 a_n6972_8799.n14 a_n6972_8799.n88 74.73
R15494 a_n6972_8799.n87 a_n6972_8799.n14 70.1674
R15495 a_n6972_8799.n87 a_n6972_8799.n141 20.9683
R15496 a_n6972_8799.n15 a_n6972_8799.n86 70.5844
R15497 a_n6972_8799.n145 a_n6972_8799.n86 20.1342
R15498 a_n6972_8799.n144 a_n6972_8799.n15 161.3
R15499 a_n6972_8799.n5 a_n6972_8799.n107 70.1674
R15500 a_n6972_8799.n171 a_n6972_8799.n107 20.9683
R15501 a_n6972_8799.n106 a_n6972_8799.n5 74.4178
R15502 a_n6972_8799.n106 a_n6972_8799.n156 12.4674
R15503 a_n6972_8799.n4 a_n6972_8799.n105 80.107
R15504 a_n6972_8799.n170 a_n6972_8799.n105 1.08907
R15505 a_n6972_8799.n104 a_n6972_8799.n4 75.3623
R15506 a_n6972_8799.n6 a_n6972_8799.n103 70.3058
R15507 a_n6972_8799.n102 a_n6972_8799.n6 70.1674
R15508 a_n6972_8799.n102 a_n6972_8799.n157 20.9683
R15509 a_n6972_8799.n7 a_n6972_8799.n101 75.0448
R15510 a_n6972_8799.n166 a_n6972_8799.n101 11.2134
R15511 a_n6972_8799.n100 a_n6972_8799.n7 80.4688
R15512 a_n6972_8799.n8 a_n6972_8799.n99 74.73
R15513 a_n6972_8799.n98 a_n6972_8799.n8 70.1674
R15514 a_n6972_8799.n98 a_n6972_8799.n158 20.9683
R15515 a_n6972_8799.n9 a_n6972_8799.n97 70.5844
R15516 a_n6972_8799.n162 a_n6972_8799.n97 20.1342
R15517 a_n6972_8799.n161 a_n6972_8799.n9 161.3
R15518 a_n6972_8799.n40 a_n6972_8799.n108 98.9633
R15519 a_n6972_8799.n228 a_n6972_8799.n41 98.9632
R15520 a_n6972_8799.n41 a_n6972_8799.n227 98.6055
R15521 a_n6972_8799.n41 a_n6972_8799.n226 98.6055
R15522 a_n6972_8799.n40 a_n6972_8799.n110 98.6055
R15523 a_n6972_8799.n40 a_n6972_8799.n109 98.6055
R15524 a_n6972_8799.n1 a_n6972_8799.n111 81.4626
R15525 a_n6972_8799.n3 a_n6972_8799.n117 81.4626
R15526 a_n6972_8799.n0 a_n6972_8799.n114 81.4626
R15527 a_n6972_8799.n2 a_n6972_8799.n120 80.9324
R15528 a_n6972_8799.n2 a_n6972_8799.n121 80.9324
R15529 a_n6972_8799.n1 a_n6972_8799.n122 80.9324
R15530 a_n6972_8799.n1 a_n6972_8799.n113 80.9324
R15531 a_n6972_8799.n1 a_n6972_8799.n112 80.9324
R15532 a_n6972_8799.n3 a_n6972_8799.n118 80.9324
R15533 a_n6972_8799.n0 a_n6972_8799.n119 80.9324
R15534 a_n6972_8799.n0 a_n6972_8799.n116 80.9324
R15535 a_n6972_8799.n0 a_n6972_8799.n115 80.9324
R15536 a_n6972_8799.n34 a_n6972_8799.n178 70.4033
R15537 a_n6972_8799.n28 a_n6972_8799.n194 70.4033
R15538 a_n6972_8799.n22 a_n6972_8799.n211 70.4033
R15539 a_n6972_8799.n21 a_n6972_8799.n127 70.4033
R15540 a_n6972_8799.n15 a_n6972_8799.n143 70.4033
R15541 a_n6972_8799.n9 a_n6972_8799.n160 70.4033
R15542 a_n6972_8799.n188 a_n6972_8799.n187 48.2005
R15543 a_n6972_8799.n44 a_n6972_8799.n185 20.9683
R15544 a_n6972_8799.n184 a_n6972_8799.n183 48.2005
R15545 a_n6972_8799.n182 a_n6972_8799.n48 20.9683
R15546 a_n6972_8799.n180 a_n6972_8799.n176 48.2005
R15547 a_n6972_8799.n204 a_n6972_8799.n203 48.2005
R15548 a_n6972_8799.n55 a_n6972_8799.n201 20.9683
R15549 a_n6972_8799.n200 a_n6972_8799.n199 48.2005
R15550 a_n6972_8799.n198 a_n6972_8799.n59 20.9683
R15551 a_n6972_8799.n196 a_n6972_8799.n192 48.2005
R15552 a_n6972_8799.n221 a_n6972_8799.n220 48.2005
R15553 a_n6972_8799.n66 a_n6972_8799.n218 20.9683
R15554 a_n6972_8799.n217 a_n6972_8799.n216 48.2005
R15555 a_n6972_8799.n215 a_n6972_8799.n70 20.9683
R15556 a_n6972_8799.n213 a_n6972_8799.n209 48.2005
R15557 a_n6972_8799.n130 a_n6972_8799.n76 20.9683
R15558 a_n6972_8799.n133 a_n6972_8799.n132 48.2005
R15559 a_n6972_8799.n134 a_n6972_8799.n80 20.9683
R15560 a_n6972_8799.n137 a_n6972_8799.n136 48.2005
R15561 a_n6972_8799.t45 a_n6972_8799.n85 485.135
R15562 a_n6972_8799.n146 a_n6972_8799.n87 20.9683
R15563 a_n6972_8799.n149 a_n6972_8799.n148 48.2005
R15564 a_n6972_8799.n150 a_n6972_8799.n91 20.9683
R15565 a_n6972_8799.n153 a_n6972_8799.n152 48.2005
R15566 a_n6972_8799.t57 a_n6972_8799.n96 485.135
R15567 a_n6972_8799.n163 a_n6972_8799.n98 20.9683
R15568 a_n6972_8799.n166 a_n6972_8799.n165 48.2005
R15569 a_n6972_8799.n167 a_n6972_8799.n102 20.9683
R15570 a_n6972_8799.n170 a_n6972_8799.n169 48.2005
R15571 a_n6972_8799.t129 a_n6972_8799.n107 485.135
R15572 a_n6972_8799.n46 a_n6972_8799.n174 47.835
R15573 a_n6972_8799.n49 a_n6972_8799.n181 20.6913
R15574 a_n6972_8799.n57 a_n6972_8799.n190 47.835
R15575 a_n6972_8799.n60 a_n6972_8799.n197 20.6913
R15576 a_n6972_8799.n68 a_n6972_8799.n207 47.835
R15577 a_n6972_8799.n71 a_n6972_8799.n214 20.6913
R15578 a_n6972_8799.n131 a_n6972_8799.n78 47.835
R15579 a_n6972_8799.n135 a_n6972_8799.n81 20.6913
R15580 a_n6972_8799.n147 a_n6972_8799.n89 47.835
R15581 a_n6972_8799.n151 a_n6972_8799.n92 20.6913
R15582 a_n6972_8799.n164 a_n6972_8799.n100 47.835
R15583 a_n6972_8799.n168 a_n6972_8799.n103 20.6913
R15584 a_n6972_8799.n186 a_n6972_8799.n43 22.3251
R15585 a_n6972_8799.n202 a_n6972_8799.n54 22.3251
R15586 a_n6972_8799.n219 a_n6972_8799.n65 22.3251
R15587 a_n6972_8799.n125 a_n6972_8799.n75 22.3251
R15588 a_n6972_8799.n141 a_n6972_8799.n86 22.3251
R15589 a_n6972_8799.n158 a_n6972_8799.n97 22.3251
R15590 a_n6972_8799.n2 a_n6972_8799.n0 34.3237
R15591 a_n6972_8799.n52 a_n6972_8799.n177 33.6462
R15592 a_n6972_8799.n63 a_n6972_8799.n193 33.6462
R15593 a_n6972_8799.n74 a_n6972_8799.n210 33.6462
R15594 a_n6972_8799.n129 a_n6972_8799.n128 27.0217
R15595 a_n6972_8799.n138 a_n6972_8799.n84 33.6462
R15596 a_n6972_8799.n145 a_n6972_8799.n144 27.0217
R15597 a_n6972_8799.n154 a_n6972_8799.n95 33.6462
R15598 a_n6972_8799.n162 a_n6972_8799.n161 27.0217
R15599 a_n6972_8799.n171 a_n6972_8799.n106 33.6462
R15600 a_n6972_8799.n45 a_n6972_8799.n174 11.843
R15601 a_n6972_8799.n181 a_n6972_8799.n50 36.139
R15602 a_n6972_8799.n56 a_n6972_8799.n190 11.843
R15603 a_n6972_8799.n197 a_n6972_8799.n61 36.139
R15604 a_n6972_8799.n67 a_n6972_8799.n207 11.843
R15605 a_n6972_8799.n214 a_n6972_8799.n72 36.139
R15606 a_n6972_8799.n131 a_n6972_8799.n77 11.843
R15607 a_n6972_8799.n135 a_n6972_8799.n82 36.139
R15608 a_n6972_8799.n147 a_n6972_8799.n88 11.843
R15609 a_n6972_8799.n151 a_n6972_8799.n93 36.139
R15610 a_n6972_8799.n164 a_n6972_8799.n99 11.843
R15611 a_n6972_8799.n168 a_n6972_8799.n104 36.139
R15612 a_n6972_8799.n47 a_n6972_8799.n175 35.3134
R15613 a_n6972_8799.n58 a_n6972_8799.n191 35.3134
R15614 a_n6972_8799.n69 a_n6972_8799.n208 35.3134
R15615 a_n6972_8799.n124 a_n6972_8799.n79 35.3134
R15616 a_n6972_8799.n140 a_n6972_8799.n90 35.3134
R15617 a_n6972_8799.n157 a_n6972_8799.n101 35.3134
R15618 a_n6972_8799.n185 a_n6972_8799.n45 34.4824
R15619 a_n6972_8799.n50 a_n6972_8799.n176 10.5784
R15620 a_n6972_8799.n201 a_n6972_8799.n56 34.4824
R15621 a_n6972_8799.n61 a_n6972_8799.n192 10.5784
R15622 a_n6972_8799.n218 a_n6972_8799.n67 34.4824
R15623 a_n6972_8799.n72 a_n6972_8799.n209 10.5784
R15624 a_n6972_8799.n77 a_n6972_8799.n130 34.4824
R15625 a_n6972_8799.n136 a_n6972_8799.n82 10.5784
R15626 a_n6972_8799.n88 a_n6972_8799.n146 34.4824
R15627 a_n6972_8799.n152 a_n6972_8799.n93 10.5784
R15628 a_n6972_8799.n99 a_n6972_8799.n163 34.4824
R15629 a_n6972_8799.n169 a_n6972_8799.n104 10.5784
R15630 a_n6972_8799.n42 a_n6972_8799.n173 36.9592
R15631 a_n6972_8799.n53 a_n6972_8799.n189 36.9592
R15632 a_n6972_8799.n64 a_n6972_8799.n206 36.9592
R15633 a_n6972_8799.n128 a_n6972_8799.n126 21.1793
R15634 a_n6972_8799.n144 a_n6972_8799.n142 21.1793
R15635 a_n6972_8799.n161 a_n6972_8799.n159 21.1793
R15636 a_n6972_8799.n178 a_n6972_8799.n177 20.9576
R15637 a_n6972_8799.n194 a_n6972_8799.n193 20.9576
R15638 a_n6972_8799.n211 a_n6972_8799.n210 20.9576
R15639 a_n6972_8799.n127 a_n6972_8799.n126 20.9576
R15640 a_n6972_8799.n143 a_n6972_8799.n142 20.9576
R15641 a_n6972_8799.n160 a_n6972_8799.n159 20.9576
R15642 a_n6972_8799.n224 a_n6972_8799.n1 12.3339
R15643 a_n6972_8799.n225 a_n6972_8799.n224 11.4887
R15644 a_n6972_8799.n205 a_n6972_8799.n39 9.07815
R15645 a_n6972_8799.n155 a_n6972_8799.n17 9.07815
R15646 a_n6972_8799.n223 a_n6972_8799.n172 6.93972
R15647 a_n6972_8799.n223 a_n6972_8799.n222 6.44309
R15648 a_n6972_8799.n205 a_n6972_8799.n33 4.9702
R15649 a_n6972_8799.n222 a_n6972_8799.n27 4.9702
R15650 a_n6972_8799.n155 a_n6972_8799.n11 4.9702
R15651 a_n6972_8799.n172 a_n6972_8799.n5 4.9702
R15652 a_n6972_8799.n222 a_n6972_8799.n205 4.10845
R15653 a_n6972_8799.n172 a_n6972_8799.n155 4.10845
R15654 a_n6972_8799.n227 a_n6972_8799.t35 3.61217
R15655 a_n6972_8799.n227 a_n6972_8799.t5 3.61217
R15656 a_n6972_8799.n226 a_n6972_8799.t34 3.61217
R15657 a_n6972_8799.n226 a_n6972_8799.t4 3.61217
R15658 a_n6972_8799.n110 a_n6972_8799.t21 3.61217
R15659 a_n6972_8799.n110 a_n6972_8799.t29 3.61217
R15660 a_n6972_8799.n109 a_n6972_8799.t17 3.61217
R15661 a_n6972_8799.n109 a_n6972_8799.t12 3.61217
R15662 a_n6972_8799.n108 a_n6972_8799.t33 3.61217
R15663 a_n6972_8799.n108 a_n6972_8799.t6 3.61217
R15664 a_n6972_8799.t3 a_n6972_8799.n228 3.61217
R15665 a_n6972_8799.n228 a_n6972_8799.t11 3.61217
R15666 a_n6972_8799.n224 a_n6972_8799.n223 3.4105
R15667 a_n6972_8799.n120 a_n6972_8799.t10 2.82907
R15668 a_n6972_8799.n120 a_n6972_8799.t13 2.82907
R15669 a_n6972_8799.n121 a_n6972_8799.t15 2.82907
R15670 a_n6972_8799.n121 a_n6972_8799.t28 2.82907
R15671 a_n6972_8799.n122 a_n6972_8799.t30 2.82907
R15672 a_n6972_8799.n122 a_n6972_8799.t31 2.82907
R15673 a_n6972_8799.n113 a_n6972_8799.t18 2.82907
R15674 a_n6972_8799.n113 a_n6972_8799.t23 2.82907
R15675 a_n6972_8799.n112 a_n6972_8799.t19 2.82907
R15676 a_n6972_8799.n112 a_n6972_8799.t2 2.82907
R15677 a_n6972_8799.n111 a_n6972_8799.t20 2.82907
R15678 a_n6972_8799.n111 a_n6972_8799.t22 2.82907
R15679 a_n6972_8799.n117 a_n6972_8799.t7 2.82907
R15680 a_n6972_8799.n117 a_n6972_8799.t8 2.82907
R15681 a_n6972_8799.n118 a_n6972_8799.t9 2.82907
R15682 a_n6972_8799.n118 a_n6972_8799.t16 2.82907
R15683 a_n6972_8799.n119 a_n6972_8799.t25 2.82907
R15684 a_n6972_8799.n119 a_n6972_8799.t24 2.82907
R15685 a_n6972_8799.n116 a_n6972_8799.t14 2.82907
R15686 a_n6972_8799.n116 a_n6972_8799.t26 2.82907
R15687 a_n6972_8799.n115 a_n6972_8799.t0 2.82907
R15688 a_n6972_8799.n115 a_n6972_8799.t1 2.82907
R15689 a_n6972_8799.n114 a_n6972_8799.t27 2.82907
R15690 a_n6972_8799.n114 a_n6972_8799.t32 2.82907
R15691 a_n6972_8799.n51 a_n6972_8799.n179 47.0982
R15692 a_n6972_8799.n62 a_n6972_8799.n195 47.0982
R15693 a_n6972_8799.n73 a_n6972_8799.n212 47.0982
R15694 a_n6972_8799.n123 a_n6972_8799.n83 47.0982
R15695 a_n6972_8799.n139 a_n6972_8799.n94 47.0982
R15696 a_n6972_8799.n156 a_n6972_8799.n105 47.0982
R15697 a_n6972_8799.n41 a_n6972_8799.n225 31.5519
R15698 a_n6972_8799.n46 a_n6972_8799.n184 0.365327
R15699 a_n6972_8799.n182 a_n6972_8799.n49 21.4216
R15700 a_n6972_8799.n57 a_n6972_8799.n200 0.365327
R15701 a_n6972_8799.n198 a_n6972_8799.n60 21.4216
R15702 a_n6972_8799.n68 a_n6972_8799.n217 0.365327
R15703 a_n6972_8799.n215 a_n6972_8799.n71 21.4216
R15704 a_n6972_8799.n132 a_n6972_8799.n78 0.365327
R15705 a_n6972_8799.n81 a_n6972_8799.n134 21.4216
R15706 a_n6972_8799.n148 a_n6972_8799.n89 0.365327
R15707 a_n6972_8799.n92 a_n6972_8799.n150 21.4216
R15708 a_n6972_8799.n165 a_n6972_8799.n100 0.365327
R15709 a_n6972_8799.n103 a_n6972_8799.n167 21.4216
R15710 a_n6972_8799.n225 a_n6972_8799.n40 17.6132
R15711 a_n6972_8799.n1 a_n6972_8799.n2 2.12119
R15712 a_n6972_8799.n0 a_n6972_8799.n3 1.59102
R15713 a_n6972_8799.n35 a_n6972_8799.n34 1.13686
R15714 a_n6972_8799.n29 a_n6972_8799.n28 1.13686
R15715 a_n6972_8799.n23 a_n6972_8799.n22 1.13686
R15716 a_n6972_8799.n17 a_n6972_8799.n16 1.13686
R15717 a_n6972_8799.n11 a_n6972_8799.n10 1.13686
R15718 a_n6972_8799.n5 a_n6972_8799.n4 1.13686
R15719 a_n6972_8799.n39 a_n6972_8799.n38 0.758076
R15720 a_n6972_8799.n36 a_n6972_8799.n38 0.758076
R15721 a_n6972_8799.n37 a_n6972_8799.n36 0.758076
R15722 a_n6972_8799.n37 a_n6972_8799.n35 0.758076
R15723 a_n6972_8799.n33 a_n6972_8799.n32 0.758076
R15724 a_n6972_8799.n30 a_n6972_8799.n32 0.758076
R15725 a_n6972_8799.n31 a_n6972_8799.n30 0.758076
R15726 a_n6972_8799.n31 a_n6972_8799.n29 0.758076
R15727 a_n6972_8799.n27 a_n6972_8799.n26 0.758076
R15728 a_n6972_8799.n24 a_n6972_8799.n26 0.758076
R15729 a_n6972_8799.n25 a_n6972_8799.n24 0.758076
R15730 a_n6972_8799.n25 a_n6972_8799.n23 0.758076
R15731 a_n6972_8799.n20 a_n6972_8799.n21 0.758076
R15732 a_n6972_8799.n19 a_n6972_8799.n20 0.758076
R15733 a_n6972_8799.n18 a_n6972_8799.n19 0.758076
R15734 a_n6972_8799.n16 a_n6972_8799.n18 0.758076
R15735 a_n6972_8799.n14 a_n6972_8799.n15 0.758076
R15736 a_n6972_8799.n13 a_n6972_8799.n14 0.758076
R15737 a_n6972_8799.n12 a_n6972_8799.n13 0.758076
R15738 a_n6972_8799.n10 a_n6972_8799.n12 0.758076
R15739 a_n6972_8799.n8 a_n6972_8799.n9 0.758076
R15740 a_n6972_8799.n7 a_n6972_8799.n8 0.758076
R15741 a_n6972_8799.n6 a_n6972_8799.n7 0.758076
R15742 a_n6972_8799.n4 a_n6972_8799.n6 0.758076
R15743 vdd.n315 vdd.n279 756.745
R15744 vdd.n260 vdd.n224 756.745
R15745 vdd.n217 vdd.n181 756.745
R15746 vdd.n162 vdd.n126 756.745
R15747 vdd.n120 vdd.n84 756.745
R15748 vdd.n65 vdd.n29 756.745
R15749 vdd.n1684 vdd.n1648 756.745
R15750 vdd.n1739 vdd.n1703 756.745
R15751 vdd.n1586 vdd.n1550 756.745
R15752 vdd.n1641 vdd.n1605 756.745
R15753 vdd.n1489 vdd.n1453 756.745
R15754 vdd.n1544 vdd.n1508 756.745
R15755 vdd.n2094 vdd.t226 640.208
R15756 vdd.n936 vdd.t211 640.208
R15757 vdd.n2068 vdd.t172 640.208
R15758 vdd.n928 vdd.t236 640.208
R15759 vdd.n2839 vdd.t198 640.208
R15760 vdd.n2559 vdd.t233 640.208
R15761 vdd.n804 vdd.t215 640.208
R15762 vdd.n2556 vdd.t219 640.208
R15763 vdd.n768 vdd.t223 640.208
R15764 vdd.n998 vdd.t229 640.208
R15765 vdd.n1148 vdd.t184 592.009
R15766 vdd.n1304 vdd.t195 592.009
R15767 vdd.n1340 vdd.t202 592.009
R15768 vdd.n2250 vdd.t191 592.009
R15769 vdd.n1887 vdd.t205 592.009
R15770 vdd.n1847 vdd.t208 592.009
R15771 vdd.n405 vdd.t180 592.009
R15772 vdd.n419 vdd.t239 592.009
R15773 vdd.n431 vdd.t245 592.009
R15774 vdd.n723 vdd.t176 592.009
R15775 vdd.n686 vdd.t188 592.009
R15776 vdd.n3013 vdd.t242 592.009
R15777 vdd.n316 vdd.n315 585
R15778 vdd.n314 vdd.n281 585
R15779 vdd.n313 vdd.n312 585
R15780 vdd.n284 vdd.n282 585
R15781 vdd.n307 vdd.n306 585
R15782 vdd.n305 vdd.n304 585
R15783 vdd.n288 vdd.n287 585
R15784 vdd.n299 vdd.n298 585
R15785 vdd.n297 vdd.n296 585
R15786 vdd.n292 vdd.n291 585
R15787 vdd.n261 vdd.n260 585
R15788 vdd.n259 vdd.n226 585
R15789 vdd.n258 vdd.n257 585
R15790 vdd.n229 vdd.n227 585
R15791 vdd.n252 vdd.n251 585
R15792 vdd.n250 vdd.n249 585
R15793 vdd.n233 vdd.n232 585
R15794 vdd.n244 vdd.n243 585
R15795 vdd.n242 vdd.n241 585
R15796 vdd.n237 vdd.n236 585
R15797 vdd.n218 vdd.n217 585
R15798 vdd.n216 vdd.n183 585
R15799 vdd.n215 vdd.n214 585
R15800 vdd.n186 vdd.n184 585
R15801 vdd.n209 vdd.n208 585
R15802 vdd.n207 vdd.n206 585
R15803 vdd.n190 vdd.n189 585
R15804 vdd.n201 vdd.n200 585
R15805 vdd.n199 vdd.n198 585
R15806 vdd.n194 vdd.n193 585
R15807 vdd.n163 vdd.n162 585
R15808 vdd.n161 vdd.n128 585
R15809 vdd.n160 vdd.n159 585
R15810 vdd.n131 vdd.n129 585
R15811 vdd.n154 vdd.n153 585
R15812 vdd.n152 vdd.n151 585
R15813 vdd.n135 vdd.n134 585
R15814 vdd.n146 vdd.n145 585
R15815 vdd.n144 vdd.n143 585
R15816 vdd.n139 vdd.n138 585
R15817 vdd.n121 vdd.n120 585
R15818 vdd.n119 vdd.n86 585
R15819 vdd.n118 vdd.n117 585
R15820 vdd.n89 vdd.n87 585
R15821 vdd.n112 vdd.n111 585
R15822 vdd.n110 vdd.n109 585
R15823 vdd.n93 vdd.n92 585
R15824 vdd.n104 vdd.n103 585
R15825 vdd.n102 vdd.n101 585
R15826 vdd.n97 vdd.n96 585
R15827 vdd.n66 vdd.n65 585
R15828 vdd.n64 vdd.n31 585
R15829 vdd.n63 vdd.n62 585
R15830 vdd.n34 vdd.n32 585
R15831 vdd.n57 vdd.n56 585
R15832 vdd.n55 vdd.n54 585
R15833 vdd.n38 vdd.n37 585
R15834 vdd.n49 vdd.n48 585
R15835 vdd.n47 vdd.n46 585
R15836 vdd.n42 vdd.n41 585
R15837 vdd.n1685 vdd.n1684 585
R15838 vdd.n1683 vdd.n1650 585
R15839 vdd.n1682 vdd.n1681 585
R15840 vdd.n1653 vdd.n1651 585
R15841 vdd.n1676 vdd.n1675 585
R15842 vdd.n1674 vdd.n1673 585
R15843 vdd.n1657 vdd.n1656 585
R15844 vdd.n1668 vdd.n1667 585
R15845 vdd.n1666 vdd.n1665 585
R15846 vdd.n1661 vdd.n1660 585
R15847 vdd.n1740 vdd.n1739 585
R15848 vdd.n1738 vdd.n1705 585
R15849 vdd.n1737 vdd.n1736 585
R15850 vdd.n1708 vdd.n1706 585
R15851 vdd.n1731 vdd.n1730 585
R15852 vdd.n1729 vdd.n1728 585
R15853 vdd.n1712 vdd.n1711 585
R15854 vdd.n1723 vdd.n1722 585
R15855 vdd.n1721 vdd.n1720 585
R15856 vdd.n1716 vdd.n1715 585
R15857 vdd.n1587 vdd.n1586 585
R15858 vdd.n1585 vdd.n1552 585
R15859 vdd.n1584 vdd.n1583 585
R15860 vdd.n1555 vdd.n1553 585
R15861 vdd.n1578 vdd.n1577 585
R15862 vdd.n1576 vdd.n1575 585
R15863 vdd.n1559 vdd.n1558 585
R15864 vdd.n1570 vdd.n1569 585
R15865 vdd.n1568 vdd.n1567 585
R15866 vdd.n1563 vdd.n1562 585
R15867 vdd.n1642 vdd.n1641 585
R15868 vdd.n1640 vdd.n1607 585
R15869 vdd.n1639 vdd.n1638 585
R15870 vdd.n1610 vdd.n1608 585
R15871 vdd.n1633 vdd.n1632 585
R15872 vdd.n1631 vdd.n1630 585
R15873 vdd.n1614 vdd.n1613 585
R15874 vdd.n1625 vdd.n1624 585
R15875 vdd.n1623 vdd.n1622 585
R15876 vdd.n1618 vdd.n1617 585
R15877 vdd.n1490 vdd.n1489 585
R15878 vdd.n1488 vdd.n1455 585
R15879 vdd.n1487 vdd.n1486 585
R15880 vdd.n1458 vdd.n1456 585
R15881 vdd.n1481 vdd.n1480 585
R15882 vdd.n1479 vdd.n1478 585
R15883 vdd.n1462 vdd.n1461 585
R15884 vdd.n1473 vdd.n1472 585
R15885 vdd.n1471 vdd.n1470 585
R15886 vdd.n1466 vdd.n1465 585
R15887 vdd.n1545 vdd.n1544 585
R15888 vdd.n1543 vdd.n1510 585
R15889 vdd.n1542 vdd.n1541 585
R15890 vdd.n1513 vdd.n1511 585
R15891 vdd.n1536 vdd.n1535 585
R15892 vdd.n1534 vdd.n1533 585
R15893 vdd.n1517 vdd.n1516 585
R15894 vdd.n1528 vdd.n1527 585
R15895 vdd.n1526 vdd.n1525 585
R15896 vdd.n1521 vdd.n1520 585
R15897 vdd.n445 vdd.n370 462.44
R15898 vdd.n3251 vdd.n372 462.44
R15899 vdd.n3146 vdd.n657 462.44
R15900 vdd.n3144 vdd.n660 462.44
R15901 vdd.n2245 vdd.n1047 462.44
R15902 vdd.n2248 vdd.n2247 462.44
R15903 vdd.n1375 vdd.n1145 462.44
R15904 vdd.n1372 vdd.n1143 462.44
R15905 vdd.n293 vdd.t148 329.043
R15906 vdd.n238 vdd.t125 329.043
R15907 vdd.n195 vdd.t137 329.043
R15908 vdd.n140 vdd.t113 329.043
R15909 vdd.n98 vdd.t70 329.043
R15910 vdd.n43 vdd.t47 329.043
R15911 vdd.n1662 vdd.t163 329.043
R15912 vdd.n1717 vdd.t73 329.043
R15913 vdd.n1564 vdd.t149 329.043
R15914 vdd.n1619 vdd.t57 329.043
R15915 vdd.n1467 vdd.t51 329.043
R15916 vdd.n1522 vdd.t72 329.043
R15917 vdd.n1148 vdd.t187 319.788
R15918 vdd.n1304 vdd.t197 319.788
R15919 vdd.n1340 vdd.t204 319.788
R15920 vdd.n2250 vdd.t193 319.788
R15921 vdd.n1887 vdd.t206 319.788
R15922 vdd.n1847 vdd.t209 319.788
R15923 vdd.n405 vdd.t182 319.788
R15924 vdd.n419 vdd.t240 319.788
R15925 vdd.n431 vdd.t246 319.788
R15926 vdd.n723 vdd.t179 319.788
R15927 vdd.n686 vdd.t190 319.788
R15928 vdd.n3013 vdd.t244 319.788
R15929 vdd.n1149 vdd.t186 303.69
R15930 vdd.n1305 vdd.t196 303.69
R15931 vdd.n1341 vdd.t203 303.69
R15932 vdd.n2251 vdd.t194 303.69
R15933 vdd.n1888 vdd.t207 303.69
R15934 vdd.n1848 vdd.t210 303.69
R15935 vdd.n406 vdd.t183 303.69
R15936 vdd.n420 vdd.t241 303.69
R15937 vdd.n432 vdd.t247 303.69
R15938 vdd.n724 vdd.t178 303.69
R15939 vdd.n687 vdd.t189 303.69
R15940 vdd.n3014 vdd.t243 303.69
R15941 vdd.n2782 vdd.n884 297.074
R15942 vdd.n2975 vdd.n778 297.074
R15943 vdd.n2912 vdd.n775 297.074
R15944 vdd.n2705 vdd.n885 297.074
R15945 vdd.n2520 vdd.n925 297.074
R15946 vdd.n2451 vdd.n2450 297.074
R15947 vdd.n2197 vdd.n1021 297.074
R15948 vdd.n2293 vdd.n1019 297.074
R15949 vdd.n2891 vdd.n776 297.074
R15950 vdd.n2978 vdd.n2977 297.074
R15951 vdd.n2554 vdd.n886 297.074
R15952 vdd.n2780 vdd.n887 297.074
R15953 vdd.n2448 vdd.n934 297.074
R15954 vdd.n932 vdd.n907 297.074
R15955 vdd.n2134 vdd.n1022 297.074
R15956 vdd.n2291 vdd.n1023 297.074
R15957 vdd.n2893 vdd.n776 185
R15958 vdd.n2976 vdd.n776 185
R15959 vdd.n2895 vdd.n2894 185
R15960 vdd.n2894 vdd.n774 185
R15961 vdd.n2896 vdd.n810 185
R15962 vdd.n2906 vdd.n810 185
R15963 vdd.n2897 vdd.n819 185
R15964 vdd.n819 vdd.n817 185
R15965 vdd.n2899 vdd.n2898 185
R15966 vdd.n2900 vdd.n2899 185
R15967 vdd.n2852 vdd.n818 185
R15968 vdd.n818 vdd.n814 185
R15969 vdd.n2851 vdd.n2850 185
R15970 vdd.n2850 vdd.n2849 185
R15971 vdd.n821 vdd.n820 185
R15972 vdd.n822 vdd.n821 185
R15973 vdd.n2842 vdd.n2841 185
R15974 vdd.n2843 vdd.n2842 185
R15975 vdd.n2838 vdd.n831 185
R15976 vdd.n831 vdd.n828 185
R15977 vdd.n2837 vdd.n2836 185
R15978 vdd.n2836 vdd.n2835 185
R15979 vdd.n833 vdd.n832 185
R15980 vdd.n841 vdd.n833 185
R15981 vdd.n2828 vdd.n2827 185
R15982 vdd.n2829 vdd.n2828 185
R15983 vdd.n2826 vdd.n842 185
R15984 vdd.n2677 vdd.n842 185
R15985 vdd.n2825 vdd.n2824 185
R15986 vdd.n2824 vdd.n2823 185
R15987 vdd.n844 vdd.n843 185
R15988 vdd.n845 vdd.n844 185
R15989 vdd.n2816 vdd.n2815 185
R15990 vdd.n2817 vdd.n2816 185
R15991 vdd.n2814 vdd.n854 185
R15992 vdd.n854 vdd.n851 185
R15993 vdd.n2813 vdd.n2812 185
R15994 vdd.n2812 vdd.n2811 185
R15995 vdd.n856 vdd.n855 185
R15996 vdd.n864 vdd.n856 185
R15997 vdd.n2804 vdd.n2803 185
R15998 vdd.n2805 vdd.n2804 185
R15999 vdd.n2802 vdd.n865 185
R16000 vdd.n871 vdd.n865 185
R16001 vdd.n2801 vdd.n2800 185
R16002 vdd.n2800 vdd.n2799 185
R16003 vdd.n867 vdd.n866 185
R16004 vdd.n868 vdd.n867 185
R16005 vdd.n2792 vdd.n2791 185
R16006 vdd.n2793 vdd.n2792 185
R16007 vdd.n2790 vdd.n877 185
R16008 vdd.n2698 vdd.n877 185
R16009 vdd.n2789 vdd.n2788 185
R16010 vdd.n2788 vdd.n2787 185
R16011 vdd.n879 vdd.n878 185
R16012 vdd.t34 vdd.n879 185
R16013 vdd.n2780 vdd.n2779 185
R16014 vdd.n2781 vdd.n2780 185
R16015 vdd.n2778 vdd.n887 185
R16016 vdd.n2777 vdd.n2776 185
R16017 vdd.n889 vdd.n888 185
R16018 vdd.n2563 vdd.n2562 185
R16019 vdd.n2565 vdd.n2564 185
R16020 vdd.n2567 vdd.n2566 185
R16021 vdd.n2569 vdd.n2568 185
R16022 vdd.n2571 vdd.n2570 185
R16023 vdd.n2573 vdd.n2572 185
R16024 vdd.n2575 vdd.n2574 185
R16025 vdd.n2577 vdd.n2576 185
R16026 vdd.n2579 vdd.n2578 185
R16027 vdd.n2581 vdd.n2580 185
R16028 vdd.n2583 vdd.n2582 185
R16029 vdd.n2585 vdd.n2584 185
R16030 vdd.n2587 vdd.n2586 185
R16031 vdd.n2589 vdd.n2588 185
R16032 vdd.n2591 vdd.n2590 185
R16033 vdd.n2593 vdd.n2592 185
R16034 vdd.n2595 vdd.n2594 185
R16035 vdd.n2597 vdd.n2596 185
R16036 vdd.n2599 vdd.n2598 185
R16037 vdd.n2601 vdd.n2600 185
R16038 vdd.n2603 vdd.n2602 185
R16039 vdd.n2605 vdd.n2604 185
R16040 vdd.n2607 vdd.n2606 185
R16041 vdd.n2609 vdd.n2608 185
R16042 vdd.n2611 vdd.n2610 185
R16043 vdd.n2613 vdd.n2612 185
R16044 vdd.n2615 vdd.n2614 185
R16045 vdd.n2617 vdd.n2616 185
R16046 vdd.n2619 vdd.n2618 185
R16047 vdd.n2621 vdd.n2620 185
R16048 vdd.n2623 vdd.n2622 185
R16049 vdd.n2624 vdd.n2554 185
R16050 vdd.n2774 vdd.n2554 185
R16051 vdd.n2979 vdd.n2978 185
R16052 vdd.n2980 vdd.n767 185
R16053 vdd.n2982 vdd.n2981 185
R16054 vdd.n2984 vdd.n765 185
R16055 vdd.n2986 vdd.n2985 185
R16056 vdd.n2987 vdd.n764 185
R16057 vdd.n2989 vdd.n2988 185
R16058 vdd.n2991 vdd.n762 185
R16059 vdd.n2993 vdd.n2992 185
R16060 vdd.n2994 vdd.n761 185
R16061 vdd.n2996 vdd.n2995 185
R16062 vdd.n2998 vdd.n759 185
R16063 vdd.n3000 vdd.n2999 185
R16064 vdd.n3001 vdd.n758 185
R16065 vdd.n3003 vdd.n3002 185
R16066 vdd.n3005 vdd.n757 185
R16067 vdd.n3006 vdd.n754 185
R16068 vdd.n3009 vdd.n3008 185
R16069 vdd.n755 vdd.n753 185
R16070 vdd.n2865 vdd.n2864 185
R16071 vdd.n2867 vdd.n2866 185
R16072 vdd.n2869 vdd.n2861 185
R16073 vdd.n2871 vdd.n2870 185
R16074 vdd.n2872 vdd.n2860 185
R16075 vdd.n2874 vdd.n2873 185
R16076 vdd.n2876 vdd.n2858 185
R16077 vdd.n2878 vdd.n2877 185
R16078 vdd.n2879 vdd.n2857 185
R16079 vdd.n2881 vdd.n2880 185
R16080 vdd.n2883 vdd.n2855 185
R16081 vdd.n2885 vdd.n2884 185
R16082 vdd.n2886 vdd.n2854 185
R16083 vdd.n2888 vdd.n2887 185
R16084 vdd.n2890 vdd.n2853 185
R16085 vdd.n2892 vdd.n2891 185
R16086 vdd.n2891 vdd.n756 185
R16087 vdd.n2977 vdd.n771 185
R16088 vdd.n2977 vdd.n2976 185
R16089 vdd.n2629 vdd.n773 185
R16090 vdd.n774 vdd.n773 185
R16091 vdd.n2630 vdd.n809 185
R16092 vdd.n2906 vdd.n809 185
R16093 vdd.n2632 vdd.n2631 185
R16094 vdd.n2631 vdd.n817 185
R16095 vdd.n2633 vdd.n816 185
R16096 vdd.n2900 vdd.n816 185
R16097 vdd.n2635 vdd.n2634 185
R16098 vdd.n2634 vdd.n814 185
R16099 vdd.n2636 vdd.n824 185
R16100 vdd.n2849 vdd.n824 185
R16101 vdd.n2638 vdd.n2637 185
R16102 vdd.n2637 vdd.n822 185
R16103 vdd.n2639 vdd.n830 185
R16104 vdd.n2843 vdd.n830 185
R16105 vdd.n2641 vdd.n2640 185
R16106 vdd.n2640 vdd.n828 185
R16107 vdd.n2642 vdd.n835 185
R16108 vdd.n2835 vdd.n835 185
R16109 vdd.n2644 vdd.n2643 185
R16110 vdd.n2643 vdd.n841 185
R16111 vdd.n2645 vdd.n840 185
R16112 vdd.n2829 vdd.n840 185
R16113 vdd.n2679 vdd.n2678 185
R16114 vdd.n2678 vdd.n2677 185
R16115 vdd.n2680 vdd.n847 185
R16116 vdd.n2823 vdd.n847 185
R16117 vdd.n2682 vdd.n2681 185
R16118 vdd.n2681 vdd.n845 185
R16119 vdd.n2683 vdd.n853 185
R16120 vdd.n2817 vdd.n853 185
R16121 vdd.n2685 vdd.n2684 185
R16122 vdd.n2684 vdd.n851 185
R16123 vdd.n2686 vdd.n858 185
R16124 vdd.n2811 vdd.n858 185
R16125 vdd.n2688 vdd.n2687 185
R16126 vdd.n2687 vdd.n864 185
R16127 vdd.n2689 vdd.n863 185
R16128 vdd.n2805 vdd.n863 185
R16129 vdd.n2691 vdd.n2690 185
R16130 vdd.n2690 vdd.n871 185
R16131 vdd.n2692 vdd.n870 185
R16132 vdd.n2799 vdd.n870 185
R16133 vdd.n2694 vdd.n2693 185
R16134 vdd.n2693 vdd.n868 185
R16135 vdd.n2695 vdd.n876 185
R16136 vdd.n2793 vdd.n876 185
R16137 vdd.n2697 vdd.n2696 185
R16138 vdd.n2698 vdd.n2697 185
R16139 vdd.n2628 vdd.n881 185
R16140 vdd.n2787 vdd.n881 185
R16141 vdd.n2627 vdd.n2626 185
R16142 vdd.n2626 vdd.t34 185
R16143 vdd.n2625 vdd.n886 185
R16144 vdd.n2781 vdd.n886 185
R16145 vdd.n2245 vdd.n2244 185
R16146 vdd.n2246 vdd.n2245 185
R16147 vdd.n1048 vdd.n1046 185
R16148 vdd.n1046 vdd.n1044 185
R16149 vdd.n1814 vdd.n1813 185
R16150 vdd.n1813 vdd.n1812 185
R16151 vdd.n1051 vdd.n1050 185
R16152 vdd.n1052 vdd.n1051 185
R16153 vdd.n1801 vdd.n1800 185
R16154 vdd.n1802 vdd.n1801 185
R16155 vdd.n1060 vdd.n1059 185
R16156 vdd.n1793 vdd.n1059 185
R16157 vdd.n1796 vdd.n1795 185
R16158 vdd.n1795 vdd.n1794 185
R16159 vdd.n1063 vdd.n1062 185
R16160 vdd.n1069 vdd.n1063 185
R16161 vdd.n1784 vdd.n1783 185
R16162 vdd.n1785 vdd.n1784 185
R16163 vdd.n1071 vdd.n1070 185
R16164 vdd.n1776 vdd.n1070 185
R16165 vdd.n1779 vdd.n1778 185
R16166 vdd.n1778 vdd.n1777 185
R16167 vdd.n1074 vdd.n1073 185
R16168 vdd.n1075 vdd.n1074 185
R16169 vdd.n1767 vdd.n1766 185
R16170 vdd.n1768 vdd.n1767 185
R16171 vdd.n1083 vdd.n1082 185
R16172 vdd.n1082 vdd.n1081 185
R16173 vdd.n1762 vdd.n1761 185
R16174 vdd.n1761 vdd.n1760 185
R16175 vdd.n1086 vdd.n1085 185
R16176 vdd.n1092 vdd.n1086 185
R16177 vdd.n1751 vdd.n1750 185
R16178 vdd.n1752 vdd.n1751 185
R16179 vdd.n1094 vdd.n1093 185
R16180 vdd.n1448 vdd.n1093 185
R16181 vdd.n1451 vdd.n1450 185
R16182 vdd.n1450 vdd.n1449 185
R16183 vdd.n1097 vdd.n1096 185
R16184 vdd.n1104 vdd.n1097 185
R16185 vdd.n1439 vdd.n1438 185
R16186 vdd.n1440 vdd.n1439 185
R16187 vdd.n1106 vdd.n1105 185
R16188 vdd.n1105 vdd.n1103 185
R16189 vdd.n1434 vdd.n1433 185
R16190 vdd.n1433 vdd.n1432 185
R16191 vdd.n1109 vdd.n1108 185
R16192 vdd.n1110 vdd.n1109 185
R16193 vdd.n1423 vdd.n1422 185
R16194 vdd.n1424 vdd.n1423 185
R16195 vdd.n1117 vdd.n1116 185
R16196 vdd.n1415 vdd.n1116 185
R16197 vdd.n1418 vdd.n1417 185
R16198 vdd.n1417 vdd.n1416 185
R16199 vdd.n1120 vdd.n1119 185
R16200 vdd.n1126 vdd.n1120 185
R16201 vdd.n1406 vdd.n1405 185
R16202 vdd.n1407 vdd.n1406 185
R16203 vdd.n1128 vdd.n1127 185
R16204 vdd.n1398 vdd.n1127 185
R16205 vdd.n1401 vdd.n1400 185
R16206 vdd.n1400 vdd.n1399 185
R16207 vdd.n1131 vdd.n1130 185
R16208 vdd.n1132 vdd.n1131 185
R16209 vdd.n1389 vdd.n1388 185
R16210 vdd.n1390 vdd.n1389 185
R16211 vdd.n1140 vdd.n1139 185
R16212 vdd.n1139 vdd.n1138 185
R16213 vdd.n1384 vdd.n1383 185
R16214 vdd.n1383 vdd.n1382 185
R16215 vdd.n1143 vdd.n1142 185
R16216 vdd.n1144 vdd.n1143 185
R16217 vdd.n1372 vdd.n1371 185
R16218 vdd.n1370 vdd.n1183 185
R16219 vdd.n1185 vdd.n1182 185
R16220 vdd.n1374 vdd.n1182 185
R16221 vdd.n1366 vdd.n1187 185
R16222 vdd.n1365 vdd.n1188 185
R16223 vdd.n1364 vdd.n1189 185
R16224 vdd.n1192 vdd.n1190 185
R16225 vdd.n1360 vdd.n1193 185
R16226 vdd.n1359 vdd.n1194 185
R16227 vdd.n1358 vdd.n1195 185
R16228 vdd.n1198 vdd.n1196 185
R16229 vdd.n1354 vdd.n1199 185
R16230 vdd.n1353 vdd.n1200 185
R16231 vdd.n1352 vdd.n1201 185
R16232 vdd.n1204 vdd.n1202 185
R16233 vdd.n1348 vdd.n1205 185
R16234 vdd.n1347 vdd.n1206 185
R16235 vdd.n1346 vdd.n1207 185
R16236 vdd.n1338 vdd.n1208 185
R16237 vdd.n1342 vdd.n1339 185
R16238 vdd.n1337 vdd.n1210 185
R16239 vdd.n1336 vdd.n1211 185
R16240 vdd.n1214 vdd.n1212 185
R16241 vdd.n1332 vdd.n1215 185
R16242 vdd.n1331 vdd.n1216 185
R16243 vdd.n1330 vdd.n1217 185
R16244 vdd.n1220 vdd.n1218 185
R16245 vdd.n1326 vdd.n1221 185
R16246 vdd.n1325 vdd.n1222 185
R16247 vdd.n1324 vdd.n1223 185
R16248 vdd.n1226 vdd.n1224 185
R16249 vdd.n1320 vdd.n1227 185
R16250 vdd.n1319 vdd.n1228 185
R16251 vdd.n1318 vdd.n1229 185
R16252 vdd.n1232 vdd.n1230 185
R16253 vdd.n1314 vdd.n1233 185
R16254 vdd.n1313 vdd.n1234 185
R16255 vdd.n1312 vdd.n1235 185
R16256 vdd.n1238 vdd.n1236 185
R16257 vdd.n1308 vdd.n1239 185
R16258 vdd.n1307 vdd.n1240 185
R16259 vdd.n1306 vdd.n1303 185
R16260 vdd.n1243 vdd.n1241 185
R16261 vdd.n1299 vdd.n1244 185
R16262 vdd.n1298 vdd.n1245 185
R16263 vdd.n1297 vdd.n1246 185
R16264 vdd.n1249 vdd.n1247 185
R16265 vdd.n1293 vdd.n1250 185
R16266 vdd.n1292 vdd.n1251 185
R16267 vdd.n1291 vdd.n1252 185
R16268 vdd.n1255 vdd.n1253 185
R16269 vdd.n1287 vdd.n1256 185
R16270 vdd.n1286 vdd.n1257 185
R16271 vdd.n1285 vdd.n1258 185
R16272 vdd.n1261 vdd.n1259 185
R16273 vdd.n1281 vdd.n1262 185
R16274 vdd.n1280 vdd.n1263 185
R16275 vdd.n1279 vdd.n1264 185
R16276 vdd.n1267 vdd.n1265 185
R16277 vdd.n1275 vdd.n1268 185
R16278 vdd.n1274 vdd.n1269 185
R16279 vdd.n1273 vdd.n1270 185
R16280 vdd.n1271 vdd.n1151 185
R16281 vdd.n1376 vdd.n1375 185
R16282 vdd.n1375 vdd.n1374 185
R16283 vdd.n2249 vdd.n2248 185
R16284 vdd.n2253 vdd.n1040 185
R16285 vdd.n1916 vdd.n1039 185
R16286 vdd.n1919 vdd.n1918 185
R16287 vdd.n1921 vdd.n1920 185
R16288 vdd.n1924 vdd.n1923 185
R16289 vdd.n1926 vdd.n1925 185
R16290 vdd.n1928 vdd.n1914 185
R16291 vdd.n1930 vdd.n1929 185
R16292 vdd.n1931 vdd.n1908 185
R16293 vdd.n1933 vdd.n1932 185
R16294 vdd.n1935 vdd.n1906 185
R16295 vdd.n1937 vdd.n1936 185
R16296 vdd.n1938 vdd.n1901 185
R16297 vdd.n1940 vdd.n1939 185
R16298 vdd.n1942 vdd.n1899 185
R16299 vdd.n1944 vdd.n1943 185
R16300 vdd.n1945 vdd.n1895 185
R16301 vdd.n1947 vdd.n1946 185
R16302 vdd.n1949 vdd.n1892 185
R16303 vdd.n1951 vdd.n1950 185
R16304 vdd.n1893 vdd.n1886 185
R16305 vdd.n1955 vdd.n1890 185
R16306 vdd.n1956 vdd.n1882 185
R16307 vdd.n1958 vdd.n1957 185
R16308 vdd.n1960 vdd.n1880 185
R16309 vdd.n1962 vdd.n1961 185
R16310 vdd.n1963 vdd.n1875 185
R16311 vdd.n1965 vdd.n1964 185
R16312 vdd.n1967 vdd.n1873 185
R16313 vdd.n1969 vdd.n1968 185
R16314 vdd.n1970 vdd.n1868 185
R16315 vdd.n1972 vdd.n1971 185
R16316 vdd.n1974 vdd.n1866 185
R16317 vdd.n1976 vdd.n1975 185
R16318 vdd.n1977 vdd.n1861 185
R16319 vdd.n1979 vdd.n1978 185
R16320 vdd.n1981 vdd.n1859 185
R16321 vdd.n1983 vdd.n1982 185
R16322 vdd.n1984 vdd.n1855 185
R16323 vdd.n1986 vdd.n1985 185
R16324 vdd.n1988 vdd.n1852 185
R16325 vdd.n1990 vdd.n1989 185
R16326 vdd.n1853 vdd.n1846 185
R16327 vdd.n1994 vdd.n1850 185
R16328 vdd.n1995 vdd.n1842 185
R16329 vdd.n1997 vdd.n1996 185
R16330 vdd.n1999 vdd.n1840 185
R16331 vdd.n2001 vdd.n2000 185
R16332 vdd.n2002 vdd.n1835 185
R16333 vdd.n2004 vdd.n2003 185
R16334 vdd.n2006 vdd.n1833 185
R16335 vdd.n2008 vdd.n2007 185
R16336 vdd.n2009 vdd.n1828 185
R16337 vdd.n2011 vdd.n2010 185
R16338 vdd.n2013 vdd.n1827 185
R16339 vdd.n2014 vdd.n1824 185
R16340 vdd.n2017 vdd.n2016 185
R16341 vdd.n1826 vdd.n1822 185
R16342 vdd.n2234 vdd.n1820 185
R16343 vdd.n2236 vdd.n2235 185
R16344 vdd.n2238 vdd.n1818 185
R16345 vdd.n2240 vdd.n2239 185
R16346 vdd.n2241 vdd.n1047 185
R16347 vdd.n2247 vdd.n1043 185
R16348 vdd.n2247 vdd.n2246 185
R16349 vdd.n1055 vdd.n1042 185
R16350 vdd.n1044 vdd.n1042 185
R16351 vdd.n1811 vdd.n1810 185
R16352 vdd.n1812 vdd.n1811 185
R16353 vdd.n1054 vdd.n1053 185
R16354 vdd.n1053 vdd.n1052 185
R16355 vdd.n1804 vdd.n1803 185
R16356 vdd.n1803 vdd.n1802 185
R16357 vdd.n1058 vdd.n1057 185
R16358 vdd.n1793 vdd.n1058 185
R16359 vdd.n1792 vdd.n1791 185
R16360 vdd.n1794 vdd.n1792 185
R16361 vdd.n1065 vdd.n1064 185
R16362 vdd.n1069 vdd.n1064 185
R16363 vdd.n1787 vdd.n1786 185
R16364 vdd.n1786 vdd.n1785 185
R16365 vdd.n1068 vdd.n1067 185
R16366 vdd.n1776 vdd.n1068 185
R16367 vdd.n1775 vdd.n1774 185
R16368 vdd.n1777 vdd.n1775 185
R16369 vdd.n1077 vdd.n1076 185
R16370 vdd.n1076 vdd.n1075 185
R16371 vdd.n1770 vdd.n1769 185
R16372 vdd.n1769 vdd.n1768 185
R16373 vdd.n1080 vdd.n1079 185
R16374 vdd.n1081 vdd.n1080 185
R16375 vdd.n1759 vdd.n1758 185
R16376 vdd.n1760 vdd.n1759 185
R16377 vdd.n1088 vdd.n1087 185
R16378 vdd.n1092 vdd.n1087 185
R16379 vdd.n1754 vdd.n1753 185
R16380 vdd.n1753 vdd.n1752 185
R16381 vdd.n1091 vdd.n1090 185
R16382 vdd.n1448 vdd.n1091 185
R16383 vdd.n1447 vdd.n1446 185
R16384 vdd.n1449 vdd.n1447 185
R16385 vdd.n1099 vdd.n1098 185
R16386 vdd.n1104 vdd.n1098 185
R16387 vdd.n1442 vdd.n1441 185
R16388 vdd.n1441 vdd.n1440 185
R16389 vdd.n1102 vdd.n1101 185
R16390 vdd.n1103 vdd.n1102 185
R16391 vdd.n1431 vdd.n1430 185
R16392 vdd.n1432 vdd.n1431 185
R16393 vdd.n1112 vdd.n1111 185
R16394 vdd.n1111 vdd.n1110 185
R16395 vdd.n1426 vdd.n1425 185
R16396 vdd.n1425 vdd.n1424 185
R16397 vdd.n1115 vdd.n1114 185
R16398 vdd.n1415 vdd.n1115 185
R16399 vdd.n1414 vdd.n1413 185
R16400 vdd.n1416 vdd.n1414 185
R16401 vdd.n1122 vdd.n1121 185
R16402 vdd.n1126 vdd.n1121 185
R16403 vdd.n1409 vdd.n1408 185
R16404 vdd.n1408 vdd.n1407 185
R16405 vdd.n1125 vdd.n1124 185
R16406 vdd.n1398 vdd.n1125 185
R16407 vdd.n1397 vdd.n1396 185
R16408 vdd.n1399 vdd.n1397 185
R16409 vdd.n1134 vdd.n1133 185
R16410 vdd.n1133 vdd.n1132 185
R16411 vdd.n1392 vdd.n1391 185
R16412 vdd.n1391 vdd.n1390 185
R16413 vdd.n1137 vdd.n1136 185
R16414 vdd.n1138 vdd.n1137 185
R16415 vdd.n1381 vdd.n1380 185
R16416 vdd.n1382 vdd.n1381 185
R16417 vdd.n1146 vdd.n1145 185
R16418 vdd.n1145 vdd.n1144 185
R16419 vdd.n927 vdd.n925 185
R16420 vdd.n2449 vdd.n925 185
R16421 vdd.n2371 vdd.n944 185
R16422 vdd.n944 vdd.t8 185
R16423 vdd.n2373 vdd.n2372 185
R16424 vdd.n2374 vdd.n2373 185
R16425 vdd.n2370 vdd.n943 185
R16426 vdd.n2073 vdd.n943 185
R16427 vdd.n2369 vdd.n2368 185
R16428 vdd.n2368 vdd.n2367 185
R16429 vdd.n946 vdd.n945 185
R16430 vdd.n947 vdd.n946 185
R16431 vdd.n2358 vdd.n2357 185
R16432 vdd.n2359 vdd.n2358 185
R16433 vdd.n2356 vdd.n957 185
R16434 vdd.n957 vdd.n954 185
R16435 vdd.n2355 vdd.n2354 185
R16436 vdd.n2354 vdd.n2353 185
R16437 vdd.n959 vdd.n958 185
R16438 vdd.n960 vdd.n959 185
R16439 vdd.n2346 vdd.n2345 185
R16440 vdd.n2347 vdd.n2346 185
R16441 vdd.n2344 vdd.n968 185
R16442 vdd.n973 vdd.n968 185
R16443 vdd.n2343 vdd.n2342 185
R16444 vdd.n2342 vdd.n2341 185
R16445 vdd.n970 vdd.n969 185
R16446 vdd.n979 vdd.n970 185
R16447 vdd.n2334 vdd.n2333 185
R16448 vdd.n2335 vdd.n2334 185
R16449 vdd.n2332 vdd.n980 185
R16450 vdd.n2174 vdd.n980 185
R16451 vdd.n2331 vdd.n2330 185
R16452 vdd.n2330 vdd.n2329 185
R16453 vdd.n982 vdd.n981 185
R16454 vdd.n983 vdd.n982 185
R16455 vdd.n2322 vdd.n2321 185
R16456 vdd.n2323 vdd.n2322 185
R16457 vdd.n2320 vdd.n992 185
R16458 vdd.n992 vdd.n989 185
R16459 vdd.n2319 vdd.n2318 185
R16460 vdd.n2318 vdd.n2317 185
R16461 vdd.n994 vdd.n993 185
R16462 vdd.n1004 vdd.n994 185
R16463 vdd.n2309 vdd.n2308 185
R16464 vdd.n2310 vdd.n2309 185
R16465 vdd.n2307 vdd.n1005 185
R16466 vdd.n1005 vdd.n1001 185
R16467 vdd.n2306 vdd.n2305 185
R16468 vdd.n2305 vdd.n2304 185
R16469 vdd.n1007 vdd.n1006 185
R16470 vdd.n1008 vdd.n1007 185
R16471 vdd.n2297 vdd.n2296 185
R16472 vdd.n2298 vdd.n2297 185
R16473 vdd.n2295 vdd.n1017 185
R16474 vdd.n1017 vdd.n1014 185
R16475 vdd.n2294 vdd.n2293 185
R16476 vdd.n2293 vdd.n2292 185
R16477 vdd.n1019 vdd.n1018 185
R16478 vdd.n2029 vdd.n2028 185
R16479 vdd.n2030 vdd.n2026 185
R16480 vdd.n2026 vdd.n1020 185
R16481 vdd.n2032 vdd.n2031 185
R16482 vdd.n2034 vdd.n2025 185
R16483 vdd.n2037 vdd.n2036 185
R16484 vdd.n2038 vdd.n2024 185
R16485 vdd.n2040 vdd.n2039 185
R16486 vdd.n2042 vdd.n2023 185
R16487 vdd.n2045 vdd.n2044 185
R16488 vdd.n2046 vdd.n2022 185
R16489 vdd.n2048 vdd.n2047 185
R16490 vdd.n2050 vdd.n2021 185
R16491 vdd.n2053 vdd.n2052 185
R16492 vdd.n2054 vdd.n2020 185
R16493 vdd.n2056 vdd.n2055 185
R16494 vdd.n2058 vdd.n2019 185
R16495 vdd.n2231 vdd.n2059 185
R16496 vdd.n2230 vdd.n2229 185
R16497 vdd.n2227 vdd.n2060 185
R16498 vdd.n2225 vdd.n2224 185
R16499 vdd.n2223 vdd.n2061 185
R16500 vdd.n2222 vdd.n2221 185
R16501 vdd.n2219 vdd.n2062 185
R16502 vdd.n2217 vdd.n2216 185
R16503 vdd.n2215 vdd.n2063 185
R16504 vdd.n2214 vdd.n2213 185
R16505 vdd.n2211 vdd.n2064 185
R16506 vdd.n2209 vdd.n2208 185
R16507 vdd.n2207 vdd.n2065 185
R16508 vdd.n2206 vdd.n2205 185
R16509 vdd.n2203 vdd.n2066 185
R16510 vdd.n2201 vdd.n2200 185
R16511 vdd.n2199 vdd.n2067 185
R16512 vdd.n2198 vdd.n2197 185
R16513 vdd.n2452 vdd.n2451 185
R16514 vdd.n2454 vdd.n2453 185
R16515 vdd.n2456 vdd.n2455 185
R16516 vdd.n2459 vdd.n2458 185
R16517 vdd.n2461 vdd.n2460 185
R16518 vdd.n2463 vdd.n2462 185
R16519 vdd.n2465 vdd.n2464 185
R16520 vdd.n2467 vdd.n2466 185
R16521 vdd.n2469 vdd.n2468 185
R16522 vdd.n2471 vdd.n2470 185
R16523 vdd.n2473 vdd.n2472 185
R16524 vdd.n2475 vdd.n2474 185
R16525 vdd.n2477 vdd.n2476 185
R16526 vdd.n2479 vdd.n2478 185
R16527 vdd.n2481 vdd.n2480 185
R16528 vdd.n2483 vdd.n2482 185
R16529 vdd.n2485 vdd.n2484 185
R16530 vdd.n2487 vdd.n2486 185
R16531 vdd.n2489 vdd.n2488 185
R16532 vdd.n2491 vdd.n2490 185
R16533 vdd.n2493 vdd.n2492 185
R16534 vdd.n2495 vdd.n2494 185
R16535 vdd.n2497 vdd.n2496 185
R16536 vdd.n2499 vdd.n2498 185
R16537 vdd.n2501 vdd.n2500 185
R16538 vdd.n2503 vdd.n2502 185
R16539 vdd.n2505 vdd.n2504 185
R16540 vdd.n2507 vdd.n2506 185
R16541 vdd.n2509 vdd.n2508 185
R16542 vdd.n2511 vdd.n2510 185
R16543 vdd.n2513 vdd.n2512 185
R16544 vdd.n2515 vdd.n2514 185
R16545 vdd.n2517 vdd.n2516 185
R16546 vdd.n2518 vdd.n926 185
R16547 vdd.n2520 vdd.n2519 185
R16548 vdd.n2521 vdd.n2520 185
R16549 vdd.n2450 vdd.n930 185
R16550 vdd.n2450 vdd.n2449 185
R16551 vdd.n2071 vdd.n931 185
R16552 vdd.t8 vdd.n931 185
R16553 vdd.n2072 vdd.n941 185
R16554 vdd.n2374 vdd.n941 185
R16555 vdd.n2075 vdd.n2074 185
R16556 vdd.n2074 vdd.n2073 185
R16557 vdd.n2076 vdd.n948 185
R16558 vdd.n2367 vdd.n948 185
R16559 vdd.n2078 vdd.n2077 185
R16560 vdd.n2077 vdd.n947 185
R16561 vdd.n2079 vdd.n955 185
R16562 vdd.n2359 vdd.n955 185
R16563 vdd.n2081 vdd.n2080 185
R16564 vdd.n2080 vdd.n954 185
R16565 vdd.n2082 vdd.n961 185
R16566 vdd.n2353 vdd.n961 185
R16567 vdd.n2084 vdd.n2083 185
R16568 vdd.n2083 vdd.n960 185
R16569 vdd.n2085 vdd.n966 185
R16570 vdd.n2347 vdd.n966 185
R16571 vdd.n2087 vdd.n2086 185
R16572 vdd.n2086 vdd.n973 185
R16573 vdd.n2088 vdd.n971 185
R16574 vdd.n2341 vdd.n971 185
R16575 vdd.n2090 vdd.n2089 185
R16576 vdd.n2089 vdd.n979 185
R16577 vdd.n2091 vdd.n977 185
R16578 vdd.n2335 vdd.n977 185
R16579 vdd.n2176 vdd.n2175 185
R16580 vdd.n2175 vdd.n2174 185
R16581 vdd.n2177 vdd.n984 185
R16582 vdd.n2329 vdd.n984 185
R16583 vdd.n2179 vdd.n2178 185
R16584 vdd.n2178 vdd.n983 185
R16585 vdd.n2180 vdd.n990 185
R16586 vdd.n2323 vdd.n990 185
R16587 vdd.n2182 vdd.n2181 185
R16588 vdd.n2181 vdd.n989 185
R16589 vdd.n2183 vdd.n995 185
R16590 vdd.n2317 vdd.n995 185
R16591 vdd.n2185 vdd.n2184 185
R16592 vdd.n2184 vdd.n1004 185
R16593 vdd.n2186 vdd.n1002 185
R16594 vdd.n2310 vdd.n1002 185
R16595 vdd.n2188 vdd.n2187 185
R16596 vdd.n2187 vdd.n1001 185
R16597 vdd.n2189 vdd.n1009 185
R16598 vdd.n2304 vdd.n1009 185
R16599 vdd.n2191 vdd.n2190 185
R16600 vdd.n2190 vdd.n1008 185
R16601 vdd.n2192 vdd.n1015 185
R16602 vdd.n2298 vdd.n1015 185
R16603 vdd.n2194 vdd.n2193 185
R16604 vdd.n2193 vdd.n1014 185
R16605 vdd.n2195 vdd.n1021 185
R16606 vdd.n2292 vdd.n1021 185
R16607 vdd.n370 vdd.n369 185
R16608 vdd.n3254 vdd.n370 185
R16609 vdd.n3257 vdd.n3256 185
R16610 vdd.n3256 vdd.n3255 185
R16611 vdd.n3258 vdd.n364 185
R16612 vdd.n364 vdd.n363 185
R16613 vdd.n3260 vdd.n3259 185
R16614 vdd.n3261 vdd.n3260 185
R16615 vdd.n359 vdd.n358 185
R16616 vdd.n3262 vdd.n359 185
R16617 vdd.n3265 vdd.n3264 185
R16618 vdd.n3264 vdd.n3263 185
R16619 vdd.n3266 vdd.n353 185
R16620 vdd.n3236 vdd.n353 185
R16621 vdd.n3268 vdd.n3267 185
R16622 vdd.n3269 vdd.n3268 185
R16623 vdd.n348 vdd.n347 185
R16624 vdd.n3270 vdd.n348 185
R16625 vdd.n3273 vdd.n3272 185
R16626 vdd.n3272 vdd.n3271 185
R16627 vdd.n3274 vdd.n342 185
R16628 vdd.n349 vdd.n342 185
R16629 vdd.n3276 vdd.n3275 185
R16630 vdd.n3277 vdd.n3276 185
R16631 vdd.n338 vdd.n337 185
R16632 vdd.n3278 vdd.n338 185
R16633 vdd.n3281 vdd.n3280 185
R16634 vdd.n3280 vdd.n3279 185
R16635 vdd.n3282 vdd.n333 185
R16636 vdd.n333 vdd.n332 185
R16637 vdd.n3284 vdd.n3283 185
R16638 vdd.n3285 vdd.n3284 185
R16639 vdd.n327 vdd.n325 185
R16640 vdd.n3286 vdd.n327 185
R16641 vdd.n3289 vdd.n3288 185
R16642 vdd.n3288 vdd.n3287 185
R16643 vdd.n326 vdd.n324 185
R16644 vdd.n328 vdd.n326 185
R16645 vdd.n3212 vdd.n3211 185
R16646 vdd.n3213 vdd.n3212 185
R16647 vdd.n615 vdd.n614 185
R16648 vdd.n614 vdd.n613 185
R16649 vdd.n3207 vdd.n3206 185
R16650 vdd.n3206 vdd.n3205 185
R16651 vdd.n618 vdd.n617 185
R16652 vdd.n624 vdd.n618 185
R16653 vdd.n3193 vdd.n3192 185
R16654 vdd.n3194 vdd.n3193 185
R16655 vdd.n626 vdd.n625 185
R16656 vdd.n3185 vdd.n625 185
R16657 vdd.n3188 vdd.n3187 185
R16658 vdd.n3187 vdd.n3186 185
R16659 vdd.n629 vdd.n628 185
R16660 vdd.n636 vdd.n629 185
R16661 vdd.n3176 vdd.n3175 185
R16662 vdd.n3177 vdd.n3176 185
R16663 vdd.n638 vdd.n637 185
R16664 vdd.n637 vdd.n635 185
R16665 vdd.n3171 vdd.n3170 185
R16666 vdd.n3170 vdd.n3169 185
R16667 vdd.n641 vdd.n640 185
R16668 vdd.n642 vdd.n641 185
R16669 vdd.n3160 vdd.n3159 185
R16670 vdd.n3161 vdd.n3160 185
R16671 vdd.n650 vdd.n649 185
R16672 vdd.n649 vdd.n648 185
R16673 vdd.n3155 vdd.n3154 185
R16674 vdd.n3154 vdd.n3153 185
R16675 vdd.n653 vdd.n652 185
R16676 vdd.n659 vdd.n653 185
R16677 vdd.n3144 vdd.n3143 185
R16678 vdd.n3145 vdd.n3144 185
R16679 vdd.n3140 vdd.n660 185
R16680 vdd.n3139 vdd.n3138 185
R16681 vdd.n3136 vdd.n662 185
R16682 vdd.n3136 vdd.n658 185
R16683 vdd.n3135 vdd.n3134 185
R16684 vdd.n3133 vdd.n3132 185
R16685 vdd.n3131 vdd.n3130 185
R16686 vdd.n3129 vdd.n3128 185
R16687 vdd.n3127 vdd.n668 185
R16688 vdd.n3125 vdd.n3124 185
R16689 vdd.n3123 vdd.n669 185
R16690 vdd.n3122 vdd.n3121 185
R16691 vdd.n3119 vdd.n674 185
R16692 vdd.n3117 vdd.n3116 185
R16693 vdd.n3115 vdd.n675 185
R16694 vdd.n3114 vdd.n3113 185
R16695 vdd.n3111 vdd.n680 185
R16696 vdd.n3109 vdd.n3108 185
R16697 vdd.n3107 vdd.n681 185
R16698 vdd.n3106 vdd.n3105 185
R16699 vdd.n3103 vdd.n688 185
R16700 vdd.n3101 vdd.n3100 185
R16701 vdd.n3099 vdd.n689 185
R16702 vdd.n3098 vdd.n3097 185
R16703 vdd.n3095 vdd.n694 185
R16704 vdd.n3093 vdd.n3092 185
R16705 vdd.n3091 vdd.n695 185
R16706 vdd.n3090 vdd.n3089 185
R16707 vdd.n3087 vdd.n700 185
R16708 vdd.n3085 vdd.n3084 185
R16709 vdd.n3083 vdd.n701 185
R16710 vdd.n3082 vdd.n3081 185
R16711 vdd.n3079 vdd.n706 185
R16712 vdd.n3077 vdd.n3076 185
R16713 vdd.n3075 vdd.n707 185
R16714 vdd.n3074 vdd.n3073 185
R16715 vdd.n3071 vdd.n712 185
R16716 vdd.n3069 vdd.n3068 185
R16717 vdd.n3067 vdd.n713 185
R16718 vdd.n3066 vdd.n3065 185
R16719 vdd.n3063 vdd.n718 185
R16720 vdd.n3061 vdd.n3060 185
R16721 vdd.n3059 vdd.n719 185
R16722 vdd.n728 vdd.n722 185
R16723 vdd.n3055 vdd.n3054 185
R16724 vdd.n3052 vdd.n726 185
R16725 vdd.n3051 vdd.n3050 185
R16726 vdd.n3049 vdd.n3048 185
R16727 vdd.n3047 vdd.n732 185
R16728 vdd.n3045 vdd.n3044 185
R16729 vdd.n3043 vdd.n733 185
R16730 vdd.n3042 vdd.n3041 185
R16731 vdd.n3039 vdd.n738 185
R16732 vdd.n3037 vdd.n3036 185
R16733 vdd.n3035 vdd.n739 185
R16734 vdd.n3034 vdd.n3033 185
R16735 vdd.n3031 vdd.n744 185
R16736 vdd.n3029 vdd.n3028 185
R16737 vdd.n3027 vdd.n745 185
R16738 vdd.n3026 vdd.n3025 185
R16739 vdd.n3023 vdd.n3022 185
R16740 vdd.n3021 vdd.n3020 185
R16741 vdd.n3019 vdd.n3018 185
R16742 vdd.n3017 vdd.n3016 185
R16743 vdd.n3012 vdd.n657 185
R16744 vdd.n658 vdd.n657 185
R16745 vdd.n3251 vdd.n3250 185
R16746 vdd.n599 vdd.n404 185
R16747 vdd.n598 vdd.n597 185
R16748 vdd.n596 vdd.n595 185
R16749 vdd.n594 vdd.n409 185
R16750 vdd.n590 vdd.n589 185
R16751 vdd.n588 vdd.n587 185
R16752 vdd.n586 vdd.n585 185
R16753 vdd.n584 vdd.n411 185
R16754 vdd.n580 vdd.n579 185
R16755 vdd.n578 vdd.n577 185
R16756 vdd.n576 vdd.n575 185
R16757 vdd.n574 vdd.n413 185
R16758 vdd.n570 vdd.n569 185
R16759 vdd.n568 vdd.n567 185
R16760 vdd.n566 vdd.n565 185
R16761 vdd.n564 vdd.n415 185
R16762 vdd.n560 vdd.n559 185
R16763 vdd.n558 vdd.n557 185
R16764 vdd.n556 vdd.n555 185
R16765 vdd.n554 vdd.n417 185
R16766 vdd.n550 vdd.n549 185
R16767 vdd.n548 vdd.n547 185
R16768 vdd.n546 vdd.n545 185
R16769 vdd.n544 vdd.n421 185
R16770 vdd.n540 vdd.n539 185
R16771 vdd.n538 vdd.n537 185
R16772 vdd.n536 vdd.n535 185
R16773 vdd.n534 vdd.n423 185
R16774 vdd.n530 vdd.n529 185
R16775 vdd.n528 vdd.n527 185
R16776 vdd.n526 vdd.n525 185
R16777 vdd.n524 vdd.n425 185
R16778 vdd.n520 vdd.n519 185
R16779 vdd.n518 vdd.n517 185
R16780 vdd.n516 vdd.n515 185
R16781 vdd.n514 vdd.n427 185
R16782 vdd.n510 vdd.n509 185
R16783 vdd.n508 vdd.n507 185
R16784 vdd.n506 vdd.n505 185
R16785 vdd.n504 vdd.n429 185
R16786 vdd.n500 vdd.n499 185
R16787 vdd.n498 vdd.n497 185
R16788 vdd.n496 vdd.n495 185
R16789 vdd.n494 vdd.n433 185
R16790 vdd.n490 vdd.n489 185
R16791 vdd.n488 vdd.n487 185
R16792 vdd.n486 vdd.n485 185
R16793 vdd.n484 vdd.n435 185
R16794 vdd.n480 vdd.n479 185
R16795 vdd.n478 vdd.n477 185
R16796 vdd.n476 vdd.n475 185
R16797 vdd.n474 vdd.n437 185
R16798 vdd.n470 vdd.n469 185
R16799 vdd.n468 vdd.n467 185
R16800 vdd.n466 vdd.n465 185
R16801 vdd.n464 vdd.n439 185
R16802 vdd.n460 vdd.n459 185
R16803 vdd.n458 vdd.n457 185
R16804 vdd.n456 vdd.n455 185
R16805 vdd.n454 vdd.n441 185
R16806 vdd.n450 vdd.n449 185
R16807 vdd.n448 vdd.n447 185
R16808 vdd.n446 vdd.n445 185
R16809 vdd.n3247 vdd.n372 185
R16810 vdd.n3254 vdd.n372 185
R16811 vdd.n3246 vdd.n371 185
R16812 vdd.n3255 vdd.n371 185
R16813 vdd.n3245 vdd.n3244 185
R16814 vdd.n3244 vdd.n363 185
R16815 vdd.n602 vdd.n362 185
R16816 vdd.n3261 vdd.n362 185
R16817 vdd.n3240 vdd.n361 185
R16818 vdd.n3262 vdd.n361 185
R16819 vdd.n3239 vdd.n360 185
R16820 vdd.n3263 vdd.n360 185
R16821 vdd.n3238 vdd.n3237 185
R16822 vdd.n3237 vdd.n3236 185
R16823 vdd.n604 vdd.n352 185
R16824 vdd.n3269 vdd.n352 185
R16825 vdd.n3232 vdd.n351 185
R16826 vdd.n3270 vdd.n351 185
R16827 vdd.n3231 vdd.n350 185
R16828 vdd.n3271 vdd.n350 185
R16829 vdd.n3230 vdd.n3229 185
R16830 vdd.n3229 vdd.n349 185
R16831 vdd.n606 vdd.n341 185
R16832 vdd.n3277 vdd.n341 185
R16833 vdd.n3225 vdd.n340 185
R16834 vdd.n3278 vdd.n340 185
R16835 vdd.n3224 vdd.n339 185
R16836 vdd.n3279 vdd.n339 185
R16837 vdd.n3223 vdd.n3222 185
R16838 vdd.n3222 vdd.n332 185
R16839 vdd.n608 vdd.n331 185
R16840 vdd.n3285 vdd.n331 185
R16841 vdd.n3218 vdd.n330 185
R16842 vdd.n3286 vdd.n330 185
R16843 vdd.n3217 vdd.n329 185
R16844 vdd.n3287 vdd.n329 185
R16845 vdd.n3216 vdd.n3215 185
R16846 vdd.n3215 vdd.n328 185
R16847 vdd.n3214 vdd.n610 185
R16848 vdd.n3214 vdd.n3213 185
R16849 vdd.n3202 vdd.n612 185
R16850 vdd.n613 vdd.n612 185
R16851 vdd.n3204 vdd.n3203 185
R16852 vdd.n3205 vdd.n3204 185
R16853 vdd.n620 vdd.n619 185
R16854 vdd.n624 vdd.n619 185
R16855 vdd.n3196 vdd.n3195 185
R16856 vdd.n3195 vdd.n3194 185
R16857 vdd.n623 vdd.n622 185
R16858 vdd.n3185 vdd.n623 185
R16859 vdd.n3184 vdd.n3183 185
R16860 vdd.n3186 vdd.n3184 185
R16861 vdd.n631 vdd.n630 185
R16862 vdd.n636 vdd.n630 185
R16863 vdd.n3179 vdd.n3178 185
R16864 vdd.n3178 vdd.n3177 185
R16865 vdd.n634 vdd.n633 185
R16866 vdd.n635 vdd.n634 185
R16867 vdd.n3168 vdd.n3167 185
R16868 vdd.n3169 vdd.n3168 185
R16869 vdd.n644 vdd.n643 185
R16870 vdd.n643 vdd.n642 185
R16871 vdd.n3163 vdd.n3162 185
R16872 vdd.n3162 vdd.n3161 185
R16873 vdd.n647 vdd.n646 185
R16874 vdd.n648 vdd.n647 185
R16875 vdd.n3152 vdd.n3151 185
R16876 vdd.n3153 vdd.n3152 185
R16877 vdd.n655 vdd.n654 185
R16878 vdd.n659 vdd.n654 185
R16879 vdd.n3147 vdd.n3146 185
R16880 vdd.n3146 vdd.n3145 185
R16881 vdd.n884 vdd.n883 185
R16882 vdd.n2772 vdd.n2771 185
R16883 vdd.n2770 vdd.n2555 185
R16884 vdd.n2774 vdd.n2555 185
R16885 vdd.n2769 vdd.n2768 185
R16886 vdd.n2767 vdd.n2766 185
R16887 vdd.n2765 vdd.n2764 185
R16888 vdd.n2763 vdd.n2762 185
R16889 vdd.n2761 vdd.n2760 185
R16890 vdd.n2759 vdd.n2758 185
R16891 vdd.n2757 vdd.n2756 185
R16892 vdd.n2755 vdd.n2754 185
R16893 vdd.n2753 vdd.n2752 185
R16894 vdd.n2751 vdd.n2750 185
R16895 vdd.n2749 vdd.n2748 185
R16896 vdd.n2747 vdd.n2746 185
R16897 vdd.n2745 vdd.n2744 185
R16898 vdd.n2743 vdd.n2742 185
R16899 vdd.n2741 vdd.n2740 185
R16900 vdd.n2739 vdd.n2738 185
R16901 vdd.n2737 vdd.n2736 185
R16902 vdd.n2735 vdd.n2734 185
R16903 vdd.n2733 vdd.n2732 185
R16904 vdd.n2731 vdd.n2730 185
R16905 vdd.n2729 vdd.n2728 185
R16906 vdd.n2727 vdd.n2726 185
R16907 vdd.n2725 vdd.n2724 185
R16908 vdd.n2723 vdd.n2722 185
R16909 vdd.n2721 vdd.n2720 185
R16910 vdd.n2719 vdd.n2718 185
R16911 vdd.n2717 vdd.n2716 185
R16912 vdd.n2715 vdd.n2714 185
R16913 vdd.n2713 vdd.n2712 185
R16914 vdd.n2710 vdd.n2709 185
R16915 vdd.n2708 vdd.n2707 185
R16916 vdd.n2706 vdd.n2705 185
R16917 vdd.n2913 vdd.n2912 185
R16918 vdd.n2914 vdd.n803 185
R16919 vdd.n2916 vdd.n2915 185
R16920 vdd.n2918 vdd.n801 185
R16921 vdd.n2920 vdd.n2919 185
R16922 vdd.n2921 vdd.n800 185
R16923 vdd.n2923 vdd.n2922 185
R16924 vdd.n2925 vdd.n798 185
R16925 vdd.n2927 vdd.n2926 185
R16926 vdd.n2928 vdd.n797 185
R16927 vdd.n2930 vdd.n2929 185
R16928 vdd.n2932 vdd.n795 185
R16929 vdd.n2934 vdd.n2933 185
R16930 vdd.n2935 vdd.n794 185
R16931 vdd.n2937 vdd.n2936 185
R16932 vdd.n2939 vdd.n792 185
R16933 vdd.n2941 vdd.n2940 185
R16934 vdd.n2943 vdd.n791 185
R16935 vdd.n2945 vdd.n2944 185
R16936 vdd.n2947 vdd.n789 185
R16937 vdd.n2949 vdd.n2948 185
R16938 vdd.n2950 vdd.n788 185
R16939 vdd.n2952 vdd.n2951 185
R16940 vdd.n2954 vdd.n786 185
R16941 vdd.n2956 vdd.n2955 185
R16942 vdd.n2957 vdd.n785 185
R16943 vdd.n2959 vdd.n2958 185
R16944 vdd.n2961 vdd.n783 185
R16945 vdd.n2963 vdd.n2962 185
R16946 vdd.n2964 vdd.n782 185
R16947 vdd.n2966 vdd.n2965 185
R16948 vdd.n2968 vdd.n781 185
R16949 vdd.n2969 vdd.n780 185
R16950 vdd.n2972 vdd.n2971 185
R16951 vdd.n2973 vdd.n778 185
R16952 vdd.n778 vdd.n756 185
R16953 vdd.n2910 vdd.n775 185
R16954 vdd.n2976 vdd.n775 185
R16955 vdd.n2909 vdd.n2908 185
R16956 vdd.n2908 vdd.n774 185
R16957 vdd.n2907 vdd.n807 185
R16958 vdd.n2907 vdd.n2906 185
R16959 vdd.n2661 vdd.n808 185
R16960 vdd.n817 vdd.n808 185
R16961 vdd.n2662 vdd.n815 185
R16962 vdd.n2900 vdd.n815 185
R16963 vdd.n2664 vdd.n2663 185
R16964 vdd.n2663 vdd.n814 185
R16965 vdd.n2665 vdd.n823 185
R16966 vdd.n2849 vdd.n823 185
R16967 vdd.n2667 vdd.n2666 185
R16968 vdd.n2666 vdd.n822 185
R16969 vdd.n2668 vdd.n829 185
R16970 vdd.n2843 vdd.n829 185
R16971 vdd.n2670 vdd.n2669 185
R16972 vdd.n2669 vdd.n828 185
R16973 vdd.n2671 vdd.n834 185
R16974 vdd.n2835 vdd.n834 185
R16975 vdd.n2673 vdd.n2672 185
R16976 vdd.n2672 vdd.n841 185
R16977 vdd.n2674 vdd.n839 185
R16978 vdd.n2829 vdd.n839 185
R16979 vdd.n2676 vdd.n2675 185
R16980 vdd.n2677 vdd.n2676 185
R16981 vdd.n2660 vdd.n846 185
R16982 vdd.n2823 vdd.n846 185
R16983 vdd.n2659 vdd.n2658 185
R16984 vdd.n2658 vdd.n845 185
R16985 vdd.n2657 vdd.n852 185
R16986 vdd.n2817 vdd.n852 185
R16987 vdd.n2656 vdd.n2655 185
R16988 vdd.n2655 vdd.n851 185
R16989 vdd.n2654 vdd.n857 185
R16990 vdd.n2811 vdd.n857 185
R16991 vdd.n2653 vdd.n2652 185
R16992 vdd.n2652 vdd.n864 185
R16993 vdd.n2651 vdd.n862 185
R16994 vdd.n2805 vdd.n862 185
R16995 vdd.n2650 vdd.n2649 185
R16996 vdd.n2649 vdd.n871 185
R16997 vdd.n2648 vdd.n869 185
R16998 vdd.n2799 vdd.n869 185
R16999 vdd.n2647 vdd.n2646 185
R17000 vdd.n2646 vdd.n868 185
R17001 vdd.n2558 vdd.n875 185
R17002 vdd.n2793 vdd.n875 185
R17003 vdd.n2700 vdd.n2699 185
R17004 vdd.n2699 vdd.n2698 185
R17005 vdd.n2701 vdd.n880 185
R17006 vdd.n2787 vdd.n880 185
R17007 vdd.n2703 vdd.n2702 185
R17008 vdd.n2702 vdd.t34 185
R17009 vdd.n2704 vdd.n885 185
R17010 vdd.n2781 vdd.n885 185
R17011 vdd.n2783 vdd.n2782 185
R17012 vdd.n2782 vdd.n2781 185
R17013 vdd.n2784 vdd.n882 185
R17014 vdd.n882 vdd.t34 185
R17015 vdd.n2786 vdd.n2785 185
R17016 vdd.n2787 vdd.n2786 185
R17017 vdd.n874 vdd.n873 185
R17018 vdd.n2698 vdd.n874 185
R17019 vdd.n2795 vdd.n2794 185
R17020 vdd.n2794 vdd.n2793 185
R17021 vdd.n2796 vdd.n872 185
R17022 vdd.n872 vdd.n868 185
R17023 vdd.n2798 vdd.n2797 185
R17024 vdd.n2799 vdd.n2798 185
R17025 vdd.n861 vdd.n860 185
R17026 vdd.n871 vdd.n861 185
R17027 vdd.n2807 vdd.n2806 185
R17028 vdd.n2806 vdd.n2805 185
R17029 vdd.n2808 vdd.n859 185
R17030 vdd.n864 vdd.n859 185
R17031 vdd.n2810 vdd.n2809 185
R17032 vdd.n2811 vdd.n2810 185
R17033 vdd.n850 vdd.n849 185
R17034 vdd.n851 vdd.n850 185
R17035 vdd.n2819 vdd.n2818 185
R17036 vdd.n2818 vdd.n2817 185
R17037 vdd.n2820 vdd.n848 185
R17038 vdd.n848 vdd.n845 185
R17039 vdd.n2822 vdd.n2821 185
R17040 vdd.n2823 vdd.n2822 185
R17041 vdd.n838 vdd.n837 185
R17042 vdd.n2677 vdd.n838 185
R17043 vdd.n2831 vdd.n2830 185
R17044 vdd.n2830 vdd.n2829 185
R17045 vdd.n2832 vdd.n836 185
R17046 vdd.n841 vdd.n836 185
R17047 vdd.n2834 vdd.n2833 185
R17048 vdd.n2835 vdd.n2834 185
R17049 vdd.n827 vdd.n826 185
R17050 vdd.n828 vdd.n827 185
R17051 vdd.n2845 vdd.n2844 185
R17052 vdd.n2844 vdd.n2843 185
R17053 vdd.n2846 vdd.n825 185
R17054 vdd.n825 vdd.n822 185
R17055 vdd.n2848 vdd.n2847 185
R17056 vdd.n2849 vdd.n2848 185
R17057 vdd.n813 vdd.n812 185
R17058 vdd.n814 vdd.n813 185
R17059 vdd.n2902 vdd.n2901 185
R17060 vdd.n2901 vdd.n2900 185
R17061 vdd.n2903 vdd.n811 185
R17062 vdd.n817 vdd.n811 185
R17063 vdd.n2905 vdd.n2904 185
R17064 vdd.n2906 vdd.n2905 185
R17065 vdd.n779 vdd.n777 185
R17066 vdd.n777 vdd.n774 185
R17067 vdd.n2975 vdd.n2974 185
R17068 vdd.n2976 vdd.n2975 185
R17069 vdd.n2448 vdd.n2447 185
R17070 vdd.n2449 vdd.n2448 185
R17071 vdd.n935 vdd.n933 185
R17072 vdd.n933 vdd.t8 185
R17073 vdd.n2363 vdd.n942 185
R17074 vdd.n2374 vdd.n942 185
R17075 vdd.n2364 vdd.n951 185
R17076 vdd.n2073 vdd.n951 185
R17077 vdd.n2366 vdd.n2365 185
R17078 vdd.n2367 vdd.n2366 185
R17079 vdd.n2362 vdd.n950 185
R17080 vdd.n950 vdd.n947 185
R17081 vdd.n2361 vdd.n2360 185
R17082 vdd.n2360 vdd.n2359 185
R17083 vdd.n953 vdd.n952 185
R17084 vdd.n954 vdd.n953 185
R17085 vdd.n2352 vdd.n2351 185
R17086 vdd.n2353 vdd.n2352 185
R17087 vdd.n2350 vdd.n963 185
R17088 vdd.n963 vdd.n960 185
R17089 vdd.n2349 vdd.n2348 185
R17090 vdd.n2348 vdd.n2347 185
R17091 vdd.n965 vdd.n964 185
R17092 vdd.n973 vdd.n965 185
R17093 vdd.n2340 vdd.n2339 185
R17094 vdd.n2341 vdd.n2340 185
R17095 vdd.n2338 vdd.n974 185
R17096 vdd.n979 vdd.n974 185
R17097 vdd.n2337 vdd.n2336 185
R17098 vdd.n2336 vdd.n2335 185
R17099 vdd.n976 vdd.n975 185
R17100 vdd.n2174 vdd.n976 185
R17101 vdd.n2328 vdd.n2327 185
R17102 vdd.n2329 vdd.n2328 185
R17103 vdd.n2326 vdd.n986 185
R17104 vdd.n986 vdd.n983 185
R17105 vdd.n2325 vdd.n2324 185
R17106 vdd.n2324 vdd.n2323 185
R17107 vdd.n988 vdd.n987 185
R17108 vdd.n989 vdd.n988 185
R17109 vdd.n2316 vdd.n2315 185
R17110 vdd.n2317 vdd.n2316 185
R17111 vdd.n2313 vdd.n997 185
R17112 vdd.n1004 vdd.n997 185
R17113 vdd.n2312 vdd.n2311 185
R17114 vdd.n2311 vdd.n2310 185
R17115 vdd.n1000 vdd.n999 185
R17116 vdd.n1001 vdd.n1000 185
R17117 vdd.n2303 vdd.n2302 185
R17118 vdd.n2304 vdd.n2303 185
R17119 vdd.n2301 vdd.n1011 185
R17120 vdd.n1011 vdd.n1008 185
R17121 vdd.n2300 vdd.n2299 185
R17122 vdd.n2299 vdd.n2298 185
R17123 vdd.n1013 vdd.n1012 185
R17124 vdd.n1014 vdd.n1013 185
R17125 vdd.n2291 vdd.n2290 185
R17126 vdd.n2292 vdd.n2291 185
R17127 vdd.n2379 vdd.n907 185
R17128 vdd.n2521 vdd.n907 185
R17129 vdd.n2381 vdd.n2380 185
R17130 vdd.n2383 vdd.n2382 185
R17131 vdd.n2385 vdd.n2384 185
R17132 vdd.n2387 vdd.n2386 185
R17133 vdd.n2389 vdd.n2388 185
R17134 vdd.n2391 vdd.n2390 185
R17135 vdd.n2393 vdd.n2392 185
R17136 vdd.n2395 vdd.n2394 185
R17137 vdd.n2397 vdd.n2396 185
R17138 vdd.n2399 vdd.n2398 185
R17139 vdd.n2401 vdd.n2400 185
R17140 vdd.n2403 vdd.n2402 185
R17141 vdd.n2405 vdd.n2404 185
R17142 vdd.n2407 vdd.n2406 185
R17143 vdd.n2409 vdd.n2408 185
R17144 vdd.n2411 vdd.n2410 185
R17145 vdd.n2413 vdd.n2412 185
R17146 vdd.n2415 vdd.n2414 185
R17147 vdd.n2417 vdd.n2416 185
R17148 vdd.n2419 vdd.n2418 185
R17149 vdd.n2421 vdd.n2420 185
R17150 vdd.n2423 vdd.n2422 185
R17151 vdd.n2425 vdd.n2424 185
R17152 vdd.n2427 vdd.n2426 185
R17153 vdd.n2429 vdd.n2428 185
R17154 vdd.n2431 vdd.n2430 185
R17155 vdd.n2433 vdd.n2432 185
R17156 vdd.n2435 vdd.n2434 185
R17157 vdd.n2437 vdd.n2436 185
R17158 vdd.n2439 vdd.n2438 185
R17159 vdd.n2441 vdd.n2440 185
R17160 vdd.n2443 vdd.n2442 185
R17161 vdd.n2445 vdd.n2444 185
R17162 vdd.n2446 vdd.n934 185
R17163 vdd.n2378 vdd.n932 185
R17164 vdd.n2449 vdd.n932 185
R17165 vdd.n2377 vdd.n2376 185
R17166 vdd.n2376 vdd.t8 185
R17167 vdd.n2375 vdd.n939 185
R17168 vdd.n2375 vdd.n2374 185
R17169 vdd.n2155 vdd.n940 185
R17170 vdd.n2073 vdd.n940 185
R17171 vdd.n2156 vdd.n949 185
R17172 vdd.n2367 vdd.n949 185
R17173 vdd.n2158 vdd.n2157 185
R17174 vdd.n2157 vdd.n947 185
R17175 vdd.n2159 vdd.n956 185
R17176 vdd.n2359 vdd.n956 185
R17177 vdd.n2161 vdd.n2160 185
R17178 vdd.n2160 vdd.n954 185
R17179 vdd.n2162 vdd.n962 185
R17180 vdd.n2353 vdd.n962 185
R17181 vdd.n2164 vdd.n2163 185
R17182 vdd.n2163 vdd.n960 185
R17183 vdd.n2165 vdd.n967 185
R17184 vdd.n2347 vdd.n967 185
R17185 vdd.n2167 vdd.n2166 185
R17186 vdd.n2166 vdd.n973 185
R17187 vdd.n2168 vdd.n972 185
R17188 vdd.n2341 vdd.n972 185
R17189 vdd.n2170 vdd.n2169 185
R17190 vdd.n2169 vdd.n979 185
R17191 vdd.n2171 vdd.n978 185
R17192 vdd.n2335 vdd.n978 185
R17193 vdd.n2173 vdd.n2172 185
R17194 vdd.n2174 vdd.n2173 185
R17195 vdd.n2154 vdd.n985 185
R17196 vdd.n2329 vdd.n985 185
R17197 vdd.n2153 vdd.n2152 185
R17198 vdd.n2152 vdd.n983 185
R17199 vdd.n2151 vdd.n991 185
R17200 vdd.n2323 vdd.n991 185
R17201 vdd.n2150 vdd.n2149 185
R17202 vdd.n2149 vdd.n989 185
R17203 vdd.n2148 vdd.n996 185
R17204 vdd.n2317 vdd.n996 185
R17205 vdd.n2147 vdd.n2146 185
R17206 vdd.n2146 vdd.n1004 185
R17207 vdd.n2145 vdd.n1003 185
R17208 vdd.n2310 vdd.n1003 185
R17209 vdd.n2144 vdd.n2143 185
R17210 vdd.n2143 vdd.n1001 185
R17211 vdd.n2142 vdd.n1010 185
R17212 vdd.n2304 vdd.n1010 185
R17213 vdd.n2141 vdd.n2140 185
R17214 vdd.n2140 vdd.n1008 185
R17215 vdd.n2139 vdd.n1016 185
R17216 vdd.n2298 vdd.n1016 185
R17217 vdd.n2138 vdd.n2137 185
R17218 vdd.n2137 vdd.n1014 185
R17219 vdd.n2136 vdd.n1022 185
R17220 vdd.n2292 vdd.n1022 185
R17221 vdd.n2289 vdd.n1023 185
R17222 vdd.n2288 vdd.n2287 185
R17223 vdd.n2285 vdd.n1024 185
R17224 vdd.n2283 vdd.n2282 185
R17225 vdd.n2281 vdd.n1025 185
R17226 vdd.n2280 vdd.n2279 185
R17227 vdd.n2277 vdd.n1026 185
R17228 vdd.n2275 vdd.n2274 185
R17229 vdd.n2273 vdd.n1027 185
R17230 vdd.n2272 vdd.n2271 185
R17231 vdd.n2269 vdd.n1028 185
R17232 vdd.n2267 vdd.n2266 185
R17233 vdd.n2265 vdd.n1029 185
R17234 vdd.n2264 vdd.n2263 185
R17235 vdd.n2261 vdd.n1030 185
R17236 vdd.n2259 vdd.n2258 185
R17237 vdd.n2257 vdd.n1031 185
R17238 vdd.n2256 vdd.n1033 185
R17239 vdd.n2101 vdd.n1034 185
R17240 vdd.n2104 vdd.n2103 185
R17241 vdd.n2106 vdd.n2105 185
R17242 vdd.n2108 vdd.n2100 185
R17243 vdd.n2111 vdd.n2110 185
R17244 vdd.n2112 vdd.n2099 185
R17245 vdd.n2114 vdd.n2113 185
R17246 vdd.n2116 vdd.n2098 185
R17247 vdd.n2119 vdd.n2118 185
R17248 vdd.n2120 vdd.n2097 185
R17249 vdd.n2122 vdd.n2121 185
R17250 vdd.n2124 vdd.n2096 185
R17251 vdd.n2127 vdd.n2126 185
R17252 vdd.n2128 vdd.n2093 185
R17253 vdd.n2131 vdd.n2130 185
R17254 vdd.n2133 vdd.n2092 185
R17255 vdd.n2135 vdd.n2134 185
R17256 vdd.n2134 vdd.n1020 185
R17257 vdd.n315 vdd.n314 171.744
R17258 vdd.n314 vdd.n313 171.744
R17259 vdd.n313 vdd.n282 171.744
R17260 vdd.n306 vdd.n282 171.744
R17261 vdd.n306 vdd.n305 171.744
R17262 vdd.n305 vdd.n287 171.744
R17263 vdd.n298 vdd.n287 171.744
R17264 vdd.n298 vdd.n297 171.744
R17265 vdd.n297 vdd.n291 171.744
R17266 vdd.n260 vdd.n259 171.744
R17267 vdd.n259 vdd.n258 171.744
R17268 vdd.n258 vdd.n227 171.744
R17269 vdd.n251 vdd.n227 171.744
R17270 vdd.n251 vdd.n250 171.744
R17271 vdd.n250 vdd.n232 171.744
R17272 vdd.n243 vdd.n232 171.744
R17273 vdd.n243 vdd.n242 171.744
R17274 vdd.n242 vdd.n236 171.744
R17275 vdd.n217 vdd.n216 171.744
R17276 vdd.n216 vdd.n215 171.744
R17277 vdd.n215 vdd.n184 171.744
R17278 vdd.n208 vdd.n184 171.744
R17279 vdd.n208 vdd.n207 171.744
R17280 vdd.n207 vdd.n189 171.744
R17281 vdd.n200 vdd.n189 171.744
R17282 vdd.n200 vdd.n199 171.744
R17283 vdd.n199 vdd.n193 171.744
R17284 vdd.n162 vdd.n161 171.744
R17285 vdd.n161 vdd.n160 171.744
R17286 vdd.n160 vdd.n129 171.744
R17287 vdd.n153 vdd.n129 171.744
R17288 vdd.n153 vdd.n152 171.744
R17289 vdd.n152 vdd.n134 171.744
R17290 vdd.n145 vdd.n134 171.744
R17291 vdd.n145 vdd.n144 171.744
R17292 vdd.n144 vdd.n138 171.744
R17293 vdd.n120 vdd.n119 171.744
R17294 vdd.n119 vdd.n118 171.744
R17295 vdd.n118 vdd.n87 171.744
R17296 vdd.n111 vdd.n87 171.744
R17297 vdd.n111 vdd.n110 171.744
R17298 vdd.n110 vdd.n92 171.744
R17299 vdd.n103 vdd.n92 171.744
R17300 vdd.n103 vdd.n102 171.744
R17301 vdd.n102 vdd.n96 171.744
R17302 vdd.n65 vdd.n64 171.744
R17303 vdd.n64 vdd.n63 171.744
R17304 vdd.n63 vdd.n32 171.744
R17305 vdd.n56 vdd.n32 171.744
R17306 vdd.n56 vdd.n55 171.744
R17307 vdd.n55 vdd.n37 171.744
R17308 vdd.n48 vdd.n37 171.744
R17309 vdd.n48 vdd.n47 171.744
R17310 vdd.n47 vdd.n41 171.744
R17311 vdd.n1684 vdd.n1683 171.744
R17312 vdd.n1683 vdd.n1682 171.744
R17313 vdd.n1682 vdd.n1651 171.744
R17314 vdd.n1675 vdd.n1651 171.744
R17315 vdd.n1675 vdd.n1674 171.744
R17316 vdd.n1674 vdd.n1656 171.744
R17317 vdd.n1667 vdd.n1656 171.744
R17318 vdd.n1667 vdd.n1666 171.744
R17319 vdd.n1666 vdd.n1660 171.744
R17320 vdd.n1739 vdd.n1738 171.744
R17321 vdd.n1738 vdd.n1737 171.744
R17322 vdd.n1737 vdd.n1706 171.744
R17323 vdd.n1730 vdd.n1706 171.744
R17324 vdd.n1730 vdd.n1729 171.744
R17325 vdd.n1729 vdd.n1711 171.744
R17326 vdd.n1722 vdd.n1711 171.744
R17327 vdd.n1722 vdd.n1721 171.744
R17328 vdd.n1721 vdd.n1715 171.744
R17329 vdd.n1586 vdd.n1585 171.744
R17330 vdd.n1585 vdd.n1584 171.744
R17331 vdd.n1584 vdd.n1553 171.744
R17332 vdd.n1577 vdd.n1553 171.744
R17333 vdd.n1577 vdd.n1576 171.744
R17334 vdd.n1576 vdd.n1558 171.744
R17335 vdd.n1569 vdd.n1558 171.744
R17336 vdd.n1569 vdd.n1568 171.744
R17337 vdd.n1568 vdd.n1562 171.744
R17338 vdd.n1641 vdd.n1640 171.744
R17339 vdd.n1640 vdd.n1639 171.744
R17340 vdd.n1639 vdd.n1608 171.744
R17341 vdd.n1632 vdd.n1608 171.744
R17342 vdd.n1632 vdd.n1631 171.744
R17343 vdd.n1631 vdd.n1613 171.744
R17344 vdd.n1624 vdd.n1613 171.744
R17345 vdd.n1624 vdd.n1623 171.744
R17346 vdd.n1623 vdd.n1617 171.744
R17347 vdd.n1489 vdd.n1488 171.744
R17348 vdd.n1488 vdd.n1487 171.744
R17349 vdd.n1487 vdd.n1456 171.744
R17350 vdd.n1480 vdd.n1456 171.744
R17351 vdd.n1480 vdd.n1479 171.744
R17352 vdd.n1479 vdd.n1461 171.744
R17353 vdd.n1472 vdd.n1461 171.744
R17354 vdd.n1472 vdd.n1471 171.744
R17355 vdd.n1471 vdd.n1465 171.744
R17356 vdd.n1544 vdd.n1543 171.744
R17357 vdd.n1543 vdd.n1542 171.744
R17358 vdd.n1542 vdd.n1511 171.744
R17359 vdd.n1535 vdd.n1511 171.744
R17360 vdd.n1535 vdd.n1534 171.744
R17361 vdd.n1534 vdd.n1516 171.744
R17362 vdd.n1527 vdd.n1516 171.744
R17363 vdd.n1527 vdd.n1526 171.744
R17364 vdd.n1526 vdd.n1520 171.744
R17365 vdd.n449 vdd.n448 146.341
R17366 vdd.n455 vdd.n454 146.341
R17367 vdd.n459 vdd.n458 146.341
R17368 vdd.n465 vdd.n464 146.341
R17369 vdd.n469 vdd.n468 146.341
R17370 vdd.n475 vdd.n474 146.341
R17371 vdd.n479 vdd.n478 146.341
R17372 vdd.n485 vdd.n484 146.341
R17373 vdd.n489 vdd.n488 146.341
R17374 vdd.n495 vdd.n494 146.341
R17375 vdd.n499 vdd.n498 146.341
R17376 vdd.n505 vdd.n504 146.341
R17377 vdd.n509 vdd.n508 146.341
R17378 vdd.n515 vdd.n514 146.341
R17379 vdd.n519 vdd.n518 146.341
R17380 vdd.n525 vdd.n524 146.341
R17381 vdd.n529 vdd.n528 146.341
R17382 vdd.n535 vdd.n534 146.341
R17383 vdd.n539 vdd.n538 146.341
R17384 vdd.n545 vdd.n544 146.341
R17385 vdd.n549 vdd.n548 146.341
R17386 vdd.n555 vdd.n554 146.341
R17387 vdd.n559 vdd.n558 146.341
R17388 vdd.n565 vdd.n564 146.341
R17389 vdd.n569 vdd.n568 146.341
R17390 vdd.n575 vdd.n574 146.341
R17391 vdd.n579 vdd.n578 146.341
R17392 vdd.n585 vdd.n584 146.341
R17393 vdd.n589 vdd.n588 146.341
R17394 vdd.n595 vdd.n594 146.341
R17395 vdd.n597 vdd.n404 146.341
R17396 vdd.n3146 vdd.n654 146.341
R17397 vdd.n3152 vdd.n654 146.341
R17398 vdd.n3152 vdd.n647 146.341
R17399 vdd.n3162 vdd.n647 146.341
R17400 vdd.n3162 vdd.n643 146.341
R17401 vdd.n3168 vdd.n643 146.341
R17402 vdd.n3168 vdd.n634 146.341
R17403 vdd.n3178 vdd.n634 146.341
R17404 vdd.n3178 vdd.n630 146.341
R17405 vdd.n3184 vdd.n630 146.341
R17406 vdd.n3184 vdd.n623 146.341
R17407 vdd.n3195 vdd.n623 146.341
R17408 vdd.n3195 vdd.n619 146.341
R17409 vdd.n3204 vdd.n619 146.341
R17410 vdd.n3204 vdd.n612 146.341
R17411 vdd.n3214 vdd.n612 146.341
R17412 vdd.n3215 vdd.n3214 146.341
R17413 vdd.n3215 vdd.n329 146.341
R17414 vdd.n330 vdd.n329 146.341
R17415 vdd.n331 vdd.n330 146.341
R17416 vdd.n3222 vdd.n331 146.341
R17417 vdd.n3222 vdd.n339 146.341
R17418 vdd.n340 vdd.n339 146.341
R17419 vdd.n341 vdd.n340 146.341
R17420 vdd.n3229 vdd.n341 146.341
R17421 vdd.n3229 vdd.n350 146.341
R17422 vdd.n351 vdd.n350 146.341
R17423 vdd.n352 vdd.n351 146.341
R17424 vdd.n3237 vdd.n352 146.341
R17425 vdd.n3237 vdd.n360 146.341
R17426 vdd.n361 vdd.n360 146.341
R17427 vdd.n362 vdd.n361 146.341
R17428 vdd.n3244 vdd.n362 146.341
R17429 vdd.n3244 vdd.n371 146.341
R17430 vdd.n372 vdd.n371 146.341
R17431 vdd.n3138 vdd.n3136 146.341
R17432 vdd.n3136 vdd.n3135 146.341
R17433 vdd.n3132 vdd.n3131 146.341
R17434 vdd.n3128 vdd.n3127 146.341
R17435 vdd.n3125 vdd.n669 146.341
R17436 vdd.n3121 vdd.n3119 146.341
R17437 vdd.n3117 vdd.n675 146.341
R17438 vdd.n3113 vdd.n3111 146.341
R17439 vdd.n3109 vdd.n681 146.341
R17440 vdd.n3105 vdd.n3103 146.341
R17441 vdd.n3101 vdd.n689 146.341
R17442 vdd.n3097 vdd.n3095 146.341
R17443 vdd.n3093 vdd.n695 146.341
R17444 vdd.n3089 vdd.n3087 146.341
R17445 vdd.n3085 vdd.n701 146.341
R17446 vdd.n3081 vdd.n3079 146.341
R17447 vdd.n3077 vdd.n707 146.341
R17448 vdd.n3073 vdd.n3071 146.341
R17449 vdd.n3069 vdd.n713 146.341
R17450 vdd.n3065 vdd.n3063 146.341
R17451 vdd.n3061 vdd.n719 146.341
R17452 vdd.n3054 vdd.n728 146.341
R17453 vdd.n3052 vdd.n3051 146.341
R17454 vdd.n3048 vdd.n3047 146.341
R17455 vdd.n3045 vdd.n733 146.341
R17456 vdd.n3041 vdd.n3039 146.341
R17457 vdd.n3037 vdd.n739 146.341
R17458 vdd.n3033 vdd.n3031 146.341
R17459 vdd.n3029 vdd.n745 146.341
R17460 vdd.n3025 vdd.n3023 146.341
R17461 vdd.n3020 vdd.n3019 146.341
R17462 vdd.n3016 vdd.n657 146.341
R17463 vdd.n3144 vdd.n653 146.341
R17464 vdd.n3154 vdd.n653 146.341
R17465 vdd.n3154 vdd.n649 146.341
R17466 vdd.n3160 vdd.n649 146.341
R17467 vdd.n3160 vdd.n641 146.341
R17468 vdd.n3170 vdd.n641 146.341
R17469 vdd.n3170 vdd.n637 146.341
R17470 vdd.n3176 vdd.n637 146.341
R17471 vdd.n3176 vdd.n629 146.341
R17472 vdd.n3187 vdd.n629 146.341
R17473 vdd.n3187 vdd.n625 146.341
R17474 vdd.n3193 vdd.n625 146.341
R17475 vdd.n3193 vdd.n618 146.341
R17476 vdd.n3206 vdd.n618 146.341
R17477 vdd.n3206 vdd.n614 146.341
R17478 vdd.n3212 vdd.n614 146.341
R17479 vdd.n3212 vdd.n326 146.341
R17480 vdd.n3288 vdd.n326 146.341
R17481 vdd.n3288 vdd.n327 146.341
R17482 vdd.n3284 vdd.n327 146.341
R17483 vdd.n3284 vdd.n333 146.341
R17484 vdd.n3280 vdd.n333 146.341
R17485 vdd.n3280 vdd.n338 146.341
R17486 vdd.n3276 vdd.n338 146.341
R17487 vdd.n3276 vdd.n342 146.341
R17488 vdd.n3272 vdd.n342 146.341
R17489 vdd.n3272 vdd.n348 146.341
R17490 vdd.n3268 vdd.n348 146.341
R17491 vdd.n3268 vdd.n353 146.341
R17492 vdd.n3264 vdd.n353 146.341
R17493 vdd.n3264 vdd.n359 146.341
R17494 vdd.n3260 vdd.n359 146.341
R17495 vdd.n3260 vdd.n364 146.341
R17496 vdd.n3256 vdd.n364 146.341
R17497 vdd.n3256 vdd.n370 146.341
R17498 vdd.n2239 vdd.n2238 146.341
R17499 vdd.n2236 vdd.n1820 146.341
R17500 vdd.n2016 vdd.n1826 146.341
R17501 vdd.n2014 vdd.n2013 146.341
R17502 vdd.n2011 vdd.n1828 146.341
R17503 vdd.n2007 vdd.n2006 146.341
R17504 vdd.n2004 vdd.n1835 146.341
R17505 vdd.n2000 vdd.n1999 146.341
R17506 vdd.n1997 vdd.n1842 146.341
R17507 vdd.n1853 vdd.n1850 146.341
R17508 vdd.n1989 vdd.n1988 146.341
R17509 vdd.n1986 vdd.n1855 146.341
R17510 vdd.n1982 vdd.n1981 146.341
R17511 vdd.n1979 vdd.n1861 146.341
R17512 vdd.n1975 vdd.n1974 146.341
R17513 vdd.n1972 vdd.n1868 146.341
R17514 vdd.n1968 vdd.n1967 146.341
R17515 vdd.n1965 vdd.n1875 146.341
R17516 vdd.n1961 vdd.n1960 146.341
R17517 vdd.n1958 vdd.n1882 146.341
R17518 vdd.n1893 vdd.n1890 146.341
R17519 vdd.n1950 vdd.n1949 146.341
R17520 vdd.n1947 vdd.n1895 146.341
R17521 vdd.n1943 vdd.n1942 146.341
R17522 vdd.n1940 vdd.n1901 146.341
R17523 vdd.n1936 vdd.n1935 146.341
R17524 vdd.n1933 vdd.n1908 146.341
R17525 vdd.n1929 vdd.n1928 146.341
R17526 vdd.n1926 vdd.n1923 146.341
R17527 vdd.n1921 vdd.n1918 146.341
R17528 vdd.n1916 vdd.n1040 146.341
R17529 vdd.n1381 vdd.n1145 146.341
R17530 vdd.n1381 vdd.n1137 146.341
R17531 vdd.n1391 vdd.n1137 146.341
R17532 vdd.n1391 vdd.n1133 146.341
R17533 vdd.n1397 vdd.n1133 146.341
R17534 vdd.n1397 vdd.n1125 146.341
R17535 vdd.n1408 vdd.n1125 146.341
R17536 vdd.n1408 vdd.n1121 146.341
R17537 vdd.n1414 vdd.n1121 146.341
R17538 vdd.n1414 vdd.n1115 146.341
R17539 vdd.n1425 vdd.n1115 146.341
R17540 vdd.n1425 vdd.n1111 146.341
R17541 vdd.n1431 vdd.n1111 146.341
R17542 vdd.n1431 vdd.n1102 146.341
R17543 vdd.n1441 vdd.n1102 146.341
R17544 vdd.n1441 vdd.n1098 146.341
R17545 vdd.n1447 vdd.n1098 146.341
R17546 vdd.n1447 vdd.n1091 146.341
R17547 vdd.n1753 vdd.n1091 146.341
R17548 vdd.n1753 vdd.n1087 146.341
R17549 vdd.n1759 vdd.n1087 146.341
R17550 vdd.n1759 vdd.n1080 146.341
R17551 vdd.n1769 vdd.n1080 146.341
R17552 vdd.n1769 vdd.n1076 146.341
R17553 vdd.n1775 vdd.n1076 146.341
R17554 vdd.n1775 vdd.n1068 146.341
R17555 vdd.n1786 vdd.n1068 146.341
R17556 vdd.n1786 vdd.n1064 146.341
R17557 vdd.n1792 vdd.n1064 146.341
R17558 vdd.n1792 vdd.n1058 146.341
R17559 vdd.n1803 vdd.n1058 146.341
R17560 vdd.n1803 vdd.n1053 146.341
R17561 vdd.n1811 vdd.n1053 146.341
R17562 vdd.n1811 vdd.n1042 146.341
R17563 vdd.n2247 vdd.n1042 146.341
R17564 vdd.n1183 vdd.n1182 146.341
R17565 vdd.n1187 vdd.n1182 146.341
R17566 vdd.n1189 vdd.n1188 146.341
R17567 vdd.n1193 vdd.n1192 146.341
R17568 vdd.n1195 vdd.n1194 146.341
R17569 vdd.n1199 vdd.n1198 146.341
R17570 vdd.n1201 vdd.n1200 146.341
R17571 vdd.n1205 vdd.n1204 146.341
R17572 vdd.n1207 vdd.n1206 146.341
R17573 vdd.n1339 vdd.n1338 146.341
R17574 vdd.n1211 vdd.n1210 146.341
R17575 vdd.n1215 vdd.n1214 146.341
R17576 vdd.n1217 vdd.n1216 146.341
R17577 vdd.n1221 vdd.n1220 146.341
R17578 vdd.n1223 vdd.n1222 146.341
R17579 vdd.n1227 vdd.n1226 146.341
R17580 vdd.n1229 vdd.n1228 146.341
R17581 vdd.n1233 vdd.n1232 146.341
R17582 vdd.n1235 vdd.n1234 146.341
R17583 vdd.n1239 vdd.n1238 146.341
R17584 vdd.n1303 vdd.n1240 146.341
R17585 vdd.n1244 vdd.n1243 146.341
R17586 vdd.n1246 vdd.n1245 146.341
R17587 vdd.n1250 vdd.n1249 146.341
R17588 vdd.n1252 vdd.n1251 146.341
R17589 vdd.n1256 vdd.n1255 146.341
R17590 vdd.n1258 vdd.n1257 146.341
R17591 vdd.n1262 vdd.n1261 146.341
R17592 vdd.n1264 vdd.n1263 146.341
R17593 vdd.n1268 vdd.n1267 146.341
R17594 vdd.n1270 vdd.n1269 146.341
R17595 vdd.n1375 vdd.n1151 146.341
R17596 vdd.n1383 vdd.n1143 146.341
R17597 vdd.n1383 vdd.n1139 146.341
R17598 vdd.n1389 vdd.n1139 146.341
R17599 vdd.n1389 vdd.n1131 146.341
R17600 vdd.n1400 vdd.n1131 146.341
R17601 vdd.n1400 vdd.n1127 146.341
R17602 vdd.n1406 vdd.n1127 146.341
R17603 vdd.n1406 vdd.n1120 146.341
R17604 vdd.n1417 vdd.n1120 146.341
R17605 vdd.n1417 vdd.n1116 146.341
R17606 vdd.n1423 vdd.n1116 146.341
R17607 vdd.n1423 vdd.n1109 146.341
R17608 vdd.n1433 vdd.n1109 146.341
R17609 vdd.n1433 vdd.n1105 146.341
R17610 vdd.n1439 vdd.n1105 146.341
R17611 vdd.n1439 vdd.n1097 146.341
R17612 vdd.n1450 vdd.n1097 146.341
R17613 vdd.n1450 vdd.n1093 146.341
R17614 vdd.n1751 vdd.n1093 146.341
R17615 vdd.n1751 vdd.n1086 146.341
R17616 vdd.n1761 vdd.n1086 146.341
R17617 vdd.n1761 vdd.n1082 146.341
R17618 vdd.n1767 vdd.n1082 146.341
R17619 vdd.n1767 vdd.n1074 146.341
R17620 vdd.n1778 vdd.n1074 146.341
R17621 vdd.n1778 vdd.n1070 146.341
R17622 vdd.n1784 vdd.n1070 146.341
R17623 vdd.n1784 vdd.n1063 146.341
R17624 vdd.n1795 vdd.n1063 146.341
R17625 vdd.n1795 vdd.n1059 146.341
R17626 vdd.n1801 vdd.n1059 146.341
R17627 vdd.n1801 vdd.n1051 146.341
R17628 vdd.n1813 vdd.n1051 146.341
R17629 vdd.n1813 vdd.n1046 146.341
R17630 vdd.n2245 vdd.n1046 146.341
R17631 vdd.n1045 vdd.n1020 141.707
R17632 vdd.n756 vdd.n658 141.707
R17633 vdd.n2094 vdd.t228 127.284
R17634 vdd.n936 vdd.t213 127.284
R17635 vdd.n2068 vdd.t175 127.284
R17636 vdd.n928 vdd.t237 127.284
R17637 vdd.n2839 vdd.t200 127.284
R17638 vdd.n2839 vdd.t201 127.284
R17639 vdd.n2559 vdd.t235 127.284
R17640 vdd.n804 vdd.t217 127.284
R17641 vdd.n2556 vdd.t222 127.284
R17642 vdd.n768 vdd.t224 127.284
R17643 vdd.n998 vdd.t231 127.284
R17644 vdd.n998 vdd.t232 127.284
R17645 vdd.n22 vdd.n20 117.314
R17646 vdd.n17 vdd.n15 117.314
R17647 vdd.n27 vdd.n26 116.927
R17648 vdd.n24 vdd.n23 116.927
R17649 vdd.n22 vdd.n21 116.927
R17650 vdd.n17 vdd.n16 116.927
R17651 vdd.n19 vdd.n18 116.927
R17652 vdd.n27 vdd.n25 116.927
R17653 vdd.n2095 vdd.t227 111.188
R17654 vdd.n937 vdd.t214 111.188
R17655 vdd.n2069 vdd.t174 111.188
R17656 vdd.n929 vdd.t238 111.188
R17657 vdd.n2560 vdd.t234 111.188
R17658 vdd.n805 vdd.t218 111.188
R17659 vdd.n2557 vdd.t221 111.188
R17660 vdd.n769 vdd.t225 111.188
R17661 vdd.n2782 vdd.n882 99.5127
R17662 vdd.n2786 vdd.n882 99.5127
R17663 vdd.n2786 vdd.n874 99.5127
R17664 vdd.n2794 vdd.n874 99.5127
R17665 vdd.n2794 vdd.n872 99.5127
R17666 vdd.n2798 vdd.n872 99.5127
R17667 vdd.n2798 vdd.n861 99.5127
R17668 vdd.n2806 vdd.n861 99.5127
R17669 vdd.n2806 vdd.n859 99.5127
R17670 vdd.n2810 vdd.n859 99.5127
R17671 vdd.n2810 vdd.n850 99.5127
R17672 vdd.n2818 vdd.n850 99.5127
R17673 vdd.n2818 vdd.n848 99.5127
R17674 vdd.n2822 vdd.n848 99.5127
R17675 vdd.n2822 vdd.n838 99.5127
R17676 vdd.n2830 vdd.n838 99.5127
R17677 vdd.n2830 vdd.n836 99.5127
R17678 vdd.n2834 vdd.n836 99.5127
R17679 vdd.n2834 vdd.n827 99.5127
R17680 vdd.n2844 vdd.n827 99.5127
R17681 vdd.n2844 vdd.n825 99.5127
R17682 vdd.n2848 vdd.n825 99.5127
R17683 vdd.n2848 vdd.n813 99.5127
R17684 vdd.n2901 vdd.n813 99.5127
R17685 vdd.n2901 vdd.n811 99.5127
R17686 vdd.n2905 vdd.n811 99.5127
R17687 vdd.n2905 vdd.n777 99.5127
R17688 vdd.n2975 vdd.n777 99.5127
R17689 vdd.n2971 vdd.n778 99.5127
R17690 vdd.n2969 vdd.n2968 99.5127
R17691 vdd.n2966 vdd.n782 99.5127
R17692 vdd.n2962 vdd.n2961 99.5127
R17693 vdd.n2959 vdd.n785 99.5127
R17694 vdd.n2955 vdd.n2954 99.5127
R17695 vdd.n2952 vdd.n788 99.5127
R17696 vdd.n2948 vdd.n2947 99.5127
R17697 vdd.n2945 vdd.n791 99.5127
R17698 vdd.n2940 vdd.n2939 99.5127
R17699 vdd.n2937 vdd.n794 99.5127
R17700 vdd.n2933 vdd.n2932 99.5127
R17701 vdd.n2930 vdd.n797 99.5127
R17702 vdd.n2926 vdd.n2925 99.5127
R17703 vdd.n2923 vdd.n800 99.5127
R17704 vdd.n2919 vdd.n2918 99.5127
R17705 vdd.n2916 vdd.n803 99.5127
R17706 vdd.n2702 vdd.n885 99.5127
R17707 vdd.n2702 vdd.n880 99.5127
R17708 vdd.n2699 vdd.n880 99.5127
R17709 vdd.n2699 vdd.n875 99.5127
R17710 vdd.n2646 vdd.n875 99.5127
R17711 vdd.n2646 vdd.n869 99.5127
R17712 vdd.n2649 vdd.n869 99.5127
R17713 vdd.n2649 vdd.n862 99.5127
R17714 vdd.n2652 vdd.n862 99.5127
R17715 vdd.n2652 vdd.n857 99.5127
R17716 vdd.n2655 vdd.n857 99.5127
R17717 vdd.n2655 vdd.n852 99.5127
R17718 vdd.n2658 vdd.n852 99.5127
R17719 vdd.n2658 vdd.n846 99.5127
R17720 vdd.n2676 vdd.n846 99.5127
R17721 vdd.n2676 vdd.n839 99.5127
R17722 vdd.n2672 vdd.n839 99.5127
R17723 vdd.n2672 vdd.n834 99.5127
R17724 vdd.n2669 vdd.n834 99.5127
R17725 vdd.n2669 vdd.n829 99.5127
R17726 vdd.n2666 vdd.n829 99.5127
R17727 vdd.n2666 vdd.n823 99.5127
R17728 vdd.n2663 vdd.n823 99.5127
R17729 vdd.n2663 vdd.n815 99.5127
R17730 vdd.n815 vdd.n808 99.5127
R17731 vdd.n2907 vdd.n808 99.5127
R17732 vdd.n2908 vdd.n2907 99.5127
R17733 vdd.n2908 vdd.n775 99.5127
R17734 vdd.n2772 vdd.n2555 99.5127
R17735 vdd.n2768 vdd.n2555 99.5127
R17736 vdd.n2766 vdd.n2765 99.5127
R17737 vdd.n2762 vdd.n2761 99.5127
R17738 vdd.n2758 vdd.n2757 99.5127
R17739 vdd.n2754 vdd.n2753 99.5127
R17740 vdd.n2750 vdd.n2749 99.5127
R17741 vdd.n2746 vdd.n2745 99.5127
R17742 vdd.n2742 vdd.n2741 99.5127
R17743 vdd.n2738 vdd.n2737 99.5127
R17744 vdd.n2734 vdd.n2733 99.5127
R17745 vdd.n2730 vdd.n2729 99.5127
R17746 vdd.n2726 vdd.n2725 99.5127
R17747 vdd.n2722 vdd.n2721 99.5127
R17748 vdd.n2718 vdd.n2717 99.5127
R17749 vdd.n2714 vdd.n2713 99.5127
R17750 vdd.n2709 vdd.n2708 99.5127
R17751 vdd.n2520 vdd.n926 99.5127
R17752 vdd.n2516 vdd.n2515 99.5127
R17753 vdd.n2512 vdd.n2511 99.5127
R17754 vdd.n2508 vdd.n2507 99.5127
R17755 vdd.n2504 vdd.n2503 99.5127
R17756 vdd.n2500 vdd.n2499 99.5127
R17757 vdd.n2496 vdd.n2495 99.5127
R17758 vdd.n2492 vdd.n2491 99.5127
R17759 vdd.n2488 vdd.n2487 99.5127
R17760 vdd.n2484 vdd.n2483 99.5127
R17761 vdd.n2480 vdd.n2479 99.5127
R17762 vdd.n2476 vdd.n2475 99.5127
R17763 vdd.n2472 vdd.n2471 99.5127
R17764 vdd.n2468 vdd.n2467 99.5127
R17765 vdd.n2464 vdd.n2463 99.5127
R17766 vdd.n2460 vdd.n2459 99.5127
R17767 vdd.n2455 vdd.n2454 99.5127
R17768 vdd.n2193 vdd.n1021 99.5127
R17769 vdd.n2193 vdd.n1015 99.5127
R17770 vdd.n2190 vdd.n1015 99.5127
R17771 vdd.n2190 vdd.n1009 99.5127
R17772 vdd.n2187 vdd.n1009 99.5127
R17773 vdd.n2187 vdd.n1002 99.5127
R17774 vdd.n2184 vdd.n1002 99.5127
R17775 vdd.n2184 vdd.n995 99.5127
R17776 vdd.n2181 vdd.n995 99.5127
R17777 vdd.n2181 vdd.n990 99.5127
R17778 vdd.n2178 vdd.n990 99.5127
R17779 vdd.n2178 vdd.n984 99.5127
R17780 vdd.n2175 vdd.n984 99.5127
R17781 vdd.n2175 vdd.n977 99.5127
R17782 vdd.n2089 vdd.n977 99.5127
R17783 vdd.n2089 vdd.n971 99.5127
R17784 vdd.n2086 vdd.n971 99.5127
R17785 vdd.n2086 vdd.n966 99.5127
R17786 vdd.n2083 vdd.n966 99.5127
R17787 vdd.n2083 vdd.n961 99.5127
R17788 vdd.n2080 vdd.n961 99.5127
R17789 vdd.n2080 vdd.n955 99.5127
R17790 vdd.n2077 vdd.n955 99.5127
R17791 vdd.n2077 vdd.n948 99.5127
R17792 vdd.n2074 vdd.n948 99.5127
R17793 vdd.n2074 vdd.n941 99.5127
R17794 vdd.n941 vdd.n931 99.5127
R17795 vdd.n2450 vdd.n931 99.5127
R17796 vdd.n2028 vdd.n2026 99.5127
R17797 vdd.n2032 vdd.n2026 99.5127
R17798 vdd.n2036 vdd.n2034 99.5127
R17799 vdd.n2040 vdd.n2024 99.5127
R17800 vdd.n2044 vdd.n2042 99.5127
R17801 vdd.n2048 vdd.n2022 99.5127
R17802 vdd.n2052 vdd.n2050 99.5127
R17803 vdd.n2056 vdd.n2020 99.5127
R17804 vdd.n2059 vdd.n2058 99.5127
R17805 vdd.n2229 vdd.n2227 99.5127
R17806 vdd.n2225 vdd.n2061 99.5127
R17807 vdd.n2221 vdd.n2219 99.5127
R17808 vdd.n2217 vdd.n2063 99.5127
R17809 vdd.n2213 vdd.n2211 99.5127
R17810 vdd.n2209 vdd.n2065 99.5127
R17811 vdd.n2205 vdd.n2203 99.5127
R17812 vdd.n2201 vdd.n2067 99.5127
R17813 vdd.n2293 vdd.n1017 99.5127
R17814 vdd.n2297 vdd.n1017 99.5127
R17815 vdd.n2297 vdd.n1007 99.5127
R17816 vdd.n2305 vdd.n1007 99.5127
R17817 vdd.n2305 vdd.n1005 99.5127
R17818 vdd.n2309 vdd.n1005 99.5127
R17819 vdd.n2309 vdd.n994 99.5127
R17820 vdd.n2318 vdd.n994 99.5127
R17821 vdd.n2318 vdd.n992 99.5127
R17822 vdd.n2322 vdd.n992 99.5127
R17823 vdd.n2322 vdd.n982 99.5127
R17824 vdd.n2330 vdd.n982 99.5127
R17825 vdd.n2330 vdd.n980 99.5127
R17826 vdd.n2334 vdd.n980 99.5127
R17827 vdd.n2334 vdd.n970 99.5127
R17828 vdd.n2342 vdd.n970 99.5127
R17829 vdd.n2342 vdd.n968 99.5127
R17830 vdd.n2346 vdd.n968 99.5127
R17831 vdd.n2346 vdd.n959 99.5127
R17832 vdd.n2354 vdd.n959 99.5127
R17833 vdd.n2354 vdd.n957 99.5127
R17834 vdd.n2358 vdd.n957 99.5127
R17835 vdd.n2358 vdd.n946 99.5127
R17836 vdd.n2368 vdd.n946 99.5127
R17837 vdd.n2368 vdd.n943 99.5127
R17838 vdd.n2373 vdd.n943 99.5127
R17839 vdd.n2373 vdd.n944 99.5127
R17840 vdd.n944 vdd.n925 99.5127
R17841 vdd.n2891 vdd.n2890 99.5127
R17842 vdd.n2888 vdd.n2854 99.5127
R17843 vdd.n2884 vdd.n2883 99.5127
R17844 vdd.n2881 vdd.n2857 99.5127
R17845 vdd.n2877 vdd.n2876 99.5127
R17846 vdd.n2874 vdd.n2860 99.5127
R17847 vdd.n2870 vdd.n2869 99.5127
R17848 vdd.n2867 vdd.n2864 99.5127
R17849 vdd.n3008 vdd.n755 99.5127
R17850 vdd.n3006 vdd.n3005 99.5127
R17851 vdd.n3003 vdd.n758 99.5127
R17852 vdd.n2999 vdd.n2998 99.5127
R17853 vdd.n2996 vdd.n761 99.5127
R17854 vdd.n2992 vdd.n2991 99.5127
R17855 vdd.n2989 vdd.n764 99.5127
R17856 vdd.n2985 vdd.n2984 99.5127
R17857 vdd.n2982 vdd.n767 99.5127
R17858 vdd.n2626 vdd.n886 99.5127
R17859 vdd.n2626 vdd.n881 99.5127
R17860 vdd.n2697 vdd.n881 99.5127
R17861 vdd.n2697 vdd.n876 99.5127
R17862 vdd.n2693 vdd.n876 99.5127
R17863 vdd.n2693 vdd.n870 99.5127
R17864 vdd.n2690 vdd.n870 99.5127
R17865 vdd.n2690 vdd.n863 99.5127
R17866 vdd.n2687 vdd.n863 99.5127
R17867 vdd.n2687 vdd.n858 99.5127
R17868 vdd.n2684 vdd.n858 99.5127
R17869 vdd.n2684 vdd.n853 99.5127
R17870 vdd.n2681 vdd.n853 99.5127
R17871 vdd.n2681 vdd.n847 99.5127
R17872 vdd.n2678 vdd.n847 99.5127
R17873 vdd.n2678 vdd.n840 99.5127
R17874 vdd.n2643 vdd.n840 99.5127
R17875 vdd.n2643 vdd.n835 99.5127
R17876 vdd.n2640 vdd.n835 99.5127
R17877 vdd.n2640 vdd.n830 99.5127
R17878 vdd.n2637 vdd.n830 99.5127
R17879 vdd.n2637 vdd.n824 99.5127
R17880 vdd.n2634 vdd.n824 99.5127
R17881 vdd.n2634 vdd.n816 99.5127
R17882 vdd.n2631 vdd.n816 99.5127
R17883 vdd.n2631 vdd.n809 99.5127
R17884 vdd.n809 vdd.n773 99.5127
R17885 vdd.n2977 vdd.n773 99.5127
R17886 vdd.n2776 vdd.n889 99.5127
R17887 vdd.n2564 vdd.n2563 99.5127
R17888 vdd.n2568 vdd.n2567 99.5127
R17889 vdd.n2572 vdd.n2571 99.5127
R17890 vdd.n2576 vdd.n2575 99.5127
R17891 vdd.n2580 vdd.n2579 99.5127
R17892 vdd.n2584 vdd.n2583 99.5127
R17893 vdd.n2588 vdd.n2587 99.5127
R17894 vdd.n2592 vdd.n2591 99.5127
R17895 vdd.n2596 vdd.n2595 99.5127
R17896 vdd.n2600 vdd.n2599 99.5127
R17897 vdd.n2604 vdd.n2603 99.5127
R17898 vdd.n2608 vdd.n2607 99.5127
R17899 vdd.n2612 vdd.n2611 99.5127
R17900 vdd.n2616 vdd.n2615 99.5127
R17901 vdd.n2620 vdd.n2619 99.5127
R17902 vdd.n2622 vdd.n2554 99.5127
R17903 vdd.n2780 vdd.n879 99.5127
R17904 vdd.n2788 vdd.n879 99.5127
R17905 vdd.n2788 vdd.n877 99.5127
R17906 vdd.n2792 vdd.n877 99.5127
R17907 vdd.n2792 vdd.n867 99.5127
R17908 vdd.n2800 vdd.n867 99.5127
R17909 vdd.n2800 vdd.n865 99.5127
R17910 vdd.n2804 vdd.n865 99.5127
R17911 vdd.n2804 vdd.n856 99.5127
R17912 vdd.n2812 vdd.n856 99.5127
R17913 vdd.n2812 vdd.n854 99.5127
R17914 vdd.n2816 vdd.n854 99.5127
R17915 vdd.n2816 vdd.n844 99.5127
R17916 vdd.n2824 vdd.n844 99.5127
R17917 vdd.n2824 vdd.n842 99.5127
R17918 vdd.n2828 vdd.n842 99.5127
R17919 vdd.n2828 vdd.n833 99.5127
R17920 vdd.n2836 vdd.n833 99.5127
R17921 vdd.n2836 vdd.n831 99.5127
R17922 vdd.n2842 vdd.n831 99.5127
R17923 vdd.n2842 vdd.n821 99.5127
R17924 vdd.n2850 vdd.n821 99.5127
R17925 vdd.n2850 vdd.n818 99.5127
R17926 vdd.n2899 vdd.n818 99.5127
R17927 vdd.n2899 vdd.n819 99.5127
R17928 vdd.n819 vdd.n810 99.5127
R17929 vdd.n2894 vdd.n810 99.5127
R17930 vdd.n2894 vdd.n776 99.5127
R17931 vdd.n2444 vdd.n2443 99.5127
R17932 vdd.n2440 vdd.n2439 99.5127
R17933 vdd.n2436 vdd.n2435 99.5127
R17934 vdd.n2432 vdd.n2431 99.5127
R17935 vdd.n2428 vdd.n2427 99.5127
R17936 vdd.n2424 vdd.n2423 99.5127
R17937 vdd.n2420 vdd.n2419 99.5127
R17938 vdd.n2416 vdd.n2415 99.5127
R17939 vdd.n2412 vdd.n2411 99.5127
R17940 vdd.n2408 vdd.n2407 99.5127
R17941 vdd.n2404 vdd.n2403 99.5127
R17942 vdd.n2400 vdd.n2399 99.5127
R17943 vdd.n2396 vdd.n2395 99.5127
R17944 vdd.n2392 vdd.n2391 99.5127
R17945 vdd.n2388 vdd.n2387 99.5127
R17946 vdd.n2384 vdd.n2383 99.5127
R17947 vdd.n2380 vdd.n907 99.5127
R17948 vdd.n2137 vdd.n1022 99.5127
R17949 vdd.n2137 vdd.n1016 99.5127
R17950 vdd.n2140 vdd.n1016 99.5127
R17951 vdd.n2140 vdd.n1010 99.5127
R17952 vdd.n2143 vdd.n1010 99.5127
R17953 vdd.n2143 vdd.n1003 99.5127
R17954 vdd.n2146 vdd.n1003 99.5127
R17955 vdd.n2146 vdd.n996 99.5127
R17956 vdd.n2149 vdd.n996 99.5127
R17957 vdd.n2149 vdd.n991 99.5127
R17958 vdd.n2152 vdd.n991 99.5127
R17959 vdd.n2152 vdd.n985 99.5127
R17960 vdd.n2173 vdd.n985 99.5127
R17961 vdd.n2173 vdd.n978 99.5127
R17962 vdd.n2169 vdd.n978 99.5127
R17963 vdd.n2169 vdd.n972 99.5127
R17964 vdd.n2166 vdd.n972 99.5127
R17965 vdd.n2166 vdd.n967 99.5127
R17966 vdd.n2163 vdd.n967 99.5127
R17967 vdd.n2163 vdd.n962 99.5127
R17968 vdd.n2160 vdd.n962 99.5127
R17969 vdd.n2160 vdd.n956 99.5127
R17970 vdd.n2157 vdd.n956 99.5127
R17971 vdd.n2157 vdd.n949 99.5127
R17972 vdd.n949 vdd.n940 99.5127
R17973 vdd.n2375 vdd.n940 99.5127
R17974 vdd.n2376 vdd.n2375 99.5127
R17975 vdd.n2376 vdd.n932 99.5127
R17976 vdd.n2287 vdd.n2285 99.5127
R17977 vdd.n2283 vdd.n1025 99.5127
R17978 vdd.n2279 vdd.n2277 99.5127
R17979 vdd.n2275 vdd.n1027 99.5127
R17980 vdd.n2271 vdd.n2269 99.5127
R17981 vdd.n2267 vdd.n1029 99.5127
R17982 vdd.n2263 vdd.n2261 99.5127
R17983 vdd.n2259 vdd.n1031 99.5127
R17984 vdd.n2101 vdd.n1033 99.5127
R17985 vdd.n2106 vdd.n2103 99.5127
R17986 vdd.n2110 vdd.n2108 99.5127
R17987 vdd.n2114 vdd.n2099 99.5127
R17988 vdd.n2118 vdd.n2116 99.5127
R17989 vdd.n2122 vdd.n2097 99.5127
R17990 vdd.n2126 vdd.n2124 99.5127
R17991 vdd.n2131 vdd.n2093 99.5127
R17992 vdd.n2134 vdd.n2133 99.5127
R17993 vdd.n2291 vdd.n1013 99.5127
R17994 vdd.n2299 vdd.n1013 99.5127
R17995 vdd.n2299 vdd.n1011 99.5127
R17996 vdd.n2303 vdd.n1011 99.5127
R17997 vdd.n2303 vdd.n1000 99.5127
R17998 vdd.n2311 vdd.n1000 99.5127
R17999 vdd.n2311 vdd.n997 99.5127
R18000 vdd.n2316 vdd.n997 99.5127
R18001 vdd.n2316 vdd.n988 99.5127
R18002 vdd.n2324 vdd.n988 99.5127
R18003 vdd.n2324 vdd.n986 99.5127
R18004 vdd.n2328 vdd.n986 99.5127
R18005 vdd.n2328 vdd.n976 99.5127
R18006 vdd.n2336 vdd.n976 99.5127
R18007 vdd.n2336 vdd.n974 99.5127
R18008 vdd.n2340 vdd.n974 99.5127
R18009 vdd.n2340 vdd.n965 99.5127
R18010 vdd.n2348 vdd.n965 99.5127
R18011 vdd.n2348 vdd.n963 99.5127
R18012 vdd.n2352 vdd.n963 99.5127
R18013 vdd.n2352 vdd.n953 99.5127
R18014 vdd.n2360 vdd.n953 99.5127
R18015 vdd.n2360 vdd.n950 99.5127
R18016 vdd.n2366 vdd.n950 99.5127
R18017 vdd.n2366 vdd.n951 99.5127
R18018 vdd.n951 vdd.n942 99.5127
R18019 vdd.n942 vdd.n933 99.5127
R18020 vdd.n2448 vdd.n933 99.5127
R18021 vdd.n9 vdd.n7 98.9633
R18022 vdd.n2 vdd.n0 98.9633
R18023 vdd.n9 vdd.n8 98.6055
R18024 vdd.n11 vdd.n10 98.6055
R18025 vdd.n13 vdd.n12 98.6055
R18026 vdd.n6 vdd.n5 98.6055
R18027 vdd.n4 vdd.n3 98.6055
R18028 vdd.n2 vdd.n1 98.6055
R18029 vdd.t148 vdd.n291 85.8723
R18030 vdd.t125 vdd.n236 85.8723
R18031 vdd.t137 vdd.n193 85.8723
R18032 vdd.t113 vdd.n138 85.8723
R18033 vdd.t70 vdd.n96 85.8723
R18034 vdd.t47 vdd.n41 85.8723
R18035 vdd.t163 vdd.n1660 85.8723
R18036 vdd.t73 vdd.n1715 85.8723
R18037 vdd.t149 vdd.n1562 85.8723
R18038 vdd.t57 vdd.n1617 85.8723
R18039 vdd.t51 vdd.n1465 85.8723
R18040 vdd.t72 vdd.n1520 85.8723
R18041 vdd.n2840 vdd.n2839 78.546
R18042 vdd.n2314 vdd.n998 78.546
R18043 vdd.n278 vdd.n277 75.1835
R18044 vdd.n276 vdd.n275 75.1835
R18045 vdd.n274 vdd.n273 75.1835
R18046 vdd.n272 vdd.n271 75.1835
R18047 vdd.n270 vdd.n269 75.1835
R18048 vdd.n268 vdd.n267 75.1835
R18049 vdd.n266 vdd.n265 75.1835
R18050 vdd.n180 vdd.n179 75.1835
R18051 vdd.n178 vdd.n177 75.1835
R18052 vdd.n176 vdd.n175 75.1835
R18053 vdd.n174 vdd.n173 75.1835
R18054 vdd.n172 vdd.n171 75.1835
R18055 vdd.n170 vdd.n169 75.1835
R18056 vdd.n168 vdd.n167 75.1835
R18057 vdd.n83 vdd.n82 75.1835
R18058 vdd.n81 vdd.n80 75.1835
R18059 vdd.n79 vdd.n78 75.1835
R18060 vdd.n77 vdd.n76 75.1835
R18061 vdd.n75 vdd.n74 75.1835
R18062 vdd.n73 vdd.n72 75.1835
R18063 vdd.n71 vdd.n70 75.1835
R18064 vdd.n1690 vdd.n1689 75.1835
R18065 vdd.n1692 vdd.n1691 75.1835
R18066 vdd.n1694 vdd.n1693 75.1835
R18067 vdd.n1696 vdd.n1695 75.1835
R18068 vdd.n1698 vdd.n1697 75.1835
R18069 vdd.n1700 vdd.n1699 75.1835
R18070 vdd.n1702 vdd.n1701 75.1835
R18071 vdd.n1592 vdd.n1591 75.1835
R18072 vdd.n1594 vdd.n1593 75.1835
R18073 vdd.n1596 vdd.n1595 75.1835
R18074 vdd.n1598 vdd.n1597 75.1835
R18075 vdd.n1600 vdd.n1599 75.1835
R18076 vdd.n1602 vdd.n1601 75.1835
R18077 vdd.n1604 vdd.n1603 75.1835
R18078 vdd.n1495 vdd.n1494 75.1835
R18079 vdd.n1497 vdd.n1496 75.1835
R18080 vdd.n1499 vdd.n1498 75.1835
R18081 vdd.n1501 vdd.n1500 75.1835
R18082 vdd.n1503 vdd.n1502 75.1835
R18083 vdd.n1505 vdd.n1504 75.1835
R18084 vdd.n1507 vdd.n1506 75.1835
R18085 vdd.n2775 vdd.n2774 72.8958
R18086 vdd.n2774 vdd.n2538 72.8958
R18087 vdd.n2774 vdd.n2539 72.8958
R18088 vdd.n2774 vdd.n2540 72.8958
R18089 vdd.n2774 vdd.n2541 72.8958
R18090 vdd.n2774 vdd.n2542 72.8958
R18091 vdd.n2774 vdd.n2543 72.8958
R18092 vdd.n2774 vdd.n2544 72.8958
R18093 vdd.n2774 vdd.n2545 72.8958
R18094 vdd.n2774 vdd.n2546 72.8958
R18095 vdd.n2774 vdd.n2547 72.8958
R18096 vdd.n2774 vdd.n2548 72.8958
R18097 vdd.n2774 vdd.n2549 72.8958
R18098 vdd.n2774 vdd.n2550 72.8958
R18099 vdd.n2774 vdd.n2551 72.8958
R18100 vdd.n2774 vdd.n2552 72.8958
R18101 vdd.n2774 vdd.n2553 72.8958
R18102 vdd.n772 vdd.n756 72.8958
R18103 vdd.n2983 vdd.n756 72.8958
R18104 vdd.n766 vdd.n756 72.8958
R18105 vdd.n2990 vdd.n756 72.8958
R18106 vdd.n763 vdd.n756 72.8958
R18107 vdd.n2997 vdd.n756 72.8958
R18108 vdd.n760 vdd.n756 72.8958
R18109 vdd.n3004 vdd.n756 72.8958
R18110 vdd.n3007 vdd.n756 72.8958
R18111 vdd.n2863 vdd.n756 72.8958
R18112 vdd.n2868 vdd.n756 72.8958
R18113 vdd.n2862 vdd.n756 72.8958
R18114 vdd.n2875 vdd.n756 72.8958
R18115 vdd.n2859 vdd.n756 72.8958
R18116 vdd.n2882 vdd.n756 72.8958
R18117 vdd.n2856 vdd.n756 72.8958
R18118 vdd.n2889 vdd.n756 72.8958
R18119 vdd.n2027 vdd.n1020 72.8958
R18120 vdd.n2033 vdd.n1020 72.8958
R18121 vdd.n2035 vdd.n1020 72.8958
R18122 vdd.n2041 vdd.n1020 72.8958
R18123 vdd.n2043 vdd.n1020 72.8958
R18124 vdd.n2049 vdd.n1020 72.8958
R18125 vdd.n2051 vdd.n1020 72.8958
R18126 vdd.n2057 vdd.n1020 72.8958
R18127 vdd.n2228 vdd.n1020 72.8958
R18128 vdd.n2226 vdd.n1020 72.8958
R18129 vdd.n2220 vdd.n1020 72.8958
R18130 vdd.n2218 vdd.n1020 72.8958
R18131 vdd.n2212 vdd.n1020 72.8958
R18132 vdd.n2210 vdd.n1020 72.8958
R18133 vdd.n2204 vdd.n1020 72.8958
R18134 vdd.n2202 vdd.n1020 72.8958
R18135 vdd.n2196 vdd.n1020 72.8958
R18136 vdd.n2521 vdd.n908 72.8958
R18137 vdd.n2521 vdd.n909 72.8958
R18138 vdd.n2521 vdd.n910 72.8958
R18139 vdd.n2521 vdd.n911 72.8958
R18140 vdd.n2521 vdd.n912 72.8958
R18141 vdd.n2521 vdd.n913 72.8958
R18142 vdd.n2521 vdd.n914 72.8958
R18143 vdd.n2521 vdd.n915 72.8958
R18144 vdd.n2521 vdd.n916 72.8958
R18145 vdd.n2521 vdd.n917 72.8958
R18146 vdd.n2521 vdd.n918 72.8958
R18147 vdd.n2521 vdd.n919 72.8958
R18148 vdd.n2521 vdd.n920 72.8958
R18149 vdd.n2521 vdd.n921 72.8958
R18150 vdd.n2521 vdd.n922 72.8958
R18151 vdd.n2521 vdd.n923 72.8958
R18152 vdd.n2521 vdd.n924 72.8958
R18153 vdd.n2774 vdd.n2773 72.8958
R18154 vdd.n2774 vdd.n2522 72.8958
R18155 vdd.n2774 vdd.n2523 72.8958
R18156 vdd.n2774 vdd.n2524 72.8958
R18157 vdd.n2774 vdd.n2525 72.8958
R18158 vdd.n2774 vdd.n2526 72.8958
R18159 vdd.n2774 vdd.n2527 72.8958
R18160 vdd.n2774 vdd.n2528 72.8958
R18161 vdd.n2774 vdd.n2529 72.8958
R18162 vdd.n2774 vdd.n2530 72.8958
R18163 vdd.n2774 vdd.n2531 72.8958
R18164 vdd.n2774 vdd.n2532 72.8958
R18165 vdd.n2774 vdd.n2533 72.8958
R18166 vdd.n2774 vdd.n2534 72.8958
R18167 vdd.n2774 vdd.n2535 72.8958
R18168 vdd.n2774 vdd.n2536 72.8958
R18169 vdd.n2774 vdd.n2537 72.8958
R18170 vdd.n2911 vdd.n756 72.8958
R18171 vdd.n2917 vdd.n756 72.8958
R18172 vdd.n802 vdd.n756 72.8958
R18173 vdd.n2924 vdd.n756 72.8958
R18174 vdd.n799 vdd.n756 72.8958
R18175 vdd.n2931 vdd.n756 72.8958
R18176 vdd.n796 vdd.n756 72.8958
R18177 vdd.n2938 vdd.n756 72.8958
R18178 vdd.n793 vdd.n756 72.8958
R18179 vdd.n2946 vdd.n756 72.8958
R18180 vdd.n790 vdd.n756 72.8958
R18181 vdd.n2953 vdd.n756 72.8958
R18182 vdd.n787 vdd.n756 72.8958
R18183 vdd.n2960 vdd.n756 72.8958
R18184 vdd.n784 vdd.n756 72.8958
R18185 vdd.n2967 vdd.n756 72.8958
R18186 vdd.n2970 vdd.n756 72.8958
R18187 vdd.n2521 vdd.n906 72.8958
R18188 vdd.n2521 vdd.n905 72.8958
R18189 vdd.n2521 vdd.n904 72.8958
R18190 vdd.n2521 vdd.n903 72.8958
R18191 vdd.n2521 vdd.n902 72.8958
R18192 vdd.n2521 vdd.n901 72.8958
R18193 vdd.n2521 vdd.n900 72.8958
R18194 vdd.n2521 vdd.n899 72.8958
R18195 vdd.n2521 vdd.n898 72.8958
R18196 vdd.n2521 vdd.n897 72.8958
R18197 vdd.n2521 vdd.n896 72.8958
R18198 vdd.n2521 vdd.n895 72.8958
R18199 vdd.n2521 vdd.n894 72.8958
R18200 vdd.n2521 vdd.n893 72.8958
R18201 vdd.n2521 vdd.n892 72.8958
R18202 vdd.n2521 vdd.n891 72.8958
R18203 vdd.n2521 vdd.n890 72.8958
R18204 vdd.n2286 vdd.n1020 72.8958
R18205 vdd.n2284 vdd.n1020 72.8958
R18206 vdd.n2278 vdd.n1020 72.8958
R18207 vdd.n2276 vdd.n1020 72.8958
R18208 vdd.n2270 vdd.n1020 72.8958
R18209 vdd.n2268 vdd.n1020 72.8958
R18210 vdd.n2262 vdd.n1020 72.8958
R18211 vdd.n2260 vdd.n1020 72.8958
R18212 vdd.n1032 vdd.n1020 72.8958
R18213 vdd.n2102 vdd.n1020 72.8958
R18214 vdd.n2107 vdd.n1020 72.8958
R18215 vdd.n2109 vdd.n1020 72.8958
R18216 vdd.n2115 vdd.n1020 72.8958
R18217 vdd.n2117 vdd.n1020 72.8958
R18218 vdd.n2123 vdd.n1020 72.8958
R18219 vdd.n2125 vdd.n1020 72.8958
R18220 vdd.n2132 vdd.n1020 72.8958
R18221 vdd.n1374 vdd.n1373 66.2847
R18222 vdd.n1374 vdd.n1152 66.2847
R18223 vdd.n1374 vdd.n1153 66.2847
R18224 vdd.n1374 vdd.n1154 66.2847
R18225 vdd.n1374 vdd.n1155 66.2847
R18226 vdd.n1374 vdd.n1156 66.2847
R18227 vdd.n1374 vdd.n1157 66.2847
R18228 vdd.n1374 vdd.n1158 66.2847
R18229 vdd.n1374 vdd.n1159 66.2847
R18230 vdd.n1374 vdd.n1160 66.2847
R18231 vdd.n1374 vdd.n1161 66.2847
R18232 vdd.n1374 vdd.n1162 66.2847
R18233 vdd.n1374 vdd.n1163 66.2847
R18234 vdd.n1374 vdd.n1164 66.2847
R18235 vdd.n1374 vdd.n1165 66.2847
R18236 vdd.n1374 vdd.n1166 66.2847
R18237 vdd.n1374 vdd.n1167 66.2847
R18238 vdd.n1374 vdd.n1168 66.2847
R18239 vdd.n1374 vdd.n1169 66.2847
R18240 vdd.n1374 vdd.n1170 66.2847
R18241 vdd.n1374 vdd.n1171 66.2847
R18242 vdd.n1374 vdd.n1172 66.2847
R18243 vdd.n1374 vdd.n1173 66.2847
R18244 vdd.n1374 vdd.n1174 66.2847
R18245 vdd.n1374 vdd.n1175 66.2847
R18246 vdd.n1374 vdd.n1176 66.2847
R18247 vdd.n1374 vdd.n1177 66.2847
R18248 vdd.n1374 vdd.n1178 66.2847
R18249 vdd.n1374 vdd.n1179 66.2847
R18250 vdd.n1374 vdd.n1180 66.2847
R18251 vdd.n1374 vdd.n1181 66.2847
R18252 vdd.n1045 vdd.n1041 66.2847
R18253 vdd.n1917 vdd.n1045 66.2847
R18254 vdd.n1922 vdd.n1045 66.2847
R18255 vdd.n1927 vdd.n1045 66.2847
R18256 vdd.n1915 vdd.n1045 66.2847
R18257 vdd.n1934 vdd.n1045 66.2847
R18258 vdd.n1907 vdd.n1045 66.2847
R18259 vdd.n1941 vdd.n1045 66.2847
R18260 vdd.n1900 vdd.n1045 66.2847
R18261 vdd.n1948 vdd.n1045 66.2847
R18262 vdd.n1894 vdd.n1045 66.2847
R18263 vdd.n1889 vdd.n1045 66.2847
R18264 vdd.n1959 vdd.n1045 66.2847
R18265 vdd.n1881 vdd.n1045 66.2847
R18266 vdd.n1966 vdd.n1045 66.2847
R18267 vdd.n1874 vdd.n1045 66.2847
R18268 vdd.n1973 vdd.n1045 66.2847
R18269 vdd.n1867 vdd.n1045 66.2847
R18270 vdd.n1980 vdd.n1045 66.2847
R18271 vdd.n1860 vdd.n1045 66.2847
R18272 vdd.n1987 vdd.n1045 66.2847
R18273 vdd.n1854 vdd.n1045 66.2847
R18274 vdd.n1849 vdd.n1045 66.2847
R18275 vdd.n1998 vdd.n1045 66.2847
R18276 vdd.n1841 vdd.n1045 66.2847
R18277 vdd.n2005 vdd.n1045 66.2847
R18278 vdd.n1834 vdd.n1045 66.2847
R18279 vdd.n2012 vdd.n1045 66.2847
R18280 vdd.n2015 vdd.n1045 66.2847
R18281 vdd.n1825 vdd.n1045 66.2847
R18282 vdd.n2237 vdd.n1045 66.2847
R18283 vdd.n1819 vdd.n1045 66.2847
R18284 vdd.n3137 vdd.n658 66.2847
R18285 vdd.n663 vdd.n658 66.2847
R18286 vdd.n666 vdd.n658 66.2847
R18287 vdd.n3126 vdd.n658 66.2847
R18288 vdd.n3120 vdd.n658 66.2847
R18289 vdd.n3118 vdd.n658 66.2847
R18290 vdd.n3112 vdd.n658 66.2847
R18291 vdd.n3110 vdd.n658 66.2847
R18292 vdd.n3104 vdd.n658 66.2847
R18293 vdd.n3102 vdd.n658 66.2847
R18294 vdd.n3096 vdd.n658 66.2847
R18295 vdd.n3094 vdd.n658 66.2847
R18296 vdd.n3088 vdd.n658 66.2847
R18297 vdd.n3086 vdd.n658 66.2847
R18298 vdd.n3080 vdd.n658 66.2847
R18299 vdd.n3078 vdd.n658 66.2847
R18300 vdd.n3072 vdd.n658 66.2847
R18301 vdd.n3070 vdd.n658 66.2847
R18302 vdd.n3064 vdd.n658 66.2847
R18303 vdd.n3062 vdd.n658 66.2847
R18304 vdd.n727 vdd.n658 66.2847
R18305 vdd.n3053 vdd.n658 66.2847
R18306 vdd.n729 vdd.n658 66.2847
R18307 vdd.n3046 vdd.n658 66.2847
R18308 vdd.n3040 vdd.n658 66.2847
R18309 vdd.n3038 vdd.n658 66.2847
R18310 vdd.n3032 vdd.n658 66.2847
R18311 vdd.n3030 vdd.n658 66.2847
R18312 vdd.n3024 vdd.n658 66.2847
R18313 vdd.n750 vdd.n658 66.2847
R18314 vdd.n752 vdd.n658 66.2847
R18315 vdd.n3253 vdd.n3252 66.2847
R18316 vdd.n3253 vdd.n403 66.2847
R18317 vdd.n3253 vdd.n402 66.2847
R18318 vdd.n3253 vdd.n401 66.2847
R18319 vdd.n3253 vdd.n400 66.2847
R18320 vdd.n3253 vdd.n399 66.2847
R18321 vdd.n3253 vdd.n398 66.2847
R18322 vdd.n3253 vdd.n397 66.2847
R18323 vdd.n3253 vdd.n396 66.2847
R18324 vdd.n3253 vdd.n395 66.2847
R18325 vdd.n3253 vdd.n394 66.2847
R18326 vdd.n3253 vdd.n393 66.2847
R18327 vdd.n3253 vdd.n392 66.2847
R18328 vdd.n3253 vdd.n391 66.2847
R18329 vdd.n3253 vdd.n390 66.2847
R18330 vdd.n3253 vdd.n389 66.2847
R18331 vdd.n3253 vdd.n388 66.2847
R18332 vdd.n3253 vdd.n387 66.2847
R18333 vdd.n3253 vdd.n386 66.2847
R18334 vdd.n3253 vdd.n385 66.2847
R18335 vdd.n3253 vdd.n384 66.2847
R18336 vdd.n3253 vdd.n383 66.2847
R18337 vdd.n3253 vdd.n382 66.2847
R18338 vdd.n3253 vdd.n381 66.2847
R18339 vdd.n3253 vdd.n380 66.2847
R18340 vdd.n3253 vdd.n379 66.2847
R18341 vdd.n3253 vdd.n378 66.2847
R18342 vdd.n3253 vdd.n377 66.2847
R18343 vdd.n3253 vdd.n376 66.2847
R18344 vdd.n3253 vdd.n375 66.2847
R18345 vdd.n3253 vdd.n374 66.2847
R18346 vdd.n3253 vdd.n373 66.2847
R18347 vdd.n448 vdd.n373 52.4337
R18348 vdd.n454 vdd.n374 52.4337
R18349 vdd.n458 vdd.n375 52.4337
R18350 vdd.n464 vdd.n376 52.4337
R18351 vdd.n468 vdd.n377 52.4337
R18352 vdd.n474 vdd.n378 52.4337
R18353 vdd.n478 vdd.n379 52.4337
R18354 vdd.n484 vdd.n380 52.4337
R18355 vdd.n488 vdd.n381 52.4337
R18356 vdd.n494 vdd.n382 52.4337
R18357 vdd.n498 vdd.n383 52.4337
R18358 vdd.n504 vdd.n384 52.4337
R18359 vdd.n508 vdd.n385 52.4337
R18360 vdd.n514 vdd.n386 52.4337
R18361 vdd.n518 vdd.n387 52.4337
R18362 vdd.n524 vdd.n388 52.4337
R18363 vdd.n528 vdd.n389 52.4337
R18364 vdd.n534 vdd.n390 52.4337
R18365 vdd.n538 vdd.n391 52.4337
R18366 vdd.n544 vdd.n392 52.4337
R18367 vdd.n548 vdd.n393 52.4337
R18368 vdd.n554 vdd.n394 52.4337
R18369 vdd.n558 vdd.n395 52.4337
R18370 vdd.n564 vdd.n396 52.4337
R18371 vdd.n568 vdd.n397 52.4337
R18372 vdd.n574 vdd.n398 52.4337
R18373 vdd.n578 vdd.n399 52.4337
R18374 vdd.n584 vdd.n400 52.4337
R18375 vdd.n588 vdd.n401 52.4337
R18376 vdd.n594 vdd.n402 52.4337
R18377 vdd.n597 vdd.n403 52.4337
R18378 vdd.n3252 vdd.n3251 52.4337
R18379 vdd.n3137 vdd.n660 52.4337
R18380 vdd.n3135 vdd.n663 52.4337
R18381 vdd.n3131 vdd.n666 52.4337
R18382 vdd.n3127 vdd.n3126 52.4337
R18383 vdd.n3120 vdd.n669 52.4337
R18384 vdd.n3119 vdd.n3118 52.4337
R18385 vdd.n3112 vdd.n675 52.4337
R18386 vdd.n3111 vdd.n3110 52.4337
R18387 vdd.n3104 vdd.n681 52.4337
R18388 vdd.n3103 vdd.n3102 52.4337
R18389 vdd.n3096 vdd.n689 52.4337
R18390 vdd.n3095 vdd.n3094 52.4337
R18391 vdd.n3088 vdd.n695 52.4337
R18392 vdd.n3087 vdd.n3086 52.4337
R18393 vdd.n3080 vdd.n701 52.4337
R18394 vdd.n3079 vdd.n3078 52.4337
R18395 vdd.n3072 vdd.n707 52.4337
R18396 vdd.n3071 vdd.n3070 52.4337
R18397 vdd.n3064 vdd.n713 52.4337
R18398 vdd.n3063 vdd.n3062 52.4337
R18399 vdd.n727 vdd.n719 52.4337
R18400 vdd.n3054 vdd.n3053 52.4337
R18401 vdd.n3051 vdd.n729 52.4337
R18402 vdd.n3047 vdd.n3046 52.4337
R18403 vdd.n3040 vdd.n733 52.4337
R18404 vdd.n3039 vdd.n3038 52.4337
R18405 vdd.n3032 vdd.n739 52.4337
R18406 vdd.n3031 vdd.n3030 52.4337
R18407 vdd.n3024 vdd.n745 52.4337
R18408 vdd.n3023 vdd.n750 52.4337
R18409 vdd.n3019 vdd.n752 52.4337
R18410 vdd.n2239 vdd.n1819 52.4337
R18411 vdd.n2237 vdd.n2236 52.4337
R18412 vdd.n1826 vdd.n1825 52.4337
R18413 vdd.n2015 vdd.n2014 52.4337
R18414 vdd.n2012 vdd.n2011 52.4337
R18415 vdd.n2007 vdd.n1834 52.4337
R18416 vdd.n2005 vdd.n2004 52.4337
R18417 vdd.n2000 vdd.n1841 52.4337
R18418 vdd.n1998 vdd.n1997 52.4337
R18419 vdd.n1850 vdd.n1849 52.4337
R18420 vdd.n1989 vdd.n1854 52.4337
R18421 vdd.n1987 vdd.n1986 52.4337
R18422 vdd.n1982 vdd.n1860 52.4337
R18423 vdd.n1980 vdd.n1979 52.4337
R18424 vdd.n1975 vdd.n1867 52.4337
R18425 vdd.n1973 vdd.n1972 52.4337
R18426 vdd.n1968 vdd.n1874 52.4337
R18427 vdd.n1966 vdd.n1965 52.4337
R18428 vdd.n1961 vdd.n1881 52.4337
R18429 vdd.n1959 vdd.n1958 52.4337
R18430 vdd.n1890 vdd.n1889 52.4337
R18431 vdd.n1950 vdd.n1894 52.4337
R18432 vdd.n1948 vdd.n1947 52.4337
R18433 vdd.n1943 vdd.n1900 52.4337
R18434 vdd.n1941 vdd.n1940 52.4337
R18435 vdd.n1936 vdd.n1907 52.4337
R18436 vdd.n1934 vdd.n1933 52.4337
R18437 vdd.n1929 vdd.n1915 52.4337
R18438 vdd.n1927 vdd.n1926 52.4337
R18439 vdd.n1922 vdd.n1921 52.4337
R18440 vdd.n1917 vdd.n1916 52.4337
R18441 vdd.n2248 vdd.n1041 52.4337
R18442 vdd.n1373 vdd.n1372 52.4337
R18443 vdd.n1187 vdd.n1152 52.4337
R18444 vdd.n1189 vdd.n1153 52.4337
R18445 vdd.n1193 vdd.n1154 52.4337
R18446 vdd.n1195 vdd.n1155 52.4337
R18447 vdd.n1199 vdd.n1156 52.4337
R18448 vdd.n1201 vdd.n1157 52.4337
R18449 vdd.n1205 vdd.n1158 52.4337
R18450 vdd.n1207 vdd.n1159 52.4337
R18451 vdd.n1339 vdd.n1160 52.4337
R18452 vdd.n1211 vdd.n1161 52.4337
R18453 vdd.n1215 vdd.n1162 52.4337
R18454 vdd.n1217 vdd.n1163 52.4337
R18455 vdd.n1221 vdd.n1164 52.4337
R18456 vdd.n1223 vdd.n1165 52.4337
R18457 vdd.n1227 vdd.n1166 52.4337
R18458 vdd.n1229 vdd.n1167 52.4337
R18459 vdd.n1233 vdd.n1168 52.4337
R18460 vdd.n1235 vdd.n1169 52.4337
R18461 vdd.n1239 vdd.n1170 52.4337
R18462 vdd.n1303 vdd.n1171 52.4337
R18463 vdd.n1244 vdd.n1172 52.4337
R18464 vdd.n1246 vdd.n1173 52.4337
R18465 vdd.n1250 vdd.n1174 52.4337
R18466 vdd.n1252 vdd.n1175 52.4337
R18467 vdd.n1256 vdd.n1176 52.4337
R18468 vdd.n1258 vdd.n1177 52.4337
R18469 vdd.n1262 vdd.n1178 52.4337
R18470 vdd.n1264 vdd.n1179 52.4337
R18471 vdd.n1268 vdd.n1180 52.4337
R18472 vdd.n1270 vdd.n1181 52.4337
R18473 vdd.n1373 vdd.n1183 52.4337
R18474 vdd.n1188 vdd.n1152 52.4337
R18475 vdd.n1192 vdd.n1153 52.4337
R18476 vdd.n1194 vdd.n1154 52.4337
R18477 vdd.n1198 vdd.n1155 52.4337
R18478 vdd.n1200 vdd.n1156 52.4337
R18479 vdd.n1204 vdd.n1157 52.4337
R18480 vdd.n1206 vdd.n1158 52.4337
R18481 vdd.n1338 vdd.n1159 52.4337
R18482 vdd.n1210 vdd.n1160 52.4337
R18483 vdd.n1214 vdd.n1161 52.4337
R18484 vdd.n1216 vdd.n1162 52.4337
R18485 vdd.n1220 vdd.n1163 52.4337
R18486 vdd.n1222 vdd.n1164 52.4337
R18487 vdd.n1226 vdd.n1165 52.4337
R18488 vdd.n1228 vdd.n1166 52.4337
R18489 vdd.n1232 vdd.n1167 52.4337
R18490 vdd.n1234 vdd.n1168 52.4337
R18491 vdd.n1238 vdd.n1169 52.4337
R18492 vdd.n1240 vdd.n1170 52.4337
R18493 vdd.n1243 vdd.n1171 52.4337
R18494 vdd.n1245 vdd.n1172 52.4337
R18495 vdd.n1249 vdd.n1173 52.4337
R18496 vdd.n1251 vdd.n1174 52.4337
R18497 vdd.n1255 vdd.n1175 52.4337
R18498 vdd.n1257 vdd.n1176 52.4337
R18499 vdd.n1261 vdd.n1177 52.4337
R18500 vdd.n1263 vdd.n1178 52.4337
R18501 vdd.n1267 vdd.n1179 52.4337
R18502 vdd.n1269 vdd.n1180 52.4337
R18503 vdd.n1181 vdd.n1151 52.4337
R18504 vdd.n1041 vdd.n1040 52.4337
R18505 vdd.n1918 vdd.n1917 52.4337
R18506 vdd.n1923 vdd.n1922 52.4337
R18507 vdd.n1928 vdd.n1927 52.4337
R18508 vdd.n1915 vdd.n1908 52.4337
R18509 vdd.n1935 vdd.n1934 52.4337
R18510 vdd.n1907 vdd.n1901 52.4337
R18511 vdd.n1942 vdd.n1941 52.4337
R18512 vdd.n1900 vdd.n1895 52.4337
R18513 vdd.n1949 vdd.n1948 52.4337
R18514 vdd.n1894 vdd.n1893 52.4337
R18515 vdd.n1889 vdd.n1882 52.4337
R18516 vdd.n1960 vdd.n1959 52.4337
R18517 vdd.n1881 vdd.n1875 52.4337
R18518 vdd.n1967 vdd.n1966 52.4337
R18519 vdd.n1874 vdd.n1868 52.4337
R18520 vdd.n1974 vdd.n1973 52.4337
R18521 vdd.n1867 vdd.n1861 52.4337
R18522 vdd.n1981 vdd.n1980 52.4337
R18523 vdd.n1860 vdd.n1855 52.4337
R18524 vdd.n1988 vdd.n1987 52.4337
R18525 vdd.n1854 vdd.n1853 52.4337
R18526 vdd.n1849 vdd.n1842 52.4337
R18527 vdd.n1999 vdd.n1998 52.4337
R18528 vdd.n1841 vdd.n1835 52.4337
R18529 vdd.n2006 vdd.n2005 52.4337
R18530 vdd.n1834 vdd.n1828 52.4337
R18531 vdd.n2013 vdd.n2012 52.4337
R18532 vdd.n2016 vdd.n2015 52.4337
R18533 vdd.n1825 vdd.n1820 52.4337
R18534 vdd.n2238 vdd.n2237 52.4337
R18535 vdd.n1819 vdd.n1047 52.4337
R18536 vdd.n3138 vdd.n3137 52.4337
R18537 vdd.n3132 vdd.n663 52.4337
R18538 vdd.n3128 vdd.n666 52.4337
R18539 vdd.n3126 vdd.n3125 52.4337
R18540 vdd.n3121 vdd.n3120 52.4337
R18541 vdd.n3118 vdd.n3117 52.4337
R18542 vdd.n3113 vdd.n3112 52.4337
R18543 vdd.n3110 vdd.n3109 52.4337
R18544 vdd.n3105 vdd.n3104 52.4337
R18545 vdd.n3102 vdd.n3101 52.4337
R18546 vdd.n3097 vdd.n3096 52.4337
R18547 vdd.n3094 vdd.n3093 52.4337
R18548 vdd.n3089 vdd.n3088 52.4337
R18549 vdd.n3086 vdd.n3085 52.4337
R18550 vdd.n3081 vdd.n3080 52.4337
R18551 vdd.n3078 vdd.n3077 52.4337
R18552 vdd.n3073 vdd.n3072 52.4337
R18553 vdd.n3070 vdd.n3069 52.4337
R18554 vdd.n3065 vdd.n3064 52.4337
R18555 vdd.n3062 vdd.n3061 52.4337
R18556 vdd.n728 vdd.n727 52.4337
R18557 vdd.n3053 vdd.n3052 52.4337
R18558 vdd.n3048 vdd.n729 52.4337
R18559 vdd.n3046 vdd.n3045 52.4337
R18560 vdd.n3041 vdd.n3040 52.4337
R18561 vdd.n3038 vdd.n3037 52.4337
R18562 vdd.n3033 vdd.n3032 52.4337
R18563 vdd.n3030 vdd.n3029 52.4337
R18564 vdd.n3025 vdd.n3024 52.4337
R18565 vdd.n3020 vdd.n750 52.4337
R18566 vdd.n3016 vdd.n752 52.4337
R18567 vdd.n3252 vdd.n404 52.4337
R18568 vdd.n595 vdd.n403 52.4337
R18569 vdd.n589 vdd.n402 52.4337
R18570 vdd.n585 vdd.n401 52.4337
R18571 vdd.n579 vdd.n400 52.4337
R18572 vdd.n575 vdd.n399 52.4337
R18573 vdd.n569 vdd.n398 52.4337
R18574 vdd.n565 vdd.n397 52.4337
R18575 vdd.n559 vdd.n396 52.4337
R18576 vdd.n555 vdd.n395 52.4337
R18577 vdd.n549 vdd.n394 52.4337
R18578 vdd.n545 vdd.n393 52.4337
R18579 vdd.n539 vdd.n392 52.4337
R18580 vdd.n535 vdd.n391 52.4337
R18581 vdd.n529 vdd.n390 52.4337
R18582 vdd.n525 vdd.n389 52.4337
R18583 vdd.n519 vdd.n388 52.4337
R18584 vdd.n515 vdd.n387 52.4337
R18585 vdd.n509 vdd.n386 52.4337
R18586 vdd.n505 vdd.n385 52.4337
R18587 vdd.n499 vdd.n384 52.4337
R18588 vdd.n495 vdd.n383 52.4337
R18589 vdd.n489 vdd.n382 52.4337
R18590 vdd.n485 vdd.n381 52.4337
R18591 vdd.n479 vdd.n380 52.4337
R18592 vdd.n475 vdd.n379 52.4337
R18593 vdd.n469 vdd.n378 52.4337
R18594 vdd.n465 vdd.n377 52.4337
R18595 vdd.n459 vdd.n376 52.4337
R18596 vdd.n455 vdd.n375 52.4337
R18597 vdd.n449 vdd.n374 52.4337
R18598 vdd.n445 vdd.n373 52.4337
R18599 vdd.t19 vdd.t248 51.4683
R18600 vdd.n266 vdd.n264 42.0461
R18601 vdd.n168 vdd.n166 42.0461
R18602 vdd.n71 vdd.n69 42.0461
R18603 vdd.n1690 vdd.n1688 42.0461
R18604 vdd.n1592 vdd.n1590 42.0461
R18605 vdd.n1495 vdd.n1493 42.0461
R18606 vdd.n320 vdd.n319 41.6884
R18607 vdd.n222 vdd.n221 41.6884
R18608 vdd.n125 vdd.n124 41.6884
R18609 vdd.n1744 vdd.n1743 41.6884
R18610 vdd.n1646 vdd.n1645 41.6884
R18611 vdd.n1549 vdd.n1548 41.6884
R18612 vdd.n1150 vdd.n1149 41.1157
R18613 vdd.n1306 vdd.n1305 41.1157
R18614 vdd.n1342 vdd.n1341 41.1157
R18615 vdd.n407 vdd.n406 41.1157
R18616 vdd.n547 vdd.n420 41.1157
R18617 vdd.n433 vdd.n432 41.1157
R18618 vdd.n2970 vdd.n2969 39.2114
R18619 vdd.n2967 vdd.n2966 39.2114
R18620 vdd.n2962 vdd.n784 39.2114
R18621 vdd.n2960 vdd.n2959 39.2114
R18622 vdd.n2955 vdd.n787 39.2114
R18623 vdd.n2953 vdd.n2952 39.2114
R18624 vdd.n2948 vdd.n790 39.2114
R18625 vdd.n2946 vdd.n2945 39.2114
R18626 vdd.n2940 vdd.n793 39.2114
R18627 vdd.n2938 vdd.n2937 39.2114
R18628 vdd.n2933 vdd.n796 39.2114
R18629 vdd.n2931 vdd.n2930 39.2114
R18630 vdd.n2926 vdd.n799 39.2114
R18631 vdd.n2924 vdd.n2923 39.2114
R18632 vdd.n2919 vdd.n802 39.2114
R18633 vdd.n2917 vdd.n2916 39.2114
R18634 vdd.n2912 vdd.n2911 39.2114
R18635 vdd.n2773 vdd.n884 39.2114
R18636 vdd.n2768 vdd.n2522 39.2114
R18637 vdd.n2765 vdd.n2523 39.2114
R18638 vdd.n2761 vdd.n2524 39.2114
R18639 vdd.n2757 vdd.n2525 39.2114
R18640 vdd.n2753 vdd.n2526 39.2114
R18641 vdd.n2749 vdd.n2527 39.2114
R18642 vdd.n2745 vdd.n2528 39.2114
R18643 vdd.n2741 vdd.n2529 39.2114
R18644 vdd.n2737 vdd.n2530 39.2114
R18645 vdd.n2733 vdd.n2531 39.2114
R18646 vdd.n2729 vdd.n2532 39.2114
R18647 vdd.n2725 vdd.n2533 39.2114
R18648 vdd.n2721 vdd.n2534 39.2114
R18649 vdd.n2717 vdd.n2535 39.2114
R18650 vdd.n2713 vdd.n2536 39.2114
R18651 vdd.n2708 vdd.n2537 39.2114
R18652 vdd.n2516 vdd.n924 39.2114
R18653 vdd.n2512 vdd.n923 39.2114
R18654 vdd.n2508 vdd.n922 39.2114
R18655 vdd.n2504 vdd.n921 39.2114
R18656 vdd.n2500 vdd.n920 39.2114
R18657 vdd.n2496 vdd.n919 39.2114
R18658 vdd.n2492 vdd.n918 39.2114
R18659 vdd.n2488 vdd.n917 39.2114
R18660 vdd.n2484 vdd.n916 39.2114
R18661 vdd.n2480 vdd.n915 39.2114
R18662 vdd.n2476 vdd.n914 39.2114
R18663 vdd.n2472 vdd.n913 39.2114
R18664 vdd.n2468 vdd.n912 39.2114
R18665 vdd.n2464 vdd.n911 39.2114
R18666 vdd.n2460 vdd.n910 39.2114
R18667 vdd.n2455 vdd.n909 39.2114
R18668 vdd.n2451 vdd.n908 39.2114
R18669 vdd.n2027 vdd.n1019 39.2114
R18670 vdd.n2033 vdd.n2032 39.2114
R18671 vdd.n2036 vdd.n2035 39.2114
R18672 vdd.n2041 vdd.n2040 39.2114
R18673 vdd.n2044 vdd.n2043 39.2114
R18674 vdd.n2049 vdd.n2048 39.2114
R18675 vdd.n2052 vdd.n2051 39.2114
R18676 vdd.n2057 vdd.n2056 39.2114
R18677 vdd.n2228 vdd.n2059 39.2114
R18678 vdd.n2227 vdd.n2226 39.2114
R18679 vdd.n2220 vdd.n2061 39.2114
R18680 vdd.n2219 vdd.n2218 39.2114
R18681 vdd.n2212 vdd.n2063 39.2114
R18682 vdd.n2211 vdd.n2210 39.2114
R18683 vdd.n2204 vdd.n2065 39.2114
R18684 vdd.n2203 vdd.n2202 39.2114
R18685 vdd.n2196 vdd.n2067 39.2114
R18686 vdd.n2889 vdd.n2888 39.2114
R18687 vdd.n2884 vdd.n2856 39.2114
R18688 vdd.n2882 vdd.n2881 39.2114
R18689 vdd.n2877 vdd.n2859 39.2114
R18690 vdd.n2875 vdd.n2874 39.2114
R18691 vdd.n2870 vdd.n2862 39.2114
R18692 vdd.n2868 vdd.n2867 39.2114
R18693 vdd.n2863 vdd.n755 39.2114
R18694 vdd.n3007 vdd.n3006 39.2114
R18695 vdd.n3004 vdd.n3003 39.2114
R18696 vdd.n2999 vdd.n760 39.2114
R18697 vdd.n2997 vdd.n2996 39.2114
R18698 vdd.n2992 vdd.n763 39.2114
R18699 vdd.n2990 vdd.n2989 39.2114
R18700 vdd.n2985 vdd.n766 39.2114
R18701 vdd.n2983 vdd.n2982 39.2114
R18702 vdd.n2978 vdd.n772 39.2114
R18703 vdd.n2775 vdd.n887 39.2114
R18704 vdd.n2538 vdd.n889 39.2114
R18705 vdd.n2564 vdd.n2539 39.2114
R18706 vdd.n2568 vdd.n2540 39.2114
R18707 vdd.n2572 vdd.n2541 39.2114
R18708 vdd.n2576 vdd.n2542 39.2114
R18709 vdd.n2580 vdd.n2543 39.2114
R18710 vdd.n2584 vdd.n2544 39.2114
R18711 vdd.n2588 vdd.n2545 39.2114
R18712 vdd.n2592 vdd.n2546 39.2114
R18713 vdd.n2596 vdd.n2547 39.2114
R18714 vdd.n2600 vdd.n2548 39.2114
R18715 vdd.n2604 vdd.n2549 39.2114
R18716 vdd.n2608 vdd.n2550 39.2114
R18717 vdd.n2612 vdd.n2551 39.2114
R18718 vdd.n2616 vdd.n2552 39.2114
R18719 vdd.n2620 vdd.n2553 39.2114
R18720 vdd.n2776 vdd.n2775 39.2114
R18721 vdd.n2563 vdd.n2538 39.2114
R18722 vdd.n2567 vdd.n2539 39.2114
R18723 vdd.n2571 vdd.n2540 39.2114
R18724 vdd.n2575 vdd.n2541 39.2114
R18725 vdd.n2579 vdd.n2542 39.2114
R18726 vdd.n2583 vdd.n2543 39.2114
R18727 vdd.n2587 vdd.n2544 39.2114
R18728 vdd.n2591 vdd.n2545 39.2114
R18729 vdd.n2595 vdd.n2546 39.2114
R18730 vdd.n2599 vdd.n2547 39.2114
R18731 vdd.n2603 vdd.n2548 39.2114
R18732 vdd.n2607 vdd.n2549 39.2114
R18733 vdd.n2611 vdd.n2550 39.2114
R18734 vdd.n2615 vdd.n2551 39.2114
R18735 vdd.n2619 vdd.n2552 39.2114
R18736 vdd.n2622 vdd.n2553 39.2114
R18737 vdd.n772 vdd.n767 39.2114
R18738 vdd.n2984 vdd.n2983 39.2114
R18739 vdd.n766 vdd.n764 39.2114
R18740 vdd.n2991 vdd.n2990 39.2114
R18741 vdd.n763 vdd.n761 39.2114
R18742 vdd.n2998 vdd.n2997 39.2114
R18743 vdd.n760 vdd.n758 39.2114
R18744 vdd.n3005 vdd.n3004 39.2114
R18745 vdd.n3008 vdd.n3007 39.2114
R18746 vdd.n2864 vdd.n2863 39.2114
R18747 vdd.n2869 vdd.n2868 39.2114
R18748 vdd.n2862 vdd.n2860 39.2114
R18749 vdd.n2876 vdd.n2875 39.2114
R18750 vdd.n2859 vdd.n2857 39.2114
R18751 vdd.n2883 vdd.n2882 39.2114
R18752 vdd.n2856 vdd.n2854 39.2114
R18753 vdd.n2890 vdd.n2889 39.2114
R18754 vdd.n2028 vdd.n2027 39.2114
R18755 vdd.n2034 vdd.n2033 39.2114
R18756 vdd.n2035 vdd.n2024 39.2114
R18757 vdd.n2042 vdd.n2041 39.2114
R18758 vdd.n2043 vdd.n2022 39.2114
R18759 vdd.n2050 vdd.n2049 39.2114
R18760 vdd.n2051 vdd.n2020 39.2114
R18761 vdd.n2058 vdd.n2057 39.2114
R18762 vdd.n2229 vdd.n2228 39.2114
R18763 vdd.n2226 vdd.n2225 39.2114
R18764 vdd.n2221 vdd.n2220 39.2114
R18765 vdd.n2218 vdd.n2217 39.2114
R18766 vdd.n2213 vdd.n2212 39.2114
R18767 vdd.n2210 vdd.n2209 39.2114
R18768 vdd.n2205 vdd.n2204 39.2114
R18769 vdd.n2202 vdd.n2201 39.2114
R18770 vdd.n2197 vdd.n2196 39.2114
R18771 vdd.n2454 vdd.n908 39.2114
R18772 vdd.n2459 vdd.n909 39.2114
R18773 vdd.n2463 vdd.n910 39.2114
R18774 vdd.n2467 vdd.n911 39.2114
R18775 vdd.n2471 vdd.n912 39.2114
R18776 vdd.n2475 vdd.n913 39.2114
R18777 vdd.n2479 vdd.n914 39.2114
R18778 vdd.n2483 vdd.n915 39.2114
R18779 vdd.n2487 vdd.n916 39.2114
R18780 vdd.n2491 vdd.n917 39.2114
R18781 vdd.n2495 vdd.n918 39.2114
R18782 vdd.n2499 vdd.n919 39.2114
R18783 vdd.n2503 vdd.n920 39.2114
R18784 vdd.n2507 vdd.n921 39.2114
R18785 vdd.n2511 vdd.n922 39.2114
R18786 vdd.n2515 vdd.n923 39.2114
R18787 vdd.n926 vdd.n924 39.2114
R18788 vdd.n2773 vdd.n2772 39.2114
R18789 vdd.n2766 vdd.n2522 39.2114
R18790 vdd.n2762 vdd.n2523 39.2114
R18791 vdd.n2758 vdd.n2524 39.2114
R18792 vdd.n2754 vdd.n2525 39.2114
R18793 vdd.n2750 vdd.n2526 39.2114
R18794 vdd.n2746 vdd.n2527 39.2114
R18795 vdd.n2742 vdd.n2528 39.2114
R18796 vdd.n2738 vdd.n2529 39.2114
R18797 vdd.n2734 vdd.n2530 39.2114
R18798 vdd.n2730 vdd.n2531 39.2114
R18799 vdd.n2726 vdd.n2532 39.2114
R18800 vdd.n2722 vdd.n2533 39.2114
R18801 vdd.n2718 vdd.n2534 39.2114
R18802 vdd.n2714 vdd.n2535 39.2114
R18803 vdd.n2709 vdd.n2536 39.2114
R18804 vdd.n2705 vdd.n2537 39.2114
R18805 vdd.n2911 vdd.n803 39.2114
R18806 vdd.n2918 vdd.n2917 39.2114
R18807 vdd.n802 vdd.n800 39.2114
R18808 vdd.n2925 vdd.n2924 39.2114
R18809 vdd.n799 vdd.n797 39.2114
R18810 vdd.n2932 vdd.n2931 39.2114
R18811 vdd.n796 vdd.n794 39.2114
R18812 vdd.n2939 vdd.n2938 39.2114
R18813 vdd.n793 vdd.n791 39.2114
R18814 vdd.n2947 vdd.n2946 39.2114
R18815 vdd.n790 vdd.n788 39.2114
R18816 vdd.n2954 vdd.n2953 39.2114
R18817 vdd.n787 vdd.n785 39.2114
R18818 vdd.n2961 vdd.n2960 39.2114
R18819 vdd.n784 vdd.n782 39.2114
R18820 vdd.n2968 vdd.n2967 39.2114
R18821 vdd.n2971 vdd.n2970 39.2114
R18822 vdd.n934 vdd.n890 39.2114
R18823 vdd.n2443 vdd.n891 39.2114
R18824 vdd.n2439 vdd.n892 39.2114
R18825 vdd.n2435 vdd.n893 39.2114
R18826 vdd.n2431 vdd.n894 39.2114
R18827 vdd.n2427 vdd.n895 39.2114
R18828 vdd.n2423 vdd.n896 39.2114
R18829 vdd.n2419 vdd.n897 39.2114
R18830 vdd.n2415 vdd.n898 39.2114
R18831 vdd.n2411 vdd.n899 39.2114
R18832 vdd.n2407 vdd.n900 39.2114
R18833 vdd.n2403 vdd.n901 39.2114
R18834 vdd.n2399 vdd.n902 39.2114
R18835 vdd.n2395 vdd.n903 39.2114
R18836 vdd.n2391 vdd.n904 39.2114
R18837 vdd.n2387 vdd.n905 39.2114
R18838 vdd.n2383 vdd.n906 39.2114
R18839 vdd.n2286 vdd.n1023 39.2114
R18840 vdd.n2285 vdd.n2284 39.2114
R18841 vdd.n2278 vdd.n1025 39.2114
R18842 vdd.n2277 vdd.n2276 39.2114
R18843 vdd.n2270 vdd.n1027 39.2114
R18844 vdd.n2269 vdd.n2268 39.2114
R18845 vdd.n2262 vdd.n1029 39.2114
R18846 vdd.n2261 vdd.n2260 39.2114
R18847 vdd.n1032 vdd.n1031 39.2114
R18848 vdd.n2102 vdd.n2101 39.2114
R18849 vdd.n2107 vdd.n2106 39.2114
R18850 vdd.n2110 vdd.n2109 39.2114
R18851 vdd.n2115 vdd.n2114 39.2114
R18852 vdd.n2118 vdd.n2117 39.2114
R18853 vdd.n2123 vdd.n2122 39.2114
R18854 vdd.n2126 vdd.n2125 39.2114
R18855 vdd.n2132 vdd.n2131 39.2114
R18856 vdd.n2380 vdd.n906 39.2114
R18857 vdd.n2384 vdd.n905 39.2114
R18858 vdd.n2388 vdd.n904 39.2114
R18859 vdd.n2392 vdd.n903 39.2114
R18860 vdd.n2396 vdd.n902 39.2114
R18861 vdd.n2400 vdd.n901 39.2114
R18862 vdd.n2404 vdd.n900 39.2114
R18863 vdd.n2408 vdd.n899 39.2114
R18864 vdd.n2412 vdd.n898 39.2114
R18865 vdd.n2416 vdd.n897 39.2114
R18866 vdd.n2420 vdd.n896 39.2114
R18867 vdd.n2424 vdd.n895 39.2114
R18868 vdd.n2428 vdd.n894 39.2114
R18869 vdd.n2432 vdd.n893 39.2114
R18870 vdd.n2436 vdd.n892 39.2114
R18871 vdd.n2440 vdd.n891 39.2114
R18872 vdd.n2444 vdd.n890 39.2114
R18873 vdd.n2287 vdd.n2286 39.2114
R18874 vdd.n2284 vdd.n2283 39.2114
R18875 vdd.n2279 vdd.n2278 39.2114
R18876 vdd.n2276 vdd.n2275 39.2114
R18877 vdd.n2271 vdd.n2270 39.2114
R18878 vdd.n2268 vdd.n2267 39.2114
R18879 vdd.n2263 vdd.n2262 39.2114
R18880 vdd.n2260 vdd.n2259 39.2114
R18881 vdd.n1033 vdd.n1032 39.2114
R18882 vdd.n2103 vdd.n2102 39.2114
R18883 vdd.n2108 vdd.n2107 39.2114
R18884 vdd.n2109 vdd.n2099 39.2114
R18885 vdd.n2116 vdd.n2115 39.2114
R18886 vdd.n2117 vdd.n2097 39.2114
R18887 vdd.n2124 vdd.n2123 39.2114
R18888 vdd.n2125 vdd.n2093 39.2114
R18889 vdd.n2133 vdd.n2132 39.2114
R18890 vdd.n2252 vdd.n2251 37.2369
R18891 vdd.n1955 vdd.n1888 37.2369
R18892 vdd.n1994 vdd.n1848 37.2369
R18893 vdd.n3059 vdd.n724 37.2369
R18894 vdd.n688 vdd.n687 37.2369
R18895 vdd.n3015 vdd.n3014 37.2369
R18896 vdd.n2294 vdd.n1018 31.6883
R18897 vdd.n2519 vdd.n927 31.6883
R18898 vdd.n2452 vdd.n930 31.6883
R18899 vdd.n2198 vdd.n2195 31.6883
R18900 vdd.n2706 vdd.n2704 31.6883
R18901 vdd.n2913 vdd.n2910 31.6883
R18902 vdd.n2783 vdd.n883 31.6883
R18903 vdd.n2974 vdd.n2973 31.6883
R18904 vdd.n2893 vdd.n2892 31.6883
R18905 vdd.n2979 vdd.n771 31.6883
R18906 vdd.n2625 vdd.n2624 31.6883
R18907 vdd.n2779 vdd.n2778 31.6883
R18908 vdd.n2290 vdd.n2289 31.6883
R18909 vdd.n2447 vdd.n2446 31.6883
R18910 vdd.n2379 vdd.n2378 31.6883
R18911 vdd.n2136 vdd.n2135 31.6883
R18912 vdd.n2129 vdd.n2095 30.449
R18913 vdd.n938 vdd.n937 30.449
R18914 vdd.n2070 vdd.n2069 30.449
R18915 vdd.n2457 vdd.n929 30.449
R18916 vdd.n2561 vdd.n2560 30.449
R18917 vdd.n806 vdd.n805 30.449
R18918 vdd.n2711 vdd.n2557 30.449
R18919 vdd.n770 vdd.n769 30.449
R18920 vdd.n1380 vdd.n1146 19.3944
R18921 vdd.n1380 vdd.n1136 19.3944
R18922 vdd.n1392 vdd.n1136 19.3944
R18923 vdd.n1392 vdd.n1134 19.3944
R18924 vdd.n1396 vdd.n1134 19.3944
R18925 vdd.n1396 vdd.n1124 19.3944
R18926 vdd.n1409 vdd.n1124 19.3944
R18927 vdd.n1409 vdd.n1122 19.3944
R18928 vdd.n1413 vdd.n1122 19.3944
R18929 vdd.n1413 vdd.n1114 19.3944
R18930 vdd.n1426 vdd.n1114 19.3944
R18931 vdd.n1426 vdd.n1112 19.3944
R18932 vdd.n1430 vdd.n1112 19.3944
R18933 vdd.n1430 vdd.n1101 19.3944
R18934 vdd.n1442 vdd.n1101 19.3944
R18935 vdd.n1442 vdd.n1099 19.3944
R18936 vdd.n1446 vdd.n1099 19.3944
R18937 vdd.n1446 vdd.n1090 19.3944
R18938 vdd.n1754 vdd.n1090 19.3944
R18939 vdd.n1754 vdd.n1088 19.3944
R18940 vdd.n1758 vdd.n1088 19.3944
R18941 vdd.n1758 vdd.n1079 19.3944
R18942 vdd.n1770 vdd.n1079 19.3944
R18943 vdd.n1770 vdd.n1077 19.3944
R18944 vdd.n1774 vdd.n1077 19.3944
R18945 vdd.n1774 vdd.n1067 19.3944
R18946 vdd.n1787 vdd.n1067 19.3944
R18947 vdd.n1787 vdd.n1065 19.3944
R18948 vdd.n1791 vdd.n1065 19.3944
R18949 vdd.n1791 vdd.n1057 19.3944
R18950 vdd.n1804 vdd.n1057 19.3944
R18951 vdd.n1804 vdd.n1054 19.3944
R18952 vdd.n1810 vdd.n1054 19.3944
R18953 vdd.n1810 vdd.n1055 19.3944
R18954 vdd.n1055 vdd.n1043 19.3944
R18955 vdd.n1299 vdd.n1241 19.3944
R18956 vdd.n1299 vdd.n1298 19.3944
R18957 vdd.n1298 vdd.n1297 19.3944
R18958 vdd.n1297 vdd.n1247 19.3944
R18959 vdd.n1293 vdd.n1247 19.3944
R18960 vdd.n1293 vdd.n1292 19.3944
R18961 vdd.n1292 vdd.n1291 19.3944
R18962 vdd.n1291 vdd.n1253 19.3944
R18963 vdd.n1287 vdd.n1253 19.3944
R18964 vdd.n1287 vdd.n1286 19.3944
R18965 vdd.n1286 vdd.n1285 19.3944
R18966 vdd.n1285 vdd.n1259 19.3944
R18967 vdd.n1281 vdd.n1259 19.3944
R18968 vdd.n1281 vdd.n1280 19.3944
R18969 vdd.n1280 vdd.n1279 19.3944
R18970 vdd.n1279 vdd.n1265 19.3944
R18971 vdd.n1275 vdd.n1265 19.3944
R18972 vdd.n1275 vdd.n1274 19.3944
R18973 vdd.n1274 vdd.n1273 19.3944
R18974 vdd.n1273 vdd.n1271 19.3944
R18975 vdd.n1337 vdd.n1336 19.3944
R18976 vdd.n1336 vdd.n1212 19.3944
R18977 vdd.n1332 vdd.n1212 19.3944
R18978 vdd.n1332 vdd.n1331 19.3944
R18979 vdd.n1331 vdd.n1330 19.3944
R18980 vdd.n1330 vdd.n1218 19.3944
R18981 vdd.n1326 vdd.n1218 19.3944
R18982 vdd.n1326 vdd.n1325 19.3944
R18983 vdd.n1325 vdd.n1324 19.3944
R18984 vdd.n1324 vdd.n1224 19.3944
R18985 vdd.n1320 vdd.n1224 19.3944
R18986 vdd.n1320 vdd.n1319 19.3944
R18987 vdd.n1319 vdd.n1318 19.3944
R18988 vdd.n1318 vdd.n1230 19.3944
R18989 vdd.n1314 vdd.n1230 19.3944
R18990 vdd.n1314 vdd.n1313 19.3944
R18991 vdd.n1313 vdd.n1312 19.3944
R18992 vdd.n1312 vdd.n1236 19.3944
R18993 vdd.n1308 vdd.n1236 19.3944
R18994 vdd.n1308 vdd.n1307 19.3944
R18995 vdd.n1371 vdd.n1370 19.3944
R18996 vdd.n1370 vdd.n1185 19.3944
R18997 vdd.n1366 vdd.n1185 19.3944
R18998 vdd.n1366 vdd.n1365 19.3944
R18999 vdd.n1365 vdd.n1364 19.3944
R19000 vdd.n1364 vdd.n1190 19.3944
R19001 vdd.n1360 vdd.n1190 19.3944
R19002 vdd.n1360 vdd.n1359 19.3944
R19003 vdd.n1359 vdd.n1358 19.3944
R19004 vdd.n1358 vdd.n1196 19.3944
R19005 vdd.n1354 vdd.n1196 19.3944
R19006 vdd.n1354 vdd.n1353 19.3944
R19007 vdd.n1353 vdd.n1352 19.3944
R19008 vdd.n1352 vdd.n1202 19.3944
R19009 vdd.n1348 vdd.n1202 19.3944
R19010 vdd.n1348 vdd.n1347 19.3944
R19011 vdd.n1347 vdd.n1346 19.3944
R19012 vdd.n1346 vdd.n1208 19.3944
R19013 vdd.n1951 vdd.n1886 19.3944
R19014 vdd.n1951 vdd.n1892 19.3944
R19015 vdd.n1946 vdd.n1892 19.3944
R19016 vdd.n1946 vdd.n1945 19.3944
R19017 vdd.n1945 vdd.n1944 19.3944
R19018 vdd.n1944 vdd.n1899 19.3944
R19019 vdd.n1939 vdd.n1899 19.3944
R19020 vdd.n1939 vdd.n1938 19.3944
R19021 vdd.n1938 vdd.n1937 19.3944
R19022 vdd.n1937 vdd.n1906 19.3944
R19023 vdd.n1932 vdd.n1906 19.3944
R19024 vdd.n1932 vdd.n1931 19.3944
R19025 vdd.n1931 vdd.n1930 19.3944
R19026 vdd.n1930 vdd.n1914 19.3944
R19027 vdd.n1925 vdd.n1914 19.3944
R19028 vdd.n1925 vdd.n1924 19.3944
R19029 vdd.n1920 vdd.n1919 19.3944
R19030 vdd.n2253 vdd.n1039 19.3944
R19031 vdd.n1990 vdd.n1846 19.3944
R19032 vdd.n1990 vdd.n1852 19.3944
R19033 vdd.n1985 vdd.n1852 19.3944
R19034 vdd.n1985 vdd.n1984 19.3944
R19035 vdd.n1984 vdd.n1983 19.3944
R19036 vdd.n1983 vdd.n1859 19.3944
R19037 vdd.n1978 vdd.n1859 19.3944
R19038 vdd.n1978 vdd.n1977 19.3944
R19039 vdd.n1977 vdd.n1976 19.3944
R19040 vdd.n1976 vdd.n1866 19.3944
R19041 vdd.n1971 vdd.n1866 19.3944
R19042 vdd.n1971 vdd.n1970 19.3944
R19043 vdd.n1970 vdd.n1969 19.3944
R19044 vdd.n1969 vdd.n1873 19.3944
R19045 vdd.n1964 vdd.n1873 19.3944
R19046 vdd.n1964 vdd.n1963 19.3944
R19047 vdd.n1963 vdd.n1962 19.3944
R19048 vdd.n1962 vdd.n1880 19.3944
R19049 vdd.n1957 vdd.n1880 19.3944
R19050 vdd.n1957 vdd.n1956 19.3944
R19051 vdd.n2241 vdd.n2240 19.3944
R19052 vdd.n2240 vdd.n1818 19.3944
R19053 vdd.n2235 vdd.n2234 19.3944
R19054 vdd.n2017 vdd.n1822 19.3944
R19055 vdd.n2017 vdd.n1824 19.3944
R19056 vdd.n1827 vdd.n1824 19.3944
R19057 vdd.n2010 vdd.n1827 19.3944
R19058 vdd.n2010 vdd.n2009 19.3944
R19059 vdd.n2009 vdd.n2008 19.3944
R19060 vdd.n2008 vdd.n1833 19.3944
R19061 vdd.n2003 vdd.n1833 19.3944
R19062 vdd.n2003 vdd.n2002 19.3944
R19063 vdd.n2002 vdd.n2001 19.3944
R19064 vdd.n2001 vdd.n1840 19.3944
R19065 vdd.n1996 vdd.n1840 19.3944
R19066 vdd.n1996 vdd.n1995 19.3944
R19067 vdd.n1384 vdd.n1142 19.3944
R19068 vdd.n1384 vdd.n1140 19.3944
R19069 vdd.n1388 vdd.n1140 19.3944
R19070 vdd.n1388 vdd.n1130 19.3944
R19071 vdd.n1401 vdd.n1130 19.3944
R19072 vdd.n1401 vdd.n1128 19.3944
R19073 vdd.n1405 vdd.n1128 19.3944
R19074 vdd.n1405 vdd.n1119 19.3944
R19075 vdd.n1418 vdd.n1119 19.3944
R19076 vdd.n1418 vdd.n1117 19.3944
R19077 vdd.n1422 vdd.n1117 19.3944
R19078 vdd.n1422 vdd.n1108 19.3944
R19079 vdd.n1434 vdd.n1108 19.3944
R19080 vdd.n1434 vdd.n1106 19.3944
R19081 vdd.n1438 vdd.n1106 19.3944
R19082 vdd.n1438 vdd.n1096 19.3944
R19083 vdd.n1451 vdd.n1096 19.3944
R19084 vdd.n1451 vdd.n1094 19.3944
R19085 vdd.n1750 vdd.n1094 19.3944
R19086 vdd.n1750 vdd.n1085 19.3944
R19087 vdd.n1762 vdd.n1085 19.3944
R19088 vdd.n1762 vdd.n1083 19.3944
R19089 vdd.n1766 vdd.n1083 19.3944
R19090 vdd.n1766 vdd.n1073 19.3944
R19091 vdd.n1779 vdd.n1073 19.3944
R19092 vdd.n1779 vdd.n1071 19.3944
R19093 vdd.n1783 vdd.n1071 19.3944
R19094 vdd.n1783 vdd.n1062 19.3944
R19095 vdd.n1796 vdd.n1062 19.3944
R19096 vdd.n1796 vdd.n1060 19.3944
R19097 vdd.n1800 vdd.n1060 19.3944
R19098 vdd.n1800 vdd.n1050 19.3944
R19099 vdd.n1814 vdd.n1050 19.3944
R19100 vdd.n1814 vdd.n1048 19.3944
R19101 vdd.n2244 vdd.n1048 19.3944
R19102 vdd.n3147 vdd.n655 19.3944
R19103 vdd.n3151 vdd.n655 19.3944
R19104 vdd.n3151 vdd.n646 19.3944
R19105 vdd.n3163 vdd.n646 19.3944
R19106 vdd.n3163 vdd.n644 19.3944
R19107 vdd.n3167 vdd.n644 19.3944
R19108 vdd.n3167 vdd.n633 19.3944
R19109 vdd.n3179 vdd.n633 19.3944
R19110 vdd.n3179 vdd.n631 19.3944
R19111 vdd.n3183 vdd.n631 19.3944
R19112 vdd.n3183 vdd.n622 19.3944
R19113 vdd.n3196 vdd.n622 19.3944
R19114 vdd.n3196 vdd.n620 19.3944
R19115 vdd.n3203 vdd.n620 19.3944
R19116 vdd.n3203 vdd.n3202 19.3944
R19117 vdd.n3202 vdd.n610 19.3944
R19118 vdd.n3216 vdd.n610 19.3944
R19119 vdd.n3217 vdd.n3216 19.3944
R19120 vdd.n3218 vdd.n3217 19.3944
R19121 vdd.n3218 vdd.n608 19.3944
R19122 vdd.n3223 vdd.n608 19.3944
R19123 vdd.n3224 vdd.n3223 19.3944
R19124 vdd.n3225 vdd.n3224 19.3944
R19125 vdd.n3225 vdd.n606 19.3944
R19126 vdd.n3230 vdd.n606 19.3944
R19127 vdd.n3231 vdd.n3230 19.3944
R19128 vdd.n3232 vdd.n3231 19.3944
R19129 vdd.n3232 vdd.n604 19.3944
R19130 vdd.n3238 vdd.n604 19.3944
R19131 vdd.n3239 vdd.n3238 19.3944
R19132 vdd.n3240 vdd.n3239 19.3944
R19133 vdd.n3240 vdd.n602 19.3944
R19134 vdd.n3245 vdd.n602 19.3944
R19135 vdd.n3246 vdd.n3245 19.3944
R19136 vdd.n3247 vdd.n3246 19.3944
R19137 vdd.n550 vdd.n417 19.3944
R19138 vdd.n556 vdd.n417 19.3944
R19139 vdd.n557 vdd.n556 19.3944
R19140 vdd.n560 vdd.n557 19.3944
R19141 vdd.n560 vdd.n415 19.3944
R19142 vdd.n566 vdd.n415 19.3944
R19143 vdd.n567 vdd.n566 19.3944
R19144 vdd.n570 vdd.n567 19.3944
R19145 vdd.n570 vdd.n413 19.3944
R19146 vdd.n576 vdd.n413 19.3944
R19147 vdd.n577 vdd.n576 19.3944
R19148 vdd.n580 vdd.n577 19.3944
R19149 vdd.n580 vdd.n411 19.3944
R19150 vdd.n586 vdd.n411 19.3944
R19151 vdd.n587 vdd.n586 19.3944
R19152 vdd.n590 vdd.n587 19.3944
R19153 vdd.n590 vdd.n409 19.3944
R19154 vdd.n596 vdd.n409 19.3944
R19155 vdd.n598 vdd.n596 19.3944
R19156 vdd.n599 vdd.n598 19.3944
R19157 vdd.n497 vdd.n496 19.3944
R19158 vdd.n500 vdd.n497 19.3944
R19159 vdd.n500 vdd.n429 19.3944
R19160 vdd.n506 vdd.n429 19.3944
R19161 vdd.n507 vdd.n506 19.3944
R19162 vdd.n510 vdd.n507 19.3944
R19163 vdd.n510 vdd.n427 19.3944
R19164 vdd.n516 vdd.n427 19.3944
R19165 vdd.n517 vdd.n516 19.3944
R19166 vdd.n520 vdd.n517 19.3944
R19167 vdd.n520 vdd.n425 19.3944
R19168 vdd.n526 vdd.n425 19.3944
R19169 vdd.n527 vdd.n526 19.3944
R19170 vdd.n530 vdd.n527 19.3944
R19171 vdd.n530 vdd.n423 19.3944
R19172 vdd.n536 vdd.n423 19.3944
R19173 vdd.n537 vdd.n536 19.3944
R19174 vdd.n540 vdd.n537 19.3944
R19175 vdd.n540 vdd.n421 19.3944
R19176 vdd.n546 vdd.n421 19.3944
R19177 vdd.n447 vdd.n446 19.3944
R19178 vdd.n450 vdd.n447 19.3944
R19179 vdd.n450 vdd.n441 19.3944
R19180 vdd.n456 vdd.n441 19.3944
R19181 vdd.n457 vdd.n456 19.3944
R19182 vdd.n460 vdd.n457 19.3944
R19183 vdd.n460 vdd.n439 19.3944
R19184 vdd.n466 vdd.n439 19.3944
R19185 vdd.n467 vdd.n466 19.3944
R19186 vdd.n470 vdd.n467 19.3944
R19187 vdd.n470 vdd.n437 19.3944
R19188 vdd.n476 vdd.n437 19.3944
R19189 vdd.n477 vdd.n476 19.3944
R19190 vdd.n480 vdd.n477 19.3944
R19191 vdd.n480 vdd.n435 19.3944
R19192 vdd.n486 vdd.n435 19.3944
R19193 vdd.n487 vdd.n486 19.3944
R19194 vdd.n490 vdd.n487 19.3944
R19195 vdd.n3143 vdd.n652 19.3944
R19196 vdd.n3155 vdd.n652 19.3944
R19197 vdd.n3155 vdd.n650 19.3944
R19198 vdd.n3159 vdd.n650 19.3944
R19199 vdd.n3159 vdd.n640 19.3944
R19200 vdd.n3171 vdd.n640 19.3944
R19201 vdd.n3171 vdd.n638 19.3944
R19202 vdd.n3175 vdd.n638 19.3944
R19203 vdd.n3175 vdd.n628 19.3944
R19204 vdd.n3188 vdd.n628 19.3944
R19205 vdd.n3188 vdd.n626 19.3944
R19206 vdd.n3192 vdd.n626 19.3944
R19207 vdd.n3192 vdd.n617 19.3944
R19208 vdd.n3207 vdd.n617 19.3944
R19209 vdd.n3207 vdd.n615 19.3944
R19210 vdd.n3211 vdd.n615 19.3944
R19211 vdd.n3211 vdd.n324 19.3944
R19212 vdd.n3289 vdd.n324 19.3944
R19213 vdd.n3289 vdd.n325 19.3944
R19214 vdd.n3283 vdd.n325 19.3944
R19215 vdd.n3283 vdd.n3282 19.3944
R19216 vdd.n3282 vdd.n3281 19.3944
R19217 vdd.n3281 vdd.n337 19.3944
R19218 vdd.n3275 vdd.n337 19.3944
R19219 vdd.n3275 vdd.n3274 19.3944
R19220 vdd.n3274 vdd.n3273 19.3944
R19221 vdd.n3273 vdd.n347 19.3944
R19222 vdd.n3267 vdd.n347 19.3944
R19223 vdd.n3267 vdd.n3266 19.3944
R19224 vdd.n3266 vdd.n3265 19.3944
R19225 vdd.n3265 vdd.n358 19.3944
R19226 vdd.n3259 vdd.n358 19.3944
R19227 vdd.n3259 vdd.n3258 19.3944
R19228 vdd.n3258 vdd.n3257 19.3944
R19229 vdd.n3257 vdd.n369 19.3944
R19230 vdd.n3100 vdd.n3099 19.3944
R19231 vdd.n3099 vdd.n3098 19.3944
R19232 vdd.n3098 vdd.n694 19.3944
R19233 vdd.n3092 vdd.n694 19.3944
R19234 vdd.n3092 vdd.n3091 19.3944
R19235 vdd.n3091 vdd.n3090 19.3944
R19236 vdd.n3090 vdd.n700 19.3944
R19237 vdd.n3084 vdd.n700 19.3944
R19238 vdd.n3084 vdd.n3083 19.3944
R19239 vdd.n3083 vdd.n3082 19.3944
R19240 vdd.n3082 vdd.n706 19.3944
R19241 vdd.n3076 vdd.n706 19.3944
R19242 vdd.n3076 vdd.n3075 19.3944
R19243 vdd.n3075 vdd.n3074 19.3944
R19244 vdd.n3074 vdd.n712 19.3944
R19245 vdd.n3068 vdd.n712 19.3944
R19246 vdd.n3068 vdd.n3067 19.3944
R19247 vdd.n3067 vdd.n3066 19.3944
R19248 vdd.n3066 vdd.n718 19.3944
R19249 vdd.n3060 vdd.n718 19.3944
R19250 vdd.n3140 vdd.n3139 19.3944
R19251 vdd.n3139 vdd.n662 19.3944
R19252 vdd.n3134 vdd.n3133 19.3944
R19253 vdd.n3130 vdd.n3129 19.3944
R19254 vdd.n3129 vdd.n668 19.3944
R19255 vdd.n3124 vdd.n668 19.3944
R19256 vdd.n3124 vdd.n3123 19.3944
R19257 vdd.n3123 vdd.n3122 19.3944
R19258 vdd.n3122 vdd.n674 19.3944
R19259 vdd.n3116 vdd.n674 19.3944
R19260 vdd.n3116 vdd.n3115 19.3944
R19261 vdd.n3115 vdd.n3114 19.3944
R19262 vdd.n3114 vdd.n680 19.3944
R19263 vdd.n3108 vdd.n680 19.3944
R19264 vdd.n3108 vdd.n3107 19.3944
R19265 vdd.n3107 vdd.n3106 19.3944
R19266 vdd.n3055 vdd.n722 19.3944
R19267 vdd.n3055 vdd.n726 19.3944
R19268 vdd.n3050 vdd.n726 19.3944
R19269 vdd.n3050 vdd.n3049 19.3944
R19270 vdd.n3049 vdd.n732 19.3944
R19271 vdd.n3044 vdd.n732 19.3944
R19272 vdd.n3044 vdd.n3043 19.3944
R19273 vdd.n3043 vdd.n3042 19.3944
R19274 vdd.n3042 vdd.n738 19.3944
R19275 vdd.n3036 vdd.n738 19.3944
R19276 vdd.n3036 vdd.n3035 19.3944
R19277 vdd.n3035 vdd.n3034 19.3944
R19278 vdd.n3034 vdd.n744 19.3944
R19279 vdd.n3028 vdd.n744 19.3944
R19280 vdd.n3028 vdd.n3027 19.3944
R19281 vdd.n3027 vdd.n3026 19.3944
R19282 vdd.n3022 vdd.n3021 19.3944
R19283 vdd.n3018 vdd.n3017 19.3944
R19284 vdd.n1306 vdd.n1241 19.0066
R19285 vdd.n1955 vdd.n1886 19.0066
R19286 vdd.n550 vdd.n547 19.0066
R19287 vdd.n3059 vdd.n722 19.0066
R19288 vdd.n1374 vdd.n1144 18.5924
R19289 vdd.n2246 vdd.n1045 18.5924
R19290 vdd.n3145 vdd.n658 18.5924
R19291 vdd.n3254 vdd.n3253 18.5924
R19292 vdd.n2095 vdd.n2094 16.0975
R19293 vdd.n937 vdd.n936 16.0975
R19294 vdd.n1149 vdd.n1148 16.0975
R19295 vdd.n1305 vdd.n1304 16.0975
R19296 vdd.n1341 vdd.n1340 16.0975
R19297 vdd.n2251 vdd.n2250 16.0975
R19298 vdd.n1888 vdd.n1887 16.0975
R19299 vdd.n1848 vdd.n1847 16.0975
R19300 vdd.n2069 vdd.n2068 16.0975
R19301 vdd.n929 vdd.n928 16.0975
R19302 vdd.n2560 vdd.n2559 16.0975
R19303 vdd.n406 vdd.n405 16.0975
R19304 vdd.n420 vdd.n419 16.0975
R19305 vdd.n432 vdd.n431 16.0975
R19306 vdd.n724 vdd.n723 16.0975
R19307 vdd.n687 vdd.n686 16.0975
R19308 vdd.n805 vdd.n804 16.0975
R19309 vdd.n2557 vdd.n2556 16.0975
R19310 vdd.n3014 vdd.n3013 16.0975
R19311 vdd.n769 vdd.n768 16.0975
R19312 vdd.t248 vdd.n2521 15.4182
R19313 vdd.n2774 vdd.t19 15.4182
R19314 vdd.n28 vdd.n27 14.7125
R19315 vdd.n2292 vdd.n1020 14.5112
R19316 vdd.n2976 vdd.n756 14.5112
R19317 vdd.n316 vdd.n281 13.1884
R19318 vdd.n261 vdd.n226 13.1884
R19319 vdd.n218 vdd.n183 13.1884
R19320 vdd.n163 vdd.n128 13.1884
R19321 vdd.n121 vdd.n86 13.1884
R19322 vdd.n66 vdd.n31 13.1884
R19323 vdd.n1685 vdd.n1650 13.1884
R19324 vdd.n1740 vdd.n1705 13.1884
R19325 vdd.n1587 vdd.n1552 13.1884
R19326 vdd.n1642 vdd.n1607 13.1884
R19327 vdd.n1490 vdd.n1455 13.1884
R19328 vdd.n1545 vdd.n1510 13.1884
R19329 vdd.n1342 vdd.n1337 12.9944
R19330 vdd.n1342 vdd.n1208 12.9944
R19331 vdd.n1994 vdd.n1846 12.9944
R19332 vdd.n1995 vdd.n1994 12.9944
R19333 vdd.n496 vdd.n433 12.9944
R19334 vdd.n490 vdd.n433 12.9944
R19335 vdd.n3100 vdd.n688 12.9944
R19336 vdd.n3106 vdd.n688 12.9944
R19337 vdd.n317 vdd.n279 12.8005
R19338 vdd.n312 vdd.n283 12.8005
R19339 vdd.n262 vdd.n224 12.8005
R19340 vdd.n257 vdd.n228 12.8005
R19341 vdd.n219 vdd.n181 12.8005
R19342 vdd.n214 vdd.n185 12.8005
R19343 vdd.n164 vdd.n126 12.8005
R19344 vdd.n159 vdd.n130 12.8005
R19345 vdd.n122 vdd.n84 12.8005
R19346 vdd.n117 vdd.n88 12.8005
R19347 vdd.n67 vdd.n29 12.8005
R19348 vdd.n62 vdd.n33 12.8005
R19349 vdd.n1686 vdd.n1648 12.8005
R19350 vdd.n1681 vdd.n1652 12.8005
R19351 vdd.n1741 vdd.n1703 12.8005
R19352 vdd.n1736 vdd.n1707 12.8005
R19353 vdd.n1588 vdd.n1550 12.8005
R19354 vdd.n1583 vdd.n1554 12.8005
R19355 vdd.n1643 vdd.n1605 12.8005
R19356 vdd.n1638 vdd.n1609 12.8005
R19357 vdd.n1491 vdd.n1453 12.8005
R19358 vdd.n1486 vdd.n1457 12.8005
R19359 vdd.n1546 vdd.n1508 12.8005
R19360 vdd.n1541 vdd.n1512 12.8005
R19361 vdd.n311 vdd.n284 12.0247
R19362 vdd.n256 vdd.n229 12.0247
R19363 vdd.n213 vdd.n186 12.0247
R19364 vdd.n158 vdd.n131 12.0247
R19365 vdd.n116 vdd.n89 12.0247
R19366 vdd.n61 vdd.n34 12.0247
R19367 vdd.n1680 vdd.n1653 12.0247
R19368 vdd.n1735 vdd.n1708 12.0247
R19369 vdd.n1582 vdd.n1555 12.0247
R19370 vdd.n1637 vdd.n1610 12.0247
R19371 vdd.n1485 vdd.n1458 12.0247
R19372 vdd.n1540 vdd.n1513 12.0247
R19373 vdd.n1382 vdd.n1144 11.337
R19374 vdd.n1390 vdd.n1138 11.337
R19375 vdd.n1390 vdd.n1132 11.337
R19376 vdd.n1399 vdd.n1132 11.337
R19377 vdd.n1407 vdd.n1126 11.337
R19378 vdd.n1416 vdd.n1415 11.337
R19379 vdd.n1432 vdd.n1110 11.337
R19380 vdd.n1440 vdd.n1103 11.337
R19381 vdd.n1449 vdd.n1448 11.337
R19382 vdd.n1752 vdd.n1092 11.337
R19383 vdd.n1768 vdd.n1081 11.337
R19384 vdd.n1777 vdd.n1075 11.337
R19385 vdd.n1785 vdd.n1069 11.337
R19386 vdd.n1794 vdd.n1793 11.337
R19387 vdd.n1802 vdd.n1052 11.337
R19388 vdd.n1812 vdd.n1052 11.337
R19389 vdd.n2246 vdd.n1044 11.337
R19390 vdd.n3145 vdd.n659 11.337
R19391 vdd.n3153 vdd.n648 11.337
R19392 vdd.n3161 vdd.n648 11.337
R19393 vdd.n3169 vdd.n642 11.337
R19394 vdd.n3177 vdd.n635 11.337
R19395 vdd.n3186 vdd.n3185 11.337
R19396 vdd.n3194 vdd.n624 11.337
R19397 vdd.n3213 vdd.n613 11.337
R19398 vdd.n3287 vdd.n328 11.337
R19399 vdd.n3285 vdd.n332 11.337
R19400 vdd.n3279 vdd.n3278 11.337
R19401 vdd.n3271 vdd.n349 11.337
R19402 vdd.n3270 vdd.n3269 11.337
R19403 vdd.n3263 vdd.n3262 11.337
R19404 vdd.n3262 vdd.n3261 11.337
R19405 vdd.n3261 vdd.n363 11.337
R19406 vdd.n3255 vdd.n3254 11.337
R19407 vdd.n308 vdd.n307 11.249
R19408 vdd.n253 vdd.n252 11.249
R19409 vdd.n210 vdd.n209 11.249
R19410 vdd.n155 vdd.n154 11.249
R19411 vdd.n113 vdd.n112 11.249
R19412 vdd.n58 vdd.n57 11.249
R19413 vdd.n1677 vdd.n1676 11.249
R19414 vdd.n1732 vdd.n1731 11.249
R19415 vdd.n1579 vdd.n1578 11.249
R19416 vdd.n1634 vdd.n1633 11.249
R19417 vdd.n1482 vdd.n1481 11.249
R19418 vdd.n1537 vdd.n1536 11.249
R19419 vdd.n2449 vdd.t10 11.1103
R19420 vdd.n2781 vdd.t36 11.1103
R19421 vdd.n1802 vdd.t50 10.7702
R19422 vdd.n3161 vdd.t46 10.7702
R19423 vdd.n293 vdd.n292 10.7238
R19424 vdd.n238 vdd.n237 10.7238
R19425 vdd.n195 vdd.n194 10.7238
R19426 vdd.n140 vdd.n139 10.7238
R19427 vdd.n98 vdd.n97 10.7238
R19428 vdd.n43 vdd.n42 10.7238
R19429 vdd.n1662 vdd.n1661 10.7238
R19430 vdd.n1717 vdd.n1716 10.7238
R19431 vdd.n1564 vdd.n1563 10.7238
R19432 vdd.n1619 vdd.n1618 10.7238
R19433 vdd.n1467 vdd.n1466 10.7238
R19434 vdd.n1522 vdd.n1521 10.7238
R19435 vdd.n2295 vdd.n2294 10.6151
R19436 vdd.n2296 vdd.n2295 10.6151
R19437 vdd.n2296 vdd.n1006 10.6151
R19438 vdd.n2306 vdd.n1006 10.6151
R19439 vdd.n2307 vdd.n2306 10.6151
R19440 vdd.n2308 vdd.n2307 10.6151
R19441 vdd.n2308 vdd.n993 10.6151
R19442 vdd.n2319 vdd.n993 10.6151
R19443 vdd.n2320 vdd.n2319 10.6151
R19444 vdd.n2321 vdd.n2320 10.6151
R19445 vdd.n2321 vdd.n981 10.6151
R19446 vdd.n2331 vdd.n981 10.6151
R19447 vdd.n2332 vdd.n2331 10.6151
R19448 vdd.n2333 vdd.n2332 10.6151
R19449 vdd.n2333 vdd.n969 10.6151
R19450 vdd.n2343 vdd.n969 10.6151
R19451 vdd.n2344 vdd.n2343 10.6151
R19452 vdd.n2345 vdd.n2344 10.6151
R19453 vdd.n2345 vdd.n958 10.6151
R19454 vdd.n2355 vdd.n958 10.6151
R19455 vdd.n2356 vdd.n2355 10.6151
R19456 vdd.n2357 vdd.n2356 10.6151
R19457 vdd.n2357 vdd.n945 10.6151
R19458 vdd.n2369 vdd.n945 10.6151
R19459 vdd.n2370 vdd.n2369 10.6151
R19460 vdd.n2372 vdd.n2370 10.6151
R19461 vdd.n2372 vdd.n2371 10.6151
R19462 vdd.n2371 vdd.n927 10.6151
R19463 vdd.n2519 vdd.n2518 10.6151
R19464 vdd.n2518 vdd.n2517 10.6151
R19465 vdd.n2517 vdd.n2514 10.6151
R19466 vdd.n2514 vdd.n2513 10.6151
R19467 vdd.n2513 vdd.n2510 10.6151
R19468 vdd.n2510 vdd.n2509 10.6151
R19469 vdd.n2509 vdd.n2506 10.6151
R19470 vdd.n2506 vdd.n2505 10.6151
R19471 vdd.n2505 vdd.n2502 10.6151
R19472 vdd.n2502 vdd.n2501 10.6151
R19473 vdd.n2501 vdd.n2498 10.6151
R19474 vdd.n2498 vdd.n2497 10.6151
R19475 vdd.n2497 vdd.n2494 10.6151
R19476 vdd.n2494 vdd.n2493 10.6151
R19477 vdd.n2493 vdd.n2490 10.6151
R19478 vdd.n2490 vdd.n2489 10.6151
R19479 vdd.n2489 vdd.n2486 10.6151
R19480 vdd.n2486 vdd.n2485 10.6151
R19481 vdd.n2485 vdd.n2482 10.6151
R19482 vdd.n2482 vdd.n2481 10.6151
R19483 vdd.n2481 vdd.n2478 10.6151
R19484 vdd.n2478 vdd.n2477 10.6151
R19485 vdd.n2477 vdd.n2474 10.6151
R19486 vdd.n2474 vdd.n2473 10.6151
R19487 vdd.n2473 vdd.n2470 10.6151
R19488 vdd.n2470 vdd.n2469 10.6151
R19489 vdd.n2469 vdd.n2466 10.6151
R19490 vdd.n2466 vdd.n2465 10.6151
R19491 vdd.n2465 vdd.n2462 10.6151
R19492 vdd.n2462 vdd.n2461 10.6151
R19493 vdd.n2461 vdd.n2458 10.6151
R19494 vdd.n2456 vdd.n2453 10.6151
R19495 vdd.n2453 vdd.n2452 10.6151
R19496 vdd.n2195 vdd.n2194 10.6151
R19497 vdd.n2194 vdd.n2192 10.6151
R19498 vdd.n2192 vdd.n2191 10.6151
R19499 vdd.n2191 vdd.n2189 10.6151
R19500 vdd.n2189 vdd.n2188 10.6151
R19501 vdd.n2188 vdd.n2186 10.6151
R19502 vdd.n2186 vdd.n2185 10.6151
R19503 vdd.n2185 vdd.n2183 10.6151
R19504 vdd.n2183 vdd.n2182 10.6151
R19505 vdd.n2182 vdd.n2180 10.6151
R19506 vdd.n2180 vdd.n2179 10.6151
R19507 vdd.n2179 vdd.n2177 10.6151
R19508 vdd.n2177 vdd.n2176 10.6151
R19509 vdd.n2176 vdd.n2091 10.6151
R19510 vdd.n2091 vdd.n2090 10.6151
R19511 vdd.n2090 vdd.n2088 10.6151
R19512 vdd.n2088 vdd.n2087 10.6151
R19513 vdd.n2087 vdd.n2085 10.6151
R19514 vdd.n2085 vdd.n2084 10.6151
R19515 vdd.n2084 vdd.n2082 10.6151
R19516 vdd.n2082 vdd.n2081 10.6151
R19517 vdd.n2081 vdd.n2079 10.6151
R19518 vdd.n2079 vdd.n2078 10.6151
R19519 vdd.n2078 vdd.n2076 10.6151
R19520 vdd.n2076 vdd.n2075 10.6151
R19521 vdd.n2075 vdd.n2072 10.6151
R19522 vdd.n2072 vdd.n2071 10.6151
R19523 vdd.n2071 vdd.n930 10.6151
R19524 vdd.n2029 vdd.n1018 10.6151
R19525 vdd.n2030 vdd.n2029 10.6151
R19526 vdd.n2031 vdd.n2030 10.6151
R19527 vdd.n2031 vdd.n2025 10.6151
R19528 vdd.n2037 vdd.n2025 10.6151
R19529 vdd.n2038 vdd.n2037 10.6151
R19530 vdd.n2039 vdd.n2038 10.6151
R19531 vdd.n2039 vdd.n2023 10.6151
R19532 vdd.n2045 vdd.n2023 10.6151
R19533 vdd.n2046 vdd.n2045 10.6151
R19534 vdd.n2047 vdd.n2046 10.6151
R19535 vdd.n2047 vdd.n2021 10.6151
R19536 vdd.n2053 vdd.n2021 10.6151
R19537 vdd.n2054 vdd.n2053 10.6151
R19538 vdd.n2055 vdd.n2054 10.6151
R19539 vdd.n2055 vdd.n2019 10.6151
R19540 vdd.n2231 vdd.n2019 10.6151
R19541 vdd.n2231 vdd.n2230 10.6151
R19542 vdd.n2230 vdd.n2060 10.6151
R19543 vdd.n2224 vdd.n2060 10.6151
R19544 vdd.n2224 vdd.n2223 10.6151
R19545 vdd.n2223 vdd.n2222 10.6151
R19546 vdd.n2222 vdd.n2062 10.6151
R19547 vdd.n2216 vdd.n2062 10.6151
R19548 vdd.n2216 vdd.n2215 10.6151
R19549 vdd.n2215 vdd.n2214 10.6151
R19550 vdd.n2214 vdd.n2064 10.6151
R19551 vdd.n2208 vdd.n2064 10.6151
R19552 vdd.n2208 vdd.n2207 10.6151
R19553 vdd.n2207 vdd.n2206 10.6151
R19554 vdd.n2206 vdd.n2066 10.6151
R19555 vdd.n2200 vdd.n2199 10.6151
R19556 vdd.n2199 vdd.n2198 10.6151
R19557 vdd.n2704 vdd.n2703 10.6151
R19558 vdd.n2703 vdd.n2701 10.6151
R19559 vdd.n2701 vdd.n2700 10.6151
R19560 vdd.n2700 vdd.n2558 10.6151
R19561 vdd.n2647 vdd.n2558 10.6151
R19562 vdd.n2648 vdd.n2647 10.6151
R19563 vdd.n2650 vdd.n2648 10.6151
R19564 vdd.n2651 vdd.n2650 10.6151
R19565 vdd.n2653 vdd.n2651 10.6151
R19566 vdd.n2654 vdd.n2653 10.6151
R19567 vdd.n2656 vdd.n2654 10.6151
R19568 vdd.n2657 vdd.n2656 10.6151
R19569 vdd.n2659 vdd.n2657 10.6151
R19570 vdd.n2660 vdd.n2659 10.6151
R19571 vdd.n2675 vdd.n2660 10.6151
R19572 vdd.n2675 vdd.n2674 10.6151
R19573 vdd.n2674 vdd.n2673 10.6151
R19574 vdd.n2673 vdd.n2671 10.6151
R19575 vdd.n2671 vdd.n2670 10.6151
R19576 vdd.n2670 vdd.n2668 10.6151
R19577 vdd.n2668 vdd.n2667 10.6151
R19578 vdd.n2667 vdd.n2665 10.6151
R19579 vdd.n2665 vdd.n2664 10.6151
R19580 vdd.n2664 vdd.n2662 10.6151
R19581 vdd.n2662 vdd.n2661 10.6151
R19582 vdd.n2661 vdd.n807 10.6151
R19583 vdd.n2909 vdd.n807 10.6151
R19584 vdd.n2910 vdd.n2909 10.6151
R19585 vdd.n2771 vdd.n883 10.6151
R19586 vdd.n2771 vdd.n2770 10.6151
R19587 vdd.n2770 vdd.n2769 10.6151
R19588 vdd.n2769 vdd.n2767 10.6151
R19589 vdd.n2767 vdd.n2764 10.6151
R19590 vdd.n2764 vdd.n2763 10.6151
R19591 vdd.n2763 vdd.n2760 10.6151
R19592 vdd.n2760 vdd.n2759 10.6151
R19593 vdd.n2759 vdd.n2756 10.6151
R19594 vdd.n2756 vdd.n2755 10.6151
R19595 vdd.n2755 vdd.n2752 10.6151
R19596 vdd.n2752 vdd.n2751 10.6151
R19597 vdd.n2751 vdd.n2748 10.6151
R19598 vdd.n2748 vdd.n2747 10.6151
R19599 vdd.n2747 vdd.n2744 10.6151
R19600 vdd.n2744 vdd.n2743 10.6151
R19601 vdd.n2743 vdd.n2740 10.6151
R19602 vdd.n2740 vdd.n2739 10.6151
R19603 vdd.n2739 vdd.n2736 10.6151
R19604 vdd.n2736 vdd.n2735 10.6151
R19605 vdd.n2735 vdd.n2732 10.6151
R19606 vdd.n2732 vdd.n2731 10.6151
R19607 vdd.n2731 vdd.n2728 10.6151
R19608 vdd.n2728 vdd.n2727 10.6151
R19609 vdd.n2727 vdd.n2724 10.6151
R19610 vdd.n2724 vdd.n2723 10.6151
R19611 vdd.n2723 vdd.n2720 10.6151
R19612 vdd.n2720 vdd.n2719 10.6151
R19613 vdd.n2719 vdd.n2716 10.6151
R19614 vdd.n2716 vdd.n2715 10.6151
R19615 vdd.n2715 vdd.n2712 10.6151
R19616 vdd.n2710 vdd.n2707 10.6151
R19617 vdd.n2707 vdd.n2706 10.6151
R19618 vdd.n2784 vdd.n2783 10.6151
R19619 vdd.n2785 vdd.n2784 10.6151
R19620 vdd.n2785 vdd.n873 10.6151
R19621 vdd.n2795 vdd.n873 10.6151
R19622 vdd.n2796 vdd.n2795 10.6151
R19623 vdd.n2797 vdd.n2796 10.6151
R19624 vdd.n2797 vdd.n860 10.6151
R19625 vdd.n2807 vdd.n860 10.6151
R19626 vdd.n2808 vdd.n2807 10.6151
R19627 vdd.n2809 vdd.n2808 10.6151
R19628 vdd.n2809 vdd.n849 10.6151
R19629 vdd.n2819 vdd.n849 10.6151
R19630 vdd.n2820 vdd.n2819 10.6151
R19631 vdd.n2821 vdd.n2820 10.6151
R19632 vdd.n2821 vdd.n837 10.6151
R19633 vdd.n2831 vdd.n837 10.6151
R19634 vdd.n2832 vdd.n2831 10.6151
R19635 vdd.n2833 vdd.n2832 10.6151
R19636 vdd.n2833 vdd.n826 10.6151
R19637 vdd.n2845 vdd.n826 10.6151
R19638 vdd.n2846 vdd.n2845 10.6151
R19639 vdd.n2847 vdd.n2846 10.6151
R19640 vdd.n2847 vdd.n812 10.6151
R19641 vdd.n2902 vdd.n812 10.6151
R19642 vdd.n2903 vdd.n2902 10.6151
R19643 vdd.n2904 vdd.n2903 10.6151
R19644 vdd.n2904 vdd.n779 10.6151
R19645 vdd.n2974 vdd.n779 10.6151
R19646 vdd.n2973 vdd.n2972 10.6151
R19647 vdd.n2972 vdd.n780 10.6151
R19648 vdd.n781 vdd.n780 10.6151
R19649 vdd.n2965 vdd.n781 10.6151
R19650 vdd.n2965 vdd.n2964 10.6151
R19651 vdd.n2964 vdd.n2963 10.6151
R19652 vdd.n2963 vdd.n783 10.6151
R19653 vdd.n2958 vdd.n783 10.6151
R19654 vdd.n2958 vdd.n2957 10.6151
R19655 vdd.n2957 vdd.n2956 10.6151
R19656 vdd.n2956 vdd.n786 10.6151
R19657 vdd.n2951 vdd.n786 10.6151
R19658 vdd.n2951 vdd.n2950 10.6151
R19659 vdd.n2950 vdd.n2949 10.6151
R19660 vdd.n2949 vdd.n789 10.6151
R19661 vdd.n2944 vdd.n789 10.6151
R19662 vdd.n2944 vdd.n2943 10.6151
R19663 vdd.n2943 vdd.n2941 10.6151
R19664 vdd.n2941 vdd.n792 10.6151
R19665 vdd.n2936 vdd.n792 10.6151
R19666 vdd.n2936 vdd.n2935 10.6151
R19667 vdd.n2935 vdd.n2934 10.6151
R19668 vdd.n2934 vdd.n795 10.6151
R19669 vdd.n2929 vdd.n795 10.6151
R19670 vdd.n2929 vdd.n2928 10.6151
R19671 vdd.n2928 vdd.n2927 10.6151
R19672 vdd.n2927 vdd.n798 10.6151
R19673 vdd.n2922 vdd.n798 10.6151
R19674 vdd.n2922 vdd.n2921 10.6151
R19675 vdd.n2921 vdd.n2920 10.6151
R19676 vdd.n2920 vdd.n801 10.6151
R19677 vdd.n2915 vdd.n2914 10.6151
R19678 vdd.n2914 vdd.n2913 10.6151
R19679 vdd.n2892 vdd.n2853 10.6151
R19680 vdd.n2887 vdd.n2853 10.6151
R19681 vdd.n2887 vdd.n2886 10.6151
R19682 vdd.n2886 vdd.n2885 10.6151
R19683 vdd.n2885 vdd.n2855 10.6151
R19684 vdd.n2880 vdd.n2855 10.6151
R19685 vdd.n2880 vdd.n2879 10.6151
R19686 vdd.n2879 vdd.n2878 10.6151
R19687 vdd.n2878 vdd.n2858 10.6151
R19688 vdd.n2873 vdd.n2858 10.6151
R19689 vdd.n2873 vdd.n2872 10.6151
R19690 vdd.n2872 vdd.n2871 10.6151
R19691 vdd.n2871 vdd.n2861 10.6151
R19692 vdd.n2866 vdd.n2861 10.6151
R19693 vdd.n2866 vdd.n2865 10.6151
R19694 vdd.n2865 vdd.n753 10.6151
R19695 vdd.n3009 vdd.n753 10.6151
R19696 vdd.n3009 vdd.n754 10.6151
R19697 vdd.n757 vdd.n754 10.6151
R19698 vdd.n3002 vdd.n757 10.6151
R19699 vdd.n3002 vdd.n3001 10.6151
R19700 vdd.n3001 vdd.n3000 10.6151
R19701 vdd.n3000 vdd.n759 10.6151
R19702 vdd.n2995 vdd.n759 10.6151
R19703 vdd.n2995 vdd.n2994 10.6151
R19704 vdd.n2994 vdd.n2993 10.6151
R19705 vdd.n2993 vdd.n762 10.6151
R19706 vdd.n2988 vdd.n762 10.6151
R19707 vdd.n2988 vdd.n2987 10.6151
R19708 vdd.n2987 vdd.n2986 10.6151
R19709 vdd.n2986 vdd.n765 10.6151
R19710 vdd.n2981 vdd.n2980 10.6151
R19711 vdd.n2980 vdd.n2979 10.6151
R19712 vdd.n2627 vdd.n2625 10.6151
R19713 vdd.n2628 vdd.n2627 10.6151
R19714 vdd.n2696 vdd.n2628 10.6151
R19715 vdd.n2696 vdd.n2695 10.6151
R19716 vdd.n2695 vdd.n2694 10.6151
R19717 vdd.n2694 vdd.n2692 10.6151
R19718 vdd.n2692 vdd.n2691 10.6151
R19719 vdd.n2691 vdd.n2689 10.6151
R19720 vdd.n2689 vdd.n2688 10.6151
R19721 vdd.n2688 vdd.n2686 10.6151
R19722 vdd.n2686 vdd.n2685 10.6151
R19723 vdd.n2685 vdd.n2683 10.6151
R19724 vdd.n2683 vdd.n2682 10.6151
R19725 vdd.n2682 vdd.n2680 10.6151
R19726 vdd.n2680 vdd.n2679 10.6151
R19727 vdd.n2679 vdd.n2645 10.6151
R19728 vdd.n2645 vdd.n2644 10.6151
R19729 vdd.n2644 vdd.n2642 10.6151
R19730 vdd.n2642 vdd.n2641 10.6151
R19731 vdd.n2641 vdd.n2639 10.6151
R19732 vdd.n2639 vdd.n2638 10.6151
R19733 vdd.n2638 vdd.n2636 10.6151
R19734 vdd.n2636 vdd.n2635 10.6151
R19735 vdd.n2635 vdd.n2633 10.6151
R19736 vdd.n2633 vdd.n2632 10.6151
R19737 vdd.n2632 vdd.n2630 10.6151
R19738 vdd.n2630 vdd.n2629 10.6151
R19739 vdd.n2629 vdd.n771 10.6151
R19740 vdd.n2778 vdd.n2777 10.6151
R19741 vdd.n2777 vdd.n888 10.6151
R19742 vdd.n2562 vdd.n888 10.6151
R19743 vdd.n2565 vdd.n2562 10.6151
R19744 vdd.n2566 vdd.n2565 10.6151
R19745 vdd.n2569 vdd.n2566 10.6151
R19746 vdd.n2570 vdd.n2569 10.6151
R19747 vdd.n2573 vdd.n2570 10.6151
R19748 vdd.n2574 vdd.n2573 10.6151
R19749 vdd.n2577 vdd.n2574 10.6151
R19750 vdd.n2578 vdd.n2577 10.6151
R19751 vdd.n2581 vdd.n2578 10.6151
R19752 vdd.n2582 vdd.n2581 10.6151
R19753 vdd.n2585 vdd.n2582 10.6151
R19754 vdd.n2586 vdd.n2585 10.6151
R19755 vdd.n2589 vdd.n2586 10.6151
R19756 vdd.n2590 vdd.n2589 10.6151
R19757 vdd.n2593 vdd.n2590 10.6151
R19758 vdd.n2594 vdd.n2593 10.6151
R19759 vdd.n2597 vdd.n2594 10.6151
R19760 vdd.n2598 vdd.n2597 10.6151
R19761 vdd.n2601 vdd.n2598 10.6151
R19762 vdd.n2602 vdd.n2601 10.6151
R19763 vdd.n2605 vdd.n2602 10.6151
R19764 vdd.n2606 vdd.n2605 10.6151
R19765 vdd.n2609 vdd.n2606 10.6151
R19766 vdd.n2610 vdd.n2609 10.6151
R19767 vdd.n2613 vdd.n2610 10.6151
R19768 vdd.n2614 vdd.n2613 10.6151
R19769 vdd.n2617 vdd.n2614 10.6151
R19770 vdd.n2618 vdd.n2617 10.6151
R19771 vdd.n2623 vdd.n2621 10.6151
R19772 vdd.n2624 vdd.n2623 10.6151
R19773 vdd.n2779 vdd.n878 10.6151
R19774 vdd.n2789 vdd.n878 10.6151
R19775 vdd.n2790 vdd.n2789 10.6151
R19776 vdd.n2791 vdd.n2790 10.6151
R19777 vdd.n2791 vdd.n866 10.6151
R19778 vdd.n2801 vdd.n866 10.6151
R19779 vdd.n2802 vdd.n2801 10.6151
R19780 vdd.n2803 vdd.n2802 10.6151
R19781 vdd.n2803 vdd.n855 10.6151
R19782 vdd.n2813 vdd.n855 10.6151
R19783 vdd.n2814 vdd.n2813 10.6151
R19784 vdd.n2815 vdd.n2814 10.6151
R19785 vdd.n2815 vdd.n843 10.6151
R19786 vdd.n2825 vdd.n843 10.6151
R19787 vdd.n2826 vdd.n2825 10.6151
R19788 vdd.n2827 vdd.n2826 10.6151
R19789 vdd.n2827 vdd.n832 10.6151
R19790 vdd.n2837 vdd.n832 10.6151
R19791 vdd.n2838 vdd.n2837 10.6151
R19792 vdd.n2841 vdd.n2838 10.6151
R19793 vdd.n2851 vdd.n820 10.6151
R19794 vdd.n2852 vdd.n2851 10.6151
R19795 vdd.n2898 vdd.n2852 10.6151
R19796 vdd.n2898 vdd.n2897 10.6151
R19797 vdd.n2897 vdd.n2896 10.6151
R19798 vdd.n2896 vdd.n2895 10.6151
R19799 vdd.n2895 vdd.n2893 10.6151
R19800 vdd.n2290 vdd.n1012 10.6151
R19801 vdd.n2300 vdd.n1012 10.6151
R19802 vdd.n2301 vdd.n2300 10.6151
R19803 vdd.n2302 vdd.n2301 10.6151
R19804 vdd.n2302 vdd.n999 10.6151
R19805 vdd.n2312 vdd.n999 10.6151
R19806 vdd.n2313 vdd.n2312 10.6151
R19807 vdd.n2315 vdd.n987 10.6151
R19808 vdd.n2325 vdd.n987 10.6151
R19809 vdd.n2326 vdd.n2325 10.6151
R19810 vdd.n2327 vdd.n2326 10.6151
R19811 vdd.n2327 vdd.n975 10.6151
R19812 vdd.n2337 vdd.n975 10.6151
R19813 vdd.n2338 vdd.n2337 10.6151
R19814 vdd.n2339 vdd.n2338 10.6151
R19815 vdd.n2339 vdd.n964 10.6151
R19816 vdd.n2349 vdd.n964 10.6151
R19817 vdd.n2350 vdd.n2349 10.6151
R19818 vdd.n2351 vdd.n2350 10.6151
R19819 vdd.n2351 vdd.n952 10.6151
R19820 vdd.n2361 vdd.n952 10.6151
R19821 vdd.n2362 vdd.n2361 10.6151
R19822 vdd.n2365 vdd.n2362 10.6151
R19823 vdd.n2365 vdd.n2364 10.6151
R19824 vdd.n2364 vdd.n2363 10.6151
R19825 vdd.n2363 vdd.n935 10.6151
R19826 vdd.n2447 vdd.n935 10.6151
R19827 vdd.n2446 vdd.n2445 10.6151
R19828 vdd.n2445 vdd.n2442 10.6151
R19829 vdd.n2442 vdd.n2441 10.6151
R19830 vdd.n2441 vdd.n2438 10.6151
R19831 vdd.n2438 vdd.n2437 10.6151
R19832 vdd.n2437 vdd.n2434 10.6151
R19833 vdd.n2434 vdd.n2433 10.6151
R19834 vdd.n2433 vdd.n2430 10.6151
R19835 vdd.n2430 vdd.n2429 10.6151
R19836 vdd.n2429 vdd.n2426 10.6151
R19837 vdd.n2426 vdd.n2425 10.6151
R19838 vdd.n2425 vdd.n2422 10.6151
R19839 vdd.n2422 vdd.n2421 10.6151
R19840 vdd.n2421 vdd.n2418 10.6151
R19841 vdd.n2418 vdd.n2417 10.6151
R19842 vdd.n2417 vdd.n2414 10.6151
R19843 vdd.n2414 vdd.n2413 10.6151
R19844 vdd.n2413 vdd.n2410 10.6151
R19845 vdd.n2410 vdd.n2409 10.6151
R19846 vdd.n2409 vdd.n2406 10.6151
R19847 vdd.n2406 vdd.n2405 10.6151
R19848 vdd.n2405 vdd.n2402 10.6151
R19849 vdd.n2402 vdd.n2401 10.6151
R19850 vdd.n2401 vdd.n2398 10.6151
R19851 vdd.n2398 vdd.n2397 10.6151
R19852 vdd.n2397 vdd.n2394 10.6151
R19853 vdd.n2394 vdd.n2393 10.6151
R19854 vdd.n2393 vdd.n2390 10.6151
R19855 vdd.n2390 vdd.n2389 10.6151
R19856 vdd.n2389 vdd.n2386 10.6151
R19857 vdd.n2386 vdd.n2385 10.6151
R19858 vdd.n2382 vdd.n2381 10.6151
R19859 vdd.n2381 vdd.n2379 10.6151
R19860 vdd.n2138 vdd.n2136 10.6151
R19861 vdd.n2139 vdd.n2138 10.6151
R19862 vdd.n2141 vdd.n2139 10.6151
R19863 vdd.n2142 vdd.n2141 10.6151
R19864 vdd.n2144 vdd.n2142 10.6151
R19865 vdd.n2145 vdd.n2144 10.6151
R19866 vdd.n2147 vdd.n2145 10.6151
R19867 vdd.n2148 vdd.n2147 10.6151
R19868 vdd.n2150 vdd.n2148 10.6151
R19869 vdd.n2151 vdd.n2150 10.6151
R19870 vdd.n2153 vdd.n2151 10.6151
R19871 vdd.n2154 vdd.n2153 10.6151
R19872 vdd.n2172 vdd.n2154 10.6151
R19873 vdd.n2172 vdd.n2171 10.6151
R19874 vdd.n2171 vdd.n2170 10.6151
R19875 vdd.n2170 vdd.n2168 10.6151
R19876 vdd.n2168 vdd.n2167 10.6151
R19877 vdd.n2167 vdd.n2165 10.6151
R19878 vdd.n2165 vdd.n2164 10.6151
R19879 vdd.n2164 vdd.n2162 10.6151
R19880 vdd.n2162 vdd.n2161 10.6151
R19881 vdd.n2161 vdd.n2159 10.6151
R19882 vdd.n2159 vdd.n2158 10.6151
R19883 vdd.n2158 vdd.n2156 10.6151
R19884 vdd.n2156 vdd.n2155 10.6151
R19885 vdd.n2155 vdd.n939 10.6151
R19886 vdd.n2377 vdd.n939 10.6151
R19887 vdd.n2378 vdd.n2377 10.6151
R19888 vdd.n2289 vdd.n2288 10.6151
R19889 vdd.n2288 vdd.n1024 10.6151
R19890 vdd.n2282 vdd.n1024 10.6151
R19891 vdd.n2282 vdd.n2281 10.6151
R19892 vdd.n2281 vdd.n2280 10.6151
R19893 vdd.n2280 vdd.n1026 10.6151
R19894 vdd.n2274 vdd.n1026 10.6151
R19895 vdd.n2274 vdd.n2273 10.6151
R19896 vdd.n2273 vdd.n2272 10.6151
R19897 vdd.n2272 vdd.n1028 10.6151
R19898 vdd.n2266 vdd.n1028 10.6151
R19899 vdd.n2266 vdd.n2265 10.6151
R19900 vdd.n2265 vdd.n2264 10.6151
R19901 vdd.n2264 vdd.n1030 10.6151
R19902 vdd.n2258 vdd.n1030 10.6151
R19903 vdd.n2258 vdd.n2257 10.6151
R19904 vdd.n2257 vdd.n2256 10.6151
R19905 vdd.n2256 vdd.n1034 10.6151
R19906 vdd.n2104 vdd.n1034 10.6151
R19907 vdd.n2105 vdd.n2104 10.6151
R19908 vdd.n2105 vdd.n2100 10.6151
R19909 vdd.n2111 vdd.n2100 10.6151
R19910 vdd.n2112 vdd.n2111 10.6151
R19911 vdd.n2113 vdd.n2112 10.6151
R19912 vdd.n2113 vdd.n2098 10.6151
R19913 vdd.n2119 vdd.n2098 10.6151
R19914 vdd.n2120 vdd.n2119 10.6151
R19915 vdd.n2121 vdd.n2120 10.6151
R19916 vdd.n2121 vdd.n2096 10.6151
R19917 vdd.n2127 vdd.n2096 10.6151
R19918 vdd.n2128 vdd.n2127 10.6151
R19919 vdd.n2130 vdd.n2092 10.6151
R19920 vdd.n2135 vdd.n2092 10.6151
R19921 vdd.t134 vdd.n1776 10.5435
R19922 vdd.n636 vdd.t52 10.5435
R19923 vdd.n304 vdd.n286 10.4732
R19924 vdd.n249 vdd.n231 10.4732
R19925 vdd.n206 vdd.n188 10.4732
R19926 vdd.n151 vdd.n133 10.4732
R19927 vdd.n109 vdd.n91 10.4732
R19928 vdd.n54 vdd.n36 10.4732
R19929 vdd.n1673 vdd.n1655 10.4732
R19930 vdd.n1728 vdd.n1710 10.4732
R19931 vdd.n1575 vdd.n1557 10.4732
R19932 vdd.n1630 vdd.n1612 10.4732
R19933 vdd.n1478 vdd.n1460 10.4732
R19934 vdd.n1533 vdd.n1515 10.4732
R19935 vdd.n1760 vdd.t102 10.3167
R19936 vdd.n3205 vdd.t44 10.3167
R19937 vdd.t58 vdd.n1104 10.09
R19938 vdd.n1812 vdd.t192 10.09
R19939 vdd.n3153 vdd.t177 10.09
R19940 vdd.n3286 vdd.t54 10.09
R19941 vdd.n1424 vdd.t76 9.86327
R19942 vdd.n3277 vdd.t110 9.86327
R19943 vdd.n303 vdd.n288 9.69747
R19944 vdd.n248 vdd.n233 9.69747
R19945 vdd.n205 vdd.n190 9.69747
R19946 vdd.n150 vdd.n135 9.69747
R19947 vdd.n108 vdd.n93 9.69747
R19948 vdd.n53 vdd.n38 9.69747
R19949 vdd.n1672 vdd.n1657 9.69747
R19950 vdd.n1727 vdd.n1712 9.69747
R19951 vdd.n1574 vdd.n1559 9.69747
R19952 vdd.n1629 vdd.n1614 9.69747
R19953 vdd.n1477 vdd.n1462 9.69747
R19954 vdd.n1532 vdd.n1517 9.69747
R19955 vdd.n2232 vdd.n2231 9.67831
R19956 vdd.n2943 vdd.n2942 9.67831
R19957 vdd.n3010 vdd.n3009 9.67831
R19958 vdd.n2256 vdd.n2255 9.67831
R19959 vdd.t56 vdd.n1398 9.63654
R19960 vdd.n3236 vdd.t69 9.63654
R19961 vdd.n319 vdd.n318 9.45567
R19962 vdd.n264 vdd.n263 9.45567
R19963 vdd.n221 vdd.n220 9.45567
R19964 vdd.n166 vdd.n165 9.45567
R19965 vdd.n124 vdd.n123 9.45567
R19966 vdd.n69 vdd.n68 9.45567
R19967 vdd.n1688 vdd.n1687 9.45567
R19968 vdd.n1743 vdd.n1742 9.45567
R19969 vdd.n1590 vdd.n1589 9.45567
R19970 vdd.n1645 vdd.n1644 9.45567
R19971 vdd.n1493 vdd.n1492 9.45567
R19972 vdd.n1548 vdd.n1547 9.45567
R19973 vdd.n1992 vdd.n1846 9.3005
R19974 vdd.n1991 vdd.n1990 9.3005
R19975 vdd.n1852 vdd.n1851 9.3005
R19976 vdd.n1985 vdd.n1856 9.3005
R19977 vdd.n1984 vdd.n1857 9.3005
R19978 vdd.n1983 vdd.n1858 9.3005
R19979 vdd.n1862 vdd.n1859 9.3005
R19980 vdd.n1978 vdd.n1863 9.3005
R19981 vdd.n1977 vdd.n1864 9.3005
R19982 vdd.n1976 vdd.n1865 9.3005
R19983 vdd.n1869 vdd.n1866 9.3005
R19984 vdd.n1971 vdd.n1870 9.3005
R19985 vdd.n1970 vdd.n1871 9.3005
R19986 vdd.n1969 vdd.n1872 9.3005
R19987 vdd.n1876 vdd.n1873 9.3005
R19988 vdd.n1964 vdd.n1877 9.3005
R19989 vdd.n1963 vdd.n1878 9.3005
R19990 vdd.n1962 vdd.n1879 9.3005
R19991 vdd.n1883 vdd.n1880 9.3005
R19992 vdd.n1957 vdd.n1884 9.3005
R19993 vdd.n1956 vdd.n1885 9.3005
R19994 vdd.n1955 vdd.n1954 9.3005
R19995 vdd.n1953 vdd.n1886 9.3005
R19996 vdd.n1952 vdd.n1951 9.3005
R19997 vdd.n1892 vdd.n1891 9.3005
R19998 vdd.n1946 vdd.n1896 9.3005
R19999 vdd.n1945 vdd.n1897 9.3005
R20000 vdd.n1944 vdd.n1898 9.3005
R20001 vdd.n1902 vdd.n1899 9.3005
R20002 vdd.n1939 vdd.n1903 9.3005
R20003 vdd.n1938 vdd.n1904 9.3005
R20004 vdd.n1937 vdd.n1905 9.3005
R20005 vdd.n1909 vdd.n1906 9.3005
R20006 vdd.n1932 vdd.n1910 9.3005
R20007 vdd.n1931 vdd.n1911 9.3005
R20008 vdd.n1930 vdd.n1912 9.3005
R20009 vdd.n1914 vdd.n1913 9.3005
R20010 vdd.n1925 vdd.n1035 9.3005
R20011 vdd.n1994 vdd.n1993 9.3005
R20012 vdd.n2018 vdd.n2017 9.3005
R20013 vdd.n1824 vdd.n1823 9.3005
R20014 vdd.n1829 vdd.n1827 9.3005
R20015 vdd.n2010 vdd.n1830 9.3005
R20016 vdd.n2009 vdd.n1831 9.3005
R20017 vdd.n2008 vdd.n1832 9.3005
R20018 vdd.n1836 vdd.n1833 9.3005
R20019 vdd.n2003 vdd.n1837 9.3005
R20020 vdd.n2002 vdd.n1838 9.3005
R20021 vdd.n2001 vdd.n1839 9.3005
R20022 vdd.n1843 vdd.n1840 9.3005
R20023 vdd.n1996 vdd.n1844 9.3005
R20024 vdd.n1995 vdd.n1845 9.3005
R20025 vdd.n2240 vdd.n1817 9.3005
R20026 vdd.n2242 vdd.n2241 9.3005
R20027 vdd.n1748 vdd.n1094 9.3005
R20028 vdd.n1750 vdd.n1749 9.3005
R20029 vdd.n1085 vdd.n1084 9.3005
R20030 vdd.n1763 vdd.n1762 9.3005
R20031 vdd.n1764 vdd.n1083 9.3005
R20032 vdd.n1766 vdd.n1765 9.3005
R20033 vdd.n1073 vdd.n1072 9.3005
R20034 vdd.n1780 vdd.n1779 9.3005
R20035 vdd.n1781 vdd.n1071 9.3005
R20036 vdd.n1783 vdd.n1782 9.3005
R20037 vdd.n1062 vdd.n1061 9.3005
R20038 vdd.n1797 vdd.n1796 9.3005
R20039 vdd.n1798 vdd.n1060 9.3005
R20040 vdd.n1800 vdd.n1799 9.3005
R20041 vdd.n1050 vdd.n1049 9.3005
R20042 vdd.n1815 vdd.n1814 9.3005
R20043 vdd.n1816 vdd.n1048 9.3005
R20044 vdd.n2244 vdd.n2243 9.3005
R20045 vdd.n295 vdd.n294 9.3005
R20046 vdd.n290 vdd.n289 9.3005
R20047 vdd.n301 vdd.n300 9.3005
R20048 vdd.n303 vdd.n302 9.3005
R20049 vdd.n286 vdd.n285 9.3005
R20050 vdd.n309 vdd.n308 9.3005
R20051 vdd.n311 vdd.n310 9.3005
R20052 vdd.n283 vdd.n280 9.3005
R20053 vdd.n318 vdd.n317 9.3005
R20054 vdd.n240 vdd.n239 9.3005
R20055 vdd.n235 vdd.n234 9.3005
R20056 vdd.n246 vdd.n245 9.3005
R20057 vdd.n248 vdd.n247 9.3005
R20058 vdd.n231 vdd.n230 9.3005
R20059 vdd.n254 vdd.n253 9.3005
R20060 vdd.n256 vdd.n255 9.3005
R20061 vdd.n228 vdd.n225 9.3005
R20062 vdd.n263 vdd.n262 9.3005
R20063 vdd.n197 vdd.n196 9.3005
R20064 vdd.n192 vdd.n191 9.3005
R20065 vdd.n203 vdd.n202 9.3005
R20066 vdd.n205 vdd.n204 9.3005
R20067 vdd.n188 vdd.n187 9.3005
R20068 vdd.n211 vdd.n210 9.3005
R20069 vdd.n213 vdd.n212 9.3005
R20070 vdd.n185 vdd.n182 9.3005
R20071 vdd.n220 vdd.n219 9.3005
R20072 vdd.n142 vdd.n141 9.3005
R20073 vdd.n137 vdd.n136 9.3005
R20074 vdd.n148 vdd.n147 9.3005
R20075 vdd.n150 vdd.n149 9.3005
R20076 vdd.n133 vdd.n132 9.3005
R20077 vdd.n156 vdd.n155 9.3005
R20078 vdd.n158 vdd.n157 9.3005
R20079 vdd.n130 vdd.n127 9.3005
R20080 vdd.n165 vdd.n164 9.3005
R20081 vdd.n100 vdd.n99 9.3005
R20082 vdd.n95 vdd.n94 9.3005
R20083 vdd.n106 vdd.n105 9.3005
R20084 vdd.n108 vdd.n107 9.3005
R20085 vdd.n91 vdd.n90 9.3005
R20086 vdd.n114 vdd.n113 9.3005
R20087 vdd.n116 vdd.n115 9.3005
R20088 vdd.n88 vdd.n85 9.3005
R20089 vdd.n123 vdd.n122 9.3005
R20090 vdd.n45 vdd.n44 9.3005
R20091 vdd.n40 vdd.n39 9.3005
R20092 vdd.n51 vdd.n50 9.3005
R20093 vdd.n53 vdd.n52 9.3005
R20094 vdd.n36 vdd.n35 9.3005
R20095 vdd.n59 vdd.n58 9.3005
R20096 vdd.n61 vdd.n60 9.3005
R20097 vdd.n33 vdd.n30 9.3005
R20098 vdd.n68 vdd.n67 9.3005
R20099 vdd.n3059 vdd.n3058 9.3005
R20100 vdd.n3060 vdd.n721 9.3005
R20101 vdd.n720 vdd.n718 9.3005
R20102 vdd.n3066 vdd.n717 9.3005
R20103 vdd.n3067 vdd.n716 9.3005
R20104 vdd.n3068 vdd.n715 9.3005
R20105 vdd.n714 vdd.n712 9.3005
R20106 vdd.n3074 vdd.n711 9.3005
R20107 vdd.n3075 vdd.n710 9.3005
R20108 vdd.n3076 vdd.n709 9.3005
R20109 vdd.n708 vdd.n706 9.3005
R20110 vdd.n3082 vdd.n705 9.3005
R20111 vdd.n3083 vdd.n704 9.3005
R20112 vdd.n3084 vdd.n703 9.3005
R20113 vdd.n702 vdd.n700 9.3005
R20114 vdd.n3090 vdd.n699 9.3005
R20115 vdd.n3091 vdd.n698 9.3005
R20116 vdd.n3092 vdd.n697 9.3005
R20117 vdd.n696 vdd.n694 9.3005
R20118 vdd.n3098 vdd.n693 9.3005
R20119 vdd.n3099 vdd.n692 9.3005
R20120 vdd.n3100 vdd.n691 9.3005
R20121 vdd.n690 vdd.n688 9.3005
R20122 vdd.n3106 vdd.n685 9.3005
R20123 vdd.n3107 vdd.n684 9.3005
R20124 vdd.n3108 vdd.n683 9.3005
R20125 vdd.n682 vdd.n680 9.3005
R20126 vdd.n3114 vdd.n679 9.3005
R20127 vdd.n3115 vdd.n678 9.3005
R20128 vdd.n3116 vdd.n677 9.3005
R20129 vdd.n676 vdd.n674 9.3005
R20130 vdd.n3122 vdd.n673 9.3005
R20131 vdd.n3123 vdd.n672 9.3005
R20132 vdd.n3124 vdd.n671 9.3005
R20133 vdd.n670 vdd.n668 9.3005
R20134 vdd.n3129 vdd.n667 9.3005
R20135 vdd.n3139 vdd.n661 9.3005
R20136 vdd.n3141 vdd.n3140 9.3005
R20137 vdd.n652 vdd.n651 9.3005
R20138 vdd.n3156 vdd.n3155 9.3005
R20139 vdd.n3157 vdd.n650 9.3005
R20140 vdd.n3159 vdd.n3158 9.3005
R20141 vdd.n640 vdd.n639 9.3005
R20142 vdd.n3172 vdd.n3171 9.3005
R20143 vdd.n3173 vdd.n638 9.3005
R20144 vdd.n3175 vdd.n3174 9.3005
R20145 vdd.n628 vdd.n627 9.3005
R20146 vdd.n3189 vdd.n3188 9.3005
R20147 vdd.n3190 vdd.n626 9.3005
R20148 vdd.n3192 vdd.n3191 9.3005
R20149 vdd.n617 vdd.n616 9.3005
R20150 vdd.n3208 vdd.n3207 9.3005
R20151 vdd.n3209 vdd.n615 9.3005
R20152 vdd.n3211 vdd.n3210 9.3005
R20153 vdd.n324 vdd.n322 9.3005
R20154 vdd.n3143 vdd.n3142 9.3005
R20155 vdd.n3290 vdd.n3289 9.3005
R20156 vdd.n325 vdd.n323 9.3005
R20157 vdd.n3283 vdd.n334 9.3005
R20158 vdd.n3282 vdd.n335 9.3005
R20159 vdd.n3281 vdd.n336 9.3005
R20160 vdd.n343 vdd.n337 9.3005
R20161 vdd.n3275 vdd.n344 9.3005
R20162 vdd.n3274 vdd.n345 9.3005
R20163 vdd.n3273 vdd.n346 9.3005
R20164 vdd.n354 vdd.n347 9.3005
R20165 vdd.n3267 vdd.n355 9.3005
R20166 vdd.n3266 vdd.n356 9.3005
R20167 vdd.n3265 vdd.n357 9.3005
R20168 vdd.n365 vdd.n358 9.3005
R20169 vdd.n3259 vdd.n366 9.3005
R20170 vdd.n3258 vdd.n367 9.3005
R20171 vdd.n3257 vdd.n368 9.3005
R20172 vdd.n443 vdd.n369 9.3005
R20173 vdd.n447 vdd.n442 9.3005
R20174 vdd.n451 vdd.n450 9.3005
R20175 vdd.n452 vdd.n441 9.3005
R20176 vdd.n456 vdd.n453 9.3005
R20177 vdd.n457 vdd.n440 9.3005
R20178 vdd.n461 vdd.n460 9.3005
R20179 vdd.n462 vdd.n439 9.3005
R20180 vdd.n466 vdd.n463 9.3005
R20181 vdd.n467 vdd.n438 9.3005
R20182 vdd.n471 vdd.n470 9.3005
R20183 vdd.n472 vdd.n437 9.3005
R20184 vdd.n476 vdd.n473 9.3005
R20185 vdd.n477 vdd.n436 9.3005
R20186 vdd.n481 vdd.n480 9.3005
R20187 vdd.n482 vdd.n435 9.3005
R20188 vdd.n486 vdd.n483 9.3005
R20189 vdd.n487 vdd.n434 9.3005
R20190 vdd.n491 vdd.n490 9.3005
R20191 vdd.n492 vdd.n433 9.3005
R20192 vdd.n496 vdd.n493 9.3005
R20193 vdd.n497 vdd.n430 9.3005
R20194 vdd.n501 vdd.n500 9.3005
R20195 vdd.n502 vdd.n429 9.3005
R20196 vdd.n506 vdd.n503 9.3005
R20197 vdd.n507 vdd.n428 9.3005
R20198 vdd.n511 vdd.n510 9.3005
R20199 vdd.n512 vdd.n427 9.3005
R20200 vdd.n516 vdd.n513 9.3005
R20201 vdd.n517 vdd.n426 9.3005
R20202 vdd.n521 vdd.n520 9.3005
R20203 vdd.n522 vdd.n425 9.3005
R20204 vdd.n526 vdd.n523 9.3005
R20205 vdd.n527 vdd.n424 9.3005
R20206 vdd.n531 vdd.n530 9.3005
R20207 vdd.n532 vdd.n423 9.3005
R20208 vdd.n536 vdd.n533 9.3005
R20209 vdd.n537 vdd.n422 9.3005
R20210 vdd.n541 vdd.n540 9.3005
R20211 vdd.n542 vdd.n421 9.3005
R20212 vdd.n546 vdd.n543 9.3005
R20213 vdd.n547 vdd.n418 9.3005
R20214 vdd.n551 vdd.n550 9.3005
R20215 vdd.n552 vdd.n417 9.3005
R20216 vdd.n556 vdd.n553 9.3005
R20217 vdd.n557 vdd.n416 9.3005
R20218 vdd.n561 vdd.n560 9.3005
R20219 vdd.n562 vdd.n415 9.3005
R20220 vdd.n566 vdd.n563 9.3005
R20221 vdd.n567 vdd.n414 9.3005
R20222 vdd.n571 vdd.n570 9.3005
R20223 vdd.n572 vdd.n413 9.3005
R20224 vdd.n576 vdd.n573 9.3005
R20225 vdd.n577 vdd.n412 9.3005
R20226 vdd.n581 vdd.n580 9.3005
R20227 vdd.n582 vdd.n411 9.3005
R20228 vdd.n586 vdd.n583 9.3005
R20229 vdd.n587 vdd.n410 9.3005
R20230 vdd.n591 vdd.n590 9.3005
R20231 vdd.n592 vdd.n409 9.3005
R20232 vdd.n596 vdd.n593 9.3005
R20233 vdd.n598 vdd.n408 9.3005
R20234 vdd.n600 vdd.n599 9.3005
R20235 vdd.n3250 vdd.n3249 9.3005
R20236 vdd.n446 vdd.n444 9.3005
R20237 vdd.n3149 vdd.n655 9.3005
R20238 vdd.n3151 vdd.n3150 9.3005
R20239 vdd.n646 vdd.n645 9.3005
R20240 vdd.n3164 vdd.n3163 9.3005
R20241 vdd.n3165 vdd.n644 9.3005
R20242 vdd.n3167 vdd.n3166 9.3005
R20243 vdd.n633 vdd.n632 9.3005
R20244 vdd.n3180 vdd.n3179 9.3005
R20245 vdd.n3181 vdd.n631 9.3005
R20246 vdd.n3183 vdd.n3182 9.3005
R20247 vdd.n622 vdd.n621 9.3005
R20248 vdd.n3197 vdd.n3196 9.3005
R20249 vdd.n3198 vdd.n620 9.3005
R20250 vdd.n3203 vdd.n3199 9.3005
R20251 vdd.n3202 vdd.n3201 9.3005
R20252 vdd.n3200 vdd.n610 9.3005
R20253 vdd.n3216 vdd.n611 9.3005
R20254 vdd.n3217 vdd.n609 9.3005
R20255 vdd.n3219 vdd.n3218 9.3005
R20256 vdd.n3220 vdd.n608 9.3005
R20257 vdd.n3223 vdd.n3221 9.3005
R20258 vdd.n3224 vdd.n607 9.3005
R20259 vdd.n3226 vdd.n3225 9.3005
R20260 vdd.n3227 vdd.n606 9.3005
R20261 vdd.n3230 vdd.n3228 9.3005
R20262 vdd.n3231 vdd.n605 9.3005
R20263 vdd.n3233 vdd.n3232 9.3005
R20264 vdd.n3234 vdd.n604 9.3005
R20265 vdd.n3238 vdd.n3235 9.3005
R20266 vdd.n3239 vdd.n603 9.3005
R20267 vdd.n3241 vdd.n3240 9.3005
R20268 vdd.n3242 vdd.n602 9.3005
R20269 vdd.n3245 vdd.n3243 9.3005
R20270 vdd.n3246 vdd.n601 9.3005
R20271 vdd.n3248 vdd.n3247 9.3005
R20272 vdd.n3148 vdd.n3147 9.3005
R20273 vdd.n3012 vdd.n656 9.3005
R20274 vdd.n3017 vdd.n3011 9.3005
R20275 vdd.n3027 vdd.n748 9.3005
R20276 vdd.n3028 vdd.n747 9.3005
R20277 vdd.n746 vdd.n744 9.3005
R20278 vdd.n3034 vdd.n743 9.3005
R20279 vdd.n3035 vdd.n742 9.3005
R20280 vdd.n3036 vdd.n741 9.3005
R20281 vdd.n740 vdd.n738 9.3005
R20282 vdd.n3042 vdd.n737 9.3005
R20283 vdd.n3043 vdd.n736 9.3005
R20284 vdd.n3044 vdd.n735 9.3005
R20285 vdd.n734 vdd.n732 9.3005
R20286 vdd.n3049 vdd.n731 9.3005
R20287 vdd.n3050 vdd.n730 9.3005
R20288 vdd.n726 vdd.n725 9.3005
R20289 vdd.n3056 vdd.n3055 9.3005
R20290 vdd.n3057 vdd.n722 9.3005
R20291 vdd.n2254 vdd.n2253 9.3005
R20292 vdd.n2249 vdd.n1038 9.3005
R20293 vdd.n1380 vdd.n1379 9.3005
R20294 vdd.n1136 vdd.n1135 9.3005
R20295 vdd.n1393 vdd.n1392 9.3005
R20296 vdd.n1394 vdd.n1134 9.3005
R20297 vdd.n1396 vdd.n1395 9.3005
R20298 vdd.n1124 vdd.n1123 9.3005
R20299 vdd.n1410 vdd.n1409 9.3005
R20300 vdd.n1411 vdd.n1122 9.3005
R20301 vdd.n1413 vdd.n1412 9.3005
R20302 vdd.n1114 vdd.n1113 9.3005
R20303 vdd.n1427 vdd.n1426 9.3005
R20304 vdd.n1428 vdd.n1112 9.3005
R20305 vdd.n1430 vdd.n1429 9.3005
R20306 vdd.n1101 vdd.n1100 9.3005
R20307 vdd.n1443 vdd.n1442 9.3005
R20308 vdd.n1444 vdd.n1099 9.3005
R20309 vdd.n1446 vdd.n1445 9.3005
R20310 vdd.n1090 vdd.n1089 9.3005
R20311 vdd.n1755 vdd.n1754 9.3005
R20312 vdd.n1756 vdd.n1088 9.3005
R20313 vdd.n1758 vdd.n1757 9.3005
R20314 vdd.n1079 vdd.n1078 9.3005
R20315 vdd.n1771 vdd.n1770 9.3005
R20316 vdd.n1772 vdd.n1077 9.3005
R20317 vdd.n1774 vdd.n1773 9.3005
R20318 vdd.n1067 vdd.n1066 9.3005
R20319 vdd.n1788 vdd.n1787 9.3005
R20320 vdd.n1789 vdd.n1065 9.3005
R20321 vdd.n1791 vdd.n1790 9.3005
R20322 vdd.n1057 vdd.n1056 9.3005
R20323 vdd.n1805 vdd.n1804 9.3005
R20324 vdd.n1806 vdd.n1054 9.3005
R20325 vdd.n1810 vdd.n1809 9.3005
R20326 vdd.n1808 vdd.n1055 9.3005
R20327 vdd.n1807 vdd.n1043 9.3005
R20328 vdd.n1378 vdd.n1146 9.3005
R20329 vdd.n1271 vdd.n1147 9.3005
R20330 vdd.n1273 vdd.n1272 9.3005
R20331 vdd.n1274 vdd.n1266 9.3005
R20332 vdd.n1276 vdd.n1275 9.3005
R20333 vdd.n1277 vdd.n1265 9.3005
R20334 vdd.n1279 vdd.n1278 9.3005
R20335 vdd.n1280 vdd.n1260 9.3005
R20336 vdd.n1282 vdd.n1281 9.3005
R20337 vdd.n1283 vdd.n1259 9.3005
R20338 vdd.n1285 vdd.n1284 9.3005
R20339 vdd.n1286 vdd.n1254 9.3005
R20340 vdd.n1288 vdd.n1287 9.3005
R20341 vdd.n1289 vdd.n1253 9.3005
R20342 vdd.n1291 vdd.n1290 9.3005
R20343 vdd.n1292 vdd.n1248 9.3005
R20344 vdd.n1294 vdd.n1293 9.3005
R20345 vdd.n1295 vdd.n1247 9.3005
R20346 vdd.n1297 vdd.n1296 9.3005
R20347 vdd.n1298 vdd.n1242 9.3005
R20348 vdd.n1300 vdd.n1299 9.3005
R20349 vdd.n1301 vdd.n1241 9.3005
R20350 vdd.n1306 vdd.n1302 9.3005
R20351 vdd.n1307 vdd.n1237 9.3005
R20352 vdd.n1309 vdd.n1308 9.3005
R20353 vdd.n1310 vdd.n1236 9.3005
R20354 vdd.n1312 vdd.n1311 9.3005
R20355 vdd.n1313 vdd.n1231 9.3005
R20356 vdd.n1315 vdd.n1314 9.3005
R20357 vdd.n1316 vdd.n1230 9.3005
R20358 vdd.n1318 vdd.n1317 9.3005
R20359 vdd.n1319 vdd.n1225 9.3005
R20360 vdd.n1321 vdd.n1320 9.3005
R20361 vdd.n1322 vdd.n1224 9.3005
R20362 vdd.n1324 vdd.n1323 9.3005
R20363 vdd.n1325 vdd.n1219 9.3005
R20364 vdd.n1327 vdd.n1326 9.3005
R20365 vdd.n1328 vdd.n1218 9.3005
R20366 vdd.n1330 vdd.n1329 9.3005
R20367 vdd.n1331 vdd.n1213 9.3005
R20368 vdd.n1333 vdd.n1332 9.3005
R20369 vdd.n1334 vdd.n1212 9.3005
R20370 vdd.n1336 vdd.n1335 9.3005
R20371 vdd.n1337 vdd.n1209 9.3005
R20372 vdd.n1343 vdd.n1342 9.3005
R20373 vdd.n1344 vdd.n1208 9.3005
R20374 vdd.n1346 vdd.n1345 9.3005
R20375 vdd.n1347 vdd.n1203 9.3005
R20376 vdd.n1349 vdd.n1348 9.3005
R20377 vdd.n1350 vdd.n1202 9.3005
R20378 vdd.n1352 vdd.n1351 9.3005
R20379 vdd.n1353 vdd.n1197 9.3005
R20380 vdd.n1355 vdd.n1354 9.3005
R20381 vdd.n1356 vdd.n1196 9.3005
R20382 vdd.n1358 vdd.n1357 9.3005
R20383 vdd.n1359 vdd.n1191 9.3005
R20384 vdd.n1361 vdd.n1360 9.3005
R20385 vdd.n1362 vdd.n1190 9.3005
R20386 vdd.n1364 vdd.n1363 9.3005
R20387 vdd.n1365 vdd.n1186 9.3005
R20388 vdd.n1367 vdd.n1366 9.3005
R20389 vdd.n1368 vdd.n1185 9.3005
R20390 vdd.n1370 vdd.n1369 9.3005
R20391 vdd.n1371 vdd.n1184 9.3005
R20392 vdd.n1377 vdd.n1376 9.3005
R20393 vdd.n1385 vdd.n1384 9.3005
R20394 vdd.n1386 vdd.n1140 9.3005
R20395 vdd.n1388 vdd.n1387 9.3005
R20396 vdd.n1130 vdd.n1129 9.3005
R20397 vdd.n1402 vdd.n1401 9.3005
R20398 vdd.n1403 vdd.n1128 9.3005
R20399 vdd.n1405 vdd.n1404 9.3005
R20400 vdd.n1119 vdd.n1118 9.3005
R20401 vdd.n1419 vdd.n1418 9.3005
R20402 vdd.n1420 vdd.n1117 9.3005
R20403 vdd.n1422 vdd.n1421 9.3005
R20404 vdd.n1108 vdd.n1107 9.3005
R20405 vdd.n1435 vdd.n1434 9.3005
R20406 vdd.n1436 vdd.n1106 9.3005
R20407 vdd.n1438 vdd.n1437 9.3005
R20408 vdd.n1096 vdd.n1095 9.3005
R20409 vdd.n1452 vdd.n1451 9.3005
R20410 vdd.n1142 vdd.n1141 9.3005
R20411 vdd.n1664 vdd.n1663 9.3005
R20412 vdd.n1659 vdd.n1658 9.3005
R20413 vdd.n1670 vdd.n1669 9.3005
R20414 vdd.n1672 vdd.n1671 9.3005
R20415 vdd.n1655 vdd.n1654 9.3005
R20416 vdd.n1678 vdd.n1677 9.3005
R20417 vdd.n1680 vdd.n1679 9.3005
R20418 vdd.n1652 vdd.n1649 9.3005
R20419 vdd.n1687 vdd.n1686 9.3005
R20420 vdd.n1719 vdd.n1718 9.3005
R20421 vdd.n1714 vdd.n1713 9.3005
R20422 vdd.n1725 vdd.n1724 9.3005
R20423 vdd.n1727 vdd.n1726 9.3005
R20424 vdd.n1710 vdd.n1709 9.3005
R20425 vdd.n1733 vdd.n1732 9.3005
R20426 vdd.n1735 vdd.n1734 9.3005
R20427 vdd.n1707 vdd.n1704 9.3005
R20428 vdd.n1742 vdd.n1741 9.3005
R20429 vdd.n1566 vdd.n1565 9.3005
R20430 vdd.n1561 vdd.n1560 9.3005
R20431 vdd.n1572 vdd.n1571 9.3005
R20432 vdd.n1574 vdd.n1573 9.3005
R20433 vdd.n1557 vdd.n1556 9.3005
R20434 vdd.n1580 vdd.n1579 9.3005
R20435 vdd.n1582 vdd.n1581 9.3005
R20436 vdd.n1554 vdd.n1551 9.3005
R20437 vdd.n1589 vdd.n1588 9.3005
R20438 vdd.n1621 vdd.n1620 9.3005
R20439 vdd.n1616 vdd.n1615 9.3005
R20440 vdd.n1627 vdd.n1626 9.3005
R20441 vdd.n1629 vdd.n1628 9.3005
R20442 vdd.n1612 vdd.n1611 9.3005
R20443 vdd.n1635 vdd.n1634 9.3005
R20444 vdd.n1637 vdd.n1636 9.3005
R20445 vdd.n1609 vdd.n1606 9.3005
R20446 vdd.n1644 vdd.n1643 9.3005
R20447 vdd.n1469 vdd.n1468 9.3005
R20448 vdd.n1464 vdd.n1463 9.3005
R20449 vdd.n1475 vdd.n1474 9.3005
R20450 vdd.n1477 vdd.n1476 9.3005
R20451 vdd.n1460 vdd.n1459 9.3005
R20452 vdd.n1483 vdd.n1482 9.3005
R20453 vdd.n1485 vdd.n1484 9.3005
R20454 vdd.n1457 vdd.n1454 9.3005
R20455 vdd.n1492 vdd.n1491 9.3005
R20456 vdd.n1524 vdd.n1523 9.3005
R20457 vdd.n1519 vdd.n1518 9.3005
R20458 vdd.n1530 vdd.n1529 9.3005
R20459 vdd.n1532 vdd.n1531 9.3005
R20460 vdd.n1515 vdd.n1514 9.3005
R20461 vdd.n1538 vdd.n1537 9.3005
R20462 vdd.n1540 vdd.n1539 9.3005
R20463 vdd.n1512 vdd.n1509 9.3005
R20464 vdd.n1547 vdd.n1546 9.3005
R20465 vdd.n1398 vdd.t118 9.18308
R20466 vdd.n3236 vdd.t62 9.18308
R20467 vdd.n1424 vdd.t66 8.95635
R20468 vdd.t64 vdd.n3277 8.95635
R20469 vdd.n300 vdd.n299 8.92171
R20470 vdd.n245 vdd.n244 8.92171
R20471 vdd.n202 vdd.n201 8.92171
R20472 vdd.n147 vdd.n146 8.92171
R20473 vdd.n105 vdd.n104 8.92171
R20474 vdd.n50 vdd.n49 8.92171
R20475 vdd.n1669 vdd.n1668 8.92171
R20476 vdd.n1724 vdd.n1723 8.92171
R20477 vdd.n1571 vdd.n1570 8.92171
R20478 vdd.n1626 vdd.n1625 8.92171
R20479 vdd.n1474 vdd.n1473 8.92171
R20480 vdd.n1529 vdd.n1528 8.92171
R20481 vdd.n223 vdd.n125 8.81535
R20482 vdd.n1647 vdd.n1549 8.81535
R20483 vdd.n1104 vdd.t123 8.72962
R20484 vdd.t91 vdd.n3286 8.72962
R20485 vdd.n1760 vdd.t48 8.50289
R20486 vdd.n3205 vdd.t121 8.50289
R20487 vdd.n28 vdd.n14 8.42249
R20488 vdd.n1776 vdd.t60 8.27616
R20489 vdd.t107 vdd.n636 8.27616
R20490 vdd.n3292 vdd.n3291 8.16225
R20491 vdd.n1747 vdd.n1746 8.16225
R20492 vdd.n296 vdd.n290 8.14595
R20493 vdd.n241 vdd.n235 8.14595
R20494 vdd.n198 vdd.n192 8.14595
R20495 vdd.n143 vdd.n137 8.14595
R20496 vdd.n101 vdd.n95 8.14595
R20497 vdd.n46 vdd.n40 8.14595
R20498 vdd.n1665 vdd.n1659 8.14595
R20499 vdd.n1720 vdd.n1714 8.14595
R20500 vdd.n1567 vdd.n1561 8.14595
R20501 vdd.n1622 vdd.n1616 8.14595
R20502 vdd.n1470 vdd.n1464 8.14595
R20503 vdd.n1525 vdd.n1519 8.14595
R20504 vdd.n2840 vdd.n820 8.11757
R20505 vdd.n2314 vdd.n2313 8.11757
R20506 vdd.t185 vdd.n1138 7.8227
R20507 vdd.t181 vdd.n363 7.8227
R20508 vdd.n2292 vdd.n1014 7.70933
R20509 vdd.n2298 vdd.n1014 7.70933
R20510 vdd.n2304 vdd.n1008 7.70933
R20511 vdd.n2304 vdd.n1001 7.70933
R20512 vdd.n2310 vdd.n1001 7.70933
R20513 vdd.n2310 vdd.n1004 7.70933
R20514 vdd.n2317 vdd.n989 7.70933
R20515 vdd.n2323 vdd.n989 7.70933
R20516 vdd.n2329 vdd.n983 7.70933
R20517 vdd.n2335 vdd.n979 7.70933
R20518 vdd.n2341 vdd.n973 7.70933
R20519 vdd.n2353 vdd.n960 7.70933
R20520 vdd.n2359 vdd.n954 7.70933
R20521 vdd.n2359 vdd.n947 7.70933
R20522 vdd.n2367 vdd.n947 7.70933
R20523 vdd.n2374 vdd.t8 7.70933
R20524 vdd.n2449 vdd.t8 7.70933
R20525 vdd.n2781 vdd.t34 7.70933
R20526 vdd.n2787 vdd.t34 7.70933
R20527 vdd.n2793 vdd.n868 7.70933
R20528 vdd.n2799 vdd.n868 7.70933
R20529 vdd.n2799 vdd.n871 7.70933
R20530 vdd.n2805 vdd.n864 7.70933
R20531 vdd.n2817 vdd.n851 7.70933
R20532 vdd.n2823 vdd.n845 7.70933
R20533 vdd.n2829 vdd.n841 7.70933
R20534 vdd.n2835 vdd.n828 7.70933
R20535 vdd.n2843 vdd.n828 7.70933
R20536 vdd.n2849 vdd.n822 7.70933
R20537 vdd.n2849 vdd.n814 7.70933
R20538 vdd.n2900 vdd.n814 7.70933
R20539 vdd.n2900 vdd.n817 7.70933
R20540 vdd.n2906 vdd.n774 7.70933
R20541 vdd.n2976 vdd.n774 7.70933
R20542 vdd.n295 vdd.n292 7.3702
R20543 vdd.n240 vdd.n237 7.3702
R20544 vdd.n197 vdd.n194 7.3702
R20545 vdd.n142 vdd.n139 7.3702
R20546 vdd.n100 vdd.n97 7.3702
R20547 vdd.n45 vdd.n42 7.3702
R20548 vdd.n1664 vdd.n1661 7.3702
R20549 vdd.n1719 vdd.n1716 7.3702
R20550 vdd.n1566 vdd.n1563 7.3702
R20551 vdd.n1621 vdd.n1618 7.3702
R20552 vdd.n1469 vdd.n1466 7.3702
R20553 vdd.n1524 vdd.n1521 7.3702
R20554 vdd.n1307 vdd.n1306 6.98232
R20555 vdd.n1956 vdd.n1955 6.98232
R20556 vdd.n547 vdd.n546 6.98232
R20557 vdd.n3060 vdd.n3059 6.98232
R20558 vdd.n1794 vdd.t151 6.91577
R20559 vdd.n3169 vdd.t114 6.91577
R20560 vdd.t81 vdd.n1075 6.68904
R20561 vdd.n3185 vdd.t79 6.68904
R20562 vdd.n1752 vdd.t132 6.46231
R20563 vdd.n3213 vdd.t89 6.46231
R20564 vdd.n3292 vdd.n321 6.32949
R20565 vdd.n1746 vdd.n1745 6.32949
R20566 vdd.t94 vdd.n1103 6.23558
R20567 vdd.t84 vdd.n332 6.23558
R20568 vdd.n1416 vdd.t116 6.00885
R20569 vdd.n2329 vdd.t39 6.00885
R20570 vdd.n2829 vdd.t25 6.00885
R20571 vdd.n3271 vdd.t87 6.00885
R20572 vdd.n1004 vdd.t230 5.89549
R20573 vdd.t199 vdd.n822 5.89549
R20574 vdd.n296 vdd.n295 5.81868
R20575 vdd.n241 vdd.n240 5.81868
R20576 vdd.n198 vdd.n197 5.81868
R20577 vdd.n143 vdd.n142 5.81868
R20578 vdd.n101 vdd.n100 5.81868
R20579 vdd.n46 vdd.n45 5.81868
R20580 vdd.n1665 vdd.n1664 5.81868
R20581 vdd.n1720 vdd.n1719 5.81868
R20582 vdd.n1567 vdd.n1566 5.81868
R20583 vdd.n1622 vdd.n1621 5.81868
R20584 vdd.n1470 vdd.n1469 5.81868
R20585 vdd.n1525 vdd.n1524 5.81868
R20586 vdd.t173 vdd.n1008 5.78212
R20587 vdd.n2073 vdd.t212 5.78212
R20588 vdd.n2698 vdd.t220 5.78212
R20589 vdd.n817 vdd.t216 5.78212
R20590 vdd.n2457 vdd.n2456 5.77611
R20591 vdd.n2200 vdd.n2070 5.77611
R20592 vdd.n2711 vdd.n2710 5.77611
R20593 vdd.n2915 vdd.n806 5.77611
R20594 vdd.n2981 vdd.n770 5.77611
R20595 vdd.n2621 vdd.n2561 5.77611
R20596 vdd.n2382 vdd.n938 5.77611
R20597 vdd.n2130 vdd.n2129 5.77611
R20598 vdd.n1376 vdd.n1150 5.62474
R20599 vdd.n2252 vdd.n2249 5.62474
R20600 vdd.n3250 vdd.n407 5.62474
R20601 vdd.n3015 vdd.n3012 5.62474
R20602 vdd.t258 vdd.n960 5.44203
R20603 vdd.n864 vdd.t4 5.44203
R20604 vdd.n1126 vdd.t116 5.32866
R20605 vdd.t87 vdd.n3270 5.32866
R20606 vdd.n1432 vdd.t94 5.10193
R20607 vdd.t18 vdd.n983 5.10193
R20608 vdd.n973 vdd.t1 5.10193
R20609 vdd.t22 vdd.n851 5.10193
R20610 vdd.n841 vdd.t13 5.10193
R20611 vdd.n3279 vdd.t84 5.10193
R20612 vdd.n299 vdd.n290 5.04292
R20613 vdd.n244 vdd.n235 5.04292
R20614 vdd.n201 vdd.n192 5.04292
R20615 vdd.n146 vdd.n137 5.04292
R20616 vdd.n104 vdd.n95 5.04292
R20617 vdd.n49 vdd.n40 5.04292
R20618 vdd.n1668 vdd.n1659 5.04292
R20619 vdd.n1723 vdd.n1714 5.04292
R20620 vdd.n1570 vdd.n1561 5.04292
R20621 vdd.n1625 vdd.n1616 5.04292
R20622 vdd.n1473 vdd.n1464 5.04292
R20623 vdd.n1528 vdd.n1519 5.04292
R20624 vdd.n1448 vdd.t132 4.8752
R20625 vdd.t21 vdd.t2 4.8752
R20626 vdd.t12 vdd.t32 4.8752
R20627 vdd.t250 vdd.t23 4.8752
R20628 vdd.t262 vdd.t38 4.8752
R20629 vdd.t89 vdd.n328 4.8752
R20630 vdd.n2458 vdd.n2457 4.83952
R20631 vdd.n2070 vdd.n2066 4.83952
R20632 vdd.n2712 vdd.n2711 4.83952
R20633 vdd.n806 vdd.n801 4.83952
R20634 vdd.n770 vdd.n765 4.83952
R20635 vdd.n2618 vdd.n2561 4.83952
R20636 vdd.n2385 vdd.n938 4.83952
R20637 vdd.n2129 vdd.n2128 4.83952
R20638 vdd.n1924 vdd.n1036 4.74817
R20639 vdd.n1919 vdd.n1037 4.74817
R20640 vdd.n1821 vdd.n1818 4.74817
R20641 vdd.n2233 vdd.n1822 4.74817
R20642 vdd.n2235 vdd.n1821 4.74817
R20643 vdd.n2234 vdd.n2233 4.74817
R20644 vdd.n664 vdd.n662 4.74817
R20645 vdd.n3130 vdd.n665 4.74817
R20646 vdd.n3133 vdd.n665 4.74817
R20647 vdd.n3134 vdd.n664 4.74817
R20648 vdd.n3022 vdd.n749 4.74817
R20649 vdd.n3018 vdd.n751 4.74817
R20650 vdd.n3021 vdd.n751 4.74817
R20651 vdd.n3026 vdd.n749 4.74817
R20652 vdd.n1920 vdd.n1036 4.74817
R20653 vdd.n1039 vdd.n1037 4.74817
R20654 vdd.n321 vdd.n320 4.7074
R20655 vdd.n223 vdd.n222 4.7074
R20656 vdd.n1745 vdd.n1744 4.7074
R20657 vdd.n1647 vdd.n1646 4.7074
R20658 vdd.n1768 vdd.t81 4.64847
R20659 vdd.n3194 vdd.t79 4.64847
R20660 vdd.n2335 vdd.t6 4.53511
R20661 vdd.n2823 vdd.t260 4.53511
R20662 vdd.n1069 vdd.t151 4.42174
R20663 vdd.t114 vdd.n635 4.42174
R20664 vdd.n2367 vdd.t41 4.30838
R20665 vdd.n2793 vdd.t256 4.30838
R20666 vdd.n300 vdd.n288 4.26717
R20667 vdd.n245 vdd.n233 4.26717
R20668 vdd.n202 vdd.n190 4.26717
R20669 vdd.n147 vdd.n135 4.26717
R20670 vdd.n105 vdd.n93 4.26717
R20671 vdd.n50 vdd.n38 4.26717
R20672 vdd.n1669 vdd.n1657 4.26717
R20673 vdd.n1724 vdd.n1712 4.26717
R20674 vdd.n1571 vdd.n1559 4.26717
R20675 vdd.n1626 vdd.n1614 4.26717
R20676 vdd.n1474 vdd.n1462 4.26717
R20677 vdd.n1529 vdd.n1517 4.26717
R20678 vdd.n321 vdd.n223 4.10845
R20679 vdd.n1745 vdd.n1647 4.10845
R20680 vdd.n277 vdd.t168 4.06363
R20681 vdd.n277 vdd.t78 4.06363
R20682 vdd.n275 vdd.t99 4.06363
R20683 vdd.n275 vdd.t167 4.06363
R20684 vdd.n273 vdd.t166 4.06363
R20685 vdd.n273 vdd.t98 4.06363
R20686 vdd.n271 vdd.t104 4.06363
R20687 vdd.n271 vdd.t106 4.06363
R20688 vdd.n269 vdd.t122 4.06363
R20689 vdd.n269 vdd.t68 4.06363
R20690 vdd.n267 vdd.t75 4.06363
R20691 vdd.n267 vdd.t126 4.06363
R20692 vdd.n265 vdd.t127 4.06363
R20693 vdd.n265 vdd.t150 4.06363
R20694 vdd.n179 vdd.t156 4.06363
R20695 vdd.n179 vdd.t63 4.06363
R20696 vdd.n177 vdd.t86 4.06363
R20697 vdd.n177 vdd.t155 4.06363
R20698 vdd.n175 vdd.t159 4.06363
R20699 vdd.n175 vdd.t85 4.06363
R20700 vdd.n173 vdd.t90 4.06363
R20701 vdd.n173 vdd.t92 4.06363
R20702 vdd.n171 vdd.t136 4.06363
R20703 vdd.n171 vdd.t45 4.06363
R20704 vdd.n169 vdd.t53 4.06363
R20705 vdd.n169 vdd.t101 4.06363
R20706 vdd.n167 vdd.t115 4.06363
R20707 vdd.n167 vdd.t139 4.06363
R20708 vdd.n82 vdd.t88 4.06363
R20709 vdd.n82 vdd.t153 4.06363
R20710 vdd.n80 vdd.t65 4.06363
R20711 vdd.n80 vdd.t111 4.06363
R20712 vdd.n78 vdd.t55 4.06363
R20713 vdd.n78 vdd.t93 4.06363
R20714 vdd.n76 vdd.t164 4.06363
R20715 vdd.n76 vdd.t143 4.06363
R20716 vdd.n74 vdd.t146 4.06363
R20717 vdd.n74 vdd.t100 4.06363
R20718 vdd.n72 vdd.t169 4.06363
R20719 vdd.n72 vdd.t80 4.06363
R20720 vdd.n70 vdd.t157 4.06363
R20721 vdd.n70 vdd.t108 4.06363
R20722 vdd.n1689 vdd.t71 4.06363
R20723 vdd.n1689 vdd.t162 4.06363
R20724 vdd.n1691 vdd.t160 4.06363
R20725 vdd.n1691 vdd.t144 4.06363
R20726 vdd.n1693 vdd.t120 4.06363
R20727 vdd.n1693 vdd.t74 4.06363
R20728 vdd.n1695 vdd.t171 4.06363
R20729 vdd.n1695 vdd.t142 4.06363
R20730 vdd.n1697 vdd.t140 4.06363
R20731 vdd.n1697 vdd.t97 4.06363
R20732 vdd.n1699 vdd.t96 4.06363
R20733 vdd.n1699 vdd.t141 4.06363
R20734 vdd.n1701 vdd.t129 4.06363
R20735 vdd.n1701 vdd.t128 4.06363
R20736 vdd.n1591 vdd.t61 4.06363
R20737 vdd.n1591 vdd.t152 4.06363
R20738 vdd.n1593 vdd.t145 4.06363
R20739 vdd.n1593 vdd.t135 4.06363
R20740 vdd.n1595 vdd.t105 4.06363
R20741 vdd.n1595 vdd.t49 4.06363
R20742 vdd.n1597 vdd.t161 4.06363
R20743 vdd.n1597 vdd.t133 4.06363
R20744 vdd.n1599 vdd.t130 4.06363
R20745 vdd.n1599 vdd.t83 4.06363
R20746 vdd.n1601 vdd.t77 4.06363
R20747 vdd.n1601 vdd.t131 4.06363
R20748 vdd.n1603 vdd.t119 4.06363
R20749 vdd.n1603 vdd.t117 4.06363
R20750 vdd.n1494 vdd.t109 4.06363
R20751 vdd.n1494 vdd.t158 4.06363
R20752 vdd.n1496 vdd.t82 4.06363
R20753 vdd.n1496 vdd.t138 4.06363
R20754 vdd.n1498 vdd.t103 4.06363
R20755 vdd.n1498 vdd.t147 4.06363
R20756 vdd.n1500 vdd.t124 4.06363
R20757 vdd.n1500 vdd.t165 4.06363
R20758 vdd.n1502 vdd.t95 4.06363
R20759 vdd.n1502 vdd.t59 4.06363
R20760 vdd.n1504 vdd.t112 4.06363
R20761 vdd.n1504 vdd.t67 4.06363
R20762 vdd.n1506 vdd.t154 4.06363
R20763 vdd.n1506 vdd.t170 4.06363
R20764 vdd.n26 vdd.t40 3.9605
R20765 vdd.n26 vdd.t27 3.9605
R20766 vdd.n23 vdd.t26 3.9605
R20767 vdd.n23 vdd.t29 3.9605
R20768 vdd.n21 vdd.t253 3.9605
R20769 vdd.n21 vdd.t30 3.9605
R20770 vdd.n20 vdd.t17 3.9605
R20771 vdd.n20 vdd.t255 3.9605
R20772 vdd.n15 vdd.t252 3.9605
R20773 vdd.n15 vdd.t254 3.9605
R20774 vdd.n16 vdd.t16 3.9605
R20775 vdd.n16 vdd.t14 3.9605
R20776 vdd.n18 vdd.t28 3.9605
R20777 vdd.n18 vdd.t43 3.9605
R20778 vdd.n25 vdd.t15 3.9605
R20779 vdd.n25 vdd.t24 3.9605
R20780 vdd.n7 vdd.t263 3.61217
R20781 vdd.n7 vdd.t261 3.61217
R20782 vdd.n8 vdd.t251 3.61217
R20783 vdd.n8 vdd.t5 3.61217
R20784 vdd.n10 vdd.t35 3.61217
R20785 vdd.n10 vdd.t257 3.61217
R20786 vdd.n12 vdd.t20 3.61217
R20787 vdd.n12 vdd.t37 3.61217
R20788 vdd.n5 vdd.t11 3.61217
R20789 vdd.n5 vdd.t249 3.61217
R20790 vdd.n3 vdd.t42 3.61217
R20791 vdd.n3 vdd.t9 3.61217
R20792 vdd.n1 vdd.t259 3.61217
R20793 vdd.n1 vdd.t33 3.61217
R20794 vdd.n0 vdd.t7 3.61217
R20795 vdd.n0 vdd.t3 3.61217
R20796 vdd.n1382 vdd.t185 3.51482
R20797 vdd.n3255 vdd.t181 3.51482
R20798 vdd.n304 vdd.n303 3.49141
R20799 vdd.n249 vdd.n248 3.49141
R20800 vdd.n206 vdd.n205 3.49141
R20801 vdd.n151 vdd.n150 3.49141
R20802 vdd.n109 vdd.n108 3.49141
R20803 vdd.n54 vdd.n53 3.49141
R20804 vdd.n1673 vdd.n1672 3.49141
R20805 vdd.n1728 vdd.n1727 3.49141
R20806 vdd.n1575 vdd.n1574 3.49141
R20807 vdd.n1630 vdd.n1629 3.49141
R20808 vdd.n1478 vdd.n1477 3.49141
R20809 vdd.n1533 vdd.n1532 3.49141
R20810 vdd.n2073 vdd.t41 3.40145
R20811 vdd.n2521 vdd.t10 3.40145
R20812 vdd.n2774 vdd.t36 3.40145
R20813 vdd.n2698 vdd.t256 3.40145
R20814 vdd.n2174 vdd.t6 3.17472
R20815 vdd.n2677 vdd.t260 3.17472
R20816 vdd.n1785 vdd.t60 3.06136
R20817 vdd.n3177 vdd.t107 3.06136
R20818 vdd.t48 vdd.n1081 2.83463
R20819 vdd.n624 vdd.t121 2.83463
R20820 vdd.n307 vdd.n286 2.71565
R20821 vdd.n252 vdd.n231 2.71565
R20822 vdd.n209 vdd.n188 2.71565
R20823 vdd.n154 vdd.n133 2.71565
R20824 vdd.n112 vdd.n91 2.71565
R20825 vdd.n57 vdd.n36 2.71565
R20826 vdd.n1676 vdd.n1655 2.71565
R20827 vdd.n1731 vdd.n1710 2.71565
R20828 vdd.n1578 vdd.n1557 2.71565
R20829 vdd.n1633 vdd.n1612 2.71565
R20830 vdd.n1481 vdd.n1460 2.71565
R20831 vdd.n1536 vdd.n1515 2.71565
R20832 vdd.n1449 vdd.t123 2.6079
R20833 vdd.n2323 vdd.t18 2.6079
R20834 vdd.n2347 vdd.t1 2.6079
R20835 vdd.n2811 vdd.t22 2.6079
R20836 vdd.n2835 vdd.t13 2.6079
R20837 vdd.n3287 vdd.t91 2.6079
R20838 vdd.n2841 vdd.n2840 2.49806
R20839 vdd.n2315 vdd.n2314 2.49806
R20840 vdd.n294 vdd.n293 2.4129
R20841 vdd.n239 vdd.n238 2.4129
R20842 vdd.n196 vdd.n195 2.4129
R20843 vdd.n141 vdd.n140 2.4129
R20844 vdd.n99 vdd.n98 2.4129
R20845 vdd.n44 vdd.n43 2.4129
R20846 vdd.n1663 vdd.n1662 2.4129
R20847 vdd.n1718 vdd.n1717 2.4129
R20848 vdd.n1565 vdd.n1564 2.4129
R20849 vdd.n1620 vdd.n1619 2.4129
R20850 vdd.n1468 vdd.n1467 2.4129
R20851 vdd.n1523 vdd.n1522 2.4129
R20852 vdd.t66 vdd.n1110 2.38117
R20853 vdd.n3278 vdd.t64 2.38117
R20854 vdd.n2232 vdd.n1821 2.27742
R20855 vdd.n2233 vdd.n2232 2.27742
R20856 vdd.n2942 vdd.n665 2.27742
R20857 vdd.n2942 vdd.n664 2.27742
R20858 vdd.n3010 vdd.n751 2.27742
R20859 vdd.n3010 vdd.n749 2.27742
R20860 vdd.n2255 vdd.n1036 2.27742
R20861 vdd.n2255 vdd.n1037 2.27742
R20862 vdd.n2347 vdd.t258 2.2678
R20863 vdd.n2811 vdd.t4 2.2678
R20864 vdd.n1407 vdd.t118 2.15444
R20865 vdd.n3269 vdd.t62 2.15444
R20866 vdd.t32 vdd.n954 2.04107
R20867 vdd.n871 vdd.t250 2.04107
R20868 vdd.n308 vdd.n284 1.93989
R20869 vdd.n253 vdd.n229 1.93989
R20870 vdd.n210 vdd.n186 1.93989
R20871 vdd.n155 vdd.n131 1.93989
R20872 vdd.n113 vdd.n89 1.93989
R20873 vdd.n58 vdd.n34 1.93989
R20874 vdd.n1677 vdd.n1653 1.93989
R20875 vdd.n1732 vdd.n1708 1.93989
R20876 vdd.n1579 vdd.n1555 1.93989
R20877 vdd.n1634 vdd.n1610 1.93989
R20878 vdd.n1482 vdd.n1458 1.93989
R20879 vdd.n1537 vdd.n1513 1.93989
R20880 vdd.n2298 vdd.t173 1.92771
R20881 vdd.n2374 vdd.t212 1.92771
R20882 vdd.n2787 vdd.t220 1.92771
R20883 vdd.n2906 vdd.t216 1.92771
R20884 vdd.n1399 vdd.t56 1.70098
R20885 vdd.n2174 vdd.t39 1.70098
R20886 vdd.n979 vdd.t21 1.70098
R20887 vdd.t38 vdd.n845 1.70098
R20888 vdd.n2677 vdd.t25 1.70098
R20889 vdd.n3263 vdd.t69 1.70098
R20890 vdd.n1415 vdd.t76 1.47425
R20891 vdd.n349 vdd.t110 1.47425
R20892 vdd.n1440 vdd.t58 1.24752
R20893 vdd.t192 vdd.n1044 1.24752
R20894 vdd.n659 vdd.t177 1.24752
R20895 vdd.t54 vdd.n3285 1.24752
R20896 vdd.n319 vdd.n279 1.16414
R20897 vdd.n312 vdd.n311 1.16414
R20898 vdd.n264 vdd.n224 1.16414
R20899 vdd.n257 vdd.n256 1.16414
R20900 vdd.n221 vdd.n181 1.16414
R20901 vdd.n214 vdd.n213 1.16414
R20902 vdd.n166 vdd.n126 1.16414
R20903 vdd.n159 vdd.n158 1.16414
R20904 vdd.n124 vdd.n84 1.16414
R20905 vdd.n117 vdd.n116 1.16414
R20906 vdd.n69 vdd.n29 1.16414
R20907 vdd.n62 vdd.n61 1.16414
R20908 vdd.n1688 vdd.n1648 1.16414
R20909 vdd.n1681 vdd.n1680 1.16414
R20910 vdd.n1743 vdd.n1703 1.16414
R20911 vdd.n1736 vdd.n1735 1.16414
R20912 vdd.n1590 vdd.n1550 1.16414
R20913 vdd.n1583 vdd.n1582 1.16414
R20914 vdd.n1645 vdd.n1605 1.16414
R20915 vdd.n1638 vdd.n1637 1.16414
R20916 vdd.n1493 vdd.n1453 1.16414
R20917 vdd.n1486 vdd.n1485 1.16414
R20918 vdd.n1548 vdd.n1508 1.16414
R20919 vdd.n1541 vdd.n1540 1.16414
R20920 vdd.n2341 vdd.t2 1.13415
R20921 vdd.n2817 vdd.t262 1.13415
R20922 vdd.n1092 vdd.t102 1.02079
R20923 vdd.t230 vdd.t31 1.02079
R20924 vdd.t0 vdd.t199 1.02079
R20925 vdd.t44 vdd.n613 1.02079
R20926 vdd.n1271 vdd.n1150 0.970197
R20927 vdd.n2253 vdd.n2252 0.970197
R20928 vdd.n599 vdd.n407 0.970197
R20929 vdd.n3017 vdd.n3015 0.970197
R20930 vdd.n1746 vdd.n28 0.852297
R20931 vdd vdd.n3292 0.844463
R20932 vdd.n1777 vdd.t134 0.794056
R20933 vdd.n2317 vdd.t31 0.794056
R20934 vdd.n2353 vdd.t12 0.794056
R20935 vdd.n2805 vdd.t23 0.794056
R20936 vdd.n2843 vdd.t0 0.794056
R20937 vdd.n3186 vdd.t52 0.794056
R20938 vdd.n1793 vdd.t50 0.567326
R20939 vdd.t46 vdd.n642 0.567326
R20940 vdd.n2243 vdd.n2242 0.482207
R20941 vdd.n3142 vdd.n3141 0.482207
R20942 vdd.n444 vdd.n443 0.482207
R20943 vdd.n3249 vdd.n3248 0.482207
R20944 vdd.n3148 vdd.n656 0.482207
R20945 vdd.n1807 vdd.n1038 0.482207
R20946 vdd.n1378 vdd.n1377 0.482207
R20947 vdd.n1184 vdd.n1141 0.482207
R20948 vdd.n4 vdd.n2 0.459552
R20949 vdd.n11 vdd.n9 0.459552
R20950 vdd.n317 vdd.n316 0.388379
R20951 vdd.n283 vdd.n281 0.388379
R20952 vdd.n262 vdd.n261 0.388379
R20953 vdd.n228 vdd.n226 0.388379
R20954 vdd.n219 vdd.n218 0.388379
R20955 vdd.n185 vdd.n183 0.388379
R20956 vdd.n164 vdd.n163 0.388379
R20957 vdd.n130 vdd.n128 0.388379
R20958 vdd.n122 vdd.n121 0.388379
R20959 vdd.n88 vdd.n86 0.388379
R20960 vdd.n67 vdd.n66 0.388379
R20961 vdd.n33 vdd.n31 0.388379
R20962 vdd.n1686 vdd.n1685 0.388379
R20963 vdd.n1652 vdd.n1650 0.388379
R20964 vdd.n1741 vdd.n1740 0.388379
R20965 vdd.n1707 vdd.n1705 0.388379
R20966 vdd.n1588 vdd.n1587 0.388379
R20967 vdd.n1554 vdd.n1552 0.388379
R20968 vdd.n1643 vdd.n1642 0.388379
R20969 vdd.n1609 vdd.n1607 0.388379
R20970 vdd.n1491 vdd.n1490 0.388379
R20971 vdd.n1457 vdd.n1455 0.388379
R20972 vdd.n1546 vdd.n1545 0.388379
R20973 vdd.n1512 vdd.n1510 0.388379
R20974 vdd.n19 vdd.n17 0.387128
R20975 vdd.n24 vdd.n22 0.387128
R20976 vdd.n6 vdd.n4 0.358259
R20977 vdd.n13 vdd.n11 0.358259
R20978 vdd.n268 vdd.n266 0.358259
R20979 vdd.n270 vdd.n268 0.358259
R20980 vdd.n272 vdd.n270 0.358259
R20981 vdd.n274 vdd.n272 0.358259
R20982 vdd.n276 vdd.n274 0.358259
R20983 vdd.n278 vdd.n276 0.358259
R20984 vdd.n320 vdd.n278 0.358259
R20985 vdd.n170 vdd.n168 0.358259
R20986 vdd.n172 vdd.n170 0.358259
R20987 vdd.n174 vdd.n172 0.358259
R20988 vdd.n176 vdd.n174 0.358259
R20989 vdd.n178 vdd.n176 0.358259
R20990 vdd.n180 vdd.n178 0.358259
R20991 vdd.n222 vdd.n180 0.358259
R20992 vdd.n73 vdd.n71 0.358259
R20993 vdd.n75 vdd.n73 0.358259
R20994 vdd.n77 vdd.n75 0.358259
R20995 vdd.n79 vdd.n77 0.358259
R20996 vdd.n81 vdd.n79 0.358259
R20997 vdd.n83 vdd.n81 0.358259
R20998 vdd.n125 vdd.n83 0.358259
R20999 vdd.n1744 vdd.n1702 0.358259
R21000 vdd.n1702 vdd.n1700 0.358259
R21001 vdd.n1700 vdd.n1698 0.358259
R21002 vdd.n1698 vdd.n1696 0.358259
R21003 vdd.n1696 vdd.n1694 0.358259
R21004 vdd.n1694 vdd.n1692 0.358259
R21005 vdd.n1692 vdd.n1690 0.358259
R21006 vdd.n1646 vdd.n1604 0.358259
R21007 vdd.n1604 vdd.n1602 0.358259
R21008 vdd.n1602 vdd.n1600 0.358259
R21009 vdd.n1600 vdd.n1598 0.358259
R21010 vdd.n1598 vdd.n1596 0.358259
R21011 vdd.n1596 vdd.n1594 0.358259
R21012 vdd.n1594 vdd.n1592 0.358259
R21013 vdd.n1549 vdd.n1507 0.358259
R21014 vdd.n1507 vdd.n1505 0.358259
R21015 vdd.n1505 vdd.n1503 0.358259
R21016 vdd.n1503 vdd.n1501 0.358259
R21017 vdd.n1501 vdd.n1499 0.358259
R21018 vdd.n1499 vdd.n1497 0.358259
R21019 vdd.n1497 vdd.n1495 0.358259
R21020 vdd.n14 vdd.n6 0.334552
R21021 vdd.n14 vdd.n13 0.334552
R21022 vdd.n27 vdd.n19 0.21707
R21023 vdd.n27 vdd.n24 0.21707
R21024 vdd.n318 vdd.n280 0.155672
R21025 vdd.n310 vdd.n280 0.155672
R21026 vdd.n310 vdd.n309 0.155672
R21027 vdd.n309 vdd.n285 0.155672
R21028 vdd.n302 vdd.n285 0.155672
R21029 vdd.n302 vdd.n301 0.155672
R21030 vdd.n301 vdd.n289 0.155672
R21031 vdd.n294 vdd.n289 0.155672
R21032 vdd.n263 vdd.n225 0.155672
R21033 vdd.n255 vdd.n225 0.155672
R21034 vdd.n255 vdd.n254 0.155672
R21035 vdd.n254 vdd.n230 0.155672
R21036 vdd.n247 vdd.n230 0.155672
R21037 vdd.n247 vdd.n246 0.155672
R21038 vdd.n246 vdd.n234 0.155672
R21039 vdd.n239 vdd.n234 0.155672
R21040 vdd.n220 vdd.n182 0.155672
R21041 vdd.n212 vdd.n182 0.155672
R21042 vdd.n212 vdd.n211 0.155672
R21043 vdd.n211 vdd.n187 0.155672
R21044 vdd.n204 vdd.n187 0.155672
R21045 vdd.n204 vdd.n203 0.155672
R21046 vdd.n203 vdd.n191 0.155672
R21047 vdd.n196 vdd.n191 0.155672
R21048 vdd.n165 vdd.n127 0.155672
R21049 vdd.n157 vdd.n127 0.155672
R21050 vdd.n157 vdd.n156 0.155672
R21051 vdd.n156 vdd.n132 0.155672
R21052 vdd.n149 vdd.n132 0.155672
R21053 vdd.n149 vdd.n148 0.155672
R21054 vdd.n148 vdd.n136 0.155672
R21055 vdd.n141 vdd.n136 0.155672
R21056 vdd.n123 vdd.n85 0.155672
R21057 vdd.n115 vdd.n85 0.155672
R21058 vdd.n115 vdd.n114 0.155672
R21059 vdd.n114 vdd.n90 0.155672
R21060 vdd.n107 vdd.n90 0.155672
R21061 vdd.n107 vdd.n106 0.155672
R21062 vdd.n106 vdd.n94 0.155672
R21063 vdd.n99 vdd.n94 0.155672
R21064 vdd.n68 vdd.n30 0.155672
R21065 vdd.n60 vdd.n30 0.155672
R21066 vdd.n60 vdd.n59 0.155672
R21067 vdd.n59 vdd.n35 0.155672
R21068 vdd.n52 vdd.n35 0.155672
R21069 vdd.n52 vdd.n51 0.155672
R21070 vdd.n51 vdd.n39 0.155672
R21071 vdd.n44 vdd.n39 0.155672
R21072 vdd.n1687 vdd.n1649 0.155672
R21073 vdd.n1679 vdd.n1649 0.155672
R21074 vdd.n1679 vdd.n1678 0.155672
R21075 vdd.n1678 vdd.n1654 0.155672
R21076 vdd.n1671 vdd.n1654 0.155672
R21077 vdd.n1671 vdd.n1670 0.155672
R21078 vdd.n1670 vdd.n1658 0.155672
R21079 vdd.n1663 vdd.n1658 0.155672
R21080 vdd.n1742 vdd.n1704 0.155672
R21081 vdd.n1734 vdd.n1704 0.155672
R21082 vdd.n1734 vdd.n1733 0.155672
R21083 vdd.n1733 vdd.n1709 0.155672
R21084 vdd.n1726 vdd.n1709 0.155672
R21085 vdd.n1726 vdd.n1725 0.155672
R21086 vdd.n1725 vdd.n1713 0.155672
R21087 vdd.n1718 vdd.n1713 0.155672
R21088 vdd.n1589 vdd.n1551 0.155672
R21089 vdd.n1581 vdd.n1551 0.155672
R21090 vdd.n1581 vdd.n1580 0.155672
R21091 vdd.n1580 vdd.n1556 0.155672
R21092 vdd.n1573 vdd.n1556 0.155672
R21093 vdd.n1573 vdd.n1572 0.155672
R21094 vdd.n1572 vdd.n1560 0.155672
R21095 vdd.n1565 vdd.n1560 0.155672
R21096 vdd.n1644 vdd.n1606 0.155672
R21097 vdd.n1636 vdd.n1606 0.155672
R21098 vdd.n1636 vdd.n1635 0.155672
R21099 vdd.n1635 vdd.n1611 0.155672
R21100 vdd.n1628 vdd.n1611 0.155672
R21101 vdd.n1628 vdd.n1627 0.155672
R21102 vdd.n1627 vdd.n1615 0.155672
R21103 vdd.n1620 vdd.n1615 0.155672
R21104 vdd.n1492 vdd.n1454 0.155672
R21105 vdd.n1484 vdd.n1454 0.155672
R21106 vdd.n1484 vdd.n1483 0.155672
R21107 vdd.n1483 vdd.n1459 0.155672
R21108 vdd.n1476 vdd.n1459 0.155672
R21109 vdd.n1476 vdd.n1475 0.155672
R21110 vdd.n1475 vdd.n1463 0.155672
R21111 vdd.n1468 vdd.n1463 0.155672
R21112 vdd.n1547 vdd.n1509 0.155672
R21113 vdd.n1539 vdd.n1509 0.155672
R21114 vdd.n1539 vdd.n1538 0.155672
R21115 vdd.n1538 vdd.n1514 0.155672
R21116 vdd.n1531 vdd.n1514 0.155672
R21117 vdd.n1531 vdd.n1530 0.155672
R21118 vdd.n1530 vdd.n1518 0.155672
R21119 vdd.n1523 vdd.n1518 0.155672
R21120 vdd.n2018 vdd.n1823 0.152939
R21121 vdd.n1829 vdd.n1823 0.152939
R21122 vdd.n1830 vdd.n1829 0.152939
R21123 vdd.n1831 vdd.n1830 0.152939
R21124 vdd.n1832 vdd.n1831 0.152939
R21125 vdd.n1836 vdd.n1832 0.152939
R21126 vdd.n1837 vdd.n1836 0.152939
R21127 vdd.n1838 vdd.n1837 0.152939
R21128 vdd.n1839 vdd.n1838 0.152939
R21129 vdd.n1843 vdd.n1839 0.152939
R21130 vdd.n1844 vdd.n1843 0.152939
R21131 vdd.n1845 vdd.n1844 0.152939
R21132 vdd.n1993 vdd.n1845 0.152939
R21133 vdd.n1993 vdd.n1992 0.152939
R21134 vdd.n1992 vdd.n1991 0.152939
R21135 vdd.n1991 vdd.n1851 0.152939
R21136 vdd.n1856 vdd.n1851 0.152939
R21137 vdd.n1857 vdd.n1856 0.152939
R21138 vdd.n1858 vdd.n1857 0.152939
R21139 vdd.n1862 vdd.n1858 0.152939
R21140 vdd.n1863 vdd.n1862 0.152939
R21141 vdd.n1864 vdd.n1863 0.152939
R21142 vdd.n1865 vdd.n1864 0.152939
R21143 vdd.n1869 vdd.n1865 0.152939
R21144 vdd.n1870 vdd.n1869 0.152939
R21145 vdd.n1871 vdd.n1870 0.152939
R21146 vdd.n1872 vdd.n1871 0.152939
R21147 vdd.n1876 vdd.n1872 0.152939
R21148 vdd.n1877 vdd.n1876 0.152939
R21149 vdd.n1878 vdd.n1877 0.152939
R21150 vdd.n1879 vdd.n1878 0.152939
R21151 vdd.n1883 vdd.n1879 0.152939
R21152 vdd.n1884 vdd.n1883 0.152939
R21153 vdd.n1885 vdd.n1884 0.152939
R21154 vdd.n1954 vdd.n1885 0.152939
R21155 vdd.n1954 vdd.n1953 0.152939
R21156 vdd.n1953 vdd.n1952 0.152939
R21157 vdd.n1952 vdd.n1891 0.152939
R21158 vdd.n1896 vdd.n1891 0.152939
R21159 vdd.n1897 vdd.n1896 0.152939
R21160 vdd.n1898 vdd.n1897 0.152939
R21161 vdd.n1902 vdd.n1898 0.152939
R21162 vdd.n1903 vdd.n1902 0.152939
R21163 vdd.n1904 vdd.n1903 0.152939
R21164 vdd.n1905 vdd.n1904 0.152939
R21165 vdd.n1909 vdd.n1905 0.152939
R21166 vdd.n1910 vdd.n1909 0.152939
R21167 vdd.n1911 vdd.n1910 0.152939
R21168 vdd.n1912 vdd.n1911 0.152939
R21169 vdd.n1913 vdd.n1912 0.152939
R21170 vdd.n1913 vdd.n1035 0.152939
R21171 vdd.n2242 vdd.n1817 0.152939
R21172 vdd.n1749 vdd.n1748 0.152939
R21173 vdd.n1749 vdd.n1084 0.152939
R21174 vdd.n1763 vdd.n1084 0.152939
R21175 vdd.n1764 vdd.n1763 0.152939
R21176 vdd.n1765 vdd.n1764 0.152939
R21177 vdd.n1765 vdd.n1072 0.152939
R21178 vdd.n1780 vdd.n1072 0.152939
R21179 vdd.n1781 vdd.n1780 0.152939
R21180 vdd.n1782 vdd.n1781 0.152939
R21181 vdd.n1782 vdd.n1061 0.152939
R21182 vdd.n1797 vdd.n1061 0.152939
R21183 vdd.n1798 vdd.n1797 0.152939
R21184 vdd.n1799 vdd.n1798 0.152939
R21185 vdd.n1799 vdd.n1049 0.152939
R21186 vdd.n1815 vdd.n1049 0.152939
R21187 vdd.n1816 vdd.n1815 0.152939
R21188 vdd.n2243 vdd.n1816 0.152939
R21189 vdd.n670 vdd.n667 0.152939
R21190 vdd.n671 vdd.n670 0.152939
R21191 vdd.n672 vdd.n671 0.152939
R21192 vdd.n673 vdd.n672 0.152939
R21193 vdd.n676 vdd.n673 0.152939
R21194 vdd.n677 vdd.n676 0.152939
R21195 vdd.n678 vdd.n677 0.152939
R21196 vdd.n679 vdd.n678 0.152939
R21197 vdd.n682 vdd.n679 0.152939
R21198 vdd.n683 vdd.n682 0.152939
R21199 vdd.n684 vdd.n683 0.152939
R21200 vdd.n685 vdd.n684 0.152939
R21201 vdd.n690 vdd.n685 0.152939
R21202 vdd.n691 vdd.n690 0.152939
R21203 vdd.n692 vdd.n691 0.152939
R21204 vdd.n693 vdd.n692 0.152939
R21205 vdd.n696 vdd.n693 0.152939
R21206 vdd.n697 vdd.n696 0.152939
R21207 vdd.n698 vdd.n697 0.152939
R21208 vdd.n699 vdd.n698 0.152939
R21209 vdd.n702 vdd.n699 0.152939
R21210 vdd.n703 vdd.n702 0.152939
R21211 vdd.n704 vdd.n703 0.152939
R21212 vdd.n705 vdd.n704 0.152939
R21213 vdd.n708 vdd.n705 0.152939
R21214 vdd.n709 vdd.n708 0.152939
R21215 vdd.n710 vdd.n709 0.152939
R21216 vdd.n711 vdd.n710 0.152939
R21217 vdd.n714 vdd.n711 0.152939
R21218 vdd.n715 vdd.n714 0.152939
R21219 vdd.n716 vdd.n715 0.152939
R21220 vdd.n717 vdd.n716 0.152939
R21221 vdd.n720 vdd.n717 0.152939
R21222 vdd.n721 vdd.n720 0.152939
R21223 vdd.n3058 vdd.n721 0.152939
R21224 vdd.n3058 vdd.n3057 0.152939
R21225 vdd.n3057 vdd.n3056 0.152939
R21226 vdd.n3056 vdd.n725 0.152939
R21227 vdd.n730 vdd.n725 0.152939
R21228 vdd.n731 vdd.n730 0.152939
R21229 vdd.n734 vdd.n731 0.152939
R21230 vdd.n735 vdd.n734 0.152939
R21231 vdd.n736 vdd.n735 0.152939
R21232 vdd.n737 vdd.n736 0.152939
R21233 vdd.n740 vdd.n737 0.152939
R21234 vdd.n741 vdd.n740 0.152939
R21235 vdd.n742 vdd.n741 0.152939
R21236 vdd.n743 vdd.n742 0.152939
R21237 vdd.n746 vdd.n743 0.152939
R21238 vdd.n747 vdd.n746 0.152939
R21239 vdd.n748 vdd.n747 0.152939
R21240 vdd.n3141 vdd.n661 0.152939
R21241 vdd.n3142 vdd.n651 0.152939
R21242 vdd.n3156 vdd.n651 0.152939
R21243 vdd.n3157 vdd.n3156 0.152939
R21244 vdd.n3158 vdd.n3157 0.152939
R21245 vdd.n3158 vdd.n639 0.152939
R21246 vdd.n3172 vdd.n639 0.152939
R21247 vdd.n3173 vdd.n3172 0.152939
R21248 vdd.n3174 vdd.n3173 0.152939
R21249 vdd.n3174 vdd.n627 0.152939
R21250 vdd.n3189 vdd.n627 0.152939
R21251 vdd.n3190 vdd.n3189 0.152939
R21252 vdd.n3191 vdd.n3190 0.152939
R21253 vdd.n3191 vdd.n616 0.152939
R21254 vdd.n3208 vdd.n616 0.152939
R21255 vdd.n3209 vdd.n3208 0.152939
R21256 vdd.n3210 vdd.n3209 0.152939
R21257 vdd.n3210 vdd.n322 0.152939
R21258 vdd.n3290 vdd.n323 0.152939
R21259 vdd.n334 vdd.n323 0.152939
R21260 vdd.n335 vdd.n334 0.152939
R21261 vdd.n336 vdd.n335 0.152939
R21262 vdd.n343 vdd.n336 0.152939
R21263 vdd.n344 vdd.n343 0.152939
R21264 vdd.n345 vdd.n344 0.152939
R21265 vdd.n346 vdd.n345 0.152939
R21266 vdd.n354 vdd.n346 0.152939
R21267 vdd.n355 vdd.n354 0.152939
R21268 vdd.n356 vdd.n355 0.152939
R21269 vdd.n357 vdd.n356 0.152939
R21270 vdd.n365 vdd.n357 0.152939
R21271 vdd.n366 vdd.n365 0.152939
R21272 vdd.n367 vdd.n366 0.152939
R21273 vdd.n368 vdd.n367 0.152939
R21274 vdd.n443 vdd.n368 0.152939
R21275 vdd.n444 vdd.n442 0.152939
R21276 vdd.n451 vdd.n442 0.152939
R21277 vdd.n452 vdd.n451 0.152939
R21278 vdd.n453 vdd.n452 0.152939
R21279 vdd.n453 vdd.n440 0.152939
R21280 vdd.n461 vdd.n440 0.152939
R21281 vdd.n462 vdd.n461 0.152939
R21282 vdd.n463 vdd.n462 0.152939
R21283 vdd.n463 vdd.n438 0.152939
R21284 vdd.n471 vdd.n438 0.152939
R21285 vdd.n472 vdd.n471 0.152939
R21286 vdd.n473 vdd.n472 0.152939
R21287 vdd.n473 vdd.n436 0.152939
R21288 vdd.n481 vdd.n436 0.152939
R21289 vdd.n482 vdd.n481 0.152939
R21290 vdd.n483 vdd.n482 0.152939
R21291 vdd.n483 vdd.n434 0.152939
R21292 vdd.n491 vdd.n434 0.152939
R21293 vdd.n492 vdd.n491 0.152939
R21294 vdd.n493 vdd.n492 0.152939
R21295 vdd.n493 vdd.n430 0.152939
R21296 vdd.n501 vdd.n430 0.152939
R21297 vdd.n502 vdd.n501 0.152939
R21298 vdd.n503 vdd.n502 0.152939
R21299 vdd.n503 vdd.n428 0.152939
R21300 vdd.n511 vdd.n428 0.152939
R21301 vdd.n512 vdd.n511 0.152939
R21302 vdd.n513 vdd.n512 0.152939
R21303 vdd.n513 vdd.n426 0.152939
R21304 vdd.n521 vdd.n426 0.152939
R21305 vdd.n522 vdd.n521 0.152939
R21306 vdd.n523 vdd.n522 0.152939
R21307 vdd.n523 vdd.n424 0.152939
R21308 vdd.n531 vdd.n424 0.152939
R21309 vdd.n532 vdd.n531 0.152939
R21310 vdd.n533 vdd.n532 0.152939
R21311 vdd.n533 vdd.n422 0.152939
R21312 vdd.n541 vdd.n422 0.152939
R21313 vdd.n542 vdd.n541 0.152939
R21314 vdd.n543 vdd.n542 0.152939
R21315 vdd.n543 vdd.n418 0.152939
R21316 vdd.n551 vdd.n418 0.152939
R21317 vdd.n552 vdd.n551 0.152939
R21318 vdd.n553 vdd.n552 0.152939
R21319 vdd.n553 vdd.n416 0.152939
R21320 vdd.n561 vdd.n416 0.152939
R21321 vdd.n562 vdd.n561 0.152939
R21322 vdd.n563 vdd.n562 0.152939
R21323 vdd.n563 vdd.n414 0.152939
R21324 vdd.n571 vdd.n414 0.152939
R21325 vdd.n572 vdd.n571 0.152939
R21326 vdd.n573 vdd.n572 0.152939
R21327 vdd.n573 vdd.n412 0.152939
R21328 vdd.n581 vdd.n412 0.152939
R21329 vdd.n582 vdd.n581 0.152939
R21330 vdd.n583 vdd.n582 0.152939
R21331 vdd.n583 vdd.n410 0.152939
R21332 vdd.n591 vdd.n410 0.152939
R21333 vdd.n592 vdd.n591 0.152939
R21334 vdd.n593 vdd.n592 0.152939
R21335 vdd.n593 vdd.n408 0.152939
R21336 vdd.n600 vdd.n408 0.152939
R21337 vdd.n3249 vdd.n600 0.152939
R21338 vdd.n3149 vdd.n3148 0.152939
R21339 vdd.n3150 vdd.n3149 0.152939
R21340 vdd.n3150 vdd.n645 0.152939
R21341 vdd.n3164 vdd.n645 0.152939
R21342 vdd.n3165 vdd.n3164 0.152939
R21343 vdd.n3166 vdd.n3165 0.152939
R21344 vdd.n3166 vdd.n632 0.152939
R21345 vdd.n3180 vdd.n632 0.152939
R21346 vdd.n3181 vdd.n3180 0.152939
R21347 vdd.n3182 vdd.n3181 0.152939
R21348 vdd.n3182 vdd.n621 0.152939
R21349 vdd.n3197 vdd.n621 0.152939
R21350 vdd.n3198 vdd.n3197 0.152939
R21351 vdd.n3199 vdd.n3198 0.152939
R21352 vdd.n3201 vdd.n3199 0.152939
R21353 vdd.n3201 vdd.n3200 0.152939
R21354 vdd.n3200 vdd.n611 0.152939
R21355 vdd.n611 vdd.n609 0.152939
R21356 vdd.n3219 vdd.n609 0.152939
R21357 vdd.n3220 vdd.n3219 0.152939
R21358 vdd.n3221 vdd.n3220 0.152939
R21359 vdd.n3221 vdd.n607 0.152939
R21360 vdd.n3226 vdd.n607 0.152939
R21361 vdd.n3227 vdd.n3226 0.152939
R21362 vdd.n3228 vdd.n3227 0.152939
R21363 vdd.n3228 vdd.n605 0.152939
R21364 vdd.n3233 vdd.n605 0.152939
R21365 vdd.n3234 vdd.n3233 0.152939
R21366 vdd.n3235 vdd.n3234 0.152939
R21367 vdd.n3235 vdd.n603 0.152939
R21368 vdd.n3241 vdd.n603 0.152939
R21369 vdd.n3242 vdd.n3241 0.152939
R21370 vdd.n3243 vdd.n3242 0.152939
R21371 vdd.n3243 vdd.n601 0.152939
R21372 vdd.n3248 vdd.n601 0.152939
R21373 vdd.n3011 vdd.n656 0.152939
R21374 vdd.n2254 vdd.n1038 0.152939
R21375 vdd.n1379 vdd.n1378 0.152939
R21376 vdd.n1379 vdd.n1135 0.152939
R21377 vdd.n1393 vdd.n1135 0.152939
R21378 vdd.n1394 vdd.n1393 0.152939
R21379 vdd.n1395 vdd.n1394 0.152939
R21380 vdd.n1395 vdd.n1123 0.152939
R21381 vdd.n1410 vdd.n1123 0.152939
R21382 vdd.n1411 vdd.n1410 0.152939
R21383 vdd.n1412 vdd.n1411 0.152939
R21384 vdd.n1412 vdd.n1113 0.152939
R21385 vdd.n1427 vdd.n1113 0.152939
R21386 vdd.n1428 vdd.n1427 0.152939
R21387 vdd.n1429 vdd.n1428 0.152939
R21388 vdd.n1429 vdd.n1100 0.152939
R21389 vdd.n1443 vdd.n1100 0.152939
R21390 vdd.n1444 vdd.n1443 0.152939
R21391 vdd.n1445 vdd.n1444 0.152939
R21392 vdd.n1445 vdd.n1089 0.152939
R21393 vdd.n1755 vdd.n1089 0.152939
R21394 vdd.n1756 vdd.n1755 0.152939
R21395 vdd.n1757 vdd.n1756 0.152939
R21396 vdd.n1757 vdd.n1078 0.152939
R21397 vdd.n1771 vdd.n1078 0.152939
R21398 vdd.n1772 vdd.n1771 0.152939
R21399 vdd.n1773 vdd.n1772 0.152939
R21400 vdd.n1773 vdd.n1066 0.152939
R21401 vdd.n1788 vdd.n1066 0.152939
R21402 vdd.n1789 vdd.n1788 0.152939
R21403 vdd.n1790 vdd.n1789 0.152939
R21404 vdd.n1790 vdd.n1056 0.152939
R21405 vdd.n1805 vdd.n1056 0.152939
R21406 vdd.n1806 vdd.n1805 0.152939
R21407 vdd.n1809 vdd.n1806 0.152939
R21408 vdd.n1809 vdd.n1808 0.152939
R21409 vdd.n1808 vdd.n1807 0.152939
R21410 vdd.n1369 vdd.n1184 0.152939
R21411 vdd.n1369 vdd.n1368 0.152939
R21412 vdd.n1368 vdd.n1367 0.152939
R21413 vdd.n1367 vdd.n1186 0.152939
R21414 vdd.n1363 vdd.n1186 0.152939
R21415 vdd.n1363 vdd.n1362 0.152939
R21416 vdd.n1362 vdd.n1361 0.152939
R21417 vdd.n1361 vdd.n1191 0.152939
R21418 vdd.n1357 vdd.n1191 0.152939
R21419 vdd.n1357 vdd.n1356 0.152939
R21420 vdd.n1356 vdd.n1355 0.152939
R21421 vdd.n1355 vdd.n1197 0.152939
R21422 vdd.n1351 vdd.n1197 0.152939
R21423 vdd.n1351 vdd.n1350 0.152939
R21424 vdd.n1350 vdd.n1349 0.152939
R21425 vdd.n1349 vdd.n1203 0.152939
R21426 vdd.n1345 vdd.n1203 0.152939
R21427 vdd.n1345 vdd.n1344 0.152939
R21428 vdd.n1344 vdd.n1343 0.152939
R21429 vdd.n1343 vdd.n1209 0.152939
R21430 vdd.n1335 vdd.n1209 0.152939
R21431 vdd.n1335 vdd.n1334 0.152939
R21432 vdd.n1334 vdd.n1333 0.152939
R21433 vdd.n1333 vdd.n1213 0.152939
R21434 vdd.n1329 vdd.n1213 0.152939
R21435 vdd.n1329 vdd.n1328 0.152939
R21436 vdd.n1328 vdd.n1327 0.152939
R21437 vdd.n1327 vdd.n1219 0.152939
R21438 vdd.n1323 vdd.n1219 0.152939
R21439 vdd.n1323 vdd.n1322 0.152939
R21440 vdd.n1322 vdd.n1321 0.152939
R21441 vdd.n1321 vdd.n1225 0.152939
R21442 vdd.n1317 vdd.n1225 0.152939
R21443 vdd.n1317 vdd.n1316 0.152939
R21444 vdd.n1316 vdd.n1315 0.152939
R21445 vdd.n1315 vdd.n1231 0.152939
R21446 vdd.n1311 vdd.n1231 0.152939
R21447 vdd.n1311 vdd.n1310 0.152939
R21448 vdd.n1310 vdd.n1309 0.152939
R21449 vdd.n1309 vdd.n1237 0.152939
R21450 vdd.n1302 vdd.n1237 0.152939
R21451 vdd.n1302 vdd.n1301 0.152939
R21452 vdd.n1301 vdd.n1300 0.152939
R21453 vdd.n1300 vdd.n1242 0.152939
R21454 vdd.n1296 vdd.n1242 0.152939
R21455 vdd.n1296 vdd.n1295 0.152939
R21456 vdd.n1295 vdd.n1294 0.152939
R21457 vdd.n1294 vdd.n1248 0.152939
R21458 vdd.n1290 vdd.n1248 0.152939
R21459 vdd.n1290 vdd.n1289 0.152939
R21460 vdd.n1289 vdd.n1288 0.152939
R21461 vdd.n1288 vdd.n1254 0.152939
R21462 vdd.n1284 vdd.n1254 0.152939
R21463 vdd.n1284 vdd.n1283 0.152939
R21464 vdd.n1283 vdd.n1282 0.152939
R21465 vdd.n1282 vdd.n1260 0.152939
R21466 vdd.n1278 vdd.n1260 0.152939
R21467 vdd.n1278 vdd.n1277 0.152939
R21468 vdd.n1277 vdd.n1276 0.152939
R21469 vdd.n1276 vdd.n1266 0.152939
R21470 vdd.n1272 vdd.n1266 0.152939
R21471 vdd.n1272 vdd.n1147 0.152939
R21472 vdd.n1377 vdd.n1147 0.152939
R21473 vdd.n1385 vdd.n1141 0.152939
R21474 vdd.n1386 vdd.n1385 0.152939
R21475 vdd.n1387 vdd.n1386 0.152939
R21476 vdd.n1387 vdd.n1129 0.152939
R21477 vdd.n1402 vdd.n1129 0.152939
R21478 vdd.n1403 vdd.n1402 0.152939
R21479 vdd.n1404 vdd.n1403 0.152939
R21480 vdd.n1404 vdd.n1118 0.152939
R21481 vdd.n1419 vdd.n1118 0.152939
R21482 vdd.n1420 vdd.n1419 0.152939
R21483 vdd.n1421 vdd.n1420 0.152939
R21484 vdd.n1421 vdd.n1107 0.152939
R21485 vdd.n1435 vdd.n1107 0.152939
R21486 vdd.n1436 vdd.n1435 0.152939
R21487 vdd.n1437 vdd.n1436 0.152939
R21488 vdd.n1437 vdd.n1095 0.152939
R21489 vdd.n1452 vdd.n1095 0.152939
R21490 vdd.n2232 vdd.n1817 0.110256
R21491 vdd.n2942 vdd.n661 0.110256
R21492 vdd.n3011 vdd.n3010 0.110256
R21493 vdd.n2255 vdd.n2254 0.110256
R21494 vdd.n1748 vdd.n1747 0.0695946
R21495 vdd.n3291 vdd.n322 0.0695946
R21496 vdd.n3291 vdd.n3290 0.0695946
R21497 vdd.n1747 vdd.n1452 0.0695946
R21498 vdd.n2232 vdd.n2018 0.0431829
R21499 vdd.n2255 vdd.n1035 0.0431829
R21500 vdd.n2942 vdd.n667 0.0431829
R21501 vdd.n3010 vdd.n748 0.0431829
R21502 vdd vdd.n28 0.00833333
R21503 CSoutput.n19 CSoutput.t206 184.661
R21504 CSoutput.n78 CSoutput.n77 165.8
R21505 CSoutput.n76 CSoutput.n0 165.8
R21506 CSoutput.n75 CSoutput.n74 165.8
R21507 CSoutput.n73 CSoutput.n72 165.8
R21508 CSoutput.n71 CSoutput.n2 165.8
R21509 CSoutput.n69 CSoutput.n68 165.8
R21510 CSoutput.n67 CSoutput.n3 165.8
R21511 CSoutput.n66 CSoutput.n65 165.8
R21512 CSoutput.n63 CSoutput.n4 165.8
R21513 CSoutput.n61 CSoutput.n60 165.8
R21514 CSoutput.n59 CSoutput.n5 165.8
R21515 CSoutput.n58 CSoutput.n57 165.8
R21516 CSoutput.n55 CSoutput.n6 165.8
R21517 CSoutput.n54 CSoutput.n53 165.8
R21518 CSoutput.n52 CSoutput.n51 165.8
R21519 CSoutput.n50 CSoutput.n8 165.8
R21520 CSoutput.n48 CSoutput.n47 165.8
R21521 CSoutput.n46 CSoutput.n9 165.8
R21522 CSoutput.n45 CSoutput.n44 165.8
R21523 CSoutput.n42 CSoutput.n10 165.8
R21524 CSoutput.n41 CSoutput.n40 165.8
R21525 CSoutput.n39 CSoutput.n38 165.8
R21526 CSoutput.n37 CSoutput.n12 165.8
R21527 CSoutput.n35 CSoutput.n34 165.8
R21528 CSoutput.n33 CSoutput.n13 165.8
R21529 CSoutput.n32 CSoutput.n31 165.8
R21530 CSoutput.n29 CSoutput.n14 165.8
R21531 CSoutput.n28 CSoutput.n27 165.8
R21532 CSoutput.n26 CSoutput.n25 165.8
R21533 CSoutput.n24 CSoutput.n16 165.8
R21534 CSoutput.n22 CSoutput.n21 165.8
R21535 CSoutput.n20 CSoutput.n17 165.8
R21536 CSoutput.n77 CSoutput.t207 162.194
R21537 CSoutput.n18 CSoutput.t208 120.501
R21538 CSoutput.n23 CSoutput.t196 120.501
R21539 CSoutput.n15 CSoutput.t194 120.501
R21540 CSoutput.n30 CSoutput.t210 120.501
R21541 CSoutput.n36 CSoutput.t198 120.501
R21542 CSoutput.n11 CSoutput.t200 120.501
R21543 CSoutput.n43 CSoutput.t213 120.501
R21544 CSoutput.n49 CSoutput.t201 120.501
R21545 CSoutput.n7 CSoutput.t203 120.501
R21546 CSoutput.n56 CSoutput.t197 120.501
R21547 CSoutput.n62 CSoutput.t211 120.501
R21548 CSoutput.n64 CSoutput.t205 120.501
R21549 CSoutput.n70 CSoutput.t199 120.501
R21550 CSoutput.n1 CSoutput.t195 120.501
R21551 CSoutput.n310 CSoutput.n308 103.469
R21552 CSoutput.n294 CSoutput.n292 103.469
R21553 CSoutput.n279 CSoutput.n277 103.469
R21554 CSoutput.n112 CSoutput.n110 103.469
R21555 CSoutput.n96 CSoutput.n94 103.469
R21556 CSoutput.n81 CSoutput.n79 103.469
R21557 CSoutput.n320 CSoutput.n319 103.111
R21558 CSoutput.n318 CSoutput.n317 103.111
R21559 CSoutput.n316 CSoutput.n315 103.111
R21560 CSoutput.n314 CSoutput.n313 103.111
R21561 CSoutput.n312 CSoutput.n311 103.111
R21562 CSoutput.n310 CSoutput.n309 103.111
R21563 CSoutput.n306 CSoutput.n305 103.111
R21564 CSoutput.n304 CSoutput.n303 103.111
R21565 CSoutput.n302 CSoutput.n301 103.111
R21566 CSoutput.n300 CSoutput.n299 103.111
R21567 CSoutput.n298 CSoutput.n297 103.111
R21568 CSoutput.n296 CSoutput.n295 103.111
R21569 CSoutput.n294 CSoutput.n293 103.111
R21570 CSoutput.n291 CSoutput.n290 103.111
R21571 CSoutput.n289 CSoutput.n288 103.111
R21572 CSoutput.n287 CSoutput.n286 103.111
R21573 CSoutput.n285 CSoutput.n284 103.111
R21574 CSoutput.n283 CSoutput.n282 103.111
R21575 CSoutput.n281 CSoutput.n280 103.111
R21576 CSoutput.n279 CSoutput.n278 103.111
R21577 CSoutput.n112 CSoutput.n111 103.111
R21578 CSoutput.n114 CSoutput.n113 103.111
R21579 CSoutput.n116 CSoutput.n115 103.111
R21580 CSoutput.n118 CSoutput.n117 103.111
R21581 CSoutput.n120 CSoutput.n119 103.111
R21582 CSoutput.n122 CSoutput.n121 103.111
R21583 CSoutput.n124 CSoutput.n123 103.111
R21584 CSoutput.n96 CSoutput.n95 103.111
R21585 CSoutput.n98 CSoutput.n97 103.111
R21586 CSoutput.n100 CSoutput.n99 103.111
R21587 CSoutput.n102 CSoutput.n101 103.111
R21588 CSoutput.n104 CSoutput.n103 103.111
R21589 CSoutput.n106 CSoutput.n105 103.111
R21590 CSoutput.n108 CSoutput.n107 103.111
R21591 CSoutput.n81 CSoutput.n80 103.111
R21592 CSoutput.n83 CSoutput.n82 103.111
R21593 CSoutput.n85 CSoutput.n84 103.111
R21594 CSoutput.n87 CSoutput.n86 103.111
R21595 CSoutput.n89 CSoutput.n88 103.111
R21596 CSoutput.n91 CSoutput.n90 103.111
R21597 CSoutput.n93 CSoutput.n92 103.111
R21598 CSoutput.n322 CSoutput.n321 103.111
R21599 CSoutput.n358 CSoutput.n356 81.5057
R21600 CSoutput.n342 CSoutput.n340 81.5057
R21601 CSoutput.n327 CSoutput.n325 81.5057
R21602 CSoutput.n406 CSoutput.n404 81.5057
R21603 CSoutput.n390 CSoutput.n388 81.5057
R21604 CSoutput.n375 CSoutput.n373 81.5057
R21605 CSoutput.n370 CSoutput.n369 80.9324
R21606 CSoutput.n368 CSoutput.n367 80.9324
R21607 CSoutput.n366 CSoutput.n365 80.9324
R21608 CSoutput.n364 CSoutput.n363 80.9324
R21609 CSoutput.n362 CSoutput.n361 80.9324
R21610 CSoutput.n360 CSoutput.n359 80.9324
R21611 CSoutput.n358 CSoutput.n357 80.9324
R21612 CSoutput.n354 CSoutput.n353 80.9324
R21613 CSoutput.n352 CSoutput.n351 80.9324
R21614 CSoutput.n350 CSoutput.n349 80.9324
R21615 CSoutput.n348 CSoutput.n347 80.9324
R21616 CSoutput.n346 CSoutput.n345 80.9324
R21617 CSoutput.n344 CSoutput.n343 80.9324
R21618 CSoutput.n342 CSoutput.n341 80.9324
R21619 CSoutput.n339 CSoutput.n338 80.9324
R21620 CSoutput.n337 CSoutput.n336 80.9324
R21621 CSoutput.n335 CSoutput.n334 80.9324
R21622 CSoutput.n333 CSoutput.n332 80.9324
R21623 CSoutput.n331 CSoutput.n330 80.9324
R21624 CSoutput.n329 CSoutput.n328 80.9324
R21625 CSoutput.n327 CSoutput.n326 80.9324
R21626 CSoutput.n406 CSoutput.n405 80.9324
R21627 CSoutput.n408 CSoutput.n407 80.9324
R21628 CSoutput.n410 CSoutput.n409 80.9324
R21629 CSoutput.n412 CSoutput.n411 80.9324
R21630 CSoutput.n414 CSoutput.n413 80.9324
R21631 CSoutput.n416 CSoutput.n415 80.9324
R21632 CSoutput.n418 CSoutput.n417 80.9324
R21633 CSoutput.n390 CSoutput.n389 80.9324
R21634 CSoutput.n392 CSoutput.n391 80.9324
R21635 CSoutput.n394 CSoutput.n393 80.9324
R21636 CSoutput.n396 CSoutput.n395 80.9324
R21637 CSoutput.n398 CSoutput.n397 80.9324
R21638 CSoutput.n400 CSoutput.n399 80.9324
R21639 CSoutput.n402 CSoutput.n401 80.9324
R21640 CSoutput.n375 CSoutput.n374 80.9324
R21641 CSoutput.n377 CSoutput.n376 80.9324
R21642 CSoutput.n379 CSoutput.n378 80.9324
R21643 CSoutput.n381 CSoutput.n380 80.9324
R21644 CSoutput.n383 CSoutput.n382 80.9324
R21645 CSoutput.n385 CSoutput.n384 80.9324
R21646 CSoutput.n387 CSoutput.n386 80.9324
R21647 CSoutput.n25 CSoutput.n24 48.1486
R21648 CSoutput.n69 CSoutput.n3 48.1486
R21649 CSoutput.n38 CSoutput.n37 48.1486
R21650 CSoutput.n42 CSoutput.n41 48.1486
R21651 CSoutput.n51 CSoutput.n50 48.1486
R21652 CSoutput.n55 CSoutput.n54 48.1486
R21653 CSoutput.n22 CSoutput.n17 46.462
R21654 CSoutput.n72 CSoutput.n71 46.462
R21655 CSoutput.n20 CSoutput.n19 44.9055
R21656 CSoutput.n29 CSoutput.n28 43.7635
R21657 CSoutput.n65 CSoutput.n63 43.7635
R21658 CSoutput.n35 CSoutput.n13 41.7396
R21659 CSoutput.n57 CSoutput.n5 41.7396
R21660 CSoutput.n44 CSoutput.n9 37.0171
R21661 CSoutput.n48 CSoutput.n9 37.0171
R21662 CSoutput.n76 CSoutput.n75 34.9932
R21663 CSoutput.n31 CSoutput.n13 32.2947
R21664 CSoutput.n61 CSoutput.n5 32.2947
R21665 CSoutput.n30 CSoutput.n29 29.6014
R21666 CSoutput.n63 CSoutput.n62 29.6014
R21667 CSoutput.n19 CSoutput.n18 28.4085
R21668 CSoutput.n18 CSoutput.n17 25.1176
R21669 CSoutput.n72 CSoutput.n1 25.1176
R21670 CSoutput.n43 CSoutput.n42 22.0922
R21671 CSoutput.n50 CSoutput.n49 22.0922
R21672 CSoutput.n77 CSoutput.n76 21.8586
R21673 CSoutput.n37 CSoutput.n36 18.9681
R21674 CSoutput.n56 CSoutput.n55 18.9681
R21675 CSoutput.n25 CSoutput.n15 17.6292
R21676 CSoutput.n64 CSoutput.n3 17.6292
R21677 CSoutput.n24 CSoutput.n23 15.844
R21678 CSoutput.n70 CSoutput.n69 15.844
R21679 CSoutput.n38 CSoutput.n11 14.5051
R21680 CSoutput.n54 CSoutput.n7 14.5051
R21681 CSoutput.n421 CSoutput.n78 11.4982
R21682 CSoutput.n41 CSoutput.n11 11.3811
R21683 CSoutput.n51 CSoutput.n7 11.3811
R21684 CSoutput.n23 CSoutput.n22 10.0422
R21685 CSoutput.n71 CSoutput.n70 10.0422
R21686 CSoutput.n307 CSoutput.n291 9.25285
R21687 CSoutput.n109 CSoutput.n93 9.25285
R21688 CSoutput.n372 CSoutput.n324 9.03201
R21689 CSoutput.n355 CSoutput.n339 8.98182
R21690 CSoutput.n403 CSoutput.n387 8.98182
R21691 CSoutput.n28 CSoutput.n15 8.25698
R21692 CSoutput.n65 CSoutput.n64 8.25698
R21693 CSoutput.n324 CSoutput.n323 7.12641
R21694 CSoutput.n126 CSoutput.n125 7.12641
R21695 CSoutput.n36 CSoutput.n35 6.91809
R21696 CSoutput.n57 CSoutput.n56 6.91809
R21697 CSoutput.n372 CSoutput.n371 6.02792
R21698 CSoutput.n420 CSoutput.n419 6.02792
R21699 CSoutput.n421 CSoutput.n126 5.43957
R21700 CSoutput.n371 CSoutput.n370 5.25266
R21701 CSoutput.n355 CSoutput.n354 5.25266
R21702 CSoutput.n419 CSoutput.n418 5.25266
R21703 CSoutput.n403 CSoutput.n402 5.25266
R21704 CSoutput.n323 CSoutput.n322 5.1449
R21705 CSoutput.n307 CSoutput.n306 5.1449
R21706 CSoutput.n125 CSoutput.n124 5.1449
R21707 CSoutput.n109 CSoutput.n108 5.1449
R21708 CSoutput.n217 CSoutput.n170 4.5005
R21709 CSoutput.n186 CSoutput.n170 4.5005
R21710 CSoutput.n181 CSoutput.n165 4.5005
R21711 CSoutput.n181 CSoutput.n167 4.5005
R21712 CSoutput.n181 CSoutput.n164 4.5005
R21713 CSoutput.n181 CSoutput.n168 4.5005
R21714 CSoutput.n181 CSoutput.n163 4.5005
R21715 CSoutput.n181 CSoutput.t209 4.5005
R21716 CSoutput.n181 CSoutput.n162 4.5005
R21717 CSoutput.n181 CSoutput.n169 4.5005
R21718 CSoutput.n181 CSoutput.n170 4.5005
R21719 CSoutput.n179 CSoutput.n165 4.5005
R21720 CSoutput.n179 CSoutput.n167 4.5005
R21721 CSoutput.n179 CSoutput.n164 4.5005
R21722 CSoutput.n179 CSoutput.n168 4.5005
R21723 CSoutput.n179 CSoutput.n163 4.5005
R21724 CSoutput.n179 CSoutput.t209 4.5005
R21725 CSoutput.n179 CSoutput.n162 4.5005
R21726 CSoutput.n179 CSoutput.n169 4.5005
R21727 CSoutput.n179 CSoutput.n170 4.5005
R21728 CSoutput.n178 CSoutput.n165 4.5005
R21729 CSoutput.n178 CSoutput.n167 4.5005
R21730 CSoutput.n178 CSoutput.n164 4.5005
R21731 CSoutput.n178 CSoutput.n168 4.5005
R21732 CSoutput.n178 CSoutput.n163 4.5005
R21733 CSoutput.n178 CSoutput.t209 4.5005
R21734 CSoutput.n178 CSoutput.n162 4.5005
R21735 CSoutput.n178 CSoutput.n169 4.5005
R21736 CSoutput.n178 CSoutput.n170 4.5005
R21737 CSoutput.n263 CSoutput.n165 4.5005
R21738 CSoutput.n263 CSoutput.n167 4.5005
R21739 CSoutput.n263 CSoutput.n164 4.5005
R21740 CSoutput.n263 CSoutput.n168 4.5005
R21741 CSoutput.n263 CSoutput.n163 4.5005
R21742 CSoutput.n263 CSoutput.t209 4.5005
R21743 CSoutput.n263 CSoutput.n162 4.5005
R21744 CSoutput.n263 CSoutput.n169 4.5005
R21745 CSoutput.n263 CSoutput.n170 4.5005
R21746 CSoutput.n261 CSoutput.n165 4.5005
R21747 CSoutput.n261 CSoutput.n167 4.5005
R21748 CSoutput.n261 CSoutput.n164 4.5005
R21749 CSoutput.n261 CSoutput.n168 4.5005
R21750 CSoutput.n261 CSoutput.n163 4.5005
R21751 CSoutput.n261 CSoutput.t209 4.5005
R21752 CSoutput.n261 CSoutput.n162 4.5005
R21753 CSoutput.n261 CSoutput.n169 4.5005
R21754 CSoutput.n259 CSoutput.n165 4.5005
R21755 CSoutput.n259 CSoutput.n167 4.5005
R21756 CSoutput.n259 CSoutput.n164 4.5005
R21757 CSoutput.n259 CSoutput.n168 4.5005
R21758 CSoutput.n259 CSoutput.n163 4.5005
R21759 CSoutput.n259 CSoutput.t209 4.5005
R21760 CSoutput.n259 CSoutput.n162 4.5005
R21761 CSoutput.n259 CSoutput.n169 4.5005
R21762 CSoutput.n189 CSoutput.n165 4.5005
R21763 CSoutput.n189 CSoutput.n167 4.5005
R21764 CSoutput.n189 CSoutput.n164 4.5005
R21765 CSoutput.n189 CSoutput.n168 4.5005
R21766 CSoutput.n189 CSoutput.n163 4.5005
R21767 CSoutput.n189 CSoutput.t209 4.5005
R21768 CSoutput.n189 CSoutput.n162 4.5005
R21769 CSoutput.n189 CSoutput.n169 4.5005
R21770 CSoutput.n189 CSoutput.n170 4.5005
R21771 CSoutput.n188 CSoutput.n165 4.5005
R21772 CSoutput.n188 CSoutput.n167 4.5005
R21773 CSoutput.n188 CSoutput.n164 4.5005
R21774 CSoutput.n188 CSoutput.n168 4.5005
R21775 CSoutput.n188 CSoutput.n163 4.5005
R21776 CSoutput.n188 CSoutput.t209 4.5005
R21777 CSoutput.n188 CSoutput.n162 4.5005
R21778 CSoutput.n188 CSoutput.n169 4.5005
R21779 CSoutput.n188 CSoutput.n170 4.5005
R21780 CSoutput.n192 CSoutput.n165 4.5005
R21781 CSoutput.n192 CSoutput.n167 4.5005
R21782 CSoutput.n192 CSoutput.n164 4.5005
R21783 CSoutput.n192 CSoutput.n168 4.5005
R21784 CSoutput.n192 CSoutput.n163 4.5005
R21785 CSoutput.n192 CSoutput.t209 4.5005
R21786 CSoutput.n192 CSoutput.n162 4.5005
R21787 CSoutput.n192 CSoutput.n169 4.5005
R21788 CSoutput.n192 CSoutput.n170 4.5005
R21789 CSoutput.n191 CSoutput.n165 4.5005
R21790 CSoutput.n191 CSoutput.n167 4.5005
R21791 CSoutput.n191 CSoutput.n164 4.5005
R21792 CSoutput.n191 CSoutput.n168 4.5005
R21793 CSoutput.n191 CSoutput.n163 4.5005
R21794 CSoutput.n191 CSoutput.t209 4.5005
R21795 CSoutput.n191 CSoutput.n162 4.5005
R21796 CSoutput.n191 CSoutput.n169 4.5005
R21797 CSoutput.n191 CSoutput.n170 4.5005
R21798 CSoutput.n174 CSoutput.n165 4.5005
R21799 CSoutput.n174 CSoutput.n167 4.5005
R21800 CSoutput.n174 CSoutput.n164 4.5005
R21801 CSoutput.n174 CSoutput.n168 4.5005
R21802 CSoutput.n174 CSoutput.n163 4.5005
R21803 CSoutput.n174 CSoutput.t209 4.5005
R21804 CSoutput.n174 CSoutput.n162 4.5005
R21805 CSoutput.n174 CSoutput.n169 4.5005
R21806 CSoutput.n174 CSoutput.n170 4.5005
R21807 CSoutput.n266 CSoutput.n165 4.5005
R21808 CSoutput.n266 CSoutput.n167 4.5005
R21809 CSoutput.n266 CSoutput.n164 4.5005
R21810 CSoutput.n266 CSoutput.n168 4.5005
R21811 CSoutput.n266 CSoutput.n163 4.5005
R21812 CSoutput.n266 CSoutput.t209 4.5005
R21813 CSoutput.n266 CSoutput.n162 4.5005
R21814 CSoutput.n266 CSoutput.n169 4.5005
R21815 CSoutput.n266 CSoutput.n170 4.5005
R21816 CSoutput.n253 CSoutput.n224 4.5005
R21817 CSoutput.n253 CSoutput.n230 4.5005
R21818 CSoutput.n211 CSoutput.n200 4.5005
R21819 CSoutput.n211 CSoutput.n202 4.5005
R21820 CSoutput.n211 CSoutput.n199 4.5005
R21821 CSoutput.n211 CSoutput.n203 4.5005
R21822 CSoutput.n211 CSoutput.n198 4.5005
R21823 CSoutput.n211 CSoutput.t202 4.5005
R21824 CSoutput.n211 CSoutput.n197 4.5005
R21825 CSoutput.n211 CSoutput.n204 4.5005
R21826 CSoutput.n253 CSoutput.n211 4.5005
R21827 CSoutput.n232 CSoutput.n200 4.5005
R21828 CSoutput.n232 CSoutput.n202 4.5005
R21829 CSoutput.n232 CSoutput.n199 4.5005
R21830 CSoutput.n232 CSoutput.n203 4.5005
R21831 CSoutput.n232 CSoutput.n198 4.5005
R21832 CSoutput.n232 CSoutput.t202 4.5005
R21833 CSoutput.n232 CSoutput.n197 4.5005
R21834 CSoutput.n232 CSoutput.n204 4.5005
R21835 CSoutput.n253 CSoutput.n232 4.5005
R21836 CSoutput.n210 CSoutput.n200 4.5005
R21837 CSoutput.n210 CSoutput.n202 4.5005
R21838 CSoutput.n210 CSoutput.n199 4.5005
R21839 CSoutput.n210 CSoutput.n203 4.5005
R21840 CSoutput.n210 CSoutput.n198 4.5005
R21841 CSoutput.n210 CSoutput.t202 4.5005
R21842 CSoutput.n210 CSoutput.n197 4.5005
R21843 CSoutput.n210 CSoutput.n204 4.5005
R21844 CSoutput.n253 CSoutput.n210 4.5005
R21845 CSoutput.n234 CSoutput.n200 4.5005
R21846 CSoutput.n234 CSoutput.n202 4.5005
R21847 CSoutput.n234 CSoutput.n199 4.5005
R21848 CSoutput.n234 CSoutput.n203 4.5005
R21849 CSoutput.n234 CSoutput.n198 4.5005
R21850 CSoutput.n234 CSoutput.t202 4.5005
R21851 CSoutput.n234 CSoutput.n197 4.5005
R21852 CSoutput.n234 CSoutput.n204 4.5005
R21853 CSoutput.n253 CSoutput.n234 4.5005
R21854 CSoutput.n200 CSoutput.n195 4.5005
R21855 CSoutput.n202 CSoutput.n195 4.5005
R21856 CSoutput.n199 CSoutput.n195 4.5005
R21857 CSoutput.n203 CSoutput.n195 4.5005
R21858 CSoutput.n198 CSoutput.n195 4.5005
R21859 CSoutput.t202 CSoutput.n195 4.5005
R21860 CSoutput.n197 CSoutput.n195 4.5005
R21861 CSoutput.n204 CSoutput.n195 4.5005
R21862 CSoutput.n256 CSoutput.n200 4.5005
R21863 CSoutput.n256 CSoutput.n202 4.5005
R21864 CSoutput.n256 CSoutput.n199 4.5005
R21865 CSoutput.n256 CSoutput.n203 4.5005
R21866 CSoutput.n256 CSoutput.n198 4.5005
R21867 CSoutput.n256 CSoutput.t202 4.5005
R21868 CSoutput.n256 CSoutput.n197 4.5005
R21869 CSoutput.n256 CSoutput.n204 4.5005
R21870 CSoutput.n254 CSoutput.n200 4.5005
R21871 CSoutput.n254 CSoutput.n202 4.5005
R21872 CSoutput.n254 CSoutput.n199 4.5005
R21873 CSoutput.n254 CSoutput.n203 4.5005
R21874 CSoutput.n254 CSoutput.n198 4.5005
R21875 CSoutput.n254 CSoutput.t202 4.5005
R21876 CSoutput.n254 CSoutput.n197 4.5005
R21877 CSoutput.n254 CSoutput.n204 4.5005
R21878 CSoutput.n254 CSoutput.n253 4.5005
R21879 CSoutput.n236 CSoutput.n200 4.5005
R21880 CSoutput.n236 CSoutput.n202 4.5005
R21881 CSoutput.n236 CSoutput.n199 4.5005
R21882 CSoutput.n236 CSoutput.n203 4.5005
R21883 CSoutput.n236 CSoutput.n198 4.5005
R21884 CSoutput.n236 CSoutput.t202 4.5005
R21885 CSoutput.n236 CSoutput.n197 4.5005
R21886 CSoutput.n236 CSoutput.n204 4.5005
R21887 CSoutput.n253 CSoutput.n236 4.5005
R21888 CSoutput.n208 CSoutput.n200 4.5005
R21889 CSoutput.n208 CSoutput.n202 4.5005
R21890 CSoutput.n208 CSoutput.n199 4.5005
R21891 CSoutput.n208 CSoutput.n203 4.5005
R21892 CSoutput.n208 CSoutput.n198 4.5005
R21893 CSoutput.n208 CSoutput.t202 4.5005
R21894 CSoutput.n208 CSoutput.n197 4.5005
R21895 CSoutput.n208 CSoutput.n204 4.5005
R21896 CSoutput.n253 CSoutput.n208 4.5005
R21897 CSoutput.n238 CSoutput.n200 4.5005
R21898 CSoutput.n238 CSoutput.n202 4.5005
R21899 CSoutput.n238 CSoutput.n199 4.5005
R21900 CSoutput.n238 CSoutput.n203 4.5005
R21901 CSoutput.n238 CSoutput.n198 4.5005
R21902 CSoutput.n238 CSoutput.t202 4.5005
R21903 CSoutput.n238 CSoutput.n197 4.5005
R21904 CSoutput.n238 CSoutput.n204 4.5005
R21905 CSoutput.n253 CSoutput.n238 4.5005
R21906 CSoutput.n207 CSoutput.n200 4.5005
R21907 CSoutput.n207 CSoutput.n202 4.5005
R21908 CSoutput.n207 CSoutput.n199 4.5005
R21909 CSoutput.n207 CSoutput.n203 4.5005
R21910 CSoutput.n207 CSoutput.n198 4.5005
R21911 CSoutput.n207 CSoutput.t202 4.5005
R21912 CSoutput.n207 CSoutput.n197 4.5005
R21913 CSoutput.n207 CSoutput.n204 4.5005
R21914 CSoutput.n253 CSoutput.n207 4.5005
R21915 CSoutput.n252 CSoutput.n200 4.5005
R21916 CSoutput.n252 CSoutput.n202 4.5005
R21917 CSoutput.n252 CSoutput.n199 4.5005
R21918 CSoutput.n252 CSoutput.n203 4.5005
R21919 CSoutput.n252 CSoutput.n198 4.5005
R21920 CSoutput.n252 CSoutput.t202 4.5005
R21921 CSoutput.n252 CSoutput.n197 4.5005
R21922 CSoutput.n252 CSoutput.n204 4.5005
R21923 CSoutput.n253 CSoutput.n252 4.5005
R21924 CSoutput.n251 CSoutput.n136 4.5005
R21925 CSoutput.n152 CSoutput.n136 4.5005
R21926 CSoutput.n147 CSoutput.n131 4.5005
R21927 CSoutput.n147 CSoutput.n133 4.5005
R21928 CSoutput.n147 CSoutput.n130 4.5005
R21929 CSoutput.n147 CSoutput.n134 4.5005
R21930 CSoutput.n147 CSoutput.n129 4.5005
R21931 CSoutput.n147 CSoutput.t192 4.5005
R21932 CSoutput.n147 CSoutput.n128 4.5005
R21933 CSoutput.n147 CSoutput.n135 4.5005
R21934 CSoutput.n147 CSoutput.n136 4.5005
R21935 CSoutput.n145 CSoutput.n131 4.5005
R21936 CSoutput.n145 CSoutput.n133 4.5005
R21937 CSoutput.n145 CSoutput.n130 4.5005
R21938 CSoutput.n145 CSoutput.n134 4.5005
R21939 CSoutput.n145 CSoutput.n129 4.5005
R21940 CSoutput.n145 CSoutput.t192 4.5005
R21941 CSoutput.n145 CSoutput.n128 4.5005
R21942 CSoutput.n145 CSoutput.n135 4.5005
R21943 CSoutput.n145 CSoutput.n136 4.5005
R21944 CSoutput.n144 CSoutput.n131 4.5005
R21945 CSoutput.n144 CSoutput.n133 4.5005
R21946 CSoutput.n144 CSoutput.n130 4.5005
R21947 CSoutput.n144 CSoutput.n134 4.5005
R21948 CSoutput.n144 CSoutput.n129 4.5005
R21949 CSoutput.n144 CSoutput.t192 4.5005
R21950 CSoutput.n144 CSoutput.n128 4.5005
R21951 CSoutput.n144 CSoutput.n135 4.5005
R21952 CSoutput.n144 CSoutput.n136 4.5005
R21953 CSoutput.n273 CSoutput.n131 4.5005
R21954 CSoutput.n273 CSoutput.n133 4.5005
R21955 CSoutput.n273 CSoutput.n130 4.5005
R21956 CSoutput.n273 CSoutput.n134 4.5005
R21957 CSoutput.n273 CSoutput.n129 4.5005
R21958 CSoutput.n273 CSoutput.t192 4.5005
R21959 CSoutput.n273 CSoutput.n128 4.5005
R21960 CSoutput.n273 CSoutput.n135 4.5005
R21961 CSoutput.n273 CSoutput.n136 4.5005
R21962 CSoutput.n271 CSoutput.n131 4.5005
R21963 CSoutput.n271 CSoutput.n133 4.5005
R21964 CSoutput.n271 CSoutput.n130 4.5005
R21965 CSoutput.n271 CSoutput.n134 4.5005
R21966 CSoutput.n271 CSoutput.n129 4.5005
R21967 CSoutput.n271 CSoutput.t192 4.5005
R21968 CSoutput.n271 CSoutput.n128 4.5005
R21969 CSoutput.n271 CSoutput.n135 4.5005
R21970 CSoutput.n269 CSoutput.n131 4.5005
R21971 CSoutput.n269 CSoutput.n133 4.5005
R21972 CSoutput.n269 CSoutput.n130 4.5005
R21973 CSoutput.n269 CSoutput.n134 4.5005
R21974 CSoutput.n269 CSoutput.n129 4.5005
R21975 CSoutput.n269 CSoutput.t192 4.5005
R21976 CSoutput.n269 CSoutput.n128 4.5005
R21977 CSoutput.n269 CSoutput.n135 4.5005
R21978 CSoutput.n155 CSoutput.n131 4.5005
R21979 CSoutput.n155 CSoutput.n133 4.5005
R21980 CSoutput.n155 CSoutput.n130 4.5005
R21981 CSoutput.n155 CSoutput.n134 4.5005
R21982 CSoutput.n155 CSoutput.n129 4.5005
R21983 CSoutput.n155 CSoutput.t192 4.5005
R21984 CSoutput.n155 CSoutput.n128 4.5005
R21985 CSoutput.n155 CSoutput.n135 4.5005
R21986 CSoutput.n155 CSoutput.n136 4.5005
R21987 CSoutput.n154 CSoutput.n131 4.5005
R21988 CSoutput.n154 CSoutput.n133 4.5005
R21989 CSoutput.n154 CSoutput.n130 4.5005
R21990 CSoutput.n154 CSoutput.n134 4.5005
R21991 CSoutput.n154 CSoutput.n129 4.5005
R21992 CSoutput.n154 CSoutput.t192 4.5005
R21993 CSoutput.n154 CSoutput.n128 4.5005
R21994 CSoutput.n154 CSoutput.n135 4.5005
R21995 CSoutput.n154 CSoutput.n136 4.5005
R21996 CSoutput.n158 CSoutput.n131 4.5005
R21997 CSoutput.n158 CSoutput.n133 4.5005
R21998 CSoutput.n158 CSoutput.n130 4.5005
R21999 CSoutput.n158 CSoutput.n134 4.5005
R22000 CSoutput.n158 CSoutput.n129 4.5005
R22001 CSoutput.n158 CSoutput.t192 4.5005
R22002 CSoutput.n158 CSoutput.n128 4.5005
R22003 CSoutput.n158 CSoutput.n135 4.5005
R22004 CSoutput.n158 CSoutput.n136 4.5005
R22005 CSoutput.n157 CSoutput.n131 4.5005
R22006 CSoutput.n157 CSoutput.n133 4.5005
R22007 CSoutput.n157 CSoutput.n130 4.5005
R22008 CSoutput.n157 CSoutput.n134 4.5005
R22009 CSoutput.n157 CSoutput.n129 4.5005
R22010 CSoutput.n157 CSoutput.t192 4.5005
R22011 CSoutput.n157 CSoutput.n128 4.5005
R22012 CSoutput.n157 CSoutput.n135 4.5005
R22013 CSoutput.n157 CSoutput.n136 4.5005
R22014 CSoutput.n140 CSoutput.n131 4.5005
R22015 CSoutput.n140 CSoutput.n133 4.5005
R22016 CSoutput.n140 CSoutput.n130 4.5005
R22017 CSoutput.n140 CSoutput.n134 4.5005
R22018 CSoutput.n140 CSoutput.n129 4.5005
R22019 CSoutput.n140 CSoutput.t192 4.5005
R22020 CSoutput.n140 CSoutput.n128 4.5005
R22021 CSoutput.n140 CSoutput.n135 4.5005
R22022 CSoutput.n140 CSoutput.n136 4.5005
R22023 CSoutput.n276 CSoutput.n131 4.5005
R22024 CSoutput.n276 CSoutput.n133 4.5005
R22025 CSoutput.n276 CSoutput.n130 4.5005
R22026 CSoutput.n276 CSoutput.n134 4.5005
R22027 CSoutput.n276 CSoutput.n129 4.5005
R22028 CSoutput.n276 CSoutput.t192 4.5005
R22029 CSoutput.n276 CSoutput.n128 4.5005
R22030 CSoutput.n276 CSoutput.n135 4.5005
R22031 CSoutput.n276 CSoutput.n136 4.5005
R22032 CSoutput.n323 CSoutput.n307 4.10845
R22033 CSoutput.n125 CSoutput.n109 4.10845
R22034 CSoutput.n321 CSoutput.t20 4.06363
R22035 CSoutput.n321 CSoutput.t73 4.06363
R22036 CSoutput.n319 CSoutput.t90 4.06363
R22037 CSoutput.n319 CSoutput.t91 4.06363
R22038 CSoutput.n317 CSoutput.t33 4.06363
R22039 CSoutput.n317 CSoutput.t34 4.06363
R22040 CSoutput.n315 CSoutput.t39 4.06363
R22041 CSoutput.n315 CSoutput.t92 4.06363
R22042 CSoutput.n313 CSoutput.t12 4.06363
R22043 CSoutput.n313 CSoutput.t37 4.06363
R22044 CSoutput.n311 CSoutput.t51 4.06363
R22045 CSoutput.n311 CSoutput.t69 4.06363
R22046 CSoutput.n309 CSoutput.t75 4.06363
R22047 CSoutput.n309 CSoutput.t16 4.06363
R22048 CSoutput.n308 CSoutput.t52 4.06363
R22049 CSoutput.n308 CSoutput.t53 4.06363
R22050 CSoutput.n305 CSoutput.t9 4.06363
R22051 CSoutput.n305 CSoutput.t61 4.06363
R22052 CSoutput.n303 CSoutput.t79 4.06363
R22053 CSoutput.n303 CSoutput.t80 4.06363
R22054 CSoutput.n301 CSoutput.t24 4.06363
R22055 CSoutput.n301 CSoutput.t25 4.06363
R22056 CSoutput.n299 CSoutput.t28 4.06363
R22057 CSoutput.n299 CSoutput.t83 4.06363
R22058 CSoutput.n297 CSoutput.t0 4.06363
R22059 CSoutput.n297 CSoutput.t27 4.06363
R22060 CSoutput.n295 CSoutput.t40 4.06363
R22061 CSoutput.n295 CSoutput.t60 4.06363
R22062 CSoutput.n293 CSoutput.t62 4.06363
R22063 CSoutput.n293 CSoutput.t4 4.06363
R22064 CSoutput.n292 CSoutput.t45 4.06363
R22065 CSoutput.n292 CSoutput.t46 4.06363
R22066 CSoutput.n290 CSoutput.t77 4.06363
R22067 CSoutput.n290 CSoutput.t13 4.06363
R22068 CSoutput.n288 CSoutput.t43 4.06363
R22069 CSoutput.n288 CSoutput.t26 4.06363
R22070 CSoutput.n286 CSoutput.t29 4.06363
R22071 CSoutput.n286 CSoutput.t10 4.06363
R22072 CSoutput.n284 CSoutput.t67 4.06363
R22073 CSoutput.n284 CSoutput.t5 4.06363
R22074 CSoutput.n282 CSoutput.t35 4.06363
R22075 CSoutput.n282 CSoutput.t88 4.06363
R22076 CSoutput.n280 CSoutput.t21 4.06363
R22077 CSoutput.n280 CSoutput.t71 4.06363
R22078 CSoutput.n278 CSoutput.t41 4.06363
R22079 CSoutput.n278 CSoutput.t93 4.06363
R22080 CSoutput.n277 CSoutput.t1 4.06363
R22081 CSoutput.n277 CSoutput.t81 4.06363
R22082 CSoutput.n110 CSoutput.t87 4.06363
R22083 CSoutput.n110 CSoutput.t86 4.06363
R22084 CSoutput.n111 CSoutput.t68 4.06363
R22085 CSoutput.n111 CSoutput.t18 4.06363
R22086 CSoutput.n113 CSoutput.t15 4.06363
R22087 CSoutput.n113 CSoutput.t84 4.06363
R22088 CSoutput.n115 CSoutput.t66 4.06363
R22089 CSoutput.n115 CSoutput.t49 4.06363
R22090 CSoutput.n117 CSoutput.t32 4.06363
R22091 CSoutput.n117 CSoutput.t95 4.06363
R22092 CSoutput.n119 CSoutput.t64 4.06363
R22093 CSoutput.n119 CSoutput.t63 4.06363
R22094 CSoutput.n121 CSoutput.t54 4.06363
R22095 CSoutput.n121 CSoutput.t31 4.06363
R22096 CSoutput.n123 CSoutput.t17 4.06363
R22097 CSoutput.n123 CSoutput.t55 4.06363
R22098 CSoutput.n94 CSoutput.t76 4.06363
R22099 CSoutput.n94 CSoutput.t74 4.06363
R22100 CSoutput.n95 CSoutput.t59 4.06363
R22101 CSoutput.n95 CSoutput.t8 4.06363
R22102 CSoutput.n97 CSoutput.t3 4.06363
R22103 CSoutput.n97 CSoutput.t70 4.06363
R22104 CSoutput.n99 CSoutput.t58 4.06363
R22105 CSoutput.n99 CSoutput.t38 4.06363
R22106 CSoutput.n101 CSoutput.t23 4.06363
R22107 CSoutput.n101 CSoutput.t85 4.06363
R22108 CSoutput.n103 CSoutput.t57 4.06363
R22109 CSoutput.n103 CSoutput.t56 4.06363
R22110 CSoutput.n105 CSoutput.t47 4.06363
R22111 CSoutput.n105 CSoutput.t19 4.06363
R22112 CSoutput.n107 CSoutput.t6 4.06363
R22113 CSoutput.n107 CSoutput.t48 4.06363
R22114 CSoutput.n79 CSoutput.t82 4.06363
R22115 CSoutput.n79 CSoutput.t2 4.06363
R22116 CSoutput.n80 CSoutput.t65 4.06363
R22117 CSoutput.n80 CSoutput.t42 4.06363
R22118 CSoutput.n82 CSoutput.t72 4.06363
R22119 CSoutput.n82 CSoutput.t22 4.06363
R22120 CSoutput.n84 CSoutput.t89 4.06363
R22121 CSoutput.n84 CSoutput.t36 4.06363
R22122 CSoutput.n86 CSoutput.t7 4.06363
R22123 CSoutput.n86 CSoutput.t50 4.06363
R22124 CSoutput.n88 CSoutput.t11 4.06363
R22125 CSoutput.n88 CSoutput.t30 4.06363
R22126 CSoutput.n90 CSoutput.t94 4.06363
R22127 CSoutput.n90 CSoutput.t44 4.06363
R22128 CSoutput.n92 CSoutput.t14 4.06363
R22129 CSoutput.n92 CSoutput.t78 4.06363
R22130 CSoutput.n44 CSoutput.n43 3.79402
R22131 CSoutput.n49 CSoutput.n48 3.79402
R22132 CSoutput.n371 CSoutput.n355 3.72967
R22133 CSoutput.n419 CSoutput.n403 3.72967
R22134 CSoutput.n421 CSoutput.n420 3.57343
R22135 CSoutput.n420 CSoutput.n372 3.3798
R22136 CSoutput.n369 CSoutput.t112 2.82907
R22137 CSoutput.n369 CSoutput.t119 2.82907
R22138 CSoutput.n367 CSoutput.t105 2.82907
R22139 CSoutput.n367 CSoutput.t185 2.82907
R22140 CSoutput.n365 CSoutput.t154 2.82907
R22141 CSoutput.n365 CSoutput.t97 2.82907
R22142 CSoutput.n363 CSoutput.t188 2.82907
R22143 CSoutput.n363 CSoutput.t174 2.82907
R22144 CSoutput.n361 CSoutput.t135 2.82907
R22145 CSoutput.n361 CSoutput.t144 2.82907
R22146 CSoutput.n359 CSoutput.t96 2.82907
R22147 CSoutput.n359 CSoutput.t181 2.82907
R22148 CSoutput.n357 CSoutput.t175 2.82907
R22149 CSoutput.n357 CSoutput.t121 2.82907
R22150 CSoutput.n356 CSoutput.t107 2.82907
R22151 CSoutput.n356 CSoutput.t187 2.82907
R22152 CSoutput.n353 CSoutput.t120 2.82907
R22153 CSoutput.n353 CSoutput.t191 2.82907
R22154 CSoutput.n351 CSoutput.t103 2.82907
R22155 CSoutput.n351 CSoutput.t186 2.82907
R22156 CSoutput.n349 CSoutput.t114 2.82907
R22157 CSoutput.n349 CSoutput.t130 2.82907
R22158 CSoutput.n347 CSoutput.t128 2.82907
R22159 CSoutput.n347 CSoutput.t106 2.82907
R22160 CSoutput.n345 CSoutput.t141 2.82907
R22161 CSoutput.n345 CSoutput.t115 2.82907
R22162 CSoutput.n343 CSoutput.t116 2.82907
R22163 CSoutput.n343 CSoutput.t129 2.82907
R22164 CSoutput.n341 CSoutput.t127 2.82907
R22165 CSoutput.n341 CSoutput.t139 2.82907
R22166 CSoutput.n340 CSoutput.t140 2.82907
R22167 CSoutput.n340 CSoutput.t117 2.82907
R22168 CSoutput.n338 CSoutput.t108 2.82907
R22169 CSoutput.n338 CSoutput.t123 2.82907
R22170 CSoutput.n336 CSoutput.t145 2.82907
R22171 CSoutput.n336 CSoutput.t173 2.82907
R22172 CSoutput.n334 CSoutput.t163 2.82907
R22173 CSoutput.n334 CSoutput.t132 2.82907
R22174 CSoutput.n332 CSoutput.t101 2.82907
R22175 CSoutput.n332 CSoutput.t149 2.82907
R22176 CSoutput.n330 CSoutput.t131 2.82907
R22177 CSoutput.n330 CSoutput.t142 2.82907
R22178 CSoutput.n328 CSoutput.t143 2.82907
R22179 CSoutput.n328 CSoutput.t180 2.82907
R22180 CSoutput.n326 CSoutput.t159 2.82907
R22181 CSoutput.n326 CSoutput.t98 2.82907
R22182 CSoutput.n325 CSoutput.t177 2.82907
R22183 CSoutput.n325 CSoutput.t109 2.82907
R22184 CSoutput.n404 CSoutput.t169 2.82907
R22185 CSoutput.n404 CSoutput.t184 2.82907
R22186 CSoutput.n405 CSoutput.t189 2.82907
R22187 CSoutput.n405 CSoutput.t158 2.82907
R22188 CSoutput.n407 CSoutput.t162 2.82907
R22189 CSoutput.n407 CSoutput.t178 2.82907
R22190 CSoutput.n409 CSoutput.t110 2.82907
R22191 CSoutput.n409 CSoutput.t152 2.82907
R22192 CSoutput.n411 CSoutput.t157 2.82907
R22193 CSoutput.n411 CSoutput.t170 2.82907
R22194 CSoutput.n413 CSoutput.t179 2.82907
R22195 CSoutput.n413 CSoutput.t161 2.82907
R22196 CSoutput.n415 CSoutput.t166 2.82907
R22197 CSoutput.n415 CSoutput.t183 2.82907
R22198 CSoutput.n417 CSoutput.t111 2.82907
R22199 CSoutput.n417 CSoutput.t122 2.82907
R22200 CSoutput.n388 CSoutput.t137 2.82907
R22201 CSoutput.n388 CSoutput.t155 2.82907
R22202 CSoutput.n389 CSoutput.t156 2.82907
R22203 CSoutput.n389 CSoutput.t146 2.82907
R22204 CSoutput.n391 CSoutput.t147 2.82907
R22205 CSoutput.n391 CSoutput.t138 2.82907
R22206 CSoutput.n393 CSoutput.t133 2.82907
R22207 CSoutput.n393 CSoutput.t125 2.82907
R22208 CSoutput.n395 CSoutput.t126 2.82907
R22209 CSoutput.n395 CSoutput.t148 2.82907
R22210 CSoutput.n397 CSoutput.t150 2.82907
R22211 CSoutput.n397 CSoutput.t99 2.82907
R22212 CSoutput.n399 CSoutput.t100 2.82907
R22213 CSoutput.n399 CSoutput.t118 2.82907
R22214 CSoutput.n401 CSoutput.t124 2.82907
R22215 CSoutput.n401 CSoutput.t113 2.82907
R22216 CSoutput.n373 CSoutput.t151 2.82907
R22217 CSoutput.n373 CSoutput.t102 2.82907
R22218 CSoutput.n374 CSoutput.t134 2.82907
R22219 CSoutput.n374 CSoutput.t182 2.82907
R22220 CSoutput.n376 CSoutput.t104 2.82907
R22221 CSoutput.n376 CSoutput.t165 2.82907
R22222 CSoutput.n378 CSoutput.t164 2.82907
R22223 CSoutput.n378 CSoutput.t153 2.82907
R22224 CSoutput.n380 CSoutput.t168 2.82907
R22225 CSoutput.n380 CSoutput.t136 2.82907
R22226 CSoutput.n382 CSoutput.t160 2.82907
R22227 CSoutput.n382 CSoutput.t176 2.82907
R22228 CSoutput.n384 CSoutput.t190 2.82907
R22229 CSoutput.n384 CSoutput.t167 2.82907
R22230 CSoutput.n386 CSoutput.t172 2.82907
R22231 CSoutput.n386 CSoutput.t171 2.82907
R22232 CSoutput.n75 CSoutput.n1 2.45513
R22233 CSoutput.n324 CSoutput.n126 2.36742
R22234 CSoutput.n217 CSoutput.n215 2.251
R22235 CSoutput.n217 CSoutput.n214 2.251
R22236 CSoutput.n217 CSoutput.n213 2.251
R22237 CSoutput.n217 CSoutput.n212 2.251
R22238 CSoutput.n186 CSoutput.n185 2.251
R22239 CSoutput.n186 CSoutput.n184 2.251
R22240 CSoutput.n186 CSoutput.n183 2.251
R22241 CSoutput.n186 CSoutput.n182 2.251
R22242 CSoutput.n259 CSoutput.n258 2.251
R22243 CSoutput.n224 CSoutput.n222 2.251
R22244 CSoutput.n224 CSoutput.n221 2.251
R22245 CSoutput.n224 CSoutput.n220 2.251
R22246 CSoutput.n242 CSoutput.n224 2.251
R22247 CSoutput.n230 CSoutput.n229 2.251
R22248 CSoutput.n230 CSoutput.n228 2.251
R22249 CSoutput.n230 CSoutput.n227 2.251
R22250 CSoutput.n230 CSoutput.n226 2.251
R22251 CSoutput.n256 CSoutput.n196 2.251
R22252 CSoutput.n251 CSoutput.n249 2.251
R22253 CSoutput.n251 CSoutput.n248 2.251
R22254 CSoutput.n251 CSoutput.n247 2.251
R22255 CSoutput.n251 CSoutput.n246 2.251
R22256 CSoutput.n152 CSoutput.n151 2.251
R22257 CSoutput.n152 CSoutput.n150 2.251
R22258 CSoutput.n152 CSoutput.n149 2.251
R22259 CSoutput.n152 CSoutput.n148 2.251
R22260 CSoutput.n269 CSoutput.n268 2.251
R22261 CSoutput.n186 CSoutput.n166 2.2505
R22262 CSoutput.n181 CSoutput.n166 2.2505
R22263 CSoutput.n179 CSoutput.n166 2.2505
R22264 CSoutput.n178 CSoutput.n166 2.2505
R22265 CSoutput.n263 CSoutput.n166 2.2505
R22266 CSoutput.n261 CSoutput.n166 2.2505
R22267 CSoutput.n259 CSoutput.n166 2.2505
R22268 CSoutput.n189 CSoutput.n166 2.2505
R22269 CSoutput.n188 CSoutput.n166 2.2505
R22270 CSoutput.n192 CSoutput.n166 2.2505
R22271 CSoutput.n191 CSoutput.n166 2.2505
R22272 CSoutput.n174 CSoutput.n166 2.2505
R22273 CSoutput.n266 CSoutput.n166 2.2505
R22274 CSoutput.n266 CSoutput.n265 2.2505
R22275 CSoutput.n230 CSoutput.n201 2.2505
R22276 CSoutput.n211 CSoutput.n201 2.2505
R22277 CSoutput.n232 CSoutput.n201 2.2505
R22278 CSoutput.n210 CSoutput.n201 2.2505
R22279 CSoutput.n234 CSoutput.n201 2.2505
R22280 CSoutput.n201 CSoutput.n195 2.2505
R22281 CSoutput.n256 CSoutput.n201 2.2505
R22282 CSoutput.n254 CSoutput.n201 2.2505
R22283 CSoutput.n236 CSoutput.n201 2.2505
R22284 CSoutput.n208 CSoutput.n201 2.2505
R22285 CSoutput.n238 CSoutput.n201 2.2505
R22286 CSoutput.n207 CSoutput.n201 2.2505
R22287 CSoutput.n252 CSoutput.n201 2.2505
R22288 CSoutput.n252 CSoutput.n205 2.2505
R22289 CSoutput.n152 CSoutput.n132 2.2505
R22290 CSoutput.n147 CSoutput.n132 2.2505
R22291 CSoutput.n145 CSoutput.n132 2.2505
R22292 CSoutput.n144 CSoutput.n132 2.2505
R22293 CSoutput.n273 CSoutput.n132 2.2505
R22294 CSoutput.n271 CSoutput.n132 2.2505
R22295 CSoutput.n269 CSoutput.n132 2.2505
R22296 CSoutput.n155 CSoutput.n132 2.2505
R22297 CSoutput.n154 CSoutput.n132 2.2505
R22298 CSoutput.n158 CSoutput.n132 2.2505
R22299 CSoutput.n157 CSoutput.n132 2.2505
R22300 CSoutput.n140 CSoutput.n132 2.2505
R22301 CSoutput.n276 CSoutput.n132 2.2505
R22302 CSoutput.n276 CSoutput.n275 2.2505
R22303 CSoutput.n194 CSoutput.n187 2.25024
R22304 CSoutput.n194 CSoutput.n180 2.25024
R22305 CSoutput.n262 CSoutput.n194 2.25024
R22306 CSoutput.n194 CSoutput.n190 2.25024
R22307 CSoutput.n194 CSoutput.n193 2.25024
R22308 CSoutput.n194 CSoutput.n161 2.25024
R22309 CSoutput.n244 CSoutput.n241 2.25024
R22310 CSoutput.n244 CSoutput.n240 2.25024
R22311 CSoutput.n244 CSoutput.n239 2.25024
R22312 CSoutput.n244 CSoutput.n206 2.25024
R22313 CSoutput.n244 CSoutput.n243 2.25024
R22314 CSoutput.n245 CSoutput.n244 2.25024
R22315 CSoutput.n160 CSoutput.n153 2.25024
R22316 CSoutput.n160 CSoutput.n146 2.25024
R22317 CSoutput.n272 CSoutput.n160 2.25024
R22318 CSoutput.n160 CSoutput.n156 2.25024
R22319 CSoutput.n160 CSoutput.n159 2.25024
R22320 CSoutput.n160 CSoutput.n127 2.25024
R22321 CSoutput.n261 CSoutput.n171 1.50111
R22322 CSoutput.n209 CSoutput.n195 1.50111
R22323 CSoutput.n271 CSoutput.n137 1.50111
R22324 CSoutput.n217 CSoutput.n216 1.501
R22325 CSoutput.n224 CSoutput.n223 1.501
R22326 CSoutput.n251 CSoutput.n250 1.501
R22327 CSoutput.n265 CSoutput.n176 1.12536
R22328 CSoutput.n265 CSoutput.n177 1.12536
R22329 CSoutput.n265 CSoutput.n264 1.12536
R22330 CSoutput.n225 CSoutput.n205 1.12536
R22331 CSoutput.n231 CSoutput.n205 1.12536
R22332 CSoutput.n233 CSoutput.n205 1.12536
R22333 CSoutput.n275 CSoutput.n142 1.12536
R22334 CSoutput.n275 CSoutput.n143 1.12536
R22335 CSoutput.n275 CSoutput.n274 1.12536
R22336 CSoutput.n265 CSoutput.n172 1.12536
R22337 CSoutput.n265 CSoutput.n173 1.12536
R22338 CSoutput.n265 CSoutput.n175 1.12536
R22339 CSoutput.n255 CSoutput.n205 1.12536
R22340 CSoutput.n235 CSoutput.n205 1.12536
R22341 CSoutput.n237 CSoutput.n205 1.12536
R22342 CSoutput.n275 CSoutput.n138 1.12536
R22343 CSoutput.n275 CSoutput.n139 1.12536
R22344 CSoutput.n275 CSoutput.n141 1.12536
R22345 CSoutput.n31 CSoutput.n30 0.669944
R22346 CSoutput.n62 CSoutput.n61 0.669944
R22347 CSoutput.n360 CSoutput.n358 0.573776
R22348 CSoutput.n362 CSoutput.n360 0.573776
R22349 CSoutput.n364 CSoutput.n362 0.573776
R22350 CSoutput.n366 CSoutput.n364 0.573776
R22351 CSoutput.n368 CSoutput.n366 0.573776
R22352 CSoutput.n370 CSoutput.n368 0.573776
R22353 CSoutput.n344 CSoutput.n342 0.573776
R22354 CSoutput.n346 CSoutput.n344 0.573776
R22355 CSoutput.n348 CSoutput.n346 0.573776
R22356 CSoutput.n350 CSoutput.n348 0.573776
R22357 CSoutput.n352 CSoutput.n350 0.573776
R22358 CSoutput.n354 CSoutput.n352 0.573776
R22359 CSoutput.n329 CSoutput.n327 0.573776
R22360 CSoutput.n331 CSoutput.n329 0.573776
R22361 CSoutput.n333 CSoutput.n331 0.573776
R22362 CSoutput.n335 CSoutput.n333 0.573776
R22363 CSoutput.n337 CSoutput.n335 0.573776
R22364 CSoutput.n339 CSoutput.n337 0.573776
R22365 CSoutput.n418 CSoutput.n416 0.573776
R22366 CSoutput.n416 CSoutput.n414 0.573776
R22367 CSoutput.n414 CSoutput.n412 0.573776
R22368 CSoutput.n412 CSoutput.n410 0.573776
R22369 CSoutput.n410 CSoutput.n408 0.573776
R22370 CSoutput.n408 CSoutput.n406 0.573776
R22371 CSoutput.n402 CSoutput.n400 0.573776
R22372 CSoutput.n400 CSoutput.n398 0.573776
R22373 CSoutput.n398 CSoutput.n396 0.573776
R22374 CSoutput.n396 CSoutput.n394 0.573776
R22375 CSoutput.n394 CSoutput.n392 0.573776
R22376 CSoutput.n392 CSoutput.n390 0.573776
R22377 CSoutput.n387 CSoutput.n385 0.573776
R22378 CSoutput.n385 CSoutput.n383 0.573776
R22379 CSoutput.n383 CSoutput.n381 0.573776
R22380 CSoutput.n381 CSoutput.n379 0.573776
R22381 CSoutput.n379 CSoutput.n377 0.573776
R22382 CSoutput.n377 CSoutput.n375 0.573776
R22383 CSoutput.n421 CSoutput.n276 0.53442
R22384 CSoutput.n312 CSoutput.n310 0.358259
R22385 CSoutput.n314 CSoutput.n312 0.358259
R22386 CSoutput.n316 CSoutput.n314 0.358259
R22387 CSoutput.n318 CSoutput.n316 0.358259
R22388 CSoutput.n320 CSoutput.n318 0.358259
R22389 CSoutput.n322 CSoutput.n320 0.358259
R22390 CSoutput.n296 CSoutput.n294 0.358259
R22391 CSoutput.n298 CSoutput.n296 0.358259
R22392 CSoutput.n300 CSoutput.n298 0.358259
R22393 CSoutput.n302 CSoutput.n300 0.358259
R22394 CSoutput.n304 CSoutput.n302 0.358259
R22395 CSoutput.n306 CSoutput.n304 0.358259
R22396 CSoutput.n281 CSoutput.n279 0.358259
R22397 CSoutput.n283 CSoutput.n281 0.358259
R22398 CSoutput.n285 CSoutput.n283 0.358259
R22399 CSoutput.n287 CSoutput.n285 0.358259
R22400 CSoutput.n289 CSoutput.n287 0.358259
R22401 CSoutput.n291 CSoutput.n289 0.358259
R22402 CSoutput.n124 CSoutput.n122 0.358259
R22403 CSoutput.n122 CSoutput.n120 0.358259
R22404 CSoutput.n120 CSoutput.n118 0.358259
R22405 CSoutput.n118 CSoutput.n116 0.358259
R22406 CSoutput.n116 CSoutput.n114 0.358259
R22407 CSoutput.n114 CSoutput.n112 0.358259
R22408 CSoutput.n108 CSoutput.n106 0.358259
R22409 CSoutput.n106 CSoutput.n104 0.358259
R22410 CSoutput.n104 CSoutput.n102 0.358259
R22411 CSoutput.n102 CSoutput.n100 0.358259
R22412 CSoutput.n100 CSoutput.n98 0.358259
R22413 CSoutput.n98 CSoutput.n96 0.358259
R22414 CSoutput.n93 CSoutput.n91 0.358259
R22415 CSoutput.n91 CSoutput.n89 0.358259
R22416 CSoutput.n89 CSoutput.n87 0.358259
R22417 CSoutput.n87 CSoutput.n85 0.358259
R22418 CSoutput.n85 CSoutput.n83 0.358259
R22419 CSoutput.n83 CSoutput.n81 0.358259
R22420 CSoutput.n21 CSoutput.n20 0.169105
R22421 CSoutput.n21 CSoutput.n16 0.169105
R22422 CSoutput.n26 CSoutput.n16 0.169105
R22423 CSoutput.n27 CSoutput.n26 0.169105
R22424 CSoutput.n27 CSoutput.n14 0.169105
R22425 CSoutput.n32 CSoutput.n14 0.169105
R22426 CSoutput.n33 CSoutput.n32 0.169105
R22427 CSoutput.n34 CSoutput.n33 0.169105
R22428 CSoutput.n34 CSoutput.n12 0.169105
R22429 CSoutput.n39 CSoutput.n12 0.169105
R22430 CSoutput.n40 CSoutput.n39 0.169105
R22431 CSoutput.n40 CSoutput.n10 0.169105
R22432 CSoutput.n45 CSoutput.n10 0.169105
R22433 CSoutput.n46 CSoutput.n45 0.169105
R22434 CSoutput.n47 CSoutput.n46 0.169105
R22435 CSoutput.n47 CSoutput.n8 0.169105
R22436 CSoutput.n52 CSoutput.n8 0.169105
R22437 CSoutput.n53 CSoutput.n52 0.169105
R22438 CSoutput.n53 CSoutput.n6 0.169105
R22439 CSoutput.n58 CSoutput.n6 0.169105
R22440 CSoutput.n59 CSoutput.n58 0.169105
R22441 CSoutput.n60 CSoutput.n59 0.169105
R22442 CSoutput.n60 CSoutput.n4 0.169105
R22443 CSoutput.n66 CSoutput.n4 0.169105
R22444 CSoutput.n67 CSoutput.n66 0.169105
R22445 CSoutput.n68 CSoutput.n67 0.169105
R22446 CSoutput.n68 CSoutput.n2 0.169105
R22447 CSoutput.n73 CSoutput.n2 0.169105
R22448 CSoutput.n74 CSoutput.n73 0.169105
R22449 CSoutput.n74 CSoutput.n0 0.169105
R22450 CSoutput.n78 CSoutput.n0 0.169105
R22451 CSoutput.n219 CSoutput.n218 0.0910737
R22452 CSoutput.n270 CSoutput.n267 0.0723685
R22453 CSoutput.n224 CSoutput.n219 0.0522944
R22454 CSoutput.n267 CSoutput.n266 0.0499135
R22455 CSoutput.n218 CSoutput.n217 0.0499135
R22456 CSoutput.n252 CSoutput.n251 0.0464294
R22457 CSoutput.n260 CSoutput.n257 0.0391444
R22458 CSoutput.n219 CSoutput.t212 0.023435
R22459 CSoutput.n267 CSoutput.t204 0.02262
R22460 CSoutput.n218 CSoutput.t193 0.02262
R22461 CSoutput CSoutput.n421 0.0052
R22462 CSoutput.n189 CSoutput.n172 0.00365111
R22463 CSoutput.n192 CSoutput.n173 0.00365111
R22464 CSoutput.n175 CSoutput.n174 0.00365111
R22465 CSoutput.n217 CSoutput.n176 0.00365111
R22466 CSoutput.n181 CSoutput.n177 0.00365111
R22467 CSoutput.n264 CSoutput.n178 0.00365111
R22468 CSoutput.n255 CSoutput.n254 0.00365111
R22469 CSoutput.n235 CSoutput.n208 0.00365111
R22470 CSoutput.n237 CSoutput.n207 0.00365111
R22471 CSoutput.n225 CSoutput.n224 0.00365111
R22472 CSoutput.n231 CSoutput.n211 0.00365111
R22473 CSoutput.n233 CSoutput.n210 0.00365111
R22474 CSoutput.n155 CSoutput.n138 0.00365111
R22475 CSoutput.n158 CSoutput.n139 0.00365111
R22476 CSoutput.n141 CSoutput.n140 0.00365111
R22477 CSoutput.n251 CSoutput.n142 0.00365111
R22478 CSoutput.n147 CSoutput.n143 0.00365111
R22479 CSoutput.n274 CSoutput.n144 0.00365111
R22480 CSoutput.n186 CSoutput.n176 0.00340054
R22481 CSoutput.n179 CSoutput.n177 0.00340054
R22482 CSoutput.n264 CSoutput.n263 0.00340054
R22483 CSoutput.n259 CSoutput.n172 0.00340054
R22484 CSoutput.n188 CSoutput.n173 0.00340054
R22485 CSoutput.n191 CSoutput.n175 0.00340054
R22486 CSoutput.n230 CSoutput.n225 0.00340054
R22487 CSoutput.n232 CSoutput.n231 0.00340054
R22488 CSoutput.n234 CSoutput.n233 0.00340054
R22489 CSoutput.n256 CSoutput.n255 0.00340054
R22490 CSoutput.n236 CSoutput.n235 0.00340054
R22491 CSoutput.n238 CSoutput.n237 0.00340054
R22492 CSoutput.n152 CSoutput.n142 0.00340054
R22493 CSoutput.n145 CSoutput.n143 0.00340054
R22494 CSoutput.n274 CSoutput.n273 0.00340054
R22495 CSoutput.n269 CSoutput.n138 0.00340054
R22496 CSoutput.n154 CSoutput.n139 0.00340054
R22497 CSoutput.n157 CSoutput.n141 0.00340054
R22498 CSoutput.n187 CSoutput.n181 0.00252698
R22499 CSoutput.n180 CSoutput.n178 0.00252698
R22500 CSoutput.n262 CSoutput.n261 0.00252698
R22501 CSoutput.n190 CSoutput.n188 0.00252698
R22502 CSoutput.n193 CSoutput.n191 0.00252698
R22503 CSoutput.n266 CSoutput.n161 0.00252698
R22504 CSoutput.n187 CSoutput.n186 0.00252698
R22505 CSoutput.n180 CSoutput.n179 0.00252698
R22506 CSoutput.n263 CSoutput.n262 0.00252698
R22507 CSoutput.n190 CSoutput.n189 0.00252698
R22508 CSoutput.n193 CSoutput.n192 0.00252698
R22509 CSoutput.n174 CSoutput.n161 0.00252698
R22510 CSoutput.n241 CSoutput.n211 0.00252698
R22511 CSoutput.n240 CSoutput.n210 0.00252698
R22512 CSoutput.n239 CSoutput.n195 0.00252698
R22513 CSoutput.n236 CSoutput.n206 0.00252698
R22514 CSoutput.n243 CSoutput.n238 0.00252698
R22515 CSoutput.n252 CSoutput.n245 0.00252698
R22516 CSoutput.n241 CSoutput.n230 0.00252698
R22517 CSoutput.n240 CSoutput.n232 0.00252698
R22518 CSoutput.n239 CSoutput.n234 0.00252698
R22519 CSoutput.n254 CSoutput.n206 0.00252698
R22520 CSoutput.n243 CSoutput.n208 0.00252698
R22521 CSoutput.n245 CSoutput.n207 0.00252698
R22522 CSoutput.n153 CSoutput.n147 0.00252698
R22523 CSoutput.n146 CSoutput.n144 0.00252698
R22524 CSoutput.n272 CSoutput.n271 0.00252698
R22525 CSoutput.n156 CSoutput.n154 0.00252698
R22526 CSoutput.n159 CSoutput.n157 0.00252698
R22527 CSoutput.n276 CSoutput.n127 0.00252698
R22528 CSoutput.n153 CSoutput.n152 0.00252698
R22529 CSoutput.n146 CSoutput.n145 0.00252698
R22530 CSoutput.n273 CSoutput.n272 0.00252698
R22531 CSoutput.n156 CSoutput.n155 0.00252698
R22532 CSoutput.n159 CSoutput.n158 0.00252698
R22533 CSoutput.n140 CSoutput.n127 0.00252698
R22534 CSoutput.n261 CSoutput.n260 0.0020275
R22535 CSoutput.n260 CSoutput.n259 0.0020275
R22536 CSoutput.n257 CSoutput.n195 0.0020275
R22537 CSoutput.n257 CSoutput.n256 0.0020275
R22538 CSoutput.n271 CSoutput.n270 0.0020275
R22539 CSoutput.n270 CSoutput.n269 0.0020275
R22540 CSoutput.n171 CSoutput.n170 0.00166668
R22541 CSoutput.n253 CSoutput.n209 0.00166668
R22542 CSoutput.n137 CSoutput.n136 0.00166668
R22543 CSoutput.n275 CSoutput.n137 0.00133328
R22544 CSoutput.n209 CSoutput.n205 0.00133328
R22545 CSoutput.n265 CSoutput.n171 0.00133328
R22546 CSoutput.n268 CSoutput.n160 0.001
R22547 CSoutput.n246 CSoutput.n160 0.001
R22548 CSoutput.n148 CSoutput.n128 0.001
R22549 CSoutput.n247 CSoutput.n128 0.001
R22550 CSoutput.n149 CSoutput.n129 0.001
R22551 CSoutput.n248 CSoutput.n129 0.001
R22552 CSoutput.n150 CSoutput.n130 0.001
R22553 CSoutput.n249 CSoutput.n130 0.001
R22554 CSoutput.n151 CSoutput.n131 0.001
R22555 CSoutput.n250 CSoutput.n131 0.001
R22556 CSoutput.n244 CSoutput.n196 0.001
R22557 CSoutput.n244 CSoutput.n242 0.001
R22558 CSoutput.n226 CSoutput.n197 0.001
R22559 CSoutput.n220 CSoutput.n197 0.001
R22560 CSoutput.n227 CSoutput.n198 0.001
R22561 CSoutput.n221 CSoutput.n198 0.001
R22562 CSoutput.n228 CSoutput.n199 0.001
R22563 CSoutput.n222 CSoutput.n199 0.001
R22564 CSoutput.n229 CSoutput.n200 0.001
R22565 CSoutput.n223 CSoutput.n200 0.001
R22566 CSoutput.n258 CSoutput.n194 0.001
R22567 CSoutput.n212 CSoutput.n194 0.001
R22568 CSoutput.n182 CSoutput.n162 0.001
R22569 CSoutput.n213 CSoutput.n162 0.001
R22570 CSoutput.n183 CSoutput.n163 0.001
R22571 CSoutput.n214 CSoutput.n163 0.001
R22572 CSoutput.n184 CSoutput.n164 0.001
R22573 CSoutput.n215 CSoutput.n164 0.001
R22574 CSoutput.n185 CSoutput.n165 0.001
R22575 CSoutput.n216 CSoutput.n165 0.001
R22576 CSoutput.n216 CSoutput.n166 0.001
R22577 CSoutput.n215 CSoutput.n167 0.001
R22578 CSoutput.n214 CSoutput.n168 0.001
R22579 CSoutput.n213 CSoutput.t209 0.001
R22580 CSoutput.n212 CSoutput.n169 0.001
R22581 CSoutput.n185 CSoutput.n167 0.001
R22582 CSoutput.n184 CSoutput.n168 0.001
R22583 CSoutput.n183 CSoutput.t209 0.001
R22584 CSoutput.n182 CSoutput.n169 0.001
R22585 CSoutput.n258 CSoutput.n170 0.001
R22586 CSoutput.n223 CSoutput.n201 0.001
R22587 CSoutput.n222 CSoutput.n202 0.001
R22588 CSoutput.n221 CSoutput.n203 0.001
R22589 CSoutput.n220 CSoutput.t202 0.001
R22590 CSoutput.n242 CSoutput.n204 0.001
R22591 CSoutput.n229 CSoutput.n202 0.001
R22592 CSoutput.n228 CSoutput.n203 0.001
R22593 CSoutput.n227 CSoutput.t202 0.001
R22594 CSoutput.n226 CSoutput.n204 0.001
R22595 CSoutput.n253 CSoutput.n196 0.001
R22596 CSoutput.n250 CSoutput.n132 0.001
R22597 CSoutput.n249 CSoutput.n133 0.001
R22598 CSoutput.n248 CSoutput.n134 0.001
R22599 CSoutput.n247 CSoutput.t192 0.001
R22600 CSoutput.n246 CSoutput.n135 0.001
R22601 CSoutput.n151 CSoutput.n133 0.001
R22602 CSoutput.n150 CSoutput.n134 0.001
R22603 CSoutput.n149 CSoutput.t192 0.001
R22604 CSoutput.n148 CSoutput.n135 0.001
R22605 CSoutput.n268 CSoutput.n136 0.001
R22606 a_n2848_n452.n10 a_n2848_n452.t74 539.01
R22607 a_n2848_n452.n93 a_n2848_n452.t57 512.366
R22608 a_n2848_n452.n92 a_n2848_n452.t61 512.366
R22609 a_n2848_n452.n66 a_n2848_n452.t51 512.366
R22610 a_n2848_n452.n91 a_n2848_n452.t66 512.366
R22611 a_n2848_n452.n6 a_n2848_n452.t25 533.058
R22612 a_n2848_n452.n97 a_n2848_n452.t23 512.366
R22613 a_n2848_n452.n96 a_n2848_n452.t11 512.366
R22614 a_n2848_n452.n65 a_n2848_n452.t3 512.366
R22615 a_n2848_n452.n94 a_n2848_n452.t5 512.366
R22616 a_n2848_n452.n24 a_n2848_n452.t9 539.01
R22617 a_n2848_n452.n74 a_n2848_n452.t17 512.366
R22618 a_n2848_n452.n75 a_n2848_n452.t13 512.366
R22619 a_n2848_n452.n69 a_n2848_n452.t15 512.366
R22620 a_n2848_n452.n76 a_n2848_n452.t7 512.366
R22621 a_n2848_n452.n28 a_n2848_n452.t69 539.01
R22622 a_n2848_n452.n71 a_n2848_n452.t70 512.366
R22623 a_n2848_n452.n72 a_n2848_n452.t49 512.366
R22624 a_n2848_n452.n70 a_n2848_n452.t56 512.366
R22625 a_n2848_n452.n73 a_n2848_n452.t64 512.366
R22626 a_n2848_n452.n88 a_n2848_n452.t63 512.366
R22627 a_n2848_n452.n78 a_n2848_n452.t54 512.366
R22628 a_n2848_n452.n89 a_n2848_n452.t48 512.366
R22629 a_n2848_n452.n86 a_n2848_n452.t71 512.366
R22630 a_n2848_n452.n79 a_n2848_n452.t60 512.366
R22631 a_n2848_n452.n87 a_n2848_n452.t59 512.366
R22632 a_n2848_n452.n84 a_n2848_n452.t67 512.366
R22633 a_n2848_n452.n80 a_n2848_n452.t52 512.366
R22634 a_n2848_n452.n85 a_n2848_n452.t53 512.366
R22635 a_n2848_n452.n82 a_n2848_n452.t55 512.366
R22636 a_n2848_n452.n81 a_n2848_n452.t65 512.366
R22637 a_n2848_n452.n83 a_n2848_n452.t75 512.366
R22638 a_n2848_n452.n51 a_n2848_n452.n8 70.3058
R22639 a_n2848_n452.n48 a_n2848_n452.n11 70.3058
R22640 a_n2848_n452.n21 a_n2848_n452.n38 70.3058
R22641 a_n2848_n452.n25 a_n2848_n452.n35 70.3058
R22642 a_n2848_n452.n34 a_n2848_n452.n26 70.1674
R22643 a_n2848_n452.n34 a_n2848_n452.n70 20.9683
R22644 a_n2848_n452.n26 a_n2848_n452.n33 75.0448
R22645 a_n2848_n452.n72 a_n2848_n452.n33 11.2134
R22646 a_n2848_n452.n27 a_n2848_n452.n28 44.8194
R22647 a_n2848_n452.n37 a_n2848_n452.n22 70.1674
R22648 a_n2848_n452.n37 a_n2848_n452.n69 20.9683
R22649 a_n2848_n452.n22 a_n2848_n452.n36 75.0448
R22650 a_n2848_n452.n75 a_n2848_n452.n36 11.2134
R22651 a_n2848_n452.n23 a_n2848_n452.n24 44.8194
R22652 a_n2848_n452.n12 a_n2848_n452.n46 70.1674
R22653 a_n2848_n452.n14 a_n2848_n452.n44 70.1674
R22654 a_n2848_n452.n16 a_n2848_n452.n42 70.1674
R22655 a_n2848_n452.n19 a_n2848_n452.n40 70.1674
R22656 a_n2848_n452.n83 a_n2848_n452.n40 20.9683
R22657 a_n2848_n452.n39 a_n2848_n452.n20 75.0448
R22658 a_n2848_n452.n39 a_n2848_n452.n81 11.2134
R22659 a_n2848_n452.n20 a_n2848_n452.n82 161.3
R22660 a_n2848_n452.n85 a_n2848_n452.n42 20.9683
R22661 a_n2848_n452.n41 a_n2848_n452.n17 75.0448
R22662 a_n2848_n452.n41 a_n2848_n452.n80 11.2134
R22663 a_n2848_n452.n17 a_n2848_n452.n84 161.3
R22664 a_n2848_n452.n87 a_n2848_n452.n44 20.9683
R22665 a_n2848_n452.n43 a_n2848_n452.n15 75.0448
R22666 a_n2848_n452.n43 a_n2848_n452.n79 11.2134
R22667 a_n2848_n452.n15 a_n2848_n452.n86 161.3
R22668 a_n2848_n452.n89 a_n2848_n452.n46 20.9683
R22669 a_n2848_n452.n45 a_n2848_n452.n13 75.0448
R22670 a_n2848_n452.n45 a_n2848_n452.n78 11.2134
R22671 a_n2848_n452.n13 a_n2848_n452.n88 161.3
R22672 a_n2848_n452.n11 a_n2848_n452.n47 70.1674
R22673 a_n2848_n452.n47 a_n2848_n452.n65 20.9683
R22674 a_n2848_n452.n95 a_n2848_n452.n5 161.3
R22675 a_n2848_n452.n9 a_n2848_n452.n50 70.1674
R22676 a_n2848_n452.n50 a_n2848_n452.n66 20.9683
R22677 a_n2848_n452.n49 a_n2848_n452.n9 75.0448
R22678 a_n2848_n452.n92 a_n2848_n452.n49 11.2134
R22679 a_n2848_n452.n7 a_n2848_n452.n10 44.8194
R22680 a_n2848_n452.n96 a_n2848_n452.n52 20.9683
R22681 a_n2848_n452.n52 a_n2848_n452.n5 70.1674
R22682 a_n2848_n452.n5 a_n2848_n452.n6 70.3058
R22683 a_n2848_n452.n3 a_n2848_n452.n62 81.4626
R22684 a_n2848_n452.n4 a_n2848_n452.n56 81.4626
R22685 a_n2848_n452.n0 a_n2848_n452.n53 81.4626
R22686 a_n2848_n452.n3 a_n2848_n452.n63 80.9324
R22687 a_n2848_n452.n2 a_n2848_n452.n64 80.9324
R22688 a_n2848_n452.n2 a_n2848_n452.n61 80.9324
R22689 a_n2848_n452.n2 a_n2848_n452.n60 80.9324
R22690 a_n2848_n452.n1 a_n2848_n452.n59 80.9324
R22691 a_n2848_n452.n4 a_n2848_n452.n57 80.9324
R22692 a_n2848_n452.n0 a_n2848_n452.n58 80.9324
R22693 a_n2848_n452.n0 a_n2848_n452.n55 80.9324
R22694 a_n2848_n452.n0 a_n2848_n452.n54 80.9324
R22695 a_n2848_n452.n32 a_n2848_n452.t20 74.6477
R22696 a_n2848_n452.n29 a_n2848_n452.t10 74.6477
R22697 a_n2848_n452.n31 a_n2848_n452.t26 74.2899
R22698 a_n2848_n452.n30 a_n2848_n452.t22 74.2897
R22699 a_n2848_n452.n32 a_n2848_n452.n99 70.6783
R22700 a_n2848_n452.n30 a_n2848_n452.n68 70.6783
R22701 a_n2848_n452.n29 a_n2848_n452.n67 70.6783
R22702 a_n2848_n452.n100 a_n2848_n452.n32 70.6782
R22703 a_n2848_n452.n93 a_n2848_n452.n92 48.2005
R22704 a_n2848_n452.n91 a_n2848_n452.n50 20.9683
R22705 a_n2848_n452.n97 a_n2848_n452.n52 20.9683
R22706 a_n2848_n452.n94 a_n2848_n452.n47 20.9683
R22707 a_n2848_n452.n75 a_n2848_n452.n74 48.2005
R22708 a_n2848_n452.n76 a_n2848_n452.n37 20.9683
R22709 a_n2848_n452.n72 a_n2848_n452.n71 48.2005
R22710 a_n2848_n452.n73 a_n2848_n452.n34 20.9683
R22711 a_n2848_n452.n88 a_n2848_n452.n78 48.2005
R22712 a_n2848_n452.t68 a_n2848_n452.n46 533.335
R22713 a_n2848_n452.n86 a_n2848_n452.n79 48.2005
R22714 a_n2848_n452.t73 a_n2848_n452.n44 533.335
R22715 a_n2848_n452.n84 a_n2848_n452.n80 48.2005
R22716 a_n2848_n452.t62 a_n2848_n452.n42 533.335
R22717 a_n2848_n452.n82 a_n2848_n452.n81 48.2005
R22718 a_n2848_n452.t58 a_n2848_n452.n40 533.335
R22719 a_n2848_n452.n51 a_n2848_n452.t72 533.058
R22720 a_n2848_n452.n48 a_n2848_n452.t19 533.058
R22721 a_n2848_n452.t21 a_n2848_n452.n38 533.058
R22722 a_n2848_n452.t50 a_n2848_n452.n35 533.058
R22723 a_n2848_n452.n1 a_n2848_n452.n0 33.585
R22724 a_n2848_n452.n49 a_n2848_n452.n66 35.3134
R22725 a_n2848_n452.n96 a_n2848_n452.n95 24.1005
R22726 a_n2848_n452.n95 a_n2848_n452.n65 24.1005
R22727 a_n2848_n452.n69 a_n2848_n452.n36 35.3134
R22728 a_n2848_n452.n70 a_n2848_n452.n33 35.3134
R22729 a_n2848_n452.n89 a_n2848_n452.n45 35.3134
R22730 a_n2848_n452.n87 a_n2848_n452.n43 35.3134
R22731 a_n2848_n452.n85 a_n2848_n452.n41 35.3134
R22732 a_n2848_n452.n83 a_n2848_n452.n39 35.3134
R22733 a_n2848_n452.n5 a_n2848_n452.n2 23.891
R22734 a_n2848_n452.n27 a_n2848_n452.n18 12.046
R22735 a_n2848_n452.n8 a_n2848_n452.n90 11.8414
R22736 a_n2848_n452.n98 a_n2848_n452.n5 10.5365
R22737 a_n2848_n452.n77 a_n2848_n452.n30 9.50122
R22738 a_n2848_n452.n20 a_n2848_n452.n18 7.47588
R22739 a_n2848_n452.n90 a_n2848_n452.n12 7.47588
R22740 a_n2848_n452.n77 a_n2848_n452.n21 6.70126
R22741 a_n2848_n452.n31 a_n2848_n452.n98 5.65783
R22742 a_n2848_n452.n90 a_n2848_n452.n77 5.3452
R22743 a_n2848_n452.n23 a_n2848_n452.n25 3.95126
R22744 a_n2848_n452.n11 a_n2848_n452.n7 3.95126
R22745 a_n2848_n452.n99 a_n2848_n452.t24 3.61217
R22746 a_n2848_n452.n99 a_n2848_n452.t12 3.61217
R22747 a_n2848_n452.n68 a_n2848_n452.t16 3.61217
R22748 a_n2848_n452.n68 a_n2848_n452.t8 3.61217
R22749 a_n2848_n452.n67 a_n2848_n452.t18 3.61217
R22750 a_n2848_n452.n67 a_n2848_n452.t14 3.61217
R22751 a_n2848_n452.t4 a_n2848_n452.n100 3.61217
R22752 a_n2848_n452.n100 a_n2848_n452.t6 3.61217
R22753 a_n2848_n452.n62 a_n2848_n452.t39 2.82907
R22754 a_n2848_n452.n62 a_n2848_n452.t45 2.82907
R22755 a_n2848_n452.n63 a_n2848_n452.t31 2.82907
R22756 a_n2848_n452.n63 a_n2848_n452.t46 2.82907
R22757 a_n2848_n452.n64 a_n2848_n452.t28 2.82907
R22758 a_n2848_n452.n64 a_n2848_n452.t42 2.82907
R22759 a_n2848_n452.n61 a_n2848_n452.t34 2.82907
R22760 a_n2848_n452.n61 a_n2848_n452.t2 2.82907
R22761 a_n2848_n452.n60 a_n2848_n452.t40 2.82907
R22762 a_n2848_n452.n60 a_n2848_n452.t41 2.82907
R22763 a_n2848_n452.n59 a_n2848_n452.t30 2.82907
R22764 a_n2848_n452.n59 a_n2848_n452.t47 2.82907
R22765 a_n2848_n452.n56 a_n2848_n452.t43 2.82907
R22766 a_n2848_n452.n56 a_n2848_n452.t33 2.82907
R22767 a_n2848_n452.n57 a_n2848_n452.t29 2.82907
R22768 a_n2848_n452.n57 a_n2848_n452.t37 2.82907
R22769 a_n2848_n452.n58 a_n2848_n452.t35 2.82907
R22770 a_n2848_n452.n58 a_n2848_n452.t36 2.82907
R22771 a_n2848_n452.n55 a_n2848_n452.t0 2.82907
R22772 a_n2848_n452.n55 a_n2848_n452.t1 2.82907
R22773 a_n2848_n452.n54 a_n2848_n452.t38 2.82907
R22774 a_n2848_n452.n54 a_n2848_n452.t32 2.82907
R22775 a_n2848_n452.n53 a_n2848_n452.t27 2.82907
R22776 a_n2848_n452.n53 a_n2848_n452.t44 2.82907
R22777 a_n2848_n452.n98 a_n2848_n452.n18 1.30542
R22778 a_n2848_n452.n15 a_n2848_n452.n16 1.04595
R22779 a_n2848_n452.n10 a_n2848_n452.n93 13.657
R22780 a_n2848_n452.n91 a_n2848_n452.n51 21.4216
R22781 a_n2848_n452.n6 a_n2848_n452.n97 21.4216
R22782 a_n2848_n452.n94 a_n2848_n452.n48 21.4216
R22783 a_n2848_n452.n74 a_n2848_n452.n24 13.657
R22784 a_n2848_n452.n38 a_n2848_n452.n76 21.4216
R22785 a_n2848_n452.n71 a_n2848_n452.n28 13.657
R22786 a_n2848_n452.n35 a_n2848_n452.n73 21.4216
R22787 a_n2848_n452.n0 a_n2848_n452.n4 1.59102
R22788 a_n2848_n452.n5 a_n2848_n452.n11 1.47777
R22789 a_n2848_n452.n2 a_n2848_n452.n3 1.06084
R22790 a_n2848_n452.n2 a_n2848_n452.n1 1.06084
R22791 a_n2848_n452.n27 a_n2848_n452.n26 0.758076
R22792 a_n2848_n452.n26 a_n2848_n452.n25 0.758076
R22793 a_n2848_n452.n23 a_n2848_n452.n22 0.758076
R22794 a_n2848_n452.n22 a_n2848_n452.n21 0.758076
R22795 a_n2848_n452.n20 a_n2848_n452.n19 0.758076
R22796 a_n2848_n452.n17 a_n2848_n452.n16 0.758076
R22797 a_n2848_n452.n15 a_n2848_n452.n14 0.758076
R22798 a_n2848_n452.n13 a_n2848_n452.n12 0.758076
R22799 a_n2848_n452.n9 a_n2848_n452.n7 0.758076
R22800 a_n2848_n452.n9 a_n2848_n452.n8 0.758076
R22801 a_n2848_n452.n32 a_n2848_n452.n31 0.716017
R22802 a_n2848_n452.n30 a_n2848_n452.n29 0.716017
R22803 a_n2848_n452.n17 a_n2848_n452.n19 0.67853
R22804 a_n2848_n452.n13 a_n2848_n452.n14 0.67853
R22805 a_n1808_13878.n17 a_n1808_13878.n16 98.9632
R22806 a_n1808_13878.n2 a_n1808_13878.n0 98.7517
R22807 a_n1808_13878.n16 a_n1808_13878.n15 98.6055
R22808 a_n1808_13878.n4 a_n1808_13878.n3 98.6055
R22809 a_n1808_13878.n2 a_n1808_13878.n1 98.6055
R22810 a_n1808_13878.n14 a_n1808_13878.n13 98.6054
R22811 a_n1808_13878.n6 a_n1808_13878.t13 74.6477
R22812 a_n1808_13878.n11 a_n1808_13878.t14 74.2899
R22813 a_n1808_13878.n8 a_n1808_13878.t15 74.2899
R22814 a_n1808_13878.n7 a_n1808_13878.t12 74.2899
R22815 a_n1808_13878.n10 a_n1808_13878.n9 70.6783
R22816 a_n1808_13878.n6 a_n1808_13878.n5 70.6783
R22817 a_n1808_13878.n12 a_n1808_13878.n4 13.5694
R22818 a_n1808_13878.n14 a_n1808_13878.n12 11.5762
R22819 a_n1808_13878.n12 a_n1808_13878.n11 6.2408
R22820 a_n1808_13878.n13 a_n1808_13878.t9 3.61217
R22821 a_n1808_13878.n13 a_n1808_13878.t10 3.61217
R22822 a_n1808_13878.n15 a_n1808_13878.t0 3.61217
R22823 a_n1808_13878.n15 a_n1808_13878.t5 3.61217
R22824 a_n1808_13878.n9 a_n1808_13878.t18 3.61217
R22825 a_n1808_13878.n9 a_n1808_13878.t19 3.61217
R22826 a_n1808_13878.n5 a_n1808_13878.t16 3.61217
R22827 a_n1808_13878.n5 a_n1808_13878.t17 3.61217
R22828 a_n1808_13878.n3 a_n1808_13878.t6 3.61217
R22829 a_n1808_13878.n3 a_n1808_13878.t1 3.61217
R22830 a_n1808_13878.n1 a_n1808_13878.t8 3.61217
R22831 a_n1808_13878.n1 a_n1808_13878.t3 3.61217
R22832 a_n1808_13878.n0 a_n1808_13878.t2 3.61217
R22833 a_n1808_13878.n0 a_n1808_13878.t4 3.61217
R22834 a_n1808_13878.n17 a_n1808_13878.t7 3.61217
R22835 a_n1808_13878.t11 a_n1808_13878.n17 3.61217
R22836 a_n1808_13878.n7 a_n1808_13878.n6 0.358259
R22837 a_n1808_13878.n10 a_n1808_13878.n8 0.358259
R22838 a_n1808_13878.n11 a_n1808_13878.n10 0.358259
R22839 a_n1808_13878.n16 a_n1808_13878.n14 0.358259
R22840 a_n1808_13878.n4 a_n1808_13878.n2 0.146627
R22841 a_n1808_13878.n8 a_n1808_13878.n7 0.101793
R22842 plus.n76 plus.t11 250.337
R22843 plus.n15 plus.t14 250.337
R22844 plus.n124 plus.t1 243.97
R22845 plus.n120 plus.t24 231.093
R22846 plus.n59 plus.t20 231.093
R22847 plus.n124 plus.n123 223.454
R22848 plus.n126 plus.n125 223.454
R22849 plus.n77 plus.t5 187.445
R22850 plus.n74 plus.t22 187.445
R22851 plus.n72 plus.t21 187.445
R22852 plus.n89 plus.t16 187.445
R22853 plus.n95 plus.t17 187.445
R22854 plus.n68 plus.t13 187.445
R22855 plus.n66 plus.t15 187.445
R22856 plus.n107 plus.t10 187.445
R22857 plus.n113 plus.t26 187.445
R22858 plus.n62 plus.t28 187.445
R22859 plus.n1 plus.t23 187.445
R22860 plus.n52 plus.t6 187.445
R22861 plus.n46 plus.t12 187.445
R22862 plus.n5 plus.t8 187.445
R22863 plus.n7 plus.t7 187.445
R22864 plus.n34 plus.t19 187.445
R22865 plus.n28 plus.t18 187.445
R22866 plus.n11 plus.t27 187.445
R22867 plus.n13 plus.t25 187.445
R22868 plus.n16 plus.t9 187.445
R22869 plus.n121 plus.n120 161.3
R22870 plus.n119 plus.n61 161.3
R22871 plus.n118 plus.n117 161.3
R22872 plus.n116 plus.n115 161.3
R22873 plus.n114 plus.n63 161.3
R22874 plus.n112 plus.n111 161.3
R22875 plus.n110 plus.n64 161.3
R22876 plus.n109 plus.n108 161.3
R22877 plus.n106 plus.n65 161.3
R22878 plus.n105 plus.n104 161.3
R22879 plus.n103 plus.n102 161.3
R22880 plus.n101 plus.n67 161.3
R22881 plus.n100 plus.n99 161.3
R22882 plus.n98 plus.n97 161.3
R22883 plus.n96 plus.n69 161.3
R22884 plus.n94 plus.n93 161.3
R22885 plus.n92 plus.n70 161.3
R22886 plus.n91 plus.n90 161.3
R22887 plus.n88 plus.n71 161.3
R22888 plus.n87 plus.n86 161.3
R22889 plus.n85 plus.n84 161.3
R22890 plus.n83 plus.n73 161.3
R22891 plus.n82 plus.n81 161.3
R22892 plus.n80 plus.n79 161.3
R22893 plus.n78 plus.n75 161.3
R22894 plus.n17 plus.n14 161.3
R22895 plus.n19 plus.n18 161.3
R22896 plus.n21 plus.n20 161.3
R22897 plus.n22 plus.n12 161.3
R22898 plus.n24 plus.n23 161.3
R22899 plus.n26 plus.n25 161.3
R22900 plus.n27 plus.n10 161.3
R22901 plus.n30 plus.n29 161.3
R22902 plus.n31 plus.n9 161.3
R22903 plus.n33 plus.n32 161.3
R22904 plus.n35 plus.n8 161.3
R22905 plus.n37 plus.n36 161.3
R22906 plus.n39 plus.n38 161.3
R22907 plus.n40 plus.n6 161.3
R22908 plus.n42 plus.n41 161.3
R22909 plus.n44 plus.n43 161.3
R22910 plus.n45 plus.n4 161.3
R22911 plus.n48 plus.n47 161.3
R22912 plus.n49 plus.n3 161.3
R22913 plus.n51 plus.n50 161.3
R22914 plus.n53 plus.n2 161.3
R22915 plus.n55 plus.n54 161.3
R22916 plus.n57 plus.n56 161.3
R22917 plus.n58 plus.n0 161.3
R22918 plus.n60 plus.n59 161.3
R22919 plus.n88 plus.n87 56.5617
R22920 plus.n97 plus.n96 56.5617
R22921 plus.n106 plus.n105 56.5617
R22922 plus.n45 plus.n44 56.5617
R22923 plus.n36 plus.n35 56.5617
R22924 plus.n27 plus.n26 56.5617
R22925 plus.n79 plus.n78 56.5617
R22926 plus.n115 plus.n114 56.5617
R22927 plus.n54 plus.n53 56.5617
R22928 plus.n18 plus.n17 56.5617
R22929 plus.n119 plus.n118 50.2647
R22930 plus.n58 plus.n57 50.2647
R22931 plus.n84 plus.n83 46.3896
R22932 plus.n108 plus.n64 46.3896
R22933 plus.n47 plus.n3 46.3896
R22934 plus.n23 plus.n22 46.3896
R22935 plus.n76 plus.n75 43.1929
R22936 plus.n15 plus.n14 43.1929
R22937 plus.n94 plus.n70 42.5146
R22938 plus.n101 plus.n100 42.5146
R22939 plus.n40 plus.n39 42.5146
R22940 plus.n33 plus.n9 42.5146
R22941 plus.n77 plus.n76 40.6041
R22942 plus.n16 plus.n15 40.6041
R22943 plus.n90 plus.n70 38.6395
R22944 plus.n102 plus.n101 38.6395
R22945 plus.n41 plus.n40 38.6395
R22946 plus.n29 plus.n9 38.6395
R22947 plus.n122 plus.n121 35.2031
R22948 plus.n83 plus.n82 34.7644
R22949 plus.n112 plus.n64 34.7644
R22950 plus.n51 plus.n3 34.7644
R22951 plus.n22 plus.n21 34.7644
R22952 plus.n79 plus.n74 21.8872
R22953 plus.n114 plus.n113 21.8872
R22954 plus.n53 plus.n52 21.8872
R22955 plus.n18 plus.n13 21.8872
R22956 plus.n89 plus.n88 19.9199
R22957 plus.n105 plus.n66 19.9199
R22958 plus.n44 plus.n5 19.9199
R22959 plus.n28 plus.n27 19.9199
R22960 plus.n123 plus.t2 19.8005
R22961 plus.n123 plus.t4 19.8005
R22962 plus.n125 plus.t3 19.8005
R22963 plus.n125 plus.t0 19.8005
R22964 plus.n96 plus.n95 17.9525
R22965 plus.n97 plus.n68 17.9525
R22966 plus.n36 plus.n7 17.9525
R22967 plus.n35 plus.n34 17.9525
R22968 plus.n87 plus.n72 15.9852
R22969 plus.n107 plus.n106 15.9852
R22970 plus.n46 plus.n45 15.9852
R22971 plus.n26 plus.n11 15.9852
R22972 plus plus.n127 15.0253
R22973 plus.n78 plus.n77 14.0178
R22974 plus.n115 plus.n62 14.0178
R22975 plus.n54 plus.n1 14.0178
R22976 plus.n17 plus.n16 14.0178
R22977 plus.n122 plus.n60 11.9342
R22978 plus.n118 plus.n62 10.575
R22979 plus.n57 plus.n1 10.575
R22980 plus.n120 plus.n119 9.49444
R22981 plus.n59 plus.n58 9.49444
R22982 plus.n84 plus.n72 8.60764
R22983 plus.n108 plus.n107 8.60764
R22984 plus.n47 plus.n46 8.60764
R22985 plus.n23 plus.n11 8.60764
R22986 plus.n95 plus.n94 6.6403
R22987 plus.n100 plus.n68 6.6403
R22988 plus.n39 plus.n7 6.6403
R22989 plus.n34 plus.n33 6.6403
R22990 plus.n127 plus.n126 5.40567
R22991 plus.n90 plus.n89 4.67295
R22992 plus.n102 plus.n66 4.67295
R22993 plus.n41 plus.n5 4.67295
R22994 plus.n29 plus.n28 4.67295
R22995 plus.n82 plus.n74 2.7056
R22996 plus.n113 plus.n112 2.7056
R22997 plus.n52 plus.n51 2.7056
R22998 plus.n21 plus.n13 2.7056
R22999 plus.n127 plus.n122 1.188
R23000 plus.n126 plus.n124 0.716017
R23001 plus.n80 plus.n75 0.189894
R23002 plus.n81 plus.n80 0.189894
R23003 plus.n81 plus.n73 0.189894
R23004 plus.n85 plus.n73 0.189894
R23005 plus.n86 plus.n85 0.189894
R23006 plus.n86 plus.n71 0.189894
R23007 plus.n91 plus.n71 0.189894
R23008 plus.n92 plus.n91 0.189894
R23009 plus.n93 plus.n92 0.189894
R23010 plus.n93 plus.n69 0.189894
R23011 plus.n98 plus.n69 0.189894
R23012 plus.n99 plus.n98 0.189894
R23013 plus.n99 plus.n67 0.189894
R23014 plus.n103 plus.n67 0.189894
R23015 plus.n104 plus.n103 0.189894
R23016 plus.n104 plus.n65 0.189894
R23017 plus.n109 plus.n65 0.189894
R23018 plus.n110 plus.n109 0.189894
R23019 plus.n111 plus.n110 0.189894
R23020 plus.n111 plus.n63 0.189894
R23021 plus.n116 plus.n63 0.189894
R23022 plus.n117 plus.n116 0.189894
R23023 plus.n117 plus.n61 0.189894
R23024 plus.n121 plus.n61 0.189894
R23025 plus.n60 plus.n0 0.189894
R23026 plus.n56 plus.n0 0.189894
R23027 plus.n56 plus.n55 0.189894
R23028 plus.n55 plus.n2 0.189894
R23029 plus.n50 plus.n2 0.189894
R23030 plus.n50 plus.n49 0.189894
R23031 plus.n49 plus.n48 0.189894
R23032 plus.n48 plus.n4 0.189894
R23033 plus.n43 plus.n4 0.189894
R23034 plus.n43 plus.n42 0.189894
R23035 plus.n42 plus.n6 0.189894
R23036 plus.n38 plus.n6 0.189894
R23037 plus.n38 plus.n37 0.189894
R23038 plus.n37 plus.n8 0.189894
R23039 plus.n32 plus.n8 0.189894
R23040 plus.n32 plus.n31 0.189894
R23041 plus.n31 plus.n30 0.189894
R23042 plus.n30 plus.n10 0.189894
R23043 plus.n25 plus.n10 0.189894
R23044 plus.n25 plus.n24 0.189894
R23045 plus.n24 plus.n12 0.189894
R23046 plus.n20 plus.n12 0.189894
R23047 plus.n20 plus.n19 0.189894
R23048 plus.n19 plus.n14 0.189894
R23049 a_n3827_n3924.n26 a_n3827_n3924.t13 214.938
R23050 a_n3827_n3924.n35 a_n3827_n3924.t7 214.409
R23051 a_n3827_n3924.n34 a_n3827_n3924.t23 214.321
R23052 a_n3827_n3924.n33 a_n3827_n3924.t3 214.321
R23053 a_n3827_n3924.n32 a_n3827_n3924.t6 214.321
R23054 a_n3827_n3924.n31 a_n3827_n3924.t28 214.321
R23055 a_n3827_n3924.n30 a_n3827_n3924.t1 214.321
R23056 a_n3827_n3924.n29 a_n3827_n3924.t22 214.321
R23057 a_n3827_n3924.n28 a_n3827_n3924.t0 214.321
R23058 a_n3827_n3924.n27 a_n3827_n3924.t20 214.321
R23059 a_n3827_n3924.n12 a_n3827_n3924.t51 55.8337
R23060 a_n3827_n3924.n13 a_n3827_n3924.t31 55.8337
R23061 a_n3827_n3924.n24 a_n3827_n3924.t11 55.8337
R23062 a_n3827_n3924.n1 a_n3827_n3924.t38 55.8335
R23063 a_n3827_n3924.n37 a_n3827_n3924.t15 55.8335
R23064 a_n3827_n3924.n48 a_n3827_n3924.t8 55.8335
R23065 a_n3827_n3924.n49 a_n3827_n3924.t48 55.8335
R23066 a_n3827_n3924.n0 a_n3827_n3924.t42 55.8335
R23067 a_n3827_n3924.n59 a_n3827_n3924.n58 53.0054
R23068 a_n3827_n3924.n3 a_n3827_n3924.n2 53.0052
R23069 a_n3827_n3924.n5 a_n3827_n3924.n4 53.0052
R23070 a_n3827_n3924.n7 a_n3827_n3924.n6 53.0052
R23071 a_n3827_n3924.n9 a_n3827_n3924.n8 53.0052
R23072 a_n3827_n3924.n11 a_n3827_n3924.n10 53.0052
R23073 a_n3827_n3924.n15 a_n3827_n3924.n14 53.0052
R23074 a_n3827_n3924.n17 a_n3827_n3924.n16 53.0052
R23075 a_n3827_n3924.n19 a_n3827_n3924.n18 53.0052
R23076 a_n3827_n3924.n21 a_n3827_n3924.n20 53.0052
R23077 a_n3827_n3924.n23 a_n3827_n3924.n22 53.0052
R23078 a_n3827_n3924.n39 a_n3827_n3924.n38 53.0051
R23079 a_n3827_n3924.n41 a_n3827_n3924.n40 53.0051
R23080 a_n3827_n3924.n43 a_n3827_n3924.n42 53.0051
R23081 a_n3827_n3924.n45 a_n3827_n3924.n44 53.0051
R23082 a_n3827_n3924.n47 a_n3827_n3924.n46 53.0051
R23083 a_n3827_n3924.n51 a_n3827_n3924.n50 53.0051
R23084 a_n3827_n3924.n53 a_n3827_n3924.n52 53.0051
R23085 a_n3827_n3924.n55 a_n3827_n3924.n54 53.0051
R23086 a_n3827_n3924.n57 a_n3827_n3924.n56 53.0051
R23087 a_n3827_n3924.n25 a_n3827_n3924.n24 12.2417
R23088 a_n3827_n3924.n36 a_n3827_n3924.n1 12.2417
R23089 a_n3827_n3924.n25 a_n3827_n3924.n0 5.16214
R23090 a_n3827_n3924.n37 a_n3827_n3924.n36 5.16214
R23091 a_n3827_n3924.n38 a_n3827_n3924.t19 2.82907
R23092 a_n3827_n3924.n38 a_n3827_n3924.t29 2.82907
R23093 a_n3827_n3924.n40 a_n3827_n3924.t18 2.82907
R23094 a_n3827_n3924.n40 a_n3827_n3924.t10 2.82907
R23095 a_n3827_n3924.n42 a_n3827_n3924.t4 2.82907
R23096 a_n3827_n3924.n42 a_n3827_n3924.t17 2.82907
R23097 a_n3827_n3924.n44 a_n3827_n3924.t14 2.82907
R23098 a_n3827_n3924.n44 a_n3827_n3924.t2 2.82907
R23099 a_n3827_n3924.n46 a_n3827_n3924.t30 2.82907
R23100 a_n3827_n3924.n46 a_n3827_n3924.t21 2.82907
R23101 a_n3827_n3924.n50 a_n3827_n3924.t37 2.82907
R23102 a_n3827_n3924.n50 a_n3827_n3924.t53 2.82907
R23103 a_n3827_n3924.n52 a_n3827_n3924.t44 2.82907
R23104 a_n3827_n3924.n52 a_n3827_n3924.t35 2.82907
R23105 a_n3827_n3924.n54 a_n3827_n3924.t55 2.82907
R23106 a_n3827_n3924.n54 a_n3827_n3924.t43 2.82907
R23107 a_n3827_n3924.n56 a_n3827_n3924.t50 2.82907
R23108 a_n3827_n3924.n56 a_n3827_n3924.t54 2.82907
R23109 a_n3827_n3924.n2 a_n3827_n3924.t36 2.82907
R23110 a_n3827_n3924.n2 a_n3827_n3924.t34 2.82907
R23111 a_n3827_n3924.n4 a_n3827_n3924.t47 2.82907
R23112 a_n3827_n3924.n4 a_n3827_n3924.t52 2.82907
R23113 a_n3827_n3924.n6 a_n3827_n3924.t45 2.82907
R23114 a_n3827_n3924.n6 a_n3827_n3924.t49 2.82907
R23115 a_n3827_n3924.n8 a_n3827_n3924.t41 2.82907
R23116 a_n3827_n3924.n8 a_n3827_n3924.t46 2.82907
R23117 a_n3827_n3924.n10 a_n3827_n3924.t57 2.82907
R23118 a_n3827_n3924.n10 a_n3827_n3924.t40 2.82907
R23119 a_n3827_n3924.n14 a_n3827_n3924.t32 2.82907
R23120 a_n3827_n3924.n14 a_n3827_n3924.t24 2.82907
R23121 a_n3827_n3924.n16 a_n3827_n3924.t27 2.82907
R23122 a_n3827_n3924.n16 a_n3827_n3924.t12 2.82907
R23123 a_n3827_n3924.n18 a_n3827_n3924.t5 2.82907
R23124 a_n3827_n3924.n18 a_n3827_n3924.t9 2.82907
R23125 a_n3827_n3924.n20 a_n3827_n3924.t26 2.82907
R23126 a_n3827_n3924.n20 a_n3827_n3924.t16 2.82907
R23127 a_n3827_n3924.n22 a_n3827_n3924.t33 2.82907
R23128 a_n3827_n3924.n22 a_n3827_n3924.t25 2.82907
R23129 a_n3827_n3924.n59 a_n3827_n3924.t39 2.82907
R23130 a_n3827_n3924.t56 a_n3827_n3924.n59 2.82907
R23131 a_n3827_n3924.n26 a_n3827_n3924.n25 1.95694
R23132 a_n3827_n3924.n36 a_n3827_n3924.n35 1.95694
R23133 a_n3827_n3924.n28 a_n3827_n3924.n27 0.672012
R23134 a_n3827_n3924.n29 a_n3827_n3924.n28 0.672012
R23135 a_n3827_n3924.n30 a_n3827_n3924.n29 0.672012
R23136 a_n3827_n3924.n31 a_n3827_n3924.n30 0.672012
R23137 a_n3827_n3924.n32 a_n3827_n3924.n31 0.672012
R23138 a_n3827_n3924.n33 a_n3827_n3924.n32 0.672012
R23139 a_n3827_n3924.n34 a_n3827_n3924.n33 0.672012
R23140 a_n3827_n3924.n35 a_n3827_n3924.n34 0.585529
R23141 a_n3827_n3924.n24 a_n3827_n3924.n23 0.530672
R23142 a_n3827_n3924.n23 a_n3827_n3924.n21 0.530672
R23143 a_n3827_n3924.n21 a_n3827_n3924.n19 0.530672
R23144 a_n3827_n3924.n19 a_n3827_n3924.n17 0.530672
R23145 a_n3827_n3924.n17 a_n3827_n3924.n15 0.530672
R23146 a_n3827_n3924.n15 a_n3827_n3924.n13 0.530672
R23147 a_n3827_n3924.n12 a_n3827_n3924.n11 0.530672
R23148 a_n3827_n3924.n11 a_n3827_n3924.n9 0.530672
R23149 a_n3827_n3924.n9 a_n3827_n3924.n7 0.530672
R23150 a_n3827_n3924.n7 a_n3827_n3924.n5 0.530672
R23151 a_n3827_n3924.n5 a_n3827_n3924.n3 0.530672
R23152 a_n3827_n3924.n3 a_n3827_n3924.n1 0.530672
R23153 a_n3827_n3924.n58 a_n3827_n3924.n0 0.530672
R23154 a_n3827_n3924.n58 a_n3827_n3924.n57 0.530672
R23155 a_n3827_n3924.n57 a_n3827_n3924.n55 0.530672
R23156 a_n3827_n3924.n55 a_n3827_n3924.n53 0.530672
R23157 a_n3827_n3924.n53 a_n3827_n3924.n51 0.530672
R23158 a_n3827_n3924.n51 a_n3827_n3924.n49 0.530672
R23159 a_n3827_n3924.n48 a_n3827_n3924.n47 0.530672
R23160 a_n3827_n3924.n47 a_n3827_n3924.n45 0.530672
R23161 a_n3827_n3924.n45 a_n3827_n3924.n43 0.530672
R23162 a_n3827_n3924.n43 a_n3827_n3924.n41 0.530672
R23163 a_n3827_n3924.n41 a_n3827_n3924.n39 0.530672
R23164 a_n3827_n3924.n39 a_n3827_n3924.n37 0.530672
R23165 a_n3827_n3924.n13 a_n3827_n3924.n12 0.235414
R23166 a_n3827_n3924.n49 a_n3827_n3924.n48 0.235414
R23167 a_n3827_n3924.n27 a_n3827_n3924.n26 0.0564593
R23168 diffpairibias.n0 diffpairibias.t27 436.822
R23169 diffpairibias.n27 diffpairibias.t24 435.479
R23170 diffpairibias.n26 diffpairibias.t21 435.479
R23171 diffpairibias.n25 diffpairibias.t22 435.479
R23172 diffpairibias.n24 diffpairibias.t26 435.479
R23173 diffpairibias.n23 diffpairibias.t20 435.479
R23174 diffpairibias.n0 diffpairibias.t23 435.479
R23175 diffpairibias.n1 diffpairibias.t28 435.479
R23176 diffpairibias.n2 diffpairibias.t25 435.479
R23177 diffpairibias.n3 diffpairibias.t29 435.479
R23178 diffpairibias.n13 diffpairibias.t14 377.536
R23179 diffpairibias.n13 diffpairibias.t0 376.193
R23180 diffpairibias.n14 diffpairibias.t10 376.193
R23181 diffpairibias.n15 diffpairibias.t12 376.193
R23182 diffpairibias.n16 diffpairibias.t6 376.193
R23183 diffpairibias.n17 diffpairibias.t2 376.193
R23184 diffpairibias.n18 diffpairibias.t16 376.193
R23185 diffpairibias.n19 diffpairibias.t4 376.193
R23186 diffpairibias.n20 diffpairibias.t18 376.193
R23187 diffpairibias.n21 diffpairibias.t8 376.193
R23188 diffpairibias.n4 diffpairibias.t15 113.368
R23189 diffpairibias.n4 diffpairibias.t1 112.698
R23190 diffpairibias.n5 diffpairibias.t11 112.698
R23191 diffpairibias.n6 diffpairibias.t13 112.698
R23192 diffpairibias.n7 diffpairibias.t7 112.698
R23193 diffpairibias.n8 diffpairibias.t3 112.698
R23194 diffpairibias.n9 diffpairibias.t17 112.698
R23195 diffpairibias.n10 diffpairibias.t5 112.698
R23196 diffpairibias.n11 diffpairibias.t19 112.698
R23197 diffpairibias.n12 diffpairibias.t9 112.698
R23198 diffpairibias.n22 diffpairibias.n21 4.77242
R23199 diffpairibias.n22 diffpairibias.n12 4.30807
R23200 diffpairibias.n23 diffpairibias.n22 4.13945
R23201 diffpairibias.n21 diffpairibias.n20 1.34352
R23202 diffpairibias.n20 diffpairibias.n19 1.34352
R23203 diffpairibias.n19 diffpairibias.n18 1.34352
R23204 diffpairibias.n18 diffpairibias.n17 1.34352
R23205 diffpairibias.n17 diffpairibias.n16 1.34352
R23206 diffpairibias.n16 diffpairibias.n15 1.34352
R23207 diffpairibias.n15 diffpairibias.n14 1.34352
R23208 diffpairibias.n14 diffpairibias.n13 1.34352
R23209 diffpairibias.n3 diffpairibias.n2 1.34352
R23210 diffpairibias.n2 diffpairibias.n1 1.34352
R23211 diffpairibias.n1 diffpairibias.n0 1.34352
R23212 diffpairibias.n24 diffpairibias.n23 1.34352
R23213 diffpairibias.n25 diffpairibias.n24 1.34352
R23214 diffpairibias.n26 diffpairibias.n25 1.34352
R23215 diffpairibias.n27 diffpairibias.n26 1.34352
R23216 diffpairibias.n28 diffpairibias.n27 0.862419
R23217 diffpairibias diffpairibias.n28 0.684875
R23218 diffpairibias.n12 diffpairibias.n11 0.672012
R23219 diffpairibias.n11 diffpairibias.n10 0.672012
R23220 diffpairibias.n10 diffpairibias.n9 0.672012
R23221 diffpairibias.n9 diffpairibias.n8 0.672012
R23222 diffpairibias.n8 diffpairibias.n7 0.672012
R23223 diffpairibias.n7 diffpairibias.n6 0.672012
R23224 diffpairibias.n6 diffpairibias.n5 0.672012
R23225 diffpairibias.n5 diffpairibias.n4 0.672012
R23226 diffpairibias.n28 diffpairibias.n3 0.190907
R23227 a_n1986_8322.n6 a_n1986_8322.t15 74.6477
R23228 a_n1986_8322.n1 a_n1986_8322.t1 74.6477
R23229 a_n1986_8322.n16 a_n1986_8322.t10 74.6474
R23230 a_n1986_8322.n14 a_n1986_8322.t3 74.2899
R23231 a_n1986_8322.n7 a_n1986_8322.t13 74.2899
R23232 a_n1986_8322.n8 a_n1986_8322.t16 74.2899
R23233 a_n1986_8322.n11 a_n1986_8322.t17 74.2899
R23234 a_n1986_8322.n4 a_n1986_8322.t0 74.2899
R23235 a_n1986_8322.n16 a_n1986_8322.n15 70.6783
R23236 a_n1986_8322.n6 a_n1986_8322.n5 70.6783
R23237 a_n1986_8322.n10 a_n1986_8322.n9 70.6783
R23238 a_n1986_8322.n1 a_n1986_8322.n0 70.6783
R23239 a_n1986_8322.n3 a_n1986_8322.n2 70.6783
R23240 a_n1986_8322.n18 a_n1986_8322.n17 70.6782
R23241 a_n1986_8322.n12 a_n1986_8322.n4 22.7556
R23242 a_n1986_8322.n13 a_n1986_8322.t20 10.109
R23243 a_n1986_8322.n12 a_n1986_8322.n11 6.2408
R23244 a_n1986_8322.n14 a_n1986_8322.n13 5.83671
R23245 a_n1986_8322.n13 a_n1986_8322.n12 5.3452
R23246 a_n1986_8322.n15 a_n1986_8322.t8 3.61217
R23247 a_n1986_8322.n15 a_n1986_8322.t5 3.61217
R23248 a_n1986_8322.n5 a_n1986_8322.t19 3.61217
R23249 a_n1986_8322.n5 a_n1986_8322.t18 3.61217
R23250 a_n1986_8322.n9 a_n1986_8322.t14 3.61217
R23251 a_n1986_8322.n9 a_n1986_8322.t12 3.61217
R23252 a_n1986_8322.n0 a_n1986_8322.t9 3.61217
R23253 a_n1986_8322.n0 a_n1986_8322.t4 3.61217
R23254 a_n1986_8322.n2 a_n1986_8322.t7 3.61217
R23255 a_n1986_8322.n2 a_n1986_8322.t6 3.61217
R23256 a_n1986_8322.n18 a_n1986_8322.t2 3.61217
R23257 a_n1986_8322.t11 a_n1986_8322.n18 3.61217
R23258 a_n1986_8322.n11 a_n1986_8322.n10 0.358259
R23259 a_n1986_8322.n10 a_n1986_8322.n8 0.358259
R23260 a_n1986_8322.n7 a_n1986_8322.n6 0.358259
R23261 a_n1986_8322.n4 a_n1986_8322.n3 0.358259
R23262 a_n1986_8322.n3 a_n1986_8322.n1 0.358259
R23263 a_n1986_8322.n17 a_n1986_8322.n14 0.358259
R23264 a_n1986_8322.n17 a_n1986_8322.n16 0.358259
R23265 a_n1986_8322.n8 a_n1986_8322.n7 0.101793
R23266 a_n1986_8322.t20 a_n1986_8322.t21 0.057021
R23267 minus.n76 minus.t28 250.337
R23268 minus.n15 minus.t20 250.337
R23269 minus.n126 minus.t1 243.255
R23270 minus.n120 minus.t8 231.093
R23271 minus.n59 minus.t10 231.093
R23272 minus.n125 minus.n123 224.169
R23273 minus.n125 minus.n124 223.454
R23274 minus.n62 minus.t12 187.445
R23275 minus.n113 minus.t18 187.445
R23276 minus.n107 minus.t25 187.445
R23277 minus.n66 minus.t22 187.445
R23278 minus.n68 minus.t19 187.445
R23279 minus.n95 minus.t7 187.445
R23280 minus.n89 minus.t6 187.445
R23281 minus.n72 minus.t16 187.445
R23282 minus.n74 minus.t15 187.445
R23283 minus.n77 minus.t23 187.445
R23284 minus.n16 minus.t14 187.445
R23285 minus.n13 minus.t9 187.445
R23286 minus.n11 minus.t5 187.445
R23287 minus.n28 minus.t26 187.445
R23288 minus.n34 minus.t27 187.445
R23289 minus.n7 minus.t21 187.445
R23290 minus.n5 minus.t24 187.445
R23291 minus.n46 minus.t17 187.445
R23292 minus.n52 minus.t11 187.445
R23293 minus.n1 minus.t13 187.445
R23294 minus.n78 minus.n75 161.3
R23295 minus.n80 minus.n79 161.3
R23296 minus.n82 minus.n81 161.3
R23297 minus.n83 minus.n73 161.3
R23298 minus.n85 minus.n84 161.3
R23299 minus.n87 minus.n86 161.3
R23300 minus.n88 minus.n71 161.3
R23301 minus.n91 minus.n90 161.3
R23302 minus.n92 minus.n70 161.3
R23303 minus.n94 minus.n93 161.3
R23304 minus.n96 minus.n69 161.3
R23305 minus.n98 minus.n97 161.3
R23306 minus.n100 minus.n99 161.3
R23307 minus.n101 minus.n67 161.3
R23308 minus.n103 minus.n102 161.3
R23309 minus.n105 minus.n104 161.3
R23310 minus.n106 minus.n65 161.3
R23311 minus.n109 minus.n108 161.3
R23312 minus.n110 minus.n64 161.3
R23313 minus.n112 minus.n111 161.3
R23314 minus.n114 minus.n63 161.3
R23315 minus.n116 minus.n115 161.3
R23316 minus.n118 minus.n117 161.3
R23317 minus.n119 minus.n61 161.3
R23318 minus.n121 minus.n120 161.3
R23319 minus.n60 minus.n59 161.3
R23320 minus.n58 minus.n0 161.3
R23321 minus.n57 minus.n56 161.3
R23322 minus.n55 minus.n54 161.3
R23323 minus.n53 minus.n2 161.3
R23324 minus.n51 minus.n50 161.3
R23325 minus.n49 minus.n3 161.3
R23326 minus.n48 minus.n47 161.3
R23327 minus.n45 minus.n4 161.3
R23328 minus.n44 minus.n43 161.3
R23329 minus.n42 minus.n41 161.3
R23330 minus.n40 minus.n6 161.3
R23331 minus.n39 minus.n38 161.3
R23332 minus.n37 minus.n36 161.3
R23333 minus.n35 minus.n8 161.3
R23334 minus.n33 minus.n32 161.3
R23335 minus.n31 minus.n9 161.3
R23336 minus.n30 minus.n29 161.3
R23337 minus.n27 minus.n10 161.3
R23338 minus.n26 minus.n25 161.3
R23339 minus.n24 minus.n23 161.3
R23340 minus.n22 minus.n12 161.3
R23341 minus.n21 minus.n20 161.3
R23342 minus.n19 minus.n18 161.3
R23343 minus.n17 minus.n14 161.3
R23344 minus.n106 minus.n105 56.5617
R23345 minus.n97 minus.n96 56.5617
R23346 minus.n88 minus.n87 56.5617
R23347 minus.n27 minus.n26 56.5617
R23348 minus.n36 minus.n35 56.5617
R23349 minus.n45 minus.n44 56.5617
R23350 minus.n115 minus.n114 56.5617
R23351 minus.n79 minus.n78 56.5617
R23352 minus.n18 minus.n17 56.5617
R23353 minus.n54 minus.n53 56.5617
R23354 minus.n119 minus.n118 50.2647
R23355 minus.n58 minus.n57 50.2647
R23356 minus.n108 minus.n64 46.3896
R23357 minus.n84 minus.n83 46.3896
R23358 minus.n23 minus.n22 46.3896
R23359 minus.n47 minus.n3 46.3896
R23360 minus.n76 minus.n75 43.1929
R23361 minus.n15 minus.n14 43.1929
R23362 minus.n101 minus.n100 42.5146
R23363 minus.n94 minus.n70 42.5146
R23364 minus.n33 minus.n9 42.5146
R23365 minus.n40 minus.n39 42.5146
R23366 minus.n77 minus.n76 40.6041
R23367 minus.n16 minus.n15 40.6041
R23368 minus.n102 minus.n101 38.6395
R23369 minus.n90 minus.n70 38.6395
R23370 minus.n29 minus.n9 38.6395
R23371 minus.n41 minus.n40 38.6395
R23372 minus.n122 minus.n121 35.4191
R23373 minus.n112 minus.n64 34.7644
R23374 minus.n83 minus.n82 34.7644
R23375 minus.n22 minus.n21 34.7644
R23376 minus.n51 minus.n3 34.7644
R23377 minus.n114 minus.n113 21.8872
R23378 minus.n79 minus.n74 21.8872
R23379 minus.n18 minus.n13 21.8872
R23380 minus.n53 minus.n52 21.8872
R23381 minus.n105 minus.n66 19.9199
R23382 minus.n89 minus.n88 19.9199
R23383 minus.n28 minus.n27 19.9199
R23384 minus.n44 minus.n5 19.9199
R23385 minus.n124 minus.t0 19.8005
R23386 minus.n124 minus.t2 19.8005
R23387 minus.n123 minus.t4 19.8005
R23388 minus.n123 minus.t3 19.8005
R23389 minus.n97 minus.n68 17.9525
R23390 minus.n96 minus.n95 17.9525
R23391 minus.n35 minus.n34 17.9525
R23392 minus.n36 minus.n7 17.9525
R23393 minus.n107 minus.n106 15.9852
R23394 minus.n87 minus.n72 15.9852
R23395 minus.n26 minus.n11 15.9852
R23396 minus.n46 minus.n45 15.9852
R23397 minus.n115 minus.n62 14.0178
R23398 minus.n78 minus.n77 14.0178
R23399 minus.n17 minus.n16 14.0178
R23400 minus.n54 minus.n1 14.0178
R23401 minus.n122 minus.n60 12.1501
R23402 minus minus.n127 11.5381
R23403 minus.n118 minus.n62 10.575
R23404 minus.n57 minus.n1 10.575
R23405 minus.n120 minus.n119 9.49444
R23406 minus.n59 minus.n58 9.49444
R23407 minus.n108 minus.n107 8.60764
R23408 minus.n84 minus.n72 8.60764
R23409 minus.n23 minus.n11 8.60764
R23410 minus.n47 minus.n46 8.60764
R23411 minus.n100 minus.n68 6.6403
R23412 minus.n95 minus.n94 6.6403
R23413 minus.n34 minus.n33 6.6403
R23414 minus.n39 minus.n7 6.6403
R23415 minus.n127 minus.n126 4.80222
R23416 minus.n102 minus.n66 4.67295
R23417 minus.n90 minus.n89 4.67295
R23418 minus.n29 minus.n28 4.67295
R23419 minus.n41 minus.n5 4.67295
R23420 minus.n113 minus.n112 2.7056
R23421 minus.n82 minus.n74 2.7056
R23422 minus.n21 minus.n13 2.7056
R23423 minus.n52 minus.n51 2.7056
R23424 minus.n127 minus.n122 0.972091
R23425 minus.n126 minus.n125 0.716017
R23426 minus.n121 minus.n61 0.189894
R23427 minus.n117 minus.n61 0.189894
R23428 minus.n117 minus.n116 0.189894
R23429 minus.n116 minus.n63 0.189894
R23430 minus.n111 minus.n63 0.189894
R23431 minus.n111 minus.n110 0.189894
R23432 minus.n110 minus.n109 0.189894
R23433 minus.n109 minus.n65 0.189894
R23434 minus.n104 minus.n65 0.189894
R23435 minus.n104 minus.n103 0.189894
R23436 minus.n103 minus.n67 0.189894
R23437 minus.n99 minus.n67 0.189894
R23438 minus.n99 minus.n98 0.189894
R23439 minus.n98 minus.n69 0.189894
R23440 minus.n93 minus.n69 0.189894
R23441 minus.n93 minus.n92 0.189894
R23442 minus.n92 minus.n91 0.189894
R23443 minus.n91 minus.n71 0.189894
R23444 minus.n86 minus.n71 0.189894
R23445 minus.n86 minus.n85 0.189894
R23446 minus.n85 minus.n73 0.189894
R23447 minus.n81 minus.n73 0.189894
R23448 minus.n81 minus.n80 0.189894
R23449 minus.n80 minus.n75 0.189894
R23450 minus.n19 minus.n14 0.189894
R23451 minus.n20 minus.n19 0.189894
R23452 minus.n20 minus.n12 0.189894
R23453 minus.n24 minus.n12 0.189894
R23454 minus.n25 minus.n24 0.189894
R23455 minus.n25 minus.n10 0.189894
R23456 minus.n30 minus.n10 0.189894
R23457 minus.n31 minus.n30 0.189894
R23458 minus.n32 minus.n31 0.189894
R23459 minus.n32 minus.n8 0.189894
R23460 minus.n37 minus.n8 0.189894
R23461 minus.n38 minus.n37 0.189894
R23462 minus.n38 minus.n6 0.189894
R23463 minus.n42 minus.n6 0.189894
R23464 minus.n43 minus.n42 0.189894
R23465 minus.n43 minus.n4 0.189894
R23466 minus.n48 minus.n4 0.189894
R23467 minus.n49 minus.n48 0.189894
R23468 minus.n50 minus.n49 0.189894
R23469 minus.n50 minus.n2 0.189894
R23470 minus.n55 minus.n2 0.189894
R23471 minus.n56 minus.n55 0.189894
R23472 minus.n56 minus.n0 0.189894
R23473 minus.n60 minus.n0 0.189894
R23474 outputibias.n27 outputibias.n1 289.615
R23475 outputibias.n58 outputibias.n32 289.615
R23476 outputibias.n90 outputibias.n64 289.615
R23477 outputibias.n122 outputibias.n96 289.615
R23478 outputibias.n28 outputibias.n27 185
R23479 outputibias.n26 outputibias.n25 185
R23480 outputibias.n5 outputibias.n4 185
R23481 outputibias.n20 outputibias.n19 185
R23482 outputibias.n18 outputibias.n17 185
R23483 outputibias.n9 outputibias.n8 185
R23484 outputibias.n12 outputibias.n11 185
R23485 outputibias.n59 outputibias.n58 185
R23486 outputibias.n57 outputibias.n56 185
R23487 outputibias.n36 outputibias.n35 185
R23488 outputibias.n51 outputibias.n50 185
R23489 outputibias.n49 outputibias.n48 185
R23490 outputibias.n40 outputibias.n39 185
R23491 outputibias.n43 outputibias.n42 185
R23492 outputibias.n91 outputibias.n90 185
R23493 outputibias.n89 outputibias.n88 185
R23494 outputibias.n68 outputibias.n67 185
R23495 outputibias.n83 outputibias.n82 185
R23496 outputibias.n81 outputibias.n80 185
R23497 outputibias.n72 outputibias.n71 185
R23498 outputibias.n75 outputibias.n74 185
R23499 outputibias.n123 outputibias.n122 185
R23500 outputibias.n121 outputibias.n120 185
R23501 outputibias.n100 outputibias.n99 185
R23502 outputibias.n115 outputibias.n114 185
R23503 outputibias.n113 outputibias.n112 185
R23504 outputibias.n104 outputibias.n103 185
R23505 outputibias.n107 outputibias.n106 185
R23506 outputibias.n0 outputibias.t9 178.945
R23507 outputibias.n133 outputibias.t8 177.018
R23508 outputibias.n132 outputibias.t11 177.018
R23509 outputibias.n0 outputibias.t10 177.018
R23510 outputibias.t5 outputibias.n10 147.661
R23511 outputibias.t7 outputibias.n41 147.661
R23512 outputibias.t1 outputibias.n73 147.661
R23513 outputibias.t3 outputibias.n105 147.661
R23514 outputibias.n128 outputibias.t4 132.363
R23515 outputibias.n128 outputibias.t6 130.436
R23516 outputibias.n129 outputibias.t0 130.436
R23517 outputibias.n130 outputibias.t2 130.436
R23518 outputibias.n27 outputibias.n26 104.615
R23519 outputibias.n26 outputibias.n4 104.615
R23520 outputibias.n19 outputibias.n4 104.615
R23521 outputibias.n19 outputibias.n18 104.615
R23522 outputibias.n18 outputibias.n8 104.615
R23523 outputibias.n11 outputibias.n8 104.615
R23524 outputibias.n58 outputibias.n57 104.615
R23525 outputibias.n57 outputibias.n35 104.615
R23526 outputibias.n50 outputibias.n35 104.615
R23527 outputibias.n50 outputibias.n49 104.615
R23528 outputibias.n49 outputibias.n39 104.615
R23529 outputibias.n42 outputibias.n39 104.615
R23530 outputibias.n90 outputibias.n89 104.615
R23531 outputibias.n89 outputibias.n67 104.615
R23532 outputibias.n82 outputibias.n67 104.615
R23533 outputibias.n82 outputibias.n81 104.615
R23534 outputibias.n81 outputibias.n71 104.615
R23535 outputibias.n74 outputibias.n71 104.615
R23536 outputibias.n122 outputibias.n121 104.615
R23537 outputibias.n121 outputibias.n99 104.615
R23538 outputibias.n114 outputibias.n99 104.615
R23539 outputibias.n114 outputibias.n113 104.615
R23540 outputibias.n113 outputibias.n103 104.615
R23541 outputibias.n106 outputibias.n103 104.615
R23542 outputibias.n63 outputibias.n31 95.6354
R23543 outputibias.n63 outputibias.n62 94.6732
R23544 outputibias.n95 outputibias.n94 94.6732
R23545 outputibias.n127 outputibias.n126 94.6732
R23546 outputibias.n11 outputibias.t5 52.3082
R23547 outputibias.n42 outputibias.t7 52.3082
R23548 outputibias.n74 outputibias.t1 52.3082
R23549 outputibias.n106 outputibias.t3 52.3082
R23550 outputibias.n12 outputibias.n10 15.6674
R23551 outputibias.n43 outputibias.n41 15.6674
R23552 outputibias.n75 outputibias.n73 15.6674
R23553 outputibias.n107 outputibias.n105 15.6674
R23554 outputibias.n13 outputibias.n9 12.8005
R23555 outputibias.n44 outputibias.n40 12.8005
R23556 outputibias.n76 outputibias.n72 12.8005
R23557 outputibias.n108 outputibias.n104 12.8005
R23558 outputibias.n17 outputibias.n16 12.0247
R23559 outputibias.n48 outputibias.n47 12.0247
R23560 outputibias.n80 outputibias.n79 12.0247
R23561 outputibias.n112 outputibias.n111 12.0247
R23562 outputibias.n20 outputibias.n7 11.249
R23563 outputibias.n51 outputibias.n38 11.249
R23564 outputibias.n83 outputibias.n70 11.249
R23565 outputibias.n115 outputibias.n102 11.249
R23566 outputibias.n21 outputibias.n5 10.4732
R23567 outputibias.n52 outputibias.n36 10.4732
R23568 outputibias.n84 outputibias.n68 10.4732
R23569 outputibias.n116 outputibias.n100 10.4732
R23570 outputibias.n25 outputibias.n24 9.69747
R23571 outputibias.n56 outputibias.n55 9.69747
R23572 outputibias.n88 outputibias.n87 9.69747
R23573 outputibias.n120 outputibias.n119 9.69747
R23574 outputibias.n31 outputibias.n30 9.45567
R23575 outputibias.n62 outputibias.n61 9.45567
R23576 outputibias.n94 outputibias.n93 9.45567
R23577 outputibias.n126 outputibias.n125 9.45567
R23578 outputibias.n30 outputibias.n29 9.3005
R23579 outputibias.n3 outputibias.n2 9.3005
R23580 outputibias.n24 outputibias.n23 9.3005
R23581 outputibias.n22 outputibias.n21 9.3005
R23582 outputibias.n7 outputibias.n6 9.3005
R23583 outputibias.n16 outputibias.n15 9.3005
R23584 outputibias.n14 outputibias.n13 9.3005
R23585 outputibias.n61 outputibias.n60 9.3005
R23586 outputibias.n34 outputibias.n33 9.3005
R23587 outputibias.n55 outputibias.n54 9.3005
R23588 outputibias.n53 outputibias.n52 9.3005
R23589 outputibias.n38 outputibias.n37 9.3005
R23590 outputibias.n47 outputibias.n46 9.3005
R23591 outputibias.n45 outputibias.n44 9.3005
R23592 outputibias.n93 outputibias.n92 9.3005
R23593 outputibias.n66 outputibias.n65 9.3005
R23594 outputibias.n87 outputibias.n86 9.3005
R23595 outputibias.n85 outputibias.n84 9.3005
R23596 outputibias.n70 outputibias.n69 9.3005
R23597 outputibias.n79 outputibias.n78 9.3005
R23598 outputibias.n77 outputibias.n76 9.3005
R23599 outputibias.n125 outputibias.n124 9.3005
R23600 outputibias.n98 outputibias.n97 9.3005
R23601 outputibias.n119 outputibias.n118 9.3005
R23602 outputibias.n117 outputibias.n116 9.3005
R23603 outputibias.n102 outputibias.n101 9.3005
R23604 outputibias.n111 outputibias.n110 9.3005
R23605 outputibias.n109 outputibias.n108 9.3005
R23606 outputibias.n28 outputibias.n3 8.92171
R23607 outputibias.n59 outputibias.n34 8.92171
R23608 outputibias.n91 outputibias.n66 8.92171
R23609 outputibias.n123 outputibias.n98 8.92171
R23610 outputibias.n29 outputibias.n1 8.14595
R23611 outputibias.n60 outputibias.n32 8.14595
R23612 outputibias.n92 outputibias.n64 8.14595
R23613 outputibias.n124 outputibias.n96 8.14595
R23614 outputibias.n31 outputibias.n1 5.81868
R23615 outputibias.n62 outputibias.n32 5.81868
R23616 outputibias.n94 outputibias.n64 5.81868
R23617 outputibias.n126 outputibias.n96 5.81868
R23618 outputibias.n131 outputibias.n130 5.20947
R23619 outputibias.n29 outputibias.n28 5.04292
R23620 outputibias.n60 outputibias.n59 5.04292
R23621 outputibias.n92 outputibias.n91 5.04292
R23622 outputibias.n124 outputibias.n123 5.04292
R23623 outputibias.n131 outputibias.n127 4.42209
R23624 outputibias.n14 outputibias.n10 4.38594
R23625 outputibias.n45 outputibias.n41 4.38594
R23626 outputibias.n77 outputibias.n73 4.38594
R23627 outputibias.n109 outputibias.n105 4.38594
R23628 outputibias.n132 outputibias.n131 4.28454
R23629 outputibias.n25 outputibias.n3 4.26717
R23630 outputibias.n56 outputibias.n34 4.26717
R23631 outputibias.n88 outputibias.n66 4.26717
R23632 outputibias.n120 outputibias.n98 4.26717
R23633 outputibias.n24 outputibias.n5 3.49141
R23634 outputibias.n55 outputibias.n36 3.49141
R23635 outputibias.n87 outputibias.n68 3.49141
R23636 outputibias.n119 outputibias.n100 3.49141
R23637 outputibias.n21 outputibias.n20 2.71565
R23638 outputibias.n52 outputibias.n51 2.71565
R23639 outputibias.n84 outputibias.n83 2.71565
R23640 outputibias.n116 outputibias.n115 2.71565
R23641 outputibias.n17 outputibias.n7 1.93989
R23642 outputibias.n48 outputibias.n38 1.93989
R23643 outputibias.n80 outputibias.n70 1.93989
R23644 outputibias.n112 outputibias.n102 1.93989
R23645 outputibias.n130 outputibias.n129 1.9266
R23646 outputibias.n129 outputibias.n128 1.9266
R23647 outputibias.n133 outputibias.n132 1.92658
R23648 outputibias.n134 outputibias.n133 1.29913
R23649 outputibias.n16 outputibias.n9 1.16414
R23650 outputibias.n47 outputibias.n40 1.16414
R23651 outputibias.n79 outputibias.n72 1.16414
R23652 outputibias.n111 outputibias.n104 1.16414
R23653 outputibias.n127 outputibias.n95 0.962709
R23654 outputibias.n95 outputibias.n63 0.962709
R23655 outputibias.n13 outputibias.n12 0.388379
R23656 outputibias.n44 outputibias.n43 0.388379
R23657 outputibias.n76 outputibias.n75 0.388379
R23658 outputibias.n108 outputibias.n107 0.388379
R23659 outputibias.n134 outputibias.n0 0.337251
R23660 outputibias outputibias.n134 0.302375
R23661 outputibias.n30 outputibias.n2 0.155672
R23662 outputibias.n23 outputibias.n2 0.155672
R23663 outputibias.n23 outputibias.n22 0.155672
R23664 outputibias.n22 outputibias.n6 0.155672
R23665 outputibias.n15 outputibias.n6 0.155672
R23666 outputibias.n15 outputibias.n14 0.155672
R23667 outputibias.n61 outputibias.n33 0.155672
R23668 outputibias.n54 outputibias.n33 0.155672
R23669 outputibias.n54 outputibias.n53 0.155672
R23670 outputibias.n53 outputibias.n37 0.155672
R23671 outputibias.n46 outputibias.n37 0.155672
R23672 outputibias.n46 outputibias.n45 0.155672
R23673 outputibias.n93 outputibias.n65 0.155672
R23674 outputibias.n86 outputibias.n65 0.155672
R23675 outputibias.n86 outputibias.n85 0.155672
R23676 outputibias.n85 outputibias.n69 0.155672
R23677 outputibias.n78 outputibias.n69 0.155672
R23678 outputibias.n78 outputibias.n77 0.155672
R23679 outputibias.n125 outputibias.n97 0.155672
R23680 outputibias.n118 outputibias.n97 0.155672
R23681 outputibias.n118 outputibias.n117 0.155672
R23682 outputibias.n117 outputibias.n101 0.155672
R23683 outputibias.n110 outputibias.n101 0.155672
R23684 outputibias.n110 outputibias.n109 0.155672
R23685 output.n41 output.n15 289.615
R23686 output.n72 output.n46 289.615
R23687 output.n104 output.n78 289.615
R23688 output.n136 output.n110 289.615
R23689 output.n77 output.n45 197.26
R23690 output.n77 output.n76 196.298
R23691 output.n109 output.n108 196.298
R23692 output.n141 output.n140 196.298
R23693 output.n42 output.n41 185
R23694 output.n40 output.n39 185
R23695 output.n19 output.n18 185
R23696 output.n34 output.n33 185
R23697 output.n32 output.n31 185
R23698 output.n23 output.n22 185
R23699 output.n26 output.n25 185
R23700 output.n73 output.n72 185
R23701 output.n71 output.n70 185
R23702 output.n50 output.n49 185
R23703 output.n65 output.n64 185
R23704 output.n63 output.n62 185
R23705 output.n54 output.n53 185
R23706 output.n57 output.n56 185
R23707 output.n105 output.n104 185
R23708 output.n103 output.n102 185
R23709 output.n82 output.n81 185
R23710 output.n97 output.n96 185
R23711 output.n95 output.n94 185
R23712 output.n86 output.n85 185
R23713 output.n89 output.n88 185
R23714 output.n137 output.n136 185
R23715 output.n135 output.n134 185
R23716 output.n114 output.n113 185
R23717 output.n129 output.n128 185
R23718 output.n127 output.n126 185
R23719 output.n118 output.n117 185
R23720 output.n121 output.n120 185
R23721 output.t2 output.n24 147.661
R23722 output.t1 output.n55 147.661
R23723 output.t3 output.n87 147.661
R23724 output.t0 output.n119 147.661
R23725 output.n41 output.n40 104.615
R23726 output.n40 output.n18 104.615
R23727 output.n33 output.n18 104.615
R23728 output.n33 output.n32 104.615
R23729 output.n32 output.n22 104.615
R23730 output.n25 output.n22 104.615
R23731 output.n72 output.n71 104.615
R23732 output.n71 output.n49 104.615
R23733 output.n64 output.n49 104.615
R23734 output.n64 output.n63 104.615
R23735 output.n63 output.n53 104.615
R23736 output.n56 output.n53 104.615
R23737 output.n104 output.n103 104.615
R23738 output.n103 output.n81 104.615
R23739 output.n96 output.n81 104.615
R23740 output.n96 output.n95 104.615
R23741 output.n95 output.n85 104.615
R23742 output.n88 output.n85 104.615
R23743 output.n136 output.n135 104.615
R23744 output.n135 output.n113 104.615
R23745 output.n128 output.n113 104.615
R23746 output.n128 output.n127 104.615
R23747 output.n127 output.n117 104.615
R23748 output.n120 output.n117 104.615
R23749 output.n1 output.t8 77.056
R23750 output.n14 output.t9 76.6694
R23751 output.n1 output.n0 72.7095
R23752 output.n3 output.n2 72.7095
R23753 output.n5 output.n4 72.7095
R23754 output.n7 output.n6 72.7095
R23755 output.n9 output.n8 72.7095
R23756 output.n11 output.n10 72.7095
R23757 output.n13 output.n12 72.7095
R23758 output.n25 output.t2 52.3082
R23759 output.n56 output.t1 52.3082
R23760 output.n88 output.t3 52.3082
R23761 output.n120 output.t0 52.3082
R23762 output.n26 output.n24 15.6674
R23763 output.n57 output.n55 15.6674
R23764 output.n89 output.n87 15.6674
R23765 output.n121 output.n119 15.6674
R23766 output.n27 output.n23 12.8005
R23767 output.n58 output.n54 12.8005
R23768 output.n90 output.n86 12.8005
R23769 output.n122 output.n118 12.8005
R23770 output.n31 output.n30 12.0247
R23771 output.n62 output.n61 12.0247
R23772 output.n94 output.n93 12.0247
R23773 output.n126 output.n125 12.0247
R23774 output.n34 output.n21 11.249
R23775 output.n65 output.n52 11.249
R23776 output.n97 output.n84 11.249
R23777 output.n129 output.n116 11.249
R23778 output.n35 output.n19 10.4732
R23779 output.n66 output.n50 10.4732
R23780 output.n98 output.n82 10.4732
R23781 output.n130 output.n114 10.4732
R23782 output.n39 output.n38 9.69747
R23783 output.n70 output.n69 9.69747
R23784 output.n102 output.n101 9.69747
R23785 output.n134 output.n133 9.69747
R23786 output.n45 output.n44 9.45567
R23787 output.n76 output.n75 9.45567
R23788 output.n108 output.n107 9.45567
R23789 output.n140 output.n139 9.45567
R23790 output.n44 output.n43 9.3005
R23791 output.n17 output.n16 9.3005
R23792 output.n38 output.n37 9.3005
R23793 output.n36 output.n35 9.3005
R23794 output.n21 output.n20 9.3005
R23795 output.n30 output.n29 9.3005
R23796 output.n28 output.n27 9.3005
R23797 output.n75 output.n74 9.3005
R23798 output.n48 output.n47 9.3005
R23799 output.n69 output.n68 9.3005
R23800 output.n67 output.n66 9.3005
R23801 output.n52 output.n51 9.3005
R23802 output.n61 output.n60 9.3005
R23803 output.n59 output.n58 9.3005
R23804 output.n107 output.n106 9.3005
R23805 output.n80 output.n79 9.3005
R23806 output.n101 output.n100 9.3005
R23807 output.n99 output.n98 9.3005
R23808 output.n84 output.n83 9.3005
R23809 output.n93 output.n92 9.3005
R23810 output.n91 output.n90 9.3005
R23811 output.n139 output.n138 9.3005
R23812 output.n112 output.n111 9.3005
R23813 output.n133 output.n132 9.3005
R23814 output.n131 output.n130 9.3005
R23815 output.n116 output.n115 9.3005
R23816 output.n125 output.n124 9.3005
R23817 output.n123 output.n122 9.3005
R23818 output.n42 output.n17 8.92171
R23819 output.n73 output.n48 8.92171
R23820 output.n105 output.n80 8.92171
R23821 output.n137 output.n112 8.92171
R23822 output output.n141 8.15037
R23823 output.n43 output.n15 8.14595
R23824 output.n74 output.n46 8.14595
R23825 output.n106 output.n78 8.14595
R23826 output.n138 output.n110 8.14595
R23827 output.n45 output.n15 5.81868
R23828 output.n76 output.n46 5.81868
R23829 output.n108 output.n78 5.81868
R23830 output.n140 output.n110 5.81868
R23831 output.n43 output.n42 5.04292
R23832 output.n74 output.n73 5.04292
R23833 output.n106 output.n105 5.04292
R23834 output.n138 output.n137 5.04292
R23835 output.n28 output.n24 4.38594
R23836 output.n59 output.n55 4.38594
R23837 output.n91 output.n87 4.38594
R23838 output.n123 output.n119 4.38594
R23839 output.n39 output.n17 4.26717
R23840 output.n70 output.n48 4.26717
R23841 output.n102 output.n80 4.26717
R23842 output.n134 output.n112 4.26717
R23843 output.n0 output.t14 3.9605
R23844 output.n0 output.t18 3.9605
R23845 output.n2 output.t5 3.9605
R23846 output.n2 output.t10 3.9605
R23847 output.n4 output.t11 3.9605
R23848 output.n4 output.t16 3.9605
R23849 output.n6 output.t4 3.9605
R23850 output.n6 output.t12 3.9605
R23851 output.n8 output.t15 3.9605
R23852 output.n8 output.t13 3.9605
R23853 output.n10 output.t19 3.9605
R23854 output.n10 output.t6 3.9605
R23855 output.n12 output.t7 3.9605
R23856 output.n12 output.t17 3.9605
R23857 output.n38 output.n19 3.49141
R23858 output.n69 output.n50 3.49141
R23859 output.n101 output.n82 3.49141
R23860 output.n133 output.n114 3.49141
R23861 output.n35 output.n34 2.71565
R23862 output.n66 output.n65 2.71565
R23863 output.n98 output.n97 2.71565
R23864 output.n130 output.n129 2.71565
R23865 output.n31 output.n21 1.93989
R23866 output.n62 output.n52 1.93989
R23867 output.n94 output.n84 1.93989
R23868 output.n126 output.n116 1.93989
R23869 output.n30 output.n23 1.16414
R23870 output.n61 output.n54 1.16414
R23871 output.n93 output.n86 1.16414
R23872 output.n125 output.n118 1.16414
R23873 output.n141 output.n109 0.962709
R23874 output.n109 output.n77 0.962709
R23875 output.n27 output.n26 0.388379
R23876 output.n58 output.n57 0.388379
R23877 output.n90 output.n89 0.388379
R23878 output.n122 output.n121 0.388379
R23879 output.n14 output.n13 0.387128
R23880 output.n13 output.n11 0.387128
R23881 output.n11 output.n9 0.387128
R23882 output.n9 output.n7 0.387128
R23883 output.n7 output.n5 0.387128
R23884 output.n5 output.n3 0.387128
R23885 output.n3 output.n1 0.387128
R23886 output.n44 output.n16 0.155672
R23887 output.n37 output.n16 0.155672
R23888 output.n37 output.n36 0.155672
R23889 output.n36 output.n20 0.155672
R23890 output.n29 output.n20 0.155672
R23891 output.n29 output.n28 0.155672
R23892 output.n75 output.n47 0.155672
R23893 output.n68 output.n47 0.155672
R23894 output.n68 output.n67 0.155672
R23895 output.n67 output.n51 0.155672
R23896 output.n60 output.n51 0.155672
R23897 output.n60 output.n59 0.155672
R23898 output.n107 output.n79 0.155672
R23899 output.n100 output.n79 0.155672
R23900 output.n100 output.n99 0.155672
R23901 output.n99 output.n83 0.155672
R23902 output.n92 output.n83 0.155672
R23903 output.n92 output.n91 0.155672
R23904 output.n139 output.n111 0.155672
R23905 output.n132 output.n111 0.155672
R23906 output.n132 output.n131 0.155672
R23907 output.n131 output.n115 0.155672
R23908 output.n124 output.n115 0.155672
R23909 output.n124 output.n123 0.155672
R23910 output output.n14 0.126227
C0 commonsourceibias output 0.006808f
C1 minus diffpairibias 5.39e-19
C2 CSoutput minus 2.76559f
C3 vdd plus 0.088406f
C4 plus diffpairibias 4.4e-19
C5 commonsourceibias outputibias 0.003832f
C6 vdd commonsourceibias 0.004218f
C7 CSoutput plus 0.912122f
C8 commonsourceibias diffpairibias 0.064336f
C9 CSoutput commonsourceibias 54.554f
C10 minus plus 10.3849f
C11 minus commonsourceibias 0.343793f
C12 plus commonsourceibias 0.290384f
C13 output outputibias 2.34152f
C14 vdd output 7.23429f
C15 CSoutput output 6.13881f
C16 CSoutput outputibias 0.032386f
C17 vdd CSoutput 0.116319p
C18 diffpairibias gnd 60.003128f
C19 outputibias gnd 32.465668f
C20 output gnd 15.47879f
C21 commonsourceibias gnd 0.184128p
C22 plus gnd 39.4907f
C23 minus gnd 31.358328f
C24 CSoutput gnd 0.126433p
C25 vdd gnd 0.407906p
C26 output.t8 gnd 0.464308f
C27 output.t14 gnd 0.044422f
C28 output.t18 gnd 0.044422f
C29 output.n0 gnd 0.364624f
C30 output.n1 gnd 0.614102f
C31 output.t5 gnd 0.044422f
C32 output.t10 gnd 0.044422f
C33 output.n2 gnd 0.364624f
C34 output.n3 gnd 0.350265f
C35 output.t11 gnd 0.044422f
C36 output.t16 gnd 0.044422f
C37 output.n4 gnd 0.364624f
C38 output.n5 gnd 0.350265f
C39 output.t4 gnd 0.044422f
C40 output.t12 gnd 0.044422f
C41 output.n6 gnd 0.364624f
C42 output.n7 gnd 0.350265f
C43 output.t15 gnd 0.044422f
C44 output.t13 gnd 0.044422f
C45 output.n8 gnd 0.364624f
C46 output.n9 gnd 0.350265f
C47 output.t19 gnd 0.044422f
C48 output.t6 gnd 0.044422f
C49 output.n10 gnd 0.364624f
C50 output.n11 gnd 0.350265f
C51 output.t7 gnd 0.044422f
C52 output.t17 gnd 0.044422f
C53 output.n12 gnd 0.364624f
C54 output.n13 gnd 0.350265f
C55 output.t9 gnd 0.462979f
C56 output.n14 gnd 0.28994f
C57 output.n15 gnd 0.015803f
C58 output.n16 gnd 0.011243f
C59 output.n17 gnd 0.006041f
C60 output.n18 gnd 0.01428f
C61 output.n19 gnd 0.006397f
C62 output.n20 gnd 0.011243f
C63 output.n21 gnd 0.006041f
C64 output.n22 gnd 0.01428f
C65 output.n23 gnd 0.006397f
C66 output.n24 gnd 0.048111f
C67 output.t2 gnd 0.023274f
C68 output.n25 gnd 0.01071f
C69 output.n26 gnd 0.008435f
C70 output.n27 gnd 0.006041f
C71 output.n28 gnd 0.267512f
C72 output.n29 gnd 0.011243f
C73 output.n30 gnd 0.006041f
C74 output.n31 gnd 0.006397f
C75 output.n32 gnd 0.01428f
C76 output.n33 gnd 0.01428f
C77 output.n34 gnd 0.006397f
C78 output.n35 gnd 0.006041f
C79 output.n36 gnd 0.011243f
C80 output.n37 gnd 0.011243f
C81 output.n38 gnd 0.006041f
C82 output.n39 gnd 0.006397f
C83 output.n40 gnd 0.01428f
C84 output.n41 gnd 0.030913f
C85 output.n42 gnd 0.006397f
C86 output.n43 gnd 0.006041f
C87 output.n44 gnd 0.025987f
C88 output.n45 gnd 0.097665f
C89 output.n46 gnd 0.015803f
C90 output.n47 gnd 0.011243f
C91 output.n48 gnd 0.006041f
C92 output.n49 gnd 0.01428f
C93 output.n50 gnd 0.006397f
C94 output.n51 gnd 0.011243f
C95 output.n52 gnd 0.006041f
C96 output.n53 gnd 0.01428f
C97 output.n54 gnd 0.006397f
C98 output.n55 gnd 0.048111f
C99 output.t1 gnd 0.023274f
C100 output.n56 gnd 0.01071f
C101 output.n57 gnd 0.008435f
C102 output.n58 gnd 0.006041f
C103 output.n59 gnd 0.267512f
C104 output.n60 gnd 0.011243f
C105 output.n61 gnd 0.006041f
C106 output.n62 gnd 0.006397f
C107 output.n63 gnd 0.01428f
C108 output.n64 gnd 0.01428f
C109 output.n65 gnd 0.006397f
C110 output.n66 gnd 0.006041f
C111 output.n67 gnd 0.011243f
C112 output.n68 gnd 0.011243f
C113 output.n69 gnd 0.006041f
C114 output.n70 gnd 0.006397f
C115 output.n71 gnd 0.01428f
C116 output.n72 gnd 0.030913f
C117 output.n73 gnd 0.006397f
C118 output.n74 gnd 0.006041f
C119 output.n75 gnd 0.025987f
C120 output.n76 gnd 0.09306f
C121 output.n77 gnd 1.65264f
C122 output.n78 gnd 0.015803f
C123 output.n79 gnd 0.011243f
C124 output.n80 gnd 0.006041f
C125 output.n81 gnd 0.01428f
C126 output.n82 gnd 0.006397f
C127 output.n83 gnd 0.011243f
C128 output.n84 gnd 0.006041f
C129 output.n85 gnd 0.01428f
C130 output.n86 gnd 0.006397f
C131 output.n87 gnd 0.048111f
C132 output.t3 gnd 0.023274f
C133 output.n88 gnd 0.01071f
C134 output.n89 gnd 0.008435f
C135 output.n90 gnd 0.006041f
C136 output.n91 gnd 0.267512f
C137 output.n92 gnd 0.011243f
C138 output.n93 gnd 0.006041f
C139 output.n94 gnd 0.006397f
C140 output.n95 gnd 0.01428f
C141 output.n96 gnd 0.01428f
C142 output.n97 gnd 0.006397f
C143 output.n98 gnd 0.006041f
C144 output.n99 gnd 0.011243f
C145 output.n100 gnd 0.011243f
C146 output.n101 gnd 0.006041f
C147 output.n102 gnd 0.006397f
C148 output.n103 gnd 0.01428f
C149 output.n104 gnd 0.030913f
C150 output.n105 gnd 0.006397f
C151 output.n106 gnd 0.006041f
C152 output.n107 gnd 0.025987f
C153 output.n108 gnd 0.09306f
C154 output.n109 gnd 0.713089f
C155 output.n110 gnd 0.015803f
C156 output.n111 gnd 0.011243f
C157 output.n112 gnd 0.006041f
C158 output.n113 gnd 0.01428f
C159 output.n114 gnd 0.006397f
C160 output.n115 gnd 0.011243f
C161 output.n116 gnd 0.006041f
C162 output.n117 gnd 0.01428f
C163 output.n118 gnd 0.006397f
C164 output.n119 gnd 0.048111f
C165 output.t0 gnd 0.023274f
C166 output.n120 gnd 0.01071f
C167 output.n121 gnd 0.008435f
C168 output.n122 gnd 0.006041f
C169 output.n123 gnd 0.267512f
C170 output.n124 gnd 0.011243f
C171 output.n125 gnd 0.006041f
C172 output.n126 gnd 0.006397f
C173 output.n127 gnd 0.01428f
C174 output.n128 gnd 0.01428f
C175 output.n129 gnd 0.006397f
C176 output.n130 gnd 0.006041f
C177 output.n131 gnd 0.011243f
C178 output.n132 gnd 0.011243f
C179 output.n133 gnd 0.006041f
C180 output.n134 gnd 0.006397f
C181 output.n135 gnd 0.01428f
C182 output.n136 gnd 0.030913f
C183 output.n137 gnd 0.006397f
C184 output.n138 gnd 0.006041f
C185 output.n139 gnd 0.025987f
C186 output.n140 gnd 0.09306f
C187 output.n141 gnd 1.67353f
C188 outputibias.t10 gnd 0.11477f
C189 outputibias.t9 gnd 0.115567f
C190 outputibias.n0 gnd 0.130108f
C191 outputibias.n1 gnd 0.001372f
C192 outputibias.n2 gnd 9.76e-19
C193 outputibias.n3 gnd 5.24e-19
C194 outputibias.n4 gnd 0.001239f
C195 outputibias.n5 gnd 5.55e-19
C196 outputibias.n6 gnd 9.76e-19
C197 outputibias.n7 gnd 5.24e-19
C198 outputibias.n8 gnd 0.001239f
C199 outputibias.n9 gnd 5.55e-19
C200 outputibias.n10 gnd 0.004176f
C201 outputibias.t5 gnd 0.00202f
C202 outputibias.n11 gnd 9.3e-19
C203 outputibias.n12 gnd 7.32e-19
C204 outputibias.n13 gnd 5.24e-19
C205 outputibias.n14 gnd 0.02322f
C206 outputibias.n15 gnd 9.76e-19
C207 outputibias.n16 gnd 5.24e-19
C208 outputibias.n17 gnd 5.55e-19
C209 outputibias.n18 gnd 0.001239f
C210 outputibias.n19 gnd 0.001239f
C211 outputibias.n20 gnd 5.55e-19
C212 outputibias.n21 gnd 5.24e-19
C213 outputibias.n22 gnd 9.76e-19
C214 outputibias.n23 gnd 9.76e-19
C215 outputibias.n24 gnd 5.24e-19
C216 outputibias.n25 gnd 5.55e-19
C217 outputibias.n26 gnd 0.001239f
C218 outputibias.n27 gnd 0.002683f
C219 outputibias.n28 gnd 5.55e-19
C220 outputibias.n29 gnd 5.24e-19
C221 outputibias.n30 gnd 0.002256f
C222 outputibias.n31 gnd 0.005781f
C223 outputibias.n32 gnd 0.001372f
C224 outputibias.n33 gnd 9.76e-19
C225 outputibias.n34 gnd 5.24e-19
C226 outputibias.n35 gnd 0.001239f
C227 outputibias.n36 gnd 5.55e-19
C228 outputibias.n37 gnd 9.76e-19
C229 outputibias.n38 gnd 5.24e-19
C230 outputibias.n39 gnd 0.001239f
C231 outputibias.n40 gnd 5.55e-19
C232 outputibias.n41 gnd 0.004176f
C233 outputibias.t7 gnd 0.00202f
C234 outputibias.n42 gnd 9.3e-19
C235 outputibias.n43 gnd 7.32e-19
C236 outputibias.n44 gnd 5.24e-19
C237 outputibias.n45 gnd 0.02322f
C238 outputibias.n46 gnd 9.76e-19
C239 outputibias.n47 gnd 5.24e-19
C240 outputibias.n48 gnd 5.55e-19
C241 outputibias.n49 gnd 0.001239f
C242 outputibias.n50 gnd 0.001239f
C243 outputibias.n51 gnd 5.55e-19
C244 outputibias.n52 gnd 5.24e-19
C245 outputibias.n53 gnd 9.76e-19
C246 outputibias.n54 gnd 9.76e-19
C247 outputibias.n55 gnd 5.24e-19
C248 outputibias.n56 gnd 5.55e-19
C249 outputibias.n57 gnd 0.001239f
C250 outputibias.n58 gnd 0.002683f
C251 outputibias.n59 gnd 5.55e-19
C252 outputibias.n60 gnd 5.24e-19
C253 outputibias.n61 gnd 0.002256f
C254 outputibias.n62 gnd 0.005197f
C255 outputibias.n63 gnd 0.121892f
C256 outputibias.n64 gnd 0.001372f
C257 outputibias.n65 gnd 9.76e-19
C258 outputibias.n66 gnd 5.24e-19
C259 outputibias.n67 gnd 0.001239f
C260 outputibias.n68 gnd 5.55e-19
C261 outputibias.n69 gnd 9.76e-19
C262 outputibias.n70 gnd 5.24e-19
C263 outputibias.n71 gnd 0.001239f
C264 outputibias.n72 gnd 5.55e-19
C265 outputibias.n73 gnd 0.004176f
C266 outputibias.t1 gnd 0.00202f
C267 outputibias.n74 gnd 9.3e-19
C268 outputibias.n75 gnd 7.32e-19
C269 outputibias.n76 gnd 5.24e-19
C270 outputibias.n77 gnd 0.02322f
C271 outputibias.n78 gnd 9.76e-19
C272 outputibias.n79 gnd 5.24e-19
C273 outputibias.n80 gnd 5.55e-19
C274 outputibias.n81 gnd 0.001239f
C275 outputibias.n82 gnd 0.001239f
C276 outputibias.n83 gnd 5.55e-19
C277 outputibias.n84 gnd 5.24e-19
C278 outputibias.n85 gnd 9.76e-19
C279 outputibias.n86 gnd 9.76e-19
C280 outputibias.n87 gnd 5.24e-19
C281 outputibias.n88 gnd 5.55e-19
C282 outputibias.n89 gnd 0.001239f
C283 outputibias.n90 gnd 0.002683f
C284 outputibias.n91 gnd 5.55e-19
C285 outputibias.n92 gnd 5.24e-19
C286 outputibias.n93 gnd 0.002256f
C287 outputibias.n94 gnd 0.005197f
C288 outputibias.n95 gnd 0.064513f
C289 outputibias.n96 gnd 0.001372f
C290 outputibias.n97 gnd 9.76e-19
C291 outputibias.n98 gnd 5.24e-19
C292 outputibias.n99 gnd 0.001239f
C293 outputibias.n100 gnd 5.55e-19
C294 outputibias.n101 gnd 9.76e-19
C295 outputibias.n102 gnd 5.24e-19
C296 outputibias.n103 gnd 0.001239f
C297 outputibias.n104 gnd 5.55e-19
C298 outputibias.n105 gnd 0.004176f
C299 outputibias.t3 gnd 0.00202f
C300 outputibias.n106 gnd 9.3e-19
C301 outputibias.n107 gnd 7.32e-19
C302 outputibias.n108 gnd 5.24e-19
C303 outputibias.n109 gnd 0.02322f
C304 outputibias.n110 gnd 9.76e-19
C305 outputibias.n111 gnd 5.24e-19
C306 outputibias.n112 gnd 5.55e-19
C307 outputibias.n113 gnd 0.001239f
C308 outputibias.n114 gnd 0.001239f
C309 outputibias.n115 gnd 5.55e-19
C310 outputibias.n116 gnd 5.24e-19
C311 outputibias.n117 gnd 9.76e-19
C312 outputibias.n118 gnd 9.76e-19
C313 outputibias.n119 gnd 5.24e-19
C314 outputibias.n120 gnd 5.55e-19
C315 outputibias.n121 gnd 0.001239f
C316 outputibias.n122 gnd 0.002683f
C317 outputibias.n123 gnd 5.55e-19
C318 outputibias.n124 gnd 5.24e-19
C319 outputibias.n125 gnd 0.002256f
C320 outputibias.n126 gnd 0.005197f
C321 outputibias.n127 gnd 0.084814f
C322 outputibias.t2 gnd 0.108319f
C323 outputibias.t0 gnd 0.108319f
C324 outputibias.t6 gnd 0.108319f
C325 outputibias.t4 gnd 0.109238f
C326 outputibias.n128 gnd 0.134674f
C327 outputibias.n129 gnd 0.07244f
C328 outputibias.n130 gnd 0.079818f
C329 outputibias.n131 gnd 0.164901f
C330 outputibias.t11 gnd 0.11477f
C331 outputibias.n132 gnd 0.067481f
C332 outputibias.t8 gnd 0.11477f
C333 outputibias.n133 gnd 0.065115f
C334 outputibias.n134 gnd 0.029159f
C335 minus.n0 gnd 0.030802f
C336 minus.t13 gnd 0.517928f
C337 minus.n1 gnd 0.209473f
C338 minus.n2 gnd 0.030802f
C339 minus.t11 gnd 0.517928f
C340 minus.n3 gnd 0.026321f
C341 minus.n4 gnd 0.030802f
C342 minus.t17 gnd 0.517928f
C343 minus.t24 gnd 0.517928f
C344 minus.n5 gnd 0.209473f
C345 minus.n6 gnd 0.030802f
C346 minus.t21 gnd 0.517928f
C347 minus.n7 gnd 0.209473f
C348 minus.n8 gnd 0.030802f
C349 minus.t27 gnd 0.517928f
C350 minus.n9 gnd 0.025035f
C351 minus.n10 gnd 0.030802f
C352 minus.t26 gnd 0.517928f
C353 minus.t5 gnd 0.517928f
C354 minus.n11 gnd 0.209473f
C355 minus.n12 gnd 0.030802f
C356 minus.t9 gnd 0.517928f
C357 minus.n13 gnd 0.209473f
C358 minus.n14 gnd 0.13072f
C359 minus.t14 gnd 0.517928f
C360 minus.t20 gnd 0.579396f
C361 minus.n15 gnd 0.244895f
C362 minus.n16 gnd 0.239886f
C363 minus.n17 gnd 0.039468f
C364 minus.n18 gnd 0.034856f
C365 minus.n19 gnd 0.030802f
C366 minus.n20 gnd 0.030802f
C367 minus.n21 gnd 0.036808f
C368 minus.n22 gnd 0.026321f
C369 minus.n23 gnd 0.040115f
C370 minus.n24 gnd 0.030802f
C371 minus.n25 gnd 0.030802f
C372 minus.n26 gnd 0.038315f
C373 minus.n27 gnd 0.036009f
C374 minus.n28 gnd 0.209473f
C375 minus.n29 gnd 0.038584f
C376 minus.n30 gnd 0.030802f
C377 minus.n31 gnd 0.030802f
C378 minus.n32 gnd 0.030802f
C379 minus.n33 gnd 0.039625f
C380 minus.n34 gnd 0.209473f
C381 minus.n35 gnd 0.037162f
C382 minus.n36 gnd 0.037162f
C383 minus.n37 gnd 0.030802f
C384 minus.n38 gnd 0.030802f
C385 minus.n39 gnd 0.039625f
C386 minus.n40 gnd 0.025035f
C387 minus.n41 gnd 0.038584f
C388 minus.n42 gnd 0.030802f
C389 minus.n43 gnd 0.030802f
C390 minus.n44 gnd 0.036009f
C391 minus.n45 gnd 0.038315f
C392 minus.n46 gnd 0.209473f
C393 minus.n47 gnd 0.040115f
C394 minus.n48 gnd 0.030802f
C395 minus.n49 gnd 0.030802f
C396 minus.n50 gnd 0.030802f
C397 minus.n51 gnd 0.036808f
C398 minus.n52 gnd 0.209473f
C399 minus.n53 gnd 0.034856f
C400 minus.n54 gnd 0.039468f
C401 minus.n55 gnd 0.030802f
C402 minus.n56 gnd 0.030802f
C403 minus.n57 gnd 0.040182f
C404 minus.n58 gnd 0.011194f
C405 minus.t10 gnd 0.560139f
C406 minus.n59 gnd 0.242535f
C407 minus.n60 gnd 0.360831f
C408 minus.n61 gnd 0.030802f
C409 minus.t8 gnd 0.560139f
C410 minus.t12 gnd 0.517928f
C411 minus.n62 gnd 0.209473f
C412 minus.n63 gnd 0.030802f
C413 minus.t18 gnd 0.517928f
C414 minus.n64 gnd 0.026321f
C415 minus.n65 gnd 0.030802f
C416 minus.t25 gnd 0.517928f
C417 minus.t22 gnd 0.517928f
C418 minus.n66 gnd 0.209473f
C419 minus.n67 gnd 0.030802f
C420 minus.t19 gnd 0.517928f
C421 minus.n68 gnd 0.209473f
C422 minus.n69 gnd 0.030802f
C423 minus.t7 gnd 0.517928f
C424 minus.n70 gnd 0.025035f
C425 minus.n71 gnd 0.030802f
C426 minus.t6 gnd 0.517928f
C427 minus.t16 gnd 0.517928f
C428 minus.n72 gnd 0.209473f
C429 minus.n73 gnd 0.030802f
C430 minus.t15 gnd 0.517928f
C431 minus.n74 gnd 0.209473f
C432 minus.n75 gnd 0.13072f
C433 minus.t23 gnd 0.517928f
C434 minus.t28 gnd 0.579396f
C435 minus.n76 gnd 0.244895f
C436 minus.n77 gnd 0.239886f
C437 minus.n78 gnd 0.039468f
C438 minus.n79 gnd 0.034856f
C439 minus.n80 gnd 0.030802f
C440 minus.n81 gnd 0.030802f
C441 minus.n82 gnd 0.036808f
C442 minus.n83 gnd 0.026321f
C443 minus.n84 gnd 0.040115f
C444 minus.n85 gnd 0.030802f
C445 minus.n86 gnd 0.030802f
C446 minus.n87 gnd 0.038315f
C447 minus.n88 gnd 0.036009f
C448 minus.n89 gnd 0.209473f
C449 minus.n90 gnd 0.038584f
C450 minus.n91 gnd 0.030802f
C451 minus.n92 gnd 0.030802f
C452 minus.n93 gnd 0.030802f
C453 minus.n94 gnd 0.039625f
C454 minus.n95 gnd 0.209473f
C455 minus.n96 gnd 0.037162f
C456 minus.n97 gnd 0.037162f
C457 minus.n98 gnd 0.030802f
C458 minus.n99 gnd 0.030802f
C459 minus.n100 gnd 0.039625f
C460 minus.n101 gnd 0.025035f
C461 minus.n102 gnd 0.038584f
C462 minus.n103 gnd 0.030802f
C463 minus.n104 gnd 0.030802f
C464 minus.n105 gnd 0.036009f
C465 minus.n106 gnd 0.038315f
C466 minus.n107 gnd 0.209473f
C467 minus.n108 gnd 0.040115f
C468 minus.n109 gnd 0.030802f
C469 minus.n110 gnd 0.030802f
C470 minus.n111 gnd 0.030802f
C471 minus.n112 gnd 0.036808f
C472 minus.n113 gnd 0.209473f
C473 minus.n114 gnd 0.034856f
C474 minus.n115 gnd 0.039468f
C475 minus.n116 gnd 0.030802f
C476 minus.n117 gnd 0.030802f
C477 minus.n118 gnd 0.040182f
C478 minus.n119 gnd 0.011194f
C479 minus.n120 gnd 0.242535f
C480 minus.n121 gnd 1.12364f
C481 minus.n122 gnd 1.65054f
C482 minus.t4 gnd 0.009495f
C483 minus.t3 gnd 0.009495f
C484 minus.n123 gnd 0.031223f
C485 minus.t0 gnd 0.009495f
C486 minus.t2 gnd 0.009495f
C487 minus.n124 gnd 0.030795f
C488 minus.n125 gnd 0.262821f
C489 minus.t1 gnd 0.05285f
C490 minus.n126 gnd 0.143419f
C491 minus.n127 gnd 1.93361f
C492 a_n1986_8322.t21 gnd 49.3316f
C493 a_n1986_8322.t20 gnd 76.0671f
C494 a_n1986_8322.t2 gnd 0.093483f
C495 a_n1986_8322.t1 gnd 0.875324f
C496 a_n1986_8322.t9 gnd 0.093483f
C497 a_n1986_8322.t4 gnd 0.093483f
C498 a_n1986_8322.n0 gnd 0.658492f
C499 a_n1986_8322.n1 gnd 0.735768f
C500 a_n1986_8322.t7 gnd 0.093483f
C501 a_n1986_8322.t6 gnd 0.093483f
C502 a_n1986_8322.n2 gnd 0.658492f
C503 a_n1986_8322.n3 gnd 0.373834f
C504 a_n1986_8322.t0 gnd 0.873581f
C505 a_n1986_8322.n4 gnd 1.39821f
C506 a_n1986_8322.t15 gnd 0.875324f
C507 a_n1986_8322.t19 gnd 0.093483f
C508 a_n1986_8322.t18 gnd 0.093483f
C509 a_n1986_8322.n5 gnd 0.658492f
C510 a_n1986_8322.n6 gnd 0.735768f
C511 a_n1986_8322.t13 gnd 0.873581f
C512 a_n1986_8322.n7 gnd 0.370248f
C513 a_n1986_8322.t16 gnd 0.873581f
C514 a_n1986_8322.n8 gnd 0.370248f
C515 a_n1986_8322.t14 gnd 0.093483f
C516 a_n1986_8322.t12 gnd 0.093483f
C517 a_n1986_8322.n9 gnd 0.658492f
C518 a_n1986_8322.n10 gnd 0.373834f
C519 a_n1986_8322.t17 gnd 0.873581f
C520 a_n1986_8322.n11 gnd 0.871851f
C521 a_n1986_8322.n12 gnd 1.58986f
C522 a_n1986_8322.n13 gnd 3.73938f
C523 a_n1986_8322.t3 gnd 0.873581f
C524 a_n1986_8322.n14 gnd 0.766111f
C525 a_n1986_8322.t10 gnd 0.875322f
C526 a_n1986_8322.t8 gnd 0.093483f
C527 a_n1986_8322.t5 gnd 0.093483f
C528 a_n1986_8322.n15 gnd 0.658492f
C529 a_n1986_8322.n16 gnd 0.73577f
C530 a_n1986_8322.n17 gnd 0.373832f
C531 a_n1986_8322.n18 gnd 0.658494f
C532 a_n1986_8322.t11 gnd 0.093483f
C533 diffpairibias.t27 gnd 0.090128f
C534 diffpairibias.t23 gnd 0.08996f
C535 diffpairibias.n0 gnd 0.105991f
C536 diffpairibias.t28 gnd 0.08996f
C537 diffpairibias.n1 gnd 0.051736f
C538 diffpairibias.t25 gnd 0.08996f
C539 diffpairibias.n2 gnd 0.051736f
C540 diffpairibias.t29 gnd 0.08996f
C541 diffpairibias.n3 gnd 0.041084f
C542 diffpairibias.t15 gnd 0.086371f
C543 diffpairibias.t1 gnd 0.085993f
C544 diffpairibias.n4 gnd 0.13579f
C545 diffpairibias.t11 gnd 0.085993f
C546 diffpairibias.n5 gnd 0.072463f
C547 diffpairibias.t13 gnd 0.085993f
C548 diffpairibias.n6 gnd 0.072463f
C549 diffpairibias.t7 gnd 0.085993f
C550 diffpairibias.n7 gnd 0.072463f
C551 diffpairibias.t3 gnd 0.085993f
C552 diffpairibias.n8 gnd 0.072463f
C553 diffpairibias.t17 gnd 0.085993f
C554 diffpairibias.n9 gnd 0.072463f
C555 diffpairibias.t5 gnd 0.085993f
C556 diffpairibias.n10 gnd 0.072463f
C557 diffpairibias.t19 gnd 0.085993f
C558 diffpairibias.n11 gnd 0.072463f
C559 diffpairibias.t9 gnd 0.085993f
C560 diffpairibias.n12 gnd 0.102883f
C561 diffpairibias.t14 gnd 0.086899f
C562 diffpairibias.t0 gnd 0.086748f
C563 diffpairibias.n13 gnd 0.094648f
C564 diffpairibias.t10 gnd 0.086748f
C565 diffpairibias.n14 gnd 0.052262f
C566 diffpairibias.t12 gnd 0.086748f
C567 diffpairibias.n15 gnd 0.052262f
C568 diffpairibias.t6 gnd 0.086748f
C569 diffpairibias.n16 gnd 0.052262f
C570 diffpairibias.t2 gnd 0.086748f
C571 diffpairibias.n17 gnd 0.052262f
C572 diffpairibias.t16 gnd 0.086748f
C573 diffpairibias.n18 gnd 0.052262f
C574 diffpairibias.t4 gnd 0.086748f
C575 diffpairibias.n19 gnd 0.052262f
C576 diffpairibias.t18 gnd 0.086748f
C577 diffpairibias.n20 gnd 0.052262f
C578 diffpairibias.t8 gnd 0.086748f
C579 diffpairibias.n21 gnd 0.061849f
C580 diffpairibias.n22 gnd 0.233513f
C581 diffpairibias.t20 gnd 0.08996f
C582 diffpairibias.n23 gnd 0.051747f
C583 diffpairibias.t26 gnd 0.08996f
C584 diffpairibias.n24 gnd 0.051736f
C585 diffpairibias.t22 gnd 0.08996f
C586 diffpairibias.n25 gnd 0.051736f
C587 diffpairibias.t21 gnd 0.08996f
C588 diffpairibias.n26 gnd 0.051736f
C589 diffpairibias.t24 gnd 0.08996f
C590 diffpairibias.n27 gnd 0.04729f
C591 diffpairibias.n28 gnd 0.047711f
C592 a_n3827_n3924.t39 gnd 0.095164f
C593 a_n3827_n3924.t42 gnd 0.989053f
C594 a_n3827_n3924.n0 gnd 0.61435f
C595 a_n3827_n3924.t38 gnd 0.989053f
C596 a_n3827_n3924.n1 gnd 0.925837f
C597 a_n3827_n3924.t36 gnd 0.095164f
C598 a_n3827_n3924.t34 gnd 0.095164f
C599 a_n3827_n3924.n2 gnd 0.777221f
C600 a_n3827_n3924.n3 gnd 0.391675f
C601 a_n3827_n3924.t47 gnd 0.095164f
C602 a_n3827_n3924.t52 gnd 0.095164f
C603 a_n3827_n3924.n4 gnd 0.777221f
C604 a_n3827_n3924.n5 gnd 0.391675f
C605 a_n3827_n3924.t45 gnd 0.095164f
C606 a_n3827_n3924.t49 gnd 0.095164f
C607 a_n3827_n3924.n6 gnd 0.777221f
C608 a_n3827_n3924.n7 gnd 0.391675f
C609 a_n3827_n3924.t41 gnd 0.095164f
C610 a_n3827_n3924.t46 gnd 0.095164f
C611 a_n3827_n3924.n8 gnd 0.777221f
C612 a_n3827_n3924.n9 gnd 0.391675f
C613 a_n3827_n3924.t57 gnd 0.095164f
C614 a_n3827_n3924.t40 gnd 0.095164f
C615 a_n3827_n3924.n10 gnd 0.777221f
C616 a_n3827_n3924.n11 gnd 0.391675f
C617 a_n3827_n3924.t51 gnd 0.989057f
C618 a_n3827_n3924.n12 gnd 0.373908f
C619 a_n3827_n3924.t31 gnd 0.989057f
C620 a_n3827_n3924.n13 gnd 0.373908f
C621 a_n3827_n3924.t32 gnd 0.095164f
C622 a_n3827_n3924.t24 gnd 0.095164f
C623 a_n3827_n3924.n14 gnd 0.777221f
C624 a_n3827_n3924.n15 gnd 0.391675f
C625 a_n3827_n3924.t27 gnd 0.095164f
C626 a_n3827_n3924.t12 gnd 0.095164f
C627 a_n3827_n3924.n16 gnd 0.777221f
C628 a_n3827_n3924.n17 gnd 0.391675f
C629 a_n3827_n3924.t5 gnd 0.095164f
C630 a_n3827_n3924.t9 gnd 0.095164f
C631 a_n3827_n3924.n18 gnd 0.777221f
C632 a_n3827_n3924.n19 gnd 0.391675f
C633 a_n3827_n3924.t26 gnd 0.095164f
C634 a_n3827_n3924.t16 gnd 0.095164f
C635 a_n3827_n3924.n20 gnd 0.777221f
C636 a_n3827_n3924.n21 gnd 0.391675f
C637 a_n3827_n3924.t33 gnd 0.095164f
C638 a_n3827_n3924.t25 gnd 0.095164f
C639 a_n3827_n3924.n22 gnd 0.777221f
C640 a_n3827_n3924.n23 gnd 0.391675f
C641 a_n3827_n3924.t11 gnd 0.989057f
C642 a_n3827_n3924.n24 gnd 0.925833f
C643 a_n3827_n3924.n25 gnd 0.897154f
C644 a_n3827_n3924.t13 gnd 1.23041f
C645 a_n3827_n3924.n26 gnd 1.00053f
C646 a_n3827_n3924.t20 gnd 1.22888f
C647 a_n3827_n3924.n27 gnd 0.565437f
C648 a_n3827_n3924.t0 gnd 1.22888f
C649 a_n3827_n3924.n28 gnd 0.865521f
C650 a_n3827_n3924.t22 gnd 1.22888f
C651 a_n3827_n3924.n29 gnd 0.865521f
C652 a_n3827_n3924.t1 gnd 1.22888f
C653 a_n3827_n3924.n30 gnd 0.865521f
C654 a_n3827_n3924.t28 gnd 1.22888f
C655 a_n3827_n3924.n31 gnd 0.865521f
C656 a_n3827_n3924.t6 gnd 1.22888f
C657 a_n3827_n3924.n32 gnd 0.865521f
C658 a_n3827_n3924.t3 gnd 1.22888f
C659 a_n3827_n3924.n33 gnd 0.865521f
C660 a_n3827_n3924.t23 gnd 1.22888f
C661 a_n3827_n3924.n34 gnd 0.823361f
C662 a_n3827_n3924.t7 gnd 1.2292f
C663 a_n3827_n3924.n35 gnd 1.25966f
C664 a_n3827_n3924.n36 gnd 0.897154f
C665 a_n3827_n3924.t15 gnd 0.989053f
C666 a_n3827_n3924.n37 gnd 0.61435f
C667 a_n3827_n3924.t19 gnd 0.095164f
C668 a_n3827_n3924.t29 gnd 0.095164f
C669 a_n3827_n3924.n38 gnd 0.777219f
C670 a_n3827_n3924.n39 gnd 0.391676f
C671 a_n3827_n3924.t18 gnd 0.095164f
C672 a_n3827_n3924.t10 gnd 0.095164f
C673 a_n3827_n3924.n40 gnd 0.777219f
C674 a_n3827_n3924.n41 gnd 0.391676f
C675 a_n3827_n3924.t4 gnd 0.095164f
C676 a_n3827_n3924.t17 gnd 0.095164f
C677 a_n3827_n3924.n42 gnd 0.777219f
C678 a_n3827_n3924.n43 gnd 0.391676f
C679 a_n3827_n3924.t14 gnd 0.095164f
C680 a_n3827_n3924.t2 gnd 0.095164f
C681 a_n3827_n3924.n44 gnd 0.777219f
C682 a_n3827_n3924.n45 gnd 0.391676f
C683 a_n3827_n3924.t30 gnd 0.095164f
C684 a_n3827_n3924.t21 gnd 0.095164f
C685 a_n3827_n3924.n46 gnd 0.777219f
C686 a_n3827_n3924.n47 gnd 0.391676f
C687 a_n3827_n3924.t8 gnd 0.989053f
C688 a_n3827_n3924.n48 gnd 0.373911f
C689 a_n3827_n3924.t48 gnd 0.989053f
C690 a_n3827_n3924.n49 gnd 0.373911f
C691 a_n3827_n3924.t37 gnd 0.095164f
C692 a_n3827_n3924.t53 gnd 0.095164f
C693 a_n3827_n3924.n50 gnd 0.777219f
C694 a_n3827_n3924.n51 gnd 0.391676f
C695 a_n3827_n3924.t44 gnd 0.095164f
C696 a_n3827_n3924.t35 gnd 0.095164f
C697 a_n3827_n3924.n52 gnd 0.777219f
C698 a_n3827_n3924.n53 gnd 0.391676f
C699 a_n3827_n3924.t55 gnd 0.095164f
C700 a_n3827_n3924.t43 gnd 0.095164f
C701 a_n3827_n3924.n54 gnd 0.777219f
C702 a_n3827_n3924.n55 gnd 0.391676f
C703 a_n3827_n3924.t50 gnd 0.095164f
C704 a_n3827_n3924.t54 gnd 0.095164f
C705 a_n3827_n3924.n56 gnd 0.777219f
C706 a_n3827_n3924.n57 gnd 0.391676f
C707 a_n3827_n3924.n58 gnd 0.39168f
C708 a_n3827_n3924.n59 gnd 0.777216f
C709 a_n3827_n3924.t56 gnd 0.095164f
C710 plus.n0 gnd 0.022919f
C711 plus.t20 gnd 0.416794f
C712 plus.t23 gnd 0.385385f
C713 plus.n1 gnd 0.155867f
C714 plus.n2 gnd 0.022919f
C715 plus.t6 gnd 0.385385f
C716 plus.n3 gnd 0.019585f
C717 plus.n4 gnd 0.022919f
C718 plus.t12 gnd 0.385385f
C719 plus.t8 gnd 0.385385f
C720 plus.n5 gnd 0.155867f
C721 plus.n6 gnd 0.022919f
C722 plus.t7 gnd 0.385385f
C723 plus.n7 gnd 0.155867f
C724 plus.n8 gnd 0.022919f
C725 plus.t19 gnd 0.385385f
C726 plus.n9 gnd 0.018628f
C727 plus.n10 gnd 0.022919f
C728 plus.t18 gnd 0.385385f
C729 plus.t27 gnd 0.385385f
C730 plus.n11 gnd 0.155867f
C731 plus.n12 gnd 0.022919f
C732 plus.t25 gnd 0.385385f
C733 plus.n13 gnd 0.155867f
C734 plus.n14 gnd 0.097267f
C735 plus.t9 gnd 0.385385f
C736 plus.t14 gnd 0.431123f
C737 plus.n15 gnd 0.182224f
C738 plus.n16 gnd 0.178497f
C739 plus.n17 gnd 0.029367f
C740 plus.n18 gnd 0.025936f
C741 plus.n19 gnd 0.022919f
C742 plus.n20 gnd 0.022919f
C743 plus.n21 gnd 0.027389f
C744 plus.n22 gnd 0.019585f
C745 plus.n23 gnd 0.029849f
C746 plus.n24 gnd 0.022919f
C747 plus.n25 gnd 0.022919f
C748 plus.n26 gnd 0.02851f
C749 plus.n27 gnd 0.026794f
C750 plus.n28 gnd 0.155867f
C751 plus.n29 gnd 0.02871f
C752 plus.n30 gnd 0.022919f
C753 plus.n31 gnd 0.022919f
C754 plus.n32 gnd 0.022919f
C755 plus.n33 gnd 0.029485f
C756 plus.n34 gnd 0.155867f
C757 plus.n35 gnd 0.027652f
C758 plus.n36 gnd 0.027652f
C759 plus.n37 gnd 0.022919f
C760 plus.n38 gnd 0.022919f
C761 plus.n39 gnd 0.029485f
C762 plus.n40 gnd 0.018628f
C763 plus.n41 gnd 0.02871f
C764 plus.n42 gnd 0.022919f
C765 plus.n43 gnd 0.022919f
C766 plus.n44 gnd 0.026794f
C767 plus.n45 gnd 0.02851f
C768 plus.n46 gnd 0.155867f
C769 plus.n47 gnd 0.029849f
C770 plus.n48 gnd 0.022919f
C771 plus.n49 gnd 0.022919f
C772 plus.n50 gnd 0.022919f
C773 plus.n51 gnd 0.027389f
C774 plus.n52 gnd 0.155867f
C775 plus.n53 gnd 0.025936f
C776 plus.n54 gnd 0.029367f
C777 plus.n55 gnd 0.022919f
C778 plus.n56 gnd 0.022919f
C779 plus.n57 gnd 0.029899f
C780 plus.n58 gnd 0.00833f
C781 plus.n59 gnd 0.180467f
C782 plus.n60 gnd 0.262595f
C783 plus.n61 gnd 0.022919f
C784 plus.t28 gnd 0.385385f
C785 plus.n62 gnd 0.155867f
C786 plus.n63 gnd 0.022919f
C787 plus.t26 gnd 0.385385f
C788 plus.n64 gnd 0.019585f
C789 plus.n65 gnd 0.022919f
C790 plus.t10 gnd 0.385385f
C791 plus.t15 gnd 0.385385f
C792 plus.n66 gnd 0.155867f
C793 plus.n67 gnd 0.022919f
C794 plus.t13 gnd 0.385385f
C795 plus.n68 gnd 0.155867f
C796 plus.n69 gnd 0.022919f
C797 plus.t17 gnd 0.385385f
C798 plus.n70 gnd 0.018628f
C799 plus.n71 gnd 0.022919f
C800 plus.t16 gnd 0.385385f
C801 plus.t21 gnd 0.385385f
C802 plus.n72 gnd 0.155867f
C803 plus.n73 gnd 0.022919f
C804 plus.t22 gnd 0.385385f
C805 plus.n74 gnd 0.155867f
C806 plus.n75 gnd 0.097267f
C807 plus.t5 gnd 0.385385f
C808 plus.t11 gnd 0.431123f
C809 plus.n76 gnd 0.182224f
C810 plus.n77 gnd 0.178497f
C811 plus.n78 gnd 0.029367f
C812 plus.n79 gnd 0.025936f
C813 plus.n80 gnd 0.022919f
C814 plus.n81 gnd 0.022919f
C815 plus.n82 gnd 0.027389f
C816 plus.n83 gnd 0.019585f
C817 plus.n84 gnd 0.029849f
C818 plus.n85 gnd 0.022919f
C819 plus.n86 gnd 0.022919f
C820 plus.n87 gnd 0.02851f
C821 plus.n88 gnd 0.026794f
C822 plus.n89 gnd 0.155867f
C823 plus.n90 gnd 0.02871f
C824 plus.n91 gnd 0.022919f
C825 plus.n92 gnd 0.022919f
C826 plus.n93 gnd 0.022919f
C827 plus.n94 gnd 0.029485f
C828 plus.n95 gnd 0.155867f
C829 plus.n96 gnd 0.027652f
C830 plus.n97 gnd 0.027652f
C831 plus.n98 gnd 0.022919f
C832 plus.n99 gnd 0.022919f
C833 plus.n100 gnd 0.029485f
C834 plus.n101 gnd 0.018628f
C835 plus.n102 gnd 0.02871f
C836 plus.n103 gnd 0.022919f
C837 plus.n104 gnd 0.022919f
C838 plus.n105 gnd 0.026794f
C839 plus.n106 gnd 0.02851f
C840 plus.n107 gnd 0.155867f
C841 plus.n108 gnd 0.029849f
C842 plus.n109 gnd 0.022919f
C843 plus.n110 gnd 0.022919f
C844 plus.n111 gnd 0.022919f
C845 plus.n112 gnd 0.027389f
C846 plus.n113 gnd 0.155867f
C847 plus.n114 gnd 0.025936f
C848 plus.n115 gnd 0.029367f
C849 plus.n116 gnd 0.022919f
C850 plus.n117 gnd 0.022919f
C851 plus.n118 gnd 0.029899f
C852 plus.n119 gnd 0.00833f
C853 plus.t24 gnd 0.416794f
C854 plus.n120 gnd 0.180467f
C855 plus.n121 gnd 0.82692f
C856 plus.n122 gnd 1.21905f
C857 plus.t1 gnd 0.039565f
C858 plus.t2 gnd 0.007065f
C859 plus.t4 gnd 0.007065f
C860 plus.n123 gnd 0.022914f
C861 plus.n124 gnd 0.177885f
C862 plus.t3 gnd 0.007065f
C863 plus.t0 gnd 0.007065f
C864 plus.n125 gnd 0.022914f
C865 plus.n126 gnd 0.133524f
C866 plus.n127 gnd 3.00933f
C867 a_n1808_13878.t7 gnd 0.185195f
C868 a_n1808_13878.t2 gnd 0.185195f
C869 a_n1808_13878.t4 gnd 0.185195f
C870 a_n1808_13878.n0 gnd 1.4598f
C871 a_n1808_13878.t8 gnd 0.185195f
C872 a_n1808_13878.t3 gnd 0.185195f
C873 a_n1808_13878.n1 gnd 1.45825f
C874 a_n1808_13878.n2 gnd 2.03762f
C875 a_n1808_13878.t6 gnd 0.185195f
C876 a_n1808_13878.t1 gnd 0.185195f
C877 a_n1808_13878.n3 gnd 1.45825f
C878 a_n1808_13878.n4 gnd 3.69301f
C879 a_n1808_13878.t13 gnd 1.73408f
C880 a_n1808_13878.t16 gnd 0.185195f
C881 a_n1808_13878.t17 gnd 0.185195f
C882 a_n1808_13878.n5 gnd 1.30452f
C883 a_n1808_13878.n6 gnd 1.4576f
C884 a_n1808_13878.t12 gnd 1.73062f
C885 a_n1808_13878.n7 gnd 0.733487f
C886 a_n1808_13878.t15 gnd 1.73062f
C887 a_n1808_13878.n8 gnd 0.733487f
C888 a_n1808_13878.t18 gnd 0.185195f
C889 a_n1808_13878.t19 gnd 0.185195f
C890 a_n1808_13878.n9 gnd 1.30452f
C891 a_n1808_13878.n10 gnd 0.74059f
C892 a_n1808_13878.t14 gnd 1.73062f
C893 a_n1808_13878.n11 gnd 1.7272f
C894 a_n1808_13878.n12 gnd 2.51438f
C895 a_n1808_13878.t9 gnd 0.185195f
C896 a_n1808_13878.t10 gnd 0.185195f
C897 a_n1808_13878.n13 gnd 1.45825f
C898 a_n1808_13878.n14 gnd 1.80025f
C899 a_n1808_13878.t0 gnd 0.185195f
C900 a_n1808_13878.t5 gnd 0.185195f
C901 a_n1808_13878.n15 gnd 1.45825f
C902 a_n1808_13878.n16 gnd 1.31079f
C903 a_n1808_13878.n17 gnd 1.46067f
C904 a_n1808_13878.t11 gnd 0.185195f
C905 a_n2848_n452.n0 gnd 4.40606f
C906 a_n2848_n452.n1 gnd 3.15028f
C907 a_n2848_n452.n2 gnd 4.02851f
C908 a_n2848_n452.n3 gnd 0.912814f
C909 a_n2848_n452.n4 gnd 0.912816f
C910 a_n2848_n452.n5 gnd 3.415f
C911 a_n2848_n452.n6 gnd 0.285666f
C912 a_n2848_n452.n7 gnd 0.492471f
C913 a_n2848_n452.n8 gnd 0.664435f
C914 a_n2848_n452.n9 gnd 0.215942f
C915 a_n2848_n452.n10 gnd 0.282512f
C916 a_n2848_n452.n11 gnd 0.546457f
C917 a_n2848_n452.n12 gnd 0.526038f
C918 a_n2848_n452.n13 gnd 0.204894f
C919 a_n2848_n452.n14 gnd 0.150908f
C920 a_n2848_n452.n15 gnd 0.23718f
C921 a_n2848_n452.n16 gnd 0.183194f
C922 a_n2848_n452.n17 gnd 0.204894f
C923 a_n2848_n452.n18 gnd 1.0063f
C924 a_n2848_n452.n19 gnd 0.150908f
C925 a_n2848_n452.n20 gnd 0.580023f
C926 a_n2848_n452.n21 gnd 0.432289f
C927 a_n2848_n452.n22 gnd 0.215942f
C928 a_n2848_n452.n23 gnd 0.492471f
C929 a_n2848_n452.n24 gnd 0.282512f
C930 a_n2848_n452.n25 gnd 0.438486f
C931 a_n2848_n452.n26 gnd 0.215942f
C932 a_n2848_n452.n27 gnd 0.731534f
C933 a_n2848_n452.n28 gnd 0.282512f
C934 a_n2848_n452.n29 gnd 1.17886f
C935 a_n2848_n452.n30 gnd 1.91568f
C936 a_n2848_n452.n31 gnd 1.14458f
C937 a_n2848_n452.n32 gnd 1.77783f
C938 a_n2848_n452.n33 gnd 0.008361f
C939 a_n2848_n452.n35 gnd 0.285666f
C940 a_n2848_n452.n36 gnd 0.008361f
C941 a_n2848_n452.n38 gnd 0.285666f
C942 a_n2848_n452.n39 gnd 0.008361f
C943 a_n2848_n452.n40 gnd 0.28526f
C944 a_n2848_n452.n41 gnd 0.008361f
C945 a_n2848_n452.n42 gnd 0.28526f
C946 a_n2848_n452.n43 gnd 0.008361f
C947 a_n2848_n452.n44 gnd 0.28526f
C948 a_n2848_n452.n45 gnd 0.008361f
C949 a_n2848_n452.n46 gnd 0.28526f
C950 a_n2848_n452.n48 gnd 0.285666f
C951 a_n2848_n452.n49 gnd 0.008361f
C952 a_n2848_n452.n51 gnd 0.285666f
C953 a_n2848_n452.t6 gnd 0.14978f
C954 a_n2848_n452.t25 gnd 0.708223f
C955 a_n2848_n452.t23 gnd 0.696704f
C956 a_n2848_n452.t11 gnd 0.696704f
C957 a_n2848_n452.t27 gnd 0.116496f
C958 a_n2848_n452.t44 gnd 0.116496f
C959 a_n2848_n452.n53 gnd 1.03243f
C960 a_n2848_n452.t38 gnd 0.116496f
C961 a_n2848_n452.t32 gnd 0.116496f
C962 a_n2848_n452.n54 gnd 1.02939f
C963 a_n2848_n452.t0 gnd 0.116496f
C964 a_n2848_n452.t1 gnd 0.116496f
C965 a_n2848_n452.n55 gnd 1.02939f
C966 a_n2848_n452.t43 gnd 0.116496f
C967 a_n2848_n452.t33 gnd 0.116496f
C968 a_n2848_n452.n56 gnd 1.03243f
C969 a_n2848_n452.t29 gnd 0.116496f
C970 a_n2848_n452.t37 gnd 0.116496f
C971 a_n2848_n452.n57 gnd 1.02939f
C972 a_n2848_n452.t35 gnd 0.116496f
C973 a_n2848_n452.t36 gnd 0.116496f
C974 a_n2848_n452.n58 gnd 1.02939f
C975 a_n2848_n452.t30 gnd 0.116496f
C976 a_n2848_n452.t47 gnd 0.116496f
C977 a_n2848_n452.n59 gnd 1.0294f
C978 a_n2848_n452.t40 gnd 0.116496f
C979 a_n2848_n452.t41 gnd 0.116496f
C980 a_n2848_n452.n60 gnd 1.0294f
C981 a_n2848_n452.t34 gnd 0.116496f
C982 a_n2848_n452.t2 gnd 0.116496f
C983 a_n2848_n452.n61 gnd 1.0294f
C984 a_n2848_n452.t39 gnd 0.116496f
C985 a_n2848_n452.t45 gnd 0.116496f
C986 a_n2848_n452.n62 gnd 1.03243f
C987 a_n2848_n452.t31 gnd 0.116496f
C988 a_n2848_n452.t46 gnd 0.116496f
C989 a_n2848_n452.n63 gnd 1.0294f
C990 a_n2848_n452.t28 gnd 0.116496f
C991 a_n2848_n452.t42 gnd 0.116496f
C992 a_n2848_n452.n64 gnd 1.0294f
C993 a_n2848_n452.t3 gnd 0.696704f
C994 a_n2848_n452.n65 gnd 0.302425f
C995 a_n2848_n452.t5 gnd 0.696704f
C996 a_n2848_n452.t19 gnd 0.708223f
C997 a_n2848_n452.t74 gnd 0.711378f
C998 a_n2848_n452.t57 gnd 0.696704f
C999 a_n2848_n452.t61 gnd 0.696704f
C1000 a_n2848_n452.t51 gnd 0.696704f
C1001 a_n2848_n452.n66 gnd 0.306315f
C1002 a_n2848_n452.t66 gnd 0.696704f
C1003 a_n2848_n452.t72 gnd 0.708223f
C1004 a_n2848_n452.t10 gnd 1.40246f
C1005 a_n2848_n452.t18 gnd 0.14978f
C1006 a_n2848_n452.t14 gnd 0.14978f
C1007 a_n2848_n452.n67 gnd 1.05505f
C1008 a_n2848_n452.t16 gnd 0.14978f
C1009 a_n2848_n452.t8 gnd 0.14978f
C1010 a_n2848_n452.n68 gnd 1.05505f
C1011 a_n2848_n452.t22 gnd 1.39967f
C1012 a_n2848_n452.t15 gnd 0.696704f
C1013 a_n2848_n452.n69 gnd 0.306315f
C1014 a_n2848_n452.t7 gnd 0.696704f
C1015 a_n2848_n452.t17 gnd 0.696704f
C1016 a_n2848_n452.t56 gnd 0.696704f
C1017 a_n2848_n452.n70 gnd 0.306315f
C1018 a_n2848_n452.t64 gnd 0.696704f
C1019 a_n2848_n452.t70 gnd 0.696704f
C1020 a_n2848_n452.t69 gnd 0.711378f
C1021 a_n2848_n452.n71 gnd 0.308932f
C1022 a_n2848_n452.t49 gnd 0.696704f
C1023 a_n2848_n452.n72 gnd 0.302425f
C1024 a_n2848_n452.n73 gnd 0.308933f
C1025 a_n2848_n452.t50 gnd 0.708223f
C1026 a_n2848_n452.t9 gnd 0.711378f
C1027 a_n2848_n452.n74 gnd 0.308932f
C1028 a_n2848_n452.t13 gnd 0.696704f
C1029 a_n2848_n452.n75 gnd 0.302425f
C1030 a_n2848_n452.n76 gnd 0.308933f
C1031 a_n2848_n452.t21 gnd 0.708223f
C1032 a_n2848_n452.n77 gnd 1.13204f
C1033 a_n2848_n452.t54 gnd 0.696704f
C1034 a_n2848_n452.n78 gnd 0.302425f
C1035 a_n2848_n452.t60 gnd 0.696704f
C1036 a_n2848_n452.n79 gnd 0.302425f
C1037 a_n2848_n452.t52 gnd 0.696704f
C1038 a_n2848_n452.n80 gnd 0.302425f
C1039 a_n2848_n452.t65 gnd 0.696704f
C1040 a_n2848_n452.n81 gnd 0.302425f
C1041 a_n2848_n452.t55 gnd 0.696704f
C1042 a_n2848_n452.n82 gnd 0.296933f
C1043 a_n2848_n452.t75 gnd 0.696704f
C1044 a_n2848_n452.n83 gnd 0.306315f
C1045 a_n2848_n452.t58 gnd 0.708378f
C1046 a_n2848_n452.t67 gnd 0.696704f
C1047 a_n2848_n452.n84 gnd 0.296933f
C1048 a_n2848_n452.t53 gnd 0.696704f
C1049 a_n2848_n452.n85 gnd 0.306315f
C1050 a_n2848_n452.t62 gnd 0.708378f
C1051 a_n2848_n452.t71 gnd 0.696704f
C1052 a_n2848_n452.n86 gnd 0.296933f
C1053 a_n2848_n452.t59 gnd 0.696704f
C1054 a_n2848_n452.n87 gnd 0.306315f
C1055 a_n2848_n452.t73 gnd 0.708378f
C1056 a_n2848_n452.t63 gnd 0.696704f
C1057 a_n2848_n452.n88 gnd 0.296933f
C1058 a_n2848_n452.t48 gnd 0.696704f
C1059 a_n2848_n452.n89 gnd 0.306315f
C1060 a_n2848_n452.t68 gnd 0.708378f
C1061 a_n2848_n452.n90 gnd 1.33845f
C1062 a_n2848_n452.n91 gnd 0.308933f
C1063 a_n2848_n452.n92 gnd 0.302425f
C1064 a_n2848_n452.n93 gnd 0.308932f
C1065 a_n2848_n452.n94 gnd 0.308933f
C1066 a_n2848_n452.n95 gnd 0.01225f
C1067 a_n2848_n452.n96 gnd 0.302425f
C1068 a_n2848_n452.n97 gnd 0.308933f
C1069 a_n2848_n452.n98 gnd 0.786935f
C1070 a_n2848_n452.t26 gnd 1.39967f
C1071 a_n2848_n452.t24 gnd 0.14978f
C1072 a_n2848_n452.t12 gnd 0.14978f
C1073 a_n2848_n452.n99 gnd 1.05505f
C1074 a_n2848_n452.t20 gnd 1.40246f
C1075 a_n2848_n452.n100 gnd 1.05505f
C1076 a_n2848_n452.t4 gnd 0.14978f
C1077 CSoutput.n0 gnd 0.04544f
C1078 CSoutput.t195 gnd 0.300579f
C1079 CSoutput.n1 gnd 0.135726f
C1080 CSoutput.n2 gnd 0.04544f
C1081 CSoutput.t199 gnd 0.300579f
C1082 CSoutput.n3 gnd 0.036015f
C1083 CSoutput.n4 gnd 0.04544f
C1084 CSoutput.t211 gnd 0.300579f
C1085 CSoutput.n5 gnd 0.031056f
C1086 CSoutput.n6 gnd 0.04544f
C1087 CSoutput.t197 gnd 0.300579f
C1088 CSoutput.t203 gnd 0.300579f
C1089 CSoutput.n7 gnd 0.134247f
C1090 CSoutput.n8 gnd 0.04544f
C1091 CSoutput.t201 gnd 0.300579f
C1092 CSoutput.n9 gnd 0.02961f
C1093 CSoutput.n10 gnd 0.04544f
C1094 CSoutput.t213 gnd 0.300579f
C1095 CSoutput.t200 gnd 0.300579f
C1096 CSoutput.n11 gnd 0.134247f
C1097 CSoutput.n12 gnd 0.04544f
C1098 CSoutput.t198 gnd 0.300579f
C1099 CSoutput.n13 gnd 0.031056f
C1100 CSoutput.n14 gnd 0.04544f
C1101 CSoutput.t210 gnd 0.300579f
C1102 CSoutput.t194 gnd 0.300579f
C1103 CSoutput.n15 gnd 0.134247f
C1104 CSoutput.n16 gnd 0.04544f
C1105 CSoutput.t196 gnd 0.300579f
C1106 CSoutput.n17 gnd 0.03317f
C1107 CSoutput.t206 gnd 0.3592f
C1108 CSoutput.t208 gnd 0.300579f
C1109 CSoutput.n18 gnd 0.171382f
C1110 CSoutput.n19 gnd 0.166299f
C1111 CSoutput.n20 gnd 0.192927f
C1112 CSoutput.n21 gnd 0.04544f
C1113 CSoutput.n22 gnd 0.037925f
C1114 CSoutput.n23 gnd 0.134247f
C1115 CSoutput.n24 gnd 0.036559f
C1116 CSoutput.n25 gnd 0.036015f
C1117 CSoutput.n26 gnd 0.04544f
C1118 CSoutput.n27 gnd 0.04544f
C1119 CSoutput.n28 gnd 0.037634f
C1120 CSoutput.n29 gnd 0.031952f
C1121 CSoutput.n30 gnd 0.137236f
C1122 CSoutput.n31 gnd 0.032392f
C1123 CSoutput.n32 gnd 0.04544f
C1124 CSoutput.n33 gnd 0.04544f
C1125 CSoutput.n34 gnd 0.04544f
C1126 CSoutput.n35 gnd 0.037233f
C1127 CSoutput.n36 gnd 0.134247f
C1128 CSoutput.n37 gnd 0.035608f
C1129 CSoutput.n38 gnd 0.036966f
C1130 CSoutput.n39 gnd 0.04544f
C1131 CSoutput.n40 gnd 0.04544f
C1132 CSoutput.n41 gnd 0.037917f
C1133 CSoutput.n42 gnd 0.034657f
C1134 CSoutput.n43 gnd 0.134247f
C1135 CSoutput.n44 gnd 0.035535f
C1136 CSoutput.n45 gnd 0.04544f
C1137 CSoutput.n46 gnd 0.04544f
C1138 CSoutput.n47 gnd 0.04544f
C1139 CSoutput.n48 gnd 0.035535f
C1140 CSoutput.n49 gnd 0.134247f
C1141 CSoutput.n50 gnd 0.034657f
C1142 CSoutput.n51 gnd 0.037917f
C1143 CSoutput.n52 gnd 0.04544f
C1144 CSoutput.n53 gnd 0.04544f
C1145 CSoutput.n54 gnd 0.036966f
C1146 CSoutput.n55 gnd 0.035608f
C1147 CSoutput.n56 gnd 0.134247f
C1148 CSoutput.n57 gnd 0.037233f
C1149 CSoutput.n58 gnd 0.04544f
C1150 CSoutput.n59 gnd 0.04544f
C1151 CSoutput.n60 gnd 0.04544f
C1152 CSoutput.n61 gnd 0.032392f
C1153 CSoutput.n62 gnd 0.137236f
C1154 CSoutput.n63 gnd 0.031952f
C1155 CSoutput.t205 gnd 0.300579f
C1156 CSoutput.n64 gnd 0.134247f
C1157 CSoutput.n65 gnd 0.037634f
C1158 CSoutput.n66 gnd 0.04544f
C1159 CSoutput.n67 gnd 0.04544f
C1160 CSoutput.n68 gnd 0.04544f
C1161 CSoutput.n69 gnd 0.036559f
C1162 CSoutput.n70 gnd 0.134247f
C1163 CSoutput.n71 gnd 0.037925f
C1164 CSoutput.n72 gnd 0.03317f
C1165 CSoutput.n73 gnd 0.04544f
C1166 CSoutput.n74 gnd 0.04544f
C1167 CSoutput.n75 gnd 0.034399f
C1168 CSoutput.n76 gnd 0.02043f
C1169 CSoutput.t207 gnd 0.337722f
C1170 CSoutput.n77 gnd 0.167767f
C1171 CSoutput.n78 gnd 0.686326f
C1172 CSoutput.t82 gnd 0.056681f
C1173 CSoutput.t2 gnd 0.056681f
C1174 CSoutput.n79 gnd 0.438841f
C1175 CSoutput.t65 gnd 0.056681f
C1176 CSoutput.t42 gnd 0.056681f
C1177 CSoutput.n80 gnd 0.438058f
C1178 CSoutput.n81 gnd 0.444628f
C1179 CSoutput.t72 gnd 0.056681f
C1180 CSoutput.t22 gnd 0.056681f
C1181 CSoutput.n82 gnd 0.438058f
C1182 CSoutput.n83 gnd 0.219094f
C1183 CSoutput.t89 gnd 0.056681f
C1184 CSoutput.t36 gnd 0.056681f
C1185 CSoutput.n84 gnd 0.438058f
C1186 CSoutput.n85 gnd 0.219094f
C1187 CSoutput.t7 gnd 0.056681f
C1188 CSoutput.t50 gnd 0.056681f
C1189 CSoutput.n86 gnd 0.438058f
C1190 CSoutput.n87 gnd 0.219094f
C1191 CSoutput.t11 gnd 0.056681f
C1192 CSoutput.t30 gnd 0.056681f
C1193 CSoutput.n88 gnd 0.438058f
C1194 CSoutput.n89 gnd 0.219094f
C1195 CSoutput.t94 gnd 0.056681f
C1196 CSoutput.t44 gnd 0.056681f
C1197 CSoutput.n90 gnd 0.438058f
C1198 CSoutput.n91 gnd 0.219094f
C1199 CSoutput.t14 gnd 0.056681f
C1200 CSoutput.t78 gnd 0.056681f
C1201 CSoutput.n92 gnd 0.438058f
C1202 CSoutput.n93 gnd 0.401768f
C1203 CSoutput.t76 gnd 0.056681f
C1204 CSoutput.t74 gnd 0.056681f
C1205 CSoutput.n94 gnd 0.438841f
C1206 CSoutput.t59 gnd 0.056681f
C1207 CSoutput.t8 gnd 0.056681f
C1208 CSoutput.n95 gnd 0.438058f
C1209 CSoutput.n96 gnd 0.444628f
C1210 CSoutput.t3 gnd 0.056681f
C1211 CSoutput.t70 gnd 0.056681f
C1212 CSoutput.n97 gnd 0.438058f
C1213 CSoutput.n98 gnd 0.219094f
C1214 CSoutput.t58 gnd 0.056681f
C1215 CSoutput.t38 gnd 0.056681f
C1216 CSoutput.n99 gnd 0.438058f
C1217 CSoutput.n100 gnd 0.219094f
C1218 CSoutput.t23 gnd 0.056681f
C1219 CSoutput.t85 gnd 0.056681f
C1220 CSoutput.n101 gnd 0.438058f
C1221 CSoutput.n102 gnd 0.219094f
C1222 CSoutput.t57 gnd 0.056681f
C1223 CSoutput.t56 gnd 0.056681f
C1224 CSoutput.n103 gnd 0.438058f
C1225 CSoutput.n104 gnd 0.219094f
C1226 CSoutput.t47 gnd 0.056681f
C1227 CSoutput.t19 gnd 0.056681f
C1228 CSoutput.n105 gnd 0.438058f
C1229 CSoutput.n106 gnd 0.219094f
C1230 CSoutput.t6 gnd 0.056681f
C1231 CSoutput.t48 gnd 0.056681f
C1232 CSoutput.n107 gnd 0.438058f
C1233 CSoutput.n108 gnd 0.326724f
C1234 CSoutput.n109 gnd 0.411997f
C1235 CSoutput.t87 gnd 0.056681f
C1236 CSoutput.t86 gnd 0.056681f
C1237 CSoutput.n110 gnd 0.438841f
C1238 CSoutput.t68 gnd 0.056681f
C1239 CSoutput.t18 gnd 0.056681f
C1240 CSoutput.n111 gnd 0.438058f
C1241 CSoutput.n112 gnd 0.444628f
C1242 CSoutput.t15 gnd 0.056681f
C1243 CSoutput.t84 gnd 0.056681f
C1244 CSoutput.n113 gnd 0.438058f
C1245 CSoutput.n114 gnd 0.219094f
C1246 CSoutput.t66 gnd 0.056681f
C1247 CSoutput.t49 gnd 0.056681f
C1248 CSoutput.n115 gnd 0.438058f
C1249 CSoutput.n116 gnd 0.219094f
C1250 CSoutput.t32 gnd 0.056681f
C1251 CSoutput.t95 gnd 0.056681f
C1252 CSoutput.n117 gnd 0.438058f
C1253 CSoutput.n118 gnd 0.219094f
C1254 CSoutput.t64 gnd 0.056681f
C1255 CSoutput.t63 gnd 0.056681f
C1256 CSoutput.n119 gnd 0.438058f
C1257 CSoutput.n120 gnd 0.219094f
C1258 CSoutput.t54 gnd 0.056681f
C1259 CSoutput.t31 gnd 0.056681f
C1260 CSoutput.n121 gnd 0.438058f
C1261 CSoutput.n122 gnd 0.219094f
C1262 CSoutput.t17 gnd 0.056681f
C1263 CSoutput.t55 gnd 0.056681f
C1264 CSoutput.n123 gnd 0.438058f
C1265 CSoutput.n124 gnd 0.326724f
C1266 CSoutput.n125 gnd 0.460508f
C1267 CSoutput.n126 gnd 8.95232f
C1268 CSoutput.n128 gnd 0.803835f
C1269 CSoutput.n129 gnd 0.602876f
C1270 CSoutput.n130 gnd 0.803835f
C1271 CSoutput.n131 gnd 0.803835f
C1272 CSoutput.n132 gnd 2.16417f
C1273 CSoutput.n133 gnd 0.803835f
C1274 CSoutput.n134 gnd 0.803835f
C1275 CSoutput.t192 gnd 1.00479f
C1276 CSoutput.n135 gnd 0.803835f
C1277 CSoutput.n136 gnd 0.803835f
C1278 CSoutput.n140 gnd 0.803835f
C1279 CSoutput.n144 gnd 0.803835f
C1280 CSoutput.n145 gnd 0.803835f
C1281 CSoutput.n147 gnd 0.803835f
C1282 CSoutput.n152 gnd 0.803835f
C1283 CSoutput.n154 gnd 0.803835f
C1284 CSoutput.n155 gnd 0.803835f
C1285 CSoutput.n157 gnd 0.803835f
C1286 CSoutput.n158 gnd 0.803835f
C1287 CSoutput.n160 gnd 0.803835f
C1288 CSoutput.t204 gnd 13.432f
C1289 CSoutput.n162 gnd 0.803835f
C1290 CSoutput.n163 gnd 0.602876f
C1291 CSoutput.n164 gnd 0.803835f
C1292 CSoutput.n165 gnd 0.803835f
C1293 CSoutput.n166 gnd 2.16417f
C1294 CSoutput.n167 gnd 0.803835f
C1295 CSoutput.n168 gnd 0.803835f
C1296 CSoutput.t209 gnd 1.00479f
C1297 CSoutput.n169 gnd 0.803835f
C1298 CSoutput.n170 gnd 0.803835f
C1299 CSoutput.n174 gnd 0.803835f
C1300 CSoutput.n178 gnd 0.803835f
C1301 CSoutput.n179 gnd 0.803835f
C1302 CSoutput.n181 gnd 0.803835f
C1303 CSoutput.n186 gnd 0.803835f
C1304 CSoutput.n188 gnd 0.803835f
C1305 CSoutput.n189 gnd 0.803835f
C1306 CSoutput.n191 gnd 0.803835f
C1307 CSoutput.n192 gnd 0.803835f
C1308 CSoutput.n194 gnd 0.803835f
C1309 CSoutput.n195 gnd 0.602876f
C1310 CSoutput.n197 gnd 0.803835f
C1311 CSoutput.n198 gnd 0.602876f
C1312 CSoutput.n199 gnd 0.803835f
C1313 CSoutput.n200 gnd 0.803835f
C1314 CSoutput.n201 gnd 2.16417f
C1315 CSoutput.n202 gnd 0.803835f
C1316 CSoutput.n203 gnd 0.803835f
C1317 CSoutput.t202 gnd 1.00479f
C1318 CSoutput.n204 gnd 0.803835f
C1319 CSoutput.n205 gnd 2.16417f
C1320 CSoutput.n207 gnd 0.803835f
C1321 CSoutput.n208 gnd 0.803835f
C1322 CSoutput.n210 gnd 0.803835f
C1323 CSoutput.n211 gnd 0.803835f
C1324 CSoutput.t212 gnd 13.213099f
C1325 CSoutput.t193 gnd 13.432f
C1326 CSoutput.n217 gnd 2.52175f
C1327 CSoutput.n218 gnd 10.2727f
C1328 CSoutput.n219 gnd 10.7025f
C1329 CSoutput.n224 gnd 2.73173f
C1330 CSoutput.n230 gnd 0.803835f
C1331 CSoutput.n232 gnd 0.803835f
C1332 CSoutput.n234 gnd 0.803835f
C1333 CSoutput.n236 gnd 0.803835f
C1334 CSoutput.n238 gnd 0.803835f
C1335 CSoutput.n244 gnd 0.803835f
C1336 CSoutput.n251 gnd 1.47473f
C1337 CSoutput.n252 gnd 1.47473f
C1338 CSoutput.n253 gnd 0.803835f
C1339 CSoutput.n254 gnd 0.803835f
C1340 CSoutput.n256 gnd 0.602876f
C1341 CSoutput.n257 gnd 0.516309f
C1342 CSoutput.n259 gnd 0.602876f
C1343 CSoutput.n260 gnd 0.516309f
C1344 CSoutput.n261 gnd 0.602876f
C1345 CSoutput.n263 gnd 0.803835f
C1346 CSoutput.n265 gnd 2.16417f
C1347 CSoutput.n266 gnd 2.52175f
C1348 CSoutput.n267 gnd 9.448231f
C1349 CSoutput.n269 gnd 0.602876f
C1350 CSoutput.n270 gnd 1.55124f
C1351 CSoutput.n271 gnd 0.602876f
C1352 CSoutput.n273 gnd 0.803835f
C1353 CSoutput.n275 gnd 2.16417f
C1354 CSoutput.n276 gnd 4.71391f
C1355 CSoutput.t1 gnd 0.056681f
C1356 CSoutput.t81 gnd 0.056681f
C1357 CSoutput.n277 gnd 0.438841f
C1358 CSoutput.t41 gnd 0.056681f
C1359 CSoutput.t93 gnd 0.056681f
C1360 CSoutput.n278 gnd 0.438058f
C1361 CSoutput.n279 gnd 0.444628f
C1362 CSoutput.t21 gnd 0.056681f
C1363 CSoutput.t71 gnd 0.056681f
C1364 CSoutput.n280 gnd 0.438058f
C1365 CSoutput.n281 gnd 0.219094f
C1366 CSoutput.t35 gnd 0.056681f
C1367 CSoutput.t88 gnd 0.056681f
C1368 CSoutput.n282 gnd 0.438058f
C1369 CSoutput.n283 gnd 0.219094f
C1370 CSoutput.t67 gnd 0.056681f
C1371 CSoutput.t5 gnd 0.056681f
C1372 CSoutput.n284 gnd 0.438058f
C1373 CSoutput.n285 gnd 0.219094f
C1374 CSoutput.t29 gnd 0.056681f
C1375 CSoutput.t10 gnd 0.056681f
C1376 CSoutput.n286 gnd 0.438058f
C1377 CSoutput.n287 gnd 0.219094f
C1378 CSoutput.t43 gnd 0.056681f
C1379 CSoutput.t26 gnd 0.056681f
C1380 CSoutput.n288 gnd 0.438058f
C1381 CSoutput.n289 gnd 0.219094f
C1382 CSoutput.t77 gnd 0.056681f
C1383 CSoutput.t13 gnd 0.056681f
C1384 CSoutput.n290 gnd 0.438058f
C1385 CSoutput.n291 gnd 0.401768f
C1386 CSoutput.t45 gnd 0.056681f
C1387 CSoutput.t46 gnd 0.056681f
C1388 CSoutput.n292 gnd 0.438841f
C1389 CSoutput.t62 gnd 0.056681f
C1390 CSoutput.t4 gnd 0.056681f
C1391 CSoutput.n293 gnd 0.438058f
C1392 CSoutput.n294 gnd 0.444628f
C1393 CSoutput.t40 gnd 0.056681f
C1394 CSoutput.t60 gnd 0.056681f
C1395 CSoutput.n295 gnd 0.438058f
C1396 CSoutput.n296 gnd 0.219094f
C1397 CSoutput.t0 gnd 0.056681f
C1398 CSoutput.t27 gnd 0.056681f
C1399 CSoutput.n297 gnd 0.438058f
C1400 CSoutput.n298 gnd 0.219094f
C1401 CSoutput.t28 gnd 0.056681f
C1402 CSoutput.t83 gnd 0.056681f
C1403 CSoutput.n299 gnd 0.438058f
C1404 CSoutput.n300 gnd 0.219094f
C1405 CSoutput.t24 gnd 0.056681f
C1406 CSoutput.t25 gnd 0.056681f
C1407 CSoutput.n301 gnd 0.438058f
C1408 CSoutput.n302 gnd 0.219094f
C1409 CSoutput.t79 gnd 0.056681f
C1410 CSoutput.t80 gnd 0.056681f
C1411 CSoutput.n303 gnd 0.438058f
C1412 CSoutput.n304 gnd 0.219094f
C1413 CSoutput.t9 gnd 0.056681f
C1414 CSoutput.t61 gnd 0.056681f
C1415 CSoutput.n305 gnd 0.438058f
C1416 CSoutput.n306 gnd 0.326724f
C1417 CSoutput.n307 gnd 0.411997f
C1418 CSoutput.t52 gnd 0.056681f
C1419 CSoutput.t53 gnd 0.056681f
C1420 CSoutput.n308 gnd 0.438841f
C1421 CSoutput.t75 gnd 0.056681f
C1422 CSoutput.t16 gnd 0.056681f
C1423 CSoutput.n309 gnd 0.438058f
C1424 CSoutput.n310 gnd 0.444628f
C1425 CSoutput.t51 gnd 0.056681f
C1426 CSoutput.t69 gnd 0.056681f
C1427 CSoutput.n311 gnd 0.438058f
C1428 CSoutput.n312 gnd 0.219094f
C1429 CSoutput.t12 gnd 0.056681f
C1430 CSoutput.t37 gnd 0.056681f
C1431 CSoutput.n313 gnd 0.438058f
C1432 CSoutput.n314 gnd 0.219094f
C1433 CSoutput.t39 gnd 0.056681f
C1434 CSoutput.t92 gnd 0.056681f
C1435 CSoutput.n315 gnd 0.438058f
C1436 CSoutput.n316 gnd 0.219094f
C1437 CSoutput.t33 gnd 0.056681f
C1438 CSoutput.t34 gnd 0.056681f
C1439 CSoutput.n317 gnd 0.438058f
C1440 CSoutput.n318 gnd 0.219094f
C1441 CSoutput.t90 gnd 0.056681f
C1442 CSoutput.t91 gnd 0.056681f
C1443 CSoutput.n319 gnd 0.438058f
C1444 CSoutput.n320 gnd 0.219094f
C1445 CSoutput.t20 gnd 0.056681f
C1446 CSoutput.t73 gnd 0.056681f
C1447 CSoutput.n321 gnd 0.438057f
C1448 CSoutput.n322 gnd 0.326726f
C1449 CSoutput.n323 gnd 0.460508f
C1450 CSoutput.n324 gnd 12.5684f
C1451 CSoutput.t177 gnd 0.049596f
C1452 CSoutput.t109 gnd 0.049596f
C1453 CSoutput.n325 gnd 0.439711f
C1454 CSoutput.t159 gnd 0.049596f
C1455 CSoutput.t98 gnd 0.049596f
C1456 CSoutput.n326 gnd 0.438244f
C1457 CSoutput.n327 gnd 0.408362f
C1458 CSoutput.t143 gnd 0.049596f
C1459 CSoutput.t180 gnd 0.049596f
C1460 CSoutput.n328 gnd 0.438244f
C1461 CSoutput.n329 gnd 0.201303f
C1462 CSoutput.t131 gnd 0.049596f
C1463 CSoutput.t142 gnd 0.049596f
C1464 CSoutput.n330 gnd 0.438244f
C1465 CSoutput.n331 gnd 0.201303f
C1466 CSoutput.t101 gnd 0.049596f
C1467 CSoutput.t149 gnd 0.049596f
C1468 CSoutput.n332 gnd 0.438244f
C1469 CSoutput.n333 gnd 0.201303f
C1470 CSoutput.t163 gnd 0.049596f
C1471 CSoutput.t132 gnd 0.049596f
C1472 CSoutput.n334 gnd 0.438244f
C1473 CSoutput.n335 gnd 0.201303f
C1474 CSoutput.t145 gnd 0.049596f
C1475 CSoutput.t173 gnd 0.049596f
C1476 CSoutput.n336 gnd 0.438244f
C1477 CSoutput.n337 gnd 0.201303f
C1478 CSoutput.t108 gnd 0.049596f
C1479 CSoutput.t123 gnd 0.049596f
C1480 CSoutput.n338 gnd 0.438244f
C1481 CSoutput.n339 gnd 0.371292f
C1482 CSoutput.t140 gnd 0.049596f
C1483 CSoutput.t117 gnd 0.049596f
C1484 CSoutput.n340 gnd 0.439711f
C1485 CSoutput.t127 gnd 0.049596f
C1486 CSoutput.t139 gnd 0.049596f
C1487 CSoutput.n341 gnd 0.438244f
C1488 CSoutput.n342 gnd 0.408362f
C1489 CSoutput.t116 gnd 0.049596f
C1490 CSoutput.t129 gnd 0.049596f
C1491 CSoutput.n343 gnd 0.438244f
C1492 CSoutput.n344 gnd 0.201303f
C1493 CSoutput.t141 gnd 0.049596f
C1494 CSoutput.t115 gnd 0.049596f
C1495 CSoutput.n345 gnd 0.438244f
C1496 CSoutput.n346 gnd 0.201303f
C1497 CSoutput.t128 gnd 0.049596f
C1498 CSoutput.t106 gnd 0.049596f
C1499 CSoutput.n347 gnd 0.438244f
C1500 CSoutput.n348 gnd 0.201303f
C1501 CSoutput.t114 gnd 0.049596f
C1502 CSoutput.t130 gnd 0.049596f
C1503 CSoutput.n349 gnd 0.438244f
C1504 CSoutput.n350 gnd 0.201303f
C1505 CSoutput.t103 gnd 0.049596f
C1506 CSoutput.t186 gnd 0.049596f
C1507 CSoutput.n351 gnd 0.438244f
C1508 CSoutput.n352 gnd 0.201303f
C1509 CSoutput.t120 gnd 0.049596f
C1510 CSoutput.t191 gnd 0.049596f
C1511 CSoutput.n353 gnd 0.438244f
C1512 CSoutput.n354 gnd 0.305621f
C1513 CSoutput.n355 gnd 0.385483f
C1514 CSoutput.t107 gnd 0.049596f
C1515 CSoutput.t187 gnd 0.049596f
C1516 CSoutput.n356 gnd 0.439711f
C1517 CSoutput.t175 gnd 0.049596f
C1518 CSoutput.t121 gnd 0.049596f
C1519 CSoutput.n357 gnd 0.438244f
C1520 CSoutput.n358 gnd 0.408362f
C1521 CSoutput.t96 gnd 0.049596f
C1522 CSoutput.t181 gnd 0.049596f
C1523 CSoutput.n359 gnd 0.438244f
C1524 CSoutput.n360 gnd 0.201303f
C1525 CSoutput.t135 gnd 0.049596f
C1526 CSoutput.t144 gnd 0.049596f
C1527 CSoutput.n361 gnd 0.438244f
C1528 CSoutput.n362 gnd 0.201303f
C1529 CSoutput.t188 gnd 0.049596f
C1530 CSoutput.t174 gnd 0.049596f
C1531 CSoutput.n363 gnd 0.438244f
C1532 CSoutput.n364 gnd 0.201303f
C1533 CSoutput.t154 gnd 0.049596f
C1534 CSoutput.t97 gnd 0.049596f
C1535 CSoutput.n365 gnd 0.438244f
C1536 CSoutput.n366 gnd 0.201303f
C1537 CSoutput.t105 gnd 0.049596f
C1538 CSoutput.t185 gnd 0.049596f
C1539 CSoutput.n367 gnd 0.438244f
C1540 CSoutput.n368 gnd 0.201303f
C1541 CSoutput.t112 gnd 0.049596f
C1542 CSoutput.t119 gnd 0.049596f
C1543 CSoutput.n369 gnd 0.438244f
C1544 CSoutput.n370 gnd 0.305621f
C1545 CSoutput.n371 gnd 0.413948f
C1546 CSoutput.n372 gnd 13.2928f
C1547 CSoutput.t151 gnd 0.049596f
C1548 CSoutput.t102 gnd 0.049596f
C1549 CSoutput.n373 gnd 0.439711f
C1550 CSoutput.t134 gnd 0.049596f
C1551 CSoutput.t182 gnd 0.049596f
C1552 CSoutput.n374 gnd 0.438244f
C1553 CSoutput.n375 gnd 0.408362f
C1554 CSoutput.t104 gnd 0.049596f
C1555 CSoutput.t165 gnd 0.049596f
C1556 CSoutput.n376 gnd 0.438244f
C1557 CSoutput.n377 gnd 0.201303f
C1558 CSoutput.t164 gnd 0.049596f
C1559 CSoutput.t153 gnd 0.049596f
C1560 CSoutput.n378 gnd 0.438244f
C1561 CSoutput.n379 gnd 0.201303f
C1562 CSoutput.t168 gnd 0.049596f
C1563 CSoutput.t136 gnd 0.049596f
C1564 CSoutput.n380 gnd 0.438244f
C1565 CSoutput.n381 gnd 0.201303f
C1566 CSoutput.t160 gnd 0.049596f
C1567 CSoutput.t176 gnd 0.049596f
C1568 CSoutput.n382 gnd 0.438244f
C1569 CSoutput.n383 gnd 0.201303f
C1570 CSoutput.t190 gnd 0.049596f
C1571 CSoutput.t167 gnd 0.049596f
C1572 CSoutput.n384 gnd 0.438244f
C1573 CSoutput.n385 gnd 0.201303f
C1574 CSoutput.t172 gnd 0.049596f
C1575 CSoutput.t171 gnd 0.049596f
C1576 CSoutput.n386 gnd 0.438244f
C1577 CSoutput.n387 gnd 0.371292f
C1578 CSoutput.t137 gnd 0.049596f
C1579 CSoutput.t155 gnd 0.049596f
C1580 CSoutput.n388 gnd 0.439711f
C1581 CSoutput.t156 gnd 0.049596f
C1582 CSoutput.t146 gnd 0.049596f
C1583 CSoutput.n389 gnd 0.438244f
C1584 CSoutput.n390 gnd 0.408362f
C1585 CSoutput.t147 gnd 0.049596f
C1586 CSoutput.t138 gnd 0.049596f
C1587 CSoutput.n391 gnd 0.438244f
C1588 CSoutput.n392 gnd 0.201303f
C1589 CSoutput.t133 gnd 0.049596f
C1590 CSoutput.t125 gnd 0.049596f
C1591 CSoutput.n393 gnd 0.438244f
C1592 CSoutput.n394 gnd 0.201303f
C1593 CSoutput.t126 gnd 0.049596f
C1594 CSoutput.t148 gnd 0.049596f
C1595 CSoutput.n395 gnd 0.438244f
C1596 CSoutput.n396 gnd 0.201303f
C1597 CSoutput.t150 gnd 0.049596f
C1598 CSoutput.t99 gnd 0.049596f
C1599 CSoutput.n397 gnd 0.438244f
C1600 CSoutput.n398 gnd 0.201303f
C1601 CSoutput.t100 gnd 0.049596f
C1602 CSoutput.t118 gnd 0.049596f
C1603 CSoutput.n399 gnd 0.438244f
C1604 CSoutput.n400 gnd 0.201303f
C1605 CSoutput.t124 gnd 0.049596f
C1606 CSoutput.t113 gnd 0.049596f
C1607 CSoutput.n401 gnd 0.438244f
C1608 CSoutput.n402 gnd 0.305621f
C1609 CSoutput.n403 gnd 0.385483f
C1610 CSoutput.t169 gnd 0.049596f
C1611 CSoutput.t184 gnd 0.049596f
C1612 CSoutput.n404 gnd 0.439711f
C1613 CSoutput.t189 gnd 0.049596f
C1614 CSoutput.t158 gnd 0.049596f
C1615 CSoutput.n405 gnd 0.438244f
C1616 CSoutput.n406 gnd 0.408362f
C1617 CSoutput.t162 gnd 0.049596f
C1618 CSoutput.t178 gnd 0.049596f
C1619 CSoutput.n407 gnd 0.438244f
C1620 CSoutput.n408 gnd 0.201303f
C1621 CSoutput.t110 gnd 0.049596f
C1622 CSoutput.t152 gnd 0.049596f
C1623 CSoutput.n409 gnd 0.438244f
C1624 CSoutput.n410 gnd 0.201303f
C1625 CSoutput.t157 gnd 0.049596f
C1626 CSoutput.t170 gnd 0.049596f
C1627 CSoutput.n411 gnd 0.438244f
C1628 CSoutput.n412 gnd 0.201303f
C1629 CSoutput.t179 gnd 0.049596f
C1630 CSoutput.t161 gnd 0.049596f
C1631 CSoutput.n413 gnd 0.438244f
C1632 CSoutput.n414 gnd 0.201303f
C1633 CSoutput.t166 gnd 0.049596f
C1634 CSoutput.t183 gnd 0.049596f
C1635 CSoutput.n415 gnd 0.438244f
C1636 CSoutput.n416 gnd 0.201303f
C1637 CSoutput.t111 gnd 0.049596f
C1638 CSoutput.t122 gnd 0.049596f
C1639 CSoutput.n417 gnd 0.438244f
C1640 CSoutput.n418 gnd 0.305621f
C1641 CSoutput.n419 gnd 0.413948f
C1642 CSoutput.n420 gnd 7.81733f
C1643 CSoutput.n421 gnd 13.9523f
C1644 vdd.t7 gnd 0.038532f
C1645 vdd.t3 gnd 0.038532f
C1646 vdd.n0 gnd 0.303904f
C1647 vdd.t259 gnd 0.038532f
C1648 vdd.t33 gnd 0.038532f
C1649 vdd.n1 gnd 0.303402f
C1650 vdd.n2 gnd 0.279795f
C1651 vdd.t42 gnd 0.038532f
C1652 vdd.t9 gnd 0.038532f
C1653 vdd.n3 gnd 0.303402f
C1654 vdd.n4 gnd 0.141503f
C1655 vdd.t11 gnd 0.038532f
C1656 vdd.t249 gnd 0.038532f
C1657 vdd.n5 gnd 0.303402f
C1658 vdd.n6 gnd 0.132774f
C1659 vdd.t263 gnd 0.038532f
C1660 vdd.t261 gnd 0.038532f
C1661 vdd.n7 gnd 0.303904f
C1662 vdd.t251 gnd 0.038532f
C1663 vdd.t5 gnd 0.038532f
C1664 vdd.n8 gnd 0.303402f
C1665 vdd.n9 gnd 0.279795f
C1666 vdd.t35 gnd 0.038532f
C1667 vdd.t257 gnd 0.038532f
C1668 vdd.n10 gnd 0.303402f
C1669 vdd.n11 gnd 0.141503f
C1670 vdd.t20 gnd 0.038532f
C1671 vdd.t37 gnd 0.038532f
C1672 vdd.n12 gnd 0.303402f
C1673 vdd.n13 gnd 0.132774f
C1674 vdd.n14 gnd 0.093869f
C1675 vdd.t252 gnd 0.021406f
C1676 vdd.t254 gnd 0.021406f
C1677 vdd.n15 gnd 0.197036f
C1678 vdd.t16 gnd 0.021406f
C1679 vdd.t14 gnd 0.021406f
C1680 vdd.n16 gnd 0.19646f
C1681 vdd.n17 gnd 0.341902f
C1682 vdd.t28 gnd 0.021406f
C1683 vdd.t43 gnd 0.021406f
C1684 vdd.n18 gnd 0.19646f
C1685 vdd.n19 gnd 0.141449f
C1686 vdd.t17 gnd 0.021406f
C1687 vdd.t255 gnd 0.021406f
C1688 vdd.n20 gnd 0.197036f
C1689 vdd.t253 gnd 0.021406f
C1690 vdd.t30 gnd 0.021406f
C1691 vdd.n21 gnd 0.19646f
C1692 vdd.n22 gnd 0.341902f
C1693 vdd.t26 gnd 0.021406f
C1694 vdd.t29 gnd 0.021406f
C1695 vdd.n23 gnd 0.19646f
C1696 vdd.n24 gnd 0.141449f
C1697 vdd.t15 gnd 0.021406f
C1698 vdd.t24 gnd 0.021406f
C1699 vdd.n25 gnd 0.19646f
C1700 vdd.t40 gnd 0.021406f
C1701 vdd.t27 gnd 0.021406f
C1702 vdd.n26 gnd 0.19646f
C1703 vdd.n27 gnd 21.7441f
C1704 vdd.n28 gnd 8.33022f
C1705 vdd.n29 gnd 0.005838f
C1706 vdd.n30 gnd 0.005418f
C1707 vdd.n31 gnd 0.002997f
C1708 vdd.n32 gnd 0.006881f
C1709 vdd.n33 gnd 0.002911f
C1710 vdd.n34 gnd 0.003083f
C1711 vdd.n35 gnd 0.005418f
C1712 vdd.n36 gnd 0.002911f
C1713 vdd.n37 gnd 0.006881f
C1714 vdd.n38 gnd 0.003083f
C1715 vdd.n39 gnd 0.005418f
C1716 vdd.n40 gnd 0.002911f
C1717 vdd.n41 gnd 0.005161f
C1718 vdd.n42 gnd 0.005176f
C1719 vdd.t47 gnd 0.014784f
C1720 vdd.n43 gnd 0.032893f
C1721 vdd.n44 gnd 0.171185f
C1722 vdd.n45 gnd 0.002911f
C1723 vdd.n46 gnd 0.003083f
C1724 vdd.n47 gnd 0.006881f
C1725 vdd.n48 gnd 0.006881f
C1726 vdd.n49 gnd 0.003083f
C1727 vdd.n50 gnd 0.002911f
C1728 vdd.n51 gnd 0.005418f
C1729 vdd.n52 gnd 0.005418f
C1730 vdd.n53 gnd 0.002911f
C1731 vdd.n54 gnd 0.003083f
C1732 vdd.n55 gnd 0.006881f
C1733 vdd.n56 gnd 0.006881f
C1734 vdd.n57 gnd 0.003083f
C1735 vdd.n58 gnd 0.002911f
C1736 vdd.n59 gnd 0.005418f
C1737 vdd.n60 gnd 0.005418f
C1738 vdd.n61 gnd 0.002911f
C1739 vdd.n62 gnd 0.003083f
C1740 vdd.n63 gnd 0.006881f
C1741 vdd.n64 gnd 0.006881f
C1742 vdd.n65 gnd 0.016268f
C1743 vdd.n66 gnd 0.002997f
C1744 vdd.n67 gnd 0.002911f
C1745 vdd.n68 gnd 0.014003f
C1746 vdd.n69 gnd 0.009776f
C1747 vdd.t157 gnd 0.03425f
C1748 vdd.t108 gnd 0.03425f
C1749 vdd.n70 gnd 0.235391f
C1750 vdd.n71 gnd 0.185099f
C1751 vdd.t169 gnd 0.03425f
C1752 vdd.t80 gnd 0.03425f
C1753 vdd.n72 gnd 0.235391f
C1754 vdd.n73 gnd 0.149374f
C1755 vdd.t146 gnd 0.03425f
C1756 vdd.t100 gnd 0.03425f
C1757 vdd.n74 gnd 0.235391f
C1758 vdd.n75 gnd 0.149374f
C1759 vdd.t164 gnd 0.03425f
C1760 vdd.t143 gnd 0.03425f
C1761 vdd.n76 gnd 0.235391f
C1762 vdd.n77 gnd 0.149374f
C1763 vdd.t55 gnd 0.03425f
C1764 vdd.t93 gnd 0.03425f
C1765 vdd.n78 gnd 0.235391f
C1766 vdd.n79 gnd 0.149374f
C1767 vdd.t65 gnd 0.03425f
C1768 vdd.t111 gnd 0.03425f
C1769 vdd.n80 gnd 0.235391f
C1770 vdd.n81 gnd 0.149374f
C1771 vdd.t88 gnd 0.03425f
C1772 vdd.t153 gnd 0.03425f
C1773 vdd.n82 gnd 0.235391f
C1774 vdd.n83 gnd 0.149374f
C1775 vdd.n84 gnd 0.005838f
C1776 vdd.n85 gnd 0.005418f
C1777 vdd.n86 gnd 0.002997f
C1778 vdd.n87 gnd 0.006881f
C1779 vdd.n88 gnd 0.002911f
C1780 vdd.n89 gnd 0.003083f
C1781 vdd.n90 gnd 0.005418f
C1782 vdd.n91 gnd 0.002911f
C1783 vdd.n92 gnd 0.006881f
C1784 vdd.n93 gnd 0.003083f
C1785 vdd.n94 gnd 0.005418f
C1786 vdd.n95 gnd 0.002911f
C1787 vdd.n96 gnd 0.005161f
C1788 vdd.n97 gnd 0.005176f
C1789 vdd.t70 gnd 0.014784f
C1790 vdd.n98 gnd 0.032893f
C1791 vdd.n99 gnd 0.171185f
C1792 vdd.n100 gnd 0.002911f
C1793 vdd.n101 gnd 0.003083f
C1794 vdd.n102 gnd 0.006881f
C1795 vdd.n103 gnd 0.006881f
C1796 vdd.n104 gnd 0.003083f
C1797 vdd.n105 gnd 0.002911f
C1798 vdd.n106 gnd 0.005418f
C1799 vdd.n107 gnd 0.005418f
C1800 vdd.n108 gnd 0.002911f
C1801 vdd.n109 gnd 0.003083f
C1802 vdd.n110 gnd 0.006881f
C1803 vdd.n111 gnd 0.006881f
C1804 vdd.n112 gnd 0.003083f
C1805 vdd.n113 gnd 0.002911f
C1806 vdd.n114 gnd 0.005418f
C1807 vdd.n115 gnd 0.005418f
C1808 vdd.n116 gnd 0.002911f
C1809 vdd.n117 gnd 0.003083f
C1810 vdd.n118 gnd 0.006881f
C1811 vdd.n119 gnd 0.006881f
C1812 vdd.n120 gnd 0.016268f
C1813 vdd.n121 gnd 0.002997f
C1814 vdd.n122 gnd 0.002911f
C1815 vdd.n123 gnd 0.014003f
C1816 vdd.n124 gnd 0.00947f
C1817 vdd.n125 gnd 0.111135f
C1818 vdd.n126 gnd 0.005838f
C1819 vdd.n127 gnd 0.005418f
C1820 vdd.n128 gnd 0.002997f
C1821 vdd.n129 gnd 0.006881f
C1822 vdd.n130 gnd 0.002911f
C1823 vdd.n131 gnd 0.003083f
C1824 vdd.n132 gnd 0.005418f
C1825 vdd.n133 gnd 0.002911f
C1826 vdd.n134 gnd 0.006881f
C1827 vdd.n135 gnd 0.003083f
C1828 vdd.n136 gnd 0.005418f
C1829 vdd.n137 gnd 0.002911f
C1830 vdd.n138 gnd 0.005161f
C1831 vdd.n139 gnd 0.005176f
C1832 vdd.t113 gnd 0.014784f
C1833 vdd.n140 gnd 0.032893f
C1834 vdd.n141 gnd 0.171185f
C1835 vdd.n142 gnd 0.002911f
C1836 vdd.n143 gnd 0.003083f
C1837 vdd.n144 gnd 0.006881f
C1838 vdd.n145 gnd 0.006881f
C1839 vdd.n146 gnd 0.003083f
C1840 vdd.n147 gnd 0.002911f
C1841 vdd.n148 gnd 0.005418f
C1842 vdd.n149 gnd 0.005418f
C1843 vdd.n150 gnd 0.002911f
C1844 vdd.n151 gnd 0.003083f
C1845 vdd.n152 gnd 0.006881f
C1846 vdd.n153 gnd 0.006881f
C1847 vdd.n154 gnd 0.003083f
C1848 vdd.n155 gnd 0.002911f
C1849 vdd.n156 gnd 0.005418f
C1850 vdd.n157 gnd 0.005418f
C1851 vdd.n158 gnd 0.002911f
C1852 vdd.n159 gnd 0.003083f
C1853 vdd.n160 gnd 0.006881f
C1854 vdd.n161 gnd 0.006881f
C1855 vdd.n162 gnd 0.016268f
C1856 vdd.n163 gnd 0.002997f
C1857 vdd.n164 gnd 0.002911f
C1858 vdd.n165 gnd 0.014003f
C1859 vdd.n166 gnd 0.009776f
C1860 vdd.t115 gnd 0.03425f
C1861 vdd.t139 gnd 0.03425f
C1862 vdd.n167 gnd 0.235391f
C1863 vdd.n168 gnd 0.185099f
C1864 vdd.t53 gnd 0.03425f
C1865 vdd.t101 gnd 0.03425f
C1866 vdd.n169 gnd 0.235391f
C1867 vdd.n170 gnd 0.149374f
C1868 vdd.t136 gnd 0.03425f
C1869 vdd.t45 gnd 0.03425f
C1870 vdd.n171 gnd 0.235391f
C1871 vdd.n172 gnd 0.149374f
C1872 vdd.t90 gnd 0.03425f
C1873 vdd.t92 gnd 0.03425f
C1874 vdd.n173 gnd 0.235391f
C1875 vdd.n174 gnd 0.149374f
C1876 vdd.t159 gnd 0.03425f
C1877 vdd.t85 gnd 0.03425f
C1878 vdd.n175 gnd 0.235391f
C1879 vdd.n176 gnd 0.149374f
C1880 vdd.t86 gnd 0.03425f
C1881 vdd.t155 gnd 0.03425f
C1882 vdd.n177 gnd 0.235391f
C1883 vdd.n178 gnd 0.149374f
C1884 vdd.t156 gnd 0.03425f
C1885 vdd.t63 gnd 0.03425f
C1886 vdd.n179 gnd 0.235391f
C1887 vdd.n180 gnd 0.149374f
C1888 vdd.n181 gnd 0.005838f
C1889 vdd.n182 gnd 0.005418f
C1890 vdd.n183 gnd 0.002997f
C1891 vdd.n184 gnd 0.006881f
C1892 vdd.n185 gnd 0.002911f
C1893 vdd.n186 gnd 0.003083f
C1894 vdd.n187 gnd 0.005418f
C1895 vdd.n188 gnd 0.002911f
C1896 vdd.n189 gnd 0.006881f
C1897 vdd.n190 gnd 0.003083f
C1898 vdd.n191 gnd 0.005418f
C1899 vdd.n192 gnd 0.002911f
C1900 vdd.n193 gnd 0.005161f
C1901 vdd.n194 gnd 0.005176f
C1902 vdd.t137 gnd 0.014784f
C1903 vdd.n195 gnd 0.032893f
C1904 vdd.n196 gnd 0.171185f
C1905 vdd.n197 gnd 0.002911f
C1906 vdd.n198 gnd 0.003083f
C1907 vdd.n199 gnd 0.006881f
C1908 vdd.n200 gnd 0.006881f
C1909 vdd.n201 gnd 0.003083f
C1910 vdd.n202 gnd 0.002911f
C1911 vdd.n203 gnd 0.005418f
C1912 vdd.n204 gnd 0.005418f
C1913 vdd.n205 gnd 0.002911f
C1914 vdd.n206 gnd 0.003083f
C1915 vdd.n207 gnd 0.006881f
C1916 vdd.n208 gnd 0.006881f
C1917 vdd.n209 gnd 0.003083f
C1918 vdd.n210 gnd 0.002911f
C1919 vdd.n211 gnd 0.005418f
C1920 vdd.n212 gnd 0.005418f
C1921 vdd.n213 gnd 0.002911f
C1922 vdd.n214 gnd 0.003083f
C1923 vdd.n215 gnd 0.006881f
C1924 vdd.n216 gnd 0.006881f
C1925 vdd.n217 gnd 0.016268f
C1926 vdd.n218 gnd 0.002997f
C1927 vdd.n219 gnd 0.002911f
C1928 vdd.n220 gnd 0.014003f
C1929 vdd.n221 gnd 0.00947f
C1930 vdd.n222 gnd 0.066114f
C1931 vdd.n223 gnd 0.238226f
C1932 vdd.n224 gnd 0.005838f
C1933 vdd.n225 gnd 0.005418f
C1934 vdd.n226 gnd 0.002997f
C1935 vdd.n227 gnd 0.006881f
C1936 vdd.n228 gnd 0.002911f
C1937 vdd.n229 gnd 0.003083f
C1938 vdd.n230 gnd 0.005418f
C1939 vdd.n231 gnd 0.002911f
C1940 vdd.n232 gnd 0.006881f
C1941 vdd.n233 gnd 0.003083f
C1942 vdd.n234 gnd 0.005418f
C1943 vdd.n235 gnd 0.002911f
C1944 vdd.n236 gnd 0.005161f
C1945 vdd.n237 gnd 0.005176f
C1946 vdd.t125 gnd 0.014784f
C1947 vdd.n238 gnd 0.032893f
C1948 vdd.n239 gnd 0.171185f
C1949 vdd.n240 gnd 0.002911f
C1950 vdd.n241 gnd 0.003083f
C1951 vdd.n242 gnd 0.006881f
C1952 vdd.n243 gnd 0.006881f
C1953 vdd.n244 gnd 0.003083f
C1954 vdd.n245 gnd 0.002911f
C1955 vdd.n246 gnd 0.005418f
C1956 vdd.n247 gnd 0.005418f
C1957 vdd.n248 gnd 0.002911f
C1958 vdd.n249 gnd 0.003083f
C1959 vdd.n250 gnd 0.006881f
C1960 vdd.n251 gnd 0.006881f
C1961 vdd.n252 gnd 0.003083f
C1962 vdd.n253 gnd 0.002911f
C1963 vdd.n254 gnd 0.005418f
C1964 vdd.n255 gnd 0.005418f
C1965 vdd.n256 gnd 0.002911f
C1966 vdd.n257 gnd 0.003083f
C1967 vdd.n258 gnd 0.006881f
C1968 vdd.n259 gnd 0.006881f
C1969 vdd.n260 gnd 0.016268f
C1970 vdd.n261 gnd 0.002997f
C1971 vdd.n262 gnd 0.002911f
C1972 vdd.n263 gnd 0.014003f
C1973 vdd.n264 gnd 0.009776f
C1974 vdd.t127 gnd 0.03425f
C1975 vdd.t150 gnd 0.03425f
C1976 vdd.n265 gnd 0.235391f
C1977 vdd.n266 gnd 0.185099f
C1978 vdd.t75 gnd 0.03425f
C1979 vdd.t126 gnd 0.03425f
C1980 vdd.n267 gnd 0.235391f
C1981 vdd.n268 gnd 0.149374f
C1982 vdd.t122 gnd 0.03425f
C1983 vdd.t68 gnd 0.03425f
C1984 vdd.n269 gnd 0.235391f
C1985 vdd.n270 gnd 0.149374f
C1986 vdd.t104 gnd 0.03425f
C1987 vdd.t106 gnd 0.03425f
C1988 vdd.n271 gnd 0.235391f
C1989 vdd.n272 gnd 0.149374f
C1990 vdd.t166 gnd 0.03425f
C1991 vdd.t98 gnd 0.03425f
C1992 vdd.n273 gnd 0.235391f
C1993 vdd.n274 gnd 0.149374f
C1994 vdd.t99 gnd 0.03425f
C1995 vdd.t167 gnd 0.03425f
C1996 vdd.n275 gnd 0.235391f
C1997 vdd.n276 gnd 0.149374f
C1998 vdd.t168 gnd 0.03425f
C1999 vdd.t78 gnd 0.03425f
C2000 vdd.n277 gnd 0.235391f
C2001 vdd.n278 gnd 0.149374f
C2002 vdd.n279 gnd 0.005838f
C2003 vdd.n280 gnd 0.005418f
C2004 vdd.n281 gnd 0.002997f
C2005 vdd.n282 gnd 0.006881f
C2006 vdd.n283 gnd 0.002911f
C2007 vdd.n284 gnd 0.003083f
C2008 vdd.n285 gnd 0.005418f
C2009 vdd.n286 gnd 0.002911f
C2010 vdd.n287 gnd 0.006881f
C2011 vdd.n288 gnd 0.003083f
C2012 vdd.n289 gnd 0.005418f
C2013 vdd.n290 gnd 0.002911f
C2014 vdd.n291 gnd 0.005161f
C2015 vdd.n292 gnd 0.005176f
C2016 vdd.t148 gnd 0.014784f
C2017 vdd.n293 gnd 0.032893f
C2018 vdd.n294 gnd 0.171185f
C2019 vdd.n295 gnd 0.002911f
C2020 vdd.n296 gnd 0.003083f
C2021 vdd.n297 gnd 0.006881f
C2022 vdd.n298 gnd 0.006881f
C2023 vdd.n299 gnd 0.003083f
C2024 vdd.n300 gnd 0.002911f
C2025 vdd.n301 gnd 0.005418f
C2026 vdd.n302 gnd 0.005418f
C2027 vdd.n303 gnd 0.002911f
C2028 vdd.n304 gnd 0.003083f
C2029 vdd.n305 gnd 0.006881f
C2030 vdd.n306 gnd 0.006881f
C2031 vdd.n307 gnd 0.003083f
C2032 vdd.n308 gnd 0.002911f
C2033 vdd.n309 gnd 0.005418f
C2034 vdd.n310 gnd 0.005418f
C2035 vdd.n311 gnd 0.002911f
C2036 vdd.n312 gnd 0.003083f
C2037 vdd.n313 gnd 0.006881f
C2038 vdd.n314 gnd 0.006881f
C2039 vdd.n315 gnd 0.016268f
C2040 vdd.n316 gnd 0.002997f
C2041 vdd.n317 gnd 0.002911f
C2042 vdd.n318 gnd 0.014003f
C2043 vdd.n319 gnd 0.00947f
C2044 vdd.n320 gnd 0.066114f
C2045 vdd.n321 gnd 0.266781f
C2046 vdd.n322 gnd 0.008176f
C2047 vdd.n323 gnd 0.010638f
C2048 vdd.n324 gnd 0.008563f
C2049 vdd.n325 gnd 0.008563f
C2050 vdd.n326 gnd 0.010638f
C2051 vdd.n327 gnd 0.010638f
C2052 vdd.n328 gnd 0.777336f
C2053 vdd.n329 gnd 0.010638f
C2054 vdd.n330 gnd 0.010638f
C2055 vdd.n331 gnd 0.010638f
C2056 vdd.n332 gnd 0.842567f
C2057 vdd.n333 gnd 0.010638f
C2058 vdd.n334 gnd 0.010638f
C2059 vdd.n335 gnd 0.010638f
C2060 vdd.n336 gnd 0.010638f
C2061 vdd.n337 gnd 0.008563f
C2062 vdd.n338 gnd 0.010638f
C2063 vdd.t84 gnd 0.543592f
C2064 vdd.n339 gnd 0.010638f
C2065 vdd.n340 gnd 0.010638f
C2066 vdd.n341 gnd 0.010638f
C2067 vdd.t110 gnd 0.543592f
C2068 vdd.n342 gnd 0.010638f
C2069 vdd.n343 gnd 0.010638f
C2070 vdd.n344 gnd 0.010638f
C2071 vdd.n345 gnd 0.010638f
C2072 vdd.n346 gnd 0.010638f
C2073 vdd.n347 gnd 0.008563f
C2074 vdd.n348 gnd 0.010638f
C2075 vdd.n349 gnd 0.614259f
C2076 vdd.n350 gnd 0.010638f
C2077 vdd.n351 gnd 0.010638f
C2078 vdd.n352 gnd 0.010638f
C2079 vdd.t62 gnd 0.543592f
C2080 vdd.n353 gnd 0.010638f
C2081 vdd.n354 gnd 0.010638f
C2082 vdd.n355 gnd 0.010638f
C2083 vdd.n356 gnd 0.010638f
C2084 vdd.n357 gnd 0.010638f
C2085 vdd.n358 gnd 0.008563f
C2086 vdd.n359 gnd 0.010638f
C2087 vdd.t69 gnd 0.543592f
C2088 vdd.n360 gnd 0.010638f
C2089 vdd.n361 gnd 0.010638f
C2090 vdd.n362 gnd 0.010638f
C2091 vdd.n363 gnd 0.91867f
C2092 vdd.n364 gnd 0.010638f
C2093 vdd.n365 gnd 0.010638f
C2094 vdd.n366 gnd 0.010638f
C2095 vdd.n367 gnd 0.010638f
C2096 vdd.n368 gnd 0.010638f
C2097 vdd.n369 gnd 0.007107f
C2098 vdd.n370 gnd 0.024226f
C2099 vdd.t181 gnd 0.543592f
C2100 vdd.n371 gnd 0.010638f
C2101 vdd.n372 gnd 0.024226f
C2102 vdd.n404 gnd 0.010638f
C2103 vdd.t183 gnd 0.130879f
C2104 vdd.t182 gnd 0.139874f
C2105 vdd.t180 gnd 0.170926f
C2106 vdd.n405 gnd 0.219103f
C2107 vdd.n406 gnd 0.184943f
C2108 vdd.n407 gnd 0.014043f
C2109 vdd.n408 gnd 0.010638f
C2110 vdd.n409 gnd 0.008563f
C2111 vdd.n410 gnd 0.010638f
C2112 vdd.n411 gnd 0.008563f
C2113 vdd.n412 gnd 0.010638f
C2114 vdd.n413 gnd 0.008563f
C2115 vdd.n414 gnd 0.010638f
C2116 vdd.n415 gnd 0.008563f
C2117 vdd.n416 gnd 0.010638f
C2118 vdd.n417 gnd 0.008563f
C2119 vdd.n418 gnd 0.010638f
C2120 vdd.t241 gnd 0.130879f
C2121 vdd.t240 gnd 0.139874f
C2122 vdd.t239 gnd 0.170926f
C2123 vdd.n419 gnd 0.219103f
C2124 vdd.n420 gnd 0.184943f
C2125 vdd.n421 gnd 0.008563f
C2126 vdd.n422 gnd 0.010638f
C2127 vdd.n423 gnd 0.008563f
C2128 vdd.n424 gnd 0.010638f
C2129 vdd.n425 gnd 0.008563f
C2130 vdd.n426 gnd 0.010638f
C2131 vdd.n427 gnd 0.008563f
C2132 vdd.n428 gnd 0.010638f
C2133 vdd.n429 gnd 0.008563f
C2134 vdd.n430 gnd 0.010638f
C2135 vdd.t247 gnd 0.130879f
C2136 vdd.t246 gnd 0.139874f
C2137 vdd.t245 gnd 0.170926f
C2138 vdd.n431 gnd 0.219103f
C2139 vdd.n432 gnd 0.184943f
C2140 vdd.n433 gnd 0.018324f
C2141 vdd.n434 gnd 0.010638f
C2142 vdd.n435 gnd 0.008563f
C2143 vdd.n436 gnd 0.010638f
C2144 vdd.n437 gnd 0.008563f
C2145 vdd.n438 gnd 0.010638f
C2146 vdd.n439 gnd 0.008563f
C2147 vdd.n440 gnd 0.010638f
C2148 vdd.n441 gnd 0.008563f
C2149 vdd.n442 gnd 0.010638f
C2150 vdd.n443 gnd 0.024226f
C2151 vdd.n444 gnd 0.024391f
C2152 vdd.n445 gnd 0.024391f
C2153 vdd.n446 gnd 0.007107f
C2154 vdd.n447 gnd 0.008563f
C2155 vdd.n448 gnd 0.010638f
C2156 vdd.n449 gnd 0.010638f
C2157 vdd.n450 gnd 0.008563f
C2158 vdd.n451 gnd 0.010638f
C2159 vdd.n452 gnd 0.010638f
C2160 vdd.n453 gnd 0.010638f
C2161 vdd.n454 gnd 0.010638f
C2162 vdd.n455 gnd 0.010638f
C2163 vdd.n456 gnd 0.008563f
C2164 vdd.n457 gnd 0.008563f
C2165 vdd.n458 gnd 0.010638f
C2166 vdd.n459 gnd 0.010638f
C2167 vdd.n460 gnd 0.008563f
C2168 vdd.n461 gnd 0.010638f
C2169 vdd.n462 gnd 0.010638f
C2170 vdd.n463 gnd 0.010638f
C2171 vdd.n464 gnd 0.010638f
C2172 vdd.n465 gnd 0.010638f
C2173 vdd.n466 gnd 0.008563f
C2174 vdd.n467 gnd 0.008563f
C2175 vdd.n468 gnd 0.010638f
C2176 vdd.n469 gnd 0.010638f
C2177 vdd.n470 gnd 0.008563f
C2178 vdd.n471 gnd 0.010638f
C2179 vdd.n472 gnd 0.010638f
C2180 vdd.n473 gnd 0.010638f
C2181 vdd.n474 gnd 0.010638f
C2182 vdd.n475 gnd 0.010638f
C2183 vdd.n476 gnd 0.008563f
C2184 vdd.n477 gnd 0.008563f
C2185 vdd.n478 gnd 0.010638f
C2186 vdd.n479 gnd 0.010638f
C2187 vdd.n480 gnd 0.008563f
C2188 vdd.n481 gnd 0.010638f
C2189 vdd.n482 gnd 0.010638f
C2190 vdd.n483 gnd 0.010638f
C2191 vdd.n484 gnd 0.010638f
C2192 vdd.n485 gnd 0.010638f
C2193 vdd.n486 gnd 0.008563f
C2194 vdd.n487 gnd 0.008563f
C2195 vdd.n488 gnd 0.010638f
C2196 vdd.n489 gnd 0.010638f
C2197 vdd.n490 gnd 0.00715f
C2198 vdd.n491 gnd 0.010638f
C2199 vdd.n492 gnd 0.010638f
C2200 vdd.n493 gnd 0.010638f
C2201 vdd.n494 gnd 0.010638f
C2202 vdd.n495 gnd 0.010638f
C2203 vdd.n496 gnd 0.00715f
C2204 vdd.n497 gnd 0.008563f
C2205 vdd.n498 gnd 0.010638f
C2206 vdd.n499 gnd 0.010638f
C2207 vdd.n500 gnd 0.008563f
C2208 vdd.n501 gnd 0.010638f
C2209 vdd.n502 gnd 0.010638f
C2210 vdd.n503 gnd 0.010638f
C2211 vdd.n504 gnd 0.010638f
C2212 vdd.n505 gnd 0.010638f
C2213 vdd.n506 gnd 0.008563f
C2214 vdd.n507 gnd 0.008563f
C2215 vdd.n508 gnd 0.010638f
C2216 vdd.n509 gnd 0.010638f
C2217 vdd.n510 gnd 0.008563f
C2218 vdd.n511 gnd 0.010638f
C2219 vdd.n512 gnd 0.010638f
C2220 vdd.n513 gnd 0.010638f
C2221 vdd.n514 gnd 0.010638f
C2222 vdd.n515 gnd 0.010638f
C2223 vdd.n516 gnd 0.008563f
C2224 vdd.n517 gnd 0.008563f
C2225 vdd.n518 gnd 0.010638f
C2226 vdd.n519 gnd 0.010638f
C2227 vdd.n520 gnd 0.008563f
C2228 vdd.n521 gnd 0.010638f
C2229 vdd.n522 gnd 0.010638f
C2230 vdd.n523 gnd 0.010638f
C2231 vdd.n524 gnd 0.010638f
C2232 vdd.n525 gnd 0.010638f
C2233 vdd.n526 gnd 0.008563f
C2234 vdd.n527 gnd 0.008563f
C2235 vdd.n528 gnd 0.010638f
C2236 vdd.n529 gnd 0.010638f
C2237 vdd.n530 gnd 0.008563f
C2238 vdd.n531 gnd 0.010638f
C2239 vdd.n532 gnd 0.010638f
C2240 vdd.n533 gnd 0.010638f
C2241 vdd.n534 gnd 0.010638f
C2242 vdd.n535 gnd 0.010638f
C2243 vdd.n536 gnd 0.008563f
C2244 vdd.n537 gnd 0.008563f
C2245 vdd.n538 gnd 0.010638f
C2246 vdd.n539 gnd 0.010638f
C2247 vdd.n540 gnd 0.008563f
C2248 vdd.n541 gnd 0.010638f
C2249 vdd.n542 gnd 0.010638f
C2250 vdd.n543 gnd 0.010638f
C2251 vdd.n544 gnd 0.010638f
C2252 vdd.n545 gnd 0.010638f
C2253 vdd.n546 gnd 0.005823f
C2254 vdd.n547 gnd 0.018324f
C2255 vdd.n548 gnd 0.010638f
C2256 vdd.n549 gnd 0.010638f
C2257 vdd.n550 gnd 0.008477f
C2258 vdd.n551 gnd 0.010638f
C2259 vdd.n552 gnd 0.010638f
C2260 vdd.n553 gnd 0.010638f
C2261 vdd.n554 gnd 0.010638f
C2262 vdd.n555 gnd 0.010638f
C2263 vdd.n556 gnd 0.008563f
C2264 vdd.n557 gnd 0.008563f
C2265 vdd.n558 gnd 0.010638f
C2266 vdd.n559 gnd 0.010638f
C2267 vdd.n560 gnd 0.008563f
C2268 vdd.n561 gnd 0.010638f
C2269 vdd.n562 gnd 0.010638f
C2270 vdd.n563 gnd 0.010638f
C2271 vdd.n564 gnd 0.010638f
C2272 vdd.n565 gnd 0.010638f
C2273 vdd.n566 gnd 0.008563f
C2274 vdd.n567 gnd 0.008563f
C2275 vdd.n568 gnd 0.010638f
C2276 vdd.n569 gnd 0.010638f
C2277 vdd.n570 gnd 0.008563f
C2278 vdd.n571 gnd 0.010638f
C2279 vdd.n572 gnd 0.010638f
C2280 vdd.n573 gnd 0.010638f
C2281 vdd.n574 gnd 0.010638f
C2282 vdd.n575 gnd 0.010638f
C2283 vdd.n576 gnd 0.008563f
C2284 vdd.n577 gnd 0.008563f
C2285 vdd.n578 gnd 0.010638f
C2286 vdd.n579 gnd 0.010638f
C2287 vdd.n580 gnd 0.008563f
C2288 vdd.n581 gnd 0.010638f
C2289 vdd.n582 gnd 0.010638f
C2290 vdd.n583 gnd 0.010638f
C2291 vdd.n584 gnd 0.010638f
C2292 vdd.n585 gnd 0.010638f
C2293 vdd.n586 gnd 0.008563f
C2294 vdd.n587 gnd 0.008563f
C2295 vdd.n588 gnd 0.010638f
C2296 vdd.n589 gnd 0.010638f
C2297 vdd.n590 gnd 0.008563f
C2298 vdd.n591 gnd 0.010638f
C2299 vdd.n592 gnd 0.010638f
C2300 vdd.n593 gnd 0.010638f
C2301 vdd.n594 gnd 0.010638f
C2302 vdd.n595 gnd 0.010638f
C2303 vdd.n596 gnd 0.008563f
C2304 vdd.n597 gnd 0.010638f
C2305 vdd.n598 gnd 0.008563f
C2306 vdd.n599 gnd 0.004495f
C2307 vdd.n600 gnd 0.010638f
C2308 vdd.n601 gnd 0.010638f
C2309 vdd.n602 gnd 0.008563f
C2310 vdd.n603 gnd 0.010638f
C2311 vdd.n604 gnd 0.008563f
C2312 vdd.n605 gnd 0.010638f
C2313 vdd.n606 gnd 0.008563f
C2314 vdd.n607 gnd 0.010638f
C2315 vdd.n608 gnd 0.008563f
C2316 vdd.n609 gnd 0.010638f
C2317 vdd.n610 gnd 0.008563f
C2318 vdd.n611 gnd 0.010638f
C2319 vdd.n612 gnd 0.010638f
C2320 vdd.n613 gnd 0.592515f
C2321 vdd.t89 gnd 0.543592f
C2322 vdd.n614 gnd 0.010638f
C2323 vdd.n615 gnd 0.008563f
C2324 vdd.n616 gnd 0.010638f
C2325 vdd.n617 gnd 0.008563f
C2326 vdd.n618 gnd 0.010638f
C2327 vdd.t121 gnd 0.543592f
C2328 vdd.n619 gnd 0.010638f
C2329 vdd.n620 gnd 0.008563f
C2330 vdd.n621 gnd 0.010638f
C2331 vdd.n622 gnd 0.008563f
C2332 vdd.n623 gnd 0.010638f
C2333 vdd.t79 gnd 0.543592f
C2334 vdd.n624 gnd 0.67949f
C2335 vdd.n625 gnd 0.010638f
C2336 vdd.n626 gnd 0.008563f
C2337 vdd.n627 gnd 0.010638f
C2338 vdd.n628 gnd 0.008563f
C2339 vdd.n629 gnd 0.010638f
C2340 vdd.t52 gnd 0.543592f
C2341 vdd.n630 gnd 0.010638f
C2342 vdd.n631 gnd 0.008563f
C2343 vdd.n632 gnd 0.010638f
C2344 vdd.n633 gnd 0.008563f
C2345 vdd.n634 gnd 0.010638f
C2346 vdd.n635 gnd 0.755593f
C2347 vdd.n636 gnd 0.902362f
C2348 vdd.t107 gnd 0.543592f
C2349 vdd.n637 gnd 0.010638f
C2350 vdd.n638 gnd 0.008563f
C2351 vdd.n639 gnd 0.010638f
C2352 vdd.n640 gnd 0.008563f
C2353 vdd.n641 gnd 0.010638f
C2354 vdd.n642 gnd 0.570771f
C2355 vdd.n643 gnd 0.010638f
C2356 vdd.n644 gnd 0.008563f
C2357 vdd.n645 gnd 0.010638f
C2358 vdd.n646 gnd 0.008563f
C2359 vdd.n647 gnd 0.010638f
C2360 vdd.n648 gnd 1.08718f
C2361 vdd.t46 gnd 0.543592f
C2362 vdd.n649 gnd 0.010638f
C2363 vdd.n650 gnd 0.008563f
C2364 vdd.n651 gnd 0.010638f
C2365 vdd.n652 gnd 0.008563f
C2366 vdd.n653 gnd 0.010638f
C2367 vdd.t177 gnd 0.543592f
C2368 vdd.n654 gnd 0.010638f
C2369 vdd.n655 gnd 0.008563f
C2370 vdd.n656 gnd 0.024391f
C2371 vdd.n657 gnd 0.024391f
C2372 vdd.n658 gnd 7.68639f
C2373 vdd.n659 gnd 0.603387f
C2374 vdd.n660 gnd 0.024391f
C2375 vdd.n661 gnd 0.009149f
C2376 vdd.n662 gnd 0.008563f
C2377 vdd.n667 gnd 0.006809f
C2378 vdd.n668 gnd 0.008563f
C2379 vdd.n669 gnd 0.010638f
C2380 vdd.n670 gnd 0.010638f
C2381 vdd.n671 gnd 0.010638f
C2382 vdd.n672 gnd 0.010638f
C2383 vdd.n673 gnd 0.010638f
C2384 vdd.n674 gnd 0.008563f
C2385 vdd.n675 gnd 0.010638f
C2386 vdd.n676 gnd 0.010638f
C2387 vdd.n677 gnd 0.010638f
C2388 vdd.n678 gnd 0.010638f
C2389 vdd.n679 gnd 0.010638f
C2390 vdd.n680 gnd 0.008563f
C2391 vdd.n681 gnd 0.010638f
C2392 vdd.n682 gnd 0.010638f
C2393 vdd.n683 gnd 0.010638f
C2394 vdd.n684 gnd 0.010638f
C2395 vdd.n685 gnd 0.010638f
C2396 vdd.t189 gnd 0.130879f
C2397 vdd.t190 gnd 0.139874f
C2398 vdd.t188 gnd 0.170926f
C2399 vdd.n686 gnd 0.219103f
C2400 vdd.n687 gnd 0.184086f
C2401 vdd.n688 gnd 0.017468f
C2402 vdd.n689 gnd 0.010638f
C2403 vdd.n690 gnd 0.010638f
C2404 vdd.n691 gnd 0.010638f
C2405 vdd.n692 gnd 0.010638f
C2406 vdd.n693 gnd 0.010638f
C2407 vdd.n694 gnd 0.008563f
C2408 vdd.n695 gnd 0.010638f
C2409 vdd.n696 gnd 0.010638f
C2410 vdd.n697 gnd 0.010638f
C2411 vdd.n698 gnd 0.010638f
C2412 vdd.n699 gnd 0.010638f
C2413 vdd.n700 gnd 0.008563f
C2414 vdd.n701 gnd 0.010638f
C2415 vdd.n702 gnd 0.010638f
C2416 vdd.n703 gnd 0.010638f
C2417 vdd.n704 gnd 0.010638f
C2418 vdd.n705 gnd 0.010638f
C2419 vdd.n706 gnd 0.008563f
C2420 vdd.n707 gnd 0.010638f
C2421 vdd.n708 gnd 0.010638f
C2422 vdd.n709 gnd 0.010638f
C2423 vdd.n710 gnd 0.010638f
C2424 vdd.n711 gnd 0.010638f
C2425 vdd.n712 gnd 0.008563f
C2426 vdd.n713 gnd 0.010638f
C2427 vdd.n714 gnd 0.010638f
C2428 vdd.n715 gnd 0.010638f
C2429 vdd.n716 gnd 0.010638f
C2430 vdd.n717 gnd 0.010638f
C2431 vdd.n718 gnd 0.008563f
C2432 vdd.n719 gnd 0.010638f
C2433 vdd.n720 gnd 0.010638f
C2434 vdd.n721 gnd 0.010638f
C2435 vdd.n722 gnd 0.008477f
C2436 vdd.t178 gnd 0.130879f
C2437 vdd.t179 gnd 0.139874f
C2438 vdd.t176 gnd 0.170926f
C2439 vdd.n723 gnd 0.219103f
C2440 vdd.n724 gnd 0.184086f
C2441 vdd.n725 gnd 0.010638f
C2442 vdd.n726 gnd 0.008563f
C2443 vdd.n728 gnd 0.010638f
C2444 vdd.n730 gnd 0.010638f
C2445 vdd.n731 gnd 0.010638f
C2446 vdd.n732 gnd 0.008563f
C2447 vdd.n733 gnd 0.010638f
C2448 vdd.n734 gnd 0.010638f
C2449 vdd.n735 gnd 0.010638f
C2450 vdd.n736 gnd 0.010638f
C2451 vdd.n737 gnd 0.010638f
C2452 vdd.n738 gnd 0.008563f
C2453 vdd.n739 gnd 0.010638f
C2454 vdd.n740 gnd 0.010638f
C2455 vdd.n741 gnd 0.010638f
C2456 vdd.n742 gnd 0.010638f
C2457 vdd.n743 gnd 0.010638f
C2458 vdd.n744 gnd 0.008563f
C2459 vdd.n745 gnd 0.010638f
C2460 vdd.n746 gnd 0.010638f
C2461 vdd.n747 gnd 0.010638f
C2462 vdd.n748 gnd 0.006809f
C2463 vdd.n753 gnd 0.007234f
C2464 vdd.n754 gnd 0.007234f
C2465 vdd.n755 gnd 0.007234f
C2466 vdd.n756 gnd 7.4907f
C2467 vdd.n757 gnd 0.007234f
C2468 vdd.n758 gnd 0.007234f
C2469 vdd.n759 gnd 0.007234f
C2470 vdd.n761 gnd 0.007234f
C2471 vdd.n762 gnd 0.007234f
C2472 vdd.n764 gnd 0.007234f
C2473 vdd.n765 gnd 0.005266f
C2474 vdd.n767 gnd 0.007234f
C2475 vdd.t225 gnd 0.292327f
C2476 vdd.t224 gnd 0.299233f
C2477 vdd.t223 gnd 0.190842f
C2478 vdd.n768 gnd 0.10314f
C2479 vdd.n769 gnd 0.058504f
C2480 vdd.n770 gnd 0.010339f
C2481 vdd.n771 gnd 0.016907f
C2482 vdd.n773 gnd 0.007234f
C2483 vdd.n774 gnd 0.739285f
C2484 vdd.n775 gnd 0.016026f
C2485 vdd.n776 gnd 0.016026f
C2486 vdd.n777 gnd 0.007234f
C2487 vdd.n778 gnd 0.017165f
C2488 vdd.n779 gnd 0.007234f
C2489 vdd.n780 gnd 0.007234f
C2490 vdd.n781 gnd 0.007234f
C2491 vdd.n782 gnd 0.007234f
C2492 vdd.n783 gnd 0.007234f
C2493 vdd.n785 gnd 0.007234f
C2494 vdd.n786 gnd 0.007234f
C2495 vdd.n788 gnd 0.007234f
C2496 vdd.n789 gnd 0.007234f
C2497 vdd.n791 gnd 0.007234f
C2498 vdd.n792 gnd 0.007234f
C2499 vdd.n794 gnd 0.007234f
C2500 vdd.n795 gnd 0.007234f
C2501 vdd.n797 gnd 0.007234f
C2502 vdd.n798 gnd 0.007234f
C2503 vdd.n800 gnd 0.007234f
C2504 vdd.n801 gnd 0.005266f
C2505 vdd.n803 gnd 0.007234f
C2506 vdd.t218 gnd 0.292327f
C2507 vdd.t217 gnd 0.299233f
C2508 vdd.t215 gnd 0.190842f
C2509 vdd.n804 gnd 0.10314f
C2510 vdd.n805 gnd 0.058504f
C2511 vdd.n806 gnd 0.010339f
C2512 vdd.n807 gnd 0.007234f
C2513 vdd.n808 gnd 0.007234f
C2514 vdd.t216 gnd 0.369642f
C2515 vdd.n809 gnd 0.007234f
C2516 vdd.n810 gnd 0.007234f
C2517 vdd.n811 gnd 0.007234f
C2518 vdd.n812 gnd 0.007234f
C2519 vdd.n813 gnd 0.007234f
C2520 vdd.n814 gnd 0.739285f
C2521 vdd.n815 gnd 0.007234f
C2522 vdd.n816 gnd 0.007234f
C2523 vdd.n817 gnd 0.646874f
C2524 vdd.n818 gnd 0.007234f
C2525 vdd.n819 gnd 0.007234f
C2526 vdd.n820 gnd 0.006383f
C2527 vdd.n821 gnd 0.007234f
C2528 vdd.n822 gnd 0.65231f
C2529 vdd.n823 gnd 0.007234f
C2530 vdd.n824 gnd 0.007234f
C2531 vdd.n825 gnd 0.007234f
C2532 vdd.n826 gnd 0.007234f
C2533 vdd.n827 gnd 0.007234f
C2534 vdd.n828 gnd 0.739285f
C2535 vdd.n829 gnd 0.007234f
C2536 vdd.n830 gnd 0.007234f
C2537 vdd.t199 gnd 0.331591f
C2538 vdd.t0 gnd 0.086975f
C2539 vdd.n831 gnd 0.007234f
C2540 vdd.n832 gnd 0.007234f
C2541 vdd.n833 gnd 0.007234f
C2542 vdd.t13 gnd 0.369642f
C2543 vdd.n834 gnd 0.007234f
C2544 vdd.n835 gnd 0.007234f
C2545 vdd.n836 gnd 0.007234f
C2546 vdd.n837 gnd 0.007234f
C2547 vdd.n838 gnd 0.007234f
C2548 vdd.t25 gnd 0.369642f
C2549 vdd.n839 gnd 0.007234f
C2550 vdd.n840 gnd 0.007234f
C2551 vdd.n841 gnd 0.614259f
C2552 vdd.n842 gnd 0.007234f
C2553 vdd.n843 gnd 0.007234f
C2554 vdd.n844 gnd 0.007234f
C2555 vdd.n845 gnd 0.451181f
C2556 vdd.n846 gnd 0.007234f
C2557 vdd.n847 gnd 0.007234f
C2558 vdd.t260 gnd 0.369642f
C2559 vdd.n848 gnd 0.007234f
C2560 vdd.n849 gnd 0.007234f
C2561 vdd.n850 gnd 0.007234f
C2562 vdd.n851 gnd 0.614259f
C2563 vdd.n852 gnd 0.007234f
C2564 vdd.n853 gnd 0.007234f
C2565 vdd.t38 gnd 0.315283f
C2566 vdd.t262 gnd 0.288104f
C2567 vdd.n854 gnd 0.007234f
C2568 vdd.n855 gnd 0.007234f
C2569 vdd.n856 gnd 0.007234f
C2570 vdd.t4 gnd 0.369642f
C2571 vdd.n857 gnd 0.007234f
C2572 vdd.n858 gnd 0.007234f
C2573 vdd.t22 gnd 0.369642f
C2574 vdd.n859 gnd 0.007234f
C2575 vdd.n860 gnd 0.007234f
C2576 vdd.n861 gnd 0.007234f
C2577 vdd.t23 gnd 0.271796f
C2578 vdd.n862 gnd 0.007234f
C2579 vdd.n863 gnd 0.007234f
C2580 vdd.n864 gnd 0.630567f
C2581 vdd.n865 gnd 0.007234f
C2582 vdd.n866 gnd 0.007234f
C2583 vdd.n867 gnd 0.007234f
C2584 vdd.n868 gnd 0.739285f
C2585 vdd.n869 gnd 0.007234f
C2586 vdd.n870 gnd 0.007234f
C2587 vdd.t250 gnd 0.331591f
C2588 vdd.n871 gnd 0.467489f
C2589 vdd.n872 gnd 0.007234f
C2590 vdd.n873 gnd 0.007234f
C2591 vdd.n874 gnd 0.007234f
C2592 vdd.t256 gnd 0.369642f
C2593 vdd.n875 gnd 0.007234f
C2594 vdd.n876 gnd 0.007234f
C2595 vdd.n877 gnd 0.007234f
C2596 vdd.n878 gnd 0.007234f
C2597 vdd.n879 gnd 0.007234f
C2598 vdd.t34 gnd 0.739285f
C2599 vdd.n880 gnd 0.007234f
C2600 vdd.n881 gnd 0.007234f
C2601 vdd.t220 gnd 0.369642f
C2602 vdd.n882 gnd 0.007234f
C2603 vdd.n883 gnd 0.017165f
C2604 vdd.n884 gnd 0.017165f
C2605 vdd.t36 gnd 0.695798f
C2606 vdd.n885 gnd 0.016026f
C2607 vdd.n886 gnd 0.016026f
C2608 vdd.n887 gnd 0.017165f
C2609 vdd.n888 gnd 0.007234f
C2610 vdd.n889 gnd 0.007234f
C2611 vdd.t10 gnd 0.695798f
C2612 vdd.n907 gnd 0.017165f
C2613 vdd.n925 gnd 0.016026f
C2614 vdd.n926 gnd 0.007234f
C2615 vdd.n927 gnd 0.016026f
C2616 vdd.t238 gnd 0.292327f
C2617 vdd.t237 gnd 0.299233f
C2618 vdd.t236 gnd 0.190842f
C2619 vdd.n928 gnd 0.10314f
C2620 vdd.n929 gnd 0.058504f
C2621 vdd.n930 gnd 0.016907f
C2622 vdd.n931 gnd 0.007234f
C2623 vdd.t8 gnd 0.739285f
C2624 vdd.n932 gnd 0.016026f
C2625 vdd.n933 gnd 0.007234f
C2626 vdd.n934 gnd 0.017165f
C2627 vdd.n935 gnd 0.007234f
C2628 vdd.t214 gnd 0.292327f
C2629 vdd.t213 gnd 0.299233f
C2630 vdd.t211 gnd 0.190842f
C2631 vdd.n936 gnd 0.10314f
C2632 vdd.n937 gnd 0.058504f
C2633 vdd.n938 gnd 0.010339f
C2634 vdd.n939 gnd 0.007234f
C2635 vdd.n940 gnd 0.007234f
C2636 vdd.t212 gnd 0.369642f
C2637 vdd.n941 gnd 0.007234f
C2638 vdd.n942 gnd 0.007234f
C2639 vdd.n943 gnd 0.007234f
C2640 vdd.n944 gnd 0.007234f
C2641 vdd.n945 gnd 0.007234f
C2642 vdd.n946 gnd 0.007234f
C2643 vdd.n947 gnd 0.739285f
C2644 vdd.n948 gnd 0.007234f
C2645 vdd.n949 gnd 0.007234f
C2646 vdd.t41 gnd 0.369642f
C2647 vdd.n950 gnd 0.007234f
C2648 vdd.n951 gnd 0.007234f
C2649 vdd.n952 gnd 0.007234f
C2650 vdd.n953 gnd 0.007234f
C2651 vdd.n954 gnd 0.467489f
C2652 vdd.n955 gnd 0.007234f
C2653 vdd.n956 gnd 0.007234f
C2654 vdd.n957 gnd 0.007234f
C2655 vdd.n958 gnd 0.007234f
C2656 vdd.n959 gnd 0.007234f
C2657 vdd.n960 gnd 0.630567f
C2658 vdd.n961 gnd 0.007234f
C2659 vdd.n962 gnd 0.007234f
C2660 vdd.t32 gnd 0.331591f
C2661 vdd.t12 gnd 0.271796f
C2662 vdd.n963 gnd 0.007234f
C2663 vdd.n964 gnd 0.007234f
C2664 vdd.n965 gnd 0.007234f
C2665 vdd.t1 gnd 0.369642f
C2666 vdd.n966 gnd 0.007234f
C2667 vdd.n967 gnd 0.007234f
C2668 vdd.t258 gnd 0.369642f
C2669 vdd.n968 gnd 0.007234f
C2670 vdd.n969 gnd 0.007234f
C2671 vdd.n970 gnd 0.007234f
C2672 vdd.t2 gnd 0.288104f
C2673 vdd.n971 gnd 0.007234f
C2674 vdd.n972 gnd 0.007234f
C2675 vdd.n973 gnd 0.614259f
C2676 vdd.n974 gnd 0.007234f
C2677 vdd.n975 gnd 0.007234f
C2678 vdd.n976 gnd 0.007234f
C2679 vdd.t6 gnd 0.369642f
C2680 vdd.n977 gnd 0.007234f
C2681 vdd.n978 gnd 0.007234f
C2682 vdd.t21 gnd 0.315283f
C2683 vdd.n979 gnd 0.451181f
C2684 vdd.n980 gnd 0.007234f
C2685 vdd.n981 gnd 0.007234f
C2686 vdd.n982 gnd 0.007234f
C2687 vdd.n983 gnd 0.614259f
C2688 vdd.n984 gnd 0.007234f
C2689 vdd.n985 gnd 0.007234f
C2690 vdd.t39 gnd 0.369642f
C2691 vdd.n986 gnd 0.007234f
C2692 vdd.n987 gnd 0.007234f
C2693 vdd.n988 gnd 0.007234f
C2694 vdd.n989 gnd 0.739285f
C2695 vdd.n990 gnd 0.007234f
C2696 vdd.n991 gnd 0.007234f
C2697 vdd.t18 gnd 0.369642f
C2698 vdd.n992 gnd 0.007234f
C2699 vdd.n993 gnd 0.007234f
C2700 vdd.n994 gnd 0.007234f
C2701 vdd.t31 gnd 0.086975f
C2702 vdd.n995 gnd 0.007234f
C2703 vdd.n996 gnd 0.007234f
C2704 vdd.n997 gnd 0.007234f
C2705 vdd.t231 gnd 0.299233f
C2706 vdd.t229 gnd 0.190842f
C2707 vdd.t232 gnd 0.299233f
C2708 vdd.n998 gnd 0.168181f
C2709 vdd.n999 gnd 0.007234f
C2710 vdd.n1000 gnd 0.007234f
C2711 vdd.n1001 gnd 0.739285f
C2712 vdd.n1002 gnd 0.007234f
C2713 vdd.n1003 gnd 0.007234f
C2714 vdd.t230 gnd 0.331591f
C2715 vdd.n1004 gnd 0.65231f
C2716 vdd.n1005 gnd 0.007234f
C2717 vdd.n1006 gnd 0.007234f
C2718 vdd.n1007 gnd 0.007234f
C2719 vdd.n1008 gnd 0.646874f
C2720 vdd.n1009 gnd 0.007234f
C2721 vdd.n1010 gnd 0.007234f
C2722 vdd.n1011 gnd 0.007234f
C2723 vdd.n1012 gnd 0.007234f
C2724 vdd.n1013 gnd 0.007234f
C2725 vdd.n1014 gnd 0.739285f
C2726 vdd.n1015 gnd 0.007234f
C2727 vdd.n1016 gnd 0.007234f
C2728 vdd.t173 gnd 0.369642f
C2729 vdd.n1017 gnd 0.007234f
C2730 vdd.n1018 gnd 0.017165f
C2731 vdd.n1019 gnd 0.017165f
C2732 vdd.n1020 gnd 7.4907f
C2733 vdd.n1021 gnd 0.016026f
C2734 vdd.n1022 gnd 0.016026f
C2735 vdd.n1023 gnd 0.017165f
C2736 vdd.n1024 gnd 0.007234f
C2737 vdd.n1025 gnd 0.007234f
C2738 vdd.n1026 gnd 0.007234f
C2739 vdd.n1027 gnd 0.007234f
C2740 vdd.n1028 gnd 0.007234f
C2741 vdd.n1029 gnd 0.007234f
C2742 vdd.n1030 gnd 0.007234f
C2743 vdd.n1031 gnd 0.007234f
C2744 vdd.n1033 gnd 0.007234f
C2745 vdd.n1034 gnd 0.007234f
C2746 vdd.n1035 gnd 0.006809f
C2747 vdd.n1038 gnd 0.024391f
C2748 vdd.n1039 gnd 0.008563f
C2749 vdd.n1040 gnd 0.010638f
C2750 vdd.n1042 gnd 0.010638f
C2751 vdd.n1043 gnd 0.007107f
C2752 vdd.n1044 gnd 0.603387f
C2753 vdd.n1045 gnd 7.68639f
C2754 vdd.n1046 gnd 0.010638f
C2755 vdd.n1047 gnd 0.024391f
C2756 vdd.n1048 gnd 0.008563f
C2757 vdd.n1049 gnd 0.010638f
C2758 vdd.n1050 gnd 0.008563f
C2759 vdd.n1051 gnd 0.010638f
C2760 vdd.n1052 gnd 1.08718f
C2761 vdd.n1053 gnd 0.010638f
C2762 vdd.n1054 gnd 0.008563f
C2763 vdd.n1055 gnd 0.008563f
C2764 vdd.n1056 gnd 0.010638f
C2765 vdd.n1057 gnd 0.008563f
C2766 vdd.n1058 gnd 0.010638f
C2767 vdd.t50 gnd 0.543592f
C2768 vdd.n1059 gnd 0.010638f
C2769 vdd.n1060 gnd 0.008563f
C2770 vdd.n1061 gnd 0.010638f
C2771 vdd.n1062 gnd 0.008563f
C2772 vdd.n1063 gnd 0.010638f
C2773 vdd.t151 gnd 0.543592f
C2774 vdd.n1064 gnd 0.010638f
C2775 vdd.n1065 gnd 0.008563f
C2776 vdd.n1066 gnd 0.010638f
C2777 vdd.n1067 gnd 0.008563f
C2778 vdd.n1068 gnd 0.010638f
C2779 vdd.t60 gnd 0.543592f
C2780 vdd.n1069 gnd 0.755593f
C2781 vdd.n1070 gnd 0.010638f
C2782 vdd.n1071 gnd 0.008563f
C2783 vdd.n1072 gnd 0.010638f
C2784 vdd.n1073 gnd 0.008563f
C2785 vdd.n1074 gnd 0.010638f
C2786 vdd.n1075 gnd 0.864311f
C2787 vdd.n1076 gnd 0.010638f
C2788 vdd.n1077 gnd 0.008563f
C2789 vdd.n1078 gnd 0.010638f
C2790 vdd.n1079 gnd 0.008563f
C2791 vdd.n1080 gnd 0.010638f
C2792 vdd.n1081 gnd 0.67949f
C2793 vdd.t81 gnd 0.543592f
C2794 vdd.n1082 gnd 0.010638f
C2795 vdd.n1083 gnd 0.008563f
C2796 vdd.n1084 gnd 0.010638f
C2797 vdd.n1085 gnd 0.008563f
C2798 vdd.n1086 gnd 0.010638f
C2799 vdd.t102 gnd 0.543592f
C2800 vdd.n1087 gnd 0.010638f
C2801 vdd.n1088 gnd 0.008563f
C2802 vdd.n1089 gnd 0.010638f
C2803 vdd.n1090 gnd 0.008563f
C2804 vdd.n1091 gnd 0.010638f
C2805 vdd.t132 gnd 0.543592f
C2806 vdd.n1092 gnd 0.592515f
C2807 vdd.n1093 gnd 0.010638f
C2808 vdd.n1094 gnd 0.008563f
C2809 vdd.n1095 gnd 0.010638f
C2810 vdd.n1096 gnd 0.008563f
C2811 vdd.n1097 gnd 0.010638f
C2812 vdd.t123 gnd 0.543592f
C2813 vdd.n1098 gnd 0.010638f
C2814 vdd.n1099 gnd 0.008563f
C2815 vdd.n1100 gnd 0.010638f
C2816 vdd.n1101 gnd 0.008563f
C2817 vdd.n1102 gnd 0.010638f
C2818 vdd.n1103 gnd 0.842567f
C2819 vdd.n1104 gnd 0.902362f
C2820 vdd.t58 gnd 0.543592f
C2821 vdd.n1105 gnd 0.010638f
C2822 vdd.n1106 gnd 0.008563f
C2823 vdd.n1107 gnd 0.010638f
C2824 vdd.n1108 gnd 0.008563f
C2825 vdd.n1109 gnd 0.010638f
C2826 vdd.n1110 gnd 0.657746f
C2827 vdd.n1111 gnd 0.010638f
C2828 vdd.n1112 gnd 0.008563f
C2829 vdd.n1113 gnd 0.010638f
C2830 vdd.n1114 gnd 0.008563f
C2831 vdd.n1115 gnd 0.010638f
C2832 vdd.t76 gnd 0.543592f
C2833 vdd.t66 gnd 0.543592f
C2834 vdd.n1116 gnd 0.010638f
C2835 vdd.n1117 gnd 0.008563f
C2836 vdd.n1118 gnd 0.010638f
C2837 vdd.n1119 gnd 0.008563f
C2838 vdd.n1120 gnd 0.010638f
C2839 vdd.t116 gnd 0.543592f
C2840 vdd.n1121 gnd 0.010638f
C2841 vdd.n1122 gnd 0.008563f
C2842 vdd.n1123 gnd 0.010638f
C2843 vdd.n1124 gnd 0.008563f
C2844 vdd.n1125 gnd 0.010638f
C2845 vdd.t118 gnd 0.543592f
C2846 vdd.n1126 gnd 0.79908f
C2847 vdd.n1127 gnd 0.010638f
C2848 vdd.n1128 gnd 0.008563f
C2849 vdd.n1129 gnd 0.010638f
C2850 vdd.n1130 gnd 0.008563f
C2851 vdd.n1131 gnd 0.010638f
C2852 vdd.n1132 gnd 1.08718f
C2853 vdd.n1133 gnd 0.010638f
C2854 vdd.n1134 gnd 0.008563f
C2855 vdd.n1135 gnd 0.010638f
C2856 vdd.n1136 gnd 0.008563f
C2857 vdd.n1137 gnd 0.010638f
C2858 vdd.n1138 gnd 0.91867f
C2859 vdd.n1139 gnd 0.010638f
C2860 vdd.n1140 gnd 0.008563f
C2861 vdd.n1141 gnd 0.024226f
C2862 vdd.n1142 gnd 0.007107f
C2863 vdd.n1143 gnd 0.024226f
C2864 vdd.n1144 gnd 1.43508f
C2865 vdd.n1145 gnd 0.024226f
C2866 vdd.n1146 gnd 0.007107f
C2867 vdd.n1147 gnd 0.010638f
C2868 vdd.t186 gnd 0.130879f
C2869 vdd.t187 gnd 0.139874f
C2870 vdd.t184 gnd 0.170926f
C2871 vdd.n1148 gnd 0.219103f
C2872 vdd.n1149 gnd 0.184943f
C2873 vdd.n1150 gnd 0.014043f
C2874 vdd.n1151 gnd 0.010638f
C2875 vdd.n1182 gnd 0.010638f
C2876 vdd.n1183 gnd 0.010638f
C2877 vdd.n1184 gnd 0.024391f
C2878 vdd.n1185 gnd 0.008563f
C2879 vdd.n1186 gnd 0.010638f
C2880 vdd.n1187 gnd 0.010638f
C2881 vdd.n1188 gnd 0.010638f
C2882 vdd.n1189 gnd 0.010638f
C2883 vdd.n1190 gnd 0.008563f
C2884 vdd.n1191 gnd 0.010638f
C2885 vdd.n1192 gnd 0.010638f
C2886 vdd.n1193 gnd 0.010638f
C2887 vdd.n1194 gnd 0.010638f
C2888 vdd.n1195 gnd 0.010638f
C2889 vdd.n1196 gnd 0.008563f
C2890 vdd.n1197 gnd 0.010638f
C2891 vdd.n1198 gnd 0.010638f
C2892 vdd.n1199 gnd 0.010638f
C2893 vdd.n1200 gnd 0.010638f
C2894 vdd.n1201 gnd 0.010638f
C2895 vdd.n1202 gnd 0.008563f
C2896 vdd.n1203 gnd 0.010638f
C2897 vdd.n1204 gnd 0.010638f
C2898 vdd.n1205 gnd 0.010638f
C2899 vdd.n1206 gnd 0.010638f
C2900 vdd.n1207 gnd 0.010638f
C2901 vdd.n1208 gnd 0.00715f
C2902 vdd.n1209 gnd 0.010638f
C2903 vdd.n1210 gnd 0.010638f
C2904 vdd.n1211 gnd 0.010638f
C2905 vdd.n1212 gnd 0.008563f
C2906 vdd.n1213 gnd 0.010638f
C2907 vdd.n1214 gnd 0.010638f
C2908 vdd.n1215 gnd 0.010638f
C2909 vdd.n1216 gnd 0.010638f
C2910 vdd.n1217 gnd 0.010638f
C2911 vdd.n1218 gnd 0.008563f
C2912 vdd.n1219 gnd 0.010638f
C2913 vdd.n1220 gnd 0.010638f
C2914 vdd.n1221 gnd 0.010638f
C2915 vdd.n1222 gnd 0.010638f
C2916 vdd.n1223 gnd 0.010638f
C2917 vdd.n1224 gnd 0.008563f
C2918 vdd.n1225 gnd 0.010638f
C2919 vdd.n1226 gnd 0.010638f
C2920 vdd.n1227 gnd 0.010638f
C2921 vdd.n1228 gnd 0.010638f
C2922 vdd.n1229 gnd 0.010638f
C2923 vdd.n1230 gnd 0.008563f
C2924 vdd.n1231 gnd 0.010638f
C2925 vdd.n1232 gnd 0.010638f
C2926 vdd.n1233 gnd 0.010638f
C2927 vdd.n1234 gnd 0.010638f
C2928 vdd.n1235 gnd 0.010638f
C2929 vdd.n1236 gnd 0.008563f
C2930 vdd.n1237 gnd 0.010638f
C2931 vdd.n1238 gnd 0.010638f
C2932 vdd.n1239 gnd 0.010638f
C2933 vdd.n1240 gnd 0.010638f
C2934 vdd.n1241 gnd 0.008477f
C2935 vdd.n1242 gnd 0.010638f
C2936 vdd.n1243 gnd 0.010638f
C2937 vdd.n1244 gnd 0.010638f
C2938 vdd.n1245 gnd 0.010638f
C2939 vdd.n1246 gnd 0.010638f
C2940 vdd.n1247 gnd 0.008563f
C2941 vdd.n1248 gnd 0.010638f
C2942 vdd.n1249 gnd 0.010638f
C2943 vdd.n1250 gnd 0.010638f
C2944 vdd.n1251 gnd 0.010638f
C2945 vdd.n1252 gnd 0.010638f
C2946 vdd.n1253 gnd 0.008563f
C2947 vdd.n1254 gnd 0.010638f
C2948 vdd.n1255 gnd 0.010638f
C2949 vdd.n1256 gnd 0.010638f
C2950 vdd.n1257 gnd 0.010638f
C2951 vdd.n1258 gnd 0.010638f
C2952 vdd.n1259 gnd 0.008563f
C2953 vdd.n1260 gnd 0.010638f
C2954 vdd.n1261 gnd 0.010638f
C2955 vdd.n1262 gnd 0.010638f
C2956 vdd.n1263 gnd 0.010638f
C2957 vdd.n1264 gnd 0.010638f
C2958 vdd.n1265 gnd 0.008563f
C2959 vdd.n1266 gnd 0.010638f
C2960 vdd.n1267 gnd 0.010638f
C2961 vdd.n1268 gnd 0.010638f
C2962 vdd.n1269 gnd 0.010638f
C2963 vdd.n1270 gnd 0.010638f
C2964 vdd.n1271 gnd 0.004495f
C2965 vdd.n1272 gnd 0.010638f
C2966 vdd.n1273 gnd 0.008563f
C2967 vdd.n1274 gnd 0.008563f
C2968 vdd.n1275 gnd 0.008563f
C2969 vdd.n1276 gnd 0.010638f
C2970 vdd.n1277 gnd 0.010638f
C2971 vdd.n1278 gnd 0.010638f
C2972 vdd.n1279 gnd 0.008563f
C2973 vdd.n1280 gnd 0.008563f
C2974 vdd.n1281 gnd 0.008563f
C2975 vdd.n1282 gnd 0.010638f
C2976 vdd.n1283 gnd 0.010638f
C2977 vdd.n1284 gnd 0.010638f
C2978 vdd.n1285 gnd 0.008563f
C2979 vdd.n1286 gnd 0.008563f
C2980 vdd.n1287 gnd 0.008563f
C2981 vdd.n1288 gnd 0.010638f
C2982 vdd.n1289 gnd 0.010638f
C2983 vdd.n1290 gnd 0.010638f
C2984 vdd.n1291 gnd 0.008563f
C2985 vdd.n1292 gnd 0.008563f
C2986 vdd.n1293 gnd 0.008563f
C2987 vdd.n1294 gnd 0.010638f
C2988 vdd.n1295 gnd 0.010638f
C2989 vdd.n1296 gnd 0.010638f
C2990 vdd.n1297 gnd 0.008563f
C2991 vdd.n1298 gnd 0.008563f
C2992 vdd.n1299 gnd 0.008563f
C2993 vdd.n1300 gnd 0.010638f
C2994 vdd.n1301 gnd 0.010638f
C2995 vdd.n1302 gnd 0.010638f
C2996 vdd.n1303 gnd 0.010638f
C2997 vdd.t196 gnd 0.130879f
C2998 vdd.t197 gnd 0.139874f
C2999 vdd.t195 gnd 0.170926f
C3000 vdd.n1304 gnd 0.219103f
C3001 vdd.n1305 gnd 0.184943f
C3002 vdd.n1306 gnd 0.018324f
C3003 vdd.n1307 gnd 0.005823f
C3004 vdd.n1308 gnd 0.008563f
C3005 vdd.n1309 gnd 0.010638f
C3006 vdd.n1310 gnd 0.010638f
C3007 vdd.n1311 gnd 0.010638f
C3008 vdd.n1312 gnd 0.008563f
C3009 vdd.n1313 gnd 0.008563f
C3010 vdd.n1314 gnd 0.008563f
C3011 vdd.n1315 gnd 0.010638f
C3012 vdd.n1316 gnd 0.010638f
C3013 vdd.n1317 gnd 0.010638f
C3014 vdd.n1318 gnd 0.008563f
C3015 vdd.n1319 gnd 0.008563f
C3016 vdd.n1320 gnd 0.008563f
C3017 vdd.n1321 gnd 0.010638f
C3018 vdd.n1322 gnd 0.010638f
C3019 vdd.n1323 gnd 0.010638f
C3020 vdd.n1324 gnd 0.008563f
C3021 vdd.n1325 gnd 0.008563f
C3022 vdd.n1326 gnd 0.008563f
C3023 vdd.n1327 gnd 0.010638f
C3024 vdd.n1328 gnd 0.010638f
C3025 vdd.n1329 gnd 0.010638f
C3026 vdd.n1330 gnd 0.008563f
C3027 vdd.n1331 gnd 0.008563f
C3028 vdd.n1332 gnd 0.008563f
C3029 vdd.n1333 gnd 0.010638f
C3030 vdd.n1334 gnd 0.010638f
C3031 vdd.n1335 gnd 0.010638f
C3032 vdd.n1336 gnd 0.008563f
C3033 vdd.n1337 gnd 0.00715f
C3034 vdd.n1338 gnd 0.010638f
C3035 vdd.n1339 gnd 0.010638f
C3036 vdd.t203 gnd 0.130879f
C3037 vdd.t204 gnd 0.139874f
C3038 vdd.t202 gnd 0.170926f
C3039 vdd.n1340 gnd 0.219103f
C3040 vdd.n1341 gnd 0.184943f
C3041 vdd.n1342 gnd 0.018324f
C3042 vdd.n1343 gnd 0.010638f
C3043 vdd.n1344 gnd 0.010638f
C3044 vdd.n1345 gnd 0.010638f
C3045 vdd.n1346 gnd 0.008563f
C3046 vdd.n1347 gnd 0.008563f
C3047 vdd.n1348 gnd 0.008563f
C3048 vdd.n1349 gnd 0.010638f
C3049 vdd.n1350 gnd 0.010638f
C3050 vdd.n1351 gnd 0.010638f
C3051 vdd.n1352 gnd 0.008563f
C3052 vdd.n1353 gnd 0.008563f
C3053 vdd.n1354 gnd 0.008563f
C3054 vdd.n1355 gnd 0.010638f
C3055 vdd.n1356 gnd 0.010638f
C3056 vdd.n1357 gnd 0.010638f
C3057 vdd.n1358 gnd 0.008563f
C3058 vdd.n1359 gnd 0.008563f
C3059 vdd.n1360 gnd 0.008563f
C3060 vdd.n1361 gnd 0.010638f
C3061 vdd.n1362 gnd 0.010638f
C3062 vdd.n1363 gnd 0.010638f
C3063 vdd.n1364 gnd 0.008563f
C3064 vdd.n1365 gnd 0.008563f
C3065 vdd.n1366 gnd 0.008563f
C3066 vdd.n1367 gnd 0.010638f
C3067 vdd.n1368 gnd 0.010638f
C3068 vdd.n1369 gnd 0.010638f
C3069 vdd.n1370 gnd 0.008563f
C3070 vdd.n1371 gnd 0.007107f
C3071 vdd.n1372 gnd 0.024391f
C3072 vdd.n1374 gnd 2.40268f
C3073 vdd.n1375 gnd 0.024391f
C3074 vdd.n1376 gnd 0.004067f
C3075 vdd.n1377 gnd 0.024391f
C3076 vdd.n1378 gnd 0.024226f
C3077 vdd.n1379 gnd 0.010638f
C3078 vdd.n1380 gnd 0.008563f
C3079 vdd.n1381 gnd 0.010638f
C3080 vdd.t185 gnd 0.543592f
C3081 vdd.n1382 gnd 0.712105f
C3082 vdd.n1383 gnd 0.010638f
C3083 vdd.n1384 gnd 0.008563f
C3084 vdd.n1385 gnd 0.010638f
C3085 vdd.n1386 gnd 0.010638f
C3086 vdd.n1387 gnd 0.010638f
C3087 vdd.n1388 gnd 0.008563f
C3088 vdd.n1389 gnd 0.010638f
C3089 vdd.n1390 gnd 1.08718f
C3090 vdd.n1391 gnd 0.010638f
C3091 vdd.n1392 gnd 0.008563f
C3092 vdd.n1393 gnd 0.010638f
C3093 vdd.n1394 gnd 0.010638f
C3094 vdd.n1395 gnd 0.010638f
C3095 vdd.n1396 gnd 0.008563f
C3096 vdd.n1397 gnd 0.010638f
C3097 vdd.n1398 gnd 0.902362f
C3098 vdd.t56 gnd 0.543592f
C3099 vdd.n1399 gnd 0.625131f
C3100 vdd.n1400 gnd 0.010638f
C3101 vdd.n1401 gnd 0.008563f
C3102 vdd.n1402 gnd 0.010638f
C3103 vdd.n1403 gnd 0.010638f
C3104 vdd.n1404 gnd 0.010638f
C3105 vdd.n1405 gnd 0.008563f
C3106 vdd.n1406 gnd 0.010638f
C3107 vdd.n1407 gnd 0.646874f
C3108 vdd.n1408 gnd 0.010638f
C3109 vdd.n1409 gnd 0.008563f
C3110 vdd.n1410 gnd 0.010638f
C3111 vdd.n1411 gnd 0.010638f
C3112 vdd.n1412 gnd 0.010638f
C3113 vdd.n1413 gnd 0.008563f
C3114 vdd.n1414 gnd 0.010638f
C3115 vdd.n1415 gnd 0.614259f
C3116 vdd.n1416 gnd 0.831696f
C3117 vdd.n1417 gnd 0.010638f
C3118 vdd.n1418 gnd 0.008563f
C3119 vdd.n1419 gnd 0.010638f
C3120 vdd.n1420 gnd 0.010638f
C3121 vdd.n1421 gnd 0.010638f
C3122 vdd.n1422 gnd 0.008563f
C3123 vdd.n1423 gnd 0.010638f
C3124 vdd.n1424 gnd 0.902362f
C3125 vdd.n1425 gnd 0.010638f
C3126 vdd.n1426 gnd 0.008563f
C3127 vdd.n1427 gnd 0.010638f
C3128 vdd.n1428 gnd 0.010638f
C3129 vdd.n1429 gnd 0.010638f
C3130 vdd.n1430 gnd 0.008563f
C3131 vdd.n1431 gnd 0.010638f
C3132 vdd.t94 gnd 0.543592f
C3133 vdd.n1432 gnd 0.788208f
C3134 vdd.n1433 gnd 0.010638f
C3135 vdd.n1434 gnd 0.008563f
C3136 vdd.n1435 gnd 0.010638f
C3137 vdd.n1436 gnd 0.010638f
C3138 vdd.n1437 gnd 0.010638f
C3139 vdd.n1438 gnd 0.008563f
C3140 vdd.n1439 gnd 0.010638f
C3141 vdd.n1440 gnd 0.603387f
C3142 vdd.n1441 gnd 0.010638f
C3143 vdd.n1442 gnd 0.008563f
C3144 vdd.n1443 gnd 0.010638f
C3145 vdd.n1444 gnd 0.010638f
C3146 vdd.n1445 gnd 0.010638f
C3147 vdd.n1446 gnd 0.008563f
C3148 vdd.n1447 gnd 0.010638f
C3149 vdd.n1448 gnd 0.777336f
C3150 vdd.n1449 gnd 0.668618f
C3151 vdd.n1450 gnd 0.010638f
C3152 vdd.n1451 gnd 0.008563f
C3153 vdd.n1452 gnd 0.008176f
C3154 vdd.n1453 gnd 0.005838f
C3155 vdd.n1454 gnd 0.005418f
C3156 vdd.n1455 gnd 0.002997f
C3157 vdd.n1456 gnd 0.006881f
C3158 vdd.n1457 gnd 0.002911f
C3159 vdd.n1458 gnd 0.003083f
C3160 vdd.n1459 gnd 0.005418f
C3161 vdd.n1460 gnd 0.002911f
C3162 vdd.n1461 gnd 0.006881f
C3163 vdd.n1462 gnd 0.003083f
C3164 vdd.n1463 gnd 0.005418f
C3165 vdd.n1464 gnd 0.002911f
C3166 vdd.n1465 gnd 0.005161f
C3167 vdd.n1466 gnd 0.005176f
C3168 vdd.t51 gnd 0.014784f
C3169 vdd.n1467 gnd 0.032893f
C3170 vdd.n1468 gnd 0.171185f
C3171 vdd.n1469 gnd 0.002911f
C3172 vdd.n1470 gnd 0.003083f
C3173 vdd.n1471 gnd 0.006881f
C3174 vdd.n1472 gnd 0.006881f
C3175 vdd.n1473 gnd 0.003083f
C3176 vdd.n1474 gnd 0.002911f
C3177 vdd.n1475 gnd 0.005418f
C3178 vdd.n1476 gnd 0.005418f
C3179 vdd.n1477 gnd 0.002911f
C3180 vdd.n1478 gnd 0.003083f
C3181 vdd.n1479 gnd 0.006881f
C3182 vdd.n1480 gnd 0.006881f
C3183 vdd.n1481 gnd 0.003083f
C3184 vdd.n1482 gnd 0.002911f
C3185 vdd.n1483 gnd 0.005418f
C3186 vdd.n1484 gnd 0.005418f
C3187 vdd.n1485 gnd 0.002911f
C3188 vdd.n1486 gnd 0.003083f
C3189 vdd.n1487 gnd 0.006881f
C3190 vdd.n1488 gnd 0.006881f
C3191 vdd.n1489 gnd 0.016268f
C3192 vdd.n1490 gnd 0.002997f
C3193 vdd.n1491 gnd 0.002911f
C3194 vdd.n1492 gnd 0.014003f
C3195 vdd.n1493 gnd 0.009776f
C3196 vdd.t109 gnd 0.03425f
C3197 vdd.t158 gnd 0.03425f
C3198 vdd.n1494 gnd 0.235391f
C3199 vdd.n1495 gnd 0.185099f
C3200 vdd.t82 gnd 0.03425f
C3201 vdd.t138 gnd 0.03425f
C3202 vdd.n1496 gnd 0.235391f
C3203 vdd.n1497 gnd 0.149374f
C3204 vdd.t103 gnd 0.03425f
C3205 vdd.t147 gnd 0.03425f
C3206 vdd.n1498 gnd 0.235391f
C3207 vdd.n1499 gnd 0.149374f
C3208 vdd.t124 gnd 0.03425f
C3209 vdd.t165 gnd 0.03425f
C3210 vdd.n1500 gnd 0.235391f
C3211 vdd.n1501 gnd 0.149374f
C3212 vdd.t95 gnd 0.03425f
C3213 vdd.t59 gnd 0.03425f
C3214 vdd.n1502 gnd 0.235391f
C3215 vdd.n1503 gnd 0.149374f
C3216 vdd.t112 gnd 0.03425f
C3217 vdd.t67 gnd 0.03425f
C3218 vdd.n1504 gnd 0.235391f
C3219 vdd.n1505 gnd 0.149374f
C3220 vdd.t154 gnd 0.03425f
C3221 vdd.t170 gnd 0.03425f
C3222 vdd.n1506 gnd 0.235391f
C3223 vdd.n1507 gnd 0.149374f
C3224 vdd.n1508 gnd 0.005838f
C3225 vdd.n1509 gnd 0.005418f
C3226 vdd.n1510 gnd 0.002997f
C3227 vdd.n1511 gnd 0.006881f
C3228 vdd.n1512 gnd 0.002911f
C3229 vdd.n1513 gnd 0.003083f
C3230 vdd.n1514 gnd 0.005418f
C3231 vdd.n1515 gnd 0.002911f
C3232 vdd.n1516 gnd 0.006881f
C3233 vdd.n1517 gnd 0.003083f
C3234 vdd.n1518 gnd 0.005418f
C3235 vdd.n1519 gnd 0.002911f
C3236 vdd.n1520 gnd 0.005161f
C3237 vdd.n1521 gnd 0.005176f
C3238 vdd.t72 gnd 0.014784f
C3239 vdd.n1522 gnd 0.032893f
C3240 vdd.n1523 gnd 0.171185f
C3241 vdd.n1524 gnd 0.002911f
C3242 vdd.n1525 gnd 0.003083f
C3243 vdd.n1526 gnd 0.006881f
C3244 vdd.n1527 gnd 0.006881f
C3245 vdd.n1528 gnd 0.003083f
C3246 vdd.n1529 gnd 0.002911f
C3247 vdd.n1530 gnd 0.005418f
C3248 vdd.n1531 gnd 0.005418f
C3249 vdd.n1532 gnd 0.002911f
C3250 vdd.n1533 gnd 0.003083f
C3251 vdd.n1534 gnd 0.006881f
C3252 vdd.n1535 gnd 0.006881f
C3253 vdd.n1536 gnd 0.003083f
C3254 vdd.n1537 gnd 0.002911f
C3255 vdd.n1538 gnd 0.005418f
C3256 vdd.n1539 gnd 0.005418f
C3257 vdd.n1540 gnd 0.002911f
C3258 vdd.n1541 gnd 0.003083f
C3259 vdd.n1542 gnd 0.006881f
C3260 vdd.n1543 gnd 0.006881f
C3261 vdd.n1544 gnd 0.016268f
C3262 vdd.n1545 gnd 0.002997f
C3263 vdd.n1546 gnd 0.002911f
C3264 vdd.n1547 gnd 0.014003f
C3265 vdd.n1548 gnd 0.00947f
C3266 vdd.n1549 gnd 0.111135f
C3267 vdd.n1550 gnd 0.005838f
C3268 vdd.n1551 gnd 0.005418f
C3269 vdd.n1552 gnd 0.002997f
C3270 vdd.n1553 gnd 0.006881f
C3271 vdd.n1554 gnd 0.002911f
C3272 vdd.n1555 gnd 0.003083f
C3273 vdd.n1556 gnd 0.005418f
C3274 vdd.n1557 gnd 0.002911f
C3275 vdd.n1558 gnd 0.006881f
C3276 vdd.n1559 gnd 0.003083f
C3277 vdd.n1560 gnd 0.005418f
C3278 vdd.n1561 gnd 0.002911f
C3279 vdd.n1562 gnd 0.005161f
C3280 vdd.n1563 gnd 0.005176f
C3281 vdd.t149 gnd 0.014784f
C3282 vdd.n1564 gnd 0.032893f
C3283 vdd.n1565 gnd 0.171185f
C3284 vdd.n1566 gnd 0.002911f
C3285 vdd.n1567 gnd 0.003083f
C3286 vdd.n1568 gnd 0.006881f
C3287 vdd.n1569 gnd 0.006881f
C3288 vdd.n1570 gnd 0.003083f
C3289 vdd.n1571 gnd 0.002911f
C3290 vdd.n1572 gnd 0.005418f
C3291 vdd.n1573 gnd 0.005418f
C3292 vdd.n1574 gnd 0.002911f
C3293 vdd.n1575 gnd 0.003083f
C3294 vdd.n1576 gnd 0.006881f
C3295 vdd.n1577 gnd 0.006881f
C3296 vdd.n1578 gnd 0.003083f
C3297 vdd.n1579 gnd 0.002911f
C3298 vdd.n1580 gnd 0.005418f
C3299 vdd.n1581 gnd 0.005418f
C3300 vdd.n1582 gnd 0.002911f
C3301 vdd.n1583 gnd 0.003083f
C3302 vdd.n1584 gnd 0.006881f
C3303 vdd.n1585 gnd 0.006881f
C3304 vdd.n1586 gnd 0.016268f
C3305 vdd.n1587 gnd 0.002997f
C3306 vdd.n1588 gnd 0.002911f
C3307 vdd.n1589 gnd 0.014003f
C3308 vdd.n1590 gnd 0.009776f
C3309 vdd.t61 gnd 0.03425f
C3310 vdd.t152 gnd 0.03425f
C3311 vdd.n1591 gnd 0.235391f
C3312 vdd.n1592 gnd 0.185099f
C3313 vdd.t145 gnd 0.03425f
C3314 vdd.t135 gnd 0.03425f
C3315 vdd.n1593 gnd 0.235391f
C3316 vdd.n1594 gnd 0.149374f
C3317 vdd.t105 gnd 0.03425f
C3318 vdd.t49 gnd 0.03425f
C3319 vdd.n1595 gnd 0.235391f
C3320 vdd.n1596 gnd 0.149374f
C3321 vdd.t161 gnd 0.03425f
C3322 vdd.t133 gnd 0.03425f
C3323 vdd.n1597 gnd 0.235391f
C3324 vdd.n1598 gnd 0.149374f
C3325 vdd.t130 gnd 0.03425f
C3326 vdd.t83 gnd 0.03425f
C3327 vdd.n1599 gnd 0.235391f
C3328 vdd.n1600 gnd 0.149374f
C3329 vdd.t77 gnd 0.03425f
C3330 vdd.t131 gnd 0.03425f
C3331 vdd.n1601 gnd 0.235391f
C3332 vdd.n1602 gnd 0.149374f
C3333 vdd.t119 gnd 0.03425f
C3334 vdd.t117 gnd 0.03425f
C3335 vdd.n1603 gnd 0.235391f
C3336 vdd.n1604 gnd 0.149374f
C3337 vdd.n1605 gnd 0.005838f
C3338 vdd.n1606 gnd 0.005418f
C3339 vdd.n1607 gnd 0.002997f
C3340 vdd.n1608 gnd 0.006881f
C3341 vdd.n1609 gnd 0.002911f
C3342 vdd.n1610 gnd 0.003083f
C3343 vdd.n1611 gnd 0.005418f
C3344 vdd.n1612 gnd 0.002911f
C3345 vdd.n1613 gnd 0.006881f
C3346 vdd.n1614 gnd 0.003083f
C3347 vdd.n1615 gnd 0.005418f
C3348 vdd.n1616 gnd 0.002911f
C3349 vdd.n1617 gnd 0.005161f
C3350 vdd.n1618 gnd 0.005176f
C3351 vdd.t57 gnd 0.014784f
C3352 vdd.n1619 gnd 0.032893f
C3353 vdd.n1620 gnd 0.171185f
C3354 vdd.n1621 gnd 0.002911f
C3355 vdd.n1622 gnd 0.003083f
C3356 vdd.n1623 gnd 0.006881f
C3357 vdd.n1624 gnd 0.006881f
C3358 vdd.n1625 gnd 0.003083f
C3359 vdd.n1626 gnd 0.002911f
C3360 vdd.n1627 gnd 0.005418f
C3361 vdd.n1628 gnd 0.005418f
C3362 vdd.n1629 gnd 0.002911f
C3363 vdd.n1630 gnd 0.003083f
C3364 vdd.n1631 gnd 0.006881f
C3365 vdd.n1632 gnd 0.006881f
C3366 vdd.n1633 gnd 0.003083f
C3367 vdd.n1634 gnd 0.002911f
C3368 vdd.n1635 gnd 0.005418f
C3369 vdd.n1636 gnd 0.005418f
C3370 vdd.n1637 gnd 0.002911f
C3371 vdd.n1638 gnd 0.003083f
C3372 vdd.n1639 gnd 0.006881f
C3373 vdd.n1640 gnd 0.006881f
C3374 vdd.n1641 gnd 0.016268f
C3375 vdd.n1642 gnd 0.002997f
C3376 vdd.n1643 gnd 0.002911f
C3377 vdd.n1644 gnd 0.014003f
C3378 vdd.n1645 gnd 0.00947f
C3379 vdd.n1646 gnd 0.066114f
C3380 vdd.n1647 gnd 0.238226f
C3381 vdd.n1648 gnd 0.005838f
C3382 vdd.n1649 gnd 0.005418f
C3383 vdd.n1650 gnd 0.002997f
C3384 vdd.n1651 gnd 0.006881f
C3385 vdd.n1652 gnd 0.002911f
C3386 vdd.n1653 gnd 0.003083f
C3387 vdd.n1654 gnd 0.005418f
C3388 vdd.n1655 gnd 0.002911f
C3389 vdd.n1656 gnd 0.006881f
C3390 vdd.n1657 gnd 0.003083f
C3391 vdd.n1658 gnd 0.005418f
C3392 vdd.n1659 gnd 0.002911f
C3393 vdd.n1660 gnd 0.005161f
C3394 vdd.n1661 gnd 0.005176f
C3395 vdd.t163 gnd 0.014784f
C3396 vdd.n1662 gnd 0.032893f
C3397 vdd.n1663 gnd 0.171185f
C3398 vdd.n1664 gnd 0.002911f
C3399 vdd.n1665 gnd 0.003083f
C3400 vdd.n1666 gnd 0.006881f
C3401 vdd.n1667 gnd 0.006881f
C3402 vdd.n1668 gnd 0.003083f
C3403 vdd.n1669 gnd 0.002911f
C3404 vdd.n1670 gnd 0.005418f
C3405 vdd.n1671 gnd 0.005418f
C3406 vdd.n1672 gnd 0.002911f
C3407 vdd.n1673 gnd 0.003083f
C3408 vdd.n1674 gnd 0.006881f
C3409 vdd.n1675 gnd 0.006881f
C3410 vdd.n1676 gnd 0.003083f
C3411 vdd.n1677 gnd 0.002911f
C3412 vdd.n1678 gnd 0.005418f
C3413 vdd.n1679 gnd 0.005418f
C3414 vdd.n1680 gnd 0.002911f
C3415 vdd.n1681 gnd 0.003083f
C3416 vdd.n1682 gnd 0.006881f
C3417 vdd.n1683 gnd 0.006881f
C3418 vdd.n1684 gnd 0.016268f
C3419 vdd.n1685 gnd 0.002997f
C3420 vdd.n1686 gnd 0.002911f
C3421 vdd.n1687 gnd 0.014003f
C3422 vdd.n1688 gnd 0.009776f
C3423 vdd.t71 gnd 0.03425f
C3424 vdd.t162 gnd 0.03425f
C3425 vdd.n1689 gnd 0.235391f
C3426 vdd.n1690 gnd 0.185099f
C3427 vdd.t160 gnd 0.03425f
C3428 vdd.t144 gnd 0.03425f
C3429 vdd.n1691 gnd 0.235391f
C3430 vdd.n1692 gnd 0.149374f
C3431 vdd.t120 gnd 0.03425f
C3432 vdd.t74 gnd 0.03425f
C3433 vdd.n1693 gnd 0.235391f
C3434 vdd.n1694 gnd 0.149374f
C3435 vdd.t171 gnd 0.03425f
C3436 vdd.t142 gnd 0.03425f
C3437 vdd.n1695 gnd 0.235391f
C3438 vdd.n1696 gnd 0.149374f
C3439 vdd.t140 gnd 0.03425f
C3440 vdd.t97 gnd 0.03425f
C3441 vdd.n1697 gnd 0.235391f
C3442 vdd.n1698 gnd 0.149374f
C3443 vdd.t96 gnd 0.03425f
C3444 vdd.t141 gnd 0.03425f
C3445 vdd.n1699 gnd 0.235391f
C3446 vdd.n1700 gnd 0.149374f
C3447 vdd.t129 gnd 0.03425f
C3448 vdd.t128 gnd 0.03425f
C3449 vdd.n1701 gnd 0.235391f
C3450 vdd.n1702 gnd 0.149374f
C3451 vdd.n1703 gnd 0.005838f
C3452 vdd.n1704 gnd 0.005418f
C3453 vdd.n1705 gnd 0.002997f
C3454 vdd.n1706 gnd 0.006881f
C3455 vdd.n1707 gnd 0.002911f
C3456 vdd.n1708 gnd 0.003083f
C3457 vdd.n1709 gnd 0.005418f
C3458 vdd.n1710 gnd 0.002911f
C3459 vdd.n1711 gnd 0.006881f
C3460 vdd.n1712 gnd 0.003083f
C3461 vdd.n1713 gnd 0.005418f
C3462 vdd.n1714 gnd 0.002911f
C3463 vdd.n1715 gnd 0.005161f
C3464 vdd.n1716 gnd 0.005176f
C3465 vdd.t73 gnd 0.014784f
C3466 vdd.n1717 gnd 0.032893f
C3467 vdd.n1718 gnd 0.171185f
C3468 vdd.n1719 gnd 0.002911f
C3469 vdd.n1720 gnd 0.003083f
C3470 vdd.n1721 gnd 0.006881f
C3471 vdd.n1722 gnd 0.006881f
C3472 vdd.n1723 gnd 0.003083f
C3473 vdd.n1724 gnd 0.002911f
C3474 vdd.n1725 gnd 0.005418f
C3475 vdd.n1726 gnd 0.005418f
C3476 vdd.n1727 gnd 0.002911f
C3477 vdd.n1728 gnd 0.003083f
C3478 vdd.n1729 gnd 0.006881f
C3479 vdd.n1730 gnd 0.006881f
C3480 vdd.n1731 gnd 0.003083f
C3481 vdd.n1732 gnd 0.002911f
C3482 vdd.n1733 gnd 0.005418f
C3483 vdd.n1734 gnd 0.005418f
C3484 vdd.n1735 gnd 0.002911f
C3485 vdd.n1736 gnd 0.003083f
C3486 vdd.n1737 gnd 0.006881f
C3487 vdd.n1738 gnd 0.006881f
C3488 vdd.n1739 gnd 0.016268f
C3489 vdd.n1740 gnd 0.002997f
C3490 vdd.n1741 gnd 0.002911f
C3491 vdd.n1742 gnd 0.014003f
C3492 vdd.n1743 gnd 0.00947f
C3493 vdd.n1744 gnd 0.066114f
C3494 vdd.n1745 gnd 0.266781f
C3495 vdd.n1746 gnd 2.54484f
C3496 vdd.n1747 gnd 0.627487f
C3497 vdd.n1748 gnd 0.008176f
C3498 vdd.n1749 gnd 0.010638f
C3499 vdd.n1750 gnd 0.008563f
C3500 vdd.n1751 gnd 0.010638f
C3501 vdd.n1752 gnd 0.853439f
C3502 vdd.n1753 gnd 0.010638f
C3503 vdd.n1754 gnd 0.008563f
C3504 vdd.n1755 gnd 0.010638f
C3505 vdd.n1756 gnd 0.010638f
C3506 vdd.n1757 gnd 0.010638f
C3507 vdd.n1758 gnd 0.008563f
C3508 vdd.n1759 gnd 0.010638f
C3509 vdd.t48 gnd 0.543592f
C3510 vdd.n1760 gnd 0.902362f
C3511 vdd.n1761 gnd 0.010638f
C3512 vdd.n1762 gnd 0.008563f
C3513 vdd.n1763 gnd 0.010638f
C3514 vdd.n1764 gnd 0.010638f
C3515 vdd.n1765 gnd 0.010638f
C3516 vdd.n1766 gnd 0.008563f
C3517 vdd.n1767 gnd 0.010638f
C3518 vdd.n1768 gnd 0.766465f
C3519 vdd.n1769 gnd 0.010638f
C3520 vdd.n1770 gnd 0.008563f
C3521 vdd.n1771 gnd 0.010638f
C3522 vdd.n1772 gnd 0.010638f
C3523 vdd.n1773 gnd 0.010638f
C3524 vdd.n1774 gnd 0.008563f
C3525 vdd.n1775 gnd 0.010638f
C3526 vdd.n1776 gnd 0.902362f
C3527 vdd.t134 gnd 0.543592f
C3528 vdd.n1777 gnd 0.581643f
C3529 vdd.n1778 gnd 0.010638f
C3530 vdd.n1779 gnd 0.008563f
C3531 vdd.n1780 gnd 0.010638f
C3532 vdd.n1781 gnd 0.010638f
C3533 vdd.n1782 gnd 0.010638f
C3534 vdd.n1783 gnd 0.008563f
C3535 vdd.n1784 gnd 0.010638f
C3536 vdd.n1785 gnd 0.690362f
C3537 vdd.n1786 gnd 0.010638f
C3538 vdd.n1787 gnd 0.008563f
C3539 vdd.n1788 gnd 0.010638f
C3540 vdd.n1789 gnd 0.010638f
C3541 vdd.n1790 gnd 0.010638f
C3542 vdd.n1791 gnd 0.008563f
C3543 vdd.n1792 gnd 0.010638f
C3544 vdd.n1793 gnd 0.570771f
C3545 vdd.n1794 gnd 0.875183f
C3546 vdd.n1795 gnd 0.010638f
C3547 vdd.n1796 gnd 0.008563f
C3548 vdd.n1797 gnd 0.010638f
C3549 vdd.n1798 gnd 0.010638f
C3550 vdd.n1799 gnd 0.010638f
C3551 vdd.n1800 gnd 0.008563f
C3552 vdd.n1801 gnd 0.010638f
C3553 vdd.n1802 gnd 1.06f
C3554 vdd.n1803 gnd 0.010638f
C3555 vdd.n1804 gnd 0.008563f
C3556 vdd.n1805 gnd 0.010638f
C3557 vdd.n1806 gnd 0.010638f
C3558 vdd.n1807 gnd 0.024226f
C3559 vdd.n1808 gnd 0.010638f
C3560 vdd.n1809 gnd 0.010638f
C3561 vdd.n1810 gnd 0.008563f
C3562 vdd.n1811 gnd 0.010638f
C3563 vdd.t192 gnd 0.543592f
C3564 vdd.n1812 gnd 1.02739f
C3565 vdd.n1813 gnd 0.010638f
C3566 vdd.n1814 gnd 0.008563f
C3567 vdd.n1815 gnd 0.010638f
C3568 vdd.n1816 gnd 0.010638f
C3569 vdd.n1817 gnd 0.009149f
C3570 vdd.n1818 gnd 0.008563f
C3571 vdd.n1820 gnd 0.010638f
C3572 vdd.n1822 gnd 0.008563f
C3573 vdd.n1823 gnd 0.010638f
C3574 vdd.n1824 gnd 0.008563f
C3575 vdd.n1826 gnd 0.010638f
C3576 vdd.n1827 gnd 0.008563f
C3577 vdd.n1828 gnd 0.010638f
C3578 vdd.n1829 gnd 0.010638f
C3579 vdd.n1830 gnd 0.010638f
C3580 vdd.n1831 gnd 0.010638f
C3581 vdd.n1832 gnd 0.010638f
C3582 vdd.n1833 gnd 0.008563f
C3583 vdd.n1835 gnd 0.010638f
C3584 vdd.n1836 gnd 0.010638f
C3585 vdd.n1837 gnd 0.010638f
C3586 vdd.n1838 gnd 0.010638f
C3587 vdd.n1839 gnd 0.010638f
C3588 vdd.n1840 gnd 0.008563f
C3589 vdd.n1842 gnd 0.010638f
C3590 vdd.n1843 gnd 0.010638f
C3591 vdd.n1844 gnd 0.010638f
C3592 vdd.n1845 gnd 0.010638f
C3593 vdd.n1846 gnd 0.00715f
C3594 vdd.t210 gnd 0.130879f
C3595 vdd.t209 gnd 0.139874f
C3596 vdd.t208 gnd 0.170926f
C3597 vdd.n1847 gnd 0.219103f
C3598 vdd.n1848 gnd 0.184086f
C3599 vdd.n1850 gnd 0.010638f
C3600 vdd.n1851 gnd 0.010638f
C3601 vdd.n1852 gnd 0.008563f
C3602 vdd.n1853 gnd 0.010638f
C3603 vdd.n1855 gnd 0.010638f
C3604 vdd.n1856 gnd 0.010638f
C3605 vdd.n1857 gnd 0.010638f
C3606 vdd.n1858 gnd 0.010638f
C3607 vdd.n1859 gnd 0.008563f
C3608 vdd.n1861 gnd 0.010638f
C3609 vdd.n1862 gnd 0.010638f
C3610 vdd.n1863 gnd 0.010638f
C3611 vdd.n1864 gnd 0.010638f
C3612 vdd.n1865 gnd 0.010638f
C3613 vdd.n1866 gnd 0.008563f
C3614 vdd.n1868 gnd 0.010638f
C3615 vdd.n1869 gnd 0.010638f
C3616 vdd.n1870 gnd 0.010638f
C3617 vdd.n1871 gnd 0.010638f
C3618 vdd.n1872 gnd 0.010638f
C3619 vdd.n1873 gnd 0.008563f
C3620 vdd.n1875 gnd 0.010638f
C3621 vdd.n1876 gnd 0.010638f
C3622 vdd.n1877 gnd 0.010638f
C3623 vdd.n1878 gnd 0.010638f
C3624 vdd.n1879 gnd 0.010638f
C3625 vdd.n1880 gnd 0.008563f
C3626 vdd.n1882 gnd 0.010638f
C3627 vdd.n1883 gnd 0.010638f
C3628 vdd.n1884 gnd 0.010638f
C3629 vdd.n1885 gnd 0.010638f
C3630 vdd.n1886 gnd 0.008477f
C3631 vdd.t207 gnd 0.130879f
C3632 vdd.t206 gnd 0.139874f
C3633 vdd.t205 gnd 0.170926f
C3634 vdd.n1887 gnd 0.219103f
C3635 vdd.n1888 gnd 0.184086f
C3636 vdd.n1890 gnd 0.010638f
C3637 vdd.n1891 gnd 0.010638f
C3638 vdd.n1892 gnd 0.008563f
C3639 vdd.n1893 gnd 0.010638f
C3640 vdd.n1895 gnd 0.010638f
C3641 vdd.n1896 gnd 0.010638f
C3642 vdd.n1897 gnd 0.010638f
C3643 vdd.n1898 gnd 0.010638f
C3644 vdd.n1899 gnd 0.008563f
C3645 vdd.n1901 gnd 0.010638f
C3646 vdd.n1902 gnd 0.010638f
C3647 vdd.n1903 gnd 0.010638f
C3648 vdd.n1904 gnd 0.010638f
C3649 vdd.n1905 gnd 0.010638f
C3650 vdd.n1906 gnd 0.008563f
C3651 vdd.n1908 gnd 0.010638f
C3652 vdd.n1909 gnd 0.010638f
C3653 vdd.n1910 gnd 0.010638f
C3654 vdd.n1911 gnd 0.010638f
C3655 vdd.n1912 gnd 0.010638f
C3656 vdd.n1913 gnd 0.010638f
C3657 vdd.n1914 gnd 0.008563f
C3658 vdd.n1916 gnd 0.010638f
C3659 vdd.n1918 gnd 0.010638f
C3660 vdd.n1919 gnd 0.008563f
C3661 vdd.n1920 gnd 0.008563f
C3662 vdd.n1921 gnd 0.010638f
C3663 vdd.n1923 gnd 0.010638f
C3664 vdd.n1924 gnd 0.008563f
C3665 vdd.n1925 gnd 0.008563f
C3666 vdd.n1926 gnd 0.010638f
C3667 vdd.n1928 gnd 0.010638f
C3668 vdd.n1929 gnd 0.010638f
C3669 vdd.n1930 gnd 0.008563f
C3670 vdd.n1931 gnd 0.008563f
C3671 vdd.n1932 gnd 0.008563f
C3672 vdd.n1933 gnd 0.010638f
C3673 vdd.n1935 gnd 0.010638f
C3674 vdd.n1936 gnd 0.010638f
C3675 vdd.n1937 gnd 0.008563f
C3676 vdd.n1938 gnd 0.008563f
C3677 vdd.n1939 gnd 0.008563f
C3678 vdd.n1940 gnd 0.010638f
C3679 vdd.n1942 gnd 0.010638f
C3680 vdd.n1943 gnd 0.010638f
C3681 vdd.n1944 gnd 0.008563f
C3682 vdd.n1945 gnd 0.008563f
C3683 vdd.n1946 gnd 0.008563f
C3684 vdd.n1947 gnd 0.010638f
C3685 vdd.n1949 gnd 0.010638f
C3686 vdd.n1950 gnd 0.010638f
C3687 vdd.n1951 gnd 0.008563f
C3688 vdd.n1952 gnd 0.010638f
C3689 vdd.n1953 gnd 0.010638f
C3690 vdd.n1954 gnd 0.010638f
C3691 vdd.n1955 gnd 0.017468f
C3692 vdd.n1956 gnd 0.005823f
C3693 vdd.n1957 gnd 0.008563f
C3694 vdd.n1958 gnd 0.010638f
C3695 vdd.n1960 gnd 0.010638f
C3696 vdd.n1961 gnd 0.010638f
C3697 vdd.n1962 gnd 0.008563f
C3698 vdd.n1963 gnd 0.008563f
C3699 vdd.n1964 gnd 0.008563f
C3700 vdd.n1965 gnd 0.010638f
C3701 vdd.n1967 gnd 0.010638f
C3702 vdd.n1968 gnd 0.010638f
C3703 vdd.n1969 gnd 0.008563f
C3704 vdd.n1970 gnd 0.008563f
C3705 vdd.n1971 gnd 0.008563f
C3706 vdd.n1972 gnd 0.010638f
C3707 vdd.n1974 gnd 0.010638f
C3708 vdd.n1975 gnd 0.010638f
C3709 vdd.n1976 gnd 0.008563f
C3710 vdd.n1977 gnd 0.008563f
C3711 vdd.n1978 gnd 0.008563f
C3712 vdd.n1979 gnd 0.010638f
C3713 vdd.n1981 gnd 0.010638f
C3714 vdd.n1982 gnd 0.010638f
C3715 vdd.n1983 gnd 0.008563f
C3716 vdd.n1984 gnd 0.008563f
C3717 vdd.n1985 gnd 0.008563f
C3718 vdd.n1986 gnd 0.010638f
C3719 vdd.n1988 gnd 0.010638f
C3720 vdd.n1989 gnd 0.010638f
C3721 vdd.n1990 gnd 0.008563f
C3722 vdd.n1991 gnd 0.010638f
C3723 vdd.n1992 gnd 0.010638f
C3724 vdd.n1993 gnd 0.010638f
C3725 vdd.n1994 gnd 0.017468f
C3726 vdd.n1995 gnd 0.00715f
C3727 vdd.n1996 gnd 0.008563f
C3728 vdd.n1997 gnd 0.010638f
C3729 vdd.n1999 gnd 0.010638f
C3730 vdd.n2000 gnd 0.010638f
C3731 vdd.n2001 gnd 0.008563f
C3732 vdd.n2002 gnd 0.008563f
C3733 vdd.n2003 gnd 0.008563f
C3734 vdd.n2004 gnd 0.010638f
C3735 vdd.n2006 gnd 0.010638f
C3736 vdd.n2007 gnd 0.010638f
C3737 vdd.n2008 gnd 0.008563f
C3738 vdd.n2009 gnd 0.008563f
C3739 vdd.n2010 gnd 0.008563f
C3740 vdd.n2011 gnd 0.010638f
C3741 vdd.n2013 gnd 0.010638f
C3742 vdd.n2014 gnd 0.010638f
C3743 vdd.n2016 gnd 0.010638f
C3744 vdd.n2017 gnd 0.008563f
C3745 vdd.n2018 gnd 0.006809f
C3746 vdd.n2019 gnd 0.007234f
C3747 vdd.n2020 gnd 0.007234f
C3748 vdd.n2021 gnd 0.007234f
C3749 vdd.n2022 gnd 0.007234f
C3750 vdd.n2023 gnd 0.007234f
C3751 vdd.n2024 gnd 0.007234f
C3752 vdd.n2025 gnd 0.007234f
C3753 vdd.n2026 gnd 0.007234f
C3754 vdd.n2028 gnd 0.007234f
C3755 vdd.n2029 gnd 0.007234f
C3756 vdd.n2030 gnd 0.007234f
C3757 vdd.n2031 gnd 0.007234f
C3758 vdd.n2032 gnd 0.007234f
C3759 vdd.n2034 gnd 0.007234f
C3760 vdd.n2036 gnd 0.007234f
C3761 vdd.n2037 gnd 0.007234f
C3762 vdd.n2038 gnd 0.007234f
C3763 vdd.n2039 gnd 0.007234f
C3764 vdd.n2040 gnd 0.007234f
C3765 vdd.n2042 gnd 0.007234f
C3766 vdd.n2044 gnd 0.007234f
C3767 vdd.n2045 gnd 0.007234f
C3768 vdd.n2046 gnd 0.007234f
C3769 vdd.n2047 gnd 0.007234f
C3770 vdd.n2048 gnd 0.007234f
C3771 vdd.n2050 gnd 0.007234f
C3772 vdd.n2052 gnd 0.007234f
C3773 vdd.n2053 gnd 0.007234f
C3774 vdd.n2054 gnd 0.007234f
C3775 vdd.n2055 gnd 0.007234f
C3776 vdd.n2056 gnd 0.007234f
C3777 vdd.n2058 gnd 0.007234f
C3778 vdd.n2059 gnd 0.007234f
C3779 vdd.n2060 gnd 0.007234f
C3780 vdd.n2061 gnd 0.007234f
C3781 vdd.n2062 gnd 0.007234f
C3782 vdd.n2063 gnd 0.007234f
C3783 vdd.n2064 gnd 0.007234f
C3784 vdd.n2065 gnd 0.007234f
C3785 vdd.n2066 gnd 0.005266f
C3786 vdd.n2067 gnd 0.007234f
C3787 vdd.t174 gnd 0.292327f
C3788 vdd.t175 gnd 0.299233f
C3789 vdd.t172 gnd 0.190842f
C3790 vdd.n2068 gnd 0.10314f
C3791 vdd.n2069 gnd 0.058504f
C3792 vdd.n2070 gnd 0.010339f
C3793 vdd.n2071 gnd 0.007234f
C3794 vdd.n2072 gnd 0.007234f
C3795 vdd.n2073 gnd 0.440309f
C3796 vdd.n2074 gnd 0.007234f
C3797 vdd.n2075 gnd 0.007234f
C3798 vdd.n2076 gnd 0.007234f
C3799 vdd.n2077 gnd 0.007234f
C3800 vdd.n2078 gnd 0.007234f
C3801 vdd.n2079 gnd 0.007234f
C3802 vdd.n2080 gnd 0.007234f
C3803 vdd.n2081 gnd 0.007234f
C3804 vdd.n2082 gnd 0.007234f
C3805 vdd.n2083 gnd 0.007234f
C3806 vdd.n2084 gnd 0.007234f
C3807 vdd.n2085 gnd 0.007234f
C3808 vdd.n2086 gnd 0.007234f
C3809 vdd.n2087 gnd 0.007234f
C3810 vdd.n2088 gnd 0.007234f
C3811 vdd.n2089 gnd 0.007234f
C3812 vdd.n2090 gnd 0.007234f
C3813 vdd.n2091 gnd 0.007234f
C3814 vdd.n2092 gnd 0.007234f
C3815 vdd.n2093 gnd 0.007234f
C3816 vdd.t227 gnd 0.292327f
C3817 vdd.t228 gnd 0.299233f
C3818 vdd.t226 gnd 0.190842f
C3819 vdd.n2094 gnd 0.10314f
C3820 vdd.n2095 gnd 0.058504f
C3821 vdd.n2096 gnd 0.007234f
C3822 vdd.n2097 gnd 0.007234f
C3823 vdd.n2098 gnd 0.007234f
C3824 vdd.n2099 gnd 0.007234f
C3825 vdd.n2100 gnd 0.007234f
C3826 vdd.n2101 gnd 0.007234f
C3827 vdd.n2103 gnd 0.007234f
C3828 vdd.n2104 gnd 0.007234f
C3829 vdd.n2105 gnd 0.007234f
C3830 vdd.n2106 gnd 0.007234f
C3831 vdd.n2108 gnd 0.007234f
C3832 vdd.n2110 gnd 0.007234f
C3833 vdd.n2111 gnd 0.007234f
C3834 vdd.n2112 gnd 0.007234f
C3835 vdd.n2113 gnd 0.007234f
C3836 vdd.n2114 gnd 0.007234f
C3837 vdd.n2116 gnd 0.007234f
C3838 vdd.n2118 gnd 0.007234f
C3839 vdd.n2119 gnd 0.007234f
C3840 vdd.n2120 gnd 0.007234f
C3841 vdd.n2121 gnd 0.007234f
C3842 vdd.n2122 gnd 0.007234f
C3843 vdd.n2124 gnd 0.007234f
C3844 vdd.n2126 gnd 0.007234f
C3845 vdd.n2127 gnd 0.007234f
C3846 vdd.n2128 gnd 0.005266f
C3847 vdd.n2129 gnd 0.010339f
C3848 vdd.n2130 gnd 0.005585f
C3849 vdd.n2131 gnd 0.007234f
C3850 vdd.n2133 gnd 0.007234f
C3851 vdd.n2134 gnd 0.017165f
C3852 vdd.n2135 gnd 0.017165f
C3853 vdd.n2136 gnd 0.016026f
C3854 vdd.n2137 gnd 0.007234f
C3855 vdd.n2138 gnd 0.007234f
C3856 vdd.n2139 gnd 0.007234f
C3857 vdd.n2140 gnd 0.007234f
C3858 vdd.n2141 gnd 0.007234f
C3859 vdd.n2142 gnd 0.007234f
C3860 vdd.n2143 gnd 0.007234f
C3861 vdd.n2144 gnd 0.007234f
C3862 vdd.n2145 gnd 0.007234f
C3863 vdd.n2146 gnd 0.007234f
C3864 vdd.n2147 gnd 0.007234f
C3865 vdd.n2148 gnd 0.007234f
C3866 vdd.n2149 gnd 0.007234f
C3867 vdd.n2150 gnd 0.007234f
C3868 vdd.n2151 gnd 0.007234f
C3869 vdd.n2152 gnd 0.007234f
C3870 vdd.n2153 gnd 0.007234f
C3871 vdd.n2154 gnd 0.007234f
C3872 vdd.n2155 gnd 0.007234f
C3873 vdd.n2156 gnd 0.007234f
C3874 vdd.n2157 gnd 0.007234f
C3875 vdd.n2158 gnd 0.007234f
C3876 vdd.n2159 gnd 0.007234f
C3877 vdd.n2160 gnd 0.007234f
C3878 vdd.n2161 gnd 0.007234f
C3879 vdd.n2162 gnd 0.007234f
C3880 vdd.n2163 gnd 0.007234f
C3881 vdd.n2164 gnd 0.007234f
C3882 vdd.n2165 gnd 0.007234f
C3883 vdd.n2166 gnd 0.007234f
C3884 vdd.n2167 gnd 0.007234f
C3885 vdd.n2168 gnd 0.007234f
C3886 vdd.n2169 gnd 0.007234f
C3887 vdd.n2170 gnd 0.007234f
C3888 vdd.n2171 gnd 0.007234f
C3889 vdd.n2172 gnd 0.007234f
C3890 vdd.n2173 gnd 0.007234f
C3891 vdd.n2174 gnd 0.233745f
C3892 vdd.n2175 gnd 0.007234f
C3893 vdd.n2176 gnd 0.007234f
C3894 vdd.n2177 gnd 0.007234f
C3895 vdd.n2178 gnd 0.007234f
C3896 vdd.n2179 gnd 0.007234f
C3897 vdd.n2180 gnd 0.007234f
C3898 vdd.n2181 gnd 0.007234f
C3899 vdd.n2182 gnd 0.007234f
C3900 vdd.n2183 gnd 0.007234f
C3901 vdd.n2184 gnd 0.007234f
C3902 vdd.n2185 gnd 0.007234f
C3903 vdd.n2186 gnd 0.007234f
C3904 vdd.n2187 gnd 0.007234f
C3905 vdd.n2188 gnd 0.007234f
C3906 vdd.n2189 gnd 0.007234f
C3907 vdd.n2190 gnd 0.007234f
C3908 vdd.n2191 gnd 0.007234f
C3909 vdd.n2192 gnd 0.007234f
C3910 vdd.n2193 gnd 0.007234f
C3911 vdd.n2194 gnd 0.007234f
C3912 vdd.n2195 gnd 0.016026f
C3913 vdd.n2197 gnd 0.017165f
C3914 vdd.n2198 gnd 0.017165f
C3915 vdd.n2199 gnd 0.007234f
C3916 vdd.n2200 gnd 0.005585f
C3917 vdd.n2201 gnd 0.007234f
C3918 vdd.n2203 gnd 0.007234f
C3919 vdd.n2205 gnd 0.007234f
C3920 vdd.n2206 gnd 0.007234f
C3921 vdd.n2207 gnd 0.007234f
C3922 vdd.n2208 gnd 0.007234f
C3923 vdd.n2209 gnd 0.007234f
C3924 vdd.n2211 gnd 0.007234f
C3925 vdd.n2213 gnd 0.007234f
C3926 vdd.n2214 gnd 0.007234f
C3927 vdd.n2215 gnd 0.007234f
C3928 vdd.n2216 gnd 0.007234f
C3929 vdd.n2217 gnd 0.007234f
C3930 vdd.n2219 gnd 0.007234f
C3931 vdd.n2221 gnd 0.007234f
C3932 vdd.n2222 gnd 0.007234f
C3933 vdd.n2223 gnd 0.007234f
C3934 vdd.n2224 gnd 0.007234f
C3935 vdd.n2225 gnd 0.007234f
C3936 vdd.n2227 gnd 0.007234f
C3937 vdd.n2229 gnd 0.007234f
C3938 vdd.n2230 gnd 0.007234f
C3939 vdd.n2231 gnd 0.021578f
C3940 vdd.n2232 gnd 0.639653f
C3941 vdd.n2234 gnd 0.008563f
C3942 vdd.n2235 gnd 0.008563f
C3943 vdd.n2236 gnd 0.010638f
C3944 vdd.n2238 gnd 0.010638f
C3945 vdd.n2239 gnd 0.010638f
C3946 vdd.n2240 gnd 0.008563f
C3947 vdd.n2241 gnd 0.007107f
C3948 vdd.n2242 gnd 0.024391f
C3949 vdd.n2243 gnd 0.024226f
C3950 vdd.n2244 gnd 0.007107f
C3951 vdd.n2245 gnd 0.024226f
C3952 vdd.n2246 gnd 1.43508f
C3953 vdd.n2247 gnd 0.024226f
C3954 vdd.n2248 gnd 0.024391f
C3955 vdd.n2249 gnd 0.004067f
C3956 vdd.t194 gnd 0.130879f
C3957 vdd.t193 gnd 0.139874f
C3958 vdd.t191 gnd 0.170926f
C3959 vdd.n2250 gnd 0.219103f
C3960 vdd.n2251 gnd 0.184086f
C3961 vdd.n2252 gnd 0.013186f
C3962 vdd.n2253 gnd 0.004495f
C3963 vdd.n2254 gnd 0.009149f
C3964 vdd.n2255 gnd 0.639653f
C3965 vdd.n2256 gnd 0.021578f
C3966 vdd.n2257 gnd 0.007234f
C3967 vdd.n2258 gnd 0.007234f
C3968 vdd.n2259 gnd 0.007234f
C3969 vdd.n2261 gnd 0.007234f
C3970 vdd.n2263 gnd 0.007234f
C3971 vdd.n2264 gnd 0.007234f
C3972 vdd.n2265 gnd 0.007234f
C3973 vdd.n2266 gnd 0.007234f
C3974 vdd.n2267 gnd 0.007234f
C3975 vdd.n2269 gnd 0.007234f
C3976 vdd.n2271 gnd 0.007234f
C3977 vdd.n2272 gnd 0.007234f
C3978 vdd.n2273 gnd 0.007234f
C3979 vdd.n2274 gnd 0.007234f
C3980 vdd.n2275 gnd 0.007234f
C3981 vdd.n2277 gnd 0.007234f
C3982 vdd.n2279 gnd 0.007234f
C3983 vdd.n2280 gnd 0.007234f
C3984 vdd.n2281 gnd 0.007234f
C3985 vdd.n2282 gnd 0.007234f
C3986 vdd.n2283 gnd 0.007234f
C3987 vdd.n2285 gnd 0.007234f
C3988 vdd.n2287 gnd 0.007234f
C3989 vdd.n2288 gnd 0.007234f
C3990 vdd.n2289 gnd 0.017165f
C3991 vdd.n2290 gnd 0.016026f
C3992 vdd.n2291 gnd 0.016026f
C3993 vdd.n2292 gnd 1.06544f
C3994 vdd.n2293 gnd 0.016026f
C3995 vdd.n2294 gnd 0.016026f
C3996 vdd.n2295 gnd 0.007234f
C3997 vdd.n2296 gnd 0.007234f
C3998 vdd.n2297 gnd 0.007234f
C3999 vdd.n2298 gnd 0.462053f
C4000 vdd.n2299 gnd 0.007234f
C4001 vdd.n2300 gnd 0.007234f
C4002 vdd.n2301 gnd 0.007234f
C4003 vdd.n2302 gnd 0.007234f
C4004 vdd.n2303 gnd 0.007234f
C4005 vdd.n2304 gnd 0.739285f
C4006 vdd.n2305 gnd 0.007234f
C4007 vdd.n2306 gnd 0.007234f
C4008 vdd.n2307 gnd 0.007234f
C4009 vdd.n2308 gnd 0.007234f
C4010 vdd.n2309 gnd 0.007234f
C4011 vdd.n2310 gnd 0.739285f
C4012 vdd.n2311 gnd 0.007234f
C4013 vdd.n2312 gnd 0.007234f
C4014 vdd.n2313 gnd 0.006383f
C4015 vdd.n2314 gnd 0.020956f
C4016 vdd.n2315 gnd 0.004468f
C4017 vdd.n2316 gnd 0.007234f
C4018 vdd.n2317 gnd 0.407694f
C4019 vdd.n2318 gnd 0.007234f
C4020 vdd.n2319 gnd 0.007234f
C4021 vdd.n2320 gnd 0.007234f
C4022 vdd.n2321 gnd 0.007234f
C4023 vdd.n2322 gnd 0.007234f
C4024 vdd.n2323 gnd 0.494669f
C4025 vdd.n2324 gnd 0.007234f
C4026 vdd.n2325 gnd 0.007234f
C4027 vdd.n2326 gnd 0.007234f
C4028 vdd.n2327 gnd 0.007234f
C4029 vdd.n2328 gnd 0.007234f
C4030 vdd.n2329 gnd 0.657746f
C4031 vdd.n2330 gnd 0.007234f
C4032 vdd.n2331 gnd 0.007234f
C4033 vdd.n2332 gnd 0.007234f
C4034 vdd.n2333 gnd 0.007234f
C4035 vdd.n2334 gnd 0.007234f
C4036 vdd.n2335 gnd 0.587079f
C4037 vdd.n2336 gnd 0.007234f
C4038 vdd.n2337 gnd 0.007234f
C4039 vdd.n2338 gnd 0.007234f
C4040 vdd.n2339 gnd 0.007234f
C4041 vdd.n2340 gnd 0.007234f
C4042 vdd.n2341 gnd 0.424002f
C4043 vdd.n2342 gnd 0.007234f
C4044 vdd.n2343 gnd 0.007234f
C4045 vdd.n2344 gnd 0.007234f
C4046 vdd.n2345 gnd 0.007234f
C4047 vdd.n2346 gnd 0.007234f
C4048 vdd.n2347 gnd 0.233745f
C4049 vdd.n2348 gnd 0.007234f
C4050 vdd.n2349 gnd 0.007234f
C4051 vdd.n2350 gnd 0.007234f
C4052 vdd.n2351 gnd 0.007234f
C4053 vdd.n2352 gnd 0.007234f
C4054 vdd.n2353 gnd 0.407694f
C4055 vdd.n2354 gnd 0.007234f
C4056 vdd.n2355 gnd 0.007234f
C4057 vdd.n2356 gnd 0.007234f
C4058 vdd.n2357 gnd 0.007234f
C4059 vdd.n2358 gnd 0.007234f
C4060 vdd.n2359 gnd 0.739285f
C4061 vdd.n2360 gnd 0.007234f
C4062 vdd.n2361 gnd 0.007234f
C4063 vdd.n2362 gnd 0.007234f
C4064 vdd.n2363 gnd 0.007234f
C4065 vdd.n2364 gnd 0.007234f
C4066 vdd.n2365 gnd 0.007234f
C4067 vdd.n2366 gnd 0.007234f
C4068 vdd.n2367 gnd 0.576207f
C4069 vdd.n2368 gnd 0.007234f
C4070 vdd.n2369 gnd 0.007234f
C4071 vdd.n2370 gnd 0.007234f
C4072 vdd.n2371 gnd 0.007234f
C4073 vdd.n2372 gnd 0.007234f
C4074 vdd.n2373 gnd 0.007234f
C4075 vdd.n2374 gnd 0.462053f
C4076 vdd.n2375 gnd 0.007234f
C4077 vdd.n2376 gnd 0.007234f
C4078 vdd.n2377 gnd 0.007234f
C4079 vdd.n2378 gnd 0.016907f
C4080 vdd.n2379 gnd 0.016284f
C4081 vdd.n2380 gnd 0.007234f
C4082 vdd.n2381 gnd 0.007234f
C4083 vdd.n2382 gnd 0.005585f
C4084 vdd.n2383 gnd 0.007234f
C4085 vdd.n2384 gnd 0.007234f
C4086 vdd.n2385 gnd 0.005266f
C4087 vdd.n2386 gnd 0.007234f
C4088 vdd.n2387 gnd 0.007234f
C4089 vdd.n2388 gnd 0.007234f
C4090 vdd.n2389 gnd 0.007234f
C4091 vdd.n2390 gnd 0.007234f
C4092 vdd.n2391 gnd 0.007234f
C4093 vdd.n2392 gnd 0.007234f
C4094 vdd.n2393 gnd 0.007234f
C4095 vdd.n2394 gnd 0.007234f
C4096 vdd.n2395 gnd 0.007234f
C4097 vdd.n2396 gnd 0.007234f
C4098 vdd.n2397 gnd 0.007234f
C4099 vdd.n2398 gnd 0.007234f
C4100 vdd.n2399 gnd 0.007234f
C4101 vdd.n2400 gnd 0.007234f
C4102 vdd.n2401 gnd 0.007234f
C4103 vdd.n2402 gnd 0.007234f
C4104 vdd.n2403 gnd 0.007234f
C4105 vdd.n2404 gnd 0.007234f
C4106 vdd.n2405 gnd 0.007234f
C4107 vdd.n2406 gnd 0.007234f
C4108 vdd.n2407 gnd 0.007234f
C4109 vdd.n2408 gnd 0.007234f
C4110 vdd.n2409 gnd 0.007234f
C4111 vdd.n2410 gnd 0.007234f
C4112 vdd.n2411 gnd 0.007234f
C4113 vdd.n2412 gnd 0.007234f
C4114 vdd.n2413 gnd 0.007234f
C4115 vdd.n2414 gnd 0.007234f
C4116 vdd.n2415 gnd 0.007234f
C4117 vdd.n2416 gnd 0.007234f
C4118 vdd.n2417 gnd 0.007234f
C4119 vdd.n2418 gnd 0.007234f
C4120 vdd.n2419 gnd 0.007234f
C4121 vdd.n2420 gnd 0.007234f
C4122 vdd.n2421 gnd 0.007234f
C4123 vdd.n2422 gnd 0.007234f
C4124 vdd.n2423 gnd 0.007234f
C4125 vdd.n2424 gnd 0.007234f
C4126 vdd.n2425 gnd 0.007234f
C4127 vdd.n2426 gnd 0.007234f
C4128 vdd.n2427 gnd 0.007234f
C4129 vdd.n2428 gnd 0.007234f
C4130 vdd.n2429 gnd 0.007234f
C4131 vdd.n2430 gnd 0.007234f
C4132 vdd.n2431 gnd 0.007234f
C4133 vdd.n2432 gnd 0.007234f
C4134 vdd.n2433 gnd 0.007234f
C4135 vdd.n2434 gnd 0.007234f
C4136 vdd.n2435 gnd 0.007234f
C4137 vdd.n2436 gnd 0.007234f
C4138 vdd.n2437 gnd 0.007234f
C4139 vdd.n2438 gnd 0.007234f
C4140 vdd.n2439 gnd 0.007234f
C4141 vdd.n2440 gnd 0.007234f
C4142 vdd.n2441 gnd 0.007234f
C4143 vdd.n2442 gnd 0.007234f
C4144 vdd.n2443 gnd 0.007234f
C4145 vdd.n2444 gnd 0.007234f
C4146 vdd.n2445 gnd 0.007234f
C4147 vdd.n2446 gnd 0.017165f
C4148 vdd.n2447 gnd 0.016026f
C4149 vdd.n2448 gnd 0.016026f
C4150 vdd.n2449 gnd 0.902362f
C4151 vdd.n2450 gnd 0.016026f
C4152 vdd.n2451 gnd 0.017165f
C4153 vdd.n2452 gnd 0.016284f
C4154 vdd.n2453 gnd 0.007234f
C4155 vdd.n2454 gnd 0.007234f
C4156 vdd.n2455 gnd 0.007234f
C4157 vdd.n2456 gnd 0.005585f
C4158 vdd.n2457 gnd 0.010339f
C4159 vdd.n2458 gnd 0.005266f
C4160 vdd.n2459 gnd 0.007234f
C4161 vdd.n2460 gnd 0.007234f
C4162 vdd.n2461 gnd 0.007234f
C4163 vdd.n2462 gnd 0.007234f
C4164 vdd.n2463 gnd 0.007234f
C4165 vdd.n2464 gnd 0.007234f
C4166 vdd.n2465 gnd 0.007234f
C4167 vdd.n2466 gnd 0.007234f
C4168 vdd.n2467 gnd 0.007234f
C4169 vdd.n2468 gnd 0.007234f
C4170 vdd.n2469 gnd 0.007234f
C4171 vdd.n2470 gnd 0.007234f
C4172 vdd.n2471 gnd 0.007234f
C4173 vdd.n2472 gnd 0.007234f
C4174 vdd.n2473 gnd 0.007234f
C4175 vdd.n2474 gnd 0.007234f
C4176 vdd.n2475 gnd 0.007234f
C4177 vdd.n2476 gnd 0.007234f
C4178 vdd.n2477 gnd 0.007234f
C4179 vdd.n2478 gnd 0.007234f
C4180 vdd.n2479 gnd 0.007234f
C4181 vdd.n2480 gnd 0.007234f
C4182 vdd.n2481 gnd 0.007234f
C4183 vdd.n2482 gnd 0.007234f
C4184 vdd.n2483 gnd 0.007234f
C4185 vdd.n2484 gnd 0.007234f
C4186 vdd.n2485 gnd 0.007234f
C4187 vdd.n2486 gnd 0.007234f
C4188 vdd.n2487 gnd 0.007234f
C4189 vdd.n2488 gnd 0.007234f
C4190 vdd.n2489 gnd 0.007234f
C4191 vdd.n2490 gnd 0.007234f
C4192 vdd.n2491 gnd 0.007234f
C4193 vdd.n2492 gnd 0.007234f
C4194 vdd.n2493 gnd 0.007234f
C4195 vdd.n2494 gnd 0.007234f
C4196 vdd.n2495 gnd 0.007234f
C4197 vdd.n2496 gnd 0.007234f
C4198 vdd.n2497 gnd 0.007234f
C4199 vdd.n2498 gnd 0.007234f
C4200 vdd.n2499 gnd 0.007234f
C4201 vdd.n2500 gnd 0.007234f
C4202 vdd.n2501 gnd 0.007234f
C4203 vdd.n2502 gnd 0.007234f
C4204 vdd.n2503 gnd 0.007234f
C4205 vdd.n2504 gnd 0.007234f
C4206 vdd.n2505 gnd 0.007234f
C4207 vdd.n2506 gnd 0.007234f
C4208 vdd.n2507 gnd 0.007234f
C4209 vdd.n2508 gnd 0.007234f
C4210 vdd.n2509 gnd 0.007234f
C4211 vdd.n2510 gnd 0.007234f
C4212 vdd.n2511 gnd 0.007234f
C4213 vdd.n2512 gnd 0.007234f
C4214 vdd.n2513 gnd 0.007234f
C4215 vdd.n2514 gnd 0.007234f
C4216 vdd.n2515 gnd 0.007234f
C4217 vdd.n2516 gnd 0.007234f
C4218 vdd.n2517 gnd 0.007234f
C4219 vdd.n2518 gnd 0.007234f
C4220 vdd.n2519 gnd 0.017165f
C4221 vdd.n2520 gnd 0.017165f
C4222 vdd.n2521 gnd 0.902362f
C4223 vdd.t248 gnd 3.20719f
C4224 vdd.t19 gnd 3.20719f
C4225 vdd.n2554 gnd 0.017165f
C4226 vdd.n2555 gnd 0.007234f
C4227 vdd.t221 gnd 0.292327f
C4228 vdd.t222 gnd 0.299233f
C4229 vdd.t219 gnd 0.190842f
C4230 vdd.n2556 gnd 0.10314f
C4231 vdd.n2557 gnd 0.058504f
C4232 vdd.n2558 gnd 0.007234f
C4233 vdd.t234 gnd 0.292327f
C4234 vdd.t235 gnd 0.299233f
C4235 vdd.t233 gnd 0.190842f
C4236 vdd.n2559 gnd 0.10314f
C4237 vdd.n2560 gnd 0.058504f
C4238 vdd.n2561 gnd 0.010339f
C4239 vdd.n2562 gnd 0.007234f
C4240 vdd.n2563 gnd 0.007234f
C4241 vdd.n2564 gnd 0.007234f
C4242 vdd.n2565 gnd 0.007234f
C4243 vdd.n2566 gnd 0.007234f
C4244 vdd.n2567 gnd 0.007234f
C4245 vdd.n2568 gnd 0.007234f
C4246 vdd.n2569 gnd 0.007234f
C4247 vdd.n2570 gnd 0.007234f
C4248 vdd.n2571 gnd 0.007234f
C4249 vdd.n2572 gnd 0.007234f
C4250 vdd.n2573 gnd 0.007234f
C4251 vdd.n2574 gnd 0.007234f
C4252 vdd.n2575 gnd 0.007234f
C4253 vdd.n2576 gnd 0.007234f
C4254 vdd.n2577 gnd 0.007234f
C4255 vdd.n2578 gnd 0.007234f
C4256 vdd.n2579 gnd 0.007234f
C4257 vdd.n2580 gnd 0.007234f
C4258 vdd.n2581 gnd 0.007234f
C4259 vdd.n2582 gnd 0.007234f
C4260 vdd.n2583 gnd 0.007234f
C4261 vdd.n2584 gnd 0.007234f
C4262 vdd.n2585 gnd 0.007234f
C4263 vdd.n2586 gnd 0.007234f
C4264 vdd.n2587 gnd 0.007234f
C4265 vdd.n2588 gnd 0.007234f
C4266 vdd.n2589 gnd 0.007234f
C4267 vdd.n2590 gnd 0.007234f
C4268 vdd.n2591 gnd 0.007234f
C4269 vdd.n2592 gnd 0.007234f
C4270 vdd.n2593 gnd 0.007234f
C4271 vdd.n2594 gnd 0.007234f
C4272 vdd.n2595 gnd 0.007234f
C4273 vdd.n2596 gnd 0.007234f
C4274 vdd.n2597 gnd 0.007234f
C4275 vdd.n2598 gnd 0.007234f
C4276 vdd.n2599 gnd 0.007234f
C4277 vdd.n2600 gnd 0.007234f
C4278 vdd.n2601 gnd 0.007234f
C4279 vdd.n2602 gnd 0.007234f
C4280 vdd.n2603 gnd 0.007234f
C4281 vdd.n2604 gnd 0.007234f
C4282 vdd.n2605 gnd 0.007234f
C4283 vdd.n2606 gnd 0.007234f
C4284 vdd.n2607 gnd 0.007234f
C4285 vdd.n2608 gnd 0.007234f
C4286 vdd.n2609 gnd 0.007234f
C4287 vdd.n2610 gnd 0.007234f
C4288 vdd.n2611 gnd 0.007234f
C4289 vdd.n2612 gnd 0.007234f
C4290 vdd.n2613 gnd 0.007234f
C4291 vdd.n2614 gnd 0.007234f
C4292 vdd.n2615 gnd 0.007234f
C4293 vdd.n2616 gnd 0.007234f
C4294 vdd.n2617 gnd 0.007234f
C4295 vdd.n2618 gnd 0.005266f
C4296 vdd.n2619 gnd 0.007234f
C4297 vdd.n2620 gnd 0.007234f
C4298 vdd.n2621 gnd 0.005585f
C4299 vdd.n2622 gnd 0.007234f
C4300 vdd.n2623 gnd 0.007234f
C4301 vdd.n2624 gnd 0.017165f
C4302 vdd.n2625 gnd 0.016026f
C4303 vdd.n2626 gnd 0.007234f
C4304 vdd.n2627 gnd 0.007234f
C4305 vdd.n2628 gnd 0.007234f
C4306 vdd.n2629 gnd 0.007234f
C4307 vdd.n2630 gnd 0.007234f
C4308 vdd.n2631 gnd 0.007234f
C4309 vdd.n2632 gnd 0.007234f
C4310 vdd.n2633 gnd 0.007234f
C4311 vdd.n2634 gnd 0.007234f
C4312 vdd.n2635 gnd 0.007234f
C4313 vdd.n2636 gnd 0.007234f
C4314 vdd.n2637 gnd 0.007234f
C4315 vdd.n2638 gnd 0.007234f
C4316 vdd.n2639 gnd 0.007234f
C4317 vdd.n2640 gnd 0.007234f
C4318 vdd.n2641 gnd 0.007234f
C4319 vdd.n2642 gnd 0.007234f
C4320 vdd.n2643 gnd 0.007234f
C4321 vdd.n2644 gnd 0.007234f
C4322 vdd.n2645 gnd 0.007234f
C4323 vdd.n2646 gnd 0.007234f
C4324 vdd.n2647 gnd 0.007234f
C4325 vdd.n2648 gnd 0.007234f
C4326 vdd.n2649 gnd 0.007234f
C4327 vdd.n2650 gnd 0.007234f
C4328 vdd.n2651 gnd 0.007234f
C4329 vdd.n2652 gnd 0.007234f
C4330 vdd.n2653 gnd 0.007234f
C4331 vdd.n2654 gnd 0.007234f
C4332 vdd.n2655 gnd 0.007234f
C4333 vdd.n2656 gnd 0.007234f
C4334 vdd.n2657 gnd 0.007234f
C4335 vdd.n2658 gnd 0.007234f
C4336 vdd.n2659 gnd 0.007234f
C4337 vdd.n2660 gnd 0.007234f
C4338 vdd.n2661 gnd 0.007234f
C4339 vdd.n2662 gnd 0.007234f
C4340 vdd.n2663 gnd 0.007234f
C4341 vdd.n2664 gnd 0.007234f
C4342 vdd.n2665 gnd 0.007234f
C4343 vdd.n2666 gnd 0.007234f
C4344 vdd.n2667 gnd 0.007234f
C4345 vdd.n2668 gnd 0.007234f
C4346 vdd.n2669 gnd 0.007234f
C4347 vdd.n2670 gnd 0.007234f
C4348 vdd.n2671 gnd 0.007234f
C4349 vdd.n2672 gnd 0.007234f
C4350 vdd.n2673 gnd 0.007234f
C4351 vdd.n2674 gnd 0.007234f
C4352 vdd.n2675 gnd 0.007234f
C4353 vdd.n2676 gnd 0.007234f
C4354 vdd.n2677 gnd 0.233745f
C4355 vdd.n2678 gnd 0.007234f
C4356 vdd.n2679 gnd 0.007234f
C4357 vdd.n2680 gnd 0.007234f
C4358 vdd.n2681 gnd 0.007234f
C4359 vdd.n2682 gnd 0.007234f
C4360 vdd.n2683 gnd 0.007234f
C4361 vdd.n2684 gnd 0.007234f
C4362 vdd.n2685 gnd 0.007234f
C4363 vdd.n2686 gnd 0.007234f
C4364 vdd.n2687 gnd 0.007234f
C4365 vdd.n2688 gnd 0.007234f
C4366 vdd.n2689 gnd 0.007234f
C4367 vdd.n2690 gnd 0.007234f
C4368 vdd.n2691 gnd 0.007234f
C4369 vdd.n2692 gnd 0.007234f
C4370 vdd.n2693 gnd 0.007234f
C4371 vdd.n2694 gnd 0.007234f
C4372 vdd.n2695 gnd 0.007234f
C4373 vdd.n2696 gnd 0.007234f
C4374 vdd.n2697 gnd 0.007234f
C4375 vdd.n2698 gnd 0.440309f
C4376 vdd.n2699 gnd 0.007234f
C4377 vdd.n2700 gnd 0.007234f
C4378 vdd.n2701 gnd 0.007234f
C4379 vdd.n2702 gnd 0.007234f
C4380 vdd.n2703 gnd 0.007234f
C4381 vdd.n2704 gnd 0.016026f
C4382 vdd.n2705 gnd 0.017165f
C4383 vdd.n2706 gnd 0.017165f
C4384 vdd.n2707 gnd 0.007234f
C4385 vdd.n2708 gnd 0.007234f
C4386 vdd.n2709 gnd 0.007234f
C4387 vdd.n2710 gnd 0.005585f
C4388 vdd.n2711 gnd 0.010339f
C4389 vdd.n2712 gnd 0.005266f
C4390 vdd.n2713 gnd 0.007234f
C4391 vdd.n2714 gnd 0.007234f
C4392 vdd.n2715 gnd 0.007234f
C4393 vdd.n2716 gnd 0.007234f
C4394 vdd.n2717 gnd 0.007234f
C4395 vdd.n2718 gnd 0.007234f
C4396 vdd.n2719 gnd 0.007234f
C4397 vdd.n2720 gnd 0.007234f
C4398 vdd.n2721 gnd 0.007234f
C4399 vdd.n2722 gnd 0.007234f
C4400 vdd.n2723 gnd 0.007234f
C4401 vdd.n2724 gnd 0.007234f
C4402 vdd.n2725 gnd 0.007234f
C4403 vdd.n2726 gnd 0.007234f
C4404 vdd.n2727 gnd 0.007234f
C4405 vdd.n2728 gnd 0.007234f
C4406 vdd.n2729 gnd 0.007234f
C4407 vdd.n2730 gnd 0.007234f
C4408 vdd.n2731 gnd 0.007234f
C4409 vdd.n2732 gnd 0.007234f
C4410 vdd.n2733 gnd 0.007234f
C4411 vdd.n2734 gnd 0.007234f
C4412 vdd.n2735 gnd 0.007234f
C4413 vdd.n2736 gnd 0.007234f
C4414 vdd.n2737 gnd 0.007234f
C4415 vdd.n2738 gnd 0.007234f
C4416 vdd.n2739 gnd 0.007234f
C4417 vdd.n2740 gnd 0.007234f
C4418 vdd.n2741 gnd 0.007234f
C4419 vdd.n2742 gnd 0.007234f
C4420 vdd.n2743 gnd 0.007234f
C4421 vdd.n2744 gnd 0.007234f
C4422 vdd.n2745 gnd 0.007234f
C4423 vdd.n2746 gnd 0.007234f
C4424 vdd.n2747 gnd 0.007234f
C4425 vdd.n2748 gnd 0.007234f
C4426 vdd.n2749 gnd 0.007234f
C4427 vdd.n2750 gnd 0.007234f
C4428 vdd.n2751 gnd 0.007234f
C4429 vdd.n2752 gnd 0.007234f
C4430 vdd.n2753 gnd 0.007234f
C4431 vdd.n2754 gnd 0.007234f
C4432 vdd.n2755 gnd 0.007234f
C4433 vdd.n2756 gnd 0.007234f
C4434 vdd.n2757 gnd 0.007234f
C4435 vdd.n2758 gnd 0.007234f
C4436 vdd.n2759 gnd 0.007234f
C4437 vdd.n2760 gnd 0.007234f
C4438 vdd.n2761 gnd 0.007234f
C4439 vdd.n2762 gnd 0.007234f
C4440 vdd.n2763 gnd 0.007234f
C4441 vdd.n2764 gnd 0.007234f
C4442 vdd.n2765 gnd 0.007234f
C4443 vdd.n2766 gnd 0.007234f
C4444 vdd.n2767 gnd 0.007234f
C4445 vdd.n2768 gnd 0.007234f
C4446 vdd.n2769 gnd 0.007234f
C4447 vdd.n2770 gnd 0.007234f
C4448 vdd.n2771 gnd 0.007234f
C4449 vdd.n2772 gnd 0.007234f
C4450 vdd.n2774 gnd 0.902362f
C4451 vdd.n2776 gnd 0.007234f
C4452 vdd.n2777 gnd 0.007234f
C4453 vdd.n2778 gnd 0.017165f
C4454 vdd.n2779 gnd 0.016026f
C4455 vdd.n2780 gnd 0.016026f
C4456 vdd.n2781 gnd 0.902362f
C4457 vdd.n2782 gnd 0.016026f
C4458 vdd.n2783 gnd 0.016026f
C4459 vdd.n2784 gnd 0.007234f
C4460 vdd.n2785 gnd 0.007234f
C4461 vdd.n2786 gnd 0.007234f
C4462 vdd.n2787 gnd 0.462053f
C4463 vdd.n2788 gnd 0.007234f
C4464 vdd.n2789 gnd 0.007234f
C4465 vdd.n2790 gnd 0.007234f
C4466 vdd.n2791 gnd 0.007234f
C4467 vdd.n2792 gnd 0.007234f
C4468 vdd.n2793 gnd 0.576207f
C4469 vdd.n2794 gnd 0.007234f
C4470 vdd.n2795 gnd 0.007234f
C4471 vdd.n2796 gnd 0.007234f
C4472 vdd.n2797 gnd 0.007234f
C4473 vdd.n2798 gnd 0.007234f
C4474 vdd.n2799 gnd 0.739285f
C4475 vdd.n2800 gnd 0.007234f
C4476 vdd.n2801 gnd 0.007234f
C4477 vdd.n2802 gnd 0.007234f
C4478 vdd.n2803 gnd 0.007234f
C4479 vdd.n2804 gnd 0.007234f
C4480 vdd.n2805 gnd 0.407694f
C4481 vdd.n2806 gnd 0.007234f
C4482 vdd.n2807 gnd 0.007234f
C4483 vdd.n2808 gnd 0.007234f
C4484 vdd.n2809 gnd 0.007234f
C4485 vdd.n2810 gnd 0.007234f
C4486 vdd.n2811 gnd 0.233745f
C4487 vdd.n2812 gnd 0.007234f
C4488 vdd.n2813 gnd 0.007234f
C4489 vdd.n2814 gnd 0.007234f
C4490 vdd.n2815 gnd 0.007234f
C4491 vdd.n2816 gnd 0.007234f
C4492 vdd.n2817 gnd 0.424002f
C4493 vdd.n2818 gnd 0.007234f
C4494 vdd.n2819 gnd 0.007234f
C4495 vdd.n2820 gnd 0.007234f
C4496 vdd.n2821 gnd 0.007234f
C4497 vdd.n2822 gnd 0.007234f
C4498 vdd.n2823 gnd 0.587079f
C4499 vdd.n2824 gnd 0.007234f
C4500 vdd.n2825 gnd 0.007234f
C4501 vdd.n2826 gnd 0.007234f
C4502 vdd.n2827 gnd 0.007234f
C4503 vdd.n2828 gnd 0.007234f
C4504 vdd.n2829 gnd 0.657746f
C4505 vdd.n2830 gnd 0.007234f
C4506 vdd.n2831 gnd 0.007234f
C4507 vdd.n2832 gnd 0.007234f
C4508 vdd.n2833 gnd 0.007234f
C4509 vdd.n2834 gnd 0.007234f
C4510 vdd.n2835 gnd 0.494669f
C4511 vdd.n2836 gnd 0.007234f
C4512 vdd.n2837 gnd 0.007234f
C4513 vdd.n2838 gnd 0.007234f
C4514 vdd.t200 gnd 0.299233f
C4515 vdd.t198 gnd 0.190842f
C4516 vdd.t201 gnd 0.299233f
C4517 vdd.n2839 gnd 0.168181f
C4518 vdd.n2840 gnd 0.020956f
C4519 vdd.n2841 gnd 0.004468f
C4520 vdd.n2842 gnd 0.007234f
C4521 vdd.n2843 gnd 0.407694f
C4522 vdd.n2844 gnd 0.007234f
C4523 vdd.n2845 gnd 0.007234f
C4524 vdd.n2846 gnd 0.007234f
C4525 vdd.n2847 gnd 0.007234f
C4526 vdd.n2848 gnd 0.007234f
C4527 vdd.n2849 gnd 0.739285f
C4528 vdd.n2850 gnd 0.007234f
C4529 vdd.n2851 gnd 0.007234f
C4530 vdd.n2852 gnd 0.007234f
C4531 vdd.n2853 gnd 0.007234f
C4532 vdd.n2854 gnd 0.007234f
C4533 vdd.n2855 gnd 0.007234f
C4534 vdd.n2857 gnd 0.007234f
C4535 vdd.n2858 gnd 0.007234f
C4536 vdd.n2860 gnd 0.007234f
C4537 vdd.n2861 gnd 0.007234f
C4538 vdd.n2864 gnd 0.007234f
C4539 vdd.n2865 gnd 0.007234f
C4540 vdd.n2866 gnd 0.007234f
C4541 vdd.n2867 gnd 0.007234f
C4542 vdd.n2869 gnd 0.007234f
C4543 vdd.n2870 gnd 0.007234f
C4544 vdd.n2871 gnd 0.007234f
C4545 vdd.n2872 gnd 0.007234f
C4546 vdd.n2873 gnd 0.007234f
C4547 vdd.n2874 gnd 0.007234f
C4548 vdd.n2876 gnd 0.007234f
C4549 vdd.n2877 gnd 0.007234f
C4550 vdd.n2878 gnd 0.007234f
C4551 vdd.n2879 gnd 0.007234f
C4552 vdd.n2880 gnd 0.007234f
C4553 vdd.n2881 gnd 0.007234f
C4554 vdd.n2883 gnd 0.007234f
C4555 vdd.n2884 gnd 0.007234f
C4556 vdd.n2885 gnd 0.007234f
C4557 vdd.n2886 gnd 0.007234f
C4558 vdd.n2887 gnd 0.007234f
C4559 vdd.n2888 gnd 0.007234f
C4560 vdd.n2890 gnd 0.007234f
C4561 vdd.n2891 gnd 0.017165f
C4562 vdd.n2892 gnd 0.017165f
C4563 vdd.n2893 gnd 0.016026f
C4564 vdd.n2894 gnd 0.007234f
C4565 vdd.n2895 gnd 0.007234f
C4566 vdd.n2896 gnd 0.007234f
C4567 vdd.n2897 gnd 0.007234f
C4568 vdd.n2898 gnd 0.007234f
C4569 vdd.n2899 gnd 0.007234f
C4570 vdd.n2900 gnd 0.739285f
C4571 vdd.n2901 gnd 0.007234f
C4572 vdd.n2902 gnd 0.007234f
C4573 vdd.n2903 gnd 0.007234f
C4574 vdd.n2904 gnd 0.007234f
C4575 vdd.n2905 gnd 0.007234f
C4576 vdd.n2906 gnd 0.462053f
C4577 vdd.n2907 gnd 0.007234f
C4578 vdd.n2908 gnd 0.007234f
C4579 vdd.n2909 gnd 0.007234f
C4580 vdd.n2910 gnd 0.016907f
C4581 vdd.n2912 gnd 0.017165f
C4582 vdd.n2913 gnd 0.016284f
C4583 vdd.n2914 gnd 0.007234f
C4584 vdd.n2915 gnd 0.005585f
C4585 vdd.n2916 gnd 0.007234f
C4586 vdd.n2918 gnd 0.007234f
C4587 vdd.n2919 gnd 0.007234f
C4588 vdd.n2920 gnd 0.007234f
C4589 vdd.n2921 gnd 0.007234f
C4590 vdd.n2922 gnd 0.007234f
C4591 vdd.n2923 gnd 0.007234f
C4592 vdd.n2925 gnd 0.007234f
C4593 vdd.n2926 gnd 0.007234f
C4594 vdd.n2927 gnd 0.007234f
C4595 vdd.n2928 gnd 0.007234f
C4596 vdd.n2929 gnd 0.007234f
C4597 vdd.n2930 gnd 0.007234f
C4598 vdd.n2932 gnd 0.007234f
C4599 vdd.n2933 gnd 0.007234f
C4600 vdd.n2934 gnd 0.007234f
C4601 vdd.n2935 gnd 0.007234f
C4602 vdd.n2936 gnd 0.007234f
C4603 vdd.n2937 gnd 0.007234f
C4604 vdd.n2939 gnd 0.007234f
C4605 vdd.n2940 gnd 0.007234f
C4606 vdd.n2941 gnd 0.007234f
C4607 vdd.n2942 gnd 0.643847f
C4608 vdd.n2943 gnd 0.017384f
C4609 vdd.n2944 gnd 0.007234f
C4610 vdd.n2945 gnd 0.007234f
C4611 vdd.n2947 gnd 0.007234f
C4612 vdd.n2948 gnd 0.007234f
C4613 vdd.n2949 gnd 0.007234f
C4614 vdd.n2950 gnd 0.007234f
C4615 vdd.n2951 gnd 0.007234f
C4616 vdd.n2952 gnd 0.007234f
C4617 vdd.n2954 gnd 0.007234f
C4618 vdd.n2955 gnd 0.007234f
C4619 vdd.n2956 gnd 0.007234f
C4620 vdd.n2957 gnd 0.007234f
C4621 vdd.n2958 gnd 0.007234f
C4622 vdd.n2959 gnd 0.007234f
C4623 vdd.n2961 gnd 0.007234f
C4624 vdd.n2962 gnd 0.007234f
C4625 vdd.n2963 gnd 0.007234f
C4626 vdd.n2964 gnd 0.007234f
C4627 vdd.n2965 gnd 0.007234f
C4628 vdd.n2966 gnd 0.007234f
C4629 vdd.n2968 gnd 0.007234f
C4630 vdd.n2969 gnd 0.007234f
C4631 vdd.n2971 gnd 0.007234f
C4632 vdd.n2972 gnd 0.007234f
C4633 vdd.n2973 gnd 0.017165f
C4634 vdd.n2974 gnd 0.016026f
C4635 vdd.n2975 gnd 0.016026f
C4636 vdd.n2976 gnd 1.06544f
C4637 vdd.n2977 gnd 0.016026f
C4638 vdd.n2978 gnd 0.017165f
C4639 vdd.n2979 gnd 0.016284f
C4640 vdd.n2980 gnd 0.007234f
C4641 vdd.n2981 gnd 0.005585f
C4642 vdd.n2982 gnd 0.007234f
C4643 vdd.n2984 gnd 0.007234f
C4644 vdd.n2985 gnd 0.007234f
C4645 vdd.n2986 gnd 0.007234f
C4646 vdd.n2987 gnd 0.007234f
C4647 vdd.n2988 gnd 0.007234f
C4648 vdd.n2989 gnd 0.007234f
C4649 vdd.n2991 gnd 0.007234f
C4650 vdd.n2992 gnd 0.007234f
C4651 vdd.n2993 gnd 0.007234f
C4652 vdd.n2994 gnd 0.007234f
C4653 vdd.n2995 gnd 0.007234f
C4654 vdd.n2996 gnd 0.007234f
C4655 vdd.n2998 gnd 0.007234f
C4656 vdd.n2999 gnd 0.007234f
C4657 vdd.n3000 gnd 0.007234f
C4658 vdd.n3001 gnd 0.007234f
C4659 vdd.n3002 gnd 0.007234f
C4660 vdd.n3003 gnd 0.007234f
C4661 vdd.n3005 gnd 0.007234f
C4662 vdd.n3006 gnd 0.007234f
C4663 vdd.n3008 gnd 0.007234f
C4664 vdd.n3009 gnd 0.017384f
C4665 vdd.n3010 gnd 0.643847f
C4666 vdd.n3011 gnd 0.009149f
C4667 vdd.n3012 gnd 0.004067f
C4668 vdd.t243 gnd 0.130879f
C4669 vdd.t244 gnd 0.139874f
C4670 vdd.t242 gnd 0.170926f
C4671 vdd.n3013 gnd 0.219103f
C4672 vdd.n3014 gnd 0.184086f
C4673 vdd.n3015 gnd 0.013186f
C4674 vdd.n3016 gnd 0.010638f
C4675 vdd.n3017 gnd 0.004495f
C4676 vdd.n3018 gnd 0.008563f
C4677 vdd.n3019 gnd 0.010638f
C4678 vdd.n3020 gnd 0.010638f
C4679 vdd.n3021 gnd 0.008563f
C4680 vdd.n3022 gnd 0.008563f
C4681 vdd.n3023 gnd 0.010638f
C4682 vdd.n3025 gnd 0.010638f
C4683 vdd.n3026 gnd 0.008563f
C4684 vdd.n3027 gnd 0.008563f
C4685 vdd.n3028 gnd 0.008563f
C4686 vdd.n3029 gnd 0.010638f
C4687 vdd.n3031 gnd 0.010638f
C4688 vdd.n3033 gnd 0.010638f
C4689 vdd.n3034 gnd 0.008563f
C4690 vdd.n3035 gnd 0.008563f
C4691 vdd.n3036 gnd 0.008563f
C4692 vdd.n3037 gnd 0.010638f
C4693 vdd.n3039 gnd 0.010638f
C4694 vdd.n3041 gnd 0.010638f
C4695 vdd.n3042 gnd 0.008563f
C4696 vdd.n3043 gnd 0.008563f
C4697 vdd.n3044 gnd 0.008563f
C4698 vdd.n3045 gnd 0.010638f
C4699 vdd.n3047 gnd 0.010638f
C4700 vdd.n3048 gnd 0.010638f
C4701 vdd.n3049 gnd 0.008563f
C4702 vdd.n3050 gnd 0.008563f
C4703 vdd.n3051 gnd 0.010638f
C4704 vdd.n3052 gnd 0.010638f
C4705 vdd.n3054 gnd 0.010638f
C4706 vdd.n3055 gnd 0.008563f
C4707 vdd.n3056 gnd 0.010638f
C4708 vdd.n3057 gnd 0.010638f
C4709 vdd.n3058 gnd 0.010638f
C4710 vdd.n3059 gnd 0.017468f
C4711 vdd.n3060 gnd 0.005823f
C4712 vdd.n3061 gnd 0.010638f
C4713 vdd.n3063 gnd 0.010638f
C4714 vdd.n3065 gnd 0.010638f
C4715 vdd.n3066 gnd 0.008563f
C4716 vdd.n3067 gnd 0.008563f
C4717 vdd.n3068 gnd 0.008563f
C4718 vdd.n3069 gnd 0.010638f
C4719 vdd.n3071 gnd 0.010638f
C4720 vdd.n3073 gnd 0.010638f
C4721 vdd.n3074 gnd 0.008563f
C4722 vdd.n3075 gnd 0.008563f
C4723 vdd.n3076 gnd 0.008563f
C4724 vdd.n3077 gnd 0.010638f
C4725 vdd.n3079 gnd 0.010638f
C4726 vdd.n3081 gnd 0.010638f
C4727 vdd.n3082 gnd 0.008563f
C4728 vdd.n3083 gnd 0.008563f
C4729 vdd.n3084 gnd 0.008563f
C4730 vdd.n3085 gnd 0.010638f
C4731 vdd.n3087 gnd 0.010638f
C4732 vdd.n3089 gnd 0.010638f
C4733 vdd.n3090 gnd 0.008563f
C4734 vdd.n3091 gnd 0.008563f
C4735 vdd.n3092 gnd 0.008563f
C4736 vdd.n3093 gnd 0.010638f
C4737 vdd.n3095 gnd 0.010638f
C4738 vdd.n3097 gnd 0.010638f
C4739 vdd.n3098 gnd 0.008563f
C4740 vdd.n3099 gnd 0.008563f
C4741 vdd.n3100 gnd 0.00715f
C4742 vdd.n3101 gnd 0.010638f
C4743 vdd.n3103 gnd 0.010638f
C4744 vdd.n3105 gnd 0.010638f
C4745 vdd.n3106 gnd 0.00715f
C4746 vdd.n3107 gnd 0.008563f
C4747 vdd.n3108 gnd 0.008563f
C4748 vdd.n3109 gnd 0.010638f
C4749 vdd.n3111 gnd 0.010638f
C4750 vdd.n3113 gnd 0.010638f
C4751 vdd.n3114 gnd 0.008563f
C4752 vdd.n3115 gnd 0.008563f
C4753 vdd.n3116 gnd 0.008563f
C4754 vdd.n3117 gnd 0.010638f
C4755 vdd.n3119 gnd 0.010638f
C4756 vdd.n3121 gnd 0.010638f
C4757 vdd.n3122 gnd 0.008563f
C4758 vdd.n3123 gnd 0.008563f
C4759 vdd.n3124 gnd 0.008563f
C4760 vdd.n3125 gnd 0.010638f
C4761 vdd.n3127 gnd 0.010638f
C4762 vdd.n3128 gnd 0.010638f
C4763 vdd.n3129 gnd 0.008563f
C4764 vdd.n3130 gnd 0.008563f
C4765 vdd.n3131 gnd 0.010638f
C4766 vdd.n3132 gnd 0.010638f
C4767 vdd.n3133 gnd 0.008563f
C4768 vdd.n3134 gnd 0.008563f
C4769 vdd.n3135 gnd 0.010638f
C4770 vdd.n3136 gnd 0.010638f
C4771 vdd.n3138 gnd 0.010638f
C4772 vdd.n3139 gnd 0.008563f
C4773 vdd.n3140 gnd 0.007107f
C4774 vdd.n3141 gnd 0.024391f
C4775 vdd.n3142 gnd 0.024226f
C4776 vdd.n3143 gnd 0.007107f
C4777 vdd.n3144 gnd 0.024226f
C4778 vdd.n3145 gnd 1.43508f
C4779 vdd.n3146 gnd 0.024226f
C4780 vdd.n3147 gnd 0.007107f
C4781 vdd.n3148 gnd 0.024226f
C4782 vdd.n3149 gnd 0.010638f
C4783 vdd.n3150 gnd 0.010638f
C4784 vdd.n3151 gnd 0.008563f
C4785 vdd.n3152 gnd 0.010638f
C4786 vdd.n3153 gnd 1.02739f
C4787 vdd.n3154 gnd 0.010638f
C4788 vdd.n3155 gnd 0.008563f
C4789 vdd.n3156 gnd 0.010638f
C4790 vdd.n3157 gnd 0.010638f
C4791 vdd.n3158 gnd 0.010638f
C4792 vdd.n3159 gnd 0.008563f
C4793 vdd.n3160 gnd 0.010638f
C4794 vdd.n3161 gnd 1.06f
C4795 vdd.n3162 gnd 0.010638f
C4796 vdd.n3163 gnd 0.008563f
C4797 vdd.n3164 gnd 0.010638f
C4798 vdd.n3165 gnd 0.010638f
C4799 vdd.n3166 gnd 0.010638f
C4800 vdd.n3167 gnd 0.008563f
C4801 vdd.n3168 gnd 0.010638f
C4802 vdd.t114 gnd 0.543592f
C4803 vdd.n3169 gnd 0.875183f
C4804 vdd.n3170 gnd 0.010638f
C4805 vdd.n3171 gnd 0.008563f
C4806 vdd.n3172 gnd 0.010638f
C4807 vdd.n3173 gnd 0.010638f
C4808 vdd.n3174 gnd 0.010638f
C4809 vdd.n3175 gnd 0.008563f
C4810 vdd.n3176 gnd 0.010638f
C4811 vdd.n3177 gnd 0.690362f
C4812 vdd.n3178 gnd 0.010638f
C4813 vdd.n3179 gnd 0.008563f
C4814 vdd.n3180 gnd 0.010638f
C4815 vdd.n3181 gnd 0.010638f
C4816 vdd.n3182 gnd 0.010638f
C4817 vdd.n3183 gnd 0.008563f
C4818 vdd.n3184 gnd 0.010638f
C4819 vdd.n3185 gnd 0.864311f
C4820 vdd.n3186 gnd 0.581643f
C4821 vdd.n3187 gnd 0.010638f
C4822 vdd.n3188 gnd 0.008563f
C4823 vdd.n3189 gnd 0.010638f
C4824 vdd.n3190 gnd 0.010638f
C4825 vdd.n3191 gnd 0.010638f
C4826 vdd.n3192 gnd 0.008563f
C4827 vdd.n3193 gnd 0.010638f
C4828 vdd.n3194 gnd 0.766465f
C4829 vdd.n3195 gnd 0.010638f
C4830 vdd.n3196 gnd 0.008563f
C4831 vdd.n3197 gnd 0.010638f
C4832 vdd.n3198 gnd 0.010638f
C4833 vdd.n3199 gnd 0.010638f
C4834 vdd.n3200 gnd 0.010638f
C4835 vdd.n3201 gnd 0.010638f
C4836 vdd.n3202 gnd 0.008563f
C4837 vdd.n3203 gnd 0.008563f
C4838 vdd.n3204 gnd 0.010638f
C4839 vdd.t44 gnd 0.543592f
C4840 vdd.n3205 gnd 0.902362f
C4841 vdd.n3206 gnd 0.010638f
C4842 vdd.n3207 gnd 0.008563f
C4843 vdd.n3208 gnd 0.010638f
C4844 vdd.n3209 gnd 0.010638f
C4845 vdd.n3210 gnd 0.010638f
C4846 vdd.n3211 gnd 0.008563f
C4847 vdd.n3212 gnd 0.010638f
C4848 vdd.n3213 gnd 0.853439f
C4849 vdd.n3214 gnd 0.010638f
C4850 vdd.n3215 gnd 0.010638f
C4851 vdd.n3216 gnd 0.008563f
C4852 vdd.n3217 gnd 0.008563f
C4853 vdd.n3218 gnd 0.008563f
C4854 vdd.n3219 gnd 0.010638f
C4855 vdd.n3220 gnd 0.010638f
C4856 vdd.n3221 gnd 0.010638f
C4857 vdd.n3222 gnd 0.010638f
C4858 vdd.n3223 gnd 0.008563f
C4859 vdd.n3224 gnd 0.008563f
C4860 vdd.n3225 gnd 0.008563f
C4861 vdd.n3226 gnd 0.010638f
C4862 vdd.n3227 gnd 0.010638f
C4863 vdd.n3228 gnd 0.010638f
C4864 vdd.n3229 gnd 0.010638f
C4865 vdd.n3230 gnd 0.008563f
C4866 vdd.n3231 gnd 0.008563f
C4867 vdd.n3232 gnd 0.008563f
C4868 vdd.n3233 gnd 0.010638f
C4869 vdd.n3234 gnd 0.010638f
C4870 vdd.n3235 gnd 0.010638f
C4871 vdd.n3236 gnd 0.902362f
C4872 vdd.n3237 gnd 0.010638f
C4873 vdd.n3238 gnd 0.008563f
C4874 vdd.n3239 gnd 0.008563f
C4875 vdd.n3240 gnd 0.008563f
C4876 vdd.n3241 gnd 0.010638f
C4877 vdd.n3242 gnd 0.010638f
C4878 vdd.n3243 gnd 0.010638f
C4879 vdd.n3244 gnd 0.010638f
C4880 vdd.n3245 gnd 0.008563f
C4881 vdd.n3246 gnd 0.008563f
C4882 vdd.n3247 gnd 0.007107f
C4883 vdd.n3248 gnd 0.024226f
C4884 vdd.n3249 gnd 0.024391f
C4885 vdd.n3250 gnd 0.004067f
C4886 vdd.n3251 gnd 0.024391f
C4887 vdd.n3253 gnd 2.40268f
C4888 vdd.n3254 gnd 1.43508f
C4889 vdd.n3255 gnd 0.712105f
C4890 vdd.n3256 gnd 0.010638f
C4891 vdd.n3257 gnd 0.008563f
C4892 vdd.n3258 gnd 0.008563f
C4893 vdd.n3259 gnd 0.008563f
C4894 vdd.n3260 gnd 0.010638f
C4895 vdd.n3261 gnd 1.08718f
C4896 vdd.n3262 gnd 1.08718f
C4897 vdd.n3263 gnd 0.625131f
C4898 vdd.n3264 gnd 0.010638f
C4899 vdd.n3265 gnd 0.008563f
C4900 vdd.n3266 gnd 0.008563f
C4901 vdd.n3267 gnd 0.008563f
C4902 vdd.n3268 gnd 0.010638f
C4903 vdd.n3269 gnd 0.646874f
C4904 vdd.n3270 gnd 0.79908f
C4905 vdd.t87 gnd 0.543592f
C4906 vdd.n3271 gnd 0.831696f
C4907 vdd.n3272 gnd 0.010638f
C4908 vdd.n3273 gnd 0.008563f
C4909 vdd.n3274 gnd 0.008563f
C4910 vdd.n3275 gnd 0.008563f
C4911 vdd.n3276 gnd 0.010638f
C4912 vdd.n3277 gnd 0.902362f
C4913 vdd.t64 gnd 0.543592f
C4914 vdd.n3278 gnd 0.657746f
C4915 vdd.n3279 gnd 0.788208f
C4916 vdd.n3280 gnd 0.010638f
C4917 vdd.n3281 gnd 0.008563f
C4918 vdd.n3282 gnd 0.008563f
C4919 vdd.n3283 gnd 0.008563f
C4920 vdd.n3284 gnd 0.010638f
C4921 vdd.n3285 gnd 0.603387f
C4922 vdd.t54 gnd 0.543592f
C4923 vdd.n3286 gnd 0.902362f
C4924 vdd.t91 gnd 0.543592f
C4925 vdd.n3287 gnd 0.668618f
C4926 vdd.n3288 gnd 0.010638f
C4927 vdd.n3289 gnd 0.008563f
C4928 vdd.n3290 gnd 0.008176f
C4929 vdd.n3291 gnd 0.627487f
C4930 vdd.n3292 gnd 2.53273f
C4931 a_n6972_8799.n0 gnd 4.28745f
C4932 a_n6972_8799.n1 gnd 2.09849f
C4933 a_n6972_8799.n2 gnd 3.52374f
C4934 a_n6972_8799.n3 gnd 0.878682f
C4935 a_n6972_8799.n4 gnd 0.207867f
C4936 a_n6972_8799.n5 gnd 0.290534f
C4937 a_n6972_8799.n6 gnd 0.207867f
C4938 a_n6972_8799.n7 gnd 0.207867f
C4939 a_n6972_8799.n8 gnd 0.207867f
C4940 a_n6972_8799.n9 gnd 0.273856f
C4941 a_n6972_8799.n10 gnd 0.207867f
C4942 a_n6972_8799.n11 gnd 0.290534f
C4943 a_n6972_8799.n12 gnd 0.207867f
C4944 a_n6972_8799.n13 gnd 0.207867f
C4945 a_n6972_8799.n14 gnd 0.207867f
C4946 a_n6972_8799.n15 gnd 0.273856f
C4947 a_n6972_8799.n16 gnd 0.207867f
C4948 a_n6972_8799.n17 gnd 0.455324f
C4949 a_n6972_8799.n18 gnd 0.207867f
C4950 a_n6972_8799.n19 gnd 0.207867f
C4951 a_n6972_8799.n20 gnd 0.207867f
C4952 a_n6972_8799.n21 gnd 0.273856f
C4953 a_n6972_8799.n22 gnd 0.325823f
C4954 a_n6972_8799.n23 gnd 0.207867f
C4955 a_n6972_8799.n24 gnd 0.207867f
C4956 a_n6972_8799.n25 gnd 0.207867f
C4957 a_n6972_8799.n26 gnd 0.207867f
C4958 a_n6972_8799.n27 gnd 0.238567f
C4959 a_n6972_8799.n28 gnd 0.325823f
C4960 a_n6972_8799.n29 gnd 0.207867f
C4961 a_n6972_8799.n30 gnd 0.207867f
C4962 a_n6972_8799.n31 gnd 0.207867f
C4963 a_n6972_8799.n32 gnd 0.207867f
C4964 a_n6972_8799.n33 gnd 0.238567f
C4965 a_n6972_8799.n34 gnd 0.325823f
C4966 a_n6972_8799.n35 gnd 0.207867f
C4967 a_n6972_8799.n36 gnd 0.207867f
C4968 a_n6972_8799.n37 gnd 0.207867f
C4969 a_n6972_8799.n38 gnd 0.207867f
C4970 a_n6972_8799.n39 gnd 0.403357f
C4971 a_n6972_8799.n40 gnd 2.79204f
C4972 a_n6972_8799.n41 gnd 4.03063f
C4973 a_n6972_8799.n42 gnd 0.008622f
C4974 a_n6972_8799.n43 gnd 0.001157f
C4975 a_n6972_8799.n45 gnd 0.007742f
C4976 a_n6972_8799.n46 gnd 0.011702f
C4977 a_n6972_8799.n47 gnd 0.008048f
C4978 a_n6972_8799.n49 gnd 4.02e-19
C4979 a_n6972_8799.n50 gnd 0.008341f
C4980 a_n6972_8799.n51 gnd 0.01152f
C4981 a_n6972_8799.n52 gnd 0.007423f
C4982 a_n6972_8799.n53 gnd 0.008622f
C4983 a_n6972_8799.n54 gnd 0.001157f
C4984 a_n6972_8799.n56 gnd 0.007742f
C4985 a_n6972_8799.n57 gnd 0.011702f
C4986 a_n6972_8799.n58 gnd 0.008048f
C4987 a_n6972_8799.n60 gnd 4.02e-19
C4988 a_n6972_8799.n61 gnd 0.008341f
C4989 a_n6972_8799.n62 gnd 0.01152f
C4990 a_n6972_8799.n63 gnd 0.007423f
C4991 a_n6972_8799.n64 gnd 0.008622f
C4992 a_n6972_8799.n65 gnd 0.001157f
C4993 a_n6972_8799.n67 gnd 0.007742f
C4994 a_n6972_8799.n68 gnd 0.011702f
C4995 a_n6972_8799.n69 gnd 0.008048f
C4996 a_n6972_8799.n71 gnd 4.02e-19
C4997 a_n6972_8799.n72 gnd 0.008341f
C4998 a_n6972_8799.n73 gnd 0.01152f
C4999 a_n6972_8799.n74 gnd 0.007423f
C5000 a_n6972_8799.n75 gnd 0.001157f
C5001 a_n6972_8799.n77 gnd 0.007742f
C5002 a_n6972_8799.n78 gnd 0.011702f
C5003 a_n6972_8799.n79 gnd 0.008048f
C5004 a_n6972_8799.n81 gnd 4.02e-19
C5005 a_n6972_8799.n82 gnd 0.008341f
C5006 a_n6972_8799.n83 gnd 0.01152f
C5007 a_n6972_8799.n84 gnd 0.007423f
C5008 a_n6972_8799.n85 gnd 0.250252f
C5009 a_n6972_8799.n86 gnd 0.001157f
C5010 a_n6972_8799.n88 gnd 0.007742f
C5011 a_n6972_8799.n89 gnd 0.011702f
C5012 a_n6972_8799.n90 gnd 0.008048f
C5013 a_n6972_8799.n92 gnd 4.02e-19
C5014 a_n6972_8799.n93 gnd 0.008341f
C5015 a_n6972_8799.n94 gnd 0.01152f
C5016 a_n6972_8799.n95 gnd 0.007423f
C5017 a_n6972_8799.n96 gnd 0.250252f
C5018 a_n6972_8799.n97 gnd 0.001157f
C5019 a_n6972_8799.n99 gnd 0.007742f
C5020 a_n6972_8799.n100 gnd 0.011702f
C5021 a_n6972_8799.n101 gnd 0.008048f
C5022 a_n6972_8799.n103 gnd 4.02e-19
C5023 a_n6972_8799.n104 gnd 0.008341f
C5024 a_n6972_8799.n105 gnd 0.01152f
C5025 a_n6972_8799.n106 gnd 0.007423f
C5026 a_n6972_8799.n107 gnd 0.250252f
C5027 a_n6972_8799.t11 gnd 0.144179f
C5028 a_n6972_8799.t33 gnd 0.144179f
C5029 a_n6972_8799.t6 gnd 0.144179f
C5030 a_n6972_8799.n108 gnd 1.13716f
C5031 a_n6972_8799.t17 gnd 0.144179f
C5032 a_n6972_8799.t12 gnd 0.144179f
C5033 a_n6972_8799.n109 gnd 1.13529f
C5034 a_n6972_8799.t21 gnd 0.144179f
C5035 a_n6972_8799.t29 gnd 0.144179f
C5036 a_n6972_8799.n110 gnd 1.13529f
C5037 a_n6972_8799.t20 gnd 0.112139f
C5038 a_n6972_8799.t22 gnd 0.112139f
C5039 a_n6972_8799.n111 gnd 0.993823f
C5040 a_n6972_8799.t19 gnd 0.112139f
C5041 a_n6972_8799.t2 gnd 0.112139f
C5042 a_n6972_8799.n112 gnd 0.990901f
C5043 a_n6972_8799.t18 gnd 0.112139f
C5044 a_n6972_8799.t23 gnd 0.112139f
C5045 a_n6972_8799.n113 gnd 0.990901f
C5046 a_n6972_8799.t27 gnd 0.112139f
C5047 a_n6972_8799.t32 gnd 0.112139f
C5048 a_n6972_8799.n114 gnd 0.993823f
C5049 a_n6972_8799.t0 gnd 0.112139f
C5050 a_n6972_8799.t1 gnd 0.112139f
C5051 a_n6972_8799.n115 gnd 0.990901f
C5052 a_n6972_8799.t14 gnd 0.112139f
C5053 a_n6972_8799.t26 gnd 0.112139f
C5054 a_n6972_8799.n116 gnd 0.990901f
C5055 a_n6972_8799.t7 gnd 0.112139f
C5056 a_n6972_8799.t8 gnd 0.112139f
C5057 a_n6972_8799.n117 gnd 0.993823f
C5058 a_n6972_8799.t9 gnd 0.112139f
C5059 a_n6972_8799.t16 gnd 0.112139f
C5060 a_n6972_8799.n118 gnd 0.990901f
C5061 a_n6972_8799.t25 gnd 0.112139f
C5062 a_n6972_8799.t24 gnd 0.112139f
C5063 a_n6972_8799.n119 gnd 0.990901f
C5064 a_n6972_8799.t10 gnd 0.112139f
C5065 a_n6972_8799.t13 gnd 0.112139f
C5066 a_n6972_8799.n120 gnd 0.990901f
C5067 a_n6972_8799.t15 gnd 0.112139f
C5068 a_n6972_8799.t28 gnd 0.112139f
C5069 a_n6972_8799.n121 gnd 0.990901f
C5070 a_n6972_8799.t30 gnd 0.112139f
C5071 a_n6972_8799.t31 gnd 0.112139f
C5072 a_n6972_8799.n122 gnd 0.990901f
C5073 a_n6972_8799.t113 gnd 0.597833f
C5074 a_n6972_8799.n123 gnd 0.267276f
C5075 a_n6972_8799.t47 gnd 0.597833f
C5076 a_n6972_8799.t65 gnd 0.597833f
C5077 a_n6972_8799.n124 gnd 0.270588f
C5078 a_n6972_8799.t82 gnd 0.597833f
C5079 a_n6972_8799.t99 gnd 0.597833f
C5080 a_n6972_8799.t100 gnd 0.597833f
C5081 a_n6972_8799.n125 gnd 0.272673f
C5082 a_n6972_8799.t67 gnd 0.597833f
C5083 a_n6972_8799.t76 gnd 0.597833f
C5084 a_n6972_8799.n126 gnd 0.266203f
C5085 a_n6972_8799.t114 gnd 0.609148f
C5086 a_n6972_8799.n127 gnd 0.250638f
C5087 a_n6972_8799.n128 gnd 0.011792f
C5088 a_n6972_8799.t77 gnd 0.597833f
C5089 a_n6972_8799.n129 gnd 0.267004f
C5090 a_n6972_8799.n130 gnd 0.270573f
C5091 a_n6972_8799.t68 gnd 0.597833f
C5092 a_n6972_8799.n131 gnd 0.267094f
C5093 a_n6972_8799.n132 gnd 0.261717f
C5094 a_n6972_8799.t36 gnd 0.597833f
C5095 a_n6972_8799.n133 gnd 0.266844f
C5096 a_n6972_8799.n134 gnd 0.273108f
C5097 a_n6972_8799.t116 gnd 0.597833f
C5098 a_n6972_8799.n135 gnd 0.270455f
C5099 a_n6972_8799.n136 gnd 0.266523f
C5100 a_n6972_8799.t63 gnd 0.597833f
C5101 a_n6972_8799.n137 gnd 0.262038f
C5102 a_n6972_8799.t44 gnd 0.597833f
C5103 a_n6972_8799.n138 gnd 0.270572f
C5104 a_n6972_8799.t45 gnd 0.609138f
C5105 a_n6972_8799.t123 gnd 0.597833f
C5106 a_n6972_8799.n139 gnd 0.267276f
C5107 a_n6972_8799.t61 gnd 0.597833f
C5108 a_n6972_8799.t73 gnd 0.597833f
C5109 a_n6972_8799.n140 gnd 0.270588f
C5110 a_n6972_8799.t93 gnd 0.597833f
C5111 a_n6972_8799.t108 gnd 0.597833f
C5112 a_n6972_8799.t112 gnd 0.597833f
C5113 a_n6972_8799.n141 gnd 0.272673f
C5114 a_n6972_8799.t74 gnd 0.597833f
C5115 a_n6972_8799.t83 gnd 0.597833f
C5116 a_n6972_8799.n142 gnd 0.266203f
C5117 a_n6972_8799.t125 gnd 0.609148f
C5118 a_n6972_8799.n143 gnd 0.250638f
C5119 a_n6972_8799.n144 gnd 0.011792f
C5120 a_n6972_8799.t84 gnd 0.597833f
C5121 a_n6972_8799.n145 gnd 0.267004f
C5122 a_n6972_8799.n146 gnd 0.270573f
C5123 a_n6972_8799.t75 gnd 0.597833f
C5124 a_n6972_8799.n147 gnd 0.267094f
C5125 a_n6972_8799.n148 gnd 0.261717f
C5126 a_n6972_8799.t46 gnd 0.597833f
C5127 a_n6972_8799.n149 gnd 0.266844f
C5128 a_n6972_8799.n150 gnd 0.273108f
C5129 a_n6972_8799.t128 gnd 0.597833f
C5130 a_n6972_8799.n151 gnd 0.270455f
C5131 a_n6972_8799.n152 gnd 0.266523f
C5132 a_n6972_8799.t72 gnd 0.597833f
C5133 a_n6972_8799.n153 gnd 0.262038f
C5134 a_n6972_8799.t55 gnd 0.597833f
C5135 a_n6972_8799.n154 gnd 0.270572f
C5136 a_n6972_8799.t57 gnd 0.609138f
C5137 a_n6972_8799.n155 gnd 0.900403f
C5138 a_n6972_8799.t89 gnd 0.597833f
C5139 a_n6972_8799.n156 gnd 0.267276f
C5140 a_n6972_8799.t109 gnd 0.597833f
C5141 a_n6972_8799.t42 gnd 0.597833f
C5142 a_n6972_8799.n157 gnd 0.270588f
C5143 a_n6972_8799.t95 gnd 0.597833f
C5144 a_n6972_8799.t124 gnd 0.597833f
C5145 a_n6972_8799.t87 gnd 0.597833f
C5146 a_n6972_8799.n158 gnd 0.272673f
C5147 a_n6972_8799.t120 gnd 0.597833f
C5148 a_n6972_8799.t53 gnd 0.597833f
C5149 a_n6972_8799.n159 gnd 0.266203f
C5150 a_n6972_8799.t117 gnd 0.609148f
C5151 a_n6972_8799.n160 gnd 0.250638f
C5152 a_n6972_8799.n161 gnd 0.011792f
C5153 a_n6972_8799.t37 gnd 0.597833f
C5154 a_n6972_8799.n162 gnd 0.267004f
C5155 a_n6972_8799.n163 gnd 0.270573f
C5156 a_n6972_8799.t101 gnd 0.597833f
C5157 a_n6972_8799.n164 gnd 0.267094f
C5158 a_n6972_8799.n165 gnd 0.261717f
C5159 a_n6972_8799.t81 gnd 0.597833f
C5160 a_n6972_8799.n166 gnd 0.266844f
C5161 a_n6972_8799.n167 gnd 0.273108f
C5162 a_n6972_8799.t59 gnd 0.597833f
C5163 a_n6972_8799.n168 gnd 0.270455f
C5164 a_n6972_8799.n169 gnd 0.266523f
C5165 a_n6972_8799.t66 gnd 0.597833f
C5166 a_n6972_8799.n170 gnd 0.262038f
C5167 a_n6972_8799.t49 gnd 0.597833f
C5168 a_n6972_8799.n171 gnd 0.270572f
C5169 a_n6972_8799.t129 gnd 0.609138f
C5170 a_n6972_8799.n172 gnd 1.53998f
C5171 a_n6972_8799.t79 gnd 0.597833f
C5172 a_n6972_8799.t78 gnd 0.597833f
C5173 a_n6972_8799.t56 gnd 0.597833f
C5174 a_n6972_8799.n173 gnd 0.270174f
C5175 a_n6972_8799.t115 gnd 0.597833f
C5176 a_n6972_8799.t80 gnd 0.597833f
C5177 a_n6972_8799.t62 gnd 0.597833f
C5178 a_n6972_8799.n174 gnd 0.267094f
C5179 a_n6972_8799.t119 gnd 0.597833f
C5180 a_n6972_8799.t94 gnd 0.597833f
C5181 a_n6972_8799.t92 gnd 0.597833f
C5182 a_n6972_8799.n175 gnd 0.270588f
C5183 a_n6972_8799.t39 gnd 0.597833f
C5184 a_n6972_8799.t98 gnd 0.597833f
C5185 a_n6972_8799.t97 gnd 0.597833f
C5186 a_n6972_8799.n176 gnd 0.266523f
C5187 a_n6972_8799.t41 gnd 0.597833f
C5188 a_n6972_8799.t40 gnd 0.597833f
C5189 a_n6972_8799.t111 gnd 0.597833f
C5190 a_n6972_8799.n177 gnd 0.270572f
C5191 a_n6972_8799.t58 gnd 0.609148f
C5192 a_n6972_8799.n178 gnd 0.250638f
C5193 a_n6972_8799.n179 gnd 0.267276f
C5194 a_n6972_8799.n180 gnd 0.262038f
C5195 a_n6972_8799.n181 gnd 0.270455f
C5196 a_n6972_8799.n182 gnd 0.273108f
C5197 a_n6972_8799.n183 gnd 0.266844f
C5198 a_n6972_8799.n184 gnd 0.261717f
C5199 a_n6972_8799.n185 gnd 0.270573f
C5200 a_n6972_8799.n186 gnd 0.272673f
C5201 a_n6972_8799.n187 gnd 0.266203f
C5202 a_n6972_8799.n188 gnd 0.261557f
C5203 a_n6972_8799.t86 gnd 0.597833f
C5204 a_n6972_8799.t85 gnd 0.597833f
C5205 a_n6972_8799.t69 gnd 0.597833f
C5206 a_n6972_8799.n189 gnd 0.270174f
C5207 a_n6972_8799.t127 gnd 0.597833f
C5208 a_n6972_8799.t91 gnd 0.597833f
C5209 a_n6972_8799.t71 gnd 0.597833f
C5210 a_n6972_8799.n190 gnd 0.267094f
C5211 a_n6972_8799.t131 gnd 0.597833f
C5212 a_n6972_8799.t104 gnd 0.597833f
C5213 a_n6972_8799.t103 gnd 0.597833f
C5214 a_n6972_8799.n191 gnd 0.270588f
C5215 a_n6972_8799.t48 gnd 0.597833f
C5216 a_n6972_8799.t107 gnd 0.597833f
C5217 a_n6972_8799.t106 gnd 0.597833f
C5218 a_n6972_8799.n192 gnd 0.266523f
C5219 a_n6972_8799.t52 gnd 0.597833f
C5220 a_n6972_8799.t51 gnd 0.597833f
C5221 a_n6972_8799.t122 gnd 0.597833f
C5222 a_n6972_8799.n193 gnd 0.270572f
C5223 a_n6972_8799.t70 gnd 0.609148f
C5224 a_n6972_8799.n194 gnd 0.250638f
C5225 a_n6972_8799.n195 gnd 0.267276f
C5226 a_n6972_8799.n196 gnd 0.262038f
C5227 a_n6972_8799.n197 gnd 0.270455f
C5228 a_n6972_8799.n198 gnd 0.273108f
C5229 a_n6972_8799.n199 gnd 0.266844f
C5230 a_n6972_8799.n200 gnd 0.261717f
C5231 a_n6972_8799.n201 gnd 0.270573f
C5232 a_n6972_8799.n202 gnd 0.272673f
C5233 a_n6972_8799.n203 gnd 0.266203f
C5234 a_n6972_8799.n204 gnd 0.261557f
C5235 a_n6972_8799.n205 gnd 0.900403f
C5236 a_n6972_8799.t130 gnd 0.597833f
C5237 a_n6972_8799.t50 gnd 0.597833f
C5238 a_n6972_8799.t90 gnd 0.597833f
C5239 a_n6972_8799.n206 gnd 0.270174f
C5240 a_n6972_8799.t38 gnd 0.597833f
C5241 a_n6972_8799.t110 gnd 0.597833f
C5242 a_n6972_8799.t60 gnd 0.597833f
C5243 a_n6972_8799.n207 gnd 0.267094f
C5244 a_n6972_8799.t96 gnd 0.597833f
C5245 a_n6972_8799.t43 gnd 0.597833f
C5246 a_n6972_8799.t64 gnd 0.597833f
C5247 a_n6972_8799.n208 gnd 0.270588f
C5248 a_n6972_8799.t126 gnd 0.597833f
C5249 a_n6972_8799.t102 gnd 0.597833f
C5250 a_n6972_8799.t121 gnd 0.597833f
C5251 a_n6972_8799.n209 gnd 0.266523f
C5252 a_n6972_8799.t88 gnd 0.597833f
C5253 a_n6972_8799.t105 gnd 0.597833f
C5254 a_n6972_8799.t54 gnd 0.597833f
C5255 a_n6972_8799.n210 gnd 0.270572f
C5256 a_n6972_8799.t118 gnd 0.609148f
C5257 a_n6972_8799.n211 gnd 0.250638f
C5258 a_n6972_8799.n212 gnd 0.267276f
C5259 a_n6972_8799.n213 gnd 0.262038f
C5260 a_n6972_8799.n214 gnd 0.270455f
C5261 a_n6972_8799.n215 gnd 0.273108f
C5262 a_n6972_8799.n216 gnd 0.266844f
C5263 a_n6972_8799.n217 gnd 0.261717f
C5264 a_n6972_8799.n218 gnd 0.270573f
C5265 a_n6972_8799.n219 gnd 0.272673f
C5266 a_n6972_8799.n220 gnd 0.266203f
C5267 a_n6972_8799.n221 gnd 0.261557f
C5268 a_n6972_8799.n222 gnd 1.08681f
C5269 a_n6972_8799.n223 gnd 12.2105f
C5270 a_n6972_8799.n224 gnd 4.37527f
C5271 a_n6972_8799.n225 gnd 5.67666f
C5272 a_n6972_8799.t34 gnd 0.144179f
C5273 a_n6972_8799.t4 gnd 0.144179f
C5274 a_n6972_8799.n226 gnd 1.13529f
C5275 a_n6972_8799.t35 gnd 0.144179f
C5276 a_n6972_8799.t5 gnd 0.144179f
C5277 a_n6972_8799.n227 gnd 1.13529f
C5278 a_n6972_8799.n228 gnd 1.13717f
C5279 a_n6972_8799.t3 gnd 0.144179f
C5280 commonsourceibias.n0 gnd 0.012626f
C5281 commonsourceibias.t78 gnd 0.191194f
C5282 commonsourceibias.t146 gnd 0.176786f
C5283 commonsourceibias.n1 gnd 0.007691f
C5284 commonsourceibias.n2 gnd 0.009462f
C5285 commonsourceibias.t96 gnd 0.176786f
C5286 commonsourceibias.n3 gnd 0.009599f
C5287 commonsourceibias.n4 gnd 0.009462f
C5288 commonsourceibias.t157 gnd 0.176786f
C5289 commonsourceibias.n5 gnd 0.070538f
C5290 commonsourceibias.t112 gnd 0.176786f
C5291 commonsourceibias.n6 gnd 0.007654f
C5292 commonsourceibias.n7 gnd 0.009462f
C5293 commonsourceibias.t75 gnd 0.176786f
C5294 commonsourceibias.n8 gnd 0.009135f
C5295 commonsourceibias.n9 gnd 0.009462f
C5296 commonsourceibias.t124 gnd 0.176786f
C5297 commonsourceibias.n10 gnd 0.070538f
C5298 commonsourceibias.t113 gnd 0.176786f
C5299 commonsourceibias.n11 gnd 0.007642f
C5300 commonsourceibias.n12 gnd 0.012626f
C5301 commonsourceibias.t20 gnd 0.191194f
C5302 commonsourceibias.t50 gnd 0.176786f
C5303 commonsourceibias.n13 gnd 0.007691f
C5304 commonsourceibias.n14 gnd 0.009462f
C5305 commonsourceibias.t4 gnd 0.176786f
C5306 commonsourceibias.n15 gnd 0.009599f
C5307 commonsourceibias.n16 gnd 0.009462f
C5308 commonsourceibias.t40 gnd 0.176786f
C5309 commonsourceibias.n17 gnd 0.070538f
C5310 commonsourceibias.t34 gnd 0.176786f
C5311 commonsourceibias.n18 gnd 0.007654f
C5312 commonsourceibias.n19 gnd 0.009462f
C5313 commonsourceibias.t22 gnd 0.176786f
C5314 commonsourceibias.n20 gnd 0.009135f
C5315 commonsourceibias.n21 gnd 0.009462f
C5316 commonsourceibias.t24 gnd 0.176786f
C5317 commonsourceibias.n22 gnd 0.070538f
C5318 commonsourceibias.t32 gnd 0.176786f
C5319 commonsourceibias.n23 gnd 0.007642f
C5320 commonsourceibias.n24 gnd 0.009462f
C5321 commonsourceibias.t42 gnd 0.176786f
C5322 commonsourceibias.t0 gnd 0.176786f
C5323 commonsourceibias.n25 gnd 0.070538f
C5324 commonsourceibias.n26 gnd 0.009462f
C5325 commonsourceibias.t8 gnd 0.176786f
C5326 commonsourceibias.n27 gnd 0.070538f
C5327 commonsourceibias.n28 gnd 0.009462f
C5328 commonsourceibias.t26 gnd 0.176786f
C5329 commonsourceibias.n29 gnd 0.070538f
C5330 commonsourceibias.n30 gnd 0.009462f
C5331 commonsourceibias.t36 gnd 0.176786f
C5332 commonsourceibias.n31 gnd 0.010756f
C5333 commonsourceibias.n32 gnd 0.009462f
C5334 commonsourceibias.t62 gnd 0.176786f
C5335 commonsourceibias.n33 gnd 0.012719f
C5336 commonsourceibias.t52 gnd 0.196936f
C5337 commonsourceibias.t48 gnd 0.176786f
C5338 commonsourceibias.n34 gnd 0.078597f
C5339 commonsourceibias.n35 gnd 0.084205f
C5340 commonsourceibias.n36 gnd 0.040277f
C5341 commonsourceibias.n37 gnd 0.009462f
C5342 commonsourceibias.n38 gnd 0.007691f
C5343 commonsourceibias.n39 gnd 0.013039f
C5344 commonsourceibias.n40 gnd 0.070538f
C5345 commonsourceibias.n41 gnd 0.013095f
C5346 commonsourceibias.n42 gnd 0.009462f
C5347 commonsourceibias.n43 gnd 0.009462f
C5348 commonsourceibias.n44 gnd 0.009462f
C5349 commonsourceibias.n45 gnd 0.009599f
C5350 commonsourceibias.n46 gnd 0.070538f
C5351 commonsourceibias.n47 gnd 0.011663f
C5352 commonsourceibias.n48 gnd 0.012902f
C5353 commonsourceibias.n49 gnd 0.009462f
C5354 commonsourceibias.n50 gnd 0.009462f
C5355 commonsourceibias.n51 gnd 0.012818f
C5356 commonsourceibias.n52 gnd 0.007654f
C5357 commonsourceibias.n53 gnd 0.012977f
C5358 commonsourceibias.n54 gnd 0.009462f
C5359 commonsourceibias.n55 gnd 0.009462f
C5360 commonsourceibias.n56 gnd 0.013056f
C5361 commonsourceibias.n57 gnd 0.011258f
C5362 commonsourceibias.n58 gnd 0.009135f
C5363 commonsourceibias.n59 gnd 0.009462f
C5364 commonsourceibias.n60 gnd 0.009462f
C5365 commonsourceibias.n61 gnd 0.011574f
C5366 commonsourceibias.n62 gnd 0.012991f
C5367 commonsourceibias.n63 gnd 0.070538f
C5368 commonsourceibias.n64 gnd 0.012903f
C5369 commonsourceibias.n65 gnd 0.009462f
C5370 commonsourceibias.n66 gnd 0.009462f
C5371 commonsourceibias.n67 gnd 0.009462f
C5372 commonsourceibias.n68 gnd 0.012903f
C5373 commonsourceibias.n69 gnd 0.070538f
C5374 commonsourceibias.n70 gnd 0.012991f
C5375 commonsourceibias.n71 gnd 0.011574f
C5376 commonsourceibias.n72 gnd 0.009462f
C5377 commonsourceibias.n73 gnd 0.009462f
C5378 commonsourceibias.n74 gnd 0.009462f
C5379 commonsourceibias.n75 gnd 0.011258f
C5380 commonsourceibias.n76 gnd 0.013056f
C5381 commonsourceibias.n77 gnd 0.070538f
C5382 commonsourceibias.n78 gnd 0.012977f
C5383 commonsourceibias.n79 gnd 0.009462f
C5384 commonsourceibias.n80 gnd 0.009462f
C5385 commonsourceibias.n81 gnd 0.009462f
C5386 commonsourceibias.n82 gnd 0.012818f
C5387 commonsourceibias.n83 gnd 0.070538f
C5388 commonsourceibias.n84 gnd 0.012902f
C5389 commonsourceibias.n85 gnd 0.011663f
C5390 commonsourceibias.n86 gnd 0.009462f
C5391 commonsourceibias.n87 gnd 0.009462f
C5392 commonsourceibias.n88 gnd 0.009462f
C5393 commonsourceibias.n89 gnd 0.010756f
C5394 commonsourceibias.n90 gnd 0.013095f
C5395 commonsourceibias.n91 gnd 0.070538f
C5396 commonsourceibias.n92 gnd 0.013039f
C5397 commonsourceibias.n93 gnd 0.009462f
C5398 commonsourceibias.n94 gnd 0.009462f
C5399 commonsourceibias.n95 gnd 0.009462f
C5400 commonsourceibias.n96 gnd 0.012719f
C5401 commonsourceibias.n97 gnd 0.070538f
C5402 commonsourceibias.n98 gnd 0.01275f
C5403 commonsourceibias.n99 gnd 0.085058f
C5404 commonsourceibias.n100 gnd 0.095108f
C5405 commonsourceibias.t21 gnd 0.020419f
C5406 commonsourceibias.t51 gnd 0.020419f
C5407 commonsourceibias.n101 gnd 0.180428f
C5408 commonsourceibias.n102 gnd 0.15629f
C5409 commonsourceibias.t5 gnd 0.020419f
C5410 commonsourceibias.t41 gnd 0.020419f
C5411 commonsourceibias.n103 gnd 0.180428f
C5412 commonsourceibias.n104 gnd 0.082878f
C5413 commonsourceibias.t35 gnd 0.020419f
C5414 commonsourceibias.t23 gnd 0.020419f
C5415 commonsourceibias.n105 gnd 0.180428f
C5416 commonsourceibias.n106 gnd 0.082878f
C5417 commonsourceibias.t25 gnd 0.020419f
C5418 commonsourceibias.t33 gnd 0.020419f
C5419 commonsourceibias.n107 gnd 0.180428f
C5420 commonsourceibias.n108 gnd 0.06924f
C5421 commonsourceibias.t49 gnd 0.020419f
C5422 commonsourceibias.t53 gnd 0.020419f
C5423 commonsourceibias.n109 gnd 0.181032f
C5424 commonsourceibias.t37 gnd 0.020419f
C5425 commonsourceibias.t63 gnd 0.020419f
C5426 commonsourceibias.n110 gnd 0.180428f
C5427 commonsourceibias.n111 gnd 0.168125f
C5428 commonsourceibias.t9 gnd 0.020419f
C5429 commonsourceibias.t27 gnd 0.020419f
C5430 commonsourceibias.n112 gnd 0.180428f
C5431 commonsourceibias.n113 gnd 0.082878f
C5432 commonsourceibias.t43 gnd 0.020419f
C5433 commonsourceibias.t1 gnd 0.020419f
C5434 commonsourceibias.n114 gnd 0.180428f
C5435 commonsourceibias.n115 gnd 0.06924f
C5436 commonsourceibias.n116 gnd 0.083843f
C5437 commonsourceibias.n117 gnd 0.009462f
C5438 commonsourceibias.t154 gnd 0.176786f
C5439 commonsourceibias.t106 gnd 0.176786f
C5440 commonsourceibias.n118 gnd 0.070538f
C5441 commonsourceibias.n119 gnd 0.009462f
C5442 commonsourceibias.t92 gnd 0.176786f
C5443 commonsourceibias.n120 gnd 0.070538f
C5444 commonsourceibias.n121 gnd 0.009462f
C5445 commonsourceibias.t123 gnd 0.176786f
C5446 commonsourceibias.n122 gnd 0.070538f
C5447 commonsourceibias.n123 gnd 0.009462f
C5448 commonsourceibias.t110 gnd 0.176786f
C5449 commonsourceibias.n124 gnd 0.010756f
C5450 commonsourceibias.n125 gnd 0.009462f
C5451 commonsourceibias.t82 gnd 0.176786f
C5452 commonsourceibias.n126 gnd 0.012719f
C5453 commonsourceibias.t132 gnd 0.196936f
C5454 commonsourceibias.t147 gnd 0.176786f
C5455 commonsourceibias.n127 gnd 0.078597f
C5456 commonsourceibias.n128 gnd 0.084205f
C5457 commonsourceibias.n129 gnd 0.040277f
C5458 commonsourceibias.n130 gnd 0.009462f
C5459 commonsourceibias.n131 gnd 0.007691f
C5460 commonsourceibias.n132 gnd 0.013039f
C5461 commonsourceibias.n133 gnd 0.070538f
C5462 commonsourceibias.n134 gnd 0.013095f
C5463 commonsourceibias.n135 gnd 0.009462f
C5464 commonsourceibias.n136 gnd 0.009462f
C5465 commonsourceibias.n137 gnd 0.009462f
C5466 commonsourceibias.n138 gnd 0.009599f
C5467 commonsourceibias.n139 gnd 0.070538f
C5468 commonsourceibias.n140 gnd 0.011663f
C5469 commonsourceibias.n141 gnd 0.012902f
C5470 commonsourceibias.n142 gnd 0.009462f
C5471 commonsourceibias.n143 gnd 0.009462f
C5472 commonsourceibias.n144 gnd 0.012818f
C5473 commonsourceibias.n145 gnd 0.007654f
C5474 commonsourceibias.n146 gnd 0.012977f
C5475 commonsourceibias.n147 gnd 0.009462f
C5476 commonsourceibias.n148 gnd 0.009462f
C5477 commonsourceibias.n149 gnd 0.013056f
C5478 commonsourceibias.n150 gnd 0.011258f
C5479 commonsourceibias.n151 gnd 0.009135f
C5480 commonsourceibias.n152 gnd 0.009462f
C5481 commonsourceibias.n153 gnd 0.009462f
C5482 commonsourceibias.n154 gnd 0.011574f
C5483 commonsourceibias.n155 gnd 0.012991f
C5484 commonsourceibias.n156 gnd 0.070538f
C5485 commonsourceibias.n157 gnd 0.012903f
C5486 commonsourceibias.n158 gnd 0.009417f
C5487 commonsourceibias.n159 gnd 0.068402f
C5488 commonsourceibias.n160 gnd 0.009417f
C5489 commonsourceibias.n161 gnd 0.012903f
C5490 commonsourceibias.n162 gnd 0.070538f
C5491 commonsourceibias.n163 gnd 0.012991f
C5492 commonsourceibias.n164 gnd 0.011574f
C5493 commonsourceibias.n165 gnd 0.009462f
C5494 commonsourceibias.n166 gnd 0.009462f
C5495 commonsourceibias.n167 gnd 0.009462f
C5496 commonsourceibias.n168 gnd 0.011258f
C5497 commonsourceibias.n169 gnd 0.013056f
C5498 commonsourceibias.n170 gnd 0.070538f
C5499 commonsourceibias.n171 gnd 0.012977f
C5500 commonsourceibias.n172 gnd 0.009462f
C5501 commonsourceibias.n173 gnd 0.009462f
C5502 commonsourceibias.n174 gnd 0.009462f
C5503 commonsourceibias.n175 gnd 0.012818f
C5504 commonsourceibias.n176 gnd 0.070538f
C5505 commonsourceibias.n177 gnd 0.012902f
C5506 commonsourceibias.n178 gnd 0.011663f
C5507 commonsourceibias.n179 gnd 0.009462f
C5508 commonsourceibias.n180 gnd 0.009462f
C5509 commonsourceibias.n181 gnd 0.009462f
C5510 commonsourceibias.n182 gnd 0.010756f
C5511 commonsourceibias.n183 gnd 0.013095f
C5512 commonsourceibias.n184 gnd 0.070538f
C5513 commonsourceibias.n185 gnd 0.013039f
C5514 commonsourceibias.n186 gnd 0.009462f
C5515 commonsourceibias.n187 gnd 0.009462f
C5516 commonsourceibias.n188 gnd 0.009462f
C5517 commonsourceibias.n189 gnd 0.012719f
C5518 commonsourceibias.n190 gnd 0.070538f
C5519 commonsourceibias.n191 gnd 0.01275f
C5520 commonsourceibias.n192 gnd 0.085058f
C5521 commonsourceibias.n193 gnd 0.056191f
C5522 commonsourceibias.n194 gnd 0.012626f
C5523 commonsourceibias.t115 gnd 0.191194f
C5524 commonsourceibias.t138 gnd 0.176786f
C5525 commonsourceibias.n195 gnd 0.007691f
C5526 commonsourceibias.n196 gnd 0.009462f
C5527 commonsourceibias.t128 gnd 0.176786f
C5528 commonsourceibias.n197 gnd 0.009599f
C5529 commonsourceibias.n198 gnd 0.009462f
C5530 commonsourceibias.t116 gnd 0.176786f
C5531 commonsourceibias.n199 gnd 0.070538f
C5532 commonsourceibias.t139 gnd 0.176786f
C5533 commonsourceibias.n200 gnd 0.007654f
C5534 commonsourceibias.n201 gnd 0.009462f
C5535 commonsourceibias.t126 gnd 0.176786f
C5536 commonsourceibias.n202 gnd 0.009135f
C5537 commonsourceibias.n203 gnd 0.009462f
C5538 commonsourceibias.t114 gnd 0.176786f
C5539 commonsourceibias.n204 gnd 0.070538f
C5540 commonsourceibias.t140 gnd 0.176786f
C5541 commonsourceibias.n205 gnd 0.007642f
C5542 commonsourceibias.n206 gnd 0.009462f
C5543 commonsourceibias.t127 gnd 0.176786f
C5544 commonsourceibias.t149 gnd 0.176786f
C5545 commonsourceibias.n207 gnd 0.070538f
C5546 commonsourceibias.n208 gnd 0.009462f
C5547 commonsourceibias.t141 gnd 0.176786f
C5548 commonsourceibias.n209 gnd 0.070538f
C5549 commonsourceibias.n210 gnd 0.009462f
C5550 commonsourceibias.t125 gnd 0.176786f
C5551 commonsourceibias.n211 gnd 0.070538f
C5552 commonsourceibias.n212 gnd 0.009462f
C5553 commonsourceibias.t152 gnd 0.176786f
C5554 commonsourceibias.n213 gnd 0.010756f
C5555 commonsourceibias.n214 gnd 0.009462f
C5556 commonsourceibias.t69 gnd 0.176786f
C5557 commonsourceibias.n215 gnd 0.012719f
C5558 commonsourceibias.t64 gnd 0.196936f
C5559 commonsourceibias.t135 gnd 0.176786f
C5560 commonsourceibias.n216 gnd 0.078597f
C5561 commonsourceibias.n217 gnd 0.084205f
C5562 commonsourceibias.n218 gnd 0.040277f
C5563 commonsourceibias.n219 gnd 0.009462f
C5564 commonsourceibias.n220 gnd 0.007691f
C5565 commonsourceibias.n221 gnd 0.013039f
C5566 commonsourceibias.n222 gnd 0.070538f
C5567 commonsourceibias.n223 gnd 0.013095f
C5568 commonsourceibias.n224 gnd 0.009462f
C5569 commonsourceibias.n225 gnd 0.009462f
C5570 commonsourceibias.n226 gnd 0.009462f
C5571 commonsourceibias.n227 gnd 0.009599f
C5572 commonsourceibias.n228 gnd 0.070538f
C5573 commonsourceibias.n229 gnd 0.011663f
C5574 commonsourceibias.n230 gnd 0.012902f
C5575 commonsourceibias.n231 gnd 0.009462f
C5576 commonsourceibias.n232 gnd 0.009462f
C5577 commonsourceibias.n233 gnd 0.012818f
C5578 commonsourceibias.n234 gnd 0.007654f
C5579 commonsourceibias.n235 gnd 0.012977f
C5580 commonsourceibias.n236 gnd 0.009462f
C5581 commonsourceibias.n237 gnd 0.009462f
C5582 commonsourceibias.n238 gnd 0.013056f
C5583 commonsourceibias.n239 gnd 0.011258f
C5584 commonsourceibias.n240 gnd 0.009135f
C5585 commonsourceibias.n241 gnd 0.009462f
C5586 commonsourceibias.n242 gnd 0.009462f
C5587 commonsourceibias.n243 gnd 0.011574f
C5588 commonsourceibias.n244 gnd 0.012991f
C5589 commonsourceibias.n245 gnd 0.070538f
C5590 commonsourceibias.n246 gnd 0.012903f
C5591 commonsourceibias.n247 gnd 0.009462f
C5592 commonsourceibias.n248 gnd 0.009462f
C5593 commonsourceibias.n249 gnd 0.009462f
C5594 commonsourceibias.n250 gnd 0.012903f
C5595 commonsourceibias.n251 gnd 0.070538f
C5596 commonsourceibias.n252 gnd 0.012991f
C5597 commonsourceibias.n253 gnd 0.011574f
C5598 commonsourceibias.n254 gnd 0.009462f
C5599 commonsourceibias.n255 gnd 0.009462f
C5600 commonsourceibias.n256 gnd 0.009462f
C5601 commonsourceibias.n257 gnd 0.011258f
C5602 commonsourceibias.n258 gnd 0.013056f
C5603 commonsourceibias.n259 gnd 0.070538f
C5604 commonsourceibias.n260 gnd 0.012977f
C5605 commonsourceibias.n261 gnd 0.009462f
C5606 commonsourceibias.n262 gnd 0.009462f
C5607 commonsourceibias.n263 gnd 0.009462f
C5608 commonsourceibias.n264 gnd 0.012818f
C5609 commonsourceibias.n265 gnd 0.070538f
C5610 commonsourceibias.n266 gnd 0.012902f
C5611 commonsourceibias.n267 gnd 0.011663f
C5612 commonsourceibias.n268 gnd 0.009462f
C5613 commonsourceibias.n269 gnd 0.009462f
C5614 commonsourceibias.n270 gnd 0.009462f
C5615 commonsourceibias.n271 gnd 0.010756f
C5616 commonsourceibias.n272 gnd 0.013095f
C5617 commonsourceibias.n273 gnd 0.070538f
C5618 commonsourceibias.n274 gnd 0.013039f
C5619 commonsourceibias.n275 gnd 0.009462f
C5620 commonsourceibias.n276 gnd 0.009462f
C5621 commonsourceibias.n277 gnd 0.009462f
C5622 commonsourceibias.n278 gnd 0.012719f
C5623 commonsourceibias.n279 gnd 0.070538f
C5624 commonsourceibias.n280 gnd 0.01275f
C5625 commonsourceibias.n281 gnd 0.085058f
C5626 commonsourceibias.n282 gnd 0.030353f
C5627 commonsourceibias.n283 gnd 0.151535f
C5628 commonsourceibias.n284 gnd 0.012626f
C5629 commonsourceibias.t68 gnd 0.176786f
C5630 commonsourceibias.n285 gnd 0.007691f
C5631 commonsourceibias.n286 gnd 0.009462f
C5632 commonsourceibias.t80 gnd 0.176786f
C5633 commonsourceibias.n287 gnd 0.009599f
C5634 commonsourceibias.n288 gnd 0.009462f
C5635 commonsourceibias.t134 gnd 0.176786f
C5636 commonsourceibias.n289 gnd 0.070538f
C5637 commonsourceibias.t159 gnd 0.176786f
C5638 commonsourceibias.n290 gnd 0.007654f
C5639 commonsourceibias.n291 gnd 0.009462f
C5640 commonsourceibias.t74 gnd 0.176786f
C5641 commonsourceibias.n292 gnd 0.009135f
C5642 commonsourceibias.n293 gnd 0.009462f
C5643 commonsourceibias.t120 gnd 0.176786f
C5644 commonsourceibias.n294 gnd 0.070538f
C5645 commonsourceibias.t111 gnd 0.176786f
C5646 commonsourceibias.n295 gnd 0.007642f
C5647 commonsourceibias.n296 gnd 0.009462f
C5648 commonsourceibias.t67 gnd 0.176786f
C5649 commonsourceibias.t81 gnd 0.176786f
C5650 commonsourceibias.n297 gnd 0.070538f
C5651 commonsourceibias.n298 gnd 0.009462f
C5652 commonsourceibias.t101 gnd 0.176786f
C5653 commonsourceibias.n299 gnd 0.070538f
C5654 commonsourceibias.n300 gnd 0.009462f
C5655 commonsourceibias.t158 gnd 0.176786f
C5656 commonsourceibias.n301 gnd 0.070538f
C5657 commonsourceibias.n302 gnd 0.009462f
C5658 commonsourceibias.t150 gnd 0.176786f
C5659 commonsourceibias.n303 gnd 0.010756f
C5660 commonsourceibias.n304 gnd 0.009462f
C5661 commonsourceibias.t70 gnd 0.176786f
C5662 commonsourceibias.n305 gnd 0.012719f
C5663 commonsourceibias.t136 gnd 0.196936f
C5664 commonsourceibias.t143 gnd 0.176786f
C5665 commonsourceibias.n306 gnd 0.078597f
C5666 commonsourceibias.n307 gnd 0.084205f
C5667 commonsourceibias.n308 gnd 0.040277f
C5668 commonsourceibias.n309 gnd 0.009462f
C5669 commonsourceibias.n310 gnd 0.007691f
C5670 commonsourceibias.n311 gnd 0.013039f
C5671 commonsourceibias.n312 gnd 0.070538f
C5672 commonsourceibias.n313 gnd 0.013095f
C5673 commonsourceibias.n314 gnd 0.009462f
C5674 commonsourceibias.n315 gnd 0.009462f
C5675 commonsourceibias.n316 gnd 0.009462f
C5676 commonsourceibias.n317 gnd 0.009599f
C5677 commonsourceibias.n318 gnd 0.070538f
C5678 commonsourceibias.n319 gnd 0.011663f
C5679 commonsourceibias.n320 gnd 0.012902f
C5680 commonsourceibias.n321 gnd 0.009462f
C5681 commonsourceibias.n322 gnd 0.009462f
C5682 commonsourceibias.n323 gnd 0.012818f
C5683 commonsourceibias.n324 gnd 0.007654f
C5684 commonsourceibias.n325 gnd 0.012977f
C5685 commonsourceibias.n326 gnd 0.009462f
C5686 commonsourceibias.n327 gnd 0.009462f
C5687 commonsourceibias.n328 gnd 0.013056f
C5688 commonsourceibias.n329 gnd 0.011258f
C5689 commonsourceibias.n330 gnd 0.009135f
C5690 commonsourceibias.n331 gnd 0.009462f
C5691 commonsourceibias.n332 gnd 0.009462f
C5692 commonsourceibias.n333 gnd 0.011574f
C5693 commonsourceibias.n334 gnd 0.012991f
C5694 commonsourceibias.n335 gnd 0.070538f
C5695 commonsourceibias.n336 gnd 0.012903f
C5696 commonsourceibias.n337 gnd 0.009462f
C5697 commonsourceibias.n338 gnd 0.009462f
C5698 commonsourceibias.n339 gnd 0.009462f
C5699 commonsourceibias.n340 gnd 0.012903f
C5700 commonsourceibias.n341 gnd 0.070538f
C5701 commonsourceibias.n342 gnd 0.012991f
C5702 commonsourceibias.n343 gnd 0.011574f
C5703 commonsourceibias.n344 gnd 0.009462f
C5704 commonsourceibias.n345 gnd 0.009462f
C5705 commonsourceibias.n346 gnd 0.009462f
C5706 commonsourceibias.n347 gnd 0.011258f
C5707 commonsourceibias.n348 gnd 0.013056f
C5708 commonsourceibias.n349 gnd 0.070538f
C5709 commonsourceibias.n350 gnd 0.012977f
C5710 commonsourceibias.n351 gnd 0.009462f
C5711 commonsourceibias.n352 gnd 0.009462f
C5712 commonsourceibias.n353 gnd 0.009462f
C5713 commonsourceibias.n354 gnd 0.012818f
C5714 commonsourceibias.n355 gnd 0.070538f
C5715 commonsourceibias.n356 gnd 0.012902f
C5716 commonsourceibias.n357 gnd 0.011663f
C5717 commonsourceibias.n358 gnd 0.009462f
C5718 commonsourceibias.n359 gnd 0.009462f
C5719 commonsourceibias.n360 gnd 0.009462f
C5720 commonsourceibias.n361 gnd 0.010756f
C5721 commonsourceibias.n362 gnd 0.013095f
C5722 commonsourceibias.n363 gnd 0.070538f
C5723 commonsourceibias.n364 gnd 0.013039f
C5724 commonsourceibias.n365 gnd 0.009462f
C5725 commonsourceibias.n366 gnd 0.009462f
C5726 commonsourceibias.n367 gnd 0.009462f
C5727 commonsourceibias.n368 gnd 0.012719f
C5728 commonsourceibias.n369 gnd 0.070538f
C5729 commonsourceibias.n370 gnd 0.01275f
C5730 commonsourceibias.t148 gnd 0.191194f
C5731 commonsourceibias.n371 gnd 0.085058f
C5732 commonsourceibias.n372 gnd 0.030353f
C5733 commonsourceibias.n373 gnd 0.53129f
C5734 commonsourceibias.n374 gnd 0.012626f
C5735 commonsourceibias.t153 gnd 0.191194f
C5736 commonsourceibias.t104 gnd 0.176786f
C5737 commonsourceibias.n375 gnd 0.007691f
C5738 commonsourceibias.n376 gnd 0.009462f
C5739 commonsourceibias.t73 gnd 0.176786f
C5740 commonsourceibias.n377 gnd 0.009599f
C5741 commonsourceibias.n378 gnd 0.009462f
C5742 commonsourceibias.t90 gnd 0.176786f
C5743 commonsourceibias.n379 gnd 0.007654f
C5744 commonsourceibias.n380 gnd 0.009462f
C5745 commonsourceibias.t151 gnd 0.176786f
C5746 commonsourceibias.n381 gnd 0.009135f
C5747 commonsourceibias.n382 gnd 0.009462f
C5748 commonsourceibias.t91 gnd 0.176786f
C5749 commonsourceibias.n383 gnd 0.007642f
C5750 commonsourceibias.n384 gnd 0.009462f
C5751 commonsourceibias.t119 gnd 0.176786f
C5752 commonsourceibias.t87 gnd 0.176786f
C5753 commonsourceibias.n385 gnd 0.070538f
C5754 commonsourceibias.n386 gnd 0.009462f
C5755 commonsourceibias.t79 gnd 0.176786f
C5756 commonsourceibias.n387 gnd 0.070538f
C5757 commonsourceibias.n388 gnd 0.009462f
C5758 commonsourceibias.t95 gnd 0.176786f
C5759 commonsourceibias.n389 gnd 0.070538f
C5760 commonsourceibias.n390 gnd 0.009462f
C5761 commonsourceibias.t88 gnd 0.176786f
C5762 commonsourceibias.n391 gnd 0.010756f
C5763 commonsourceibias.n392 gnd 0.009462f
C5764 commonsourceibias.t65 gnd 0.176786f
C5765 commonsourceibias.n393 gnd 0.012719f
C5766 commonsourceibias.t83 gnd 0.196936f
C5767 commonsourceibias.t84 gnd 0.176786f
C5768 commonsourceibias.n394 gnd 0.078597f
C5769 commonsourceibias.n395 gnd 0.084205f
C5770 commonsourceibias.n396 gnd 0.040277f
C5771 commonsourceibias.n397 gnd 0.009462f
C5772 commonsourceibias.n398 gnd 0.007691f
C5773 commonsourceibias.n399 gnd 0.013039f
C5774 commonsourceibias.n400 gnd 0.070538f
C5775 commonsourceibias.n401 gnd 0.013095f
C5776 commonsourceibias.n402 gnd 0.009462f
C5777 commonsourceibias.n403 gnd 0.009462f
C5778 commonsourceibias.n404 gnd 0.009462f
C5779 commonsourceibias.n405 gnd 0.009599f
C5780 commonsourceibias.n406 gnd 0.070538f
C5781 commonsourceibias.n407 gnd 0.011663f
C5782 commonsourceibias.n408 gnd 0.012902f
C5783 commonsourceibias.n409 gnd 0.009462f
C5784 commonsourceibias.n410 gnd 0.009462f
C5785 commonsourceibias.n411 gnd 0.012818f
C5786 commonsourceibias.n412 gnd 0.007654f
C5787 commonsourceibias.n413 gnd 0.012977f
C5788 commonsourceibias.n414 gnd 0.009462f
C5789 commonsourceibias.n415 gnd 0.009462f
C5790 commonsourceibias.n416 gnd 0.013056f
C5791 commonsourceibias.n417 gnd 0.011258f
C5792 commonsourceibias.n418 gnd 0.009135f
C5793 commonsourceibias.n419 gnd 0.009462f
C5794 commonsourceibias.n420 gnd 0.009462f
C5795 commonsourceibias.n421 gnd 0.011574f
C5796 commonsourceibias.n422 gnd 0.012991f
C5797 commonsourceibias.n423 gnd 0.070538f
C5798 commonsourceibias.n424 gnd 0.012903f
C5799 commonsourceibias.n425 gnd 0.009417f
C5800 commonsourceibias.t61 gnd 0.020419f
C5801 commonsourceibias.t59 gnd 0.020419f
C5802 commonsourceibias.n426 gnd 0.181032f
C5803 commonsourceibias.t39 gnd 0.020419f
C5804 commonsourceibias.t55 gnd 0.020419f
C5805 commonsourceibias.n427 gnd 0.180428f
C5806 commonsourceibias.n428 gnd 0.168125f
C5807 commonsourceibias.t7 gnd 0.020419f
C5808 commonsourceibias.t19 gnd 0.020419f
C5809 commonsourceibias.n429 gnd 0.180428f
C5810 commonsourceibias.n430 gnd 0.082878f
C5811 commonsourceibias.t57 gnd 0.020419f
C5812 commonsourceibias.t31 gnd 0.020419f
C5813 commonsourceibias.n431 gnd 0.180428f
C5814 commonsourceibias.n432 gnd 0.06924f
C5815 commonsourceibias.n433 gnd 0.012626f
C5816 commonsourceibias.t2 gnd 0.176786f
C5817 commonsourceibias.n434 gnd 0.007691f
C5818 commonsourceibias.n435 gnd 0.009462f
C5819 commonsourceibias.t14 gnd 0.176786f
C5820 commonsourceibias.n436 gnd 0.009599f
C5821 commonsourceibias.n437 gnd 0.009462f
C5822 commonsourceibias.t12 gnd 0.176786f
C5823 commonsourceibias.n438 gnd 0.007654f
C5824 commonsourceibias.n439 gnd 0.009462f
C5825 commonsourceibias.t46 gnd 0.176786f
C5826 commonsourceibias.n440 gnd 0.009135f
C5827 commonsourceibias.n441 gnd 0.009462f
C5828 commonsourceibias.t10 gnd 0.176786f
C5829 commonsourceibias.n442 gnd 0.007642f
C5830 commonsourceibias.n443 gnd 0.009462f
C5831 commonsourceibias.t30 gnd 0.176786f
C5832 commonsourceibias.t56 gnd 0.176786f
C5833 commonsourceibias.n444 gnd 0.070538f
C5834 commonsourceibias.n445 gnd 0.009462f
C5835 commonsourceibias.t18 gnd 0.176786f
C5836 commonsourceibias.n446 gnd 0.070538f
C5837 commonsourceibias.n447 gnd 0.009462f
C5838 commonsourceibias.t6 gnd 0.176786f
C5839 commonsourceibias.n448 gnd 0.070538f
C5840 commonsourceibias.n449 gnd 0.009462f
C5841 commonsourceibias.t54 gnd 0.176786f
C5842 commonsourceibias.n450 gnd 0.010756f
C5843 commonsourceibias.n451 gnd 0.009462f
C5844 commonsourceibias.t38 gnd 0.176786f
C5845 commonsourceibias.n452 gnd 0.012719f
C5846 commonsourceibias.t60 gnd 0.196936f
C5847 commonsourceibias.t58 gnd 0.176786f
C5848 commonsourceibias.n453 gnd 0.078597f
C5849 commonsourceibias.n454 gnd 0.084205f
C5850 commonsourceibias.n455 gnd 0.040277f
C5851 commonsourceibias.n456 gnd 0.009462f
C5852 commonsourceibias.n457 gnd 0.007691f
C5853 commonsourceibias.n458 gnd 0.013039f
C5854 commonsourceibias.n459 gnd 0.070538f
C5855 commonsourceibias.n460 gnd 0.013095f
C5856 commonsourceibias.n461 gnd 0.009462f
C5857 commonsourceibias.n462 gnd 0.009462f
C5858 commonsourceibias.n463 gnd 0.009462f
C5859 commonsourceibias.n464 gnd 0.009599f
C5860 commonsourceibias.n465 gnd 0.070538f
C5861 commonsourceibias.n466 gnd 0.011663f
C5862 commonsourceibias.n467 gnd 0.012902f
C5863 commonsourceibias.n468 gnd 0.009462f
C5864 commonsourceibias.n469 gnd 0.009462f
C5865 commonsourceibias.n470 gnd 0.012818f
C5866 commonsourceibias.n471 gnd 0.007654f
C5867 commonsourceibias.n472 gnd 0.012977f
C5868 commonsourceibias.n473 gnd 0.009462f
C5869 commonsourceibias.n474 gnd 0.009462f
C5870 commonsourceibias.n475 gnd 0.013056f
C5871 commonsourceibias.n476 gnd 0.011258f
C5872 commonsourceibias.n477 gnd 0.009135f
C5873 commonsourceibias.n478 gnd 0.009462f
C5874 commonsourceibias.n479 gnd 0.009462f
C5875 commonsourceibias.n480 gnd 0.011574f
C5876 commonsourceibias.n481 gnd 0.012991f
C5877 commonsourceibias.n482 gnd 0.070538f
C5878 commonsourceibias.n483 gnd 0.012903f
C5879 commonsourceibias.n484 gnd 0.009462f
C5880 commonsourceibias.n485 gnd 0.009462f
C5881 commonsourceibias.n486 gnd 0.009462f
C5882 commonsourceibias.n487 gnd 0.012903f
C5883 commonsourceibias.n488 gnd 0.070538f
C5884 commonsourceibias.n489 gnd 0.012991f
C5885 commonsourceibias.t16 gnd 0.176786f
C5886 commonsourceibias.n490 gnd 0.070538f
C5887 commonsourceibias.n491 gnd 0.011574f
C5888 commonsourceibias.n492 gnd 0.009462f
C5889 commonsourceibias.n493 gnd 0.009462f
C5890 commonsourceibias.n494 gnd 0.009462f
C5891 commonsourceibias.n495 gnd 0.011258f
C5892 commonsourceibias.n496 gnd 0.013056f
C5893 commonsourceibias.n497 gnd 0.070538f
C5894 commonsourceibias.n498 gnd 0.012977f
C5895 commonsourceibias.n499 gnd 0.009462f
C5896 commonsourceibias.n500 gnd 0.009462f
C5897 commonsourceibias.n501 gnd 0.009462f
C5898 commonsourceibias.n502 gnd 0.012818f
C5899 commonsourceibias.n503 gnd 0.070538f
C5900 commonsourceibias.n504 gnd 0.012902f
C5901 commonsourceibias.t28 gnd 0.176786f
C5902 commonsourceibias.n505 gnd 0.070538f
C5903 commonsourceibias.n506 gnd 0.011663f
C5904 commonsourceibias.n507 gnd 0.009462f
C5905 commonsourceibias.n508 gnd 0.009462f
C5906 commonsourceibias.n509 gnd 0.009462f
C5907 commonsourceibias.n510 gnd 0.010756f
C5908 commonsourceibias.n511 gnd 0.013095f
C5909 commonsourceibias.n512 gnd 0.070538f
C5910 commonsourceibias.n513 gnd 0.013039f
C5911 commonsourceibias.n514 gnd 0.009462f
C5912 commonsourceibias.n515 gnd 0.009462f
C5913 commonsourceibias.n516 gnd 0.009462f
C5914 commonsourceibias.n517 gnd 0.012719f
C5915 commonsourceibias.n518 gnd 0.070538f
C5916 commonsourceibias.n519 gnd 0.01275f
C5917 commonsourceibias.t44 gnd 0.191194f
C5918 commonsourceibias.n520 gnd 0.085058f
C5919 commonsourceibias.n521 gnd 0.095108f
C5920 commonsourceibias.t3 gnd 0.020419f
C5921 commonsourceibias.t45 gnd 0.020419f
C5922 commonsourceibias.n522 gnd 0.180428f
C5923 commonsourceibias.n523 gnd 0.15629f
C5924 commonsourceibias.t29 gnd 0.020419f
C5925 commonsourceibias.t15 gnd 0.020419f
C5926 commonsourceibias.n524 gnd 0.180428f
C5927 commonsourceibias.n525 gnd 0.082878f
C5928 commonsourceibias.t47 gnd 0.020419f
C5929 commonsourceibias.t13 gnd 0.020419f
C5930 commonsourceibias.n526 gnd 0.180428f
C5931 commonsourceibias.n527 gnd 0.082878f
C5932 commonsourceibias.t11 gnd 0.020419f
C5933 commonsourceibias.t17 gnd 0.020419f
C5934 commonsourceibias.n528 gnd 0.180428f
C5935 commonsourceibias.n529 gnd 0.06924f
C5936 commonsourceibias.n530 gnd 0.083843f
C5937 commonsourceibias.n531 gnd 0.068402f
C5938 commonsourceibias.n532 gnd 0.009417f
C5939 commonsourceibias.n533 gnd 0.012903f
C5940 commonsourceibias.n534 gnd 0.070538f
C5941 commonsourceibias.n535 gnd 0.012991f
C5942 commonsourceibias.t102 gnd 0.176786f
C5943 commonsourceibias.n536 gnd 0.070538f
C5944 commonsourceibias.n537 gnd 0.011574f
C5945 commonsourceibias.n538 gnd 0.009462f
C5946 commonsourceibias.n539 gnd 0.009462f
C5947 commonsourceibias.n540 gnd 0.009462f
C5948 commonsourceibias.n541 gnd 0.011258f
C5949 commonsourceibias.n542 gnd 0.013056f
C5950 commonsourceibias.n543 gnd 0.070538f
C5951 commonsourceibias.n544 gnd 0.012977f
C5952 commonsourceibias.n545 gnd 0.009462f
C5953 commonsourceibias.n546 gnd 0.009462f
C5954 commonsourceibias.n547 gnd 0.009462f
C5955 commonsourceibias.n548 gnd 0.012818f
C5956 commonsourceibias.n549 gnd 0.070538f
C5957 commonsourceibias.n550 gnd 0.012902f
C5958 commonsourceibias.t121 gnd 0.176786f
C5959 commonsourceibias.n551 gnd 0.070538f
C5960 commonsourceibias.n552 gnd 0.011663f
C5961 commonsourceibias.n553 gnd 0.009462f
C5962 commonsourceibias.n554 gnd 0.009462f
C5963 commonsourceibias.n555 gnd 0.009462f
C5964 commonsourceibias.n556 gnd 0.010756f
C5965 commonsourceibias.n557 gnd 0.013095f
C5966 commonsourceibias.n558 gnd 0.070538f
C5967 commonsourceibias.n559 gnd 0.013039f
C5968 commonsourceibias.n560 gnd 0.009462f
C5969 commonsourceibias.n561 gnd 0.009462f
C5970 commonsourceibias.n562 gnd 0.009462f
C5971 commonsourceibias.n563 gnd 0.012719f
C5972 commonsourceibias.n564 gnd 0.070538f
C5973 commonsourceibias.n565 gnd 0.01275f
C5974 commonsourceibias.n566 gnd 0.085058f
C5975 commonsourceibias.n567 gnd 0.056191f
C5976 commonsourceibias.n568 gnd 0.012626f
C5977 commonsourceibias.t118 gnd 0.176786f
C5978 commonsourceibias.n569 gnd 0.007691f
C5979 commonsourceibias.n570 gnd 0.009462f
C5980 commonsourceibias.t109 gnd 0.176786f
C5981 commonsourceibias.n571 gnd 0.009599f
C5982 commonsourceibias.n572 gnd 0.009462f
C5983 commonsourceibias.t117 gnd 0.176786f
C5984 commonsourceibias.n573 gnd 0.007654f
C5985 commonsourceibias.n574 gnd 0.009462f
C5986 commonsourceibias.t108 gnd 0.176786f
C5987 commonsourceibias.n575 gnd 0.009135f
C5988 commonsourceibias.n576 gnd 0.009462f
C5989 commonsourceibias.t122 gnd 0.176786f
C5990 commonsourceibias.n577 gnd 0.007642f
C5991 commonsourceibias.n578 gnd 0.009462f
C5992 commonsourceibias.t107 gnd 0.176786f
C5993 commonsourceibias.t129 gnd 0.176786f
C5994 commonsourceibias.n579 gnd 0.070538f
C5995 commonsourceibias.n580 gnd 0.009462f
C5996 commonsourceibias.t156 gnd 0.176786f
C5997 commonsourceibias.n581 gnd 0.070538f
C5998 commonsourceibias.n582 gnd 0.009462f
C5999 commonsourceibias.t105 gnd 0.176786f
C6000 commonsourceibias.n583 gnd 0.070538f
C6001 commonsourceibias.n584 gnd 0.009462f
C6002 commonsourceibias.t137 gnd 0.176786f
C6003 commonsourceibias.n585 gnd 0.010756f
C6004 commonsourceibias.n586 gnd 0.009462f
C6005 commonsourceibias.t155 gnd 0.176786f
C6006 commonsourceibias.n587 gnd 0.012719f
C6007 commonsourceibias.t131 gnd 0.196936f
C6008 commonsourceibias.t142 gnd 0.176786f
C6009 commonsourceibias.n588 gnd 0.078597f
C6010 commonsourceibias.n589 gnd 0.084205f
C6011 commonsourceibias.n590 gnd 0.040277f
C6012 commonsourceibias.n591 gnd 0.009462f
C6013 commonsourceibias.n592 gnd 0.007691f
C6014 commonsourceibias.n593 gnd 0.013039f
C6015 commonsourceibias.n594 gnd 0.070538f
C6016 commonsourceibias.n595 gnd 0.013095f
C6017 commonsourceibias.n596 gnd 0.009462f
C6018 commonsourceibias.n597 gnd 0.009462f
C6019 commonsourceibias.n598 gnd 0.009462f
C6020 commonsourceibias.n599 gnd 0.009599f
C6021 commonsourceibias.n600 gnd 0.070538f
C6022 commonsourceibias.n601 gnd 0.011663f
C6023 commonsourceibias.n602 gnd 0.012902f
C6024 commonsourceibias.n603 gnd 0.009462f
C6025 commonsourceibias.n604 gnd 0.009462f
C6026 commonsourceibias.n605 gnd 0.012818f
C6027 commonsourceibias.n606 gnd 0.007654f
C6028 commonsourceibias.n607 gnd 0.012977f
C6029 commonsourceibias.n608 gnd 0.009462f
C6030 commonsourceibias.n609 gnd 0.009462f
C6031 commonsourceibias.n610 gnd 0.013056f
C6032 commonsourceibias.n611 gnd 0.011258f
C6033 commonsourceibias.n612 gnd 0.009135f
C6034 commonsourceibias.n613 gnd 0.009462f
C6035 commonsourceibias.n614 gnd 0.009462f
C6036 commonsourceibias.n615 gnd 0.011574f
C6037 commonsourceibias.n616 gnd 0.012991f
C6038 commonsourceibias.n617 gnd 0.070538f
C6039 commonsourceibias.n618 gnd 0.012903f
C6040 commonsourceibias.n619 gnd 0.009462f
C6041 commonsourceibias.n620 gnd 0.009462f
C6042 commonsourceibias.n621 gnd 0.009462f
C6043 commonsourceibias.n622 gnd 0.012903f
C6044 commonsourceibias.n623 gnd 0.070538f
C6045 commonsourceibias.n624 gnd 0.012991f
C6046 commonsourceibias.t130 gnd 0.176786f
C6047 commonsourceibias.n625 gnd 0.070538f
C6048 commonsourceibias.n626 gnd 0.011574f
C6049 commonsourceibias.n627 gnd 0.009462f
C6050 commonsourceibias.n628 gnd 0.009462f
C6051 commonsourceibias.n629 gnd 0.009462f
C6052 commonsourceibias.n630 gnd 0.011258f
C6053 commonsourceibias.n631 gnd 0.013056f
C6054 commonsourceibias.n632 gnd 0.070538f
C6055 commonsourceibias.n633 gnd 0.012977f
C6056 commonsourceibias.n634 gnd 0.009462f
C6057 commonsourceibias.n635 gnd 0.009462f
C6058 commonsourceibias.n636 gnd 0.009462f
C6059 commonsourceibias.n637 gnd 0.012818f
C6060 commonsourceibias.n638 gnd 0.070538f
C6061 commonsourceibias.n639 gnd 0.012902f
C6062 commonsourceibias.t99 gnd 0.176786f
C6063 commonsourceibias.n640 gnd 0.070538f
C6064 commonsourceibias.n641 gnd 0.011663f
C6065 commonsourceibias.n642 gnd 0.009462f
C6066 commonsourceibias.n643 gnd 0.009462f
C6067 commonsourceibias.n644 gnd 0.009462f
C6068 commonsourceibias.n645 gnd 0.010756f
C6069 commonsourceibias.n646 gnd 0.013095f
C6070 commonsourceibias.n647 gnd 0.070538f
C6071 commonsourceibias.n648 gnd 0.013039f
C6072 commonsourceibias.n649 gnd 0.009462f
C6073 commonsourceibias.n650 gnd 0.009462f
C6074 commonsourceibias.n651 gnd 0.009462f
C6075 commonsourceibias.n652 gnd 0.012719f
C6076 commonsourceibias.n653 gnd 0.070538f
C6077 commonsourceibias.n654 gnd 0.01275f
C6078 commonsourceibias.t100 gnd 0.191194f
C6079 commonsourceibias.n655 gnd 0.085058f
C6080 commonsourceibias.n656 gnd 0.030353f
C6081 commonsourceibias.n657 gnd 0.151535f
C6082 commonsourceibias.n658 gnd 0.012626f
C6083 commonsourceibias.t86 gnd 0.176786f
C6084 commonsourceibias.n659 gnd 0.007691f
C6085 commonsourceibias.n660 gnd 0.009462f
C6086 commonsourceibias.t97 gnd 0.176786f
C6087 commonsourceibias.n661 gnd 0.009599f
C6088 commonsourceibias.n662 gnd 0.009462f
C6089 commonsourceibias.t77 gnd 0.176786f
C6090 commonsourceibias.n663 gnd 0.007654f
C6091 commonsourceibias.n664 gnd 0.009462f
C6092 commonsourceibias.t93 gnd 0.176786f
C6093 commonsourceibias.n665 gnd 0.009135f
C6094 commonsourceibias.n666 gnd 0.009462f
C6095 commonsourceibias.t145 gnd 0.176786f
C6096 commonsourceibias.n667 gnd 0.007642f
C6097 commonsourceibias.n668 gnd 0.009462f
C6098 commonsourceibias.t85 gnd 0.176786f
C6099 commonsourceibias.t98 gnd 0.176786f
C6100 commonsourceibias.n669 gnd 0.070538f
C6101 commonsourceibias.n670 gnd 0.009462f
C6102 commonsourceibias.t94 gnd 0.176786f
C6103 commonsourceibias.n671 gnd 0.070538f
C6104 commonsourceibias.n672 gnd 0.009462f
C6105 commonsourceibias.t76 gnd 0.176786f
C6106 commonsourceibias.n673 gnd 0.070538f
C6107 commonsourceibias.n674 gnd 0.009462f
C6108 commonsourceibias.t72 gnd 0.176786f
C6109 commonsourceibias.n675 gnd 0.010756f
C6110 commonsourceibias.n676 gnd 0.009462f
C6111 commonsourceibias.t89 gnd 0.176786f
C6112 commonsourceibias.n677 gnd 0.012719f
C6113 commonsourceibias.t144 gnd 0.196936f
C6114 commonsourceibias.t133 gnd 0.176786f
C6115 commonsourceibias.n678 gnd 0.078597f
C6116 commonsourceibias.n679 gnd 0.084205f
C6117 commonsourceibias.n680 gnd 0.040277f
C6118 commonsourceibias.n681 gnd 0.009462f
C6119 commonsourceibias.n682 gnd 0.007691f
C6120 commonsourceibias.n683 gnd 0.013039f
C6121 commonsourceibias.n684 gnd 0.070538f
C6122 commonsourceibias.n685 gnd 0.013095f
C6123 commonsourceibias.n686 gnd 0.009462f
C6124 commonsourceibias.n687 gnd 0.009462f
C6125 commonsourceibias.n688 gnd 0.009462f
C6126 commonsourceibias.n689 gnd 0.009599f
C6127 commonsourceibias.n690 gnd 0.070538f
C6128 commonsourceibias.n691 gnd 0.011663f
C6129 commonsourceibias.n692 gnd 0.012902f
C6130 commonsourceibias.n693 gnd 0.009462f
C6131 commonsourceibias.n694 gnd 0.009462f
C6132 commonsourceibias.n695 gnd 0.012818f
C6133 commonsourceibias.n696 gnd 0.007654f
C6134 commonsourceibias.n697 gnd 0.012977f
C6135 commonsourceibias.n698 gnd 0.009462f
C6136 commonsourceibias.n699 gnd 0.009462f
C6137 commonsourceibias.n700 gnd 0.013056f
C6138 commonsourceibias.n701 gnd 0.011258f
C6139 commonsourceibias.n702 gnd 0.009135f
C6140 commonsourceibias.n703 gnd 0.009462f
C6141 commonsourceibias.n704 gnd 0.009462f
C6142 commonsourceibias.n705 gnd 0.011574f
C6143 commonsourceibias.n706 gnd 0.012991f
C6144 commonsourceibias.n707 gnd 0.070538f
C6145 commonsourceibias.n708 gnd 0.012903f
C6146 commonsourceibias.n709 gnd 0.009462f
C6147 commonsourceibias.n710 gnd 0.009462f
C6148 commonsourceibias.n711 gnd 0.009462f
C6149 commonsourceibias.n712 gnd 0.012903f
C6150 commonsourceibias.n713 gnd 0.070538f
C6151 commonsourceibias.n714 gnd 0.012991f
C6152 commonsourceibias.t103 gnd 0.176786f
C6153 commonsourceibias.n715 gnd 0.070538f
C6154 commonsourceibias.n716 gnd 0.011574f
C6155 commonsourceibias.n717 gnd 0.009462f
C6156 commonsourceibias.n718 gnd 0.009462f
C6157 commonsourceibias.n719 gnd 0.009462f
C6158 commonsourceibias.n720 gnd 0.011258f
C6159 commonsourceibias.n721 gnd 0.013056f
C6160 commonsourceibias.n722 gnd 0.070538f
C6161 commonsourceibias.n723 gnd 0.012977f
C6162 commonsourceibias.n724 gnd 0.009462f
C6163 commonsourceibias.n725 gnd 0.009462f
C6164 commonsourceibias.n726 gnd 0.009462f
C6165 commonsourceibias.n727 gnd 0.012818f
C6166 commonsourceibias.n728 gnd 0.070538f
C6167 commonsourceibias.n729 gnd 0.012902f
C6168 commonsourceibias.t66 gnd 0.176786f
C6169 commonsourceibias.n730 gnd 0.070538f
C6170 commonsourceibias.n731 gnd 0.011663f
C6171 commonsourceibias.n732 gnd 0.009462f
C6172 commonsourceibias.n733 gnd 0.009462f
C6173 commonsourceibias.n734 gnd 0.009462f
C6174 commonsourceibias.n735 gnd 0.010756f
C6175 commonsourceibias.n736 gnd 0.013095f
C6176 commonsourceibias.n737 gnd 0.070538f
C6177 commonsourceibias.n738 gnd 0.013039f
C6178 commonsourceibias.n739 gnd 0.009462f
C6179 commonsourceibias.n740 gnd 0.009462f
C6180 commonsourceibias.n741 gnd 0.009462f
C6181 commonsourceibias.n742 gnd 0.012719f
C6182 commonsourceibias.n743 gnd 0.070538f
C6183 commonsourceibias.n744 gnd 0.01275f
C6184 commonsourceibias.t71 gnd 0.191194f
C6185 commonsourceibias.n745 gnd 0.085058f
C6186 commonsourceibias.n746 gnd 0.030353f
C6187 commonsourceibias.n747 gnd 0.199689f
C6188 commonsourceibias.n748 gnd 5.4246f
.ends

