* NGSPICE file created from opamp297.ext - technology: sky130A

.subckt opamp297 gnd CSoutput output vdd plus minus commonsourceibias outputibias
+ diffpairibias
X0 gnd.t310 commonsourceibias.t64 CSoutput.t162 gnd.t191 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X1 CSoutput.t71 a_n8964_8799.t44 vdd.t292 vdd.t232 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=3.12 ps=16.78 w=8 l=0.5
X2 a_n2472_13878.t19 a_n2650_13878.t34 a_n2650_13878.t35 vdd.t9 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X3 commonsourceibias.t63 commonsourceibias.t62 gnd.t309 gnd.t279 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X4 a_n2472_13878.t27 a_n2650_13878.t64 vdd.t15 vdd.t14 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X5 CSoutput.t184 a_n2650_8322.t33 sky130_fd_pr__cap_mim_m3_1 l=12 w=12
X6 vdd.t291 a_n8964_8799.t45 CSoutput.t9 vdd.t226 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X7 CSoutput.t42 a_n8964_8799.t46 vdd.t290 vdd.t149 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X8 CSoutput.t40 a_n8964_8799.t47 vdd.t289 vdd.t141 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X9 gnd.t308 commonsourceibias.t65 CSoutput.t161 gnd.t274 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X10 gnd.t181 gnd.t179 gnd.t180 gnd.t79 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=0 ps=0 w=7 l=1
X11 gnd.t307 commonsourceibias.t60 commonsourceibias.t61 gnd.t185 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X12 vdd.t288 a_n8964_8799.t48 CSoutput.t174 vdd.t214 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X13 gnd.t306 commonsourceibias.t66 CSoutput.t160 gnd.t185 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X14 a_n2650_8322.t27 a_n2650_13878.t65 a_n8964_8799.t17 vdd.t16 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X15 CSoutput.t49 a_n8964_8799.t49 vdd.t287 vdd.t175 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X16 output.t17 CSoutput.t185 vdd.t36 gnd.t59 sky130_fd_pr__nfet_01v8 ad=0.825 pd=5.33 as=0.825 ps=5.33 w=5 l=1
X17 vdd.t286 a_n8964_8799.t50 CSoutput.t29 vdd.t272 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X18 gnd.t178 gnd.t176 gnd.t177 gnd.t126 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=0 ps=0 w=7 l=0.5
X19 CSoutput.t169 a_n8964_8799.t51 vdd.t285 vdd.t184 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X20 gnd.t175 gnd.t173 gnd.t174 gnd.t119 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=0 ps=0 w=7 l=0.5
X21 gnd.t172 gnd.t171 plus.t4 gnd.t126 sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.5
X22 a_n8964_8799.t30 plus.t5 a_n2903_n3924.t33 gnd.t68 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.5
X23 gnd.t305 commonsourceibias.t67 CSoutput.t159 gnd.t216 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X24 vdd.t284 a_n8964_8799.t52 CSoutput.t58 vdd.t272 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X25 vdd.t283 a_n8964_8799.t53 CSoutput.t167 vdd.t219 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X26 minus.t4 gnd.t168 gnd.t170 gnd.t169 sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.5
X27 gnd.t304 commonsourceibias.t8 commonsourceibias.t9 gnd.t228 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X28 a_n8964_8799.t36 a_n2650_13878.t66 a_n2650_8322.t26 vdd.t56 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X29 vdd.t282 a_n8964_8799.t54 CSoutput.t17 vdd.t137 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X30 vdd.t281 a_n8964_8799.t55 CSoutput.t166 vdd.t248 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X31 a_n8964_8799.t37 a_n2650_13878.t67 a_n2650_8322.t25 vdd.t293 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=3.51 ps=18.78 w=9 l=0.5
X32 output.t0 outputibias.t8 gnd.t37 gnd.t36 sky130_fd_pr__nfet_01v8 ad=2.34 pd=12.78 as=2.34 ps=12.78 w=6 l=2
X33 CSoutput.t186 a_n2650_8322.t32 sky130_fd_pr__cap_mim_m3_1 l=12 w=12
X34 a_n8964_8799.t38 plus.t6 a_n2903_n3924.t32 gnd.t9 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.5
X35 CSoutput.t106 commonsourceibias.t68 gnd.t303 gnd.t202 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X36 gnd.t167 gnd.t165 gnd.t166 gnd.t111 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=0 ps=0 w=7 l=1
X37 gnd.t302 commonsourceibias.t6 commonsourceibias.t7 gnd.t270 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X38 output.t1 outputibias.t9 gnd.t40 gnd.t39 sky130_fd_pr__nfet_01v8 ad=2.34 pd=12.78 as=2.34 ps=12.78 w=6 l=2
X39 CSoutput.t36 a_n8964_8799.t56 vdd.t280 vdd.t232 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=3.12 ps=16.78 w=8 l=0.5
X40 vdd.t33 CSoutput.t187 output.t16 gnd.t58 sky130_fd_pr__nfet_01v8 ad=0.825 pd=5.33 as=0.825 ps=5.33 w=5 l=1
X41 CSoutput.t105 commonsourceibias.t69 gnd.t301 gnd.t197 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X42 a_n2903_n3924.t4 diffpairibias.t16 gnd.t5 gnd.t4 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=2.73 ps=14.78 w=7 l=1
X43 a_n2903_n3924.t1 minus.t5 a_n2650_13878.t1 gnd.t1 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.5
X44 CSoutput.t12 a_n8964_8799.t57 vdd.t279 vdd.t198 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X45 a_n2903_n3924.t31 plus.t7 a_n8964_8799.t18 gnd.t38 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.5
X46 vdd.t278 a_n8964_8799.t58 CSoutput.t93 vdd.t137 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X47 a_n2650_13878.t57 minus.t6 a_n2903_n3924.t47 gnd.t43 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.5
X48 output.t19 outputibias.t10 gnd.t316 gnd.t315 sky130_fd_pr__nfet_01v8 ad=2.34 pd=12.78 as=2.34 ps=12.78 w=6 l=2
X49 CSoutput.t104 commonsourceibias.t70 gnd.t300 gnd.t193 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X50 a_n2903_n3924.t30 plus.t8 a_n8964_8799.t33 gnd.t31 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.5
X51 a_n2903_n3924.t42 minus.t7 a_n2650_13878.t55 gnd.t33 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.5
X52 CSoutput.t164 a_n8964_8799.t59 vdd.t277 vdd.t141 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X53 vdd.t276 a_n8964_8799.t60 CSoutput.t64 vdd.t214 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X54 vdd.t132 vdd.t130 vdd.t131 vdd.t66 sky130_fd_pr__pfet_01v8 ad=3.51 pd=18.78 as=0 ps=0 w=9 l=0.5
X55 output.t15 CSoutput.t188 vdd.t22 gnd.t57 sky130_fd_pr__nfet_01v8 ad=1.95 pd=10.78 as=0.825 ps=5.33 w=5 l=1
X56 gnd.t299 commonsourceibias.t4 commonsourceibias.t5 gnd.t236 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=1.155 ps=7.33 w=7 l=1
X57 a_n2472_13878.t18 a_n2650_13878.t8 a_n2650_13878.t9 vdd.t20 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X58 CSoutput.t103 commonsourceibias.t71 gnd.t298 gnd.t279 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X59 a_n2650_13878.t15 a_n2650_13878.t14 a_n2472_13878.t17 vdd.t39 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X60 CSoutput.t2 a_n8964_8799.t61 vdd.t275 vdd.t184 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X61 vdd.t129 vdd.t127 vdd.t128 vdd.t104 sky130_fd_pr__pfet_01v8 ad=3.51 pd=18.78 as=0 ps=0 w=9 l=0.5
X62 a_n2903_n3924.t37 minus.t8 a_n2650_13878.t50 gnd.t30 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.5
X63 vdd.t274 a_n8964_8799.t62 CSoutput.t74 vdd.t219 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X64 vdd.t273 a_n8964_8799.t63 CSoutput.t1 vdd.t272 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X65 diffpairibias.t15 diffpairibias.t14 gnd.t312 gnd.t311 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=2.73 ps=14.78 w=7 l=1
X66 a_n2650_13878.t11 a_n2650_13878.t10 a_n2472_13878.t16 vdd.t6 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X67 CSoutput.t35 a_n8964_8799.t64 vdd.t271 vdd.t245 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X68 vdd.t270 a_n8964_8799.t65 CSoutput.t91 vdd.t181 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X69 a_n8964_8799.t40 a_n2650_13878.t68 a_n2650_8322.t24 vdd.t4 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X70 CSoutput.t62 a_n8964_8799.t66 vdd.t269 vdd.t230 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X71 a_n2650_13878.t48 minus.t9 a_n2903_n3924.t35 gnd.t26 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=2.73 ps=14.78 w=7 l=0.5
X72 a_n2650_13878.t45 a_n2650_13878.t44 a_n2472_13878.t15 vdd.t18 sky130_fd_pr__pfet_01v8 ad=3.51 pd=18.78 as=1.485 ps=9.33 w=9 l=0.5
X73 gnd.t164 gnd.t162 plus.t3 gnd.t163 sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.39 ps=2.78 w=1 l=0.5
X74 vdd.t268 a_n8964_8799.t67 CSoutput.t46 vdd.t153 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X75 vdd.t267 a_n8964_8799.t68 CSoutput.t54 vdd.t248 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X76 a_n8964_8799.t41 a_n2650_13878.t69 a_n2650_8322.t23 vdd.t55 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=3.51 ps=18.78 w=9 l=0.5
X77 gnd.t297 commonsourceibias.t72 CSoutput.t102 gnd.t274 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X78 diffpairibias.t13 diffpairibias.t12 gnd.t35 gnd.t34 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=2.73 ps=14.78 w=7 l=1
X79 gnd.t296 commonsourceibias.t73 CSoutput.t101 gnd.t183 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X80 CSoutput.t72 a_n8964_8799.t69 vdd.t266 vdd.t160 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X81 output.t14 CSoutput.t189 vdd.t34 gnd.t56 sky130_fd_pr__nfet_01v8 ad=0.825 pd=5.33 as=0.825 ps=5.33 w=5 l=1
X82 commonsourceibias.t3 commonsourceibias.t2 gnd.t295 gnd.t202 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X83 vdd.t24 CSoutput.t190 output.t13 gnd.t55 sky130_fd_pr__nfet_01v8 ad=0.825 pd=5.33 as=1.95 ps=10.78 w=5 l=1
X84 gnd.t294 commonsourceibias.t74 CSoutput.t100 gnd.t270 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X85 a_n2650_8322.t22 a_n2650_13878.t70 a_n8964_8799.t20 vdd.t18 sky130_fd_pr__pfet_01v8 ad=3.51 pd=18.78 as=1.485 ps=9.33 w=9 l=0.5
X86 CSoutput.t7 a_n8964_8799.t70 vdd.t265 vdd.t202 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X87 commonsourceibias.t1 commonsourceibias.t0 gnd.t293 gnd.t230 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X88 gnd.t292 commonsourceibias.t75 CSoutput.t99 gnd.t216 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X89 CSoutput.t191 a_n2650_8322.t31 sky130_fd_pr__cap_mim_m3_1 l=12 w=12
X90 plus.t2 gnd.t159 gnd.t161 gnd.t160 sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.5
X91 commonsourceibias.t59 commonsourceibias.t58 gnd.t291 gnd.t218 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X92 a_n8964_8799.t1 plus.t9 a_n2903_n3924.t29 gnd.t13 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.5
X93 gnd.t290 commonsourceibias.t76 CSoutput.t158 gnd.t267 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X94 CSoutput.t157 commonsourceibias.t77 gnd.t289 gnd.t264 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=2.73 ps=14.78 w=7 l=1
X95 vdd.t126 vdd.t124 vdd.t125 vdd.t100 sky130_fd_pr__pfet_01v8 ad=3.12 pd=16.78 as=0 ps=0 w=8 l=0.5
X96 gnd.t288 commonsourceibias.t56 commonsourceibias.t57 gnd.t267 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X97 a_n2903_n3924.t9 diffpairibias.t17 gnd.t12 gnd.t11 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=2.73 ps=14.78 w=7 l=1
X98 vdd.t264 a_n8964_8799.t71 CSoutput.t52 vdd.t217 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X99 a_n2903_n3924.t3 minus.t10 a_n2650_13878.t3 gnd.t3 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.5
X100 vdd.t263 a_n8964_8799.t72 CSoutput.t97 vdd.t252 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X101 a_n2650_13878.t27 a_n2650_13878.t26 a_n2472_13878.t14 vdd.t16 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X102 vdd.t262 a_n8964_8799.t73 CSoutput.t45 vdd.t192 sky130_fd_pr__pfet_01v8 ad=3.12 pd=16.78 as=1.32 ps=8.33 w=8 l=0.5
X103 vdd.t261 a_n8964_8799.t74 CSoutput.t5 vdd.t224 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X104 a_n8964_8799.t21 a_n2650_13878.t71 a_n2650_8322.t21 vdd.t5 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X105 a_n2650_13878.t31 a_n2650_13878.t30 a_n2472_13878.t13 vdd.t11 sky130_fd_pr__pfet_01v8 ad=3.51 pd=18.78 as=1.485 ps=9.33 w=9 l=0.5
X106 gnd.t287 commonsourceibias.t54 commonsourceibias.t55 gnd.t257 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=1.155 ps=7.33 w=7 l=1
X107 a_n2650_13878.t54 minus.t11 a_n2903_n3924.t41 gnd.t15 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.5
X108 gnd.t158 gnd.t156 gnd.t157 gnd.t111 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=0 ps=0 w=7 l=1
X109 a_n2903_n3924.t28 plus.t10 a_n8964_8799.t4 gnd.t7 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.5
X110 commonsourceibias.t53 commonsourceibias.t52 gnd.t286 gnd.t193 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X111 CSoutput.t156 commonsourceibias.t78 gnd.t285 gnd.t197 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X112 vdd.t260 a_n8964_8799.t75 CSoutput.t6 vdd.t158 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X113 CSoutput.t10 a_n8964_8799.t76 vdd.t259 vdd.t245 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X114 CSoutput.t21 a_n8964_8799.t77 vdd.t258 vdd.t196 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X115 CSoutput.t155 commonsourceibias.t79 gnd.t284 gnd.t254 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X116 vdd.t35 CSoutput.t192 output.t12 gnd.t54 sky130_fd_pr__nfet_01v8 ad=0.825 pd=5.33 as=0.825 ps=5.33 w=5 l=1
X117 a_n2903_n3924.t0 minus.t12 a_n2650_13878.t0 gnd.t0 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=1.155 ps=7.33 w=7 l=0.5
X118 vdd.t123 vdd.t121 vdd.t122 vdd.t108 sky130_fd_pr__pfet_01v8 ad=3.51 pd=18.78 as=0 ps=0 w=9 l=0.5
X119 CSoutput.t154 commonsourceibias.t80 gnd.t283 gnd.t259 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X120 CSoutput.t171 a_n8964_8799.t78 vdd.t257 vdd.t160 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X121 vdd.t120 vdd.t117 vdd.t119 vdd.t118 sky130_fd_pr__pfet_01v8 ad=3.51 pd=18.78 as=0 ps=0 w=9 l=0.5
X122 gnd.t282 commonsourceibias.t81 CSoutput.t153 gnd.t257 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=1.155 ps=7.33 w=7 l=1
X123 commonsourceibias.t51 commonsourceibias.t50 gnd.t281 gnd.t214 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X124 CSoutput.t152 commonsourceibias.t82 gnd.t280 gnd.t279 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X125 CSoutput.t32 a_n8964_8799.t79 vdd.t256 vdd.t133 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X126 CSoutput.t193 a_n2650_8322.t30 sky130_fd_pr__cap_mim_m3_1 l=12 w=12
X127 vdd.t255 a_n8964_8799.t80 CSoutput.t11 vdd.t252 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X128 vdd.t295 a_n2650_13878.t72 a_n2650_8322.t7 vdd.t294 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X129 a_n2650_13878.t29 a_n2650_13878.t28 a_n2472_13878.t12 vdd.t17 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X130 vdd.t116 vdd.t114 vdd.t115 vdd.t84 sky130_fd_pr__pfet_01v8 ad=3.12 pd=16.78 as=0 ps=0 w=8 l=0.5
X131 a_n2650_8322.t6 a_n2650_13878.t73 vdd.t297 vdd.t296 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X132 a_n2903_n3924.t34 diffpairibias.t18 gnd.t17 gnd.t16 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=2.73 ps=14.78 w=7 l=1
X133 CSoutput.t56 a_n8964_8799.t81 vdd.t254 vdd.t202 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X134 output.t18 outputibias.t11 gnd.t70 gnd.t69 sky130_fd_pr__nfet_01v8 ad=2.34 pd=12.78 as=2.34 ps=12.78 w=6 l=2
X135 a_n2650_13878.t53 minus.t13 a_n2903_n3924.t40 gnd.t10 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.5
X136 gnd.t278 commonsourceibias.t83 CSoutput.t113 gnd.t234 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X137 CSoutput.t194 a_n2650_8322.t29 sky130_fd_pr__cap_mim_m3_1 l=12 w=12
X138 commonsourceibias.t17 commonsourceibias.t16 gnd.t277 gnd.t259 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X139 a_n2903_n3924.t27 plus.t11 a_n8964_8799.t12 gnd.t27 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.5
X140 vdd.t1 a_n2650_13878.t74 a_n2472_13878.t26 vdd.t0 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X141 gnd.t155 gnd.t153 minus.t3 gnd.t154 sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.39 ps=2.78 w=1 l=0.5
X142 vdd.t113 vdd.t111 vdd.t112 vdd.t100 sky130_fd_pr__pfet_01v8 ad=3.12 pd=16.78 as=0 ps=0 w=8 l=0.5
X143 vdd.t110 vdd.t107 vdd.t109 vdd.t108 sky130_fd_pr__pfet_01v8 ad=3.51 pd=18.78 as=0 ps=0 w=9 l=0.5
X144 vdd.t253 a_n8964_8799.t82 CSoutput.t94 vdd.t252 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X145 vdd.t251 a_n8964_8799.t83 CSoutput.t30 vdd.t224 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X146 gnd.t276 commonsourceibias.t84 CSoutput.t112 gnd.t183 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X147 gnd.t275 commonsourceibias.t14 commonsourceibias.t15 gnd.t274 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X148 a_n8964_8799.t11 plus.t12 a_n2903_n3924.t26 gnd.t21 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=2.73 ps=14.78 w=7 l=0.5
X149 vdd.t106 vdd.t103 vdd.t105 vdd.t104 sky130_fd_pr__pfet_01v8 ad=3.51 pd=18.78 as=0 ps=0 w=9 l=0.5
X150 a_n2650_8322.t5 a_n2650_13878.t75 vdd.t3 vdd.t2 sky130_fd_pr__pfet_01v8 ad=3.51 pd=18.78 as=1.485 ps=9.33 w=9 l=0.5
X151 commonsourceibias.t13 commonsourceibias.t12 gnd.t273 gnd.t222 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X152 gnd.t272 commonsourceibias.t85 CSoutput.t111 gnd.t225 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X153 a_n2650_13878.t63 minus.t14 a_n2903_n3924.t55 gnd.t14 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.5
X154 gnd.t271 commonsourceibias.t86 CSoutput.t110 gnd.t270 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X155 a_n8964_8799.t6 a_n2650_13878.t76 a_n2650_8322.t20 vdd.t8 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X156 CSoutput.t165 a_n8964_8799.t84 vdd.t250 vdd.t168 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X157 diffpairibias.t11 diffpairibias.t10 gnd.t322 gnd.t321 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=2.73 ps=14.78 w=7 l=1
X158 vdd.t249 a_n8964_8799.t85 CSoutput.t61 vdd.t248 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X159 a_n2650_13878.t41 a_n2650_13878.t40 a_n2472_13878.t11 vdd.t42 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X160 vdd.t247 a_n8964_8799.t86 CSoutput.t175 vdd.t158 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X161 a_n8964_8799.t7 a_n2650_13878.t77 a_n2650_8322.t19 vdd.t9 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X162 CSoutput.t83 a_n8964_8799.t87 vdd.t246 vdd.t245 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X163 CSoutput.t177 a_n8964_8799.t88 vdd.t244 vdd.t196 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X164 CSoutput.t179 a_n8964_8799.t89 vdd.t243 vdd.t211 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X165 gnd.t152 gnd.t149 gnd.t151 gnd.t150 sky130_fd_pr__nfet_01v8 ad=2.34 pd=12.78 as=0 ps=0 w=6 l=2
X166 gnd.t269 commonsourceibias.t87 CSoutput.t109 gnd.t243 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X167 a_n2472_13878.t10 a_n2650_13878.t22 a_n2650_13878.t23 vdd.t5 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X168 gnd.t268 commonsourceibias.t88 CSoutput.t108 gnd.t267 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X169 CSoutput.t107 commonsourceibias.t89 gnd.t266 gnd.t264 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=2.73 ps=14.78 w=7 l=1
X170 commonsourceibias.t11 commonsourceibias.t10 gnd.t265 gnd.t264 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=2.73 ps=14.78 w=7 l=1
X171 a_n8964_8799.t31 plus.t13 a_n2903_n3924.t25 gnd.t8 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.5
X172 vdd.t102 vdd.t99 vdd.t101 vdd.t100 sky130_fd_pr__pfet_01v8 ad=3.12 pd=16.78 as=0 ps=0 w=8 l=0.5
X173 a_n2903_n3924.t52 minus.t15 a_n2650_13878.t60 gnd.t182 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.5
X174 vdd.t98 vdd.t96 vdd.t97 vdd.t70 sky130_fd_pr__pfet_01v8 ad=3.12 pd=16.78 as=0 ps=0 w=8 l=0.5
X175 a_n2903_n3924.t2 minus.t16 a_n2650_13878.t2 gnd.t2 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=1.155 ps=7.33 w=7 l=0.5
X176 CSoutput.t57 a_n8964_8799.t90 vdd.t242 vdd.t230 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X177 a_n2650_13878.t4 minus.t17 a_n2903_n3924.t5 gnd.t6 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.5
X178 vdd.t38 a_n2650_13878.t78 a_n2650_8322.t4 vdd.t37 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=3.51 ps=18.78 w=9 l=0.5
X179 a_n2472_13878.t9 a_n2650_13878.t18 a_n2650_13878.t19 vdd.t56 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X180 CSoutput.t138 commonsourceibias.t90 gnd.t263 gnd.t206 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X181 vdd.t241 a_n8964_8799.t91 CSoutput.t69 vdd.t228 sky130_fd_pr__pfet_01v8 ad=3.12 pd=16.78 as=1.32 ps=8.33 w=8 l=0.5
X182 vdd.t240 a_n8964_8799.t92 CSoutput.t182 vdd.t226 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X183 vdd.t95 vdd.t93 vdd.t94 vdd.t84 sky130_fd_pr__pfet_01v8 ad=3.12 pd=16.78 as=0 ps=0 w=8 l=0.5
X184 a_n2650_13878.t25 a_n2650_13878.t24 a_n2472_13878.t8 vdd.t7 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X185 vdd.t239 a_n8964_8799.t93 CSoutput.t19 vdd.t170 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X186 CSoutput.t137 commonsourceibias.t91 gnd.t262 gnd.t254 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X187 a_n2903_n3924.t45 diffpairibias.t19 gnd.t63 gnd.t62 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=2.73 ps=14.78 w=7 l=1
X188 gnd.t148 gnd.t145 gnd.t147 gnd.t146 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=0 ps=0 w=7 l=1
X189 a_n2903_n3924.t44 diffpairibias.t20 gnd.t61 gnd.t60 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=2.73 ps=14.78 w=7 l=1
X190 a_n2650_13878.t62 minus.t18 a_n2903_n3924.t54 gnd.t68 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.5
X191 vdd.t26 CSoutput.t195 output.t11 gnd.t53 sky130_fd_pr__nfet_01v8 ad=0.825 pd=5.33 as=0.825 ps=5.33 w=5 l=1
X192 vdd.t238 a_n8964_8799.t94 CSoutput.t3 vdd.t228 sky130_fd_pr__pfet_01v8 ad=3.12 pd=16.78 as=1.32 ps=8.33 w=8 l=0.5
X193 CSoutput.t136 commonsourceibias.t92 gnd.t261 gnd.t189 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X194 CSoutput.t135 commonsourceibias.t93 gnd.t260 gnd.t259 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X195 vdd.t237 a_n8964_8799.t95 CSoutput.t84 vdd.t217 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X196 CSoutput.t79 a_n8964_8799.t96 vdd.t236 vdd.t151 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=3.12 ps=16.78 w=8 l=0.5
X197 gnd.t258 commonsourceibias.t94 CSoutput.t134 gnd.t257 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=1.155 ps=7.33 w=7 l=1
X198 gnd.t256 commonsourceibias.t95 CSoutput.t133 gnd.t236 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=1.155 ps=7.33 w=7 l=1
X199 gnd.t144 gnd.t142 minus.t2 gnd.t143 sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.5
X200 commonsourceibias.t29 commonsourceibias.t28 gnd.t255 gnd.t254 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X201 CSoutput.t132 commonsourceibias.t96 gnd.t253 gnd.t212 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X202 a_n2472_13878.t7 a_n2650_13878.t12 a_n2650_13878.t13 vdd.t10 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X203 vdd.t92 vdd.t90 vdd.t91 vdd.t62 sky130_fd_pr__pfet_01v8 ad=3.51 pd=18.78 as=0 ps=0 w=9 l=0.5
X204 a_n2650_8322.t18 a_n2650_13878.t79 a_n8964_8799.t25 vdd.t6 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X205 CSoutput.t172 a_n8964_8799.t97 vdd.t235 vdd.t211 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X206 CSoutput.t183 a_n8964_8799.t98 vdd.t234 vdd.t135 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X207 gnd.t252 commonsourceibias.t97 CSoutput.t131 gnd.t234 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X208 CSoutput.t55 a_n8964_8799.t99 vdd.t233 vdd.t232 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=3.12 ps=16.78 w=8 l=0.5
X209 a_n2650_13878.t7 minus.t19 a_n2903_n3924.t8 gnd.t9 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.5
X210 gnd.t141 gnd.t139 gnd.t140 gnd.t97 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=0 ps=0 w=7 l=1
X211 CSoutput.t130 commonsourceibias.t98 gnd.t251 gnd.t230 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X212 diffpairibias.t9 diffpairibias.t8 gnd.t42 gnd.t41 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=2.73 ps=14.78 w=7 l=1
X213 a_n2472_13878.t25 a_n2650_13878.t80 vdd.t52 vdd.t51 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X214 vdd.t54 a_n2650_13878.t81 a_n2472_13878.t24 vdd.t53 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X215 CSoutput.t85 a_n8964_8799.t100 vdd.t231 vdd.t230 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X216 a_n2903_n3924.t24 plus.t14 a_n8964_8799.t16 gnd.t1 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.5
X217 vdd.t229 a_n8964_8799.t101 CSoutput.t67 vdd.t228 sky130_fd_pr__pfet_01v8 ad=3.12 pd=16.78 as=1.32 ps=8.33 w=8 l=0.5
X218 vdd.t227 a_n8964_8799.t102 CSoutput.t37 vdd.t226 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X219 vdd.t225 a_n8964_8799.t103 CSoutput.t60 vdd.t224 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X220 gnd.t250 commonsourceibias.t99 CSoutput.t122 gnd.t228 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X221 CSoutput.t121 commonsourceibias.t100 gnd.t249 gnd.t187 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=2.73 ps=14.78 w=7 l=1
X222 CSoutput.t68 a_n8964_8799.t104 vdd.t223 vdd.t190 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X223 a_n2903_n3924.t38 minus.t20 a_n2650_13878.t51 gnd.t31 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.5
X224 a_n2472_13878.t6 a_n2650_13878.t36 a_n2650_13878.t37 vdd.t4 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X225 gnd.t248 commonsourceibias.t22 commonsourceibias.t23 gnd.t204 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X226 a_n2903_n3924.t23 plus.t15 a_n8964_8799.t32 gnd.t33 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.5
X227 gnd.t247 commonsourceibias.t101 CSoutput.t120 gnd.t225 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X228 a_n2903_n3924.t36 minus.t21 a_n2650_13878.t49 gnd.t20 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.5
X229 a_n8964_8799.t13 plus.t16 a_n2903_n3924.t22 gnd.t32 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.5
X230 vdd.t222 a_n8964_8799.t105 CSoutput.t176 vdd.t170 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X231 gnd.t245 commonsourceibias.t102 CSoutput.t118 gnd.t243 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X232 a_n2650_8322.t17 a_n2650_13878.t82 a_n8964_8799.t29 vdd.t19 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X233 vdd.t31 CSoutput.t196 output.t10 gnd.t52 sky130_fd_pr__nfet_01v8 ad=0.825 pd=5.33 as=0.825 ps=5.33 w=5 l=1
X234 CSoutput.t70 a_n8964_8799.t106 vdd.t221 vdd.t173 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X235 diffpairibias.t7 diffpairibias.t6 gnd.t67 gnd.t66 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=2.73 ps=14.78 w=7 l=1
X236 CSoutput.t119 commonsourceibias.t103 gnd.t246 gnd.t222 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X237 vdd.t220 a_n8964_8799.t107 CSoutput.t178 vdd.t219 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X238 a_n2472_13878.t5 a_n2650_13878.t20 a_n2650_13878.t21 vdd.t55 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=3.51 ps=18.78 w=9 l=0.5
X239 vdd.t44 a_n2650_13878.t83 a_n2650_8322.t3 vdd.t43 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=3.51 ps=18.78 w=9 l=0.5
X240 gnd.t244 commonsourceibias.t20 commonsourceibias.t21 gnd.t243 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X241 gnd.t138 gnd.t135 gnd.t137 gnd.t136 sky130_fd_pr__nfet_01v8 ad=1.95 pd=10.78 as=0 ps=0 w=5 l=1
X242 vdd.t218 a_n8964_8799.t108 CSoutput.t44 vdd.t217 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X243 gnd.t134 gnd.t132 gnd.t133 gnd.t97 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=0 ps=0 w=7 l=1
X244 CSoutput.t117 commonsourceibias.t104 gnd.t242 gnd.t218 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X245 CSoutput.t116 commonsourceibias.t105 gnd.t241 gnd.t206 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X246 CSoutput.t20 a_n8964_8799.t109 vdd.t216 vdd.t198 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X247 a_n2472_13878.t23 a_n2650_13878.t84 vdd.t48 vdd.t47 sky130_fd_pr__pfet_01v8 ad=3.51 pd=18.78 as=1.485 ps=9.33 w=9 l=0.5
X248 vdd.t89 vdd.t87 vdd.t88 vdd.t70 sky130_fd_pr__pfet_01v8 ad=3.12 pd=16.78 as=0 ps=0 w=8 l=0.5
X249 plus.t1 gnd.t129 gnd.t131 gnd.t130 sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.5
X250 vdd.t215 a_n8964_8799.t110 CSoutput.t180 vdd.t214 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X251 vdd.t213 a_n8964_8799.t111 CSoutput.t78 vdd.t192 sky130_fd_pr__pfet_01v8 ad=3.12 pd=16.78 as=1.32 ps=8.33 w=8 l=0.5
X252 CSoutput.t80 a_n8964_8799.t112 vdd.t212 vdd.t211 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X253 CSoutput.t95 a_n8964_8799.t113 vdd.t210 vdd.t190 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X254 gnd.t128 gnd.t125 gnd.t127 gnd.t126 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=0 ps=0 w=7 l=0.5
X255 gnd.t240 commonsourceibias.t18 commonsourceibias.t19 gnd.t209 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X256 gnd.t124 gnd.t122 minus.t1 gnd.t123 sky130_fd_pr__nfet_01v8 ad=0.39 pd=2.78 as=0.165 ps=1.33 w=1 l=0.5
X257 gnd.t121 gnd.t118 gnd.t120 gnd.t119 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=0 ps=0 w=7 l=0.5
X258 gnd.t117 gnd.t114 gnd.t116 gnd.t115 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=0 ps=0 w=7 l=1
X259 vdd.t209 a_n8964_8799.t114 CSoutput.t96 vdd.t186 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X260 a_n2903_n3924.t49 diffpairibias.t21 gnd.t74 gnd.t73 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=2.73 ps=14.78 w=7 l=1
X261 gnd.t113 gnd.t110 gnd.t112 gnd.t111 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=0 ps=0 w=7 l=1
X262 CSoutput.t115 commonsourceibias.t106 gnd.t239 gnd.t214 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X263 vdd.t50 a_n2650_13878.t85 a_n2650_8322.t2 vdd.t49 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X264 a_n2650_8322.t16 a_n2650_13878.t86 a_n8964_8799.t27 vdd.t42 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X265 CSoutput.t87 a_n8964_8799.t115 vdd.t208 vdd.t155 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X266 CSoutput.t114 commonsourceibias.t107 gnd.t238 gnd.t189 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X267 vdd.t86 vdd.t83 vdd.t85 vdd.t84 sky130_fd_pr__pfet_01v8 ad=3.12 pd=16.78 as=0 ps=0 w=8 l=0.5
X268 vdd.t207 a_n8964_8799.t116 CSoutput.t98 vdd.t181 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X269 vdd.t82 vdd.t80 vdd.t81 vdd.t58 sky130_fd_pr__pfet_01v8 ad=3.12 pd=16.78 as=0 ps=0 w=8 l=0.5
X270 vdd.t206 a_n8964_8799.t117 CSoutput.t33 vdd.t179 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X271 gnd.t237 commonsourceibias.t108 CSoutput.t145 gnd.t236 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=1.155 ps=7.33 w=7 l=1
X272 vdd.t205 a_n8964_8799.t118 CSoutput.t38 vdd.t145 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X273 gnd.t235 commonsourceibias.t32 commonsourceibias.t33 gnd.t234 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X274 gnd.t109 gnd.t106 gnd.t108 gnd.t107 sky130_fd_pr__nfet_01v8 ad=2.34 pd=12.78 as=0 ps=0 w=6 l=2
X275 CSoutput.t144 commonsourceibias.t109 gnd.t233 gnd.t212 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X276 output.t9 CSoutput.t197 vdd.t29 gnd.t51 sky130_fd_pr__nfet_01v8 ad=0.825 pd=5.33 as=0.825 ps=5.33 w=5 l=1
X277 gnd.t232 commonsourceibias.t110 CSoutput.t143 gnd.t209 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X278 a_n2903_n3924.t21 plus.t17 a_n8964_8799.t19 gnd.t3 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.5
X279 vdd.t79 vdd.t76 vdd.t78 vdd.t77 sky130_fd_pr__pfet_01v8 ad=3.51 pd=18.78 as=0 ps=0 w=9 l=0.5
X280 gnd.t105 gnd.t103 gnd.t104 gnd.t86 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=0 ps=0 w=7 l=1
X281 vdd.t204 a_n8964_8799.t119 CSoutput.t89 vdd.t139 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X282 a_n8964_8799.t5 plus.t18 a_n2903_n3924.t20 gnd.t15 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.5
X283 CSoutput.t50 a_n8964_8799.t120 vdd.t203 vdd.t202 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X284 outputibias.t7 outputibias.t6 gnd.t320 gnd.t319 sky130_fd_pr__nfet_01v8 ad=2.34 pd=12.78 as=2.34 ps=12.78 w=6 l=2
X285 a_n2903_n3924.t6 minus.t22 a_n2650_13878.t5 gnd.t7 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.5
X286 a_n2472_13878.t4 a_n2650_13878.t16 a_n2650_13878.t17 vdd.t45 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X287 CSoutput.t48 a_n8964_8799.t121 vdd.t201 vdd.t175 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X288 CSoutput.t168 a_n8964_8799.t122 vdd.t200 vdd.t173 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X289 gnd.t102 gnd.t100 gnd.t101 gnd.t86 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=0 ps=0 w=7 l=1
X290 CSoutput.t142 commonsourceibias.t111 gnd.t231 gnd.t230 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X291 a_n2650_8322.t15 a_n2650_13878.t87 a_n8964_8799.t28 vdd.t39 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X292 vdd.t75 vdd.t73 vdd.t74 vdd.t58 sky130_fd_pr__pfet_01v8 ad=3.12 pd=16.78 as=0 ps=0 w=8 l=0.5
X293 diffpairibias.t5 diffpairibias.t4 gnd.t25 gnd.t24 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=2.73 ps=14.78 w=7 l=1
X294 a_n2903_n3924.t50 minus.t23 a_n2650_13878.t58 gnd.t38 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.5
X295 a_n8964_8799.t22 plus.t19 a_n2903_n3924.t19 gnd.t43 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.5
X296 outputibias.t5 outputibias.t4 gnd.t23 gnd.t22 sky130_fd_pr__nfet_01v8 ad=2.34 pd=12.78 as=2.34 ps=12.78 w=6 l=2
X297 CSoutput.t31 a_n8964_8799.t123 vdd.t199 vdd.t198 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X298 CSoutput.t28 a_n8964_8799.t124 vdd.t197 vdd.t196 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X299 CSoutput.t163 a_n8964_8799.t125 vdd.t195 vdd.t168 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X300 vdd.t194 a_n8964_8799.t126 CSoutput.t16 vdd.t179 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X301 gnd.t229 commonsourceibias.t112 CSoutput.t141 gnd.t228 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X302 vdd.t72 vdd.t69 vdd.t71 vdd.t70 sky130_fd_pr__pfet_01v8 ad=3.12 pd=16.78 as=0 ps=0 w=8 l=0.5
X303 CSoutput.t140 commonsourceibias.t113 gnd.t227 gnd.t187 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=2.73 ps=14.78 w=7 l=1
X304 vdd.t193 a_n8964_8799.t127 CSoutput.t27 vdd.t192 sky130_fd_pr__pfet_01v8 ad=3.12 pd=16.78 as=1.32 ps=8.33 w=8 l=0.5
X305 outputibias.t3 outputibias.t2 gnd.t29 gnd.t28 sky130_fd_pr__nfet_01v8 ad=2.34 pd=12.78 as=2.34 ps=12.78 w=6 l=2
X306 output.t8 CSoutput.t198 vdd.t21 gnd.t50 sky130_fd_pr__nfet_01v8 ad=0.825 pd=5.33 as=0.825 ps=5.33 w=5 l=1
X307 a_n2650_8322.t1 a_n2650_13878.t88 vdd.t301 vdd.t300 sky130_fd_pr__pfet_01v8 ad=3.51 pd=18.78 as=1.485 ps=9.33 w=9 l=0.5
X308 gnd.t226 commonsourceibias.t30 commonsourceibias.t31 gnd.t225 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X309 outputibias.t1 outputibias.t0 gnd.t318 gnd.t317 sky130_fd_pr__nfet_01v8 ad=2.34 pd=12.78 as=2.34 ps=12.78 w=6 l=2
X310 gnd.t224 commonsourceibias.t114 CSoutput.t139 gnd.t204 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X311 CSoutput.t13 a_n8964_8799.t128 vdd.t191 vdd.t190 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X312 a_n2903_n3924.t18 plus.t20 a_n8964_8799.t15 gnd.t30 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.5
X313 vdd.t189 a_n8964_8799.t129 CSoutput.t51 vdd.t186 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X314 CSoutput.t24 a_n8964_8799.t130 vdd.t188 vdd.t149 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X315 CSoutput.t129 commonsourceibias.t115 gnd.t223 gnd.t222 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X316 vdd.t303 a_n2650_13878.t89 a_n2472_13878.t22 vdd.t302 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=3.51 ps=18.78 w=9 l=0.5
X317 vdd.t187 a_n8964_8799.t131 CSoutput.t82 vdd.t186 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X318 CSoutput.t23 a_n8964_8799.t132 vdd.t185 vdd.t184 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X319 output.t7 CSoutput.t199 vdd.t27 gnd.t49 sky130_fd_pr__nfet_01v8 ad=0.825 pd=5.33 as=0.825 ps=5.33 w=5 l=1
X320 CSoutput.t88 a_n8964_8799.t133 vdd.t183 vdd.t155 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X321 gnd.t99 gnd.t96 gnd.t98 gnd.t97 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=0 ps=0 w=7 l=1
X322 vdd.t30 CSoutput.t200 output.t6 gnd.t48 sky130_fd_pr__nfet_01v8 ad=0.825 pd=5.33 as=0.825 ps=5.33 w=5 l=1
X323 gnd.t221 commonsourceibias.t116 CSoutput.t128 gnd.t195 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X324 vdd.t182 a_n8964_8799.t134 CSoutput.t8 vdd.t181 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X325 CSoutput.t127 commonsourceibias.t117 gnd.t220 gnd.t199 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X326 CSoutput.t126 commonsourceibias.t118 gnd.t219 gnd.t218 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X327 vdd.t180 a_n8964_8799.t135 CSoutput.t173 vdd.t179 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X328 gnd.t217 commonsourceibias.t26 commonsourceibias.t27 gnd.t216 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X329 a_n8964_8799.t39 plus.t21 a_n2903_n3924.t17 gnd.t26 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=2.73 ps=14.78 w=7 l=0.5
X330 vdd.t178 a_n8964_8799.t136 CSoutput.t0 vdd.t145 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X331 a_n2903_n3924.t43 minus.t24 a_n2650_13878.t56 gnd.t27 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.5
X332 a_n2650_8322.t14 a_n2650_13878.t90 a_n8964_8799.t34 vdd.t46 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X333 a_n8964_8799.t35 a_n2650_13878.t91 a_n2650_8322.t13 vdd.t45 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X334 a_n2472_13878.t21 a_n2650_13878.t92 vdd.t299 vdd.t298 sky130_fd_pr__pfet_01v8 ad=3.51 pd=18.78 as=1.485 ps=9.33 w=9 l=0.5
X335 vdd.t68 vdd.t65 vdd.t67 vdd.t66 sky130_fd_pr__pfet_01v8 ad=3.51 pd=18.78 as=0 ps=0 w=9 l=0.5
X336 vdd.t177 a_n8964_8799.t137 CSoutput.t4 vdd.t153 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X337 vdd.t64 vdd.t61 vdd.t63 vdd.t62 sky130_fd_pr__pfet_01v8 ad=3.51 pd=18.78 as=0 ps=0 w=9 l=0.5
X338 CSoutput.t76 a_n8964_8799.t138 vdd.t176 vdd.t175 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X339 CSoutput.t75 a_n8964_8799.t139 vdd.t174 vdd.t173 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X340 CSoutput.t26 a_n8964_8799.t140 vdd.t172 vdd.t151 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=3.12 ps=16.78 w=8 l=0.5
X341 vdd.t60 vdd.t57 vdd.t59 vdd.t58 sky130_fd_pr__pfet_01v8 ad=3.12 pd=16.78 as=0 ps=0 w=8 l=0.5
X342 a_n8964_8799.t3 plus.t22 a_n2903_n3924.t16 gnd.t14 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.5
X343 a_n8964_8799.t42 a_n2650_13878.t93 a_n2650_8322.t12 vdd.t10 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X344 CSoutput.t125 commonsourceibias.t119 gnd.t215 gnd.t214 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X345 a_n2650_8322.t11 a_n2650_13878.t94 a_n8964_8799.t23 vdd.t17 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X346 a_n2650_13878.t52 minus.t25 a_n2903_n3924.t39 gnd.t13 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.5
X347 vdd.t171 a_n8964_8799.t141 CSoutput.t90 vdd.t170 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X348 CSoutput.t22 a_n8964_8799.t142 vdd.t169 vdd.t168 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X349 CSoutput.t181 a_n8964_8799.t143 vdd.t167 vdd.t147 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X350 CSoutput.t92 a_n8964_8799.t144 vdd.t166 vdd.t147 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X351 output.t5 CSoutput.t201 vdd.t28 gnd.t47 sky130_fd_pr__nfet_01v8 ad=0.825 pd=5.33 as=0.825 ps=5.33 w=5 l=1
X352 a_n2472_13878.t3 a_n2650_13878.t46 a_n2650_13878.t47 vdd.t8 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X353 commonsourceibias.t25 commonsourceibias.t24 gnd.t213 gnd.t212 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X354 gnd.t211 commonsourceibias.t120 CSoutput.t124 gnd.t191 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X355 vdd.t165 a_n8964_8799.t145 CSoutput.t25 vdd.t143 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X356 gnd.t95 gnd.t92 gnd.t94 gnd.t93 sky130_fd_pr__nfet_01v8 ad=1.95 pd=10.78 as=0 ps=0 w=5 l=1
X357 gnd.t210 commonsourceibias.t121 CSoutput.t123 gnd.t209 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X358 a_n2903_n3924.t15 plus.t23 a_n8964_8799.t2 gnd.t2 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=1.155 ps=7.33 w=7 l=0.5
X359 a_n8964_8799.t10 plus.t24 a_n2903_n3924.t14 gnd.t6 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.5
X360 output.t4 CSoutput.t202 vdd.t25 gnd.t46 sky130_fd_pr__nfet_01v8 ad=0.825 pd=5.33 as=0.825 ps=5.33 w=5 l=1
X361 gnd.t91 gnd.t89 gnd.t90 gnd.t79 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=0 ps=0 w=7 l=1
X362 a_n2903_n3924.t46 diffpairibias.t22 gnd.t65 gnd.t64 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=2.73 ps=14.78 w=7 l=1
X363 vdd.t164 a_n8964_8799.t146 CSoutput.t39 vdd.t139 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X364 gnd.t88 gnd.t85 gnd.t87 gnd.t86 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=0 ps=0 w=7 l=1
X365 gnd.t186 commonsourceibias.t122 CSoutput.t150 gnd.t185 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X366 CSoutput.t53 a_n8964_8799.t147 vdd.t163 vdd.t135 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X367 a_n2650_13878.t39 a_n2650_13878.t38 a_n2472_13878.t2 vdd.t46 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X368 commonsourceibias.t41 commonsourceibias.t40 gnd.t208 gnd.t199 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X369 a_n8964_8799.t24 a_n2650_13878.t95 a_n2650_8322.t10 vdd.t20 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X370 vdd.t162 a_n8964_8799.t148 CSoutput.t47 vdd.t143 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X371 CSoutput.t86 a_n8964_8799.t149 vdd.t161 vdd.t160 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X372 a_n2903_n3924.t13 plus.t25 a_n8964_8799.t14 gnd.t0 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=1.155 ps=7.33 w=7 l=0.5
X373 diffpairibias.t3 diffpairibias.t2 gnd.t19 gnd.t18 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=2.73 ps=14.78 w=7 l=1
X374 vdd.t159 a_n8964_8799.t150 CSoutput.t170 vdd.t158 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X375 CSoutput.t14 a_n8964_8799.t151 vdd.t157 vdd.t133 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X376 CSoutput.t203 a_n2650_8322.t28 sky130_fd_pr__cap_mim_m3_1 l=12 w=12
X377 CSoutput.t81 a_n8964_8799.t152 vdd.t156 vdd.t155 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X378 a_n2650_8322.t9 a_n2650_13878.t96 a_n8964_8799.t26 vdd.t7 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X379 commonsourceibias.t39 commonsourceibias.t38 gnd.t207 gnd.t206 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X380 vdd.t154 a_n8964_8799.t153 CSoutput.t34 vdd.t153 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X381 gnd.t205 commonsourceibias.t123 CSoutput.t149 gnd.t204 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X382 CSoutput.t66 a_n8964_8799.t154 vdd.t152 vdd.t151 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=3.12 ps=16.78 w=8 l=0.5
X383 CSoutput.t59 a_n8964_8799.t155 vdd.t150 vdd.t149 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X384 gnd.t81 gnd.t78 gnd.t80 gnd.t79 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=0 ps=0 w=7 l=1
X385 diffpairibias.t1 diffpairibias.t0 gnd.t314 gnd.t313 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=2.73 ps=14.78 w=7 l=1
X386 gnd.t84 gnd.t82 plus.t0 gnd.t83 sky130_fd_pr__nfet_01v8 ad=0.39 pd=2.78 as=0.165 ps=1.33 w=1 l=0.5
X387 a_n8964_8799.t0 plus.t26 a_n2903_n3924.t12 gnd.t10 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.5
X388 vdd.t32 CSoutput.t204 output.t3 gnd.t45 sky130_fd_pr__nfet_01v8 ad=0.825 pd=5.33 as=0.825 ps=5.33 w=5 l=1
X389 CSoutput.t148 commonsourceibias.t124 gnd.t203 gnd.t202 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X390 minus.t0 gnd.t75 gnd.t77 gnd.t76 sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.5
X391 vdd.t41 a_n2650_13878.t97 a_n2472_13878.t20 vdd.t40 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=3.51 ps=18.78 w=9 l=0.5
X392 CSoutput.t73 a_n8964_8799.t156 vdd.t148 vdd.t147 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X393 gnd.t201 commonsourceibias.t125 CSoutput.t147 gnd.t195 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X394 CSoutput.t146 commonsourceibias.t126 gnd.t200 gnd.t199 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X395 vdd.t146 a_n8964_8799.t157 CSoutput.t15 vdd.t145 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X396 commonsourceibias.t37 commonsourceibias.t36 gnd.t198 gnd.t197 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X397 vdd.t144 a_n8964_8799.t158 CSoutput.t41 vdd.t143 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X398 CSoutput.t77 a_n8964_8799.t159 vdd.t142 vdd.t141 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X399 gnd.t196 commonsourceibias.t34 commonsourceibias.t35 gnd.t195 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X400 vdd.t23 CSoutput.t205 output.t2 gnd.t44 sky130_fd_pr__nfet_01v8 ad=0.825 pd=5.33 as=0.825 ps=5.33 w=5 l=1
X401 a_n2650_13878.t59 minus.t26 a_n2903_n3924.t51 gnd.t21 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=2.73 ps=14.78 w=7 l=0.5
X402 CSoutput.t151 commonsourceibias.t127 gnd.t194 gnd.t193 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X403 a_n2650_8322.t8 a_n2650_13878.t98 a_n8964_8799.t8 vdd.t11 sky130_fd_pr__pfet_01v8 ad=3.51 pd=18.78 as=1.485 ps=9.33 w=9 l=0.5
X404 gnd.t192 commonsourceibias.t48 commonsourceibias.t49 gnd.t191 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X405 vdd.t140 a_n8964_8799.t160 CSoutput.t18 vdd.t139 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X406 vdd.t138 a_n8964_8799.t161 CSoutput.t43 vdd.t137 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X407 CSoutput.t65 a_n8964_8799.t162 vdd.t136 vdd.t135 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X408 commonsourceibias.t47 commonsourceibias.t46 gnd.t190 gnd.t189 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X409 a_n2903_n3924.t11 plus.t27 a_n8964_8799.t9 gnd.t20 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.5
X410 a_n2650_8322.t0 a_n2650_13878.t99 vdd.t13 vdd.t12 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X411 a_n2650_13878.t61 minus.t27 a_n2903_n3924.t53 gnd.t32 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.5
X412 a_n2472_13878.t1 a_n2650_13878.t42 a_n2650_13878.t43 vdd.t293 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=3.51 ps=18.78 w=9 l=0.5
X413 commonsourceibias.t45 commonsourceibias.t44 gnd.t188 gnd.t187 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=2.73 ps=14.78 w=7 l=1
X414 a_n2903_n3924.t48 diffpairibias.t23 gnd.t72 gnd.t71 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=2.73 ps=14.78 w=7 l=1
X415 a_n2650_13878.t6 minus.t28 a_n2903_n3924.t7 gnd.t8 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.5
X416 CSoutput.t63 a_n8964_8799.t163 vdd.t134 vdd.t133 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X417 gnd.t184 commonsourceibias.t42 commonsourceibias.t43 gnd.t183 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X418 a_n2650_13878.t33 a_n2650_13878.t32 a_n2472_13878.t0 vdd.t19 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X419 a_n2903_n3924.t10 plus.t28 a_n8964_8799.t43 gnd.t182 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.5
R0 commonsourceibias.n35 commonsourceibias.t10 223.028
R1 commonsourceibias.n128 commonsourceibias.t89 223.028
R2 commonsourceibias.n217 commonsourceibias.t77 223.028
R3 commonsourceibias.n364 commonsourceibias.t4 223.028
R4 commonsourceibias.n305 commonsourceibias.t108 223.028
R5 commonsourceibias.n499 commonsourceibias.t95 223.028
R6 commonsourceibias.n99 commonsourceibias.t54 207.983
R7 commonsourceibias.n192 commonsourceibias.t94 207.983
R8 commonsourceibias.n281 commonsourceibias.t81 207.983
R9 commonsourceibias.n430 commonsourceibias.t44 207.983
R10 commonsourceibias.n476 commonsourceibias.t113 207.983
R11 commonsourceibias.n565 commonsourceibias.t100 207.983
R12 commonsourceibias.n97 commonsourceibias.t24 168.701
R13 commonsourceibias.n91 commonsourceibias.t14 168.701
R14 commonsourceibias.n17 commonsourceibias.t52 168.701
R15 commonsourceibias.n83 commonsourceibias.t20 168.701
R16 commonsourceibias.n77 commonsourceibias.t58 168.701
R17 commonsourceibias.n22 commonsourceibias.t60 168.701
R18 commonsourceibias.n69 commonsourceibias.t16 168.701
R19 commonsourceibias.n63 commonsourceibias.t56 168.701
R20 commonsourceibias.n25 commonsourceibias.t38 168.701
R21 commonsourceibias.n27 commonsourceibias.t6 168.701
R22 commonsourceibias.n29 commonsourceibias.t62 168.701
R23 commonsourceibias.n46 commonsourceibias.t32 168.701
R24 commonsourceibias.n40 commonsourceibias.t0 168.701
R25 commonsourceibias.n34 commonsourceibias.t26 168.701
R26 commonsourceibias.n190 commonsourceibias.t109 168.701
R27 commonsourceibias.n184 commonsourceibias.t72 168.701
R28 commonsourceibias.n5 commonsourceibias.t70 168.701
R29 commonsourceibias.n176 commonsourceibias.t102 168.701
R30 commonsourceibias.n170 commonsourceibias.t118 168.701
R31 commonsourceibias.n10 commonsourceibias.t66 168.701
R32 commonsourceibias.n162 commonsourceibias.t93 168.701
R33 commonsourceibias.n156 commonsourceibias.t88 168.701
R34 commonsourceibias.n118 commonsourceibias.t105 168.701
R35 commonsourceibias.n120 commonsourceibias.t86 168.701
R36 commonsourceibias.n122 commonsourceibias.t82 168.701
R37 commonsourceibias.n139 commonsourceibias.t97 168.701
R38 commonsourceibias.n133 commonsourceibias.t111 168.701
R39 commonsourceibias.n127 commonsourceibias.t75 168.701
R40 commonsourceibias.n216 commonsourceibias.t67 168.701
R41 commonsourceibias.n222 commonsourceibias.t98 168.701
R42 commonsourceibias.n228 commonsourceibias.t83 168.701
R43 commonsourceibias.n211 commonsourceibias.t71 168.701
R44 commonsourceibias.n209 commonsourceibias.t74 168.701
R45 commonsourceibias.n207 commonsourceibias.t90 168.701
R46 commonsourceibias.n245 commonsourceibias.t76 168.701
R47 commonsourceibias.n251 commonsourceibias.t80 168.701
R48 commonsourceibias.n204 commonsourceibias.t122 168.701
R49 commonsourceibias.n259 commonsourceibias.t104 168.701
R50 commonsourceibias.n265 commonsourceibias.t87 168.701
R51 commonsourceibias.n199 commonsourceibias.t127 168.701
R52 commonsourceibias.n273 commonsourceibias.t65 168.701
R53 commonsourceibias.n279 commonsourceibias.t96 168.701
R54 commonsourceibias.n363 commonsourceibias.t28 168.701
R55 commonsourceibias.n369 commonsourceibias.t34 168.701
R56 commonsourceibias.n375 commonsourceibias.t12 168.701
R57 commonsourceibias.n358 commonsourceibias.t30 168.701
R58 commonsourceibias.n356 commonsourceibias.t36 168.701
R59 commonsourceibias.n354 commonsourceibias.t18 168.701
R60 commonsourceibias.n392 commonsourceibias.t46 168.701
R61 commonsourceibias.n398 commonsourceibias.t8 168.701
R62 commonsourceibias.n400 commonsourceibias.t40 168.701
R63 commonsourceibias.n407 commonsourceibias.t48 168.701
R64 commonsourceibias.n413 commonsourceibias.t50 168.701
R65 commonsourceibias.n415 commonsourceibias.t42 168.701
R66 commonsourceibias.n422 commonsourceibias.t2 168.701
R67 commonsourceibias.n428 commonsourceibias.t22 168.701
R68 commonsourceibias.n474 commonsourceibias.t123 168.701
R69 commonsourceibias.n468 commonsourceibias.t68 168.701
R70 commonsourceibias.n461 commonsourceibias.t84 168.701
R71 commonsourceibias.n459 commonsourceibias.t119 168.701
R72 commonsourceibias.n453 commonsourceibias.t64 168.701
R73 commonsourceibias.n446 commonsourceibias.t126 168.701
R74 commonsourceibias.n444 commonsourceibias.t112 168.701
R75 commonsourceibias.n304 commonsourceibias.t91 168.701
R76 commonsourceibias.n310 commonsourceibias.t125 168.701
R77 commonsourceibias.n316 commonsourceibias.t115 168.701
R78 commonsourceibias.n299 commonsourceibias.t101 168.701
R79 commonsourceibias.n297 commonsourceibias.t78 168.701
R80 commonsourceibias.n295 commonsourceibias.t121 168.701
R81 commonsourceibias.n333 commonsourceibias.t107 168.701
R82 commonsourceibias.n498 commonsourceibias.t79 168.701
R83 commonsourceibias.n504 commonsourceibias.t116 168.701
R84 commonsourceibias.n510 commonsourceibias.t103 168.701
R85 commonsourceibias.n493 commonsourceibias.t85 168.701
R86 commonsourceibias.n491 commonsourceibias.t69 168.701
R87 commonsourceibias.n489 commonsourceibias.t110 168.701
R88 commonsourceibias.n527 commonsourceibias.t92 168.701
R89 commonsourceibias.n533 commonsourceibias.t99 168.701
R90 commonsourceibias.n535 commonsourceibias.t117 168.701
R91 commonsourceibias.n542 commonsourceibias.t120 168.701
R92 commonsourceibias.n548 commonsourceibias.t106 168.701
R93 commonsourceibias.n550 commonsourceibias.t73 168.701
R94 commonsourceibias.n557 commonsourceibias.t124 168.701
R95 commonsourceibias.n563 commonsourceibias.t114 168.701
R96 commonsourceibias.n36 commonsourceibias.n33 161.3
R97 commonsourceibias.n38 commonsourceibias.n37 161.3
R98 commonsourceibias.n39 commonsourceibias.n32 161.3
R99 commonsourceibias.n42 commonsourceibias.n41 161.3
R100 commonsourceibias.n43 commonsourceibias.n31 161.3
R101 commonsourceibias.n45 commonsourceibias.n44 161.3
R102 commonsourceibias.n47 commonsourceibias.n30 161.3
R103 commonsourceibias.n49 commonsourceibias.n48 161.3
R104 commonsourceibias.n51 commonsourceibias.n50 161.3
R105 commonsourceibias.n52 commonsourceibias.n28 161.3
R106 commonsourceibias.n54 commonsourceibias.n53 161.3
R107 commonsourceibias.n56 commonsourceibias.n55 161.3
R108 commonsourceibias.n57 commonsourceibias.n26 161.3
R109 commonsourceibias.n59 commonsourceibias.n58 161.3
R110 commonsourceibias.n61 commonsourceibias.n60 161.3
R111 commonsourceibias.n62 commonsourceibias.n24 161.3
R112 commonsourceibias.n65 commonsourceibias.n64 161.3
R113 commonsourceibias.n66 commonsourceibias.n23 161.3
R114 commonsourceibias.n68 commonsourceibias.n67 161.3
R115 commonsourceibias.n70 commonsourceibias.n21 161.3
R116 commonsourceibias.n72 commonsourceibias.n71 161.3
R117 commonsourceibias.n73 commonsourceibias.n20 161.3
R118 commonsourceibias.n75 commonsourceibias.n74 161.3
R119 commonsourceibias.n76 commonsourceibias.n19 161.3
R120 commonsourceibias.n79 commonsourceibias.n78 161.3
R121 commonsourceibias.n80 commonsourceibias.n18 161.3
R122 commonsourceibias.n82 commonsourceibias.n81 161.3
R123 commonsourceibias.n84 commonsourceibias.n16 161.3
R124 commonsourceibias.n86 commonsourceibias.n85 161.3
R125 commonsourceibias.n87 commonsourceibias.n15 161.3
R126 commonsourceibias.n89 commonsourceibias.n88 161.3
R127 commonsourceibias.n90 commonsourceibias.n14 161.3
R128 commonsourceibias.n93 commonsourceibias.n92 161.3
R129 commonsourceibias.n94 commonsourceibias.n13 161.3
R130 commonsourceibias.n96 commonsourceibias.n95 161.3
R131 commonsourceibias.n98 commonsourceibias.n12 161.3
R132 commonsourceibias.n129 commonsourceibias.n126 161.3
R133 commonsourceibias.n131 commonsourceibias.n130 161.3
R134 commonsourceibias.n132 commonsourceibias.n125 161.3
R135 commonsourceibias.n135 commonsourceibias.n134 161.3
R136 commonsourceibias.n136 commonsourceibias.n124 161.3
R137 commonsourceibias.n138 commonsourceibias.n137 161.3
R138 commonsourceibias.n140 commonsourceibias.n123 161.3
R139 commonsourceibias.n142 commonsourceibias.n141 161.3
R140 commonsourceibias.n144 commonsourceibias.n143 161.3
R141 commonsourceibias.n145 commonsourceibias.n121 161.3
R142 commonsourceibias.n147 commonsourceibias.n146 161.3
R143 commonsourceibias.n149 commonsourceibias.n148 161.3
R144 commonsourceibias.n150 commonsourceibias.n119 161.3
R145 commonsourceibias.n152 commonsourceibias.n151 161.3
R146 commonsourceibias.n154 commonsourceibias.n153 161.3
R147 commonsourceibias.n155 commonsourceibias.n117 161.3
R148 commonsourceibias.n158 commonsourceibias.n157 161.3
R149 commonsourceibias.n159 commonsourceibias.n11 161.3
R150 commonsourceibias.n161 commonsourceibias.n160 161.3
R151 commonsourceibias.n163 commonsourceibias.n9 161.3
R152 commonsourceibias.n165 commonsourceibias.n164 161.3
R153 commonsourceibias.n166 commonsourceibias.n8 161.3
R154 commonsourceibias.n168 commonsourceibias.n167 161.3
R155 commonsourceibias.n169 commonsourceibias.n7 161.3
R156 commonsourceibias.n172 commonsourceibias.n171 161.3
R157 commonsourceibias.n173 commonsourceibias.n6 161.3
R158 commonsourceibias.n175 commonsourceibias.n174 161.3
R159 commonsourceibias.n177 commonsourceibias.n4 161.3
R160 commonsourceibias.n179 commonsourceibias.n178 161.3
R161 commonsourceibias.n180 commonsourceibias.n3 161.3
R162 commonsourceibias.n182 commonsourceibias.n181 161.3
R163 commonsourceibias.n183 commonsourceibias.n2 161.3
R164 commonsourceibias.n186 commonsourceibias.n185 161.3
R165 commonsourceibias.n187 commonsourceibias.n1 161.3
R166 commonsourceibias.n189 commonsourceibias.n188 161.3
R167 commonsourceibias.n191 commonsourceibias.n0 161.3
R168 commonsourceibias.n280 commonsourceibias.n194 161.3
R169 commonsourceibias.n278 commonsourceibias.n277 161.3
R170 commonsourceibias.n276 commonsourceibias.n195 161.3
R171 commonsourceibias.n275 commonsourceibias.n274 161.3
R172 commonsourceibias.n272 commonsourceibias.n196 161.3
R173 commonsourceibias.n271 commonsourceibias.n270 161.3
R174 commonsourceibias.n269 commonsourceibias.n197 161.3
R175 commonsourceibias.n268 commonsourceibias.n267 161.3
R176 commonsourceibias.n266 commonsourceibias.n198 161.3
R177 commonsourceibias.n264 commonsourceibias.n263 161.3
R178 commonsourceibias.n262 commonsourceibias.n200 161.3
R179 commonsourceibias.n261 commonsourceibias.n260 161.3
R180 commonsourceibias.n258 commonsourceibias.n201 161.3
R181 commonsourceibias.n257 commonsourceibias.n256 161.3
R182 commonsourceibias.n255 commonsourceibias.n202 161.3
R183 commonsourceibias.n254 commonsourceibias.n253 161.3
R184 commonsourceibias.n252 commonsourceibias.n203 161.3
R185 commonsourceibias.n250 commonsourceibias.n249 161.3
R186 commonsourceibias.n248 commonsourceibias.n205 161.3
R187 commonsourceibias.n247 commonsourceibias.n246 161.3
R188 commonsourceibias.n244 commonsourceibias.n206 161.3
R189 commonsourceibias.n243 commonsourceibias.n242 161.3
R190 commonsourceibias.n241 commonsourceibias.n240 161.3
R191 commonsourceibias.n239 commonsourceibias.n208 161.3
R192 commonsourceibias.n238 commonsourceibias.n237 161.3
R193 commonsourceibias.n236 commonsourceibias.n235 161.3
R194 commonsourceibias.n234 commonsourceibias.n210 161.3
R195 commonsourceibias.n233 commonsourceibias.n232 161.3
R196 commonsourceibias.n231 commonsourceibias.n230 161.3
R197 commonsourceibias.n229 commonsourceibias.n212 161.3
R198 commonsourceibias.n227 commonsourceibias.n226 161.3
R199 commonsourceibias.n225 commonsourceibias.n213 161.3
R200 commonsourceibias.n224 commonsourceibias.n223 161.3
R201 commonsourceibias.n221 commonsourceibias.n214 161.3
R202 commonsourceibias.n220 commonsourceibias.n219 161.3
R203 commonsourceibias.n218 commonsourceibias.n215 161.3
R204 commonsourceibias.n429 commonsourceibias.n343 161.3
R205 commonsourceibias.n427 commonsourceibias.n426 161.3
R206 commonsourceibias.n425 commonsourceibias.n344 161.3
R207 commonsourceibias.n424 commonsourceibias.n423 161.3
R208 commonsourceibias.n421 commonsourceibias.n345 161.3
R209 commonsourceibias.n420 commonsourceibias.n419 161.3
R210 commonsourceibias.n418 commonsourceibias.n346 161.3
R211 commonsourceibias.n417 commonsourceibias.n416 161.3
R212 commonsourceibias.n414 commonsourceibias.n347 161.3
R213 commonsourceibias.n412 commonsourceibias.n411 161.3
R214 commonsourceibias.n410 commonsourceibias.n348 161.3
R215 commonsourceibias.n409 commonsourceibias.n408 161.3
R216 commonsourceibias.n406 commonsourceibias.n349 161.3
R217 commonsourceibias.n405 commonsourceibias.n404 161.3
R218 commonsourceibias.n403 commonsourceibias.n350 161.3
R219 commonsourceibias.n402 commonsourceibias.n401 161.3
R220 commonsourceibias.n399 commonsourceibias.n351 161.3
R221 commonsourceibias.n397 commonsourceibias.n396 161.3
R222 commonsourceibias.n395 commonsourceibias.n352 161.3
R223 commonsourceibias.n394 commonsourceibias.n393 161.3
R224 commonsourceibias.n391 commonsourceibias.n353 161.3
R225 commonsourceibias.n390 commonsourceibias.n389 161.3
R226 commonsourceibias.n388 commonsourceibias.n387 161.3
R227 commonsourceibias.n386 commonsourceibias.n355 161.3
R228 commonsourceibias.n385 commonsourceibias.n384 161.3
R229 commonsourceibias.n383 commonsourceibias.n382 161.3
R230 commonsourceibias.n381 commonsourceibias.n357 161.3
R231 commonsourceibias.n380 commonsourceibias.n379 161.3
R232 commonsourceibias.n378 commonsourceibias.n377 161.3
R233 commonsourceibias.n376 commonsourceibias.n359 161.3
R234 commonsourceibias.n374 commonsourceibias.n373 161.3
R235 commonsourceibias.n372 commonsourceibias.n360 161.3
R236 commonsourceibias.n371 commonsourceibias.n370 161.3
R237 commonsourceibias.n368 commonsourceibias.n361 161.3
R238 commonsourceibias.n367 commonsourceibias.n366 161.3
R239 commonsourceibias.n365 commonsourceibias.n362 161.3
R240 commonsourceibias.n335 commonsourceibias.n334 161.3
R241 commonsourceibias.n332 commonsourceibias.n294 161.3
R242 commonsourceibias.n331 commonsourceibias.n330 161.3
R243 commonsourceibias.n329 commonsourceibias.n328 161.3
R244 commonsourceibias.n327 commonsourceibias.n296 161.3
R245 commonsourceibias.n326 commonsourceibias.n325 161.3
R246 commonsourceibias.n324 commonsourceibias.n323 161.3
R247 commonsourceibias.n322 commonsourceibias.n298 161.3
R248 commonsourceibias.n321 commonsourceibias.n320 161.3
R249 commonsourceibias.n319 commonsourceibias.n318 161.3
R250 commonsourceibias.n317 commonsourceibias.n300 161.3
R251 commonsourceibias.n315 commonsourceibias.n314 161.3
R252 commonsourceibias.n313 commonsourceibias.n301 161.3
R253 commonsourceibias.n312 commonsourceibias.n311 161.3
R254 commonsourceibias.n309 commonsourceibias.n302 161.3
R255 commonsourceibias.n308 commonsourceibias.n307 161.3
R256 commonsourceibias.n306 commonsourceibias.n303 161.3
R257 commonsourceibias.n441 commonsourceibias.n293 161.3
R258 commonsourceibias.n475 commonsourceibias.n284 161.3
R259 commonsourceibias.n473 commonsourceibias.n472 161.3
R260 commonsourceibias.n471 commonsourceibias.n285 161.3
R261 commonsourceibias.n470 commonsourceibias.n469 161.3
R262 commonsourceibias.n467 commonsourceibias.n286 161.3
R263 commonsourceibias.n466 commonsourceibias.n465 161.3
R264 commonsourceibias.n464 commonsourceibias.n287 161.3
R265 commonsourceibias.n463 commonsourceibias.n462 161.3
R266 commonsourceibias.n460 commonsourceibias.n288 161.3
R267 commonsourceibias.n458 commonsourceibias.n457 161.3
R268 commonsourceibias.n456 commonsourceibias.n289 161.3
R269 commonsourceibias.n455 commonsourceibias.n454 161.3
R270 commonsourceibias.n452 commonsourceibias.n290 161.3
R271 commonsourceibias.n451 commonsourceibias.n450 161.3
R272 commonsourceibias.n449 commonsourceibias.n291 161.3
R273 commonsourceibias.n448 commonsourceibias.n447 161.3
R274 commonsourceibias.n445 commonsourceibias.n292 161.3
R275 commonsourceibias.n443 commonsourceibias.n442 161.3
R276 commonsourceibias.n564 commonsourceibias.n478 161.3
R277 commonsourceibias.n562 commonsourceibias.n561 161.3
R278 commonsourceibias.n560 commonsourceibias.n479 161.3
R279 commonsourceibias.n559 commonsourceibias.n558 161.3
R280 commonsourceibias.n556 commonsourceibias.n480 161.3
R281 commonsourceibias.n555 commonsourceibias.n554 161.3
R282 commonsourceibias.n553 commonsourceibias.n481 161.3
R283 commonsourceibias.n552 commonsourceibias.n551 161.3
R284 commonsourceibias.n549 commonsourceibias.n482 161.3
R285 commonsourceibias.n547 commonsourceibias.n546 161.3
R286 commonsourceibias.n545 commonsourceibias.n483 161.3
R287 commonsourceibias.n544 commonsourceibias.n543 161.3
R288 commonsourceibias.n541 commonsourceibias.n484 161.3
R289 commonsourceibias.n540 commonsourceibias.n539 161.3
R290 commonsourceibias.n538 commonsourceibias.n485 161.3
R291 commonsourceibias.n537 commonsourceibias.n536 161.3
R292 commonsourceibias.n534 commonsourceibias.n486 161.3
R293 commonsourceibias.n532 commonsourceibias.n531 161.3
R294 commonsourceibias.n530 commonsourceibias.n487 161.3
R295 commonsourceibias.n529 commonsourceibias.n528 161.3
R296 commonsourceibias.n526 commonsourceibias.n488 161.3
R297 commonsourceibias.n525 commonsourceibias.n524 161.3
R298 commonsourceibias.n523 commonsourceibias.n522 161.3
R299 commonsourceibias.n521 commonsourceibias.n490 161.3
R300 commonsourceibias.n520 commonsourceibias.n519 161.3
R301 commonsourceibias.n518 commonsourceibias.n517 161.3
R302 commonsourceibias.n516 commonsourceibias.n492 161.3
R303 commonsourceibias.n515 commonsourceibias.n514 161.3
R304 commonsourceibias.n513 commonsourceibias.n512 161.3
R305 commonsourceibias.n511 commonsourceibias.n494 161.3
R306 commonsourceibias.n509 commonsourceibias.n508 161.3
R307 commonsourceibias.n507 commonsourceibias.n495 161.3
R308 commonsourceibias.n506 commonsourceibias.n505 161.3
R309 commonsourceibias.n503 commonsourceibias.n496 161.3
R310 commonsourceibias.n502 commonsourceibias.n501 161.3
R311 commonsourceibias.n500 commonsourceibias.n497 161.3
R312 commonsourceibias.n111 commonsourceibias.n109 81.5057
R313 commonsourceibias.n338 commonsourceibias.n336 81.5057
R314 commonsourceibias.n111 commonsourceibias.n110 80.9324
R315 commonsourceibias.n113 commonsourceibias.n112 80.9324
R316 commonsourceibias.n115 commonsourceibias.n114 80.9324
R317 commonsourceibias.n108 commonsourceibias.n107 80.9324
R318 commonsourceibias.n106 commonsourceibias.n105 80.9324
R319 commonsourceibias.n104 commonsourceibias.n103 80.9324
R320 commonsourceibias.n102 commonsourceibias.n101 80.9324
R321 commonsourceibias.n433 commonsourceibias.n432 80.9324
R322 commonsourceibias.n435 commonsourceibias.n434 80.9324
R323 commonsourceibias.n437 commonsourceibias.n436 80.9324
R324 commonsourceibias.n439 commonsourceibias.n438 80.9324
R325 commonsourceibias.n342 commonsourceibias.n341 80.9324
R326 commonsourceibias.n340 commonsourceibias.n339 80.9324
R327 commonsourceibias.n338 commonsourceibias.n337 80.9324
R328 commonsourceibias.n100 commonsourceibias.n99 80.6037
R329 commonsourceibias.n193 commonsourceibias.n192 80.6037
R330 commonsourceibias.n282 commonsourceibias.n281 80.6037
R331 commonsourceibias.n431 commonsourceibias.n430 80.6037
R332 commonsourceibias.n477 commonsourceibias.n476 80.6037
R333 commonsourceibias.n566 commonsourceibias.n565 80.6037
R334 commonsourceibias.n85 commonsourceibias.n84 56.5617
R335 commonsourceibias.n71 commonsourceibias.n70 56.5617
R336 commonsourceibias.n62 commonsourceibias.n61 56.5617
R337 commonsourceibias.n48 commonsourceibias.n47 56.5617
R338 commonsourceibias.n178 commonsourceibias.n177 56.5617
R339 commonsourceibias.n164 commonsourceibias.n163 56.5617
R340 commonsourceibias.n155 commonsourceibias.n154 56.5617
R341 commonsourceibias.n141 commonsourceibias.n140 56.5617
R342 commonsourceibias.n230 commonsourceibias.n229 56.5617
R343 commonsourceibias.n244 commonsourceibias.n243 56.5617
R344 commonsourceibias.n253 commonsourceibias.n252 56.5617
R345 commonsourceibias.n267 commonsourceibias.n266 56.5617
R346 commonsourceibias.n377 commonsourceibias.n376 56.5617
R347 commonsourceibias.n391 commonsourceibias.n390 56.5617
R348 commonsourceibias.n401 commonsourceibias.n399 56.5617
R349 commonsourceibias.n416 commonsourceibias.n414 56.5617
R350 commonsourceibias.n462 commonsourceibias.n460 56.5617
R351 commonsourceibias.n447 commonsourceibias.n445 56.5617
R352 commonsourceibias.n318 commonsourceibias.n317 56.5617
R353 commonsourceibias.n332 commonsourceibias.n331 56.5617
R354 commonsourceibias.n512 commonsourceibias.n511 56.5617
R355 commonsourceibias.n526 commonsourceibias.n525 56.5617
R356 commonsourceibias.n536 commonsourceibias.n534 56.5617
R357 commonsourceibias.n551 commonsourceibias.n549 56.5617
R358 commonsourceibias.n76 commonsourceibias.n75 56.0773
R359 commonsourceibias.n57 commonsourceibias.n56 56.0773
R360 commonsourceibias.n169 commonsourceibias.n168 56.0773
R361 commonsourceibias.n150 commonsourceibias.n149 56.0773
R362 commonsourceibias.n239 commonsourceibias.n238 56.0773
R363 commonsourceibias.n258 commonsourceibias.n257 56.0773
R364 commonsourceibias.n386 commonsourceibias.n385 56.0773
R365 commonsourceibias.n406 commonsourceibias.n405 56.0773
R366 commonsourceibias.n452 commonsourceibias.n451 56.0773
R367 commonsourceibias.n327 commonsourceibias.n326 56.0773
R368 commonsourceibias.n521 commonsourceibias.n520 56.0773
R369 commonsourceibias.n541 commonsourceibias.n540 56.0773
R370 commonsourceibias.n99 commonsourceibias.n98 55.3321
R371 commonsourceibias.n192 commonsourceibias.n191 55.3321
R372 commonsourceibias.n281 commonsourceibias.n280 55.3321
R373 commonsourceibias.n430 commonsourceibias.n429 55.3321
R374 commonsourceibias.n476 commonsourceibias.n475 55.3321
R375 commonsourceibias.n565 commonsourceibias.n564 55.3321
R376 commonsourceibias.n90 commonsourceibias.n89 55.1086
R377 commonsourceibias.n41 commonsourceibias.n31 55.1086
R378 commonsourceibias.n183 commonsourceibias.n182 55.1086
R379 commonsourceibias.n134 commonsourceibias.n124 55.1086
R380 commonsourceibias.n223 commonsourceibias.n213 55.1086
R381 commonsourceibias.n272 commonsourceibias.n271 55.1086
R382 commonsourceibias.n370 commonsourceibias.n360 55.1086
R383 commonsourceibias.n421 commonsourceibias.n420 55.1086
R384 commonsourceibias.n467 commonsourceibias.n466 55.1086
R385 commonsourceibias.n311 commonsourceibias.n301 55.1086
R386 commonsourceibias.n505 commonsourceibias.n495 55.1086
R387 commonsourceibias.n556 commonsourceibias.n555 55.1086
R388 commonsourceibias.n35 commonsourceibias.n34 47.4592
R389 commonsourceibias.n128 commonsourceibias.n127 47.4592
R390 commonsourceibias.n217 commonsourceibias.n216 47.4592
R391 commonsourceibias.n364 commonsourceibias.n363 47.4592
R392 commonsourceibias.n305 commonsourceibias.n304 47.4592
R393 commonsourceibias.n499 commonsourceibias.n498 47.4592
R394 commonsourceibias.n218 commonsourceibias.n217 44.0436
R395 commonsourceibias.n365 commonsourceibias.n364 44.0436
R396 commonsourceibias.n306 commonsourceibias.n305 44.0436
R397 commonsourceibias.n500 commonsourceibias.n499 44.0436
R398 commonsourceibias.n36 commonsourceibias.n35 44.0436
R399 commonsourceibias.n129 commonsourceibias.n128 44.0436
R400 commonsourceibias.n92 commonsourceibias.n13 42.5146
R401 commonsourceibias.n39 commonsourceibias.n38 42.5146
R402 commonsourceibias.n185 commonsourceibias.n1 42.5146
R403 commonsourceibias.n132 commonsourceibias.n131 42.5146
R404 commonsourceibias.n221 commonsourceibias.n220 42.5146
R405 commonsourceibias.n274 commonsourceibias.n195 42.5146
R406 commonsourceibias.n368 commonsourceibias.n367 42.5146
R407 commonsourceibias.n423 commonsourceibias.n344 42.5146
R408 commonsourceibias.n469 commonsourceibias.n285 42.5146
R409 commonsourceibias.n309 commonsourceibias.n308 42.5146
R410 commonsourceibias.n503 commonsourceibias.n502 42.5146
R411 commonsourceibias.n558 commonsourceibias.n479 42.5146
R412 commonsourceibias.n78 commonsourceibias.n18 41.5458
R413 commonsourceibias.n53 commonsourceibias.n52 41.5458
R414 commonsourceibias.n171 commonsourceibias.n6 41.5458
R415 commonsourceibias.n146 commonsourceibias.n145 41.5458
R416 commonsourceibias.n235 commonsourceibias.n234 41.5458
R417 commonsourceibias.n260 commonsourceibias.n200 41.5458
R418 commonsourceibias.n382 commonsourceibias.n381 41.5458
R419 commonsourceibias.n408 commonsourceibias.n348 41.5458
R420 commonsourceibias.n454 commonsourceibias.n289 41.5458
R421 commonsourceibias.n323 commonsourceibias.n322 41.5458
R422 commonsourceibias.n517 commonsourceibias.n516 41.5458
R423 commonsourceibias.n543 commonsourceibias.n483 41.5458
R424 commonsourceibias.n68 commonsourceibias.n23 40.577
R425 commonsourceibias.n64 commonsourceibias.n23 40.577
R426 commonsourceibias.n161 commonsourceibias.n11 40.577
R427 commonsourceibias.n157 commonsourceibias.n11 40.577
R428 commonsourceibias.n246 commonsourceibias.n205 40.577
R429 commonsourceibias.n250 commonsourceibias.n205 40.577
R430 commonsourceibias.n393 commonsourceibias.n352 40.577
R431 commonsourceibias.n397 commonsourceibias.n352 40.577
R432 commonsourceibias.n443 commonsourceibias.n293 40.577
R433 commonsourceibias.n334 commonsourceibias.n293 40.577
R434 commonsourceibias.n528 commonsourceibias.n487 40.577
R435 commonsourceibias.n532 commonsourceibias.n487 40.577
R436 commonsourceibias.n82 commonsourceibias.n18 39.6083
R437 commonsourceibias.n52 commonsourceibias.n51 39.6083
R438 commonsourceibias.n175 commonsourceibias.n6 39.6083
R439 commonsourceibias.n145 commonsourceibias.n144 39.6083
R440 commonsourceibias.n234 commonsourceibias.n233 39.6083
R441 commonsourceibias.n264 commonsourceibias.n200 39.6083
R442 commonsourceibias.n381 commonsourceibias.n380 39.6083
R443 commonsourceibias.n412 commonsourceibias.n348 39.6083
R444 commonsourceibias.n458 commonsourceibias.n289 39.6083
R445 commonsourceibias.n322 commonsourceibias.n321 39.6083
R446 commonsourceibias.n516 commonsourceibias.n515 39.6083
R447 commonsourceibias.n547 commonsourceibias.n483 39.6083
R448 commonsourceibias.n96 commonsourceibias.n13 38.6395
R449 commonsourceibias.n38 commonsourceibias.n33 38.6395
R450 commonsourceibias.n189 commonsourceibias.n1 38.6395
R451 commonsourceibias.n131 commonsourceibias.n126 38.6395
R452 commonsourceibias.n220 commonsourceibias.n215 38.6395
R453 commonsourceibias.n278 commonsourceibias.n195 38.6395
R454 commonsourceibias.n367 commonsourceibias.n362 38.6395
R455 commonsourceibias.n427 commonsourceibias.n344 38.6395
R456 commonsourceibias.n473 commonsourceibias.n285 38.6395
R457 commonsourceibias.n308 commonsourceibias.n303 38.6395
R458 commonsourceibias.n502 commonsourceibias.n497 38.6395
R459 commonsourceibias.n562 commonsourceibias.n479 38.6395
R460 commonsourceibias.n89 commonsourceibias.n15 26.0455
R461 commonsourceibias.n45 commonsourceibias.n31 26.0455
R462 commonsourceibias.n182 commonsourceibias.n3 26.0455
R463 commonsourceibias.n138 commonsourceibias.n124 26.0455
R464 commonsourceibias.n227 commonsourceibias.n213 26.0455
R465 commonsourceibias.n271 commonsourceibias.n197 26.0455
R466 commonsourceibias.n374 commonsourceibias.n360 26.0455
R467 commonsourceibias.n420 commonsourceibias.n346 26.0455
R468 commonsourceibias.n466 commonsourceibias.n287 26.0455
R469 commonsourceibias.n315 commonsourceibias.n301 26.0455
R470 commonsourceibias.n509 commonsourceibias.n495 26.0455
R471 commonsourceibias.n555 commonsourceibias.n481 26.0455
R472 commonsourceibias.n75 commonsourceibias.n20 25.0767
R473 commonsourceibias.n58 commonsourceibias.n57 25.0767
R474 commonsourceibias.n168 commonsourceibias.n8 25.0767
R475 commonsourceibias.n151 commonsourceibias.n150 25.0767
R476 commonsourceibias.n240 commonsourceibias.n239 25.0767
R477 commonsourceibias.n257 commonsourceibias.n202 25.0767
R478 commonsourceibias.n387 commonsourceibias.n386 25.0767
R479 commonsourceibias.n405 commonsourceibias.n350 25.0767
R480 commonsourceibias.n451 commonsourceibias.n291 25.0767
R481 commonsourceibias.n328 commonsourceibias.n327 25.0767
R482 commonsourceibias.n522 commonsourceibias.n521 25.0767
R483 commonsourceibias.n540 commonsourceibias.n485 25.0767
R484 commonsourceibias.n71 commonsourceibias.n22 24.3464
R485 commonsourceibias.n61 commonsourceibias.n25 24.3464
R486 commonsourceibias.n164 commonsourceibias.n10 24.3464
R487 commonsourceibias.n154 commonsourceibias.n118 24.3464
R488 commonsourceibias.n243 commonsourceibias.n207 24.3464
R489 commonsourceibias.n253 commonsourceibias.n204 24.3464
R490 commonsourceibias.n390 commonsourceibias.n354 24.3464
R491 commonsourceibias.n401 commonsourceibias.n400 24.3464
R492 commonsourceibias.n447 commonsourceibias.n446 24.3464
R493 commonsourceibias.n331 commonsourceibias.n295 24.3464
R494 commonsourceibias.n525 commonsourceibias.n489 24.3464
R495 commonsourceibias.n536 commonsourceibias.n535 24.3464
R496 commonsourceibias.n85 commonsourceibias.n17 23.8546
R497 commonsourceibias.n47 commonsourceibias.n46 23.8546
R498 commonsourceibias.n178 commonsourceibias.n5 23.8546
R499 commonsourceibias.n140 commonsourceibias.n139 23.8546
R500 commonsourceibias.n229 commonsourceibias.n228 23.8546
R501 commonsourceibias.n267 commonsourceibias.n199 23.8546
R502 commonsourceibias.n376 commonsourceibias.n375 23.8546
R503 commonsourceibias.n416 commonsourceibias.n415 23.8546
R504 commonsourceibias.n462 commonsourceibias.n461 23.8546
R505 commonsourceibias.n317 commonsourceibias.n316 23.8546
R506 commonsourceibias.n511 commonsourceibias.n510 23.8546
R507 commonsourceibias.n551 commonsourceibias.n550 23.8546
R508 commonsourceibias.n98 commonsourceibias.n97 17.4607
R509 commonsourceibias.n191 commonsourceibias.n190 17.4607
R510 commonsourceibias.n280 commonsourceibias.n279 17.4607
R511 commonsourceibias.n429 commonsourceibias.n428 17.4607
R512 commonsourceibias.n475 commonsourceibias.n474 17.4607
R513 commonsourceibias.n564 commonsourceibias.n563 17.4607
R514 commonsourceibias.n84 commonsourceibias.n83 16.9689
R515 commonsourceibias.n48 commonsourceibias.n29 16.9689
R516 commonsourceibias.n177 commonsourceibias.n176 16.9689
R517 commonsourceibias.n141 commonsourceibias.n122 16.9689
R518 commonsourceibias.n230 commonsourceibias.n211 16.9689
R519 commonsourceibias.n266 commonsourceibias.n265 16.9689
R520 commonsourceibias.n377 commonsourceibias.n358 16.9689
R521 commonsourceibias.n414 commonsourceibias.n413 16.9689
R522 commonsourceibias.n460 commonsourceibias.n459 16.9689
R523 commonsourceibias.n318 commonsourceibias.n299 16.9689
R524 commonsourceibias.n512 commonsourceibias.n493 16.9689
R525 commonsourceibias.n549 commonsourceibias.n548 16.9689
R526 commonsourceibias.n70 commonsourceibias.n69 16.477
R527 commonsourceibias.n63 commonsourceibias.n62 16.477
R528 commonsourceibias.n163 commonsourceibias.n162 16.477
R529 commonsourceibias.n156 commonsourceibias.n155 16.477
R530 commonsourceibias.n245 commonsourceibias.n244 16.477
R531 commonsourceibias.n252 commonsourceibias.n251 16.477
R532 commonsourceibias.n392 commonsourceibias.n391 16.477
R533 commonsourceibias.n399 commonsourceibias.n398 16.477
R534 commonsourceibias.n445 commonsourceibias.n444 16.477
R535 commonsourceibias.n333 commonsourceibias.n332 16.477
R536 commonsourceibias.n527 commonsourceibias.n526 16.477
R537 commonsourceibias.n534 commonsourceibias.n533 16.477
R538 commonsourceibias.n77 commonsourceibias.n76 15.9852
R539 commonsourceibias.n56 commonsourceibias.n27 15.9852
R540 commonsourceibias.n170 commonsourceibias.n169 15.9852
R541 commonsourceibias.n149 commonsourceibias.n120 15.9852
R542 commonsourceibias.n238 commonsourceibias.n209 15.9852
R543 commonsourceibias.n259 commonsourceibias.n258 15.9852
R544 commonsourceibias.n385 commonsourceibias.n356 15.9852
R545 commonsourceibias.n407 commonsourceibias.n406 15.9852
R546 commonsourceibias.n453 commonsourceibias.n452 15.9852
R547 commonsourceibias.n326 commonsourceibias.n297 15.9852
R548 commonsourceibias.n520 commonsourceibias.n491 15.9852
R549 commonsourceibias.n542 commonsourceibias.n541 15.9852
R550 commonsourceibias.n91 commonsourceibias.n90 15.4934
R551 commonsourceibias.n41 commonsourceibias.n40 15.4934
R552 commonsourceibias.n184 commonsourceibias.n183 15.4934
R553 commonsourceibias.n134 commonsourceibias.n133 15.4934
R554 commonsourceibias.n223 commonsourceibias.n222 15.4934
R555 commonsourceibias.n273 commonsourceibias.n272 15.4934
R556 commonsourceibias.n370 commonsourceibias.n369 15.4934
R557 commonsourceibias.n422 commonsourceibias.n421 15.4934
R558 commonsourceibias.n468 commonsourceibias.n467 15.4934
R559 commonsourceibias.n311 commonsourceibias.n310 15.4934
R560 commonsourceibias.n505 commonsourceibias.n504 15.4934
R561 commonsourceibias.n557 commonsourceibias.n556 15.4934
R562 commonsourceibias.n102 commonsourceibias.n100 13.2663
R563 commonsourceibias.n433 commonsourceibias.n431 13.2663
R564 commonsourceibias.n568 commonsourceibias.n283 11.9876
R565 commonsourceibias.n568 commonsourceibias.n567 10.3347
R566 commonsourceibias.n159 commonsourceibias.n116 9.50363
R567 commonsourceibias.n441 commonsourceibias.n440 9.50363
R568 commonsourceibias.n92 commonsourceibias.n91 9.09948
R569 commonsourceibias.n40 commonsourceibias.n39 9.09948
R570 commonsourceibias.n185 commonsourceibias.n184 9.09948
R571 commonsourceibias.n133 commonsourceibias.n132 9.09948
R572 commonsourceibias.n222 commonsourceibias.n221 9.09948
R573 commonsourceibias.n274 commonsourceibias.n273 9.09948
R574 commonsourceibias.n369 commonsourceibias.n368 9.09948
R575 commonsourceibias.n423 commonsourceibias.n422 9.09948
R576 commonsourceibias.n469 commonsourceibias.n468 9.09948
R577 commonsourceibias.n310 commonsourceibias.n309 9.09948
R578 commonsourceibias.n504 commonsourceibias.n503 9.09948
R579 commonsourceibias.n558 commonsourceibias.n557 9.09948
R580 commonsourceibias.n283 commonsourceibias.n193 8.79261
R581 commonsourceibias.n567 commonsourceibias.n477 8.79261
R582 commonsourceibias.n78 commonsourceibias.n77 8.60764
R583 commonsourceibias.n53 commonsourceibias.n27 8.60764
R584 commonsourceibias.n171 commonsourceibias.n170 8.60764
R585 commonsourceibias.n146 commonsourceibias.n120 8.60764
R586 commonsourceibias.n235 commonsourceibias.n209 8.60764
R587 commonsourceibias.n260 commonsourceibias.n259 8.60764
R588 commonsourceibias.n382 commonsourceibias.n356 8.60764
R589 commonsourceibias.n408 commonsourceibias.n407 8.60764
R590 commonsourceibias.n454 commonsourceibias.n453 8.60764
R591 commonsourceibias.n323 commonsourceibias.n297 8.60764
R592 commonsourceibias.n517 commonsourceibias.n491 8.60764
R593 commonsourceibias.n543 commonsourceibias.n542 8.60764
R594 commonsourceibias.n69 commonsourceibias.n68 8.11581
R595 commonsourceibias.n64 commonsourceibias.n63 8.11581
R596 commonsourceibias.n162 commonsourceibias.n161 8.11581
R597 commonsourceibias.n157 commonsourceibias.n156 8.11581
R598 commonsourceibias.n246 commonsourceibias.n245 8.11581
R599 commonsourceibias.n251 commonsourceibias.n250 8.11581
R600 commonsourceibias.n393 commonsourceibias.n392 8.11581
R601 commonsourceibias.n398 commonsourceibias.n397 8.11581
R602 commonsourceibias.n444 commonsourceibias.n443 8.11581
R603 commonsourceibias.n334 commonsourceibias.n333 8.11581
R604 commonsourceibias.n528 commonsourceibias.n527 8.11581
R605 commonsourceibias.n533 commonsourceibias.n532 8.11581
R606 commonsourceibias.n83 commonsourceibias.n82 7.62397
R607 commonsourceibias.n51 commonsourceibias.n29 7.62397
R608 commonsourceibias.n176 commonsourceibias.n175 7.62397
R609 commonsourceibias.n144 commonsourceibias.n122 7.62397
R610 commonsourceibias.n233 commonsourceibias.n211 7.62397
R611 commonsourceibias.n265 commonsourceibias.n264 7.62397
R612 commonsourceibias.n380 commonsourceibias.n358 7.62397
R613 commonsourceibias.n413 commonsourceibias.n412 7.62397
R614 commonsourceibias.n459 commonsourceibias.n458 7.62397
R615 commonsourceibias.n321 commonsourceibias.n299 7.62397
R616 commonsourceibias.n515 commonsourceibias.n493 7.62397
R617 commonsourceibias.n548 commonsourceibias.n547 7.62397
R618 commonsourceibias.n97 commonsourceibias.n96 7.13213
R619 commonsourceibias.n34 commonsourceibias.n33 7.13213
R620 commonsourceibias.n190 commonsourceibias.n189 7.13213
R621 commonsourceibias.n127 commonsourceibias.n126 7.13213
R622 commonsourceibias.n216 commonsourceibias.n215 7.13213
R623 commonsourceibias.n279 commonsourceibias.n278 7.13213
R624 commonsourceibias.n363 commonsourceibias.n362 7.13213
R625 commonsourceibias.n428 commonsourceibias.n427 7.13213
R626 commonsourceibias.n474 commonsourceibias.n473 7.13213
R627 commonsourceibias.n304 commonsourceibias.n303 7.13213
R628 commonsourceibias.n498 commonsourceibias.n497 7.13213
R629 commonsourceibias.n563 commonsourceibias.n562 7.13213
R630 commonsourceibias.n283 commonsourceibias.n282 5.06534
R631 commonsourceibias.n567 commonsourceibias.n566 5.06534
R632 commonsourceibias commonsourceibias.n568 4.04308
R633 commonsourceibias.n109 commonsourceibias.t27 2.82907
R634 commonsourceibias.n109 commonsourceibias.t11 2.82907
R635 commonsourceibias.n110 commonsourceibias.t33 2.82907
R636 commonsourceibias.n110 commonsourceibias.t1 2.82907
R637 commonsourceibias.n112 commonsourceibias.t7 2.82907
R638 commonsourceibias.n112 commonsourceibias.t63 2.82907
R639 commonsourceibias.n114 commonsourceibias.t57 2.82907
R640 commonsourceibias.n114 commonsourceibias.t39 2.82907
R641 commonsourceibias.n107 commonsourceibias.t61 2.82907
R642 commonsourceibias.n107 commonsourceibias.t17 2.82907
R643 commonsourceibias.n105 commonsourceibias.t21 2.82907
R644 commonsourceibias.n105 commonsourceibias.t59 2.82907
R645 commonsourceibias.n103 commonsourceibias.t15 2.82907
R646 commonsourceibias.n103 commonsourceibias.t53 2.82907
R647 commonsourceibias.n101 commonsourceibias.t55 2.82907
R648 commonsourceibias.n101 commonsourceibias.t25 2.82907
R649 commonsourceibias.n432 commonsourceibias.t23 2.82907
R650 commonsourceibias.n432 commonsourceibias.t45 2.82907
R651 commonsourceibias.n434 commonsourceibias.t43 2.82907
R652 commonsourceibias.n434 commonsourceibias.t3 2.82907
R653 commonsourceibias.n436 commonsourceibias.t49 2.82907
R654 commonsourceibias.n436 commonsourceibias.t51 2.82907
R655 commonsourceibias.n438 commonsourceibias.t9 2.82907
R656 commonsourceibias.n438 commonsourceibias.t41 2.82907
R657 commonsourceibias.n341 commonsourceibias.t19 2.82907
R658 commonsourceibias.n341 commonsourceibias.t47 2.82907
R659 commonsourceibias.n339 commonsourceibias.t31 2.82907
R660 commonsourceibias.n339 commonsourceibias.t37 2.82907
R661 commonsourceibias.n337 commonsourceibias.t35 2.82907
R662 commonsourceibias.n337 commonsourceibias.t13 2.82907
R663 commonsourceibias.n336 commonsourceibias.t5 2.82907
R664 commonsourceibias.n336 commonsourceibias.t29 2.82907
R665 commonsourceibias.n17 commonsourceibias.n15 0.738255
R666 commonsourceibias.n46 commonsourceibias.n45 0.738255
R667 commonsourceibias.n5 commonsourceibias.n3 0.738255
R668 commonsourceibias.n139 commonsourceibias.n138 0.738255
R669 commonsourceibias.n228 commonsourceibias.n227 0.738255
R670 commonsourceibias.n199 commonsourceibias.n197 0.738255
R671 commonsourceibias.n375 commonsourceibias.n374 0.738255
R672 commonsourceibias.n415 commonsourceibias.n346 0.738255
R673 commonsourceibias.n461 commonsourceibias.n287 0.738255
R674 commonsourceibias.n316 commonsourceibias.n315 0.738255
R675 commonsourceibias.n510 commonsourceibias.n509 0.738255
R676 commonsourceibias.n550 commonsourceibias.n481 0.738255
R677 commonsourceibias.n104 commonsourceibias.n102 0.573776
R678 commonsourceibias.n106 commonsourceibias.n104 0.573776
R679 commonsourceibias.n108 commonsourceibias.n106 0.573776
R680 commonsourceibias.n115 commonsourceibias.n113 0.573776
R681 commonsourceibias.n113 commonsourceibias.n111 0.573776
R682 commonsourceibias.n340 commonsourceibias.n338 0.573776
R683 commonsourceibias.n342 commonsourceibias.n340 0.573776
R684 commonsourceibias.n439 commonsourceibias.n437 0.573776
R685 commonsourceibias.n437 commonsourceibias.n435 0.573776
R686 commonsourceibias.n435 commonsourceibias.n433 0.573776
R687 commonsourceibias.n116 commonsourceibias.n108 0.287138
R688 commonsourceibias.n116 commonsourceibias.n115 0.287138
R689 commonsourceibias.n440 commonsourceibias.n342 0.287138
R690 commonsourceibias.n440 commonsourceibias.n439 0.287138
R691 commonsourceibias.n100 commonsourceibias.n12 0.285035
R692 commonsourceibias.n193 commonsourceibias.n0 0.285035
R693 commonsourceibias.n282 commonsourceibias.n194 0.285035
R694 commonsourceibias.n431 commonsourceibias.n343 0.285035
R695 commonsourceibias.n477 commonsourceibias.n284 0.285035
R696 commonsourceibias.n566 commonsourceibias.n478 0.285035
R697 commonsourceibias.n22 commonsourceibias.n20 0.246418
R698 commonsourceibias.n58 commonsourceibias.n25 0.246418
R699 commonsourceibias.n10 commonsourceibias.n8 0.246418
R700 commonsourceibias.n151 commonsourceibias.n118 0.246418
R701 commonsourceibias.n240 commonsourceibias.n207 0.246418
R702 commonsourceibias.n204 commonsourceibias.n202 0.246418
R703 commonsourceibias.n387 commonsourceibias.n354 0.246418
R704 commonsourceibias.n400 commonsourceibias.n350 0.246418
R705 commonsourceibias.n446 commonsourceibias.n291 0.246418
R706 commonsourceibias.n328 commonsourceibias.n295 0.246418
R707 commonsourceibias.n522 commonsourceibias.n489 0.246418
R708 commonsourceibias.n535 commonsourceibias.n485 0.246418
R709 commonsourceibias.n95 commonsourceibias.n12 0.189894
R710 commonsourceibias.n95 commonsourceibias.n94 0.189894
R711 commonsourceibias.n94 commonsourceibias.n93 0.189894
R712 commonsourceibias.n93 commonsourceibias.n14 0.189894
R713 commonsourceibias.n88 commonsourceibias.n14 0.189894
R714 commonsourceibias.n88 commonsourceibias.n87 0.189894
R715 commonsourceibias.n87 commonsourceibias.n86 0.189894
R716 commonsourceibias.n86 commonsourceibias.n16 0.189894
R717 commonsourceibias.n81 commonsourceibias.n16 0.189894
R718 commonsourceibias.n81 commonsourceibias.n80 0.189894
R719 commonsourceibias.n80 commonsourceibias.n79 0.189894
R720 commonsourceibias.n79 commonsourceibias.n19 0.189894
R721 commonsourceibias.n74 commonsourceibias.n19 0.189894
R722 commonsourceibias.n74 commonsourceibias.n73 0.189894
R723 commonsourceibias.n73 commonsourceibias.n72 0.189894
R724 commonsourceibias.n72 commonsourceibias.n21 0.189894
R725 commonsourceibias.n67 commonsourceibias.n21 0.189894
R726 commonsourceibias.n67 commonsourceibias.n66 0.189894
R727 commonsourceibias.n66 commonsourceibias.n65 0.189894
R728 commonsourceibias.n65 commonsourceibias.n24 0.189894
R729 commonsourceibias.n60 commonsourceibias.n24 0.189894
R730 commonsourceibias.n60 commonsourceibias.n59 0.189894
R731 commonsourceibias.n59 commonsourceibias.n26 0.189894
R732 commonsourceibias.n55 commonsourceibias.n26 0.189894
R733 commonsourceibias.n55 commonsourceibias.n54 0.189894
R734 commonsourceibias.n54 commonsourceibias.n28 0.189894
R735 commonsourceibias.n50 commonsourceibias.n28 0.189894
R736 commonsourceibias.n50 commonsourceibias.n49 0.189894
R737 commonsourceibias.n49 commonsourceibias.n30 0.189894
R738 commonsourceibias.n44 commonsourceibias.n30 0.189894
R739 commonsourceibias.n44 commonsourceibias.n43 0.189894
R740 commonsourceibias.n43 commonsourceibias.n42 0.189894
R741 commonsourceibias.n42 commonsourceibias.n32 0.189894
R742 commonsourceibias.n37 commonsourceibias.n32 0.189894
R743 commonsourceibias.n37 commonsourceibias.n36 0.189894
R744 commonsourceibias.n158 commonsourceibias.n117 0.189894
R745 commonsourceibias.n153 commonsourceibias.n117 0.189894
R746 commonsourceibias.n153 commonsourceibias.n152 0.189894
R747 commonsourceibias.n152 commonsourceibias.n119 0.189894
R748 commonsourceibias.n148 commonsourceibias.n119 0.189894
R749 commonsourceibias.n148 commonsourceibias.n147 0.189894
R750 commonsourceibias.n147 commonsourceibias.n121 0.189894
R751 commonsourceibias.n143 commonsourceibias.n121 0.189894
R752 commonsourceibias.n143 commonsourceibias.n142 0.189894
R753 commonsourceibias.n142 commonsourceibias.n123 0.189894
R754 commonsourceibias.n137 commonsourceibias.n123 0.189894
R755 commonsourceibias.n137 commonsourceibias.n136 0.189894
R756 commonsourceibias.n136 commonsourceibias.n135 0.189894
R757 commonsourceibias.n135 commonsourceibias.n125 0.189894
R758 commonsourceibias.n130 commonsourceibias.n125 0.189894
R759 commonsourceibias.n130 commonsourceibias.n129 0.189894
R760 commonsourceibias.n188 commonsourceibias.n0 0.189894
R761 commonsourceibias.n188 commonsourceibias.n187 0.189894
R762 commonsourceibias.n187 commonsourceibias.n186 0.189894
R763 commonsourceibias.n186 commonsourceibias.n2 0.189894
R764 commonsourceibias.n181 commonsourceibias.n2 0.189894
R765 commonsourceibias.n181 commonsourceibias.n180 0.189894
R766 commonsourceibias.n180 commonsourceibias.n179 0.189894
R767 commonsourceibias.n179 commonsourceibias.n4 0.189894
R768 commonsourceibias.n174 commonsourceibias.n4 0.189894
R769 commonsourceibias.n174 commonsourceibias.n173 0.189894
R770 commonsourceibias.n173 commonsourceibias.n172 0.189894
R771 commonsourceibias.n172 commonsourceibias.n7 0.189894
R772 commonsourceibias.n167 commonsourceibias.n7 0.189894
R773 commonsourceibias.n167 commonsourceibias.n166 0.189894
R774 commonsourceibias.n166 commonsourceibias.n165 0.189894
R775 commonsourceibias.n165 commonsourceibias.n9 0.189894
R776 commonsourceibias.n160 commonsourceibias.n9 0.189894
R777 commonsourceibias.n277 commonsourceibias.n194 0.189894
R778 commonsourceibias.n277 commonsourceibias.n276 0.189894
R779 commonsourceibias.n276 commonsourceibias.n275 0.189894
R780 commonsourceibias.n275 commonsourceibias.n196 0.189894
R781 commonsourceibias.n270 commonsourceibias.n196 0.189894
R782 commonsourceibias.n270 commonsourceibias.n269 0.189894
R783 commonsourceibias.n269 commonsourceibias.n268 0.189894
R784 commonsourceibias.n268 commonsourceibias.n198 0.189894
R785 commonsourceibias.n263 commonsourceibias.n198 0.189894
R786 commonsourceibias.n263 commonsourceibias.n262 0.189894
R787 commonsourceibias.n262 commonsourceibias.n261 0.189894
R788 commonsourceibias.n261 commonsourceibias.n201 0.189894
R789 commonsourceibias.n256 commonsourceibias.n201 0.189894
R790 commonsourceibias.n256 commonsourceibias.n255 0.189894
R791 commonsourceibias.n255 commonsourceibias.n254 0.189894
R792 commonsourceibias.n254 commonsourceibias.n203 0.189894
R793 commonsourceibias.n249 commonsourceibias.n203 0.189894
R794 commonsourceibias.n249 commonsourceibias.n248 0.189894
R795 commonsourceibias.n248 commonsourceibias.n247 0.189894
R796 commonsourceibias.n247 commonsourceibias.n206 0.189894
R797 commonsourceibias.n242 commonsourceibias.n206 0.189894
R798 commonsourceibias.n242 commonsourceibias.n241 0.189894
R799 commonsourceibias.n241 commonsourceibias.n208 0.189894
R800 commonsourceibias.n237 commonsourceibias.n208 0.189894
R801 commonsourceibias.n237 commonsourceibias.n236 0.189894
R802 commonsourceibias.n236 commonsourceibias.n210 0.189894
R803 commonsourceibias.n232 commonsourceibias.n210 0.189894
R804 commonsourceibias.n232 commonsourceibias.n231 0.189894
R805 commonsourceibias.n231 commonsourceibias.n212 0.189894
R806 commonsourceibias.n226 commonsourceibias.n212 0.189894
R807 commonsourceibias.n226 commonsourceibias.n225 0.189894
R808 commonsourceibias.n225 commonsourceibias.n224 0.189894
R809 commonsourceibias.n224 commonsourceibias.n214 0.189894
R810 commonsourceibias.n219 commonsourceibias.n214 0.189894
R811 commonsourceibias.n219 commonsourceibias.n218 0.189894
R812 commonsourceibias.n366 commonsourceibias.n365 0.189894
R813 commonsourceibias.n366 commonsourceibias.n361 0.189894
R814 commonsourceibias.n371 commonsourceibias.n361 0.189894
R815 commonsourceibias.n372 commonsourceibias.n371 0.189894
R816 commonsourceibias.n373 commonsourceibias.n372 0.189894
R817 commonsourceibias.n373 commonsourceibias.n359 0.189894
R818 commonsourceibias.n378 commonsourceibias.n359 0.189894
R819 commonsourceibias.n379 commonsourceibias.n378 0.189894
R820 commonsourceibias.n379 commonsourceibias.n357 0.189894
R821 commonsourceibias.n383 commonsourceibias.n357 0.189894
R822 commonsourceibias.n384 commonsourceibias.n383 0.189894
R823 commonsourceibias.n384 commonsourceibias.n355 0.189894
R824 commonsourceibias.n388 commonsourceibias.n355 0.189894
R825 commonsourceibias.n389 commonsourceibias.n388 0.189894
R826 commonsourceibias.n389 commonsourceibias.n353 0.189894
R827 commonsourceibias.n394 commonsourceibias.n353 0.189894
R828 commonsourceibias.n395 commonsourceibias.n394 0.189894
R829 commonsourceibias.n396 commonsourceibias.n395 0.189894
R830 commonsourceibias.n396 commonsourceibias.n351 0.189894
R831 commonsourceibias.n402 commonsourceibias.n351 0.189894
R832 commonsourceibias.n403 commonsourceibias.n402 0.189894
R833 commonsourceibias.n404 commonsourceibias.n403 0.189894
R834 commonsourceibias.n404 commonsourceibias.n349 0.189894
R835 commonsourceibias.n409 commonsourceibias.n349 0.189894
R836 commonsourceibias.n410 commonsourceibias.n409 0.189894
R837 commonsourceibias.n411 commonsourceibias.n410 0.189894
R838 commonsourceibias.n411 commonsourceibias.n347 0.189894
R839 commonsourceibias.n417 commonsourceibias.n347 0.189894
R840 commonsourceibias.n418 commonsourceibias.n417 0.189894
R841 commonsourceibias.n419 commonsourceibias.n418 0.189894
R842 commonsourceibias.n419 commonsourceibias.n345 0.189894
R843 commonsourceibias.n424 commonsourceibias.n345 0.189894
R844 commonsourceibias.n425 commonsourceibias.n424 0.189894
R845 commonsourceibias.n426 commonsourceibias.n425 0.189894
R846 commonsourceibias.n426 commonsourceibias.n343 0.189894
R847 commonsourceibias.n307 commonsourceibias.n306 0.189894
R848 commonsourceibias.n307 commonsourceibias.n302 0.189894
R849 commonsourceibias.n312 commonsourceibias.n302 0.189894
R850 commonsourceibias.n313 commonsourceibias.n312 0.189894
R851 commonsourceibias.n314 commonsourceibias.n313 0.189894
R852 commonsourceibias.n314 commonsourceibias.n300 0.189894
R853 commonsourceibias.n319 commonsourceibias.n300 0.189894
R854 commonsourceibias.n320 commonsourceibias.n319 0.189894
R855 commonsourceibias.n320 commonsourceibias.n298 0.189894
R856 commonsourceibias.n324 commonsourceibias.n298 0.189894
R857 commonsourceibias.n325 commonsourceibias.n324 0.189894
R858 commonsourceibias.n325 commonsourceibias.n296 0.189894
R859 commonsourceibias.n329 commonsourceibias.n296 0.189894
R860 commonsourceibias.n330 commonsourceibias.n329 0.189894
R861 commonsourceibias.n330 commonsourceibias.n294 0.189894
R862 commonsourceibias.n335 commonsourceibias.n294 0.189894
R863 commonsourceibias.n442 commonsourceibias.n292 0.189894
R864 commonsourceibias.n448 commonsourceibias.n292 0.189894
R865 commonsourceibias.n449 commonsourceibias.n448 0.189894
R866 commonsourceibias.n450 commonsourceibias.n449 0.189894
R867 commonsourceibias.n450 commonsourceibias.n290 0.189894
R868 commonsourceibias.n455 commonsourceibias.n290 0.189894
R869 commonsourceibias.n456 commonsourceibias.n455 0.189894
R870 commonsourceibias.n457 commonsourceibias.n456 0.189894
R871 commonsourceibias.n457 commonsourceibias.n288 0.189894
R872 commonsourceibias.n463 commonsourceibias.n288 0.189894
R873 commonsourceibias.n464 commonsourceibias.n463 0.189894
R874 commonsourceibias.n465 commonsourceibias.n464 0.189894
R875 commonsourceibias.n465 commonsourceibias.n286 0.189894
R876 commonsourceibias.n470 commonsourceibias.n286 0.189894
R877 commonsourceibias.n471 commonsourceibias.n470 0.189894
R878 commonsourceibias.n472 commonsourceibias.n471 0.189894
R879 commonsourceibias.n472 commonsourceibias.n284 0.189894
R880 commonsourceibias.n501 commonsourceibias.n500 0.189894
R881 commonsourceibias.n501 commonsourceibias.n496 0.189894
R882 commonsourceibias.n506 commonsourceibias.n496 0.189894
R883 commonsourceibias.n507 commonsourceibias.n506 0.189894
R884 commonsourceibias.n508 commonsourceibias.n507 0.189894
R885 commonsourceibias.n508 commonsourceibias.n494 0.189894
R886 commonsourceibias.n513 commonsourceibias.n494 0.189894
R887 commonsourceibias.n514 commonsourceibias.n513 0.189894
R888 commonsourceibias.n514 commonsourceibias.n492 0.189894
R889 commonsourceibias.n518 commonsourceibias.n492 0.189894
R890 commonsourceibias.n519 commonsourceibias.n518 0.189894
R891 commonsourceibias.n519 commonsourceibias.n490 0.189894
R892 commonsourceibias.n523 commonsourceibias.n490 0.189894
R893 commonsourceibias.n524 commonsourceibias.n523 0.189894
R894 commonsourceibias.n524 commonsourceibias.n488 0.189894
R895 commonsourceibias.n529 commonsourceibias.n488 0.189894
R896 commonsourceibias.n530 commonsourceibias.n529 0.189894
R897 commonsourceibias.n531 commonsourceibias.n530 0.189894
R898 commonsourceibias.n531 commonsourceibias.n486 0.189894
R899 commonsourceibias.n537 commonsourceibias.n486 0.189894
R900 commonsourceibias.n538 commonsourceibias.n537 0.189894
R901 commonsourceibias.n539 commonsourceibias.n538 0.189894
R902 commonsourceibias.n539 commonsourceibias.n484 0.189894
R903 commonsourceibias.n544 commonsourceibias.n484 0.189894
R904 commonsourceibias.n545 commonsourceibias.n544 0.189894
R905 commonsourceibias.n546 commonsourceibias.n545 0.189894
R906 commonsourceibias.n546 commonsourceibias.n482 0.189894
R907 commonsourceibias.n552 commonsourceibias.n482 0.189894
R908 commonsourceibias.n553 commonsourceibias.n552 0.189894
R909 commonsourceibias.n554 commonsourceibias.n553 0.189894
R910 commonsourceibias.n554 commonsourceibias.n480 0.189894
R911 commonsourceibias.n559 commonsourceibias.n480 0.189894
R912 commonsourceibias.n560 commonsourceibias.n559 0.189894
R913 commonsourceibias.n561 commonsourceibias.n560 0.189894
R914 commonsourceibias.n561 commonsourceibias.n478 0.189894
R915 commonsourceibias.n159 commonsourceibias.n158 0.170955
R916 commonsourceibias.n160 commonsourceibias.n159 0.170955
R917 commonsourceibias.n441 commonsourceibias.n335 0.170955
R918 commonsourceibias.n442 commonsourceibias.n441 0.170955
R919 CSoutput.n19 CSoutput.t188 184.661
R920 CSoutput.n78 CSoutput.n77 165.8
R921 CSoutput.n76 CSoutput.n0 165.8
R922 CSoutput.n75 CSoutput.n74 165.8
R923 CSoutput.n73 CSoutput.n72 165.8
R924 CSoutput.n71 CSoutput.n2 165.8
R925 CSoutput.n69 CSoutput.n68 165.8
R926 CSoutput.n67 CSoutput.n3 165.8
R927 CSoutput.n66 CSoutput.n65 165.8
R928 CSoutput.n63 CSoutput.n4 165.8
R929 CSoutput.n61 CSoutput.n60 165.8
R930 CSoutput.n59 CSoutput.n5 165.8
R931 CSoutput.n58 CSoutput.n57 165.8
R932 CSoutput.n55 CSoutput.n6 165.8
R933 CSoutput.n54 CSoutput.n53 165.8
R934 CSoutput.n52 CSoutput.n51 165.8
R935 CSoutput.n50 CSoutput.n8 165.8
R936 CSoutput.n48 CSoutput.n47 165.8
R937 CSoutput.n46 CSoutput.n9 165.8
R938 CSoutput.n45 CSoutput.n44 165.8
R939 CSoutput.n42 CSoutput.n10 165.8
R940 CSoutput.n41 CSoutput.n40 165.8
R941 CSoutput.n39 CSoutput.n38 165.8
R942 CSoutput.n37 CSoutput.n12 165.8
R943 CSoutput.n35 CSoutput.n34 165.8
R944 CSoutput.n33 CSoutput.n13 165.8
R945 CSoutput.n32 CSoutput.n31 165.8
R946 CSoutput.n29 CSoutput.n14 165.8
R947 CSoutput.n28 CSoutput.n27 165.8
R948 CSoutput.n26 CSoutput.n25 165.8
R949 CSoutput.n24 CSoutput.n16 165.8
R950 CSoutput.n22 CSoutput.n21 165.8
R951 CSoutput.n20 CSoutput.n17 165.8
R952 CSoutput.n77 CSoutput.t190 162.194
R953 CSoutput.n18 CSoutput.t205 120.501
R954 CSoutput.n23 CSoutput.t199 120.501
R955 CSoutput.n15 CSoutput.t196 120.501
R956 CSoutput.n30 CSoutput.t185 120.501
R957 CSoutput.n36 CSoutput.t187 120.501
R958 CSoutput.n11 CSoutput.t197 120.501
R959 CSoutput.n43 CSoutput.t195 120.501
R960 CSoutput.n49 CSoutput.t189 120.501
R961 CSoutput.n7 CSoutput.t200 120.501
R962 CSoutput.n56 CSoutput.t201 120.501
R963 CSoutput.n62 CSoutput.t192 120.501
R964 CSoutput.n64 CSoutput.t202 120.501
R965 CSoutput.n70 CSoutput.t204 120.501
R966 CSoutput.n1 CSoutput.t198 120.501
R967 CSoutput.n330 CSoutput.n328 103.469
R968 CSoutput.n310 CSoutput.n308 103.469
R969 CSoutput.n291 CSoutput.n289 103.469
R970 CSoutput.n120 CSoutput.n118 103.469
R971 CSoutput.n100 CSoutput.n98 103.469
R972 CSoutput.n81 CSoutput.n79 103.469
R973 CSoutput.n344 CSoutput.n343 103.111
R974 CSoutput.n342 CSoutput.n341 103.111
R975 CSoutput.n340 CSoutput.n339 103.111
R976 CSoutput.n338 CSoutput.n337 103.111
R977 CSoutput.n336 CSoutput.n335 103.111
R978 CSoutput.n334 CSoutput.n333 103.111
R979 CSoutput.n332 CSoutput.n331 103.111
R980 CSoutput.n330 CSoutput.n329 103.111
R981 CSoutput.n326 CSoutput.n325 103.111
R982 CSoutput.n324 CSoutput.n323 103.111
R983 CSoutput.n322 CSoutput.n321 103.111
R984 CSoutput.n320 CSoutput.n319 103.111
R985 CSoutput.n318 CSoutput.n317 103.111
R986 CSoutput.n316 CSoutput.n315 103.111
R987 CSoutput.n314 CSoutput.n313 103.111
R988 CSoutput.n312 CSoutput.n311 103.111
R989 CSoutput.n310 CSoutput.n309 103.111
R990 CSoutput.n307 CSoutput.n306 103.111
R991 CSoutput.n305 CSoutput.n304 103.111
R992 CSoutput.n303 CSoutput.n302 103.111
R993 CSoutput.n301 CSoutput.n300 103.111
R994 CSoutput.n299 CSoutput.n298 103.111
R995 CSoutput.n297 CSoutput.n296 103.111
R996 CSoutput.n295 CSoutput.n294 103.111
R997 CSoutput.n293 CSoutput.n292 103.111
R998 CSoutput.n291 CSoutput.n290 103.111
R999 CSoutput.n120 CSoutput.n119 103.111
R1000 CSoutput.n122 CSoutput.n121 103.111
R1001 CSoutput.n124 CSoutput.n123 103.111
R1002 CSoutput.n126 CSoutput.n125 103.111
R1003 CSoutput.n128 CSoutput.n127 103.111
R1004 CSoutput.n130 CSoutput.n129 103.111
R1005 CSoutput.n132 CSoutput.n131 103.111
R1006 CSoutput.n134 CSoutput.n133 103.111
R1007 CSoutput.n136 CSoutput.n135 103.111
R1008 CSoutput.n100 CSoutput.n99 103.111
R1009 CSoutput.n102 CSoutput.n101 103.111
R1010 CSoutput.n104 CSoutput.n103 103.111
R1011 CSoutput.n106 CSoutput.n105 103.111
R1012 CSoutput.n108 CSoutput.n107 103.111
R1013 CSoutput.n110 CSoutput.n109 103.111
R1014 CSoutput.n112 CSoutput.n111 103.111
R1015 CSoutput.n114 CSoutput.n113 103.111
R1016 CSoutput.n116 CSoutput.n115 103.111
R1017 CSoutput.n81 CSoutput.n80 103.111
R1018 CSoutput.n83 CSoutput.n82 103.111
R1019 CSoutput.n85 CSoutput.n84 103.111
R1020 CSoutput.n87 CSoutput.n86 103.111
R1021 CSoutput.n89 CSoutput.n88 103.111
R1022 CSoutput.n91 CSoutput.n90 103.111
R1023 CSoutput.n93 CSoutput.n92 103.111
R1024 CSoutput.n95 CSoutput.n94 103.111
R1025 CSoutput.n97 CSoutput.n96 103.111
R1026 CSoutput.n346 CSoutput.n345 103.111
R1027 CSoutput.n366 CSoutput.n364 81.5057
R1028 CSoutput.n351 CSoutput.n349 81.5057
R1029 CSoutput.n398 CSoutput.n396 81.5057
R1030 CSoutput.n383 CSoutput.n381 81.5057
R1031 CSoutput.n378 CSoutput.n377 80.9324
R1032 CSoutput.n376 CSoutput.n375 80.9324
R1033 CSoutput.n374 CSoutput.n373 80.9324
R1034 CSoutput.n372 CSoutput.n371 80.9324
R1035 CSoutput.n370 CSoutput.n369 80.9324
R1036 CSoutput.n368 CSoutput.n367 80.9324
R1037 CSoutput.n366 CSoutput.n365 80.9324
R1038 CSoutput.n363 CSoutput.n362 80.9324
R1039 CSoutput.n361 CSoutput.n360 80.9324
R1040 CSoutput.n359 CSoutput.n358 80.9324
R1041 CSoutput.n357 CSoutput.n356 80.9324
R1042 CSoutput.n355 CSoutput.n354 80.9324
R1043 CSoutput.n353 CSoutput.n352 80.9324
R1044 CSoutput.n351 CSoutput.n350 80.9324
R1045 CSoutput.n398 CSoutput.n397 80.9324
R1046 CSoutput.n400 CSoutput.n399 80.9324
R1047 CSoutput.n402 CSoutput.n401 80.9324
R1048 CSoutput.n404 CSoutput.n403 80.9324
R1049 CSoutput.n406 CSoutput.n405 80.9324
R1050 CSoutput.n408 CSoutput.n407 80.9324
R1051 CSoutput.n410 CSoutput.n409 80.9324
R1052 CSoutput.n383 CSoutput.n382 80.9324
R1053 CSoutput.n385 CSoutput.n384 80.9324
R1054 CSoutput.n387 CSoutput.n386 80.9324
R1055 CSoutput.n389 CSoutput.n388 80.9324
R1056 CSoutput.n391 CSoutput.n390 80.9324
R1057 CSoutput.n393 CSoutput.n392 80.9324
R1058 CSoutput.n395 CSoutput.n394 80.9324
R1059 CSoutput.n25 CSoutput.n24 48.1486
R1060 CSoutput.n69 CSoutput.n3 48.1486
R1061 CSoutput.n38 CSoutput.n37 48.1486
R1062 CSoutput.n42 CSoutput.n41 48.1486
R1063 CSoutput.n51 CSoutput.n50 48.1486
R1064 CSoutput.n55 CSoutput.n54 48.1486
R1065 CSoutput.n22 CSoutput.n17 46.462
R1066 CSoutput.n72 CSoutput.n71 46.462
R1067 CSoutput.n20 CSoutput.n19 44.9055
R1068 CSoutput.n29 CSoutput.n28 43.7635
R1069 CSoutput.n65 CSoutput.n63 43.7635
R1070 CSoutput.n35 CSoutput.n13 41.7396
R1071 CSoutput.n57 CSoutput.n5 41.7396
R1072 CSoutput.n44 CSoutput.n9 37.0171
R1073 CSoutput.n48 CSoutput.n9 37.0171
R1074 CSoutput.n76 CSoutput.n75 34.9932
R1075 CSoutput.n31 CSoutput.n13 32.2947
R1076 CSoutput.n61 CSoutput.n5 32.2947
R1077 CSoutput.n30 CSoutput.n29 29.6014
R1078 CSoutput.n63 CSoutput.n62 29.6014
R1079 CSoutput.n19 CSoutput.n18 28.4085
R1080 CSoutput.n18 CSoutput.n17 25.1176
R1081 CSoutput.n72 CSoutput.n1 25.1176
R1082 CSoutput.n43 CSoutput.n42 22.0922
R1083 CSoutput.n50 CSoutput.n49 22.0922
R1084 CSoutput.n77 CSoutput.n76 21.8586
R1085 CSoutput.n37 CSoutput.n36 18.9681
R1086 CSoutput.n56 CSoutput.n55 18.9681
R1087 CSoutput.n25 CSoutput.n15 17.6292
R1088 CSoutput.n64 CSoutput.n3 17.6292
R1089 CSoutput.n24 CSoutput.n23 15.844
R1090 CSoutput.n70 CSoutput.n69 15.844
R1091 CSoutput.n38 CSoutput.n11 14.5051
R1092 CSoutput.n54 CSoutput.n7 14.5051
R1093 CSoutput.n413 CSoutput.n78 11.6139
R1094 CSoutput.n41 CSoutput.n11 11.3811
R1095 CSoutput.n51 CSoutput.n7 11.3811
R1096 CSoutput.n23 CSoutput.n22 10.0422
R1097 CSoutput.n71 CSoutput.n70 10.0422
R1098 CSoutput.n327 CSoutput.n307 9.25285
R1099 CSoutput.n117 CSoutput.n97 9.25285
R1100 CSoutput.n379 CSoutput.n363 8.97993
R1101 CSoutput.n411 CSoutput.n395 8.97993
R1102 CSoutput.n380 CSoutput.n348 8.57485
R1103 CSoutput.n28 CSoutput.n15 8.25698
R1104 CSoutput.n65 CSoutput.n64 8.25698
R1105 CSoutput.n380 CSoutput.n379 7.89345
R1106 CSoutput.n412 CSoutput.n411 7.89345
R1107 CSoutput.n348 CSoutput.n347 7.12641
R1108 CSoutput.n138 CSoutput.n137 7.12641
R1109 CSoutput.n36 CSoutput.n35 6.91809
R1110 CSoutput.n57 CSoutput.n56 6.91809
R1111 CSoutput.n379 CSoutput.n378 5.25266
R1112 CSoutput.n411 CSoutput.n410 5.25266
R1113 CSoutput.n347 CSoutput.n346 5.1449
R1114 CSoutput.n327 CSoutput.n326 5.1449
R1115 CSoutput.n137 CSoutput.n136 5.1449
R1116 CSoutput.n117 CSoutput.n116 5.1449
R1117 CSoutput.n413 CSoutput.n138 4.98241
R1118 CSoutput.n229 CSoutput.n182 4.5005
R1119 CSoutput.n198 CSoutput.n182 4.5005
R1120 CSoutput.n193 CSoutput.n177 4.5005
R1121 CSoutput.n193 CSoutput.n179 4.5005
R1122 CSoutput.n193 CSoutput.n176 4.5005
R1123 CSoutput.n193 CSoutput.n180 4.5005
R1124 CSoutput.n193 CSoutput.n175 4.5005
R1125 CSoutput.n193 CSoutput.t203 4.5005
R1126 CSoutput.n193 CSoutput.n174 4.5005
R1127 CSoutput.n193 CSoutput.n181 4.5005
R1128 CSoutput.n193 CSoutput.n182 4.5005
R1129 CSoutput.n191 CSoutput.n177 4.5005
R1130 CSoutput.n191 CSoutput.n179 4.5005
R1131 CSoutput.n191 CSoutput.n176 4.5005
R1132 CSoutput.n191 CSoutput.n180 4.5005
R1133 CSoutput.n191 CSoutput.n175 4.5005
R1134 CSoutput.n191 CSoutput.t203 4.5005
R1135 CSoutput.n191 CSoutput.n174 4.5005
R1136 CSoutput.n191 CSoutput.n181 4.5005
R1137 CSoutput.n191 CSoutput.n182 4.5005
R1138 CSoutput.n190 CSoutput.n177 4.5005
R1139 CSoutput.n190 CSoutput.n179 4.5005
R1140 CSoutput.n190 CSoutput.n176 4.5005
R1141 CSoutput.n190 CSoutput.n180 4.5005
R1142 CSoutput.n190 CSoutput.n175 4.5005
R1143 CSoutput.n190 CSoutput.t203 4.5005
R1144 CSoutput.n190 CSoutput.n174 4.5005
R1145 CSoutput.n190 CSoutput.n181 4.5005
R1146 CSoutput.n190 CSoutput.n182 4.5005
R1147 CSoutput.n275 CSoutput.n177 4.5005
R1148 CSoutput.n275 CSoutput.n179 4.5005
R1149 CSoutput.n275 CSoutput.n176 4.5005
R1150 CSoutput.n275 CSoutput.n180 4.5005
R1151 CSoutput.n275 CSoutput.n175 4.5005
R1152 CSoutput.n275 CSoutput.t203 4.5005
R1153 CSoutput.n275 CSoutput.n174 4.5005
R1154 CSoutput.n275 CSoutput.n181 4.5005
R1155 CSoutput.n275 CSoutput.n182 4.5005
R1156 CSoutput.n273 CSoutput.n177 4.5005
R1157 CSoutput.n273 CSoutput.n179 4.5005
R1158 CSoutput.n273 CSoutput.n176 4.5005
R1159 CSoutput.n273 CSoutput.n180 4.5005
R1160 CSoutput.n273 CSoutput.n175 4.5005
R1161 CSoutput.n273 CSoutput.t203 4.5005
R1162 CSoutput.n273 CSoutput.n174 4.5005
R1163 CSoutput.n273 CSoutput.n181 4.5005
R1164 CSoutput.n271 CSoutput.n177 4.5005
R1165 CSoutput.n271 CSoutput.n179 4.5005
R1166 CSoutput.n271 CSoutput.n176 4.5005
R1167 CSoutput.n271 CSoutput.n180 4.5005
R1168 CSoutput.n271 CSoutput.n175 4.5005
R1169 CSoutput.n271 CSoutput.t203 4.5005
R1170 CSoutput.n271 CSoutput.n174 4.5005
R1171 CSoutput.n271 CSoutput.n181 4.5005
R1172 CSoutput.n201 CSoutput.n177 4.5005
R1173 CSoutput.n201 CSoutput.n179 4.5005
R1174 CSoutput.n201 CSoutput.n176 4.5005
R1175 CSoutput.n201 CSoutput.n180 4.5005
R1176 CSoutput.n201 CSoutput.n175 4.5005
R1177 CSoutput.n201 CSoutput.t203 4.5005
R1178 CSoutput.n201 CSoutput.n174 4.5005
R1179 CSoutput.n201 CSoutput.n181 4.5005
R1180 CSoutput.n201 CSoutput.n182 4.5005
R1181 CSoutput.n200 CSoutput.n177 4.5005
R1182 CSoutput.n200 CSoutput.n179 4.5005
R1183 CSoutput.n200 CSoutput.n176 4.5005
R1184 CSoutput.n200 CSoutput.n180 4.5005
R1185 CSoutput.n200 CSoutput.n175 4.5005
R1186 CSoutput.n200 CSoutput.t203 4.5005
R1187 CSoutput.n200 CSoutput.n174 4.5005
R1188 CSoutput.n200 CSoutput.n181 4.5005
R1189 CSoutput.n200 CSoutput.n182 4.5005
R1190 CSoutput.n204 CSoutput.n177 4.5005
R1191 CSoutput.n204 CSoutput.n179 4.5005
R1192 CSoutput.n204 CSoutput.n176 4.5005
R1193 CSoutput.n204 CSoutput.n180 4.5005
R1194 CSoutput.n204 CSoutput.n175 4.5005
R1195 CSoutput.n204 CSoutput.t203 4.5005
R1196 CSoutput.n204 CSoutput.n174 4.5005
R1197 CSoutput.n204 CSoutput.n181 4.5005
R1198 CSoutput.n204 CSoutput.n182 4.5005
R1199 CSoutput.n203 CSoutput.n177 4.5005
R1200 CSoutput.n203 CSoutput.n179 4.5005
R1201 CSoutput.n203 CSoutput.n176 4.5005
R1202 CSoutput.n203 CSoutput.n180 4.5005
R1203 CSoutput.n203 CSoutput.n175 4.5005
R1204 CSoutput.n203 CSoutput.t203 4.5005
R1205 CSoutput.n203 CSoutput.n174 4.5005
R1206 CSoutput.n203 CSoutput.n181 4.5005
R1207 CSoutput.n203 CSoutput.n182 4.5005
R1208 CSoutput.n186 CSoutput.n177 4.5005
R1209 CSoutput.n186 CSoutput.n179 4.5005
R1210 CSoutput.n186 CSoutput.n176 4.5005
R1211 CSoutput.n186 CSoutput.n180 4.5005
R1212 CSoutput.n186 CSoutput.n175 4.5005
R1213 CSoutput.n186 CSoutput.t203 4.5005
R1214 CSoutput.n186 CSoutput.n174 4.5005
R1215 CSoutput.n186 CSoutput.n181 4.5005
R1216 CSoutput.n186 CSoutput.n182 4.5005
R1217 CSoutput.n278 CSoutput.n177 4.5005
R1218 CSoutput.n278 CSoutput.n179 4.5005
R1219 CSoutput.n278 CSoutput.n176 4.5005
R1220 CSoutput.n278 CSoutput.n180 4.5005
R1221 CSoutput.n278 CSoutput.n175 4.5005
R1222 CSoutput.n278 CSoutput.t203 4.5005
R1223 CSoutput.n278 CSoutput.n174 4.5005
R1224 CSoutput.n278 CSoutput.n181 4.5005
R1225 CSoutput.n278 CSoutput.n182 4.5005
R1226 CSoutput.n265 CSoutput.n236 4.5005
R1227 CSoutput.n265 CSoutput.n242 4.5005
R1228 CSoutput.n223 CSoutput.n212 4.5005
R1229 CSoutput.n223 CSoutput.n214 4.5005
R1230 CSoutput.n223 CSoutput.n211 4.5005
R1231 CSoutput.n223 CSoutput.n215 4.5005
R1232 CSoutput.n223 CSoutput.n210 4.5005
R1233 CSoutput.n223 CSoutput.t184 4.5005
R1234 CSoutput.n223 CSoutput.n209 4.5005
R1235 CSoutput.n223 CSoutput.n216 4.5005
R1236 CSoutput.n265 CSoutput.n223 4.5005
R1237 CSoutput.n244 CSoutput.n212 4.5005
R1238 CSoutput.n244 CSoutput.n214 4.5005
R1239 CSoutput.n244 CSoutput.n211 4.5005
R1240 CSoutput.n244 CSoutput.n215 4.5005
R1241 CSoutput.n244 CSoutput.n210 4.5005
R1242 CSoutput.n244 CSoutput.t184 4.5005
R1243 CSoutput.n244 CSoutput.n209 4.5005
R1244 CSoutput.n244 CSoutput.n216 4.5005
R1245 CSoutput.n265 CSoutput.n244 4.5005
R1246 CSoutput.n222 CSoutput.n212 4.5005
R1247 CSoutput.n222 CSoutput.n214 4.5005
R1248 CSoutput.n222 CSoutput.n211 4.5005
R1249 CSoutput.n222 CSoutput.n215 4.5005
R1250 CSoutput.n222 CSoutput.n210 4.5005
R1251 CSoutput.n222 CSoutput.t184 4.5005
R1252 CSoutput.n222 CSoutput.n209 4.5005
R1253 CSoutput.n222 CSoutput.n216 4.5005
R1254 CSoutput.n265 CSoutput.n222 4.5005
R1255 CSoutput.n246 CSoutput.n212 4.5005
R1256 CSoutput.n246 CSoutput.n214 4.5005
R1257 CSoutput.n246 CSoutput.n211 4.5005
R1258 CSoutput.n246 CSoutput.n215 4.5005
R1259 CSoutput.n246 CSoutput.n210 4.5005
R1260 CSoutput.n246 CSoutput.t184 4.5005
R1261 CSoutput.n246 CSoutput.n209 4.5005
R1262 CSoutput.n246 CSoutput.n216 4.5005
R1263 CSoutput.n265 CSoutput.n246 4.5005
R1264 CSoutput.n212 CSoutput.n207 4.5005
R1265 CSoutput.n214 CSoutput.n207 4.5005
R1266 CSoutput.n211 CSoutput.n207 4.5005
R1267 CSoutput.n215 CSoutput.n207 4.5005
R1268 CSoutput.n210 CSoutput.n207 4.5005
R1269 CSoutput.t184 CSoutput.n207 4.5005
R1270 CSoutput.n209 CSoutput.n207 4.5005
R1271 CSoutput.n216 CSoutput.n207 4.5005
R1272 CSoutput.n268 CSoutput.n212 4.5005
R1273 CSoutput.n268 CSoutput.n214 4.5005
R1274 CSoutput.n268 CSoutput.n211 4.5005
R1275 CSoutput.n268 CSoutput.n215 4.5005
R1276 CSoutput.n268 CSoutput.n210 4.5005
R1277 CSoutput.n268 CSoutput.t184 4.5005
R1278 CSoutput.n268 CSoutput.n209 4.5005
R1279 CSoutput.n268 CSoutput.n216 4.5005
R1280 CSoutput.n266 CSoutput.n212 4.5005
R1281 CSoutput.n266 CSoutput.n214 4.5005
R1282 CSoutput.n266 CSoutput.n211 4.5005
R1283 CSoutput.n266 CSoutput.n215 4.5005
R1284 CSoutput.n266 CSoutput.n210 4.5005
R1285 CSoutput.n266 CSoutput.t184 4.5005
R1286 CSoutput.n266 CSoutput.n209 4.5005
R1287 CSoutput.n266 CSoutput.n216 4.5005
R1288 CSoutput.n266 CSoutput.n265 4.5005
R1289 CSoutput.n248 CSoutput.n212 4.5005
R1290 CSoutput.n248 CSoutput.n214 4.5005
R1291 CSoutput.n248 CSoutput.n211 4.5005
R1292 CSoutput.n248 CSoutput.n215 4.5005
R1293 CSoutput.n248 CSoutput.n210 4.5005
R1294 CSoutput.n248 CSoutput.t184 4.5005
R1295 CSoutput.n248 CSoutput.n209 4.5005
R1296 CSoutput.n248 CSoutput.n216 4.5005
R1297 CSoutput.n265 CSoutput.n248 4.5005
R1298 CSoutput.n220 CSoutput.n212 4.5005
R1299 CSoutput.n220 CSoutput.n214 4.5005
R1300 CSoutput.n220 CSoutput.n211 4.5005
R1301 CSoutput.n220 CSoutput.n215 4.5005
R1302 CSoutput.n220 CSoutput.n210 4.5005
R1303 CSoutput.n220 CSoutput.t184 4.5005
R1304 CSoutput.n220 CSoutput.n209 4.5005
R1305 CSoutput.n220 CSoutput.n216 4.5005
R1306 CSoutput.n265 CSoutput.n220 4.5005
R1307 CSoutput.n250 CSoutput.n212 4.5005
R1308 CSoutput.n250 CSoutput.n214 4.5005
R1309 CSoutput.n250 CSoutput.n211 4.5005
R1310 CSoutput.n250 CSoutput.n215 4.5005
R1311 CSoutput.n250 CSoutput.n210 4.5005
R1312 CSoutput.n250 CSoutput.t184 4.5005
R1313 CSoutput.n250 CSoutput.n209 4.5005
R1314 CSoutput.n250 CSoutput.n216 4.5005
R1315 CSoutput.n265 CSoutput.n250 4.5005
R1316 CSoutput.n219 CSoutput.n212 4.5005
R1317 CSoutput.n219 CSoutput.n214 4.5005
R1318 CSoutput.n219 CSoutput.n211 4.5005
R1319 CSoutput.n219 CSoutput.n215 4.5005
R1320 CSoutput.n219 CSoutput.n210 4.5005
R1321 CSoutput.n219 CSoutput.t184 4.5005
R1322 CSoutput.n219 CSoutput.n209 4.5005
R1323 CSoutput.n219 CSoutput.n216 4.5005
R1324 CSoutput.n265 CSoutput.n219 4.5005
R1325 CSoutput.n264 CSoutput.n212 4.5005
R1326 CSoutput.n264 CSoutput.n214 4.5005
R1327 CSoutput.n264 CSoutput.n211 4.5005
R1328 CSoutput.n264 CSoutput.n215 4.5005
R1329 CSoutput.n264 CSoutput.n210 4.5005
R1330 CSoutput.n264 CSoutput.t184 4.5005
R1331 CSoutput.n264 CSoutput.n209 4.5005
R1332 CSoutput.n264 CSoutput.n216 4.5005
R1333 CSoutput.n265 CSoutput.n264 4.5005
R1334 CSoutput.n263 CSoutput.n148 4.5005
R1335 CSoutput.n164 CSoutput.n148 4.5005
R1336 CSoutput.n159 CSoutput.n143 4.5005
R1337 CSoutput.n159 CSoutput.n145 4.5005
R1338 CSoutput.n159 CSoutput.n142 4.5005
R1339 CSoutput.n159 CSoutput.n146 4.5005
R1340 CSoutput.n159 CSoutput.n141 4.5005
R1341 CSoutput.n159 CSoutput.t193 4.5005
R1342 CSoutput.n159 CSoutput.n140 4.5005
R1343 CSoutput.n159 CSoutput.n147 4.5005
R1344 CSoutput.n159 CSoutput.n148 4.5005
R1345 CSoutput.n157 CSoutput.n143 4.5005
R1346 CSoutput.n157 CSoutput.n145 4.5005
R1347 CSoutput.n157 CSoutput.n142 4.5005
R1348 CSoutput.n157 CSoutput.n146 4.5005
R1349 CSoutput.n157 CSoutput.n141 4.5005
R1350 CSoutput.n157 CSoutput.t193 4.5005
R1351 CSoutput.n157 CSoutput.n140 4.5005
R1352 CSoutput.n157 CSoutput.n147 4.5005
R1353 CSoutput.n157 CSoutput.n148 4.5005
R1354 CSoutput.n156 CSoutput.n143 4.5005
R1355 CSoutput.n156 CSoutput.n145 4.5005
R1356 CSoutput.n156 CSoutput.n142 4.5005
R1357 CSoutput.n156 CSoutput.n146 4.5005
R1358 CSoutput.n156 CSoutput.n141 4.5005
R1359 CSoutput.n156 CSoutput.t193 4.5005
R1360 CSoutput.n156 CSoutput.n140 4.5005
R1361 CSoutput.n156 CSoutput.n147 4.5005
R1362 CSoutput.n156 CSoutput.n148 4.5005
R1363 CSoutput.n285 CSoutput.n143 4.5005
R1364 CSoutput.n285 CSoutput.n145 4.5005
R1365 CSoutput.n285 CSoutput.n142 4.5005
R1366 CSoutput.n285 CSoutput.n146 4.5005
R1367 CSoutput.n285 CSoutput.n141 4.5005
R1368 CSoutput.n285 CSoutput.t193 4.5005
R1369 CSoutput.n285 CSoutput.n140 4.5005
R1370 CSoutput.n285 CSoutput.n147 4.5005
R1371 CSoutput.n285 CSoutput.n148 4.5005
R1372 CSoutput.n283 CSoutput.n143 4.5005
R1373 CSoutput.n283 CSoutput.n145 4.5005
R1374 CSoutput.n283 CSoutput.n142 4.5005
R1375 CSoutput.n283 CSoutput.n146 4.5005
R1376 CSoutput.n283 CSoutput.n141 4.5005
R1377 CSoutput.n283 CSoutput.t193 4.5005
R1378 CSoutput.n283 CSoutput.n140 4.5005
R1379 CSoutput.n283 CSoutput.n147 4.5005
R1380 CSoutput.n281 CSoutput.n143 4.5005
R1381 CSoutput.n281 CSoutput.n145 4.5005
R1382 CSoutput.n281 CSoutput.n142 4.5005
R1383 CSoutput.n281 CSoutput.n146 4.5005
R1384 CSoutput.n281 CSoutput.n141 4.5005
R1385 CSoutput.n281 CSoutput.t193 4.5005
R1386 CSoutput.n281 CSoutput.n140 4.5005
R1387 CSoutput.n281 CSoutput.n147 4.5005
R1388 CSoutput.n167 CSoutput.n143 4.5005
R1389 CSoutput.n167 CSoutput.n145 4.5005
R1390 CSoutput.n167 CSoutput.n142 4.5005
R1391 CSoutput.n167 CSoutput.n146 4.5005
R1392 CSoutput.n167 CSoutput.n141 4.5005
R1393 CSoutput.n167 CSoutput.t193 4.5005
R1394 CSoutput.n167 CSoutput.n140 4.5005
R1395 CSoutput.n167 CSoutput.n147 4.5005
R1396 CSoutput.n167 CSoutput.n148 4.5005
R1397 CSoutput.n166 CSoutput.n143 4.5005
R1398 CSoutput.n166 CSoutput.n145 4.5005
R1399 CSoutput.n166 CSoutput.n142 4.5005
R1400 CSoutput.n166 CSoutput.n146 4.5005
R1401 CSoutput.n166 CSoutput.n141 4.5005
R1402 CSoutput.n166 CSoutput.t193 4.5005
R1403 CSoutput.n166 CSoutput.n140 4.5005
R1404 CSoutput.n166 CSoutput.n147 4.5005
R1405 CSoutput.n166 CSoutput.n148 4.5005
R1406 CSoutput.n170 CSoutput.n143 4.5005
R1407 CSoutput.n170 CSoutput.n145 4.5005
R1408 CSoutput.n170 CSoutput.n142 4.5005
R1409 CSoutput.n170 CSoutput.n146 4.5005
R1410 CSoutput.n170 CSoutput.n141 4.5005
R1411 CSoutput.n170 CSoutput.t193 4.5005
R1412 CSoutput.n170 CSoutput.n140 4.5005
R1413 CSoutput.n170 CSoutput.n147 4.5005
R1414 CSoutput.n170 CSoutput.n148 4.5005
R1415 CSoutput.n169 CSoutput.n143 4.5005
R1416 CSoutput.n169 CSoutput.n145 4.5005
R1417 CSoutput.n169 CSoutput.n142 4.5005
R1418 CSoutput.n169 CSoutput.n146 4.5005
R1419 CSoutput.n169 CSoutput.n141 4.5005
R1420 CSoutput.n169 CSoutput.t193 4.5005
R1421 CSoutput.n169 CSoutput.n140 4.5005
R1422 CSoutput.n169 CSoutput.n147 4.5005
R1423 CSoutput.n169 CSoutput.n148 4.5005
R1424 CSoutput.n152 CSoutput.n143 4.5005
R1425 CSoutput.n152 CSoutput.n145 4.5005
R1426 CSoutput.n152 CSoutput.n142 4.5005
R1427 CSoutput.n152 CSoutput.n146 4.5005
R1428 CSoutput.n152 CSoutput.n141 4.5005
R1429 CSoutput.n152 CSoutput.t193 4.5005
R1430 CSoutput.n152 CSoutput.n140 4.5005
R1431 CSoutput.n152 CSoutput.n147 4.5005
R1432 CSoutput.n152 CSoutput.n148 4.5005
R1433 CSoutput.n288 CSoutput.n143 4.5005
R1434 CSoutput.n288 CSoutput.n145 4.5005
R1435 CSoutput.n288 CSoutput.n142 4.5005
R1436 CSoutput.n288 CSoutput.n146 4.5005
R1437 CSoutput.n288 CSoutput.n141 4.5005
R1438 CSoutput.n288 CSoutput.t193 4.5005
R1439 CSoutput.n288 CSoutput.n140 4.5005
R1440 CSoutput.n288 CSoutput.n147 4.5005
R1441 CSoutput.n288 CSoutput.n148 4.5005
R1442 CSoutput.n347 CSoutput.n327 4.10845
R1443 CSoutput.n137 CSoutput.n117 4.10845
R1444 CSoutput.n345 CSoutput.t58 4.06363
R1445 CSoutput.n345 CSoutput.t26 4.06363
R1446 CSoutput.n343 CSoutput.t98 4.06363
R1447 CSoutput.n343 CSoutput.t179 4.06363
R1448 CSoutput.n341 CSoutput.t97 4.06363
R1449 CSoutput.n341 CSoutput.t59 4.06363
R1450 CSoutput.n339 CSoutput.t43 4.06363
R1451 CSoutput.n339 CSoutput.t95 4.06363
R1452 CSoutput.n337 CSoutput.t84 4.06363
R1453 CSoutput.n337 CSoutput.t7 4.06363
R1454 CSoutput.n335 CSoutput.t166 4.06363
R1455 CSoutput.n335 CSoutput.t181 4.06363
R1456 CSoutput.n333 CSoutput.t4 4.06363
R1457 CSoutput.n333 CSoutput.t72 4.06363
R1458 CSoutput.n331 CSoutput.t167 4.06363
R1459 CSoutput.n331 CSoutput.t169 4.06363
R1460 CSoutput.n329 CSoutput.t33 4.06363
R1461 CSoutput.n329 CSoutput.t87 4.06363
R1462 CSoutput.n328 CSoutput.t78 4.06363
R1463 CSoutput.n328 CSoutput.t40 4.06363
R1464 CSoutput.n325 CSoutput.t1 4.06363
R1465 CSoutput.n325 CSoutput.t66 4.06363
R1466 CSoutput.n323 CSoutput.t8 4.06363
R1467 CSoutput.n323 CSoutput.t172 4.06363
R1468 CSoutput.n321 CSoutput.t94 4.06363
R1469 CSoutput.n321 CSoutput.t42 4.06363
R1470 CSoutput.n319 CSoutput.t17 4.06363
R1471 CSoutput.n319 CSoutput.t13 4.06363
R1472 CSoutput.n317 CSoutput.t44 4.06363
R1473 CSoutput.n317 CSoutput.t56 4.06363
R1474 CSoutput.n315 CSoutput.t54 4.06363
R1475 CSoutput.n315 CSoutput.t73 4.06363
R1476 CSoutput.n313 CSoutput.t34 4.06363
R1477 CSoutput.n313 CSoutput.t171 4.06363
R1478 CSoutput.n311 CSoutput.t74 4.06363
R1479 CSoutput.n311 CSoutput.t2 4.06363
R1480 CSoutput.n309 CSoutput.t173 4.06363
R1481 CSoutput.n309 CSoutput.t88 4.06363
R1482 CSoutput.n308 CSoutput.t27 4.06363
R1483 CSoutput.n308 CSoutput.t164 4.06363
R1484 CSoutput.n306 CSoutput.t29 4.06363
R1485 CSoutput.n306 CSoutput.t79 4.06363
R1486 CSoutput.n304 CSoutput.t91 4.06363
R1487 CSoutput.n304 CSoutput.t80 4.06363
R1488 CSoutput.n302 CSoutput.t11 4.06363
R1489 CSoutput.n302 CSoutput.t24 4.06363
R1490 CSoutput.n300 CSoutput.t93 4.06363
R1491 CSoutput.n300 CSoutput.t68 4.06363
R1492 CSoutput.n298 CSoutput.t52 4.06363
R1493 CSoutput.n298 CSoutput.t50 4.06363
R1494 CSoutput.n296 CSoutput.t61 4.06363
R1495 CSoutput.n296 CSoutput.t92 4.06363
R1496 CSoutput.n294 CSoutput.t46 4.06363
R1497 CSoutput.n294 CSoutput.t86 4.06363
R1498 CSoutput.n292 CSoutput.t178 4.06363
R1499 CSoutput.n292 CSoutput.t23 4.06363
R1500 CSoutput.n290 CSoutput.t16 4.06363
R1501 CSoutput.n290 CSoutput.t81 4.06363
R1502 CSoutput.n289 CSoutput.t45 4.06363
R1503 CSoutput.n289 CSoutput.t77 4.06363
R1504 CSoutput.n118 CSoutput.t38 4.06363
R1505 CSoutput.n118 CSoutput.t71 4.06363
R1506 CSoutput.n119 CSoutput.t6 4.06363
R1507 CSoutput.n119 CSoutput.t21 4.06363
R1508 CSoutput.n121 CSoutput.t182 4.06363
R1509 CSoutput.n121 CSoutput.t168 4.06363
R1510 CSoutput.n123 CSoutput.t25 4.06363
R1511 CSoutput.n123 CSoutput.t57 4.06363
R1512 CSoutput.n125 CSoutput.t19 4.06363
R1513 CSoutput.n125 CSoutput.t163 4.06363
R1514 CSoutput.n127 CSoutput.t39 4.06363
R1515 CSoutput.n127 CSoutput.t53 4.06363
R1516 CSoutput.n129 CSoutput.t5 4.06363
R1517 CSoutput.n129 CSoutput.t20 4.06363
R1518 CSoutput.n131 CSoutput.t96 4.06363
R1519 CSoutput.n131 CSoutput.t14 4.06363
R1520 CSoutput.n133 CSoutput.t174 4.06363
R1521 CSoutput.n133 CSoutput.t10 4.06363
R1522 CSoutput.n135 CSoutput.t69 4.06363
R1523 CSoutput.n135 CSoutput.t48 4.06363
R1524 CSoutput.n98 CSoutput.t0 4.06363
R1525 CSoutput.n98 CSoutput.t36 4.06363
R1526 CSoutput.n99 CSoutput.t175 4.06363
R1527 CSoutput.n99 CSoutput.t177 4.06363
R1528 CSoutput.n101 CSoutput.t37 4.06363
R1529 CSoutput.n101 CSoutput.t75 4.06363
R1530 CSoutput.n103 CSoutput.t41 4.06363
R1531 CSoutput.n103 CSoutput.t85 4.06363
R1532 CSoutput.n105 CSoutput.t176 4.06363
R1533 CSoutput.n105 CSoutput.t22 4.06363
R1534 CSoutput.n107 CSoutput.t18 4.06363
R1535 CSoutput.n107 CSoutput.t65 4.06363
R1536 CSoutput.n109 CSoutput.t30 4.06363
R1537 CSoutput.n109 CSoutput.t31 4.06363
R1538 CSoutput.n111 CSoutput.t51 4.06363
R1539 CSoutput.n111 CSoutput.t63 4.06363
R1540 CSoutput.n113 CSoutput.t64 4.06363
R1541 CSoutput.n113 CSoutput.t83 4.06363
R1542 CSoutput.n115 CSoutput.t67 4.06363
R1543 CSoutput.n115 CSoutput.t76 4.06363
R1544 CSoutput.n79 CSoutput.t15 4.06363
R1545 CSoutput.n79 CSoutput.t55 4.06363
R1546 CSoutput.n80 CSoutput.t170 4.06363
R1547 CSoutput.n80 CSoutput.t28 4.06363
R1548 CSoutput.n82 CSoutput.t9 4.06363
R1549 CSoutput.n82 CSoutput.t70 4.06363
R1550 CSoutput.n84 CSoutput.t47 4.06363
R1551 CSoutput.n84 CSoutput.t62 4.06363
R1552 CSoutput.n86 CSoutput.t90 4.06363
R1553 CSoutput.n86 CSoutput.t165 4.06363
R1554 CSoutput.n88 CSoutput.t89 4.06363
R1555 CSoutput.n88 CSoutput.t183 4.06363
R1556 CSoutput.n90 CSoutput.t60 4.06363
R1557 CSoutput.n90 CSoutput.t12 4.06363
R1558 CSoutput.n92 CSoutput.t82 4.06363
R1559 CSoutput.n92 CSoutput.t32 4.06363
R1560 CSoutput.n94 CSoutput.t180 4.06363
R1561 CSoutput.n94 CSoutput.t35 4.06363
R1562 CSoutput.n96 CSoutput.t3 4.06363
R1563 CSoutput.n96 CSoutput.t49 4.06363
R1564 CSoutput.n44 CSoutput.n43 3.79402
R1565 CSoutput.n49 CSoutput.n48 3.79402
R1566 CSoutput.n413 CSoutput.n412 3.57343
R1567 CSoutput.n412 CSoutput.n380 3.08965
R1568 CSoutput.n348 CSoutput.n138 2.99158
R1569 CSoutput.n377 CSoutput.t159 2.82907
R1570 CSoutput.n377 CSoutput.t157 2.82907
R1571 CSoutput.n375 CSoutput.t113 2.82907
R1572 CSoutput.n375 CSoutput.t130 2.82907
R1573 CSoutput.n373 CSoutput.t100 2.82907
R1574 CSoutput.n373 CSoutput.t103 2.82907
R1575 CSoutput.n371 CSoutput.t158 2.82907
R1576 CSoutput.n371 CSoutput.t138 2.82907
R1577 CSoutput.n369 CSoutput.t150 2.82907
R1578 CSoutput.n369 CSoutput.t154 2.82907
R1579 CSoutput.n367 CSoutput.t109 2.82907
R1580 CSoutput.n367 CSoutput.t117 2.82907
R1581 CSoutput.n365 CSoutput.t161 2.82907
R1582 CSoutput.n365 CSoutput.t151 2.82907
R1583 CSoutput.n364 CSoutput.t153 2.82907
R1584 CSoutput.n364 CSoutput.t132 2.82907
R1585 CSoutput.n362 CSoutput.t99 2.82907
R1586 CSoutput.n362 CSoutput.t107 2.82907
R1587 CSoutput.n360 CSoutput.t131 2.82907
R1588 CSoutput.n360 CSoutput.t142 2.82907
R1589 CSoutput.n358 CSoutput.t110 2.82907
R1590 CSoutput.n358 CSoutput.t152 2.82907
R1591 CSoutput.n356 CSoutput.t108 2.82907
R1592 CSoutput.n356 CSoutput.t116 2.82907
R1593 CSoutput.n354 CSoutput.t160 2.82907
R1594 CSoutput.n354 CSoutput.t135 2.82907
R1595 CSoutput.n352 CSoutput.t118 2.82907
R1596 CSoutput.n352 CSoutput.t126 2.82907
R1597 CSoutput.n350 CSoutput.t102 2.82907
R1598 CSoutput.n350 CSoutput.t104 2.82907
R1599 CSoutput.n349 CSoutput.t134 2.82907
R1600 CSoutput.n349 CSoutput.t144 2.82907
R1601 CSoutput.n396 CSoutput.t139 2.82907
R1602 CSoutput.n396 CSoutput.t121 2.82907
R1603 CSoutput.n397 CSoutput.t101 2.82907
R1604 CSoutput.n397 CSoutput.t148 2.82907
R1605 CSoutput.n399 CSoutput.t124 2.82907
R1606 CSoutput.n399 CSoutput.t115 2.82907
R1607 CSoutput.n401 CSoutput.t122 2.82907
R1608 CSoutput.n401 CSoutput.t127 2.82907
R1609 CSoutput.n403 CSoutput.t143 2.82907
R1610 CSoutput.n403 CSoutput.t136 2.82907
R1611 CSoutput.n405 CSoutput.t111 2.82907
R1612 CSoutput.n405 CSoutput.t105 2.82907
R1613 CSoutput.n407 CSoutput.t128 2.82907
R1614 CSoutput.n407 CSoutput.t119 2.82907
R1615 CSoutput.n409 CSoutput.t133 2.82907
R1616 CSoutput.n409 CSoutput.t155 2.82907
R1617 CSoutput.n381 CSoutput.t149 2.82907
R1618 CSoutput.n381 CSoutput.t140 2.82907
R1619 CSoutput.n382 CSoutput.t112 2.82907
R1620 CSoutput.n382 CSoutput.t106 2.82907
R1621 CSoutput.n384 CSoutput.t162 2.82907
R1622 CSoutput.n384 CSoutput.t125 2.82907
R1623 CSoutput.n386 CSoutput.t141 2.82907
R1624 CSoutput.n386 CSoutput.t146 2.82907
R1625 CSoutput.n388 CSoutput.t123 2.82907
R1626 CSoutput.n388 CSoutput.t114 2.82907
R1627 CSoutput.n390 CSoutput.t120 2.82907
R1628 CSoutput.n390 CSoutput.t156 2.82907
R1629 CSoutput.n392 CSoutput.t147 2.82907
R1630 CSoutput.n392 CSoutput.t129 2.82907
R1631 CSoutput.n394 CSoutput.t145 2.82907
R1632 CSoutput.n394 CSoutput.t137 2.82907
R1633 CSoutput.n75 CSoutput.n1 2.45513
R1634 CSoutput.n229 CSoutput.n227 2.251
R1635 CSoutput.n229 CSoutput.n226 2.251
R1636 CSoutput.n229 CSoutput.n225 2.251
R1637 CSoutput.n229 CSoutput.n224 2.251
R1638 CSoutput.n198 CSoutput.n197 2.251
R1639 CSoutput.n198 CSoutput.n196 2.251
R1640 CSoutput.n198 CSoutput.n195 2.251
R1641 CSoutput.n198 CSoutput.n194 2.251
R1642 CSoutput.n271 CSoutput.n270 2.251
R1643 CSoutput.n236 CSoutput.n234 2.251
R1644 CSoutput.n236 CSoutput.n233 2.251
R1645 CSoutput.n236 CSoutput.n232 2.251
R1646 CSoutput.n254 CSoutput.n236 2.251
R1647 CSoutput.n242 CSoutput.n241 2.251
R1648 CSoutput.n242 CSoutput.n240 2.251
R1649 CSoutput.n242 CSoutput.n239 2.251
R1650 CSoutput.n242 CSoutput.n238 2.251
R1651 CSoutput.n268 CSoutput.n208 2.251
R1652 CSoutput.n263 CSoutput.n261 2.251
R1653 CSoutput.n263 CSoutput.n260 2.251
R1654 CSoutput.n263 CSoutput.n259 2.251
R1655 CSoutput.n263 CSoutput.n258 2.251
R1656 CSoutput.n164 CSoutput.n163 2.251
R1657 CSoutput.n164 CSoutput.n162 2.251
R1658 CSoutput.n164 CSoutput.n161 2.251
R1659 CSoutput.n164 CSoutput.n160 2.251
R1660 CSoutput.n281 CSoutput.n280 2.251
R1661 CSoutput.n198 CSoutput.n178 2.2505
R1662 CSoutput.n193 CSoutput.n178 2.2505
R1663 CSoutput.n191 CSoutput.n178 2.2505
R1664 CSoutput.n190 CSoutput.n178 2.2505
R1665 CSoutput.n275 CSoutput.n178 2.2505
R1666 CSoutput.n273 CSoutput.n178 2.2505
R1667 CSoutput.n271 CSoutput.n178 2.2505
R1668 CSoutput.n201 CSoutput.n178 2.2505
R1669 CSoutput.n200 CSoutput.n178 2.2505
R1670 CSoutput.n204 CSoutput.n178 2.2505
R1671 CSoutput.n203 CSoutput.n178 2.2505
R1672 CSoutput.n186 CSoutput.n178 2.2505
R1673 CSoutput.n278 CSoutput.n178 2.2505
R1674 CSoutput.n278 CSoutput.n277 2.2505
R1675 CSoutput.n242 CSoutput.n213 2.2505
R1676 CSoutput.n223 CSoutput.n213 2.2505
R1677 CSoutput.n244 CSoutput.n213 2.2505
R1678 CSoutput.n222 CSoutput.n213 2.2505
R1679 CSoutput.n246 CSoutput.n213 2.2505
R1680 CSoutput.n213 CSoutput.n207 2.2505
R1681 CSoutput.n268 CSoutput.n213 2.2505
R1682 CSoutput.n266 CSoutput.n213 2.2505
R1683 CSoutput.n248 CSoutput.n213 2.2505
R1684 CSoutput.n220 CSoutput.n213 2.2505
R1685 CSoutput.n250 CSoutput.n213 2.2505
R1686 CSoutput.n219 CSoutput.n213 2.2505
R1687 CSoutput.n264 CSoutput.n213 2.2505
R1688 CSoutput.n264 CSoutput.n217 2.2505
R1689 CSoutput.n164 CSoutput.n144 2.2505
R1690 CSoutput.n159 CSoutput.n144 2.2505
R1691 CSoutput.n157 CSoutput.n144 2.2505
R1692 CSoutput.n156 CSoutput.n144 2.2505
R1693 CSoutput.n285 CSoutput.n144 2.2505
R1694 CSoutput.n283 CSoutput.n144 2.2505
R1695 CSoutput.n281 CSoutput.n144 2.2505
R1696 CSoutput.n167 CSoutput.n144 2.2505
R1697 CSoutput.n166 CSoutput.n144 2.2505
R1698 CSoutput.n170 CSoutput.n144 2.2505
R1699 CSoutput.n169 CSoutput.n144 2.2505
R1700 CSoutput.n152 CSoutput.n144 2.2505
R1701 CSoutput.n288 CSoutput.n144 2.2505
R1702 CSoutput.n288 CSoutput.n287 2.2505
R1703 CSoutput.n206 CSoutput.n199 2.25024
R1704 CSoutput.n206 CSoutput.n192 2.25024
R1705 CSoutput.n274 CSoutput.n206 2.25024
R1706 CSoutput.n206 CSoutput.n202 2.25024
R1707 CSoutput.n206 CSoutput.n205 2.25024
R1708 CSoutput.n206 CSoutput.n173 2.25024
R1709 CSoutput.n256 CSoutput.n253 2.25024
R1710 CSoutput.n256 CSoutput.n252 2.25024
R1711 CSoutput.n256 CSoutput.n251 2.25024
R1712 CSoutput.n256 CSoutput.n218 2.25024
R1713 CSoutput.n256 CSoutput.n255 2.25024
R1714 CSoutput.n257 CSoutput.n256 2.25024
R1715 CSoutput.n172 CSoutput.n165 2.25024
R1716 CSoutput.n172 CSoutput.n158 2.25024
R1717 CSoutput.n284 CSoutput.n172 2.25024
R1718 CSoutput.n172 CSoutput.n168 2.25024
R1719 CSoutput.n172 CSoutput.n171 2.25024
R1720 CSoutput.n172 CSoutput.n139 2.25024
R1721 CSoutput.n273 CSoutput.n183 1.50111
R1722 CSoutput.n221 CSoutput.n207 1.50111
R1723 CSoutput.n283 CSoutput.n149 1.50111
R1724 CSoutput.n229 CSoutput.n228 1.501
R1725 CSoutput.n236 CSoutput.n235 1.501
R1726 CSoutput.n263 CSoutput.n262 1.501
R1727 CSoutput.n277 CSoutput.n188 1.12536
R1728 CSoutput.n277 CSoutput.n189 1.12536
R1729 CSoutput.n277 CSoutput.n276 1.12536
R1730 CSoutput.n237 CSoutput.n217 1.12536
R1731 CSoutput.n243 CSoutput.n217 1.12536
R1732 CSoutput.n245 CSoutput.n217 1.12536
R1733 CSoutput.n287 CSoutput.n154 1.12536
R1734 CSoutput.n287 CSoutput.n155 1.12536
R1735 CSoutput.n287 CSoutput.n286 1.12536
R1736 CSoutput.n277 CSoutput.n184 1.12536
R1737 CSoutput.n277 CSoutput.n185 1.12536
R1738 CSoutput.n277 CSoutput.n187 1.12536
R1739 CSoutput.n267 CSoutput.n217 1.12536
R1740 CSoutput.n247 CSoutput.n217 1.12536
R1741 CSoutput.n249 CSoutput.n217 1.12536
R1742 CSoutput.n287 CSoutput.n150 1.12536
R1743 CSoutput.n287 CSoutput.n151 1.12536
R1744 CSoutput.n287 CSoutput.n153 1.12536
R1745 CSoutput.n31 CSoutput.n30 0.669944
R1746 CSoutput.n62 CSoutput.n61 0.669944
R1747 CSoutput.n368 CSoutput.n366 0.573776
R1748 CSoutput.n370 CSoutput.n368 0.573776
R1749 CSoutput.n372 CSoutput.n370 0.573776
R1750 CSoutput.n374 CSoutput.n372 0.573776
R1751 CSoutput.n376 CSoutput.n374 0.573776
R1752 CSoutput.n378 CSoutput.n376 0.573776
R1753 CSoutput.n353 CSoutput.n351 0.573776
R1754 CSoutput.n355 CSoutput.n353 0.573776
R1755 CSoutput.n357 CSoutput.n355 0.573776
R1756 CSoutput.n359 CSoutput.n357 0.573776
R1757 CSoutput.n361 CSoutput.n359 0.573776
R1758 CSoutput.n363 CSoutput.n361 0.573776
R1759 CSoutput.n410 CSoutput.n408 0.573776
R1760 CSoutput.n408 CSoutput.n406 0.573776
R1761 CSoutput.n406 CSoutput.n404 0.573776
R1762 CSoutput.n404 CSoutput.n402 0.573776
R1763 CSoutput.n402 CSoutput.n400 0.573776
R1764 CSoutput.n400 CSoutput.n398 0.573776
R1765 CSoutput.n395 CSoutput.n393 0.573776
R1766 CSoutput.n393 CSoutput.n391 0.573776
R1767 CSoutput.n391 CSoutput.n389 0.573776
R1768 CSoutput.n389 CSoutput.n387 0.573776
R1769 CSoutput.n387 CSoutput.n385 0.573776
R1770 CSoutput.n385 CSoutput.n383 0.573776
R1771 CSoutput.n413 CSoutput.n288 0.53442
R1772 CSoutput.n332 CSoutput.n330 0.358259
R1773 CSoutput.n334 CSoutput.n332 0.358259
R1774 CSoutput.n336 CSoutput.n334 0.358259
R1775 CSoutput.n338 CSoutput.n336 0.358259
R1776 CSoutput.n340 CSoutput.n338 0.358259
R1777 CSoutput.n342 CSoutput.n340 0.358259
R1778 CSoutput.n344 CSoutput.n342 0.358259
R1779 CSoutput.n346 CSoutput.n344 0.358259
R1780 CSoutput.n312 CSoutput.n310 0.358259
R1781 CSoutput.n314 CSoutput.n312 0.358259
R1782 CSoutput.n316 CSoutput.n314 0.358259
R1783 CSoutput.n318 CSoutput.n316 0.358259
R1784 CSoutput.n320 CSoutput.n318 0.358259
R1785 CSoutput.n322 CSoutput.n320 0.358259
R1786 CSoutput.n324 CSoutput.n322 0.358259
R1787 CSoutput.n326 CSoutput.n324 0.358259
R1788 CSoutput.n293 CSoutput.n291 0.358259
R1789 CSoutput.n295 CSoutput.n293 0.358259
R1790 CSoutput.n297 CSoutput.n295 0.358259
R1791 CSoutput.n299 CSoutput.n297 0.358259
R1792 CSoutput.n301 CSoutput.n299 0.358259
R1793 CSoutput.n303 CSoutput.n301 0.358259
R1794 CSoutput.n305 CSoutput.n303 0.358259
R1795 CSoutput.n307 CSoutput.n305 0.358259
R1796 CSoutput.n136 CSoutput.n134 0.358259
R1797 CSoutput.n134 CSoutput.n132 0.358259
R1798 CSoutput.n132 CSoutput.n130 0.358259
R1799 CSoutput.n130 CSoutput.n128 0.358259
R1800 CSoutput.n128 CSoutput.n126 0.358259
R1801 CSoutput.n126 CSoutput.n124 0.358259
R1802 CSoutput.n124 CSoutput.n122 0.358259
R1803 CSoutput.n122 CSoutput.n120 0.358259
R1804 CSoutput.n116 CSoutput.n114 0.358259
R1805 CSoutput.n114 CSoutput.n112 0.358259
R1806 CSoutput.n112 CSoutput.n110 0.358259
R1807 CSoutput.n110 CSoutput.n108 0.358259
R1808 CSoutput.n108 CSoutput.n106 0.358259
R1809 CSoutput.n106 CSoutput.n104 0.358259
R1810 CSoutput.n104 CSoutput.n102 0.358259
R1811 CSoutput.n102 CSoutput.n100 0.358259
R1812 CSoutput.n97 CSoutput.n95 0.358259
R1813 CSoutput.n95 CSoutput.n93 0.358259
R1814 CSoutput.n93 CSoutput.n91 0.358259
R1815 CSoutput.n91 CSoutput.n89 0.358259
R1816 CSoutput.n89 CSoutput.n87 0.358259
R1817 CSoutput.n87 CSoutput.n85 0.358259
R1818 CSoutput.n85 CSoutput.n83 0.358259
R1819 CSoutput.n83 CSoutput.n81 0.358259
R1820 CSoutput.n21 CSoutput.n20 0.169105
R1821 CSoutput.n21 CSoutput.n16 0.169105
R1822 CSoutput.n26 CSoutput.n16 0.169105
R1823 CSoutput.n27 CSoutput.n26 0.169105
R1824 CSoutput.n27 CSoutput.n14 0.169105
R1825 CSoutput.n32 CSoutput.n14 0.169105
R1826 CSoutput.n33 CSoutput.n32 0.169105
R1827 CSoutput.n34 CSoutput.n33 0.169105
R1828 CSoutput.n34 CSoutput.n12 0.169105
R1829 CSoutput.n39 CSoutput.n12 0.169105
R1830 CSoutput.n40 CSoutput.n39 0.169105
R1831 CSoutput.n40 CSoutput.n10 0.169105
R1832 CSoutput.n45 CSoutput.n10 0.169105
R1833 CSoutput.n46 CSoutput.n45 0.169105
R1834 CSoutput.n47 CSoutput.n46 0.169105
R1835 CSoutput.n47 CSoutput.n8 0.169105
R1836 CSoutput.n52 CSoutput.n8 0.169105
R1837 CSoutput.n53 CSoutput.n52 0.169105
R1838 CSoutput.n53 CSoutput.n6 0.169105
R1839 CSoutput.n58 CSoutput.n6 0.169105
R1840 CSoutput.n59 CSoutput.n58 0.169105
R1841 CSoutput.n60 CSoutput.n59 0.169105
R1842 CSoutput.n60 CSoutput.n4 0.169105
R1843 CSoutput.n66 CSoutput.n4 0.169105
R1844 CSoutput.n67 CSoutput.n66 0.169105
R1845 CSoutput.n68 CSoutput.n67 0.169105
R1846 CSoutput.n68 CSoutput.n2 0.169105
R1847 CSoutput.n73 CSoutput.n2 0.169105
R1848 CSoutput.n74 CSoutput.n73 0.169105
R1849 CSoutput.n74 CSoutput.n0 0.169105
R1850 CSoutput.n78 CSoutput.n0 0.169105
R1851 CSoutput.n231 CSoutput.n230 0.0910737
R1852 CSoutput.n282 CSoutput.n279 0.0723685
R1853 CSoutput.n236 CSoutput.n231 0.0522944
R1854 CSoutput.n279 CSoutput.n278 0.0499135
R1855 CSoutput.n230 CSoutput.n229 0.0499135
R1856 CSoutput.n264 CSoutput.n263 0.0464294
R1857 CSoutput.n272 CSoutput.n269 0.0391444
R1858 CSoutput.n231 CSoutput.t194 0.023435
R1859 CSoutput.n279 CSoutput.t186 0.02262
R1860 CSoutput.n230 CSoutput.t191 0.02262
R1861 CSoutput CSoutput.n413 0.0052
R1862 CSoutput.n201 CSoutput.n184 0.00365111
R1863 CSoutput.n204 CSoutput.n185 0.00365111
R1864 CSoutput.n187 CSoutput.n186 0.00365111
R1865 CSoutput.n229 CSoutput.n188 0.00365111
R1866 CSoutput.n193 CSoutput.n189 0.00365111
R1867 CSoutput.n276 CSoutput.n190 0.00365111
R1868 CSoutput.n267 CSoutput.n266 0.00365111
R1869 CSoutput.n247 CSoutput.n220 0.00365111
R1870 CSoutput.n249 CSoutput.n219 0.00365111
R1871 CSoutput.n237 CSoutput.n236 0.00365111
R1872 CSoutput.n243 CSoutput.n223 0.00365111
R1873 CSoutput.n245 CSoutput.n222 0.00365111
R1874 CSoutput.n167 CSoutput.n150 0.00365111
R1875 CSoutput.n170 CSoutput.n151 0.00365111
R1876 CSoutput.n153 CSoutput.n152 0.00365111
R1877 CSoutput.n263 CSoutput.n154 0.00365111
R1878 CSoutput.n159 CSoutput.n155 0.00365111
R1879 CSoutput.n286 CSoutput.n156 0.00365111
R1880 CSoutput.n198 CSoutput.n188 0.00340054
R1881 CSoutput.n191 CSoutput.n189 0.00340054
R1882 CSoutput.n276 CSoutput.n275 0.00340054
R1883 CSoutput.n271 CSoutput.n184 0.00340054
R1884 CSoutput.n200 CSoutput.n185 0.00340054
R1885 CSoutput.n203 CSoutput.n187 0.00340054
R1886 CSoutput.n242 CSoutput.n237 0.00340054
R1887 CSoutput.n244 CSoutput.n243 0.00340054
R1888 CSoutput.n246 CSoutput.n245 0.00340054
R1889 CSoutput.n268 CSoutput.n267 0.00340054
R1890 CSoutput.n248 CSoutput.n247 0.00340054
R1891 CSoutput.n250 CSoutput.n249 0.00340054
R1892 CSoutput.n164 CSoutput.n154 0.00340054
R1893 CSoutput.n157 CSoutput.n155 0.00340054
R1894 CSoutput.n286 CSoutput.n285 0.00340054
R1895 CSoutput.n281 CSoutput.n150 0.00340054
R1896 CSoutput.n166 CSoutput.n151 0.00340054
R1897 CSoutput.n169 CSoutput.n153 0.00340054
R1898 CSoutput.n199 CSoutput.n193 0.00252698
R1899 CSoutput.n192 CSoutput.n190 0.00252698
R1900 CSoutput.n274 CSoutput.n273 0.00252698
R1901 CSoutput.n202 CSoutput.n200 0.00252698
R1902 CSoutput.n205 CSoutput.n203 0.00252698
R1903 CSoutput.n278 CSoutput.n173 0.00252698
R1904 CSoutput.n199 CSoutput.n198 0.00252698
R1905 CSoutput.n192 CSoutput.n191 0.00252698
R1906 CSoutput.n275 CSoutput.n274 0.00252698
R1907 CSoutput.n202 CSoutput.n201 0.00252698
R1908 CSoutput.n205 CSoutput.n204 0.00252698
R1909 CSoutput.n186 CSoutput.n173 0.00252698
R1910 CSoutput.n253 CSoutput.n223 0.00252698
R1911 CSoutput.n252 CSoutput.n222 0.00252698
R1912 CSoutput.n251 CSoutput.n207 0.00252698
R1913 CSoutput.n248 CSoutput.n218 0.00252698
R1914 CSoutput.n255 CSoutput.n250 0.00252698
R1915 CSoutput.n264 CSoutput.n257 0.00252698
R1916 CSoutput.n253 CSoutput.n242 0.00252698
R1917 CSoutput.n252 CSoutput.n244 0.00252698
R1918 CSoutput.n251 CSoutput.n246 0.00252698
R1919 CSoutput.n266 CSoutput.n218 0.00252698
R1920 CSoutput.n255 CSoutput.n220 0.00252698
R1921 CSoutput.n257 CSoutput.n219 0.00252698
R1922 CSoutput.n165 CSoutput.n159 0.00252698
R1923 CSoutput.n158 CSoutput.n156 0.00252698
R1924 CSoutput.n284 CSoutput.n283 0.00252698
R1925 CSoutput.n168 CSoutput.n166 0.00252698
R1926 CSoutput.n171 CSoutput.n169 0.00252698
R1927 CSoutput.n288 CSoutput.n139 0.00252698
R1928 CSoutput.n165 CSoutput.n164 0.00252698
R1929 CSoutput.n158 CSoutput.n157 0.00252698
R1930 CSoutput.n285 CSoutput.n284 0.00252698
R1931 CSoutput.n168 CSoutput.n167 0.00252698
R1932 CSoutput.n171 CSoutput.n170 0.00252698
R1933 CSoutput.n152 CSoutput.n139 0.00252698
R1934 CSoutput.n273 CSoutput.n272 0.0020275
R1935 CSoutput.n272 CSoutput.n271 0.0020275
R1936 CSoutput.n269 CSoutput.n207 0.0020275
R1937 CSoutput.n269 CSoutput.n268 0.0020275
R1938 CSoutput.n283 CSoutput.n282 0.0020275
R1939 CSoutput.n282 CSoutput.n281 0.0020275
R1940 CSoutput.n183 CSoutput.n182 0.00166668
R1941 CSoutput.n265 CSoutput.n221 0.00166668
R1942 CSoutput.n149 CSoutput.n148 0.00166668
R1943 CSoutput.n287 CSoutput.n149 0.00133328
R1944 CSoutput.n221 CSoutput.n217 0.00133328
R1945 CSoutput.n277 CSoutput.n183 0.00133328
R1946 CSoutput.n280 CSoutput.n172 0.001
R1947 CSoutput.n258 CSoutput.n172 0.001
R1948 CSoutput.n160 CSoutput.n140 0.001
R1949 CSoutput.n259 CSoutput.n140 0.001
R1950 CSoutput.n161 CSoutput.n141 0.001
R1951 CSoutput.n260 CSoutput.n141 0.001
R1952 CSoutput.n162 CSoutput.n142 0.001
R1953 CSoutput.n261 CSoutput.n142 0.001
R1954 CSoutput.n163 CSoutput.n143 0.001
R1955 CSoutput.n262 CSoutput.n143 0.001
R1956 CSoutput.n256 CSoutput.n208 0.001
R1957 CSoutput.n256 CSoutput.n254 0.001
R1958 CSoutput.n238 CSoutput.n209 0.001
R1959 CSoutput.n232 CSoutput.n209 0.001
R1960 CSoutput.n239 CSoutput.n210 0.001
R1961 CSoutput.n233 CSoutput.n210 0.001
R1962 CSoutput.n240 CSoutput.n211 0.001
R1963 CSoutput.n234 CSoutput.n211 0.001
R1964 CSoutput.n241 CSoutput.n212 0.001
R1965 CSoutput.n235 CSoutput.n212 0.001
R1966 CSoutput.n270 CSoutput.n206 0.001
R1967 CSoutput.n224 CSoutput.n206 0.001
R1968 CSoutput.n194 CSoutput.n174 0.001
R1969 CSoutput.n225 CSoutput.n174 0.001
R1970 CSoutput.n195 CSoutput.n175 0.001
R1971 CSoutput.n226 CSoutput.n175 0.001
R1972 CSoutput.n196 CSoutput.n176 0.001
R1973 CSoutput.n227 CSoutput.n176 0.001
R1974 CSoutput.n197 CSoutput.n177 0.001
R1975 CSoutput.n228 CSoutput.n177 0.001
R1976 CSoutput.n228 CSoutput.n178 0.001
R1977 CSoutput.n227 CSoutput.n179 0.001
R1978 CSoutput.n226 CSoutput.n180 0.001
R1979 CSoutput.n225 CSoutput.t203 0.001
R1980 CSoutput.n224 CSoutput.n181 0.001
R1981 CSoutput.n197 CSoutput.n179 0.001
R1982 CSoutput.n196 CSoutput.n180 0.001
R1983 CSoutput.n195 CSoutput.t203 0.001
R1984 CSoutput.n194 CSoutput.n181 0.001
R1985 CSoutput.n270 CSoutput.n182 0.001
R1986 CSoutput.n235 CSoutput.n213 0.001
R1987 CSoutput.n234 CSoutput.n214 0.001
R1988 CSoutput.n233 CSoutput.n215 0.001
R1989 CSoutput.n232 CSoutput.t184 0.001
R1990 CSoutput.n254 CSoutput.n216 0.001
R1991 CSoutput.n241 CSoutput.n214 0.001
R1992 CSoutput.n240 CSoutput.n215 0.001
R1993 CSoutput.n239 CSoutput.t184 0.001
R1994 CSoutput.n238 CSoutput.n216 0.001
R1995 CSoutput.n265 CSoutput.n208 0.001
R1996 CSoutput.n262 CSoutput.n144 0.001
R1997 CSoutput.n261 CSoutput.n145 0.001
R1998 CSoutput.n260 CSoutput.n146 0.001
R1999 CSoutput.n259 CSoutput.t193 0.001
R2000 CSoutput.n258 CSoutput.n147 0.001
R2001 CSoutput.n163 CSoutput.n145 0.001
R2002 CSoutput.n162 CSoutput.n146 0.001
R2003 CSoutput.n161 CSoutput.t193 0.001
R2004 CSoutput.n160 CSoutput.n147 0.001
R2005 CSoutput.n280 CSoutput.n148 0.001
R2006 gnd.n6913 gnd.n506 2229.06
R2007 gnd.n6195 gnd.n6148 939.716
R2008 gnd.n7279 gnd.n103 795.207
R2009 gnd.n7443 gnd.n99 795.207
R2010 gnd.n2873 gnd.n2820 795.207
R2011 gnd.n5693 gnd.n2875 795.207
R2012 gnd.n5909 gnd.n2673 795.207
R2013 gnd.n4592 gnd.n2671 795.207
R2014 gnd.n3810 gnd.n2350 795.207
R2015 gnd.n4035 gnd.n3974 795.207
R2016 gnd.n7441 gnd.n105 775.989
R2017 gnd.n173 gnd.n101 775.989
R2018 gnd.n5696 gnd.n5695 775.989
R2019 gnd.n5768 gnd.n2824 775.989
R2020 gnd.n5911 gnd.n2668 775.989
R2021 gnd.n3726 gnd.n2670 775.989
R2022 gnd.n6070 gnd.n6069 775.989
R2023 gnd.n6146 gnd.n2354 775.989
R2024 gnd.n3599 gnd.n2678 771.183
R2025 gnd.n5780 gnd.n2781 771.183
R2026 gnd.n4623 gnd.n3520 771.183
R2027 gnd.n5452 gnd.n2784 771.183
R2028 gnd.n6210 gnd.n1045 766.379
R2029 gnd.n2321 gnd.n1042 766.379
R2030 gnd.n1613 gnd.n1516 766.379
R2031 gnd.n1609 gnd.n1514 766.379
R2032 gnd.n6194 gnd.n1039 756.769
R2033 gnd.n6205 gnd.n6204 756.769
R2034 gnd.n1706 gnd.n1423 756.769
R2035 gnd.n1704 gnd.n1426 756.769
R2036 gnd.n6421 gnd.n798 703.915
R2037 gnd.n6912 gnd.n507 703.915
R2038 gnd.n7125 gnd.n7124 703.915
R2039 gnd.n3972 gnd.n3811 703.915
R2040 gnd.n6421 gnd.n6420 585
R2041 gnd.n6422 gnd.n6421 585
R2042 gnd.n6419 gnd.n800 585
R2043 gnd.n800 gnd.n799 585
R2044 gnd.n6418 gnd.n6417 585
R2045 gnd.n6417 gnd.n6416 585
R2046 gnd.n805 gnd.n804 585
R2047 gnd.n6415 gnd.n805 585
R2048 gnd.n6413 gnd.n6412 585
R2049 gnd.n6414 gnd.n6413 585
R2050 gnd.n6411 gnd.n807 585
R2051 gnd.n807 gnd.n806 585
R2052 gnd.n6410 gnd.n6409 585
R2053 gnd.n6409 gnd.n6408 585
R2054 gnd.n813 gnd.n812 585
R2055 gnd.n6407 gnd.n813 585
R2056 gnd.n6405 gnd.n6404 585
R2057 gnd.n6406 gnd.n6405 585
R2058 gnd.n6403 gnd.n815 585
R2059 gnd.n815 gnd.n814 585
R2060 gnd.n6402 gnd.n6401 585
R2061 gnd.n6401 gnd.n6400 585
R2062 gnd.n821 gnd.n820 585
R2063 gnd.n6399 gnd.n821 585
R2064 gnd.n6397 gnd.n6396 585
R2065 gnd.n6398 gnd.n6397 585
R2066 gnd.n6395 gnd.n823 585
R2067 gnd.n823 gnd.n822 585
R2068 gnd.n6394 gnd.n6393 585
R2069 gnd.n6393 gnd.n6392 585
R2070 gnd.n829 gnd.n828 585
R2071 gnd.n6391 gnd.n829 585
R2072 gnd.n6389 gnd.n6388 585
R2073 gnd.n6390 gnd.n6389 585
R2074 gnd.n6387 gnd.n831 585
R2075 gnd.n831 gnd.n830 585
R2076 gnd.n6386 gnd.n6385 585
R2077 gnd.n6385 gnd.n6384 585
R2078 gnd.n837 gnd.n836 585
R2079 gnd.n6383 gnd.n837 585
R2080 gnd.n6381 gnd.n6380 585
R2081 gnd.n6382 gnd.n6381 585
R2082 gnd.n6379 gnd.n839 585
R2083 gnd.n839 gnd.n838 585
R2084 gnd.n6378 gnd.n6377 585
R2085 gnd.n6377 gnd.n6376 585
R2086 gnd.n845 gnd.n844 585
R2087 gnd.n6375 gnd.n845 585
R2088 gnd.n6373 gnd.n6372 585
R2089 gnd.n6374 gnd.n6373 585
R2090 gnd.n6371 gnd.n847 585
R2091 gnd.n847 gnd.n846 585
R2092 gnd.n6370 gnd.n6369 585
R2093 gnd.n6369 gnd.n6368 585
R2094 gnd.n853 gnd.n852 585
R2095 gnd.n6367 gnd.n853 585
R2096 gnd.n6365 gnd.n6364 585
R2097 gnd.n6366 gnd.n6365 585
R2098 gnd.n6363 gnd.n855 585
R2099 gnd.n855 gnd.n854 585
R2100 gnd.n6362 gnd.n6361 585
R2101 gnd.n6361 gnd.n6360 585
R2102 gnd.n861 gnd.n860 585
R2103 gnd.n6359 gnd.n861 585
R2104 gnd.n6357 gnd.n6356 585
R2105 gnd.n6358 gnd.n6357 585
R2106 gnd.n6355 gnd.n863 585
R2107 gnd.n863 gnd.n862 585
R2108 gnd.n6354 gnd.n6353 585
R2109 gnd.n6353 gnd.n6352 585
R2110 gnd.n869 gnd.n868 585
R2111 gnd.n6351 gnd.n869 585
R2112 gnd.n6349 gnd.n6348 585
R2113 gnd.n6350 gnd.n6349 585
R2114 gnd.n6347 gnd.n871 585
R2115 gnd.n871 gnd.n870 585
R2116 gnd.n6346 gnd.n6345 585
R2117 gnd.n6345 gnd.n6344 585
R2118 gnd.n877 gnd.n876 585
R2119 gnd.n6343 gnd.n877 585
R2120 gnd.n6341 gnd.n6340 585
R2121 gnd.n6342 gnd.n6341 585
R2122 gnd.n6339 gnd.n879 585
R2123 gnd.n879 gnd.n878 585
R2124 gnd.n6338 gnd.n6337 585
R2125 gnd.n6337 gnd.n6336 585
R2126 gnd.n885 gnd.n884 585
R2127 gnd.n6335 gnd.n885 585
R2128 gnd.n6333 gnd.n6332 585
R2129 gnd.n6334 gnd.n6333 585
R2130 gnd.n6331 gnd.n887 585
R2131 gnd.n887 gnd.n886 585
R2132 gnd.n6330 gnd.n6329 585
R2133 gnd.n6329 gnd.n6328 585
R2134 gnd.n893 gnd.n892 585
R2135 gnd.n6327 gnd.n893 585
R2136 gnd.n6325 gnd.n6324 585
R2137 gnd.n6326 gnd.n6325 585
R2138 gnd.n6323 gnd.n895 585
R2139 gnd.n895 gnd.n894 585
R2140 gnd.n6322 gnd.n6321 585
R2141 gnd.n6321 gnd.n6320 585
R2142 gnd.n901 gnd.n900 585
R2143 gnd.n6319 gnd.n901 585
R2144 gnd.n6317 gnd.n6316 585
R2145 gnd.n6318 gnd.n6317 585
R2146 gnd.n6315 gnd.n903 585
R2147 gnd.n903 gnd.n902 585
R2148 gnd.n6314 gnd.n6313 585
R2149 gnd.n6313 gnd.n6312 585
R2150 gnd.n909 gnd.n908 585
R2151 gnd.n6311 gnd.n909 585
R2152 gnd.n6309 gnd.n6308 585
R2153 gnd.n6310 gnd.n6309 585
R2154 gnd.n6307 gnd.n911 585
R2155 gnd.n911 gnd.n910 585
R2156 gnd.n6306 gnd.n6305 585
R2157 gnd.n6305 gnd.n6304 585
R2158 gnd.n917 gnd.n916 585
R2159 gnd.n6303 gnd.n917 585
R2160 gnd.n6301 gnd.n6300 585
R2161 gnd.n6302 gnd.n6301 585
R2162 gnd.n6299 gnd.n919 585
R2163 gnd.n919 gnd.n918 585
R2164 gnd.n6298 gnd.n6297 585
R2165 gnd.n6297 gnd.n6296 585
R2166 gnd.n925 gnd.n924 585
R2167 gnd.n6295 gnd.n925 585
R2168 gnd.n6293 gnd.n6292 585
R2169 gnd.n6294 gnd.n6293 585
R2170 gnd.n6291 gnd.n927 585
R2171 gnd.n927 gnd.n926 585
R2172 gnd.n6290 gnd.n6289 585
R2173 gnd.n6289 gnd.n6288 585
R2174 gnd.n933 gnd.n932 585
R2175 gnd.n6287 gnd.n933 585
R2176 gnd.n6285 gnd.n6284 585
R2177 gnd.n6286 gnd.n6285 585
R2178 gnd.n6283 gnd.n935 585
R2179 gnd.n935 gnd.n934 585
R2180 gnd.n6282 gnd.n6281 585
R2181 gnd.n6281 gnd.n6280 585
R2182 gnd.n941 gnd.n940 585
R2183 gnd.n6279 gnd.n941 585
R2184 gnd.n6277 gnd.n6276 585
R2185 gnd.n6278 gnd.n6277 585
R2186 gnd.n6275 gnd.n943 585
R2187 gnd.n943 gnd.n942 585
R2188 gnd.n6274 gnd.n6273 585
R2189 gnd.n6273 gnd.n6272 585
R2190 gnd.n949 gnd.n948 585
R2191 gnd.n6271 gnd.n949 585
R2192 gnd.n6269 gnd.n6268 585
R2193 gnd.n6270 gnd.n6269 585
R2194 gnd.n6267 gnd.n951 585
R2195 gnd.n951 gnd.n950 585
R2196 gnd.n6266 gnd.n6265 585
R2197 gnd.n6265 gnd.n6264 585
R2198 gnd.n957 gnd.n956 585
R2199 gnd.n6263 gnd.n957 585
R2200 gnd.n6261 gnd.n6260 585
R2201 gnd.n6262 gnd.n6261 585
R2202 gnd.n6259 gnd.n959 585
R2203 gnd.n959 gnd.n958 585
R2204 gnd.n6258 gnd.n6257 585
R2205 gnd.n6257 gnd.n6256 585
R2206 gnd.n965 gnd.n964 585
R2207 gnd.n6255 gnd.n965 585
R2208 gnd.n798 gnd.n797 585
R2209 gnd.n6423 gnd.n798 585
R2210 gnd.n6426 gnd.n6425 585
R2211 gnd.n6425 gnd.n6424 585
R2212 gnd.n795 gnd.n794 585
R2213 gnd.n794 gnd.n793 585
R2214 gnd.n6431 gnd.n6430 585
R2215 gnd.n6432 gnd.n6431 585
R2216 gnd.n792 gnd.n791 585
R2217 gnd.n6433 gnd.n792 585
R2218 gnd.n6436 gnd.n6435 585
R2219 gnd.n6435 gnd.n6434 585
R2220 gnd.n789 gnd.n788 585
R2221 gnd.n788 gnd.n787 585
R2222 gnd.n6441 gnd.n6440 585
R2223 gnd.n6442 gnd.n6441 585
R2224 gnd.n786 gnd.n785 585
R2225 gnd.n6443 gnd.n786 585
R2226 gnd.n6446 gnd.n6445 585
R2227 gnd.n6445 gnd.n6444 585
R2228 gnd.n783 gnd.n782 585
R2229 gnd.n782 gnd.n781 585
R2230 gnd.n6451 gnd.n6450 585
R2231 gnd.n6452 gnd.n6451 585
R2232 gnd.n780 gnd.n779 585
R2233 gnd.n6453 gnd.n780 585
R2234 gnd.n6456 gnd.n6455 585
R2235 gnd.n6455 gnd.n6454 585
R2236 gnd.n777 gnd.n776 585
R2237 gnd.n776 gnd.n775 585
R2238 gnd.n6461 gnd.n6460 585
R2239 gnd.n6462 gnd.n6461 585
R2240 gnd.n774 gnd.n773 585
R2241 gnd.n6463 gnd.n774 585
R2242 gnd.n6466 gnd.n6465 585
R2243 gnd.n6465 gnd.n6464 585
R2244 gnd.n771 gnd.n770 585
R2245 gnd.n770 gnd.n769 585
R2246 gnd.n6471 gnd.n6470 585
R2247 gnd.n6472 gnd.n6471 585
R2248 gnd.n768 gnd.n767 585
R2249 gnd.n6473 gnd.n768 585
R2250 gnd.n6476 gnd.n6475 585
R2251 gnd.n6475 gnd.n6474 585
R2252 gnd.n765 gnd.n764 585
R2253 gnd.n764 gnd.n763 585
R2254 gnd.n6481 gnd.n6480 585
R2255 gnd.n6482 gnd.n6481 585
R2256 gnd.n762 gnd.n761 585
R2257 gnd.n6483 gnd.n762 585
R2258 gnd.n6486 gnd.n6485 585
R2259 gnd.n6485 gnd.n6484 585
R2260 gnd.n759 gnd.n758 585
R2261 gnd.n758 gnd.n757 585
R2262 gnd.n6491 gnd.n6490 585
R2263 gnd.n6492 gnd.n6491 585
R2264 gnd.n756 gnd.n755 585
R2265 gnd.n6493 gnd.n756 585
R2266 gnd.n6496 gnd.n6495 585
R2267 gnd.n6495 gnd.n6494 585
R2268 gnd.n753 gnd.n752 585
R2269 gnd.n752 gnd.n751 585
R2270 gnd.n6501 gnd.n6500 585
R2271 gnd.n6502 gnd.n6501 585
R2272 gnd.n750 gnd.n749 585
R2273 gnd.n6503 gnd.n750 585
R2274 gnd.n6506 gnd.n6505 585
R2275 gnd.n6505 gnd.n6504 585
R2276 gnd.n747 gnd.n746 585
R2277 gnd.n746 gnd.n745 585
R2278 gnd.n6511 gnd.n6510 585
R2279 gnd.n6512 gnd.n6511 585
R2280 gnd.n744 gnd.n743 585
R2281 gnd.n6513 gnd.n744 585
R2282 gnd.n6516 gnd.n6515 585
R2283 gnd.n6515 gnd.n6514 585
R2284 gnd.n741 gnd.n740 585
R2285 gnd.n740 gnd.n739 585
R2286 gnd.n6521 gnd.n6520 585
R2287 gnd.n6522 gnd.n6521 585
R2288 gnd.n738 gnd.n737 585
R2289 gnd.n6523 gnd.n738 585
R2290 gnd.n6526 gnd.n6525 585
R2291 gnd.n6525 gnd.n6524 585
R2292 gnd.n735 gnd.n734 585
R2293 gnd.n734 gnd.n733 585
R2294 gnd.n6531 gnd.n6530 585
R2295 gnd.n6532 gnd.n6531 585
R2296 gnd.n732 gnd.n731 585
R2297 gnd.n6533 gnd.n732 585
R2298 gnd.n6536 gnd.n6535 585
R2299 gnd.n6535 gnd.n6534 585
R2300 gnd.n729 gnd.n728 585
R2301 gnd.n728 gnd.n727 585
R2302 gnd.n6541 gnd.n6540 585
R2303 gnd.n6542 gnd.n6541 585
R2304 gnd.n726 gnd.n725 585
R2305 gnd.n6543 gnd.n726 585
R2306 gnd.n6546 gnd.n6545 585
R2307 gnd.n6545 gnd.n6544 585
R2308 gnd.n723 gnd.n722 585
R2309 gnd.n722 gnd.n721 585
R2310 gnd.n6551 gnd.n6550 585
R2311 gnd.n6552 gnd.n6551 585
R2312 gnd.n720 gnd.n719 585
R2313 gnd.n6553 gnd.n720 585
R2314 gnd.n6556 gnd.n6555 585
R2315 gnd.n6555 gnd.n6554 585
R2316 gnd.n717 gnd.n716 585
R2317 gnd.n716 gnd.n715 585
R2318 gnd.n6561 gnd.n6560 585
R2319 gnd.n6562 gnd.n6561 585
R2320 gnd.n714 gnd.n713 585
R2321 gnd.n6563 gnd.n714 585
R2322 gnd.n6566 gnd.n6565 585
R2323 gnd.n6565 gnd.n6564 585
R2324 gnd.n711 gnd.n710 585
R2325 gnd.n710 gnd.n709 585
R2326 gnd.n6571 gnd.n6570 585
R2327 gnd.n6572 gnd.n6571 585
R2328 gnd.n708 gnd.n707 585
R2329 gnd.n6573 gnd.n708 585
R2330 gnd.n6576 gnd.n6575 585
R2331 gnd.n6575 gnd.n6574 585
R2332 gnd.n705 gnd.n704 585
R2333 gnd.n704 gnd.n703 585
R2334 gnd.n6581 gnd.n6580 585
R2335 gnd.n6582 gnd.n6581 585
R2336 gnd.n702 gnd.n701 585
R2337 gnd.n6583 gnd.n702 585
R2338 gnd.n6586 gnd.n6585 585
R2339 gnd.n6585 gnd.n6584 585
R2340 gnd.n699 gnd.n698 585
R2341 gnd.n698 gnd.n697 585
R2342 gnd.n6591 gnd.n6590 585
R2343 gnd.n6592 gnd.n6591 585
R2344 gnd.n696 gnd.n695 585
R2345 gnd.n6593 gnd.n696 585
R2346 gnd.n6596 gnd.n6595 585
R2347 gnd.n6595 gnd.n6594 585
R2348 gnd.n693 gnd.n692 585
R2349 gnd.n692 gnd.n691 585
R2350 gnd.n6601 gnd.n6600 585
R2351 gnd.n6602 gnd.n6601 585
R2352 gnd.n690 gnd.n689 585
R2353 gnd.n6603 gnd.n690 585
R2354 gnd.n6606 gnd.n6605 585
R2355 gnd.n6605 gnd.n6604 585
R2356 gnd.n687 gnd.n686 585
R2357 gnd.n686 gnd.n685 585
R2358 gnd.n6611 gnd.n6610 585
R2359 gnd.n6612 gnd.n6611 585
R2360 gnd.n684 gnd.n683 585
R2361 gnd.n6613 gnd.n684 585
R2362 gnd.n6616 gnd.n6615 585
R2363 gnd.n6615 gnd.n6614 585
R2364 gnd.n681 gnd.n680 585
R2365 gnd.n680 gnd.n679 585
R2366 gnd.n6621 gnd.n6620 585
R2367 gnd.n6622 gnd.n6621 585
R2368 gnd.n678 gnd.n677 585
R2369 gnd.n6623 gnd.n678 585
R2370 gnd.n6626 gnd.n6625 585
R2371 gnd.n6625 gnd.n6624 585
R2372 gnd.n675 gnd.n674 585
R2373 gnd.n674 gnd.n673 585
R2374 gnd.n6631 gnd.n6630 585
R2375 gnd.n6632 gnd.n6631 585
R2376 gnd.n672 gnd.n671 585
R2377 gnd.n6633 gnd.n672 585
R2378 gnd.n6636 gnd.n6635 585
R2379 gnd.n6635 gnd.n6634 585
R2380 gnd.n669 gnd.n668 585
R2381 gnd.n668 gnd.n667 585
R2382 gnd.n6641 gnd.n6640 585
R2383 gnd.n6642 gnd.n6641 585
R2384 gnd.n666 gnd.n665 585
R2385 gnd.n6643 gnd.n666 585
R2386 gnd.n6646 gnd.n6645 585
R2387 gnd.n6645 gnd.n6644 585
R2388 gnd.n663 gnd.n662 585
R2389 gnd.n662 gnd.n661 585
R2390 gnd.n6651 gnd.n6650 585
R2391 gnd.n6652 gnd.n6651 585
R2392 gnd.n660 gnd.n659 585
R2393 gnd.n6653 gnd.n660 585
R2394 gnd.n6656 gnd.n6655 585
R2395 gnd.n6655 gnd.n6654 585
R2396 gnd.n657 gnd.n656 585
R2397 gnd.n656 gnd.n655 585
R2398 gnd.n6661 gnd.n6660 585
R2399 gnd.n6662 gnd.n6661 585
R2400 gnd.n654 gnd.n653 585
R2401 gnd.n6663 gnd.n654 585
R2402 gnd.n6666 gnd.n6665 585
R2403 gnd.n6665 gnd.n6664 585
R2404 gnd.n651 gnd.n650 585
R2405 gnd.n650 gnd.n649 585
R2406 gnd.n6671 gnd.n6670 585
R2407 gnd.n6672 gnd.n6671 585
R2408 gnd.n648 gnd.n647 585
R2409 gnd.n6673 gnd.n648 585
R2410 gnd.n6676 gnd.n6675 585
R2411 gnd.n6675 gnd.n6674 585
R2412 gnd.n645 gnd.n644 585
R2413 gnd.n644 gnd.n643 585
R2414 gnd.n6681 gnd.n6680 585
R2415 gnd.n6682 gnd.n6681 585
R2416 gnd.n642 gnd.n641 585
R2417 gnd.n6683 gnd.n642 585
R2418 gnd.n6686 gnd.n6685 585
R2419 gnd.n6685 gnd.n6684 585
R2420 gnd.n639 gnd.n638 585
R2421 gnd.n638 gnd.n637 585
R2422 gnd.n6691 gnd.n6690 585
R2423 gnd.n6692 gnd.n6691 585
R2424 gnd.n636 gnd.n635 585
R2425 gnd.n6693 gnd.n636 585
R2426 gnd.n6696 gnd.n6695 585
R2427 gnd.n6695 gnd.n6694 585
R2428 gnd.n633 gnd.n632 585
R2429 gnd.n632 gnd.n631 585
R2430 gnd.n6701 gnd.n6700 585
R2431 gnd.n6702 gnd.n6701 585
R2432 gnd.n630 gnd.n629 585
R2433 gnd.n6703 gnd.n630 585
R2434 gnd.n6706 gnd.n6705 585
R2435 gnd.n6705 gnd.n6704 585
R2436 gnd.n627 gnd.n626 585
R2437 gnd.n626 gnd.n625 585
R2438 gnd.n6711 gnd.n6710 585
R2439 gnd.n6712 gnd.n6711 585
R2440 gnd.n624 gnd.n623 585
R2441 gnd.n6713 gnd.n624 585
R2442 gnd.n6716 gnd.n6715 585
R2443 gnd.n6715 gnd.n6714 585
R2444 gnd.n621 gnd.n620 585
R2445 gnd.n620 gnd.n619 585
R2446 gnd.n6721 gnd.n6720 585
R2447 gnd.n6722 gnd.n6721 585
R2448 gnd.n618 gnd.n617 585
R2449 gnd.n6723 gnd.n618 585
R2450 gnd.n6726 gnd.n6725 585
R2451 gnd.n6725 gnd.n6724 585
R2452 gnd.n615 gnd.n614 585
R2453 gnd.n614 gnd.n613 585
R2454 gnd.n6731 gnd.n6730 585
R2455 gnd.n6732 gnd.n6731 585
R2456 gnd.n612 gnd.n611 585
R2457 gnd.n6733 gnd.n612 585
R2458 gnd.n6736 gnd.n6735 585
R2459 gnd.n6735 gnd.n6734 585
R2460 gnd.n609 gnd.n608 585
R2461 gnd.n608 gnd.n607 585
R2462 gnd.n6741 gnd.n6740 585
R2463 gnd.n6742 gnd.n6741 585
R2464 gnd.n606 gnd.n605 585
R2465 gnd.n6743 gnd.n606 585
R2466 gnd.n6746 gnd.n6745 585
R2467 gnd.n6745 gnd.n6744 585
R2468 gnd.n603 gnd.n602 585
R2469 gnd.n602 gnd.n601 585
R2470 gnd.n6751 gnd.n6750 585
R2471 gnd.n6752 gnd.n6751 585
R2472 gnd.n600 gnd.n599 585
R2473 gnd.n6753 gnd.n600 585
R2474 gnd.n6756 gnd.n6755 585
R2475 gnd.n6755 gnd.n6754 585
R2476 gnd.n597 gnd.n596 585
R2477 gnd.n596 gnd.n595 585
R2478 gnd.n6761 gnd.n6760 585
R2479 gnd.n6762 gnd.n6761 585
R2480 gnd.n594 gnd.n593 585
R2481 gnd.n6763 gnd.n594 585
R2482 gnd.n6766 gnd.n6765 585
R2483 gnd.n6765 gnd.n6764 585
R2484 gnd.n591 gnd.n590 585
R2485 gnd.n590 gnd.n589 585
R2486 gnd.n6771 gnd.n6770 585
R2487 gnd.n6772 gnd.n6771 585
R2488 gnd.n588 gnd.n587 585
R2489 gnd.n6773 gnd.n588 585
R2490 gnd.n6776 gnd.n6775 585
R2491 gnd.n6775 gnd.n6774 585
R2492 gnd.n585 gnd.n584 585
R2493 gnd.n584 gnd.n583 585
R2494 gnd.n6781 gnd.n6780 585
R2495 gnd.n6782 gnd.n6781 585
R2496 gnd.n582 gnd.n581 585
R2497 gnd.n6783 gnd.n582 585
R2498 gnd.n6786 gnd.n6785 585
R2499 gnd.n6785 gnd.n6784 585
R2500 gnd.n579 gnd.n578 585
R2501 gnd.n578 gnd.n577 585
R2502 gnd.n6791 gnd.n6790 585
R2503 gnd.n6792 gnd.n6791 585
R2504 gnd.n576 gnd.n575 585
R2505 gnd.n6793 gnd.n576 585
R2506 gnd.n6796 gnd.n6795 585
R2507 gnd.n6795 gnd.n6794 585
R2508 gnd.n573 gnd.n572 585
R2509 gnd.n572 gnd.n571 585
R2510 gnd.n6801 gnd.n6800 585
R2511 gnd.n6802 gnd.n6801 585
R2512 gnd.n570 gnd.n569 585
R2513 gnd.n6803 gnd.n570 585
R2514 gnd.n6806 gnd.n6805 585
R2515 gnd.n6805 gnd.n6804 585
R2516 gnd.n567 gnd.n566 585
R2517 gnd.n566 gnd.n565 585
R2518 gnd.n6811 gnd.n6810 585
R2519 gnd.n6812 gnd.n6811 585
R2520 gnd.n564 gnd.n563 585
R2521 gnd.n6813 gnd.n564 585
R2522 gnd.n6816 gnd.n6815 585
R2523 gnd.n6815 gnd.n6814 585
R2524 gnd.n561 gnd.n560 585
R2525 gnd.n560 gnd.n559 585
R2526 gnd.n6821 gnd.n6820 585
R2527 gnd.n6822 gnd.n6821 585
R2528 gnd.n558 gnd.n557 585
R2529 gnd.n6823 gnd.n558 585
R2530 gnd.n6826 gnd.n6825 585
R2531 gnd.n6825 gnd.n6824 585
R2532 gnd.n555 gnd.n554 585
R2533 gnd.n554 gnd.n553 585
R2534 gnd.n6831 gnd.n6830 585
R2535 gnd.n6832 gnd.n6831 585
R2536 gnd.n552 gnd.n551 585
R2537 gnd.n6833 gnd.n552 585
R2538 gnd.n6836 gnd.n6835 585
R2539 gnd.n6835 gnd.n6834 585
R2540 gnd.n549 gnd.n548 585
R2541 gnd.n548 gnd.n547 585
R2542 gnd.n6841 gnd.n6840 585
R2543 gnd.n6842 gnd.n6841 585
R2544 gnd.n546 gnd.n545 585
R2545 gnd.n6843 gnd.n546 585
R2546 gnd.n6846 gnd.n6845 585
R2547 gnd.n6845 gnd.n6844 585
R2548 gnd.n543 gnd.n542 585
R2549 gnd.n542 gnd.n541 585
R2550 gnd.n6851 gnd.n6850 585
R2551 gnd.n6852 gnd.n6851 585
R2552 gnd.n540 gnd.n539 585
R2553 gnd.n6853 gnd.n540 585
R2554 gnd.n6856 gnd.n6855 585
R2555 gnd.n6855 gnd.n6854 585
R2556 gnd.n537 gnd.n536 585
R2557 gnd.n536 gnd.n535 585
R2558 gnd.n6861 gnd.n6860 585
R2559 gnd.n6862 gnd.n6861 585
R2560 gnd.n534 gnd.n533 585
R2561 gnd.n6863 gnd.n534 585
R2562 gnd.n6866 gnd.n6865 585
R2563 gnd.n6865 gnd.n6864 585
R2564 gnd.n531 gnd.n530 585
R2565 gnd.n530 gnd.n529 585
R2566 gnd.n6871 gnd.n6870 585
R2567 gnd.n6872 gnd.n6871 585
R2568 gnd.n528 gnd.n527 585
R2569 gnd.n6873 gnd.n528 585
R2570 gnd.n6876 gnd.n6875 585
R2571 gnd.n6875 gnd.n6874 585
R2572 gnd.n525 gnd.n524 585
R2573 gnd.n524 gnd.n523 585
R2574 gnd.n6881 gnd.n6880 585
R2575 gnd.n6882 gnd.n6881 585
R2576 gnd.n522 gnd.n521 585
R2577 gnd.n6883 gnd.n522 585
R2578 gnd.n6886 gnd.n6885 585
R2579 gnd.n6885 gnd.n6884 585
R2580 gnd.n519 gnd.n518 585
R2581 gnd.n518 gnd.n517 585
R2582 gnd.n6891 gnd.n6890 585
R2583 gnd.n6892 gnd.n6891 585
R2584 gnd.n516 gnd.n515 585
R2585 gnd.n6893 gnd.n516 585
R2586 gnd.n6896 gnd.n6895 585
R2587 gnd.n6895 gnd.n6894 585
R2588 gnd.n513 gnd.n512 585
R2589 gnd.n512 gnd.n511 585
R2590 gnd.n6902 gnd.n6901 585
R2591 gnd.n6903 gnd.n6902 585
R2592 gnd.n510 gnd.n509 585
R2593 gnd.n6904 gnd.n510 585
R2594 gnd.n6907 gnd.n6906 585
R2595 gnd.n6906 gnd.n6905 585
R2596 gnd.n6908 gnd.n507 585
R2597 gnd.n507 gnd.n506 585
R2598 gnd.n382 gnd.n381 585
R2599 gnd.n7115 gnd.n381 585
R2600 gnd.n7118 gnd.n7117 585
R2601 gnd.n7117 gnd.n7116 585
R2602 gnd.n385 gnd.n384 585
R2603 gnd.n7114 gnd.n385 585
R2604 gnd.n7112 gnd.n7111 585
R2605 gnd.n7113 gnd.n7112 585
R2606 gnd.n388 gnd.n387 585
R2607 gnd.n387 gnd.n386 585
R2608 gnd.n7107 gnd.n7106 585
R2609 gnd.n7106 gnd.n7105 585
R2610 gnd.n391 gnd.n390 585
R2611 gnd.n7104 gnd.n391 585
R2612 gnd.n7102 gnd.n7101 585
R2613 gnd.n7103 gnd.n7102 585
R2614 gnd.n394 gnd.n393 585
R2615 gnd.n393 gnd.n392 585
R2616 gnd.n7097 gnd.n7096 585
R2617 gnd.n7096 gnd.n7095 585
R2618 gnd.n397 gnd.n396 585
R2619 gnd.n7094 gnd.n397 585
R2620 gnd.n7092 gnd.n7091 585
R2621 gnd.n7093 gnd.n7092 585
R2622 gnd.n400 gnd.n399 585
R2623 gnd.n399 gnd.n398 585
R2624 gnd.n7087 gnd.n7086 585
R2625 gnd.n7086 gnd.n7085 585
R2626 gnd.n403 gnd.n402 585
R2627 gnd.n7084 gnd.n403 585
R2628 gnd.n7082 gnd.n7081 585
R2629 gnd.n7083 gnd.n7082 585
R2630 gnd.n406 gnd.n405 585
R2631 gnd.n405 gnd.n404 585
R2632 gnd.n7077 gnd.n7076 585
R2633 gnd.n7076 gnd.n7075 585
R2634 gnd.n409 gnd.n408 585
R2635 gnd.n7074 gnd.n409 585
R2636 gnd.n7072 gnd.n7071 585
R2637 gnd.n7073 gnd.n7072 585
R2638 gnd.n412 gnd.n411 585
R2639 gnd.n411 gnd.n410 585
R2640 gnd.n7067 gnd.n7066 585
R2641 gnd.n7066 gnd.n7065 585
R2642 gnd.n415 gnd.n414 585
R2643 gnd.n7064 gnd.n415 585
R2644 gnd.n7062 gnd.n7061 585
R2645 gnd.n7063 gnd.n7062 585
R2646 gnd.n418 gnd.n417 585
R2647 gnd.n417 gnd.n416 585
R2648 gnd.n7057 gnd.n7056 585
R2649 gnd.n7056 gnd.n7055 585
R2650 gnd.n421 gnd.n420 585
R2651 gnd.n7054 gnd.n421 585
R2652 gnd.n7052 gnd.n7051 585
R2653 gnd.n7053 gnd.n7052 585
R2654 gnd.n424 gnd.n423 585
R2655 gnd.n423 gnd.n422 585
R2656 gnd.n7047 gnd.n7046 585
R2657 gnd.n7046 gnd.n7045 585
R2658 gnd.n427 gnd.n426 585
R2659 gnd.n7044 gnd.n427 585
R2660 gnd.n7042 gnd.n7041 585
R2661 gnd.n7043 gnd.n7042 585
R2662 gnd.n430 gnd.n429 585
R2663 gnd.n429 gnd.n428 585
R2664 gnd.n7037 gnd.n7036 585
R2665 gnd.n7036 gnd.n7035 585
R2666 gnd.n433 gnd.n432 585
R2667 gnd.n7034 gnd.n433 585
R2668 gnd.n7032 gnd.n7031 585
R2669 gnd.n7033 gnd.n7032 585
R2670 gnd.n436 gnd.n435 585
R2671 gnd.n435 gnd.n434 585
R2672 gnd.n7027 gnd.n7026 585
R2673 gnd.n7026 gnd.n7025 585
R2674 gnd.n439 gnd.n438 585
R2675 gnd.n7024 gnd.n439 585
R2676 gnd.n7022 gnd.n7021 585
R2677 gnd.n7023 gnd.n7022 585
R2678 gnd.n442 gnd.n441 585
R2679 gnd.n441 gnd.n440 585
R2680 gnd.n7017 gnd.n7016 585
R2681 gnd.n7016 gnd.n7015 585
R2682 gnd.n445 gnd.n444 585
R2683 gnd.n7014 gnd.n445 585
R2684 gnd.n7012 gnd.n7011 585
R2685 gnd.n7013 gnd.n7012 585
R2686 gnd.n448 gnd.n447 585
R2687 gnd.n447 gnd.n446 585
R2688 gnd.n7007 gnd.n7006 585
R2689 gnd.n7006 gnd.n7005 585
R2690 gnd.n451 gnd.n450 585
R2691 gnd.n7004 gnd.n451 585
R2692 gnd.n7002 gnd.n7001 585
R2693 gnd.n7003 gnd.n7002 585
R2694 gnd.n454 gnd.n453 585
R2695 gnd.n453 gnd.n452 585
R2696 gnd.n6997 gnd.n6996 585
R2697 gnd.n6996 gnd.n6995 585
R2698 gnd.n457 gnd.n456 585
R2699 gnd.n6994 gnd.n457 585
R2700 gnd.n6992 gnd.n6991 585
R2701 gnd.n6993 gnd.n6992 585
R2702 gnd.n460 gnd.n459 585
R2703 gnd.n459 gnd.n458 585
R2704 gnd.n6987 gnd.n6986 585
R2705 gnd.n6986 gnd.n6985 585
R2706 gnd.n463 gnd.n462 585
R2707 gnd.n6984 gnd.n463 585
R2708 gnd.n6982 gnd.n6981 585
R2709 gnd.n6983 gnd.n6982 585
R2710 gnd.n466 gnd.n465 585
R2711 gnd.n465 gnd.n464 585
R2712 gnd.n6977 gnd.n6976 585
R2713 gnd.n6976 gnd.n6975 585
R2714 gnd.n469 gnd.n468 585
R2715 gnd.n6974 gnd.n469 585
R2716 gnd.n6972 gnd.n6971 585
R2717 gnd.n6973 gnd.n6972 585
R2718 gnd.n472 gnd.n471 585
R2719 gnd.n471 gnd.n470 585
R2720 gnd.n6967 gnd.n6966 585
R2721 gnd.n6966 gnd.n6965 585
R2722 gnd.n475 gnd.n474 585
R2723 gnd.n6964 gnd.n475 585
R2724 gnd.n6962 gnd.n6961 585
R2725 gnd.n6963 gnd.n6962 585
R2726 gnd.n478 gnd.n477 585
R2727 gnd.n477 gnd.n476 585
R2728 gnd.n6957 gnd.n6956 585
R2729 gnd.n6956 gnd.n6955 585
R2730 gnd.n481 gnd.n480 585
R2731 gnd.n6954 gnd.n481 585
R2732 gnd.n6952 gnd.n6951 585
R2733 gnd.n6953 gnd.n6952 585
R2734 gnd.n484 gnd.n483 585
R2735 gnd.n483 gnd.n482 585
R2736 gnd.n6947 gnd.n6946 585
R2737 gnd.n6946 gnd.n6945 585
R2738 gnd.n487 gnd.n486 585
R2739 gnd.n6944 gnd.n487 585
R2740 gnd.n6942 gnd.n6941 585
R2741 gnd.n6943 gnd.n6942 585
R2742 gnd.n490 gnd.n489 585
R2743 gnd.n489 gnd.n488 585
R2744 gnd.n6937 gnd.n6936 585
R2745 gnd.n6936 gnd.n6935 585
R2746 gnd.n493 gnd.n492 585
R2747 gnd.n6934 gnd.n493 585
R2748 gnd.n6932 gnd.n6931 585
R2749 gnd.n6933 gnd.n6932 585
R2750 gnd.n496 gnd.n495 585
R2751 gnd.n495 gnd.n494 585
R2752 gnd.n6927 gnd.n6926 585
R2753 gnd.n6926 gnd.n6925 585
R2754 gnd.n499 gnd.n498 585
R2755 gnd.n6924 gnd.n499 585
R2756 gnd.n6922 gnd.n6921 585
R2757 gnd.n6923 gnd.n6922 585
R2758 gnd.n502 gnd.n501 585
R2759 gnd.n501 gnd.n500 585
R2760 gnd.n6917 gnd.n6916 585
R2761 gnd.n6916 gnd.n6915 585
R2762 gnd.n505 gnd.n504 585
R2763 gnd.n6914 gnd.n505 585
R2764 gnd.n6912 gnd.n6911 585
R2765 gnd.n6913 gnd.n6912 585
R2766 gnd.n5909 gnd.n5908 585
R2767 gnd.n5910 gnd.n5909 585
R2768 gnd.n2659 gnd.n2658 585
R2769 gnd.n4256 gnd.n2659 585
R2770 gnd.n5918 gnd.n5917 585
R2771 gnd.n5917 gnd.n5916 585
R2772 gnd.n5919 gnd.n2653 585
R2773 gnd.n4248 gnd.n2653 585
R2774 gnd.n5921 gnd.n5920 585
R2775 gnd.n5922 gnd.n5921 585
R2776 gnd.n2637 gnd.n2636 585
R2777 gnd.n4239 gnd.n2637 585
R2778 gnd.n5930 gnd.n5929 585
R2779 gnd.n5929 gnd.n5928 585
R2780 gnd.n5931 gnd.n2631 585
R2781 gnd.n4231 gnd.n2631 585
R2782 gnd.n5933 gnd.n5932 585
R2783 gnd.n5934 gnd.n5933 585
R2784 gnd.n2615 gnd.n2614 585
R2785 gnd.n4223 gnd.n2615 585
R2786 gnd.n5942 gnd.n5941 585
R2787 gnd.n5941 gnd.n5940 585
R2788 gnd.n5943 gnd.n2609 585
R2789 gnd.n4215 gnd.n2609 585
R2790 gnd.n5945 gnd.n5944 585
R2791 gnd.n5946 gnd.n5945 585
R2792 gnd.n2594 gnd.n2593 585
R2793 gnd.n4207 gnd.n2594 585
R2794 gnd.n5954 gnd.n5953 585
R2795 gnd.n5953 gnd.n5952 585
R2796 gnd.n5955 gnd.n2588 585
R2797 gnd.n4199 gnd.n2588 585
R2798 gnd.n5957 gnd.n5956 585
R2799 gnd.n5958 gnd.n5957 585
R2800 gnd.n2572 gnd.n2571 585
R2801 gnd.n4191 gnd.n2572 585
R2802 gnd.n5966 gnd.n5965 585
R2803 gnd.n5965 gnd.n5964 585
R2804 gnd.n5967 gnd.n2566 585
R2805 gnd.n4183 gnd.n2566 585
R2806 gnd.n5969 gnd.n5968 585
R2807 gnd.n5970 gnd.n5969 585
R2808 gnd.n2552 gnd.n2551 585
R2809 gnd.n4175 gnd.n2552 585
R2810 gnd.n5978 gnd.n5977 585
R2811 gnd.n5977 gnd.n5976 585
R2812 gnd.n5979 gnd.n2546 585
R2813 gnd.n4167 gnd.n2546 585
R2814 gnd.n5981 gnd.n5980 585
R2815 gnd.n5982 gnd.n5981 585
R2816 gnd.n2533 gnd.n2532 585
R2817 gnd.n4159 gnd.n2533 585
R2818 gnd.n5991 gnd.n5990 585
R2819 gnd.n5990 gnd.n5989 585
R2820 gnd.n5992 gnd.n2527 585
R2821 gnd.n4150 gnd.n2527 585
R2822 gnd.n5994 gnd.n5993 585
R2823 gnd.n5995 gnd.n5994 585
R2824 gnd.n2514 gnd.n2513 585
R2825 gnd.n4140 gnd.n2514 585
R2826 gnd.n6003 gnd.n6002 585
R2827 gnd.n6002 gnd.n6001 585
R2828 gnd.n6004 gnd.n2508 585
R2829 gnd.n4132 gnd.n2508 585
R2830 gnd.n6006 gnd.n6005 585
R2831 gnd.n6007 gnd.n6006 585
R2832 gnd.n2492 gnd.n2491 585
R2833 gnd.n4124 gnd.n2492 585
R2834 gnd.n6015 gnd.n6014 585
R2835 gnd.n6014 gnd.n6013 585
R2836 gnd.n6016 gnd.n2486 585
R2837 gnd.n4116 gnd.n2486 585
R2838 gnd.n6018 gnd.n6017 585
R2839 gnd.n6019 gnd.n6018 585
R2840 gnd.n2471 gnd.n2470 585
R2841 gnd.n4108 gnd.n2471 585
R2842 gnd.n6027 gnd.n6026 585
R2843 gnd.n6026 gnd.n6025 585
R2844 gnd.n6028 gnd.n2465 585
R2845 gnd.n4100 gnd.n2465 585
R2846 gnd.n6030 gnd.n6029 585
R2847 gnd.n6031 gnd.n6030 585
R2848 gnd.n2449 gnd.n2448 585
R2849 gnd.n4092 gnd.n2449 585
R2850 gnd.n6039 gnd.n6038 585
R2851 gnd.n6038 gnd.n6037 585
R2852 gnd.n6040 gnd.n2443 585
R2853 gnd.n4084 gnd.n2443 585
R2854 gnd.n6042 gnd.n6041 585
R2855 gnd.n6043 gnd.n6042 585
R2856 gnd.n2428 gnd.n2427 585
R2857 gnd.n4076 gnd.n2428 585
R2858 gnd.n6051 gnd.n6050 585
R2859 gnd.n6050 gnd.n6049 585
R2860 gnd.n6052 gnd.n2422 585
R2861 gnd.n4068 gnd.n2422 585
R2862 gnd.n6054 gnd.n6053 585
R2863 gnd.n6055 gnd.n6054 585
R2864 gnd.n2423 gnd.n2421 585
R2865 gnd.n4059 gnd.n2421 585
R2866 gnd.n4040 gnd.n2408 585
R2867 gnd.n6061 gnd.n2408 585
R2868 gnd.n3977 gnd.n3975 585
R2869 gnd.n3975 gnd.n2405 585
R2870 gnd.n4045 gnd.n4044 585
R2871 gnd.n4052 gnd.n4045 585
R2872 gnd.n3976 gnd.n3974 585
R2873 gnd.n3974 gnd.n2351 585
R2874 gnd.n4036 gnd.n4035 585
R2875 gnd.n4034 gnd.n4033 585
R2876 gnd.n4032 gnd.n4031 585
R2877 gnd.n4030 gnd.n4029 585
R2878 gnd.n4028 gnd.n4027 585
R2879 gnd.n4026 gnd.n4025 585
R2880 gnd.n4024 gnd.n4023 585
R2881 gnd.n4022 gnd.n4021 585
R2882 gnd.n4020 gnd.n4019 585
R2883 gnd.n4018 gnd.n4017 585
R2884 gnd.n4016 gnd.n4015 585
R2885 gnd.n4014 gnd.n4013 585
R2886 gnd.n4012 gnd.n4011 585
R2887 gnd.n4010 gnd.n4009 585
R2888 gnd.n4008 gnd.n4007 585
R2889 gnd.n4006 gnd.n4005 585
R2890 gnd.n4004 gnd.n4003 585
R2891 gnd.n3996 gnd.n3993 585
R2892 gnd.n3999 gnd.n2350 585
R2893 gnd.n6148 gnd.n2350 585
R2894 gnd.n4593 gnd.n4592 585
R2895 gnd.n3563 gnd.n3562 585
R2896 gnd.n3664 gnd.n3663 585
R2897 gnd.n3573 gnd.n3572 585
R2898 gnd.n3653 gnd.n3652 585
R2899 gnd.n3651 gnd.n3579 585
R2900 gnd.n3578 gnd.n3577 585
R2901 gnd.n3642 gnd.n3641 585
R2902 gnd.n3640 gnd.n3639 585
R2903 gnd.n3628 gnd.n3585 585
R2904 gnd.n3630 gnd.n3629 585
R2905 gnd.n3627 gnd.n3591 585
R2906 gnd.n3590 gnd.n3589 585
R2907 gnd.n3618 gnd.n3617 585
R2908 gnd.n3616 gnd.n3615 585
R2909 gnd.n3604 gnd.n3597 585
R2910 gnd.n3606 gnd.n3605 585
R2911 gnd.n3603 gnd.n3602 585
R2912 gnd.n2675 gnd.n2673 585
R2913 gnd.n4590 gnd.n2673 585
R2914 gnd.n3734 gnd.n2671 585
R2915 gnd.n5910 gnd.n2671 585
R2916 gnd.n4255 gnd.n4254 585
R2917 gnd.n4256 gnd.n4255 585
R2918 gnd.n3733 gnd.n2662 585
R2919 gnd.n5916 gnd.n2662 585
R2920 gnd.n4250 gnd.n4249 585
R2921 gnd.n4249 gnd.n4248 585
R2922 gnd.n3736 gnd.n2651 585
R2923 gnd.n5922 gnd.n2651 585
R2924 gnd.n4238 gnd.n4237 585
R2925 gnd.n4239 gnd.n4238 585
R2926 gnd.n3740 gnd.n2640 585
R2927 gnd.n5928 gnd.n2640 585
R2928 gnd.n4233 gnd.n4232 585
R2929 gnd.n4232 gnd.n4231 585
R2930 gnd.n3742 gnd.n2629 585
R2931 gnd.n5934 gnd.n2629 585
R2932 gnd.n4222 gnd.n4221 585
R2933 gnd.n4223 gnd.n4222 585
R2934 gnd.n3746 gnd.n2618 585
R2935 gnd.n5940 gnd.n2618 585
R2936 gnd.n4217 gnd.n4216 585
R2937 gnd.n4216 gnd.n4215 585
R2938 gnd.n3748 gnd.n2608 585
R2939 gnd.n5946 gnd.n2608 585
R2940 gnd.n4206 gnd.n4205 585
R2941 gnd.n4207 gnd.n4206 585
R2942 gnd.n3753 gnd.n2597 585
R2943 gnd.n5952 gnd.n2597 585
R2944 gnd.n4201 gnd.n4200 585
R2945 gnd.n4200 gnd.n4199 585
R2946 gnd.n3755 gnd.n2586 585
R2947 gnd.n5958 gnd.n2586 585
R2948 gnd.n4190 gnd.n4189 585
R2949 gnd.n4191 gnd.n4190 585
R2950 gnd.n3759 gnd.n2575 585
R2951 gnd.n5964 gnd.n2575 585
R2952 gnd.n4185 gnd.n4184 585
R2953 gnd.n4184 gnd.n4183 585
R2954 gnd.n3761 gnd.n2565 585
R2955 gnd.n5970 gnd.n2565 585
R2956 gnd.n4174 gnd.n4173 585
R2957 gnd.n4175 gnd.n4174 585
R2958 gnd.n3766 gnd.n2555 585
R2959 gnd.n5976 gnd.n2555 585
R2960 gnd.n4169 gnd.n4168 585
R2961 gnd.n4168 gnd.n4167 585
R2962 gnd.n3768 gnd.n2544 585
R2963 gnd.n5982 gnd.n2544 585
R2964 gnd.n4158 gnd.n4157 585
R2965 gnd.n4159 gnd.n4158 585
R2966 gnd.n3772 gnd.n2536 585
R2967 gnd.n5989 gnd.n2536 585
R2968 gnd.n4152 gnd.n4151 585
R2969 gnd.n4151 gnd.n4150 585
R2970 gnd.n3774 gnd.n2526 585
R2971 gnd.n5995 gnd.n2526 585
R2972 gnd.n4139 gnd.n4138 585
R2973 gnd.n4140 gnd.n4139 585
R2974 gnd.n3779 gnd.n2517 585
R2975 gnd.n6001 gnd.n2517 585
R2976 gnd.n4134 gnd.n4133 585
R2977 gnd.n4133 gnd.n4132 585
R2978 gnd.n3781 gnd.n2506 585
R2979 gnd.n6007 gnd.n2506 585
R2980 gnd.n4123 gnd.n4122 585
R2981 gnd.n4124 gnd.n4123 585
R2982 gnd.n3785 gnd.n2495 585
R2983 gnd.n6013 gnd.n2495 585
R2984 gnd.n4118 gnd.n4117 585
R2985 gnd.n4117 gnd.n4116 585
R2986 gnd.n3787 gnd.n2485 585
R2987 gnd.n6019 gnd.n2485 585
R2988 gnd.n4107 gnd.n4106 585
R2989 gnd.n4108 gnd.n4107 585
R2990 gnd.n3792 gnd.n2474 585
R2991 gnd.n6025 gnd.n2474 585
R2992 gnd.n4102 gnd.n4101 585
R2993 gnd.n4101 gnd.n4100 585
R2994 gnd.n3794 gnd.n2463 585
R2995 gnd.n6031 gnd.n2463 585
R2996 gnd.n4091 gnd.n4090 585
R2997 gnd.n4092 gnd.n4091 585
R2998 gnd.n3798 gnd.n2452 585
R2999 gnd.n6037 gnd.n2452 585
R3000 gnd.n4086 gnd.n4085 585
R3001 gnd.n4085 gnd.n4084 585
R3002 gnd.n3800 gnd.n2442 585
R3003 gnd.n6043 gnd.n2442 585
R3004 gnd.n4075 gnd.n4074 585
R3005 gnd.n4076 gnd.n4075 585
R3006 gnd.n3805 gnd.n2431 585
R3007 gnd.n6049 gnd.n2431 585
R3008 gnd.n4070 gnd.n4069 585
R3009 gnd.n4069 gnd.n4068 585
R3010 gnd.n4062 gnd.n2419 585
R3011 gnd.n6055 gnd.n2419 585
R3012 gnd.n4061 gnd.n4060 585
R3013 gnd.n4060 gnd.n4059 585
R3014 gnd.n3807 gnd.n2406 585
R3015 gnd.n6061 gnd.n2406 585
R3016 gnd.n4055 gnd.n4054 585
R3017 gnd.n4054 gnd.n2405 585
R3018 gnd.n4053 gnd.n3809 585
R3019 gnd.n4053 gnd.n4052 585
R3020 gnd.n3997 gnd.n3810 585
R3021 gnd.n3810 gnd.n2351 585
R3022 gnd.n7346 gnd.n103 585
R3023 gnd.n7442 gnd.n103 585
R3024 gnd.n7347 gnd.n7277 585
R3025 gnd.n7277 gnd.n100 585
R3026 gnd.n7348 gnd.n183 585
R3027 gnd.n7362 gnd.n183 585
R3028 gnd.n195 gnd.n193 585
R3029 gnd.n193 gnd.n181 585
R3030 gnd.n7353 gnd.n7352 585
R3031 gnd.n7354 gnd.n7353 585
R3032 gnd.n194 gnd.n192 585
R3033 gnd.n359 gnd.n192 585
R3034 gnd.n7273 gnd.n7272 585
R3035 gnd.n7272 gnd.n7271 585
R3036 gnd.n198 gnd.n197 585
R3037 gnd.n7132 gnd.n198 585
R3038 gnd.n7262 gnd.n7261 585
R3039 gnd.n7263 gnd.n7262 585
R3040 gnd.n210 gnd.n209 585
R3041 gnd.n7136 gnd.n209 585
R3042 gnd.n7257 gnd.n7256 585
R3043 gnd.n7256 gnd.n7255 585
R3044 gnd.n213 gnd.n212 585
R3045 gnd.n7143 gnd.n213 585
R3046 gnd.n7246 gnd.n7245 585
R3047 gnd.n7247 gnd.n7246 585
R3048 gnd.n225 gnd.n224 585
R3049 gnd.n342 gnd.n224 585
R3050 gnd.n7241 gnd.n7240 585
R3051 gnd.n7240 gnd.n7239 585
R3052 gnd.n228 gnd.n227 585
R3053 gnd.n7152 gnd.n228 585
R3054 gnd.n7230 gnd.n7229 585
R3055 gnd.n7231 gnd.n7230 585
R3056 gnd.n240 gnd.n239 585
R3057 gnd.n7156 gnd.n239 585
R3058 gnd.n7225 gnd.n7224 585
R3059 gnd.n7224 gnd.n7223 585
R3060 gnd.n243 gnd.n242 585
R3061 gnd.n7163 gnd.n243 585
R3062 gnd.n7214 gnd.n7213 585
R3063 gnd.n7215 gnd.n7214 585
R3064 gnd.n255 gnd.n254 585
R3065 gnd.n310 gnd.n254 585
R3066 gnd.n7209 gnd.n7208 585
R3067 gnd.n7208 gnd.n7207 585
R3068 gnd.n258 gnd.n257 585
R3069 gnd.n7173 gnd.n258 585
R3070 gnd.n7186 gnd.n7185 585
R3071 gnd.n7185 gnd.n7184 585
R3072 gnd.n7187 gnd.n289 585
R3073 gnd.n7179 gnd.n289 585
R3074 gnd.n5619 gnd.n286 585
R3075 gnd.n5620 gnd.n5619 585
R3076 gnd.n7192 gnd.n285 585
R3077 gnd.n5632 gnd.n285 585
R3078 gnd.n7193 gnd.n284 585
R3079 gnd.n5636 gnd.n284 585
R3080 gnd.n7194 gnd.n283 585
R3081 gnd.n2926 gnd.n283 585
R3082 gnd.n280 gnd.n278 585
R3083 gnd.n5609 gnd.n278 585
R3084 gnd.n7199 gnd.n7198 585
R3085 gnd.n7200 gnd.n7199 585
R3086 gnd.n279 gnd.n277 585
R3087 gnd.n5597 gnd.n277 585
R3088 gnd.n5662 gnd.n5660 585
R3089 gnd.n5660 gnd.n5659 585
R3090 gnd.n5663 gnd.n2901 585
R3091 gnd.n2913 gnd.n2901 585
R3092 gnd.n5664 gnd.n2900 585
R3093 gnd.n5651 gnd.n2900 585
R3094 gnd.n5583 gnd.n2898 585
R3095 gnd.n5584 gnd.n5583 585
R3096 gnd.n5668 gnd.n2897 585
R3097 gnd.n2956 gnd.n2897 585
R3098 gnd.n5669 gnd.n2896 585
R3099 gnd.n5571 gnd.n2896 585
R3100 gnd.n5670 gnd.n2895 585
R3101 gnd.n2965 gnd.n2895 585
R3102 gnd.n5560 gnd.n2893 585
R3103 gnd.n5561 gnd.n5560 585
R3104 gnd.n5674 gnd.n2892 585
R3105 gnd.n5541 gnd.n2892 585
R3106 gnd.n5675 gnd.n2891 585
R3107 gnd.n2973 gnd.n2891 585
R3108 gnd.n5676 gnd.n2890 585
R3109 gnd.n5532 gnd.n2890 585
R3110 gnd.n2993 gnd.n2888 585
R3111 gnd.n2994 gnd.n2993 585
R3112 gnd.n5680 gnd.n2887 585
R3113 gnd.n5522 gnd.n2887 585
R3114 gnd.n5681 gnd.n2886 585
R3115 gnd.n5510 gnd.n2886 585
R3116 gnd.n5682 gnd.n2885 585
R3117 gnd.n3001 gnd.n2885 585
R3118 gnd.n3012 gnd.n2883 585
R3119 gnd.n5501 gnd.n3012 585
R3120 gnd.n5686 gnd.n2882 585
R3121 gnd.n3022 gnd.n2882 585
R3122 gnd.n5687 gnd.n2881 585
R3123 gnd.n5491 gnd.n2881 585
R3124 gnd.n5688 gnd.n2880 585
R3125 gnd.n5479 gnd.n2880 585
R3126 gnd.n2877 gnd.n2876 585
R3127 gnd.n3041 gnd.n2876 585
R3128 gnd.n5693 gnd.n5692 585
R3129 gnd.n5694 gnd.n5693 585
R3130 gnd.n3126 gnd.n2875 585
R3131 gnd.n3130 gnd.n3129 585
R3132 gnd.n3132 gnd.n3131 585
R3133 gnd.n3121 gnd.n3120 585
R3134 gnd.n3144 gnd.n3122 585
R3135 gnd.n3146 gnd.n3145 585
R3136 gnd.n3148 gnd.n3147 585
R3137 gnd.n3112 gnd.n3111 585
R3138 gnd.n3161 gnd.n3113 585
R3139 gnd.n3163 gnd.n3162 585
R3140 gnd.n3165 gnd.n3164 585
R3141 gnd.n3103 gnd.n3102 585
R3142 gnd.n3178 gnd.n3104 585
R3143 gnd.n3180 gnd.n3179 585
R3144 gnd.n3182 gnd.n3181 585
R3145 gnd.n3094 gnd.n3093 585
R3146 gnd.n3195 gnd.n3095 585
R3147 gnd.n3196 gnd.n3090 585
R3148 gnd.n3197 gnd.n2820 585
R3149 gnd.n5770 gnd.n2820 585
R3150 gnd.n7317 gnd.n99 585
R3151 gnd.n7318 gnd.n7315 585
R3152 gnd.n7319 gnd.n7311 585
R3153 gnd.n7309 gnd.n7307 585
R3154 gnd.n7323 gnd.n7306 585
R3155 gnd.n7324 gnd.n7304 585
R3156 gnd.n7325 gnd.n7303 585
R3157 gnd.n7301 gnd.n7299 585
R3158 gnd.n7329 gnd.n7298 585
R3159 gnd.n7330 gnd.n7296 585
R3160 gnd.n7331 gnd.n7295 585
R3161 gnd.n7293 gnd.n7291 585
R3162 gnd.n7335 gnd.n7290 585
R3163 gnd.n7336 gnd.n7288 585
R3164 gnd.n7337 gnd.n7287 585
R3165 gnd.n7285 gnd.n7283 585
R3166 gnd.n7341 gnd.n7282 585
R3167 gnd.n7342 gnd.n7280 585
R3168 gnd.n7343 gnd.n7279 585
R3169 gnd.n7279 gnd.n102 585
R3170 gnd.n7444 gnd.n7443 585
R3171 gnd.n7443 gnd.n7442 585
R3172 gnd.n7445 gnd.n97 585
R3173 gnd.n100 gnd.n97 585
R3174 gnd.n7446 gnd.n96 585
R3175 gnd.n7362 gnd.n96 585
R3176 gnd.n180 gnd.n94 585
R3177 gnd.n181 gnd.n180 585
R3178 gnd.n7450 gnd.n93 585
R3179 gnd.n7354 gnd.n93 585
R3180 gnd.n7451 gnd.n92 585
R3181 gnd.n359 gnd.n92 585
R3182 gnd.n7452 gnd.n91 585
R3183 gnd.n7271 gnd.n91 585
R3184 gnd.n363 gnd.n89 585
R3185 gnd.n7132 gnd.n363 585
R3186 gnd.n7456 gnd.n88 585
R3187 gnd.n7263 gnd.n88 585
R3188 gnd.n7457 gnd.n87 585
R3189 gnd.n7136 gnd.n87 585
R3190 gnd.n7458 gnd.n86 585
R3191 gnd.n7255 gnd.n86 585
R3192 gnd.n7142 gnd.n84 585
R3193 gnd.n7143 gnd.n7142 585
R3194 gnd.n7462 gnd.n83 585
R3195 gnd.n7247 gnd.n83 585
R3196 gnd.n7463 gnd.n82 585
R3197 gnd.n342 gnd.n82 585
R3198 gnd.n7464 gnd.n81 585
R3199 gnd.n7239 gnd.n81 585
R3200 gnd.n321 gnd.n79 585
R3201 gnd.n7152 gnd.n321 585
R3202 gnd.n7468 gnd.n78 585
R3203 gnd.n7231 gnd.n78 585
R3204 gnd.n7469 gnd.n77 585
R3205 gnd.n7156 gnd.n77 585
R3206 gnd.n7470 gnd.n76 585
R3207 gnd.n7223 gnd.n76 585
R3208 gnd.n7162 gnd.n74 585
R3209 gnd.n7163 gnd.n7162 585
R3210 gnd.n7474 gnd.n73 585
R3211 gnd.n7215 gnd.n73 585
R3212 gnd.n7475 gnd.n72 585
R3213 gnd.n310 gnd.n72 585
R3214 gnd.n7476 gnd.n71 585
R3215 gnd.n7207 gnd.n71 585
R3216 gnd.n301 gnd.n69 585
R3217 gnd.n7173 gnd.n301 585
R3218 gnd.n7480 gnd.n68 585
R3219 gnd.n7184 gnd.n68 585
R3220 gnd.n7481 gnd.n67 585
R3221 gnd.n7179 gnd.n67 585
R3222 gnd.n7482 gnd.n66 585
R3223 gnd.n5620 gnd.n66 585
R3224 gnd.n5618 gnd.n65 585
R3225 gnd.n5632 gnd.n5618 585
R3226 gnd.n5602 gnd.n2928 585
R3227 gnd.n5636 gnd.n2928 585
R3228 gnd.n2938 gnd.n2936 585
R3229 gnd.n2936 gnd.n2926 585
R3230 gnd.n5607 gnd.n5606 585
R3231 gnd.n5609 gnd.n5607 585
R3232 gnd.n2937 gnd.n275 585
R3233 gnd.n7200 gnd.n275 585
R3234 gnd.n5599 gnd.n5598 585
R3235 gnd.n5598 gnd.n5597 585
R3236 gnd.n2940 gnd.n2903 585
R3237 gnd.n5659 gnd.n2903 585
R3238 gnd.n5577 gnd.n5576 585
R3239 gnd.n5576 gnd.n2913 585
R3240 gnd.n2949 gnd.n2912 585
R3241 gnd.n5651 gnd.n2912 585
R3242 gnd.n5582 gnd.n5581 585
R3243 gnd.n5584 gnd.n5582 585
R3244 gnd.n2948 gnd.n2947 585
R3245 gnd.n2956 gnd.n2947 585
R3246 gnd.n5573 gnd.n5572 585
R3247 gnd.n5572 gnd.n5571 585
R3248 gnd.n2952 gnd.n2951 585
R3249 gnd.n2965 gnd.n2952 585
R3250 gnd.n2977 gnd.n2964 585
R3251 gnd.n5561 gnd.n2964 585
R3252 gnd.n5540 gnd.n5539 585
R3253 gnd.n5541 gnd.n5540 585
R3254 gnd.n2976 gnd.n2975 585
R3255 gnd.n2975 gnd.n2973 585
R3256 gnd.n5534 gnd.n5533 585
R3257 gnd.n5533 gnd.n5532 585
R3258 gnd.n2980 gnd.n2979 585
R3259 gnd.n2994 gnd.n2980 585
R3260 gnd.n3005 gnd.n2992 585
R3261 gnd.n5522 gnd.n2992 585
R3262 gnd.n5509 gnd.n5508 585
R3263 gnd.n5510 gnd.n5509 585
R3264 gnd.n3004 gnd.n3003 585
R3265 gnd.n3003 gnd.n3001 585
R3266 gnd.n5503 gnd.n5502 585
R3267 gnd.n5502 gnd.n5501 585
R3268 gnd.n3008 gnd.n3007 585
R3269 gnd.n3022 gnd.n3008 585
R3270 gnd.n3081 gnd.n3021 585
R3271 gnd.n5491 gnd.n3021 585
R3272 gnd.n5478 gnd.n5477 585
R3273 gnd.n5479 gnd.n5478 585
R3274 gnd.n3080 gnd.n3079 585
R3275 gnd.n3079 gnd.n3041 585
R3276 gnd.n5472 gnd.n2873 585
R3277 gnd.n5694 gnd.n2873 585
R3278 gnd.n6210 gnd.n6209 585
R3279 gnd.n6211 gnd.n6210 585
R3280 gnd.n1046 gnd.n1044 585
R3281 gnd.n1044 gnd.n1040 585
R3282 gnd.n1026 gnd.n1025 585
R3283 gnd.n2313 gnd.n1026 585
R3284 gnd.n6221 gnd.n6220 585
R3285 gnd.n6220 gnd.n6219 585
R3286 gnd.n6222 gnd.n1020 585
R3287 gnd.n1968 gnd.n1020 585
R3288 gnd.n6224 gnd.n6223 585
R3289 gnd.n6225 gnd.n6224 585
R3290 gnd.n1021 gnd.n1019 585
R3291 gnd.n1019 gnd.n1015 585
R3292 gnd.n1000 gnd.n999 585
R3293 gnd.n1004 gnd.n1000 585
R3294 gnd.n6235 gnd.n6234 585
R3295 gnd.n6234 gnd.n6233 585
R3296 gnd.n6236 gnd.n994 585
R3297 gnd.n1977 gnd.n994 585
R3298 gnd.n6238 gnd.n6237 585
R3299 gnd.n6239 gnd.n6238 585
R3300 gnd.n995 gnd.n993 585
R3301 gnd.n993 gnd.n989 585
R3302 gnd.n976 gnd.n975 585
R3303 gnd.n980 gnd.n976 585
R3304 gnd.n6249 gnd.n6248 585
R3305 gnd.n6248 gnd.n6247 585
R3306 gnd.n6250 gnd.n970 585
R3307 gnd.n1986 gnd.n970 585
R3308 gnd.n6252 gnd.n6251 585
R3309 gnd.n6253 gnd.n6252 585
R3310 gnd.n971 gnd.n969 585
R3311 gnd.n1167 gnd.n969 585
R3312 gnd.n2013 gnd.n2012 585
R3313 gnd.n2012 gnd.n2011 585
R3314 gnd.n1164 gnd.n1163 585
R3315 gnd.n1995 gnd.n1164 585
R3316 gnd.n1942 gnd.n1184 585
R3317 gnd.n1184 gnd.n1174 585
R3318 gnd.n1944 gnd.n1943 585
R3319 gnd.n1945 gnd.n1944 585
R3320 gnd.n1185 gnd.n1183 585
R3321 gnd.n1193 gnd.n1183 585
R3322 gnd.n1918 gnd.n1205 585
R3323 gnd.n1205 gnd.n1192 585
R3324 gnd.n1920 gnd.n1919 585
R3325 gnd.n1921 gnd.n1920 585
R3326 gnd.n1206 gnd.n1204 585
R3327 gnd.n1204 gnd.n1200 585
R3328 gnd.n1906 gnd.n1905 585
R3329 gnd.n1905 gnd.n1904 585
R3330 gnd.n1211 gnd.n1210 585
R3331 gnd.n1220 gnd.n1211 585
R3332 gnd.n1895 gnd.n1894 585
R3333 gnd.n1894 gnd.n1893 585
R3334 gnd.n1218 gnd.n1217 585
R3335 gnd.n1881 gnd.n1218 585
R3336 gnd.n1319 gnd.n1318 585
R3337 gnd.n1319 gnd.n1227 585
R3338 gnd.n1838 gnd.n1837 585
R3339 gnd.n1837 gnd.n1836 585
R3340 gnd.n1839 gnd.n1313 585
R3341 gnd.n1324 gnd.n1313 585
R3342 gnd.n1841 gnd.n1840 585
R3343 gnd.n1842 gnd.n1841 585
R3344 gnd.n1314 gnd.n1312 585
R3345 gnd.n1337 gnd.n1312 585
R3346 gnd.n1297 gnd.n1296 585
R3347 gnd.n1300 gnd.n1297 585
R3348 gnd.n1852 gnd.n1851 585
R3349 gnd.n1851 gnd.n1850 585
R3350 gnd.n1853 gnd.n1291 585
R3351 gnd.n1812 gnd.n1291 585
R3352 gnd.n1855 gnd.n1854 585
R3353 gnd.n1856 gnd.n1855 585
R3354 gnd.n1292 gnd.n1290 585
R3355 gnd.n1351 gnd.n1290 585
R3356 gnd.n1804 gnd.n1803 585
R3357 gnd.n1803 gnd.n1802 585
R3358 gnd.n1348 gnd.n1347 585
R3359 gnd.n1786 gnd.n1348 585
R3360 gnd.n1773 gnd.n1367 585
R3361 gnd.n1367 gnd.n1366 585
R3362 gnd.n1775 gnd.n1774 585
R3363 gnd.n1776 gnd.n1775 585
R3364 gnd.n1368 gnd.n1365 585
R3365 gnd.n1374 gnd.n1365 585
R3366 gnd.n1754 gnd.n1753 585
R3367 gnd.n1755 gnd.n1754 585
R3368 gnd.n1385 gnd.n1384 585
R3369 gnd.n1384 gnd.n1380 585
R3370 gnd.n1744 gnd.n1743 585
R3371 gnd.n1745 gnd.n1744 585
R3372 gnd.n1395 gnd.n1394 585
R3373 gnd.n1400 gnd.n1394 585
R3374 gnd.n1722 gnd.n1413 585
R3375 gnd.n1413 gnd.n1399 585
R3376 gnd.n1724 gnd.n1723 585
R3377 gnd.n1725 gnd.n1724 585
R3378 gnd.n1414 gnd.n1412 585
R3379 gnd.n1412 gnd.n1408 585
R3380 gnd.n1713 gnd.n1712 585
R3381 gnd.n1714 gnd.n1713 585
R3382 gnd.n1421 gnd.n1420 585
R3383 gnd.n1425 gnd.n1420 585
R3384 gnd.n1690 gnd.n1442 585
R3385 gnd.n1442 gnd.n1424 585
R3386 gnd.n1692 gnd.n1691 585
R3387 gnd.n1693 gnd.n1692 585
R3388 gnd.n1443 gnd.n1441 585
R3389 gnd.n1441 gnd.n1432 585
R3390 gnd.n1685 gnd.n1684 585
R3391 gnd.n1684 gnd.n1683 585
R3392 gnd.n1490 gnd.n1489 585
R3393 gnd.n1491 gnd.n1490 585
R3394 gnd.n1644 gnd.n1643 585
R3395 gnd.n1645 gnd.n1644 585
R3396 gnd.n1500 gnd.n1499 585
R3397 gnd.n1499 gnd.n1498 585
R3398 gnd.n1639 gnd.n1638 585
R3399 gnd.n1638 gnd.n1637 585
R3400 gnd.n1503 gnd.n1502 585
R3401 gnd.n1504 gnd.n1503 585
R3402 gnd.n1628 gnd.n1627 585
R3403 gnd.n1629 gnd.n1628 585
R3404 gnd.n1511 gnd.n1510 585
R3405 gnd.n1620 gnd.n1510 585
R3406 gnd.n1623 gnd.n1622 585
R3407 gnd.n1622 gnd.n1621 585
R3408 gnd.n1514 gnd.n1513 585
R3409 gnd.n1515 gnd.n1514 585
R3410 gnd.n1609 gnd.n1608 585
R3411 gnd.n1607 gnd.n1533 585
R3412 gnd.n1606 gnd.n1532 585
R3413 gnd.n1611 gnd.n1532 585
R3414 gnd.n1605 gnd.n1604 585
R3415 gnd.n1603 gnd.n1602 585
R3416 gnd.n1601 gnd.n1600 585
R3417 gnd.n1599 gnd.n1598 585
R3418 gnd.n1597 gnd.n1596 585
R3419 gnd.n1595 gnd.n1594 585
R3420 gnd.n1593 gnd.n1592 585
R3421 gnd.n1591 gnd.n1590 585
R3422 gnd.n1589 gnd.n1588 585
R3423 gnd.n1587 gnd.n1586 585
R3424 gnd.n1585 gnd.n1584 585
R3425 gnd.n1583 gnd.n1582 585
R3426 gnd.n1581 gnd.n1580 585
R3427 gnd.n1579 gnd.n1578 585
R3428 gnd.n1577 gnd.n1576 585
R3429 gnd.n1575 gnd.n1574 585
R3430 gnd.n1573 gnd.n1572 585
R3431 gnd.n1571 gnd.n1570 585
R3432 gnd.n1569 gnd.n1568 585
R3433 gnd.n1567 gnd.n1566 585
R3434 gnd.n1565 gnd.n1564 585
R3435 gnd.n1563 gnd.n1562 585
R3436 gnd.n1520 gnd.n1519 585
R3437 gnd.n1614 gnd.n1613 585
R3438 gnd.n2321 gnd.n2320 585
R3439 gnd.n1070 gnd.n1069 585
R3440 gnd.n1146 gnd.n1145 585
R3441 gnd.n1144 gnd.n1143 585
R3442 gnd.n1142 gnd.n1141 585
R3443 gnd.n1135 gnd.n1075 585
R3444 gnd.n1137 gnd.n1136 585
R3445 gnd.n1134 gnd.n1133 585
R3446 gnd.n1132 gnd.n1131 585
R3447 gnd.n1125 gnd.n1077 585
R3448 gnd.n1127 gnd.n1126 585
R3449 gnd.n1124 gnd.n1123 585
R3450 gnd.n1122 gnd.n1121 585
R3451 gnd.n1115 gnd.n1079 585
R3452 gnd.n1117 gnd.n1116 585
R3453 gnd.n1114 gnd.n1113 585
R3454 gnd.n1112 gnd.n1111 585
R3455 gnd.n1105 gnd.n1081 585
R3456 gnd.n1107 gnd.n1106 585
R3457 gnd.n1104 gnd.n1103 585
R3458 gnd.n1102 gnd.n1101 585
R3459 gnd.n1095 gnd.n1083 585
R3460 gnd.n1097 gnd.n1096 585
R3461 gnd.n1094 gnd.n1093 585
R3462 gnd.n1092 gnd.n1091 585
R3463 gnd.n1086 gnd.n1085 585
R3464 gnd.n1087 gnd.n1045 585
R3465 gnd.n6195 gnd.n1045 585
R3466 gnd.n2317 gnd.n1042 585
R3467 gnd.n6211 gnd.n1042 585
R3468 gnd.n2316 gnd.n2315 585
R3469 gnd.n2315 gnd.n1040 585
R3470 gnd.n2314 gnd.n1150 585
R3471 gnd.n2314 gnd.n2313 585
R3472 gnd.n1967 gnd.n1028 585
R3473 gnd.n6219 gnd.n1028 585
R3474 gnd.n1970 gnd.n1969 585
R3475 gnd.n1969 gnd.n1968 585
R3476 gnd.n1971 gnd.n1017 585
R3477 gnd.n6225 gnd.n1017 585
R3478 gnd.n1973 gnd.n1972 585
R3479 gnd.n1973 gnd.n1015 585
R3480 gnd.n1975 gnd.n1974 585
R3481 gnd.n1974 gnd.n1004 585
R3482 gnd.n1976 gnd.n1002 585
R3483 gnd.n6233 gnd.n1002 585
R3484 gnd.n1979 gnd.n1978 585
R3485 gnd.n1978 gnd.n1977 585
R3486 gnd.n1980 gnd.n991 585
R3487 gnd.n6239 gnd.n991 585
R3488 gnd.n1982 gnd.n1981 585
R3489 gnd.n1982 gnd.n989 585
R3490 gnd.n1984 gnd.n1983 585
R3491 gnd.n1983 gnd.n980 585
R3492 gnd.n1985 gnd.n978 585
R3493 gnd.n6247 gnd.n978 585
R3494 gnd.n1988 gnd.n1987 585
R3495 gnd.n1987 gnd.n1986 585
R3496 gnd.n1989 gnd.n967 585
R3497 gnd.n6253 gnd.n967 585
R3498 gnd.n1991 gnd.n1990 585
R3499 gnd.n1990 gnd.n1167 585
R3500 gnd.n1992 gnd.n1166 585
R3501 gnd.n2011 gnd.n1166 585
R3502 gnd.n1994 gnd.n1993 585
R3503 gnd.n1995 gnd.n1994 585
R3504 gnd.n1177 gnd.n1176 585
R3505 gnd.n1176 gnd.n1174 585
R3506 gnd.n1947 gnd.n1946 585
R3507 gnd.n1946 gnd.n1945 585
R3508 gnd.n1180 gnd.n1179 585
R3509 gnd.n1193 gnd.n1180 585
R3510 gnd.n1869 gnd.n1868 585
R3511 gnd.n1868 gnd.n1192 585
R3512 gnd.n1870 gnd.n1202 585
R3513 gnd.n1921 gnd.n1202 585
R3514 gnd.n1872 gnd.n1871 585
R3515 gnd.n1871 gnd.n1200 585
R3516 gnd.n1873 gnd.n1213 585
R3517 gnd.n1904 gnd.n1213 585
R3518 gnd.n1875 gnd.n1874 585
R3519 gnd.n1874 gnd.n1220 585
R3520 gnd.n1876 gnd.n1219 585
R3521 gnd.n1893 gnd.n1219 585
R3522 gnd.n1878 gnd.n1877 585
R3523 gnd.n1881 gnd.n1878 585
R3524 gnd.n1230 gnd.n1229 585
R3525 gnd.n1229 gnd.n1227 585
R3526 gnd.n1321 gnd.n1320 585
R3527 gnd.n1836 gnd.n1320 585
R3528 gnd.n1323 gnd.n1322 585
R3529 gnd.n1324 gnd.n1323 585
R3530 gnd.n1334 gnd.n1310 585
R3531 gnd.n1842 gnd.n1310 585
R3532 gnd.n1336 gnd.n1335 585
R3533 gnd.n1337 gnd.n1336 585
R3534 gnd.n1333 gnd.n1332 585
R3535 gnd.n1333 gnd.n1300 585
R3536 gnd.n1331 gnd.n1298 585
R3537 gnd.n1850 gnd.n1298 585
R3538 gnd.n1287 gnd.n1285 585
R3539 gnd.n1812 gnd.n1287 585
R3540 gnd.n1858 gnd.n1857 585
R3541 gnd.n1857 gnd.n1856 585
R3542 gnd.n1286 gnd.n1284 585
R3543 gnd.n1351 gnd.n1286 585
R3544 gnd.n1783 gnd.n1350 585
R3545 gnd.n1802 gnd.n1350 585
R3546 gnd.n1785 gnd.n1784 585
R3547 gnd.n1786 gnd.n1785 585
R3548 gnd.n1360 gnd.n1359 585
R3549 gnd.n1366 gnd.n1359 585
R3550 gnd.n1778 gnd.n1777 585
R3551 gnd.n1777 gnd.n1776 585
R3552 gnd.n1363 gnd.n1362 585
R3553 gnd.n1374 gnd.n1363 585
R3554 gnd.n1663 gnd.n1382 585
R3555 gnd.n1755 gnd.n1382 585
R3556 gnd.n1665 gnd.n1664 585
R3557 gnd.n1664 gnd.n1380 585
R3558 gnd.n1666 gnd.n1393 585
R3559 gnd.n1745 gnd.n1393 585
R3560 gnd.n1668 gnd.n1667 585
R3561 gnd.n1668 gnd.n1400 585
R3562 gnd.n1670 gnd.n1669 585
R3563 gnd.n1669 gnd.n1399 585
R3564 gnd.n1671 gnd.n1410 585
R3565 gnd.n1725 gnd.n1410 585
R3566 gnd.n1673 gnd.n1672 585
R3567 gnd.n1672 gnd.n1408 585
R3568 gnd.n1674 gnd.n1419 585
R3569 gnd.n1714 gnd.n1419 585
R3570 gnd.n1676 gnd.n1675 585
R3571 gnd.n1676 gnd.n1425 585
R3572 gnd.n1678 gnd.n1677 585
R3573 gnd.n1677 gnd.n1424 585
R3574 gnd.n1679 gnd.n1440 585
R3575 gnd.n1693 gnd.n1440 585
R3576 gnd.n1680 gnd.n1493 585
R3577 gnd.n1493 gnd.n1432 585
R3578 gnd.n1682 gnd.n1681 585
R3579 gnd.n1683 gnd.n1682 585
R3580 gnd.n1494 gnd.n1492 585
R3581 gnd.n1492 gnd.n1491 585
R3582 gnd.n1647 gnd.n1646 585
R3583 gnd.n1646 gnd.n1645 585
R3584 gnd.n1497 gnd.n1496 585
R3585 gnd.n1498 gnd.n1497 585
R3586 gnd.n1636 gnd.n1635 585
R3587 gnd.n1637 gnd.n1636 585
R3588 gnd.n1506 gnd.n1505 585
R3589 gnd.n1505 gnd.n1504 585
R3590 gnd.n1631 gnd.n1630 585
R3591 gnd.n1630 gnd.n1629 585
R3592 gnd.n1509 gnd.n1508 585
R3593 gnd.n1620 gnd.n1509 585
R3594 gnd.n1619 gnd.n1618 585
R3595 gnd.n1621 gnd.n1619 585
R3596 gnd.n1517 gnd.n1516 585
R3597 gnd.n1516 gnd.n1515 585
R3598 gnd.n1039 gnd.n1038 585
R3599 gnd.n1043 gnd.n1039 585
R3600 gnd.n6214 gnd.n6213 585
R3601 gnd.n6213 gnd.n6212 585
R3602 gnd.n6215 gnd.n1031 585
R3603 gnd.n2312 gnd.n1031 585
R3604 gnd.n6217 gnd.n6216 585
R3605 gnd.n6218 gnd.n6217 585
R3606 gnd.n1032 gnd.n1030 585
R3607 gnd.n1030 gnd.n1027 585
R3608 gnd.n1014 gnd.n1013 585
R3609 gnd.n1018 gnd.n1014 585
R3610 gnd.n6228 gnd.n6227 585
R3611 gnd.n6227 gnd.n6226 585
R3612 gnd.n6229 gnd.n1006 585
R3613 gnd.n1151 gnd.n1006 585
R3614 gnd.n6231 gnd.n6230 585
R3615 gnd.n6232 gnd.n6231 585
R3616 gnd.n1007 gnd.n1005 585
R3617 gnd.n1005 gnd.n1001 585
R3618 gnd.n988 gnd.n987 585
R3619 gnd.n992 gnd.n988 585
R3620 gnd.n6242 gnd.n6241 585
R3621 gnd.n6241 gnd.n6240 585
R3622 gnd.n6243 gnd.n982 585
R3623 gnd.n1154 gnd.n982 585
R3624 gnd.n6245 gnd.n6244 585
R3625 gnd.n6246 gnd.n6245 585
R3626 gnd.n983 gnd.n981 585
R3627 gnd.n981 gnd.n977 585
R3628 gnd.n2006 gnd.n2005 585
R3629 gnd.n2005 gnd.n968 585
R3630 gnd.n2007 gnd.n1169 585
R3631 gnd.n1169 gnd.n966 585
R3632 gnd.n2009 gnd.n2008 585
R3633 gnd.n2010 gnd.n2009 585
R3634 gnd.n1170 gnd.n1168 585
R3635 gnd.n1168 gnd.n1165 585
R3636 gnd.n1998 gnd.n1997 585
R3637 gnd.n1997 gnd.n1996 585
R3638 gnd.n1173 gnd.n1172 585
R3639 gnd.n1182 gnd.n1173 585
R3640 gnd.n1929 gnd.n1195 585
R3641 gnd.n1195 gnd.n1181 585
R3642 gnd.n1931 gnd.n1930 585
R3643 gnd.n1932 gnd.n1931 585
R3644 gnd.n1196 gnd.n1194 585
R3645 gnd.n1203 gnd.n1194 585
R3646 gnd.n1924 gnd.n1923 585
R3647 gnd.n1923 gnd.n1922 585
R3648 gnd.n1199 gnd.n1198 585
R3649 gnd.n1903 gnd.n1199 585
R3650 gnd.n1889 gnd.n1222 585
R3651 gnd.n1222 gnd.n1212 585
R3652 gnd.n1891 gnd.n1890 585
R3653 gnd.n1892 gnd.n1891 585
R3654 gnd.n1223 gnd.n1221 585
R3655 gnd.n1880 gnd.n1221 585
R3656 gnd.n1884 gnd.n1883 585
R3657 gnd.n1883 gnd.n1882 585
R3658 gnd.n1226 gnd.n1225 585
R3659 gnd.n1835 gnd.n1226 585
R3660 gnd.n1328 gnd.n1327 585
R3661 gnd.n1329 gnd.n1328 585
R3662 gnd.n1308 gnd.n1307 585
R3663 gnd.n1311 gnd.n1308 585
R3664 gnd.n1845 gnd.n1844 585
R3665 gnd.n1844 gnd.n1843 585
R3666 gnd.n1846 gnd.n1302 585
R3667 gnd.n1338 gnd.n1302 585
R3668 gnd.n1848 gnd.n1847 585
R3669 gnd.n1849 gnd.n1848 585
R3670 gnd.n1303 gnd.n1301 585
R3671 gnd.n1813 gnd.n1301 585
R3672 gnd.n1797 gnd.n1796 585
R3673 gnd.n1796 gnd.n1289 585
R3674 gnd.n1798 gnd.n1353 585
R3675 gnd.n1353 gnd.n1288 585
R3676 gnd.n1800 gnd.n1799 585
R3677 gnd.n1801 gnd.n1800 585
R3678 gnd.n1354 gnd.n1352 585
R3679 gnd.n1352 gnd.n1349 585
R3680 gnd.n1789 gnd.n1788 585
R3681 gnd.n1788 gnd.n1787 585
R3682 gnd.n1357 gnd.n1356 585
R3683 gnd.n1364 gnd.n1357 585
R3684 gnd.n1763 gnd.n1762 585
R3685 gnd.n1764 gnd.n1763 585
R3686 gnd.n1376 gnd.n1375 585
R3687 gnd.n1383 gnd.n1375 585
R3688 gnd.n1758 gnd.n1757 585
R3689 gnd.n1757 gnd.n1756 585
R3690 gnd.n1379 gnd.n1378 585
R3691 gnd.n1746 gnd.n1379 585
R3692 gnd.n1733 gnd.n1403 585
R3693 gnd.n1403 gnd.n1402 585
R3694 gnd.n1735 gnd.n1734 585
R3695 gnd.n1736 gnd.n1735 585
R3696 gnd.n1404 gnd.n1401 585
R3697 gnd.n1411 gnd.n1401 585
R3698 gnd.n1728 gnd.n1727 585
R3699 gnd.n1727 gnd.n1726 585
R3700 gnd.n1407 gnd.n1406 585
R3701 gnd.n1715 gnd.n1407 585
R3702 gnd.n1702 gnd.n1428 585
R3703 gnd.n1428 gnd.n1427 585
R3704 gnd.n1704 gnd.n1703 585
R3705 gnd.n1705 gnd.n1704 585
R3706 gnd.n1698 gnd.n1426 585
R3707 gnd.n1697 gnd.n1696 585
R3708 gnd.n1431 gnd.n1430 585
R3709 gnd.n1694 gnd.n1431 585
R3710 gnd.n1453 gnd.n1452 585
R3711 gnd.n1456 gnd.n1455 585
R3712 gnd.n1454 gnd.n1449 585
R3713 gnd.n1461 gnd.n1460 585
R3714 gnd.n1463 gnd.n1462 585
R3715 gnd.n1466 gnd.n1465 585
R3716 gnd.n1464 gnd.n1447 585
R3717 gnd.n1471 gnd.n1470 585
R3718 gnd.n1473 gnd.n1472 585
R3719 gnd.n1476 gnd.n1475 585
R3720 gnd.n1474 gnd.n1445 585
R3721 gnd.n1481 gnd.n1480 585
R3722 gnd.n1485 gnd.n1482 585
R3723 gnd.n1486 gnd.n1423 585
R3724 gnd.n6204 gnd.n6203 585
R3725 gnd.n6197 gnd.n1053 585
R3726 gnd.n6199 gnd.n6198 585
R3727 gnd.n1056 gnd.n1055 585
R3728 gnd.n6169 gnd.n6168 585
R3729 gnd.n6171 gnd.n6170 585
R3730 gnd.n6173 gnd.n6172 585
R3731 gnd.n6175 gnd.n6174 585
R3732 gnd.n6177 gnd.n6176 585
R3733 gnd.n6179 gnd.n6178 585
R3734 gnd.n6181 gnd.n6180 585
R3735 gnd.n6183 gnd.n6182 585
R3736 gnd.n6185 gnd.n6184 585
R3737 gnd.n6188 gnd.n6187 585
R3738 gnd.n6186 gnd.n6158 585
R3739 gnd.n6192 gnd.n6155 585
R3740 gnd.n6194 gnd.n6193 585
R3741 gnd.n6195 gnd.n6194 585
R3742 gnd.n6206 gnd.n6205 585
R3743 gnd.n6205 gnd.n1043 585
R3744 gnd.n1049 gnd.n1041 585
R3745 gnd.n6212 gnd.n1041 585
R3746 gnd.n2311 gnd.n2310 585
R3747 gnd.n2312 gnd.n2311 585
R3748 gnd.n2305 gnd.n1029 585
R3749 gnd.n6218 gnd.n1029 585
R3750 gnd.n2304 gnd.n2303 585
R3751 gnd.n2303 gnd.n1027 585
R3752 gnd.n2302 gnd.n2300 585
R3753 gnd.n2302 gnd.n1018 585
R3754 gnd.n2042 gnd.n1016 585
R3755 gnd.n6226 gnd.n1016 585
R3756 gnd.n1153 gnd.n1152 585
R3757 gnd.n1152 gnd.n1151 585
R3758 gnd.n2036 gnd.n1003 585
R3759 gnd.n6232 gnd.n1003 585
R3760 gnd.n2035 gnd.n2034 585
R3761 gnd.n2034 gnd.n1001 585
R3762 gnd.n2033 gnd.n2031 585
R3763 gnd.n2033 gnd.n992 585
R3764 gnd.n2029 gnd.n990 585
R3765 gnd.n6240 gnd.n990 585
R3766 gnd.n1156 gnd.n1155 585
R3767 gnd.n1155 gnd.n1154 585
R3768 gnd.n2023 gnd.n979 585
R3769 gnd.n6246 gnd.n979 585
R3770 gnd.n2022 gnd.n2021 585
R3771 gnd.n2021 gnd.n977 585
R3772 gnd.n2020 gnd.n1158 585
R3773 gnd.n2020 gnd.n968 585
R3774 gnd.n2019 gnd.n2018 585
R3775 gnd.n2019 gnd.n966 585
R3776 gnd.n1161 gnd.n1160 585
R3777 gnd.n2010 gnd.n1160 585
R3778 gnd.n1938 gnd.n1937 585
R3779 gnd.n1937 gnd.n1165 585
R3780 gnd.n1939 gnd.n1175 585
R3781 gnd.n1996 gnd.n1175 585
R3782 gnd.n1936 gnd.n1935 585
R3783 gnd.n1935 gnd.n1182 585
R3784 gnd.n1934 gnd.n1189 585
R3785 gnd.n1934 gnd.n1181 585
R3786 gnd.n1933 gnd.n1191 585
R3787 gnd.n1933 gnd.n1932 585
R3788 gnd.n1912 gnd.n1190 585
R3789 gnd.n1203 gnd.n1190 585
R3790 gnd.n1911 gnd.n1201 585
R3791 gnd.n1922 gnd.n1201 585
R3792 gnd.n1902 gnd.n1208 585
R3793 gnd.n1903 gnd.n1902 585
R3794 gnd.n1901 gnd.n1900 585
R3795 gnd.n1901 gnd.n1212 585
R3796 gnd.n1899 gnd.n1214 585
R3797 gnd.n1892 gnd.n1214 585
R3798 gnd.n1879 gnd.n1215 585
R3799 gnd.n1880 gnd.n1879 585
R3800 gnd.n1832 gnd.n1228 585
R3801 gnd.n1882 gnd.n1228 585
R3802 gnd.n1834 gnd.n1833 585
R3803 gnd.n1835 gnd.n1834 585
R3804 gnd.n1827 gnd.n1330 585
R3805 gnd.n1330 gnd.n1329 585
R3806 gnd.n1825 gnd.n1824 585
R3807 gnd.n1824 gnd.n1311 585
R3808 gnd.n1822 gnd.n1309 585
R3809 gnd.n1843 gnd.n1309 585
R3810 gnd.n1340 gnd.n1339 585
R3811 gnd.n1339 gnd.n1338 585
R3812 gnd.n1816 gnd.n1299 585
R3813 gnd.n1849 gnd.n1299 585
R3814 gnd.n1815 gnd.n1814 585
R3815 gnd.n1814 gnd.n1813 585
R3816 gnd.n1811 gnd.n1342 585
R3817 gnd.n1811 gnd.n1289 585
R3818 gnd.n1810 gnd.n1809 585
R3819 gnd.n1810 gnd.n1288 585
R3820 gnd.n1345 gnd.n1344 585
R3821 gnd.n1801 gnd.n1344 585
R3822 gnd.n1769 gnd.n1768 585
R3823 gnd.n1768 gnd.n1349 585
R3824 gnd.n1770 gnd.n1358 585
R3825 gnd.n1787 gnd.n1358 585
R3826 gnd.n1767 gnd.n1766 585
R3827 gnd.n1766 gnd.n1364 585
R3828 gnd.n1765 gnd.n1372 585
R3829 gnd.n1765 gnd.n1764 585
R3830 gnd.n1750 gnd.n1373 585
R3831 gnd.n1383 gnd.n1373 585
R3832 gnd.n1749 gnd.n1381 585
R3833 gnd.n1756 gnd.n1381 585
R3834 gnd.n1748 gnd.n1747 585
R3835 gnd.n1747 gnd.n1746 585
R3836 gnd.n1392 gnd.n1389 585
R3837 gnd.n1402 gnd.n1392 585
R3838 gnd.n1738 gnd.n1737 585
R3839 gnd.n1737 gnd.n1736 585
R3840 gnd.n1398 gnd.n1397 585
R3841 gnd.n1411 gnd.n1398 585
R3842 gnd.n1718 gnd.n1409 585
R3843 gnd.n1726 gnd.n1409 585
R3844 gnd.n1717 gnd.n1716 585
R3845 gnd.n1716 gnd.n1715 585
R3846 gnd.n1418 gnd.n1416 585
R3847 gnd.n1427 gnd.n1418 585
R3848 gnd.n1707 gnd.n1706 585
R3849 gnd.n1706 gnd.n1705 585
R3850 gnd.n5912 gnd.n5911 585
R3851 gnd.n5911 gnd.n5910 585
R3852 gnd.n5913 gnd.n2663 585
R3853 gnd.n4256 gnd.n2663 585
R3854 gnd.n5915 gnd.n5914 585
R3855 gnd.n5916 gnd.n5915 585
R3856 gnd.n2648 gnd.n2647 585
R3857 gnd.n4248 gnd.n2648 585
R3858 gnd.n5924 gnd.n5923 585
R3859 gnd.n5923 gnd.n5922 585
R3860 gnd.n5925 gnd.n2642 585
R3861 gnd.n4239 gnd.n2642 585
R3862 gnd.n5927 gnd.n5926 585
R3863 gnd.n5928 gnd.n5927 585
R3864 gnd.n2626 gnd.n2625 585
R3865 gnd.n4231 gnd.n2626 585
R3866 gnd.n5936 gnd.n5935 585
R3867 gnd.n5935 gnd.n5934 585
R3868 gnd.n5937 gnd.n2620 585
R3869 gnd.n4223 gnd.n2620 585
R3870 gnd.n5939 gnd.n5938 585
R3871 gnd.n5940 gnd.n5939 585
R3872 gnd.n2605 gnd.n2604 585
R3873 gnd.n4215 gnd.n2605 585
R3874 gnd.n5948 gnd.n5947 585
R3875 gnd.n5947 gnd.n5946 585
R3876 gnd.n5949 gnd.n2599 585
R3877 gnd.n4207 gnd.n2599 585
R3878 gnd.n5951 gnd.n5950 585
R3879 gnd.n5952 gnd.n5951 585
R3880 gnd.n2583 gnd.n2582 585
R3881 gnd.n4199 gnd.n2583 585
R3882 gnd.n5960 gnd.n5959 585
R3883 gnd.n5959 gnd.n5958 585
R3884 gnd.n5961 gnd.n2577 585
R3885 gnd.n4191 gnd.n2577 585
R3886 gnd.n5963 gnd.n5962 585
R3887 gnd.n5964 gnd.n5963 585
R3888 gnd.n2562 gnd.n2561 585
R3889 gnd.n4183 gnd.n2562 585
R3890 gnd.n5972 gnd.n5971 585
R3891 gnd.n5971 gnd.n5970 585
R3892 gnd.n5973 gnd.n2557 585
R3893 gnd.n4175 gnd.n2557 585
R3894 gnd.n5975 gnd.n5974 585
R3895 gnd.n5976 gnd.n5975 585
R3896 gnd.n2558 gnd.n2541 585
R3897 gnd.n4167 gnd.n2541 585
R3898 gnd.n5984 gnd.n5983 585
R3899 gnd.n5983 gnd.n5982 585
R3900 gnd.n5985 gnd.n2538 585
R3901 gnd.n4159 gnd.n2538 585
R3902 gnd.n5988 gnd.n5987 585
R3903 gnd.n5989 gnd.n5988 585
R3904 gnd.n2539 gnd.n2523 585
R3905 gnd.n4150 gnd.n2523 585
R3906 gnd.n5997 gnd.n5996 585
R3907 gnd.n5996 gnd.n5995 585
R3908 gnd.n5998 gnd.n2519 585
R3909 gnd.n4140 gnd.n2519 585
R3910 gnd.n6000 gnd.n5999 585
R3911 gnd.n6001 gnd.n6000 585
R3912 gnd.n2503 gnd.n2502 585
R3913 gnd.n4132 gnd.n2503 585
R3914 gnd.n6009 gnd.n6008 585
R3915 gnd.n6008 gnd.n6007 585
R3916 gnd.n6010 gnd.n2497 585
R3917 gnd.n4124 gnd.n2497 585
R3918 gnd.n6012 gnd.n6011 585
R3919 gnd.n6013 gnd.n6012 585
R3920 gnd.n2482 gnd.n2481 585
R3921 gnd.n4116 gnd.n2482 585
R3922 gnd.n6021 gnd.n6020 585
R3923 gnd.n6020 gnd.n6019 585
R3924 gnd.n6022 gnd.n2476 585
R3925 gnd.n4108 gnd.n2476 585
R3926 gnd.n6024 gnd.n6023 585
R3927 gnd.n6025 gnd.n6024 585
R3928 gnd.n2460 gnd.n2459 585
R3929 gnd.n4100 gnd.n2460 585
R3930 gnd.n6033 gnd.n6032 585
R3931 gnd.n6032 gnd.n6031 585
R3932 gnd.n6034 gnd.n2454 585
R3933 gnd.n4092 gnd.n2454 585
R3934 gnd.n6036 gnd.n6035 585
R3935 gnd.n6037 gnd.n6036 585
R3936 gnd.n2439 gnd.n2438 585
R3937 gnd.n4084 gnd.n2439 585
R3938 gnd.n6045 gnd.n6044 585
R3939 gnd.n6044 gnd.n6043 585
R3940 gnd.n6046 gnd.n2433 585
R3941 gnd.n4076 gnd.n2433 585
R3942 gnd.n6048 gnd.n6047 585
R3943 gnd.n6049 gnd.n6048 585
R3944 gnd.n2416 gnd.n2415 585
R3945 gnd.n4068 gnd.n2416 585
R3946 gnd.n6057 gnd.n6056 585
R3947 gnd.n6056 gnd.n6055 585
R3948 gnd.n6058 gnd.n2410 585
R3949 gnd.n4059 gnd.n2410 585
R3950 gnd.n6060 gnd.n6059 585
R3951 gnd.n6061 gnd.n6060 585
R3952 gnd.n2411 gnd.n2409 585
R3953 gnd.n2409 gnd.n2405 585
R3954 gnd.n4051 gnd.n4050 585
R3955 gnd.n4052 gnd.n4051 585
R3956 gnd.n4046 gnd.n2354 585
R3957 gnd.n2354 gnd.n2351 585
R3958 gnd.n6146 gnd.n6145 585
R3959 gnd.n6144 gnd.n2353 585
R3960 gnd.n6143 gnd.n2352 585
R3961 gnd.n6148 gnd.n2352 585
R3962 gnd.n6142 gnd.n6141 585
R3963 gnd.n6140 gnd.n6139 585
R3964 gnd.n6138 gnd.n6137 585
R3965 gnd.n6136 gnd.n6135 585
R3966 gnd.n6134 gnd.n6133 585
R3967 gnd.n6132 gnd.n6131 585
R3968 gnd.n6130 gnd.n6129 585
R3969 gnd.n6128 gnd.n6127 585
R3970 gnd.n6126 gnd.n6125 585
R3971 gnd.n6124 gnd.n6123 585
R3972 gnd.n6122 gnd.n6121 585
R3973 gnd.n6120 gnd.n6119 585
R3974 gnd.n6118 gnd.n6117 585
R3975 gnd.n6116 gnd.n6115 585
R3976 gnd.n6114 gnd.n6113 585
R3977 gnd.n6111 gnd.n6110 585
R3978 gnd.n6109 gnd.n6108 585
R3979 gnd.n6107 gnd.n6106 585
R3980 gnd.n6105 gnd.n6104 585
R3981 gnd.n6103 gnd.n6102 585
R3982 gnd.n6101 gnd.n6100 585
R3983 gnd.n6099 gnd.n6098 585
R3984 gnd.n6097 gnd.n6096 585
R3985 gnd.n6095 gnd.n6094 585
R3986 gnd.n6093 gnd.n6092 585
R3987 gnd.n6091 gnd.n6090 585
R3988 gnd.n6089 gnd.n6088 585
R3989 gnd.n6087 gnd.n6086 585
R3990 gnd.n6085 gnd.n6084 585
R3991 gnd.n6083 gnd.n6082 585
R3992 gnd.n6081 gnd.n6080 585
R3993 gnd.n6079 gnd.n6078 585
R3994 gnd.n6077 gnd.n6076 585
R3995 gnd.n6075 gnd.n2393 585
R3996 gnd.n2397 gnd.n2394 585
R3997 gnd.n6071 gnd.n6070 585
R3998 gnd.n3727 gnd.n3726 585
R3999 gnd.n4264 gnd.n4263 585
R4000 gnd.n4266 gnd.n4265 585
R4001 gnd.n4268 gnd.n4267 585
R4002 gnd.n4270 gnd.n4269 585
R4003 gnd.n4272 gnd.n4271 585
R4004 gnd.n4274 gnd.n4273 585
R4005 gnd.n4276 gnd.n4275 585
R4006 gnd.n4278 gnd.n4277 585
R4007 gnd.n4280 gnd.n4279 585
R4008 gnd.n4282 gnd.n4281 585
R4009 gnd.n4284 gnd.n4283 585
R4010 gnd.n4286 gnd.n4285 585
R4011 gnd.n4288 gnd.n4287 585
R4012 gnd.n4290 gnd.n4289 585
R4013 gnd.n4292 gnd.n4291 585
R4014 gnd.n4294 gnd.n4293 585
R4015 gnd.n4296 gnd.n4295 585
R4016 gnd.n4298 gnd.n4297 585
R4017 gnd.n4301 gnd.n4300 585
R4018 gnd.n4299 gnd.n3705 585
R4019 gnd.n4563 gnd.n4562 585
R4020 gnd.n4565 gnd.n4564 585
R4021 gnd.n4567 gnd.n4566 585
R4022 gnd.n4569 gnd.n4568 585
R4023 gnd.n4571 gnd.n4570 585
R4024 gnd.n4573 gnd.n4572 585
R4025 gnd.n4575 gnd.n4574 585
R4026 gnd.n4577 gnd.n4576 585
R4027 gnd.n4579 gnd.n4578 585
R4028 gnd.n4581 gnd.n4580 585
R4029 gnd.n4583 gnd.n4582 585
R4030 gnd.n4585 gnd.n4584 585
R4031 gnd.n4586 gnd.n3686 585
R4032 gnd.n4588 gnd.n4587 585
R4033 gnd.n3687 gnd.n3685 585
R4034 gnd.n3688 gnd.n2668 585
R4035 gnd.n4590 gnd.n2668 585
R4036 gnd.n4259 gnd.n2670 585
R4037 gnd.n5910 gnd.n2670 585
R4038 gnd.n4258 gnd.n4257 585
R4039 gnd.n4257 gnd.n4256 585
R4040 gnd.n3731 gnd.n2661 585
R4041 gnd.n5916 gnd.n2661 585
R4042 gnd.n4247 gnd.n4246 585
R4043 gnd.n4248 gnd.n4247 585
R4044 gnd.n3737 gnd.n2650 585
R4045 gnd.n5922 gnd.n2650 585
R4046 gnd.n4241 gnd.n4240 585
R4047 gnd.n4240 gnd.n4239 585
R4048 gnd.n3739 gnd.n2639 585
R4049 gnd.n5928 gnd.n2639 585
R4050 gnd.n4230 gnd.n4229 585
R4051 gnd.n4231 gnd.n4230 585
R4052 gnd.n3743 gnd.n2628 585
R4053 gnd.n5934 gnd.n2628 585
R4054 gnd.n4225 gnd.n4224 585
R4055 gnd.n4224 gnd.n4223 585
R4056 gnd.n3745 gnd.n2617 585
R4057 gnd.n5940 gnd.n2617 585
R4058 gnd.n4214 gnd.n4213 585
R4059 gnd.n4215 gnd.n4214 585
R4060 gnd.n3750 gnd.n2607 585
R4061 gnd.n5946 gnd.n2607 585
R4062 gnd.n4209 gnd.n4208 585
R4063 gnd.n4208 gnd.n4207 585
R4064 gnd.n3752 gnd.n2596 585
R4065 gnd.n5952 gnd.n2596 585
R4066 gnd.n4198 gnd.n4197 585
R4067 gnd.n4199 gnd.n4198 585
R4068 gnd.n3756 gnd.n2585 585
R4069 gnd.n5958 gnd.n2585 585
R4070 gnd.n4193 gnd.n4192 585
R4071 gnd.n4192 gnd.n4191 585
R4072 gnd.n3758 gnd.n2574 585
R4073 gnd.n5964 gnd.n2574 585
R4074 gnd.n4182 gnd.n4181 585
R4075 gnd.n4183 gnd.n4182 585
R4076 gnd.n3763 gnd.n2564 585
R4077 gnd.n5970 gnd.n2564 585
R4078 gnd.n4177 gnd.n4176 585
R4079 gnd.n4176 gnd.n4175 585
R4080 gnd.n3765 gnd.n2554 585
R4081 gnd.n5976 gnd.n2554 585
R4082 gnd.n4166 gnd.n4165 585
R4083 gnd.n4167 gnd.n4166 585
R4084 gnd.n3769 gnd.n2543 585
R4085 gnd.n5982 gnd.n2543 585
R4086 gnd.n4161 gnd.n4160 585
R4087 gnd.n4160 gnd.n4159 585
R4088 gnd.n3771 gnd.n2535 585
R4089 gnd.n5989 gnd.n2535 585
R4090 gnd.n4149 gnd.n4148 585
R4091 gnd.n4150 gnd.n4149 585
R4092 gnd.n3776 gnd.n2525 585
R4093 gnd.n5995 gnd.n2525 585
R4094 gnd.n4142 gnd.n4141 585
R4095 gnd.n4141 gnd.n4140 585
R4096 gnd.n3778 gnd.n2516 585
R4097 gnd.n6001 gnd.n2516 585
R4098 gnd.n4131 gnd.n4130 585
R4099 gnd.n4132 gnd.n4131 585
R4100 gnd.n3782 gnd.n2505 585
R4101 gnd.n6007 gnd.n2505 585
R4102 gnd.n4126 gnd.n4125 585
R4103 gnd.n4125 gnd.n4124 585
R4104 gnd.n3784 gnd.n2494 585
R4105 gnd.n6013 gnd.n2494 585
R4106 gnd.n4115 gnd.n4114 585
R4107 gnd.n4116 gnd.n4115 585
R4108 gnd.n3789 gnd.n2484 585
R4109 gnd.n6019 gnd.n2484 585
R4110 gnd.n4110 gnd.n4109 585
R4111 gnd.n4109 gnd.n4108 585
R4112 gnd.n3791 gnd.n2473 585
R4113 gnd.n6025 gnd.n2473 585
R4114 gnd.n4099 gnd.n4098 585
R4115 gnd.n4100 gnd.n4099 585
R4116 gnd.n3795 gnd.n2462 585
R4117 gnd.n6031 gnd.n2462 585
R4118 gnd.n4094 gnd.n4093 585
R4119 gnd.n4093 gnd.n4092 585
R4120 gnd.n3797 gnd.n2451 585
R4121 gnd.n6037 gnd.n2451 585
R4122 gnd.n4083 gnd.n4082 585
R4123 gnd.n4084 gnd.n4083 585
R4124 gnd.n3802 gnd.n2441 585
R4125 gnd.n6043 gnd.n2441 585
R4126 gnd.n4078 gnd.n4077 585
R4127 gnd.n4077 gnd.n4076 585
R4128 gnd.n3804 gnd.n2430 585
R4129 gnd.n6049 gnd.n2430 585
R4130 gnd.n4067 gnd.n4066 585
R4131 gnd.n4068 gnd.n4067 585
R4132 gnd.n4063 gnd.n2418 585
R4133 gnd.n6055 gnd.n2418 585
R4134 gnd.n2404 gnd.n2402 585
R4135 gnd.n4059 gnd.n2404 585
R4136 gnd.n6063 gnd.n6062 585
R4137 gnd.n6062 gnd.n6061 585
R4138 gnd.n2403 gnd.n2400 585
R4139 gnd.n2405 gnd.n2403 585
R4140 gnd.n6067 gnd.n2399 585
R4141 gnd.n4052 gnd.n2399 585
R4142 gnd.n6069 gnd.n6068 585
R4143 gnd.n6069 gnd.n2351 585
R4144 gnd.n7441 gnd.n7440 585
R4145 gnd.n7442 gnd.n7441 585
R4146 gnd.n106 gnd.n104 585
R4147 gnd.n104 gnd.n100 585
R4148 gnd.n7361 gnd.n7360 585
R4149 gnd.n7362 gnd.n7361 585
R4150 gnd.n185 gnd.n184 585
R4151 gnd.n184 gnd.n181 585
R4152 gnd.n7356 gnd.n7355 585
R4153 gnd.n7355 gnd.n7354 585
R4154 gnd.n188 gnd.n187 585
R4155 gnd.n359 gnd.n188 585
R4156 gnd.n7270 gnd.n7269 585
R4157 gnd.n7271 gnd.n7270 585
R4158 gnd.n202 gnd.n201 585
R4159 gnd.n7132 gnd.n201 585
R4160 gnd.n7265 gnd.n7264 585
R4161 gnd.n7264 gnd.n7263 585
R4162 gnd.n205 gnd.n204 585
R4163 gnd.n7136 gnd.n205 585
R4164 gnd.n7254 gnd.n7253 585
R4165 gnd.n7255 gnd.n7254 585
R4166 gnd.n218 gnd.n217 585
R4167 gnd.n7143 gnd.n217 585
R4168 gnd.n7249 gnd.n7248 585
R4169 gnd.n7248 gnd.n7247 585
R4170 gnd.n221 gnd.n220 585
R4171 gnd.n342 gnd.n221 585
R4172 gnd.n7238 gnd.n7237 585
R4173 gnd.n7239 gnd.n7238 585
R4174 gnd.n232 gnd.n231 585
R4175 gnd.n7152 gnd.n231 585
R4176 gnd.n7233 gnd.n7232 585
R4177 gnd.n7232 gnd.n7231 585
R4178 gnd.n235 gnd.n234 585
R4179 gnd.n7156 gnd.n235 585
R4180 gnd.n7222 gnd.n7221 585
R4181 gnd.n7223 gnd.n7222 585
R4182 gnd.n248 gnd.n247 585
R4183 gnd.n7163 gnd.n247 585
R4184 gnd.n7217 gnd.n7216 585
R4185 gnd.n7216 gnd.n7215 585
R4186 gnd.n251 gnd.n250 585
R4187 gnd.n310 gnd.n251 585
R4188 gnd.n7206 gnd.n7205 585
R4189 gnd.n7207 gnd.n7206 585
R4190 gnd.n262 gnd.n261 585
R4191 gnd.n7173 gnd.n261 585
R4192 gnd.n7183 gnd.n7182 585
R4193 gnd.n7184 gnd.n7183 585
R4194 gnd.n7181 gnd.n7180 585
R4195 gnd.n7180 gnd.n7179 585
R4196 gnd.n2930 gnd.n293 585
R4197 gnd.n5620 gnd.n293 585
R4198 gnd.n5633 gnd.n2931 585
R4199 gnd.n5633 gnd.n5632 585
R4200 gnd.n5635 gnd.n5634 585
R4201 gnd.n5636 gnd.n5635 585
R4202 gnd.n2929 gnd.n268 585
R4203 gnd.n2929 gnd.n2926 585
R4204 gnd.n272 gnd.n269 585
R4205 gnd.n5609 gnd.n272 585
R4206 gnd.n7202 gnd.n7201 585
R4207 gnd.n7201 gnd.n7200 585
R4208 gnd.n271 gnd.n270 585
R4209 gnd.n5597 gnd.n271 585
R4210 gnd.n5658 gnd.n5657 585
R4211 gnd.n5659 gnd.n5658 585
R4212 gnd.n2906 gnd.n2905 585
R4213 gnd.n2913 gnd.n2905 585
R4214 gnd.n5653 gnd.n5652 585
R4215 gnd.n5652 gnd.n5651 585
R4216 gnd.n2909 gnd.n2908 585
R4217 gnd.n5584 gnd.n2909 585
R4218 gnd.n5568 gnd.n2957 585
R4219 gnd.n2957 gnd.n2956 585
R4220 gnd.n5570 gnd.n5569 585
R4221 gnd.n5571 gnd.n5570 585
R4222 gnd.n2958 gnd.n2955 585
R4223 gnd.n2965 gnd.n2955 585
R4224 gnd.n5563 gnd.n5562 585
R4225 gnd.n5562 gnd.n5561 585
R4226 gnd.n2961 gnd.n2960 585
R4227 gnd.n5541 gnd.n2961 585
R4228 gnd.n5529 gnd.n2985 585
R4229 gnd.n2985 gnd.n2973 585
R4230 gnd.n5531 gnd.n5530 585
R4231 gnd.n5532 gnd.n5531 585
R4232 gnd.n2986 gnd.n2984 585
R4233 gnd.n2994 gnd.n2984 585
R4234 gnd.n5524 gnd.n5523 585
R4235 gnd.n5523 gnd.n5522 585
R4236 gnd.n2989 gnd.n2988 585
R4237 gnd.n5510 gnd.n2989 585
R4238 gnd.n5498 gnd.n3014 585
R4239 gnd.n3014 gnd.n3001 585
R4240 gnd.n5500 gnd.n5499 585
R4241 gnd.n5501 gnd.n5500 585
R4242 gnd.n3015 gnd.n3013 585
R4243 gnd.n3022 gnd.n3013 585
R4244 gnd.n5493 gnd.n5492 585
R4245 gnd.n5492 gnd.n5491 585
R4246 gnd.n3018 gnd.n3017 585
R4247 gnd.n5479 gnd.n3018 585
R4248 gnd.n3040 gnd.n3039 585
R4249 gnd.n3041 gnd.n3040 585
R4250 gnd.n3036 gnd.n2824 585
R4251 gnd.n5694 gnd.n2824 585
R4252 gnd.n5768 gnd.n5767 585
R4253 gnd.n5766 gnd.n2823 585
R4254 gnd.n5765 gnd.n2822 585
R4255 gnd.n5770 gnd.n2822 585
R4256 gnd.n5764 gnd.n5763 585
R4257 gnd.n5762 gnd.n5761 585
R4258 gnd.n5760 gnd.n5759 585
R4259 gnd.n5758 gnd.n5757 585
R4260 gnd.n5756 gnd.n5755 585
R4261 gnd.n5754 gnd.n5753 585
R4262 gnd.n5752 gnd.n5751 585
R4263 gnd.n5750 gnd.n5749 585
R4264 gnd.n5748 gnd.n5747 585
R4265 gnd.n5746 gnd.n5745 585
R4266 gnd.n5744 gnd.n5743 585
R4267 gnd.n5742 gnd.n5741 585
R4268 gnd.n5740 gnd.n5739 585
R4269 gnd.n5737 gnd.n5736 585
R4270 gnd.n5735 gnd.n5734 585
R4271 gnd.n5733 gnd.n5732 585
R4272 gnd.n5731 gnd.n5730 585
R4273 gnd.n5729 gnd.n5728 585
R4274 gnd.n5727 gnd.n5726 585
R4275 gnd.n5725 gnd.n5724 585
R4276 gnd.n5723 gnd.n5722 585
R4277 gnd.n5721 gnd.n5720 585
R4278 gnd.n5719 gnd.n5718 585
R4279 gnd.n5717 gnd.n5716 585
R4280 gnd.n5715 gnd.n5714 585
R4281 gnd.n5713 gnd.n5712 585
R4282 gnd.n5711 gnd.n5710 585
R4283 gnd.n5709 gnd.n5708 585
R4284 gnd.n5707 gnd.n5706 585
R4285 gnd.n5705 gnd.n5704 585
R4286 gnd.n5703 gnd.n5702 585
R4287 gnd.n5701 gnd.n2864 585
R4288 gnd.n2868 gnd.n2865 585
R4289 gnd.n5697 gnd.n5696 585
R4290 gnd.n174 gnd.n173 585
R4291 gnd.n7370 gnd.n169 585
R4292 gnd.n7372 gnd.n7371 585
R4293 gnd.n7374 gnd.n167 585
R4294 gnd.n7376 gnd.n7375 585
R4295 gnd.n7377 gnd.n162 585
R4296 gnd.n7379 gnd.n7378 585
R4297 gnd.n7381 gnd.n160 585
R4298 gnd.n7383 gnd.n7382 585
R4299 gnd.n7384 gnd.n155 585
R4300 gnd.n7386 gnd.n7385 585
R4301 gnd.n7388 gnd.n153 585
R4302 gnd.n7390 gnd.n7389 585
R4303 gnd.n7391 gnd.n148 585
R4304 gnd.n7393 gnd.n7392 585
R4305 gnd.n7395 gnd.n146 585
R4306 gnd.n7397 gnd.n7396 585
R4307 gnd.n7398 gnd.n141 585
R4308 gnd.n7400 gnd.n7399 585
R4309 gnd.n7402 gnd.n139 585
R4310 gnd.n7404 gnd.n7403 585
R4311 gnd.n7408 gnd.n134 585
R4312 gnd.n7410 gnd.n7409 585
R4313 gnd.n7412 gnd.n132 585
R4314 gnd.n7414 gnd.n7413 585
R4315 gnd.n7415 gnd.n127 585
R4316 gnd.n7417 gnd.n7416 585
R4317 gnd.n7419 gnd.n125 585
R4318 gnd.n7421 gnd.n7420 585
R4319 gnd.n7422 gnd.n120 585
R4320 gnd.n7424 gnd.n7423 585
R4321 gnd.n7426 gnd.n118 585
R4322 gnd.n7428 gnd.n7427 585
R4323 gnd.n7429 gnd.n113 585
R4324 gnd.n7431 gnd.n7430 585
R4325 gnd.n7433 gnd.n111 585
R4326 gnd.n7435 gnd.n7434 585
R4327 gnd.n7436 gnd.n109 585
R4328 gnd.n7437 gnd.n105 585
R4329 gnd.n105 gnd.n102 585
R4330 gnd.n7366 gnd.n101 585
R4331 gnd.n7442 gnd.n101 585
R4332 gnd.n7365 gnd.n7364 585
R4333 gnd.n7364 gnd.n100 585
R4334 gnd.n7363 gnd.n178 585
R4335 gnd.n7363 gnd.n7362 585
R4336 gnd.n357 gnd.n179 585
R4337 gnd.n181 gnd.n179 585
R4338 gnd.n358 gnd.n190 585
R4339 gnd.n7354 gnd.n190 585
R4340 gnd.n361 gnd.n360 585
R4341 gnd.n360 gnd.n359 585
R4342 gnd.n362 gnd.n199 585
R4343 gnd.n7271 gnd.n199 585
R4344 gnd.n7134 gnd.n7133 585
R4345 gnd.n7133 gnd.n7132 585
R4346 gnd.n7135 gnd.n207 585
R4347 gnd.n7263 gnd.n207 585
R4348 gnd.n7138 gnd.n7137 585
R4349 gnd.n7137 gnd.n7136 585
R4350 gnd.n7139 gnd.n215 585
R4351 gnd.n7255 gnd.n215 585
R4352 gnd.n7141 gnd.n7140 585
R4353 gnd.n7143 gnd.n7141 585
R4354 gnd.n340 gnd.n223 585
R4355 gnd.n7247 gnd.n223 585
R4356 gnd.n344 gnd.n343 585
R4357 gnd.n343 gnd.n342 585
R4358 gnd.n320 gnd.n229 585
R4359 gnd.n7239 gnd.n229 585
R4360 gnd.n7154 gnd.n7153 585
R4361 gnd.n7153 gnd.n7152 585
R4362 gnd.n7155 gnd.n237 585
R4363 gnd.n7231 gnd.n237 585
R4364 gnd.n7158 gnd.n7157 585
R4365 gnd.n7157 gnd.n7156 585
R4366 gnd.n7159 gnd.n245 585
R4367 gnd.n7223 gnd.n245 585
R4368 gnd.n7161 gnd.n7160 585
R4369 gnd.n7163 gnd.n7161 585
R4370 gnd.n308 gnd.n253 585
R4371 gnd.n7215 gnd.n253 585
R4372 gnd.n312 gnd.n311 585
R4373 gnd.n311 gnd.n310 585
R4374 gnd.n300 gnd.n259 585
R4375 gnd.n7207 gnd.n259 585
R4376 gnd.n7175 gnd.n7174 585
R4377 gnd.n7174 gnd.n7173 585
R4378 gnd.n7176 gnd.n291 585
R4379 gnd.n7184 gnd.n291 585
R4380 gnd.n7178 gnd.n7177 585
R4381 gnd.n7179 gnd.n7178 585
R4382 gnd.n295 gnd.n294 585
R4383 gnd.n5620 gnd.n294 585
R4384 gnd.n5617 gnd.n5616 585
R4385 gnd.n5632 gnd.n5617 585
R4386 gnd.n2933 gnd.n2927 585
R4387 gnd.n5636 gnd.n2927 585
R4388 gnd.n5612 gnd.n5611 585
R4389 gnd.n5611 gnd.n2926 585
R4390 gnd.n5610 gnd.n2935 585
R4391 gnd.n5610 gnd.n5609 585
R4392 gnd.n5594 gnd.n274 585
R4393 gnd.n7200 gnd.n274 585
R4394 gnd.n5596 gnd.n5595 585
R4395 gnd.n5597 gnd.n5596 585
R4396 gnd.n2941 gnd.n2902 585
R4397 gnd.n5659 gnd.n2902 585
R4398 gnd.n5589 gnd.n5588 585
R4399 gnd.n5588 gnd.n2913 585
R4400 gnd.n5587 gnd.n2911 585
R4401 gnd.n5651 gnd.n2911 585
R4402 gnd.n5586 gnd.n5585 585
R4403 gnd.n5585 gnd.n5584 585
R4404 gnd.n2945 gnd.n2943 585
R4405 gnd.n2956 gnd.n2945 585
R4406 gnd.n3059 gnd.n2953 585
R4407 gnd.n5571 gnd.n2953 585
R4408 gnd.n3061 gnd.n3060 585
R4409 gnd.n3060 gnd.n2965 585
R4410 gnd.n3062 gnd.n2963 585
R4411 gnd.n5561 gnd.n2963 585
R4412 gnd.n3063 gnd.n2974 585
R4413 gnd.n5541 gnd.n2974 585
R4414 gnd.n3065 gnd.n3064 585
R4415 gnd.n3064 gnd.n2973 585
R4416 gnd.n3066 gnd.n2982 585
R4417 gnd.n5532 gnd.n2982 585
R4418 gnd.n3068 gnd.n3067 585
R4419 gnd.n3067 gnd.n2994 585
R4420 gnd.n3069 gnd.n2991 585
R4421 gnd.n5522 gnd.n2991 585
R4422 gnd.n3070 gnd.n3002 585
R4423 gnd.n5510 gnd.n3002 585
R4424 gnd.n3072 gnd.n3071 585
R4425 gnd.n3071 gnd.n3001 585
R4426 gnd.n3073 gnd.n3010 585
R4427 gnd.n5501 gnd.n3010 585
R4428 gnd.n3075 gnd.n3074 585
R4429 gnd.n3074 gnd.n3022 585
R4430 gnd.n3076 gnd.n3020 585
R4431 gnd.n5491 gnd.n3020 585
R4432 gnd.n3078 gnd.n3077 585
R4433 gnd.n5479 gnd.n3078 585
R4434 gnd.n3042 gnd.n2870 585
R4435 gnd.n3041 gnd.n2870 585
R4436 gnd.n5695 gnd.n2871 585
R4437 gnd.n5695 gnd.n5694 585
R4438 gnd.n5310 gnd.n5309 585
R4439 gnd.n5309 gnd.n3262 585
R4440 gnd.n5311 gnd.n5111 585
R4441 gnd.n5111 gnd.n5110 585
R4442 gnd.n5313 gnd.n5312 585
R4443 gnd.n5314 gnd.n5313 585
R4444 gnd.n5113 gnd.n5109 585
R4445 gnd.n5109 gnd.t143 585
R4446 gnd.n5112 gnd.n5101 585
R4447 gnd.n5101 gnd.n3268 585
R4448 gnd.n5323 gnd.n5100 585
R4449 gnd.n5323 gnd.n5322 585
R4450 gnd.n5325 gnd.n5324 585
R4451 gnd.n5324 gnd.n3275 585
R4452 gnd.n5326 gnd.n5098 585
R4453 gnd.n5098 gnd.n3274 585
R4454 gnd.n5328 gnd.n5327 585
R4455 gnd.n5329 gnd.n5328 585
R4456 gnd.n5099 gnd.n5097 585
R4457 gnd.n5097 gnd.n3281 585
R4458 gnd.n5089 gnd.n5088 585
R4459 gnd.n5335 gnd.n5089 585
R4460 gnd.n5339 gnd.n5338 585
R4461 gnd.n5338 gnd.n5337 585
R4462 gnd.n5340 gnd.n3304 585
R4463 gnd.n3304 gnd.n3287 585
R4464 gnd.n5342 gnd.n5341 585
R4465 gnd.n5343 gnd.n5342 585
R4466 gnd.n5087 gnd.n3303 585
R4467 gnd.n3303 gnd.n3294 585
R4468 gnd.n5086 gnd.n3293 585
R4469 gnd.n5349 gnd.n3293 585
R4470 gnd.n5085 gnd.n5084 585
R4471 gnd.n5084 gnd.n5083 585
R4472 gnd.n3306 gnd.n3305 585
R4473 gnd.n3307 gnd.n3306 585
R4474 gnd.n4959 gnd.n4950 585
R4475 gnd.n4959 gnd.n4958 585
R4476 gnd.n4961 gnd.n4960 585
R4477 gnd.n4960 gnd.n3316 585
R4478 gnd.n4962 gnd.n4947 585
R4479 gnd.n4947 gnd.n3314 585
R4480 gnd.n4964 gnd.n4963 585
R4481 gnd.n4965 gnd.n4964 585
R4482 gnd.n4949 gnd.n4946 585
R4483 gnd.n4946 gnd.n3323 585
R4484 gnd.n4948 gnd.n4936 585
R4485 gnd.n4971 gnd.n4936 585
R4486 gnd.n4974 gnd.n4935 585
R4487 gnd.n4974 gnd.n4973 585
R4488 gnd.n4976 gnd.n4975 585
R4489 gnd.n4975 gnd.n3331 585
R4490 gnd.n4977 gnd.n4932 585
R4491 gnd.n4932 gnd.n3329 585
R4492 gnd.n4979 gnd.n4978 585
R4493 gnd.n4980 gnd.n4979 585
R4494 gnd.n4934 gnd.n4931 585
R4495 gnd.n4931 gnd.n3338 585
R4496 gnd.n4933 gnd.n4924 585
R4497 gnd.n4924 gnd.n3337 585
R4498 gnd.n4989 gnd.n4923 585
R4499 gnd.n4989 gnd.n4988 585
R4500 gnd.n4991 gnd.n4990 585
R4501 gnd.n4990 gnd.n3346 585
R4502 gnd.n4992 gnd.n4921 585
R4503 gnd.n4921 gnd.n3344 585
R4504 gnd.n4994 gnd.n4993 585
R4505 gnd.n4995 gnd.n4994 585
R4506 gnd.n4922 gnd.n4920 585
R4507 gnd.n4920 gnd.n3352 585
R4508 gnd.n4913 gnd.n4912 585
R4509 gnd.n5001 gnd.n4913 585
R4510 gnd.n5005 gnd.n5004 585
R4511 gnd.n5004 gnd.n5003 585
R4512 gnd.n5006 gnd.n3376 585
R4513 gnd.n3376 gnd.n3359 585
R4514 gnd.n5008 gnd.n5007 585
R4515 gnd.n5009 gnd.n5008 585
R4516 gnd.n4911 gnd.n3375 585
R4517 gnd.n3375 gnd.n3367 585
R4518 gnd.n4910 gnd.n3366 585
R4519 gnd.n5015 gnd.n3366 585
R4520 gnd.n4909 gnd.n4908 585
R4521 gnd.n4908 gnd.n3365 585
R4522 gnd.n4907 gnd.n3377 585
R4523 gnd.n4907 gnd.n4906 585
R4524 gnd.n4764 gnd.n3378 585
R4525 gnd.n4779 gnd.n3378 585
R4526 gnd.n4766 gnd.n4765 585
R4527 gnd.n4766 gnd.n3387 585
R4528 gnd.n4767 gnd.n4763 585
R4529 gnd.n4767 gnd.n3386 585
R4530 gnd.n4789 gnd.n4788 585
R4531 gnd.n4788 gnd.n4787 585
R4532 gnd.n4790 gnd.n4762 585
R4533 gnd.n4762 gnd.n3394 585
R4534 gnd.n4792 gnd.n4791 585
R4535 gnd.n4793 gnd.n4792 585
R4536 gnd.n4757 gnd.n4756 585
R4537 gnd.n4795 gnd.n4757 585
R4538 gnd.n4798 gnd.n4797 585
R4539 gnd.n4797 gnd.n4796 585
R4540 gnd.n4799 gnd.n4753 585
R4541 gnd.n4753 gnd.n3400 585
R4542 gnd.n4801 gnd.n4800 585
R4543 gnd.n4802 gnd.n4801 585
R4544 gnd.n4755 gnd.n4752 585
R4545 gnd.n4752 gnd.n3407 585
R4546 gnd.n4754 gnd.n4745 585
R4547 gnd.n4745 gnd.n3406 585
R4548 gnd.n4812 gnd.n4744 585
R4549 gnd.n4812 gnd.n4811 585
R4550 gnd.n4814 gnd.n4813 585
R4551 gnd.n4813 gnd.n3413 585
R4552 gnd.n4815 gnd.n4742 585
R4553 gnd.n4742 gnd.n4741 585
R4554 gnd.n4817 gnd.n4816 585
R4555 gnd.n4818 gnd.n4817 585
R4556 gnd.n4743 gnd.n4740 585
R4557 gnd.n4740 gnd.n3419 585
R4558 gnd.n4732 gnd.n4731 585
R4559 gnd.n4824 gnd.n4732 585
R4560 gnd.n4828 gnd.n4827 585
R4561 gnd.n4827 gnd.n4826 585
R4562 gnd.n4829 gnd.n3442 585
R4563 gnd.n3442 gnd.n3425 585
R4564 gnd.n4831 gnd.n4830 585
R4565 gnd.n4832 gnd.n4831 585
R4566 gnd.n4730 gnd.n3441 585
R4567 gnd.n3441 gnd.n3440 585
R4568 gnd.n4729 gnd.n3432 585
R4569 gnd.n4838 gnd.n3432 585
R4570 gnd.n4728 gnd.n4727 585
R4571 gnd.n4727 gnd.n3431 585
R4572 gnd.n4726 gnd.n3443 585
R4573 gnd.n4726 gnd.n4725 585
R4574 gnd.n4450 gnd.n3444 585
R4575 gnd.n4461 gnd.n3444 585
R4576 gnd.n4451 gnd.n4449 585
R4577 gnd.n4449 gnd.n3453 585
R4578 gnd.n4453 gnd.n4452 585
R4579 gnd.n4467 gnd.n4453 585
R4580 gnd.n4470 gnd.n4448 585
R4581 gnd.n4470 gnd.n4469 585
R4582 gnd.n4472 gnd.n4471 585
R4583 gnd.n4471 gnd.n3461 585
R4584 gnd.n4473 gnd.n4445 585
R4585 gnd.n4445 gnd.n4444 585
R4586 gnd.n4475 gnd.n4474 585
R4587 gnd.n4476 gnd.n4475 585
R4588 gnd.n4447 gnd.n4443 585
R4589 gnd.n4443 gnd.n3467 585
R4590 gnd.n4446 gnd.n4433 585
R4591 gnd.n4482 gnd.n4433 585
R4592 gnd.n4485 gnd.n4432 585
R4593 gnd.n4485 gnd.n4484 585
R4594 gnd.n4487 gnd.n4486 585
R4595 gnd.n4486 gnd.n3475 585
R4596 gnd.n4488 gnd.n4329 585
R4597 gnd.n4329 gnd.n3473 585
R4598 gnd.n4490 gnd.n4489 585
R4599 gnd.n4491 gnd.n4490 585
R4600 gnd.n4430 gnd.n4328 585
R4601 gnd.n4429 gnd.n4428 585
R4602 gnd.n4426 gnd.n4350 585
R4603 gnd.n4426 gnd.n3481 585
R4604 gnd.n4425 gnd.n4424 585
R4605 gnd.n4423 gnd.n4422 585
R4606 gnd.n4421 gnd.n4352 585
R4607 gnd.n4419 gnd.n4418 585
R4608 gnd.n4417 gnd.n4353 585
R4609 gnd.n4416 gnd.n4415 585
R4610 gnd.n4413 gnd.n4354 585
R4611 gnd.n4411 gnd.n4410 585
R4612 gnd.n4409 gnd.n4355 585
R4613 gnd.n4408 gnd.n4407 585
R4614 gnd.n4405 gnd.n4356 585
R4615 gnd.n4403 gnd.n4402 585
R4616 gnd.n4401 gnd.n4357 585
R4617 gnd.n4400 gnd.n4399 585
R4618 gnd.n4397 gnd.n4358 585
R4619 gnd.n4395 gnd.n4394 585
R4620 gnd.n4393 gnd.n4359 585
R4621 gnd.n4392 gnd.n4391 585
R4622 gnd.n4389 gnd.n4360 585
R4623 gnd.n4387 gnd.n4386 585
R4624 gnd.n4385 gnd.n4361 585
R4625 gnd.n4384 gnd.n4383 585
R4626 gnd.n4381 gnd.n4362 585
R4627 gnd.n4379 gnd.n4378 585
R4628 gnd.n4377 gnd.n4363 585
R4629 gnd.n4376 gnd.n4375 585
R4630 gnd.n4373 gnd.n4372 585
R4631 gnd.n4371 gnd.n4370 585
R4632 gnd.n4369 gnd.n4306 585
R4633 gnd.n4560 gnd.n4559 585
R4634 gnd.n4557 gnd.n4305 585
R4635 gnd.n4555 gnd.n4554 585
R4636 gnd.n4553 gnd.n4308 585
R4637 gnd.n4551 gnd.n4550 585
R4638 gnd.n4548 gnd.n4311 585
R4639 gnd.n4546 gnd.n4545 585
R4640 gnd.n4544 gnd.n4312 585
R4641 gnd.n4543 gnd.n4542 585
R4642 gnd.n4540 gnd.n4313 585
R4643 gnd.n4538 gnd.n4537 585
R4644 gnd.n4536 gnd.n4314 585
R4645 gnd.n4535 gnd.n4534 585
R4646 gnd.n4532 gnd.n4315 585
R4647 gnd.n4530 gnd.n4529 585
R4648 gnd.n4528 gnd.n4316 585
R4649 gnd.n4527 gnd.n4526 585
R4650 gnd.n4524 gnd.n4317 585
R4651 gnd.n4522 gnd.n4521 585
R4652 gnd.n4520 gnd.n4318 585
R4653 gnd.n4519 gnd.n4518 585
R4654 gnd.n4516 gnd.n4319 585
R4655 gnd.n4514 gnd.n4513 585
R4656 gnd.n4512 gnd.n4320 585
R4657 gnd.n4511 gnd.n4510 585
R4658 gnd.n4508 gnd.n4321 585
R4659 gnd.n4506 gnd.n4505 585
R4660 gnd.n4504 gnd.n4322 585
R4661 gnd.n4503 gnd.n4502 585
R4662 gnd.n4500 gnd.n4323 585
R4663 gnd.n4498 gnd.n4497 585
R4664 gnd.n4496 gnd.n4324 585
R4665 gnd.n4495 gnd.n4494 585
R4666 gnd.n5193 gnd.n5192 585
R4667 gnd.n5194 gnd.n5187 585
R4668 gnd.n5196 gnd.n5195 585
R4669 gnd.n5198 gnd.n5185 585
R4670 gnd.n5200 gnd.n5199 585
R4671 gnd.n5201 gnd.n5184 585
R4672 gnd.n5203 gnd.n5202 585
R4673 gnd.n5205 gnd.n5182 585
R4674 gnd.n5207 gnd.n5206 585
R4675 gnd.n5208 gnd.n5181 585
R4676 gnd.n5210 gnd.n5209 585
R4677 gnd.n5212 gnd.n5179 585
R4678 gnd.n5214 gnd.n5213 585
R4679 gnd.n5215 gnd.n5178 585
R4680 gnd.n5217 gnd.n5216 585
R4681 gnd.n5219 gnd.n5176 585
R4682 gnd.n5221 gnd.n5220 585
R4683 gnd.n5222 gnd.n5175 585
R4684 gnd.n5224 gnd.n5223 585
R4685 gnd.n5226 gnd.n5173 585
R4686 gnd.n5228 gnd.n5227 585
R4687 gnd.n5229 gnd.n5172 585
R4688 gnd.n5231 gnd.n5230 585
R4689 gnd.n5233 gnd.n5170 585
R4690 gnd.n5235 gnd.n5234 585
R4691 gnd.n5236 gnd.n5169 585
R4692 gnd.n5238 gnd.n5237 585
R4693 gnd.n5240 gnd.n5167 585
R4694 gnd.n5242 gnd.n5241 585
R4695 gnd.n5244 gnd.n5164 585
R4696 gnd.n5246 gnd.n5245 585
R4697 gnd.n5248 gnd.n5163 585
R4698 gnd.n5249 gnd.n5136 585
R4699 gnd.n5252 gnd.n2841 585
R4700 gnd.n5254 gnd.n5253 585
R4701 gnd.n5255 gnd.n5158 585
R4702 gnd.n5257 gnd.n5256 585
R4703 gnd.n5259 gnd.n5156 585
R4704 gnd.n5261 gnd.n5260 585
R4705 gnd.n5262 gnd.n5155 585
R4706 gnd.n5264 gnd.n5263 585
R4707 gnd.n5266 gnd.n5153 585
R4708 gnd.n5268 gnd.n5267 585
R4709 gnd.n5269 gnd.n5152 585
R4710 gnd.n5271 gnd.n5270 585
R4711 gnd.n5273 gnd.n5150 585
R4712 gnd.n5275 gnd.n5274 585
R4713 gnd.n5276 gnd.n5149 585
R4714 gnd.n5278 gnd.n5277 585
R4715 gnd.n5280 gnd.n5147 585
R4716 gnd.n5282 gnd.n5281 585
R4717 gnd.n5283 gnd.n5146 585
R4718 gnd.n5285 gnd.n5284 585
R4719 gnd.n5287 gnd.n5144 585
R4720 gnd.n5289 gnd.n5288 585
R4721 gnd.n5290 gnd.n5143 585
R4722 gnd.n5292 gnd.n5291 585
R4723 gnd.n5294 gnd.n5141 585
R4724 gnd.n5296 gnd.n5295 585
R4725 gnd.n5297 gnd.n5140 585
R4726 gnd.n5299 gnd.n5298 585
R4727 gnd.n5301 gnd.n5138 585
R4728 gnd.n5303 gnd.n5302 585
R4729 gnd.n5304 gnd.n5137 585
R4730 gnd.n5306 gnd.n5305 585
R4731 gnd.n5308 gnd.n5134 585
R4732 gnd.n5191 gnd.n5189 585
R4733 gnd.n5191 gnd.n3262 585
R4734 gnd.n5188 gnd.n5106 585
R4735 gnd.n5110 gnd.n5106 585
R4736 gnd.n5315 gnd.n5105 585
R4737 gnd.n5315 gnd.n5314 585
R4738 gnd.n5317 gnd.n5316 585
R4739 gnd.n5316 gnd.t143 585
R4740 gnd.n5318 gnd.n5103 585
R4741 gnd.n5103 gnd.n3268 585
R4742 gnd.n5320 gnd.n5319 585
R4743 gnd.n5322 gnd.n5320 585
R4744 gnd.n5104 gnd.n5102 585
R4745 gnd.n5102 gnd.n3275 585
R4746 gnd.n5094 gnd.n5093 585
R4747 gnd.n5094 gnd.n3274 585
R4748 gnd.n5331 gnd.n5330 585
R4749 gnd.n5330 gnd.n5329 585
R4750 gnd.n5332 gnd.n5091 585
R4751 gnd.n5091 gnd.n3281 585
R4752 gnd.n5334 gnd.n5333 585
R4753 gnd.n5335 gnd.n5334 585
R4754 gnd.n5092 gnd.n5090 585
R4755 gnd.n5337 gnd.n5090 585
R4756 gnd.n3300 gnd.n3299 585
R4757 gnd.n3300 gnd.n3287 585
R4758 gnd.n5345 gnd.n5344 585
R4759 gnd.n5344 gnd.n5343 585
R4760 gnd.n5346 gnd.n3297 585
R4761 gnd.n3297 gnd.n3294 585
R4762 gnd.n5348 gnd.n5347 585
R4763 gnd.n5349 gnd.n5348 585
R4764 gnd.n3298 gnd.n3296 585
R4765 gnd.n5083 gnd.n3296 585
R4766 gnd.n4954 gnd.n4952 585
R4767 gnd.n4952 gnd.n3307 585
R4768 gnd.n4956 gnd.n4955 585
R4769 gnd.n4958 gnd.n4956 585
R4770 gnd.n4953 gnd.n4951 585
R4771 gnd.n4951 gnd.n3316 585
R4772 gnd.n4944 gnd.n4943 585
R4773 gnd.n4944 gnd.n3314 585
R4774 gnd.n4967 gnd.n4966 585
R4775 gnd.n4966 gnd.n4965 585
R4776 gnd.n4968 gnd.n4938 585
R4777 gnd.n4938 gnd.n3323 585
R4778 gnd.n4970 gnd.n4969 585
R4779 gnd.n4971 gnd.n4970 585
R4780 gnd.n4942 gnd.n4937 585
R4781 gnd.n4973 gnd.n4937 585
R4782 gnd.n4941 gnd.n4940 585
R4783 gnd.n4940 gnd.n3331 585
R4784 gnd.n4939 gnd.n4929 585
R4785 gnd.n4929 gnd.n3329 585
R4786 gnd.n4981 gnd.n4928 585
R4787 gnd.n4981 gnd.n4980 585
R4788 gnd.n4983 gnd.n4982 585
R4789 gnd.n4982 gnd.n3338 585
R4790 gnd.n4984 gnd.n4926 585
R4791 gnd.n4926 gnd.n3337 585
R4792 gnd.n4986 gnd.n4985 585
R4793 gnd.n4988 gnd.n4986 585
R4794 gnd.n4927 gnd.n4925 585
R4795 gnd.n4925 gnd.n3346 585
R4796 gnd.n4918 gnd.n4917 585
R4797 gnd.n4918 gnd.n3344 585
R4798 gnd.n4997 gnd.n4996 585
R4799 gnd.n4996 gnd.n4995 585
R4800 gnd.n4998 gnd.n4915 585
R4801 gnd.n4915 gnd.n3352 585
R4802 gnd.n5000 gnd.n4999 585
R4803 gnd.n5001 gnd.n5000 585
R4804 gnd.n4916 gnd.n4914 585
R4805 gnd.n5003 gnd.n4914 585
R4806 gnd.n3373 gnd.n3372 585
R4807 gnd.n3373 gnd.n3359 585
R4808 gnd.n5011 gnd.n5010 585
R4809 gnd.n5010 gnd.n5009 585
R4810 gnd.n5012 gnd.n3370 585
R4811 gnd.n3370 gnd.n3367 585
R4812 gnd.n5014 gnd.n5013 585
R4813 gnd.n5015 gnd.n5014 585
R4814 gnd.n3371 gnd.n3369 585
R4815 gnd.n3369 gnd.n3365 585
R4816 gnd.n4775 gnd.n3379 585
R4817 gnd.n4906 gnd.n3379 585
R4818 gnd.n4780 gnd.n4776 585
R4819 gnd.n4780 gnd.n4779 585
R4820 gnd.n4782 gnd.n4781 585
R4821 gnd.n4781 gnd.n3387 585
R4822 gnd.n4783 gnd.n4769 585
R4823 gnd.n4769 gnd.n3386 585
R4824 gnd.n4785 gnd.n4784 585
R4825 gnd.n4787 gnd.n4785 585
R4826 gnd.n4774 gnd.n4768 585
R4827 gnd.n4768 gnd.n3394 585
R4828 gnd.n4773 gnd.n4761 585
R4829 gnd.n4793 gnd.n4761 585
R4830 gnd.n4772 gnd.n4759 585
R4831 gnd.n4795 gnd.n4759 585
R4832 gnd.n4771 gnd.n4758 585
R4833 gnd.n4796 gnd.n4758 585
R4834 gnd.n4770 gnd.n4750 585
R4835 gnd.n4750 gnd.n3400 585
R4836 gnd.n4803 gnd.n4749 585
R4837 gnd.n4803 gnd.n4802 585
R4838 gnd.n4805 gnd.n4804 585
R4839 gnd.n4804 gnd.n3407 585
R4840 gnd.n4806 gnd.n4747 585
R4841 gnd.n4747 gnd.n3406 585
R4842 gnd.n4808 gnd.n4807 585
R4843 gnd.n4811 gnd.n4808 585
R4844 gnd.n4748 gnd.n4746 585
R4845 gnd.n4746 gnd.n3413 585
R4846 gnd.n4738 gnd.n4737 585
R4847 gnd.n4741 gnd.n4738 585
R4848 gnd.n4820 gnd.n4819 585
R4849 gnd.n4819 gnd.n4818 585
R4850 gnd.n4821 gnd.n4735 585
R4851 gnd.n4735 gnd.n3419 585
R4852 gnd.n4823 gnd.n4822 585
R4853 gnd.n4824 gnd.n4823 585
R4854 gnd.n4736 gnd.n4733 585
R4855 gnd.n4826 gnd.n4733 585
R4856 gnd.n3438 gnd.n3437 585
R4857 gnd.n3438 gnd.n3425 585
R4858 gnd.n4834 gnd.n4833 585
R4859 gnd.n4833 gnd.n4832 585
R4860 gnd.n4835 gnd.n3435 585
R4861 gnd.n3440 gnd.n3435 585
R4862 gnd.n4837 gnd.n4836 585
R4863 gnd.n4838 gnd.n4837 585
R4864 gnd.n3436 gnd.n3434 585
R4865 gnd.n3434 gnd.n3431 585
R4866 gnd.n4459 gnd.n3445 585
R4867 gnd.n4725 gnd.n3445 585
R4868 gnd.n4463 gnd.n4462 585
R4869 gnd.n4462 gnd.n4461 585
R4870 gnd.n4464 gnd.n4455 585
R4871 gnd.n4455 gnd.n3453 585
R4872 gnd.n4466 gnd.n4465 585
R4873 gnd.n4467 gnd.n4466 585
R4874 gnd.n4458 gnd.n4454 585
R4875 gnd.n4469 gnd.n4454 585
R4876 gnd.n4457 gnd.n4456 585
R4877 gnd.n4456 gnd.n3461 585
R4878 gnd.n4441 gnd.n4440 585
R4879 gnd.n4444 gnd.n4441 585
R4880 gnd.n4478 gnd.n4477 585
R4881 gnd.n4477 gnd.n4476 585
R4882 gnd.n4479 gnd.n4435 585
R4883 gnd.n4435 gnd.n3467 585
R4884 gnd.n4481 gnd.n4480 585
R4885 gnd.n4482 gnd.n4481 585
R4886 gnd.n4439 gnd.n4434 585
R4887 gnd.n4484 gnd.n4434 585
R4888 gnd.n4438 gnd.n4437 585
R4889 gnd.n4437 gnd.n3475 585
R4890 gnd.n4436 gnd.n4326 585
R4891 gnd.n4326 gnd.n3473 585
R4892 gnd.n4492 gnd.n4325 585
R4893 gnd.n4492 gnd.n4491 585
R4894 gnd.n3972 gnd.n3971 585
R4895 gnd.n3973 gnd.n3972 585
R4896 gnd.n7124 gnd.n7123 585
R4897 gnd.n7124 gnd.n182 585
R4898 gnd.n7125 gnd.n380 585
R4899 gnd.n7125 gnd.n191 585
R4900 gnd.n7127 gnd.n7126 585
R4901 gnd.n7126 gnd.n189 585
R4902 gnd.n7128 gnd.n365 585
R4903 gnd.n365 gnd.n200 585
R4904 gnd.n7130 gnd.n7129 585
R4905 gnd.n7131 gnd.n7130 585
R4906 gnd.n366 gnd.n364 585
R4907 gnd.n364 gnd.n208 585
R4908 gnd.n374 gnd.n373 585
R4909 gnd.n373 gnd.n206 585
R4910 gnd.n372 gnd.n371 585
R4911 gnd.n372 gnd.n216 585
R4912 gnd.n370 gnd.n339 585
R4913 gnd.n339 gnd.n214 585
R4914 gnd.n7145 gnd.n338 585
R4915 gnd.n7145 gnd.n7144 585
R4916 gnd.n7147 gnd.n7146 585
R4917 gnd.n7146 gnd.n222 585
R4918 gnd.n7148 gnd.n323 585
R4919 gnd.n323 gnd.n230 585
R4920 gnd.n7150 gnd.n7149 585
R4921 gnd.n7151 gnd.n7150 585
R4922 gnd.n324 gnd.n322 585
R4923 gnd.n322 gnd.n238 585
R4924 gnd.n332 gnd.n331 585
R4925 gnd.n331 gnd.n236 585
R4926 gnd.n330 gnd.n329 585
R4927 gnd.n330 gnd.n246 585
R4928 gnd.n328 gnd.n307 585
R4929 gnd.n307 gnd.n244 585
R4930 gnd.n7165 gnd.n306 585
R4931 gnd.n7165 gnd.n7164 585
R4932 gnd.n7167 gnd.n7166 585
R4933 gnd.n7166 gnd.n252 585
R4934 gnd.n7168 gnd.n303 585
R4935 gnd.n303 gnd.n260 585
R4936 gnd.n7171 gnd.n7170 585
R4937 gnd.n7172 gnd.n7171 585
R4938 gnd.n304 gnd.n302 585
R4939 gnd.n302 gnd.n292 585
R4940 gnd.n5626 gnd.n5625 585
R4941 gnd.n5625 gnd.n290 585
R4942 gnd.n5627 gnd.n5622 585
R4943 gnd.n5622 gnd.n5621 585
R4944 gnd.n5630 gnd.n5629 585
R4945 gnd.n5631 gnd.n5630 585
R4946 gnd.n5623 gnd.n2925 585
R4947 gnd.n2932 gnd.n2925 585
R4948 gnd.n5639 gnd.n5638 585
R4949 gnd.n5638 gnd.n5637 585
R4950 gnd.n5640 gnd.n2923 585
R4951 gnd.n5608 gnd.n2923 585
R4952 gnd.n5643 gnd.n5642 585
R4953 gnd.n5643 gnd.n276 585
R4954 gnd.n5644 gnd.n2922 585
R4955 gnd.n5644 gnd.n273 585
R4956 gnd.n5646 gnd.n5645 585
R4957 gnd.n5645 gnd.n2904 585
R4958 gnd.n5647 gnd.n2916 585
R4959 gnd.n2916 gnd.n2915 585
R4960 gnd.n5649 gnd.n5648 585
R4961 gnd.n5650 gnd.n5649 585
R4962 gnd.n2917 gnd.n2914 585
R4963 gnd.n2914 gnd.n2910 585
R4964 gnd.n5553 gnd.n5552 585
R4965 gnd.n5553 gnd.n2946 585
R4966 gnd.n5555 gnd.n5554 585
R4967 gnd.n5554 gnd.n2954 585
R4968 gnd.n5556 gnd.n2968 585
R4969 gnd.n2968 gnd.n2967 585
R4970 gnd.n5558 gnd.n5557 585
R4971 gnd.n5559 gnd.n5558 585
R4972 gnd.n2969 gnd.n2966 585
R4973 gnd.n2966 gnd.n2962 585
R4974 gnd.n5544 gnd.n5543 585
R4975 gnd.n5543 gnd.n5542 585
R4976 gnd.n2972 gnd.n2971 585
R4977 gnd.n2983 gnd.n2972 585
R4978 gnd.n5518 gnd.n2996 585
R4979 gnd.n2996 gnd.n2981 585
R4980 gnd.n5520 gnd.n5519 585
R4981 gnd.n5521 gnd.n5520 585
R4982 gnd.n2997 gnd.n2995 585
R4983 gnd.n2995 gnd.n2990 585
R4984 gnd.n5513 gnd.n5512 585
R4985 gnd.n5512 gnd.n5511 585
R4986 gnd.n3000 gnd.n2999 585
R4987 gnd.n3011 gnd.n3000 585
R4988 gnd.n5487 gnd.n3024 585
R4989 gnd.n3024 gnd.n3009 585
R4990 gnd.n5489 gnd.n5488 585
R4991 gnd.n5490 gnd.n5489 585
R4992 gnd.n3025 gnd.n3023 585
R4993 gnd.n3023 gnd.n3019 585
R4994 gnd.n5482 gnd.n5481 585
R4995 gnd.n5481 gnd.n5480 585
R4996 gnd.n3035 gnd.n3027 585
R4997 gnd.n3035 gnd.n2874 585
R4998 gnd.n3034 gnd.n3033 585
R4999 gnd.n3034 gnd.n2872 585
R5000 gnd.n3029 gnd.n3028 585
R5001 gnd.n3028 gnd.n2821 585
R5002 gnd.n2792 gnd.n2791 585
R5003 gnd.n5771 gnd.n2792 585
R5004 gnd.n5774 gnd.n5773 585
R5005 gnd.n5773 gnd.n5772 585
R5006 gnd.n5775 gnd.n2786 585
R5007 gnd.n2786 gnd.n2785 585
R5008 gnd.n5777 gnd.n5776 585
R5009 gnd.n5778 gnd.n5777 585
R5010 gnd.n2787 gnd.n2783 585
R5011 gnd.n5779 gnd.n2783 585
R5012 gnd.n5439 gnd.n3225 585
R5013 gnd.n3225 gnd.n2782 585
R5014 gnd.n5441 gnd.n5440 585
R5015 gnd.n5442 gnd.n5441 585
R5016 gnd.n3226 gnd.n3224 585
R5017 gnd.n3224 gnd.n3223 585
R5018 gnd.n5433 gnd.n5432 585
R5019 gnd.n5432 gnd.n5431 585
R5020 gnd.n3229 gnd.n3228 585
R5021 gnd.n3230 gnd.n3229 585
R5022 gnd.n5420 gnd.n5419 585
R5023 gnd.n5421 gnd.n5420 585
R5024 gnd.n3238 gnd.n3237 585
R5025 gnd.n3244 gnd.n3237 585
R5026 gnd.n5415 gnd.n5414 585
R5027 gnd.n5414 gnd.n5413 585
R5028 gnd.n3241 gnd.n3240 585
R5029 gnd.n3242 gnd.n3241 585
R5030 gnd.n5404 gnd.n5403 585
R5031 gnd.n5405 gnd.n5404 585
R5032 gnd.n3251 gnd.n3250 585
R5033 gnd.n3256 gnd.n3250 585
R5034 gnd.n5399 gnd.n5398 585
R5035 gnd.n5398 gnd.n5397 585
R5036 gnd.n3254 gnd.n3253 585
R5037 gnd.n5135 gnd.n3254 585
R5038 gnd.n5388 gnd.n5387 585
R5039 gnd.n5389 gnd.n5388 585
R5040 gnd.n3264 gnd.n3263 585
R5041 gnd.n5108 gnd.n3263 585
R5042 gnd.n5383 gnd.n5382 585
R5043 gnd.n5382 gnd.n5381 585
R5044 gnd.n3267 gnd.n3266 585
R5045 gnd.n5321 gnd.n3267 585
R5046 gnd.n5372 gnd.n5371 585
R5047 gnd.n5373 gnd.n5372 585
R5048 gnd.n3277 gnd.n3276 585
R5049 gnd.n5096 gnd.n3276 585
R5050 gnd.n5367 gnd.n5366 585
R5051 gnd.n5366 gnd.n5365 585
R5052 gnd.n3280 gnd.n3279 585
R5053 gnd.n5336 gnd.n3280 585
R5054 gnd.n5356 gnd.n5355 585
R5055 gnd.n5357 gnd.n5356 585
R5056 gnd.n3289 gnd.n3288 585
R5057 gnd.n3302 gnd.n3288 585
R5058 gnd.n5351 gnd.n5350 585
R5059 gnd.n5350 gnd.n5349 585
R5060 gnd.n3292 gnd.n3291 585
R5061 gnd.n5082 gnd.n3292 585
R5062 gnd.n5070 gnd.n3318 585
R5063 gnd.n4957 gnd.n3318 585
R5064 gnd.n5072 gnd.n5071 585
R5065 gnd.n5073 gnd.n5072 585
R5066 gnd.n3319 gnd.n3317 585
R5067 gnd.n4945 gnd.n3317 585
R5068 gnd.n5065 gnd.n5064 585
R5069 gnd.n5064 gnd.n5063 585
R5070 gnd.n3322 gnd.n3321 585
R5071 gnd.n4972 gnd.n3322 585
R5072 gnd.n5054 gnd.n5053 585
R5073 gnd.n5055 gnd.n5054 585
R5074 gnd.n3333 gnd.n3332 585
R5075 gnd.n4930 gnd.n3332 585
R5076 gnd.n5049 gnd.n5048 585
R5077 gnd.n5048 gnd.n5047 585
R5078 gnd.n3336 gnd.n3335 585
R5079 gnd.n4987 gnd.n3336 585
R5080 gnd.n5038 gnd.n5037 585
R5081 gnd.n5039 gnd.n5038 585
R5082 gnd.n3348 gnd.n3347 585
R5083 gnd.n4919 gnd.n3347 585
R5084 gnd.n5033 gnd.n5032 585
R5085 gnd.n5032 gnd.n5031 585
R5086 gnd.n3351 gnd.n3350 585
R5087 gnd.n5002 gnd.n3351 585
R5088 gnd.n5022 gnd.n5021 585
R5089 gnd.n5023 gnd.n5022 585
R5090 gnd.n3361 gnd.n3360 585
R5091 gnd.n3374 gnd.n3360 585
R5092 gnd.n5017 gnd.n5016 585
R5093 gnd.n5016 gnd.n5015 585
R5094 gnd.n3364 gnd.n3363 585
R5095 gnd.n4905 gnd.n3364 585
R5096 gnd.n4893 gnd.n3389 585
R5097 gnd.n4778 gnd.n3389 585
R5098 gnd.n4895 gnd.n4894 585
R5099 gnd.n4896 gnd.n4895 585
R5100 gnd.n3390 gnd.n3388 585
R5101 gnd.n4786 gnd.n3388 585
R5102 gnd.n4888 gnd.n4887 585
R5103 gnd.n4887 gnd.n4886 585
R5104 gnd.n3393 gnd.n3392 585
R5105 gnd.n4794 gnd.n3393 585
R5106 gnd.n4877 gnd.n4876 585
R5107 gnd.n4878 gnd.n4877 585
R5108 gnd.n3402 gnd.n3401 585
R5109 gnd.n4751 gnd.n3401 585
R5110 gnd.n4872 gnd.n4871 585
R5111 gnd.n4871 gnd.n4870 585
R5112 gnd.n3405 gnd.n3404 585
R5113 gnd.n4810 gnd.n3405 585
R5114 gnd.n4861 gnd.n4860 585
R5115 gnd.n4862 gnd.n4861 585
R5116 gnd.n3415 gnd.n3414 585
R5117 gnd.n4739 gnd.n3414 585
R5118 gnd.n4856 gnd.n4855 585
R5119 gnd.n4855 gnd.n4854 585
R5120 gnd.n3418 gnd.n3417 585
R5121 gnd.n4825 gnd.n3418 585
R5122 gnd.n4845 gnd.n4844 585
R5123 gnd.n4846 gnd.n4845 585
R5124 gnd.n3427 gnd.n3426 585
R5125 gnd.n3439 gnd.n3426 585
R5126 gnd.n4840 gnd.n4839 585
R5127 gnd.n4839 gnd.n4838 585
R5128 gnd.n3430 gnd.n3429 585
R5129 gnd.n4724 gnd.n3430 585
R5130 gnd.n4712 gnd.n3455 585
R5131 gnd.n4460 gnd.n3455 585
R5132 gnd.n4714 gnd.n4713 585
R5133 gnd.n4715 gnd.n4714 585
R5134 gnd.n3456 gnd.n3454 585
R5135 gnd.n4468 gnd.n3454 585
R5136 gnd.n4707 gnd.n4706 585
R5137 gnd.n4706 gnd.n4705 585
R5138 gnd.n3459 gnd.n3458 585
R5139 gnd.n4442 gnd.n3459 585
R5140 gnd.n4696 gnd.n4695 585
R5141 gnd.n4697 gnd.n4696 585
R5142 gnd.n3469 gnd.n3468 585
R5143 gnd.n4483 gnd.n3468 585
R5144 gnd.n4691 gnd.n4690 585
R5145 gnd.n4690 gnd.n4689 585
R5146 gnd.n3472 gnd.n3471 585
R5147 gnd.n4327 gnd.n3472 585
R5148 gnd.n4680 gnd.n4679 585
R5149 gnd.n4681 gnd.n4680 585
R5150 gnd.n3483 gnd.n3482 585
R5151 gnd.n3488 gnd.n3482 585
R5152 gnd.n4675 gnd.n4674 585
R5153 gnd.n4674 gnd.n4673 585
R5154 gnd.n3486 gnd.n3485 585
R5155 gnd.n3495 gnd.n3486 585
R5156 gnd.n4664 gnd.n4663 585
R5157 gnd.n4665 gnd.n4664 585
R5158 gnd.n3497 gnd.n3496 585
R5159 gnd.n3496 gnd.n3494 585
R5160 gnd.n4659 gnd.n4658 585
R5161 gnd.n4658 gnd.n4657 585
R5162 gnd.n3500 gnd.n3499 585
R5163 gnd.n3508 gnd.n3500 585
R5164 gnd.n4648 gnd.n4647 585
R5165 gnd.n4649 gnd.n4648 585
R5166 gnd.n3510 gnd.n3509 585
R5167 gnd.n3509 gnd.n3507 585
R5168 gnd.n4643 gnd.n4642 585
R5169 gnd.n4642 gnd.n4641 585
R5170 gnd.n3513 gnd.n3512 585
R5171 gnd.n3514 gnd.n3513 585
R5172 gnd.n4632 gnd.n4631 585
R5173 gnd.n4633 gnd.n4632 585
R5174 gnd.n3523 gnd.n3522 585
R5175 gnd.n3522 gnd.n3521 585
R5176 gnd.n4627 gnd.n4626 585
R5177 gnd.n4626 gnd.n4625 585
R5178 gnd.n3526 gnd.n3525 585
R5179 gnd.n4624 gnd.n3526 585
R5180 gnd.n3886 gnd.n3885 585
R5181 gnd.n3885 gnd.n3527 585
R5182 gnd.n3887 gnd.n3880 585
R5183 gnd.n3880 gnd.n3666 585
R5184 gnd.n3889 gnd.n3888 585
R5185 gnd.n3889 gnd.n3564 585
R5186 gnd.n3890 gnd.n3879 585
R5187 gnd.n3890 gnd.n2672 585
R5188 gnd.n3892 gnd.n3891 585
R5189 gnd.n3891 gnd.n2669 585
R5190 gnd.n3893 gnd.n3874 585
R5191 gnd.n3874 gnd.n3732 585
R5192 gnd.n3895 gnd.n3894 585
R5193 gnd.n3895 gnd.n2660 585
R5194 gnd.n3896 gnd.n3873 585
R5195 gnd.n3896 gnd.n2652 585
R5196 gnd.n3898 gnd.n3897 585
R5197 gnd.n3897 gnd.n2649 585
R5198 gnd.n3899 gnd.n3868 585
R5199 gnd.n3868 gnd.n2641 585
R5200 gnd.n3901 gnd.n3900 585
R5201 gnd.n3901 gnd.n2638 585
R5202 gnd.n3902 gnd.n3867 585
R5203 gnd.n3902 gnd.n2630 585
R5204 gnd.n3904 gnd.n3903 585
R5205 gnd.n3903 gnd.n2627 585
R5206 gnd.n3905 gnd.n3862 585
R5207 gnd.n3862 gnd.n2619 585
R5208 gnd.n3907 gnd.n3906 585
R5209 gnd.n3907 gnd.n2616 585
R5210 gnd.n3908 gnd.n3861 585
R5211 gnd.n3908 gnd.n3749 585
R5212 gnd.n3910 gnd.n3909 585
R5213 gnd.n3909 gnd.n2606 585
R5214 gnd.n3911 gnd.n3856 585
R5215 gnd.n3856 gnd.n2598 585
R5216 gnd.n3913 gnd.n3912 585
R5217 gnd.n3913 gnd.n2595 585
R5218 gnd.n3914 gnd.n3855 585
R5219 gnd.n3914 gnd.n2587 585
R5220 gnd.n3916 gnd.n3915 585
R5221 gnd.n3915 gnd.n2584 585
R5222 gnd.n3917 gnd.n3850 585
R5223 gnd.n3850 gnd.n2576 585
R5224 gnd.n3919 gnd.n3918 585
R5225 gnd.n3919 gnd.n2573 585
R5226 gnd.n3920 gnd.n3849 585
R5227 gnd.n3920 gnd.n3762 585
R5228 gnd.n3922 gnd.n3921 585
R5229 gnd.n3921 gnd.n2563 585
R5230 gnd.n3923 gnd.n3847 585
R5231 gnd.n3847 gnd.n2556 585
R5232 gnd.n3925 gnd.n3924 585
R5233 gnd.n3925 gnd.n2553 585
R5234 gnd.n3927 gnd.n3926 585
R5235 gnd.n3926 gnd.n2545 585
R5236 gnd.n3929 gnd.n3928 585
R5237 gnd.n3929 gnd.n2542 585
R5238 gnd.n3931 gnd.n3930 585
R5239 gnd.n3931 gnd.n2537 585
R5240 gnd.n3932 gnd.n3845 585
R5241 gnd.n3932 gnd.n2534 585
R5242 gnd.n3934 gnd.n3933 585
R5243 gnd.n3933 gnd.n3775 585
R5244 gnd.n3846 gnd.n3841 585
R5245 gnd.n3846 gnd.n2524 585
R5246 gnd.n3938 gnd.n3839 585
R5247 gnd.n3839 gnd.n2518 585
R5248 gnd.n3940 gnd.n3939 585
R5249 gnd.n3940 gnd.n2515 585
R5250 gnd.n3941 gnd.n3838 585
R5251 gnd.n3941 gnd.n2507 585
R5252 gnd.n3943 gnd.n3942 585
R5253 gnd.n3942 gnd.n2504 585
R5254 gnd.n3944 gnd.n3833 585
R5255 gnd.n3833 gnd.n2496 585
R5256 gnd.n3946 gnd.n3945 585
R5257 gnd.n3946 gnd.n2493 585
R5258 gnd.n3947 gnd.n3832 585
R5259 gnd.n3947 gnd.n3788 585
R5260 gnd.n3949 gnd.n3948 585
R5261 gnd.n3948 gnd.n2483 585
R5262 gnd.n3950 gnd.n3827 585
R5263 gnd.n3827 gnd.n2475 585
R5264 gnd.n3952 gnd.n3951 585
R5265 gnd.n3952 gnd.n2472 585
R5266 gnd.n3953 gnd.n3826 585
R5267 gnd.n3953 gnd.n2464 585
R5268 gnd.n3955 gnd.n3954 585
R5269 gnd.n3954 gnd.n2461 585
R5270 gnd.n3956 gnd.n3821 585
R5271 gnd.n3821 gnd.n2453 585
R5272 gnd.n3958 gnd.n3957 585
R5273 gnd.n3958 gnd.n2450 585
R5274 gnd.n3959 gnd.n3820 585
R5275 gnd.n3959 gnd.n3801 585
R5276 gnd.n3961 gnd.n3960 585
R5277 gnd.n3960 gnd.n2440 585
R5278 gnd.n3962 gnd.n3815 585
R5279 gnd.n3815 gnd.n2432 585
R5280 gnd.n3964 gnd.n3963 585
R5281 gnd.n3964 gnd.n2429 585
R5282 gnd.n3965 gnd.n3814 585
R5283 gnd.n3965 gnd.n2420 585
R5284 gnd.n3967 gnd.n3966 585
R5285 gnd.n3966 gnd.n2417 585
R5286 gnd.n3968 gnd.n3811 585
R5287 gnd.n3811 gnd.n2407 585
R5288 gnd.n5781 gnd.n5780 585
R5289 gnd.n5780 gnd.n5779 585
R5290 gnd.n5782 gnd.n2779 585
R5291 gnd.n2782 gnd.n2779 585
R5292 gnd.n5783 gnd.n2778 585
R5293 gnd.n5442 gnd.n2778 585
R5294 gnd.n3222 gnd.n2776 585
R5295 gnd.n3223 gnd.n3222 585
R5296 gnd.n5787 gnd.n2775 585
R5297 gnd.n5431 gnd.n2775 585
R5298 gnd.n5788 gnd.n2774 585
R5299 gnd.n3230 gnd.n2774 585
R5300 gnd.n5789 gnd.n2773 585
R5301 gnd.n5421 gnd.n2773 585
R5302 gnd.n3243 gnd.n2771 585
R5303 gnd.n3244 gnd.n3243 585
R5304 gnd.n5793 gnd.n2770 585
R5305 gnd.n5413 gnd.n2770 585
R5306 gnd.n5794 gnd.n2769 585
R5307 gnd.n3242 gnd.n2769 585
R5308 gnd.n5795 gnd.n2768 585
R5309 gnd.n5405 gnd.n2768 585
R5310 gnd.n3255 gnd.n2766 585
R5311 gnd.n3256 gnd.n3255 585
R5312 gnd.n5799 gnd.n2765 585
R5313 gnd.n5397 gnd.n2765 585
R5314 gnd.n5800 gnd.n2764 585
R5315 gnd.n5135 gnd.n2764 585
R5316 gnd.n5801 gnd.n2763 585
R5317 gnd.n5389 gnd.n2763 585
R5318 gnd.n5107 gnd.n2761 585
R5319 gnd.n5108 gnd.n5107 585
R5320 gnd.n5805 gnd.n2760 585
R5321 gnd.n5381 gnd.n2760 585
R5322 gnd.n5806 gnd.n2759 585
R5323 gnd.n5321 gnd.n2759 585
R5324 gnd.n5807 gnd.n2758 585
R5325 gnd.n5373 gnd.n2758 585
R5326 gnd.n5095 gnd.n2756 585
R5327 gnd.n5096 gnd.n5095 585
R5328 gnd.n5811 gnd.n2755 585
R5329 gnd.n5365 gnd.n2755 585
R5330 gnd.n5812 gnd.n2754 585
R5331 gnd.n5336 gnd.n2754 585
R5332 gnd.n5813 gnd.n2753 585
R5333 gnd.n5357 gnd.n2753 585
R5334 gnd.n3301 gnd.n2751 585
R5335 gnd.n3302 gnd.n3301 585
R5336 gnd.n5817 gnd.n2750 585
R5337 gnd.n5349 gnd.n2750 585
R5338 gnd.n5818 gnd.n2749 585
R5339 gnd.n5082 gnd.n2749 585
R5340 gnd.n5819 gnd.n2748 585
R5341 gnd.n4957 gnd.n2748 585
R5342 gnd.n3315 gnd.n2746 585
R5343 gnd.n5073 gnd.n3315 585
R5344 gnd.n5823 gnd.n2745 585
R5345 gnd.n4945 gnd.n2745 585
R5346 gnd.n5824 gnd.n2744 585
R5347 gnd.n5063 gnd.n2744 585
R5348 gnd.n5825 gnd.n2743 585
R5349 gnd.n4972 gnd.n2743 585
R5350 gnd.n3330 gnd.n2741 585
R5351 gnd.n5055 gnd.n3330 585
R5352 gnd.n5829 gnd.n2740 585
R5353 gnd.n4930 gnd.n2740 585
R5354 gnd.n5830 gnd.n2739 585
R5355 gnd.n5047 gnd.n2739 585
R5356 gnd.n5831 gnd.n2738 585
R5357 gnd.n4987 gnd.n2738 585
R5358 gnd.n3345 gnd.n2736 585
R5359 gnd.n5039 gnd.n3345 585
R5360 gnd.n5835 gnd.n2735 585
R5361 gnd.n4919 gnd.n2735 585
R5362 gnd.n5836 gnd.n2734 585
R5363 gnd.n5031 gnd.n2734 585
R5364 gnd.n5837 gnd.n2733 585
R5365 gnd.n5002 gnd.n2733 585
R5366 gnd.n3358 gnd.n2731 585
R5367 gnd.n5023 gnd.n3358 585
R5368 gnd.n5841 gnd.n2730 585
R5369 gnd.n3374 gnd.n2730 585
R5370 gnd.n5842 gnd.n2729 585
R5371 gnd.n5015 gnd.n2729 585
R5372 gnd.n5843 gnd.n2728 585
R5373 gnd.n4905 gnd.n2728 585
R5374 gnd.n4777 gnd.n2726 585
R5375 gnd.n4778 gnd.n4777 585
R5376 gnd.n5847 gnd.n2725 585
R5377 gnd.n4896 gnd.n2725 585
R5378 gnd.n5848 gnd.n2724 585
R5379 gnd.n4786 gnd.n2724 585
R5380 gnd.n5849 gnd.n2723 585
R5381 gnd.n4886 gnd.n2723 585
R5382 gnd.n4760 gnd.n2721 585
R5383 gnd.n4794 gnd.n4760 585
R5384 gnd.n5853 gnd.n2720 585
R5385 gnd.n4878 gnd.n2720 585
R5386 gnd.n5854 gnd.n2719 585
R5387 gnd.n4751 gnd.n2719 585
R5388 gnd.n5855 gnd.n2718 585
R5389 gnd.n4870 gnd.n2718 585
R5390 gnd.n4809 gnd.n2716 585
R5391 gnd.n4810 gnd.n4809 585
R5392 gnd.n5859 gnd.n2715 585
R5393 gnd.n4862 gnd.n2715 585
R5394 gnd.n5860 gnd.n2714 585
R5395 gnd.n4739 gnd.n2714 585
R5396 gnd.n5861 gnd.n2713 585
R5397 gnd.n4854 gnd.n2713 585
R5398 gnd.n4734 gnd.n2711 585
R5399 gnd.n4825 gnd.n4734 585
R5400 gnd.n5865 gnd.n2710 585
R5401 gnd.n4846 gnd.n2710 585
R5402 gnd.n5866 gnd.n2709 585
R5403 gnd.n3439 gnd.n2709 585
R5404 gnd.n5867 gnd.n2708 585
R5405 gnd.n4838 gnd.n2708 585
R5406 gnd.n3446 gnd.n2706 585
R5407 gnd.n4724 gnd.n3446 585
R5408 gnd.n5871 gnd.n2705 585
R5409 gnd.n4460 gnd.n2705 585
R5410 gnd.n5872 gnd.n2704 585
R5411 gnd.n4715 gnd.n2704 585
R5412 gnd.n5873 gnd.n2703 585
R5413 gnd.n4468 gnd.n2703 585
R5414 gnd.n3460 gnd.n2701 585
R5415 gnd.n4705 gnd.n3460 585
R5416 gnd.n5877 gnd.n2700 585
R5417 gnd.n4442 gnd.n2700 585
R5418 gnd.n5878 gnd.n2699 585
R5419 gnd.n4697 gnd.n2699 585
R5420 gnd.n5879 gnd.n2698 585
R5421 gnd.n4483 gnd.n2698 585
R5422 gnd.n3474 gnd.n2696 585
R5423 gnd.n4689 gnd.n3474 585
R5424 gnd.n5883 gnd.n2695 585
R5425 gnd.n4327 gnd.n2695 585
R5426 gnd.n5884 gnd.n2694 585
R5427 gnd.n4681 gnd.n2694 585
R5428 gnd.n5885 gnd.n2693 585
R5429 gnd.n3488 gnd.n2693 585
R5430 gnd.n3487 gnd.n2691 585
R5431 gnd.n4673 gnd.n3487 585
R5432 gnd.n5889 gnd.n2690 585
R5433 gnd.n3495 gnd.n2690 585
R5434 gnd.n5890 gnd.n2689 585
R5435 gnd.n4665 gnd.n2689 585
R5436 gnd.n5891 gnd.n2688 585
R5437 gnd.n3494 gnd.n2688 585
R5438 gnd.n3501 gnd.n2686 585
R5439 gnd.n4657 gnd.n3501 585
R5440 gnd.n5895 gnd.n2685 585
R5441 gnd.n3508 gnd.n2685 585
R5442 gnd.n5896 gnd.n2684 585
R5443 gnd.n4649 gnd.n2684 585
R5444 gnd.n5897 gnd.n2683 585
R5445 gnd.n3507 gnd.n2683 585
R5446 gnd.n3515 gnd.n2681 585
R5447 gnd.n4641 gnd.n3515 585
R5448 gnd.n5901 gnd.n2680 585
R5449 gnd.n3514 gnd.n2680 585
R5450 gnd.n5902 gnd.n2679 585
R5451 gnd.n4633 gnd.n2679 585
R5452 gnd.n5903 gnd.n2678 585
R5453 gnd.n3521 gnd.n2678 585
R5454 gnd.n3600 gnd.n3599 585
R5455 gnd.n3610 gnd.n3609 585
R5456 gnd.n3612 gnd.n3611 585
R5457 gnd.n3594 gnd.n3593 585
R5458 gnd.n3621 gnd.n3595 585
R5459 gnd.n3624 gnd.n3623 585
R5460 gnd.n3622 gnd.n3587 585
R5461 gnd.n3634 gnd.n3633 585
R5462 gnd.n3636 gnd.n3635 585
R5463 gnd.n3582 gnd.n3581 585
R5464 gnd.n3645 gnd.n3583 585
R5465 gnd.n3648 gnd.n3647 585
R5466 gnd.n3646 gnd.n3575 585
R5467 gnd.n3657 gnd.n3656 585
R5468 gnd.n3659 gnd.n3658 585
R5469 gnd.n3557 gnd.n3556 585
R5470 gnd.n4596 gnd.n3558 585
R5471 gnd.n4598 gnd.n4597 585
R5472 gnd.n4600 gnd.n4599 585
R5473 gnd.n3552 gnd.n3551 585
R5474 gnd.n4605 gnd.n3553 585
R5475 gnd.n4607 gnd.n4606 585
R5476 gnd.n4609 gnd.n4608 585
R5477 gnd.n3548 gnd.n3547 585
R5478 gnd.n4613 gnd.n3549 585
R5479 gnd.n4616 gnd.n4615 585
R5480 gnd.n4618 gnd.n4617 585
R5481 gnd.n3543 gnd.n3542 585
R5482 gnd.n4623 gnd.n4622 585
R5483 gnd.n4624 gnd.n4623 585
R5484 gnd.n5446 gnd.n2784 585
R5485 gnd.n5779 gnd.n2784 585
R5486 gnd.n5445 gnd.n5444 585
R5487 gnd.n5444 gnd.n2782 585
R5488 gnd.n5443 gnd.n3220 585
R5489 gnd.n5443 gnd.n5442 585
R5490 gnd.n3233 gnd.n3221 585
R5491 gnd.n3223 gnd.n3221 585
R5492 gnd.n5430 gnd.n5429 585
R5493 gnd.n5431 gnd.n5430 585
R5494 gnd.n3232 gnd.n3231 585
R5495 gnd.n3231 gnd.n3230 585
R5496 gnd.n5423 gnd.n5422 585
R5497 gnd.n5422 gnd.n5421 585
R5498 gnd.n3236 gnd.n3235 585
R5499 gnd.n3244 gnd.n3236 585
R5500 gnd.n5412 gnd.n5411 585
R5501 gnd.n5413 gnd.n5412 585
R5502 gnd.n3246 gnd.n3245 585
R5503 gnd.n3245 gnd.n3242 585
R5504 gnd.n5407 gnd.n5406 585
R5505 gnd.n5406 gnd.n5405 585
R5506 gnd.n3249 gnd.n3248 585
R5507 gnd.n3256 gnd.n3249 585
R5508 gnd.n5396 gnd.n5395 585
R5509 gnd.n5397 gnd.n5396 585
R5510 gnd.n3258 gnd.n3257 585
R5511 gnd.n5135 gnd.n3257 585
R5512 gnd.n5391 gnd.n5390 585
R5513 gnd.n5390 gnd.n5389 585
R5514 gnd.n3261 gnd.n3260 585
R5515 gnd.n5108 gnd.n3261 585
R5516 gnd.n5380 gnd.n5379 585
R5517 gnd.n5381 gnd.n5380 585
R5518 gnd.n3270 gnd.n3269 585
R5519 gnd.n5321 gnd.n3269 585
R5520 gnd.n5375 gnd.n5374 585
R5521 gnd.n5374 gnd.n5373 585
R5522 gnd.n3273 gnd.n3272 585
R5523 gnd.n5096 gnd.n3273 585
R5524 gnd.n5364 gnd.n5363 585
R5525 gnd.n5365 gnd.n5364 585
R5526 gnd.n3283 gnd.n3282 585
R5527 gnd.n5336 gnd.n3282 585
R5528 gnd.n5359 gnd.n5358 585
R5529 gnd.n5358 gnd.n5357 585
R5530 gnd.n3286 gnd.n3285 585
R5531 gnd.n3302 gnd.n3286 585
R5532 gnd.n3310 gnd.n3295 585
R5533 gnd.n5349 gnd.n3295 585
R5534 gnd.n5081 gnd.n5080 585
R5535 gnd.n5082 gnd.n5081 585
R5536 gnd.n3309 gnd.n3308 585
R5537 gnd.n4957 gnd.n3308 585
R5538 gnd.n5075 gnd.n5074 585
R5539 gnd.n5074 gnd.n5073 585
R5540 gnd.n3313 gnd.n3312 585
R5541 gnd.n4945 gnd.n3313 585
R5542 gnd.n5062 gnd.n5061 585
R5543 gnd.n5063 gnd.n5062 585
R5544 gnd.n3325 gnd.n3324 585
R5545 gnd.n4972 gnd.n3324 585
R5546 gnd.n5057 gnd.n5056 585
R5547 gnd.n5056 gnd.n5055 585
R5548 gnd.n3328 gnd.n3327 585
R5549 gnd.n4930 gnd.n3328 585
R5550 gnd.n5046 gnd.n5045 585
R5551 gnd.n5047 gnd.n5046 585
R5552 gnd.n3340 gnd.n3339 585
R5553 gnd.n4987 gnd.n3339 585
R5554 gnd.n5041 gnd.n5040 585
R5555 gnd.n5040 gnd.n5039 585
R5556 gnd.n3343 gnd.n3342 585
R5557 gnd.n4919 gnd.n3343 585
R5558 gnd.n5030 gnd.n5029 585
R5559 gnd.n5031 gnd.n5030 585
R5560 gnd.n3354 gnd.n3353 585
R5561 gnd.n5002 gnd.n3353 585
R5562 gnd.n5025 gnd.n5024 585
R5563 gnd.n5024 gnd.n5023 585
R5564 gnd.n3357 gnd.n3356 585
R5565 gnd.n3374 gnd.n3357 585
R5566 gnd.n3382 gnd.n3368 585
R5567 gnd.n5015 gnd.n3368 585
R5568 gnd.n4904 gnd.n4903 585
R5569 gnd.n4905 gnd.n4904 585
R5570 gnd.n3381 gnd.n3380 585
R5571 gnd.n4778 gnd.n3380 585
R5572 gnd.n4898 gnd.n4897 585
R5573 gnd.n4897 gnd.n4896 585
R5574 gnd.n3385 gnd.n3384 585
R5575 gnd.n4786 gnd.n3385 585
R5576 gnd.n4885 gnd.n4884 585
R5577 gnd.n4886 gnd.n4885 585
R5578 gnd.n3396 gnd.n3395 585
R5579 gnd.n4794 gnd.n3395 585
R5580 gnd.n4880 gnd.n4879 585
R5581 gnd.n4879 gnd.n4878 585
R5582 gnd.n3399 gnd.n3398 585
R5583 gnd.n4751 gnd.n3399 585
R5584 gnd.n4869 gnd.n4868 585
R5585 gnd.n4870 gnd.n4869 585
R5586 gnd.n3409 gnd.n3408 585
R5587 gnd.n4810 gnd.n3408 585
R5588 gnd.n4864 gnd.n4863 585
R5589 gnd.n4863 gnd.n4862 585
R5590 gnd.n3412 gnd.n3411 585
R5591 gnd.n4739 gnd.n3412 585
R5592 gnd.n4853 gnd.n4852 585
R5593 gnd.n4854 gnd.n4853 585
R5594 gnd.n3421 gnd.n3420 585
R5595 gnd.n4825 gnd.n3420 585
R5596 gnd.n4848 gnd.n4847 585
R5597 gnd.n4847 gnd.n4846 585
R5598 gnd.n3424 gnd.n3423 585
R5599 gnd.n3439 gnd.n3424 585
R5600 gnd.n3449 gnd.n3433 585
R5601 gnd.n4838 gnd.n3433 585
R5602 gnd.n4723 gnd.n4722 585
R5603 gnd.n4724 gnd.n4723 585
R5604 gnd.n3448 gnd.n3447 585
R5605 gnd.n4460 gnd.n3447 585
R5606 gnd.n4717 gnd.n4716 585
R5607 gnd.n4716 gnd.n4715 585
R5608 gnd.n3452 gnd.n3451 585
R5609 gnd.n4468 gnd.n3452 585
R5610 gnd.n4704 gnd.n4703 585
R5611 gnd.n4705 gnd.n4704 585
R5612 gnd.n3463 gnd.n3462 585
R5613 gnd.n4442 gnd.n3462 585
R5614 gnd.n4699 gnd.n4698 585
R5615 gnd.n4698 gnd.n4697 585
R5616 gnd.n3466 gnd.n3465 585
R5617 gnd.n4483 gnd.n3466 585
R5618 gnd.n4688 gnd.n4687 585
R5619 gnd.n4689 gnd.n4688 585
R5620 gnd.n3477 gnd.n3476 585
R5621 gnd.n4327 gnd.n3476 585
R5622 gnd.n4683 gnd.n4682 585
R5623 gnd.n4682 gnd.n4681 585
R5624 gnd.n3480 gnd.n3479 585
R5625 gnd.n3488 gnd.n3480 585
R5626 gnd.n4672 gnd.n4671 585
R5627 gnd.n4673 gnd.n4672 585
R5628 gnd.n3490 gnd.n3489 585
R5629 gnd.n3495 gnd.n3489 585
R5630 gnd.n4667 gnd.n4666 585
R5631 gnd.n4666 gnd.n4665 585
R5632 gnd.n3493 gnd.n3492 585
R5633 gnd.n3494 gnd.n3493 585
R5634 gnd.n4656 gnd.n4655 585
R5635 gnd.n4657 gnd.n4656 585
R5636 gnd.n3503 gnd.n3502 585
R5637 gnd.n3508 gnd.n3502 585
R5638 gnd.n4651 gnd.n4650 585
R5639 gnd.n4650 gnd.n4649 585
R5640 gnd.n3506 gnd.n3505 585
R5641 gnd.n3507 gnd.n3506 585
R5642 gnd.n4640 gnd.n4639 585
R5643 gnd.n4641 gnd.n4640 585
R5644 gnd.n3517 gnd.n3516 585
R5645 gnd.n3516 gnd.n3514 585
R5646 gnd.n4635 gnd.n4634 585
R5647 gnd.n4634 gnd.n4633 585
R5648 gnd.n3520 gnd.n3519 585
R5649 gnd.n3521 gnd.n3520 585
R5650 gnd.n5453 gnd.n5452 585
R5651 gnd.n5452 gnd.n2785 585
R5652 gnd.n5454 gnd.n5451 585
R5653 gnd.n5449 gnd.n3218 585
R5654 gnd.n5458 gnd.n3217 585
R5655 gnd.n5462 gnd.n3215 585
R5656 gnd.n5463 gnd.n3214 585
R5657 gnd.n3212 gnd.n3210 585
R5658 gnd.n5467 gnd.n3209 585
R5659 gnd.n5468 gnd.n3207 585
R5660 gnd.n5469 gnd.n3206 585
R5661 gnd.n3204 gnd.n3084 585
R5662 gnd.n3203 gnd.n3085 585
R5663 gnd.n3201 gnd.n3200 585
R5664 gnd.n3087 gnd.n3086 585
R5665 gnd.n3191 gnd.n3190 585
R5666 gnd.n3188 gnd.n3097 585
R5667 gnd.n3186 gnd.n3185 585
R5668 gnd.n3099 gnd.n3098 585
R5669 gnd.n3174 gnd.n3173 585
R5670 gnd.n3171 gnd.n3106 585
R5671 gnd.n3169 gnd.n3168 585
R5672 gnd.n3108 gnd.n3107 585
R5673 gnd.n3157 gnd.n3156 585
R5674 gnd.n3154 gnd.n3115 585
R5675 gnd.n3152 gnd.n3151 585
R5676 gnd.n3117 gnd.n3116 585
R5677 gnd.n3140 gnd.n3139 585
R5678 gnd.n3137 gnd.n3135 585
R5679 gnd.n3124 gnd.n2781 585
R5680 gnd.n4309 gnd.t176 543.808
R5681 gnd.n5165 gnd.t173 543.808
R5682 gnd.n4364 gnd.t125 543.808
R5683 gnd.n5159 gnd.t118 543.808
R5684 gnd.n6423 gnd.n6422 491.447
R5685 gnd.n5309 gnd.n5308 458.866
R5686 gnd.n5192 gnd.n5191 458.866
R5687 gnd.n4494 gnd.n4492 458.866
R5688 gnd.n4490 gnd.n4328 458.866
R5689 gnd.n3545 gnd.t145 371.625
R5690 gnd.n7312 gnd.t78 371.625
R5691 gnd.n3091 gnd.t103 371.625
R5692 gnd.n3560 gnd.t139 371.625
R5693 gnd.n2844 gnd.t100 371.625
R5694 gnd.n2866 gnd.t85 371.625
R5695 gnd.n175 gnd.t179 371.625
R5696 gnd.n7405 gnd.t89 371.625
R5697 gnd.n2373 gnd.t165 371.625
R5698 gnd.n2395 gnd.t156 371.625
R5699 gnd.n3728 gnd.t96 371.625
R5700 gnd.n3706 gnd.t132 371.625
R5701 gnd.n3994 gnd.t110 371.625
R5702 gnd.n5459 gnd.t114 371.625
R5703 gnd.n1483 gnd.t92 323.425
R5704 gnd.n1051 gnd.t135 323.425
R5705 gnd.n2291 gnd.n2265 289.615
R5706 gnd.n2259 gnd.n2233 289.615
R5707 gnd.n2227 gnd.n2201 289.615
R5708 gnd.n2196 gnd.n2170 289.615
R5709 gnd.n2164 gnd.n2138 289.615
R5710 gnd.n2132 gnd.n2106 289.615
R5711 gnd.n2100 gnd.n2074 289.615
R5712 gnd.n2069 gnd.n2043 289.615
R5713 gnd.n1557 gnd.t106 279.217
R5714 gnd.n1072 gnd.t149 279.217
R5715 gnd.n7115 gnd.n102 275.24
R5716 gnd.n4336 gnd.t84 260.649
R5717 gnd.n5125 gnd.t124 260.649
R5718 gnd.n4427 gnd.n3481 256.663
R5719 gnd.n4351 gnd.n3481 256.663
R5720 gnd.n4420 gnd.n3481 256.663
R5721 gnd.n4414 gnd.n3481 256.663
R5722 gnd.n4412 gnd.n3481 256.663
R5723 gnd.n4406 gnd.n3481 256.663
R5724 gnd.n4404 gnd.n3481 256.663
R5725 gnd.n4398 gnd.n3481 256.663
R5726 gnd.n4396 gnd.n3481 256.663
R5727 gnd.n4390 gnd.n3481 256.663
R5728 gnd.n4388 gnd.n3481 256.663
R5729 gnd.n4382 gnd.n3481 256.663
R5730 gnd.n4380 gnd.n3481 256.663
R5731 gnd.n4374 gnd.n3481 256.663
R5732 gnd.n4367 gnd.n3481 256.663
R5733 gnd.n4368 gnd.n3481 256.663
R5734 gnd.n4560 gnd.n4307 256.663
R5735 gnd.n4558 gnd.n3481 256.663
R5736 gnd.n4556 gnd.n3481 256.663
R5737 gnd.n4549 gnd.n3481 256.663
R5738 gnd.n4547 gnd.n3481 256.663
R5739 gnd.n4541 gnd.n3481 256.663
R5740 gnd.n4539 gnd.n3481 256.663
R5741 gnd.n4533 gnd.n3481 256.663
R5742 gnd.n4531 gnd.n3481 256.663
R5743 gnd.n4525 gnd.n3481 256.663
R5744 gnd.n4523 gnd.n3481 256.663
R5745 gnd.n4517 gnd.n3481 256.663
R5746 gnd.n4515 gnd.n3481 256.663
R5747 gnd.n4509 gnd.n3481 256.663
R5748 gnd.n4507 gnd.n3481 256.663
R5749 gnd.n4501 gnd.n3481 256.663
R5750 gnd.n4499 gnd.n3481 256.663
R5751 gnd.n4493 gnd.n3481 256.663
R5752 gnd.n5190 gnd.n5136 256.663
R5753 gnd.n5197 gnd.n5136 256.663
R5754 gnd.n5186 gnd.n5136 256.663
R5755 gnd.n5204 gnd.n5136 256.663
R5756 gnd.n5183 gnd.n5136 256.663
R5757 gnd.n5211 gnd.n5136 256.663
R5758 gnd.n5180 gnd.n5136 256.663
R5759 gnd.n5218 gnd.n5136 256.663
R5760 gnd.n5177 gnd.n5136 256.663
R5761 gnd.n5225 gnd.n5136 256.663
R5762 gnd.n5174 gnd.n5136 256.663
R5763 gnd.n5232 gnd.n5136 256.663
R5764 gnd.n5171 gnd.n5136 256.663
R5765 gnd.n5239 gnd.n5136 256.663
R5766 gnd.n5168 gnd.n5136 256.663
R5767 gnd.n5247 gnd.n5136 256.663
R5768 gnd.n5250 gnd.n2841 256.663
R5769 gnd.n5251 gnd.n5136 256.663
R5770 gnd.n5162 gnd.n5136 256.663
R5771 gnd.n5258 gnd.n5136 256.663
R5772 gnd.n5157 gnd.n5136 256.663
R5773 gnd.n5265 gnd.n5136 256.663
R5774 gnd.n5154 gnd.n5136 256.663
R5775 gnd.n5272 gnd.n5136 256.663
R5776 gnd.n5151 gnd.n5136 256.663
R5777 gnd.n5279 gnd.n5136 256.663
R5778 gnd.n5148 gnd.n5136 256.663
R5779 gnd.n5286 gnd.n5136 256.663
R5780 gnd.n5145 gnd.n5136 256.663
R5781 gnd.n5293 gnd.n5136 256.663
R5782 gnd.n5142 gnd.n5136 256.663
R5783 gnd.n5300 gnd.n5136 256.663
R5784 gnd.n5139 gnd.n5136 256.663
R5785 gnd.n5307 gnd.n5136 256.663
R5786 gnd.n6148 gnd.n2341 242.672
R5787 gnd.n6148 gnd.n2342 242.672
R5788 gnd.n6148 gnd.n2343 242.672
R5789 gnd.n6148 gnd.n2344 242.672
R5790 gnd.n6148 gnd.n2345 242.672
R5791 gnd.n6148 gnd.n2346 242.672
R5792 gnd.n6148 gnd.n2347 242.672
R5793 gnd.n6148 gnd.n2348 242.672
R5794 gnd.n6148 gnd.n2349 242.672
R5795 gnd.n4591 gnd.n4590 242.672
R5796 gnd.n4590 gnd.n3665 242.672
R5797 gnd.n4590 gnd.n3571 242.672
R5798 gnd.n4590 gnd.n3570 242.672
R5799 gnd.n4590 gnd.n3569 242.672
R5800 gnd.n4590 gnd.n3568 242.672
R5801 gnd.n4590 gnd.n3567 242.672
R5802 gnd.n4590 gnd.n3566 242.672
R5803 gnd.n4590 gnd.n3565 242.672
R5804 gnd.n5770 gnd.n2811 242.672
R5805 gnd.n5770 gnd.n2812 242.672
R5806 gnd.n5770 gnd.n2813 242.672
R5807 gnd.n5770 gnd.n2814 242.672
R5808 gnd.n5770 gnd.n2815 242.672
R5809 gnd.n5770 gnd.n2816 242.672
R5810 gnd.n5770 gnd.n2817 242.672
R5811 gnd.n5770 gnd.n2818 242.672
R5812 gnd.n5770 gnd.n2819 242.672
R5813 gnd.n7314 gnd.n102 242.672
R5814 gnd.n7310 gnd.n102 242.672
R5815 gnd.n7305 gnd.n102 242.672
R5816 gnd.n7302 gnd.n102 242.672
R5817 gnd.n7297 gnd.n102 242.672
R5818 gnd.n7294 gnd.n102 242.672
R5819 gnd.n7289 gnd.n102 242.672
R5820 gnd.n7286 gnd.n102 242.672
R5821 gnd.n7281 gnd.n102 242.672
R5822 gnd.n1611 gnd.n1610 242.672
R5823 gnd.n1611 gnd.n1521 242.672
R5824 gnd.n1611 gnd.n1522 242.672
R5825 gnd.n1611 gnd.n1523 242.672
R5826 gnd.n1611 gnd.n1524 242.672
R5827 gnd.n1611 gnd.n1525 242.672
R5828 gnd.n1611 gnd.n1526 242.672
R5829 gnd.n1611 gnd.n1527 242.672
R5830 gnd.n1611 gnd.n1528 242.672
R5831 gnd.n1611 gnd.n1529 242.672
R5832 gnd.n1611 gnd.n1530 242.672
R5833 gnd.n1611 gnd.n1531 242.672
R5834 gnd.n1612 gnd.n1611 242.672
R5835 gnd.n6195 gnd.n2322 242.672
R5836 gnd.n6195 gnd.n1068 242.672
R5837 gnd.n6195 gnd.n1067 242.672
R5838 gnd.n6195 gnd.n1066 242.672
R5839 gnd.n6195 gnd.n1065 242.672
R5840 gnd.n6195 gnd.n1064 242.672
R5841 gnd.n6195 gnd.n1063 242.672
R5842 gnd.n6195 gnd.n1062 242.672
R5843 gnd.n6195 gnd.n1061 242.672
R5844 gnd.n6195 gnd.n1060 242.672
R5845 gnd.n6195 gnd.n1059 242.672
R5846 gnd.n6195 gnd.n1058 242.672
R5847 gnd.n6195 gnd.n1057 242.672
R5848 gnd.n1695 gnd.n1694 242.672
R5849 gnd.n1694 gnd.n1433 242.672
R5850 gnd.n1694 gnd.n1434 242.672
R5851 gnd.n1694 gnd.n1435 242.672
R5852 gnd.n1694 gnd.n1436 242.672
R5853 gnd.n1694 gnd.n1437 242.672
R5854 gnd.n1694 gnd.n1438 242.672
R5855 gnd.n1694 gnd.n1439 242.672
R5856 gnd.n6195 gnd.n1050 242.672
R5857 gnd.n6196 gnd.n6195 242.672
R5858 gnd.n6195 gnd.n6149 242.672
R5859 gnd.n6195 gnd.n6150 242.672
R5860 gnd.n6195 gnd.n6151 242.672
R5861 gnd.n6195 gnd.n6152 242.672
R5862 gnd.n6195 gnd.n6153 242.672
R5863 gnd.n6195 gnd.n6154 242.672
R5864 gnd.n6148 gnd.n6147 242.672
R5865 gnd.n6148 gnd.n2323 242.672
R5866 gnd.n6148 gnd.n2324 242.672
R5867 gnd.n6148 gnd.n2325 242.672
R5868 gnd.n6148 gnd.n2326 242.672
R5869 gnd.n6148 gnd.n2327 242.672
R5870 gnd.n6148 gnd.n2328 242.672
R5871 gnd.n6148 gnd.n2329 242.672
R5872 gnd.n6148 gnd.n2330 242.672
R5873 gnd.n6148 gnd.n2331 242.672
R5874 gnd.n6148 gnd.n2332 242.672
R5875 gnd.n6148 gnd.n2333 242.672
R5876 gnd.n6148 gnd.n2334 242.672
R5877 gnd.n6148 gnd.n2335 242.672
R5878 gnd.n6148 gnd.n2336 242.672
R5879 gnd.n6148 gnd.n2337 242.672
R5880 gnd.n6148 gnd.n2338 242.672
R5881 gnd.n6148 gnd.n2339 242.672
R5882 gnd.n6148 gnd.n2340 242.672
R5883 gnd.n4590 gnd.n3667 242.672
R5884 gnd.n4590 gnd.n3668 242.672
R5885 gnd.n4590 gnd.n3669 242.672
R5886 gnd.n4590 gnd.n3670 242.672
R5887 gnd.n4590 gnd.n3671 242.672
R5888 gnd.n4590 gnd.n3672 242.672
R5889 gnd.n4590 gnd.n3673 242.672
R5890 gnd.n4590 gnd.n3674 242.672
R5891 gnd.n4590 gnd.n3675 242.672
R5892 gnd.n4590 gnd.n3676 242.672
R5893 gnd.n4590 gnd.n3677 242.672
R5894 gnd.n4561 gnd.n3708 242.672
R5895 gnd.n4590 gnd.n3678 242.672
R5896 gnd.n4590 gnd.n3679 242.672
R5897 gnd.n4590 gnd.n3680 242.672
R5898 gnd.n4590 gnd.n3681 242.672
R5899 gnd.n4590 gnd.n3682 242.672
R5900 gnd.n4590 gnd.n3683 242.672
R5901 gnd.n4590 gnd.n3684 242.672
R5902 gnd.n4590 gnd.n4589 242.672
R5903 gnd.n5770 gnd.n5769 242.672
R5904 gnd.n5770 gnd.n2793 242.672
R5905 gnd.n5770 gnd.n2794 242.672
R5906 gnd.n5770 gnd.n2795 242.672
R5907 gnd.n5770 gnd.n2796 242.672
R5908 gnd.n5770 gnd.n2797 242.672
R5909 gnd.n5770 gnd.n2798 242.672
R5910 gnd.n5770 gnd.n2799 242.672
R5911 gnd.n5738 gnd.n2842 242.672
R5912 gnd.n5770 gnd.n2800 242.672
R5913 gnd.n5770 gnd.n2801 242.672
R5914 gnd.n5770 gnd.n2802 242.672
R5915 gnd.n5770 gnd.n2803 242.672
R5916 gnd.n5770 gnd.n2804 242.672
R5917 gnd.n5770 gnd.n2805 242.672
R5918 gnd.n5770 gnd.n2806 242.672
R5919 gnd.n5770 gnd.n2807 242.672
R5920 gnd.n5770 gnd.n2808 242.672
R5921 gnd.n5770 gnd.n2809 242.672
R5922 gnd.n5770 gnd.n2810 242.672
R5923 gnd.n172 gnd.n102 242.672
R5924 gnd.n7373 gnd.n102 242.672
R5925 gnd.n168 gnd.n102 242.672
R5926 gnd.n7380 gnd.n102 242.672
R5927 gnd.n161 gnd.n102 242.672
R5928 gnd.n7387 gnd.n102 242.672
R5929 gnd.n154 gnd.n102 242.672
R5930 gnd.n7394 gnd.n102 242.672
R5931 gnd.n147 gnd.n102 242.672
R5932 gnd.n7401 gnd.n102 242.672
R5933 gnd.n140 gnd.n102 242.672
R5934 gnd.n7411 gnd.n102 242.672
R5935 gnd.n133 gnd.n102 242.672
R5936 gnd.n7418 gnd.n102 242.672
R5937 gnd.n126 gnd.n102 242.672
R5938 gnd.n7425 gnd.n102 242.672
R5939 gnd.n119 gnd.n102 242.672
R5940 gnd.n7432 gnd.n102 242.672
R5941 gnd.n112 gnd.n102 242.672
R5942 gnd.n4624 gnd.n3528 242.672
R5943 gnd.n4624 gnd.n3529 242.672
R5944 gnd.n4624 gnd.n3530 242.672
R5945 gnd.n4624 gnd.n3531 242.672
R5946 gnd.n4624 gnd.n3532 242.672
R5947 gnd.n4624 gnd.n3533 242.672
R5948 gnd.n4624 gnd.n3534 242.672
R5949 gnd.n4624 gnd.n3535 242.672
R5950 gnd.n4624 gnd.n3536 242.672
R5951 gnd.n4624 gnd.n3537 242.672
R5952 gnd.n4624 gnd.n3538 242.672
R5953 gnd.n4624 gnd.n3539 242.672
R5954 gnd.n4624 gnd.n3540 242.672
R5955 gnd.n4624 gnd.n3541 242.672
R5956 gnd.n5450 gnd.n2785 242.672
R5957 gnd.n3216 gnd.n2785 242.672
R5958 gnd.n3213 gnd.n2785 242.672
R5959 gnd.n3208 gnd.n2785 242.672
R5960 gnd.n3205 gnd.n2785 242.672
R5961 gnd.n3202 gnd.n2785 242.672
R5962 gnd.n3189 gnd.n2785 242.672
R5963 gnd.n3187 gnd.n2785 242.672
R5964 gnd.n3172 gnd.n2785 242.672
R5965 gnd.n3170 gnd.n2785 242.672
R5966 gnd.n3155 gnd.n2785 242.672
R5967 gnd.n3153 gnd.n2785 242.672
R5968 gnd.n3138 gnd.n2785 242.672
R5969 gnd.n3136 gnd.n2785 242.672
R5970 gnd.n109 gnd.n105 240.244
R5971 gnd.n7434 gnd.n7433 240.244
R5972 gnd.n7431 gnd.n113 240.244
R5973 gnd.n7427 gnd.n7426 240.244
R5974 gnd.n7424 gnd.n120 240.244
R5975 gnd.n7420 gnd.n7419 240.244
R5976 gnd.n7417 gnd.n127 240.244
R5977 gnd.n7413 gnd.n7412 240.244
R5978 gnd.n7410 gnd.n134 240.244
R5979 gnd.n7403 gnd.n7402 240.244
R5980 gnd.n7400 gnd.n141 240.244
R5981 gnd.n7396 gnd.n7395 240.244
R5982 gnd.n7393 gnd.n148 240.244
R5983 gnd.n7389 gnd.n7388 240.244
R5984 gnd.n7386 gnd.n155 240.244
R5985 gnd.n7382 gnd.n7381 240.244
R5986 gnd.n7379 gnd.n162 240.244
R5987 gnd.n7375 gnd.n7374 240.244
R5988 gnd.n7372 gnd.n169 240.244
R5989 gnd.n5695 gnd.n2870 240.244
R5990 gnd.n3078 gnd.n2870 240.244
R5991 gnd.n3078 gnd.n3020 240.244
R5992 gnd.n3074 gnd.n3020 240.244
R5993 gnd.n3074 gnd.n3010 240.244
R5994 gnd.n3071 gnd.n3010 240.244
R5995 gnd.n3071 gnd.n3002 240.244
R5996 gnd.n3002 gnd.n2991 240.244
R5997 gnd.n3067 gnd.n2991 240.244
R5998 gnd.n3067 gnd.n2982 240.244
R5999 gnd.n3064 gnd.n2982 240.244
R6000 gnd.n3064 gnd.n2974 240.244
R6001 gnd.n2974 gnd.n2963 240.244
R6002 gnd.n3060 gnd.n2963 240.244
R6003 gnd.n3060 gnd.n2953 240.244
R6004 gnd.n2953 gnd.n2945 240.244
R6005 gnd.n5585 gnd.n2945 240.244
R6006 gnd.n5585 gnd.n2911 240.244
R6007 gnd.n5588 gnd.n2911 240.244
R6008 gnd.n5588 gnd.n2902 240.244
R6009 gnd.n5596 gnd.n2902 240.244
R6010 gnd.n5596 gnd.n274 240.244
R6011 gnd.n5610 gnd.n274 240.244
R6012 gnd.n5611 gnd.n5610 240.244
R6013 gnd.n5611 gnd.n2927 240.244
R6014 gnd.n5617 gnd.n2927 240.244
R6015 gnd.n5617 gnd.n294 240.244
R6016 gnd.n7178 gnd.n294 240.244
R6017 gnd.n7178 gnd.n291 240.244
R6018 gnd.n7174 gnd.n291 240.244
R6019 gnd.n7174 gnd.n259 240.244
R6020 gnd.n311 gnd.n259 240.244
R6021 gnd.n311 gnd.n253 240.244
R6022 gnd.n7161 gnd.n253 240.244
R6023 gnd.n7161 gnd.n245 240.244
R6024 gnd.n7157 gnd.n245 240.244
R6025 gnd.n7157 gnd.n237 240.244
R6026 gnd.n7153 gnd.n237 240.244
R6027 gnd.n7153 gnd.n229 240.244
R6028 gnd.n343 gnd.n229 240.244
R6029 gnd.n343 gnd.n223 240.244
R6030 gnd.n7141 gnd.n223 240.244
R6031 gnd.n7141 gnd.n215 240.244
R6032 gnd.n7137 gnd.n215 240.244
R6033 gnd.n7137 gnd.n207 240.244
R6034 gnd.n7133 gnd.n207 240.244
R6035 gnd.n7133 gnd.n199 240.244
R6036 gnd.n360 gnd.n199 240.244
R6037 gnd.n360 gnd.n190 240.244
R6038 gnd.n190 gnd.n179 240.244
R6039 gnd.n7363 gnd.n179 240.244
R6040 gnd.n7364 gnd.n7363 240.244
R6041 gnd.n7364 gnd.n101 240.244
R6042 gnd.n2823 gnd.n2822 240.244
R6043 gnd.n5763 gnd.n2822 240.244
R6044 gnd.n5761 gnd.n5760 240.244
R6045 gnd.n5757 gnd.n5756 240.244
R6046 gnd.n5753 gnd.n5752 240.244
R6047 gnd.n5749 gnd.n5748 240.244
R6048 gnd.n5745 gnd.n5744 240.244
R6049 gnd.n5741 gnd.n5740 240.244
R6050 gnd.n5736 gnd.n5735 240.244
R6051 gnd.n5732 gnd.n5731 240.244
R6052 gnd.n5728 gnd.n5727 240.244
R6053 gnd.n5724 gnd.n5723 240.244
R6054 gnd.n5720 gnd.n5719 240.244
R6055 gnd.n5716 gnd.n5715 240.244
R6056 gnd.n5712 gnd.n5711 240.244
R6057 gnd.n5708 gnd.n5707 240.244
R6058 gnd.n5704 gnd.n5703 240.244
R6059 gnd.n2865 gnd.n2864 240.244
R6060 gnd.n3040 gnd.n2824 240.244
R6061 gnd.n3040 gnd.n3018 240.244
R6062 gnd.n5492 gnd.n3018 240.244
R6063 gnd.n5492 gnd.n3013 240.244
R6064 gnd.n5500 gnd.n3013 240.244
R6065 gnd.n5500 gnd.n3014 240.244
R6066 gnd.n3014 gnd.n2989 240.244
R6067 gnd.n5523 gnd.n2989 240.244
R6068 gnd.n5523 gnd.n2984 240.244
R6069 gnd.n5531 gnd.n2984 240.244
R6070 gnd.n5531 gnd.n2985 240.244
R6071 gnd.n2985 gnd.n2961 240.244
R6072 gnd.n5562 gnd.n2961 240.244
R6073 gnd.n5562 gnd.n2955 240.244
R6074 gnd.n5570 gnd.n2955 240.244
R6075 gnd.n5570 gnd.n2957 240.244
R6076 gnd.n2957 gnd.n2909 240.244
R6077 gnd.n5652 gnd.n2909 240.244
R6078 gnd.n5652 gnd.n2905 240.244
R6079 gnd.n5658 gnd.n2905 240.244
R6080 gnd.n5658 gnd.n271 240.244
R6081 gnd.n7201 gnd.n271 240.244
R6082 gnd.n7201 gnd.n272 240.244
R6083 gnd.n2929 gnd.n272 240.244
R6084 gnd.n5635 gnd.n2929 240.244
R6085 gnd.n5635 gnd.n5633 240.244
R6086 gnd.n5633 gnd.n293 240.244
R6087 gnd.n7180 gnd.n293 240.244
R6088 gnd.n7183 gnd.n7180 240.244
R6089 gnd.n7183 gnd.n261 240.244
R6090 gnd.n7206 gnd.n261 240.244
R6091 gnd.n7206 gnd.n251 240.244
R6092 gnd.n7216 gnd.n251 240.244
R6093 gnd.n7216 gnd.n247 240.244
R6094 gnd.n7222 gnd.n247 240.244
R6095 gnd.n7222 gnd.n235 240.244
R6096 gnd.n7232 gnd.n235 240.244
R6097 gnd.n7232 gnd.n231 240.244
R6098 gnd.n7238 gnd.n231 240.244
R6099 gnd.n7238 gnd.n221 240.244
R6100 gnd.n7248 gnd.n221 240.244
R6101 gnd.n7248 gnd.n217 240.244
R6102 gnd.n7254 gnd.n217 240.244
R6103 gnd.n7254 gnd.n205 240.244
R6104 gnd.n7264 gnd.n205 240.244
R6105 gnd.n7264 gnd.n201 240.244
R6106 gnd.n7270 gnd.n201 240.244
R6107 gnd.n7270 gnd.n188 240.244
R6108 gnd.n7355 gnd.n188 240.244
R6109 gnd.n7355 gnd.n184 240.244
R6110 gnd.n7361 gnd.n184 240.244
R6111 gnd.n7361 gnd.n104 240.244
R6112 gnd.n7441 gnd.n104 240.244
R6113 gnd.n3685 gnd.n2668 240.244
R6114 gnd.n4588 gnd.n3686 240.244
R6115 gnd.n4584 gnd.n4583 240.244
R6116 gnd.n4580 gnd.n4579 240.244
R6117 gnd.n4576 gnd.n4575 240.244
R6118 gnd.n4572 gnd.n4571 240.244
R6119 gnd.n4568 gnd.n4567 240.244
R6120 gnd.n4564 gnd.n4563 240.244
R6121 gnd.n4300 gnd.n4299 240.244
R6122 gnd.n4297 gnd.n4296 240.244
R6123 gnd.n4293 gnd.n4292 240.244
R6124 gnd.n4289 gnd.n4288 240.244
R6125 gnd.n4285 gnd.n4284 240.244
R6126 gnd.n4281 gnd.n4280 240.244
R6127 gnd.n4277 gnd.n4276 240.244
R6128 gnd.n4273 gnd.n4272 240.244
R6129 gnd.n4269 gnd.n4268 240.244
R6130 gnd.n4265 gnd.n4264 240.244
R6131 gnd.n6069 gnd.n2399 240.244
R6132 gnd.n2403 gnd.n2399 240.244
R6133 gnd.n6062 gnd.n2403 240.244
R6134 gnd.n6062 gnd.n2404 240.244
R6135 gnd.n2418 gnd.n2404 240.244
R6136 gnd.n4067 gnd.n2418 240.244
R6137 gnd.n4067 gnd.n2430 240.244
R6138 gnd.n4077 gnd.n2430 240.244
R6139 gnd.n4077 gnd.n2441 240.244
R6140 gnd.n4083 gnd.n2441 240.244
R6141 gnd.n4083 gnd.n2451 240.244
R6142 gnd.n4093 gnd.n2451 240.244
R6143 gnd.n4093 gnd.n2462 240.244
R6144 gnd.n4099 gnd.n2462 240.244
R6145 gnd.n4099 gnd.n2473 240.244
R6146 gnd.n4109 gnd.n2473 240.244
R6147 gnd.n4109 gnd.n2484 240.244
R6148 gnd.n4115 gnd.n2484 240.244
R6149 gnd.n4115 gnd.n2494 240.244
R6150 gnd.n4125 gnd.n2494 240.244
R6151 gnd.n4125 gnd.n2505 240.244
R6152 gnd.n4131 gnd.n2505 240.244
R6153 gnd.n4131 gnd.n2516 240.244
R6154 gnd.n4141 gnd.n2516 240.244
R6155 gnd.n4141 gnd.n2525 240.244
R6156 gnd.n4149 gnd.n2525 240.244
R6157 gnd.n4149 gnd.n2535 240.244
R6158 gnd.n4160 gnd.n2535 240.244
R6159 gnd.n4160 gnd.n2543 240.244
R6160 gnd.n4166 gnd.n2543 240.244
R6161 gnd.n4166 gnd.n2554 240.244
R6162 gnd.n4176 gnd.n2554 240.244
R6163 gnd.n4176 gnd.n2564 240.244
R6164 gnd.n4182 gnd.n2564 240.244
R6165 gnd.n4182 gnd.n2574 240.244
R6166 gnd.n4192 gnd.n2574 240.244
R6167 gnd.n4192 gnd.n2585 240.244
R6168 gnd.n4198 gnd.n2585 240.244
R6169 gnd.n4198 gnd.n2596 240.244
R6170 gnd.n4208 gnd.n2596 240.244
R6171 gnd.n4208 gnd.n2607 240.244
R6172 gnd.n4214 gnd.n2607 240.244
R6173 gnd.n4214 gnd.n2617 240.244
R6174 gnd.n4224 gnd.n2617 240.244
R6175 gnd.n4224 gnd.n2628 240.244
R6176 gnd.n4230 gnd.n2628 240.244
R6177 gnd.n4230 gnd.n2639 240.244
R6178 gnd.n4240 gnd.n2639 240.244
R6179 gnd.n4240 gnd.n2650 240.244
R6180 gnd.n4247 gnd.n2650 240.244
R6181 gnd.n4247 gnd.n2661 240.244
R6182 gnd.n4257 gnd.n2661 240.244
R6183 gnd.n4257 gnd.n2670 240.244
R6184 gnd.n2353 gnd.n2352 240.244
R6185 gnd.n6141 gnd.n2352 240.244
R6186 gnd.n6139 gnd.n6138 240.244
R6187 gnd.n6135 gnd.n6134 240.244
R6188 gnd.n6131 gnd.n6130 240.244
R6189 gnd.n6127 gnd.n6126 240.244
R6190 gnd.n6123 gnd.n6122 240.244
R6191 gnd.n6119 gnd.n6118 240.244
R6192 gnd.n6115 gnd.n6114 240.244
R6193 gnd.n6110 gnd.n6109 240.244
R6194 gnd.n6106 gnd.n6105 240.244
R6195 gnd.n6102 gnd.n6101 240.244
R6196 gnd.n6098 gnd.n6097 240.244
R6197 gnd.n6094 gnd.n6093 240.244
R6198 gnd.n6090 gnd.n6089 240.244
R6199 gnd.n6086 gnd.n6085 240.244
R6200 gnd.n6082 gnd.n6081 240.244
R6201 gnd.n6078 gnd.n6077 240.244
R6202 gnd.n2394 gnd.n2393 240.244
R6203 gnd.n4051 gnd.n2354 240.244
R6204 gnd.n4051 gnd.n2409 240.244
R6205 gnd.n6060 gnd.n2409 240.244
R6206 gnd.n6060 gnd.n2410 240.244
R6207 gnd.n6056 gnd.n2410 240.244
R6208 gnd.n6056 gnd.n2416 240.244
R6209 gnd.n6048 gnd.n2416 240.244
R6210 gnd.n6048 gnd.n2433 240.244
R6211 gnd.n6044 gnd.n2433 240.244
R6212 gnd.n6044 gnd.n2439 240.244
R6213 gnd.n6036 gnd.n2439 240.244
R6214 gnd.n6036 gnd.n2454 240.244
R6215 gnd.n6032 gnd.n2454 240.244
R6216 gnd.n6032 gnd.n2460 240.244
R6217 gnd.n6024 gnd.n2460 240.244
R6218 gnd.n6024 gnd.n2476 240.244
R6219 gnd.n6020 gnd.n2476 240.244
R6220 gnd.n6020 gnd.n2482 240.244
R6221 gnd.n6012 gnd.n2482 240.244
R6222 gnd.n6012 gnd.n2497 240.244
R6223 gnd.n6008 gnd.n2497 240.244
R6224 gnd.n6008 gnd.n2503 240.244
R6225 gnd.n6000 gnd.n2503 240.244
R6226 gnd.n6000 gnd.n2519 240.244
R6227 gnd.n5996 gnd.n2519 240.244
R6228 gnd.n5996 gnd.n2523 240.244
R6229 gnd.n5988 gnd.n2523 240.244
R6230 gnd.n5988 gnd.n2538 240.244
R6231 gnd.n5983 gnd.n2538 240.244
R6232 gnd.n5983 gnd.n2541 240.244
R6233 gnd.n5975 gnd.n2541 240.244
R6234 gnd.n5975 gnd.n2557 240.244
R6235 gnd.n5971 gnd.n2557 240.244
R6236 gnd.n5971 gnd.n2562 240.244
R6237 gnd.n5963 gnd.n2562 240.244
R6238 gnd.n5963 gnd.n2577 240.244
R6239 gnd.n5959 gnd.n2577 240.244
R6240 gnd.n5959 gnd.n2583 240.244
R6241 gnd.n5951 gnd.n2583 240.244
R6242 gnd.n5951 gnd.n2599 240.244
R6243 gnd.n5947 gnd.n2599 240.244
R6244 gnd.n5947 gnd.n2605 240.244
R6245 gnd.n5939 gnd.n2605 240.244
R6246 gnd.n5939 gnd.n2620 240.244
R6247 gnd.n5935 gnd.n2620 240.244
R6248 gnd.n5935 gnd.n2626 240.244
R6249 gnd.n5927 gnd.n2626 240.244
R6250 gnd.n5927 gnd.n2642 240.244
R6251 gnd.n5923 gnd.n2642 240.244
R6252 gnd.n5923 gnd.n2648 240.244
R6253 gnd.n5915 gnd.n2648 240.244
R6254 gnd.n5915 gnd.n2663 240.244
R6255 gnd.n5911 gnd.n2663 240.244
R6256 gnd.n6194 gnd.n6155 240.244
R6257 gnd.n6187 gnd.n6186 240.244
R6258 gnd.n6184 gnd.n6183 240.244
R6259 gnd.n6180 gnd.n6179 240.244
R6260 gnd.n6176 gnd.n6175 240.244
R6261 gnd.n6172 gnd.n6171 240.244
R6262 gnd.n6168 gnd.n1056 240.244
R6263 gnd.n6198 gnd.n6197 240.244
R6264 gnd.n1706 gnd.n1418 240.244
R6265 gnd.n1716 gnd.n1418 240.244
R6266 gnd.n1716 gnd.n1409 240.244
R6267 gnd.n1409 gnd.n1398 240.244
R6268 gnd.n1737 gnd.n1398 240.244
R6269 gnd.n1737 gnd.n1392 240.244
R6270 gnd.n1747 gnd.n1392 240.244
R6271 gnd.n1747 gnd.n1381 240.244
R6272 gnd.n1381 gnd.n1373 240.244
R6273 gnd.n1765 gnd.n1373 240.244
R6274 gnd.n1766 gnd.n1765 240.244
R6275 gnd.n1766 gnd.n1358 240.244
R6276 gnd.n1768 gnd.n1358 240.244
R6277 gnd.n1768 gnd.n1344 240.244
R6278 gnd.n1810 gnd.n1344 240.244
R6279 gnd.n1811 gnd.n1810 240.244
R6280 gnd.n1814 gnd.n1811 240.244
R6281 gnd.n1814 gnd.n1299 240.244
R6282 gnd.n1339 gnd.n1299 240.244
R6283 gnd.n1339 gnd.n1309 240.244
R6284 gnd.n1824 gnd.n1309 240.244
R6285 gnd.n1824 gnd.n1330 240.244
R6286 gnd.n1834 gnd.n1330 240.244
R6287 gnd.n1834 gnd.n1228 240.244
R6288 gnd.n1879 gnd.n1228 240.244
R6289 gnd.n1879 gnd.n1214 240.244
R6290 gnd.n1901 gnd.n1214 240.244
R6291 gnd.n1902 gnd.n1901 240.244
R6292 gnd.n1902 gnd.n1201 240.244
R6293 gnd.n1201 gnd.n1190 240.244
R6294 gnd.n1933 gnd.n1190 240.244
R6295 gnd.n1934 gnd.n1933 240.244
R6296 gnd.n1935 gnd.n1934 240.244
R6297 gnd.n1935 gnd.n1175 240.244
R6298 gnd.n1937 gnd.n1175 240.244
R6299 gnd.n1937 gnd.n1160 240.244
R6300 gnd.n2019 gnd.n1160 240.244
R6301 gnd.n2020 gnd.n2019 240.244
R6302 gnd.n2021 gnd.n2020 240.244
R6303 gnd.n2021 gnd.n979 240.244
R6304 gnd.n1155 gnd.n979 240.244
R6305 gnd.n1155 gnd.n990 240.244
R6306 gnd.n2033 gnd.n990 240.244
R6307 gnd.n2034 gnd.n2033 240.244
R6308 gnd.n2034 gnd.n1003 240.244
R6309 gnd.n1152 gnd.n1003 240.244
R6310 gnd.n1152 gnd.n1016 240.244
R6311 gnd.n2302 gnd.n1016 240.244
R6312 gnd.n2303 gnd.n2302 240.244
R6313 gnd.n2303 gnd.n1029 240.244
R6314 gnd.n2311 gnd.n1029 240.244
R6315 gnd.n2311 gnd.n1041 240.244
R6316 gnd.n6205 gnd.n1041 240.244
R6317 gnd.n1696 gnd.n1431 240.244
R6318 gnd.n1452 gnd.n1431 240.244
R6319 gnd.n1455 gnd.n1454 240.244
R6320 gnd.n1462 gnd.n1461 240.244
R6321 gnd.n1465 gnd.n1464 240.244
R6322 gnd.n1472 gnd.n1471 240.244
R6323 gnd.n1475 gnd.n1474 240.244
R6324 gnd.n1482 gnd.n1481 240.244
R6325 gnd.n1704 gnd.n1428 240.244
R6326 gnd.n1428 gnd.n1407 240.244
R6327 gnd.n1727 gnd.n1407 240.244
R6328 gnd.n1727 gnd.n1401 240.244
R6329 gnd.n1735 gnd.n1401 240.244
R6330 gnd.n1735 gnd.n1403 240.244
R6331 gnd.n1403 gnd.n1379 240.244
R6332 gnd.n1757 gnd.n1379 240.244
R6333 gnd.n1757 gnd.n1375 240.244
R6334 gnd.n1763 gnd.n1375 240.244
R6335 gnd.n1763 gnd.n1357 240.244
R6336 gnd.n1788 gnd.n1357 240.244
R6337 gnd.n1788 gnd.n1352 240.244
R6338 gnd.n1800 gnd.n1352 240.244
R6339 gnd.n1800 gnd.n1353 240.244
R6340 gnd.n1796 gnd.n1353 240.244
R6341 gnd.n1796 gnd.n1301 240.244
R6342 gnd.n1848 gnd.n1301 240.244
R6343 gnd.n1848 gnd.n1302 240.244
R6344 gnd.n1844 gnd.n1302 240.244
R6345 gnd.n1844 gnd.n1308 240.244
R6346 gnd.n1328 gnd.n1308 240.244
R6347 gnd.n1328 gnd.n1226 240.244
R6348 gnd.n1883 gnd.n1226 240.244
R6349 gnd.n1883 gnd.n1221 240.244
R6350 gnd.n1891 gnd.n1221 240.244
R6351 gnd.n1891 gnd.n1222 240.244
R6352 gnd.n1222 gnd.n1199 240.244
R6353 gnd.n1923 gnd.n1199 240.244
R6354 gnd.n1923 gnd.n1194 240.244
R6355 gnd.n1931 gnd.n1194 240.244
R6356 gnd.n1931 gnd.n1195 240.244
R6357 gnd.n1195 gnd.n1173 240.244
R6358 gnd.n1997 gnd.n1173 240.244
R6359 gnd.n1997 gnd.n1168 240.244
R6360 gnd.n2009 gnd.n1168 240.244
R6361 gnd.n2009 gnd.n1169 240.244
R6362 gnd.n2005 gnd.n1169 240.244
R6363 gnd.n2005 gnd.n981 240.244
R6364 gnd.n6245 gnd.n981 240.244
R6365 gnd.n6245 gnd.n982 240.244
R6366 gnd.n6241 gnd.n982 240.244
R6367 gnd.n6241 gnd.n988 240.244
R6368 gnd.n1005 gnd.n988 240.244
R6369 gnd.n6231 gnd.n1005 240.244
R6370 gnd.n6231 gnd.n1006 240.244
R6371 gnd.n6227 gnd.n1006 240.244
R6372 gnd.n6227 gnd.n1014 240.244
R6373 gnd.n1030 gnd.n1014 240.244
R6374 gnd.n6217 gnd.n1030 240.244
R6375 gnd.n6217 gnd.n1031 240.244
R6376 gnd.n6213 gnd.n1031 240.244
R6377 gnd.n6213 gnd.n1039 240.244
R6378 gnd.n1085 gnd.n1045 240.244
R6379 gnd.n1093 gnd.n1092 240.244
R6380 gnd.n1096 gnd.n1095 240.244
R6381 gnd.n1103 gnd.n1102 240.244
R6382 gnd.n1106 gnd.n1105 240.244
R6383 gnd.n1113 gnd.n1112 240.244
R6384 gnd.n1116 gnd.n1115 240.244
R6385 gnd.n1123 gnd.n1122 240.244
R6386 gnd.n1126 gnd.n1125 240.244
R6387 gnd.n1133 gnd.n1132 240.244
R6388 gnd.n1136 gnd.n1135 240.244
R6389 gnd.n1143 gnd.n1142 240.244
R6390 gnd.n1145 gnd.n1069 240.244
R6391 gnd.n1619 gnd.n1516 240.244
R6392 gnd.n1619 gnd.n1509 240.244
R6393 gnd.n1630 gnd.n1509 240.244
R6394 gnd.n1630 gnd.n1505 240.244
R6395 gnd.n1636 gnd.n1505 240.244
R6396 gnd.n1636 gnd.n1497 240.244
R6397 gnd.n1646 gnd.n1497 240.244
R6398 gnd.n1646 gnd.n1492 240.244
R6399 gnd.n1682 gnd.n1492 240.244
R6400 gnd.n1682 gnd.n1493 240.244
R6401 gnd.n1493 gnd.n1440 240.244
R6402 gnd.n1677 gnd.n1440 240.244
R6403 gnd.n1677 gnd.n1676 240.244
R6404 gnd.n1676 gnd.n1419 240.244
R6405 gnd.n1672 gnd.n1419 240.244
R6406 gnd.n1672 gnd.n1410 240.244
R6407 gnd.n1669 gnd.n1410 240.244
R6408 gnd.n1669 gnd.n1668 240.244
R6409 gnd.n1668 gnd.n1393 240.244
R6410 gnd.n1664 gnd.n1393 240.244
R6411 gnd.n1664 gnd.n1382 240.244
R6412 gnd.n1382 gnd.n1363 240.244
R6413 gnd.n1777 gnd.n1363 240.244
R6414 gnd.n1777 gnd.n1359 240.244
R6415 gnd.n1785 gnd.n1359 240.244
R6416 gnd.n1785 gnd.n1350 240.244
R6417 gnd.n1350 gnd.n1286 240.244
R6418 gnd.n1857 gnd.n1286 240.244
R6419 gnd.n1857 gnd.n1287 240.244
R6420 gnd.n1298 gnd.n1287 240.244
R6421 gnd.n1333 gnd.n1298 240.244
R6422 gnd.n1336 gnd.n1333 240.244
R6423 gnd.n1336 gnd.n1310 240.244
R6424 gnd.n1323 gnd.n1310 240.244
R6425 gnd.n1323 gnd.n1320 240.244
R6426 gnd.n1320 gnd.n1229 240.244
R6427 gnd.n1878 gnd.n1229 240.244
R6428 gnd.n1878 gnd.n1219 240.244
R6429 gnd.n1874 gnd.n1219 240.244
R6430 gnd.n1874 gnd.n1213 240.244
R6431 gnd.n1871 gnd.n1213 240.244
R6432 gnd.n1871 gnd.n1202 240.244
R6433 gnd.n1868 gnd.n1202 240.244
R6434 gnd.n1868 gnd.n1180 240.244
R6435 gnd.n1946 gnd.n1180 240.244
R6436 gnd.n1946 gnd.n1176 240.244
R6437 gnd.n1994 gnd.n1176 240.244
R6438 gnd.n1994 gnd.n1166 240.244
R6439 gnd.n1990 gnd.n1166 240.244
R6440 gnd.n1990 gnd.n967 240.244
R6441 gnd.n1987 gnd.n967 240.244
R6442 gnd.n1987 gnd.n978 240.244
R6443 gnd.n1983 gnd.n978 240.244
R6444 gnd.n1983 gnd.n1982 240.244
R6445 gnd.n1982 gnd.n991 240.244
R6446 gnd.n1978 gnd.n991 240.244
R6447 gnd.n1978 gnd.n1002 240.244
R6448 gnd.n1974 gnd.n1002 240.244
R6449 gnd.n1974 gnd.n1973 240.244
R6450 gnd.n1973 gnd.n1017 240.244
R6451 gnd.n1969 gnd.n1017 240.244
R6452 gnd.n1969 gnd.n1028 240.244
R6453 gnd.n2314 gnd.n1028 240.244
R6454 gnd.n2315 gnd.n2314 240.244
R6455 gnd.n2315 gnd.n1042 240.244
R6456 gnd.n1533 gnd.n1532 240.244
R6457 gnd.n1604 gnd.n1532 240.244
R6458 gnd.n1602 gnd.n1601 240.244
R6459 gnd.n1598 gnd.n1597 240.244
R6460 gnd.n1594 gnd.n1593 240.244
R6461 gnd.n1590 gnd.n1589 240.244
R6462 gnd.n1586 gnd.n1585 240.244
R6463 gnd.n1582 gnd.n1581 240.244
R6464 gnd.n1578 gnd.n1577 240.244
R6465 gnd.n1574 gnd.n1573 240.244
R6466 gnd.n1570 gnd.n1569 240.244
R6467 gnd.n1566 gnd.n1565 240.244
R6468 gnd.n1562 gnd.n1520 240.244
R6469 gnd.n1622 gnd.n1514 240.244
R6470 gnd.n1622 gnd.n1510 240.244
R6471 gnd.n1628 gnd.n1510 240.244
R6472 gnd.n1628 gnd.n1503 240.244
R6473 gnd.n1638 gnd.n1503 240.244
R6474 gnd.n1638 gnd.n1499 240.244
R6475 gnd.n1644 gnd.n1499 240.244
R6476 gnd.n1644 gnd.n1490 240.244
R6477 gnd.n1684 gnd.n1490 240.244
R6478 gnd.n1684 gnd.n1441 240.244
R6479 gnd.n1692 gnd.n1441 240.244
R6480 gnd.n1692 gnd.n1442 240.244
R6481 gnd.n1442 gnd.n1420 240.244
R6482 gnd.n1713 gnd.n1420 240.244
R6483 gnd.n1713 gnd.n1412 240.244
R6484 gnd.n1724 gnd.n1412 240.244
R6485 gnd.n1724 gnd.n1413 240.244
R6486 gnd.n1413 gnd.n1394 240.244
R6487 gnd.n1744 gnd.n1394 240.244
R6488 gnd.n1744 gnd.n1384 240.244
R6489 gnd.n1754 gnd.n1384 240.244
R6490 gnd.n1754 gnd.n1365 240.244
R6491 gnd.n1775 gnd.n1365 240.244
R6492 gnd.n1775 gnd.n1367 240.244
R6493 gnd.n1367 gnd.n1348 240.244
R6494 gnd.n1803 gnd.n1348 240.244
R6495 gnd.n1803 gnd.n1290 240.244
R6496 gnd.n1855 gnd.n1290 240.244
R6497 gnd.n1855 gnd.n1291 240.244
R6498 gnd.n1851 gnd.n1291 240.244
R6499 gnd.n1851 gnd.n1297 240.244
R6500 gnd.n1312 gnd.n1297 240.244
R6501 gnd.n1841 gnd.n1312 240.244
R6502 gnd.n1841 gnd.n1313 240.244
R6503 gnd.n1837 gnd.n1313 240.244
R6504 gnd.n1837 gnd.n1319 240.244
R6505 gnd.n1319 gnd.n1218 240.244
R6506 gnd.n1894 gnd.n1218 240.244
R6507 gnd.n1894 gnd.n1211 240.244
R6508 gnd.n1905 gnd.n1211 240.244
R6509 gnd.n1905 gnd.n1204 240.244
R6510 gnd.n1920 gnd.n1204 240.244
R6511 gnd.n1920 gnd.n1205 240.244
R6512 gnd.n1205 gnd.n1183 240.244
R6513 gnd.n1944 gnd.n1183 240.244
R6514 gnd.n1944 gnd.n1184 240.244
R6515 gnd.n1184 gnd.n1164 240.244
R6516 gnd.n2012 gnd.n1164 240.244
R6517 gnd.n2012 gnd.n969 240.244
R6518 gnd.n6252 gnd.n969 240.244
R6519 gnd.n6252 gnd.n970 240.244
R6520 gnd.n6248 gnd.n970 240.244
R6521 gnd.n6248 gnd.n976 240.244
R6522 gnd.n993 gnd.n976 240.244
R6523 gnd.n6238 gnd.n993 240.244
R6524 gnd.n6238 gnd.n994 240.244
R6525 gnd.n6234 gnd.n994 240.244
R6526 gnd.n6234 gnd.n1000 240.244
R6527 gnd.n1019 gnd.n1000 240.244
R6528 gnd.n6224 gnd.n1019 240.244
R6529 gnd.n6224 gnd.n1020 240.244
R6530 gnd.n6220 gnd.n1020 240.244
R6531 gnd.n6220 gnd.n1026 240.244
R6532 gnd.n1044 gnd.n1026 240.244
R6533 gnd.n6210 gnd.n1044 240.244
R6534 gnd.n7280 gnd.n7279 240.244
R6535 gnd.n7285 gnd.n7282 240.244
R6536 gnd.n7288 gnd.n7287 240.244
R6537 gnd.n7293 gnd.n7290 240.244
R6538 gnd.n7296 gnd.n7295 240.244
R6539 gnd.n7301 gnd.n7298 240.244
R6540 gnd.n7304 gnd.n7303 240.244
R6541 gnd.n7309 gnd.n7306 240.244
R6542 gnd.n7315 gnd.n7311 240.244
R6543 gnd.n3079 gnd.n2873 240.244
R6544 gnd.n5478 gnd.n3079 240.244
R6545 gnd.n5478 gnd.n3021 240.244
R6546 gnd.n3021 gnd.n3008 240.244
R6547 gnd.n5502 gnd.n3008 240.244
R6548 gnd.n5502 gnd.n3003 240.244
R6549 gnd.n5509 gnd.n3003 240.244
R6550 gnd.n5509 gnd.n2992 240.244
R6551 gnd.n2992 gnd.n2980 240.244
R6552 gnd.n5533 gnd.n2980 240.244
R6553 gnd.n5533 gnd.n2975 240.244
R6554 gnd.n5540 gnd.n2975 240.244
R6555 gnd.n5540 gnd.n2964 240.244
R6556 gnd.n2964 gnd.n2952 240.244
R6557 gnd.n5572 gnd.n2952 240.244
R6558 gnd.n5572 gnd.n2947 240.244
R6559 gnd.n5582 gnd.n2947 240.244
R6560 gnd.n5582 gnd.n2912 240.244
R6561 gnd.n5576 gnd.n2912 240.244
R6562 gnd.n5576 gnd.n2903 240.244
R6563 gnd.n5598 gnd.n2903 240.244
R6564 gnd.n5598 gnd.n275 240.244
R6565 gnd.n5607 gnd.n275 240.244
R6566 gnd.n5607 gnd.n2936 240.244
R6567 gnd.n2936 gnd.n2928 240.244
R6568 gnd.n5618 gnd.n2928 240.244
R6569 gnd.n5618 gnd.n66 240.244
R6570 gnd.n67 gnd.n66 240.244
R6571 gnd.n68 gnd.n67 240.244
R6572 gnd.n301 gnd.n68 240.244
R6573 gnd.n301 gnd.n71 240.244
R6574 gnd.n72 gnd.n71 240.244
R6575 gnd.n73 gnd.n72 240.244
R6576 gnd.n7162 gnd.n73 240.244
R6577 gnd.n7162 gnd.n76 240.244
R6578 gnd.n77 gnd.n76 240.244
R6579 gnd.n78 gnd.n77 240.244
R6580 gnd.n321 gnd.n78 240.244
R6581 gnd.n321 gnd.n81 240.244
R6582 gnd.n82 gnd.n81 240.244
R6583 gnd.n83 gnd.n82 240.244
R6584 gnd.n7142 gnd.n83 240.244
R6585 gnd.n7142 gnd.n86 240.244
R6586 gnd.n87 gnd.n86 240.244
R6587 gnd.n88 gnd.n87 240.244
R6588 gnd.n363 gnd.n88 240.244
R6589 gnd.n363 gnd.n91 240.244
R6590 gnd.n92 gnd.n91 240.244
R6591 gnd.n93 gnd.n92 240.244
R6592 gnd.n180 gnd.n93 240.244
R6593 gnd.n180 gnd.n96 240.244
R6594 gnd.n97 gnd.n96 240.244
R6595 gnd.n7443 gnd.n97 240.244
R6596 gnd.n3131 gnd.n3130 240.244
R6597 gnd.n3122 gnd.n3121 240.244
R6598 gnd.n3147 gnd.n3146 240.244
R6599 gnd.n3113 gnd.n3112 240.244
R6600 gnd.n3164 gnd.n3163 240.244
R6601 gnd.n3104 gnd.n3103 240.244
R6602 gnd.n3181 gnd.n3180 240.244
R6603 gnd.n3095 gnd.n3094 240.244
R6604 gnd.n3090 gnd.n2820 240.244
R6605 gnd.n5693 gnd.n2876 240.244
R6606 gnd.n2880 gnd.n2876 240.244
R6607 gnd.n2881 gnd.n2880 240.244
R6608 gnd.n2882 gnd.n2881 240.244
R6609 gnd.n3012 gnd.n2882 240.244
R6610 gnd.n3012 gnd.n2885 240.244
R6611 gnd.n2886 gnd.n2885 240.244
R6612 gnd.n2887 gnd.n2886 240.244
R6613 gnd.n2993 gnd.n2887 240.244
R6614 gnd.n2993 gnd.n2890 240.244
R6615 gnd.n2891 gnd.n2890 240.244
R6616 gnd.n2892 gnd.n2891 240.244
R6617 gnd.n5560 gnd.n2892 240.244
R6618 gnd.n5560 gnd.n2895 240.244
R6619 gnd.n2896 gnd.n2895 240.244
R6620 gnd.n2897 gnd.n2896 240.244
R6621 gnd.n5583 gnd.n2897 240.244
R6622 gnd.n5583 gnd.n2900 240.244
R6623 gnd.n2901 gnd.n2900 240.244
R6624 gnd.n5660 gnd.n2901 240.244
R6625 gnd.n5660 gnd.n277 240.244
R6626 gnd.n7199 gnd.n277 240.244
R6627 gnd.n7199 gnd.n278 240.244
R6628 gnd.n283 gnd.n278 240.244
R6629 gnd.n284 gnd.n283 240.244
R6630 gnd.n285 gnd.n284 240.244
R6631 gnd.n5619 gnd.n285 240.244
R6632 gnd.n5619 gnd.n289 240.244
R6633 gnd.n7185 gnd.n289 240.244
R6634 gnd.n7185 gnd.n258 240.244
R6635 gnd.n7208 gnd.n258 240.244
R6636 gnd.n7208 gnd.n254 240.244
R6637 gnd.n7214 gnd.n254 240.244
R6638 gnd.n7214 gnd.n243 240.244
R6639 gnd.n7224 gnd.n243 240.244
R6640 gnd.n7224 gnd.n239 240.244
R6641 gnd.n7230 gnd.n239 240.244
R6642 gnd.n7230 gnd.n228 240.244
R6643 gnd.n7240 gnd.n228 240.244
R6644 gnd.n7240 gnd.n224 240.244
R6645 gnd.n7246 gnd.n224 240.244
R6646 gnd.n7246 gnd.n213 240.244
R6647 gnd.n7256 gnd.n213 240.244
R6648 gnd.n7256 gnd.n209 240.244
R6649 gnd.n7262 gnd.n209 240.244
R6650 gnd.n7262 gnd.n198 240.244
R6651 gnd.n7272 gnd.n198 240.244
R6652 gnd.n7272 gnd.n192 240.244
R6653 gnd.n7353 gnd.n192 240.244
R6654 gnd.n7353 gnd.n193 240.244
R6655 gnd.n193 gnd.n183 240.244
R6656 gnd.n7277 gnd.n183 240.244
R6657 gnd.n7277 gnd.n103 240.244
R6658 gnd.n3602 gnd.n2673 240.244
R6659 gnd.n3605 gnd.n3604 240.244
R6660 gnd.n3617 gnd.n3616 240.244
R6661 gnd.n3591 gnd.n3590 240.244
R6662 gnd.n3629 gnd.n3628 240.244
R6663 gnd.n3641 gnd.n3640 240.244
R6664 gnd.n3579 gnd.n3578 240.244
R6665 gnd.n3652 gnd.n3572 240.244
R6666 gnd.n3664 gnd.n3563 240.244
R6667 gnd.n4053 gnd.n3810 240.244
R6668 gnd.n4054 gnd.n4053 240.244
R6669 gnd.n4054 gnd.n2406 240.244
R6670 gnd.n4060 gnd.n2406 240.244
R6671 gnd.n4060 gnd.n2419 240.244
R6672 gnd.n4069 gnd.n2419 240.244
R6673 gnd.n4069 gnd.n2431 240.244
R6674 gnd.n4075 gnd.n2431 240.244
R6675 gnd.n4075 gnd.n2442 240.244
R6676 gnd.n4085 gnd.n2442 240.244
R6677 gnd.n4085 gnd.n2452 240.244
R6678 gnd.n4091 gnd.n2452 240.244
R6679 gnd.n4091 gnd.n2463 240.244
R6680 gnd.n4101 gnd.n2463 240.244
R6681 gnd.n4101 gnd.n2474 240.244
R6682 gnd.n4107 gnd.n2474 240.244
R6683 gnd.n4107 gnd.n2485 240.244
R6684 gnd.n4117 gnd.n2485 240.244
R6685 gnd.n4117 gnd.n2495 240.244
R6686 gnd.n4123 gnd.n2495 240.244
R6687 gnd.n4123 gnd.n2506 240.244
R6688 gnd.n4133 gnd.n2506 240.244
R6689 gnd.n4133 gnd.n2517 240.244
R6690 gnd.n4139 gnd.n2517 240.244
R6691 gnd.n4139 gnd.n2526 240.244
R6692 gnd.n4151 gnd.n2526 240.244
R6693 gnd.n4151 gnd.n2536 240.244
R6694 gnd.n4158 gnd.n2536 240.244
R6695 gnd.n4158 gnd.n2544 240.244
R6696 gnd.n4168 gnd.n2544 240.244
R6697 gnd.n4168 gnd.n2555 240.244
R6698 gnd.n4174 gnd.n2555 240.244
R6699 gnd.n4174 gnd.n2565 240.244
R6700 gnd.n4184 gnd.n2565 240.244
R6701 gnd.n4184 gnd.n2575 240.244
R6702 gnd.n4190 gnd.n2575 240.244
R6703 gnd.n4190 gnd.n2586 240.244
R6704 gnd.n4200 gnd.n2586 240.244
R6705 gnd.n4200 gnd.n2597 240.244
R6706 gnd.n4206 gnd.n2597 240.244
R6707 gnd.n4206 gnd.n2608 240.244
R6708 gnd.n4216 gnd.n2608 240.244
R6709 gnd.n4216 gnd.n2618 240.244
R6710 gnd.n4222 gnd.n2618 240.244
R6711 gnd.n4222 gnd.n2629 240.244
R6712 gnd.n4232 gnd.n2629 240.244
R6713 gnd.n4232 gnd.n2640 240.244
R6714 gnd.n4238 gnd.n2640 240.244
R6715 gnd.n4238 gnd.n2651 240.244
R6716 gnd.n4249 gnd.n2651 240.244
R6717 gnd.n4249 gnd.n2662 240.244
R6718 gnd.n4255 gnd.n2662 240.244
R6719 gnd.n4255 gnd.n2671 240.244
R6720 gnd.n4033 gnd.n4032 240.244
R6721 gnd.n4029 gnd.n4028 240.244
R6722 gnd.n4025 gnd.n4024 240.244
R6723 gnd.n4021 gnd.n4020 240.244
R6724 gnd.n4017 gnd.n4016 240.244
R6725 gnd.n4013 gnd.n4012 240.244
R6726 gnd.n4009 gnd.n4008 240.244
R6727 gnd.n4005 gnd.n4004 240.244
R6728 gnd.n3993 gnd.n2350 240.244
R6729 gnd.n4045 gnd.n3974 240.244
R6730 gnd.n4045 gnd.n3975 240.244
R6731 gnd.n3975 gnd.n2408 240.244
R6732 gnd.n2421 gnd.n2408 240.244
R6733 gnd.n6054 gnd.n2421 240.244
R6734 gnd.n6054 gnd.n2422 240.244
R6735 gnd.n6050 gnd.n2422 240.244
R6736 gnd.n6050 gnd.n2428 240.244
R6737 gnd.n6042 gnd.n2428 240.244
R6738 gnd.n6042 gnd.n2443 240.244
R6739 gnd.n6038 gnd.n2443 240.244
R6740 gnd.n6038 gnd.n2449 240.244
R6741 gnd.n6030 gnd.n2449 240.244
R6742 gnd.n6030 gnd.n2465 240.244
R6743 gnd.n6026 gnd.n2465 240.244
R6744 gnd.n6026 gnd.n2471 240.244
R6745 gnd.n6018 gnd.n2471 240.244
R6746 gnd.n6018 gnd.n2486 240.244
R6747 gnd.n6014 gnd.n2486 240.244
R6748 gnd.n6014 gnd.n2492 240.244
R6749 gnd.n6006 gnd.n2492 240.244
R6750 gnd.n6006 gnd.n2508 240.244
R6751 gnd.n6002 gnd.n2508 240.244
R6752 gnd.n6002 gnd.n2514 240.244
R6753 gnd.n5994 gnd.n2514 240.244
R6754 gnd.n5994 gnd.n2527 240.244
R6755 gnd.n5990 gnd.n2527 240.244
R6756 gnd.n5990 gnd.n2533 240.244
R6757 gnd.n5981 gnd.n2533 240.244
R6758 gnd.n5981 gnd.n2546 240.244
R6759 gnd.n5977 gnd.n2546 240.244
R6760 gnd.n5977 gnd.n2552 240.244
R6761 gnd.n5969 gnd.n2552 240.244
R6762 gnd.n5969 gnd.n2566 240.244
R6763 gnd.n5965 gnd.n2566 240.244
R6764 gnd.n5965 gnd.n2572 240.244
R6765 gnd.n5957 gnd.n2572 240.244
R6766 gnd.n5957 gnd.n2588 240.244
R6767 gnd.n5953 gnd.n2588 240.244
R6768 gnd.n5953 gnd.n2594 240.244
R6769 gnd.n5945 gnd.n2594 240.244
R6770 gnd.n5945 gnd.n2609 240.244
R6771 gnd.n5941 gnd.n2609 240.244
R6772 gnd.n5941 gnd.n2615 240.244
R6773 gnd.n5933 gnd.n2615 240.244
R6774 gnd.n5933 gnd.n2631 240.244
R6775 gnd.n5929 gnd.n2631 240.244
R6776 gnd.n5929 gnd.n2637 240.244
R6777 gnd.n5921 gnd.n2637 240.244
R6778 gnd.n5921 gnd.n2653 240.244
R6779 gnd.n5917 gnd.n2653 240.244
R6780 gnd.n5917 gnd.n2659 240.244
R6781 gnd.n5909 gnd.n2659 240.244
R6782 gnd.n6425 gnd.n798 240.244
R6783 gnd.n6425 gnd.n794 240.244
R6784 gnd.n6431 gnd.n794 240.244
R6785 gnd.n6431 gnd.n792 240.244
R6786 gnd.n6435 gnd.n792 240.244
R6787 gnd.n6435 gnd.n788 240.244
R6788 gnd.n6441 gnd.n788 240.244
R6789 gnd.n6441 gnd.n786 240.244
R6790 gnd.n6445 gnd.n786 240.244
R6791 gnd.n6445 gnd.n782 240.244
R6792 gnd.n6451 gnd.n782 240.244
R6793 gnd.n6451 gnd.n780 240.244
R6794 gnd.n6455 gnd.n780 240.244
R6795 gnd.n6455 gnd.n776 240.244
R6796 gnd.n6461 gnd.n776 240.244
R6797 gnd.n6461 gnd.n774 240.244
R6798 gnd.n6465 gnd.n774 240.244
R6799 gnd.n6465 gnd.n770 240.244
R6800 gnd.n6471 gnd.n770 240.244
R6801 gnd.n6471 gnd.n768 240.244
R6802 gnd.n6475 gnd.n768 240.244
R6803 gnd.n6475 gnd.n764 240.244
R6804 gnd.n6481 gnd.n764 240.244
R6805 gnd.n6481 gnd.n762 240.244
R6806 gnd.n6485 gnd.n762 240.244
R6807 gnd.n6485 gnd.n758 240.244
R6808 gnd.n6491 gnd.n758 240.244
R6809 gnd.n6491 gnd.n756 240.244
R6810 gnd.n6495 gnd.n756 240.244
R6811 gnd.n6495 gnd.n752 240.244
R6812 gnd.n6501 gnd.n752 240.244
R6813 gnd.n6501 gnd.n750 240.244
R6814 gnd.n6505 gnd.n750 240.244
R6815 gnd.n6505 gnd.n746 240.244
R6816 gnd.n6511 gnd.n746 240.244
R6817 gnd.n6511 gnd.n744 240.244
R6818 gnd.n6515 gnd.n744 240.244
R6819 gnd.n6515 gnd.n740 240.244
R6820 gnd.n6521 gnd.n740 240.244
R6821 gnd.n6521 gnd.n738 240.244
R6822 gnd.n6525 gnd.n738 240.244
R6823 gnd.n6525 gnd.n734 240.244
R6824 gnd.n6531 gnd.n734 240.244
R6825 gnd.n6531 gnd.n732 240.244
R6826 gnd.n6535 gnd.n732 240.244
R6827 gnd.n6535 gnd.n728 240.244
R6828 gnd.n6541 gnd.n728 240.244
R6829 gnd.n6541 gnd.n726 240.244
R6830 gnd.n6545 gnd.n726 240.244
R6831 gnd.n6545 gnd.n722 240.244
R6832 gnd.n6551 gnd.n722 240.244
R6833 gnd.n6551 gnd.n720 240.244
R6834 gnd.n6555 gnd.n720 240.244
R6835 gnd.n6555 gnd.n716 240.244
R6836 gnd.n6561 gnd.n716 240.244
R6837 gnd.n6561 gnd.n714 240.244
R6838 gnd.n6565 gnd.n714 240.244
R6839 gnd.n6565 gnd.n710 240.244
R6840 gnd.n6571 gnd.n710 240.244
R6841 gnd.n6571 gnd.n708 240.244
R6842 gnd.n6575 gnd.n708 240.244
R6843 gnd.n6575 gnd.n704 240.244
R6844 gnd.n6581 gnd.n704 240.244
R6845 gnd.n6581 gnd.n702 240.244
R6846 gnd.n6585 gnd.n702 240.244
R6847 gnd.n6585 gnd.n698 240.244
R6848 gnd.n6591 gnd.n698 240.244
R6849 gnd.n6591 gnd.n696 240.244
R6850 gnd.n6595 gnd.n696 240.244
R6851 gnd.n6595 gnd.n692 240.244
R6852 gnd.n6601 gnd.n692 240.244
R6853 gnd.n6601 gnd.n690 240.244
R6854 gnd.n6605 gnd.n690 240.244
R6855 gnd.n6605 gnd.n686 240.244
R6856 gnd.n6611 gnd.n686 240.244
R6857 gnd.n6611 gnd.n684 240.244
R6858 gnd.n6615 gnd.n684 240.244
R6859 gnd.n6615 gnd.n680 240.244
R6860 gnd.n6621 gnd.n680 240.244
R6861 gnd.n6621 gnd.n678 240.244
R6862 gnd.n6625 gnd.n678 240.244
R6863 gnd.n6625 gnd.n674 240.244
R6864 gnd.n6631 gnd.n674 240.244
R6865 gnd.n6631 gnd.n672 240.244
R6866 gnd.n6635 gnd.n672 240.244
R6867 gnd.n6635 gnd.n668 240.244
R6868 gnd.n6641 gnd.n668 240.244
R6869 gnd.n6641 gnd.n666 240.244
R6870 gnd.n6645 gnd.n666 240.244
R6871 gnd.n6645 gnd.n662 240.244
R6872 gnd.n6651 gnd.n662 240.244
R6873 gnd.n6651 gnd.n660 240.244
R6874 gnd.n6655 gnd.n660 240.244
R6875 gnd.n6655 gnd.n656 240.244
R6876 gnd.n6661 gnd.n656 240.244
R6877 gnd.n6661 gnd.n654 240.244
R6878 gnd.n6665 gnd.n654 240.244
R6879 gnd.n6665 gnd.n650 240.244
R6880 gnd.n6671 gnd.n650 240.244
R6881 gnd.n6671 gnd.n648 240.244
R6882 gnd.n6675 gnd.n648 240.244
R6883 gnd.n6675 gnd.n644 240.244
R6884 gnd.n6681 gnd.n644 240.244
R6885 gnd.n6681 gnd.n642 240.244
R6886 gnd.n6685 gnd.n642 240.244
R6887 gnd.n6685 gnd.n638 240.244
R6888 gnd.n6691 gnd.n638 240.244
R6889 gnd.n6691 gnd.n636 240.244
R6890 gnd.n6695 gnd.n636 240.244
R6891 gnd.n6695 gnd.n632 240.244
R6892 gnd.n6701 gnd.n632 240.244
R6893 gnd.n6701 gnd.n630 240.244
R6894 gnd.n6705 gnd.n630 240.244
R6895 gnd.n6705 gnd.n626 240.244
R6896 gnd.n6711 gnd.n626 240.244
R6897 gnd.n6711 gnd.n624 240.244
R6898 gnd.n6715 gnd.n624 240.244
R6899 gnd.n6715 gnd.n620 240.244
R6900 gnd.n6721 gnd.n620 240.244
R6901 gnd.n6721 gnd.n618 240.244
R6902 gnd.n6725 gnd.n618 240.244
R6903 gnd.n6725 gnd.n614 240.244
R6904 gnd.n6731 gnd.n614 240.244
R6905 gnd.n6731 gnd.n612 240.244
R6906 gnd.n6735 gnd.n612 240.244
R6907 gnd.n6735 gnd.n608 240.244
R6908 gnd.n6741 gnd.n608 240.244
R6909 gnd.n6741 gnd.n606 240.244
R6910 gnd.n6745 gnd.n606 240.244
R6911 gnd.n6745 gnd.n602 240.244
R6912 gnd.n6751 gnd.n602 240.244
R6913 gnd.n6751 gnd.n600 240.244
R6914 gnd.n6755 gnd.n600 240.244
R6915 gnd.n6755 gnd.n596 240.244
R6916 gnd.n6761 gnd.n596 240.244
R6917 gnd.n6761 gnd.n594 240.244
R6918 gnd.n6765 gnd.n594 240.244
R6919 gnd.n6765 gnd.n590 240.244
R6920 gnd.n6771 gnd.n590 240.244
R6921 gnd.n6771 gnd.n588 240.244
R6922 gnd.n6775 gnd.n588 240.244
R6923 gnd.n6775 gnd.n584 240.244
R6924 gnd.n6781 gnd.n584 240.244
R6925 gnd.n6781 gnd.n582 240.244
R6926 gnd.n6785 gnd.n582 240.244
R6927 gnd.n6785 gnd.n578 240.244
R6928 gnd.n6791 gnd.n578 240.244
R6929 gnd.n6791 gnd.n576 240.244
R6930 gnd.n6795 gnd.n576 240.244
R6931 gnd.n6795 gnd.n572 240.244
R6932 gnd.n6801 gnd.n572 240.244
R6933 gnd.n6801 gnd.n570 240.244
R6934 gnd.n6805 gnd.n570 240.244
R6935 gnd.n6805 gnd.n566 240.244
R6936 gnd.n6811 gnd.n566 240.244
R6937 gnd.n6811 gnd.n564 240.244
R6938 gnd.n6815 gnd.n564 240.244
R6939 gnd.n6815 gnd.n560 240.244
R6940 gnd.n6821 gnd.n560 240.244
R6941 gnd.n6821 gnd.n558 240.244
R6942 gnd.n6825 gnd.n558 240.244
R6943 gnd.n6825 gnd.n554 240.244
R6944 gnd.n6831 gnd.n554 240.244
R6945 gnd.n6831 gnd.n552 240.244
R6946 gnd.n6835 gnd.n552 240.244
R6947 gnd.n6835 gnd.n548 240.244
R6948 gnd.n6841 gnd.n548 240.244
R6949 gnd.n6841 gnd.n546 240.244
R6950 gnd.n6845 gnd.n546 240.244
R6951 gnd.n6845 gnd.n542 240.244
R6952 gnd.n6851 gnd.n542 240.244
R6953 gnd.n6851 gnd.n540 240.244
R6954 gnd.n6855 gnd.n540 240.244
R6955 gnd.n6855 gnd.n536 240.244
R6956 gnd.n6861 gnd.n536 240.244
R6957 gnd.n6861 gnd.n534 240.244
R6958 gnd.n6865 gnd.n534 240.244
R6959 gnd.n6865 gnd.n530 240.244
R6960 gnd.n6871 gnd.n530 240.244
R6961 gnd.n6871 gnd.n528 240.244
R6962 gnd.n6875 gnd.n528 240.244
R6963 gnd.n6875 gnd.n524 240.244
R6964 gnd.n6881 gnd.n524 240.244
R6965 gnd.n6881 gnd.n522 240.244
R6966 gnd.n6885 gnd.n522 240.244
R6967 gnd.n6885 gnd.n518 240.244
R6968 gnd.n6891 gnd.n518 240.244
R6969 gnd.n6891 gnd.n516 240.244
R6970 gnd.n6895 gnd.n516 240.244
R6971 gnd.n6895 gnd.n512 240.244
R6972 gnd.n6902 gnd.n512 240.244
R6973 gnd.n6902 gnd.n510 240.244
R6974 gnd.n6906 gnd.n510 240.244
R6975 gnd.n6906 gnd.n507 240.244
R6976 gnd.n6912 gnd.n505 240.244
R6977 gnd.n6916 gnd.n505 240.244
R6978 gnd.n6916 gnd.n501 240.244
R6979 gnd.n6922 gnd.n501 240.244
R6980 gnd.n6922 gnd.n499 240.244
R6981 gnd.n6926 gnd.n499 240.244
R6982 gnd.n6926 gnd.n495 240.244
R6983 gnd.n6932 gnd.n495 240.244
R6984 gnd.n6932 gnd.n493 240.244
R6985 gnd.n6936 gnd.n493 240.244
R6986 gnd.n6936 gnd.n489 240.244
R6987 gnd.n6942 gnd.n489 240.244
R6988 gnd.n6942 gnd.n487 240.244
R6989 gnd.n6946 gnd.n487 240.244
R6990 gnd.n6946 gnd.n483 240.244
R6991 gnd.n6952 gnd.n483 240.244
R6992 gnd.n6952 gnd.n481 240.244
R6993 gnd.n6956 gnd.n481 240.244
R6994 gnd.n6956 gnd.n477 240.244
R6995 gnd.n6962 gnd.n477 240.244
R6996 gnd.n6962 gnd.n475 240.244
R6997 gnd.n6966 gnd.n475 240.244
R6998 gnd.n6966 gnd.n471 240.244
R6999 gnd.n6972 gnd.n471 240.244
R7000 gnd.n6972 gnd.n469 240.244
R7001 gnd.n6976 gnd.n469 240.244
R7002 gnd.n6976 gnd.n465 240.244
R7003 gnd.n6982 gnd.n465 240.244
R7004 gnd.n6982 gnd.n463 240.244
R7005 gnd.n6986 gnd.n463 240.244
R7006 gnd.n6986 gnd.n459 240.244
R7007 gnd.n6992 gnd.n459 240.244
R7008 gnd.n6992 gnd.n457 240.244
R7009 gnd.n6996 gnd.n457 240.244
R7010 gnd.n6996 gnd.n453 240.244
R7011 gnd.n7002 gnd.n453 240.244
R7012 gnd.n7002 gnd.n451 240.244
R7013 gnd.n7006 gnd.n451 240.244
R7014 gnd.n7006 gnd.n447 240.244
R7015 gnd.n7012 gnd.n447 240.244
R7016 gnd.n7012 gnd.n445 240.244
R7017 gnd.n7016 gnd.n445 240.244
R7018 gnd.n7016 gnd.n441 240.244
R7019 gnd.n7022 gnd.n441 240.244
R7020 gnd.n7022 gnd.n439 240.244
R7021 gnd.n7026 gnd.n439 240.244
R7022 gnd.n7026 gnd.n435 240.244
R7023 gnd.n7032 gnd.n435 240.244
R7024 gnd.n7032 gnd.n433 240.244
R7025 gnd.n7036 gnd.n433 240.244
R7026 gnd.n7036 gnd.n429 240.244
R7027 gnd.n7042 gnd.n429 240.244
R7028 gnd.n7042 gnd.n427 240.244
R7029 gnd.n7046 gnd.n427 240.244
R7030 gnd.n7046 gnd.n423 240.244
R7031 gnd.n7052 gnd.n423 240.244
R7032 gnd.n7052 gnd.n421 240.244
R7033 gnd.n7056 gnd.n421 240.244
R7034 gnd.n7056 gnd.n417 240.244
R7035 gnd.n7062 gnd.n417 240.244
R7036 gnd.n7062 gnd.n415 240.244
R7037 gnd.n7066 gnd.n415 240.244
R7038 gnd.n7066 gnd.n411 240.244
R7039 gnd.n7072 gnd.n411 240.244
R7040 gnd.n7072 gnd.n409 240.244
R7041 gnd.n7076 gnd.n409 240.244
R7042 gnd.n7076 gnd.n405 240.244
R7043 gnd.n7082 gnd.n405 240.244
R7044 gnd.n7082 gnd.n403 240.244
R7045 gnd.n7086 gnd.n403 240.244
R7046 gnd.n7086 gnd.n399 240.244
R7047 gnd.n7092 gnd.n399 240.244
R7048 gnd.n7092 gnd.n397 240.244
R7049 gnd.n7096 gnd.n397 240.244
R7050 gnd.n7096 gnd.n393 240.244
R7051 gnd.n7102 gnd.n393 240.244
R7052 gnd.n7102 gnd.n391 240.244
R7053 gnd.n7106 gnd.n391 240.244
R7054 gnd.n7106 gnd.n387 240.244
R7055 gnd.n7112 gnd.n387 240.244
R7056 gnd.n7112 gnd.n385 240.244
R7057 gnd.n7117 gnd.n385 240.244
R7058 gnd.n7117 gnd.n381 240.244
R7059 gnd.n7124 gnd.n381 240.244
R7060 gnd.n3966 gnd.n3811 240.244
R7061 gnd.n3966 gnd.n3965 240.244
R7062 gnd.n3965 gnd.n3964 240.244
R7063 gnd.n3964 gnd.n3815 240.244
R7064 gnd.n3960 gnd.n3815 240.244
R7065 gnd.n3960 gnd.n3959 240.244
R7066 gnd.n3959 gnd.n3958 240.244
R7067 gnd.n3958 gnd.n3821 240.244
R7068 gnd.n3954 gnd.n3821 240.244
R7069 gnd.n3954 gnd.n3953 240.244
R7070 gnd.n3953 gnd.n3952 240.244
R7071 gnd.n3952 gnd.n3827 240.244
R7072 gnd.n3948 gnd.n3827 240.244
R7073 gnd.n3948 gnd.n3947 240.244
R7074 gnd.n3947 gnd.n3946 240.244
R7075 gnd.n3946 gnd.n3833 240.244
R7076 gnd.n3942 gnd.n3833 240.244
R7077 gnd.n3942 gnd.n3941 240.244
R7078 gnd.n3941 gnd.n3940 240.244
R7079 gnd.n3940 gnd.n3839 240.244
R7080 gnd.n3846 gnd.n3839 240.244
R7081 gnd.n3933 gnd.n3846 240.244
R7082 gnd.n3933 gnd.n3932 240.244
R7083 gnd.n3932 gnd.n3931 240.244
R7084 gnd.n3931 gnd.n3929 240.244
R7085 gnd.n3929 gnd.n3926 240.244
R7086 gnd.n3926 gnd.n3925 240.244
R7087 gnd.n3925 gnd.n3847 240.244
R7088 gnd.n3921 gnd.n3847 240.244
R7089 gnd.n3921 gnd.n3920 240.244
R7090 gnd.n3920 gnd.n3919 240.244
R7091 gnd.n3919 gnd.n3850 240.244
R7092 gnd.n3915 gnd.n3850 240.244
R7093 gnd.n3915 gnd.n3914 240.244
R7094 gnd.n3914 gnd.n3913 240.244
R7095 gnd.n3913 gnd.n3856 240.244
R7096 gnd.n3909 gnd.n3856 240.244
R7097 gnd.n3909 gnd.n3908 240.244
R7098 gnd.n3908 gnd.n3907 240.244
R7099 gnd.n3907 gnd.n3862 240.244
R7100 gnd.n3903 gnd.n3862 240.244
R7101 gnd.n3903 gnd.n3902 240.244
R7102 gnd.n3902 gnd.n3901 240.244
R7103 gnd.n3901 gnd.n3868 240.244
R7104 gnd.n3897 gnd.n3868 240.244
R7105 gnd.n3897 gnd.n3896 240.244
R7106 gnd.n3896 gnd.n3895 240.244
R7107 gnd.n3895 gnd.n3874 240.244
R7108 gnd.n3891 gnd.n3874 240.244
R7109 gnd.n3891 gnd.n3890 240.244
R7110 gnd.n3890 gnd.n3889 240.244
R7111 gnd.n3889 gnd.n3880 240.244
R7112 gnd.n3885 gnd.n3880 240.244
R7113 gnd.n3885 gnd.n3526 240.244
R7114 gnd.n4626 gnd.n3526 240.244
R7115 gnd.n4626 gnd.n3522 240.244
R7116 gnd.n4632 gnd.n3522 240.244
R7117 gnd.n4632 gnd.n3513 240.244
R7118 gnd.n4642 gnd.n3513 240.244
R7119 gnd.n4642 gnd.n3509 240.244
R7120 gnd.n4648 gnd.n3509 240.244
R7121 gnd.n4648 gnd.n3500 240.244
R7122 gnd.n4658 gnd.n3500 240.244
R7123 gnd.n4658 gnd.n3496 240.244
R7124 gnd.n4664 gnd.n3496 240.244
R7125 gnd.n4664 gnd.n3486 240.244
R7126 gnd.n4674 gnd.n3486 240.244
R7127 gnd.n4674 gnd.n3482 240.244
R7128 gnd.n4680 gnd.n3482 240.244
R7129 gnd.n4680 gnd.n3472 240.244
R7130 gnd.n4690 gnd.n3472 240.244
R7131 gnd.n4690 gnd.n3468 240.244
R7132 gnd.n4696 gnd.n3468 240.244
R7133 gnd.n4696 gnd.n3459 240.244
R7134 gnd.n4706 gnd.n3459 240.244
R7135 gnd.n4706 gnd.n3454 240.244
R7136 gnd.n4714 gnd.n3454 240.244
R7137 gnd.n4714 gnd.n3455 240.244
R7138 gnd.n3455 gnd.n3430 240.244
R7139 gnd.n4839 gnd.n3430 240.244
R7140 gnd.n4839 gnd.n3426 240.244
R7141 gnd.n4845 gnd.n3426 240.244
R7142 gnd.n4845 gnd.n3418 240.244
R7143 gnd.n4855 gnd.n3418 240.244
R7144 gnd.n4855 gnd.n3414 240.244
R7145 gnd.n4861 gnd.n3414 240.244
R7146 gnd.n4861 gnd.n3405 240.244
R7147 gnd.n4871 gnd.n3405 240.244
R7148 gnd.n4871 gnd.n3401 240.244
R7149 gnd.n4877 gnd.n3401 240.244
R7150 gnd.n4877 gnd.n3393 240.244
R7151 gnd.n4887 gnd.n3393 240.244
R7152 gnd.n4887 gnd.n3388 240.244
R7153 gnd.n4895 gnd.n3388 240.244
R7154 gnd.n4895 gnd.n3389 240.244
R7155 gnd.n3389 gnd.n3364 240.244
R7156 gnd.n5016 gnd.n3364 240.244
R7157 gnd.n5016 gnd.n3360 240.244
R7158 gnd.n5022 gnd.n3360 240.244
R7159 gnd.n5022 gnd.n3351 240.244
R7160 gnd.n5032 gnd.n3351 240.244
R7161 gnd.n5032 gnd.n3347 240.244
R7162 gnd.n5038 gnd.n3347 240.244
R7163 gnd.n5038 gnd.n3336 240.244
R7164 gnd.n5048 gnd.n3336 240.244
R7165 gnd.n5048 gnd.n3332 240.244
R7166 gnd.n5054 gnd.n3332 240.244
R7167 gnd.n5054 gnd.n3322 240.244
R7168 gnd.n5064 gnd.n3322 240.244
R7169 gnd.n5064 gnd.n3317 240.244
R7170 gnd.n5072 gnd.n3317 240.244
R7171 gnd.n5072 gnd.n3318 240.244
R7172 gnd.n3318 gnd.n3292 240.244
R7173 gnd.n5350 gnd.n3292 240.244
R7174 gnd.n5350 gnd.n3288 240.244
R7175 gnd.n5356 gnd.n3288 240.244
R7176 gnd.n5356 gnd.n3280 240.244
R7177 gnd.n5366 gnd.n3280 240.244
R7178 gnd.n5366 gnd.n3276 240.244
R7179 gnd.n5372 gnd.n3276 240.244
R7180 gnd.n5372 gnd.n3267 240.244
R7181 gnd.n5382 gnd.n3267 240.244
R7182 gnd.n5382 gnd.n3263 240.244
R7183 gnd.n5388 gnd.n3263 240.244
R7184 gnd.n5388 gnd.n3254 240.244
R7185 gnd.n5398 gnd.n3254 240.244
R7186 gnd.n5398 gnd.n3250 240.244
R7187 gnd.n5404 gnd.n3250 240.244
R7188 gnd.n5404 gnd.n3241 240.244
R7189 gnd.n5414 gnd.n3241 240.244
R7190 gnd.n5414 gnd.n3237 240.244
R7191 gnd.n5420 gnd.n3237 240.244
R7192 gnd.n5420 gnd.n3229 240.244
R7193 gnd.n5432 gnd.n3229 240.244
R7194 gnd.n5432 gnd.n3224 240.244
R7195 gnd.n5441 gnd.n3224 240.244
R7196 gnd.n5441 gnd.n3225 240.244
R7197 gnd.n3225 gnd.n2783 240.244
R7198 gnd.n5777 gnd.n2783 240.244
R7199 gnd.n5777 gnd.n2786 240.244
R7200 gnd.n5773 gnd.n2786 240.244
R7201 gnd.n5773 gnd.n2792 240.244
R7202 gnd.n3028 gnd.n2792 240.244
R7203 gnd.n3034 gnd.n3028 240.244
R7204 gnd.n3035 gnd.n3034 240.244
R7205 gnd.n5481 gnd.n3035 240.244
R7206 gnd.n5481 gnd.n3023 240.244
R7207 gnd.n5489 gnd.n3023 240.244
R7208 gnd.n5489 gnd.n3024 240.244
R7209 gnd.n3024 gnd.n3000 240.244
R7210 gnd.n5512 gnd.n3000 240.244
R7211 gnd.n5512 gnd.n2995 240.244
R7212 gnd.n5520 gnd.n2995 240.244
R7213 gnd.n5520 gnd.n2996 240.244
R7214 gnd.n2996 gnd.n2972 240.244
R7215 gnd.n5543 gnd.n2972 240.244
R7216 gnd.n5543 gnd.n2966 240.244
R7217 gnd.n5558 gnd.n2966 240.244
R7218 gnd.n5558 gnd.n2968 240.244
R7219 gnd.n5554 gnd.n2968 240.244
R7220 gnd.n5554 gnd.n5553 240.244
R7221 gnd.n5553 gnd.n2914 240.244
R7222 gnd.n5649 gnd.n2914 240.244
R7223 gnd.n5649 gnd.n2916 240.244
R7224 gnd.n5645 gnd.n2916 240.244
R7225 gnd.n5645 gnd.n5644 240.244
R7226 gnd.n5644 gnd.n5643 240.244
R7227 gnd.n5643 gnd.n2923 240.244
R7228 gnd.n5638 gnd.n2923 240.244
R7229 gnd.n5638 gnd.n2925 240.244
R7230 gnd.n5630 gnd.n2925 240.244
R7231 gnd.n5630 gnd.n5622 240.244
R7232 gnd.n5625 gnd.n5622 240.244
R7233 gnd.n5625 gnd.n302 240.244
R7234 gnd.n7171 gnd.n302 240.244
R7235 gnd.n7171 gnd.n303 240.244
R7236 gnd.n7166 gnd.n303 240.244
R7237 gnd.n7166 gnd.n7165 240.244
R7238 gnd.n7165 gnd.n307 240.244
R7239 gnd.n330 gnd.n307 240.244
R7240 gnd.n331 gnd.n330 240.244
R7241 gnd.n331 gnd.n322 240.244
R7242 gnd.n7150 gnd.n322 240.244
R7243 gnd.n7150 gnd.n323 240.244
R7244 gnd.n7146 gnd.n323 240.244
R7245 gnd.n7146 gnd.n7145 240.244
R7246 gnd.n7145 gnd.n339 240.244
R7247 gnd.n372 gnd.n339 240.244
R7248 gnd.n373 gnd.n372 240.244
R7249 gnd.n373 gnd.n364 240.244
R7250 gnd.n7130 gnd.n364 240.244
R7251 gnd.n7130 gnd.n365 240.244
R7252 gnd.n7126 gnd.n365 240.244
R7253 gnd.n7126 gnd.n7125 240.244
R7254 gnd.n6421 gnd.n800 240.244
R7255 gnd.n6417 gnd.n800 240.244
R7256 gnd.n6417 gnd.n805 240.244
R7257 gnd.n6413 gnd.n805 240.244
R7258 gnd.n6413 gnd.n807 240.244
R7259 gnd.n6409 gnd.n807 240.244
R7260 gnd.n6409 gnd.n813 240.244
R7261 gnd.n6405 gnd.n813 240.244
R7262 gnd.n6405 gnd.n815 240.244
R7263 gnd.n6401 gnd.n815 240.244
R7264 gnd.n6401 gnd.n821 240.244
R7265 gnd.n6397 gnd.n821 240.244
R7266 gnd.n6397 gnd.n823 240.244
R7267 gnd.n6393 gnd.n823 240.244
R7268 gnd.n6393 gnd.n829 240.244
R7269 gnd.n6389 gnd.n829 240.244
R7270 gnd.n6389 gnd.n831 240.244
R7271 gnd.n6385 gnd.n831 240.244
R7272 gnd.n6385 gnd.n837 240.244
R7273 gnd.n6381 gnd.n837 240.244
R7274 gnd.n6381 gnd.n839 240.244
R7275 gnd.n6377 gnd.n839 240.244
R7276 gnd.n6377 gnd.n845 240.244
R7277 gnd.n6373 gnd.n845 240.244
R7278 gnd.n6373 gnd.n847 240.244
R7279 gnd.n6369 gnd.n847 240.244
R7280 gnd.n6369 gnd.n853 240.244
R7281 gnd.n6365 gnd.n853 240.244
R7282 gnd.n6365 gnd.n855 240.244
R7283 gnd.n6361 gnd.n855 240.244
R7284 gnd.n6361 gnd.n861 240.244
R7285 gnd.n6357 gnd.n861 240.244
R7286 gnd.n6357 gnd.n863 240.244
R7287 gnd.n6353 gnd.n863 240.244
R7288 gnd.n6353 gnd.n869 240.244
R7289 gnd.n6349 gnd.n869 240.244
R7290 gnd.n6349 gnd.n871 240.244
R7291 gnd.n6345 gnd.n871 240.244
R7292 gnd.n6345 gnd.n877 240.244
R7293 gnd.n6341 gnd.n877 240.244
R7294 gnd.n6341 gnd.n879 240.244
R7295 gnd.n6337 gnd.n879 240.244
R7296 gnd.n6337 gnd.n885 240.244
R7297 gnd.n6333 gnd.n885 240.244
R7298 gnd.n6333 gnd.n887 240.244
R7299 gnd.n6329 gnd.n887 240.244
R7300 gnd.n6329 gnd.n893 240.244
R7301 gnd.n6325 gnd.n893 240.244
R7302 gnd.n6325 gnd.n895 240.244
R7303 gnd.n6321 gnd.n895 240.244
R7304 gnd.n6321 gnd.n901 240.244
R7305 gnd.n6317 gnd.n901 240.244
R7306 gnd.n6317 gnd.n903 240.244
R7307 gnd.n6313 gnd.n903 240.244
R7308 gnd.n6313 gnd.n909 240.244
R7309 gnd.n6309 gnd.n909 240.244
R7310 gnd.n6309 gnd.n911 240.244
R7311 gnd.n6305 gnd.n911 240.244
R7312 gnd.n6305 gnd.n917 240.244
R7313 gnd.n6301 gnd.n917 240.244
R7314 gnd.n6301 gnd.n919 240.244
R7315 gnd.n6297 gnd.n919 240.244
R7316 gnd.n6297 gnd.n925 240.244
R7317 gnd.n6293 gnd.n925 240.244
R7318 gnd.n6293 gnd.n927 240.244
R7319 gnd.n6289 gnd.n927 240.244
R7320 gnd.n6289 gnd.n933 240.244
R7321 gnd.n6285 gnd.n933 240.244
R7322 gnd.n6285 gnd.n935 240.244
R7323 gnd.n6281 gnd.n935 240.244
R7324 gnd.n6281 gnd.n941 240.244
R7325 gnd.n6277 gnd.n941 240.244
R7326 gnd.n6277 gnd.n943 240.244
R7327 gnd.n6273 gnd.n943 240.244
R7328 gnd.n6273 gnd.n949 240.244
R7329 gnd.n6269 gnd.n949 240.244
R7330 gnd.n6269 gnd.n951 240.244
R7331 gnd.n6265 gnd.n951 240.244
R7332 gnd.n6265 gnd.n957 240.244
R7333 gnd.n6261 gnd.n957 240.244
R7334 gnd.n6261 gnd.n959 240.244
R7335 gnd.n6257 gnd.n959 240.244
R7336 gnd.n6257 gnd.n965 240.244
R7337 gnd.n3972 gnd.n965 240.244
R7338 gnd.n2679 gnd.n2678 240.244
R7339 gnd.n2680 gnd.n2679 240.244
R7340 gnd.n3515 gnd.n2680 240.244
R7341 gnd.n3515 gnd.n2683 240.244
R7342 gnd.n2684 gnd.n2683 240.244
R7343 gnd.n2685 gnd.n2684 240.244
R7344 gnd.n3501 gnd.n2685 240.244
R7345 gnd.n3501 gnd.n2688 240.244
R7346 gnd.n2689 gnd.n2688 240.244
R7347 gnd.n2690 gnd.n2689 240.244
R7348 gnd.n3487 gnd.n2690 240.244
R7349 gnd.n3487 gnd.n2693 240.244
R7350 gnd.n2694 gnd.n2693 240.244
R7351 gnd.n2695 gnd.n2694 240.244
R7352 gnd.n3474 gnd.n2695 240.244
R7353 gnd.n3474 gnd.n2698 240.244
R7354 gnd.n2699 gnd.n2698 240.244
R7355 gnd.n2700 gnd.n2699 240.244
R7356 gnd.n3460 gnd.n2700 240.244
R7357 gnd.n3460 gnd.n2703 240.244
R7358 gnd.n2704 gnd.n2703 240.244
R7359 gnd.n2705 gnd.n2704 240.244
R7360 gnd.n3446 gnd.n2705 240.244
R7361 gnd.n3446 gnd.n2708 240.244
R7362 gnd.n2709 gnd.n2708 240.244
R7363 gnd.n2710 gnd.n2709 240.244
R7364 gnd.n4734 gnd.n2710 240.244
R7365 gnd.n4734 gnd.n2713 240.244
R7366 gnd.n2714 gnd.n2713 240.244
R7367 gnd.n2715 gnd.n2714 240.244
R7368 gnd.n4809 gnd.n2715 240.244
R7369 gnd.n4809 gnd.n2718 240.244
R7370 gnd.n2719 gnd.n2718 240.244
R7371 gnd.n2720 gnd.n2719 240.244
R7372 gnd.n4760 gnd.n2720 240.244
R7373 gnd.n4760 gnd.n2723 240.244
R7374 gnd.n2724 gnd.n2723 240.244
R7375 gnd.n2725 gnd.n2724 240.244
R7376 gnd.n4777 gnd.n2725 240.244
R7377 gnd.n4777 gnd.n2728 240.244
R7378 gnd.n2729 gnd.n2728 240.244
R7379 gnd.n2730 gnd.n2729 240.244
R7380 gnd.n3358 gnd.n2730 240.244
R7381 gnd.n3358 gnd.n2733 240.244
R7382 gnd.n2734 gnd.n2733 240.244
R7383 gnd.n2735 gnd.n2734 240.244
R7384 gnd.n3345 gnd.n2735 240.244
R7385 gnd.n3345 gnd.n2738 240.244
R7386 gnd.n2739 gnd.n2738 240.244
R7387 gnd.n2740 gnd.n2739 240.244
R7388 gnd.n3330 gnd.n2740 240.244
R7389 gnd.n3330 gnd.n2743 240.244
R7390 gnd.n2744 gnd.n2743 240.244
R7391 gnd.n2745 gnd.n2744 240.244
R7392 gnd.n3315 gnd.n2745 240.244
R7393 gnd.n3315 gnd.n2748 240.244
R7394 gnd.n2749 gnd.n2748 240.244
R7395 gnd.n2750 gnd.n2749 240.244
R7396 gnd.n3301 gnd.n2750 240.244
R7397 gnd.n3301 gnd.n2753 240.244
R7398 gnd.n2754 gnd.n2753 240.244
R7399 gnd.n2755 gnd.n2754 240.244
R7400 gnd.n5095 gnd.n2755 240.244
R7401 gnd.n5095 gnd.n2758 240.244
R7402 gnd.n2759 gnd.n2758 240.244
R7403 gnd.n2760 gnd.n2759 240.244
R7404 gnd.n5107 gnd.n2760 240.244
R7405 gnd.n5107 gnd.n2763 240.244
R7406 gnd.n2764 gnd.n2763 240.244
R7407 gnd.n2765 gnd.n2764 240.244
R7408 gnd.n3255 gnd.n2765 240.244
R7409 gnd.n3255 gnd.n2768 240.244
R7410 gnd.n2769 gnd.n2768 240.244
R7411 gnd.n2770 gnd.n2769 240.244
R7412 gnd.n3243 gnd.n2770 240.244
R7413 gnd.n3243 gnd.n2773 240.244
R7414 gnd.n2774 gnd.n2773 240.244
R7415 gnd.n2775 gnd.n2774 240.244
R7416 gnd.n3222 gnd.n2775 240.244
R7417 gnd.n3222 gnd.n2778 240.244
R7418 gnd.n2779 gnd.n2778 240.244
R7419 gnd.n5780 gnd.n2779 240.244
R7420 gnd.n3611 gnd.n3610 240.244
R7421 gnd.n3595 gnd.n3594 240.244
R7422 gnd.n3623 gnd.n3622 240.244
R7423 gnd.n3635 gnd.n3634 240.244
R7424 gnd.n3583 gnd.n3582 240.244
R7425 gnd.n3647 gnd.n3646 240.244
R7426 gnd.n3658 gnd.n3657 240.244
R7427 gnd.n3558 gnd.n3557 240.244
R7428 gnd.n4599 gnd.n4598 240.244
R7429 gnd.n3553 gnd.n3552 240.244
R7430 gnd.n4608 gnd.n4607 240.244
R7431 gnd.n3549 gnd.n3548 240.244
R7432 gnd.n4617 gnd.n4616 240.244
R7433 gnd.n4623 gnd.n3542 240.244
R7434 gnd.n4634 gnd.n3520 240.244
R7435 gnd.n4634 gnd.n3516 240.244
R7436 gnd.n4640 gnd.n3516 240.244
R7437 gnd.n4640 gnd.n3506 240.244
R7438 gnd.n4650 gnd.n3506 240.244
R7439 gnd.n4650 gnd.n3502 240.244
R7440 gnd.n4656 gnd.n3502 240.244
R7441 gnd.n4656 gnd.n3493 240.244
R7442 gnd.n4666 gnd.n3493 240.244
R7443 gnd.n4666 gnd.n3489 240.244
R7444 gnd.n4672 gnd.n3489 240.244
R7445 gnd.n4672 gnd.n3480 240.244
R7446 gnd.n4682 gnd.n3480 240.244
R7447 gnd.n4682 gnd.n3476 240.244
R7448 gnd.n4688 gnd.n3476 240.244
R7449 gnd.n4688 gnd.n3466 240.244
R7450 gnd.n4698 gnd.n3466 240.244
R7451 gnd.n4698 gnd.n3462 240.244
R7452 gnd.n4704 gnd.n3462 240.244
R7453 gnd.n4704 gnd.n3452 240.244
R7454 gnd.n4716 gnd.n3452 240.244
R7455 gnd.n4716 gnd.n3447 240.244
R7456 gnd.n4723 gnd.n3447 240.244
R7457 gnd.n4723 gnd.n3433 240.244
R7458 gnd.n3433 gnd.n3424 240.244
R7459 gnd.n4847 gnd.n3424 240.244
R7460 gnd.n4847 gnd.n3420 240.244
R7461 gnd.n4853 gnd.n3420 240.244
R7462 gnd.n4853 gnd.n3412 240.244
R7463 gnd.n4863 gnd.n3412 240.244
R7464 gnd.n4863 gnd.n3408 240.244
R7465 gnd.n4869 gnd.n3408 240.244
R7466 gnd.n4869 gnd.n3399 240.244
R7467 gnd.n4879 gnd.n3399 240.244
R7468 gnd.n4879 gnd.n3395 240.244
R7469 gnd.n4885 gnd.n3395 240.244
R7470 gnd.n4885 gnd.n3385 240.244
R7471 gnd.n4897 gnd.n3385 240.244
R7472 gnd.n4897 gnd.n3380 240.244
R7473 gnd.n4904 gnd.n3380 240.244
R7474 gnd.n4904 gnd.n3368 240.244
R7475 gnd.n3368 gnd.n3357 240.244
R7476 gnd.n5024 gnd.n3357 240.244
R7477 gnd.n5024 gnd.n3353 240.244
R7478 gnd.n5030 gnd.n3353 240.244
R7479 gnd.n5030 gnd.n3343 240.244
R7480 gnd.n5040 gnd.n3343 240.244
R7481 gnd.n5040 gnd.n3339 240.244
R7482 gnd.n5046 gnd.n3339 240.244
R7483 gnd.n5046 gnd.n3328 240.244
R7484 gnd.n5056 gnd.n3328 240.244
R7485 gnd.n5056 gnd.n3324 240.244
R7486 gnd.n5062 gnd.n3324 240.244
R7487 gnd.n5062 gnd.n3313 240.244
R7488 gnd.n5074 gnd.n3313 240.244
R7489 gnd.n5074 gnd.n3308 240.244
R7490 gnd.n5081 gnd.n3308 240.244
R7491 gnd.n5081 gnd.n3295 240.244
R7492 gnd.n3295 gnd.n3286 240.244
R7493 gnd.n5358 gnd.n3286 240.244
R7494 gnd.n5358 gnd.n3282 240.244
R7495 gnd.n5364 gnd.n3282 240.244
R7496 gnd.n5364 gnd.n3273 240.244
R7497 gnd.n5374 gnd.n3273 240.244
R7498 gnd.n5374 gnd.n3269 240.244
R7499 gnd.n5380 gnd.n3269 240.244
R7500 gnd.n5380 gnd.n3261 240.244
R7501 gnd.n5390 gnd.n3261 240.244
R7502 gnd.n5390 gnd.n3257 240.244
R7503 gnd.n5396 gnd.n3257 240.244
R7504 gnd.n5396 gnd.n3249 240.244
R7505 gnd.n5406 gnd.n3249 240.244
R7506 gnd.n5406 gnd.n3245 240.244
R7507 gnd.n5412 gnd.n3245 240.244
R7508 gnd.n5412 gnd.n3236 240.244
R7509 gnd.n5422 gnd.n3236 240.244
R7510 gnd.n5422 gnd.n3231 240.244
R7511 gnd.n5430 gnd.n3231 240.244
R7512 gnd.n5430 gnd.n3221 240.244
R7513 gnd.n5443 gnd.n3221 240.244
R7514 gnd.n5444 gnd.n5443 240.244
R7515 gnd.n5444 gnd.n2784 240.244
R7516 gnd.n3139 gnd.n3137 240.244
R7517 gnd.n3152 gnd.n3116 240.244
R7518 gnd.n3156 gnd.n3154 240.244
R7519 gnd.n3169 gnd.n3107 240.244
R7520 gnd.n3173 gnd.n3171 240.244
R7521 gnd.n3186 gnd.n3098 240.244
R7522 gnd.n3190 gnd.n3188 240.244
R7523 gnd.n3201 gnd.n3086 240.244
R7524 gnd.n3204 gnd.n3203 240.244
R7525 gnd.n3207 gnd.n3206 240.244
R7526 gnd.n3212 gnd.n3209 240.244
R7527 gnd.n3215 gnd.n3214 240.244
R7528 gnd.n5449 gnd.n3217 240.244
R7529 gnd.n5452 gnd.n5451 240.244
R7530 gnd.n4336 gnd.n4335 240.132
R7531 gnd.n5125 gnd.n5124 240.132
R7532 gnd.n6914 gnd.n6913 235.673
R7533 gnd.n6915 gnd.n6914 235.673
R7534 gnd.n6915 gnd.n500 235.673
R7535 gnd.n6923 gnd.n500 235.673
R7536 gnd.n6924 gnd.n6923 235.673
R7537 gnd.n6925 gnd.n6924 235.673
R7538 gnd.n6925 gnd.n494 235.673
R7539 gnd.n6933 gnd.n494 235.673
R7540 gnd.n6934 gnd.n6933 235.673
R7541 gnd.n6935 gnd.n6934 235.673
R7542 gnd.n6935 gnd.n488 235.673
R7543 gnd.n6943 gnd.n488 235.673
R7544 gnd.n6944 gnd.n6943 235.673
R7545 gnd.n6945 gnd.n6944 235.673
R7546 gnd.n6945 gnd.n482 235.673
R7547 gnd.n6953 gnd.n482 235.673
R7548 gnd.n6954 gnd.n6953 235.673
R7549 gnd.n6955 gnd.n6954 235.673
R7550 gnd.n6955 gnd.n476 235.673
R7551 gnd.n6963 gnd.n476 235.673
R7552 gnd.n6964 gnd.n6963 235.673
R7553 gnd.n6965 gnd.n6964 235.673
R7554 gnd.n6965 gnd.n470 235.673
R7555 gnd.n6973 gnd.n470 235.673
R7556 gnd.n6974 gnd.n6973 235.673
R7557 gnd.n6975 gnd.n6974 235.673
R7558 gnd.n6975 gnd.n464 235.673
R7559 gnd.n6983 gnd.n464 235.673
R7560 gnd.n6984 gnd.n6983 235.673
R7561 gnd.n6985 gnd.n6984 235.673
R7562 gnd.n6985 gnd.n458 235.673
R7563 gnd.n6993 gnd.n458 235.673
R7564 gnd.n6994 gnd.n6993 235.673
R7565 gnd.n6995 gnd.n6994 235.673
R7566 gnd.n6995 gnd.n452 235.673
R7567 gnd.n7003 gnd.n452 235.673
R7568 gnd.n7004 gnd.n7003 235.673
R7569 gnd.n7005 gnd.n7004 235.673
R7570 gnd.n7005 gnd.n446 235.673
R7571 gnd.n7013 gnd.n446 235.673
R7572 gnd.n7014 gnd.n7013 235.673
R7573 gnd.n7015 gnd.n7014 235.673
R7574 gnd.n7015 gnd.n440 235.673
R7575 gnd.n7023 gnd.n440 235.673
R7576 gnd.n7024 gnd.n7023 235.673
R7577 gnd.n7025 gnd.n7024 235.673
R7578 gnd.n7025 gnd.n434 235.673
R7579 gnd.n7033 gnd.n434 235.673
R7580 gnd.n7034 gnd.n7033 235.673
R7581 gnd.n7035 gnd.n7034 235.673
R7582 gnd.n7035 gnd.n428 235.673
R7583 gnd.n7043 gnd.n428 235.673
R7584 gnd.n7044 gnd.n7043 235.673
R7585 gnd.n7045 gnd.n7044 235.673
R7586 gnd.n7045 gnd.n422 235.673
R7587 gnd.n7053 gnd.n422 235.673
R7588 gnd.n7054 gnd.n7053 235.673
R7589 gnd.n7055 gnd.n7054 235.673
R7590 gnd.n7055 gnd.n416 235.673
R7591 gnd.n7063 gnd.n416 235.673
R7592 gnd.n7064 gnd.n7063 235.673
R7593 gnd.n7065 gnd.n7064 235.673
R7594 gnd.n7065 gnd.n410 235.673
R7595 gnd.n7073 gnd.n410 235.673
R7596 gnd.n7074 gnd.n7073 235.673
R7597 gnd.n7075 gnd.n7074 235.673
R7598 gnd.n7075 gnd.n404 235.673
R7599 gnd.n7083 gnd.n404 235.673
R7600 gnd.n7084 gnd.n7083 235.673
R7601 gnd.n7085 gnd.n7084 235.673
R7602 gnd.n7085 gnd.n398 235.673
R7603 gnd.n7093 gnd.n398 235.673
R7604 gnd.n7094 gnd.n7093 235.673
R7605 gnd.n7095 gnd.n7094 235.673
R7606 gnd.n7095 gnd.n392 235.673
R7607 gnd.n7103 gnd.n392 235.673
R7608 gnd.n7104 gnd.n7103 235.673
R7609 gnd.n7105 gnd.n7104 235.673
R7610 gnd.n7105 gnd.n386 235.673
R7611 gnd.n7113 gnd.n386 235.673
R7612 gnd.n7114 gnd.n7113 235.673
R7613 gnd.n7116 gnd.n7114 235.673
R7614 gnd.n7116 gnd.n7115 235.673
R7615 gnd.n6424 gnd.n6423 225.874
R7616 gnd.n6424 gnd.n793 225.874
R7617 gnd.n6432 gnd.n793 225.874
R7618 gnd.n6433 gnd.n6432 225.874
R7619 gnd.n6434 gnd.n6433 225.874
R7620 gnd.n6434 gnd.n787 225.874
R7621 gnd.n6442 gnd.n787 225.874
R7622 gnd.n6443 gnd.n6442 225.874
R7623 gnd.n6444 gnd.n6443 225.874
R7624 gnd.n6444 gnd.n781 225.874
R7625 gnd.n6452 gnd.n781 225.874
R7626 gnd.n6453 gnd.n6452 225.874
R7627 gnd.n6454 gnd.n6453 225.874
R7628 gnd.n6454 gnd.n775 225.874
R7629 gnd.n6462 gnd.n775 225.874
R7630 gnd.n6463 gnd.n6462 225.874
R7631 gnd.n6464 gnd.n6463 225.874
R7632 gnd.n6464 gnd.n769 225.874
R7633 gnd.n6472 gnd.n769 225.874
R7634 gnd.n6473 gnd.n6472 225.874
R7635 gnd.n6474 gnd.n6473 225.874
R7636 gnd.n6474 gnd.n763 225.874
R7637 gnd.n6482 gnd.n763 225.874
R7638 gnd.n6483 gnd.n6482 225.874
R7639 gnd.n6484 gnd.n6483 225.874
R7640 gnd.n6484 gnd.n757 225.874
R7641 gnd.n6492 gnd.n757 225.874
R7642 gnd.n6493 gnd.n6492 225.874
R7643 gnd.n6494 gnd.n6493 225.874
R7644 gnd.n6494 gnd.n751 225.874
R7645 gnd.n6502 gnd.n751 225.874
R7646 gnd.n6503 gnd.n6502 225.874
R7647 gnd.n6504 gnd.n6503 225.874
R7648 gnd.n6504 gnd.n745 225.874
R7649 gnd.n6512 gnd.n745 225.874
R7650 gnd.n6513 gnd.n6512 225.874
R7651 gnd.n6514 gnd.n6513 225.874
R7652 gnd.n6514 gnd.n739 225.874
R7653 gnd.n6522 gnd.n739 225.874
R7654 gnd.n6523 gnd.n6522 225.874
R7655 gnd.n6524 gnd.n6523 225.874
R7656 gnd.n6524 gnd.n733 225.874
R7657 gnd.n6532 gnd.n733 225.874
R7658 gnd.n6533 gnd.n6532 225.874
R7659 gnd.n6534 gnd.n6533 225.874
R7660 gnd.n6534 gnd.n727 225.874
R7661 gnd.n6542 gnd.n727 225.874
R7662 gnd.n6543 gnd.n6542 225.874
R7663 gnd.n6544 gnd.n6543 225.874
R7664 gnd.n6544 gnd.n721 225.874
R7665 gnd.n6552 gnd.n721 225.874
R7666 gnd.n6553 gnd.n6552 225.874
R7667 gnd.n6554 gnd.n6553 225.874
R7668 gnd.n6554 gnd.n715 225.874
R7669 gnd.n6562 gnd.n715 225.874
R7670 gnd.n6563 gnd.n6562 225.874
R7671 gnd.n6564 gnd.n6563 225.874
R7672 gnd.n6564 gnd.n709 225.874
R7673 gnd.n6572 gnd.n709 225.874
R7674 gnd.n6573 gnd.n6572 225.874
R7675 gnd.n6574 gnd.n6573 225.874
R7676 gnd.n6574 gnd.n703 225.874
R7677 gnd.n6582 gnd.n703 225.874
R7678 gnd.n6583 gnd.n6582 225.874
R7679 gnd.n6584 gnd.n6583 225.874
R7680 gnd.n6584 gnd.n697 225.874
R7681 gnd.n6592 gnd.n697 225.874
R7682 gnd.n6593 gnd.n6592 225.874
R7683 gnd.n6594 gnd.n6593 225.874
R7684 gnd.n6594 gnd.n691 225.874
R7685 gnd.n6602 gnd.n691 225.874
R7686 gnd.n6603 gnd.n6602 225.874
R7687 gnd.n6604 gnd.n6603 225.874
R7688 gnd.n6604 gnd.n685 225.874
R7689 gnd.n6612 gnd.n685 225.874
R7690 gnd.n6613 gnd.n6612 225.874
R7691 gnd.n6614 gnd.n6613 225.874
R7692 gnd.n6614 gnd.n679 225.874
R7693 gnd.n6622 gnd.n679 225.874
R7694 gnd.n6623 gnd.n6622 225.874
R7695 gnd.n6624 gnd.n6623 225.874
R7696 gnd.n6624 gnd.n673 225.874
R7697 gnd.n6632 gnd.n673 225.874
R7698 gnd.n6633 gnd.n6632 225.874
R7699 gnd.n6634 gnd.n6633 225.874
R7700 gnd.n6634 gnd.n667 225.874
R7701 gnd.n6642 gnd.n667 225.874
R7702 gnd.n6643 gnd.n6642 225.874
R7703 gnd.n6644 gnd.n6643 225.874
R7704 gnd.n6644 gnd.n661 225.874
R7705 gnd.n6652 gnd.n661 225.874
R7706 gnd.n6653 gnd.n6652 225.874
R7707 gnd.n6654 gnd.n6653 225.874
R7708 gnd.n6654 gnd.n655 225.874
R7709 gnd.n6662 gnd.n655 225.874
R7710 gnd.n6663 gnd.n6662 225.874
R7711 gnd.n6664 gnd.n6663 225.874
R7712 gnd.n6664 gnd.n649 225.874
R7713 gnd.n6672 gnd.n649 225.874
R7714 gnd.n6673 gnd.n6672 225.874
R7715 gnd.n6674 gnd.n6673 225.874
R7716 gnd.n6674 gnd.n643 225.874
R7717 gnd.n6682 gnd.n643 225.874
R7718 gnd.n6683 gnd.n6682 225.874
R7719 gnd.n6684 gnd.n6683 225.874
R7720 gnd.n6684 gnd.n637 225.874
R7721 gnd.n6692 gnd.n637 225.874
R7722 gnd.n6693 gnd.n6692 225.874
R7723 gnd.n6694 gnd.n6693 225.874
R7724 gnd.n6694 gnd.n631 225.874
R7725 gnd.n6702 gnd.n631 225.874
R7726 gnd.n6703 gnd.n6702 225.874
R7727 gnd.n6704 gnd.n6703 225.874
R7728 gnd.n6704 gnd.n625 225.874
R7729 gnd.n6712 gnd.n625 225.874
R7730 gnd.n6713 gnd.n6712 225.874
R7731 gnd.n6714 gnd.n6713 225.874
R7732 gnd.n6714 gnd.n619 225.874
R7733 gnd.n6722 gnd.n619 225.874
R7734 gnd.n6723 gnd.n6722 225.874
R7735 gnd.n6724 gnd.n6723 225.874
R7736 gnd.n6724 gnd.n613 225.874
R7737 gnd.n6732 gnd.n613 225.874
R7738 gnd.n6733 gnd.n6732 225.874
R7739 gnd.n6734 gnd.n6733 225.874
R7740 gnd.n6734 gnd.n607 225.874
R7741 gnd.n6742 gnd.n607 225.874
R7742 gnd.n6743 gnd.n6742 225.874
R7743 gnd.n6744 gnd.n6743 225.874
R7744 gnd.n6744 gnd.n601 225.874
R7745 gnd.n6752 gnd.n601 225.874
R7746 gnd.n6753 gnd.n6752 225.874
R7747 gnd.n6754 gnd.n6753 225.874
R7748 gnd.n6754 gnd.n595 225.874
R7749 gnd.n6762 gnd.n595 225.874
R7750 gnd.n6763 gnd.n6762 225.874
R7751 gnd.n6764 gnd.n6763 225.874
R7752 gnd.n6764 gnd.n589 225.874
R7753 gnd.n6772 gnd.n589 225.874
R7754 gnd.n6773 gnd.n6772 225.874
R7755 gnd.n6774 gnd.n6773 225.874
R7756 gnd.n6774 gnd.n583 225.874
R7757 gnd.n6782 gnd.n583 225.874
R7758 gnd.n6783 gnd.n6782 225.874
R7759 gnd.n6784 gnd.n6783 225.874
R7760 gnd.n6784 gnd.n577 225.874
R7761 gnd.n6792 gnd.n577 225.874
R7762 gnd.n6793 gnd.n6792 225.874
R7763 gnd.n6794 gnd.n6793 225.874
R7764 gnd.n6794 gnd.n571 225.874
R7765 gnd.n6802 gnd.n571 225.874
R7766 gnd.n6803 gnd.n6802 225.874
R7767 gnd.n6804 gnd.n6803 225.874
R7768 gnd.n6804 gnd.n565 225.874
R7769 gnd.n6812 gnd.n565 225.874
R7770 gnd.n6813 gnd.n6812 225.874
R7771 gnd.n6814 gnd.n6813 225.874
R7772 gnd.n6814 gnd.n559 225.874
R7773 gnd.n6822 gnd.n559 225.874
R7774 gnd.n6823 gnd.n6822 225.874
R7775 gnd.n6824 gnd.n6823 225.874
R7776 gnd.n6824 gnd.n553 225.874
R7777 gnd.n6832 gnd.n553 225.874
R7778 gnd.n6833 gnd.n6832 225.874
R7779 gnd.n6834 gnd.n6833 225.874
R7780 gnd.n6834 gnd.n547 225.874
R7781 gnd.n6842 gnd.n547 225.874
R7782 gnd.n6843 gnd.n6842 225.874
R7783 gnd.n6844 gnd.n6843 225.874
R7784 gnd.n6844 gnd.n541 225.874
R7785 gnd.n6852 gnd.n541 225.874
R7786 gnd.n6853 gnd.n6852 225.874
R7787 gnd.n6854 gnd.n6853 225.874
R7788 gnd.n6854 gnd.n535 225.874
R7789 gnd.n6862 gnd.n535 225.874
R7790 gnd.n6863 gnd.n6862 225.874
R7791 gnd.n6864 gnd.n6863 225.874
R7792 gnd.n6864 gnd.n529 225.874
R7793 gnd.n6872 gnd.n529 225.874
R7794 gnd.n6873 gnd.n6872 225.874
R7795 gnd.n6874 gnd.n6873 225.874
R7796 gnd.n6874 gnd.n523 225.874
R7797 gnd.n6882 gnd.n523 225.874
R7798 gnd.n6883 gnd.n6882 225.874
R7799 gnd.n6884 gnd.n6883 225.874
R7800 gnd.n6884 gnd.n517 225.874
R7801 gnd.n6892 gnd.n517 225.874
R7802 gnd.n6893 gnd.n6892 225.874
R7803 gnd.n6894 gnd.n6893 225.874
R7804 gnd.n6894 gnd.n511 225.874
R7805 gnd.n6903 gnd.n511 225.874
R7806 gnd.n6904 gnd.n6903 225.874
R7807 gnd.n6905 gnd.n6904 225.874
R7808 gnd.n6905 gnd.n506 225.874
R7809 gnd.n1557 gnd.t109 224.174
R7810 gnd.n1072 gnd.t151 224.174
R7811 gnd.n2842 gnd.n2799 199.319
R7812 gnd.n2842 gnd.n2800 199.319
R7813 gnd.n3708 gnd.n3678 199.319
R7814 gnd.n3708 gnd.n3677 199.319
R7815 gnd.n4337 gnd.n4334 186.49
R7816 gnd.n5126 gnd.n5123 186.49
R7817 gnd.n2292 gnd.n2291 185
R7818 gnd.n2290 gnd.n2289 185
R7819 gnd.n2269 gnd.n2268 185
R7820 gnd.n2284 gnd.n2283 185
R7821 gnd.n2282 gnd.n2281 185
R7822 gnd.n2273 gnd.n2272 185
R7823 gnd.n2276 gnd.n2275 185
R7824 gnd.n2260 gnd.n2259 185
R7825 gnd.n2258 gnd.n2257 185
R7826 gnd.n2237 gnd.n2236 185
R7827 gnd.n2252 gnd.n2251 185
R7828 gnd.n2250 gnd.n2249 185
R7829 gnd.n2241 gnd.n2240 185
R7830 gnd.n2244 gnd.n2243 185
R7831 gnd.n2228 gnd.n2227 185
R7832 gnd.n2226 gnd.n2225 185
R7833 gnd.n2205 gnd.n2204 185
R7834 gnd.n2220 gnd.n2219 185
R7835 gnd.n2218 gnd.n2217 185
R7836 gnd.n2209 gnd.n2208 185
R7837 gnd.n2212 gnd.n2211 185
R7838 gnd.n2197 gnd.n2196 185
R7839 gnd.n2195 gnd.n2194 185
R7840 gnd.n2174 gnd.n2173 185
R7841 gnd.n2189 gnd.n2188 185
R7842 gnd.n2187 gnd.n2186 185
R7843 gnd.n2178 gnd.n2177 185
R7844 gnd.n2181 gnd.n2180 185
R7845 gnd.n2165 gnd.n2164 185
R7846 gnd.n2163 gnd.n2162 185
R7847 gnd.n2142 gnd.n2141 185
R7848 gnd.n2157 gnd.n2156 185
R7849 gnd.n2155 gnd.n2154 185
R7850 gnd.n2146 gnd.n2145 185
R7851 gnd.n2149 gnd.n2148 185
R7852 gnd.n2133 gnd.n2132 185
R7853 gnd.n2131 gnd.n2130 185
R7854 gnd.n2110 gnd.n2109 185
R7855 gnd.n2125 gnd.n2124 185
R7856 gnd.n2123 gnd.n2122 185
R7857 gnd.n2114 gnd.n2113 185
R7858 gnd.n2117 gnd.n2116 185
R7859 gnd.n2101 gnd.n2100 185
R7860 gnd.n2099 gnd.n2098 185
R7861 gnd.n2078 gnd.n2077 185
R7862 gnd.n2093 gnd.n2092 185
R7863 gnd.n2091 gnd.n2090 185
R7864 gnd.n2082 gnd.n2081 185
R7865 gnd.n2085 gnd.n2084 185
R7866 gnd.n2070 gnd.n2069 185
R7867 gnd.n2068 gnd.n2067 185
R7868 gnd.n2047 gnd.n2046 185
R7869 gnd.n2062 gnd.n2061 185
R7870 gnd.n2060 gnd.n2059 185
R7871 gnd.n2051 gnd.n2050 185
R7872 gnd.n2054 gnd.n2053 185
R7873 gnd.n1558 gnd.t108 178.987
R7874 gnd.n1073 gnd.t152 178.987
R7875 gnd.n1 gnd.t74 170.774
R7876 gnd.n7 gnd.t17 170.103
R7877 gnd.n6 gnd.t65 170.103
R7878 gnd.n5 gnd.t61 170.103
R7879 gnd.n4 gnd.t72 170.103
R7880 gnd.n3 gnd.t63 170.103
R7881 gnd.n2 gnd.t5 170.103
R7882 gnd.n1 gnd.t12 170.103
R7883 gnd.n5306 gnd.n5137 163.367
R7884 gnd.n5302 gnd.n5301 163.367
R7885 gnd.n5299 gnd.n5140 163.367
R7886 gnd.n5295 gnd.n5294 163.367
R7887 gnd.n5292 gnd.n5143 163.367
R7888 gnd.n5288 gnd.n5287 163.367
R7889 gnd.n5285 gnd.n5146 163.367
R7890 gnd.n5281 gnd.n5280 163.367
R7891 gnd.n5278 gnd.n5149 163.367
R7892 gnd.n5274 gnd.n5273 163.367
R7893 gnd.n5271 gnd.n5152 163.367
R7894 gnd.n5267 gnd.n5266 163.367
R7895 gnd.n5264 gnd.n5155 163.367
R7896 gnd.n5260 gnd.n5259 163.367
R7897 gnd.n5257 gnd.n5158 163.367
R7898 gnd.n5253 gnd.n5252 163.367
R7899 gnd.n5249 gnd.n5248 163.367
R7900 gnd.n5246 gnd.n5164 163.367
R7901 gnd.n5241 gnd.n5240 163.367
R7902 gnd.n5238 gnd.n5169 163.367
R7903 gnd.n5234 gnd.n5233 163.367
R7904 gnd.n5231 gnd.n5172 163.367
R7905 gnd.n5227 gnd.n5226 163.367
R7906 gnd.n5224 gnd.n5175 163.367
R7907 gnd.n5220 gnd.n5219 163.367
R7908 gnd.n5217 gnd.n5178 163.367
R7909 gnd.n5213 gnd.n5212 163.367
R7910 gnd.n5210 gnd.n5181 163.367
R7911 gnd.n5206 gnd.n5205 163.367
R7912 gnd.n5203 gnd.n5184 163.367
R7913 gnd.n5199 gnd.n5198 163.367
R7914 gnd.n5196 gnd.n5187 163.367
R7915 gnd.n4492 gnd.n4326 163.367
R7916 gnd.n4437 gnd.n4326 163.367
R7917 gnd.n4437 gnd.n4434 163.367
R7918 gnd.n4481 gnd.n4434 163.367
R7919 gnd.n4481 gnd.n4435 163.367
R7920 gnd.n4477 gnd.n4435 163.367
R7921 gnd.n4477 gnd.n4441 163.367
R7922 gnd.n4456 gnd.n4441 163.367
R7923 gnd.n4456 gnd.n4454 163.367
R7924 gnd.n4466 gnd.n4454 163.367
R7925 gnd.n4466 gnd.n4455 163.367
R7926 gnd.n4462 gnd.n4455 163.367
R7927 gnd.n4462 gnd.n3445 163.367
R7928 gnd.n3445 gnd.n3434 163.367
R7929 gnd.n4837 gnd.n3434 163.367
R7930 gnd.n4837 gnd.n3435 163.367
R7931 gnd.n4833 gnd.n3435 163.367
R7932 gnd.n4833 gnd.n3438 163.367
R7933 gnd.n4733 gnd.n3438 163.367
R7934 gnd.n4823 gnd.n4733 163.367
R7935 gnd.n4823 gnd.n4735 163.367
R7936 gnd.n4819 gnd.n4735 163.367
R7937 gnd.n4819 gnd.n4738 163.367
R7938 gnd.n4746 gnd.n4738 163.367
R7939 gnd.n4808 gnd.n4746 163.367
R7940 gnd.n4808 gnd.n4747 163.367
R7941 gnd.n4804 gnd.n4747 163.367
R7942 gnd.n4804 gnd.n4803 163.367
R7943 gnd.n4803 gnd.n4750 163.367
R7944 gnd.n4758 gnd.n4750 163.367
R7945 gnd.n4759 gnd.n4758 163.367
R7946 gnd.n4761 gnd.n4759 163.367
R7947 gnd.n4768 gnd.n4761 163.367
R7948 gnd.n4785 gnd.n4768 163.367
R7949 gnd.n4785 gnd.n4769 163.367
R7950 gnd.n4781 gnd.n4769 163.367
R7951 gnd.n4781 gnd.n4780 163.367
R7952 gnd.n4780 gnd.n3379 163.367
R7953 gnd.n3379 gnd.n3369 163.367
R7954 gnd.n5014 gnd.n3369 163.367
R7955 gnd.n5014 gnd.n3370 163.367
R7956 gnd.n5010 gnd.n3370 163.367
R7957 gnd.n5010 gnd.n3373 163.367
R7958 gnd.n4914 gnd.n3373 163.367
R7959 gnd.n5000 gnd.n4914 163.367
R7960 gnd.n5000 gnd.n4915 163.367
R7961 gnd.n4996 gnd.n4915 163.367
R7962 gnd.n4996 gnd.n4918 163.367
R7963 gnd.n4925 gnd.n4918 163.367
R7964 gnd.n4986 gnd.n4925 163.367
R7965 gnd.n4986 gnd.n4926 163.367
R7966 gnd.n4982 gnd.n4926 163.367
R7967 gnd.n4982 gnd.n4981 163.367
R7968 gnd.n4981 gnd.n4929 163.367
R7969 gnd.n4940 gnd.n4929 163.367
R7970 gnd.n4940 gnd.n4937 163.367
R7971 gnd.n4970 gnd.n4937 163.367
R7972 gnd.n4970 gnd.n4938 163.367
R7973 gnd.n4966 gnd.n4938 163.367
R7974 gnd.n4966 gnd.n4944 163.367
R7975 gnd.n4951 gnd.n4944 163.367
R7976 gnd.n4956 gnd.n4951 163.367
R7977 gnd.n4956 gnd.n4952 163.367
R7978 gnd.n4952 gnd.n3296 163.367
R7979 gnd.n5348 gnd.n3296 163.367
R7980 gnd.n5348 gnd.n3297 163.367
R7981 gnd.n5344 gnd.n3297 163.367
R7982 gnd.n5344 gnd.n3300 163.367
R7983 gnd.n5090 gnd.n3300 163.367
R7984 gnd.n5334 gnd.n5090 163.367
R7985 gnd.n5334 gnd.n5091 163.367
R7986 gnd.n5330 gnd.n5091 163.367
R7987 gnd.n5330 gnd.n5094 163.367
R7988 gnd.n5102 gnd.n5094 163.367
R7989 gnd.n5320 gnd.n5102 163.367
R7990 gnd.n5320 gnd.n5103 163.367
R7991 gnd.n5316 gnd.n5103 163.367
R7992 gnd.n5316 gnd.n5315 163.367
R7993 gnd.n5315 gnd.n5106 163.367
R7994 gnd.n5191 gnd.n5106 163.367
R7995 gnd.n4428 gnd.n4426 163.367
R7996 gnd.n4426 gnd.n4425 163.367
R7997 gnd.n4422 gnd.n4421 163.367
R7998 gnd.n4419 gnd.n4353 163.367
R7999 gnd.n4415 gnd.n4413 163.367
R8000 gnd.n4411 gnd.n4355 163.367
R8001 gnd.n4407 gnd.n4405 163.367
R8002 gnd.n4403 gnd.n4357 163.367
R8003 gnd.n4399 gnd.n4397 163.367
R8004 gnd.n4395 gnd.n4359 163.367
R8005 gnd.n4391 gnd.n4389 163.367
R8006 gnd.n4387 gnd.n4361 163.367
R8007 gnd.n4383 gnd.n4381 163.367
R8008 gnd.n4379 gnd.n4363 163.367
R8009 gnd.n4375 gnd.n4373 163.367
R8010 gnd.n4370 gnd.n4369 163.367
R8011 gnd.n4559 gnd.n4557 163.367
R8012 gnd.n4555 gnd.n4308 163.367
R8013 gnd.n4550 gnd.n4548 163.367
R8014 gnd.n4546 gnd.n4312 163.367
R8015 gnd.n4542 gnd.n4540 163.367
R8016 gnd.n4538 gnd.n4314 163.367
R8017 gnd.n4534 gnd.n4532 163.367
R8018 gnd.n4530 gnd.n4316 163.367
R8019 gnd.n4526 gnd.n4524 163.367
R8020 gnd.n4522 gnd.n4318 163.367
R8021 gnd.n4518 gnd.n4516 163.367
R8022 gnd.n4514 gnd.n4320 163.367
R8023 gnd.n4510 gnd.n4508 163.367
R8024 gnd.n4506 gnd.n4322 163.367
R8025 gnd.n4502 gnd.n4500 163.367
R8026 gnd.n4498 gnd.n4324 163.367
R8027 gnd.n4490 gnd.n4329 163.367
R8028 gnd.n4486 gnd.n4329 163.367
R8029 gnd.n4486 gnd.n4485 163.367
R8030 gnd.n4485 gnd.n4433 163.367
R8031 gnd.n4443 gnd.n4433 163.367
R8032 gnd.n4475 gnd.n4443 163.367
R8033 gnd.n4475 gnd.n4445 163.367
R8034 gnd.n4471 gnd.n4445 163.367
R8035 gnd.n4471 gnd.n4470 163.367
R8036 gnd.n4470 gnd.n4453 163.367
R8037 gnd.n4453 gnd.n4449 163.367
R8038 gnd.n4449 gnd.n3444 163.367
R8039 gnd.n4726 gnd.n3444 163.367
R8040 gnd.n4727 gnd.n4726 163.367
R8041 gnd.n4727 gnd.n3432 163.367
R8042 gnd.n3441 gnd.n3432 163.367
R8043 gnd.n4831 gnd.n3441 163.367
R8044 gnd.n4831 gnd.n3442 163.367
R8045 gnd.n4827 gnd.n3442 163.367
R8046 gnd.n4827 gnd.n4732 163.367
R8047 gnd.n4740 gnd.n4732 163.367
R8048 gnd.n4817 gnd.n4740 163.367
R8049 gnd.n4817 gnd.n4742 163.367
R8050 gnd.n4813 gnd.n4742 163.367
R8051 gnd.n4813 gnd.n4812 163.367
R8052 gnd.n4812 gnd.n4745 163.367
R8053 gnd.n4752 gnd.n4745 163.367
R8054 gnd.n4801 gnd.n4752 163.367
R8055 gnd.n4801 gnd.n4753 163.367
R8056 gnd.n4797 gnd.n4753 163.367
R8057 gnd.n4797 gnd.n4757 163.367
R8058 gnd.n4792 gnd.n4757 163.367
R8059 gnd.n4792 gnd.n4762 163.367
R8060 gnd.n4788 gnd.n4762 163.367
R8061 gnd.n4788 gnd.n4767 163.367
R8062 gnd.n4767 gnd.n4766 163.367
R8063 gnd.n4766 gnd.n3378 163.367
R8064 gnd.n4907 gnd.n3378 163.367
R8065 gnd.n4908 gnd.n4907 163.367
R8066 gnd.n4908 gnd.n3366 163.367
R8067 gnd.n3375 gnd.n3366 163.367
R8068 gnd.n5008 gnd.n3375 163.367
R8069 gnd.n5008 gnd.n3376 163.367
R8070 gnd.n5004 gnd.n3376 163.367
R8071 gnd.n5004 gnd.n4913 163.367
R8072 gnd.n4920 gnd.n4913 163.367
R8073 gnd.n4994 gnd.n4920 163.367
R8074 gnd.n4994 gnd.n4921 163.367
R8075 gnd.n4990 gnd.n4921 163.367
R8076 gnd.n4990 gnd.n4989 163.367
R8077 gnd.n4989 gnd.n4924 163.367
R8078 gnd.n4931 gnd.n4924 163.367
R8079 gnd.n4979 gnd.n4931 163.367
R8080 gnd.n4979 gnd.n4932 163.367
R8081 gnd.n4975 gnd.n4932 163.367
R8082 gnd.n4975 gnd.n4974 163.367
R8083 gnd.n4974 gnd.n4936 163.367
R8084 gnd.n4946 gnd.n4936 163.367
R8085 gnd.n4964 gnd.n4946 163.367
R8086 gnd.n4964 gnd.n4947 163.367
R8087 gnd.n4960 gnd.n4947 163.367
R8088 gnd.n4960 gnd.n4959 163.367
R8089 gnd.n4959 gnd.n3306 163.367
R8090 gnd.n5084 gnd.n3306 163.367
R8091 gnd.n5084 gnd.n3293 163.367
R8092 gnd.n3303 gnd.n3293 163.367
R8093 gnd.n5342 gnd.n3303 163.367
R8094 gnd.n5342 gnd.n3304 163.367
R8095 gnd.n5338 gnd.n3304 163.367
R8096 gnd.n5338 gnd.n5089 163.367
R8097 gnd.n5097 gnd.n5089 163.367
R8098 gnd.n5328 gnd.n5097 163.367
R8099 gnd.n5328 gnd.n5098 163.367
R8100 gnd.n5324 gnd.n5098 163.367
R8101 gnd.n5324 gnd.n5323 163.367
R8102 gnd.n5323 gnd.n5101 163.367
R8103 gnd.n5109 gnd.n5101 163.367
R8104 gnd.n5313 gnd.n5109 163.367
R8105 gnd.n5313 gnd.n5111 163.367
R8106 gnd.n5309 gnd.n5111 163.367
R8107 gnd.n5132 gnd.n5131 156.462
R8108 gnd.n2232 gnd.n2200 153.042
R8109 gnd.n2296 gnd.n2295 152.079
R8110 gnd.n2264 gnd.n2263 152.079
R8111 gnd.n2232 gnd.n2231 152.079
R8112 gnd.n4342 gnd.n4341 152
R8113 gnd.n4343 gnd.n4332 152
R8114 gnd.n4345 gnd.n4344 152
R8115 gnd.n4347 gnd.n4330 152
R8116 gnd.n4349 gnd.n4348 152
R8117 gnd.n5130 gnd.n5114 152
R8118 gnd.n5122 gnd.n5115 152
R8119 gnd.n5121 gnd.n5120 152
R8120 gnd.n5119 gnd.n5116 152
R8121 gnd.n5117 gnd.t122 150.546
R8122 gnd.t37 gnd.n2274 147.661
R8123 gnd.t70 gnd.n2242 147.661
R8124 gnd.t40 gnd.n2210 147.661
R8125 gnd.t316 gnd.n2179 147.661
R8126 gnd.t320 gnd.n2147 147.661
R8127 gnd.t23 gnd.n2115 147.661
R8128 gnd.t318 gnd.n2083 147.661
R8129 gnd.t29 gnd.n2052 147.661
R8130 gnd.n5251 gnd.n5250 143.351
R8131 gnd.n4368 gnd.n4307 143.351
R8132 gnd.n4558 gnd.n4307 143.351
R8133 gnd.n4339 gnd.t162 130.484
R8134 gnd.n4348 gnd.t82 126.766
R8135 gnd.n4346 gnd.t159 126.766
R8136 gnd.n4332 gnd.t171 126.766
R8137 gnd.n4340 gnd.t129 126.766
R8138 gnd.n5118 gnd.t168 126.766
R8139 gnd.n5120 gnd.t142 126.766
R8140 gnd.n5129 gnd.t75 126.766
R8141 gnd.n5131 gnd.t153 126.766
R8142 gnd.n5738 gnd.n2841 112.192
R8143 gnd.n4561 gnd.n4560 112.192
R8144 gnd.n2291 gnd.n2290 104.615
R8145 gnd.n2290 gnd.n2268 104.615
R8146 gnd.n2283 gnd.n2268 104.615
R8147 gnd.n2283 gnd.n2282 104.615
R8148 gnd.n2282 gnd.n2272 104.615
R8149 gnd.n2275 gnd.n2272 104.615
R8150 gnd.n2259 gnd.n2258 104.615
R8151 gnd.n2258 gnd.n2236 104.615
R8152 gnd.n2251 gnd.n2236 104.615
R8153 gnd.n2251 gnd.n2250 104.615
R8154 gnd.n2250 gnd.n2240 104.615
R8155 gnd.n2243 gnd.n2240 104.615
R8156 gnd.n2227 gnd.n2226 104.615
R8157 gnd.n2226 gnd.n2204 104.615
R8158 gnd.n2219 gnd.n2204 104.615
R8159 gnd.n2219 gnd.n2218 104.615
R8160 gnd.n2218 gnd.n2208 104.615
R8161 gnd.n2211 gnd.n2208 104.615
R8162 gnd.n2196 gnd.n2195 104.615
R8163 gnd.n2195 gnd.n2173 104.615
R8164 gnd.n2188 gnd.n2173 104.615
R8165 gnd.n2188 gnd.n2187 104.615
R8166 gnd.n2187 gnd.n2177 104.615
R8167 gnd.n2180 gnd.n2177 104.615
R8168 gnd.n2164 gnd.n2163 104.615
R8169 gnd.n2163 gnd.n2141 104.615
R8170 gnd.n2156 gnd.n2141 104.615
R8171 gnd.n2156 gnd.n2155 104.615
R8172 gnd.n2155 gnd.n2145 104.615
R8173 gnd.n2148 gnd.n2145 104.615
R8174 gnd.n2132 gnd.n2131 104.615
R8175 gnd.n2131 gnd.n2109 104.615
R8176 gnd.n2124 gnd.n2109 104.615
R8177 gnd.n2124 gnd.n2123 104.615
R8178 gnd.n2123 gnd.n2113 104.615
R8179 gnd.n2116 gnd.n2113 104.615
R8180 gnd.n2100 gnd.n2099 104.615
R8181 gnd.n2099 gnd.n2077 104.615
R8182 gnd.n2092 gnd.n2077 104.615
R8183 gnd.n2092 gnd.n2091 104.615
R8184 gnd.n2091 gnd.n2081 104.615
R8185 gnd.n2084 gnd.n2081 104.615
R8186 gnd.n2069 gnd.n2068 104.615
R8187 gnd.n2068 gnd.n2046 104.615
R8188 gnd.n2061 gnd.n2046 104.615
R8189 gnd.n2061 gnd.n2060 104.615
R8190 gnd.n2060 gnd.n2050 104.615
R8191 gnd.n2053 gnd.n2050 104.615
R8192 gnd.n1483 gnd.t95 100.632
R8193 gnd.n1051 gnd.t137 100.632
R8194 gnd.n7434 gnd.n112 99.6594
R8195 gnd.n7432 gnd.n7431 99.6594
R8196 gnd.n7427 gnd.n119 99.6594
R8197 gnd.n7425 gnd.n7424 99.6594
R8198 gnd.n7420 gnd.n126 99.6594
R8199 gnd.n7418 gnd.n7417 99.6594
R8200 gnd.n7413 gnd.n133 99.6594
R8201 gnd.n7411 gnd.n7410 99.6594
R8202 gnd.n7403 gnd.n140 99.6594
R8203 gnd.n7401 gnd.n7400 99.6594
R8204 gnd.n7396 gnd.n147 99.6594
R8205 gnd.n7394 gnd.n7393 99.6594
R8206 gnd.n7389 gnd.n154 99.6594
R8207 gnd.n7387 gnd.n7386 99.6594
R8208 gnd.n7382 gnd.n161 99.6594
R8209 gnd.n7380 gnd.n7379 99.6594
R8210 gnd.n7375 gnd.n168 99.6594
R8211 gnd.n7373 gnd.n7372 99.6594
R8212 gnd.n173 gnd.n172 99.6594
R8213 gnd.n5769 gnd.n5768 99.6594
R8214 gnd.n5763 gnd.n2793 99.6594
R8215 gnd.n5760 gnd.n2794 99.6594
R8216 gnd.n5756 gnd.n2795 99.6594
R8217 gnd.n5752 gnd.n2796 99.6594
R8218 gnd.n5748 gnd.n2797 99.6594
R8219 gnd.n5744 gnd.n2798 99.6594
R8220 gnd.n5740 gnd.n2799 99.6594
R8221 gnd.n5735 gnd.n2801 99.6594
R8222 gnd.n5731 gnd.n2802 99.6594
R8223 gnd.n5727 gnd.n2803 99.6594
R8224 gnd.n5723 gnd.n2804 99.6594
R8225 gnd.n5719 gnd.n2805 99.6594
R8226 gnd.n5715 gnd.n2806 99.6594
R8227 gnd.n5711 gnd.n2807 99.6594
R8228 gnd.n5707 gnd.n2808 99.6594
R8229 gnd.n5703 gnd.n2809 99.6594
R8230 gnd.n2865 gnd.n2810 99.6594
R8231 gnd.n4589 gnd.n4588 99.6594
R8232 gnd.n4584 gnd.n3684 99.6594
R8233 gnd.n4580 gnd.n3683 99.6594
R8234 gnd.n4576 gnd.n3682 99.6594
R8235 gnd.n4572 gnd.n3681 99.6594
R8236 gnd.n4568 gnd.n3680 99.6594
R8237 gnd.n4564 gnd.n3679 99.6594
R8238 gnd.n4299 gnd.n3677 99.6594
R8239 gnd.n4297 gnd.n3676 99.6594
R8240 gnd.n4293 gnd.n3675 99.6594
R8241 gnd.n4289 gnd.n3674 99.6594
R8242 gnd.n4285 gnd.n3673 99.6594
R8243 gnd.n4281 gnd.n3672 99.6594
R8244 gnd.n4277 gnd.n3671 99.6594
R8245 gnd.n4273 gnd.n3670 99.6594
R8246 gnd.n4269 gnd.n3669 99.6594
R8247 gnd.n4265 gnd.n3668 99.6594
R8248 gnd.n3726 gnd.n3667 99.6594
R8249 gnd.n6147 gnd.n6146 99.6594
R8250 gnd.n6141 gnd.n2323 99.6594
R8251 gnd.n6138 gnd.n2324 99.6594
R8252 gnd.n6134 gnd.n2325 99.6594
R8253 gnd.n6130 gnd.n2326 99.6594
R8254 gnd.n6126 gnd.n2327 99.6594
R8255 gnd.n6122 gnd.n2328 99.6594
R8256 gnd.n6118 gnd.n2329 99.6594
R8257 gnd.n6114 gnd.n2330 99.6594
R8258 gnd.n6109 gnd.n2331 99.6594
R8259 gnd.n6105 gnd.n2332 99.6594
R8260 gnd.n6101 gnd.n2333 99.6594
R8261 gnd.n6097 gnd.n2334 99.6594
R8262 gnd.n6093 gnd.n2335 99.6594
R8263 gnd.n6089 gnd.n2336 99.6594
R8264 gnd.n6085 gnd.n2337 99.6594
R8265 gnd.n6081 gnd.n2338 99.6594
R8266 gnd.n6077 gnd.n2339 99.6594
R8267 gnd.n2394 gnd.n2340 99.6594
R8268 gnd.n6186 gnd.n6154 99.6594
R8269 gnd.n6184 gnd.n6153 99.6594
R8270 gnd.n6180 gnd.n6152 99.6594
R8271 gnd.n6176 gnd.n6151 99.6594
R8272 gnd.n6172 gnd.n6150 99.6594
R8273 gnd.n6168 gnd.n6149 99.6594
R8274 gnd.n6198 gnd.n6196 99.6594
R8275 gnd.n6204 gnd.n1050 99.6594
R8276 gnd.n1695 gnd.n1426 99.6594
R8277 gnd.n1452 gnd.n1433 99.6594
R8278 gnd.n1454 gnd.n1434 99.6594
R8279 gnd.n1462 gnd.n1435 99.6594
R8280 gnd.n1464 gnd.n1436 99.6594
R8281 gnd.n1472 gnd.n1437 99.6594
R8282 gnd.n1474 gnd.n1438 99.6594
R8283 gnd.n1482 gnd.n1439 99.6594
R8284 gnd.n1092 gnd.n1057 99.6594
R8285 gnd.n1096 gnd.n1058 99.6594
R8286 gnd.n1102 gnd.n1059 99.6594
R8287 gnd.n1106 gnd.n1060 99.6594
R8288 gnd.n1112 gnd.n1061 99.6594
R8289 gnd.n1116 gnd.n1062 99.6594
R8290 gnd.n1122 gnd.n1063 99.6594
R8291 gnd.n1126 gnd.n1064 99.6594
R8292 gnd.n1132 gnd.n1065 99.6594
R8293 gnd.n1136 gnd.n1066 99.6594
R8294 gnd.n1142 gnd.n1067 99.6594
R8295 gnd.n1145 gnd.n1068 99.6594
R8296 gnd.n2322 gnd.n2321 99.6594
R8297 gnd.n1610 gnd.n1609 99.6594
R8298 gnd.n1604 gnd.n1521 99.6594
R8299 gnd.n1601 gnd.n1522 99.6594
R8300 gnd.n1597 gnd.n1523 99.6594
R8301 gnd.n1593 gnd.n1524 99.6594
R8302 gnd.n1589 gnd.n1525 99.6594
R8303 gnd.n1585 gnd.n1526 99.6594
R8304 gnd.n1581 gnd.n1527 99.6594
R8305 gnd.n1577 gnd.n1528 99.6594
R8306 gnd.n1573 gnd.n1529 99.6594
R8307 gnd.n1569 gnd.n1530 99.6594
R8308 gnd.n1565 gnd.n1531 99.6594
R8309 gnd.n1612 gnd.n1520 99.6594
R8310 gnd.n7282 gnd.n7281 99.6594
R8311 gnd.n7287 gnd.n7286 99.6594
R8312 gnd.n7290 gnd.n7289 99.6594
R8313 gnd.n7295 gnd.n7294 99.6594
R8314 gnd.n7298 gnd.n7297 99.6594
R8315 gnd.n7303 gnd.n7302 99.6594
R8316 gnd.n7306 gnd.n7305 99.6594
R8317 gnd.n7311 gnd.n7310 99.6594
R8318 gnd.n7314 gnd.n99 99.6594
R8319 gnd.n2875 gnd.n2811 99.6594
R8320 gnd.n3131 gnd.n2812 99.6594
R8321 gnd.n3122 gnd.n2813 99.6594
R8322 gnd.n3147 gnd.n2814 99.6594
R8323 gnd.n3113 gnd.n2815 99.6594
R8324 gnd.n3164 gnd.n2816 99.6594
R8325 gnd.n3104 gnd.n2817 99.6594
R8326 gnd.n3181 gnd.n2818 99.6594
R8327 gnd.n3095 gnd.n2819 99.6594
R8328 gnd.n3605 gnd.n3565 99.6594
R8329 gnd.n3616 gnd.n3566 99.6594
R8330 gnd.n3590 gnd.n3567 99.6594
R8331 gnd.n3629 gnd.n3568 99.6594
R8332 gnd.n3640 gnd.n3569 99.6594
R8333 gnd.n3578 gnd.n3570 99.6594
R8334 gnd.n3652 gnd.n3571 99.6594
R8335 gnd.n3665 gnd.n3664 99.6594
R8336 gnd.n4592 gnd.n4591 99.6594
R8337 gnd.n4035 gnd.n2341 99.6594
R8338 gnd.n4032 gnd.n2342 99.6594
R8339 gnd.n4028 gnd.n2343 99.6594
R8340 gnd.n4024 gnd.n2344 99.6594
R8341 gnd.n4020 gnd.n2345 99.6594
R8342 gnd.n4016 gnd.n2346 99.6594
R8343 gnd.n4012 gnd.n2347 99.6594
R8344 gnd.n4008 gnd.n2348 99.6594
R8345 gnd.n4004 gnd.n2349 99.6594
R8346 gnd.n4033 gnd.n2341 99.6594
R8347 gnd.n4029 gnd.n2342 99.6594
R8348 gnd.n4025 gnd.n2343 99.6594
R8349 gnd.n4021 gnd.n2344 99.6594
R8350 gnd.n4017 gnd.n2345 99.6594
R8351 gnd.n4013 gnd.n2346 99.6594
R8352 gnd.n4009 gnd.n2347 99.6594
R8353 gnd.n4005 gnd.n2348 99.6594
R8354 gnd.n3993 gnd.n2349 99.6594
R8355 gnd.n4591 gnd.n3563 99.6594
R8356 gnd.n3665 gnd.n3572 99.6594
R8357 gnd.n3579 gnd.n3571 99.6594
R8358 gnd.n3641 gnd.n3570 99.6594
R8359 gnd.n3628 gnd.n3569 99.6594
R8360 gnd.n3591 gnd.n3568 99.6594
R8361 gnd.n3617 gnd.n3567 99.6594
R8362 gnd.n3604 gnd.n3566 99.6594
R8363 gnd.n3602 gnd.n3565 99.6594
R8364 gnd.n3130 gnd.n2811 99.6594
R8365 gnd.n3121 gnd.n2812 99.6594
R8366 gnd.n3146 gnd.n2813 99.6594
R8367 gnd.n3112 gnd.n2814 99.6594
R8368 gnd.n3163 gnd.n2815 99.6594
R8369 gnd.n3103 gnd.n2816 99.6594
R8370 gnd.n3180 gnd.n2817 99.6594
R8371 gnd.n3094 gnd.n2818 99.6594
R8372 gnd.n3090 gnd.n2819 99.6594
R8373 gnd.n7315 gnd.n7314 99.6594
R8374 gnd.n7310 gnd.n7309 99.6594
R8375 gnd.n7305 gnd.n7304 99.6594
R8376 gnd.n7302 gnd.n7301 99.6594
R8377 gnd.n7297 gnd.n7296 99.6594
R8378 gnd.n7294 gnd.n7293 99.6594
R8379 gnd.n7289 gnd.n7288 99.6594
R8380 gnd.n7286 gnd.n7285 99.6594
R8381 gnd.n7281 gnd.n7280 99.6594
R8382 gnd.n1610 gnd.n1533 99.6594
R8383 gnd.n1602 gnd.n1521 99.6594
R8384 gnd.n1598 gnd.n1522 99.6594
R8385 gnd.n1594 gnd.n1523 99.6594
R8386 gnd.n1590 gnd.n1524 99.6594
R8387 gnd.n1586 gnd.n1525 99.6594
R8388 gnd.n1582 gnd.n1526 99.6594
R8389 gnd.n1578 gnd.n1527 99.6594
R8390 gnd.n1574 gnd.n1528 99.6594
R8391 gnd.n1570 gnd.n1529 99.6594
R8392 gnd.n1566 gnd.n1530 99.6594
R8393 gnd.n1562 gnd.n1531 99.6594
R8394 gnd.n1613 gnd.n1612 99.6594
R8395 gnd.n2322 gnd.n1069 99.6594
R8396 gnd.n1143 gnd.n1068 99.6594
R8397 gnd.n1135 gnd.n1067 99.6594
R8398 gnd.n1133 gnd.n1066 99.6594
R8399 gnd.n1125 gnd.n1065 99.6594
R8400 gnd.n1123 gnd.n1064 99.6594
R8401 gnd.n1115 gnd.n1063 99.6594
R8402 gnd.n1113 gnd.n1062 99.6594
R8403 gnd.n1105 gnd.n1061 99.6594
R8404 gnd.n1103 gnd.n1060 99.6594
R8405 gnd.n1095 gnd.n1059 99.6594
R8406 gnd.n1093 gnd.n1058 99.6594
R8407 gnd.n1085 gnd.n1057 99.6594
R8408 gnd.n1696 gnd.n1695 99.6594
R8409 gnd.n1455 gnd.n1433 99.6594
R8410 gnd.n1461 gnd.n1434 99.6594
R8411 gnd.n1465 gnd.n1435 99.6594
R8412 gnd.n1471 gnd.n1436 99.6594
R8413 gnd.n1475 gnd.n1437 99.6594
R8414 gnd.n1481 gnd.n1438 99.6594
R8415 gnd.n1439 gnd.n1423 99.6594
R8416 gnd.n6197 gnd.n1050 99.6594
R8417 gnd.n6196 gnd.n1056 99.6594
R8418 gnd.n6171 gnd.n6149 99.6594
R8419 gnd.n6175 gnd.n6150 99.6594
R8420 gnd.n6179 gnd.n6151 99.6594
R8421 gnd.n6183 gnd.n6152 99.6594
R8422 gnd.n6187 gnd.n6153 99.6594
R8423 gnd.n6155 gnd.n6154 99.6594
R8424 gnd.n6147 gnd.n2353 99.6594
R8425 gnd.n6139 gnd.n2323 99.6594
R8426 gnd.n6135 gnd.n2324 99.6594
R8427 gnd.n6131 gnd.n2325 99.6594
R8428 gnd.n6127 gnd.n2326 99.6594
R8429 gnd.n6123 gnd.n2327 99.6594
R8430 gnd.n6119 gnd.n2328 99.6594
R8431 gnd.n6115 gnd.n2329 99.6594
R8432 gnd.n6110 gnd.n2330 99.6594
R8433 gnd.n6106 gnd.n2331 99.6594
R8434 gnd.n6102 gnd.n2332 99.6594
R8435 gnd.n6098 gnd.n2333 99.6594
R8436 gnd.n6094 gnd.n2334 99.6594
R8437 gnd.n6090 gnd.n2335 99.6594
R8438 gnd.n6086 gnd.n2336 99.6594
R8439 gnd.n6082 gnd.n2337 99.6594
R8440 gnd.n6078 gnd.n2338 99.6594
R8441 gnd.n2393 gnd.n2339 99.6594
R8442 gnd.n6070 gnd.n2340 99.6594
R8443 gnd.n4264 gnd.n3667 99.6594
R8444 gnd.n4268 gnd.n3668 99.6594
R8445 gnd.n4272 gnd.n3669 99.6594
R8446 gnd.n4276 gnd.n3670 99.6594
R8447 gnd.n4280 gnd.n3671 99.6594
R8448 gnd.n4284 gnd.n3672 99.6594
R8449 gnd.n4288 gnd.n3673 99.6594
R8450 gnd.n4292 gnd.n3674 99.6594
R8451 gnd.n4296 gnd.n3675 99.6594
R8452 gnd.n4300 gnd.n3676 99.6594
R8453 gnd.n4563 gnd.n3678 99.6594
R8454 gnd.n4567 gnd.n3679 99.6594
R8455 gnd.n4571 gnd.n3680 99.6594
R8456 gnd.n4575 gnd.n3681 99.6594
R8457 gnd.n4579 gnd.n3682 99.6594
R8458 gnd.n4583 gnd.n3683 99.6594
R8459 gnd.n3686 gnd.n3684 99.6594
R8460 gnd.n4589 gnd.n3685 99.6594
R8461 gnd.n5769 gnd.n2823 99.6594
R8462 gnd.n5761 gnd.n2793 99.6594
R8463 gnd.n5757 gnd.n2794 99.6594
R8464 gnd.n5753 gnd.n2795 99.6594
R8465 gnd.n5749 gnd.n2796 99.6594
R8466 gnd.n5745 gnd.n2797 99.6594
R8467 gnd.n5741 gnd.n2798 99.6594
R8468 gnd.n5736 gnd.n2800 99.6594
R8469 gnd.n5732 gnd.n2801 99.6594
R8470 gnd.n5728 gnd.n2802 99.6594
R8471 gnd.n5724 gnd.n2803 99.6594
R8472 gnd.n5720 gnd.n2804 99.6594
R8473 gnd.n5716 gnd.n2805 99.6594
R8474 gnd.n5712 gnd.n2806 99.6594
R8475 gnd.n5708 gnd.n2807 99.6594
R8476 gnd.n5704 gnd.n2808 99.6594
R8477 gnd.n2864 gnd.n2809 99.6594
R8478 gnd.n5696 gnd.n2810 99.6594
R8479 gnd.n172 gnd.n169 99.6594
R8480 gnd.n7374 gnd.n7373 99.6594
R8481 gnd.n168 gnd.n162 99.6594
R8482 gnd.n7381 gnd.n7380 99.6594
R8483 gnd.n161 gnd.n155 99.6594
R8484 gnd.n7388 gnd.n7387 99.6594
R8485 gnd.n154 gnd.n148 99.6594
R8486 gnd.n7395 gnd.n7394 99.6594
R8487 gnd.n147 gnd.n141 99.6594
R8488 gnd.n7402 gnd.n7401 99.6594
R8489 gnd.n140 gnd.n134 99.6594
R8490 gnd.n7412 gnd.n7411 99.6594
R8491 gnd.n133 gnd.n127 99.6594
R8492 gnd.n7419 gnd.n7418 99.6594
R8493 gnd.n126 gnd.n120 99.6594
R8494 gnd.n7426 gnd.n7425 99.6594
R8495 gnd.n119 gnd.n113 99.6594
R8496 gnd.n7433 gnd.n7432 99.6594
R8497 gnd.n112 gnd.n109 99.6594
R8498 gnd.n3599 gnd.n3528 99.6594
R8499 gnd.n3611 gnd.n3529 99.6594
R8500 gnd.n3595 gnd.n3530 99.6594
R8501 gnd.n3622 gnd.n3531 99.6594
R8502 gnd.n3635 gnd.n3532 99.6594
R8503 gnd.n3583 gnd.n3533 99.6594
R8504 gnd.n3646 gnd.n3534 99.6594
R8505 gnd.n3658 gnd.n3535 99.6594
R8506 gnd.n3558 gnd.n3536 99.6594
R8507 gnd.n4599 gnd.n3537 99.6594
R8508 gnd.n3553 gnd.n3538 99.6594
R8509 gnd.n4608 gnd.n3539 99.6594
R8510 gnd.n3549 gnd.n3540 99.6594
R8511 gnd.n4617 gnd.n3541 99.6594
R8512 gnd.n3610 gnd.n3528 99.6594
R8513 gnd.n3594 gnd.n3529 99.6594
R8514 gnd.n3623 gnd.n3530 99.6594
R8515 gnd.n3634 gnd.n3531 99.6594
R8516 gnd.n3582 gnd.n3532 99.6594
R8517 gnd.n3647 gnd.n3533 99.6594
R8518 gnd.n3657 gnd.n3534 99.6594
R8519 gnd.n3557 gnd.n3535 99.6594
R8520 gnd.n4598 gnd.n3536 99.6594
R8521 gnd.n3552 gnd.n3537 99.6594
R8522 gnd.n4607 gnd.n3538 99.6594
R8523 gnd.n3548 gnd.n3539 99.6594
R8524 gnd.n4616 gnd.n3540 99.6594
R8525 gnd.n3542 gnd.n3541 99.6594
R8526 gnd.n3136 gnd.n2781 99.6594
R8527 gnd.n3139 gnd.n3138 99.6594
R8528 gnd.n3153 gnd.n3152 99.6594
R8529 gnd.n3156 gnd.n3155 99.6594
R8530 gnd.n3170 gnd.n3169 99.6594
R8531 gnd.n3173 gnd.n3172 99.6594
R8532 gnd.n3187 gnd.n3186 99.6594
R8533 gnd.n3190 gnd.n3189 99.6594
R8534 gnd.n3202 gnd.n3201 99.6594
R8535 gnd.n3205 gnd.n3204 99.6594
R8536 gnd.n3208 gnd.n3207 99.6594
R8537 gnd.n3213 gnd.n3212 99.6594
R8538 gnd.n3216 gnd.n3215 99.6594
R8539 gnd.n5450 gnd.n5449 99.6594
R8540 gnd.n5451 gnd.n5450 99.6594
R8541 gnd.n3217 gnd.n3216 99.6594
R8542 gnd.n3214 gnd.n3213 99.6594
R8543 gnd.n3209 gnd.n3208 99.6594
R8544 gnd.n3206 gnd.n3205 99.6594
R8545 gnd.n3203 gnd.n3202 99.6594
R8546 gnd.n3189 gnd.n3086 99.6594
R8547 gnd.n3188 gnd.n3187 99.6594
R8548 gnd.n3172 gnd.n3098 99.6594
R8549 gnd.n3171 gnd.n3170 99.6594
R8550 gnd.n3155 gnd.n3107 99.6594
R8551 gnd.n3154 gnd.n3153 99.6594
R8552 gnd.n3138 gnd.n3116 99.6594
R8553 gnd.n3137 gnd.n3136 99.6594
R8554 gnd.n3545 gnd.t148 98.63
R8555 gnd.n7312 gnd.t80 98.63
R8556 gnd.n3091 gnd.t105 98.63
R8557 gnd.n3560 gnd.t140 98.63
R8558 gnd.n2844 gnd.t102 98.63
R8559 gnd.n2866 gnd.t88 98.63
R8560 gnd.n175 gnd.t180 98.63
R8561 gnd.n7405 gnd.t90 98.63
R8562 gnd.n2373 gnd.t167 98.63
R8563 gnd.n2395 gnd.t158 98.63
R8564 gnd.n3728 gnd.t98 98.63
R8565 gnd.n3706 gnd.t133 98.63
R8566 gnd.n3994 gnd.t113 98.63
R8567 gnd.n5459 gnd.t116 98.63
R8568 gnd.n4309 gnd.t178 88.9408
R8569 gnd.n5165 gnd.t174 88.9408
R8570 gnd.n4364 gnd.t128 88.933
R8571 gnd.n5159 gnd.t120 88.933
R8572 gnd.n4339 gnd.n4338 81.8399
R8573 gnd.n1484 gnd.t94 74.8376
R8574 gnd.n1052 gnd.t138 74.8376
R8575 gnd.n4310 gnd.t177 72.8438
R8576 gnd.n5166 gnd.t175 72.8438
R8577 gnd.n4340 gnd.n4333 72.8411
R8578 gnd.n4346 gnd.n4331 72.8411
R8579 gnd.n5129 gnd.n5128 72.8411
R8580 gnd.n3546 gnd.t147 72.836
R8581 gnd.n4365 gnd.t127 72.836
R8582 gnd.n5160 gnd.t121 72.836
R8583 gnd.n7313 gnd.t81 72.836
R8584 gnd.n3092 gnd.t104 72.836
R8585 gnd.n3561 gnd.t141 72.836
R8586 gnd.n2845 gnd.t101 72.836
R8587 gnd.n2867 gnd.t87 72.836
R8588 gnd.n176 gnd.t181 72.836
R8589 gnd.n7406 gnd.t91 72.836
R8590 gnd.n2374 gnd.t166 72.836
R8591 gnd.n2396 gnd.t157 72.836
R8592 gnd.n3729 gnd.t99 72.836
R8593 gnd.n3707 gnd.t134 72.836
R8594 gnd.n3995 gnd.t112 72.836
R8595 gnd.n5460 gnd.t117 72.836
R8596 gnd.n5307 gnd.n5306 71.676
R8597 gnd.n5302 gnd.n5139 71.676
R8598 gnd.n5300 gnd.n5299 71.676
R8599 gnd.n5295 gnd.n5142 71.676
R8600 gnd.n5293 gnd.n5292 71.676
R8601 gnd.n5288 gnd.n5145 71.676
R8602 gnd.n5286 gnd.n5285 71.676
R8603 gnd.n5281 gnd.n5148 71.676
R8604 gnd.n5279 gnd.n5278 71.676
R8605 gnd.n5274 gnd.n5151 71.676
R8606 gnd.n5272 gnd.n5271 71.676
R8607 gnd.n5267 gnd.n5154 71.676
R8608 gnd.n5265 gnd.n5264 71.676
R8609 gnd.n5260 gnd.n5157 71.676
R8610 gnd.n5258 gnd.n5257 71.676
R8611 gnd.n5253 gnd.n5162 71.676
R8612 gnd.n5250 gnd.n5249 71.676
R8613 gnd.n5247 gnd.n5246 71.676
R8614 gnd.n5241 gnd.n5168 71.676
R8615 gnd.n5239 gnd.n5238 71.676
R8616 gnd.n5234 gnd.n5171 71.676
R8617 gnd.n5232 gnd.n5231 71.676
R8618 gnd.n5227 gnd.n5174 71.676
R8619 gnd.n5225 gnd.n5224 71.676
R8620 gnd.n5220 gnd.n5177 71.676
R8621 gnd.n5218 gnd.n5217 71.676
R8622 gnd.n5213 gnd.n5180 71.676
R8623 gnd.n5211 gnd.n5210 71.676
R8624 gnd.n5206 gnd.n5183 71.676
R8625 gnd.n5204 gnd.n5203 71.676
R8626 gnd.n5199 gnd.n5186 71.676
R8627 gnd.n5197 gnd.n5196 71.676
R8628 gnd.n5192 gnd.n5190 71.676
R8629 gnd.n4427 gnd.n4328 71.676
R8630 gnd.n4425 gnd.n4351 71.676
R8631 gnd.n4421 gnd.n4420 71.676
R8632 gnd.n4414 gnd.n4353 71.676
R8633 gnd.n4413 gnd.n4412 71.676
R8634 gnd.n4406 gnd.n4355 71.676
R8635 gnd.n4405 gnd.n4404 71.676
R8636 gnd.n4398 gnd.n4357 71.676
R8637 gnd.n4397 gnd.n4396 71.676
R8638 gnd.n4390 gnd.n4359 71.676
R8639 gnd.n4389 gnd.n4388 71.676
R8640 gnd.n4382 gnd.n4361 71.676
R8641 gnd.n4381 gnd.n4380 71.676
R8642 gnd.n4374 gnd.n4363 71.676
R8643 gnd.n4373 gnd.n4367 71.676
R8644 gnd.n4369 gnd.n4368 71.676
R8645 gnd.n4557 gnd.n4556 71.676
R8646 gnd.n4549 gnd.n4308 71.676
R8647 gnd.n4548 gnd.n4547 71.676
R8648 gnd.n4541 gnd.n4312 71.676
R8649 gnd.n4540 gnd.n4539 71.676
R8650 gnd.n4533 gnd.n4314 71.676
R8651 gnd.n4532 gnd.n4531 71.676
R8652 gnd.n4525 gnd.n4316 71.676
R8653 gnd.n4524 gnd.n4523 71.676
R8654 gnd.n4517 gnd.n4318 71.676
R8655 gnd.n4516 gnd.n4515 71.676
R8656 gnd.n4509 gnd.n4320 71.676
R8657 gnd.n4508 gnd.n4507 71.676
R8658 gnd.n4501 gnd.n4322 71.676
R8659 gnd.n4500 gnd.n4499 71.676
R8660 gnd.n4493 gnd.n4324 71.676
R8661 gnd.n4428 gnd.n4427 71.676
R8662 gnd.n4422 gnd.n4351 71.676
R8663 gnd.n4420 gnd.n4419 71.676
R8664 gnd.n4415 gnd.n4414 71.676
R8665 gnd.n4412 gnd.n4411 71.676
R8666 gnd.n4407 gnd.n4406 71.676
R8667 gnd.n4404 gnd.n4403 71.676
R8668 gnd.n4399 gnd.n4398 71.676
R8669 gnd.n4396 gnd.n4395 71.676
R8670 gnd.n4391 gnd.n4390 71.676
R8671 gnd.n4388 gnd.n4387 71.676
R8672 gnd.n4383 gnd.n4382 71.676
R8673 gnd.n4380 gnd.n4379 71.676
R8674 gnd.n4375 gnd.n4374 71.676
R8675 gnd.n4370 gnd.n4367 71.676
R8676 gnd.n4559 gnd.n4558 71.676
R8677 gnd.n4556 gnd.n4555 71.676
R8678 gnd.n4550 gnd.n4549 71.676
R8679 gnd.n4547 gnd.n4546 71.676
R8680 gnd.n4542 gnd.n4541 71.676
R8681 gnd.n4539 gnd.n4538 71.676
R8682 gnd.n4534 gnd.n4533 71.676
R8683 gnd.n4531 gnd.n4530 71.676
R8684 gnd.n4526 gnd.n4525 71.676
R8685 gnd.n4523 gnd.n4522 71.676
R8686 gnd.n4518 gnd.n4517 71.676
R8687 gnd.n4515 gnd.n4514 71.676
R8688 gnd.n4510 gnd.n4509 71.676
R8689 gnd.n4507 gnd.n4506 71.676
R8690 gnd.n4502 gnd.n4501 71.676
R8691 gnd.n4499 gnd.n4498 71.676
R8692 gnd.n4494 gnd.n4493 71.676
R8693 gnd.n5190 gnd.n5187 71.676
R8694 gnd.n5198 gnd.n5197 71.676
R8695 gnd.n5186 gnd.n5184 71.676
R8696 gnd.n5205 gnd.n5204 71.676
R8697 gnd.n5183 gnd.n5181 71.676
R8698 gnd.n5212 gnd.n5211 71.676
R8699 gnd.n5180 gnd.n5178 71.676
R8700 gnd.n5219 gnd.n5218 71.676
R8701 gnd.n5177 gnd.n5175 71.676
R8702 gnd.n5226 gnd.n5225 71.676
R8703 gnd.n5174 gnd.n5172 71.676
R8704 gnd.n5233 gnd.n5232 71.676
R8705 gnd.n5171 gnd.n5169 71.676
R8706 gnd.n5240 gnd.n5239 71.676
R8707 gnd.n5168 gnd.n5164 71.676
R8708 gnd.n5248 gnd.n5247 71.676
R8709 gnd.n5252 gnd.n5251 71.676
R8710 gnd.n5162 gnd.n5158 71.676
R8711 gnd.n5259 gnd.n5258 71.676
R8712 gnd.n5157 gnd.n5155 71.676
R8713 gnd.n5266 gnd.n5265 71.676
R8714 gnd.n5154 gnd.n5152 71.676
R8715 gnd.n5273 gnd.n5272 71.676
R8716 gnd.n5151 gnd.n5149 71.676
R8717 gnd.n5280 gnd.n5279 71.676
R8718 gnd.n5148 gnd.n5146 71.676
R8719 gnd.n5287 gnd.n5286 71.676
R8720 gnd.n5145 gnd.n5143 71.676
R8721 gnd.n5294 gnd.n5293 71.676
R8722 gnd.n5142 gnd.n5140 71.676
R8723 gnd.n5301 gnd.n5300 71.676
R8724 gnd.n5139 gnd.n5137 71.676
R8725 gnd.n5308 gnd.n5307 71.676
R8726 gnd.n8 gnd.t312 69.1507
R8727 gnd.n14 gnd.t314 68.4792
R8728 gnd.n13 gnd.t42 68.4792
R8729 gnd.n12 gnd.t322 68.4792
R8730 gnd.n11 gnd.t67 68.4792
R8731 gnd.n10 gnd.t19 68.4792
R8732 gnd.n9 gnd.t35 68.4792
R8733 gnd.n8 gnd.t25 68.4792
R8734 gnd.n1611 gnd.n1515 64.369
R8735 gnd.n4552 gnd.n4310 59.5399
R8736 gnd.n5243 gnd.n5166 59.5399
R8737 gnd.n4366 gnd.n4365 59.5399
R8738 gnd.n5161 gnd.n5160 59.5399
R8739 gnd.n4431 gnd.n4349 59.1804
R8740 gnd.n6195 gnd.n1043 57.3586
R8741 gnd.n6148 gnd.n2351 57.3586
R8742 gnd.n7442 gnd.n102 57.3586
R8743 gnd.n1266 gnd.t188 56.607
R8744 gnd.n48 gnd.t287 56.607
R8745 gnd.n1235 gnd.t249 56.407
R8746 gnd.n1250 gnd.t227 56.407
R8747 gnd.n17 gnd.t282 56.407
R8748 gnd.n32 gnd.t258 56.407
R8749 gnd.n1279 gnd.t299 55.8337
R8750 gnd.n1248 gnd.t256 55.8337
R8751 gnd.n1263 gnd.t237 55.8337
R8752 gnd.n61 gnd.t265 55.8337
R8753 gnd.n30 gnd.t289 55.8337
R8754 gnd.n45 gnd.t266 55.8337
R8755 gnd.n4337 gnd.n4336 54.358
R8756 gnd.n5126 gnd.n5125 54.358
R8757 gnd.n1266 gnd.n1265 53.0052
R8758 gnd.n1268 gnd.n1267 53.0052
R8759 gnd.n1270 gnd.n1269 53.0052
R8760 gnd.n1272 gnd.n1271 53.0052
R8761 gnd.n1274 gnd.n1273 53.0052
R8762 gnd.n1276 gnd.n1275 53.0052
R8763 gnd.n1278 gnd.n1277 53.0052
R8764 gnd.n1235 gnd.n1234 53.0052
R8765 gnd.n1237 gnd.n1236 53.0052
R8766 gnd.n1239 gnd.n1238 53.0052
R8767 gnd.n1241 gnd.n1240 53.0052
R8768 gnd.n1243 gnd.n1242 53.0052
R8769 gnd.n1245 gnd.n1244 53.0052
R8770 gnd.n1247 gnd.n1246 53.0052
R8771 gnd.n1250 gnd.n1249 53.0052
R8772 gnd.n1252 gnd.n1251 53.0052
R8773 gnd.n1254 gnd.n1253 53.0052
R8774 gnd.n1256 gnd.n1255 53.0052
R8775 gnd.n1258 gnd.n1257 53.0052
R8776 gnd.n1260 gnd.n1259 53.0052
R8777 gnd.n1262 gnd.n1261 53.0052
R8778 gnd.n60 gnd.n59 53.0052
R8779 gnd.n58 gnd.n57 53.0052
R8780 gnd.n56 gnd.n55 53.0052
R8781 gnd.n54 gnd.n53 53.0052
R8782 gnd.n52 gnd.n51 53.0052
R8783 gnd.n50 gnd.n49 53.0052
R8784 gnd.n48 gnd.n47 53.0052
R8785 gnd.n29 gnd.n28 53.0052
R8786 gnd.n27 gnd.n26 53.0052
R8787 gnd.n25 gnd.n24 53.0052
R8788 gnd.n23 gnd.n22 53.0052
R8789 gnd.n21 gnd.n20 53.0052
R8790 gnd.n19 gnd.n18 53.0052
R8791 gnd.n17 gnd.n16 53.0052
R8792 gnd.n44 gnd.n43 53.0052
R8793 gnd.n42 gnd.n41 53.0052
R8794 gnd.n40 gnd.n39 53.0052
R8795 gnd.n38 gnd.n37 53.0052
R8796 gnd.n36 gnd.n35 53.0052
R8797 gnd.n34 gnd.n33 53.0052
R8798 gnd.n32 gnd.n31 53.0052
R8799 gnd.n5117 gnd.n5116 52.4801
R8800 gnd.n2275 gnd.t37 52.3082
R8801 gnd.n2243 gnd.t70 52.3082
R8802 gnd.n2211 gnd.t40 52.3082
R8803 gnd.n2180 gnd.t316 52.3082
R8804 gnd.n2148 gnd.t320 52.3082
R8805 gnd.n2116 gnd.t23 52.3082
R8806 gnd.n2084 gnd.t318 52.3082
R8807 gnd.n2053 gnd.t29 52.3082
R8808 gnd.n2105 gnd.n2073 51.4173
R8809 gnd.n2169 gnd.n2168 50.455
R8810 gnd.n2137 gnd.n2136 50.455
R8811 gnd.n2105 gnd.n2104 50.455
R8812 gnd.n1558 gnd.n1557 45.1884
R8813 gnd.n1073 gnd.n1072 45.1884
R8814 gnd.n5133 gnd.n5132 44.3322
R8815 gnd.n4340 gnd.n4339 44.3189
R8816 gnd.n4614 gnd.n3546 42.2793
R8817 gnd.n1559 gnd.n1558 42.2793
R8818 gnd.n1074 gnd.n1073 42.2793
R8819 gnd.n1485 gnd.n1484 42.2793
R8820 gnd.n1053 gnd.n1052 42.2793
R8821 gnd.n7318 gnd.n7313 42.2793
R8822 gnd.n3196 gnd.n3092 42.2793
R8823 gnd.n3562 gnd.n3561 42.2793
R8824 gnd.n2868 gnd.n2867 42.2793
R8825 gnd.n7370 gnd.n176 42.2793
R8826 gnd.n7407 gnd.n7406 42.2793
R8827 gnd.n6112 gnd.n2374 42.2793
R8828 gnd.n2397 gnd.n2396 42.2793
R8829 gnd.n4263 gnd.n3729 42.2793
R8830 gnd.n3996 gnd.n3995 42.2793
R8831 gnd.n5461 gnd.n5460 42.2793
R8832 gnd.n6422 gnd.n799 42.1703
R8833 gnd.n6416 gnd.n799 42.1703
R8834 gnd.n6416 gnd.n6415 42.1703
R8835 gnd.n6415 gnd.n6414 42.1703
R8836 gnd.n6414 gnd.n806 42.1703
R8837 gnd.n6408 gnd.n806 42.1703
R8838 gnd.n6408 gnd.n6407 42.1703
R8839 gnd.n6407 gnd.n6406 42.1703
R8840 gnd.n6406 gnd.n814 42.1703
R8841 gnd.n6400 gnd.n814 42.1703
R8842 gnd.n6400 gnd.n6399 42.1703
R8843 gnd.n6399 gnd.n6398 42.1703
R8844 gnd.n6398 gnd.n822 42.1703
R8845 gnd.n6392 gnd.n822 42.1703
R8846 gnd.n6392 gnd.n6391 42.1703
R8847 gnd.n6391 gnd.n6390 42.1703
R8848 gnd.n6390 gnd.n830 42.1703
R8849 gnd.n6384 gnd.n830 42.1703
R8850 gnd.n6384 gnd.n6383 42.1703
R8851 gnd.n6383 gnd.n6382 42.1703
R8852 gnd.n6382 gnd.n838 42.1703
R8853 gnd.n6376 gnd.n838 42.1703
R8854 gnd.n6376 gnd.n6375 42.1703
R8855 gnd.n6375 gnd.n6374 42.1703
R8856 gnd.n6374 gnd.n846 42.1703
R8857 gnd.n6368 gnd.n846 42.1703
R8858 gnd.n6368 gnd.n6367 42.1703
R8859 gnd.n6367 gnd.n6366 42.1703
R8860 gnd.n6366 gnd.n854 42.1703
R8861 gnd.n6360 gnd.n854 42.1703
R8862 gnd.n6360 gnd.n6359 42.1703
R8863 gnd.n6359 gnd.n6358 42.1703
R8864 gnd.n6358 gnd.n862 42.1703
R8865 gnd.n6352 gnd.n862 42.1703
R8866 gnd.n6352 gnd.n6351 42.1703
R8867 gnd.n6351 gnd.n6350 42.1703
R8868 gnd.n6350 gnd.n870 42.1703
R8869 gnd.n6344 gnd.n870 42.1703
R8870 gnd.n6344 gnd.n6343 42.1703
R8871 gnd.n6343 gnd.n6342 42.1703
R8872 gnd.n6342 gnd.n878 42.1703
R8873 gnd.n6336 gnd.n878 42.1703
R8874 gnd.n6336 gnd.n6335 42.1703
R8875 gnd.n6335 gnd.n6334 42.1703
R8876 gnd.n6334 gnd.n886 42.1703
R8877 gnd.n6328 gnd.n886 42.1703
R8878 gnd.n6328 gnd.n6327 42.1703
R8879 gnd.n6327 gnd.n6326 42.1703
R8880 gnd.n6326 gnd.n894 42.1703
R8881 gnd.n6320 gnd.n894 42.1703
R8882 gnd.n6320 gnd.n6319 42.1703
R8883 gnd.n6319 gnd.n6318 42.1703
R8884 gnd.n6318 gnd.n902 42.1703
R8885 gnd.n6312 gnd.n902 42.1703
R8886 gnd.n6312 gnd.n6311 42.1703
R8887 gnd.n6311 gnd.n6310 42.1703
R8888 gnd.n6310 gnd.n910 42.1703
R8889 gnd.n6304 gnd.n910 42.1703
R8890 gnd.n6304 gnd.n6303 42.1703
R8891 gnd.n6303 gnd.n6302 42.1703
R8892 gnd.n6302 gnd.n918 42.1703
R8893 gnd.n6296 gnd.n918 42.1703
R8894 gnd.n6296 gnd.n6295 42.1703
R8895 gnd.n6295 gnd.n6294 42.1703
R8896 gnd.n6294 gnd.n926 42.1703
R8897 gnd.n6288 gnd.n926 42.1703
R8898 gnd.n6288 gnd.n6287 42.1703
R8899 gnd.n6287 gnd.n6286 42.1703
R8900 gnd.n6286 gnd.n934 42.1703
R8901 gnd.n6280 gnd.n934 42.1703
R8902 gnd.n6280 gnd.n6279 42.1703
R8903 gnd.n6279 gnd.n6278 42.1703
R8904 gnd.n6278 gnd.n942 42.1703
R8905 gnd.n6272 gnd.n942 42.1703
R8906 gnd.n6272 gnd.n6271 42.1703
R8907 gnd.n6271 gnd.n6270 42.1703
R8908 gnd.n6270 gnd.n950 42.1703
R8909 gnd.n6264 gnd.n950 42.1703
R8910 gnd.n6264 gnd.n6263 42.1703
R8911 gnd.n6263 gnd.n6262 42.1703
R8912 gnd.n6262 gnd.n958 42.1703
R8913 gnd.n6256 gnd.n958 42.1703
R8914 gnd.n6256 gnd.n6255 42.1703
R8915 gnd.n4338 gnd.n4337 41.6274
R8916 gnd.n5127 gnd.n5126 41.6274
R8917 gnd.n4347 gnd.n4346 40.8975
R8918 gnd.n5130 gnd.n5129 40.8975
R8919 gnd.n5738 gnd.n2845 36.9518
R8920 gnd.n4561 gnd.n3707 36.9518
R8921 gnd.n4346 gnd.n4345 35.055
R8922 gnd.n4341 gnd.n4340 35.055
R8923 gnd.n5119 gnd.n5118 35.055
R8924 gnd.n5129 gnd.n5115 35.055
R8925 gnd.n1621 gnd.n1515 31.8661
R8926 gnd.n1621 gnd.n1620 31.8661
R8927 gnd.n1629 gnd.n1504 31.8661
R8928 gnd.n1637 gnd.n1504 31.8661
R8929 gnd.n1637 gnd.n1498 31.8661
R8930 gnd.n1645 gnd.n1498 31.8661
R8931 gnd.n1645 gnd.n1491 31.8661
R8932 gnd.n1683 gnd.n1491 31.8661
R8933 gnd.n1693 gnd.n1424 31.8661
R8934 gnd.n4052 gnd.n2351 31.8661
R8935 gnd.n6061 gnd.n2405 31.8661
R8936 gnd.n3564 gnd.n2672 31.8661
R8937 gnd.n3666 gnd.n3527 31.8661
R8938 gnd.n4624 gnd.n3527 31.8661
R8939 gnd.n4625 gnd.n4624 31.8661
R8940 gnd.n4625 gnd.n3521 31.8661
R8941 gnd.n4633 gnd.n3521 31.8661
R8942 gnd.n4641 gnd.n3514 31.8661
R8943 gnd.n4641 gnd.n3507 31.8661
R8944 gnd.n4649 gnd.n3507 31.8661
R8945 gnd.n4649 gnd.n3508 31.8661
R8946 gnd.n4657 gnd.n3494 31.8661
R8947 gnd.n4665 gnd.n3494 31.8661
R8948 gnd.n4665 gnd.n3495 31.8661
R8949 gnd.n4673 gnd.n3488 31.8661
R8950 gnd.n5397 gnd.n3256 31.8661
R8951 gnd.n5405 gnd.n3242 31.8661
R8952 gnd.n5413 gnd.n3242 31.8661
R8953 gnd.n5413 gnd.n3244 31.8661
R8954 gnd.n5421 gnd.n3230 31.8661
R8955 gnd.n5431 gnd.n3230 31.8661
R8956 gnd.n5431 gnd.n3223 31.8661
R8957 gnd.n5442 gnd.n3223 31.8661
R8958 gnd.n5779 gnd.n2782 31.8661
R8959 gnd.n5779 gnd.n5778 31.8661
R8960 gnd.n5778 gnd.n2785 31.8661
R8961 gnd.n5772 gnd.n2785 31.8661
R8962 gnd.n5772 gnd.n5771 31.8661
R8963 gnd.n2872 gnd.n2821 31.8661
R8964 gnd.n7362 gnd.n181 31.8661
R8965 gnd.n7442 gnd.n100 31.8661
R8966 gnd.n3495 gnd.t311 30.9101
R8967 gnd.n5405 gnd.t16 30.9101
R8968 gnd.n5193 gnd.n5189 29.8151
R8969 gnd.n4495 gnd.n4325 29.8151
R8970 gnd.n4590 gnd.n3666 27.4049
R8971 gnd.n5771 gnd.n5770 27.4049
R8972 gnd.n3546 gnd.n3545 25.7944
R8973 gnd.n1484 gnd.n1483 25.7944
R8974 gnd.n1052 gnd.n1051 25.7944
R8975 gnd.n7313 gnd.n7312 25.7944
R8976 gnd.n3092 gnd.n3091 25.7944
R8977 gnd.n3561 gnd.n3560 25.7944
R8978 gnd.n2845 gnd.n2844 25.7944
R8979 gnd.n2867 gnd.n2866 25.7944
R8980 gnd.n176 gnd.n175 25.7944
R8981 gnd.n7406 gnd.n7405 25.7944
R8982 gnd.n2374 gnd.n2373 25.7944
R8983 gnd.n2396 gnd.n2395 25.7944
R8984 gnd.n3729 gnd.n3728 25.7944
R8985 gnd.n3707 gnd.n3706 25.7944
R8986 gnd.n3995 gnd.n3994 25.7944
R8987 gnd.n5460 gnd.n5459 25.7944
R8988 gnd.n5135 gnd.n3262 25.493
R8989 gnd.n6255 gnd.n6254 25.3024
R8990 gnd.n1705 gnd.n1425 24.8557
R8991 gnd.n1715 gnd.n1408 24.8557
R8992 gnd.n1411 gnd.n1399 24.8557
R8993 gnd.n1736 gnd.n1400 24.8557
R8994 gnd.n1746 gnd.n1380 24.8557
R8995 gnd.n1756 gnd.n1755 24.8557
R8996 gnd.n1366 gnd.n1364 24.8557
R8997 gnd.n1787 gnd.n1786 24.8557
R8998 gnd.n1802 gnd.n1349 24.8557
R8999 gnd.n1856 gnd.n1288 24.8557
R9000 gnd.n1812 gnd.n1289 24.8557
R9001 gnd.n1849 gnd.n1300 24.8557
R9002 gnd.n1338 gnd.n1337 24.8557
R9003 gnd.n1843 gnd.n1842 24.8557
R9004 gnd.n1324 gnd.n1311 24.8557
R9005 gnd.n1882 gnd.n1881 24.8557
R9006 gnd.n1892 gnd.n1220 24.8557
R9007 gnd.n1904 gnd.n1212 24.8557
R9008 gnd.n1903 gnd.n1200 24.8557
R9009 gnd.n1922 gnd.n1921 24.8557
R9010 gnd.n1932 gnd.n1193 24.8557
R9011 gnd.n1945 gnd.n1181 24.8557
R9012 gnd.n1996 gnd.n1995 24.8557
R9013 gnd.n2011 gnd.n1165 24.8557
R9014 gnd.n2010 gnd.n1167 24.8557
R9015 gnd.n6247 gnd.n977 24.8557
R9016 gnd.n6246 gnd.n980 24.8557
R9017 gnd.n6240 gnd.n6239 24.8557
R9018 gnd.n6233 gnd.n1001 24.8557
R9019 gnd.n6232 gnd.n1004 24.8557
R9020 gnd.n6226 gnd.n6225 24.8557
R9021 gnd.n1968 gnd.n1018 24.8557
R9022 gnd.n6219 gnd.n1027 24.8557
R9023 gnd.n6212 gnd.n6211 24.8557
R9024 gnd.n1726 gnd.t28 23.2624
R9025 gnd.n1427 gnd.t93 22.6251
R9026 gnd.n4052 gnd.t111 22.6251
R9027 gnd.t79 gnd.n100 22.6251
R9028 gnd.n4476 gnd.n3467 21.6691
R9029 gnd.n4469 gnd.n3461 21.6691
R9030 gnd.n4461 gnd.n3453 21.6691
R9031 gnd.n4838 gnd.n3431 21.6691
R9032 gnd.n4826 gnd.n3425 21.6691
R9033 gnd.n4818 gnd.n3419 21.6691
R9034 gnd.n4796 gnd.n4795 21.6691
R9035 gnd.n4787 gnd.n3394 21.6691
R9036 gnd.n5015 gnd.n3365 21.6691
R9037 gnd.n5015 gnd.n3367 21.6691
R9038 gnd.n4995 gnd.n3352 21.6691
R9039 gnd.n4988 gnd.n3346 21.6691
R9040 gnd.n4965 gnd.n3323 21.6691
R9041 gnd.n4958 gnd.n3316 21.6691
R9042 gnd.n5349 gnd.n3294 21.6691
R9043 gnd.n5337 gnd.n3287 21.6691
R9044 gnd.n5329 gnd.n3281 21.6691
R9045 gnd.t315 gnd.n1432 21.3504
R9046 gnd.n3488 gnd.n3481 21.3504
R9047 gnd.n6061 gnd.n2407 21.0318
R9048 gnd.n4059 gnd.n2417 21.0318
R9049 gnd.n6055 gnd.n2420 21.0318
R9050 gnd.n6049 gnd.n2432 21.0318
R9051 gnd.n4076 gnd.n2440 21.0318
R9052 gnd.n4084 gnd.n2450 21.0318
R9053 gnd.n6037 gnd.n2453 21.0318
R9054 gnd.n4092 gnd.n2461 21.0318
R9055 gnd.n6031 gnd.n2464 21.0318
R9056 gnd.n6025 gnd.n2475 21.0318
R9057 gnd.n4108 gnd.n2483 21.0318
R9058 gnd.n4116 gnd.n2493 21.0318
R9059 gnd.n6013 gnd.n2496 21.0318
R9060 gnd.n4124 gnd.n2504 21.0318
R9061 gnd.n6007 gnd.n2507 21.0318
R9062 gnd.n6001 gnd.n2518 21.0318
R9063 gnd.n4140 gnd.n2524 21.0318
R9064 gnd.n4150 gnd.n2534 21.0318
R9065 gnd.n5989 gnd.n2537 21.0318
R9066 gnd.n4159 gnd.n2542 21.0318
R9067 gnd.n5982 gnd.n2545 21.0318
R9068 gnd.n5976 gnd.n2556 21.0318
R9069 gnd.n4175 gnd.n2563 21.0318
R9070 gnd.n4183 gnd.n2573 21.0318
R9071 gnd.n5964 gnd.n2576 21.0318
R9072 gnd.n4191 gnd.n2584 21.0318
R9073 gnd.n5958 gnd.n2587 21.0318
R9074 gnd.n5952 gnd.n2598 21.0318
R9075 gnd.n4207 gnd.n2606 21.0318
R9076 gnd.n4215 gnd.n2616 21.0318
R9077 gnd.n5940 gnd.n2619 21.0318
R9078 gnd.n4223 gnd.n2627 21.0318
R9079 gnd.n5934 gnd.n2630 21.0318
R9080 gnd.n5928 gnd.n2641 21.0318
R9081 gnd.n4239 gnd.n2649 21.0318
R9082 gnd.n5922 gnd.n2652 21.0318
R9083 gnd.n4248 gnd.n2660 21.0318
R9084 gnd.n4256 gnd.n2669 21.0318
R9085 gnd.n5910 gnd.n2672 21.0318
R9086 gnd.n4681 gnd.t83 21.0318
R9087 gnd.t1 gnd.n3413 21.0318
R9088 gnd.n4973 gnd.t9 21.0318
R9089 gnd.n5694 gnd.n2872 21.0318
R9090 gnd.n3041 gnd.n2874 21.0318
R9091 gnd.n5491 gnd.n3019 21.0318
R9092 gnd.n5490 gnd.n3022 21.0318
R9093 gnd.n5501 gnd.n3009 21.0318
R9094 gnd.n3011 gnd.n3001 21.0318
R9095 gnd.n5522 gnd.n2990 21.0318
R9096 gnd.n5521 gnd.n2994 21.0318
R9097 gnd.n5532 gnd.n2981 21.0318
R9098 gnd.n2983 gnd.n2973 21.0318
R9099 gnd.n5561 gnd.n2962 21.0318
R9100 gnd.n5559 gnd.n2965 21.0318
R9101 gnd.n2956 gnd.n2954 21.0318
R9102 gnd.n5584 gnd.n2946 21.0318
R9103 gnd.n5651 gnd.n2910 21.0318
R9104 gnd.n5650 gnd.n2913 21.0318
R9105 gnd.n5597 gnd.n2904 21.0318
R9106 gnd.n7200 gnd.n273 21.0318
R9107 gnd.n5608 gnd.n2926 21.0318
R9108 gnd.n5637 gnd.n5636 21.0318
R9109 gnd.n5632 gnd.n2932 21.0318
R9110 gnd.n5631 gnd.n5620 21.0318
R9111 gnd.n7184 gnd.n290 21.0318
R9112 gnd.n7173 gnd.n292 21.0318
R9113 gnd.n310 gnd.n260 21.0318
R9114 gnd.n7215 gnd.n252 21.0318
R9115 gnd.n7164 gnd.n7163 21.0318
R9116 gnd.n7223 gnd.n244 21.0318
R9117 gnd.n7231 gnd.n236 21.0318
R9118 gnd.n7152 gnd.n238 21.0318
R9119 gnd.n342 gnd.n230 21.0318
R9120 gnd.n7247 gnd.n222 21.0318
R9121 gnd.n7144 gnd.n7143 21.0318
R9122 gnd.n7255 gnd.n214 21.0318
R9123 gnd.n7263 gnd.n206 21.0318
R9124 gnd.n7132 gnd.n208 21.0318
R9125 gnd.n359 gnd.n200 21.0318
R9126 gnd.n7354 gnd.n189 21.0318
R9127 gnd.n191 gnd.n181 21.0318
R9128 gnd.t45 gnd.n989 20.7131
R9129 gnd.n4657 gnd.t73 20.7131
R9130 gnd.n3244 gnd.t313 20.7131
R9131 gnd.t47 gnd.n1174 20.0758
R9132 gnd.n4334 gnd.t131 19.8005
R9133 gnd.n4334 gnd.t164 19.8005
R9134 gnd.n4335 gnd.t161 19.8005
R9135 gnd.n4335 gnd.t172 19.8005
R9136 gnd.n5123 gnd.t77 19.8005
R9137 gnd.n5123 gnd.t155 19.8005
R9138 gnd.n5124 gnd.t170 19.8005
R9139 gnd.n5124 gnd.t144 19.8005
R9140 gnd.n4331 gnd.n4330 19.5087
R9141 gnd.n4344 gnd.n4331 19.5087
R9142 gnd.n4342 gnd.n4333 19.5087
R9143 gnd.n5128 gnd.n5122 19.5087
R9144 gnd.n1893 gnd.t53 19.4385
R9145 gnd.n4635 gnd.n3519 19.3944
R9146 gnd.n4635 gnd.n3517 19.3944
R9147 gnd.n4639 gnd.n3517 19.3944
R9148 gnd.n4639 gnd.n3505 19.3944
R9149 gnd.n4651 gnd.n3505 19.3944
R9150 gnd.n4651 gnd.n3503 19.3944
R9151 gnd.n4655 gnd.n3503 19.3944
R9152 gnd.n4655 gnd.n3492 19.3944
R9153 gnd.n4667 gnd.n3492 19.3944
R9154 gnd.n4667 gnd.n3490 19.3944
R9155 gnd.n4671 gnd.n3490 19.3944
R9156 gnd.n4671 gnd.n3479 19.3944
R9157 gnd.n4683 gnd.n3479 19.3944
R9158 gnd.n4683 gnd.n3477 19.3944
R9159 gnd.n4687 gnd.n3477 19.3944
R9160 gnd.n4687 gnd.n3465 19.3944
R9161 gnd.n4699 gnd.n3465 19.3944
R9162 gnd.n4699 gnd.n3463 19.3944
R9163 gnd.n4703 gnd.n3463 19.3944
R9164 gnd.n4703 gnd.n3451 19.3944
R9165 gnd.n4717 gnd.n3451 19.3944
R9166 gnd.n4717 gnd.n3448 19.3944
R9167 gnd.n4722 gnd.n3448 19.3944
R9168 gnd.n4722 gnd.n3449 19.3944
R9169 gnd.n3449 gnd.n3423 19.3944
R9170 gnd.n4848 gnd.n3423 19.3944
R9171 gnd.n4848 gnd.n3421 19.3944
R9172 gnd.n4852 gnd.n3421 19.3944
R9173 gnd.n4852 gnd.n3411 19.3944
R9174 gnd.n4864 gnd.n3411 19.3944
R9175 gnd.n4864 gnd.n3409 19.3944
R9176 gnd.n4868 gnd.n3409 19.3944
R9177 gnd.n4868 gnd.n3398 19.3944
R9178 gnd.n4880 gnd.n3398 19.3944
R9179 gnd.n4880 gnd.n3396 19.3944
R9180 gnd.n4884 gnd.n3396 19.3944
R9181 gnd.n4884 gnd.n3384 19.3944
R9182 gnd.n4898 gnd.n3384 19.3944
R9183 gnd.n4898 gnd.n3381 19.3944
R9184 gnd.n4903 gnd.n3381 19.3944
R9185 gnd.n4903 gnd.n3382 19.3944
R9186 gnd.n3382 gnd.n3356 19.3944
R9187 gnd.n5025 gnd.n3356 19.3944
R9188 gnd.n5025 gnd.n3354 19.3944
R9189 gnd.n5029 gnd.n3354 19.3944
R9190 gnd.n5029 gnd.n3342 19.3944
R9191 gnd.n5041 gnd.n3342 19.3944
R9192 gnd.n5041 gnd.n3340 19.3944
R9193 gnd.n5045 gnd.n3340 19.3944
R9194 gnd.n5045 gnd.n3327 19.3944
R9195 gnd.n5057 gnd.n3327 19.3944
R9196 gnd.n5057 gnd.n3325 19.3944
R9197 gnd.n5061 gnd.n3325 19.3944
R9198 gnd.n5061 gnd.n3312 19.3944
R9199 gnd.n5075 gnd.n3312 19.3944
R9200 gnd.n5075 gnd.n3309 19.3944
R9201 gnd.n5080 gnd.n3309 19.3944
R9202 gnd.n5080 gnd.n3310 19.3944
R9203 gnd.n3310 gnd.n3285 19.3944
R9204 gnd.n5359 gnd.n3285 19.3944
R9205 gnd.n5359 gnd.n3283 19.3944
R9206 gnd.n5363 gnd.n3283 19.3944
R9207 gnd.n5363 gnd.n3272 19.3944
R9208 gnd.n5375 gnd.n3272 19.3944
R9209 gnd.n5375 gnd.n3270 19.3944
R9210 gnd.n5379 gnd.n3270 19.3944
R9211 gnd.n5379 gnd.n3260 19.3944
R9212 gnd.n5391 gnd.n3260 19.3944
R9213 gnd.n5391 gnd.n3258 19.3944
R9214 gnd.n5395 gnd.n3258 19.3944
R9215 gnd.n5395 gnd.n3248 19.3944
R9216 gnd.n5407 gnd.n3248 19.3944
R9217 gnd.n5407 gnd.n3246 19.3944
R9218 gnd.n5411 gnd.n3246 19.3944
R9219 gnd.n5411 gnd.n3235 19.3944
R9220 gnd.n5423 gnd.n3235 19.3944
R9221 gnd.n5423 gnd.n3232 19.3944
R9222 gnd.n5429 gnd.n3232 19.3944
R9223 gnd.n5429 gnd.n3233 19.3944
R9224 gnd.n3233 gnd.n3220 19.3944
R9225 gnd.n5445 gnd.n3220 19.3944
R9226 gnd.n5446 gnd.n5445 19.3944
R9227 gnd.n4618 gnd.n4615 19.3944
R9228 gnd.n4618 gnd.n3543 19.3944
R9229 gnd.n4622 gnd.n3543 19.3944
R9230 gnd.n3609 gnd.n3600 19.3944
R9231 gnd.n3612 gnd.n3609 19.3944
R9232 gnd.n3612 gnd.n3593 19.3944
R9233 gnd.n3621 gnd.n3593 19.3944
R9234 gnd.n3624 gnd.n3621 19.3944
R9235 gnd.n3624 gnd.n3587 19.3944
R9236 gnd.n3633 gnd.n3587 19.3944
R9237 gnd.n3636 gnd.n3633 19.3944
R9238 gnd.n3636 gnd.n3581 19.3944
R9239 gnd.n3645 gnd.n3581 19.3944
R9240 gnd.n3648 gnd.n3645 19.3944
R9241 gnd.n3648 gnd.n3575 19.3944
R9242 gnd.n3656 gnd.n3575 19.3944
R9243 gnd.n3659 gnd.n3656 19.3944
R9244 gnd.n3659 gnd.n3556 19.3944
R9245 gnd.n4596 gnd.n3556 19.3944
R9246 gnd.n4597 gnd.n4596 19.3944
R9247 gnd.n4600 gnd.n4597 19.3944
R9248 gnd.n4600 gnd.n3551 19.3944
R9249 gnd.n4605 gnd.n3551 19.3944
R9250 gnd.n4606 gnd.n4605 19.3944
R9251 gnd.n4609 gnd.n4606 19.3944
R9252 gnd.n4609 gnd.n3547 19.3944
R9253 gnd.n4613 gnd.n3547 19.3944
R9254 gnd.n1608 gnd.n1607 19.3944
R9255 gnd.n1607 gnd.n1606 19.3944
R9256 gnd.n1606 gnd.n1605 19.3944
R9257 gnd.n1605 gnd.n1603 19.3944
R9258 gnd.n1603 gnd.n1600 19.3944
R9259 gnd.n1600 gnd.n1599 19.3944
R9260 gnd.n1599 gnd.n1596 19.3944
R9261 gnd.n1596 gnd.n1595 19.3944
R9262 gnd.n1595 gnd.n1592 19.3944
R9263 gnd.n1592 gnd.n1591 19.3944
R9264 gnd.n1591 gnd.n1588 19.3944
R9265 gnd.n1588 gnd.n1587 19.3944
R9266 gnd.n1587 gnd.n1584 19.3944
R9267 gnd.n1584 gnd.n1583 19.3944
R9268 gnd.n1583 gnd.n1580 19.3944
R9269 gnd.n1580 gnd.n1579 19.3944
R9270 gnd.n1579 gnd.n1576 19.3944
R9271 gnd.n1576 gnd.n1575 19.3944
R9272 gnd.n1575 gnd.n1572 19.3944
R9273 gnd.n1572 gnd.n1571 19.3944
R9274 gnd.n1571 gnd.n1568 19.3944
R9275 gnd.n1568 gnd.n1567 19.3944
R9276 gnd.n1564 gnd.n1563 19.3944
R9277 gnd.n1563 gnd.n1519 19.3944
R9278 gnd.n1614 gnd.n1519 19.3944
R9279 gnd.n1146 gnd.n1144 19.3944
R9280 gnd.n1146 gnd.n1070 19.3944
R9281 gnd.n2320 gnd.n1070 19.3944
R9282 gnd.n1087 gnd.n1086 19.3944
R9283 gnd.n1091 gnd.n1086 19.3944
R9284 gnd.n1094 gnd.n1091 19.3944
R9285 gnd.n1097 gnd.n1094 19.3944
R9286 gnd.n1097 gnd.n1083 19.3944
R9287 gnd.n1101 gnd.n1083 19.3944
R9288 gnd.n1104 gnd.n1101 19.3944
R9289 gnd.n1107 gnd.n1104 19.3944
R9290 gnd.n1107 gnd.n1081 19.3944
R9291 gnd.n1111 gnd.n1081 19.3944
R9292 gnd.n1114 gnd.n1111 19.3944
R9293 gnd.n1117 gnd.n1114 19.3944
R9294 gnd.n1117 gnd.n1079 19.3944
R9295 gnd.n1121 gnd.n1079 19.3944
R9296 gnd.n1124 gnd.n1121 19.3944
R9297 gnd.n1127 gnd.n1124 19.3944
R9298 gnd.n1127 gnd.n1077 19.3944
R9299 gnd.n1131 gnd.n1077 19.3944
R9300 gnd.n1134 gnd.n1131 19.3944
R9301 gnd.n1137 gnd.n1134 19.3944
R9302 gnd.n1137 gnd.n1075 19.3944
R9303 gnd.n1141 gnd.n1075 19.3944
R9304 gnd.n1707 gnd.n1416 19.3944
R9305 gnd.n1717 gnd.n1416 19.3944
R9306 gnd.n1718 gnd.n1717 19.3944
R9307 gnd.n1718 gnd.n1397 19.3944
R9308 gnd.n1738 gnd.n1397 19.3944
R9309 gnd.n1738 gnd.n1389 19.3944
R9310 gnd.n1748 gnd.n1389 19.3944
R9311 gnd.n1749 gnd.n1748 19.3944
R9312 gnd.n1750 gnd.n1749 19.3944
R9313 gnd.n1750 gnd.n1372 19.3944
R9314 gnd.n1767 gnd.n1372 19.3944
R9315 gnd.n1770 gnd.n1767 19.3944
R9316 gnd.n1770 gnd.n1769 19.3944
R9317 gnd.n1769 gnd.n1345 19.3944
R9318 gnd.n1809 gnd.n1345 19.3944
R9319 gnd.n1809 gnd.n1342 19.3944
R9320 gnd.n1815 gnd.n1342 19.3944
R9321 gnd.n1816 gnd.n1815 19.3944
R9322 gnd.n1816 gnd.n1340 19.3944
R9323 gnd.n1822 gnd.n1340 19.3944
R9324 gnd.n1825 gnd.n1822 19.3944
R9325 gnd.n1827 gnd.n1825 19.3944
R9326 gnd.n1833 gnd.n1827 19.3944
R9327 gnd.n1833 gnd.n1832 19.3944
R9328 gnd.n1832 gnd.n1215 19.3944
R9329 gnd.n1899 gnd.n1215 19.3944
R9330 gnd.n1900 gnd.n1899 19.3944
R9331 gnd.n1900 gnd.n1208 19.3944
R9332 gnd.n1911 gnd.n1208 19.3944
R9333 gnd.n1912 gnd.n1911 19.3944
R9334 gnd.n1912 gnd.n1191 19.3944
R9335 gnd.n1191 gnd.n1189 19.3944
R9336 gnd.n1936 gnd.n1189 19.3944
R9337 gnd.n1939 gnd.n1936 19.3944
R9338 gnd.n1939 gnd.n1938 19.3944
R9339 gnd.n1938 gnd.n1161 19.3944
R9340 gnd.n2018 gnd.n1161 19.3944
R9341 gnd.n2018 gnd.n1158 19.3944
R9342 gnd.n2022 gnd.n1158 19.3944
R9343 gnd.n2023 gnd.n2022 19.3944
R9344 gnd.n2023 gnd.n1156 19.3944
R9345 gnd.n2029 gnd.n1156 19.3944
R9346 gnd.n2031 gnd.n2029 19.3944
R9347 gnd.n2035 gnd.n2031 19.3944
R9348 gnd.n2036 gnd.n2035 19.3944
R9349 gnd.n2036 gnd.n1153 19.3944
R9350 gnd.n2042 gnd.n1153 19.3944
R9351 gnd.n2300 gnd.n2042 19.3944
R9352 gnd.n2304 gnd.n2300 19.3944
R9353 gnd.n2305 gnd.n2304 19.3944
R9354 gnd.n2310 gnd.n2305 19.3944
R9355 gnd.n2310 gnd.n1049 19.3944
R9356 gnd.n6206 gnd.n1049 19.3944
R9357 gnd.n1698 gnd.n1697 19.3944
R9358 gnd.n1697 gnd.n1430 19.3944
R9359 gnd.n1453 gnd.n1430 19.3944
R9360 gnd.n1456 gnd.n1453 19.3944
R9361 gnd.n1456 gnd.n1449 19.3944
R9362 gnd.n1460 gnd.n1449 19.3944
R9363 gnd.n1463 gnd.n1460 19.3944
R9364 gnd.n1466 gnd.n1463 19.3944
R9365 gnd.n1466 gnd.n1447 19.3944
R9366 gnd.n1470 gnd.n1447 19.3944
R9367 gnd.n1473 gnd.n1470 19.3944
R9368 gnd.n1476 gnd.n1473 19.3944
R9369 gnd.n1476 gnd.n1445 19.3944
R9370 gnd.n1480 gnd.n1445 19.3944
R9371 gnd.n1703 gnd.n1702 19.3944
R9372 gnd.n1702 gnd.n1406 19.3944
R9373 gnd.n1728 gnd.n1406 19.3944
R9374 gnd.n1728 gnd.n1404 19.3944
R9375 gnd.n1734 gnd.n1404 19.3944
R9376 gnd.n1734 gnd.n1733 19.3944
R9377 gnd.n1733 gnd.n1378 19.3944
R9378 gnd.n1758 gnd.n1378 19.3944
R9379 gnd.n1758 gnd.n1376 19.3944
R9380 gnd.n1762 gnd.n1376 19.3944
R9381 gnd.n1762 gnd.n1356 19.3944
R9382 gnd.n1789 gnd.n1356 19.3944
R9383 gnd.n1789 gnd.n1354 19.3944
R9384 gnd.n1799 gnd.n1354 19.3944
R9385 gnd.n1799 gnd.n1798 19.3944
R9386 gnd.n1798 gnd.n1797 19.3944
R9387 gnd.n1797 gnd.n1303 19.3944
R9388 gnd.n1847 gnd.n1303 19.3944
R9389 gnd.n1847 gnd.n1846 19.3944
R9390 gnd.n1846 gnd.n1845 19.3944
R9391 gnd.n1845 gnd.n1307 19.3944
R9392 gnd.n1327 gnd.n1307 19.3944
R9393 gnd.n1327 gnd.n1225 19.3944
R9394 gnd.n1884 gnd.n1225 19.3944
R9395 gnd.n1884 gnd.n1223 19.3944
R9396 gnd.n1890 gnd.n1223 19.3944
R9397 gnd.n1890 gnd.n1889 19.3944
R9398 gnd.n1889 gnd.n1198 19.3944
R9399 gnd.n1924 gnd.n1198 19.3944
R9400 gnd.n1924 gnd.n1196 19.3944
R9401 gnd.n1930 gnd.n1196 19.3944
R9402 gnd.n1930 gnd.n1929 19.3944
R9403 gnd.n1929 gnd.n1172 19.3944
R9404 gnd.n1998 gnd.n1172 19.3944
R9405 gnd.n1998 gnd.n1170 19.3944
R9406 gnd.n2008 gnd.n1170 19.3944
R9407 gnd.n2008 gnd.n2007 19.3944
R9408 gnd.n2007 gnd.n2006 19.3944
R9409 gnd.n2006 gnd.n983 19.3944
R9410 gnd.n6244 gnd.n983 19.3944
R9411 gnd.n6244 gnd.n6243 19.3944
R9412 gnd.n6243 gnd.n6242 19.3944
R9413 gnd.n6242 gnd.n987 19.3944
R9414 gnd.n1007 gnd.n987 19.3944
R9415 gnd.n6230 gnd.n1007 19.3944
R9416 gnd.n6230 gnd.n6229 19.3944
R9417 gnd.n6229 gnd.n6228 19.3944
R9418 gnd.n6228 gnd.n1013 19.3944
R9419 gnd.n1032 gnd.n1013 19.3944
R9420 gnd.n6216 gnd.n1032 19.3944
R9421 gnd.n6216 gnd.n6215 19.3944
R9422 gnd.n6215 gnd.n6214 19.3944
R9423 gnd.n6214 gnd.n1038 19.3944
R9424 gnd.n6193 gnd.n6192 19.3944
R9425 gnd.n6192 gnd.n6158 19.3944
R9426 gnd.n6188 gnd.n6158 19.3944
R9427 gnd.n6188 gnd.n6185 19.3944
R9428 gnd.n6185 gnd.n6182 19.3944
R9429 gnd.n6182 gnd.n6181 19.3944
R9430 gnd.n6181 gnd.n6178 19.3944
R9431 gnd.n6178 gnd.n6177 19.3944
R9432 gnd.n6177 gnd.n6174 19.3944
R9433 gnd.n6174 gnd.n6173 19.3944
R9434 gnd.n6173 gnd.n6170 19.3944
R9435 gnd.n6170 gnd.n6169 19.3944
R9436 gnd.n6169 gnd.n1055 19.3944
R9437 gnd.n6199 gnd.n1055 19.3944
R9438 gnd.n1618 gnd.n1517 19.3944
R9439 gnd.n1618 gnd.n1508 19.3944
R9440 gnd.n1631 gnd.n1508 19.3944
R9441 gnd.n1631 gnd.n1506 19.3944
R9442 gnd.n1635 gnd.n1506 19.3944
R9443 gnd.n1635 gnd.n1496 19.3944
R9444 gnd.n1647 gnd.n1496 19.3944
R9445 gnd.n1647 gnd.n1494 19.3944
R9446 gnd.n1681 gnd.n1494 19.3944
R9447 gnd.n1681 gnd.n1680 19.3944
R9448 gnd.n1680 gnd.n1679 19.3944
R9449 gnd.n1679 gnd.n1678 19.3944
R9450 gnd.n1678 gnd.n1675 19.3944
R9451 gnd.n1675 gnd.n1674 19.3944
R9452 gnd.n1674 gnd.n1673 19.3944
R9453 gnd.n1673 gnd.n1671 19.3944
R9454 gnd.n1671 gnd.n1670 19.3944
R9455 gnd.n1670 gnd.n1667 19.3944
R9456 gnd.n1667 gnd.n1666 19.3944
R9457 gnd.n1666 gnd.n1665 19.3944
R9458 gnd.n1665 gnd.n1663 19.3944
R9459 gnd.n1663 gnd.n1362 19.3944
R9460 gnd.n1778 gnd.n1362 19.3944
R9461 gnd.n1778 gnd.n1360 19.3944
R9462 gnd.n1784 gnd.n1360 19.3944
R9463 gnd.n1784 gnd.n1783 19.3944
R9464 gnd.n1783 gnd.n1284 19.3944
R9465 gnd.n1858 gnd.n1284 19.3944
R9466 gnd.n1858 gnd.n1285 19.3944
R9467 gnd.n1332 gnd.n1331 19.3944
R9468 gnd.n1335 gnd.n1334 19.3944
R9469 gnd.n1322 gnd.n1321 19.3944
R9470 gnd.n1877 gnd.n1230 19.3944
R9471 gnd.n1877 gnd.n1876 19.3944
R9472 gnd.n1876 gnd.n1875 19.3944
R9473 gnd.n1875 gnd.n1873 19.3944
R9474 gnd.n1873 gnd.n1872 19.3944
R9475 gnd.n1872 gnd.n1870 19.3944
R9476 gnd.n1870 gnd.n1869 19.3944
R9477 gnd.n1869 gnd.n1179 19.3944
R9478 gnd.n1947 gnd.n1179 19.3944
R9479 gnd.n1947 gnd.n1177 19.3944
R9480 gnd.n1993 gnd.n1177 19.3944
R9481 gnd.n1993 gnd.n1992 19.3944
R9482 gnd.n1992 gnd.n1991 19.3944
R9483 gnd.n1991 gnd.n1989 19.3944
R9484 gnd.n1989 gnd.n1988 19.3944
R9485 gnd.n1988 gnd.n1985 19.3944
R9486 gnd.n1985 gnd.n1984 19.3944
R9487 gnd.n1984 gnd.n1981 19.3944
R9488 gnd.n1981 gnd.n1980 19.3944
R9489 gnd.n1980 gnd.n1979 19.3944
R9490 gnd.n1979 gnd.n1976 19.3944
R9491 gnd.n1976 gnd.n1975 19.3944
R9492 gnd.n1975 gnd.n1972 19.3944
R9493 gnd.n1972 gnd.n1971 19.3944
R9494 gnd.n1971 gnd.n1970 19.3944
R9495 gnd.n1970 gnd.n1967 19.3944
R9496 gnd.n1967 gnd.n1150 19.3944
R9497 gnd.n2316 gnd.n1150 19.3944
R9498 gnd.n2317 gnd.n2316 19.3944
R9499 gnd.n1623 gnd.n1513 19.3944
R9500 gnd.n1623 gnd.n1511 19.3944
R9501 gnd.n1627 gnd.n1511 19.3944
R9502 gnd.n1627 gnd.n1502 19.3944
R9503 gnd.n1639 gnd.n1502 19.3944
R9504 gnd.n1639 gnd.n1500 19.3944
R9505 gnd.n1643 gnd.n1500 19.3944
R9506 gnd.n1643 gnd.n1489 19.3944
R9507 gnd.n1685 gnd.n1489 19.3944
R9508 gnd.n1685 gnd.n1443 19.3944
R9509 gnd.n1691 gnd.n1443 19.3944
R9510 gnd.n1691 gnd.n1690 19.3944
R9511 gnd.n1690 gnd.n1421 19.3944
R9512 gnd.n1712 gnd.n1421 19.3944
R9513 gnd.n1712 gnd.n1414 19.3944
R9514 gnd.n1723 gnd.n1414 19.3944
R9515 gnd.n1723 gnd.n1722 19.3944
R9516 gnd.n1722 gnd.n1395 19.3944
R9517 gnd.n1743 gnd.n1395 19.3944
R9518 gnd.n1743 gnd.n1385 19.3944
R9519 gnd.n1753 gnd.n1385 19.3944
R9520 gnd.n1753 gnd.n1368 19.3944
R9521 gnd.n1774 gnd.n1368 19.3944
R9522 gnd.n1774 gnd.n1773 19.3944
R9523 gnd.n1773 gnd.n1347 19.3944
R9524 gnd.n1804 gnd.n1347 19.3944
R9525 gnd.n1804 gnd.n1292 19.3944
R9526 gnd.n1854 gnd.n1292 19.3944
R9527 gnd.n1854 gnd.n1853 19.3944
R9528 gnd.n1853 gnd.n1852 19.3944
R9529 gnd.n1852 gnd.n1296 19.3944
R9530 gnd.n1314 gnd.n1296 19.3944
R9531 gnd.n1840 gnd.n1314 19.3944
R9532 gnd.n1840 gnd.n1839 19.3944
R9533 gnd.n1839 gnd.n1838 19.3944
R9534 gnd.n1838 gnd.n1318 19.3944
R9535 gnd.n1318 gnd.n1217 19.3944
R9536 gnd.n1895 gnd.n1217 19.3944
R9537 gnd.n1895 gnd.n1210 19.3944
R9538 gnd.n1906 gnd.n1210 19.3944
R9539 gnd.n1906 gnd.n1206 19.3944
R9540 gnd.n1919 gnd.n1206 19.3944
R9541 gnd.n1919 gnd.n1918 19.3944
R9542 gnd.n1918 gnd.n1185 19.3944
R9543 gnd.n1943 gnd.n1185 19.3944
R9544 gnd.n1943 gnd.n1942 19.3944
R9545 gnd.n1942 gnd.n1163 19.3944
R9546 gnd.n2013 gnd.n1163 19.3944
R9547 gnd.n2013 gnd.n971 19.3944
R9548 gnd.n6251 gnd.n971 19.3944
R9549 gnd.n6251 gnd.n6250 19.3944
R9550 gnd.n6250 gnd.n6249 19.3944
R9551 gnd.n6249 gnd.n975 19.3944
R9552 gnd.n995 gnd.n975 19.3944
R9553 gnd.n6237 gnd.n995 19.3944
R9554 gnd.n6237 gnd.n6236 19.3944
R9555 gnd.n6236 gnd.n6235 19.3944
R9556 gnd.n6235 gnd.n999 19.3944
R9557 gnd.n1021 gnd.n999 19.3944
R9558 gnd.n6223 gnd.n1021 19.3944
R9559 gnd.n6223 gnd.n6222 19.3944
R9560 gnd.n6222 gnd.n6221 19.3944
R9561 gnd.n6221 gnd.n1025 19.3944
R9562 gnd.n1046 gnd.n1025 19.3944
R9563 gnd.n6209 gnd.n1046 19.3944
R9564 gnd.n5472 gnd.n3080 19.3944
R9565 gnd.n5477 gnd.n3080 19.3944
R9566 gnd.n5477 gnd.n3081 19.3944
R9567 gnd.n3081 gnd.n3007 19.3944
R9568 gnd.n5503 gnd.n3007 19.3944
R9569 gnd.n5503 gnd.n3004 19.3944
R9570 gnd.n5508 gnd.n3004 19.3944
R9571 gnd.n5508 gnd.n3005 19.3944
R9572 gnd.n3005 gnd.n2979 19.3944
R9573 gnd.n5534 gnd.n2979 19.3944
R9574 gnd.n5534 gnd.n2976 19.3944
R9575 gnd.n5539 gnd.n2976 19.3944
R9576 gnd.n5539 gnd.n2977 19.3944
R9577 gnd.n2977 gnd.n2951 19.3944
R9578 gnd.n5573 gnd.n2951 19.3944
R9579 gnd.n5573 gnd.n2948 19.3944
R9580 gnd.n5581 gnd.n2948 19.3944
R9581 gnd.n5581 gnd.n2949 19.3944
R9582 gnd.n5577 gnd.n2949 19.3944
R9583 gnd.n5577 gnd.n2940 19.3944
R9584 gnd.n5599 gnd.n2940 19.3944
R9585 gnd.n5599 gnd.n2937 19.3944
R9586 gnd.n5606 gnd.n2937 19.3944
R9587 gnd.n5606 gnd.n2938 19.3944
R9588 gnd.n5602 gnd.n2938 19.3944
R9589 gnd.n5602 gnd.n65 19.3944
R9590 gnd.n7482 gnd.n65 19.3944
R9591 gnd.n7482 gnd.n7481 19.3944
R9592 gnd.n7481 gnd.n7480 19.3944
R9593 gnd.n7480 gnd.n69 19.3944
R9594 gnd.n7476 gnd.n69 19.3944
R9595 gnd.n7476 gnd.n7475 19.3944
R9596 gnd.n7475 gnd.n7474 19.3944
R9597 gnd.n7474 gnd.n74 19.3944
R9598 gnd.n7470 gnd.n74 19.3944
R9599 gnd.n7470 gnd.n7469 19.3944
R9600 gnd.n7469 gnd.n7468 19.3944
R9601 gnd.n7468 gnd.n79 19.3944
R9602 gnd.n7464 gnd.n79 19.3944
R9603 gnd.n7464 gnd.n7463 19.3944
R9604 gnd.n7463 gnd.n7462 19.3944
R9605 gnd.n7462 gnd.n84 19.3944
R9606 gnd.n7458 gnd.n84 19.3944
R9607 gnd.n7458 gnd.n7457 19.3944
R9608 gnd.n7457 gnd.n7456 19.3944
R9609 gnd.n7456 gnd.n89 19.3944
R9610 gnd.n7452 gnd.n89 19.3944
R9611 gnd.n7452 gnd.n7451 19.3944
R9612 gnd.n7451 gnd.n7450 19.3944
R9613 gnd.n7450 gnd.n94 19.3944
R9614 gnd.n7446 gnd.n94 19.3944
R9615 gnd.n7446 gnd.n7445 19.3944
R9616 gnd.n7445 gnd.n7444 19.3944
R9617 gnd.n7343 gnd.n7342 19.3944
R9618 gnd.n7342 gnd.n7341 19.3944
R9619 gnd.n7341 gnd.n7283 19.3944
R9620 gnd.n7337 gnd.n7283 19.3944
R9621 gnd.n7337 gnd.n7336 19.3944
R9622 gnd.n7336 gnd.n7335 19.3944
R9623 gnd.n7335 gnd.n7291 19.3944
R9624 gnd.n7331 gnd.n7291 19.3944
R9625 gnd.n7331 gnd.n7330 19.3944
R9626 gnd.n7330 gnd.n7329 19.3944
R9627 gnd.n7329 gnd.n7299 19.3944
R9628 gnd.n7325 gnd.n7299 19.3944
R9629 gnd.n7325 gnd.n7324 19.3944
R9630 gnd.n7324 gnd.n7323 19.3944
R9631 gnd.n7323 gnd.n7307 19.3944
R9632 gnd.n7319 gnd.n7307 19.3944
R9633 gnd.n3129 gnd.n3126 19.3944
R9634 gnd.n3132 gnd.n3129 19.3944
R9635 gnd.n3132 gnd.n3120 19.3944
R9636 gnd.n3144 gnd.n3120 19.3944
R9637 gnd.n3145 gnd.n3144 19.3944
R9638 gnd.n3148 gnd.n3145 19.3944
R9639 gnd.n3148 gnd.n3111 19.3944
R9640 gnd.n3161 gnd.n3111 19.3944
R9641 gnd.n3162 gnd.n3161 19.3944
R9642 gnd.n3165 gnd.n3162 19.3944
R9643 gnd.n3165 gnd.n3102 19.3944
R9644 gnd.n3178 gnd.n3102 19.3944
R9645 gnd.n3179 gnd.n3178 19.3944
R9646 gnd.n3182 gnd.n3179 19.3944
R9647 gnd.n3182 gnd.n3093 19.3944
R9648 gnd.n3195 gnd.n3093 19.3944
R9649 gnd.n5692 gnd.n2877 19.3944
R9650 gnd.n5688 gnd.n2877 19.3944
R9651 gnd.n5688 gnd.n5687 19.3944
R9652 gnd.n5687 gnd.n5686 19.3944
R9653 gnd.n5686 gnd.n2883 19.3944
R9654 gnd.n5682 gnd.n2883 19.3944
R9655 gnd.n5682 gnd.n5681 19.3944
R9656 gnd.n5681 gnd.n5680 19.3944
R9657 gnd.n5680 gnd.n2888 19.3944
R9658 gnd.n5676 gnd.n2888 19.3944
R9659 gnd.n5676 gnd.n5675 19.3944
R9660 gnd.n5675 gnd.n5674 19.3944
R9661 gnd.n5674 gnd.n2893 19.3944
R9662 gnd.n5670 gnd.n2893 19.3944
R9663 gnd.n5670 gnd.n5669 19.3944
R9664 gnd.n5669 gnd.n5668 19.3944
R9665 gnd.n5668 gnd.n2898 19.3944
R9666 gnd.n5664 gnd.n2898 19.3944
R9667 gnd.n5664 gnd.n5663 19.3944
R9668 gnd.n5663 gnd.n5662 19.3944
R9669 gnd.n5662 gnd.n279 19.3944
R9670 gnd.n7198 gnd.n279 19.3944
R9671 gnd.n7198 gnd.n280 19.3944
R9672 gnd.n7194 gnd.n280 19.3944
R9673 gnd.n7194 gnd.n7193 19.3944
R9674 gnd.n7193 gnd.n7192 19.3944
R9675 gnd.n7192 gnd.n286 19.3944
R9676 gnd.n7187 gnd.n286 19.3944
R9677 gnd.n7187 gnd.n7186 19.3944
R9678 gnd.n7186 gnd.n257 19.3944
R9679 gnd.n7209 gnd.n257 19.3944
R9680 gnd.n7209 gnd.n255 19.3944
R9681 gnd.n7213 gnd.n255 19.3944
R9682 gnd.n7213 gnd.n242 19.3944
R9683 gnd.n7225 gnd.n242 19.3944
R9684 gnd.n7225 gnd.n240 19.3944
R9685 gnd.n7229 gnd.n240 19.3944
R9686 gnd.n7229 gnd.n227 19.3944
R9687 gnd.n7241 gnd.n227 19.3944
R9688 gnd.n7241 gnd.n225 19.3944
R9689 gnd.n7245 gnd.n225 19.3944
R9690 gnd.n7245 gnd.n212 19.3944
R9691 gnd.n7257 gnd.n212 19.3944
R9692 gnd.n7257 gnd.n210 19.3944
R9693 gnd.n7261 gnd.n210 19.3944
R9694 gnd.n7261 gnd.n197 19.3944
R9695 gnd.n7273 gnd.n197 19.3944
R9696 gnd.n7273 gnd.n194 19.3944
R9697 gnd.n7352 gnd.n194 19.3944
R9698 gnd.n7352 gnd.n195 19.3944
R9699 gnd.n7348 gnd.n195 19.3944
R9700 gnd.n7348 gnd.n7347 19.3944
R9701 gnd.n7347 gnd.n7346 19.3944
R9702 gnd.n3603 gnd.n2675 19.3944
R9703 gnd.n3606 gnd.n3603 19.3944
R9704 gnd.n3606 gnd.n3597 19.3944
R9705 gnd.n3615 gnd.n3597 19.3944
R9706 gnd.n3618 gnd.n3615 19.3944
R9707 gnd.n3618 gnd.n3589 19.3944
R9708 gnd.n3627 gnd.n3589 19.3944
R9709 gnd.n3630 gnd.n3627 19.3944
R9710 gnd.n3630 gnd.n3585 19.3944
R9711 gnd.n3639 gnd.n3585 19.3944
R9712 gnd.n3642 gnd.n3639 19.3944
R9713 gnd.n3642 gnd.n3577 19.3944
R9714 gnd.n3651 gnd.n3577 19.3944
R9715 gnd.n3653 gnd.n3651 19.3944
R9716 gnd.n3653 gnd.n3573 19.3944
R9717 gnd.n3663 gnd.n3573 19.3944
R9718 gnd.n6911 gnd.n504 19.3944
R9719 gnd.n6917 gnd.n504 19.3944
R9720 gnd.n6917 gnd.n502 19.3944
R9721 gnd.n6921 gnd.n502 19.3944
R9722 gnd.n6921 gnd.n498 19.3944
R9723 gnd.n6927 gnd.n498 19.3944
R9724 gnd.n6927 gnd.n496 19.3944
R9725 gnd.n6931 gnd.n496 19.3944
R9726 gnd.n6931 gnd.n492 19.3944
R9727 gnd.n6937 gnd.n492 19.3944
R9728 gnd.n6937 gnd.n490 19.3944
R9729 gnd.n6941 gnd.n490 19.3944
R9730 gnd.n6941 gnd.n486 19.3944
R9731 gnd.n6947 gnd.n486 19.3944
R9732 gnd.n6947 gnd.n484 19.3944
R9733 gnd.n6951 gnd.n484 19.3944
R9734 gnd.n6951 gnd.n480 19.3944
R9735 gnd.n6957 gnd.n480 19.3944
R9736 gnd.n6957 gnd.n478 19.3944
R9737 gnd.n6961 gnd.n478 19.3944
R9738 gnd.n6961 gnd.n474 19.3944
R9739 gnd.n6967 gnd.n474 19.3944
R9740 gnd.n6967 gnd.n472 19.3944
R9741 gnd.n6971 gnd.n472 19.3944
R9742 gnd.n6971 gnd.n468 19.3944
R9743 gnd.n6977 gnd.n468 19.3944
R9744 gnd.n6977 gnd.n466 19.3944
R9745 gnd.n6981 gnd.n466 19.3944
R9746 gnd.n6981 gnd.n462 19.3944
R9747 gnd.n6987 gnd.n462 19.3944
R9748 gnd.n6987 gnd.n460 19.3944
R9749 gnd.n6991 gnd.n460 19.3944
R9750 gnd.n6991 gnd.n456 19.3944
R9751 gnd.n6997 gnd.n456 19.3944
R9752 gnd.n6997 gnd.n454 19.3944
R9753 gnd.n7001 gnd.n454 19.3944
R9754 gnd.n7001 gnd.n450 19.3944
R9755 gnd.n7007 gnd.n450 19.3944
R9756 gnd.n7007 gnd.n448 19.3944
R9757 gnd.n7011 gnd.n448 19.3944
R9758 gnd.n7011 gnd.n444 19.3944
R9759 gnd.n7017 gnd.n444 19.3944
R9760 gnd.n7017 gnd.n442 19.3944
R9761 gnd.n7021 gnd.n442 19.3944
R9762 gnd.n7021 gnd.n438 19.3944
R9763 gnd.n7027 gnd.n438 19.3944
R9764 gnd.n7027 gnd.n436 19.3944
R9765 gnd.n7031 gnd.n436 19.3944
R9766 gnd.n7031 gnd.n432 19.3944
R9767 gnd.n7037 gnd.n432 19.3944
R9768 gnd.n7037 gnd.n430 19.3944
R9769 gnd.n7041 gnd.n430 19.3944
R9770 gnd.n7041 gnd.n426 19.3944
R9771 gnd.n7047 gnd.n426 19.3944
R9772 gnd.n7047 gnd.n424 19.3944
R9773 gnd.n7051 gnd.n424 19.3944
R9774 gnd.n7051 gnd.n420 19.3944
R9775 gnd.n7057 gnd.n420 19.3944
R9776 gnd.n7057 gnd.n418 19.3944
R9777 gnd.n7061 gnd.n418 19.3944
R9778 gnd.n7061 gnd.n414 19.3944
R9779 gnd.n7067 gnd.n414 19.3944
R9780 gnd.n7067 gnd.n412 19.3944
R9781 gnd.n7071 gnd.n412 19.3944
R9782 gnd.n7071 gnd.n408 19.3944
R9783 gnd.n7077 gnd.n408 19.3944
R9784 gnd.n7077 gnd.n406 19.3944
R9785 gnd.n7081 gnd.n406 19.3944
R9786 gnd.n7081 gnd.n402 19.3944
R9787 gnd.n7087 gnd.n402 19.3944
R9788 gnd.n7087 gnd.n400 19.3944
R9789 gnd.n7091 gnd.n400 19.3944
R9790 gnd.n7091 gnd.n396 19.3944
R9791 gnd.n7097 gnd.n396 19.3944
R9792 gnd.n7097 gnd.n394 19.3944
R9793 gnd.n7101 gnd.n394 19.3944
R9794 gnd.n7101 gnd.n390 19.3944
R9795 gnd.n7107 gnd.n390 19.3944
R9796 gnd.n7107 gnd.n388 19.3944
R9797 gnd.n7111 gnd.n388 19.3944
R9798 gnd.n7111 gnd.n384 19.3944
R9799 gnd.n7118 gnd.n384 19.3944
R9800 gnd.n7118 gnd.n382 19.3944
R9801 gnd.n7123 gnd.n382 19.3944
R9802 gnd.n6426 gnd.n797 19.3944
R9803 gnd.n6426 gnd.n795 19.3944
R9804 gnd.n6430 gnd.n795 19.3944
R9805 gnd.n6430 gnd.n791 19.3944
R9806 gnd.n6436 gnd.n791 19.3944
R9807 gnd.n6436 gnd.n789 19.3944
R9808 gnd.n6440 gnd.n789 19.3944
R9809 gnd.n6440 gnd.n785 19.3944
R9810 gnd.n6446 gnd.n785 19.3944
R9811 gnd.n6446 gnd.n783 19.3944
R9812 gnd.n6450 gnd.n783 19.3944
R9813 gnd.n6450 gnd.n779 19.3944
R9814 gnd.n6456 gnd.n779 19.3944
R9815 gnd.n6456 gnd.n777 19.3944
R9816 gnd.n6460 gnd.n777 19.3944
R9817 gnd.n6460 gnd.n773 19.3944
R9818 gnd.n6466 gnd.n773 19.3944
R9819 gnd.n6466 gnd.n771 19.3944
R9820 gnd.n6470 gnd.n771 19.3944
R9821 gnd.n6470 gnd.n767 19.3944
R9822 gnd.n6476 gnd.n767 19.3944
R9823 gnd.n6476 gnd.n765 19.3944
R9824 gnd.n6480 gnd.n765 19.3944
R9825 gnd.n6480 gnd.n761 19.3944
R9826 gnd.n6486 gnd.n761 19.3944
R9827 gnd.n6486 gnd.n759 19.3944
R9828 gnd.n6490 gnd.n759 19.3944
R9829 gnd.n6490 gnd.n755 19.3944
R9830 gnd.n6496 gnd.n755 19.3944
R9831 gnd.n6496 gnd.n753 19.3944
R9832 gnd.n6500 gnd.n753 19.3944
R9833 gnd.n6500 gnd.n749 19.3944
R9834 gnd.n6506 gnd.n749 19.3944
R9835 gnd.n6506 gnd.n747 19.3944
R9836 gnd.n6510 gnd.n747 19.3944
R9837 gnd.n6510 gnd.n743 19.3944
R9838 gnd.n6516 gnd.n743 19.3944
R9839 gnd.n6516 gnd.n741 19.3944
R9840 gnd.n6520 gnd.n741 19.3944
R9841 gnd.n6520 gnd.n737 19.3944
R9842 gnd.n6526 gnd.n737 19.3944
R9843 gnd.n6526 gnd.n735 19.3944
R9844 gnd.n6530 gnd.n735 19.3944
R9845 gnd.n6530 gnd.n731 19.3944
R9846 gnd.n6536 gnd.n731 19.3944
R9847 gnd.n6536 gnd.n729 19.3944
R9848 gnd.n6540 gnd.n729 19.3944
R9849 gnd.n6540 gnd.n725 19.3944
R9850 gnd.n6546 gnd.n725 19.3944
R9851 gnd.n6546 gnd.n723 19.3944
R9852 gnd.n6550 gnd.n723 19.3944
R9853 gnd.n6550 gnd.n719 19.3944
R9854 gnd.n6556 gnd.n719 19.3944
R9855 gnd.n6556 gnd.n717 19.3944
R9856 gnd.n6560 gnd.n717 19.3944
R9857 gnd.n6560 gnd.n713 19.3944
R9858 gnd.n6566 gnd.n713 19.3944
R9859 gnd.n6566 gnd.n711 19.3944
R9860 gnd.n6570 gnd.n711 19.3944
R9861 gnd.n6570 gnd.n707 19.3944
R9862 gnd.n6576 gnd.n707 19.3944
R9863 gnd.n6576 gnd.n705 19.3944
R9864 gnd.n6580 gnd.n705 19.3944
R9865 gnd.n6580 gnd.n701 19.3944
R9866 gnd.n6586 gnd.n701 19.3944
R9867 gnd.n6586 gnd.n699 19.3944
R9868 gnd.n6590 gnd.n699 19.3944
R9869 gnd.n6590 gnd.n695 19.3944
R9870 gnd.n6596 gnd.n695 19.3944
R9871 gnd.n6596 gnd.n693 19.3944
R9872 gnd.n6600 gnd.n693 19.3944
R9873 gnd.n6600 gnd.n689 19.3944
R9874 gnd.n6606 gnd.n689 19.3944
R9875 gnd.n6606 gnd.n687 19.3944
R9876 gnd.n6610 gnd.n687 19.3944
R9877 gnd.n6610 gnd.n683 19.3944
R9878 gnd.n6616 gnd.n683 19.3944
R9879 gnd.n6616 gnd.n681 19.3944
R9880 gnd.n6620 gnd.n681 19.3944
R9881 gnd.n6620 gnd.n677 19.3944
R9882 gnd.n6626 gnd.n677 19.3944
R9883 gnd.n6626 gnd.n675 19.3944
R9884 gnd.n6630 gnd.n675 19.3944
R9885 gnd.n6630 gnd.n671 19.3944
R9886 gnd.n6636 gnd.n671 19.3944
R9887 gnd.n6636 gnd.n669 19.3944
R9888 gnd.n6640 gnd.n669 19.3944
R9889 gnd.n6640 gnd.n665 19.3944
R9890 gnd.n6646 gnd.n665 19.3944
R9891 gnd.n6646 gnd.n663 19.3944
R9892 gnd.n6650 gnd.n663 19.3944
R9893 gnd.n6650 gnd.n659 19.3944
R9894 gnd.n6656 gnd.n659 19.3944
R9895 gnd.n6656 gnd.n657 19.3944
R9896 gnd.n6660 gnd.n657 19.3944
R9897 gnd.n6660 gnd.n653 19.3944
R9898 gnd.n6666 gnd.n653 19.3944
R9899 gnd.n6666 gnd.n651 19.3944
R9900 gnd.n6670 gnd.n651 19.3944
R9901 gnd.n6670 gnd.n647 19.3944
R9902 gnd.n6676 gnd.n647 19.3944
R9903 gnd.n6676 gnd.n645 19.3944
R9904 gnd.n6680 gnd.n645 19.3944
R9905 gnd.n6680 gnd.n641 19.3944
R9906 gnd.n6686 gnd.n641 19.3944
R9907 gnd.n6686 gnd.n639 19.3944
R9908 gnd.n6690 gnd.n639 19.3944
R9909 gnd.n6690 gnd.n635 19.3944
R9910 gnd.n6696 gnd.n635 19.3944
R9911 gnd.n6696 gnd.n633 19.3944
R9912 gnd.n6700 gnd.n633 19.3944
R9913 gnd.n6700 gnd.n629 19.3944
R9914 gnd.n6706 gnd.n629 19.3944
R9915 gnd.n6706 gnd.n627 19.3944
R9916 gnd.n6710 gnd.n627 19.3944
R9917 gnd.n6710 gnd.n623 19.3944
R9918 gnd.n6716 gnd.n623 19.3944
R9919 gnd.n6716 gnd.n621 19.3944
R9920 gnd.n6720 gnd.n621 19.3944
R9921 gnd.n6720 gnd.n617 19.3944
R9922 gnd.n6726 gnd.n617 19.3944
R9923 gnd.n6726 gnd.n615 19.3944
R9924 gnd.n6730 gnd.n615 19.3944
R9925 gnd.n6730 gnd.n611 19.3944
R9926 gnd.n6736 gnd.n611 19.3944
R9927 gnd.n6736 gnd.n609 19.3944
R9928 gnd.n6740 gnd.n609 19.3944
R9929 gnd.n6740 gnd.n605 19.3944
R9930 gnd.n6746 gnd.n605 19.3944
R9931 gnd.n6746 gnd.n603 19.3944
R9932 gnd.n6750 gnd.n603 19.3944
R9933 gnd.n6750 gnd.n599 19.3944
R9934 gnd.n6756 gnd.n599 19.3944
R9935 gnd.n6756 gnd.n597 19.3944
R9936 gnd.n6760 gnd.n597 19.3944
R9937 gnd.n6760 gnd.n593 19.3944
R9938 gnd.n6766 gnd.n593 19.3944
R9939 gnd.n6766 gnd.n591 19.3944
R9940 gnd.n6770 gnd.n591 19.3944
R9941 gnd.n6770 gnd.n587 19.3944
R9942 gnd.n6776 gnd.n587 19.3944
R9943 gnd.n6776 gnd.n585 19.3944
R9944 gnd.n6780 gnd.n585 19.3944
R9945 gnd.n6780 gnd.n581 19.3944
R9946 gnd.n6786 gnd.n581 19.3944
R9947 gnd.n6786 gnd.n579 19.3944
R9948 gnd.n6790 gnd.n579 19.3944
R9949 gnd.n6790 gnd.n575 19.3944
R9950 gnd.n6796 gnd.n575 19.3944
R9951 gnd.n6796 gnd.n573 19.3944
R9952 gnd.n6800 gnd.n573 19.3944
R9953 gnd.n6800 gnd.n569 19.3944
R9954 gnd.n6806 gnd.n569 19.3944
R9955 gnd.n6806 gnd.n567 19.3944
R9956 gnd.n6810 gnd.n567 19.3944
R9957 gnd.n6810 gnd.n563 19.3944
R9958 gnd.n6816 gnd.n563 19.3944
R9959 gnd.n6816 gnd.n561 19.3944
R9960 gnd.n6820 gnd.n561 19.3944
R9961 gnd.n6820 gnd.n557 19.3944
R9962 gnd.n6826 gnd.n557 19.3944
R9963 gnd.n6826 gnd.n555 19.3944
R9964 gnd.n6830 gnd.n555 19.3944
R9965 gnd.n6830 gnd.n551 19.3944
R9966 gnd.n6836 gnd.n551 19.3944
R9967 gnd.n6836 gnd.n549 19.3944
R9968 gnd.n6840 gnd.n549 19.3944
R9969 gnd.n6840 gnd.n545 19.3944
R9970 gnd.n6846 gnd.n545 19.3944
R9971 gnd.n6846 gnd.n543 19.3944
R9972 gnd.n6850 gnd.n543 19.3944
R9973 gnd.n6850 gnd.n539 19.3944
R9974 gnd.n6856 gnd.n539 19.3944
R9975 gnd.n6856 gnd.n537 19.3944
R9976 gnd.n6860 gnd.n537 19.3944
R9977 gnd.n6860 gnd.n533 19.3944
R9978 gnd.n6866 gnd.n533 19.3944
R9979 gnd.n6866 gnd.n531 19.3944
R9980 gnd.n6870 gnd.n531 19.3944
R9981 gnd.n6870 gnd.n527 19.3944
R9982 gnd.n6876 gnd.n527 19.3944
R9983 gnd.n6876 gnd.n525 19.3944
R9984 gnd.n6880 gnd.n525 19.3944
R9985 gnd.n6880 gnd.n521 19.3944
R9986 gnd.n6886 gnd.n521 19.3944
R9987 gnd.n6886 gnd.n519 19.3944
R9988 gnd.n6890 gnd.n519 19.3944
R9989 gnd.n6890 gnd.n515 19.3944
R9990 gnd.n6896 gnd.n515 19.3944
R9991 gnd.n6896 gnd.n513 19.3944
R9992 gnd.n6901 gnd.n513 19.3944
R9993 gnd.n6901 gnd.n509 19.3944
R9994 gnd.n6907 gnd.n509 19.3944
R9995 gnd.n6908 gnd.n6907 19.3944
R9996 gnd.n5767 gnd.n5766 19.3944
R9997 gnd.n5766 gnd.n5765 19.3944
R9998 gnd.n5765 gnd.n5764 19.3944
R9999 gnd.n5764 gnd.n5762 19.3944
R10000 gnd.n5762 gnd.n5759 19.3944
R10001 gnd.n5759 gnd.n5758 19.3944
R10002 gnd.n5758 gnd.n5755 19.3944
R10003 gnd.n5755 gnd.n5754 19.3944
R10004 gnd.n5754 gnd.n5751 19.3944
R10005 gnd.n5751 gnd.n5750 19.3944
R10006 gnd.n5750 gnd.n5747 19.3944
R10007 gnd.n5747 gnd.n5746 19.3944
R10008 gnd.n5746 gnd.n5743 19.3944
R10009 gnd.n5743 gnd.n5742 19.3944
R10010 gnd.n5742 gnd.n5739 19.3944
R10011 gnd.n5737 gnd.n5734 19.3944
R10012 gnd.n5734 gnd.n5733 19.3944
R10013 gnd.n5733 gnd.n5730 19.3944
R10014 gnd.n5730 gnd.n5729 19.3944
R10015 gnd.n5729 gnd.n5726 19.3944
R10016 gnd.n5726 gnd.n5725 19.3944
R10017 gnd.n5725 gnd.n5722 19.3944
R10018 gnd.n5722 gnd.n5721 19.3944
R10019 gnd.n5721 gnd.n5718 19.3944
R10020 gnd.n5718 gnd.n5717 19.3944
R10021 gnd.n5717 gnd.n5714 19.3944
R10022 gnd.n5714 gnd.n5713 19.3944
R10023 gnd.n5713 gnd.n5710 19.3944
R10024 gnd.n5710 gnd.n5709 19.3944
R10025 gnd.n5709 gnd.n5706 19.3944
R10026 gnd.n5706 gnd.n5705 19.3944
R10027 gnd.n5705 gnd.n5702 19.3944
R10028 gnd.n5702 gnd.n5701 19.3944
R10029 gnd.n3042 gnd.n2871 19.3944
R10030 gnd.n3077 gnd.n3042 19.3944
R10031 gnd.n3077 gnd.n3076 19.3944
R10032 gnd.n3076 gnd.n3075 19.3944
R10033 gnd.n3075 gnd.n3073 19.3944
R10034 gnd.n3073 gnd.n3072 19.3944
R10035 gnd.n3072 gnd.n3070 19.3944
R10036 gnd.n3070 gnd.n3069 19.3944
R10037 gnd.n3069 gnd.n3068 19.3944
R10038 gnd.n3068 gnd.n3066 19.3944
R10039 gnd.n3066 gnd.n3065 19.3944
R10040 gnd.n3065 gnd.n3063 19.3944
R10041 gnd.n3063 gnd.n3062 19.3944
R10042 gnd.n3062 gnd.n3061 19.3944
R10043 gnd.n3061 gnd.n3059 19.3944
R10044 gnd.n3059 gnd.n2943 19.3944
R10045 gnd.n5586 gnd.n2943 19.3944
R10046 gnd.n5587 gnd.n5586 19.3944
R10047 gnd.n5589 gnd.n5587 19.3944
R10048 gnd.n5589 gnd.n2941 19.3944
R10049 gnd.n5595 gnd.n2941 19.3944
R10050 gnd.n5595 gnd.n5594 19.3944
R10051 gnd.n5594 gnd.n2935 19.3944
R10052 gnd.n5612 gnd.n2935 19.3944
R10053 gnd.n5612 gnd.n2933 19.3944
R10054 gnd.n5616 gnd.n2933 19.3944
R10055 gnd.n5616 gnd.n295 19.3944
R10056 gnd.n7177 gnd.n295 19.3944
R10057 gnd.n7177 gnd.n7176 19.3944
R10058 gnd.n7176 gnd.n7175 19.3944
R10059 gnd.n7175 gnd.n300 19.3944
R10060 gnd.n312 gnd.n300 19.3944
R10061 gnd.n312 gnd.n308 19.3944
R10062 gnd.n7160 gnd.n308 19.3944
R10063 gnd.n7160 gnd.n7159 19.3944
R10064 gnd.n7159 gnd.n7158 19.3944
R10065 gnd.n7158 gnd.n7155 19.3944
R10066 gnd.n7155 gnd.n7154 19.3944
R10067 gnd.n7154 gnd.n320 19.3944
R10068 gnd.n344 gnd.n320 19.3944
R10069 gnd.n344 gnd.n340 19.3944
R10070 gnd.n7140 gnd.n340 19.3944
R10071 gnd.n7140 gnd.n7139 19.3944
R10072 gnd.n7139 gnd.n7138 19.3944
R10073 gnd.n7138 gnd.n7135 19.3944
R10074 gnd.n7135 gnd.n7134 19.3944
R10075 gnd.n7134 gnd.n362 19.3944
R10076 gnd.n362 gnd.n361 19.3944
R10077 gnd.n361 gnd.n358 19.3944
R10078 gnd.n358 gnd.n357 19.3944
R10079 gnd.n357 gnd.n178 19.3944
R10080 gnd.n7365 gnd.n178 19.3944
R10081 gnd.n7366 gnd.n7365 19.3944
R10082 gnd.n7404 gnd.n139 19.3944
R10083 gnd.n7399 gnd.n139 19.3944
R10084 gnd.n7399 gnd.n7398 19.3944
R10085 gnd.n7398 gnd.n7397 19.3944
R10086 gnd.n7397 gnd.n146 19.3944
R10087 gnd.n7392 gnd.n146 19.3944
R10088 gnd.n7392 gnd.n7391 19.3944
R10089 gnd.n7391 gnd.n7390 19.3944
R10090 gnd.n7390 gnd.n153 19.3944
R10091 gnd.n7385 gnd.n153 19.3944
R10092 gnd.n7385 gnd.n7384 19.3944
R10093 gnd.n7384 gnd.n7383 19.3944
R10094 gnd.n7383 gnd.n160 19.3944
R10095 gnd.n7378 gnd.n160 19.3944
R10096 gnd.n7378 gnd.n7377 19.3944
R10097 gnd.n7377 gnd.n7376 19.3944
R10098 gnd.n7376 gnd.n167 19.3944
R10099 gnd.n7371 gnd.n167 19.3944
R10100 gnd.n7437 gnd.n7436 19.3944
R10101 gnd.n7436 gnd.n7435 19.3944
R10102 gnd.n7435 gnd.n111 19.3944
R10103 gnd.n7430 gnd.n111 19.3944
R10104 gnd.n7430 gnd.n7429 19.3944
R10105 gnd.n7429 gnd.n7428 19.3944
R10106 gnd.n7428 gnd.n118 19.3944
R10107 gnd.n7423 gnd.n118 19.3944
R10108 gnd.n7423 gnd.n7422 19.3944
R10109 gnd.n7422 gnd.n7421 19.3944
R10110 gnd.n7421 gnd.n125 19.3944
R10111 gnd.n7416 gnd.n125 19.3944
R10112 gnd.n7416 gnd.n7415 19.3944
R10113 gnd.n7415 gnd.n7414 19.3944
R10114 gnd.n7414 gnd.n132 19.3944
R10115 gnd.n7409 gnd.n132 19.3944
R10116 gnd.n7409 gnd.n7408 19.3944
R10117 gnd.n3039 gnd.n3036 19.3944
R10118 gnd.n3039 gnd.n3017 19.3944
R10119 gnd.n5493 gnd.n3017 19.3944
R10120 gnd.n5493 gnd.n3015 19.3944
R10121 gnd.n5499 gnd.n3015 19.3944
R10122 gnd.n5499 gnd.n5498 19.3944
R10123 gnd.n5498 gnd.n2988 19.3944
R10124 gnd.n5524 gnd.n2988 19.3944
R10125 gnd.n5524 gnd.n2986 19.3944
R10126 gnd.n5530 gnd.n2986 19.3944
R10127 gnd.n5530 gnd.n5529 19.3944
R10128 gnd.n5529 gnd.n2960 19.3944
R10129 gnd.n5563 gnd.n2960 19.3944
R10130 gnd.n5563 gnd.n2958 19.3944
R10131 gnd.n5569 gnd.n2958 19.3944
R10132 gnd.n5569 gnd.n5568 19.3944
R10133 gnd.n5568 gnd.n2908 19.3944
R10134 gnd.n5653 gnd.n2908 19.3944
R10135 gnd.n5653 gnd.n2906 19.3944
R10136 gnd.n5657 gnd.n2906 19.3944
R10137 gnd.n5657 gnd.n270 19.3944
R10138 gnd.n7202 gnd.n270 19.3944
R10139 gnd.n269 gnd.n268 19.3944
R10140 gnd.n5634 gnd.n268 19.3944
R10141 gnd.n2931 gnd.n2930 19.3944
R10142 gnd.n7182 gnd.n7181 19.3944
R10143 gnd.n7205 gnd.n262 19.3944
R10144 gnd.n7205 gnd.n250 19.3944
R10145 gnd.n7217 gnd.n250 19.3944
R10146 gnd.n7217 gnd.n248 19.3944
R10147 gnd.n7221 gnd.n248 19.3944
R10148 gnd.n7221 gnd.n234 19.3944
R10149 gnd.n7233 gnd.n234 19.3944
R10150 gnd.n7233 gnd.n232 19.3944
R10151 gnd.n7237 gnd.n232 19.3944
R10152 gnd.n7237 gnd.n220 19.3944
R10153 gnd.n7249 gnd.n220 19.3944
R10154 gnd.n7249 gnd.n218 19.3944
R10155 gnd.n7253 gnd.n218 19.3944
R10156 gnd.n7253 gnd.n204 19.3944
R10157 gnd.n7265 gnd.n204 19.3944
R10158 gnd.n7265 gnd.n202 19.3944
R10159 gnd.n7269 gnd.n202 19.3944
R10160 gnd.n7269 gnd.n187 19.3944
R10161 gnd.n7356 gnd.n187 19.3944
R10162 gnd.n7356 gnd.n185 19.3944
R10163 gnd.n7360 gnd.n185 19.3944
R10164 gnd.n7360 gnd.n106 19.3944
R10165 gnd.n7440 gnd.n106 19.3944
R10166 gnd.n3968 gnd.n3967 19.3944
R10167 gnd.n3967 gnd.n3814 19.3944
R10168 gnd.n3963 gnd.n3814 19.3944
R10169 gnd.n3963 gnd.n3962 19.3944
R10170 gnd.n3962 gnd.n3961 19.3944
R10171 gnd.n3961 gnd.n3820 19.3944
R10172 gnd.n3957 gnd.n3820 19.3944
R10173 gnd.n3957 gnd.n3956 19.3944
R10174 gnd.n3956 gnd.n3955 19.3944
R10175 gnd.n3955 gnd.n3826 19.3944
R10176 gnd.n3951 gnd.n3826 19.3944
R10177 gnd.n3951 gnd.n3950 19.3944
R10178 gnd.n3950 gnd.n3949 19.3944
R10179 gnd.n3949 gnd.n3832 19.3944
R10180 gnd.n3945 gnd.n3832 19.3944
R10181 gnd.n3945 gnd.n3944 19.3944
R10182 gnd.n3944 gnd.n3943 19.3944
R10183 gnd.n3943 gnd.n3838 19.3944
R10184 gnd.n3939 gnd.n3938 19.3944
R10185 gnd.n3934 gnd.n3841 19.3944
R10186 gnd.n3930 gnd.n3845 19.3944
R10187 gnd.n3928 gnd.n3927 19.3944
R10188 gnd.n3924 gnd.n3923 19.3944
R10189 gnd.n3923 gnd.n3922 19.3944
R10190 gnd.n3922 gnd.n3849 19.3944
R10191 gnd.n3918 gnd.n3849 19.3944
R10192 gnd.n3918 gnd.n3917 19.3944
R10193 gnd.n3917 gnd.n3916 19.3944
R10194 gnd.n3916 gnd.n3855 19.3944
R10195 gnd.n3912 gnd.n3855 19.3944
R10196 gnd.n3912 gnd.n3911 19.3944
R10197 gnd.n3911 gnd.n3910 19.3944
R10198 gnd.n3910 gnd.n3861 19.3944
R10199 gnd.n3906 gnd.n3861 19.3944
R10200 gnd.n3906 gnd.n3905 19.3944
R10201 gnd.n3905 gnd.n3904 19.3944
R10202 gnd.n3904 gnd.n3867 19.3944
R10203 gnd.n3900 gnd.n3867 19.3944
R10204 gnd.n3900 gnd.n3899 19.3944
R10205 gnd.n3899 gnd.n3898 19.3944
R10206 gnd.n3898 gnd.n3873 19.3944
R10207 gnd.n3894 gnd.n3873 19.3944
R10208 gnd.n3894 gnd.n3893 19.3944
R10209 gnd.n3893 gnd.n3892 19.3944
R10210 gnd.n3892 gnd.n3879 19.3944
R10211 gnd.n3888 gnd.n3879 19.3944
R10212 gnd.n3888 gnd.n3887 19.3944
R10213 gnd.n3887 gnd.n3886 19.3944
R10214 gnd.n3886 gnd.n3525 19.3944
R10215 gnd.n4627 gnd.n3525 19.3944
R10216 gnd.n4627 gnd.n3523 19.3944
R10217 gnd.n4631 gnd.n3523 19.3944
R10218 gnd.n4631 gnd.n3512 19.3944
R10219 gnd.n4643 gnd.n3512 19.3944
R10220 gnd.n4643 gnd.n3510 19.3944
R10221 gnd.n4647 gnd.n3510 19.3944
R10222 gnd.n4647 gnd.n3499 19.3944
R10223 gnd.n4659 gnd.n3499 19.3944
R10224 gnd.n4659 gnd.n3497 19.3944
R10225 gnd.n4663 gnd.n3497 19.3944
R10226 gnd.n4663 gnd.n3485 19.3944
R10227 gnd.n4675 gnd.n3485 19.3944
R10228 gnd.n4675 gnd.n3483 19.3944
R10229 gnd.n4679 gnd.n3483 19.3944
R10230 gnd.n4679 gnd.n3471 19.3944
R10231 gnd.n4691 gnd.n3471 19.3944
R10232 gnd.n4691 gnd.n3469 19.3944
R10233 gnd.n4695 gnd.n3469 19.3944
R10234 gnd.n4695 gnd.n3458 19.3944
R10235 gnd.n4707 gnd.n3458 19.3944
R10236 gnd.n4707 gnd.n3456 19.3944
R10237 gnd.n4713 gnd.n3456 19.3944
R10238 gnd.n4713 gnd.n4712 19.3944
R10239 gnd.n4712 gnd.n3429 19.3944
R10240 gnd.n4840 gnd.n3429 19.3944
R10241 gnd.n4840 gnd.n3427 19.3944
R10242 gnd.n4844 gnd.n3427 19.3944
R10243 gnd.n4844 gnd.n3417 19.3944
R10244 gnd.n4856 gnd.n3417 19.3944
R10245 gnd.n4856 gnd.n3415 19.3944
R10246 gnd.n4860 gnd.n3415 19.3944
R10247 gnd.n4860 gnd.n3404 19.3944
R10248 gnd.n4872 gnd.n3404 19.3944
R10249 gnd.n4872 gnd.n3402 19.3944
R10250 gnd.n4876 gnd.n3402 19.3944
R10251 gnd.n4876 gnd.n3392 19.3944
R10252 gnd.n4888 gnd.n3392 19.3944
R10253 gnd.n4888 gnd.n3390 19.3944
R10254 gnd.n4894 gnd.n3390 19.3944
R10255 gnd.n4894 gnd.n4893 19.3944
R10256 gnd.n4893 gnd.n3363 19.3944
R10257 gnd.n5017 gnd.n3363 19.3944
R10258 gnd.n5017 gnd.n3361 19.3944
R10259 gnd.n5021 gnd.n3361 19.3944
R10260 gnd.n5021 gnd.n3350 19.3944
R10261 gnd.n5033 gnd.n3350 19.3944
R10262 gnd.n5033 gnd.n3348 19.3944
R10263 gnd.n5037 gnd.n3348 19.3944
R10264 gnd.n5037 gnd.n3335 19.3944
R10265 gnd.n5049 gnd.n3335 19.3944
R10266 gnd.n5049 gnd.n3333 19.3944
R10267 gnd.n5053 gnd.n3333 19.3944
R10268 gnd.n5053 gnd.n3321 19.3944
R10269 gnd.n5065 gnd.n3321 19.3944
R10270 gnd.n5065 gnd.n3319 19.3944
R10271 gnd.n5071 gnd.n3319 19.3944
R10272 gnd.n5071 gnd.n5070 19.3944
R10273 gnd.n5070 gnd.n3291 19.3944
R10274 gnd.n5351 gnd.n3291 19.3944
R10275 gnd.n5351 gnd.n3289 19.3944
R10276 gnd.n5355 gnd.n3289 19.3944
R10277 gnd.n5355 gnd.n3279 19.3944
R10278 gnd.n5367 gnd.n3279 19.3944
R10279 gnd.n5367 gnd.n3277 19.3944
R10280 gnd.n5371 gnd.n3277 19.3944
R10281 gnd.n5371 gnd.n3266 19.3944
R10282 gnd.n5383 gnd.n3266 19.3944
R10283 gnd.n5383 gnd.n3264 19.3944
R10284 gnd.n5387 gnd.n3264 19.3944
R10285 gnd.n5387 gnd.n3253 19.3944
R10286 gnd.n5399 gnd.n3253 19.3944
R10287 gnd.n5399 gnd.n3251 19.3944
R10288 gnd.n5403 gnd.n3251 19.3944
R10289 gnd.n5403 gnd.n3240 19.3944
R10290 gnd.n5415 gnd.n3240 19.3944
R10291 gnd.n5415 gnd.n3238 19.3944
R10292 gnd.n5419 gnd.n3238 19.3944
R10293 gnd.n5419 gnd.n3228 19.3944
R10294 gnd.n5433 gnd.n3228 19.3944
R10295 gnd.n5433 gnd.n3226 19.3944
R10296 gnd.n5440 gnd.n3226 19.3944
R10297 gnd.n5440 gnd.n5439 19.3944
R10298 gnd.n5439 gnd.n2787 19.3944
R10299 gnd.n5776 gnd.n2787 19.3944
R10300 gnd.n5776 gnd.n5775 19.3944
R10301 gnd.n5775 gnd.n5774 19.3944
R10302 gnd.n5774 gnd.n2791 19.3944
R10303 gnd.n3029 gnd.n2791 19.3944
R10304 gnd.n3033 gnd.n3029 19.3944
R10305 gnd.n3033 gnd.n3027 19.3944
R10306 gnd.n5482 gnd.n3027 19.3944
R10307 gnd.n5482 gnd.n3025 19.3944
R10308 gnd.n5488 gnd.n3025 19.3944
R10309 gnd.n5488 gnd.n5487 19.3944
R10310 gnd.n5487 gnd.n2999 19.3944
R10311 gnd.n5513 gnd.n2999 19.3944
R10312 gnd.n5513 gnd.n2997 19.3944
R10313 gnd.n5519 gnd.n2997 19.3944
R10314 gnd.n5519 gnd.n5518 19.3944
R10315 gnd.n5518 gnd.n2971 19.3944
R10316 gnd.n5544 gnd.n2971 19.3944
R10317 gnd.n5544 gnd.n2969 19.3944
R10318 gnd.n5557 gnd.n2969 19.3944
R10319 gnd.n5557 gnd.n5556 19.3944
R10320 gnd.n5556 gnd.n5555 19.3944
R10321 gnd.n5555 gnd.n5552 19.3944
R10322 gnd.n5552 gnd.n2917 19.3944
R10323 gnd.n5648 gnd.n2917 19.3944
R10324 gnd.n5648 gnd.n5647 19.3944
R10325 gnd.n5647 gnd.n5646 19.3944
R10326 gnd.n5646 gnd.n2922 19.3944
R10327 gnd.n5642 gnd.n2922 19.3944
R10328 gnd.n5640 gnd.n5639 19.3944
R10329 gnd.n5629 gnd.n5623 19.3944
R10330 gnd.n5627 gnd.n5626 19.3944
R10331 gnd.n7170 gnd.n304 19.3944
R10332 gnd.n7168 gnd.n7167 19.3944
R10333 gnd.n7167 gnd.n306 19.3944
R10334 gnd.n328 gnd.n306 19.3944
R10335 gnd.n329 gnd.n328 19.3944
R10336 gnd.n332 gnd.n329 19.3944
R10337 gnd.n332 gnd.n324 19.3944
R10338 gnd.n7149 gnd.n324 19.3944
R10339 gnd.n7149 gnd.n7148 19.3944
R10340 gnd.n7148 gnd.n7147 19.3944
R10341 gnd.n7147 gnd.n338 19.3944
R10342 gnd.n370 gnd.n338 19.3944
R10343 gnd.n371 gnd.n370 19.3944
R10344 gnd.n374 gnd.n371 19.3944
R10345 gnd.n374 gnd.n366 19.3944
R10346 gnd.n7129 gnd.n366 19.3944
R10347 gnd.n7129 gnd.n7128 19.3944
R10348 gnd.n7128 gnd.n7127 19.3944
R10349 gnd.n7127 gnd.n380 19.3944
R10350 gnd.n6145 gnd.n6144 19.3944
R10351 gnd.n6144 gnd.n6143 19.3944
R10352 gnd.n6143 gnd.n6142 19.3944
R10353 gnd.n6142 gnd.n6140 19.3944
R10354 gnd.n6140 gnd.n6137 19.3944
R10355 gnd.n6137 gnd.n6136 19.3944
R10356 gnd.n6136 gnd.n6133 19.3944
R10357 gnd.n6133 gnd.n6132 19.3944
R10358 gnd.n6132 gnd.n6129 19.3944
R10359 gnd.n6129 gnd.n6128 19.3944
R10360 gnd.n6128 gnd.n6125 19.3944
R10361 gnd.n6125 gnd.n6124 19.3944
R10362 gnd.n6124 gnd.n6121 19.3944
R10363 gnd.n6121 gnd.n6120 19.3944
R10364 gnd.n6120 gnd.n6117 19.3944
R10365 gnd.n6117 gnd.n6116 19.3944
R10366 gnd.n6116 gnd.n6113 19.3944
R10367 gnd.n6111 gnd.n6108 19.3944
R10368 gnd.n6108 gnd.n6107 19.3944
R10369 gnd.n6107 gnd.n6104 19.3944
R10370 gnd.n6104 gnd.n6103 19.3944
R10371 gnd.n6103 gnd.n6100 19.3944
R10372 gnd.n6100 gnd.n6099 19.3944
R10373 gnd.n6099 gnd.n6096 19.3944
R10374 gnd.n6096 gnd.n6095 19.3944
R10375 gnd.n6095 gnd.n6092 19.3944
R10376 gnd.n6092 gnd.n6091 19.3944
R10377 gnd.n6091 gnd.n6088 19.3944
R10378 gnd.n6088 gnd.n6087 19.3944
R10379 gnd.n6087 gnd.n6084 19.3944
R10380 gnd.n6084 gnd.n6083 19.3944
R10381 gnd.n6083 gnd.n6080 19.3944
R10382 gnd.n6080 gnd.n6079 19.3944
R10383 gnd.n6079 gnd.n6076 19.3944
R10384 gnd.n6076 gnd.n6075 19.3944
R10385 gnd.n6068 gnd.n6067 19.3944
R10386 gnd.n6067 gnd.n2400 19.3944
R10387 gnd.n6063 gnd.n2400 19.3944
R10388 gnd.n6063 gnd.n2402 19.3944
R10389 gnd.n4063 gnd.n2402 19.3944
R10390 gnd.n4066 gnd.n4063 19.3944
R10391 gnd.n4066 gnd.n3804 19.3944
R10392 gnd.n4078 gnd.n3804 19.3944
R10393 gnd.n4078 gnd.n3802 19.3944
R10394 gnd.n4082 gnd.n3802 19.3944
R10395 gnd.n4082 gnd.n3797 19.3944
R10396 gnd.n4094 gnd.n3797 19.3944
R10397 gnd.n4094 gnd.n3795 19.3944
R10398 gnd.n4098 gnd.n3795 19.3944
R10399 gnd.n4098 gnd.n3791 19.3944
R10400 gnd.n4110 gnd.n3791 19.3944
R10401 gnd.n4110 gnd.n3789 19.3944
R10402 gnd.n4114 gnd.n3789 19.3944
R10403 gnd.n4114 gnd.n3784 19.3944
R10404 gnd.n4126 gnd.n3784 19.3944
R10405 gnd.n4126 gnd.n3782 19.3944
R10406 gnd.n4130 gnd.n3782 19.3944
R10407 gnd.n4130 gnd.n3778 19.3944
R10408 gnd.n4142 gnd.n3778 19.3944
R10409 gnd.n4142 gnd.n3776 19.3944
R10410 gnd.n4148 gnd.n3776 19.3944
R10411 gnd.n4148 gnd.n3771 19.3944
R10412 gnd.n4161 gnd.n3771 19.3944
R10413 gnd.n4161 gnd.n3769 19.3944
R10414 gnd.n4165 gnd.n3769 19.3944
R10415 gnd.n4165 gnd.n3765 19.3944
R10416 gnd.n4177 gnd.n3765 19.3944
R10417 gnd.n4177 gnd.n3763 19.3944
R10418 gnd.n4181 gnd.n3763 19.3944
R10419 gnd.n4181 gnd.n3758 19.3944
R10420 gnd.n4193 gnd.n3758 19.3944
R10421 gnd.n4193 gnd.n3756 19.3944
R10422 gnd.n4197 gnd.n3756 19.3944
R10423 gnd.n4197 gnd.n3752 19.3944
R10424 gnd.n4209 gnd.n3752 19.3944
R10425 gnd.n4209 gnd.n3750 19.3944
R10426 gnd.n4213 gnd.n3750 19.3944
R10427 gnd.n4213 gnd.n3745 19.3944
R10428 gnd.n4225 gnd.n3745 19.3944
R10429 gnd.n4225 gnd.n3743 19.3944
R10430 gnd.n4229 gnd.n3743 19.3944
R10431 gnd.n4229 gnd.n3739 19.3944
R10432 gnd.n4241 gnd.n3739 19.3944
R10433 gnd.n4241 gnd.n3737 19.3944
R10434 gnd.n4246 gnd.n3737 19.3944
R10435 gnd.n4246 gnd.n3731 19.3944
R10436 gnd.n4258 gnd.n3731 19.3944
R10437 gnd.n4259 gnd.n4258 19.3944
R10438 gnd.n4301 gnd.n3705 19.3944
R10439 gnd.n4301 gnd.n4298 19.3944
R10440 gnd.n4298 gnd.n4295 19.3944
R10441 gnd.n4295 gnd.n4294 19.3944
R10442 gnd.n4294 gnd.n4291 19.3944
R10443 gnd.n4291 gnd.n4290 19.3944
R10444 gnd.n4290 gnd.n4287 19.3944
R10445 gnd.n4287 gnd.n4286 19.3944
R10446 gnd.n4286 gnd.n4283 19.3944
R10447 gnd.n4283 gnd.n4282 19.3944
R10448 gnd.n4282 gnd.n4279 19.3944
R10449 gnd.n4279 gnd.n4278 19.3944
R10450 gnd.n4278 gnd.n4275 19.3944
R10451 gnd.n4275 gnd.n4274 19.3944
R10452 gnd.n4274 gnd.n4271 19.3944
R10453 gnd.n4271 gnd.n4270 19.3944
R10454 gnd.n4270 gnd.n4267 19.3944
R10455 gnd.n4267 gnd.n4266 19.3944
R10456 gnd.n3688 gnd.n3687 19.3944
R10457 gnd.n4587 gnd.n3687 19.3944
R10458 gnd.n4587 gnd.n4586 19.3944
R10459 gnd.n4586 gnd.n4585 19.3944
R10460 gnd.n4585 gnd.n4582 19.3944
R10461 gnd.n4582 gnd.n4581 19.3944
R10462 gnd.n4581 gnd.n4578 19.3944
R10463 gnd.n4578 gnd.n4577 19.3944
R10464 gnd.n4577 gnd.n4574 19.3944
R10465 gnd.n4574 gnd.n4573 19.3944
R10466 gnd.n4573 gnd.n4570 19.3944
R10467 gnd.n4570 gnd.n4569 19.3944
R10468 gnd.n4569 gnd.n4566 19.3944
R10469 gnd.n4566 gnd.n4565 19.3944
R10470 gnd.n4565 gnd.n4562 19.3944
R10471 gnd.n4044 gnd.n3976 19.3944
R10472 gnd.n4044 gnd.n3977 19.3944
R10473 gnd.n4040 gnd.n3977 19.3944
R10474 gnd.n4040 gnd.n2423 19.3944
R10475 gnd.n6053 gnd.n2423 19.3944
R10476 gnd.n6053 gnd.n6052 19.3944
R10477 gnd.n6052 gnd.n6051 19.3944
R10478 gnd.n6051 gnd.n2427 19.3944
R10479 gnd.n6041 gnd.n2427 19.3944
R10480 gnd.n6041 gnd.n6040 19.3944
R10481 gnd.n6040 gnd.n6039 19.3944
R10482 gnd.n6039 gnd.n2448 19.3944
R10483 gnd.n6029 gnd.n2448 19.3944
R10484 gnd.n6029 gnd.n6028 19.3944
R10485 gnd.n6028 gnd.n6027 19.3944
R10486 gnd.n6027 gnd.n2470 19.3944
R10487 gnd.n6017 gnd.n2470 19.3944
R10488 gnd.n6017 gnd.n6016 19.3944
R10489 gnd.n6016 gnd.n6015 19.3944
R10490 gnd.n6015 gnd.n2491 19.3944
R10491 gnd.n6005 gnd.n2491 19.3944
R10492 gnd.n6005 gnd.n6004 19.3944
R10493 gnd.n6004 gnd.n6003 19.3944
R10494 gnd.n6003 gnd.n2513 19.3944
R10495 gnd.n5993 gnd.n2513 19.3944
R10496 gnd.n5993 gnd.n5992 19.3944
R10497 gnd.n5992 gnd.n5991 19.3944
R10498 gnd.n5991 gnd.n2532 19.3944
R10499 gnd.n5980 gnd.n2532 19.3944
R10500 gnd.n5980 gnd.n5979 19.3944
R10501 gnd.n5979 gnd.n5978 19.3944
R10502 gnd.n5978 gnd.n2551 19.3944
R10503 gnd.n5968 gnd.n2551 19.3944
R10504 gnd.n5968 gnd.n5967 19.3944
R10505 gnd.n5967 gnd.n5966 19.3944
R10506 gnd.n5966 gnd.n2571 19.3944
R10507 gnd.n5956 gnd.n2571 19.3944
R10508 gnd.n5956 gnd.n5955 19.3944
R10509 gnd.n5955 gnd.n5954 19.3944
R10510 gnd.n5954 gnd.n2593 19.3944
R10511 gnd.n5944 gnd.n2593 19.3944
R10512 gnd.n5944 gnd.n5943 19.3944
R10513 gnd.n5943 gnd.n5942 19.3944
R10514 gnd.n5942 gnd.n2614 19.3944
R10515 gnd.n5932 gnd.n2614 19.3944
R10516 gnd.n5932 gnd.n5931 19.3944
R10517 gnd.n5931 gnd.n5930 19.3944
R10518 gnd.n5930 gnd.n2636 19.3944
R10519 gnd.n5920 gnd.n2636 19.3944
R10520 gnd.n5920 gnd.n5919 19.3944
R10521 gnd.n5919 gnd.n5918 19.3944
R10522 gnd.n5918 gnd.n2658 19.3944
R10523 gnd.n5908 gnd.n2658 19.3944
R10524 gnd.n4036 gnd.n4034 19.3944
R10525 gnd.n4034 gnd.n4031 19.3944
R10526 gnd.n4031 gnd.n4030 19.3944
R10527 gnd.n4030 gnd.n4027 19.3944
R10528 gnd.n4027 gnd.n4026 19.3944
R10529 gnd.n4026 gnd.n4023 19.3944
R10530 gnd.n4023 gnd.n4022 19.3944
R10531 gnd.n4022 gnd.n4019 19.3944
R10532 gnd.n4019 gnd.n4018 19.3944
R10533 gnd.n4018 gnd.n4015 19.3944
R10534 gnd.n4015 gnd.n4014 19.3944
R10535 gnd.n4014 gnd.n4011 19.3944
R10536 gnd.n4011 gnd.n4010 19.3944
R10537 gnd.n4010 gnd.n4007 19.3944
R10538 gnd.n4007 gnd.n4006 19.3944
R10539 gnd.n4006 gnd.n4003 19.3944
R10540 gnd.n3997 gnd.n3809 19.3944
R10541 gnd.n4055 gnd.n3809 19.3944
R10542 gnd.n4055 gnd.n3807 19.3944
R10543 gnd.n4061 gnd.n3807 19.3944
R10544 gnd.n4062 gnd.n4061 19.3944
R10545 gnd.n4070 gnd.n4062 19.3944
R10546 gnd.n4070 gnd.n3805 19.3944
R10547 gnd.n4074 gnd.n3805 19.3944
R10548 gnd.n4074 gnd.n3800 19.3944
R10549 gnd.n4086 gnd.n3800 19.3944
R10550 gnd.n4086 gnd.n3798 19.3944
R10551 gnd.n4090 gnd.n3798 19.3944
R10552 gnd.n4090 gnd.n3794 19.3944
R10553 gnd.n4102 gnd.n3794 19.3944
R10554 gnd.n4102 gnd.n3792 19.3944
R10555 gnd.n4106 gnd.n3792 19.3944
R10556 gnd.n4106 gnd.n3787 19.3944
R10557 gnd.n4118 gnd.n3787 19.3944
R10558 gnd.n4118 gnd.n3785 19.3944
R10559 gnd.n4122 gnd.n3785 19.3944
R10560 gnd.n4122 gnd.n3781 19.3944
R10561 gnd.n4134 gnd.n3781 19.3944
R10562 gnd.n4134 gnd.n3779 19.3944
R10563 gnd.n4138 gnd.n3779 19.3944
R10564 gnd.n4138 gnd.n3774 19.3944
R10565 gnd.n4152 gnd.n3774 19.3944
R10566 gnd.n4152 gnd.n3772 19.3944
R10567 gnd.n4157 gnd.n3772 19.3944
R10568 gnd.n4157 gnd.n3768 19.3944
R10569 gnd.n4169 gnd.n3768 19.3944
R10570 gnd.n4169 gnd.n3766 19.3944
R10571 gnd.n4173 gnd.n3766 19.3944
R10572 gnd.n4173 gnd.n3761 19.3944
R10573 gnd.n4185 gnd.n3761 19.3944
R10574 gnd.n4185 gnd.n3759 19.3944
R10575 gnd.n4189 gnd.n3759 19.3944
R10576 gnd.n4189 gnd.n3755 19.3944
R10577 gnd.n4201 gnd.n3755 19.3944
R10578 gnd.n4201 gnd.n3753 19.3944
R10579 gnd.n4205 gnd.n3753 19.3944
R10580 gnd.n4205 gnd.n3748 19.3944
R10581 gnd.n4217 gnd.n3748 19.3944
R10582 gnd.n4217 gnd.n3746 19.3944
R10583 gnd.n4221 gnd.n3746 19.3944
R10584 gnd.n4221 gnd.n3742 19.3944
R10585 gnd.n4233 gnd.n3742 19.3944
R10586 gnd.n4233 gnd.n3740 19.3944
R10587 gnd.n4237 gnd.n3740 19.3944
R10588 gnd.n4237 gnd.n3736 19.3944
R10589 gnd.n4250 gnd.n3736 19.3944
R10590 gnd.n4250 gnd.n3733 19.3944
R10591 gnd.n4254 gnd.n3733 19.3944
R10592 gnd.n4254 gnd.n3734 19.3944
R10593 gnd.n4050 gnd.n4046 19.3944
R10594 gnd.n4050 gnd.n2411 19.3944
R10595 gnd.n6059 gnd.n2411 19.3944
R10596 gnd.n6059 gnd.n6058 19.3944
R10597 gnd.n6058 gnd.n6057 19.3944
R10598 gnd.n6057 gnd.n2415 19.3944
R10599 gnd.n6047 gnd.n2415 19.3944
R10600 gnd.n6047 gnd.n6046 19.3944
R10601 gnd.n6046 gnd.n6045 19.3944
R10602 gnd.n6045 gnd.n2438 19.3944
R10603 gnd.n6035 gnd.n2438 19.3944
R10604 gnd.n6035 gnd.n6034 19.3944
R10605 gnd.n6034 gnd.n6033 19.3944
R10606 gnd.n6033 gnd.n2459 19.3944
R10607 gnd.n6023 gnd.n2459 19.3944
R10608 gnd.n6023 gnd.n6022 19.3944
R10609 gnd.n6022 gnd.n6021 19.3944
R10610 gnd.n6021 gnd.n2481 19.3944
R10611 gnd.n6011 gnd.n2481 19.3944
R10612 gnd.n6011 gnd.n6010 19.3944
R10613 gnd.n6010 gnd.n6009 19.3944
R10614 gnd.n6009 gnd.n2502 19.3944
R10615 gnd.n5999 gnd.n5998 19.3944
R10616 gnd.n5998 gnd.n5997 19.3944
R10617 gnd.n5987 gnd.n2539 19.3944
R10618 gnd.n5985 gnd.n5984 19.3944
R10619 gnd.n5974 gnd.n2558 19.3944
R10620 gnd.n5974 gnd.n5973 19.3944
R10621 gnd.n5973 gnd.n5972 19.3944
R10622 gnd.n5972 gnd.n2561 19.3944
R10623 gnd.n5962 gnd.n2561 19.3944
R10624 gnd.n5962 gnd.n5961 19.3944
R10625 gnd.n5961 gnd.n5960 19.3944
R10626 gnd.n5960 gnd.n2582 19.3944
R10627 gnd.n5950 gnd.n2582 19.3944
R10628 gnd.n5950 gnd.n5949 19.3944
R10629 gnd.n5949 gnd.n5948 19.3944
R10630 gnd.n5948 gnd.n2604 19.3944
R10631 gnd.n5938 gnd.n2604 19.3944
R10632 gnd.n5938 gnd.n5937 19.3944
R10633 gnd.n5937 gnd.n5936 19.3944
R10634 gnd.n5936 gnd.n2625 19.3944
R10635 gnd.n5926 gnd.n2625 19.3944
R10636 gnd.n5926 gnd.n5925 19.3944
R10637 gnd.n5925 gnd.n5924 19.3944
R10638 gnd.n5924 gnd.n2647 19.3944
R10639 gnd.n5914 gnd.n2647 19.3944
R10640 gnd.n5914 gnd.n5913 19.3944
R10641 gnd.n5913 gnd.n5912 19.3944
R10642 gnd.n6420 gnd.n6419 19.3944
R10643 gnd.n6419 gnd.n6418 19.3944
R10644 gnd.n6418 gnd.n804 19.3944
R10645 gnd.n6412 gnd.n804 19.3944
R10646 gnd.n6412 gnd.n6411 19.3944
R10647 gnd.n6411 gnd.n6410 19.3944
R10648 gnd.n6410 gnd.n812 19.3944
R10649 gnd.n6404 gnd.n812 19.3944
R10650 gnd.n6404 gnd.n6403 19.3944
R10651 gnd.n6403 gnd.n6402 19.3944
R10652 gnd.n6402 gnd.n820 19.3944
R10653 gnd.n6396 gnd.n820 19.3944
R10654 gnd.n6396 gnd.n6395 19.3944
R10655 gnd.n6395 gnd.n6394 19.3944
R10656 gnd.n6394 gnd.n828 19.3944
R10657 gnd.n6388 gnd.n828 19.3944
R10658 gnd.n6388 gnd.n6387 19.3944
R10659 gnd.n6387 gnd.n6386 19.3944
R10660 gnd.n6386 gnd.n836 19.3944
R10661 gnd.n6380 gnd.n836 19.3944
R10662 gnd.n6380 gnd.n6379 19.3944
R10663 gnd.n6379 gnd.n6378 19.3944
R10664 gnd.n6378 gnd.n844 19.3944
R10665 gnd.n6372 gnd.n844 19.3944
R10666 gnd.n6372 gnd.n6371 19.3944
R10667 gnd.n6371 gnd.n6370 19.3944
R10668 gnd.n6370 gnd.n852 19.3944
R10669 gnd.n6364 gnd.n852 19.3944
R10670 gnd.n6364 gnd.n6363 19.3944
R10671 gnd.n6363 gnd.n6362 19.3944
R10672 gnd.n6362 gnd.n860 19.3944
R10673 gnd.n6356 gnd.n860 19.3944
R10674 gnd.n6356 gnd.n6355 19.3944
R10675 gnd.n6355 gnd.n6354 19.3944
R10676 gnd.n6354 gnd.n868 19.3944
R10677 gnd.n6348 gnd.n868 19.3944
R10678 gnd.n6348 gnd.n6347 19.3944
R10679 gnd.n6347 gnd.n6346 19.3944
R10680 gnd.n6346 gnd.n876 19.3944
R10681 gnd.n6340 gnd.n876 19.3944
R10682 gnd.n6340 gnd.n6339 19.3944
R10683 gnd.n6339 gnd.n6338 19.3944
R10684 gnd.n6338 gnd.n884 19.3944
R10685 gnd.n6332 gnd.n884 19.3944
R10686 gnd.n6332 gnd.n6331 19.3944
R10687 gnd.n6331 gnd.n6330 19.3944
R10688 gnd.n6330 gnd.n892 19.3944
R10689 gnd.n6324 gnd.n892 19.3944
R10690 gnd.n6324 gnd.n6323 19.3944
R10691 gnd.n6323 gnd.n6322 19.3944
R10692 gnd.n6322 gnd.n900 19.3944
R10693 gnd.n6316 gnd.n900 19.3944
R10694 gnd.n6316 gnd.n6315 19.3944
R10695 gnd.n6315 gnd.n6314 19.3944
R10696 gnd.n6314 gnd.n908 19.3944
R10697 gnd.n6308 gnd.n908 19.3944
R10698 gnd.n6308 gnd.n6307 19.3944
R10699 gnd.n6307 gnd.n6306 19.3944
R10700 gnd.n6306 gnd.n916 19.3944
R10701 gnd.n6300 gnd.n916 19.3944
R10702 gnd.n6300 gnd.n6299 19.3944
R10703 gnd.n6299 gnd.n6298 19.3944
R10704 gnd.n6298 gnd.n924 19.3944
R10705 gnd.n6292 gnd.n924 19.3944
R10706 gnd.n6292 gnd.n6291 19.3944
R10707 gnd.n6291 gnd.n6290 19.3944
R10708 gnd.n6290 gnd.n932 19.3944
R10709 gnd.n6284 gnd.n932 19.3944
R10710 gnd.n6284 gnd.n6283 19.3944
R10711 gnd.n6283 gnd.n6282 19.3944
R10712 gnd.n6282 gnd.n940 19.3944
R10713 gnd.n6276 gnd.n940 19.3944
R10714 gnd.n6276 gnd.n6275 19.3944
R10715 gnd.n6275 gnd.n6274 19.3944
R10716 gnd.n6274 gnd.n948 19.3944
R10717 gnd.n6268 gnd.n948 19.3944
R10718 gnd.n6268 gnd.n6267 19.3944
R10719 gnd.n6267 gnd.n6266 19.3944
R10720 gnd.n6266 gnd.n956 19.3944
R10721 gnd.n6260 gnd.n956 19.3944
R10722 gnd.n6260 gnd.n6259 19.3944
R10723 gnd.n6259 gnd.n6258 19.3944
R10724 gnd.n6258 gnd.n964 19.3944
R10725 gnd.n3971 gnd.n964 19.3944
R10726 gnd.n5903 gnd.n5902 19.3944
R10727 gnd.n5902 gnd.n5901 19.3944
R10728 gnd.n5901 gnd.n2681 19.3944
R10729 gnd.n5897 gnd.n2681 19.3944
R10730 gnd.n5897 gnd.n5896 19.3944
R10731 gnd.n5896 gnd.n5895 19.3944
R10732 gnd.n5895 gnd.n2686 19.3944
R10733 gnd.n5891 gnd.n2686 19.3944
R10734 gnd.n5891 gnd.n5890 19.3944
R10735 gnd.n5890 gnd.n5889 19.3944
R10736 gnd.n5889 gnd.n2691 19.3944
R10737 gnd.n5885 gnd.n2691 19.3944
R10738 gnd.n5885 gnd.n5884 19.3944
R10739 gnd.n5884 gnd.n5883 19.3944
R10740 gnd.n5883 gnd.n2696 19.3944
R10741 gnd.n5879 gnd.n2696 19.3944
R10742 gnd.n5879 gnd.n5878 19.3944
R10743 gnd.n5878 gnd.n5877 19.3944
R10744 gnd.n5877 gnd.n2701 19.3944
R10745 gnd.n5873 gnd.n2701 19.3944
R10746 gnd.n5873 gnd.n5872 19.3944
R10747 gnd.n5872 gnd.n5871 19.3944
R10748 gnd.n5871 gnd.n2706 19.3944
R10749 gnd.n5867 gnd.n2706 19.3944
R10750 gnd.n5867 gnd.n5866 19.3944
R10751 gnd.n5866 gnd.n5865 19.3944
R10752 gnd.n5865 gnd.n2711 19.3944
R10753 gnd.n5861 gnd.n2711 19.3944
R10754 gnd.n5861 gnd.n5860 19.3944
R10755 gnd.n5860 gnd.n5859 19.3944
R10756 gnd.n5859 gnd.n2716 19.3944
R10757 gnd.n5855 gnd.n2716 19.3944
R10758 gnd.n5855 gnd.n5854 19.3944
R10759 gnd.n5854 gnd.n5853 19.3944
R10760 gnd.n5853 gnd.n2721 19.3944
R10761 gnd.n5849 gnd.n2721 19.3944
R10762 gnd.n5849 gnd.n5848 19.3944
R10763 gnd.n5848 gnd.n5847 19.3944
R10764 gnd.n5847 gnd.n2726 19.3944
R10765 gnd.n5843 gnd.n2726 19.3944
R10766 gnd.n5843 gnd.n5842 19.3944
R10767 gnd.n5842 gnd.n5841 19.3944
R10768 gnd.n5841 gnd.n2731 19.3944
R10769 gnd.n5837 gnd.n2731 19.3944
R10770 gnd.n5837 gnd.n5836 19.3944
R10771 gnd.n5836 gnd.n5835 19.3944
R10772 gnd.n5835 gnd.n2736 19.3944
R10773 gnd.n5831 gnd.n2736 19.3944
R10774 gnd.n5831 gnd.n5830 19.3944
R10775 gnd.n5830 gnd.n5829 19.3944
R10776 gnd.n5829 gnd.n2741 19.3944
R10777 gnd.n5825 gnd.n2741 19.3944
R10778 gnd.n5825 gnd.n5824 19.3944
R10779 gnd.n5824 gnd.n5823 19.3944
R10780 gnd.n5823 gnd.n2746 19.3944
R10781 gnd.n5819 gnd.n2746 19.3944
R10782 gnd.n5819 gnd.n5818 19.3944
R10783 gnd.n5818 gnd.n5817 19.3944
R10784 gnd.n5817 gnd.n2751 19.3944
R10785 gnd.n5813 gnd.n2751 19.3944
R10786 gnd.n5813 gnd.n5812 19.3944
R10787 gnd.n5812 gnd.n5811 19.3944
R10788 gnd.n5811 gnd.n2756 19.3944
R10789 gnd.n5807 gnd.n2756 19.3944
R10790 gnd.n5807 gnd.n5806 19.3944
R10791 gnd.n5806 gnd.n5805 19.3944
R10792 gnd.n5805 gnd.n2761 19.3944
R10793 gnd.n5801 gnd.n2761 19.3944
R10794 gnd.n5801 gnd.n5800 19.3944
R10795 gnd.n5800 gnd.n5799 19.3944
R10796 gnd.n5799 gnd.n2766 19.3944
R10797 gnd.n5795 gnd.n2766 19.3944
R10798 gnd.n5795 gnd.n5794 19.3944
R10799 gnd.n5794 gnd.n5793 19.3944
R10800 gnd.n5793 gnd.n2771 19.3944
R10801 gnd.n5789 gnd.n2771 19.3944
R10802 gnd.n5789 gnd.n5788 19.3944
R10803 gnd.n5788 gnd.n5787 19.3944
R10804 gnd.n5787 gnd.n2776 19.3944
R10805 gnd.n5783 gnd.n2776 19.3944
R10806 gnd.n5783 gnd.n5782 19.3944
R10807 gnd.n5782 gnd.n5781 19.3944
R10808 gnd.n5458 gnd.n3218 19.3944
R10809 gnd.n5454 gnd.n3218 19.3944
R10810 gnd.n5454 gnd.n5453 19.3944
R10811 gnd.n3135 gnd.n3124 19.3944
R10812 gnd.n3140 gnd.n3135 19.3944
R10813 gnd.n3140 gnd.n3117 19.3944
R10814 gnd.n3151 gnd.n3117 19.3944
R10815 gnd.n3151 gnd.n3115 19.3944
R10816 gnd.n3157 gnd.n3115 19.3944
R10817 gnd.n3157 gnd.n3108 19.3944
R10818 gnd.n3168 gnd.n3108 19.3944
R10819 gnd.n3168 gnd.n3106 19.3944
R10820 gnd.n3174 gnd.n3106 19.3944
R10821 gnd.n3174 gnd.n3099 19.3944
R10822 gnd.n3185 gnd.n3099 19.3944
R10823 gnd.n3185 gnd.n3097 19.3944
R10824 gnd.n3191 gnd.n3097 19.3944
R10825 gnd.n3191 gnd.n3087 19.3944
R10826 gnd.n3200 gnd.n3087 19.3944
R10827 gnd.n3200 gnd.n3085 19.3944
R10828 gnd.n3085 gnd.n3084 19.3944
R10829 gnd.n5469 gnd.n3084 19.3944
R10830 gnd.n5469 gnd.n5468 19.3944
R10831 gnd.n5468 gnd.n5467 19.3944
R10832 gnd.n5467 gnd.n3210 19.3944
R10833 gnd.n5463 gnd.n3210 19.3944
R10834 gnd.n5463 gnd.n5462 19.3944
R10835 gnd.n1850 gnd.t59 18.8012
R10836 gnd.n1835 gnd.t69 18.8012
R10837 gnd.n1694 gnd.n1693 18.4825
R10838 gnd.n5739 gnd.n5738 18.4247
R10839 gnd.n4562 gnd.n4561 18.4247
R10840 gnd.n7319 gnd.n7318 18.2308
R10841 gnd.n3196 gnd.n3195 18.2308
R10842 gnd.n3663 gnd.n3562 18.2308
R10843 gnd.n4003 gnd.n3996 18.2308
R10844 gnd.t44 gnd.n1374 18.1639
R10845 gnd.n4444 gnd.n4442 17.8452
R10846 gnd.n4794 gnd.n4793 17.8452
R10847 gnd.n4906 gnd.t21 17.8452
R10848 gnd.n5009 gnd.t0 17.8452
R10849 gnd.n5039 gnd.n3344 17.8452
R10850 gnd.n5373 gnd.n3274 17.8452
R10851 gnd.n4489 gnd.n4431 17.6395
R10852 gnd.n5310 gnd.n5133 17.6395
R10853 gnd.n1402 gnd.t57 17.5266
R10854 gnd.n4068 gnd.t236 17.5266
R10855 gnd.n4862 gnd.t34 17.5266
R10856 gnd.n4972 gnd.t60 17.5266
R10857 gnd.n7271 gnd.t264 17.5266
R10858 gnd.n3440 gnd.t20 17.2079
R10859 gnd.n4854 gnd.t38 17.2079
R10860 gnd.n4945 gnd.t43 17.2079
R10861 gnd.n5083 gnd.t32 17.2079
R10862 gnd.n1801 gnd.t52 16.8893
R10863 gnd.n4100 gnd.t222 16.8893
R10864 gnd.n3749 gnd.t202 16.8893
R10865 gnd.n5542 gnd.t274 16.8893
R10866 gnd.n7239 gnd.t234 16.8893
R10867 gnd.n6254 gnd.n6253 16.5706
R10868 gnd.n4689 gnd.n3473 16.5706
R10869 gnd.n4483 gnd.n4482 16.5706
R10870 gnd.n4870 gnd.n3406 16.5706
R10871 gnd.n4751 gnd.n3400 16.5706
R10872 gnd.n5047 gnd.n3337 16.5706
R10873 gnd.n4930 gnd.n3329 16.5706
R10874 gnd.n5381 gnd.n3268 16.5706
R10875 gnd.n5110 gnd.n5108 16.5706
R10876 gnd.n5397 gnd.t154 16.5706
R10877 gnd.n1629 gnd.t107 16.2519
R10878 gnd.n1329 gnd.t51 16.2519
R10879 gnd.n4132 gnd.t209 16.2519
R10880 gnd.n3762 gnd.t191 16.2519
R10881 gnd.n4633 gnd.t146 16.2519
R10882 gnd.t115 gnd.n2782 16.2519
R10883 gnd.n2915 gnd.t218 16.2519
R10884 gnd.n7207 gnd.t206 16.2519
R10885 gnd.n4310 gnd.n4309 16.0975
R10886 gnd.n5166 gnd.n5165 16.0975
R10887 gnd.n4365 gnd.n4364 16.0975
R10888 gnd.n5160 gnd.n5159 16.0975
R10889 gnd.n2276 gnd.n2274 15.6674
R10890 gnd.n2244 gnd.n2242 15.6674
R10891 gnd.n2212 gnd.n2210 15.6674
R10892 gnd.n2181 gnd.n2179 15.6674
R10893 gnd.n2149 gnd.n2147 15.6674
R10894 gnd.n2117 gnd.n2115 15.6674
R10895 gnd.n2085 gnd.n2083 15.6674
R10896 gnd.n2054 gnd.n2052 15.6674
R10897 gnd.n1620 gnd.t107 15.6146
R10898 gnd.n2313 gnd.t150 15.6146
R10899 gnd.t136 gnd.n1040 15.6146
R10900 gnd.n3775 gnd.t189 15.6146
R10901 gnd.n4167 gnd.t199 15.6146
R10902 gnd.t146 gnd.n3514 15.6146
R10903 gnd.n5442 gnd.t115 15.6146
R10904 gnd.n5609 gnd.t185 15.6146
R10905 gnd.n5621 gnd.t267 15.6146
R10906 gnd.n4327 gnd.n3473 15.296
R10907 gnd.n4460 gnd.t8 15.296
R10908 gnd.n4810 gnd.n3406 15.296
R10909 gnd.n4878 gnd.n3400 15.296
R10910 gnd.n4987 gnd.n3337 15.296
R10911 gnd.n5055 gnd.n3329 15.296
R10912 gnd.n5357 gnd.t182 15.296
R10913 gnd.n5118 gnd.n5117 15.0827
R10914 gnd.n4338 gnd.n4333 15.0481
R10915 gnd.n5128 gnd.n5127 15.0481
R10916 gnd.t46 gnd.n968 14.9773
R10917 gnd.n3788 gnd.t225 14.9773
R10918 gnd.n4199 gnd.t183 14.9773
R10919 gnd.n5571 gnd.t193 14.9773
R10920 gnd.t279 gnd.n246 14.9773
R10921 gnd.n4482 gnd.t126 14.6587
R10922 gnd.t119 gnd.n3268 14.6587
R10923 gnd.t319 gnd.n992 14.34
R10924 gnd.n1151 gnd.t55 14.34
R10925 gnd.n3801 gnd.t254 14.34
R10926 gnd.n4231 gnd.t187 14.34
R10927 gnd.t257 gnd.n5510 14.34
R10928 gnd.t216 gnd.n216 14.34
R10929 gnd.n4832 gnd.t14 14.0214
R10930 gnd.t31 gnd.n3307 14.0214
R10931 gnd.n5096 gnd.n3274 14.0214
R10932 gnd.n1776 gnd.t39 13.7027
R10933 gnd.n5314 gnd.t41 13.7027
R10934 gnd.n1486 gnd.n1485 13.5763
R10935 gnd.n6203 gnd.n1053 13.5763
R10936 gnd.n5701 gnd.n2868 13.5763
R10937 gnd.n7371 gnd.n7370 13.5763
R10938 gnd.n6075 gnd.n2397 13.5763
R10939 gnd.n4266 gnd.n4263 13.5763
R10940 gnd.n1694 gnd.n1432 13.384
R10941 gnd.n4786 gnd.t33 13.384
R10942 gnd.n5031 gnd.t68 13.384
R10943 gnd.n4349 gnd.n4330 13.1884
R10944 gnd.n4344 gnd.n4343 13.1884
R10945 gnd.n4343 gnd.n4342 13.1884
R10946 gnd.n5121 gnd.n5116 13.1884
R10947 gnd.n5122 gnd.n5121 13.1884
R10948 gnd.n4345 gnd.n4332 13.146
R10949 gnd.n4341 gnd.n4332 13.146
R10950 gnd.n5120 gnd.n5119 13.146
R10951 gnd.n5120 gnd.n5115 13.146
R10952 gnd.t18 gnd.n3387 13.0654
R10953 gnd.n5003 gnd.t71 13.0654
R10954 gnd.n2277 gnd.n2273 12.8005
R10955 gnd.n2245 gnd.n2241 12.8005
R10956 gnd.n2213 gnd.n2209 12.8005
R10957 gnd.n2182 gnd.n2178 12.8005
R10958 gnd.n2150 gnd.n2146 12.8005
R10959 gnd.n2118 gnd.n2114 12.8005
R10960 gnd.n2086 gnd.n2082 12.8005
R10961 gnd.n2055 gnd.n2051 12.8005
R10962 gnd.n4825 gnd.n4824 12.7467
R10963 gnd.n4802 gnd.t6 12.7467
R10964 gnd.n4896 gnd.n3386 12.7467
R10965 gnd.n5002 gnd.n5001 12.7467
R10966 gnd.t27 gnd.n3338 12.7467
R10967 gnd.n5073 gnd.n3314 12.7467
R10968 gnd.n5335 gnd.t64 12.4281
R10969 gnd.n1485 gnd.n1480 12.4126
R10970 gnd.n6199 gnd.n1053 12.4126
R10971 gnd.n5697 gnd.n2868 12.4126
R10972 gnd.n7370 gnd.n174 12.4126
R10973 gnd.n6071 gnd.n2397 12.4126
R10974 gnd.n4263 gnd.n3727 12.4126
R10975 gnd.n4431 gnd.n4430 12.1761
R10976 gnd.n5134 gnd.n5133 12.1761
R10977 gnd.t169 gnd.n3275 12.1094
R10978 gnd.n2281 gnd.n2280 12.0247
R10979 gnd.n2249 gnd.n2248 12.0247
R10980 gnd.n2217 gnd.n2216 12.0247
R10981 gnd.n2186 gnd.n2185 12.0247
R10982 gnd.n2154 gnd.n2153 12.0247
R10983 gnd.n2122 gnd.n2121 12.0247
R10984 gnd.n2090 gnd.n2089 12.0247
R10985 gnd.n2059 gnd.n2058 12.0247
R10986 gnd.n3732 gnd.t97 11.7908
R10987 gnd.n5480 gnd.t86 11.7908
R10988 gnd.n4705 gnd.t130 11.4721
R10989 gnd.n4725 gnd.n4724 11.4721
R10990 gnd.n4832 gnd.n3439 11.4721
R10991 gnd.n4906 gnd.n4905 11.4721
R10992 gnd.n5009 gnd.n3374 11.4721
R10993 gnd.n5082 gnd.n3307 11.4721
R10994 gnd.n5343 gnd.n3302 11.4721
R10995 gnd.n2284 gnd.n2271 11.249
R10996 gnd.n2252 gnd.n2239 11.249
R10997 gnd.n2220 gnd.n2207 11.249
R10998 gnd.n2189 gnd.n2176 11.249
R10999 gnd.n2157 gnd.n2144 11.249
R11000 gnd.n2125 gnd.n2112 11.249
R11001 gnd.n2093 gnd.n2080 11.249
R11002 gnd.n2062 gnd.n2049 11.249
R11003 gnd.n1764 gnd.t39 11.1535
R11004 gnd.n3508 gnd.t73 11.1535
R11005 gnd.n5421 gnd.t313 11.1535
R11006 gnd.n4059 gnd.n2407 10.8348
R11007 gnd.n6055 gnd.n2417 10.8348
R11008 gnd.n4068 gnd.n2420 10.8348
R11009 gnd.n6049 gnd.n2429 10.8348
R11010 gnd.n4076 gnd.n2432 10.8348
R11011 gnd.n6043 gnd.n2440 10.8348
R11012 gnd.n4084 gnd.n3801 10.8348
R11013 gnd.n6037 gnd.n2450 10.8348
R11014 gnd.n6031 gnd.n2461 10.8348
R11015 gnd.n4100 gnd.n2464 10.8348
R11016 gnd.n6025 gnd.n2472 10.8348
R11017 gnd.n4108 gnd.n2475 10.8348
R11018 gnd.n6019 gnd.n2483 10.8348
R11019 gnd.n4116 gnd.n3788 10.8348
R11020 gnd.n6013 gnd.n2493 10.8348
R11021 gnd.n6007 gnd.n2504 10.8348
R11022 gnd.n4132 gnd.n2507 10.8348
R11023 gnd.n6001 gnd.n2515 10.8348
R11024 gnd.n4140 gnd.n2518 10.8348
R11025 gnd.n5995 gnd.n2524 10.8348
R11026 gnd.n4150 gnd.n3775 10.8348
R11027 gnd.n5989 gnd.n2534 10.8348
R11028 gnd.n5982 gnd.n2542 10.8348
R11029 gnd.n4167 gnd.n2545 10.8348
R11030 gnd.n5976 gnd.n2553 10.8348
R11031 gnd.n4175 gnd.n2556 10.8348
R11032 gnd.n5970 gnd.n2563 10.8348
R11033 gnd.n4183 gnd.n3762 10.8348
R11034 gnd.n5964 gnd.n2573 10.8348
R11035 gnd.n5958 gnd.n2584 10.8348
R11036 gnd.n4199 gnd.n2587 10.8348
R11037 gnd.n5952 gnd.n2595 10.8348
R11038 gnd.n4207 gnd.n2598 10.8348
R11039 gnd.n5946 gnd.n2606 10.8348
R11040 gnd.n4215 gnd.n3749 10.8348
R11041 gnd.n5940 gnd.n2616 10.8348
R11042 gnd.n5934 gnd.n2627 10.8348
R11043 gnd.n4231 gnd.n2630 10.8348
R11044 gnd.n5928 gnd.n2638 10.8348
R11045 gnd.n4239 gnd.n2641 10.8348
R11046 gnd.n5922 gnd.n2649 10.8348
R11047 gnd.n4248 gnd.n2652 10.8348
R11048 gnd.n5916 gnd.n2660 10.8348
R11049 gnd.n4256 gnd.n3732 10.8348
R11050 gnd.n5910 gnd.n2669 10.8348
R11051 gnd.n5694 gnd.n2874 10.8348
R11052 gnd.n5480 gnd.n3041 10.8348
R11053 gnd.n5479 gnd.n3019 10.8348
R11054 gnd.n5491 gnd.n5490 10.8348
R11055 gnd.n3022 gnd.n3009 10.8348
R11056 gnd.n5501 gnd.n3011 10.8348
R11057 gnd.n5511 gnd.n3001 10.8348
R11058 gnd.n5510 gnd.n2990 10.8348
R11059 gnd.n5522 gnd.n5521 10.8348
R11060 gnd.n5532 gnd.n2983 10.8348
R11061 gnd.n5542 gnd.n2973 10.8348
R11062 gnd.n5541 gnd.n2962 10.8348
R11063 gnd.n5561 gnd.n5559 10.8348
R11064 gnd.n2967 gnd.n2965 10.8348
R11065 gnd.n5571 gnd.n2954 10.8348
R11066 gnd.n2956 gnd.n2946 10.8348
R11067 gnd.n5651 gnd.n5650 10.8348
R11068 gnd.n2915 gnd.n2913 10.8348
R11069 gnd.n5659 gnd.n2904 10.8348
R11070 gnd.n5597 gnd.n273 10.8348
R11071 gnd.n7200 gnd.n276 10.8348
R11072 gnd.n5609 gnd.n5608 10.8348
R11073 gnd.n5637 gnd.n2926 10.8348
R11074 gnd.n5632 gnd.n5631 10.8348
R11075 gnd.n5621 gnd.n5620 10.8348
R11076 gnd.n7179 gnd.n290 10.8348
R11077 gnd.n7184 gnd.n292 10.8348
R11078 gnd.n7173 gnd.n7172 10.8348
R11079 gnd.n7207 gnd.n260 10.8348
R11080 gnd.n310 gnd.n252 10.8348
R11081 gnd.n7163 gnd.n244 10.8348
R11082 gnd.n7223 gnd.n246 10.8348
R11083 gnd.n7156 gnd.n236 10.8348
R11084 gnd.n7231 gnd.n238 10.8348
R11085 gnd.n7152 gnd.n7151 10.8348
R11086 gnd.n7239 gnd.n230 10.8348
R11087 gnd.n342 gnd.n222 10.8348
R11088 gnd.n7143 gnd.n214 10.8348
R11089 gnd.n7255 gnd.n216 10.8348
R11090 gnd.n7136 gnd.n206 10.8348
R11091 gnd.n7263 gnd.n208 10.8348
R11092 gnd.n7132 gnd.n7131 10.8348
R11093 gnd.n7271 gnd.n200 10.8348
R11094 gnd.n359 gnd.n189 10.8348
R11095 gnd.n7354 gnd.n191 10.8348
R11096 gnd.n5245 gnd.n5163 10.6151
R11097 gnd.n5245 gnd.n5244 10.6151
R11098 gnd.n5242 gnd.n5167 10.6151
R11099 gnd.n5237 gnd.n5167 10.6151
R11100 gnd.n5237 gnd.n5236 10.6151
R11101 gnd.n5236 gnd.n5235 10.6151
R11102 gnd.n5235 gnd.n5170 10.6151
R11103 gnd.n5230 gnd.n5170 10.6151
R11104 gnd.n5230 gnd.n5229 10.6151
R11105 gnd.n5229 gnd.n5228 10.6151
R11106 gnd.n5228 gnd.n5173 10.6151
R11107 gnd.n5223 gnd.n5173 10.6151
R11108 gnd.n5223 gnd.n5222 10.6151
R11109 gnd.n5222 gnd.n5221 10.6151
R11110 gnd.n5221 gnd.n5176 10.6151
R11111 gnd.n5216 gnd.n5176 10.6151
R11112 gnd.n5216 gnd.n5215 10.6151
R11113 gnd.n5215 gnd.n5214 10.6151
R11114 gnd.n5214 gnd.n5179 10.6151
R11115 gnd.n5209 gnd.n5179 10.6151
R11116 gnd.n5209 gnd.n5208 10.6151
R11117 gnd.n5208 gnd.n5207 10.6151
R11118 gnd.n5207 gnd.n5182 10.6151
R11119 gnd.n5202 gnd.n5182 10.6151
R11120 gnd.n5202 gnd.n5201 10.6151
R11121 gnd.n5201 gnd.n5200 10.6151
R11122 gnd.n5200 gnd.n5185 10.6151
R11123 gnd.n5195 gnd.n5185 10.6151
R11124 gnd.n5195 gnd.n5194 10.6151
R11125 gnd.n5194 gnd.n5193 10.6151
R11126 gnd.n4436 gnd.n4325 10.6151
R11127 gnd.n4438 gnd.n4436 10.6151
R11128 gnd.n4439 gnd.n4438 10.6151
R11129 gnd.n4480 gnd.n4439 10.6151
R11130 gnd.n4480 gnd.n4479 10.6151
R11131 gnd.n4479 gnd.n4478 10.6151
R11132 gnd.n4478 gnd.n4440 10.6151
R11133 gnd.n4457 gnd.n4440 10.6151
R11134 gnd.n4458 gnd.n4457 10.6151
R11135 gnd.n4465 gnd.n4458 10.6151
R11136 gnd.n4465 gnd.n4464 10.6151
R11137 gnd.n4464 gnd.n4463 10.6151
R11138 gnd.n4463 gnd.n4459 10.6151
R11139 gnd.n4459 gnd.n3436 10.6151
R11140 gnd.n4836 gnd.n3436 10.6151
R11141 gnd.n4836 gnd.n4835 10.6151
R11142 gnd.n4835 gnd.n4834 10.6151
R11143 gnd.n4834 gnd.n3437 10.6151
R11144 gnd.n4736 gnd.n3437 10.6151
R11145 gnd.n4822 gnd.n4736 10.6151
R11146 gnd.n4822 gnd.n4821 10.6151
R11147 gnd.n4821 gnd.n4820 10.6151
R11148 gnd.n4820 gnd.n4737 10.6151
R11149 gnd.n4748 gnd.n4737 10.6151
R11150 gnd.n4807 gnd.n4748 10.6151
R11151 gnd.n4807 gnd.n4806 10.6151
R11152 gnd.n4806 gnd.n4805 10.6151
R11153 gnd.n4805 gnd.n4749 10.6151
R11154 gnd.n4770 gnd.n4749 10.6151
R11155 gnd.n4771 gnd.n4770 10.6151
R11156 gnd.n4772 gnd.n4771 10.6151
R11157 gnd.n4773 gnd.n4772 10.6151
R11158 gnd.n4774 gnd.n4773 10.6151
R11159 gnd.n4784 gnd.n4774 10.6151
R11160 gnd.n4784 gnd.n4783 10.6151
R11161 gnd.n4783 gnd.n4782 10.6151
R11162 gnd.n4782 gnd.n4776 10.6151
R11163 gnd.n4776 gnd.n4775 10.6151
R11164 gnd.n4775 gnd.n3371 10.6151
R11165 gnd.n5013 gnd.n3371 10.6151
R11166 gnd.n5013 gnd.n5012 10.6151
R11167 gnd.n5012 gnd.n5011 10.6151
R11168 gnd.n5011 gnd.n3372 10.6151
R11169 gnd.n4916 gnd.n3372 10.6151
R11170 gnd.n4999 gnd.n4916 10.6151
R11171 gnd.n4999 gnd.n4998 10.6151
R11172 gnd.n4998 gnd.n4997 10.6151
R11173 gnd.n4997 gnd.n4917 10.6151
R11174 gnd.n4927 gnd.n4917 10.6151
R11175 gnd.n4985 gnd.n4927 10.6151
R11176 gnd.n4985 gnd.n4984 10.6151
R11177 gnd.n4984 gnd.n4983 10.6151
R11178 gnd.n4983 gnd.n4928 10.6151
R11179 gnd.n4939 gnd.n4928 10.6151
R11180 gnd.n4941 gnd.n4939 10.6151
R11181 gnd.n4942 gnd.n4941 10.6151
R11182 gnd.n4969 gnd.n4942 10.6151
R11183 gnd.n4969 gnd.n4968 10.6151
R11184 gnd.n4968 gnd.n4967 10.6151
R11185 gnd.n4967 gnd.n4943 10.6151
R11186 gnd.n4953 gnd.n4943 10.6151
R11187 gnd.n4955 gnd.n4953 10.6151
R11188 gnd.n4955 gnd.n4954 10.6151
R11189 gnd.n4954 gnd.n3298 10.6151
R11190 gnd.n5347 gnd.n3298 10.6151
R11191 gnd.n5347 gnd.n5346 10.6151
R11192 gnd.n5346 gnd.n5345 10.6151
R11193 gnd.n5345 gnd.n3299 10.6151
R11194 gnd.n5092 gnd.n3299 10.6151
R11195 gnd.n5333 gnd.n5092 10.6151
R11196 gnd.n5333 gnd.n5332 10.6151
R11197 gnd.n5332 gnd.n5331 10.6151
R11198 gnd.n5331 gnd.n5093 10.6151
R11199 gnd.n5104 gnd.n5093 10.6151
R11200 gnd.n5319 gnd.n5104 10.6151
R11201 gnd.n5319 gnd.n5318 10.6151
R11202 gnd.n5318 gnd.n5317 10.6151
R11203 gnd.n5317 gnd.n5105 10.6151
R11204 gnd.n5188 gnd.n5105 10.6151
R11205 gnd.n5189 gnd.n5188 10.6151
R11206 gnd.n4554 gnd.n4305 10.6151
R11207 gnd.n4554 gnd.n4553 10.6151
R11208 gnd.n4551 gnd.n4311 10.6151
R11209 gnd.n4545 gnd.n4311 10.6151
R11210 gnd.n4545 gnd.n4544 10.6151
R11211 gnd.n4544 gnd.n4543 10.6151
R11212 gnd.n4543 gnd.n4313 10.6151
R11213 gnd.n4537 gnd.n4313 10.6151
R11214 gnd.n4537 gnd.n4536 10.6151
R11215 gnd.n4536 gnd.n4535 10.6151
R11216 gnd.n4535 gnd.n4315 10.6151
R11217 gnd.n4529 gnd.n4315 10.6151
R11218 gnd.n4529 gnd.n4528 10.6151
R11219 gnd.n4528 gnd.n4527 10.6151
R11220 gnd.n4527 gnd.n4317 10.6151
R11221 gnd.n4521 gnd.n4317 10.6151
R11222 gnd.n4521 gnd.n4520 10.6151
R11223 gnd.n4520 gnd.n4519 10.6151
R11224 gnd.n4519 gnd.n4319 10.6151
R11225 gnd.n4513 gnd.n4319 10.6151
R11226 gnd.n4513 gnd.n4512 10.6151
R11227 gnd.n4512 gnd.n4511 10.6151
R11228 gnd.n4511 gnd.n4321 10.6151
R11229 gnd.n4505 gnd.n4321 10.6151
R11230 gnd.n4505 gnd.n4504 10.6151
R11231 gnd.n4504 gnd.n4503 10.6151
R11232 gnd.n4503 gnd.n4323 10.6151
R11233 gnd.n4497 gnd.n4323 10.6151
R11234 gnd.n4497 gnd.n4496 10.6151
R11235 gnd.n4496 gnd.n4495 10.6151
R11236 gnd.n4430 gnd.n4429 10.6151
R11237 gnd.n4429 gnd.n4350 10.6151
R11238 gnd.n4424 gnd.n4350 10.6151
R11239 gnd.n4424 gnd.n4423 10.6151
R11240 gnd.n4423 gnd.n4352 10.6151
R11241 gnd.n4418 gnd.n4352 10.6151
R11242 gnd.n4418 gnd.n4417 10.6151
R11243 gnd.n4417 gnd.n4416 10.6151
R11244 gnd.n4416 gnd.n4354 10.6151
R11245 gnd.n4410 gnd.n4354 10.6151
R11246 gnd.n4410 gnd.n4409 10.6151
R11247 gnd.n4409 gnd.n4408 10.6151
R11248 gnd.n4408 gnd.n4356 10.6151
R11249 gnd.n4402 gnd.n4356 10.6151
R11250 gnd.n4402 gnd.n4401 10.6151
R11251 gnd.n4401 gnd.n4400 10.6151
R11252 gnd.n4400 gnd.n4358 10.6151
R11253 gnd.n4394 gnd.n4358 10.6151
R11254 gnd.n4394 gnd.n4393 10.6151
R11255 gnd.n4393 gnd.n4392 10.6151
R11256 gnd.n4392 gnd.n4360 10.6151
R11257 gnd.n4386 gnd.n4360 10.6151
R11258 gnd.n4386 gnd.n4385 10.6151
R11259 gnd.n4385 gnd.n4384 10.6151
R11260 gnd.n4384 gnd.n4362 10.6151
R11261 gnd.n4378 gnd.n4362 10.6151
R11262 gnd.n4378 gnd.n4377 10.6151
R11263 gnd.n4377 gnd.n4376 10.6151
R11264 gnd.n4372 gnd.n4371 10.6151
R11265 gnd.n4371 gnd.n4306 10.6151
R11266 gnd.n5305 gnd.n5134 10.6151
R11267 gnd.n5305 gnd.n5304 10.6151
R11268 gnd.n5304 gnd.n5303 10.6151
R11269 gnd.n5303 gnd.n5138 10.6151
R11270 gnd.n5298 gnd.n5138 10.6151
R11271 gnd.n5298 gnd.n5297 10.6151
R11272 gnd.n5297 gnd.n5296 10.6151
R11273 gnd.n5296 gnd.n5141 10.6151
R11274 gnd.n5291 gnd.n5141 10.6151
R11275 gnd.n5291 gnd.n5290 10.6151
R11276 gnd.n5290 gnd.n5289 10.6151
R11277 gnd.n5289 gnd.n5144 10.6151
R11278 gnd.n5284 gnd.n5144 10.6151
R11279 gnd.n5284 gnd.n5283 10.6151
R11280 gnd.n5283 gnd.n5282 10.6151
R11281 gnd.n5282 gnd.n5147 10.6151
R11282 gnd.n5277 gnd.n5147 10.6151
R11283 gnd.n5277 gnd.n5276 10.6151
R11284 gnd.n5276 gnd.n5275 10.6151
R11285 gnd.n5275 gnd.n5150 10.6151
R11286 gnd.n5270 gnd.n5150 10.6151
R11287 gnd.n5270 gnd.n5269 10.6151
R11288 gnd.n5269 gnd.n5268 10.6151
R11289 gnd.n5268 gnd.n5153 10.6151
R11290 gnd.n5263 gnd.n5153 10.6151
R11291 gnd.n5263 gnd.n5262 10.6151
R11292 gnd.n5262 gnd.n5261 10.6151
R11293 gnd.n5261 gnd.n5156 10.6151
R11294 gnd.n5256 gnd.n5255 10.6151
R11295 gnd.n5255 gnd.n5254 10.6151
R11296 gnd.n4489 gnd.n4488 10.6151
R11297 gnd.n4488 gnd.n4487 10.6151
R11298 gnd.n4487 gnd.n4432 10.6151
R11299 gnd.n4446 gnd.n4432 10.6151
R11300 gnd.n4447 gnd.n4446 10.6151
R11301 gnd.n4474 gnd.n4447 10.6151
R11302 gnd.n4474 gnd.n4473 10.6151
R11303 gnd.n4473 gnd.n4472 10.6151
R11304 gnd.n4472 gnd.n4448 10.6151
R11305 gnd.n4452 gnd.n4448 10.6151
R11306 gnd.n4452 gnd.n4451 10.6151
R11307 gnd.n4451 gnd.n4450 10.6151
R11308 gnd.n4450 gnd.n3443 10.6151
R11309 gnd.n4728 gnd.n3443 10.6151
R11310 gnd.n4729 gnd.n4728 10.6151
R11311 gnd.n4730 gnd.n4729 10.6151
R11312 gnd.n4830 gnd.n4730 10.6151
R11313 gnd.n4830 gnd.n4829 10.6151
R11314 gnd.n4829 gnd.n4828 10.6151
R11315 gnd.n4828 gnd.n4731 10.6151
R11316 gnd.n4743 gnd.n4731 10.6151
R11317 gnd.n4816 gnd.n4743 10.6151
R11318 gnd.n4816 gnd.n4815 10.6151
R11319 gnd.n4815 gnd.n4814 10.6151
R11320 gnd.n4814 gnd.n4744 10.6151
R11321 gnd.n4754 gnd.n4744 10.6151
R11322 gnd.n4755 gnd.n4754 10.6151
R11323 gnd.n4800 gnd.n4755 10.6151
R11324 gnd.n4800 gnd.n4799 10.6151
R11325 gnd.n4799 gnd.n4798 10.6151
R11326 gnd.n4798 gnd.n4756 10.6151
R11327 gnd.n4791 gnd.n4756 10.6151
R11328 gnd.n4791 gnd.n4790 10.6151
R11329 gnd.n4790 gnd.n4789 10.6151
R11330 gnd.n4789 gnd.n4763 10.6151
R11331 gnd.n4765 gnd.n4763 10.6151
R11332 gnd.n4765 gnd.n4764 10.6151
R11333 gnd.n4764 gnd.n3377 10.6151
R11334 gnd.n4909 gnd.n3377 10.6151
R11335 gnd.n4910 gnd.n4909 10.6151
R11336 gnd.n4911 gnd.n4910 10.6151
R11337 gnd.n5007 gnd.n4911 10.6151
R11338 gnd.n5007 gnd.n5006 10.6151
R11339 gnd.n5006 gnd.n5005 10.6151
R11340 gnd.n5005 gnd.n4912 10.6151
R11341 gnd.n4922 gnd.n4912 10.6151
R11342 gnd.n4993 gnd.n4922 10.6151
R11343 gnd.n4993 gnd.n4992 10.6151
R11344 gnd.n4992 gnd.n4991 10.6151
R11345 gnd.n4991 gnd.n4923 10.6151
R11346 gnd.n4933 gnd.n4923 10.6151
R11347 gnd.n4934 gnd.n4933 10.6151
R11348 gnd.n4978 gnd.n4934 10.6151
R11349 gnd.n4978 gnd.n4977 10.6151
R11350 gnd.n4977 gnd.n4976 10.6151
R11351 gnd.n4976 gnd.n4935 10.6151
R11352 gnd.n4948 gnd.n4935 10.6151
R11353 gnd.n4949 gnd.n4948 10.6151
R11354 gnd.n4963 gnd.n4949 10.6151
R11355 gnd.n4963 gnd.n4962 10.6151
R11356 gnd.n4962 gnd.n4961 10.6151
R11357 gnd.n4961 gnd.n4950 10.6151
R11358 gnd.n4950 gnd.n3305 10.6151
R11359 gnd.n5085 gnd.n3305 10.6151
R11360 gnd.n5086 gnd.n5085 10.6151
R11361 gnd.n5087 gnd.n5086 10.6151
R11362 gnd.n5341 gnd.n5087 10.6151
R11363 gnd.n5341 gnd.n5340 10.6151
R11364 gnd.n5340 gnd.n5339 10.6151
R11365 gnd.n5339 gnd.n5088 10.6151
R11366 gnd.n5099 gnd.n5088 10.6151
R11367 gnd.n5327 gnd.n5099 10.6151
R11368 gnd.n5327 gnd.n5326 10.6151
R11369 gnd.n5326 gnd.n5325 10.6151
R11370 gnd.n5325 gnd.n5100 10.6151
R11371 gnd.n5112 gnd.n5100 10.6151
R11372 gnd.n5113 gnd.n5112 10.6151
R11373 gnd.n5312 gnd.n5113 10.6151
R11374 gnd.n5312 gnd.n5311 10.6151
R11375 gnd.n5311 gnd.n5310 10.6151
R11376 gnd.n1683 gnd.t315 10.5161
R11377 gnd.n1977 gnd.t319 10.5161
R11378 gnd.t55 gnd.n1015 10.5161
R11379 gnd.n4681 gnd.n3481 10.5161
R11380 gnd.n5136 gnd.n5135 10.5161
R11381 gnd.n2285 gnd.n2269 10.4732
R11382 gnd.n2253 gnd.n2237 10.4732
R11383 gnd.n2221 gnd.n2205 10.4732
R11384 gnd.n2190 gnd.n2174 10.4732
R11385 gnd.n2158 gnd.n2142 10.4732
R11386 gnd.n2126 gnd.n2110 10.4732
R11387 gnd.n2094 gnd.n2078 10.4732
R11388 gnd.n2063 gnd.n2047 10.4732
R11389 gnd.n4724 gnd.n3431 10.1975
R11390 gnd.n4741 gnd.t15 10.1975
R11391 gnd.n4905 gnd.n3365 10.1975
R11392 gnd.n3374 gnd.n3367 10.1975
R11393 gnd.n4971 gnd.t7 10.1975
R11394 gnd.n3302 gnd.n3294 10.1975
R11395 gnd.n1986 gnd.t46 9.87883
R11396 gnd.n7485 gnd.n62 9.73455
R11397 gnd.n2289 gnd.n2288 9.69747
R11398 gnd.n2257 gnd.n2256 9.69747
R11399 gnd.n2225 gnd.n2224 9.69747
R11400 gnd.n2194 gnd.n2193 9.69747
R11401 gnd.n2162 gnd.n2161 9.69747
R11402 gnd.n2130 gnd.n2129 9.69747
R11403 gnd.n2098 gnd.n2097 9.69747
R11404 gnd.n2067 gnd.n2066 9.69747
R11405 gnd.t163 gnd.n4467 9.56018
R11406 gnd.n5322 gnd.t169 9.56018
R11407 gnd.n5110 gnd.t76 9.56018
R11408 gnd.n5906 gnd.n2675 9.45599
R11409 gnd.n3126 gnd.n2878 9.45599
R11410 gnd.n2295 gnd.n2294 9.45567
R11411 gnd.n2263 gnd.n2262 9.45567
R11412 gnd.n2231 gnd.n2230 9.45567
R11413 gnd.n2200 gnd.n2199 9.45567
R11414 gnd.n2168 gnd.n2167 9.45567
R11415 gnd.n2136 gnd.n2135 9.45567
R11416 gnd.n2104 gnd.n2103 9.45567
R11417 gnd.n2073 gnd.n2072 9.45567
R11418 gnd.n1281 gnd.n1280 9.39724
R11419 gnd.n2294 gnd.n2293 9.3005
R11420 gnd.n2267 gnd.n2266 9.3005
R11421 gnd.n2288 gnd.n2287 9.3005
R11422 gnd.n2286 gnd.n2285 9.3005
R11423 gnd.n2271 gnd.n2270 9.3005
R11424 gnd.n2280 gnd.n2279 9.3005
R11425 gnd.n2278 gnd.n2277 9.3005
R11426 gnd.n2262 gnd.n2261 9.3005
R11427 gnd.n2235 gnd.n2234 9.3005
R11428 gnd.n2256 gnd.n2255 9.3005
R11429 gnd.n2254 gnd.n2253 9.3005
R11430 gnd.n2239 gnd.n2238 9.3005
R11431 gnd.n2248 gnd.n2247 9.3005
R11432 gnd.n2246 gnd.n2245 9.3005
R11433 gnd.n2230 gnd.n2229 9.3005
R11434 gnd.n2203 gnd.n2202 9.3005
R11435 gnd.n2224 gnd.n2223 9.3005
R11436 gnd.n2222 gnd.n2221 9.3005
R11437 gnd.n2207 gnd.n2206 9.3005
R11438 gnd.n2216 gnd.n2215 9.3005
R11439 gnd.n2214 gnd.n2213 9.3005
R11440 gnd.n2199 gnd.n2198 9.3005
R11441 gnd.n2172 gnd.n2171 9.3005
R11442 gnd.n2193 gnd.n2192 9.3005
R11443 gnd.n2191 gnd.n2190 9.3005
R11444 gnd.n2176 gnd.n2175 9.3005
R11445 gnd.n2185 gnd.n2184 9.3005
R11446 gnd.n2183 gnd.n2182 9.3005
R11447 gnd.n2167 gnd.n2166 9.3005
R11448 gnd.n2140 gnd.n2139 9.3005
R11449 gnd.n2161 gnd.n2160 9.3005
R11450 gnd.n2159 gnd.n2158 9.3005
R11451 gnd.n2144 gnd.n2143 9.3005
R11452 gnd.n2153 gnd.n2152 9.3005
R11453 gnd.n2151 gnd.n2150 9.3005
R11454 gnd.n2135 gnd.n2134 9.3005
R11455 gnd.n2108 gnd.n2107 9.3005
R11456 gnd.n2129 gnd.n2128 9.3005
R11457 gnd.n2127 gnd.n2126 9.3005
R11458 gnd.n2112 gnd.n2111 9.3005
R11459 gnd.n2121 gnd.n2120 9.3005
R11460 gnd.n2119 gnd.n2118 9.3005
R11461 gnd.n2103 gnd.n2102 9.3005
R11462 gnd.n2076 gnd.n2075 9.3005
R11463 gnd.n2097 gnd.n2096 9.3005
R11464 gnd.n2095 gnd.n2094 9.3005
R11465 gnd.n2080 gnd.n2079 9.3005
R11466 gnd.n2089 gnd.n2088 9.3005
R11467 gnd.n2087 gnd.n2086 9.3005
R11468 gnd.n2072 gnd.n2071 9.3005
R11469 gnd.n2045 gnd.n2044 9.3005
R11470 gnd.n2066 gnd.n2065 9.3005
R11471 gnd.n2064 gnd.n2063 9.3005
R11472 gnd.n2049 gnd.n2048 9.3005
R11473 gnd.n2058 gnd.n2057 9.3005
R11474 gnd.n2056 gnd.n2055 9.3005
R11475 gnd.n6192 gnd.n6191 9.3005
R11476 gnd.n6190 gnd.n6158 9.3005
R11477 gnd.n6189 gnd.n6188 9.3005
R11478 gnd.n6185 gnd.n6159 9.3005
R11479 gnd.n6182 gnd.n6160 9.3005
R11480 gnd.n6181 gnd.n6161 9.3005
R11481 gnd.n6178 gnd.n6162 9.3005
R11482 gnd.n6177 gnd.n6163 9.3005
R11483 gnd.n6174 gnd.n6164 9.3005
R11484 gnd.n6173 gnd.n6165 9.3005
R11485 gnd.n6170 gnd.n6166 9.3005
R11486 gnd.n6169 gnd.n6167 9.3005
R11487 gnd.n1055 gnd.n1054 9.3005
R11488 gnd.n6200 gnd.n6199 9.3005
R11489 gnd.n6201 gnd.n1053 9.3005
R11490 gnd.n6203 gnd.n6202 9.3005
R11491 gnd.n6193 gnd.n6157 9.3005
R11492 gnd.n1702 gnd.n1701 9.3005
R11493 gnd.n1406 gnd.n1405 9.3005
R11494 gnd.n1729 gnd.n1728 9.3005
R11495 gnd.n1730 gnd.n1404 9.3005
R11496 gnd.n1734 gnd.n1731 9.3005
R11497 gnd.n1733 gnd.n1732 9.3005
R11498 gnd.n1378 gnd.n1377 9.3005
R11499 gnd.n1759 gnd.n1758 9.3005
R11500 gnd.n1760 gnd.n1376 9.3005
R11501 gnd.n1762 gnd.n1761 9.3005
R11502 gnd.n1356 gnd.n1355 9.3005
R11503 gnd.n1790 gnd.n1789 9.3005
R11504 gnd.n1791 gnd.n1354 9.3005
R11505 gnd.n1799 gnd.n1792 9.3005
R11506 gnd.n1798 gnd.n1793 9.3005
R11507 gnd.n1797 gnd.n1795 9.3005
R11508 gnd.n1794 gnd.n1303 9.3005
R11509 gnd.n1847 gnd.n1304 9.3005
R11510 gnd.n1846 gnd.n1305 9.3005
R11511 gnd.n1845 gnd.n1306 9.3005
R11512 gnd.n1325 gnd.n1307 9.3005
R11513 gnd.n1327 gnd.n1326 9.3005
R11514 gnd.n1225 gnd.n1224 9.3005
R11515 gnd.n1885 gnd.n1884 9.3005
R11516 gnd.n1886 gnd.n1223 9.3005
R11517 gnd.n1890 gnd.n1887 9.3005
R11518 gnd.n1889 gnd.n1888 9.3005
R11519 gnd.n1198 gnd.n1197 9.3005
R11520 gnd.n1925 gnd.n1924 9.3005
R11521 gnd.n1926 gnd.n1196 9.3005
R11522 gnd.n1930 gnd.n1927 9.3005
R11523 gnd.n1929 gnd.n1928 9.3005
R11524 gnd.n1172 gnd.n1171 9.3005
R11525 gnd.n1999 gnd.n1998 9.3005
R11526 gnd.n2000 gnd.n1170 9.3005
R11527 gnd.n2008 gnd.n2001 9.3005
R11528 gnd.n2007 gnd.n2002 9.3005
R11529 gnd.n2006 gnd.n2004 9.3005
R11530 gnd.n2003 gnd.n983 9.3005
R11531 gnd.n6244 gnd.n984 9.3005
R11532 gnd.n6243 gnd.n985 9.3005
R11533 gnd.n6242 gnd.n986 9.3005
R11534 gnd.n1008 gnd.n987 9.3005
R11535 gnd.n1009 gnd.n1007 9.3005
R11536 gnd.n6230 gnd.n1010 9.3005
R11537 gnd.n6229 gnd.n1011 9.3005
R11538 gnd.n6228 gnd.n1012 9.3005
R11539 gnd.n1033 gnd.n1013 9.3005
R11540 gnd.n1034 gnd.n1032 9.3005
R11541 gnd.n6216 gnd.n1035 9.3005
R11542 gnd.n6215 gnd.n1036 9.3005
R11543 gnd.n6214 gnd.n1037 9.3005
R11544 gnd.n6156 gnd.n1038 9.3005
R11545 gnd.n1703 gnd.n1700 9.3005
R11546 gnd.n1485 gnd.n1444 9.3005
R11547 gnd.n1480 gnd.n1479 9.3005
R11548 gnd.n1478 gnd.n1445 9.3005
R11549 gnd.n1477 gnd.n1476 9.3005
R11550 gnd.n1473 gnd.n1446 9.3005
R11551 gnd.n1470 gnd.n1469 9.3005
R11552 gnd.n1468 gnd.n1447 9.3005
R11553 gnd.n1467 gnd.n1466 9.3005
R11554 gnd.n1463 gnd.n1448 9.3005
R11555 gnd.n1460 gnd.n1459 9.3005
R11556 gnd.n1458 gnd.n1449 9.3005
R11557 gnd.n1457 gnd.n1456 9.3005
R11558 gnd.n1453 gnd.n1451 9.3005
R11559 gnd.n1450 gnd.n1430 9.3005
R11560 gnd.n1697 gnd.n1429 9.3005
R11561 gnd.n1699 gnd.n1698 9.3005
R11562 gnd.n1487 gnd.n1486 9.3005
R11563 gnd.n1710 gnd.n1416 9.3005
R11564 gnd.n1717 gnd.n1417 9.3005
R11565 gnd.n1719 gnd.n1718 9.3005
R11566 gnd.n1720 gnd.n1397 9.3005
R11567 gnd.n1739 gnd.n1738 9.3005
R11568 gnd.n1741 gnd.n1389 9.3005
R11569 gnd.n1748 gnd.n1391 9.3005
R11570 gnd.n1749 gnd.n1386 9.3005
R11571 gnd.n1751 gnd.n1750 9.3005
R11572 gnd.n1387 gnd.n1372 9.3005
R11573 gnd.n1767 gnd.n1370 9.3005
R11574 gnd.n1771 gnd.n1770 9.3005
R11575 gnd.n1769 gnd.n1346 9.3005
R11576 gnd.n1806 gnd.n1345 9.3005
R11577 gnd.n1809 gnd.n1808 9.3005
R11578 gnd.n1342 gnd.n1341 9.3005
R11579 gnd.n1815 gnd.n1343 9.3005
R11580 gnd.n1817 gnd.n1816 9.3005
R11581 gnd.n1819 gnd.n1340 9.3005
R11582 gnd.n1822 gnd.n1821 9.3005
R11583 gnd.n1825 gnd.n1823 9.3005
R11584 gnd.n1827 gnd.n1826 9.3005
R11585 gnd.n1833 gnd.n1828 9.3005
R11586 gnd.n1832 gnd.n1831 9.3005
R11587 gnd.n1216 gnd.n1215 9.3005
R11588 gnd.n1899 gnd.n1898 9.3005
R11589 gnd.n1900 gnd.n1209 9.3005
R11590 gnd.n1908 gnd.n1208 9.3005
R11591 gnd.n1911 gnd.n1910 9.3005
R11592 gnd.n1913 gnd.n1912 9.3005
R11593 gnd.n1916 gnd.n1191 9.3005
R11594 gnd.n1914 gnd.n1189 9.3005
R11595 gnd.n1936 gnd.n1187 9.3005
R11596 gnd.n1940 gnd.n1939 9.3005
R11597 gnd.n1938 gnd.n1162 9.3005
R11598 gnd.n2015 gnd.n1161 9.3005
R11599 gnd.n2018 gnd.n2017 9.3005
R11600 gnd.n1158 gnd.n1157 9.3005
R11601 gnd.n2022 gnd.n1159 9.3005
R11602 gnd.n2024 gnd.n2023 9.3005
R11603 gnd.n2026 gnd.n1156 9.3005
R11604 gnd.n2029 gnd.n2028 9.3005
R11605 gnd.n2031 gnd.n2030 9.3005
R11606 gnd.n2035 gnd.n2032 9.3005
R11607 gnd.n2037 gnd.n2036 9.3005
R11608 gnd.n2039 gnd.n1153 9.3005
R11609 gnd.n2042 gnd.n2041 9.3005
R11610 gnd.n2300 gnd.n2299 9.3005
R11611 gnd.n2304 gnd.n2301 9.3005
R11612 gnd.n2306 gnd.n2305 9.3005
R11613 gnd.n2310 gnd.n2309 9.3005
R11614 gnd.n1049 gnd.n1047 9.3005
R11615 gnd.n6207 gnd.n6206 9.3005
R11616 gnd.n1708 gnd.n1707 9.3005
R11617 gnd.n1089 gnd.n1086 9.3005
R11618 gnd.n1091 gnd.n1090 9.3005
R11619 gnd.n1094 gnd.n1084 9.3005
R11620 gnd.n1098 gnd.n1097 9.3005
R11621 gnd.n1099 gnd.n1083 9.3005
R11622 gnd.n1101 gnd.n1100 9.3005
R11623 gnd.n1104 gnd.n1082 9.3005
R11624 gnd.n1108 gnd.n1107 9.3005
R11625 gnd.n1109 gnd.n1081 9.3005
R11626 gnd.n1111 gnd.n1110 9.3005
R11627 gnd.n1114 gnd.n1080 9.3005
R11628 gnd.n1118 gnd.n1117 9.3005
R11629 gnd.n1119 gnd.n1079 9.3005
R11630 gnd.n1121 gnd.n1120 9.3005
R11631 gnd.n1124 gnd.n1078 9.3005
R11632 gnd.n1128 gnd.n1127 9.3005
R11633 gnd.n1129 gnd.n1077 9.3005
R11634 gnd.n1131 gnd.n1130 9.3005
R11635 gnd.n1134 gnd.n1076 9.3005
R11636 gnd.n1138 gnd.n1137 9.3005
R11637 gnd.n1139 gnd.n1075 9.3005
R11638 gnd.n1141 gnd.n1140 9.3005
R11639 gnd.n1144 gnd.n1071 9.3005
R11640 gnd.n1147 gnd.n1146 9.3005
R11641 gnd.n1148 gnd.n1070 9.3005
R11642 gnd.n2320 gnd.n2319 9.3005
R11643 gnd.n1088 gnd.n1087 9.3005
R11644 gnd.n1877 gnd.n1861 9.3005
R11645 gnd.n1876 gnd.n1862 9.3005
R11646 gnd.n1875 gnd.n1863 9.3005
R11647 gnd.n1873 gnd.n1864 9.3005
R11648 gnd.n1872 gnd.n1865 9.3005
R11649 gnd.n1870 gnd.n1866 9.3005
R11650 gnd.n1869 gnd.n1867 9.3005
R11651 gnd.n1179 gnd.n1178 9.3005
R11652 gnd.n1948 gnd.n1947 9.3005
R11653 gnd.n1949 gnd.n1177 9.3005
R11654 gnd.n1993 gnd.n1950 9.3005
R11655 gnd.n1992 gnd.n1951 9.3005
R11656 gnd.n1991 gnd.n1952 9.3005
R11657 gnd.n1989 gnd.n1953 9.3005
R11658 gnd.n1988 gnd.n1954 9.3005
R11659 gnd.n1985 gnd.n1955 9.3005
R11660 gnd.n1984 gnd.n1956 9.3005
R11661 gnd.n1981 gnd.n1957 9.3005
R11662 gnd.n1980 gnd.n1958 9.3005
R11663 gnd.n1979 gnd.n1959 9.3005
R11664 gnd.n1976 gnd.n1960 9.3005
R11665 gnd.n1975 gnd.n1961 9.3005
R11666 gnd.n1972 gnd.n1962 9.3005
R11667 gnd.n1971 gnd.n1963 9.3005
R11668 gnd.n1970 gnd.n1964 9.3005
R11669 gnd.n1967 gnd.n1966 9.3005
R11670 gnd.n1965 gnd.n1150 9.3005
R11671 gnd.n2316 gnd.n1149 9.3005
R11672 gnd.n2318 gnd.n2317 9.3005
R11673 gnd.n1618 gnd.n1617 9.3005
R11674 gnd.n1508 gnd.n1507 9.3005
R11675 gnd.n1632 gnd.n1631 9.3005
R11676 gnd.n1633 gnd.n1506 9.3005
R11677 gnd.n1635 gnd.n1634 9.3005
R11678 gnd.n1496 gnd.n1495 9.3005
R11679 gnd.n1648 gnd.n1647 9.3005
R11680 gnd.n1649 gnd.n1494 9.3005
R11681 gnd.n1681 gnd.n1650 9.3005
R11682 gnd.n1680 gnd.n1651 9.3005
R11683 gnd.n1679 gnd.n1652 9.3005
R11684 gnd.n1678 gnd.n1653 9.3005
R11685 gnd.n1675 gnd.n1654 9.3005
R11686 gnd.n1674 gnd.n1655 9.3005
R11687 gnd.n1673 gnd.n1656 9.3005
R11688 gnd.n1671 gnd.n1657 9.3005
R11689 gnd.n1670 gnd.n1658 9.3005
R11690 gnd.n1667 gnd.n1659 9.3005
R11691 gnd.n1666 gnd.n1660 9.3005
R11692 gnd.n1665 gnd.n1661 9.3005
R11693 gnd.n1663 gnd.n1662 9.3005
R11694 gnd.n1362 gnd.n1361 9.3005
R11695 gnd.n1779 gnd.n1778 9.3005
R11696 gnd.n1780 gnd.n1360 9.3005
R11697 gnd.n1784 gnd.n1781 9.3005
R11698 gnd.n1783 gnd.n1782 9.3005
R11699 gnd.n1284 gnd.n1283 9.3005
R11700 gnd.n1859 gnd.n1858 9.3005
R11701 gnd.n1616 gnd.n1517 9.3005
R11702 gnd.n1519 gnd.n1518 9.3005
R11703 gnd.n1563 gnd.n1561 9.3005
R11704 gnd.n1564 gnd.n1560 9.3005
R11705 gnd.n1567 gnd.n1556 9.3005
R11706 gnd.n1568 gnd.n1555 9.3005
R11707 gnd.n1571 gnd.n1554 9.3005
R11708 gnd.n1572 gnd.n1553 9.3005
R11709 gnd.n1575 gnd.n1552 9.3005
R11710 gnd.n1576 gnd.n1551 9.3005
R11711 gnd.n1579 gnd.n1550 9.3005
R11712 gnd.n1580 gnd.n1549 9.3005
R11713 gnd.n1583 gnd.n1548 9.3005
R11714 gnd.n1584 gnd.n1547 9.3005
R11715 gnd.n1587 gnd.n1546 9.3005
R11716 gnd.n1588 gnd.n1545 9.3005
R11717 gnd.n1591 gnd.n1544 9.3005
R11718 gnd.n1592 gnd.n1543 9.3005
R11719 gnd.n1595 gnd.n1542 9.3005
R11720 gnd.n1596 gnd.n1541 9.3005
R11721 gnd.n1599 gnd.n1540 9.3005
R11722 gnd.n1600 gnd.n1539 9.3005
R11723 gnd.n1603 gnd.n1538 9.3005
R11724 gnd.n1605 gnd.n1537 9.3005
R11725 gnd.n1606 gnd.n1536 9.3005
R11726 gnd.n1607 gnd.n1535 9.3005
R11727 gnd.n1608 gnd.n1534 9.3005
R11728 gnd.n1615 gnd.n1614 9.3005
R11729 gnd.n1624 gnd.n1623 9.3005
R11730 gnd.n1625 gnd.n1511 9.3005
R11731 gnd.n1627 gnd.n1626 9.3005
R11732 gnd.n1502 gnd.n1501 9.3005
R11733 gnd.n1640 gnd.n1639 9.3005
R11734 gnd.n1641 gnd.n1500 9.3005
R11735 gnd.n1643 gnd.n1642 9.3005
R11736 gnd.n1489 gnd.n1488 9.3005
R11737 gnd.n1686 gnd.n1685 9.3005
R11738 gnd.n1687 gnd.n1443 9.3005
R11739 gnd.n1691 gnd.n1689 9.3005
R11740 gnd.n1690 gnd.n1422 9.3005
R11741 gnd.n1709 gnd.n1421 9.3005
R11742 gnd.n1712 gnd.n1711 9.3005
R11743 gnd.n1415 gnd.n1414 9.3005
R11744 gnd.n1723 gnd.n1721 9.3005
R11745 gnd.n1722 gnd.n1396 9.3005
R11746 gnd.n1740 gnd.n1395 9.3005
R11747 gnd.n1743 gnd.n1742 9.3005
R11748 gnd.n1390 gnd.n1385 9.3005
R11749 gnd.n1753 gnd.n1752 9.3005
R11750 gnd.n1388 gnd.n1368 9.3005
R11751 gnd.n1774 gnd.n1369 9.3005
R11752 gnd.n1773 gnd.n1772 9.3005
R11753 gnd.n1371 gnd.n1347 9.3005
R11754 gnd.n1805 gnd.n1804 9.3005
R11755 gnd.n1807 gnd.n1292 9.3005
R11756 gnd.n1854 gnd.n1293 9.3005
R11757 gnd.n1853 gnd.n1294 9.3005
R11758 gnd.n1852 gnd.n1295 9.3005
R11759 gnd.n1818 gnd.n1296 9.3005
R11760 gnd.n1820 gnd.n1314 9.3005
R11761 gnd.n1840 gnd.n1315 9.3005
R11762 gnd.n1839 gnd.n1316 9.3005
R11763 gnd.n1838 gnd.n1317 9.3005
R11764 gnd.n1829 gnd.n1318 9.3005
R11765 gnd.n1830 gnd.n1217 9.3005
R11766 gnd.n1896 gnd.n1895 9.3005
R11767 gnd.n1897 gnd.n1210 9.3005
R11768 gnd.n1907 gnd.n1906 9.3005
R11769 gnd.n1909 gnd.n1206 9.3005
R11770 gnd.n1919 gnd.n1207 9.3005
R11771 gnd.n1918 gnd.n1917 9.3005
R11772 gnd.n1915 gnd.n1185 9.3005
R11773 gnd.n1943 gnd.n1186 9.3005
R11774 gnd.n1942 gnd.n1941 9.3005
R11775 gnd.n1188 gnd.n1163 9.3005
R11776 gnd.n2014 gnd.n2013 9.3005
R11777 gnd.n2016 gnd.n971 9.3005
R11778 gnd.n6251 gnd.n972 9.3005
R11779 gnd.n6250 gnd.n973 9.3005
R11780 gnd.n6249 gnd.n974 9.3005
R11781 gnd.n2025 gnd.n975 9.3005
R11782 gnd.n2027 gnd.n995 9.3005
R11783 gnd.n6237 gnd.n996 9.3005
R11784 gnd.n6236 gnd.n997 9.3005
R11785 gnd.n6235 gnd.n998 9.3005
R11786 gnd.n2038 gnd.n999 9.3005
R11787 gnd.n2040 gnd.n1021 9.3005
R11788 gnd.n6223 gnd.n1022 9.3005
R11789 gnd.n6222 gnd.n1023 9.3005
R11790 gnd.n6221 gnd.n1024 9.3005
R11791 gnd.n2307 gnd.n1025 9.3005
R11792 gnd.n2308 gnd.n1046 9.3005
R11793 gnd.n6209 gnd.n6208 9.3005
R11794 gnd.n1513 gnd.n1512 9.3005
R11795 gnd.n797 gnd.n796 9.3005
R11796 gnd.n6427 gnd.n6426 9.3005
R11797 gnd.n6428 gnd.n795 9.3005
R11798 gnd.n6430 gnd.n6429 9.3005
R11799 gnd.n791 gnd.n790 9.3005
R11800 gnd.n6437 gnd.n6436 9.3005
R11801 gnd.n6438 gnd.n789 9.3005
R11802 gnd.n6440 gnd.n6439 9.3005
R11803 gnd.n785 gnd.n784 9.3005
R11804 gnd.n6447 gnd.n6446 9.3005
R11805 gnd.n6448 gnd.n783 9.3005
R11806 gnd.n6450 gnd.n6449 9.3005
R11807 gnd.n779 gnd.n778 9.3005
R11808 gnd.n6457 gnd.n6456 9.3005
R11809 gnd.n6458 gnd.n777 9.3005
R11810 gnd.n6460 gnd.n6459 9.3005
R11811 gnd.n773 gnd.n772 9.3005
R11812 gnd.n6467 gnd.n6466 9.3005
R11813 gnd.n6468 gnd.n771 9.3005
R11814 gnd.n6470 gnd.n6469 9.3005
R11815 gnd.n767 gnd.n766 9.3005
R11816 gnd.n6477 gnd.n6476 9.3005
R11817 gnd.n6478 gnd.n765 9.3005
R11818 gnd.n6480 gnd.n6479 9.3005
R11819 gnd.n761 gnd.n760 9.3005
R11820 gnd.n6487 gnd.n6486 9.3005
R11821 gnd.n6488 gnd.n759 9.3005
R11822 gnd.n6490 gnd.n6489 9.3005
R11823 gnd.n755 gnd.n754 9.3005
R11824 gnd.n6497 gnd.n6496 9.3005
R11825 gnd.n6498 gnd.n753 9.3005
R11826 gnd.n6500 gnd.n6499 9.3005
R11827 gnd.n749 gnd.n748 9.3005
R11828 gnd.n6507 gnd.n6506 9.3005
R11829 gnd.n6508 gnd.n747 9.3005
R11830 gnd.n6510 gnd.n6509 9.3005
R11831 gnd.n743 gnd.n742 9.3005
R11832 gnd.n6517 gnd.n6516 9.3005
R11833 gnd.n6518 gnd.n741 9.3005
R11834 gnd.n6520 gnd.n6519 9.3005
R11835 gnd.n737 gnd.n736 9.3005
R11836 gnd.n6527 gnd.n6526 9.3005
R11837 gnd.n6528 gnd.n735 9.3005
R11838 gnd.n6530 gnd.n6529 9.3005
R11839 gnd.n731 gnd.n730 9.3005
R11840 gnd.n6537 gnd.n6536 9.3005
R11841 gnd.n6538 gnd.n729 9.3005
R11842 gnd.n6540 gnd.n6539 9.3005
R11843 gnd.n725 gnd.n724 9.3005
R11844 gnd.n6547 gnd.n6546 9.3005
R11845 gnd.n6548 gnd.n723 9.3005
R11846 gnd.n6550 gnd.n6549 9.3005
R11847 gnd.n719 gnd.n718 9.3005
R11848 gnd.n6557 gnd.n6556 9.3005
R11849 gnd.n6558 gnd.n717 9.3005
R11850 gnd.n6560 gnd.n6559 9.3005
R11851 gnd.n713 gnd.n712 9.3005
R11852 gnd.n6567 gnd.n6566 9.3005
R11853 gnd.n6568 gnd.n711 9.3005
R11854 gnd.n6570 gnd.n6569 9.3005
R11855 gnd.n707 gnd.n706 9.3005
R11856 gnd.n6577 gnd.n6576 9.3005
R11857 gnd.n6578 gnd.n705 9.3005
R11858 gnd.n6580 gnd.n6579 9.3005
R11859 gnd.n701 gnd.n700 9.3005
R11860 gnd.n6587 gnd.n6586 9.3005
R11861 gnd.n6588 gnd.n699 9.3005
R11862 gnd.n6590 gnd.n6589 9.3005
R11863 gnd.n695 gnd.n694 9.3005
R11864 gnd.n6597 gnd.n6596 9.3005
R11865 gnd.n6598 gnd.n693 9.3005
R11866 gnd.n6600 gnd.n6599 9.3005
R11867 gnd.n689 gnd.n688 9.3005
R11868 gnd.n6607 gnd.n6606 9.3005
R11869 gnd.n6608 gnd.n687 9.3005
R11870 gnd.n6610 gnd.n6609 9.3005
R11871 gnd.n683 gnd.n682 9.3005
R11872 gnd.n6617 gnd.n6616 9.3005
R11873 gnd.n6618 gnd.n681 9.3005
R11874 gnd.n6620 gnd.n6619 9.3005
R11875 gnd.n677 gnd.n676 9.3005
R11876 gnd.n6627 gnd.n6626 9.3005
R11877 gnd.n6628 gnd.n675 9.3005
R11878 gnd.n6630 gnd.n6629 9.3005
R11879 gnd.n671 gnd.n670 9.3005
R11880 gnd.n6637 gnd.n6636 9.3005
R11881 gnd.n6638 gnd.n669 9.3005
R11882 gnd.n6640 gnd.n6639 9.3005
R11883 gnd.n665 gnd.n664 9.3005
R11884 gnd.n6647 gnd.n6646 9.3005
R11885 gnd.n6648 gnd.n663 9.3005
R11886 gnd.n6650 gnd.n6649 9.3005
R11887 gnd.n659 gnd.n658 9.3005
R11888 gnd.n6657 gnd.n6656 9.3005
R11889 gnd.n6658 gnd.n657 9.3005
R11890 gnd.n6660 gnd.n6659 9.3005
R11891 gnd.n653 gnd.n652 9.3005
R11892 gnd.n6667 gnd.n6666 9.3005
R11893 gnd.n6668 gnd.n651 9.3005
R11894 gnd.n6670 gnd.n6669 9.3005
R11895 gnd.n647 gnd.n646 9.3005
R11896 gnd.n6677 gnd.n6676 9.3005
R11897 gnd.n6678 gnd.n645 9.3005
R11898 gnd.n6680 gnd.n6679 9.3005
R11899 gnd.n641 gnd.n640 9.3005
R11900 gnd.n6687 gnd.n6686 9.3005
R11901 gnd.n6688 gnd.n639 9.3005
R11902 gnd.n6690 gnd.n6689 9.3005
R11903 gnd.n635 gnd.n634 9.3005
R11904 gnd.n6697 gnd.n6696 9.3005
R11905 gnd.n6698 gnd.n633 9.3005
R11906 gnd.n6700 gnd.n6699 9.3005
R11907 gnd.n629 gnd.n628 9.3005
R11908 gnd.n6707 gnd.n6706 9.3005
R11909 gnd.n6708 gnd.n627 9.3005
R11910 gnd.n6710 gnd.n6709 9.3005
R11911 gnd.n623 gnd.n622 9.3005
R11912 gnd.n6717 gnd.n6716 9.3005
R11913 gnd.n6718 gnd.n621 9.3005
R11914 gnd.n6720 gnd.n6719 9.3005
R11915 gnd.n617 gnd.n616 9.3005
R11916 gnd.n6727 gnd.n6726 9.3005
R11917 gnd.n6728 gnd.n615 9.3005
R11918 gnd.n6730 gnd.n6729 9.3005
R11919 gnd.n611 gnd.n610 9.3005
R11920 gnd.n6737 gnd.n6736 9.3005
R11921 gnd.n6738 gnd.n609 9.3005
R11922 gnd.n6740 gnd.n6739 9.3005
R11923 gnd.n605 gnd.n604 9.3005
R11924 gnd.n6747 gnd.n6746 9.3005
R11925 gnd.n6748 gnd.n603 9.3005
R11926 gnd.n6750 gnd.n6749 9.3005
R11927 gnd.n599 gnd.n598 9.3005
R11928 gnd.n6757 gnd.n6756 9.3005
R11929 gnd.n6758 gnd.n597 9.3005
R11930 gnd.n6760 gnd.n6759 9.3005
R11931 gnd.n593 gnd.n592 9.3005
R11932 gnd.n6767 gnd.n6766 9.3005
R11933 gnd.n6768 gnd.n591 9.3005
R11934 gnd.n6770 gnd.n6769 9.3005
R11935 gnd.n587 gnd.n586 9.3005
R11936 gnd.n6777 gnd.n6776 9.3005
R11937 gnd.n6778 gnd.n585 9.3005
R11938 gnd.n6780 gnd.n6779 9.3005
R11939 gnd.n581 gnd.n580 9.3005
R11940 gnd.n6787 gnd.n6786 9.3005
R11941 gnd.n6788 gnd.n579 9.3005
R11942 gnd.n6790 gnd.n6789 9.3005
R11943 gnd.n575 gnd.n574 9.3005
R11944 gnd.n6797 gnd.n6796 9.3005
R11945 gnd.n6798 gnd.n573 9.3005
R11946 gnd.n6800 gnd.n6799 9.3005
R11947 gnd.n569 gnd.n568 9.3005
R11948 gnd.n6807 gnd.n6806 9.3005
R11949 gnd.n6808 gnd.n567 9.3005
R11950 gnd.n6810 gnd.n6809 9.3005
R11951 gnd.n563 gnd.n562 9.3005
R11952 gnd.n6817 gnd.n6816 9.3005
R11953 gnd.n6818 gnd.n561 9.3005
R11954 gnd.n6820 gnd.n6819 9.3005
R11955 gnd.n557 gnd.n556 9.3005
R11956 gnd.n6827 gnd.n6826 9.3005
R11957 gnd.n6828 gnd.n555 9.3005
R11958 gnd.n6830 gnd.n6829 9.3005
R11959 gnd.n551 gnd.n550 9.3005
R11960 gnd.n6837 gnd.n6836 9.3005
R11961 gnd.n6838 gnd.n549 9.3005
R11962 gnd.n6840 gnd.n6839 9.3005
R11963 gnd.n545 gnd.n544 9.3005
R11964 gnd.n6847 gnd.n6846 9.3005
R11965 gnd.n6848 gnd.n543 9.3005
R11966 gnd.n6850 gnd.n6849 9.3005
R11967 gnd.n539 gnd.n538 9.3005
R11968 gnd.n6857 gnd.n6856 9.3005
R11969 gnd.n6858 gnd.n537 9.3005
R11970 gnd.n6860 gnd.n6859 9.3005
R11971 gnd.n533 gnd.n532 9.3005
R11972 gnd.n6867 gnd.n6866 9.3005
R11973 gnd.n6868 gnd.n531 9.3005
R11974 gnd.n6870 gnd.n6869 9.3005
R11975 gnd.n527 gnd.n526 9.3005
R11976 gnd.n6877 gnd.n6876 9.3005
R11977 gnd.n6878 gnd.n525 9.3005
R11978 gnd.n6880 gnd.n6879 9.3005
R11979 gnd.n521 gnd.n520 9.3005
R11980 gnd.n6887 gnd.n6886 9.3005
R11981 gnd.n6888 gnd.n519 9.3005
R11982 gnd.n6890 gnd.n6889 9.3005
R11983 gnd.n515 gnd.n514 9.3005
R11984 gnd.n6897 gnd.n6896 9.3005
R11985 gnd.n6898 gnd.n513 9.3005
R11986 gnd.n6901 gnd.n6900 9.3005
R11987 gnd.n6899 gnd.n509 9.3005
R11988 gnd.n6907 gnd.n508 9.3005
R11989 gnd.n6909 gnd.n6908 9.3005
R11990 gnd.n504 gnd.n503 9.3005
R11991 gnd.n6918 gnd.n6917 9.3005
R11992 gnd.n6919 gnd.n502 9.3005
R11993 gnd.n6921 gnd.n6920 9.3005
R11994 gnd.n498 gnd.n497 9.3005
R11995 gnd.n6928 gnd.n6927 9.3005
R11996 gnd.n6929 gnd.n496 9.3005
R11997 gnd.n6931 gnd.n6930 9.3005
R11998 gnd.n492 gnd.n491 9.3005
R11999 gnd.n6938 gnd.n6937 9.3005
R12000 gnd.n6939 gnd.n490 9.3005
R12001 gnd.n6941 gnd.n6940 9.3005
R12002 gnd.n486 gnd.n485 9.3005
R12003 gnd.n6948 gnd.n6947 9.3005
R12004 gnd.n6949 gnd.n484 9.3005
R12005 gnd.n6951 gnd.n6950 9.3005
R12006 gnd.n480 gnd.n479 9.3005
R12007 gnd.n6958 gnd.n6957 9.3005
R12008 gnd.n6959 gnd.n478 9.3005
R12009 gnd.n6961 gnd.n6960 9.3005
R12010 gnd.n474 gnd.n473 9.3005
R12011 gnd.n6968 gnd.n6967 9.3005
R12012 gnd.n6969 gnd.n472 9.3005
R12013 gnd.n6971 gnd.n6970 9.3005
R12014 gnd.n468 gnd.n467 9.3005
R12015 gnd.n6978 gnd.n6977 9.3005
R12016 gnd.n6979 gnd.n466 9.3005
R12017 gnd.n6981 gnd.n6980 9.3005
R12018 gnd.n462 gnd.n461 9.3005
R12019 gnd.n6988 gnd.n6987 9.3005
R12020 gnd.n6989 gnd.n460 9.3005
R12021 gnd.n6991 gnd.n6990 9.3005
R12022 gnd.n456 gnd.n455 9.3005
R12023 gnd.n6998 gnd.n6997 9.3005
R12024 gnd.n6999 gnd.n454 9.3005
R12025 gnd.n7001 gnd.n7000 9.3005
R12026 gnd.n450 gnd.n449 9.3005
R12027 gnd.n7008 gnd.n7007 9.3005
R12028 gnd.n7009 gnd.n448 9.3005
R12029 gnd.n7011 gnd.n7010 9.3005
R12030 gnd.n444 gnd.n443 9.3005
R12031 gnd.n7018 gnd.n7017 9.3005
R12032 gnd.n7019 gnd.n442 9.3005
R12033 gnd.n7021 gnd.n7020 9.3005
R12034 gnd.n438 gnd.n437 9.3005
R12035 gnd.n7028 gnd.n7027 9.3005
R12036 gnd.n7029 gnd.n436 9.3005
R12037 gnd.n7031 gnd.n7030 9.3005
R12038 gnd.n432 gnd.n431 9.3005
R12039 gnd.n7038 gnd.n7037 9.3005
R12040 gnd.n7039 gnd.n430 9.3005
R12041 gnd.n7041 gnd.n7040 9.3005
R12042 gnd.n426 gnd.n425 9.3005
R12043 gnd.n7048 gnd.n7047 9.3005
R12044 gnd.n7049 gnd.n424 9.3005
R12045 gnd.n7051 gnd.n7050 9.3005
R12046 gnd.n420 gnd.n419 9.3005
R12047 gnd.n7058 gnd.n7057 9.3005
R12048 gnd.n7059 gnd.n418 9.3005
R12049 gnd.n7061 gnd.n7060 9.3005
R12050 gnd.n414 gnd.n413 9.3005
R12051 gnd.n7068 gnd.n7067 9.3005
R12052 gnd.n7069 gnd.n412 9.3005
R12053 gnd.n7071 gnd.n7070 9.3005
R12054 gnd.n408 gnd.n407 9.3005
R12055 gnd.n7078 gnd.n7077 9.3005
R12056 gnd.n7079 gnd.n406 9.3005
R12057 gnd.n7081 gnd.n7080 9.3005
R12058 gnd.n402 gnd.n401 9.3005
R12059 gnd.n7088 gnd.n7087 9.3005
R12060 gnd.n7089 gnd.n400 9.3005
R12061 gnd.n7091 gnd.n7090 9.3005
R12062 gnd.n396 gnd.n395 9.3005
R12063 gnd.n7098 gnd.n7097 9.3005
R12064 gnd.n7099 gnd.n394 9.3005
R12065 gnd.n7101 gnd.n7100 9.3005
R12066 gnd.n390 gnd.n389 9.3005
R12067 gnd.n7108 gnd.n7107 9.3005
R12068 gnd.n7109 gnd.n388 9.3005
R12069 gnd.n7111 gnd.n7110 9.3005
R12070 gnd.n384 gnd.n383 9.3005
R12071 gnd.n7119 gnd.n7118 9.3005
R12072 gnd.n7120 gnd.n382 9.3005
R12073 gnd.n7123 gnd.n7122 9.3005
R12074 gnd.n6911 gnd.n6910 9.3005
R12075 gnd.n7436 gnd.n108 9.3005
R12076 gnd.n7435 gnd.n110 9.3005
R12077 gnd.n114 gnd.n111 9.3005
R12078 gnd.n7430 gnd.n115 9.3005
R12079 gnd.n7429 gnd.n116 9.3005
R12080 gnd.n7428 gnd.n117 9.3005
R12081 gnd.n121 gnd.n118 9.3005
R12082 gnd.n7423 gnd.n122 9.3005
R12083 gnd.n7422 gnd.n123 9.3005
R12084 gnd.n7421 gnd.n124 9.3005
R12085 gnd.n128 gnd.n125 9.3005
R12086 gnd.n7416 gnd.n129 9.3005
R12087 gnd.n7415 gnd.n130 9.3005
R12088 gnd.n7414 gnd.n131 9.3005
R12089 gnd.n135 gnd.n132 9.3005
R12090 gnd.n7409 gnd.n136 9.3005
R12091 gnd.n7408 gnd.n137 9.3005
R12092 gnd.n7404 gnd.n138 9.3005
R12093 gnd.n142 gnd.n139 9.3005
R12094 gnd.n7399 gnd.n143 9.3005
R12095 gnd.n7398 gnd.n144 9.3005
R12096 gnd.n7397 gnd.n145 9.3005
R12097 gnd.n149 gnd.n146 9.3005
R12098 gnd.n7392 gnd.n150 9.3005
R12099 gnd.n7391 gnd.n151 9.3005
R12100 gnd.n7390 gnd.n152 9.3005
R12101 gnd.n156 gnd.n153 9.3005
R12102 gnd.n7385 gnd.n157 9.3005
R12103 gnd.n7384 gnd.n158 9.3005
R12104 gnd.n7383 gnd.n159 9.3005
R12105 gnd.n163 gnd.n160 9.3005
R12106 gnd.n7378 gnd.n164 9.3005
R12107 gnd.n7377 gnd.n165 9.3005
R12108 gnd.n7376 gnd.n166 9.3005
R12109 gnd.n170 gnd.n167 9.3005
R12110 gnd.n7371 gnd.n171 9.3005
R12111 gnd.n7370 gnd.n7369 9.3005
R12112 gnd.n7368 gnd.n174 9.3005
R12113 gnd.n7438 gnd.n7437 9.3005
R12114 gnd.n3043 gnd.n3042 9.3005
R12115 gnd.n3077 gnd.n3044 9.3005
R12116 gnd.n3076 gnd.n3045 9.3005
R12117 gnd.n3075 gnd.n3046 9.3005
R12118 gnd.n3073 gnd.n3047 9.3005
R12119 gnd.n3072 gnd.n3048 9.3005
R12120 gnd.n3070 gnd.n3049 9.3005
R12121 gnd.n3069 gnd.n3050 9.3005
R12122 gnd.n3068 gnd.n3051 9.3005
R12123 gnd.n3066 gnd.n3052 9.3005
R12124 gnd.n3065 gnd.n3053 9.3005
R12125 gnd.n3063 gnd.n3054 9.3005
R12126 gnd.n3062 gnd.n3055 9.3005
R12127 gnd.n3061 gnd.n3056 9.3005
R12128 gnd.n3059 gnd.n3058 9.3005
R12129 gnd.n3057 gnd.n2943 9.3005
R12130 gnd.n5586 gnd.n2944 9.3005
R12131 gnd.n5587 gnd.n2942 9.3005
R12132 gnd.n5590 gnd.n5589 9.3005
R12133 gnd.n5591 gnd.n2941 9.3005
R12134 gnd.n5595 gnd.n5592 9.3005
R12135 gnd.n5594 gnd.n5593 9.3005
R12136 gnd.n2935 gnd.n2934 9.3005
R12137 gnd.n5613 gnd.n5612 9.3005
R12138 gnd.n5614 gnd.n2933 9.3005
R12139 gnd.n5616 gnd.n5615 9.3005
R12140 gnd.n296 gnd.n295 9.3005
R12141 gnd.n7177 gnd.n297 9.3005
R12142 gnd.n7176 gnd.n298 9.3005
R12143 gnd.n7175 gnd.n299 9.3005
R12144 gnd.n309 gnd.n300 9.3005
R12145 gnd.n313 gnd.n312 9.3005
R12146 gnd.n314 gnd.n308 9.3005
R12147 gnd.n7160 gnd.n315 9.3005
R12148 gnd.n7159 gnd.n316 9.3005
R12149 gnd.n7158 gnd.n317 9.3005
R12150 gnd.n7155 gnd.n318 9.3005
R12151 gnd.n7154 gnd.n319 9.3005
R12152 gnd.n341 gnd.n320 9.3005
R12153 gnd.n345 gnd.n344 9.3005
R12154 gnd.n346 gnd.n340 9.3005
R12155 gnd.n7140 gnd.n347 9.3005
R12156 gnd.n7139 gnd.n348 9.3005
R12157 gnd.n7138 gnd.n349 9.3005
R12158 gnd.n7135 gnd.n350 9.3005
R12159 gnd.n7134 gnd.n351 9.3005
R12160 gnd.n362 gnd.n352 9.3005
R12161 gnd.n361 gnd.n353 9.3005
R12162 gnd.n358 gnd.n354 9.3005
R12163 gnd.n357 gnd.n356 9.3005
R12164 gnd.n355 gnd.n178 9.3005
R12165 gnd.n7365 gnd.n177 9.3005
R12166 gnd.n7367 gnd.n7366 9.3005
R12167 gnd.n2871 gnd.n2869 9.3005
R12168 gnd.n5701 gnd.n5700 9.3005
R12169 gnd.n5702 gnd.n2863 9.3005
R12170 gnd.n5705 gnd.n2862 9.3005
R12171 gnd.n5706 gnd.n2861 9.3005
R12172 gnd.n5709 gnd.n2860 9.3005
R12173 gnd.n5710 gnd.n2859 9.3005
R12174 gnd.n5713 gnd.n2858 9.3005
R12175 gnd.n5714 gnd.n2857 9.3005
R12176 gnd.n5717 gnd.n2856 9.3005
R12177 gnd.n5718 gnd.n2855 9.3005
R12178 gnd.n5721 gnd.n2854 9.3005
R12179 gnd.n5722 gnd.n2853 9.3005
R12180 gnd.n5725 gnd.n2852 9.3005
R12181 gnd.n5726 gnd.n2851 9.3005
R12182 gnd.n5729 gnd.n2850 9.3005
R12183 gnd.n5730 gnd.n2849 9.3005
R12184 gnd.n5733 gnd.n2848 9.3005
R12185 gnd.n5734 gnd.n2847 9.3005
R12186 gnd.n5737 gnd.n2846 9.3005
R12187 gnd.n5739 gnd.n2840 9.3005
R12188 gnd.n5742 gnd.n2839 9.3005
R12189 gnd.n5743 gnd.n2838 9.3005
R12190 gnd.n5746 gnd.n2837 9.3005
R12191 gnd.n5747 gnd.n2836 9.3005
R12192 gnd.n5750 gnd.n2835 9.3005
R12193 gnd.n5751 gnd.n2834 9.3005
R12194 gnd.n5754 gnd.n2833 9.3005
R12195 gnd.n5755 gnd.n2832 9.3005
R12196 gnd.n5758 gnd.n2831 9.3005
R12197 gnd.n5759 gnd.n2830 9.3005
R12198 gnd.n5762 gnd.n2829 9.3005
R12199 gnd.n5764 gnd.n2828 9.3005
R12200 gnd.n5765 gnd.n2827 9.3005
R12201 gnd.n5766 gnd.n2826 9.3005
R12202 gnd.n5767 gnd.n2825 9.3005
R12203 gnd.n5699 gnd.n2868 9.3005
R12204 gnd.n5698 gnd.n5697 9.3005
R12205 gnd.n3039 gnd.n3038 9.3005
R12206 gnd.n3017 gnd.n3016 9.3005
R12207 gnd.n5494 gnd.n5493 9.3005
R12208 gnd.n5495 gnd.n3015 9.3005
R12209 gnd.n5499 gnd.n5496 9.3005
R12210 gnd.n5498 gnd.n5497 9.3005
R12211 gnd.n2988 gnd.n2987 9.3005
R12212 gnd.n5525 gnd.n5524 9.3005
R12213 gnd.n5526 gnd.n2986 9.3005
R12214 gnd.n5530 gnd.n5527 9.3005
R12215 gnd.n5529 gnd.n5528 9.3005
R12216 gnd.n2960 gnd.n2959 9.3005
R12217 gnd.n5564 gnd.n5563 9.3005
R12218 gnd.n5565 gnd.n2958 9.3005
R12219 gnd.n5569 gnd.n5566 9.3005
R12220 gnd.n5568 gnd.n5567 9.3005
R12221 gnd.n2908 gnd.n2907 9.3005
R12222 gnd.n5654 gnd.n5653 9.3005
R12223 gnd.n5655 gnd.n2906 9.3005
R12224 gnd.n5657 gnd.n5656 9.3005
R12225 gnd.n270 gnd.n263 9.3005
R12226 gnd.n250 gnd.n249 9.3005
R12227 gnd.n7218 gnd.n7217 9.3005
R12228 gnd.n7219 gnd.n248 9.3005
R12229 gnd.n7221 gnd.n7220 9.3005
R12230 gnd.n234 gnd.n233 9.3005
R12231 gnd.n7234 gnd.n7233 9.3005
R12232 gnd.n7235 gnd.n232 9.3005
R12233 gnd.n7237 gnd.n7236 9.3005
R12234 gnd.n220 gnd.n219 9.3005
R12235 gnd.n7250 gnd.n7249 9.3005
R12236 gnd.n7251 gnd.n218 9.3005
R12237 gnd.n7253 gnd.n7252 9.3005
R12238 gnd.n204 gnd.n203 9.3005
R12239 gnd.n7266 gnd.n7265 9.3005
R12240 gnd.n7267 gnd.n202 9.3005
R12241 gnd.n7269 gnd.n7268 9.3005
R12242 gnd.n187 gnd.n186 9.3005
R12243 gnd.n7357 gnd.n7356 9.3005
R12244 gnd.n7358 gnd.n185 9.3005
R12245 gnd.n7360 gnd.n7359 9.3005
R12246 gnd.n107 gnd.n106 9.3005
R12247 gnd.n7440 gnd.n7439 9.3005
R12248 gnd.n3037 gnd.n3036 9.3005
R12249 gnd.n7204 gnd.n268 9.3005
R12250 gnd.n7205 gnd.n7204 9.3005
R12251 gnd.n3923 gnd.n3842 9.3005
R12252 gnd.n3922 gnd.n3848 9.3005
R12253 gnd.n3851 gnd.n3849 9.3005
R12254 gnd.n3918 gnd.n3852 9.3005
R12255 gnd.n3917 gnd.n3853 9.3005
R12256 gnd.n3916 gnd.n3854 9.3005
R12257 gnd.n3857 gnd.n3855 9.3005
R12258 gnd.n3912 gnd.n3858 9.3005
R12259 gnd.n3911 gnd.n3859 9.3005
R12260 gnd.n3910 gnd.n3860 9.3005
R12261 gnd.n3863 gnd.n3861 9.3005
R12262 gnd.n3906 gnd.n3864 9.3005
R12263 gnd.n3905 gnd.n3865 9.3005
R12264 gnd.n3904 gnd.n3866 9.3005
R12265 gnd.n3869 gnd.n3867 9.3005
R12266 gnd.n3900 gnd.n3870 9.3005
R12267 gnd.n3899 gnd.n3871 9.3005
R12268 gnd.n3898 gnd.n3872 9.3005
R12269 gnd.n3875 gnd.n3873 9.3005
R12270 gnd.n3894 gnd.n3876 9.3005
R12271 gnd.n3893 gnd.n3877 9.3005
R12272 gnd.n3892 gnd.n3878 9.3005
R12273 gnd.n3881 gnd.n3879 9.3005
R12274 gnd.n3888 gnd.n3882 9.3005
R12275 gnd.n3887 gnd.n3883 9.3005
R12276 gnd.n3886 gnd.n3884 9.3005
R12277 gnd.n3525 gnd.n3524 9.3005
R12278 gnd.n4628 gnd.n4627 9.3005
R12279 gnd.n4629 gnd.n3523 9.3005
R12280 gnd.n4631 gnd.n4630 9.3005
R12281 gnd.n3512 gnd.n3511 9.3005
R12282 gnd.n4644 gnd.n4643 9.3005
R12283 gnd.n4645 gnd.n3510 9.3005
R12284 gnd.n4647 gnd.n4646 9.3005
R12285 gnd.n3499 gnd.n3498 9.3005
R12286 gnd.n4660 gnd.n4659 9.3005
R12287 gnd.n4661 gnd.n3497 9.3005
R12288 gnd.n4663 gnd.n4662 9.3005
R12289 gnd.n3485 gnd.n3484 9.3005
R12290 gnd.n4676 gnd.n4675 9.3005
R12291 gnd.n4677 gnd.n3483 9.3005
R12292 gnd.n4679 gnd.n4678 9.3005
R12293 gnd.n3471 gnd.n3470 9.3005
R12294 gnd.n4692 gnd.n4691 9.3005
R12295 gnd.n4693 gnd.n3469 9.3005
R12296 gnd.n4695 gnd.n4694 9.3005
R12297 gnd.n3458 gnd.n3457 9.3005
R12298 gnd.n4708 gnd.n4707 9.3005
R12299 gnd.n4709 gnd.n3456 9.3005
R12300 gnd.n4713 gnd.n4710 9.3005
R12301 gnd.n4712 gnd.n4711 9.3005
R12302 gnd.n3429 gnd.n3428 9.3005
R12303 gnd.n4841 gnd.n4840 9.3005
R12304 gnd.n4842 gnd.n3427 9.3005
R12305 gnd.n4844 gnd.n4843 9.3005
R12306 gnd.n3417 gnd.n3416 9.3005
R12307 gnd.n4857 gnd.n4856 9.3005
R12308 gnd.n4858 gnd.n3415 9.3005
R12309 gnd.n4860 gnd.n4859 9.3005
R12310 gnd.n3404 gnd.n3403 9.3005
R12311 gnd.n4873 gnd.n4872 9.3005
R12312 gnd.n4874 gnd.n3402 9.3005
R12313 gnd.n4876 gnd.n4875 9.3005
R12314 gnd.n3392 gnd.n3391 9.3005
R12315 gnd.n4889 gnd.n4888 9.3005
R12316 gnd.n4890 gnd.n3390 9.3005
R12317 gnd.n4894 gnd.n4891 9.3005
R12318 gnd.n4893 gnd.n4892 9.3005
R12319 gnd.n3363 gnd.n3362 9.3005
R12320 gnd.n5018 gnd.n5017 9.3005
R12321 gnd.n5019 gnd.n3361 9.3005
R12322 gnd.n5021 gnd.n5020 9.3005
R12323 gnd.n3350 gnd.n3349 9.3005
R12324 gnd.n5034 gnd.n5033 9.3005
R12325 gnd.n5035 gnd.n3348 9.3005
R12326 gnd.n5037 gnd.n5036 9.3005
R12327 gnd.n3335 gnd.n3334 9.3005
R12328 gnd.n5050 gnd.n5049 9.3005
R12329 gnd.n5051 gnd.n3333 9.3005
R12330 gnd.n5053 gnd.n5052 9.3005
R12331 gnd.n3321 gnd.n3320 9.3005
R12332 gnd.n5066 gnd.n5065 9.3005
R12333 gnd.n5067 gnd.n3319 9.3005
R12334 gnd.n5071 gnd.n5068 9.3005
R12335 gnd.n5070 gnd.n5069 9.3005
R12336 gnd.n3291 gnd.n3290 9.3005
R12337 gnd.n5352 gnd.n5351 9.3005
R12338 gnd.n5353 gnd.n3289 9.3005
R12339 gnd.n5355 gnd.n5354 9.3005
R12340 gnd.n3279 gnd.n3278 9.3005
R12341 gnd.n5368 gnd.n5367 9.3005
R12342 gnd.n5369 gnd.n3277 9.3005
R12343 gnd.n5371 gnd.n5370 9.3005
R12344 gnd.n3266 gnd.n3265 9.3005
R12345 gnd.n5384 gnd.n5383 9.3005
R12346 gnd.n5385 gnd.n3264 9.3005
R12347 gnd.n5387 gnd.n5386 9.3005
R12348 gnd.n3253 gnd.n3252 9.3005
R12349 gnd.n5400 gnd.n5399 9.3005
R12350 gnd.n5401 gnd.n3251 9.3005
R12351 gnd.n5403 gnd.n5402 9.3005
R12352 gnd.n3240 gnd.n3239 9.3005
R12353 gnd.n5416 gnd.n5415 9.3005
R12354 gnd.n5417 gnd.n3238 9.3005
R12355 gnd.n5419 gnd.n5418 9.3005
R12356 gnd.n3228 gnd.n3227 9.3005
R12357 gnd.n5434 gnd.n5433 9.3005
R12358 gnd.n5435 gnd.n3226 9.3005
R12359 gnd.n5440 gnd.n5436 9.3005
R12360 gnd.n5439 gnd.n5438 9.3005
R12361 gnd.n5437 gnd.n2787 9.3005
R12362 gnd.n5776 gnd.n2788 9.3005
R12363 gnd.n5775 gnd.n2789 9.3005
R12364 gnd.n5774 gnd.n2790 9.3005
R12365 gnd.n3030 gnd.n2791 9.3005
R12366 gnd.n3031 gnd.n3029 9.3005
R12367 gnd.n3033 gnd.n3032 9.3005
R12368 gnd.n3027 gnd.n3026 9.3005
R12369 gnd.n5483 gnd.n5482 9.3005
R12370 gnd.n5484 gnd.n3025 9.3005
R12371 gnd.n5488 gnd.n5485 9.3005
R12372 gnd.n5487 gnd.n5486 9.3005
R12373 gnd.n2999 gnd.n2998 9.3005
R12374 gnd.n5514 gnd.n5513 9.3005
R12375 gnd.n5515 gnd.n2997 9.3005
R12376 gnd.n5519 gnd.n5516 9.3005
R12377 gnd.n5518 gnd.n5517 9.3005
R12378 gnd.n2971 gnd.n2970 9.3005
R12379 gnd.n5545 gnd.n5544 9.3005
R12380 gnd.n5546 gnd.n2969 9.3005
R12381 gnd.n5557 gnd.n5547 9.3005
R12382 gnd.n5556 gnd.n5548 9.3005
R12383 gnd.n5555 gnd.n5549 9.3005
R12384 gnd.n5552 gnd.n5551 9.3005
R12385 gnd.n5550 gnd.n2917 9.3005
R12386 gnd.n5648 gnd.n2918 9.3005
R12387 gnd.n5647 gnd.n2919 9.3005
R12388 gnd.n5646 gnd.n2920 9.3005
R12389 gnd.n2922 gnd.n2921 9.3005
R12390 gnd.n7167 gnd.n305 9.3005
R12391 gnd.n326 gnd.n306 9.3005
R12392 gnd.n328 gnd.n327 9.3005
R12393 gnd.n329 gnd.n325 9.3005
R12394 gnd.n333 gnd.n332 9.3005
R12395 gnd.n334 gnd.n324 9.3005
R12396 gnd.n7149 gnd.n335 9.3005
R12397 gnd.n7148 gnd.n336 9.3005
R12398 gnd.n7147 gnd.n337 9.3005
R12399 gnd.n368 gnd.n338 9.3005
R12400 gnd.n370 gnd.n369 9.3005
R12401 gnd.n371 gnd.n367 9.3005
R12402 gnd.n375 gnd.n374 9.3005
R12403 gnd.n376 gnd.n366 9.3005
R12404 gnd.n7129 gnd.n377 9.3005
R12405 gnd.n7128 gnd.n378 9.3005
R12406 gnd.n7127 gnd.n379 9.3005
R12407 gnd.n7121 gnd.n380 9.3005
R12408 gnd.n4562 gnd.n3704 9.3005
R12409 gnd.n4565 gnd.n3703 9.3005
R12410 gnd.n4566 gnd.n3702 9.3005
R12411 gnd.n4569 gnd.n3701 9.3005
R12412 gnd.n4570 gnd.n3700 9.3005
R12413 gnd.n4573 gnd.n3699 9.3005
R12414 gnd.n4574 gnd.n3698 9.3005
R12415 gnd.n4577 gnd.n3697 9.3005
R12416 gnd.n4578 gnd.n3696 9.3005
R12417 gnd.n4581 gnd.n3695 9.3005
R12418 gnd.n4582 gnd.n3694 9.3005
R12419 gnd.n4585 gnd.n3693 9.3005
R12420 gnd.n4586 gnd.n3692 9.3005
R12421 gnd.n4587 gnd.n3691 9.3005
R12422 gnd.n3690 gnd.n3687 9.3005
R12423 gnd.n3689 gnd.n3688 9.3005
R12424 gnd.n4302 gnd.n4301 9.3005
R12425 gnd.n4298 gnd.n3709 9.3005
R12426 gnd.n4295 gnd.n3710 9.3005
R12427 gnd.n4294 gnd.n3711 9.3005
R12428 gnd.n4291 gnd.n3712 9.3005
R12429 gnd.n4290 gnd.n3713 9.3005
R12430 gnd.n4287 gnd.n3714 9.3005
R12431 gnd.n4286 gnd.n3715 9.3005
R12432 gnd.n4283 gnd.n3716 9.3005
R12433 gnd.n4282 gnd.n3717 9.3005
R12434 gnd.n4279 gnd.n3718 9.3005
R12435 gnd.n4278 gnd.n3719 9.3005
R12436 gnd.n4275 gnd.n3720 9.3005
R12437 gnd.n4274 gnd.n3721 9.3005
R12438 gnd.n4271 gnd.n3722 9.3005
R12439 gnd.n4270 gnd.n3723 9.3005
R12440 gnd.n4267 gnd.n3724 9.3005
R12441 gnd.n4266 gnd.n3725 9.3005
R12442 gnd.n4263 gnd.n4262 9.3005
R12443 gnd.n4261 gnd.n3727 9.3005
R12444 gnd.n4303 gnd.n3705 9.3005
R12445 gnd.n3809 gnd.n3808 9.3005
R12446 gnd.n4056 gnd.n4055 9.3005
R12447 gnd.n4057 gnd.n3807 9.3005
R12448 gnd.n4061 gnd.n4058 9.3005
R12449 gnd.n4062 gnd.n3806 9.3005
R12450 gnd.n4071 gnd.n4070 9.3005
R12451 gnd.n4072 gnd.n3805 9.3005
R12452 gnd.n4074 gnd.n4073 9.3005
R12453 gnd.n3800 gnd.n3799 9.3005
R12454 gnd.n4087 gnd.n4086 9.3005
R12455 gnd.n4088 gnd.n3798 9.3005
R12456 gnd.n4090 gnd.n4089 9.3005
R12457 gnd.n3794 gnd.n3793 9.3005
R12458 gnd.n4103 gnd.n4102 9.3005
R12459 gnd.n4104 gnd.n3792 9.3005
R12460 gnd.n4106 gnd.n4105 9.3005
R12461 gnd.n3787 gnd.n3786 9.3005
R12462 gnd.n4119 gnd.n4118 9.3005
R12463 gnd.n4120 gnd.n3785 9.3005
R12464 gnd.n4122 gnd.n4121 9.3005
R12465 gnd.n3781 gnd.n3780 9.3005
R12466 gnd.n4135 gnd.n4134 9.3005
R12467 gnd.n4136 gnd.n3779 9.3005
R12468 gnd.n4138 gnd.n4137 9.3005
R12469 gnd.n3774 gnd.n3773 9.3005
R12470 gnd.n4153 gnd.n4152 9.3005
R12471 gnd.n3998 gnd.n3997 9.3005
R12472 gnd.n4003 gnd.n4002 9.3005
R12473 gnd.n4006 gnd.n3992 9.3005
R12474 gnd.n4007 gnd.n3991 9.3005
R12475 gnd.n4010 gnd.n3990 9.3005
R12476 gnd.n4011 gnd.n3989 9.3005
R12477 gnd.n4014 gnd.n3988 9.3005
R12478 gnd.n4015 gnd.n3987 9.3005
R12479 gnd.n4018 gnd.n3986 9.3005
R12480 gnd.n4019 gnd.n3985 9.3005
R12481 gnd.n4022 gnd.n3984 9.3005
R12482 gnd.n4023 gnd.n3983 9.3005
R12483 gnd.n4026 gnd.n3982 9.3005
R12484 gnd.n4027 gnd.n3981 9.3005
R12485 gnd.n4030 gnd.n3980 9.3005
R12486 gnd.n4031 gnd.n3979 9.3005
R12487 gnd.n4034 gnd.n3978 9.3005
R12488 gnd.n4037 gnd.n4036 9.3005
R12489 gnd.n4001 gnd.n3996 9.3005
R12490 gnd.n4000 gnd.n3999 9.3005
R12491 gnd.n4044 gnd.n4043 9.3005
R12492 gnd.n4042 gnd.n3977 9.3005
R12493 gnd.n4041 gnd.n4040 9.3005
R12494 gnd.n4039 gnd.n2423 9.3005
R12495 gnd.n6053 gnd.n2424 9.3005
R12496 gnd.n6052 gnd.n2425 9.3005
R12497 gnd.n6051 gnd.n2426 9.3005
R12498 gnd.n2444 gnd.n2427 9.3005
R12499 gnd.n6041 gnd.n2445 9.3005
R12500 gnd.n6040 gnd.n2446 9.3005
R12501 gnd.n6039 gnd.n2447 9.3005
R12502 gnd.n2466 gnd.n2448 9.3005
R12503 gnd.n6029 gnd.n2467 9.3005
R12504 gnd.n6028 gnd.n2468 9.3005
R12505 gnd.n6027 gnd.n2469 9.3005
R12506 gnd.n2487 gnd.n2470 9.3005
R12507 gnd.n6017 gnd.n2488 9.3005
R12508 gnd.n6016 gnd.n2489 9.3005
R12509 gnd.n6015 gnd.n2490 9.3005
R12510 gnd.n2509 gnd.n2491 9.3005
R12511 gnd.n6005 gnd.n2510 9.3005
R12512 gnd.n6004 gnd.n2511 9.3005
R12513 gnd.n6003 gnd.n2512 9.3005
R12514 gnd.n2528 gnd.n2513 9.3005
R12515 gnd.n5993 gnd.n2529 9.3005
R12516 gnd.n5992 gnd.n2530 9.3005
R12517 gnd.n5991 gnd.n2531 9.3005
R12518 gnd.n2547 gnd.n2532 9.3005
R12519 gnd.n5980 gnd.n2548 9.3005
R12520 gnd.n5979 gnd.n2549 9.3005
R12521 gnd.n5978 gnd.n2550 9.3005
R12522 gnd.n2567 gnd.n2551 9.3005
R12523 gnd.n5968 gnd.n2568 9.3005
R12524 gnd.n5967 gnd.n2569 9.3005
R12525 gnd.n5966 gnd.n2570 9.3005
R12526 gnd.n2589 gnd.n2571 9.3005
R12527 gnd.n5956 gnd.n2590 9.3005
R12528 gnd.n5955 gnd.n2591 9.3005
R12529 gnd.n5954 gnd.n2592 9.3005
R12530 gnd.n2610 gnd.n2593 9.3005
R12531 gnd.n5944 gnd.n2611 9.3005
R12532 gnd.n5943 gnd.n2612 9.3005
R12533 gnd.n5942 gnd.n2613 9.3005
R12534 gnd.n2632 gnd.n2614 9.3005
R12535 gnd.n5932 gnd.n2633 9.3005
R12536 gnd.n5931 gnd.n2634 9.3005
R12537 gnd.n5930 gnd.n2635 9.3005
R12538 gnd.n2654 gnd.n2636 9.3005
R12539 gnd.n5920 gnd.n2655 9.3005
R12540 gnd.n5919 gnd.n2656 9.3005
R12541 gnd.n5918 gnd.n2657 9.3005
R12542 gnd.n2674 gnd.n2658 9.3005
R12543 gnd.n5908 gnd.n5907 9.3005
R12544 gnd.n4038 gnd.n3976 9.3005
R12545 gnd.n6067 gnd.n6066 9.3005
R12546 gnd.n6065 gnd.n2400 9.3005
R12547 gnd.n6064 gnd.n6063 9.3005
R12548 gnd.n2402 gnd.n2401 9.3005
R12549 gnd.n4064 gnd.n4063 9.3005
R12550 gnd.n4066 gnd.n4065 9.3005
R12551 gnd.n3804 gnd.n3803 9.3005
R12552 gnd.n4079 gnd.n4078 9.3005
R12553 gnd.n4080 gnd.n3802 9.3005
R12554 gnd.n4082 gnd.n4081 9.3005
R12555 gnd.n3797 gnd.n3796 9.3005
R12556 gnd.n4095 gnd.n4094 9.3005
R12557 gnd.n4096 gnd.n3795 9.3005
R12558 gnd.n4098 gnd.n4097 9.3005
R12559 gnd.n3791 gnd.n3790 9.3005
R12560 gnd.n4111 gnd.n4110 9.3005
R12561 gnd.n4112 gnd.n3789 9.3005
R12562 gnd.n4114 gnd.n4113 9.3005
R12563 gnd.n3784 gnd.n3783 9.3005
R12564 gnd.n4127 gnd.n4126 9.3005
R12565 gnd.n4128 gnd.n3782 9.3005
R12566 gnd.n4130 gnd.n4129 9.3005
R12567 gnd.n3778 gnd.n3777 9.3005
R12568 gnd.n4143 gnd.n4142 9.3005
R12569 gnd.n4144 gnd.n3776 9.3005
R12570 gnd.n4148 gnd.n4147 9.3005
R12571 gnd.n3771 gnd.n3770 9.3005
R12572 gnd.n4162 gnd.n4161 9.3005
R12573 gnd.n4163 gnd.n3769 9.3005
R12574 gnd.n4165 gnd.n4164 9.3005
R12575 gnd.n3765 gnd.n3764 9.3005
R12576 gnd.n4178 gnd.n4177 9.3005
R12577 gnd.n4179 gnd.n3763 9.3005
R12578 gnd.n4181 gnd.n4180 9.3005
R12579 gnd.n3758 gnd.n3757 9.3005
R12580 gnd.n4194 gnd.n4193 9.3005
R12581 gnd.n4195 gnd.n3756 9.3005
R12582 gnd.n4197 gnd.n4196 9.3005
R12583 gnd.n3752 gnd.n3751 9.3005
R12584 gnd.n4210 gnd.n4209 9.3005
R12585 gnd.n4211 gnd.n3750 9.3005
R12586 gnd.n4213 gnd.n4212 9.3005
R12587 gnd.n3745 gnd.n3744 9.3005
R12588 gnd.n4226 gnd.n4225 9.3005
R12589 gnd.n4227 gnd.n3743 9.3005
R12590 gnd.n4229 gnd.n4228 9.3005
R12591 gnd.n3739 gnd.n3738 9.3005
R12592 gnd.n4242 gnd.n4241 9.3005
R12593 gnd.n4243 gnd.n3737 9.3005
R12594 gnd.n4246 gnd.n4245 9.3005
R12595 gnd.n4244 gnd.n3731 9.3005
R12596 gnd.n4258 gnd.n3730 9.3005
R12597 gnd.n4260 gnd.n4259 9.3005
R12598 gnd.n6068 gnd.n2398 9.3005
R12599 gnd.n6075 gnd.n6074 9.3005
R12600 gnd.n6076 gnd.n2392 9.3005
R12601 gnd.n6079 gnd.n2391 9.3005
R12602 gnd.n6080 gnd.n2390 9.3005
R12603 gnd.n6083 gnd.n2389 9.3005
R12604 gnd.n6084 gnd.n2388 9.3005
R12605 gnd.n6087 gnd.n2387 9.3005
R12606 gnd.n6088 gnd.n2386 9.3005
R12607 gnd.n6091 gnd.n2385 9.3005
R12608 gnd.n6092 gnd.n2384 9.3005
R12609 gnd.n6095 gnd.n2383 9.3005
R12610 gnd.n6096 gnd.n2382 9.3005
R12611 gnd.n6099 gnd.n2381 9.3005
R12612 gnd.n6100 gnd.n2380 9.3005
R12613 gnd.n6103 gnd.n2379 9.3005
R12614 gnd.n6104 gnd.n2378 9.3005
R12615 gnd.n6107 gnd.n2377 9.3005
R12616 gnd.n6108 gnd.n2376 9.3005
R12617 gnd.n6111 gnd.n2375 9.3005
R12618 gnd.n6113 gnd.n2372 9.3005
R12619 gnd.n6116 gnd.n2371 9.3005
R12620 gnd.n6117 gnd.n2370 9.3005
R12621 gnd.n6120 gnd.n2369 9.3005
R12622 gnd.n6121 gnd.n2368 9.3005
R12623 gnd.n6124 gnd.n2367 9.3005
R12624 gnd.n6125 gnd.n2366 9.3005
R12625 gnd.n6128 gnd.n2365 9.3005
R12626 gnd.n6129 gnd.n2364 9.3005
R12627 gnd.n6132 gnd.n2363 9.3005
R12628 gnd.n6133 gnd.n2362 9.3005
R12629 gnd.n6136 gnd.n2361 9.3005
R12630 gnd.n6137 gnd.n2360 9.3005
R12631 gnd.n6140 gnd.n2359 9.3005
R12632 gnd.n6142 gnd.n2358 9.3005
R12633 gnd.n6143 gnd.n2357 9.3005
R12634 gnd.n6144 gnd.n2356 9.3005
R12635 gnd.n6145 gnd.n2355 9.3005
R12636 gnd.n6073 gnd.n2397 9.3005
R12637 gnd.n6072 gnd.n6071 9.3005
R12638 gnd.n4050 gnd.n4049 9.3005
R12639 gnd.n4048 gnd.n2411 9.3005
R12640 gnd.n6059 gnd.n2412 9.3005
R12641 gnd.n6058 gnd.n2413 9.3005
R12642 gnd.n6057 gnd.n2414 9.3005
R12643 gnd.n2434 gnd.n2415 9.3005
R12644 gnd.n6047 gnd.n2435 9.3005
R12645 gnd.n6046 gnd.n2436 9.3005
R12646 gnd.n6045 gnd.n2437 9.3005
R12647 gnd.n2455 gnd.n2438 9.3005
R12648 gnd.n6035 gnd.n2456 9.3005
R12649 gnd.n6034 gnd.n2457 9.3005
R12650 gnd.n6033 gnd.n2458 9.3005
R12651 gnd.n2477 gnd.n2459 9.3005
R12652 gnd.n6023 gnd.n2478 9.3005
R12653 gnd.n6022 gnd.n2479 9.3005
R12654 gnd.n6021 gnd.n2480 9.3005
R12655 gnd.n2498 gnd.n2481 9.3005
R12656 gnd.n6011 gnd.n2499 9.3005
R12657 gnd.n6010 gnd.n2500 9.3005
R12658 gnd.n6009 gnd.n2501 9.3005
R12659 gnd.n5973 gnd.n2559 9.3005
R12660 gnd.n5972 gnd.n2560 9.3005
R12661 gnd.n2578 gnd.n2561 9.3005
R12662 gnd.n5962 gnd.n2579 9.3005
R12663 gnd.n5961 gnd.n2580 9.3005
R12664 gnd.n5960 gnd.n2581 9.3005
R12665 gnd.n2600 gnd.n2582 9.3005
R12666 gnd.n5950 gnd.n2601 9.3005
R12667 gnd.n5949 gnd.n2602 9.3005
R12668 gnd.n5948 gnd.n2603 9.3005
R12669 gnd.n2621 gnd.n2604 9.3005
R12670 gnd.n5938 gnd.n2622 9.3005
R12671 gnd.n5937 gnd.n2623 9.3005
R12672 gnd.n5936 gnd.n2624 9.3005
R12673 gnd.n2643 gnd.n2625 9.3005
R12674 gnd.n5926 gnd.n2644 9.3005
R12675 gnd.n5925 gnd.n2645 9.3005
R12676 gnd.n5924 gnd.n2646 9.3005
R12677 gnd.n2664 gnd.n2647 9.3005
R12678 gnd.n5914 gnd.n2665 9.3005
R12679 gnd.n5913 gnd.n2666 9.3005
R12680 gnd.n5912 gnd.n2667 9.3005
R12681 gnd.n4047 gnd.n4046 9.3005
R12682 gnd.n5998 gnd.n2521 9.3005
R12683 gnd.n5974 gnd.n2521 9.3005
R12684 gnd.n3967 gnd.n3813 9.3005
R12685 gnd.n3816 gnd.n3814 9.3005
R12686 gnd.n3963 gnd.n3817 9.3005
R12687 gnd.n3962 gnd.n3818 9.3005
R12688 gnd.n3961 gnd.n3819 9.3005
R12689 gnd.n3822 gnd.n3820 9.3005
R12690 gnd.n3957 gnd.n3823 9.3005
R12691 gnd.n3956 gnd.n3824 9.3005
R12692 gnd.n3955 gnd.n3825 9.3005
R12693 gnd.n3828 gnd.n3826 9.3005
R12694 gnd.n3951 gnd.n3829 9.3005
R12695 gnd.n3950 gnd.n3830 9.3005
R12696 gnd.n3949 gnd.n3831 9.3005
R12697 gnd.n3834 gnd.n3832 9.3005
R12698 gnd.n3945 gnd.n3835 9.3005
R12699 gnd.n3944 gnd.n3836 9.3005
R12700 gnd.n3943 gnd.n3837 9.3005
R12701 gnd.n3969 gnd.n3968 9.3005
R12702 gnd.n3812 gnd.n964 9.3005
R12703 gnd.n6258 gnd.n963 9.3005
R12704 gnd.n6259 gnd.n962 9.3005
R12705 gnd.n6260 gnd.n961 9.3005
R12706 gnd.n960 gnd.n956 9.3005
R12707 gnd.n6266 gnd.n955 9.3005
R12708 gnd.n6267 gnd.n954 9.3005
R12709 gnd.n6268 gnd.n953 9.3005
R12710 gnd.n952 gnd.n948 9.3005
R12711 gnd.n6274 gnd.n947 9.3005
R12712 gnd.n6275 gnd.n946 9.3005
R12713 gnd.n6276 gnd.n945 9.3005
R12714 gnd.n944 gnd.n940 9.3005
R12715 gnd.n6282 gnd.n939 9.3005
R12716 gnd.n6283 gnd.n938 9.3005
R12717 gnd.n6284 gnd.n937 9.3005
R12718 gnd.n936 gnd.n932 9.3005
R12719 gnd.n6290 gnd.n931 9.3005
R12720 gnd.n6291 gnd.n930 9.3005
R12721 gnd.n6292 gnd.n929 9.3005
R12722 gnd.n928 gnd.n924 9.3005
R12723 gnd.n6298 gnd.n923 9.3005
R12724 gnd.n6299 gnd.n922 9.3005
R12725 gnd.n6300 gnd.n921 9.3005
R12726 gnd.n920 gnd.n916 9.3005
R12727 gnd.n6306 gnd.n915 9.3005
R12728 gnd.n6307 gnd.n914 9.3005
R12729 gnd.n6308 gnd.n913 9.3005
R12730 gnd.n912 gnd.n908 9.3005
R12731 gnd.n6314 gnd.n907 9.3005
R12732 gnd.n6315 gnd.n906 9.3005
R12733 gnd.n6316 gnd.n905 9.3005
R12734 gnd.n904 gnd.n900 9.3005
R12735 gnd.n6322 gnd.n899 9.3005
R12736 gnd.n6323 gnd.n898 9.3005
R12737 gnd.n6324 gnd.n897 9.3005
R12738 gnd.n896 gnd.n892 9.3005
R12739 gnd.n6330 gnd.n891 9.3005
R12740 gnd.n6331 gnd.n890 9.3005
R12741 gnd.n6332 gnd.n889 9.3005
R12742 gnd.n888 gnd.n884 9.3005
R12743 gnd.n6338 gnd.n883 9.3005
R12744 gnd.n6339 gnd.n882 9.3005
R12745 gnd.n6340 gnd.n881 9.3005
R12746 gnd.n880 gnd.n876 9.3005
R12747 gnd.n6346 gnd.n875 9.3005
R12748 gnd.n6347 gnd.n874 9.3005
R12749 gnd.n6348 gnd.n873 9.3005
R12750 gnd.n872 gnd.n868 9.3005
R12751 gnd.n6354 gnd.n867 9.3005
R12752 gnd.n6355 gnd.n866 9.3005
R12753 gnd.n6356 gnd.n865 9.3005
R12754 gnd.n864 gnd.n860 9.3005
R12755 gnd.n6362 gnd.n859 9.3005
R12756 gnd.n6363 gnd.n858 9.3005
R12757 gnd.n6364 gnd.n857 9.3005
R12758 gnd.n856 gnd.n852 9.3005
R12759 gnd.n6370 gnd.n851 9.3005
R12760 gnd.n6371 gnd.n850 9.3005
R12761 gnd.n6372 gnd.n849 9.3005
R12762 gnd.n848 gnd.n844 9.3005
R12763 gnd.n6378 gnd.n843 9.3005
R12764 gnd.n6379 gnd.n842 9.3005
R12765 gnd.n6380 gnd.n841 9.3005
R12766 gnd.n840 gnd.n836 9.3005
R12767 gnd.n6386 gnd.n835 9.3005
R12768 gnd.n6387 gnd.n834 9.3005
R12769 gnd.n6388 gnd.n833 9.3005
R12770 gnd.n832 gnd.n828 9.3005
R12771 gnd.n6394 gnd.n827 9.3005
R12772 gnd.n6395 gnd.n826 9.3005
R12773 gnd.n6396 gnd.n825 9.3005
R12774 gnd.n824 gnd.n820 9.3005
R12775 gnd.n6402 gnd.n819 9.3005
R12776 gnd.n6403 gnd.n818 9.3005
R12777 gnd.n6404 gnd.n817 9.3005
R12778 gnd.n816 gnd.n812 9.3005
R12779 gnd.n6410 gnd.n811 9.3005
R12780 gnd.n6411 gnd.n810 9.3005
R12781 gnd.n6412 gnd.n809 9.3005
R12782 gnd.n808 gnd.n804 9.3005
R12783 gnd.n6418 gnd.n803 9.3005
R12784 gnd.n6419 gnd.n802 9.3005
R12785 gnd.n6420 gnd.n801 9.3005
R12786 gnd.n3971 gnd.n3970 9.3005
R12787 gnd.n3135 gnd.n3134 9.3005
R12788 gnd.n3141 gnd.n3140 9.3005
R12789 gnd.n3142 gnd.n3117 9.3005
R12790 gnd.n3151 gnd.n3150 9.3005
R12791 gnd.n3119 gnd.n3115 9.3005
R12792 gnd.n3158 gnd.n3157 9.3005
R12793 gnd.n3159 gnd.n3108 9.3005
R12794 gnd.n3168 gnd.n3167 9.3005
R12795 gnd.n3110 gnd.n3106 9.3005
R12796 gnd.n3175 gnd.n3174 9.3005
R12797 gnd.n3176 gnd.n3099 9.3005
R12798 gnd.n3185 gnd.n3184 9.3005
R12799 gnd.n3101 gnd.n3097 9.3005
R12800 gnd.n3192 gnd.n3191 9.3005
R12801 gnd.n3193 gnd.n3087 9.3005
R12802 gnd.n3200 gnd.n3199 9.3005
R12803 gnd.n3089 gnd.n3085 9.3005
R12804 gnd.n3084 gnd.n3082 9.3005
R12805 gnd.n3125 gnd.n3124 9.3005
R12806 gnd.n3195 gnd.n3194 9.3005
R12807 gnd.n3096 gnd.n3093 9.3005
R12808 gnd.n3183 gnd.n3182 9.3005
R12809 gnd.n3179 gnd.n3100 9.3005
R12810 gnd.n3178 gnd.n3177 9.3005
R12811 gnd.n3105 gnd.n3102 9.3005
R12812 gnd.n3166 gnd.n3165 9.3005
R12813 gnd.n3162 gnd.n3109 9.3005
R12814 gnd.n3161 gnd.n3160 9.3005
R12815 gnd.n3114 gnd.n3111 9.3005
R12816 gnd.n3149 gnd.n3148 9.3005
R12817 gnd.n3145 gnd.n3118 9.3005
R12818 gnd.n3144 gnd.n3143 9.3005
R12819 gnd.n3123 gnd.n3120 9.3005
R12820 gnd.n3133 gnd.n3132 9.3005
R12821 gnd.n3129 gnd.n3128 9.3005
R12822 gnd.n3196 gnd.n3088 9.3005
R12823 gnd.n3198 gnd.n3197 9.3005
R12824 gnd.n5470 gnd.n5469 9.3005
R12825 gnd.n5468 gnd.n3083 9.3005
R12826 gnd.n5467 gnd.n5466 9.3005
R12827 gnd.n5465 gnd.n3210 9.3005
R12828 gnd.n5464 gnd.n5463 9.3005
R12829 gnd.n5462 gnd.n3211 9.3005
R12830 gnd.n5458 gnd.n5457 9.3005
R12831 gnd.n5456 gnd.n3218 9.3005
R12832 gnd.n5455 gnd.n5454 9.3005
R12833 gnd.n5453 gnd.n5448 9.3005
R12834 gnd.n4636 gnd.n4635 9.3005
R12835 gnd.n4637 gnd.n3517 9.3005
R12836 gnd.n4639 gnd.n4638 9.3005
R12837 gnd.n3505 gnd.n3504 9.3005
R12838 gnd.n4652 gnd.n4651 9.3005
R12839 gnd.n4653 gnd.n3503 9.3005
R12840 gnd.n4655 gnd.n4654 9.3005
R12841 gnd.n3492 gnd.n3491 9.3005
R12842 gnd.n4668 gnd.n4667 9.3005
R12843 gnd.n4669 gnd.n3490 9.3005
R12844 gnd.n4671 gnd.n4670 9.3005
R12845 gnd.n3479 gnd.n3478 9.3005
R12846 gnd.n4684 gnd.n4683 9.3005
R12847 gnd.n4685 gnd.n3477 9.3005
R12848 gnd.n4687 gnd.n4686 9.3005
R12849 gnd.n3465 gnd.n3464 9.3005
R12850 gnd.n4700 gnd.n4699 9.3005
R12851 gnd.n4701 gnd.n3463 9.3005
R12852 gnd.n4703 gnd.n4702 9.3005
R12853 gnd.n3451 gnd.n3450 9.3005
R12854 gnd.n4718 gnd.n4717 9.3005
R12855 gnd.n4719 gnd.n3448 9.3005
R12856 gnd.n4722 gnd.n4721 9.3005
R12857 gnd.n4720 gnd.n3449 9.3005
R12858 gnd.n3423 gnd.n3422 9.3005
R12859 gnd.n4849 gnd.n4848 9.3005
R12860 gnd.n4850 gnd.n3421 9.3005
R12861 gnd.n4852 gnd.n4851 9.3005
R12862 gnd.n3411 gnd.n3410 9.3005
R12863 gnd.n4865 gnd.n4864 9.3005
R12864 gnd.n4866 gnd.n3409 9.3005
R12865 gnd.n4868 gnd.n4867 9.3005
R12866 gnd.n3398 gnd.n3397 9.3005
R12867 gnd.n4881 gnd.n4880 9.3005
R12868 gnd.n4882 gnd.n3396 9.3005
R12869 gnd.n4884 gnd.n4883 9.3005
R12870 gnd.n3384 gnd.n3383 9.3005
R12871 gnd.n4899 gnd.n4898 9.3005
R12872 gnd.n4900 gnd.n3381 9.3005
R12873 gnd.n4903 gnd.n4902 9.3005
R12874 gnd.n4901 gnd.n3382 9.3005
R12875 gnd.n3356 gnd.n3355 9.3005
R12876 gnd.n5026 gnd.n5025 9.3005
R12877 gnd.n5027 gnd.n3354 9.3005
R12878 gnd.n5029 gnd.n5028 9.3005
R12879 gnd.n3342 gnd.n3341 9.3005
R12880 gnd.n5042 gnd.n5041 9.3005
R12881 gnd.n5043 gnd.n3340 9.3005
R12882 gnd.n5045 gnd.n5044 9.3005
R12883 gnd.n3327 gnd.n3326 9.3005
R12884 gnd.n5058 gnd.n5057 9.3005
R12885 gnd.n5059 gnd.n3325 9.3005
R12886 gnd.n5061 gnd.n5060 9.3005
R12887 gnd.n3312 gnd.n3311 9.3005
R12888 gnd.n5076 gnd.n5075 9.3005
R12889 gnd.n5077 gnd.n3309 9.3005
R12890 gnd.n5080 gnd.n5079 9.3005
R12891 gnd.n5078 gnd.n3310 9.3005
R12892 gnd.n3285 gnd.n3284 9.3005
R12893 gnd.n5360 gnd.n5359 9.3005
R12894 gnd.n5361 gnd.n3283 9.3005
R12895 gnd.n5363 gnd.n5362 9.3005
R12896 gnd.n3272 gnd.n3271 9.3005
R12897 gnd.n5376 gnd.n5375 9.3005
R12898 gnd.n5377 gnd.n3270 9.3005
R12899 gnd.n5379 gnd.n5378 9.3005
R12900 gnd.n3260 gnd.n3259 9.3005
R12901 gnd.n5392 gnd.n5391 9.3005
R12902 gnd.n5393 gnd.n3258 9.3005
R12903 gnd.n5395 gnd.n5394 9.3005
R12904 gnd.n3248 gnd.n3247 9.3005
R12905 gnd.n5408 gnd.n5407 9.3005
R12906 gnd.n5409 gnd.n3246 9.3005
R12907 gnd.n5411 gnd.n5410 9.3005
R12908 gnd.n3235 gnd.n3234 9.3005
R12909 gnd.n5424 gnd.n5423 9.3005
R12910 gnd.n5425 gnd.n3232 9.3005
R12911 gnd.n5429 gnd.n5428 9.3005
R12912 gnd.n5427 gnd.n3233 9.3005
R12913 gnd.n5426 gnd.n3220 9.3005
R12914 gnd.n5445 gnd.n3219 9.3005
R12915 gnd.n5447 gnd.n5446 9.3005
R12916 gnd.n3519 gnd.n3518 9.3005
R12917 gnd.n4620 gnd.n3543 9.3005
R12918 gnd.n4619 gnd.n4618 9.3005
R12919 gnd.n4615 gnd.n3544 9.3005
R12920 gnd.n4613 gnd.n4612 9.3005
R12921 gnd.n4611 gnd.n3547 9.3005
R12922 gnd.n4610 gnd.n4609 9.3005
R12923 gnd.n4606 gnd.n3550 9.3005
R12924 gnd.n4605 gnd.n4604 9.3005
R12925 gnd.n4603 gnd.n3551 9.3005
R12926 gnd.n4622 gnd.n4621 9.3005
R12927 gnd.n4155 gnd.n3772 9.3005
R12928 gnd.n4157 gnd.n4156 9.3005
R12929 gnd.n3768 gnd.n3767 9.3005
R12930 gnd.n4170 gnd.n4169 9.3005
R12931 gnd.n4171 gnd.n3766 9.3005
R12932 gnd.n4173 gnd.n4172 9.3005
R12933 gnd.n3761 gnd.n3760 9.3005
R12934 gnd.n4186 gnd.n4185 9.3005
R12935 gnd.n4187 gnd.n3759 9.3005
R12936 gnd.n4189 gnd.n4188 9.3005
R12937 gnd.n3755 gnd.n3754 9.3005
R12938 gnd.n4202 gnd.n4201 9.3005
R12939 gnd.n4203 gnd.n3753 9.3005
R12940 gnd.n4205 gnd.n4204 9.3005
R12941 gnd.n3748 gnd.n3747 9.3005
R12942 gnd.n4218 gnd.n4217 9.3005
R12943 gnd.n4219 gnd.n3746 9.3005
R12944 gnd.n4221 gnd.n4220 9.3005
R12945 gnd.n3742 gnd.n3741 9.3005
R12946 gnd.n4234 gnd.n4233 9.3005
R12947 gnd.n4235 gnd.n3740 9.3005
R12948 gnd.n4237 gnd.n4236 9.3005
R12949 gnd.n3736 gnd.n3735 9.3005
R12950 gnd.n4251 gnd.n4250 9.3005
R12951 gnd.n4252 gnd.n3733 9.3005
R12952 gnd.n4254 gnd.n4253 9.3005
R12953 gnd.n3734 gnd.n3554 9.3005
R12954 gnd.n4601 gnd.n4600 9.3005
R12955 gnd.n4597 gnd.n3555 9.3005
R12956 gnd.n4596 gnd.n4595 9.3005
R12957 gnd.n3661 gnd.n3556 9.3005
R12958 gnd.n3660 gnd.n3659 9.3005
R12959 gnd.n3656 gnd.n3655 9.3005
R12960 gnd.n3576 gnd.n3575 9.3005
R12961 gnd.n3649 gnd.n3648 9.3005
R12962 gnd.n3645 gnd.n3644 9.3005
R12963 gnd.n3584 gnd.n3581 9.3005
R12964 gnd.n3637 gnd.n3636 9.3005
R12965 gnd.n3633 gnd.n3632 9.3005
R12966 gnd.n3588 gnd.n3587 9.3005
R12967 gnd.n3625 gnd.n3624 9.3005
R12968 gnd.n3621 gnd.n3620 9.3005
R12969 gnd.n3596 gnd.n3593 9.3005
R12970 gnd.n3613 gnd.n3612 9.3005
R12971 gnd.n3609 gnd.n3608 9.3005
R12972 gnd.n3601 gnd.n3600 9.3005
R12973 gnd.n3603 gnd.n2676 9.3005
R12974 gnd.n3607 gnd.n3606 9.3005
R12975 gnd.n3598 gnd.n3597 9.3005
R12976 gnd.n3615 gnd.n3614 9.3005
R12977 gnd.n3619 gnd.n3618 9.3005
R12978 gnd.n3592 gnd.n3589 9.3005
R12979 gnd.n3627 gnd.n3626 9.3005
R12980 gnd.n3631 gnd.n3630 9.3005
R12981 gnd.n3586 gnd.n3585 9.3005
R12982 gnd.n3639 gnd.n3638 9.3005
R12983 gnd.n3643 gnd.n3642 9.3005
R12984 gnd.n3580 gnd.n3577 9.3005
R12985 gnd.n3651 gnd.n3650 9.3005
R12986 gnd.n3654 gnd.n3653 9.3005
R12987 gnd.n3574 gnd.n3573 9.3005
R12988 gnd.n3663 gnd.n3662 9.3005
R12989 gnd.n3562 gnd.n3559 9.3005
R12990 gnd.n4594 gnd.n4593 9.3005
R12991 gnd.n5902 gnd.n2677 9.3005
R12992 gnd.n5901 gnd.n5900 9.3005
R12993 gnd.n5899 gnd.n2681 9.3005
R12994 gnd.n5898 gnd.n5897 9.3005
R12995 gnd.n5896 gnd.n2682 9.3005
R12996 gnd.n5895 gnd.n5894 9.3005
R12997 gnd.n5893 gnd.n2686 9.3005
R12998 gnd.n5892 gnd.n5891 9.3005
R12999 gnd.n5890 gnd.n2687 9.3005
R13000 gnd.n5889 gnd.n5888 9.3005
R13001 gnd.n5887 gnd.n2691 9.3005
R13002 gnd.n5886 gnd.n5885 9.3005
R13003 gnd.n5884 gnd.n2692 9.3005
R13004 gnd.n5883 gnd.n5882 9.3005
R13005 gnd.n5881 gnd.n2696 9.3005
R13006 gnd.n5880 gnd.n5879 9.3005
R13007 gnd.n5878 gnd.n2697 9.3005
R13008 gnd.n5877 gnd.n5876 9.3005
R13009 gnd.n5875 gnd.n2701 9.3005
R13010 gnd.n5874 gnd.n5873 9.3005
R13011 gnd.n5872 gnd.n2702 9.3005
R13012 gnd.n5871 gnd.n5870 9.3005
R13013 gnd.n5869 gnd.n2706 9.3005
R13014 gnd.n5868 gnd.n5867 9.3005
R13015 gnd.n5866 gnd.n2707 9.3005
R13016 gnd.n5865 gnd.n5864 9.3005
R13017 gnd.n5863 gnd.n2711 9.3005
R13018 gnd.n5862 gnd.n5861 9.3005
R13019 gnd.n5860 gnd.n2712 9.3005
R13020 gnd.n5859 gnd.n5858 9.3005
R13021 gnd.n5857 gnd.n2716 9.3005
R13022 gnd.n5856 gnd.n5855 9.3005
R13023 gnd.n5854 gnd.n2717 9.3005
R13024 gnd.n5853 gnd.n5852 9.3005
R13025 gnd.n5851 gnd.n2721 9.3005
R13026 gnd.n5850 gnd.n5849 9.3005
R13027 gnd.n5848 gnd.n2722 9.3005
R13028 gnd.n5847 gnd.n5846 9.3005
R13029 gnd.n5845 gnd.n2726 9.3005
R13030 gnd.n5844 gnd.n5843 9.3005
R13031 gnd.n5842 gnd.n2727 9.3005
R13032 gnd.n5841 gnd.n5840 9.3005
R13033 gnd.n5839 gnd.n2731 9.3005
R13034 gnd.n5838 gnd.n5837 9.3005
R13035 gnd.n5836 gnd.n2732 9.3005
R13036 gnd.n5835 gnd.n5834 9.3005
R13037 gnd.n5833 gnd.n2736 9.3005
R13038 gnd.n5832 gnd.n5831 9.3005
R13039 gnd.n5830 gnd.n2737 9.3005
R13040 gnd.n5829 gnd.n5828 9.3005
R13041 gnd.n5827 gnd.n2741 9.3005
R13042 gnd.n5826 gnd.n5825 9.3005
R13043 gnd.n5824 gnd.n2742 9.3005
R13044 gnd.n5823 gnd.n5822 9.3005
R13045 gnd.n5821 gnd.n2746 9.3005
R13046 gnd.n5820 gnd.n5819 9.3005
R13047 gnd.n5818 gnd.n2747 9.3005
R13048 gnd.n5817 gnd.n5816 9.3005
R13049 gnd.n5815 gnd.n2751 9.3005
R13050 gnd.n5814 gnd.n5813 9.3005
R13051 gnd.n5812 gnd.n2752 9.3005
R13052 gnd.n5811 gnd.n5810 9.3005
R13053 gnd.n5809 gnd.n2756 9.3005
R13054 gnd.n5808 gnd.n5807 9.3005
R13055 gnd.n5806 gnd.n2757 9.3005
R13056 gnd.n5805 gnd.n5804 9.3005
R13057 gnd.n5803 gnd.n2761 9.3005
R13058 gnd.n5802 gnd.n5801 9.3005
R13059 gnd.n5800 gnd.n2762 9.3005
R13060 gnd.n5799 gnd.n5798 9.3005
R13061 gnd.n5797 gnd.n2766 9.3005
R13062 gnd.n5796 gnd.n5795 9.3005
R13063 gnd.n5794 gnd.n2767 9.3005
R13064 gnd.n5793 gnd.n5792 9.3005
R13065 gnd.n5791 gnd.n2771 9.3005
R13066 gnd.n5790 gnd.n5789 9.3005
R13067 gnd.n5788 gnd.n2772 9.3005
R13068 gnd.n5787 gnd.n5786 9.3005
R13069 gnd.n5785 gnd.n2776 9.3005
R13070 gnd.n5784 gnd.n5783 9.3005
R13071 gnd.n5782 gnd.n2777 9.3005
R13072 gnd.n5781 gnd.n2780 9.3005
R13073 gnd.n5904 gnd.n5903 9.3005
R13074 gnd.n5690 gnd.n2877 9.3005
R13075 gnd.n5689 gnd.n5688 9.3005
R13076 gnd.n5687 gnd.n2879 9.3005
R13077 gnd.n5686 gnd.n5685 9.3005
R13078 gnd.n5684 gnd.n2883 9.3005
R13079 gnd.n5683 gnd.n5682 9.3005
R13080 gnd.n5681 gnd.n2884 9.3005
R13081 gnd.n5680 gnd.n5679 9.3005
R13082 gnd.n5678 gnd.n2888 9.3005
R13083 gnd.n5677 gnd.n5676 9.3005
R13084 gnd.n5675 gnd.n2889 9.3005
R13085 gnd.n5674 gnd.n5673 9.3005
R13086 gnd.n5672 gnd.n2893 9.3005
R13087 gnd.n5671 gnd.n5670 9.3005
R13088 gnd.n5669 gnd.n2894 9.3005
R13089 gnd.n5668 gnd.n5667 9.3005
R13090 gnd.n5666 gnd.n2898 9.3005
R13091 gnd.n5665 gnd.n5664 9.3005
R13092 gnd.n5663 gnd.n2899 9.3005
R13093 gnd.n5662 gnd.n5661 9.3005
R13094 gnd.n281 gnd.n279 9.3005
R13095 gnd.n7198 gnd.n7197 9.3005
R13096 gnd.n7196 gnd.n280 9.3005
R13097 gnd.n7195 gnd.n7194 9.3005
R13098 gnd.n7193 gnd.n282 9.3005
R13099 gnd.n7192 gnd.n7191 9.3005
R13100 gnd.n7189 gnd.n286 9.3005
R13101 gnd.n7188 gnd.n7187 9.3005
R13102 gnd.n7186 gnd.n288 9.3005
R13103 gnd.n257 gnd.n256 9.3005
R13104 gnd.n7210 gnd.n7209 9.3005
R13105 gnd.n7211 gnd.n255 9.3005
R13106 gnd.n7213 gnd.n7212 9.3005
R13107 gnd.n242 gnd.n241 9.3005
R13108 gnd.n7226 gnd.n7225 9.3005
R13109 gnd.n7227 gnd.n240 9.3005
R13110 gnd.n7229 gnd.n7228 9.3005
R13111 gnd.n227 gnd.n226 9.3005
R13112 gnd.n7242 gnd.n7241 9.3005
R13113 gnd.n7243 gnd.n225 9.3005
R13114 gnd.n7245 gnd.n7244 9.3005
R13115 gnd.n212 gnd.n211 9.3005
R13116 gnd.n7258 gnd.n7257 9.3005
R13117 gnd.n7259 gnd.n210 9.3005
R13118 gnd.n7261 gnd.n7260 9.3005
R13119 gnd.n197 gnd.n196 9.3005
R13120 gnd.n7274 gnd.n7273 9.3005
R13121 gnd.n7275 gnd.n194 9.3005
R13122 gnd.n7352 gnd.n7351 9.3005
R13123 gnd.n7350 gnd.n195 9.3005
R13124 gnd.n7349 gnd.n7348 9.3005
R13125 gnd.n7347 gnd.n7276 9.3005
R13126 gnd.n7346 gnd.n7345 9.3005
R13127 gnd.n5692 gnd.n5691 9.3005
R13128 gnd.n7342 gnd.n7278 9.3005
R13129 gnd.n7341 gnd.n7340 9.3005
R13130 gnd.n7339 gnd.n7283 9.3005
R13131 gnd.n7338 gnd.n7337 9.3005
R13132 gnd.n7336 gnd.n7284 9.3005
R13133 gnd.n7335 gnd.n7334 9.3005
R13134 gnd.n7333 gnd.n7291 9.3005
R13135 gnd.n7332 gnd.n7331 9.3005
R13136 gnd.n7330 gnd.n7292 9.3005
R13137 gnd.n7329 gnd.n7328 9.3005
R13138 gnd.n7327 gnd.n7299 9.3005
R13139 gnd.n7326 gnd.n7325 9.3005
R13140 gnd.n7324 gnd.n7300 9.3005
R13141 gnd.n7323 gnd.n7322 9.3005
R13142 gnd.n7321 gnd.n7307 9.3005
R13143 gnd.n7320 gnd.n7319 9.3005
R13144 gnd.n7318 gnd.n7308 9.3005
R13145 gnd.n7317 gnd.n7316 9.3005
R13146 gnd.n7344 gnd.n7343 9.3005
R13147 gnd.n5474 gnd.n3080 9.3005
R13148 gnd.n5477 gnd.n5476 9.3005
R13149 gnd.n5475 gnd.n3081 9.3005
R13150 gnd.n3007 gnd.n3006 9.3005
R13151 gnd.n5504 gnd.n5503 9.3005
R13152 gnd.n5505 gnd.n3004 9.3005
R13153 gnd.n5508 gnd.n5507 9.3005
R13154 gnd.n5506 gnd.n3005 9.3005
R13155 gnd.n2979 gnd.n2978 9.3005
R13156 gnd.n5535 gnd.n5534 9.3005
R13157 gnd.n5536 gnd.n2976 9.3005
R13158 gnd.n5539 gnd.n5538 9.3005
R13159 gnd.n5537 gnd.n2977 9.3005
R13160 gnd.n2951 gnd.n2950 9.3005
R13161 gnd.n5574 gnd.n5573 9.3005
R13162 gnd.n5575 gnd.n2948 9.3005
R13163 gnd.n5581 gnd.n5580 9.3005
R13164 gnd.n5579 gnd.n2949 9.3005
R13165 gnd.n5578 gnd.n5577 9.3005
R13166 gnd.n2940 gnd.n2939 9.3005
R13167 gnd.n5600 gnd.n5599 9.3005
R13168 gnd.n5601 gnd.n2937 9.3005
R13169 gnd.n5606 gnd.n5605 9.3005
R13170 gnd.n5604 gnd.n2938 9.3005
R13171 gnd.n5603 gnd.n5602 9.3005
R13172 gnd.n65 gnd.n63 9.3005
R13173 gnd.n7483 gnd.n7482 9.3005
R13174 gnd.n7481 gnd.n64 9.3005
R13175 gnd.n7480 gnd.n7479 9.3005
R13176 gnd.n7478 gnd.n69 9.3005
R13177 gnd.n7477 gnd.n7476 9.3005
R13178 gnd.n7475 gnd.n70 9.3005
R13179 gnd.n7474 gnd.n7473 9.3005
R13180 gnd.n7472 gnd.n74 9.3005
R13181 gnd.n7471 gnd.n7470 9.3005
R13182 gnd.n7469 gnd.n75 9.3005
R13183 gnd.n7468 gnd.n7467 9.3005
R13184 gnd.n7466 gnd.n79 9.3005
R13185 gnd.n7465 gnd.n7464 9.3005
R13186 gnd.n7463 gnd.n80 9.3005
R13187 gnd.n7462 gnd.n7461 9.3005
R13188 gnd.n7460 gnd.n84 9.3005
R13189 gnd.n7459 gnd.n7458 9.3005
R13190 gnd.n7457 gnd.n85 9.3005
R13191 gnd.n7456 gnd.n7455 9.3005
R13192 gnd.n7454 gnd.n89 9.3005
R13193 gnd.n7453 gnd.n7452 9.3005
R13194 gnd.n7451 gnd.n90 9.3005
R13195 gnd.n7450 gnd.n7449 9.3005
R13196 gnd.n7448 gnd.n94 9.3005
R13197 gnd.n7447 gnd.n7446 9.3005
R13198 gnd.n7445 gnd.n95 9.3005
R13199 gnd.n7444 gnd.n98 9.3005
R13200 gnd.n5473 gnd.n5472 9.3005
R13201 gnd.t48 gnd.n1192 9.24152
R13202 gnd.n6218 gnd.t150 9.24152
R13203 gnd.n2312 gnd.t136 9.24152
R13204 gnd.n5916 gnd.t97 9.24152
R13205 gnd.t86 gnd.n5479 9.24152
R13206 gnd.t22 gnd.t48 8.92286
R13207 gnd.n4715 gnd.n3453 8.92286
R13208 gnd.n4826 gnd.n4825 8.92286
R13209 gnd.t6 gnd.n3407 8.92286
R13210 gnd.n4896 gnd.n3387 8.92286
R13211 gnd.n5003 gnd.n5002 8.92286
R13212 gnd.n4980 gnd.t27 8.92286
R13213 gnd.n5073 gnd.n3316 8.92286
R13214 gnd.n5337 gnd.n5336 8.92286
R13215 gnd.n2292 gnd.n2267 8.92171
R13216 gnd.n2260 gnd.n2235 8.92171
R13217 gnd.n2228 gnd.n2203 8.92171
R13218 gnd.n2197 gnd.n2172 8.92171
R13219 gnd.n2165 gnd.n2140 8.92171
R13220 gnd.n2133 gnd.n2108 8.92171
R13221 gnd.n2101 gnd.n2076 8.92171
R13222 gnd.n2070 gnd.n2045 8.92171
R13223 gnd.n5132 gnd.n5114 8.72777
R13224 gnd.n1836 gnd.t51 8.60421
R13225 gnd.t11 gnd.t160 8.60421
R13226 gnd.n4779 gnd.t18 8.60421
R13227 gnd.t71 gnd.n3359 8.60421
R13228 gnd.n1264 gnd.n1248 8.43467
R13229 gnd.n46 gnd.n30 8.43467
R13230 gnd.n4154 gnd.n0 8.41456
R13231 gnd.n7485 gnd.n7484 8.41456
R13232 gnd.n6254 gnd.n966 8.28555
R13233 gnd.n2293 gnd.n2265 8.14595
R13234 gnd.n2261 gnd.n2233 8.14595
R13235 gnd.n2229 gnd.n2201 8.14595
R13236 gnd.n2198 gnd.n2170 8.14595
R13237 gnd.n2166 gnd.n2138 8.14595
R13238 gnd.n2134 gnd.n2106 8.14595
R13239 gnd.n2102 gnd.n2074 8.14595
R13240 gnd.n2071 gnd.n2043 8.14595
R13241 gnd.n2298 gnd.n2297 7.97301
R13242 gnd.t52 gnd.n1351 7.9669
R13243 gnd.n4484 gnd.t11 7.9669
R13244 gnd.t41 gnd.t143 7.9669
R13245 gnd.n7318 gnd.n7317 7.75808
R13246 gnd.n3197 gnd.n3196 7.75808
R13247 gnd.n4593 gnd.n3562 7.75808
R13248 gnd.n3999 gnd.n3996 7.75808
R13249 gnd.n4705 gnd.n3461 7.64824
R13250 gnd.n4818 gnd.n4739 7.64824
R13251 gnd.n4886 gnd.t13 7.64824
R13252 gnd.n4886 gnd.n3394 7.64824
R13253 gnd.n4995 gnd.n4919 7.64824
R13254 gnd.n4919 gnd.t30 7.64824
R13255 gnd.n5063 gnd.n3323 7.64824
R13256 gnd.n1745 gnd.t57 7.32958
R13257 gnd.n4348 gnd.n4347 7.30353
R13258 gnd.n5131 gnd.n5130 7.30353
R13259 gnd.n1705 gnd.n1424 7.01093
R13260 gnd.n1427 gnd.n1425 7.01093
R13261 gnd.n1715 gnd.n1714 7.01093
R13262 gnd.n1726 gnd.n1408 7.01093
R13263 gnd.n1725 gnd.n1411 7.01093
R13264 gnd.n1736 gnd.n1399 7.01093
R13265 gnd.n1402 gnd.n1400 7.01093
R13266 gnd.n1746 gnd.n1745 7.01093
R13267 gnd.n1756 gnd.n1380 7.01093
R13268 gnd.n1755 gnd.n1383 7.01093
R13269 gnd.n1764 gnd.n1374 7.01093
R13270 gnd.n1776 gnd.n1364 7.01093
R13271 gnd.n1786 gnd.n1349 7.01093
R13272 gnd.n1802 gnd.n1801 7.01093
R13273 gnd.n1351 gnd.n1288 7.01093
R13274 gnd.n1856 gnd.n1289 7.01093
R13275 gnd.n1850 gnd.n1849 7.01093
R13276 gnd.n1338 gnd.n1300 7.01093
R13277 gnd.n1842 gnd.n1311 7.01093
R13278 gnd.n1329 gnd.n1324 7.01093
R13279 gnd.n1836 gnd.n1835 7.01093
R13280 gnd.n1882 gnd.n1227 7.01093
R13281 gnd.n1881 gnd.n1880 7.01093
R13282 gnd.n1893 gnd.n1892 7.01093
R13283 gnd.n1220 gnd.n1212 7.01093
R13284 gnd.n1922 gnd.n1200 7.01093
R13285 gnd.n1921 gnd.n1203 7.01093
R13286 gnd.n1932 gnd.n1192 7.01093
R13287 gnd.n1193 gnd.n1181 7.01093
R13288 gnd.n1945 gnd.n1182 7.01093
R13289 gnd.n1996 gnd.n1174 7.01093
R13290 gnd.n1995 gnd.n1165 7.01093
R13291 gnd.n6253 gnd.n968 7.01093
R13292 gnd.n1986 gnd.n977 7.01093
R13293 gnd.n6247 gnd.n6246 7.01093
R13294 gnd.n1154 gnd.n980 7.01093
R13295 gnd.n6240 gnd.n989 7.01093
R13296 gnd.n6239 gnd.n992 7.01093
R13297 gnd.n6233 gnd.n6232 7.01093
R13298 gnd.n1151 gnd.n1004 7.01093
R13299 gnd.n6226 gnd.n1015 7.01093
R13300 gnd.n6225 gnd.n1018 7.01093
R13301 gnd.n1968 gnd.n1027 7.01093
R13302 gnd.n6219 gnd.n6218 7.01093
R13303 gnd.n2313 gnd.n2312 7.01093
R13304 gnd.n6212 gnd.n1040 7.01093
R13305 gnd.n6211 gnd.n1043 7.01093
R13306 gnd.t111 gnd.n3973 7.01093
R13307 gnd.n4467 gnd.t2 7.01093
R13308 gnd.t26 gnd.n5335 7.01093
R13309 gnd.n182 gnd.t79 7.01093
R13310 gnd.n1383 gnd.t44 6.69227
R13311 gnd.n1203 gnd.t22 6.69227
R13312 gnd.t50 gnd.n1001 6.69227
R13313 gnd.n6043 gnd.t254 6.69227
R13314 gnd.t195 gnd.n2453 6.69227
R13315 gnd.n4223 gnd.t204 6.69227
R13316 gnd.t187 gnd.n2638 6.69227
R13317 gnd.n4468 gnd.t24 6.69227
R13318 gnd.n5365 gnd.t64 6.69227
R13319 gnd.n5511 gnd.t257 6.69227
R13320 gnd.n2994 gnd.t212 6.69227
R13321 gnd.n7144 gnd.t230 6.69227
R13322 gnd.n7136 gnd.t216 6.69227
R13323 gnd.n5244 gnd.n5243 6.5566
R13324 gnd.n4553 gnd.n4552 6.5566
R13325 gnd.n4372 gnd.n4366 6.5566
R13326 gnd.n5256 gnd.n5161 6.5566
R13327 gnd.n4491 gnd.n4327 6.37362
R13328 gnd.n4697 gnd.n3467 6.37362
R13329 gnd.n4846 gnd.t14 6.37362
R13330 gnd.n4811 gnd.n4810 6.37362
R13331 gnd.n4793 gnd.t13 6.37362
R13332 gnd.t30 gnd.n3344 6.37362
R13333 gnd.n5055 gnd.n3331 6.37362
R13334 gnd.n4957 gnd.t31 6.37362
R13335 gnd.n5322 gnd.n5321 6.37362
R13336 gnd.n5389 gnd.n3262 6.37362
R13337 gnd.n4615 gnd.n4614 6.20656
R13338 gnd.n7407 gnd.n7404 6.20656
R13339 gnd.n6112 gnd.n6111 6.20656
R13340 gnd.n5461 gnd.n5458 6.20656
R13341 gnd.t317 gnd.n1812 6.05496
R13342 gnd.n1813 gnd.t59 6.05496
R13343 gnd.t69 gnd.n1227 6.05496
R13344 gnd.t54 gnd.n2010 6.05496
R13345 gnd.n6019 gnd.t225 6.05496
R13346 gnd.t197 gnd.n2496 6.05496
R13347 gnd.n4191 gnd.t214 6.05496
R13348 gnd.t183 gnd.n2595 6.05496
R13349 gnd.n2967 gnd.t193 6.05496
R13350 gnd.n5584 gnd.t243 6.05496
R13351 gnd.n7164 gnd.t270 6.05496
R13352 gnd.n7156 gnd.t279 6.05496
R13353 gnd.n2295 gnd.n2265 5.81868
R13354 gnd.n2263 gnd.n2233 5.81868
R13355 gnd.n2231 gnd.n2201 5.81868
R13356 gnd.n2200 gnd.n2170 5.81868
R13357 gnd.n2168 gnd.n2138 5.81868
R13358 gnd.n2136 gnd.n2106 5.81868
R13359 gnd.n2104 gnd.n2074 5.81868
R13360 gnd.n2073 gnd.n2043 5.81868
R13361 gnd.n4715 gnd.t2 5.73631
R13362 gnd.t33 gnd.n3386 5.73631
R13363 gnd.n5001 gnd.t68 5.73631
R13364 gnd.n5336 gnd.t26 5.73631
R13365 gnd.n5389 gnd.t76 5.73631
R13366 gnd.n5163 gnd.n2841 5.62001
R13367 gnd.n4560 gnd.n4305 5.62001
R13368 gnd.n4560 gnd.n4306 5.62001
R13369 gnd.n5254 gnd.n2841 5.62001
R13370 gnd.n1564 gnd.n1559 5.4308
R13371 gnd.n1144 gnd.n1074 5.4308
R13372 gnd.n1880 gnd.t53 5.41765
R13373 gnd.t56 gnd.n1903 5.41765
R13374 gnd.t36 gnd.n966 5.41765
R13375 gnd.n5995 gnd.t189 5.41765
R13376 gnd.t228 gnd.n2537 5.41765
R13377 gnd.n4159 gnd.t228 5.41765
R13378 gnd.t199 gnd.n2553 5.41765
R13379 gnd.t4 gnd.n3439 5.41765
R13380 gnd.t321 gnd.n5082 5.41765
R13381 gnd.t185 gnd.n276 5.41765
R13382 gnd.n5636 gnd.t259 5.41765
R13383 gnd.n2932 gnd.t259 5.41765
R13384 gnd.n7179 gnd.t267 5.41765
R13385 gnd.n4689 gnd.n3475 5.09899
R13386 gnd.t160 gnd.n3475 5.09899
R13387 gnd.n4484 gnd.n4483 5.09899
R13388 gnd.n4725 gnd.t8 5.09899
R13389 gnd.n4870 gnd.n3407 5.09899
R13390 gnd.n4802 gnd.n4751 5.09899
R13391 gnd.n5047 gnd.n3338 5.09899
R13392 gnd.n4980 gnd.n4930 5.09899
R13393 gnd.n5343 gnd.t182 5.09899
R13394 gnd.t123 gnd.n5096 5.09899
R13395 gnd.n5381 gnd.t143 5.09899
R13396 gnd.n5314 gnd.n5108 5.09899
R13397 gnd.n2293 gnd.n2292 5.04292
R13398 gnd.n2261 gnd.n2260 5.04292
R13399 gnd.n2229 gnd.n2228 5.04292
R13400 gnd.n2198 gnd.n2197 5.04292
R13401 gnd.n2166 gnd.n2165 5.04292
R13402 gnd.n2134 gnd.n2133 5.04292
R13403 gnd.n2102 gnd.n2101 5.04292
R13404 gnd.n2071 gnd.n2070 5.04292
R13405 gnd.n1280 gnd.n1279 4.82753
R13406 gnd.n62 gnd.n61 4.82753
R13407 gnd.n1843 gnd.t58 4.78034
R13408 gnd.n1182 gnd.t47 4.78034
R13409 gnd.n4124 gnd.t197 4.78034
R13410 gnd.t209 gnd.n2515 4.78034
R13411 gnd.n5970 gnd.t191 4.78034
R13412 gnd.t214 gnd.n2576 4.78034
R13413 gnd.n3440 gnd.t4 4.78034
R13414 gnd.n5083 gnd.t321 4.78034
R13415 gnd.n5136 gnd.t154 4.78034
R13416 gnd.t243 gnd.n2910 4.78034
R13417 gnd.n5659 gnd.t218 4.78034
R13418 gnd.n7172 gnd.t206 4.78034
R13419 gnd.n7215 gnd.t270 4.78034
R13420 gnd.n1285 gnd.n1282 4.74817
R13421 gnd.n1335 gnd.n1233 4.74817
R13422 gnd.n1322 gnd.n1232 4.74817
R13423 gnd.n1231 gnd.n1230 4.74817
R13424 gnd.n1331 gnd.n1282 4.74817
R13425 gnd.n1332 gnd.n1233 4.74817
R13426 gnd.n1334 gnd.n1232 4.74817
R13427 gnd.n1321 gnd.n1231 4.74817
R13428 gnd.n7203 gnd.n7202 4.74817
R13429 gnd.n2931 gnd.n267 4.74817
R13430 gnd.n7181 gnd.n266 4.74817
R13431 gnd.n265 gnd.n262 4.74817
R13432 gnd.n7203 gnd.n269 4.74817
R13433 gnd.n5634 gnd.n267 4.74817
R13434 gnd.n2930 gnd.n266 4.74817
R13435 gnd.n7182 gnd.n265 4.74817
R13436 gnd.n3840 gnd.n3838 4.74817
R13437 gnd.n3937 gnd.n3841 4.74817
R13438 gnd.n3935 gnd.n3845 4.74817
R13439 gnd.n3928 gnd.n3844 4.74817
R13440 gnd.n3924 gnd.n3843 4.74817
R13441 gnd.n5641 gnd.n5640 4.74817
R13442 gnd.n5623 gnd.n2924 4.74817
R13443 gnd.n5628 gnd.n5627 4.74817
R13444 gnd.n5624 gnd.n304 4.74817
R13445 gnd.n7169 gnd.n7168 4.74817
R13446 gnd.n5642 gnd.n5641 4.74817
R13447 gnd.n5639 gnd.n2924 4.74817
R13448 gnd.n5629 gnd.n5628 4.74817
R13449 gnd.n5626 gnd.n5624 4.74817
R13450 gnd.n7170 gnd.n7169 4.74817
R13451 gnd.n2520 gnd.n2502 4.74817
R13452 gnd.n2539 gnd.n2522 4.74817
R13453 gnd.n5986 gnd.n5985 4.74817
R13454 gnd.n2558 gnd.n2540 4.74817
R13455 gnd.n5999 gnd.n2520 4.74817
R13456 gnd.n5997 gnd.n2522 4.74817
R13457 gnd.n5987 gnd.n5986 4.74817
R13458 gnd.n5984 gnd.n2540 4.74817
R13459 gnd.n3939 gnd.n3840 4.74817
R13460 gnd.n3938 gnd.n3937 4.74817
R13461 gnd.n3935 gnd.n3934 4.74817
R13462 gnd.n3930 gnd.n3844 4.74817
R13463 gnd.n3927 gnd.n3843 4.74817
R13464 gnd.n1264 gnd.n1263 4.7074
R13465 gnd.n46 gnd.n45 4.7074
R13466 gnd.n1280 gnd.n1264 4.65959
R13467 gnd.n62 gnd.n46 4.65959
R13468 gnd.n5738 gnd.n2843 4.6132
R13469 gnd.n4561 gnd.n4304 4.6132
R13470 gnd.n4590 gnd.n3564 4.46168
R13471 gnd.n4491 gnd.t83 4.46168
R13472 gnd.n4838 gnd.t20 4.46168
R13473 gnd.n5349 gnd.t32 4.46168
R13474 gnd.n5770 gnd.n2821 4.46168
R13475 gnd.n5127 gnd.n5114 4.46111
R13476 gnd.n2278 gnd.n2274 4.38594
R13477 gnd.n2246 gnd.n2242 4.38594
R13478 gnd.n2214 gnd.n2210 4.38594
R13479 gnd.n2183 gnd.n2179 4.38594
R13480 gnd.n2151 gnd.n2147 4.38594
R13481 gnd.n2119 gnd.n2115 4.38594
R13482 gnd.n2087 gnd.n2083 4.38594
R13483 gnd.n2056 gnd.n2052 4.38594
R13484 gnd.n2289 gnd.n2267 4.26717
R13485 gnd.n2257 gnd.n2235 4.26717
R13486 gnd.n2225 gnd.n2203 4.26717
R13487 gnd.n2194 gnd.n2172 4.26717
R13488 gnd.n2162 gnd.n2140 4.26717
R13489 gnd.n2130 gnd.n2108 4.26717
R13490 gnd.n2098 gnd.n2076 4.26717
R13491 gnd.n2067 gnd.n2045 4.26717
R13492 gnd.n1787 gnd.t49 4.14303
R13493 gnd.n1154 gnd.t45 4.14303
R13494 gnd.n4092 gnd.t195 4.14303
R13495 gnd.t222 gnd.n2472 4.14303
R13496 gnd.n5946 gnd.t202 4.14303
R13497 gnd.t204 gnd.n2619 4.14303
R13498 gnd.t212 gnd.n2981 4.14303
R13499 gnd.t274 gnd.n5541 4.14303
R13500 gnd.n7151 gnd.t234 4.14303
R13501 gnd.n7247 gnd.t230 4.14303
R13502 gnd.n2297 gnd.n2296 4.08274
R13503 gnd.n5243 gnd.n5242 4.05904
R13504 gnd.n4552 gnd.n4551 4.05904
R13505 gnd.n4376 gnd.n4366 4.05904
R13506 gnd.n5161 gnd.n5156 4.05904
R13507 gnd.n15 gnd.n7 3.99943
R13508 gnd.n4476 gnd.n4442 3.82437
R13509 gnd.t15 gnd.n4739 3.82437
R13510 gnd.n4862 gnd.n3413 3.82437
R13511 gnd.n4795 gnd.n4794 3.82437
R13512 gnd.n5039 gnd.n3346 3.82437
R13513 gnd.n4973 gnd.n4972 3.82437
R13514 gnd.n5063 gnd.t7 3.82437
R13515 gnd.n5373 gnd.n3275 3.82437
R13516 gnd.n2297 gnd.n2169 3.70378
R13517 gnd.n1860 gnd.n1281 3.65935
R13518 gnd.n15 gnd.n14 3.60163
R13519 gnd.t236 gnd.n2429 3.50571
R13520 gnd.n7131 gnd.t264 3.50571
R13521 gnd.n2288 gnd.n2269 3.49141
R13522 gnd.n2256 gnd.n2237 3.49141
R13523 gnd.n2224 gnd.n2205 3.49141
R13524 gnd.n2193 gnd.n2174 3.49141
R13525 gnd.n2161 gnd.n2142 3.49141
R13526 gnd.n2129 gnd.n2110 3.49141
R13527 gnd.n2097 gnd.n2078 3.49141
R13528 gnd.n2066 gnd.n2047 3.49141
R13529 gnd.n4796 gnd.t3 3.18706
R13530 gnd.n4988 gnd.t10 3.18706
R13531 gnd.n1366 gnd.t49 2.8684
R13532 gnd.t24 gnd.t163 2.8684
R13533 gnd.n1265 gnd.t295 2.82907
R13534 gnd.n1265 gnd.t248 2.82907
R13535 gnd.n1267 gnd.t281 2.82907
R13536 gnd.n1267 gnd.t184 2.82907
R13537 gnd.n1269 gnd.t208 2.82907
R13538 gnd.n1269 gnd.t192 2.82907
R13539 gnd.n1271 gnd.t190 2.82907
R13540 gnd.n1271 gnd.t304 2.82907
R13541 gnd.n1273 gnd.t198 2.82907
R13542 gnd.n1273 gnd.t240 2.82907
R13543 gnd.n1275 gnd.t273 2.82907
R13544 gnd.n1275 gnd.t226 2.82907
R13545 gnd.n1277 gnd.t255 2.82907
R13546 gnd.n1277 gnd.t196 2.82907
R13547 gnd.n1234 gnd.t203 2.82907
R13548 gnd.n1234 gnd.t224 2.82907
R13549 gnd.n1236 gnd.t239 2.82907
R13550 gnd.n1236 gnd.t296 2.82907
R13551 gnd.n1238 gnd.t220 2.82907
R13552 gnd.n1238 gnd.t211 2.82907
R13553 gnd.n1240 gnd.t261 2.82907
R13554 gnd.n1240 gnd.t250 2.82907
R13555 gnd.n1242 gnd.t301 2.82907
R13556 gnd.n1242 gnd.t232 2.82907
R13557 gnd.n1244 gnd.t246 2.82907
R13558 gnd.n1244 gnd.t272 2.82907
R13559 gnd.n1246 gnd.t284 2.82907
R13560 gnd.n1246 gnd.t221 2.82907
R13561 gnd.n1249 gnd.t303 2.82907
R13562 gnd.n1249 gnd.t205 2.82907
R13563 gnd.n1251 gnd.t215 2.82907
R13564 gnd.n1251 gnd.t276 2.82907
R13565 gnd.n1253 gnd.t200 2.82907
R13566 gnd.n1253 gnd.t310 2.82907
R13567 gnd.n1255 gnd.t238 2.82907
R13568 gnd.n1255 gnd.t229 2.82907
R13569 gnd.n1257 gnd.t285 2.82907
R13570 gnd.n1257 gnd.t210 2.82907
R13571 gnd.n1259 gnd.t223 2.82907
R13572 gnd.n1259 gnd.t247 2.82907
R13573 gnd.n1261 gnd.t262 2.82907
R13574 gnd.n1261 gnd.t201 2.82907
R13575 gnd.n59 gnd.t293 2.82907
R13576 gnd.n59 gnd.t217 2.82907
R13577 gnd.n57 gnd.t309 2.82907
R13578 gnd.n57 gnd.t235 2.82907
R13579 gnd.n55 gnd.t207 2.82907
R13580 gnd.n55 gnd.t302 2.82907
R13581 gnd.n53 gnd.t277 2.82907
R13582 gnd.n53 gnd.t288 2.82907
R13583 gnd.n51 gnd.t291 2.82907
R13584 gnd.n51 gnd.t307 2.82907
R13585 gnd.n49 gnd.t286 2.82907
R13586 gnd.n49 gnd.t244 2.82907
R13587 gnd.n47 gnd.t213 2.82907
R13588 gnd.n47 gnd.t275 2.82907
R13589 gnd.n28 gnd.t251 2.82907
R13590 gnd.n28 gnd.t305 2.82907
R13591 gnd.n26 gnd.t298 2.82907
R13592 gnd.n26 gnd.t278 2.82907
R13593 gnd.n24 gnd.t263 2.82907
R13594 gnd.n24 gnd.t294 2.82907
R13595 gnd.n22 gnd.t283 2.82907
R13596 gnd.n22 gnd.t290 2.82907
R13597 gnd.n20 gnd.t242 2.82907
R13598 gnd.n20 gnd.t186 2.82907
R13599 gnd.n18 gnd.t194 2.82907
R13600 gnd.n18 gnd.t269 2.82907
R13601 gnd.n16 gnd.t253 2.82907
R13602 gnd.n16 gnd.t308 2.82907
R13603 gnd.n43 gnd.t231 2.82907
R13604 gnd.n43 gnd.t292 2.82907
R13605 gnd.n41 gnd.t280 2.82907
R13606 gnd.n41 gnd.t252 2.82907
R13607 gnd.n39 gnd.t241 2.82907
R13608 gnd.n39 gnd.t271 2.82907
R13609 gnd.n37 gnd.t260 2.82907
R13610 gnd.n37 gnd.t268 2.82907
R13611 gnd.n35 gnd.t219 2.82907
R13612 gnd.n35 gnd.t306 2.82907
R13613 gnd.n33 gnd.t300 2.82907
R13614 gnd.n33 gnd.t245 2.82907
R13615 gnd.n31 gnd.t233 2.82907
R13616 gnd.n31 gnd.t297 2.82907
R13617 gnd.n2285 gnd.n2284 2.71565
R13618 gnd.n2253 gnd.n2252 2.71565
R13619 gnd.n2221 gnd.n2220 2.71565
R13620 gnd.n2190 gnd.n2189 2.71565
R13621 gnd.n2158 gnd.n2157 2.71565
R13622 gnd.n2126 gnd.n2125 2.71565
R13623 gnd.n2094 gnd.n2093 2.71565
R13624 gnd.n2063 gnd.n2062 2.71565
R13625 gnd.n4444 gnd.t130 2.54975
R13626 gnd.n4469 gnd.n4468 2.54975
R13627 gnd.n4854 gnd.n3419 2.54975
R13628 gnd.n4787 gnd.n4786 2.54975
R13629 gnd.n4778 gnd.t21 2.54975
R13630 gnd.n5023 gnd.t0 2.54975
R13631 gnd.n5031 gnd.n3352 2.54975
R13632 gnd.n4965 gnd.n4945 2.54975
R13633 gnd.n5365 gnd.n3281 2.54975
R13634 gnd.n5329 gnd.t123 2.54975
R13635 gnd.n1860 gnd.n1282 2.27742
R13636 gnd.n1860 gnd.n1233 2.27742
R13637 gnd.n1860 gnd.n1232 2.27742
R13638 gnd.n1860 gnd.n1231 2.27742
R13639 gnd.n7204 gnd.n7203 2.27742
R13640 gnd.n7204 gnd.n267 2.27742
R13641 gnd.n7204 gnd.n266 2.27742
R13642 gnd.n7204 gnd.n265 2.27742
R13643 gnd.n5641 gnd.n264 2.27742
R13644 gnd.n2924 gnd.n264 2.27742
R13645 gnd.n5628 gnd.n264 2.27742
R13646 gnd.n5624 gnd.n264 2.27742
R13647 gnd.n7169 gnd.n264 2.27742
R13648 gnd.n2521 gnd.n2520 2.27742
R13649 gnd.n2522 gnd.n2521 2.27742
R13650 gnd.n5986 gnd.n2521 2.27742
R13651 gnd.n2540 gnd.n2521 2.27742
R13652 gnd.n3936 gnd.n3840 2.27742
R13653 gnd.n3937 gnd.n3936 2.27742
R13654 gnd.n3936 gnd.n3935 2.27742
R13655 gnd.n3936 gnd.n3844 2.27742
R13656 gnd.n3936 gnd.n3843 2.27742
R13657 gnd.n1714 gnd.t93 2.23109
R13658 gnd.n1337 gnd.t58 2.23109
R13659 gnd.n3973 gnd.n2405 2.23109
R13660 gnd.n4878 gnd.t62 2.23109
R13661 gnd.t66 gnd.n4987 2.23109
R13662 gnd.n7362 gnd.n182 2.23109
R13663 gnd.n2281 gnd.n2271 1.93989
R13664 gnd.n2249 gnd.n2239 1.93989
R13665 gnd.n2217 gnd.n2207 1.93989
R13666 gnd.n2186 gnd.n2176 1.93989
R13667 gnd.n2154 gnd.n2144 1.93989
R13668 gnd.n2122 gnd.n2112 1.93989
R13669 gnd.n2090 gnd.n2080 1.93989
R13670 gnd.n2059 gnd.n2049 1.93989
R13671 gnd.n4824 gnd.t38 1.91244
R13672 gnd.t43 gnd.n3314 1.91244
R13673 gnd.t28 gnd.n1725 1.59378
R13674 gnd.n1904 gnd.t56 1.59378
R13675 gnd.n1167 gnd.t36 1.59378
R13676 gnd.n4461 gnd.n4460 1.27512
R13677 gnd.n4846 gnd.n3425 1.27512
R13678 gnd.n4779 gnd.n4778 1.27512
R13679 gnd.n5023 gnd.n3359 1.27512
R13680 gnd.n4958 gnd.n4957 1.27512
R13681 gnd.n5357 gnd.n3287 1.27512
R13682 gnd.n1567 gnd.n1559 1.16414
R13683 gnd.n1141 gnd.n1074 1.16414
R13684 gnd.n2280 gnd.n2273 1.16414
R13685 gnd.n2248 gnd.n2241 1.16414
R13686 gnd.n2216 gnd.n2209 1.16414
R13687 gnd.n2185 gnd.n2178 1.16414
R13688 gnd.n2153 gnd.n2146 1.16414
R13689 gnd.n2121 gnd.n2114 1.16414
R13690 gnd.n2089 gnd.n2082 1.16414
R13691 gnd.n2058 gnd.n2051 1.16414
R13692 gnd.n5738 gnd.n5737 0.970197
R13693 gnd.n4561 gnd.n3705 0.970197
R13694 gnd.n2264 gnd.n2232 0.962709
R13695 gnd.n2296 gnd.n2264 0.962709
R13696 gnd.n2137 gnd.n2105 0.962709
R13697 gnd.n2169 gnd.n2137 0.962709
R13698 gnd.n1813 gnd.t317 0.956468
R13699 gnd.n2011 gnd.t54 0.956468
R13700 gnd.n4673 gnd.t311 0.956468
R13701 gnd.t3 gnd.t62 0.956468
R13702 gnd.t10 gnd.t66 0.956468
R13703 gnd.n3256 gnd.t16 0.956468
R13704 gnd.n1274 gnd.n1272 0.773756
R13705 gnd.n56 gnd.n54 0.773756
R13706 gnd.n1279 gnd.n1278 0.773756
R13707 gnd.n1278 gnd.n1276 0.773756
R13708 gnd.n1276 gnd.n1274 0.773756
R13709 gnd.n1272 gnd.n1270 0.773756
R13710 gnd.n1270 gnd.n1268 0.773756
R13711 gnd.n1268 gnd.n1266 0.773756
R13712 gnd.n50 gnd.n48 0.773756
R13713 gnd.n52 gnd.n50 0.773756
R13714 gnd.n54 gnd.n52 0.773756
R13715 gnd.n58 gnd.n56 0.773756
R13716 gnd.n60 gnd.n58 0.773756
R13717 gnd.n61 gnd.n60 0.773756
R13718 gnd.n2 gnd.n1 0.672012
R13719 gnd.n3 gnd.n2 0.672012
R13720 gnd.n4 gnd.n3 0.672012
R13721 gnd.n5 gnd.n4 0.672012
R13722 gnd.n6 gnd.n5 0.672012
R13723 gnd.n7 gnd.n6 0.672012
R13724 gnd.n9 gnd.n8 0.672012
R13725 gnd.n10 gnd.n9 0.672012
R13726 gnd.n11 gnd.n10 0.672012
R13727 gnd.n12 gnd.n11 0.672012
R13728 gnd.n13 gnd.n12 0.672012
R13729 gnd.n14 gnd.n13 0.672012
R13730 gnd.n4697 gnd.t126 0.637812
R13731 gnd.n4811 gnd.t1 0.637812
R13732 gnd.t9 gnd.n3331 0.637812
R13733 gnd.n5321 gnd.t119 0.637812
R13734 gnd gnd.n0 0.59317
R13735 gnd.n1248 gnd.n1247 0.573776
R13736 gnd.n1247 gnd.n1245 0.573776
R13737 gnd.n1245 gnd.n1243 0.573776
R13738 gnd.n1243 gnd.n1241 0.573776
R13739 gnd.n1241 gnd.n1239 0.573776
R13740 gnd.n1239 gnd.n1237 0.573776
R13741 gnd.n1237 gnd.n1235 0.573776
R13742 gnd.n1263 gnd.n1262 0.573776
R13743 gnd.n1262 gnd.n1260 0.573776
R13744 gnd.n1260 gnd.n1258 0.573776
R13745 gnd.n1258 gnd.n1256 0.573776
R13746 gnd.n1256 gnd.n1254 0.573776
R13747 gnd.n1254 gnd.n1252 0.573776
R13748 gnd.n1252 gnd.n1250 0.573776
R13749 gnd.n19 gnd.n17 0.573776
R13750 gnd.n21 gnd.n19 0.573776
R13751 gnd.n23 gnd.n21 0.573776
R13752 gnd.n25 gnd.n23 0.573776
R13753 gnd.n27 gnd.n25 0.573776
R13754 gnd.n29 gnd.n27 0.573776
R13755 gnd.n30 gnd.n29 0.573776
R13756 gnd.n34 gnd.n32 0.573776
R13757 gnd.n36 gnd.n34 0.573776
R13758 gnd.n38 gnd.n36 0.573776
R13759 gnd.n40 gnd.n38 0.573776
R13760 gnd.n42 gnd.n40 0.573776
R13761 gnd.n44 gnd.n42 0.573776
R13762 gnd.n45 gnd.n44 0.573776
R13763 gnd.n7486 gnd.n7485 0.553533
R13764 gnd.n7204 gnd.n264 0.548625
R13765 gnd.n3936 gnd.n2521 0.548625
R13766 gnd.n5905 gnd.n5904 0.523366
R13767 gnd.n3127 gnd.n2780 0.523366
R13768 gnd.n4000 gnd.n3998 0.505073
R13769 gnd.n4038 gnd.n4037 0.505073
R13770 gnd.n7345 gnd.n7344 0.505073
R13771 gnd.n7316 gnd.n98 0.505073
R13772 gnd.n7439 gnd.n7438 0.492878
R13773 gnd.n7368 gnd.n7367 0.492878
R13774 gnd.n5698 gnd.n2869 0.492878
R13775 gnd.n3037 gnd.n2825 0.492878
R13776 gnd.n3689 gnd.n2667 0.492878
R13777 gnd.n4261 gnd.n4260 0.492878
R13778 gnd.n6072 gnd.n2398 0.492878
R13779 gnd.n4047 gnd.n2355 0.492878
R13780 gnd.n5448 gnd.n5447 0.489829
R13781 gnd.n4621 gnd.n3518 0.489829
R13782 gnd.n2319 gnd.n2318 0.486781
R13783 gnd.n1616 gnd.n1615 0.48678
R13784 gnd.n6157 gnd.n6156 0.480683
R13785 gnd.n1700 gnd.n1699 0.480683
R13786 gnd.n801 gnd.n796 0.447146
R13787 gnd.n6910 gnd.n6909 0.447146
R13788 gnd.n7122 gnd.n7121 0.447146
R13789 gnd.n3970 gnd.n3969 0.447146
R13790 gnd.n5907 gnd.n5906 0.404992
R13791 gnd.n5691 gnd.n2878 0.404992
R13792 gnd.n4614 gnd.n4613 0.388379
R13793 gnd.n2277 gnd.n2276 0.388379
R13794 gnd.n2245 gnd.n2244 0.388379
R13795 gnd.n2213 gnd.n2212 0.388379
R13796 gnd.n2182 gnd.n2181 0.388379
R13797 gnd.n2150 gnd.n2149 0.388379
R13798 gnd.n2118 gnd.n2117 0.388379
R13799 gnd.n2086 gnd.n2085 0.388379
R13800 gnd.n2055 gnd.n2054 0.388379
R13801 gnd.n7408 gnd.n7407 0.388379
R13802 gnd.n6113 gnd.n6112 0.388379
R13803 gnd.n5462 gnd.n5461 0.388379
R13804 gnd.n7486 gnd.n15 0.374463
R13805 gnd.n1977 gnd.t50 0.319156
R13806 gnd.n4741 gnd.t34 0.319156
R13807 gnd.t60 gnd.n4971 0.319156
R13808 gnd.n1534 gnd.n1512 0.311721
R13809 gnd gnd.n7486 0.295112
R13810 gnd.n4602 gnd.n3554 0.27489
R13811 gnd.n5473 gnd.n5471 0.27489
R13812 gnd.n6202 gnd.n1048 0.268793
R13813 gnd.n1088 gnd.n1048 0.241354
R13814 gnd.n2843 gnd.n2840 0.229039
R13815 gnd.n2846 gnd.n2843 0.229039
R13816 gnd.n4304 gnd.n3704 0.229039
R13817 gnd.n4304 gnd.n4303 0.229039
R13818 gnd.n1688 gnd.n1487 0.206293
R13819 gnd.n1281 gnd.n0 0.169152
R13820 gnd.n2294 gnd.n2266 0.155672
R13821 gnd.n2287 gnd.n2266 0.155672
R13822 gnd.n2287 gnd.n2286 0.155672
R13823 gnd.n2286 gnd.n2270 0.155672
R13824 gnd.n2279 gnd.n2270 0.155672
R13825 gnd.n2279 gnd.n2278 0.155672
R13826 gnd.n2262 gnd.n2234 0.155672
R13827 gnd.n2255 gnd.n2234 0.155672
R13828 gnd.n2255 gnd.n2254 0.155672
R13829 gnd.n2254 gnd.n2238 0.155672
R13830 gnd.n2247 gnd.n2238 0.155672
R13831 gnd.n2247 gnd.n2246 0.155672
R13832 gnd.n2230 gnd.n2202 0.155672
R13833 gnd.n2223 gnd.n2202 0.155672
R13834 gnd.n2223 gnd.n2222 0.155672
R13835 gnd.n2222 gnd.n2206 0.155672
R13836 gnd.n2215 gnd.n2206 0.155672
R13837 gnd.n2215 gnd.n2214 0.155672
R13838 gnd.n2199 gnd.n2171 0.155672
R13839 gnd.n2192 gnd.n2171 0.155672
R13840 gnd.n2192 gnd.n2191 0.155672
R13841 gnd.n2191 gnd.n2175 0.155672
R13842 gnd.n2184 gnd.n2175 0.155672
R13843 gnd.n2184 gnd.n2183 0.155672
R13844 gnd.n2167 gnd.n2139 0.155672
R13845 gnd.n2160 gnd.n2139 0.155672
R13846 gnd.n2160 gnd.n2159 0.155672
R13847 gnd.n2159 gnd.n2143 0.155672
R13848 gnd.n2152 gnd.n2143 0.155672
R13849 gnd.n2152 gnd.n2151 0.155672
R13850 gnd.n2135 gnd.n2107 0.155672
R13851 gnd.n2128 gnd.n2107 0.155672
R13852 gnd.n2128 gnd.n2127 0.155672
R13853 gnd.n2127 gnd.n2111 0.155672
R13854 gnd.n2120 gnd.n2111 0.155672
R13855 gnd.n2120 gnd.n2119 0.155672
R13856 gnd.n2103 gnd.n2075 0.155672
R13857 gnd.n2096 gnd.n2075 0.155672
R13858 gnd.n2096 gnd.n2095 0.155672
R13859 gnd.n2095 gnd.n2079 0.155672
R13860 gnd.n2088 gnd.n2079 0.155672
R13861 gnd.n2088 gnd.n2087 0.155672
R13862 gnd.n2072 gnd.n2044 0.155672
R13863 gnd.n2065 gnd.n2044 0.155672
R13864 gnd.n2065 gnd.n2064 0.155672
R13865 gnd.n2064 gnd.n2048 0.155672
R13866 gnd.n2057 gnd.n2048 0.155672
R13867 gnd.n2057 gnd.n2056 0.155672
R13868 gnd.n6191 gnd.n6157 0.152939
R13869 gnd.n6191 gnd.n6190 0.152939
R13870 gnd.n6190 gnd.n6189 0.152939
R13871 gnd.n6189 gnd.n6159 0.152939
R13872 gnd.n6160 gnd.n6159 0.152939
R13873 gnd.n6161 gnd.n6160 0.152939
R13874 gnd.n6162 gnd.n6161 0.152939
R13875 gnd.n6163 gnd.n6162 0.152939
R13876 gnd.n6164 gnd.n6163 0.152939
R13877 gnd.n6165 gnd.n6164 0.152939
R13878 gnd.n6166 gnd.n6165 0.152939
R13879 gnd.n6167 gnd.n6166 0.152939
R13880 gnd.n6167 gnd.n1054 0.152939
R13881 gnd.n6200 gnd.n1054 0.152939
R13882 gnd.n6201 gnd.n6200 0.152939
R13883 gnd.n6202 gnd.n6201 0.152939
R13884 gnd.n1701 gnd.n1700 0.152939
R13885 gnd.n1701 gnd.n1405 0.152939
R13886 gnd.n1729 gnd.n1405 0.152939
R13887 gnd.n1730 gnd.n1729 0.152939
R13888 gnd.n1731 gnd.n1730 0.152939
R13889 gnd.n1732 gnd.n1731 0.152939
R13890 gnd.n1732 gnd.n1377 0.152939
R13891 gnd.n1759 gnd.n1377 0.152939
R13892 gnd.n1760 gnd.n1759 0.152939
R13893 gnd.n1761 gnd.n1760 0.152939
R13894 gnd.n1761 gnd.n1355 0.152939
R13895 gnd.n1790 gnd.n1355 0.152939
R13896 gnd.n1791 gnd.n1790 0.152939
R13897 gnd.n1792 gnd.n1791 0.152939
R13898 gnd.n1793 gnd.n1792 0.152939
R13899 gnd.n1795 gnd.n1793 0.152939
R13900 gnd.n1795 gnd.n1794 0.152939
R13901 gnd.n1794 gnd.n1304 0.152939
R13902 gnd.n1305 gnd.n1304 0.152939
R13903 gnd.n1306 gnd.n1305 0.152939
R13904 gnd.n1325 gnd.n1306 0.152939
R13905 gnd.n1326 gnd.n1325 0.152939
R13906 gnd.n1326 gnd.n1224 0.152939
R13907 gnd.n1885 gnd.n1224 0.152939
R13908 gnd.n1886 gnd.n1885 0.152939
R13909 gnd.n1887 gnd.n1886 0.152939
R13910 gnd.n1888 gnd.n1887 0.152939
R13911 gnd.n1888 gnd.n1197 0.152939
R13912 gnd.n1925 gnd.n1197 0.152939
R13913 gnd.n1926 gnd.n1925 0.152939
R13914 gnd.n1927 gnd.n1926 0.152939
R13915 gnd.n1928 gnd.n1927 0.152939
R13916 gnd.n1928 gnd.n1171 0.152939
R13917 gnd.n1999 gnd.n1171 0.152939
R13918 gnd.n2000 gnd.n1999 0.152939
R13919 gnd.n2001 gnd.n2000 0.152939
R13920 gnd.n2002 gnd.n2001 0.152939
R13921 gnd.n2004 gnd.n2002 0.152939
R13922 gnd.n2004 gnd.n2003 0.152939
R13923 gnd.n2003 gnd.n984 0.152939
R13924 gnd.n985 gnd.n984 0.152939
R13925 gnd.n986 gnd.n985 0.152939
R13926 gnd.n1008 gnd.n986 0.152939
R13927 gnd.n1009 gnd.n1008 0.152939
R13928 gnd.n1010 gnd.n1009 0.152939
R13929 gnd.n1011 gnd.n1010 0.152939
R13930 gnd.n1012 gnd.n1011 0.152939
R13931 gnd.n1033 gnd.n1012 0.152939
R13932 gnd.n1034 gnd.n1033 0.152939
R13933 gnd.n1035 gnd.n1034 0.152939
R13934 gnd.n1036 gnd.n1035 0.152939
R13935 gnd.n1037 gnd.n1036 0.152939
R13936 gnd.n6156 gnd.n1037 0.152939
R13937 gnd.n1699 gnd.n1429 0.152939
R13938 gnd.n1450 gnd.n1429 0.152939
R13939 gnd.n1451 gnd.n1450 0.152939
R13940 gnd.n1457 gnd.n1451 0.152939
R13941 gnd.n1458 gnd.n1457 0.152939
R13942 gnd.n1459 gnd.n1458 0.152939
R13943 gnd.n1459 gnd.n1448 0.152939
R13944 gnd.n1467 gnd.n1448 0.152939
R13945 gnd.n1468 gnd.n1467 0.152939
R13946 gnd.n1469 gnd.n1468 0.152939
R13947 gnd.n1469 gnd.n1446 0.152939
R13948 gnd.n1477 gnd.n1446 0.152939
R13949 gnd.n1478 gnd.n1477 0.152939
R13950 gnd.n1479 gnd.n1478 0.152939
R13951 gnd.n1479 gnd.n1444 0.152939
R13952 gnd.n1487 gnd.n1444 0.152939
R13953 gnd.n1089 gnd.n1088 0.152939
R13954 gnd.n1090 gnd.n1089 0.152939
R13955 gnd.n1090 gnd.n1084 0.152939
R13956 gnd.n1098 gnd.n1084 0.152939
R13957 gnd.n1099 gnd.n1098 0.152939
R13958 gnd.n1100 gnd.n1099 0.152939
R13959 gnd.n1100 gnd.n1082 0.152939
R13960 gnd.n1108 gnd.n1082 0.152939
R13961 gnd.n1109 gnd.n1108 0.152939
R13962 gnd.n1110 gnd.n1109 0.152939
R13963 gnd.n1110 gnd.n1080 0.152939
R13964 gnd.n1118 gnd.n1080 0.152939
R13965 gnd.n1119 gnd.n1118 0.152939
R13966 gnd.n1120 gnd.n1119 0.152939
R13967 gnd.n1120 gnd.n1078 0.152939
R13968 gnd.n1128 gnd.n1078 0.152939
R13969 gnd.n1129 gnd.n1128 0.152939
R13970 gnd.n1130 gnd.n1129 0.152939
R13971 gnd.n1130 gnd.n1076 0.152939
R13972 gnd.n1138 gnd.n1076 0.152939
R13973 gnd.n1139 gnd.n1138 0.152939
R13974 gnd.n1140 gnd.n1139 0.152939
R13975 gnd.n1140 gnd.n1071 0.152939
R13976 gnd.n1147 gnd.n1071 0.152939
R13977 gnd.n1148 gnd.n1147 0.152939
R13978 gnd.n2319 gnd.n1148 0.152939
R13979 gnd.n1862 gnd.n1861 0.152939
R13980 gnd.n1863 gnd.n1862 0.152939
R13981 gnd.n1864 gnd.n1863 0.152939
R13982 gnd.n1865 gnd.n1864 0.152939
R13983 gnd.n1866 gnd.n1865 0.152939
R13984 gnd.n1867 gnd.n1866 0.152939
R13985 gnd.n1867 gnd.n1178 0.152939
R13986 gnd.n1948 gnd.n1178 0.152939
R13987 gnd.n1949 gnd.n1948 0.152939
R13988 gnd.n1950 gnd.n1949 0.152939
R13989 gnd.n1951 gnd.n1950 0.152939
R13990 gnd.n1952 gnd.n1951 0.152939
R13991 gnd.n1953 gnd.n1952 0.152939
R13992 gnd.n1954 gnd.n1953 0.152939
R13993 gnd.n1955 gnd.n1954 0.152939
R13994 gnd.n1956 gnd.n1955 0.152939
R13995 gnd.n1957 gnd.n1956 0.152939
R13996 gnd.n1958 gnd.n1957 0.152939
R13997 gnd.n1959 gnd.n1958 0.152939
R13998 gnd.n1960 gnd.n1959 0.152939
R13999 gnd.n1961 gnd.n1960 0.152939
R14000 gnd.n1962 gnd.n1961 0.152939
R14001 gnd.n1963 gnd.n1962 0.152939
R14002 gnd.n1964 gnd.n1963 0.152939
R14003 gnd.n1966 gnd.n1964 0.152939
R14004 gnd.n1966 gnd.n1965 0.152939
R14005 gnd.n1965 gnd.n1149 0.152939
R14006 gnd.n2318 gnd.n1149 0.152939
R14007 gnd.n1617 gnd.n1616 0.152939
R14008 gnd.n1617 gnd.n1507 0.152939
R14009 gnd.n1632 gnd.n1507 0.152939
R14010 gnd.n1633 gnd.n1632 0.152939
R14011 gnd.n1634 gnd.n1633 0.152939
R14012 gnd.n1634 gnd.n1495 0.152939
R14013 gnd.n1648 gnd.n1495 0.152939
R14014 gnd.n1649 gnd.n1648 0.152939
R14015 gnd.n1650 gnd.n1649 0.152939
R14016 gnd.n1651 gnd.n1650 0.152939
R14017 gnd.n1652 gnd.n1651 0.152939
R14018 gnd.n1653 gnd.n1652 0.152939
R14019 gnd.n1654 gnd.n1653 0.152939
R14020 gnd.n1655 gnd.n1654 0.152939
R14021 gnd.n1656 gnd.n1655 0.152939
R14022 gnd.n1657 gnd.n1656 0.152939
R14023 gnd.n1658 gnd.n1657 0.152939
R14024 gnd.n1659 gnd.n1658 0.152939
R14025 gnd.n1660 gnd.n1659 0.152939
R14026 gnd.n1661 gnd.n1660 0.152939
R14027 gnd.n1662 gnd.n1661 0.152939
R14028 gnd.n1662 gnd.n1361 0.152939
R14029 gnd.n1779 gnd.n1361 0.152939
R14030 gnd.n1780 gnd.n1779 0.152939
R14031 gnd.n1781 gnd.n1780 0.152939
R14032 gnd.n1782 gnd.n1781 0.152939
R14033 gnd.n1782 gnd.n1283 0.152939
R14034 gnd.n1859 gnd.n1283 0.152939
R14035 gnd.n1535 gnd.n1534 0.152939
R14036 gnd.n1536 gnd.n1535 0.152939
R14037 gnd.n1537 gnd.n1536 0.152939
R14038 gnd.n1538 gnd.n1537 0.152939
R14039 gnd.n1539 gnd.n1538 0.152939
R14040 gnd.n1540 gnd.n1539 0.152939
R14041 gnd.n1541 gnd.n1540 0.152939
R14042 gnd.n1542 gnd.n1541 0.152939
R14043 gnd.n1543 gnd.n1542 0.152939
R14044 gnd.n1544 gnd.n1543 0.152939
R14045 gnd.n1545 gnd.n1544 0.152939
R14046 gnd.n1546 gnd.n1545 0.152939
R14047 gnd.n1547 gnd.n1546 0.152939
R14048 gnd.n1548 gnd.n1547 0.152939
R14049 gnd.n1549 gnd.n1548 0.152939
R14050 gnd.n1550 gnd.n1549 0.152939
R14051 gnd.n1551 gnd.n1550 0.152939
R14052 gnd.n1552 gnd.n1551 0.152939
R14053 gnd.n1553 gnd.n1552 0.152939
R14054 gnd.n1554 gnd.n1553 0.152939
R14055 gnd.n1555 gnd.n1554 0.152939
R14056 gnd.n1556 gnd.n1555 0.152939
R14057 gnd.n1560 gnd.n1556 0.152939
R14058 gnd.n1561 gnd.n1560 0.152939
R14059 gnd.n1561 gnd.n1518 0.152939
R14060 gnd.n1615 gnd.n1518 0.152939
R14061 gnd.n6427 gnd.n796 0.152939
R14062 gnd.n6428 gnd.n6427 0.152939
R14063 gnd.n6429 gnd.n6428 0.152939
R14064 gnd.n6429 gnd.n790 0.152939
R14065 gnd.n6437 gnd.n790 0.152939
R14066 gnd.n6438 gnd.n6437 0.152939
R14067 gnd.n6439 gnd.n6438 0.152939
R14068 gnd.n6439 gnd.n784 0.152939
R14069 gnd.n6447 gnd.n784 0.152939
R14070 gnd.n6448 gnd.n6447 0.152939
R14071 gnd.n6449 gnd.n6448 0.152939
R14072 gnd.n6449 gnd.n778 0.152939
R14073 gnd.n6457 gnd.n778 0.152939
R14074 gnd.n6458 gnd.n6457 0.152939
R14075 gnd.n6459 gnd.n6458 0.152939
R14076 gnd.n6459 gnd.n772 0.152939
R14077 gnd.n6467 gnd.n772 0.152939
R14078 gnd.n6468 gnd.n6467 0.152939
R14079 gnd.n6469 gnd.n6468 0.152939
R14080 gnd.n6469 gnd.n766 0.152939
R14081 gnd.n6477 gnd.n766 0.152939
R14082 gnd.n6478 gnd.n6477 0.152939
R14083 gnd.n6479 gnd.n6478 0.152939
R14084 gnd.n6479 gnd.n760 0.152939
R14085 gnd.n6487 gnd.n760 0.152939
R14086 gnd.n6488 gnd.n6487 0.152939
R14087 gnd.n6489 gnd.n6488 0.152939
R14088 gnd.n6489 gnd.n754 0.152939
R14089 gnd.n6497 gnd.n754 0.152939
R14090 gnd.n6498 gnd.n6497 0.152939
R14091 gnd.n6499 gnd.n6498 0.152939
R14092 gnd.n6499 gnd.n748 0.152939
R14093 gnd.n6507 gnd.n748 0.152939
R14094 gnd.n6508 gnd.n6507 0.152939
R14095 gnd.n6509 gnd.n6508 0.152939
R14096 gnd.n6509 gnd.n742 0.152939
R14097 gnd.n6517 gnd.n742 0.152939
R14098 gnd.n6518 gnd.n6517 0.152939
R14099 gnd.n6519 gnd.n6518 0.152939
R14100 gnd.n6519 gnd.n736 0.152939
R14101 gnd.n6527 gnd.n736 0.152939
R14102 gnd.n6528 gnd.n6527 0.152939
R14103 gnd.n6529 gnd.n6528 0.152939
R14104 gnd.n6529 gnd.n730 0.152939
R14105 gnd.n6537 gnd.n730 0.152939
R14106 gnd.n6538 gnd.n6537 0.152939
R14107 gnd.n6539 gnd.n6538 0.152939
R14108 gnd.n6539 gnd.n724 0.152939
R14109 gnd.n6547 gnd.n724 0.152939
R14110 gnd.n6548 gnd.n6547 0.152939
R14111 gnd.n6549 gnd.n6548 0.152939
R14112 gnd.n6549 gnd.n718 0.152939
R14113 gnd.n6557 gnd.n718 0.152939
R14114 gnd.n6558 gnd.n6557 0.152939
R14115 gnd.n6559 gnd.n6558 0.152939
R14116 gnd.n6559 gnd.n712 0.152939
R14117 gnd.n6567 gnd.n712 0.152939
R14118 gnd.n6568 gnd.n6567 0.152939
R14119 gnd.n6569 gnd.n6568 0.152939
R14120 gnd.n6569 gnd.n706 0.152939
R14121 gnd.n6577 gnd.n706 0.152939
R14122 gnd.n6578 gnd.n6577 0.152939
R14123 gnd.n6579 gnd.n6578 0.152939
R14124 gnd.n6579 gnd.n700 0.152939
R14125 gnd.n6587 gnd.n700 0.152939
R14126 gnd.n6588 gnd.n6587 0.152939
R14127 gnd.n6589 gnd.n6588 0.152939
R14128 gnd.n6589 gnd.n694 0.152939
R14129 gnd.n6597 gnd.n694 0.152939
R14130 gnd.n6598 gnd.n6597 0.152939
R14131 gnd.n6599 gnd.n6598 0.152939
R14132 gnd.n6599 gnd.n688 0.152939
R14133 gnd.n6607 gnd.n688 0.152939
R14134 gnd.n6608 gnd.n6607 0.152939
R14135 gnd.n6609 gnd.n6608 0.152939
R14136 gnd.n6609 gnd.n682 0.152939
R14137 gnd.n6617 gnd.n682 0.152939
R14138 gnd.n6618 gnd.n6617 0.152939
R14139 gnd.n6619 gnd.n6618 0.152939
R14140 gnd.n6619 gnd.n676 0.152939
R14141 gnd.n6627 gnd.n676 0.152939
R14142 gnd.n6628 gnd.n6627 0.152939
R14143 gnd.n6629 gnd.n6628 0.152939
R14144 gnd.n6629 gnd.n670 0.152939
R14145 gnd.n6637 gnd.n670 0.152939
R14146 gnd.n6638 gnd.n6637 0.152939
R14147 gnd.n6639 gnd.n6638 0.152939
R14148 gnd.n6639 gnd.n664 0.152939
R14149 gnd.n6647 gnd.n664 0.152939
R14150 gnd.n6648 gnd.n6647 0.152939
R14151 gnd.n6649 gnd.n6648 0.152939
R14152 gnd.n6649 gnd.n658 0.152939
R14153 gnd.n6657 gnd.n658 0.152939
R14154 gnd.n6658 gnd.n6657 0.152939
R14155 gnd.n6659 gnd.n6658 0.152939
R14156 gnd.n6659 gnd.n652 0.152939
R14157 gnd.n6667 gnd.n652 0.152939
R14158 gnd.n6668 gnd.n6667 0.152939
R14159 gnd.n6669 gnd.n6668 0.152939
R14160 gnd.n6669 gnd.n646 0.152939
R14161 gnd.n6677 gnd.n646 0.152939
R14162 gnd.n6678 gnd.n6677 0.152939
R14163 gnd.n6679 gnd.n6678 0.152939
R14164 gnd.n6679 gnd.n640 0.152939
R14165 gnd.n6687 gnd.n640 0.152939
R14166 gnd.n6688 gnd.n6687 0.152939
R14167 gnd.n6689 gnd.n6688 0.152939
R14168 gnd.n6689 gnd.n634 0.152939
R14169 gnd.n6697 gnd.n634 0.152939
R14170 gnd.n6698 gnd.n6697 0.152939
R14171 gnd.n6699 gnd.n6698 0.152939
R14172 gnd.n6699 gnd.n628 0.152939
R14173 gnd.n6707 gnd.n628 0.152939
R14174 gnd.n6708 gnd.n6707 0.152939
R14175 gnd.n6709 gnd.n6708 0.152939
R14176 gnd.n6709 gnd.n622 0.152939
R14177 gnd.n6717 gnd.n622 0.152939
R14178 gnd.n6718 gnd.n6717 0.152939
R14179 gnd.n6719 gnd.n6718 0.152939
R14180 gnd.n6719 gnd.n616 0.152939
R14181 gnd.n6727 gnd.n616 0.152939
R14182 gnd.n6728 gnd.n6727 0.152939
R14183 gnd.n6729 gnd.n6728 0.152939
R14184 gnd.n6729 gnd.n610 0.152939
R14185 gnd.n6737 gnd.n610 0.152939
R14186 gnd.n6738 gnd.n6737 0.152939
R14187 gnd.n6739 gnd.n6738 0.152939
R14188 gnd.n6739 gnd.n604 0.152939
R14189 gnd.n6747 gnd.n604 0.152939
R14190 gnd.n6748 gnd.n6747 0.152939
R14191 gnd.n6749 gnd.n6748 0.152939
R14192 gnd.n6749 gnd.n598 0.152939
R14193 gnd.n6757 gnd.n598 0.152939
R14194 gnd.n6758 gnd.n6757 0.152939
R14195 gnd.n6759 gnd.n6758 0.152939
R14196 gnd.n6759 gnd.n592 0.152939
R14197 gnd.n6767 gnd.n592 0.152939
R14198 gnd.n6768 gnd.n6767 0.152939
R14199 gnd.n6769 gnd.n6768 0.152939
R14200 gnd.n6769 gnd.n586 0.152939
R14201 gnd.n6777 gnd.n586 0.152939
R14202 gnd.n6778 gnd.n6777 0.152939
R14203 gnd.n6779 gnd.n6778 0.152939
R14204 gnd.n6779 gnd.n580 0.152939
R14205 gnd.n6787 gnd.n580 0.152939
R14206 gnd.n6788 gnd.n6787 0.152939
R14207 gnd.n6789 gnd.n6788 0.152939
R14208 gnd.n6789 gnd.n574 0.152939
R14209 gnd.n6797 gnd.n574 0.152939
R14210 gnd.n6798 gnd.n6797 0.152939
R14211 gnd.n6799 gnd.n6798 0.152939
R14212 gnd.n6799 gnd.n568 0.152939
R14213 gnd.n6807 gnd.n568 0.152939
R14214 gnd.n6808 gnd.n6807 0.152939
R14215 gnd.n6809 gnd.n6808 0.152939
R14216 gnd.n6809 gnd.n562 0.152939
R14217 gnd.n6817 gnd.n562 0.152939
R14218 gnd.n6818 gnd.n6817 0.152939
R14219 gnd.n6819 gnd.n6818 0.152939
R14220 gnd.n6819 gnd.n556 0.152939
R14221 gnd.n6827 gnd.n556 0.152939
R14222 gnd.n6828 gnd.n6827 0.152939
R14223 gnd.n6829 gnd.n6828 0.152939
R14224 gnd.n6829 gnd.n550 0.152939
R14225 gnd.n6837 gnd.n550 0.152939
R14226 gnd.n6838 gnd.n6837 0.152939
R14227 gnd.n6839 gnd.n6838 0.152939
R14228 gnd.n6839 gnd.n544 0.152939
R14229 gnd.n6847 gnd.n544 0.152939
R14230 gnd.n6848 gnd.n6847 0.152939
R14231 gnd.n6849 gnd.n6848 0.152939
R14232 gnd.n6849 gnd.n538 0.152939
R14233 gnd.n6857 gnd.n538 0.152939
R14234 gnd.n6858 gnd.n6857 0.152939
R14235 gnd.n6859 gnd.n6858 0.152939
R14236 gnd.n6859 gnd.n532 0.152939
R14237 gnd.n6867 gnd.n532 0.152939
R14238 gnd.n6868 gnd.n6867 0.152939
R14239 gnd.n6869 gnd.n6868 0.152939
R14240 gnd.n6869 gnd.n526 0.152939
R14241 gnd.n6877 gnd.n526 0.152939
R14242 gnd.n6878 gnd.n6877 0.152939
R14243 gnd.n6879 gnd.n6878 0.152939
R14244 gnd.n6879 gnd.n520 0.152939
R14245 gnd.n6887 gnd.n520 0.152939
R14246 gnd.n6888 gnd.n6887 0.152939
R14247 gnd.n6889 gnd.n6888 0.152939
R14248 gnd.n6889 gnd.n514 0.152939
R14249 gnd.n6897 gnd.n514 0.152939
R14250 gnd.n6898 gnd.n6897 0.152939
R14251 gnd.n6900 gnd.n6898 0.152939
R14252 gnd.n6900 gnd.n6899 0.152939
R14253 gnd.n6899 gnd.n508 0.152939
R14254 gnd.n6909 gnd.n508 0.152939
R14255 gnd.n6910 gnd.n503 0.152939
R14256 gnd.n6918 gnd.n503 0.152939
R14257 gnd.n6919 gnd.n6918 0.152939
R14258 gnd.n6920 gnd.n6919 0.152939
R14259 gnd.n6920 gnd.n497 0.152939
R14260 gnd.n6928 gnd.n497 0.152939
R14261 gnd.n6929 gnd.n6928 0.152939
R14262 gnd.n6930 gnd.n6929 0.152939
R14263 gnd.n6930 gnd.n491 0.152939
R14264 gnd.n6938 gnd.n491 0.152939
R14265 gnd.n6939 gnd.n6938 0.152939
R14266 gnd.n6940 gnd.n6939 0.152939
R14267 gnd.n6940 gnd.n485 0.152939
R14268 gnd.n6948 gnd.n485 0.152939
R14269 gnd.n6949 gnd.n6948 0.152939
R14270 gnd.n6950 gnd.n6949 0.152939
R14271 gnd.n6950 gnd.n479 0.152939
R14272 gnd.n6958 gnd.n479 0.152939
R14273 gnd.n6959 gnd.n6958 0.152939
R14274 gnd.n6960 gnd.n6959 0.152939
R14275 gnd.n6960 gnd.n473 0.152939
R14276 gnd.n6968 gnd.n473 0.152939
R14277 gnd.n6969 gnd.n6968 0.152939
R14278 gnd.n6970 gnd.n6969 0.152939
R14279 gnd.n6970 gnd.n467 0.152939
R14280 gnd.n6978 gnd.n467 0.152939
R14281 gnd.n6979 gnd.n6978 0.152939
R14282 gnd.n6980 gnd.n6979 0.152939
R14283 gnd.n6980 gnd.n461 0.152939
R14284 gnd.n6988 gnd.n461 0.152939
R14285 gnd.n6989 gnd.n6988 0.152939
R14286 gnd.n6990 gnd.n6989 0.152939
R14287 gnd.n6990 gnd.n455 0.152939
R14288 gnd.n6998 gnd.n455 0.152939
R14289 gnd.n6999 gnd.n6998 0.152939
R14290 gnd.n7000 gnd.n6999 0.152939
R14291 gnd.n7000 gnd.n449 0.152939
R14292 gnd.n7008 gnd.n449 0.152939
R14293 gnd.n7009 gnd.n7008 0.152939
R14294 gnd.n7010 gnd.n7009 0.152939
R14295 gnd.n7010 gnd.n443 0.152939
R14296 gnd.n7018 gnd.n443 0.152939
R14297 gnd.n7019 gnd.n7018 0.152939
R14298 gnd.n7020 gnd.n7019 0.152939
R14299 gnd.n7020 gnd.n437 0.152939
R14300 gnd.n7028 gnd.n437 0.152939
R14301 gnd.n7029 gnd.n7028 0.152939
R14302 gnd.n7030 gnd.n7029 0.152939
R14303 gnd.n7030 gnd.n431 0.152939
R14304 gnd.n7038 gnd.n431 0.152939
R14305 gnd.n7039 gnd.n7038 0.152939
R14306 gnd.n7040 gnd.n7039 0.152939
R14307 gnd.n7040 gnd.n425 0.152939
R14308 gnd.n7048 gnd.n425 0.152939
R14309 gnd.n7049 gnd.n7048 0.152939
R14310 gnd.n7050 gnd.n7049 0.152939
R14311 gnd.n7050 gnd.n419 0.152939
R14312 gnd.n7058 gnd.n419 0.152939
R14313 gnd.n7059 gnd.n7058 0.152939
R14314 gnd.n7060 gnd.n7059 0.152939
R14315 gnd.n7060 gnd.n413 0.152939
R14316 gnd.n7068 gnd.n413 0.152939
R14317 gnd.n7069 gnd.n7068 0.152939
R14318 gnd.n7070 gnd.n7069 0.152939
R14319 gnd.n7070 gnd.n407 0.152939
R14320 gnd.n7078 gnd.n407 0.152939
R14321 gnd.n7079 gnd.n7078 0.152939
R14322 gnd.n7080 gnd.n7079 0.152939
R14323 gnd.n7080 gnd.n401 0.152939
R14324 gnd.n7088 gnd.n401 0.152939
R14325 gnd.n7089 gnd.n7088 0.152939
R14326 gnd.n7090 gnd.n7089 0.152939
R14327 gnd.n7090 gnd.n395 0.152939
R14328 gnd.n7098 gnd.n395 0.152939
R14329 gnd.n7099 gnd.n7098 0.152939
R14330 gnd.n7100 gnd.n7099 0.152939
R14331 gnd.n7100 gnd.n389 0.152939
R14332 gnd.n7108 gnd.n389 0.152939
R14333 gnd.n7109 gnd.n7108 0.152939
R14334 gnd.n7110 gnd.n7109 0.152939
R14335 gnd.n7110 gnd.n383 0.152939
R14336 gnd.n7119 gnd.n383 0.152939
R14337 gnd.n7120 gnd.n7119 0.152939
R14338 gnd.n7122 gnd.n7120 0.152939
R14339 gnd.n326 gnd.n305 0.152939
R14340 gnd.n327 gnd.n326 0.152939
R14341 gnd.n327 gnd.n325 0.152939
R14342 gnd.n333 gnd.n325 0.152939
R14343 gnd.n334 gnd.n333 0.152939
R14344 gnd.n335 gnd.n334 0.152939
R14345 gnd.n336 gnd.n335 0.152939
R14346 gnd.n337 gnd.n336 0.152939
R14347 gnd.n368 gnd.n337 0.152939
R14348 gnd.n369 gnd.n368 0.152939
R14349 gnd.n369 gnd.n367 0.152939
R14350 gnd.n375 gnd.n367 0.152939
R14351 gnd.n376 gnd.n375 0.152939
R14352 gnd.n377 gnd.n376 0.152939
R14353 gnd.n378 gnd.n377 0.152939
R14354 gnd.n379 gnd.n378 0.152939
R14355 gnd.n7121 gnd.n379 0.152939
R14356 gnd.n7218 gnd.n249 0.152939
R14357 gnd.n7219 gnd.n7218 0.152939
R14358 gnd.n7220 gnd.n7219 0.152939
R14359 gnd.n7220 gnd.n233 0.152939
R14360 gnd.n7234 gnd.n233 0.152939
R14361 gnd.n7235 gnd.n7234 0.152939
R14362 gnd.n7236 gnd.n7235 0.152939
R14363 gnd.n7236 gnd.n219 0.152939
R14364 gnd.n7250 gnd.n219 0.152939
R14365 gnd.n7251 gnd.n7250 0.152939
R14366 gnd.n7252 gnd.n7251 0.152939
R14367 gnd.n7252 gnd.n203 0.152939
R14368 gnd.n7266 gnd.n203 0.152939
R14369 gnd.n7267 gnd.n7266 0.152939
R14370 gnd.n7268 gnd.n7267 0.152939
R14371 gnd.n7268 gnd.n186 0.152939
R14372 gnd.n7357 gnd.n186 0.152939
R14373 gnd.n7358 gnd.n7357 0.152939
R14374 gnd.n7359 gnd.n7358 0.152939
R14375 gnd.n7359 gnd.n107 0.152939
R14376 gnd.n7439 gnd.n107 0.152939
R14377 gnd.n7438 gnd.n108 0.152939
R14378 gnd.n110 gnd.n108 0.152939
R14379 gnd.n114 gnd.n110 0.152939
R14380 gnd.n115 gnd.n114 0.152939
R14381 gnd.n116 gnd.n115 0.152939
R14382 gnd.n117 gnd.n116 0.152939
R14383 gnd.n121 gnd.n117 0.152939
R14384 gnd.n122 gnd.n121 0.152939
R14385 gnd.n123 gnd.n122 0.152939
R14386 gnd.n124 gnd.n123 0.152939
R14387 gnd.n128 gnd.n124 0.152939
R14388 gnd.n129 gnd.n128 0.152939
R14389 gnd.n130 gnd.n129 0.152939
R14390 gnd.n131 gnd.n130 0.152939
R14391 gnd.n135 gnd.n131 0.152939
R14392 gnd.n136 gnd.n135 0.152939
R14393 gnd.n137 gnd.n136 0.152939
R14394 gnd.n138 gnd.n137 0.152939
R14395 gnd.n142 gnd.n138 0.152939
R14396 gnd.n143 gnd.n142 0.152939
R14397 gnd.n144 gnd.n143 0.152939
R14398 gnd.n145 gnd.n144 0.152939
R14399 gnd.n149 gnd.n145 0.152939
R14400 gnd.n150 gnd.n149 0.152939
R14401 gnd.n151 gnd.n150 0.152939
R14402 gnd.n152 gnd.n151 0.152939
R14403 gnd.n156 gnd.n152 0.152939
R14404 gnd.n157 gnd.n156 0.152939
R14405 gnd.n158 gnd.n157 0.152939
R14406 gnd.n159 gnd.n158 0.152939
R14407 gnd.n163 gnd.n159 0.152939
R14408 gnd.n164 gnd.n163 0.152939
R14409 gnd.n165 gnd.n164 0.152939
R14410 gnd.n166 gnd.n165 0.152939
R14411 gnd.n170 gnd.n166 0.152939
R14412 gnd.n171 gnd.n170 0.152939
R14413 gnd.n7369 gnd.n171 0.152939
R14414 gnd.n7369 gnd.n7368 0.152939
R14415 gnd.n3043 gnd.n2869 0.152939
R14416 gnd.n3044 gnd.n3043 0.152939
R14417 gnd.n3045 gnd.n3044 0.152939
R14418 gnd.n3046 gnd.n3045 0.152939
R14419 gnd.n3047 gnd.n3046 0.152939
R14420 gnd.n3048 gnd.n3047 0.152939
R14421 gnd.n3049 gnd.n3048 0.152939
R14422 gnd.n3050 gnd.n3049 0.152939
R14423 gnd.n3051 gnd.n3050 0.152939
R14424 gnd.n3052 gnd.n3051 0.152939
R14425 gnd.n3053 gnd.n3052 0.152939
R14426 gnd.n3054 gnd.n3053 0.152939
R14427 gnd.n3055 gnd.n3054 0.152939
R14428 gnd.n3056 gnd.n3055 0.152939
R14429 gnd.n3058 gnd.n3056 0.152939
R14430 gnd.n3058 gnd.n3057 0.152939
R14431 gnd.n3057 gnd.n2944 0.152939
R14432 gnd.n2944 gnd.n2942 0.152939
R14433 gnd.n5590 gnd.n2942 0.152939
R14434 gnd.n5591 gnd.n5590 0.152939
R14435 gnd.n5592 gnd.n5591 0.152939
R14436 gnd.n5593 gnd.n5592 0.152939
R14437 gnd.n5593 gnd.n2934 0.152939
R14438 gnd.n5613 gnd.n2934 0.152939
R14439 gnd.n5614 gnd.n5613 0.152939
R14440 gnd.n5615 gnd.n5614 0.152939
R14441 gnd.n297 gnd.n296 0.152939
R14442 gnd.n298 gnd.n297 0.152939
R14443 gnd.n299 gnd.n298 0.152939
R14444 gnd.n309 gnd.n299 0.152939
R14445 gnd.n313 gnd.n309 0.152939
R14446 gnd.n314 gnd.n313 0.152939
R14447 gnd.n315 gnd.n314 0.152939
R14448 gnd.n316 gnd.n315 0.152939
R14449 gnd.n317 gnd.n316 0.152939
R14450 gnd.n318 gnd.n317 0.152939
R14451 gnd.n319 gnd.n318 0.152939
R14452 gnd.n341 gnd.n319 0.152939
R14453 gnd.n345 gnd.n341 0.152939
R14454 gnd.n346 gnd.n345 0.152939
R14455 gnd.n347 gnd.n346 0.152939
R14456 gnd.n348 gnd.n347 0.152939
R14457 gnd.n349 gnd.n348 0.152939
R14458 gnd.n350 gnd.n349 0.152939
R14459 gnd.n351 gnd.n350 0.152939
R14460 gnd.n352 gnd.n351 0.152939
R14461 gnd.n353 gnd.n352 0.152939
R14462 gnd.n354 gnd.n353 0.152939
R14463 gnd.n356 gnd.n354 0.152939
R14464 gnd.n356 gnd.n355 0.152939
R14465 gnd.n355 gnd.n177 0.152939
R14466 gnd.n7367 gnd.n177 0.152939
R14467 gnd.n2826 gnd.n2825 0.152939
R14468 gnd.n2827 gnd.n2826 0.152939
R14469 gnd.n2828 gnd.n2827 0.152939
R14470 gnd.n2829 gnd.n2828 0.152939
R14471 gnd.n2830 gnd.n2829 0.152939
R14472 gnd.n2831 gnd.n2830 0.152939
R14473 gnd.n2832 gnd.n2831 0.152939
R14474 gnd.n2833 gnd.n2832 0.152939
R14475 gnd.n2834 gnd.n2833 0.152939
R14476 gnd.n2835 gnd.n2834 0.152939
R14477 gnd.n2836 gnd.n2835 0.152939
R14478 gnd.n2837 gnd.n2836 0.152939
R14479 gnd.n2838 gnd.n2837 0.152939
R14480 gnd.n2839 gnd.n2838 0.152939
R14481 gnd.n2840 gnd.n2839 0.152939
R14482 gnd.n2847 gnd.n2846 0.152939
R14483 gnd.n2848 gnd.n2847 0.152939
R14484 gnd.n2849 gnd.n2848 0.152939
R14485 gnd.n2850 gnd.n2849 0.152939
R14486 gnd.n2851 gnd.n2850 0.152939
R14487 gnd.n2852 gnd.n2851 0.152939
R14488 gnd.n2853 gnd.n2852 0.152939
R14489 gnd.n2854 gnd.n2853 0.152939
R14490 gnd.n2855 gnd.n2854 0.152939
R14491 gnd.n2856 gnd.n2855 0.152939
R14492 gnd.n2857 gnd.n2856 0.152939
R14493 gnd.n2858 gnd.n2857 0.152939
R14494 gnd.n2859 gnd.n2858 0.152939
R14495 gnd.n2860 gnd.n2859 0.152939
R14496 gnd.n2861 gnd.n2860 0.152939
R14497 gnd.n2862 gnd.n2861 0.152939
R14498 gnd.n2863 gnd.n2862 0.152939
R14499 gnd.n5700 gnd.n2863 0.152939
R14500 gnd.n5700 gnd.n5699 0.152939
R14501 gnd.n5699 gnd.n5698 0.152939
R14502 gnd.n3038 gnd.n3037 0.152939
R14503 gnd.n3038 gnd.n3016 0.152939
R14504 gnd.n5494 gnd.n3016 0.152939
R14505 gnd.n5495 gnd.n5494 0.152939
R14506 gnd.n5496 gnd.n5495 0.152939
R14507 gnd.n5497 gnd.n5496 0.152939
R14508 gnd.n5497 gnd.n2987 0.152939
R14509 gnd.n5525 gnd.n2987 0.152939
R14510 gnd.n5526 gnd.n5525 0.152939
R14511 gnd.n5527 gnd.n5526 0.152939
R14512 gnd.n5528 gnd.n5527 0.152939
R14513 gnd.n5528 gnd.n2959 0.152939
R14514 gnd.n5564 gnd.n2959 0.152939
R14515 gnd.n5565 gnd.n5564 0.152939
R14516 gnd.n5566 gnd.n5565 0.152939
R14517 gnd.n5567 gnd.n5566 0.152939
R14518 gnd.n5567 gnd.n2907 0.152939
R14519 gnd.n5654 gnd.n2907 0.152939
R14520 gnd.n5655 gnd.n5654 0.152939
R14521 gnd.n5656 gnd.n5655 0.152939
R14522 gnd.n5656 gnd.n263 0.152939
R14523 gnd.n3848 gnd.n3842 0.152939
R14524 gnd.n3851 gnd.n3848 0.152939
R14525 gnd.n3852 gnd.n3851 0.152939
R14526 gnd.n3853 gnd.n3852 0.152939
R14527 gnd.n3854 gnd.n3853 0.152939
R14528 gnd.n3857 gnd.n3854 0.152939
R14529 gnd.n3858 gnd.n3857 0.152939
R14530 gnd.n3859 gnd.n3858 0.152939
R14531 gnd.n3860 gnd.n3859 0.152939
R14532 gnd.n3863 gnd.n3860 0.152939
R14533 gnd.n3864 gnd.n3863 0.152939
R14534 gnd.n3865 gnd.n3864 0.152939
R14535 gnd.n3866 gnd.n3865 0.152939
R14536 gnd.n3869 gnd.n3866 0.152939
R14537 gnd.n3870 gnd.n3869 0.152939
R14538 gnd.n3871 gnd.n3870 0.152939
R14539 gnd.n3872 gnd.n3871 0.152939
R14540 gnd.n3875 gnd.n3872 0.152939
R14541 gnd.n3876 gnd.n3875 0.152939
R14542 gnd.n3877 gnd.n3876 0.152939
R14543 gnd.n3878 gnd.n3877 0.152939
R14544 gnd.n3881 gnd.n3878 0.152939
R14545 gnd.n3882 gnd.n3881 0.152939
R14546 gnd.n3883 gnd.n3882 0.152939
R14547 gnd.n3884 gnd.n3883 0.152939
R14548 gnd.n3884 gnd.n3524 0.152939
R14549 gnd.n4628 gnd.n3524 0.152939
R14550 gnd.n4629 gnd.n4628 0.152939
R14551 gnd.n4630 gnd.n4629 0.152939
R14552 gnd.n4630 gnd.n3511 0.152939
R14553 gnd.n4644 gnd.n3511 0.152939
R14554 gnd.n4645 gnd.n4644 0.152939
R14555 gnd.n4646 gnd.n4645 0.152939
R14556 gnd.n4646 gnd.n3498 0.152939
R14557 gnd.n4660 gnd.n3498 0.152939
R14558 gnd.n4661 gnd.n4660 0.152939
R14559 gnd.n4662 gnd.n4661 0.152939
R14560 gnd.n4662 gnd.n3484 0.152939
R14561 gnd.n4676 gnd.n3484 0.152939
R14562 gnd.n4677 gnd.n4676 0.152939
R14563 gnd.n4678 gnd.n4677 0.152939
R14564 gnd.n4678 gnd.n3470 0.152939
R14565 gnd.n4692 gnd.n3470 0.152939
R14566 gnd.n4693 gnd.n4692 0.152939
R14567 gnd.n4694 gnd.n4693 0.152939
R14568 gnd.n4694 gnd.n3457 0.152939
R14569 gnd.n4708 gnd.n3457 0.152939
R14570 gnd.n4709 gnd.n4708 0.152939
R14571 gnd.n4710 gnd.n4709 0.152939
R14572 gnd.n4711 gnd.n4710 0.152939
R14573 gnd.n4711 gnd.n3428 0.152939
R14574 gnd.n4841 gnd.n3428 0.152939
R14575 gnd.n4842 gnd.n4841 0.152939
R14576 gnd.n4843 gnd.n4842 0.152939
R14577 gnd.n4843 gnd.n3416 0.152939
R14578 gnd.n4857 gnd.n3416 0.152939
R14579 gnd.n4858 gnd.n4857 0.152939
R14580 gnd.n4859 gnd.n4858 0.152939
R14581 gnd.n4859 gnd.n3403 0.152939
R14582 gnd.n4873 gnd.n3403 0.152939
R14583 gnd.n4874 gnd.n4873 0.152939
R14584 gnd.n4875 gnd.n4874 0.152939
R14585 gnd.n4875 gnd.n3391 0.152939
R14586 gnd.n4889 gnd.n3391 0.152939
R14587 gnd.n4890 gnd.n4889 0.152939
R14588 gnd.n4891 gnd.n4890 0.152939
R14589 gnd.n4892 gnd.n4891 0.152939
R14590 gnd.n4892 gnd.n3362 0.152939
R14591 gnd.n5018 gnd.n3362 0.152939
R14592 gnd.n5019 gnd.n5018 0.152939
R14593 gnd.n5020 gnd.n5019 0.152939
R14594 gnd.n5020 gnd.n3349 0.152939
R14595 gnd.n5034 gnd.n3349 0.152939
R14596 gnd.n5035 gnd.n5034 0.152939
R14597 gnd.n5036 gnd.n5035 0.152939
R14598 gnd.n5036 gnd.n3334 0.152939
R14599 gnd.n5050 gnd.n3334 0.152939
R14600 gnd.n5051 gnd.n5050 0.152939
R14601 gnd.n5052 gnd.n5051 0.152939
R14602 gnd.n5052 gnd.n3320 0.152939
R14603 gnd.n5066 gnd.n3320 0.152939
R14604 gnd.n5067 gnd.n5066 0.152939
R14605 gnd.n5068 gnd.n5067 0.152939
R14606 gnd.n5069 gnd.n5068 0.152939
R14607 gnd.n5069 gnd.n3290 0.152939
R14608 gnd.n5352 gnd.n3290 0.152939
R14609 gnd.n5353 gnd.n5352 0.152939
R14610 gnd.n5354 gnd.n5353 0.152939
R14611 gnd.n5354 gnd.n3278 0.152939
R14612 gnd.n5368 gnd.n3278 0.152939
R14613 gnd.n5369 gnd.n5368 0.152939
R14614 gnd.n5370 gnd.n5369 0.152939
R14615 gnd.n5370 gnd.n3265 0.152939
R14616 gnd.n5384 gnd.n3265 0.152939
R14617 gnd.n5385 gnd.n5384 0.152939
R14618 gnd.n5386 gnd.n5385 0.152939
R14619 gnd.n5386 gnd.n3252 0.152939
R14620 gnd.n5400 gnd.n3252 0.152939
R14621 gnd.n5401 gnd.n5400 0.152939
R14622 gnd.n5402 gnd.n5401 0.152939
R14623 gnd.n5402 gnd.n3239 0.152939
R14624 gnd.n5416 gnd.n3239 0.152939
R14625 gnd.n5417 gnd.n5416 0.152939
R14626 gnd.n5418 gnd.n5417 0.152939
R14627 gnd.n5418 gnd.n3227 0.152939
R14628 gnd.n5434 gnd.n3227 0.152939
R14629 gnd.n5435 gnd.n5434 0.152939
R14630 gnd.n5436 gnd.n5435 0.152939
R14631 gnd.n5438 gnd.n5436 0.152939
R14632 gnd.n5438 gnd.n5437 0.152939
R14633 gnd.n5437 gnd.n2788 0.152939
R14634 gnd.n2789 gnd.n2788 0.152939
R14635 gnd.n2790 gnd.n2789 0.152939
R14636 gnd.n3030 gnd.n2790 0.152939
R14637 gnd.n3031 gnd.n3030 0.152939
R14638 gnd.n3032 gnd.n3031 0.152939
R14639 gnd.n3032 gnd.n3026 0.152939
R14640 gnd.n5483 gnd.n3026 0.152939
R14641 gnd.n5484 gnd.n5483 0.152939
R14642 gnd.n5485 gnd.n5484 0.152939
R14643 gnd.n5486 gnd.n5485 0.152939
R14644 gnd.n5486 gnd.n2998 0.152939
R14645 gnd.n5514 gnd.n2998 0.152939
R14646 gnd.n5515 gnd.n5514 0.152939
R14647 gnd.n5516 gnd.n5515 0.152939
R14648 gnd.n5517 gnd.n5516 0.152939
R14649 gnd.n5517 gnd.n2970 0.152939
R14650 gnd.n5545 gnd.n2970 0.152939
R14651 gnd.n5546 gnd.n5545 0.152939
R14652 gnd.n5547 gnd.n5546 0.152939
R14653 gnd.n5548 gnd.n5547 0.152939
R14654 gnd.n5549 gnd.n5548 0.152939
R14655 gnd.n5551 gnd.n5549 0.152939
R14656 gnd.n5551 gnd.n5550 0.152939
R14657 gnd.n5550 gnd.n2918 0.152939
R14658 gnd.n2919 gnd.n2918 0.152939
R14659 gnd.n2920 gnd.n2919 0.152939
R14660 gnd.n2921 gnd.n2920 0.152939
R14661 gnd.n2560 gnd.n2559 0.152939
R14662 gnd.n2578 gnd.n2560 0.152939
R14663 gnd.n2579 gnd.n2578 0.152939
R14664 gnd.n2580 gnd.n2579 0.152939
R14665 gnd.n2581 gnd.n2580 0.152939
R14666 gnd.n2600 gnd.n2581 0.152939
R14667 gnd.n2601 gnd.n2600 0.152939
R14668 gnd.n2602 gnd.n2601 0.152939
R14669 gnd.n2603 gnd.n2602 0.152939
R14670 gnd.n2621 gnd.n2603 0.152939
R14671 gnd.n2622 gnd.n2621 0.152939
R14672 gnd.n2623 gnd.n2622 0.152939
R14673 gnd.n2624 gnd.n2623 0.152939
R14674 gnd.n2643 gnd.n2624 0.152939
R14675 gnd.n2644 gnd.n2643 0.152939
R14676 gnd.n2645 gnd.n2644 0.152939
R14677 gnd.n2646 gnd.n2645 0.152939
R14678 gnd.n2664 gnd.n2646 0.152939
R14679 gnd.n2665 gnd.n2664 0.152939
R14680 gnd.n2666 gnd.n2665 0.152939
R14681 gnd.n2667 gnd.n2666 0.152939
R14682 gnd.n3690 gnd.n3689 0.152939
R14683 gnd.n3691 gnd.n3690 0.152939
R14684 gnd.n3692 gnd.n3691 0.152939
R14685 gnd.n3693 gnd.n3692 0.152939
R14686 gnd.n3694 gnd.n3693 0.152939
R14687 gnd.n3695 gnd.n3694 0.152939
R14688 gnd.n3696 gnd.n3695 0.152939
R14689 gnd.n3697 gnd.n3696 0.152939
R14690 gnd.n3698 gnd.n3697 0.152939
R14691 gnd.n3699 gnd.n3698 0.152939
R14692 gnd.n3700 gnd.n3699 0.152939
R14693 gnd.n3701 gnd.n3700 0.152939
R14694 gnd.n3702 gnd.n3701 0.152939
R14695 gnd.n3703 gnd.n3702 0.152939
R14696 gnd.n3704 gnd.n3703 0.152939
R14697 gnd.n4303 gnd.n4302 0.152939
R14698 gnd.n4302 gnd.n3709 0.152939
R14699 gnd.n3710 gnd.n3709 0.152939
R14700 gnd.n3711 gnd.n3710 0.152939
R14701 gnd.n3712 gnd.n3711 0.152939
R14702 gnd.n3713 gnd.n3712 0.152939
R14703 gnd.n3714 gnd.n3713 0.152939
R14704 gnd.n3715 gnd.n3714 0.152939
R14705 gnd.n3716 gnd.n3715 0.152939
R14706 gnd.n3717 gnd.n3716 0.152939
R14707 gnd.n3718 gnd.n3717 0.152939
R14708 gnd.n3719 gnd.n3718 0.152939
R14709 gnd.n3720 gnd.n3719 0.152939
R14710 gnd.n3721 gnd.n3720 0.152939
R14711 gnd.n3722 gnd.n3721 0.152939
R14712 gnd.n3723 gnd.n3722 0.152939
R14713 gnd.n3724 gnd.n3723 0.152939
R14714 gnd.n3725 gnd.n3724 0.152939
R14715 gnd.n4262 gnd.n3725 0.152939
R14716 gnd.n4262 gnd.n4261 0.152939
R14717 gnd.n3998 gnd.n3808 0.152939
R14718 gnd.n4056 gnd.n3808 0.152939
R14719 gnd.n4057 gnd.n4056 0.152939
R14720 gnd.n4058 gnd.n4057 0.152939
R14721 gnd.n4058 gnd.n3806 0.152939
R14722 gnd.n4071 gnd.n3806 0.152939
R14723 gnd.n4072 gnd.n4071 0.152939
R14724 gnd.n4073 gnd.n4072 0.152939
R14725 gnd.n4073 gnd.n3799 0.152939
R14726 gnd.n4087 gnd.n3799 0.152939
R14727 gnd.n4088 gnd.n4087 0.152939
R14728 gnd.n4089 gnd.n4088 0.152939
R14729 gnd.n4089 gnd.n3793 0.152939
R14730 gnd.n4103 gnd.n3793 0.152939
R14731 gnd.n4104 gnd.n4103 0.152939
R14732 gnd.n4105 gnd.n4104 0.152939
R14733 gnd.n4105 gnd.n3786 0.152939
R14734 gnd.n4119 gnd.n3786 0.152939
R14735 gnd.n4120 gnd.n4119 0.152939
R14736 gnd.n4121 gnd.n4120 0.152939
R14737 gnd.n4121 gnd.n3780 0.152939
R14738 gnd.n4135 gnd.n3780 0.152939
R14739 gnd.n4136 gnd.n4135 0.152939
R14740 gnd.n4137 gnd.n4136 0.152939
R14741 gnd.n4137 gnd.n3773 0.152939
R14742 gnd.n4153 gnd.n3773 0.152939
R14743 gnd.n4037 gnd.n3978 0.152939
R14744 gnd.n3979 gnd.n3978 0.152939
R14745 gnd.n3980 gnd.n3979 0.152939
R14746 gnd.n3981 gnd.n3980 0.152939
R14747 gnd.n3982 gnd.n3981 0.152939
R14748 gnd.n3983 gnd.n3982 0.152939
R14749 gnd.n3984 gnd.n3983 0.152939
R14750 gnd.n3985 gnd.n3984 0.152939
R14751 gnd.n3986 gnd.n3985 0.152939
R14752 gnd.n3987 gnd.n3986 0.152939
R14753 gnd.n3988 gnd.n3987 0.152939
R14754 gnd.n3989 gnd.n3988 0.152939
R14755 gnd.n3990 gnd.n3989 0.152939
R14756 gnd.n3991 gnd.n3990 0.152939
R14757 gnd.n3992 gnd.n3991 0.152939
R14758 gnd.n4002 gnd.n3992 0.152939
R14759 gnd.n4002 gnd.n4001 0.152939
R14760 gnd.n4001 gnd.n4000 0.152939
R14761 gnd.n4043 gnd.n4038 0.152939
R14762 gnd.n4043 gnd.n4042 0.152939
R14763 gnd.n4042 gnd.n4041 0.152939
R14764 gnd.n4041 gnd.n4039 0.152939
R14765 gnd.n4039 gnd.n2424 0.152939
R14766 gnd.n2425 gnd.n2424 0.152939
R14767 gnd.n2426 gnd.n2425 0.152939
R14768 gnd.n2444 gnd.n2426 0.152939
R14769 gnd.n2445 gnd.n2444 0.152939
R14770 gnd.n2446 gnd.n2445 0.152939
R14771 gnd.n2447 gnd.n2446 0.152939
R14772 gnd.n2466 gnd.n2447 0.152939
R14773 gnd.n2467 gnd.n2466 0.152939
R14774 gnd.n2468 gnd.n2467 0.152939
R14775 gnd.n2469 gnd.n2468 0.152939
R14776 gnd.n2487 gnd.n2469 0.152939
R14777 gnd.n2488 gnd.n2487 0.152939
R14778 gnd.n2489 gnd.n2488 0.152939
R14779 gnd.n2490 gnd.n2489 0.152939
R14780 gnd.n2509 gnd.n2490 0.152939
R14781 gnd.n2510 gnd.n2509 0.152939
R14782 gnd.n2511 gnd.n2510 0.152939
R14783 gnd.n2512 gnd.n2511 0.152939
R14784 gnd.n2528 gnd.n2512 0.152939
R14785 gnd.n2529 gnd.n2528 0.152939
R14786 gnd.n2530 gnd.n2529 0.152939
R14787 gnd.n2547 gnd.n2531 0.152939
R14788 gnd.n2548 gnd.n2547 0.152939
R14789 gnd.n2549 gnd.n2548 0.152939
R14790 gnd.n2550 gnd.n2549 0.152939
R14791 gnd.n2567 gnd.n2550 0.152939
R14792 gnd.n2568 gnd.n2567 0.152939
R14793 gnd.n2569 gnd.n2568 0.152939
R14794 gnd.n2570 gnd.n2569 0.152939
R14795 gnd.n2589 gnd.n2570 0.152939
R14796 gnd.n2590 gnd.n2589 0.152939
R14797 gnd.n2591 gnd.n2590 0.152939
R14798 gnd.n2592 gnd.n2591 0.152939
R14799 gnd.n2610 gnd.n2592 0.152939
R14800 gnd.n2611 gnd.n2610 0.152939
R14801 gnd.n2612 gnd.n2611 0.152939
R14802 gnd.n2613 gnd.n2612 0.152939
R14803 gnd.n2632 gnd.n2613 0.152939
R14804 gnd.n2633 gnd.n2632 0.152939
R14805 gnd.n2634 gnd.n2633 0.152939
R14806 gnd.n2635 gnd.n2634 0.152939
R14807 gnd.n2654 gnd.n2635 0.152939
R14808 gnd.n2655 gnd.n2654 0.152939
R14809 gnd.n2656 gnd.n2655 0.152939
R14810 gnd.n2657 gnd.n2656 0.152939
R14811 gnd.n2674 gnd.n2657 0.152939
R14812 gnd.n5907 gnd.n2674 0.152939
R14813 gnd.n6066 gnd.n2398 0.152939
R14814 gnd.n6066 gnd.n6065 0.152939
R14815 gnd.n6065 gnd.n6064 0.152939
R14816 gnd.n6064 gnd.n2401 0.152939
R14817 gnd.n4064 gnd.n2401 0.152939
R14818 gnd.n4065 gnd.n4064 0.152939
R14819 gnd.n4065 gnd.n3803 0.152939
R14820 gnd.n4079 gnd.n3803 0.152939
R14821 gnd.n4080 gnd.n4079 0.152939
R14822 gnd.n4081 gnd.n4080 0.152939
R14823 gnd.n4081 gnd.n3796 0.152939
R14824 gnd.n4095 gnd.n3796 0.152939
R14825 gnd.n4096 gnd.n4095 0.152939
R14826 gnd.n4097 gnd.n4096 0.152939
R14827 gnd.n4097 gnd.n3790 0.152939
R14828 gnd.n4111 gnd.n3790 0.152939
R14829 gnd.n4112 gnd.n4111 0.152939
R14830 gnd.n4113 gnd.n4112 0.152939
R14831 gnd.n4113 gnd.n3783 0.152939
R14832 gnd.n4127 gnd.n3783 0.152939
R14833 gnd.n4128 gnd.n4127 0.152939
R14834 gnd.n4129 gnd.n4128 0.152939
R14835 gnd.n4129 gnd.n3777 0.152939
R14836 gnd.n4143 gnd.n3777 0.152939
R14837 gnd.n4144 gnd.n4143 0.152939
R14838 gnd.n4147 gnd.n4144 0.152939
R14839 gnd.n4162 gnd.n3770 0.152939
R14840 gnd.n4163 gnd.n4162 0.152939
R14841 gnd.n4164 gnd.n4163 0.152939
R14842 gnd.n4164 gnd.n3764 0.152939
R14843 gnd.n4178 gnd.n3764 0.152939
R14844 gnd.n4179 gnd.n4178 0.152939
R14845 gnd.n4180 gnd.n4179 0.152939
R14846 gnd.n4180 gnd.n3757 0.152939
R14847 gnd.n4194 gnd.n3757 0.152939
R14848 gnd.n4195 gnd.n4194 0.152939
R14849 gnd.n4196 gnd.n4195 0.152939
R14850 gnd.n4196 gnd.n3751 0.152939
R14851 gnd.n4210 gnd.n3751 0.152939
R14852 gnd.n4211 gnd.n4210 0.152939
R14853 gnd.n4212 gnd.n4211 0.152939
R14854 gnd.n4212 gnd.n3744 0.152939
R14855 gnd.n4226 gnd.n3744 0.152939
R14856 gnd.n4227 gnd.n4226 0.152939
R14857 gnd.n4228 gnd.n4227 0.152939
R14858 gnd.n4228 gnd.n3738 0.152939
R14859 gnd.n4242 gnd.n3738 0.152939
R14860 gnd.n4243 gnd.n4242 0.152939
R14861 gnd.n4245 gnd.n4243 0.152939
R14862 gnd.n4245 gnd.n4244 0.152939
R14863 gnd.n4244 gnd.n3730 0.152939
R14864 gnd.n4260 gnd.n3730 0.152939
R14865 gnd.n2356 gnd.n2355 0.152939
R14866 gnd.n2357 gnd.n2356 0.152939
R14867 gnd.n2358 gnd.n2357 0.152939
R14868 gnd.n2359 gnd.n2358 0.152939
R14869 gnd.n2360 gnd.n2359 0.152939
R14870 gnd.n2361 gnd.n2360 0.152939
R14871 gnd.n2362 gnd.n2361 0.152939
R14872 gnd.n2363 gnd.n2362 0.152939
R14873 gnd.n2364 gnd.n2363 0.152939
R14874 gnd.n2365 gnd.n2364 0.152939
R14875 gnd.n2366 gnd.n2365 0.152939
R14876 gnd.n2367 gnd.n2366 0.152939
R14877 gnd.n2368 gnd.n2367 0.152939
R14878 gnd.n2369 gnd.n2368 0.152939
R14879 gnd.n2370 gnd.n2369 0.152939
R14880 gnd.n2371 gnd.n2370 0.152939
R14881 gnd.n2372 gnd.n2371 0.152939
R14882 gnd.n2375 gnd.n2372 0.152939
R14883 gnd.n2376 gnd.n2375 0.152939
R14884 gnd.n2377 gnd.n2376 0.152939
R14885 gnd.n2378 gnd.n2377 0.152939
R14886 gnd.n2379 gnd.n2378 0.152939
R14887 gnd.n2380 gnd.n2379 0.152939
R14888 gnd.n2381 gnd.n2380 0.152939
R14889 gnd.n2382 gnd.n2381 0.152939
R14890 gnd.n2383 gnd.n2382 0.152939
R14891 gnd.n2384 gnd.n2383 0.152939
R14892 gnd.n2385 gnd.n2384 0.152939
R14893 gnd.n2386 gnd.n2385 0.152939
R14894 gnd.n2387 gnd.n2386 0.152939
R14895 gnd.n2388 gnd.n2387 0.152939
R14896 gnd.n2389 gnd.n2388 0.152939
R14897 gnd.n2390 gnd.n2389 0.152939
R14898 gnd.n2391 gnd.n2390 0.152939
R14899 gnd.n2392 gnd.n2391 0.152939
R14900 gnd.n6074 gnd.n2392 0.152939
R14901 gnd.n6074 gnd.n6073 0.152939
R14902 gnd.n6073 gnd.n6072 0.152939
R14903 gnd.n4049 gnd.n4047 0.152939
R14904 gnd.n4049 gnd.n4048 0.152939
R14905 gnd.n4048 gnd.n2412 0.152939
R14906 gnd.n2413 gnd.n2412 0.152939
R14907 gnd.n2414 gnd.n2413 0.152939
R14908 gnd.n2434 gnd.n2414 0.152939
R14909 gnd.n2435 gnd.n2434 0.152939
R14910 gnd.n2436 gnd.n2435 0.152939
R14911 gnd.n2437 gnd.n2436 0.152939
R14912 gnd.n2455 gnd.n2437 0.152939
R14913 gnd.n2456 gnd.n2455 0.152939
R14914 gnd.n2457 gnd.n2456 0.152939
R14915 gnd.n2458 gnd.n2457 0.152939
R14916 gnd.n2477 gnd.n2458 0.152939
R14917 gnd.n2478 gnd.n2477 0.152939
R14918 gnd.n2479 gnd.n2478 0.152939
R14919 gnd.n2480 gnd.n2479 0.152939
R14920 gnd.n2498 gnd.n2480 0.152939
R14921 gnd.n2499 gnd.n2498 0.152939
R14922 gnd.n2500 gnd.n2499 0.152939
R14923 gnd.n2501 gnd.n2500 0.152939
R14924 gnd.n3969 gnd.n3813 0.152939
R14925 gnd.n3816 gnd.n3813 0.152939
R14926 gnd.n3817 gnd.n3816 0.152939
R14927 gnd.n3818 gnd.n3817 0.152939
R14928 gnd.n3819 gnd.n3818 0.152939
R14929 gnd.n3822 gnd.n3819 0.152939
R14930 gnd.n3823 gnd.n3822 0.152939
R14931 gnd.n3824 gnd.n3823 0.152939
R14932 gnd.n3825 gnd.n3824 0.152939
R14933 gnd.n3828 gnd.n3825 0.152939
R14934 gnd.n3829 gnd.n3828 0.152939
R14935 gnd.n3830 gnd.n3829 0.152939
R14936 gnd.n3831 gnd.n3830 0.152939
R14937 gnd.n3834 gnd.n3831 0.152939
R14938 gnd.n3835 gnd.n3834 0.152939
R14939 gnd.n3836 gnd.n3835 0.152939
R14940 gnd.n3837 gnd.n3836 0.152939
R14941 gnd.n802 gnd.n801 0.152939
R14942 gnd.n803 gnd.n802 0.152939
R14943 gnd.n808 gnd.n803 0.152939
R14944 gnd.n809 gnd.n808 0.152939
R14945 gnd.n810 gnd.n809 0.152939
R14946 gnd.n811 gnd.n810 0.152939
R14947 gnd.n816 gnd.n811 0.152939
R14948 gnd.n817 gnd.n816 0.152939
R14949 gnd.n818 gnd.n817 0.152939
R14950 gnd.n819 gnd.n818 0.152939
R14951 gnd.n824 gnd.n819 0.152939
R14952 gnd.n825 gnd.n824 0.152939
R14953 gnd.n826 gnd.n825 0.152939
R14954 gnd.n827 gnd.n826 0.152939
R14955 gnd.n832 gnd.n827 0.152939
R14956 gnd.n833 gnd.n832 0.152939
R14957 gnd.n834 gnd.n833 0.152939
R14958 gnd.n835 gnd.n834 0.152939
R14959 gnd.n840 gnd.n835 0.152939
R14960 gnd.n841 gnd.n840 0.152939
R14961 gnd.n842 gnd.n841 0.152939
R14962 gnd.n843 gnd.n842 0.152939
R14963 gnd.n848 gnd.n843 0.152939
R14964 gnd.n849 gnd.n848 0.152939
R14965 gnd.n850 gnd.n849 0.152939
R14966 gnd.n851 gnd.n850 0.152939
R14967 gnd.n856 gnd.n851 0.152939
R14968 gnd.n857 gnd.n856 0.152939
R14969 gnd.n858 gnd.n857 0.152939
R14970 gnd.n859 gnd.n858 0.152939
R14971 gnd.n864 gnd.n859 0.152939
R14972 gnd.n865 gnd.n864 0.152939
R14973 gnd.n866 gnd.n865 0.152939
R14974 gnd.n867 gnd.n866 0.152939
R14975 gnd.n872 gnd.n867 0.152939
R14976 gnd.n873 gnd.n872 0.152939
R14977 gnd.n874 gnd.n873 0.152939
R14978 gnd.n875 gnd.n874 0.152939
R14979 gnd.n880 gnd.n875 0.152939
R14980 gnd.n881 gnd.n880 0.152939
R14981 gnd.n882 gnd.n881 0.152939
R14982 gnd.n883 gnd.n882 0.152939
R14983 gnd.n888 gnd.n883 0.152939
R14984 gnd.n889 gnd.n888 0.152939
R14985 gnd.n890 gnd.n889 0.152939
R14986 gnd.n891 gnd.n890 0.152939
R14987 gnd.n896 gnd.n891 0.152939
R14988 gnd.n897 gnd.n896 0.152939
R14989 gnd.n898 gnd.n897 0.152939
R14990 gnd.n899 gnd.n898 0.152939
R14991 gnd.n904 gnd.n899 0.152939
R14992 gnd.n905 gnd.n904 0.152939
R14993 gnd.n906 gnd.n905 0.152939
R14994 gnd.n907 gnd.n906 0.152939
R14995 gnd.n912 gnd.n907 0.152939
R14996 gnd.n913 gnd.n912 0.152939
R14997 gnd.n914 gnd.n913 0.152939
R14998 gnd.n915 gnd.n914 0.152939
R14999 gnd.n920 gnd.n915 0.152939
R15000 gnd.n921 gnd.n920 0.152939
R15001 gnd.n922 gnd.n921 0.152939
R15002 gnd.n923 gnd.n922 0.152939
R15003 gnd.n928 gnd.n923 0.152939
R15004 gnd.n929 gnd.n928 0.152939
R15005 gnd.n930 gnd.n929 0.152939
R15006 gnd.n931 gnd.n930 0.152939
R15007 gnd.n936 gnd.n931 0.152939
R15008 gnd.n937 gnd.n936 0.152939
R15009 gnd.n938 gnd.n937 0.152939
R15010 gnd.n939 gnd.n938 0.152939
R15011 gnd.n944 gnd.n939 0.152939
R15012 gnd.n945 gnd.n944 0.152939
R15013 gnd.n946 gnd.n945 0.152939
R15014 gnd.n947 gnd.n946 0.152939
R15015 gnd.n952 gnd.n947 0.152939
R15016 gnd.n953 gnd.n952 0.152939
R15017 gnd.n954 gnd.n953 0.152939
R15018 gnd.n955 gnd.n954 0.152939
R15019 gnd.n960 gnd.n955 0.152939
R15020 gnd.n961 gnd.n960 0.152939
R15021 gnd.n962 gnd.n961 0.152939
R15022 gnd.n963 gnd.n962 0.152939
R15023 gnd.n3812 gnd.n963 0.152939
R15024 gnd.n3970 gnd.n3812 0.152939
R15025 gnd.n5470 gnd.n3083 0.152939
R15026 gnd.n5466 gnd.n3083 0.152939
R15027 gnd.n5466 gnd.n5465 0.152939
R15028 gnd.n5465 gnd.n5464 0.152939
R15029 gnd.n5464 gnd.n3211 0.152939
R15030 gnd.n5457 gnd.n3211 0.152939
R15031 gnd.n5457 gnd.n5456 0.152939
R15032 gnd.n5456 gnd.n5455 0.152939
R15033 gnd.n5455 gnd.n5448 0.152939
R15034 gnd.n4636 gnd.n3518 0.152939
R15035 gnd.n4637 gnd.n4636 0.152939
R15036 gnd.n4638 gnd.n4637 0.152939
R15037 gnd.n4638 gnd.n3504 0.152939
R15038 gnd.n4652 gnd.n3504 0.152939
R15039 gnd.n4653 gnd.n4652 0.152939
R15040 gnd.n4654 gnd.n4653 0.152939
R15041 gnd.n4654 gnd.n3491 0.152939
R15042 gnd.n4668 gnd.n3491 0.152939
R15043 gnd.n4669 gnd.n4668 0.152939
R15044 gnd.n4670 gnd.n4669 0.152939
R15045 gnd.n4670 gnd.n3478 0.152939
R15046 gnd.n4684 gnd.n3478 0.152939
R15047 gnd.n4685 gnd.n4684 0.152939
R15048 gnd.n4686 gnd.n4685 0.152939
R15049 gnd.n4686 gnd.n3464 0.152939
R15050 gnd.n4700 gnd.n3464 0.152939
R15051 gnd.n4701 gnd.n4700 0.152939
R15052 gnd.n4702 gnd.n4701 0.152939
R15053 gnd.n4702 gnd.n3450 0.152939
R15054 gnd.n4718 gnd.n3450 0.152939
R15055 gnd.n4719 gnd.n4718 0.152939
R15056 gnd.n4721 gnd.n4719 0.152939
R15057 gnd.n4721 gnd.n4720 0.152939
R15058 gnd.n4720 gnd.n3422 0.152939
R15059 gnd.n4849 gnd.n3422 0.152939
R15060 gnd.n4850 gnd.n4849 0.152939
R15061 gnd.n4851 gnd.n4850 0.152939
R15062 gnd.n4851 gnd.n3410 0.152939
R15063 gnd.n4865 gnd.n3410 0.152939
R15064 gnd.n4866 gnd.n4865 0.152939
R15065 gnd.n4867 gnd.n4866 0.152939
R15066 gnd.n4867 gnd.n3397 0.152939
R15067 gnd.n4881 gnd.n3397 0.152939
R15068 gnd.n4882 gnd.n4881 0.152939
R15069 gnd.n4883 gnd.n4882 0.152939
R15070 gnd.n4883 gnd.n3383 0.152939
R15071 gnd.n4899 gnd.n3383 0.152939
R15072 gnd.n4900 gnd.n4899 0.152939
R15073 gnd.n4902 gnd.n4900 0.152939
R15074 gnd.n4902 gnd.n4901 0.152939
R15075 gnd.n4901 gnd.n3355 0.152939
R15076 gnd.n5026 gnd.n3355 0.152939
R15077 gnd.n5027 gnd.n5026 0.152939
R15078 gnd.n5028 gnd.n5027 0.152939
R15079 gnd.n5028 gnd.n3341 0.152939
R15080 gnd.n5042 gnd.n3341 0.152939
R15081 gnd.n5043 gnd.n5042 0.152939
R15082 gnd.n5044 gnd.n5043 0.152939
R15083 gnd.n5044 gnd.n3326 0.152939
R15084 gnd.n5058 gnd.n3326 0.152939
R15085 gnd.n5059 gnd.n5058 0.152939
R15086 gnd.n5060 gnd.n5059 0.152939
R15087 gnd.n5060 gnd.n3311 0.152939
R15088 gnd.n5076 gnd.n3311 0.152939
R15089 gnd.n5077 gnd.n5076 0.152939
R15090 gnd.n5079 gnd.n5077 0.152939
R15091 gnd.n5079 gnd.n5078 0.152939
R15092 gnd.n5078 gnd.n3284 0.152939
R15093 gnd.n5360 gnd.n3284 0.152939
R15094 gnd.n5361 gnd.n5360 0.152939
R15095 gnd.n5362 gnd.n5361 0.152939
R15096 gnd.n5362 gnd.n3271 0.152939
R15097 gnd.n5376 gnd.n3271 0.152939
R15098 gnd.n5377 gnd.n5376 0.152939
R15099 gnd.n5378 gnd.n5377 0.152939
R15100 gnd.n5378 gnd.n3259 0.152939
R15101 gnd.n5392 gnd.n3259 0.152939
R15102 gnd.n5393 gnd.n5392 0.152939
R15103 gnd.n5394 gnd.n5393 0.152939
R15104 gnd.n5394 gnd.n3247 0.152939
R15105 gnd.n5408 gnd.n3247 0.152939
R15106 gnd.n5409 gnd.n5408 0.152939
R15107 gnd.n5410 gnd.n5409 0.152939
R15108 gnd.n5410 gnd.n3234 0.152939
R15109 gnd.n5424 gnd.n3234 0.152939
R15110 gnd.n5425 gnd.n5424 0.152939
R15111 gnd.n5428 gnd.n5425 0.152939
R15112 gnd.n5428 gnd.n5427 0.152939
R15113 gnd.n5427 gnd.n5426 0.152939
R15114 gnd.n5426 gnd.n3219 0.152939
R15115 gnd.n5447 gnd.n3219 0.152939
R15116 gnd.n4604 gnd.n4603 0.152939
R15117 gnd.n4604 gnd.n3550 0.152939
R15118 gnd.n4610 gnd.n3550 0.152939
R15119 gnd.n4611 gnd.n4610 0.152939
R15120 gnd.n4612 gnd.n4611 0.152939
R15121 gnd.n4612 gnd.n3544 0.152939
R15122 gnd.n4619 gnd.n3544 0.152939
R15123 gnd.n4620 gnd.n4619 0.152939
R15124 gnd.n4621 gnd.n4620 0.152939
R15125 gnd.n4156 gnd.n4155 0.152939
R15126 gnd.n4156 gnd.n3767 0.152939
R15127 gnd.n4170 gnd.n3767 0.152939
R15128 gnd.n4171 gnd.n4170 0.152939
R15129 gnd.n4172 gnd.n4171 0.152939
R15130 gnd.n4172 gnd.n3760 0.152939
R15131 gnd.n4186 gnd.n3760 0.152939
R15132 gnd.n4187 gnd.n4186 0.152939
R15133 gnd.n4188 gnd.n4187 0.152939
R15134 gnd.n4188 gnd.n3754 0.152939
R15135 gnd.n4202 gnd.n3754 0.152939
R15136 gnd.n4203 gnd.n4202 0.152939
R15137 gnd.n4204 gnd.n4203 0.152939
R15138 gnd.n4204 gnd.n3747 0.152939
R15139 gnd.n4218 gnd.n3747 0.152939
R15140 gnd.n4219 gnd.n4218 0.152939
R15141 gnd.n4220 gnd.n4219 0.152939
R15142 gnd.n4220 gnd.n3741 0.152939
R15143 gnd.n4234 gnd.n3741 0.152939
R15144 gnd.n4235 gnd.n4234 0.152939
R15145 gnd.n4236 gnd.n4235 0.152939
R15146 gnd.n4236 gnd.n3735 0.152939
R15147 gnd.n4251 gnd.n3735 0.152939
R15148 gnd.n4252 gnd.n4251 0.152939
R15149 gnd.n4253 gnd.n4252 0.152939
R15150 gnd.n4253 gnd.n3554 0.152939
R15151 gnd.n5904 gnd.n2677 0.152939
R15152 gnd.n5900 gnd.n2677 0.152939
R15153 gnd.n5900 gnd.n5899 0.152939
R15154 gnd.n5899 gnd.n5898 0.152939
R15155 gnd.n5898 gnd.n2682 0.152939
R15156 gnd.n5894 gnd.n2682 0.152939
R15157 gnd.n5894 gnd.n5893 0.152939
R15158 gnd.n5893 gnd.n5892 0.152939
R15159 gnd.n5892 gnd.n2687 0.152939
R15160 gnd.n5888 gnd.n2687 0.152939
R15161 gnd.n5888 gnd.n5887 0.152939
R15162 gnd.n5887 gnd.n5886 0.152939
R15163 gnd.n5886 gnd.n2692 0.152939
R15164 gnd.n5882 gnd.n2692 0.152939
R15165 gnd.n5882 gnd.n5881 0.152939
R15166 gnd.n5881 gnd.n5880 0.152939
R15167 gnd.n5880 gnd.n2697 0.152939
R15168 gnd.n5876 gnd.n2697 0.152939
R15169 gnd.n5876 gnd.n5875 0.152939
R15170 gnd.n5875 gnd.n5874 0.152939
R15171 gnd.n5874 gnd.n2702 0.152939
R15172 gnd.n5870 gnd.n2702 0.152939
R15173 gnd.n5870 gnd.n5869 0.152939
R15174 gnd.n5869 gnd.n5868 0.152939
R15175 gnd.n5868 gnd.n2707 0.152939
R15176 gnd.n5864 gnd.n2707 0.152939
R15177 gnd.n5864 gnd.n5863 0.152939
R15178 gnd.n5863 gnd.n5862 0.152939
R15179 gnd.n5862 gnd.n2712 0.152939
R15180 gnd.n5858 gnd.n2712 0.152939
R15181 gnd.n5858 gnd.n5857 0.152939
R15182 gnd.n5857 gnd.n5856 0.152939
R15183 gnd.n5856 gnd.n2717 0.152939
R15184 gnd.n5852 gnd.n2717 0.152939
R15185 gnd.n5852 gnd.n5851 0.152939
R15186 gnd.n5851 gnd.n5850 0.152939
R15187 gnd.n5850 gnd.n2722 0.152939
R15188 gnd.n5846 gnd.n2722 0.152939
R15189 gnd.n5846 gnd.n5845 0.152939
R15190 gnd.n5845 gnd.n5844 0.152939
R15191 gnd.n5844 gnd.n2727 0.152939
R15192 gnd.n5840 gnd.n2727 0.152939
R15193 gnd.n5840 gnd.n5839 0.152939
R15194 gnd.n5839 gnd.n5838 0.152939
R15195 gnd.n5838 gnd.n2732 0.152939
R15196 gnd.n5834 gnd.n2732 0.152939
R15197 gnd.n5834 gnd.n5833 0.152939
R15198 gnd.n5833 gnd.n5832 0.152939
R15199 gnd.n5832 gnd.n2737 0.152939
R15200 gnd.n5828 gnd.n2737 0.152939
R15201 gnd.n5828 gnd.n5827 0.152939
R15202 gnd.n5827 gnd.n5826 0.152939
R15203 gnd.n5826 gnd.n2742 0.152939
R15204 gnd.n5822 gnd.n2742 0.152939
R15205 gnd.n5822 gnd.n5821 0.152939
R15206 gnd.n5821 gnd.n5820 0.152939
R15207 gnd.n5820 gnd.n2747 0.152939
R15208 gnd.n5816 gnd.n2747 0.152939
R15209 gnd.n5816 gnd.n5815 0.152939
R15210 gnd.n5815 gnd.n5814 0.152939
R15211 gnd.n5814 gnd.n2752 0.152939
R15212 gnd.n5810 gnd.n2752 0.152939
R15213 gnd.n5810 gnd.n5809 0.152939
R15214 gnd.n5809 gnd.n5808 0.152939
R15215 gnd.n5808 gnd.n2757 0.152939
R15216 gnd.n5804 gnd.n2757 0.152939
R15217 gnd.n5804 gnd.n5803 0.152939
R15218 gnd.n5803 gnd.n5802 0.152939
R15219 gnd.n5802 gnd.n2762 0.152939
R15220 gnd.n5798 gnd.n2762 0.152939
R15221 gnd.n5798 gnd.n5797 0.152939
R15222 gnd.n5797 gnd.n5796 0.152939
R15223 gnd.n5796 gnd.n2767 0.152939
R15224 gnd.n5792 gnd.n2767 0.152939
R15225 gnd.n5792 gnd.n5791 0.152939
R15226 gnd.n5791 gnd.n5790 0.152939
R15227 gnd.n5790 gnd.n2772 0.152939
R15228 gnd.n5786 gnd.n2772 0.152939
R15229 gnd.n5786 gnd.n5785 0.152939
R15230 gnd.n5785 gnd.n5784 0.152939
R15231 gnd.n5784 gnd.n2777 0.152939
R15232 gnd.n2780 gnd.n2777 0.152939
R15233 gnd.n5691 gnd.n5690 0.152939
R15234 gnd.n5690 gnd.n5689 0.152939
R15235 gnd.n5689 gnd.n2879 0.152939
R15236 gnd.n5685 gnd.n2879 0.152939
R15237 gnd.n5685 gnd.n5684 0.152939
R15238 gnd.n5684 gnd.n5683 0.152939
R15239 gnd.n5683 gnd.n2884 0.152939
R15240 gnd.n5679 gnd.n2884 0.152939
R15241 gnd.n5679 gnd.n5678 0.152939
R15242 gnd.n5678 gnd.n5677 0.152939
R15243 gnd.n5677 gnd.n2889 0.152939
R15244 gnd.n5673 gnd.n2889 0.152939
R15245 gnd.n5673 gnd.n5672 0.152939
R15246 gnd.n5672 gnd.n5671 0.152939
R15247 gnd.n5671 gnd.n2894 0.152939
R15248 gnd.n5667 gnd.n2894 0.152939
R15249 gnd.n5667 gnd.n5666 0.152939
R15250 gnd.n5666 gnd.n5665 0.152939
R15251 gnd.n5665 gnd.n2899 0.152939
R15252 gnd.n5661 gnd.n2899 0.152939
R15253 gnd.n5661 gnd.n281 0.152939
R15254 gnd.n7197 gnd.n281 0.152939
R15255 gnd.n7197 gnd.n7196 0.152939
R15256 gnd.n7196 gnd.n7195 0.152939
R15257 gnd.n7195 gnd.n282 0.152939
R15258 gnd.n7191 gnd.n282 0.152939
R15259 gnd.n7189 gnd.n7188 0.152939
R15260 gnd.n7188 gnd.n288 0.152939
R15261 gnd.n288 gnd.n256 0.152939
R15262 gnd.n7210 gnd.n256 0.152939
R15263 gnd.n7211 gnd.n7210 0.152939
R15264 gnd.n7212 gnd.n7211 0.152939
R15265 gnd.n7212 gnd.n241 0.152939
R15266 gnd.n7226 gnd.n241 0.152939
R15267 gnd.n7227 gnd.n7226 0.152939
R15268 gnd.n7228 gnd.n7227 0.152939
R15269 gnd.n7228 gnd.n226 0.152939
R15270 gnd.n7242 gnd.n226 0.152939
R15271 gnd.n7243 gnd.n7242 0.152939
R15272 gnd.n7244 gnd.n7243 0.152939
R15273 gnd.n7244 gnd.n211 0.152939
R15274 gnd.n7258 gnd.n211 0.152939
R15275 gnd.n7259 gnd.n7258 0.152939
R15276 gnd.n7260 gnd.n7259 0.152939
R15277 gnd.n7260 gnd.n196 0.152939
R15278 gnd.n7274 gnd.n196 0.152939
R15279 gnd.n7275 gnd.n7274 0.152939
R15280 gnd.n7351 gnd.n7275 0.152939
R15281 gnd.n7351 gnd.n7350 0.152939
R15282 gnd.n7350 gnd.n7349 0.152939
R15283 gnd.n7349 gnd.n7276 0.152939
R15284 gnd.n7345 gnd.n7276 0.152939
R15285 gnd.n7344 gnd.n7278 0.152939
R15286 gnd.n7340 gnd.n7278 0.152939
R15287 gnd.n7340 gnd.n7339 0.152939
R15288 gnd.n7339 gnd.n7338 0.152939
R15289 gnd.n7338 gnd.n7284 0.152939
R15290 gnd.n7334 gnd.n7284 0.152939
R15291 gnd.n7334 gnd.n7333 0.152939
R15292 gnd.n7333 gnd.n7332 0.152939
R15293 gnd.n7332 gnd.n7292 0.152939
R15294 gnd.n7328 gnd.n7292 0.152939
R15295 gnd.n7328 gnd.n7327 0.152939
R15296 gnd.n7327 gnd.n7326 0.152939
R15297 gnd.n7326 gnd.n7300 0.152939
R15298 gnd.n7322 gnd.n7300 0.152939
R15299 gnd.n7322 gnd.n7321 0.152939
R15300 gnd.n7321 gnd.n7320 0.152939
R15301 gnd.n7320 gnd.n7308 0.152939
R15302 gnd.n7316 gnd.n7308 0.152939
R15303 gnd.n5474 gnd.n5473 0.152939
R15304 gnd.n5476 gnd.n5474 0.152939
R15305 gnd.n5476 gnd.n5475 0.152939
R15306 gnd.n5475 gnd.n3006 0.152939
R15307 gnd.n5504 gnd.n3006 0.152939
R15308 gnd.n5505 gnd.n5504 0.152939
R15309 gnd.n5507 gnd.n5505 0.152939
R15310 gnd.n5507 gnd.n5506 0.152939
R15311 gnd.n5506 gnd.n2978 0.152939
R15312 gnd.n5535 gnd.n2978 0.152939
R15313 gnd.n5536 gnd.n5535 0.152939
R15314 gnd.n5538 gnd.n5536 0.152939
R15315 gnd.n5538 gnd.n5537 0.152939
R15316 gnd.n5537 gnd.n2950 0.152939
R15317 gnd.n5574 gnd.n2950 0.152939
R15318 gnd.n5575 gnd.n5574 0.152939
R15319 gnd.n5580 gnd.n5575 0.152939
R15320 gnd.n5580 gnd.n5579 0.152939
R15321 gnd.n5579 gnd.n5578 0.152939
R15322 gnd.n5578 gnd.n2939 0.152939
R15323 gnd.n5600 gnd.n2939 0.152939
R15324 gnd.n5601 gnd.n5600 0.152939
R15325 gnd.n5605 gnd.n5601 0.152939
R15326 gnd.n5605 gnd.n5604 0.152939
R15327 gnd.n5604 gnd.n5603 0.152939
R15328 gnd.n5603 gnd.n63 0.152939
R15329 gnd.n7483 gnd.n64 0.152939
R15330 gnd.n7479 gnd.n64 0.152939
R15331 gnd.n7479 gnd.n7478 0.152939
R15332 gnd.n7478 gnd.n7477 0.152939
R15333 gnd.n7477 gnd.n70 0.152939
R15334 gnd.n7473 gnd.n70 0.152939
R15335 gnd.n7473 gnd.n7472 0.152939
R15336 gnd.n7472 gnd.n7471 0.152939
R15337 gnd.n7471 gnd.n75 0.152939
R15338 gnd.n7467 gnd.n75 0.152939
R15339 gnd.n7467 gnd.n7466 0.152939
R15340 gnd.n7466 gnd.n7465 0.152939
R15341 gnd.n7465 gnd.n80 0.152939
R15342 gnd.n7461 gnd.n80 0.152939
R15343 gnd.n7461 gnd.n7460 0.152939
R15344 gnd.n7460 gnd.n7459 0.152939
R15345 gnd.n7459 gnd.n85 0.152939
R15346 gnd.n7455 gnd.n85 0.152939
R15347 gnd.n7455 gnd.n7454 0.152939
R15348 gnd.n7454 gnd.n7453 0.152939
R15349 gnd.n7453 gnd.n90 0.152939
R15350 gnd.n7449 gnd.n90 0.152939
R15351 gnd.n7449 gnd.n7448 0.152939
R15352 gnd.n7448 gnd.n7447 0.152939
R15353 gnd.n7447 gnd.n95 0.152939
R15354 gnd.n98 gnd.n95 0.152939
R15355 gnd.n5471 gnd.n5470 0.151415
R15356 gnd.n4603 gnd.n4602 0.151415
R15357 gnd.n305 gnd.n264 0.128549
R15358 gnd.n3936 gnd.n3837 0.128549
R15359 gnd.n1861 gnd.n1860 0.0767195
R15360 gnd.n1860 gnd.n1859 0.0767195
R15361 gnd.n7204 gnd.n249 0.0767195
R15362 gnd.n5615 gnd.n287 0.0767195
R15363 gnd.n296 gnd.n287 0.0767195
R15364 gnd.n7204 gnd.n263 0.0767195
R15365 gnd.n2559 gnd.n2521 0.0767195
R15366 gnd.n4145 gnd.n2530 0.0767195
R15367 gnd.n4145 gnd.n2531 0.0767195
R15368 gnd.n4147 gnd.n4146 0.0767195
R15369 gnd.n4146 gnd.n3770 0.0767195
R15370 gnd.n2521 gnd.n2501 0.0767195
R15371 gnd.n7191 gnd.n7190 0.0767195
R15372 gnd.n7190 gnd.n7189 0.0767195
R15373 gnd.n7484 gnd.n63 0.0767195
R15374 gnd.n7484 gnd.n7483 0.0767195
R15375 gnd.n4154 gnd.n4153 0.0695946
R15376 gnd.n4155 gnd.n4154 0.0695946
R15377 gnd.n5906 gnd.n5905 0.063
R15378 gnd.n3127 gnd.n2878 0.063
R15379 gnd.n6207 gnd.n1048 0.0477147
R15380 gnd.n1624 gnd.n1512 0.0442063
R15381 gnd.n1625 gnd.n1624 0.0442063
R15382 gnd.n1626 gnd.n1625 0.0442063
R15383 gnd.n1626 gnd.n1501 0.0442063
R15384 gnd.n1640 gnd.n1501 0.0442063
R15385 gnd.n1641 gnd.n1640 0.0442063
R15386 gnd.n1642 gnd.n1641 0.0442063
R15387 gnd.n1642 gnd.n1488 0.0442063
R15388 gnd.n1686 gnd.n1488 0.0442063
R15389 gnd.n1687 gnd.n1686 0.0442063
R15390 gnd.n1689 gnd.n1422 0.0344674
R15391 gnd.n3089 gnd.n3082 0.0344674
R15392 gnd.n4601 gnd.n3555 0.0344674
R15393 gnd.n1709 gnd.n1708 0.0269946
R15394 gnd.n1711 gnd.n1710 0.0269946
R15395 gnd.n1417 gnd.n1415 0.0269946
R15396 gnd.n1721 gnd.n1719 0.0269946
R15397 gnd.n1720 gnd.n1396 0.0269946
R15398 gnd.n1740 gnd.n1739 0.0269946
R15399 gnd.n1742 gnd.n1741 0.0269946
R15400 gnd.n1391 gnd.n1390 0.0269946
R15401 gnd.n1752 gnd.n1386 0.0269946
R15402 gnd.n1751 gnd.n1388 0.0269946
R15403 gnd.n1387 gnd.n1369 0.0269946
R15404 gnd.n1772 gnd.n1370 0.0269946
R15405 gnd.n1771 gnd.n1371 0.0269946
R15406 gnd.n1805 gnd.n1346 0.0269946
R15407 gnd.n1807 gnd.n1806 0.0269946
R15408 gnd.n1808 gnd.n1293 0.0269946
R15409 gnd.n1341 gnd.n1294 0.0269946
R15410 gnd.n1343 gnd.n1295 0.0269946
R15411 gnd.n1818 gnd.n1817 0.0269946
R15412 gnd.n1820 gnd.n1819 0.0269946
R15413 gnd.n1821 gnd.n1315 0.0269946
R15414 gnd.n1823 gnd.n1316 0.0269946
R15415 gnd.n1826 gnd.n1317 0.0269946
R15416 gnd.n1829 gnd.n1828 0.0269946
R15417 gnd.n1831 gnd.n1830 0.0269946
R15418 gnd.n1896 gnd.n1216 0.0269946
R15419 gnd.n1898 gnd.n1897 0.0269946
R15420 gnd.n1907 gnd.n1209 0.0269946
R15421 gnd.n1909 gnd.n1908 0.0269946
R15422 gnd.n1910 gnd.n1207 0.0269946
R15423 gnd.n1917 gnd.n1913 0.0269946
R15424 gnd.n1916 gnd.n1915 0.0269946
R15425 gnd.n1914 gnd.n1186 0.0269946
R15426 gnd.n1941 gnd.n1187 0.0269946
R15427 gnd.n1940 gnd.n1188 0.0269946
R15428 gnd.n2014 gnd.n1162 0.0269946
R15429 gnd.n2016 gnd.n2015 0.0269946
R15430 gnd.n2017 gnd.n972 0.0269946
R15431 gnd.n1157 gnd.n973 0.0269946
R15432 gnd.n1159 gnd.n974 0.0269946
R15433 gnd.n2025 gnd.n2024 0.0269946
R15434 gnd.n2027 gnd.n2026 0.0269946
R15435 gnd.n2028 gnd.n996 0.0269946
R15436 gnd.n2030 gnd.n997 0.0269946
R15437 gnd.n2032 gnd.n998 0.0269946
R15438 gnd.n2038 gnd.n2037 0.0269946
R15439 gnd.n2040 gnd.n2039 0.0269946
R15440 gnd.n2041 gnd.n1022 0.0269946
R15441 gnd.n2301 gnd.n1024 0.0269946
R15442 gnd.n2307 gnd.n2306 0.0269946
R15443 gnd.n2309 gnd.n2308 0.0269946
R15444 gnd.n6208 gnd.n1047 0.0269946
R15445 gnd.n3936 gnd.n3842 0.0248902
R15446 gnd.n2921 gnd.n264 0.0248902
R15447 gnd.n3128 gnd.n3127 0.0246168
R15448 gnd.n5905 gnd.n2676 0.0246168
R15449 gnd.n1689 gnd.n1688 0.0202011
R15450 gnd.n3128 gnd.n3125 0.0174837
R15451 gnd.n3133 gnd.n3125 0.0174837
R15452 gnd.n3134 gnd.n3133 0.0174837
R15453 gnd.n3134 gnd.n3123 0.0174837
R15454 gnd.n3141 gnd.n3123 0.0174837
R15455 gnd.n3143 gnd.n3141 0.0174837
R15456 gnd.n3143 gnd.n3142 0.0174837
R15457 gnd.n3142 gnd.n3118 0.0174837
R15458 gnd.n3150 gnd.n3118 0.0174837
R15459 gnd.n3150 gnd.n3149 0.0174837
R15460 gnd.n3149 gnd.n3119 0.0174837
R15461 gnd.n3119 gnd.n3114 0.0174837
R15462 gnd.n3158 gnd.n3114 0.0174837
R15463 gnd.n3160 gnd.n3158 0.0174837
R15464 gnd.n3160 gnd.n3159 0.0174837
R15465 gnd.n3159 gnd.n3109 0.0174837
R15466 gnd.n3167 gnd.n3109 0.0174837
R15467 gnd.n3167 gnd.n3166 0.0174837
R15468 gnd.n3166 gnd.n3110 0.0174837
R15469 gnd.n3110 gnd.n3105 0.0174837
R15470 gnd.n3175 gnd.n3105 0.0174837
R15471 gnd.n3177 gnd.n3175 0.0174837
R15472 gnd.n3177 gnd.n3176 0.0174837
R15473 gnd.n3176 gnd.n3100 0.0174837
R15474 gnd.n3184 gnd.n3100 0.0174837
R15475 gnd.n3184 gnd.n3183 0.0174837
R15476 gnd.n3183 gnd.n3101 0.0174837
R15477 gnd.n3101 gnd.n3096 0.0174837
R15478 gnd.n3192 gnd.n3096 0.0174837
R15479 gnd.n3194 gnd.n3192 0.0174837
R15480 gnd.n3194 gnd.n3193 0.0174837
R15481 gnd.n3193 gnd.n3088 0.0174837
R15482 gnd.n3199 gnd.n3088 0.0174837
R15483 gnd.n3199 gnd.n3198 0.0174837
R15484 gnd.n3198 gnd.n3089 0.0174837
R15485 gnd.n3601 gnd.n2676 0.0174837
R15486 gnd.n3607 gnd.n3601 0.0174837
R15487 gnd.n3608 gnd.n3607 0.0174837
R15488 gnd.n3608 gnd.n3598 0.0174837
R15489 gnd.n3613 gnd.n3598 0.0174837
R15490 gnd.n3614 gnd.n3613 0.0174837
R15491 gnd.n3614 gnd.n3596 0.0174837
R15492 gnd.n3619 gnd.n3596 0.0174837
R15493 gnd.n3620 gnd.n3619 0.0174837
R15494 gnd.n3620 gnd.n3592 0.0174837
R15495 gnd.n3625 gnd.n3592 0.0174837
R15496 gnd.n3626 gnd.n3625 0.0174837
R15497 gnd.n3626 gnd.n3588 0.0174837
R15498 gnd.n3631 gnd.n3588 0.0174837
R15499 gnd.n3632 gnd.n3631 0.0174837
R15500 gnd.n3632 gnd.n3586 0.0174837
R15501 gnd.n3637 gnd.n3586 0.0174837
R15502 gnd.n3638 gnd.n3637 0.0174837
R15503 gnd.n3638 gnd.n3584 0.0174837
R15504 gnd.n3643 gnd.n3584 0.0174837
R15505 gnd.n3644 gnd.n3643 0.0174837
R15506 gnd.n3644 gnd.n3580 0.0174837
R15507 gnd.n3649 gnd.n3580 0.0174837
R15508 gnd.n3650 gnd.n3649 0.0174837
R15509 gnd.n3650 gnd.n3576 0.0174837
R15510 gnd.n3654 gnd.n3576 0.0174837
R15511 gnd.n3655 gnd.n3654 0.0174837
R15512 gnd.n3655 gnd.n3574 0.0174837
R15513 gnd.n3660 gnd.n3574 0.0174837
R15514 gnd.n3662 gnd.n3660 0.0174837
R15515 gnd.n3662 gnd.n3661 0.0174837
R15516 gnd.n3661 gnd.n3559 0.0174837
R15517 gnd.n4595 gnd.n3559 0.0174837
R15518 gnd.n4595 gnd.n4594 0.0174837
R15519 gnd.n4594 gnd.n3555 0.0174837
R15520 gnd.n1688 gnd.n1687 0.0148637
R15521 gnd.n2299 gnd.n2298 0.0144266
R15522 gnd.n2298 gnd.n1023 0.0130679
R15523 gnd.n1708 gnd.n1422 0.00797283
R15524 gnd.n1710 gnd.n1709 0.00797283
R15525 gnd.n1711 gnd.n1417 0.00797283
R15526 gnd.n1719 gnd.n1415 0.00797283
R15527 gnd.n1721 gnd.n1720 0.00797283
R15528 gnd.n1739 gnd.n1396 0.00797283
R15529 gnd.n1741 gnd.n1740 0.00797283
R15530 gnd.n1742 gnd.n1391 0.00797283
R15531 gnd.n1390 gnd.n1386 0.00797283
R15532 gnd.n1752 gnd.n1751 0.00797283
R15533 gnd.n1388 gnd.n1387 0.00797283
R15534 gnd.n1370 gnd.n1369 0.00797283
R15535 gnd.n1772 gnd.n1771 0.00797283
R15536 gnd.n1371 gnd.n1346 0.00797283
R15537 gnd.n1806 gnd.n1805 0.00797283
R15538 gnd.n1808 gnd.n1807 0.00797283
R15539 gnd.n1341 gnd.n1293 0.00797283
R15540 gnd.n1343 gnd.n1294 0.00797283
R15541 gnd.n1817 gnd.n1295 0.00797283
R15542 gnd.n1819 gnd.n1818 0.00797283
R15543 gnd.n1821 gnd.n1820 0.00797283
R15544 gnd.n1823 gnd.n1315 0.00797283
R15545 gnd.n1826 gnd.n1316 0.00797283
R15546 gnd.n1828 gnd.n1317 0.00797283
R15547 gnd.n1831 gnd.n1829 0.00797283
R15548 gnd.n1830 gnd.n1216 0.00797283
R15549 gnd.n1898 gnd.n1896 0.00797283
R15550 gnd.n1897 gnd.n1209 0.00797283
R15551 gnd.n1908 gnd.n1907 0.00797283
R15552 gnd.n1910 gnd.n1909 0.00797283
R15553 gnd.n1913 gnd.n1207 0.00797283
R15554 gnd.n1917 gnd.n1916 0.00797283
R15555 gnd.n1915 gnd.n1914 0.00797283
R15556 gnd.n1187 gnd.n1186 0.00797283
R15557 gnd.n1941 gnd.n1940 0.00797283
R15558 gnd.n1188 gnd.n1162 0.00797283
R15559 gnd.n2015 gnd.n2014 0.00797283
R15560 gnd.n2017 gnd.n2016 0.00797283
R15561 gnd.n1157 gnd.n972 0.00797283
R15562 gnd.n1159 gnd.n973 0.00797283
R15563 gnd.n2024 gnd.n974 0.00797283
R15564 gnd.n2026 gnd.n2025 0.00797283
R15565 gnd.n2028 gnd.n2027 0.00797283
R15566 gnd.n2030 gnd.n996 0.00797283
R15567 gnd.n2032 gnd.n997 0.00797283
R15568 gnd.n2037 gnd.n998 0.00797283
R15569 gnd.n2039 gnd.n2038 0.00797283
R15570 gnd.n2041 gnd.n2040 0.00797283
R15571 gnd.n2299 gnd.n1022 0.00797283
R15572 gnd.n2301 gnd.n1023 0.00797283
R15573 gnd.n2306 gnd.n1024 0.00797283
R15574 gnd.n2309 gnd.n2307 0.00797283
R15575 gnd.n2308 gnd.n1047 0.00797283
R15576 gnd.n6208 gnd.n6207 0.00797283
R15577 gnd.n7190 gnd.n287 0.00507153
R15578 gnd.n4146 gnd.n4145 0.00507153
R15579 gnd.n5471 gnd.n3082 0.000839674
R15580 gnd.n4602 gnd.n4601 0.000839674
R15581 a_n8964_8799.n228 a_n8964_8799.t140 485.149
R15582 a_n8964_8799.n247 a_n8964_8799.t154 485.149
R15583 a_n8964_8799.n267 a_n8964_8799.t96 485.149
R15584 a_n8964_8799.n167 a_n8964_8799.t91 485.149
R15585 a_n8964_8799.n186 a_n8964_8799.t101 485.149
R15586 a_n8964_8799.n206 a_n8964_8799.t94 485.149
R15587 a_n8964_8799.n56 a_n8964_8799.t111 485.135
R15588 a_n8964_8799.n240 a_n8964_8799.t47 464.166
R15589 a_n8964_8799.n222 a_n8964_8799.t117 464.166
R15590 a_n8964_8799.n239 a_n8964_8799.t115 464.166
R15591 a_n8964_8799.n238 a_n8964_8799.t53 464.166
R15592 a_n8964_8799.n223 a_n8964_8799.t51 464.166
R15593 a_n8964_8799.n237 a_n8964_8799.t137 464.166
R15594 a_n8964_8799.n236 a_n8964_8799.t69 464.166
R15595 a_n8964_8799.n224 a_n8964_8799.t55 464.166
R15596 a_n8964_8799.n235 a_n8964_8799.t143 464.166
R15597 a_n8964_8799.n234 a_n8964_8799.t95 464.166
R15598 a_n8964_8799.n225 a_n8964_8799.t70 464.166
R15599 a_n8964_8799.n233 a_n8964_8799.t161 464.166
R15600 a_n8964_8799.n232 a_n8964_8799.t113 464.166
R15601 a_n8964_8799.n226 a_n8964_8799.t72 464.166
R15602 a_n8964_8799.n231 a_n8964_8799.t155 464.166
R15603 a_n8964_8799.n230 a_n8964_8799.t116 464.166
R15604 a_n8964_8799.n227 a_n8964_8799.t89 464.166
R15605 a_n8964_8799.n229 a_n8964_8799.t52 464.166
R15606 a_n8964_8799.n71 a_n8964_8799.t127 485.135
R15607 a_n8964_8799.n259 a_n8964_8799.t59 464.166
R15608 a_n8964_8799.n241 a_n8964_8799.t135 464.166
R15609 a_n8964_8799.n258 a_n8964_8799.t133 464.166
R15610 a_n8964_8799.n257 a_n8964_8799.t62 464.166
R15611 a_n8964_8799.n242 a_n8964_8799.t61 464.166
R15612 a_n8964_8799.n256 a_n8964_8799.t153 464.166
R15613 a_n8964_8799.n255 a_n8964_8799.t78 464.166
R15614 a_n8964_8799.n243 a_n8964_8799.t68 464.166
R15615 a_n8964_8799.n254 a_n8964_8799.t156 464.166
R15616 a_n8964_8799.n253 a_n8964_8799.t108 464.166
R15617 a_n8964_8799.n244 a_n8964_8799.t81 464.166
R15618 a_n8964_8799.n252 a_n8964_8799.t54 464.166
R15619 a_n8964_8799.n251 a_n8964_8799.t128 464.166
R15620 a_n8964_8799.n245 a_n8964_8799.t82 464.166
R15621 a_n8964_8799.n250 a_n8964_8799.t46 464.166
R15622 a_n8964_8799.n249 a_n8964_8799.t134 464.166
R15623 a_n8964_8799.n246 a_n8964_8799.t97 464.166
R15624 a_n8964_8799.n248 a_n8964_8799.t63 464.166
R15625 a_n8964_8799.n86 a_n8964_8799.t73 485.135
R15626 a_n8964_8799.n279 a_n8964_8799.t159 464.166
R15627 a_n8964_8799.n261 a_n8964_8799.t126 464.166
R15628 a_n8964_8799.n278 a_n8964_8799.t152 464.166
R15629 a_n8964_8799.n277 a_n8964_8799.t107 464.166
R15630 a_n8964_8799.n262 a_n8964_8799.t132 464.166
R15631 a_n8964_8799.n276 a_n8964_8799.t67 464.166
R15632 a_n8964_8799.n275 a_n8964_8799.t149 464.166
R15633 a_n8964_8799.n263 a_n8964_8799.t85 464.166
R15634 a_n8964_8799.n274 a_n8964_8799.t144 464.166
R15635 a_n8964_8799.n273 a_n8964_8799.t71 464.166
R15636 a_n8964_8799.n264 a_n8964_8799.t120 464.166
R15637 a_n8964_8799.n272 a_n8964_8799.t58 464.166
R15638 a_n8964_8799.n271 a_n8964_8799.t104 464.166
R15639 a_n8964_8799.n265 a_n8964_8799.t80 464.166
R15640 a_n8964_8799.n270 a_n8964_8799.t130 464.166
R15641 a_n8964_8799.n269 a_n8964_8799.t65 464.166
R15642 a_n8964_8799.n266 a_n8964_8799.t112 464.166
R15643 a_n8964_8799.n268 a_n8964_8799.t50 464.166
R15644 a_n8964_8799.n168 a_n8964_8799.t121 464.166
R15645 a_n8964_8799.n169 a_n8964_8799.t48 464.166
R15646 a_n8964_8799.n170 a_n8964_8799.t76 464.166
R15647 a_n8964_8799.n171 a_n8964_8799.t114 464.166
R15648 a_n8964_8799.n166 a_n8964_8799.t151 464.166
R15649 a_n8964_8799.n172 a_n8964_8799.t74 464.166
R15650 a_n8964_8799.n173 a_n8964_8799.t109 464.166
R15651 a_n8964_8799.n174 a_n8964_8799.t146 464.166
R15652 a_n8964_8799.n175 a_n8964_8799.t147 464.166
R15653 a_n8964_8799.n165 a_n8964_8799.t93 464.166
R15654 a_n8964_8799.n176 a_n8964_8799.t125 464.166
R15655 a_n8964_8799.n164 a_n8964_8799.t145 464.166
R15656 a_n8964_8799.n177 a_n8964_8799.t90 464.166
R15657 a_n8964_8799.n178 a_n8964_8799.t92 464.166
R15658 a_n8964_8799.n179 a_n8964_8799.t122 464.166
R15659 a_n8964_8799.n180 a_n8964_8799.t75 464.166
R15660 a_n8964_8799.n163 a_n8964_8799.t77 464.166
R15661 a_n8964_8799.n181 a_n8964_8799.t118 464.166
R15662 a_n8964_8799.n187 a_n8964_8799.t138 464.166
R15663 a_n8964_8799.n188 a_n8964_8799.t60 464.166
R15664 a_n8964_8799.n189 a_n8964_8799.t87 464.166
R15665 a_n8964_8799.n190 a_n8964_8799.t129 464.166
R15666 a_n8964_8799.n185 a_n8964_8799.t163 464.166
R15667 a_n8964_8799.n191 a_n8964_8799.t83 464.166
R15668 a_n8964_8799.n192 a_n8964_8799.t123 464.166
R15669 a_n8964_8799.n193 a_n8964_8799.t160 464.166
R15670 a_n8964_8799.n194 a_n8964_8799.t162 464.166
R15671 a_n8964_8799.n184 a_n8964_8799.t105 464.166
R15672 a_n8964_8799.n195 a_n8964_8799.t142 464.166
R15673 a_n8964_8799.n183 a_n8964_8799.t158 464.166
R15674 a_n8964_8799.n196 a_n8964_8799.t100 464.166
R15675 a_n8964_8799.n197 a_n8964_8799.t102 464.166
R15676 a_n8964_8799.n198 a_n8964_8799.t139 464.166
R15677 a_n8964_8799.n199 a_n8964_8799.t86 464.166
R15678 a_n8964_8799.n182 a_n8964_8799.t88 464.166
R15679 a_n8964_8799.n200 a_n8964_8799.t136 464.166
R15680 a_n8964_8799.n207 a_n8964_8799.t49 464.166
R15681 a_n8964_8799.n208 a_n8964_8799.t110 464.166
R15682 a_n8964_8799.n209 a_n8964_8799.t64 464.166
R15683 a_n8964_8799.n210 a_n8964_8799.t131 464.166
R15684 a_n8964_8799.n205 a_n8964_8799.t79 464.166
R15685 a_n8964_8799.n211 a_n8964_8799.t103 464.166
R15686 a_n8964_8799.n212 a_n8964_8799.t57 464.166
R15687 a_n8964_8799.n213 a_n8964_8799.t119 464.166
R15688 a_n8964_8799.n214 a_n8964_8799.t98 464.166
R15689 a_n8964_8799.n204 a_n8964_8799.t141 464.166
R15690 a_n8964_8799.n215 a_n8964_8799.t84 464.166
R15691 a_n8964_8799.n203 a_n8964_8799.t148 464.166
R15692 a_n8964_8799.n216 a_n8964_8799.t66 464.166
R15693 a_n8964_8799.n217 a_n8964_8799.t45 464.166
R15694 a_n8964_8799.n218 a_n8964_8799.t106 464.166
R15695 a_n8964_8799.n219 a_n8964_8799.t150 464.166
R15696 a_n8964_8799.n202 a_n8964_8799.t124 464.166
R15697 a_n8964_8799.n220 a_n8964_8799.t157 464.166
R15698 a_n8964_8799.n41 a_n8964_8799.n70 71.7212
R15699 a_n8964_8799.n70 a_n8964_8799.n227 17.8606
R15700 a_n8964_8799.n69 a_n8964_8799.n41 76.9909
R15701 a_n8964_8799.n230 a_n8964_8799.n69 7.32118
R15702 a_n8964_8799.n68 a_n8964_8799.n40 78.3454
R15703 a_n8964_8799.n40 a_n8964_8799.n67 72.8951
R15704 a_n8964_8799.n66 a_n8964_8799.n42 70.1674
R15705 a_n8964_8799.n233 a_n8964_8799.n66 20.9683
R15706 a_n8964_8799.n42 a_n8964_8799.n65 72.3034
R15707 a_n8964_8799.n65 a_n8964_8799.n225 16.6962
R15708 a_n8964_8799.n64 a_n8964_8799.n43 77.6622
R15709 a_n8964_8799.n234 a_n8964_8799.n64 5.97853
R15710 a_n8964_8799.n63 a_n8964_8799.n43 77.6622
R15711 a_n8964_8799.n44 a_n8964_8799.n62 72.3034
R15712 a_n8964_8799.n61 a_n8964_8799.n44 70.1674
R15713 a_n8964_8799.n237 a_n8964_8799.n61 20.9683
R15714 a_n8964_8799.n46 a_n8964_8799.n60 72.8951
R15715 a_n8964_8799.n60 a_n8964_8799.n223 15.5127
R15716 a_n8964_8799.n59 a_n8964_8799.n46 78.3454
R15717 a_n8964_8799.n238 a_n8964_8799.n59 4.61226
R15718 a_n8964_8799.n58 a_n8964_8799.n45 76.9909
R15719 a_n8964_8799.n45 a_n8964_8799.n57 71.7212
R15720 a_n8964_8799.n240 a_n8964_8799.n56 20.9683
R15721 a_n8964_8799.n47 a_n8964_8799.n56 70.1674
R15722 a_n8964_8799.n33 a_n8964_8799.n85 71.7212
R15723 a_n8964_8799.n85 a_n8964_8799.n246 17.8606
R15724 a_n8964_8799.n84 a_n8964_8799.n33 76.9909
R15725 a_n8964_8799.n249 a_n8964_8799.n84 7.32118
R15726 a_n8964_8799.n83 a_n8964_8799.n32 78.3454
R15727 a_n8964_8799.n32 a_n8964_8799.n82 72.8951
R15728 a_n8964_8799.n81 a_n8964_8799.n34 70.1674
R15729 a_n8964_8799.n252 a_n8964_8799.n81 20.9683
R15730 a_n8964_8799.n34 a_n8964_8799.n80 72.3034
R15731 a_n8964_8799.n80 a_n8964_8799.n244 16.6962
R15732 a_n8964_8799.n79 a_n8964_8799.n35 77.6622
R15733 a_n8964_8799.n253 a_n8964_8799.n79 5.97853
R15734 a_n8964_8799.n78 a_n8964_8799.n35 77.6622
R15735 a_n8964_8799.n36 a_n8964_8799.n77 72.3034
R15736 a_n8964_8799.n76 a_n8964_8799.n36 70.1674
R15737 a_n8964_8799.n256 a_n8964_8799.n76 20.9683
R15738 a_n8964_8799.n38 a_n8964_8799.n75 72.8951
R15739 a_n8964_8799.n75 a_n8964_8799.n242 15.5127
R15740 a_n8964_8799.n74 a_n8964_8799.n38 78.3454
R15741 a_n8964_8799.n257 a_n8964_8799.n74 4.61226
R15742 a_n8964_8799.n73 a_n8964_8799.n37 76.9909
R15743 a_n8964_8799.n37 a_n8964_8799.n72 71.7212
R15744 a_n8964_8799.n259 a_n8964_8799.n71 20.9683
R15745 a_n8964_8799.n39 a_n8964_8799.n71 70.1674
R15746 a_n8964_8799.n25 a_n8964_8799.n100 71.7212
R15747 a_n8964_8799.n100 a_n8964_8799.n266 17.8606
R15748 a_n8964_8799.n99 a_n8964_8799.n25 76.9909
R15749 a_n8964_8799.n269 a_n8964_8799.n99 7.32118
R15750 a_n8964_8799.n98 a_n8964_8799.n24 78.3454
R15751 a_n8964_8799.n24 a_n8964_8799.n97 72.8951
R15752 a_n8964_8799.n96 a_n8964_8799.n26 70.1674
R15753 a_n8964_8799.n272 a_n8964_8799.n96 20.9683
R15754 a_n8964_8799.n26 a_n8964_8799.n95 72.3034
R15755 a_n8964_8799.n95 a_n8964_8799.n264 16.6962
R15756 a_n8964_8799.n94 a_n8964_8799.n27 77.6622
R15757 a_n8964_8799.n273 a_n8964_8799.n94 5.97853
R15758 a_n8964_8799.n93 a_n8964_8799.n27 77.6622
R15759 a_n8964_8799.n28 a_n8964_8799.n92 72.3034
R15760 a_n8964_8799.n91 a_n8964_8799.n28 70.1674
R15761 a_n8964_8799.n276 a_n8964_8799.n91 20.9683
R15762 a_n8964_8799.n30 a_n8964_8799.n90 72.8951
R15763 a_n8964_8799.n90 a_n8964_8799.n262 15.5127
R15764 a_n8964_8799.n89 a_n8964_8799.n30 78.3454
R15765 a_n8964_8799.n277 a_n8964_8799.n89 4.61226
R15766 a_n8964_8799.n88 a_n8964_8799.n29 76.9909
R15767 a_n8964_8799.n29 a_n8964_8799.n87 71.7212
R15768 a_n8964_8799.n279 a_n8964_8799.n86 20.9683
R15769 a_n8964_8799.n31 a_n8964_8799.n86 70.1674
R15770 a_n8964_8799.n17 a_n8964_8799.n115 70.1674
R15771 a_n8964_8799.n181 a_n8964_8799.n115 20.9683
R15772 a_n8964_8799.n114 a_n8964_8799.n17 71.7212
R15773 a_n8964_8799.n114 a_n8964_8799.n163 17.8606
R15774 a_n8964_8799.n16 a_n8964_8799.n113 76.9909
R15775 a_n8964_8799.n180 a_n8964_8799.n113 7.32118
R15776 a_n8964_8799.n112 a_n8964_8799.n16 78.3454
R15777 a_n8964_8799.n18 a_n8964_8799.n111 72.8951
R15778 a_n8964_8799.n110 a_n8964_8799.n18 70.1674
R15779 a_n8964_8799.n110 a_n8964_8799.n164 20.9683
R15780 a_n8964_8799.n19 a_n8964_8799.n109 72.3034
R15781 a_n8964_8799.n176 a_n8964_8799.n109 16.6962
R15782 a_n8964_8799.n108 a_n8964_8799.n19 77.6622
R15783 a_n8964_8799.n108 a_n8964_8799.n165 5.97853
R15784 a_n8964_8799.n20 a_n8964_8799.n107 77.6622
R15785 a_n8964_8799.n106 a_n8964_8799.n20 72.3034
R15786 a_n8964_8799.n21 a_n8964_8799.n105 70.1674
R15787 a_n8964_8799.n172 a_n8964_8799.n105 20.9683
R15788 a_n8964_8799.n104 a_n8964_8799.n21 72.8951
R15789 a_n8964_8799.n104 a_n8964_8799.n166 15.5127
R15790 a_n8964_8799.n22 a_n8964_8799.n103 78.3454
R15791 a_n8964_8799.n171 a_n8964_8799.n103 4.61226
R15792 a_n8964_8799.n102 a_n8964_8799.n22 76.9909
R15793 a_n8964_8799.n101 a_n8964_8799.n169 17.8606
R15794 a_n8964_8799.n101 a_n8964_8799.n23 71.7212
R15795 a_n8964_8799.n9 a_n8964_8799.n130 70.1674
R15796 a_n8964_8799.n200 a_n8964_8799.n130 20.9683
R15797 a_n8964_8799.n129 a_n8964_8799.n9 71.7212
R15798 a_n8964_8799.n129 a_n8964_8799.n182 17.8606
R15799 a_n8964_8799.n8 a_n8964_8799.n128 76.9909
R15800 a_n8964_8799.n199 a_n8964_8799.n128 7.32118
R15801 a_n8964_8799.n127 a_n8964_8799.n8 78.3454
R15802 a_n8964_8799.n10 a_n8964_8799.n126 72.8951
R15803 a_n8964_8799.n125 a_n8964_8799.n10 70.1674
R15804 a_n8964_8799.n125 a_n8964_8799.n183 20.9683
R15805 a_n8964_8799.n11 a_n8964_8799.n124 72.3034
R15806 a_n8964_8799.n195 a_n8964_8799.n124 16.6962
R15807 a_n8964_8799.n123 a_n8964_8799.n11 77.6622
R15808 a_n8964_8799.n123 a_n8964_8799.n184 5.97853
R15809 a_n8964_8799.n12 a_n8964_8799.n122 77.6622
R15810 a_n8964_8799.n121 a_n8964_8799.n12 72.3034
R15811 a_n8964_8799.n13 a_n8964_8799.n120 70.1674
R15812 a_n8964_8799.n191 a_n8964_8799.n120 20.9683
R15813 a_n8964_8799.n119 a_n8964_8799.n13 72.8951
R15814 a_n8964_8799.n119 a_n8964_8799.n185 15.5127
R15815 a_n8964_8799.n14 a_n8964_8799.n118 78.3454
R15816 a_n8964_8799.n190 a_n8964_8799.n118 4.61226
R15817 a_n8964_8799.n117 a_n8964_8799.n14 76.9909
R15818 a_n8964_8799.n116 a_n8964_8799.n188 17.8606
R15819 a_n8964_8799.n116 a_n8964_8799.n15 71.7212
R15820 a_n8964_8799.n1 a_n8964_8799.n145 70.1674
R15821 a_n8964_8799.n220 a_n8964_8799.n145 20.9683
R15822 a_n8964_8799.n144 a_n8964_8799.n1 71.7212
R15823 a_n8964_8799.n144 a_n8964_8799.n202 17.8606
R15824 a_n8964_8799.n0 a_n8964_8799.n143 76.9909
R15825 a_n8964_8799.n219 a_n8964_8799.n143 7.32118
R15826 a_n8964_8799.n142 a_n8964_8799.n0 78.3454
R15827 a_n8964_8799.n2 a_n8964_8799.n141 72.8951
R15828 a_n8964_8799.n140 a_n8964_8799.n2 70.1674
R15829 a_n8964_8799.n140 a_n8964_8799.n203 20.9683
R15830 a_n8964_8799.n3 a_n8964_8799.n139 72.3034
R15831 a_n8964_8799.n215 a_n8964_8799.n139 16.6962
R15832 a_n8964_8799.n138 a_n8964_8799.n3 77.6622
R15833 a_n8964_8799.n138 a_n8964_8799.n204 5.97853
R15834 a_n8964_8799.n4 a_n8964_8799.n137 77.6622
R15835 a_n8964_8799.n136 a_n8964_8799.n4 72.3034
R15836 a_n8964_8799.n5 a_n8964_8799.n135 70.1674
R15837 a_n8964_8799.n211 a_n8964_8799.n135 20.9683
R15838 a_n8964_8799.n134 a_n8964_8799.n5 72.8951
R15839 a_n8964_8799.n134 a_n8964_8799.n205 15.5127
R15840 a_n8964_8799.n6 a_n8964_8799.n133 78.3454
R15841 a_n8964_8799.n210 a_n8964_8799.n133 4.61226
R15842 a_n8964_8799.n132 a_n8964_8799.n6 76.9909
R15843 a_n8964_8799.n131 a_n8964_8799.n208 17.8606
R15844 a_n8964_8799.n131 a_n8964_8799.n7 71.7212
R15845 a_n8964_8799.n51 a_n8964_8799.n146 98.9633
R15846 a_n8964_8799.n54 a_n8964_8799.n287 98.9631
R15847 a_n8964_8799.n54 a_n8964_8799.n286 98.6055
R15848 a_n8964_8799.n53 a_n8964_8799.n285 98.6055
R15849 a_n8964_8799.n53 a_n8964_8799.n284 98.6055
R15850 a_n8964_8799.n52 a_n8964_8799.n150 98.6055
R15851 a_n8964_8799.n52 a_n8964_8799.n149 98.6055
R15852 a_n8964_8799.n51 a_n8964_8799.n148 98.6055
R15853 a_n8964_8799.n51 a_n8964_8799.n147 98.6055
R15854 a_n8964_8799.n288 a_n8964_8799.n54 98.6054
R15855 a_n8964_8799.n49 a_n8964_8799.n151 81.2902
R15856 a_n8964_8799.n55 a_n8964_8799.n157 81.2902
R15857 a_n8964_8799.n48 a_n8964_8799.n154 81.2902
R15858 a_n8964_8799.n50 a_n8964_8799.n160 80.9324
R15859 a_n8964_8799.n50 a_n8964_8799.n161 80.9324
R15860 a_n8964_8799.n49 a_n8964_8799.n162 80.9324
R15861 a_n8964_8799.n49 a_n8964_8799.n153 80.9324
R15862 a_n8964_8799.n49 a_n8964_8799.n152 80.9324
R15863 a_n8964_8799.n55 a_n8964_8799.n158 80.9324
R15864 a_n8964_8799.n48 a_n8964_8799.n159 80.9324
R15865 a_n8964_8799.n48 a_n8964_8799.n156 80.9324
R15866 a_n8964_8799.n48 a_n8964_8799.n155 80.9324
R15867 a_n8964_8799.n41 a_n8964_8799.n228 70.4033
R15868 a_n8964_8799.n33 a_n8964_8799.n247 70.4033
R15869 a_n8964_8799.n25 a_n8964_8799.n267 70.4033
R15870 a_n8964_8799.n167 a_n8964_8799.n23 70.4033
R15871 a_n8964_8799.n186 a_n8964_8799.n15 70.4033
R15872 a_n8964_8799.n206 a_n8964_8799.n7 70.4033
R15873 a_n8964_8799.n239 a_n8964_8799.n238 48.2005
R15874 a_n8964_8799.n61 a_n8964_8799.n236 20.9683
R15875 a_n8964_8799.n235 a_n8964_8799.n234 48.2005
R15876 a_n8964_8799.n66 a_n8964_8799.n232 20.9683
R15877 a_n8964_8799.n231 a_n8964_8799.n230 48.2005
R15878 a_n8964_8799.n258 a_n8964_8799.n257 48.2005
R15879 a_n8964_8799.n76 a_n8964_8799.n255 20.9683
R15880 a_n8964_8799.n254 a_n8964_8799.n253 48.2005
R15881 a_n8964_8799.n81 a_n8964_8799.n251 20.9683
R15882 a_n8964_8799.n250 a_n8964_8799.n249 48.2005
R15883 a_n8964_8799.n278 a_n8964_8799.n277 48.2005
R15884 a_n8964_8799.n91 a_n8964_8799.n275 20.9683
R15885 a_n8964_8799.n274 a_n8964_8799.n273 48.2005
R15886 a_n8964_8799.n96 a_n8964_8799.n271 20.9683
R15887 a_n8964_8799.n270 a_n8964_8799.n269 48.2005
R15888 a_n8964_8799.n171 a_n8964_8799.n170 48.2005
R15889 a_n8964_8799.n173 a_n8964_8799.n105 20.9683
R15890 a_n8964_8799.n175 a_n8964_8799.n165 48.2005
R15891 a_n8964_8799.n177 a_n8964_8799.n110 20.9683
R15892 a_n8964_8799.n180 a_n8964_8799.n179 48.2005
R15893 a_n8964_8799.t44 a_n8964_8799.n115 485.135
R15894 a_n8964_8799.n190 a_n8964_8799.n189 48.2005
R15895 a_n8964_8799.n192 a_n8964_8799.n120 20.9683
R15896 a_n8964_8799.n194 a_n8964_8799.n184 48.2005
R15897 a_n8964_8799.n196 a_n8964_8799.n125 20.9683
R15898 a_n8964_8799.n199 a_n8964_8799.n198 48.2005
R15899 a_n8964_8799.t56 a_n8964_8799.n130 485.135
R15900 a_n8964_8799.n210 a_n8964_8799.n209 48.2005
R15901 a_n8964_8799.n212 a_n8964_8799.n135 20.9683
R15902 a_n8964_8799.n214 a_n8964_8799.n204 48.2005
R15903 a_n8964_8799.n216 a_n8964_8799.n140 20.9683
R15904 a_n8964_8799.n219 a_n8964_8799.n218 48.2005
R15905 a_n8964_8799.t99 a_n8964_8799.n145 485.135
R15906 a_n8964_8799.n57 a_n8964_8799.n222 17.8606
R15907 a_n8964_8799.n229 a_n8964_8799.n70 25.894
R15908 a_n8964_8799.n72 a_n8964_8799.n241 17.8606
R15909 a_n8964_8799.n248 a_n8964_8799.n85 25.894
R15910 a_n8964_8799.n87 a_n8964_8799.n261 17.8606
R15911 a_n8964_8799.n268 a_n8964_8799.n100 25.894
R15912 a_n8964_8799.n181 a_n8964_8799.n114 25.894
R15913 a_n8964_8799.n200 a_n8964_8799.n129 25.894
R15914 a_n8964_8799.n220 a_n8964_8799.n144 25.894
R15915 a_n8964_8799.n68 a_n8964_8799.n226 43.3183
R15916 a_n8964_8799.n83 a_n8964_8799.n245 43.3183
R15917 a_n8964_8799.n98 a_n8964_8799.n265 43.3183
R15918 a_n8964_8799.n178 a_n8964_8799.n112 43.3183
R15919 a_n8964_8799.n197 a_n8964_8799.n127 43.3183
R15920 a_n8964_8799.n217 a_n8964_8799.n142 43.3183
R15921 a_n8964_8799.n62 a_n8964_8799.n224 16.6962
R15922 a_n8964_8799.n233 a_n8964_8799.n65 27.6507
R15923 a_n8964_8799.n77 a_n8964_8799.n243 16.6962
R15924 a_n8964_8799.n252 a_n8964_8799.n80 27.6507
R15925 a_n8964_8799.n92 a_n8964_8799.n263 16.6962
R15926 a_n8964_8799.n272 a_n8964_8799.n95 27.6507
R15927 a_n8964_8799.n174 a_n8964_8799.n106 16.6962
R15928 a_n8964_8799.n164 a_n8964_8799.n109 27.6507
R15929 a_n8964_8799.n193 a_n8964_8799.n121 16.6962
R15930 a_n8964_8799.n183 a_n8964_8799.n124 27.6507
R15931 a_n8964_8799.n213 a_n8964_8799.n136 16.6962
R15932 a_n8964_8799.n203 a_n8964_8799.n139 27.6507
R15933 a_n8964_8799.n63 a_n8964_8799.n224 41.7634
R15934 a_n8964_8799.n78 a_n8964_8799.n243 41.7634
R15935 a_n8964_8799.n93 a_n8964_8799.n263 41.7634
R15936 a_n8964_8799.n107 a_n8964_8799.n174 41.7634
R15937 a_n8964_8799.n122 a_n8964_8799.n193 41.7634
R15938 a_n8964_8799.n137 a_n8964_8799.n213 41.7634
R15939 a_n8964_8799.n237 a_n8964_8799.n60 29.3885
R15940 a_n8964_8799.n67 a_n8964_8799.n226 15.5127
R15941 a_n8964_8799.n256 a_n8964_8799.n75 29.3885
R15942 a_n8964_8799.n82 a_n8964_8799.n245 15.5127
R15943 a_n8964_8799.n276 a_n8964_8799.n90 29.3885
R15944 a_n8964_8799.n97 a_n8964_8799.n265 15.5127
R15945 a_n8964_8799.n172 a_n8964_8799.n104 29.3885
R15946 a_n8964_8799.n178 a_n8964_8799.n111 15.5127
R15947 a_n8964_8799.n191 a_n8964_8799.n119 29.3885
R15948 a_n8964_8799.n197 a_n8964_8799.n126 15.5127
R15949 a_n8964_8799.n211 a_n8964_8799.n134 29.3885
R15950 a_n8964_8799.n217 a_n8964_8799.n141 15.5127
R15951 a_n8964_8799.n58 a_n8964_8799.n222 40.1848
R15952 a_n8964_8799.n73 a_n8964_8799.n241 40.1848
R15953 a_n8964_8799.n88 a_n8964_8799.n261 40.1848
R15954 a_n8964_8799.n169 a_n8964_8799.n102 40.1848
R15955 a_n8964_8799.n188 a_n8964_8799.n117 40.1848
R15956 a_n8964_8799.n208 a_n8964_8799.n132 40.1848
R15957 a_n8964_8799.n53 a_n8964_8799.n283 32.8234
R15958 a_n8964_8799.n50 a_n8964_8799.n48 32.5134
R15959 a_n8964_8799.n229 a_n8964_8799.n228 20.9576
R15960 a_n8964_8799.n248 a_n8964_8799.n247 20.9576
R15961 a_n8964_8799.n268 a_n8964_8799.n267 20.9576
R15962 a_n8964_8799.n168 a_n8964_8799.n167 20.9576
R15963 a_n8964_8799.n187 a_n8964_8799.n186 20.9576
R15964 a_n8964_8799.n207 a_n8964_8799.n206 20.9576
R15965 a_n8964_8799.n283 a_n8964_8799.n52 19.9193
R15966 a_n8964_8799.n58 a_n8964_8799.n239 7.32118
R15967 a_n8964_8799.n69 a_n8964_8799.n227 40.1848
R15968 a_n8964_8799.n73 a_n8964_8799.n258 7.32118
R15969 a_n8964_8799.n84 a_n8964_8799.n246 40.1848
R15970 a_n8964_8799.n88 a_n8964_8799.n278 7.32118
R15971 a_n8964_8799.n99 a_n8964_8799.n266 40.1848
R15972 a_n8964_8799.n170 a_n8964_8799.n102 7.32118
R15973 a_n8964_8799.n163 a_n8964_8799.n113 40.1848
R15974 a_n8964_8799.n189 a_n8964_8799.n117 7.32118
R15975 a_n8964_8799.n182 a_n8964_8799.n128 40.1848
R15976 a_n8964_8799.n209 a_n8964_8799.n132 7.32118
R15977 a_n8964_8799.n202 a_n8964_8799.n143 40.1848
R15978 a_n8964_8799.n232 a_n8964_8799.n67 29.3885
R15979 a_n8964_8799.n251 a_n8964_8799.n82 29.3885
R15980 a_n8964_8799.n271 a_n8964_8799.n97 29.3885
R15981 a_n8964_8799.n111 a_n8964_8799.n177 29.3885
R15982 a_n8964_8799.n126 a_n8964_8799.n196 29.3885
R15983 a_n8964_8799.n141 a_n8964_8799.n216 29.3885
R15984 a_n8964_8799.n63 a_n8964_8799.n235 5.97853
R15985 a_n8964_8799.n64 a_n8964_8799.n225 41.7634
R15986 a_n8964_8799.n78 a_n8964_8799.n254 5.97853
R15987 a_n8964_8799.n79 a_n8964_8799.n244 41.7634
R15988 a_n8964_8799.n93 a_n8964_8799.n274 5.97853
R15989 a_n8964_8799.n94 a_n8964_8799.n264 41.7634
R15990 a_n8964_8799.n175 a_n8964_8799.n107 5.97853
R15991 a_n8964_8799.n176 a_n8964_8799.n108 41.7634
R15992 a_n8964_8799.n194 a_n8964_8799.n122 5.97853
R15993 a_n8964_8799.n195 a_n8964_8799.n123 41.7634
R15994 a_n8964_8799.n214 a_n8964_8799.n137 5.97853
R15995 a_n8964_8799.n215 a_n8964_8799.n138 41.7634
R15996 a_n8964_8799.n282 a_n8964_8799.n49 12.3339
R15997 a_n8964_8799.n283 a_n8964_8799.n282 11.4887
R15998 a_n8964_8799.n236 a_n8964_8799.n62 27.6507
R15999 a_n8964_8799.n255 a_n8964_8799.n77 27.6507
R16000 a_n8964_8799.n275 a_n8964_8799.n92 27.6507
R16001 a_n8964_8799.n173 a_n8964_8799.n106 27.6507
R16002 a_n8964_8799.n192 a_n8964_8799.n121 27.6507
R16003 a_n8964_8799.n212 a_n8964_8799.n136 27.6507
R16004 a_n8964_8799.n59 a_n8964_8799.n223 43.3183
R16005 a_n8964_8799.n68 a_n8964_8799.n231 4.61226
R16006 a_n8964_8799.n74 a_n8964_8799.n242 43.3183
R16007 a_n8964_8799.n83 a_n8964_8799.n250 4.61226
R16008 a_n8964_8799.n89 a_n8964_8799.n262 43.3183
R16009 a_n8964_8799.n98 a_n8964_8799.n270 4.61226
R16010 a_n8964_8799.n166 a_n8964_8799.n103 43.3183
R16011 a_n8964_8799.n179 a_n8964_8799.n112 4.61226
R16012 a_n8964_8799.n185 a_n8964_8799.n118 43.3183
R16013 a_n8964_8799.n198 a_n8964_8799.n127 4.61226
R16014 a_n8964_8799.n205 a_n8964_8799.n133 43.3183
R16015 a_n8964_8799.n218 a_n8964_8799.n142 4.61226
R16016 a_n8964_8799.n260 a_n8964_8799.n47 9.04406
R16017 a_n8964_8799.n201 a_n8964_8799.n17 9.04406
R16018 a_n8964_8799.n240 a_n8964_8799.n57 25.894
R16019 a_n8964_8799.n259 a_n8964_8799.n72 25.894
R16020 a_n8964_8799.n279 a_n8964_8799.n87 25.894
R16021 a_n8964_8799.n101 a_n8964_8799.n168 25.894
R16022 a_n8964_8799.n116 a_n8964_8799.n187 25.894
R16023 a_n8964_8799.n131 a_n8964_8799.n207 25.894
R16024 a_n8964_8799.n281 a_n8964_8799.n221 7.07257
R16025 a_n8964_8799.n281 a_n8964_8799.n280 6.72634
R16026 a_n8964_8799.n260 a_n8964_8799.n39 4.93611
R16027 a_n8964_8799.n280 a_n8964_8799.n31 4.93611
R16028 a_n8964_8799.n201 a_n8964_8799.n9 4.93611
R16029 a_n8964_8799.n221 a_n8964_8799.n1 4.93611
R16030 a_n8964_8799.n280 a_n8964_8799.n260 4.10845
R16031 a_n8964_8799.n221 a_n8964_8799.n201 4.10845
R16032 a_n8964_8799.n287 a_n8964_8799.t27 3.61217
R16033 a_n8964_8799.n287 a_n8964_8799.t37 3.61217
R16034 a_n8964_8799.n286 a_n8964_8799.t34 3.61217
R16035 a_n8964_8799.n286 a_n8964_8799.t35 3.61217
R16036 a_n8964_8799.n285 a_n8964_8799.t23 3.61217
R16037 a_n8964_8799.n285 a_n8964_8799.t40 3.61217
R16038 a_n8964_8799.n284 a_n8964_8799.t20 3.61217
R16039 a_n8964_8799.n284 a_n8964_8799.t42 3.61217
R16040 a_n8964_8799.n150 a_n8964_8799.t25 3.61217
R16041 a_n8964_8799.n150 a_n8964_8799.t41 3.61217
R16042 a_n8964_8799.n149 a_n8964_8799.t26 3.61217
R16043 a_n8964_8799.n149 a_n8964_8799.t36 3.61217
R16044 a_n8964_8799.n148 a_n8964_8799.t28 3.61217
R16045 a_n8964_8799.n148 a_n8964_8799.t24 3.61217
R16046 a_n8964_8799.n147 a_n8964_8799.t29 3.61217
R16047 a_n8964_8799.n147 a_n8964_8799.t21 3.61217
R16048 a_n8964_8799.n146 a_n8964_8799.t8 3.61217
R16049 a_n8964_8799.n146 a_n8964_8799.t7 3.61217
R16050 a_n8964_8799.n288 a_n8964_8799.t17 3.61217
R16051 a_n8964_8799.t6 a_n8964_8799.n288 3.61217
R16052 a_n8964_8799.n282 a_n8964_8799.n281 3.4105
R16053 a_n8964_8799.n160 a_n8964_8799.t43 2.82907
R16054 a_n8964_8799.n160 a_n8964_8799.t39 2.82907
R16055 a_n8964_8799.n161 a_n8964_8799.t33 2.82907
R16056 a_n8964_8799.n161 a_n8964_8799.t13 2.82907
R16057 a_n8964_8799.n162 a_n8964_8799.t4 2.82907
R16058 a_n8964_8799.n162 a_n8964_8799.t22 2.82907
R16059 a_n8964_8799.n153 a_n8964_8799.t12 2.82907
R16060 a_n8964_8799.n153 a_n8964_8799.t38 2.82907
R16061 a_n8964_8799.n152 a_n8964_8799.t15 2.82907
R16062 a_n8964_8799.n152 a_n8964_8799.t0 2.82907
R16063 a_n8964_8799.n151 a_n8964_8799.t14 2.82907
R16064 a_n8964_8799.n151 a_n8964_8799.t30 2.82907
R16065 a_n8964_8799.n157 a_n8964_8799.t32 2.82907
R16066 a_n8964_8799.n157 a_n8964_8799.t11 2.82907
R16067 a_n8964_8799.n158 a_n8964_8799.t19 2.82907
R16068 a_n8964_8799.n158 a_n8964_8799.t1 2.82907
R16069 a_n8964_8799.n159 a_n8964_8799.t16 2.82907
R16070 a_n8964_8799.n159 a_n8964_8799.t10 2.82907
R16071 a_n8964_8799.n156 a_n8964_8799.t18 2.82907
R16072 a_n8964_8799.n156 a_n8964_8799.t5 2.82907
R16073 a_n8964_8799.n155 a_n8964_8799.t9 2.82907
R16074 a_n8964_8799.n155 a_n8964_8799.t3 2.82907
R16075 a_n8964_8799.n154 a_n8964_8799.t2 2.82907
R16076 a_n8964_8799.n154 a_n8964_8799.t31 2.82907
R16077 a_n8964_8799.n49 a_n8964_8799.n50 1.43153
R16078 a_n8964_8799.n41 a_n8964_8799.n40 1.13686
R16079 a_n8964_8799.n33 a_n8964_8799.n32 1.13686
R16080 a_n8964_8799.n25 a_n8964_8799.n24 1.13686
R16081 a_n8964_8799.n17 a_n8964_8799.n16 1.13686
R16082 a_n8964_8799.n9 a_n8964_8799.n8 1.13686
R16083 a_n8964_8799.n1 a_n8964_8799.n0 1.13686
R16084 a_n8964_8799.n54 a_n8964_8799.n53 1.07378
R16085 a_n8964_8799.n52 a_n8964_8799.n51 1.07378
R16086 a_n8964_8799.n48 a_n8964_8799.n55 1.07378
R16087 a_n8964_8799.n46 a_n8964_8799.n45 0.758076
R16088 a_n8964_8799.n46 a_n8964_8799.n44 0.758076
R16089 a_n8964_8799.n44 a_n8964_8799.n43 0.758076
R16090 a_n8964_8799.n43 a_n8964_8799.n42 0.758076
R16091 a_n8964_8799.n40 a_n8964_8799.n42 0.758076
R16092 a_n8964_8799.n38 a_n8964_8799.n37 0.758076
R16093 a_n8964_8799.n38 a_n8964_8799.n36 0.758076
R16094 a_n8964_8799.n36 a_n8964_8799.n35 0.758076
R16095 a_n8964_8799.n35 a_n8964_8799.n34 0.758076
R16096 a_n8964_8799.n32 a_n8964_8799.n34 0.758076
R16097 a_n8964_8799.n30 a_n8964_8799.n29 0.758076
R16098 a_n8964_8799.n30 a_n8964_8799.n28 0.758076
R16099 a_n8964_8799.n28 a_n8964_8799.n27 0.758076
R16100 a_n8964_8799.n27 a_n8964_8799.n26 0.758076
R16101 a_n8964_8799.n24 a_n8964_8799.n26 0.758076
R16102 a_n8964_8799.n21 a_n8964_8799.n22 0.758076
R16103 a_n8964_8799.n20 a_n8964_8799.n21 0.758076
R16104 a_n8964_8799.n19 a_n8964_8799.n20 0.758076
R16105 a_n8964_8799.n18 a_n8964_8799.n19 0.758076
R16106 a_n8964_8799.n16 a_n8964_8799.n18 0.758076
R16107 a_n8964_8799.n13 a_n8964_8799.n14 0.758076
R16108 a_n8964_8799.n12 a_n8964_8799.n13 0.758076
R16109 a_n8964_8799.n11 a_n8964_8799.n12 0.758076
R16110 a_n8964_8799.n10 a_n8964_8799.n11 0.758076
R16111 a_n8964_8799.n8 a_n8964_8799.n10 0.758076
R16112 a_n8964_8799.n5 a_n8964_8799.n6 0.758076
R16113 a_n8964_8799.n4 a_n8964_8799.n5 0.758076
R16114 a_n8964_8799.n3 a_n8964_8799.n4 0.758076
R16115 a_n8964_8799.n2 a_n8964_8799.n3 0.758076
R16116 a_n8964_8799.n0 a_n8964_8799.n2 0.758076
R16117 a_n8964_8799.n6 a_n8964_8799.n7 0.568682
R16118 a_n8964_8799.n14 a_n8964_8799.n15 0.568682
R16119 a_n8964_8799.n22 a_n8964_8799.n23 0.568682
R16120 a_n8964_8799.n29 a_n8964_8799.n31 0.568682
R16121 a_n8964_8799.n37 a_n8964_8799.n39 0.568682
R16122 a_n8964_8799.n45 a_n8964_8799.n47 0.568682
R16123 vdd.n327 vdd.n291 756.745
R16124 vdd.n268 vdd.n232 756.745
R16125 vdd.n225 vdd.n189 756.745
R16126 vdd.n166 vdd.n130 756.745
R16127 vdd.n124 vdd.n88 756.745
R16128 vdd.n65 vdd.n29 756.745
R16129 vdd.n1826 vdd.n1790 756.745
R16130 vdd.n1885 vdd.n1849 756.745
R16131 vdd.n1724 vdd.n1688 756.745
R16132 vdd.n1783 vdd.n1747 756.745
R16133 vdd.n1623 vdd.n1587 756.745
R16134 vdd.n1682 vdd.n1646 756.745
R16135 vdd.n1136 vdd.t65 640.208
R16136 vdd.n997 vdd.t103 640.208
R16137 vdd.n1130 vdd.t130 640.208
R16138 vdd.n988 vdd.t127 640.208
R16139 vdd.n885 vdd.t76 640.208
R16140 vdd.n2761 vdd.t121 640.208
R16141 vdd.n832 vdd.t90 640.208
R16142 vdd.n2830 vdd.t107 640.208
R16143 vdd.n799 vdd.t61 640.208
R16144 vdd.n1058 vdd.t117 640.208
R16145 vdd.n1397 vdd.t99 592.009
R16146 vdd.n1435 vdd.t111 592.009
R16147 vdd.n1331 vdd.t124 592.009
R16148 vdd.n2200 vdd.t83 592.009
R16149 vdd.n2050 vdd.t93 592.009
R16150 vdd.n2010 vdd.t114 592.009
R16151 vdd.n426 vdd.t96 592.009
R16152 vdd.n440 vdd.t69 592.009
R16153 vdd.n452 vdd.t87 592.009
R16154 vdd.n768 vdd.t57 592.009
R16155 vdd.n3366 vdd.t73 592.009
R16156 vdd.n688 vdd.t80 592.009
R16157 vdd.n328 vdd.n327 585
R16158 vdd.n326 vdd.n293 585
R16159 vdd.n325 vdd.n324 585
R16160 vdd.n296 vdd.n294 585
R16161 vdd.n319 vdd.n318 585
R16162 vdd.n317 vdd.n316 585
R16163 vdd.n300 vdd.n299 585
R16164 vdd.n311 vdd.n310 585
R16165 vdd.n309 vdd.n308 585
R16166 vdd.n304 vdd.n303 585
R16167 vdd.n269 vdd.n268 585
R16168 vdd.n267 vdd.n234 585
R16169 vdd.n266 vdd.n265 585
R16170 vdd.n237 vdd.n235 585
R16171 vdd.n260 vdd.n259 585
R16172 vdd.n258 vdd.n257 585
R16173 vdd.n241 vdd.n240 585
R16174 vdd.n252 vdd.n251 585
R16175 vdd.n250 vdd.n249 585
R16176 vdd.n245 vdd.n244 585
R16177 vdd.n226 vdd.n225 585
R16178 vdd.n224 vdd.n191 585
R16179 vdd.n223 vdd.n222 585
R16180 vdd.n194 vdd.n192 585
R16181 vdd.n217 vdd.n216 585
R16182 vdd.n215 vdd.n214 585
R16183 vdd.n198 vdd.n197 585
R16184 vdd.n209 vdd.n208 585
R16185 vdd.n207 vdd.n206 585
R16186 vdd.n202 vdd.n201 585
R16187 vdd.n167 vdd.n166 585
R16188 vdd.n165 vdd.n132 585
R16189 vdd.n164 vdd.n163 585
R16190 vdd.n135 vdd.n133 585
R16191 vdd.n158 vdd.n157 585
R16192 vdd.n156 vdd.n155 585
R16193 vdd.n139 vdd.n138 585
R16194 vdd.n150 vdd.n149 585
R16195 vdd.n148 vdd.n147 585
R16196 vdd.n143 vdd.n142 585
R16197 vdd.n125 vdd.n124 585
R16198 vdd.n123 vdd.n90 585
R16199 vdd.n122 vdd.n121 585
R16200 vdd.n93 vdd.n91 585
R16201 vdd.n116 vdd.n115 585
R16202 vdd.n114 vdd.n113 585
R16203 vdd.n97 vdd.n96 585
R16204 vdd.n108 vdd.n107 585
R16205 vdd.n106 vdd.n105 585
R16206 vdd.n101 vdd.n100 585
R16207 vdd.n66 vdd.n65 585
R16208 vdd.n64 vdd.n31 585
R16209 vdd.n63 vdd.n62 585
R16210 vdd.n34 vdd.n32 585
R16211 vdd.n57 vdd.n56 585
R16212 vdd.n55 vdd.n54 585
R16213 vdd.n38 vdd.n37 585
R16214 vdd.n49 vdd.n48 585
R16215 vdd.n47 vdd.n46 585
R16216 vdd.n42 vdd.n41 585
R16217 vdd.n1827 vdd.n1826 585
R16218 vdd.n1825 vdd.n1792 585
R16219 vdd.n1824 vdd.n1823 585
R16220 vdd.n1795 vdd.n1793 585
R16221 vdd.n1818 vdd.n1817 585
R16222 vdd.n1816 vdd.n1815 585
R16223 vdd.n1799 vdd.n1798 585
R16224 vdd.n1810 vdd.n1809 585
R16225 vdd.n1808 vdd.n1807 585
R16226 vdd.n1803 vdd.n1802 585
R16227 vdd.n1886 vdd.n1885 585
R16228 vdd.n1884 vdd.n1851 585
R16229 vdd.n1883 vdd.n1882 585
R16230 vdd.n1854 vdd.n1852 585
R16231 vdd.n1877 vdd.n1876 585
R16232 vdd.n1875 vdd.n1874 585
R16233 vdd.n1858 vdd.n1857 585
R16234 vdd.n1869 vdd.n1868 585
R16235 vdd.n1867 vdd.n1866 585
R16236 vdd.n1862 vdd.n1861 585
R16237 vdd.n1725 vdd.n1724 585
R16238 vdd.n1723 vdd.n1690 585
R16239 vdd.n1722 vdd.n1721 585
R16240 vdd.n1693 vdd.n1691 585
R16241 vdd.n1716 vdd.n1715 585
R16242 vdd.n1714 vdd.n1713 585
R16243 vdd.n1697 vdd.n1696 585
R16244 vdd.n1708 vdd.n1707 585
R16245 vdd.n1706 vdd.n1705 585
R16246 vdd.n1701 vdd.n1700 585
R16247 vdd.n1784 vdd.n1783 585
R16248 vdd.n1782 vdd.n1749 585
R16249 vdd.n1781 vdd.n1780 585
R16250 vdd.n1752 vdd.n1750 585
R16251 vdd.n1775 vdd.n1774 585
R16252 vdd.n1773 vdd.n1772 585
R16253 vdd.n1756 vdd.n1755 585
R16254 vdd.n1767 vdd.n1766 585
R16255 vdd.n1765 vdd.n1764 585
R16256 vdd.n1760 vdd.n1759 585
R16257 vdd.n1624 vdd.n1623 585
R16258 vdd.n1622 vdd.n1589 585
R16259 vdd.n1621 vdd.n1620 585
R16260 vdd.n1592 vdd.n1590 585
R16261 vdd.n1615 vdd.n1614 585
R16262 vdd.n1613 vdd.n1612 585
R16263 vdd.n1596 vdd.n1595 585
R16264 vdd.n1607 vdd.n1606 585
R16265 vdd.n1605 vdd.n1604 585
R16266 vdd.n1600 vdd.n1599 585
R16267 vdd.n1683 vdd.n1682 585
R16268 vdd.n1681 vdd.n1648 585
R16269 vdd.n1680 vdd.n1679 585
R16270 vdd.n1651 vdd.n1649 585
R16271 vdd.n1674 vdd.n1673 585
R16272 vdd.n1672 vdd.n1671 585
R16273 vdd.n1655 vdd.n1654 585
R16274 vdd.n1666 vdd.n1665 585
R16275 vdd.n1664 vdd.n1663 585
R16276 vdd.n1659 vdd.n1658 585
R16277 vdd.n3538 vdd.n392 509.269
R16278 vdd.n3534 vdd.n393 509.269
R16279 vdd.n3406 vdd.n685 509.269
R16280 vdd.n3403 vdd.n684 509.269
R16281 vdd.n2195 vdd.n1155 509.269
R16282 vdd.n2198 vdd.n2197 509.269
R16283 vdd.n1304 vdd.n1268 509.269
R16284 vdd.n1500 vdd.n1269 509.269
R16285 vdd.n305 vdd.t172 329.043
R16286 vdd.n246 vdd.t213 329.043
R16287 vdd.n203 vdd.t152 329.043
R16288 vdd.n144 vdd.t193 329.043
R16289 vdd.n102 vdd.t236 329.043
R16290 vdd.n43 vdd.t262 329.043
R16291 vdd.n1804 vdd.t292 329.043
R16292 vdd.n1863 vdd.t241 329.043
R16293 vdd.n1702 vdd.t280 329.043
R16294 vdd.n1761 vdd.t229 329.043
R16295 vdd.n1601 vdd.t233 329.043
R16296 vdd.n1660 vdd.t238 329.043
R16297 vdd.n1397 vdd.t102 319.788
R16298 vdd.n1435 vdd.t113 319.788
R16299 vdd.n1331 vdd.t126 319.788
R16300 vdd.n2200 vdd.t85 319.788
R16301 vdd.n2050 vdd.t94 319.788
R16302 vdd.n2010 vdd.t115 319.788
R16303 vdd.n426 vdd.t97 319.788
R16304 vdd.n440 vdd.t71 319.788
R16305 vdd.n452 vdd.t88 319.788
R16306 vdd.n768 vdd.t60 319.788
R16307 vdd.n3366 vdd.t75 319.788
R16308 vdd.n688 vdd.t82 319.788
R16309 vdd.n1398 vdd.t101 303.69
R16310 vdd.n1436 vdd.t112 303.69
R16311 vdd.n1332 vdd.t125 303.69
R16312 vdd.n2201 vdd.t86 303.69
R16313 vdd.n2051 vdd.t95 303.69
R16314 vdd.n2011 vdd.t116 303.69
R16315 vdd.n427 vdd.t98 303.69
R16316 vdd.n441 vdd.t72 303.69
R16317 vdd.n453 vdd.t89 303.69
R16318 vdd.n769 vdd.t59 303.69
R16319 vdd.n3367 vdd.t74 303.69
R16320 vdd.n689 vdd.t81 303.69
R16321 vdd.n3016 vdd.n947 285.366
R16322 vdd.n3240 vdd.n809 285.366
R16323 vdd.n3177 vdd.n806 285.366
R16324 vdd.n2895 vdd.n944 285.366
R16325 vdd.n2725 vdd.n985 285.366
R16326 vdd.n2656 vdd.n2655 285.366
R16327 vdd.n2396 vdd.n1111 285.366
R16328 vdd.n2466 vdd.n1113 285.366
R16329 vdd.n3156 vdd.n807 285.366
R16330 vdd.n3243 vdd.n3242 285.366
R16331 vdd.n3009 vdd.n945 285.366
R16332 vdd.n3018 vdd.n943 285.366
R16333 vdd.n2653 vdd.n995 285.366
R16334 vdd.n993 vdd.n967 285.366
R16335 vdd.n2282 vdd.n1112 285.366
R16336 vdd.n2468 vdd.n1109 285.366
R16337 vdd.n1153 vdd.n1110 216.982
R16338 vdd.n3405 vdd.n692 216.982
R16339 vdd.n3158 vdd.n807 185
R16340 vdd.n3241 vdd.n807 185
R16341 vdd.n3160 vdd.n3159 185
R16342 vdd.n3159 vdd.n805 185
R16343 vdd.n3161 vdd.n839 185
R16344 vdd.n3171 vdd.n839 185
R16345 vdd.n3162 vdd.n848 185
R16346 vdd.n848 vdd.n846 185
R16347 vdd.n3164 vdd.n3163 185
R16348 vdd.n3165 vdd.n3164 185
R16349 vdd.n3117 vdd.n847 185
R16350 vdd.n847 vdd.n843 185
R16351 vdd.n3116 vdd.n3115 185
R16352 vdd.n3115 vdd.n3114 185
R16353 vdd.n850 vdd.n849 185
R16354 vdd.n851 vdd.n850 185
R16355 vdd.n3107 vdd.n3106 185
R16356 vdd.n3108 vdd.n3107 185
R16357 vdd.n3105 vdd.n859 185
R16358 vdd.n864 vdd.n859 185
R16359 vdd.n3104 vdd.n3103 185
R16360 vdd.n3103 vdd.n3102 185
R16361 vdd.n861 vdd.n860 185
R16362 vdd.n870 vdd.n861 185
R16363 vdd.n3095 vdd.n3094 185
R16364 vdd.n3096 vdd.n3095 185
R16365 vdd.n3093 vdd.n871 185
R16366 vdd.n877 vdd.n871 185
R16367 vdd.n3092 vdd.n3091 185
R16368 vdd.n3091 vdd.n3090 185
R16369 vdd.n873 vdd.n872 185
R16370 vdd.n874 vdd.n873 185
R16371 vdd.n3083 vdd.n3082 185
R16372 vdd.n3084 vdd.n3083 185
R16373 vdd.n3081 vdd.n884 185
R16374 vdd.n884 vdd.n881 185
R16375 vdd.n3079 vdd.n3078 185
R16376 vdd.n3078 vdd.n3077 185
R16377 vdd.n887 vdd.n886 185
R16378 vdd.n888 vdd.n887 185
R16379 vdd.n3070 vdd.n3069 185
R16380 vdd.n3071 vdd.n3070 185
R16381 vdd.n3068 vdd.n896 185
R16382 vdd.n901 vdd.n896 185
R16383 vdd.n3067 vdd.n3066 185
R16384 vdd.n3066 vdd.n3065 185
R16385 vdd.n898 vdd.n897 185
R16386 vdd.n2977 vdd.n898 185
R16387 vdd.n3058 vdd.n3057 185
R16388 vdd.n3059 vdd.n3058 185
R16389 vdd.n3056 vdd.n908 185
R16390 vdd.n908 vdd.n905 185
R16391 vdd.n3055 vdd.n3054 185
R16392 vdd.n3054 vdd.n3053 185
R16393 vdd.n910 vdd.n909 185
R16394 vdd.n911 vdd.n910 185
R16395 vdd.n3046 vdd.n3045 185
R16396 vdd.n3047 vdd.n3046 185
R16397 vdd.n3044 vdd.n919 185
R16398 vdd.n2989 vdd.n919 185
R16399 vdd.n3043 vdd.n3042 185
R16400 vdd.n3042 vdd.n3041 185
R16401 vdd.n921 vdd.n920 185
R16402 vdd.n930 vdd.n921 185
R16403 vdd.n3034 vdd.n3033 185
R16404 vdd.n3035 vdd.n3034 185
R16405 vdd.n3032 vdd.n931 185
R16406 vdd.n931 vdd.n927 185
R16407 vdd.n3031 vdd.n3030 185
R16408 vdd.n3030 vdd.n3029 185
R16409 vdd.n933 vdd.n932 185
R16410 vdd.n3001 vdd.n933 185
R16411 vdd.n3022 vdd.n3021 185
R16412 vdd.n3023 vdd.n3022 185
R16413 vdd.n3020 vdd.n941 185
R16414 vdd.n946 vdd.n941 185
R16415 vdd.n3019 vdd.n3018 185
R16416 vdd.n3018 vdd.n3017 185
R16417 vdd.n943 vdd.n942 185
R16418 vdd.n2765 vdd.n2764 185
R16419 vdd.n2767 vdd.n2766 185
R16420 vdd.n2769 vdd.n2768 185
R16421 vdd.n2771 vdd.n2770 185
R16422 vdd.n2773 vdd.n2772 185
R16423 vdd.n2775 vdd.n2774 185
R16424 vdd.n2777 vdd.n2776 185
R16425 vdd.n2779 vdd.n2778 185
R16426 vdd.n2781 vdd.n2780 185
R16427 vdd.n2783 vdd.n2782 185
R16428 vdd.n2785 vdd.n2784 185
R16429 vdd.n2787 vdd.n2786 185
R16430 vdd.n2789 vdd.n2788 185
R16431 vdd.n2791 vdd.n2790 185
R16432 vdd.n2793 vdd.n2792 185
R16433 vdd.n2795 vdd.n2794 185
R16434 vdd.n2797 vdd.n2796 185
R16435 vdd.n2799 vdd.n2798 185
R16436 vdd.n2801 vdd.n2800 185
R16437 vdd.n2803 vdd.n2802 185
R16438 vdd.n2805 vdd.n2804 185
R16439 vdd.n2807 vdd.n2806 185
R16440 vdd.n2809 vdd.n2808 185
R16441 vdd.n2811 vdd.n2810 185
R16442 vdd.n2813 vdd.n2812 185
R16443 vdd.n2815 vdd.n2814 185
R16444 vdd.n2817 vdd.n2816 185
R16445 vdd.n2819 vdd.n2818 185
R16446 vdd.n2821 vdd.n2820 185
R16447 vdd.n2823 vdd.n2822 185
R16448 vdd.n2825 vdd.n2824 185
R16449 vdd.n2827 vdd.n2826 185
R16450 vdd.n2828 vdd.n2760 185
R16451 vdd.n3009 vdd.n3008 185
R16452 vdd.n3010 vdd.n3009 185
R16453 vdd.n3244 vdd.n3243 185
R16454 vdd.n3245 vdd.n798 185
R16455 vdd.n3247 vdd.n3246 185
R16456 vdd.n3249 vdd.n796 185
R16457 vdd.n3251 vdd.n3250 185
R16458 vdd.n3252 vdd.n795 185
R16459 vdd.n3254 vdd.n3253 185
R16460 vdd.n3256 vdd.n793 185
R16461 vdd.n3258 vdd.n3257 185
R16462 vdd.n3259 vdd.n792 185
R16463 vdd.n3261 vdd.n3260 185
R16464 vdd.n3263 vdd.n790 185
R16465 vdd.n3265 vdd.n3264 185
R16466 vdd.n3266 vdd.n789 185
R16467 vdd.n3268 vdd.n3267 185
R16468 vdd.n3270 vdd.n788 185
R16469 vdd.n3271 vdd.n786 185
R16470 vdd.n3274 vdd.n3273 185
R16471 vdd.n787 vdd.n785 185
R16472 vdd.n3130 vdd.n3129 185
R16473 vdd.n3132 vdd.n3131 185
R16474 vdd.n3134 vdd.n3126 185
R16475 vdd.n3136 vdd.n3135 185
R16476 vdd.n3137 vdd.n3125 185
R16477 vdd.n3139 vdd.n3138 185
R16478 vdd.n3141 vdd.n3123 185
R16479 vdd.n3143 vdd.n3142 185
R16480 vdd.n3144 vdd.n3122 185
R16481 vdd.n3146 vdd.n3145 185
R16482 vdd.n3148 vdd.n3120 185
R16483 vdd.n3150 vdd.n3149 185
R16484 vdd.n3151 vdd.n3119 185
R16485 vdd.n3153 vdd.n3152 185
R16486 vdd.n3155 vdd.n3118 185
R16487 vdd.n3157 vdd.n3156 185
R16488 vdd.n3156 vdd.n692 185
R16489 vdd.n3242 vdd.n802 185
R16490 vdd.n3242 vdd.n3241 185
R16491 vdd.n2908 vdd.n804 185
R16492 vdd.n805 vdd.n804 185
R16493 vdd.n2909 vdd.n838 185
R16494 vdd.n3171 vdd.n838 185
R16495 vdd.n2911 vdd.n2910 185
R16496 vdd.n2910 vdd.n846 185
R16497 vdd.n2912 vdd.n845 185
R16498 vdd.n3165 vdd.n845 185
R16499 vdd.n2914 vdd.n2913 185
R16500 vdd.n2913 vdd.n843 185
R16501 vdd.n2915 vdd.n853 185
R16502 vdd.n3114 vdd.n853 185
R16503 vdd.n2917 vdd.n2916 185
R16504 vdd.n2916 vdd.n851 185
R16505 vdd.n2918 vdd.n858 185
R16506 vdd.n3108 vdd.n858 185
R16507 vdd.n2920 vdd.n2919 185
R16508 vdd.n2919 vdd.n864 185
R16509 vdd.n2921 vdd.n863 185
R16510 vdd.n3102 vdd.n863 185
R16511 vdd.n2923 vdd.n2922 185
R16512 vdd.n2922 vdd.n870 185
R16513 vdd.n2924 vdd.n869 185
R16514 vdd.n3096 vdd.n869 185
R16515 vdd.n2926 vdd.n2925 185
R16516 vdd.n2925 vdd.n877 185
R16517 vdd.n2927 vdd.n876 185
R16518 vdd.n3090 vdd.n876 185
R16519 vdd.n2929 vdd.n2928 185
R16520 vdd.n2928 vdd.n874 185
R16521 vdd.n2930 vdd.n883 185
R16522 vdd.n3084 vdd.n883 185
R16523 vdd.n2932 vdd.n2931 185
R16524 vdd.n2931 vdd.n881 185
R16525 vdd.n2933 vdd.n890 185
R16526 vdd.n3077 vdd.n890 185
R16527 vdd.n2935 vdd.n2934 185
R16528 vdd.n2934 vdd.n888 185
R16529 vdd.n2936 vdd.n895 185
R16530 vdd.n3071 vdd.n895 185
R16531 vdd.n2938 vdd.n2937 185
R16532 vdd.n2937 vdd.n901 185
R16533 vdd.n2939 vdd.n900 185
R16534 vdd.n3065 vdd.n900 185
R16535 vdd.n2979 vdd.n2978 185
R16536 vdd.n2978 vdd.n2977 185
R16537 vdd.n2980 vdd.n907 185
R16538 vdd.n3059 vdd.n907 185
R16539 vdd.n2982 vdd.n2981 185
R16540 vdd.n2981 vdd.n905 185
R16541 vdd.n2983 vdd.n913 185
R16542 vdd.n3053 vdd.n913 185
R16543 vdd.n2985 vdd.n2984 185
R16544 vdd.n2984 vdd.n911 185
R16545 vdd.n2986 vdd.n918 185
R16546 vdd.n3047 vdd.n918 185
R16547 vdd.n2988 vdd.n2987 185
R16548 vdd.n2989 vdd.n2988 185
R16549 vdd.n2907 vdd.n923 185
R16550 vdd.n3041 vdd.n923 185
R16551 vdd.n2906 vdd.n2905 185
R16552 vdd.n2905 vdd.n930 185
R16553 vdd.n2904 vdd.n929 185
R16554 vdd.n3035 vdd.n929 185
R16555 vdd.n2903 vdd.n2902 185
R16556 vdd.n2902 vdd.n927 185
R16557 vdd.n2829 vdd.n935 185
R16558 vdd.n3029 vdd.n935 185
R16559 vdd.n3003 vdd.n3002 185
R16560 vdd.n3002 vdd.n3001 185
R16561 vdd.n3004 vdd.n940 185
R16562 vdd.n3023 vdd.n940 185
R16563 vdd.n3006 vdd.n3005 185
R16564 vdd.n3005 vdd.n946 185
R16565 vdd.n3007 vdd.n945 185
R16566 vdd.n3017 vdd.n945 185
R16567 vdd.n2195 vdd.n2194 185
R16568 vdd.n2196 vdd.n2195 185
R16569 vdd.n1156 vdd.n1154 185
R16570 vdd.n1974 vdd.n1154 185
R16571 vdd.n1977 vdd.n1976 185
R16572 vdd.n1976 vdd.n1975 185
R16573 vdd.n1159 vdd.n1158 185
R16574 vdd.n1160 vdd.n1159 185
R16575 vdd.n1963 vdd.n1962 185
R16576 vdd.n1964 vdd.n1963 185
R16577 vdd.n1168 vdd.n1167 185
R16578 vdd.n1955 vdd.n1167 185
R16579 vdd.n1958 vdd.n1957 185
R16580 vdd.n1957 vdd.n1956 185
R16581 vdd.n1171 vdd.n1170 185
R16582 vdd.n1178 vdd.n1171 185
R16583 vdd.n1946 vdd.n1945 185
R16584 vdd.n1947 vdd.n1946 185
R16585 vdd.n1180 vdd.n1179 185
R16586 vdd.n1179 vdd.n1177 185
R16587 vdd.n1941 vdd.n1940 185
R16588 vdd.n1940 vdd.n1939 185
R16589 vdd.n1183 vdd.n1182 185
R16590 vdd.n1184 vdd.n1183 185
R16591 vdd.n1930 vdd.n1929 185
R16592 vdd.n1931 vdd.n1930 185
R16593 vdd.n1191 vdd.n1190 185
R16594 vdd.n1922 vdd.n1190 185
R16595 vdd.n1925 vdd.n1924 185
R16596 vdd.n1924 vdd.n1923 185
R16597 vdd.n1194 vdd.n1193 185
R16598 vdd.n1200 vdd.n1194 185
R16599 vdd.n1913 vdd.n1912 185
R16600 vdd.n1914 vdd.n1913 185
R16601 vdd.n1202 vdd.n1201 185
R16602 vdd.n1905 vdd.n1201 185
R16603 vdd.n1908 vdd.n1907 185
R16604 vdd.n1907 vdd.n1906 185
R16605 vdd.n1205 vdd.n1204 185
R16606 vdd.n1206 vdd.n1205 185
R16607 vdd.n1896 vdd.n1895 185
R16608 vdd.n1897 vdd.n1896 185
R16609 vdd.n1214 vdd.n1213 185
R16610 vdd.n1213 vdd.n1212 185
R16611 vdd.n1584 vdd.n1583 185
R16612 vdd.n1583 vdd.n1582 185
R16613 vdd.n1217 vdd.n1216 185
R16614 vdd.n1223 vdd.n1217 185
R16615 vdd.n1573 vdd.n1572 185
R16616 vdd.n1574 vdd.n1573 185
R16617 vdd.n1225 vdd.n1224 185
R16618 vdd.n1565 vdd.n1224 185
R16619 vdd.n1568 vdd.n1567 185
R16620 vdd.n1567 vdd.n1566 185
R16621 vdd.n1228 vdd.n1227 185
R16622 vdd.n1235 vdd.n1228 185
R16623 vdd.n1556 vdd.n1555 185
R16624 vdd.n1557 vdd.n1556 185
R16625 vdd.n1237 vdd.n1236 185
R16626 vdd.n1236 vdd.n1234 185
R16627 vdd.n1551 vdd.n1550 185
R16628 vdd.n1550 vdd.n1549 185
R16629 vdd.n1240 vdd.n1239 185
R16630 vdd.n1241 vdd.n1240 185
R16631 vdd.n1540 vdd.n1539 185
R16632 vdd.n1541 vdd.n1540 185
R16633 vdd.n1248 vdd.n1247 185
R16634 vdd.n1532 vdd.n1247 185
R16635 vdd.n1535 vdd.n1534 185
R16636 vdd.n1534 vdd.n1533 185
R16637 vdd.n1251 vdd.n1250 185
R16638 vdd.n1257 vdd.n1251 185
R16639 vdd.n1523 vdd.n1522 185
R16640 vdd.n1524 vdd.n1523 185
R16641 vdd.n1259 vdd.n1258 185
R16642 vdd.n1515 vdd.n1258 185
R16643 vdd.n1518 vdd.n1517 185
R16644 vdd.n1517 vdd.n1516 185
R16645 vdd.n1262 vdd.n1261 185
R16646 vdd.n1263 vdd.n1262 185
R16647 vdd.n1506 vdd.n1505 185
R16648 vdd.n1507 vdd.n1506 185
R16649 vdd.n1270 vdd.n1269 185
R16650 vdd.n1305 vdd.n1269 185
R16651 vdd.n1501 vdd.n1500 185
R16652 vdd.n1273 vdd.n1272 185
R16653 vdd.n1497 vdd.n1496 185
R16654 vdd.n1498 vdd.n1497 185
R16655 vdd.n1307 vdd.n1306 185
R16656 vdd.n1492 vdd.n1309 185
R16657 vdd.n1491 vdd.n1310 185
R16658 vdd.n1490 vdd.n1311 185
R16659 vdd.n1313 vdd.n1312 185
R16660 vdd.n1486 vdd.n1315 185
R16661 vdd.n1485 vdd.n1316 185
R16662 vdd.n1484 vdd.n1317 185
R16663 vdd.n1319 vdd.n1318 185
R16664 vdd.n1480 vdd.n1321 185
R16665 vdd.n1479 vdd.n1322 185
R16666 vdd.n1478 vdd.n1323 185
R16667 vdd.n1325 vdd.n1324 185
R16668 vdd.n1474 vdd.n1327 185
R16669 vdd.n1473 vdd.n1328 185
R16670 vdd.n1472 vdd.n1329 185
R16671 vdd.n1333 vdd.n1330 185
R16672 vdd.n1468 vdd.n1335 185
R16673 vdd.n1467 vdd.n1336 185
R16674 vdd.n1466 vdd.n1337 185
R16675 vdd.n1339 vdd.n1338 185
R16676 vdd.n1462 vdd.n1341 185
R16677 vdd.n1461 vdd.n1342 185
R16678 vdd.n1460 vdd.n1343 185
R16679 vdd.n1345 vdd.n1344 185
R16680 vdd.n1456 vdd.n1347 185
R16681 vdd.n1455 vdd.n1348 185
R16682 vdd.n1454 vdd.n1349 185
R16683 vdd.n1351 vdd.n1350 185
R16684 vdd.n1450 vdd.n1353 185
R16685 vdd.n1449 vdd.n1354 185
R16686 vdd.n1448 vdd.n1355 185
R16687 vdd.n1357 vdd.n1356 185
R16688 vdd.n1444 vdd.n1359 185
R16689 vdd.n1443 vdd.n1360 185
R16690 vdd.n1442 vdd.n1361 185
R16691 vdd.n1363 vdd.n1362 185
R16692 vdd.n1438 vdd.n1365 185
R16693 vdd.n1437 vdd.n1434 185
R16694 vdd.n1433 vdd.n1366 185
R16695 vdd.n1368 vdd.n1367 185
R16696 vdd.n1429 vdd.n1370 185
R16697 vdd.n1428 vdd.n1371 185
R16698 vdd.n1427 vdd.n1372 185
R16699 vdd.n1374 vdd.n1373 185
R16700 vdd.n1423 vdd.n1376 185
R16701 vdd.n1422 vdd.n1377 185
R16702 vdd.n1421 vdd.n1378 185
R16703 vdd.n1380 vdd.n1379 185
R16704 vdd.n1417 vdd.n1382 185
R16705 vdd.n1416 vdd.n1383 185
R16706 vdd.n1415 vdd.n1384 185
R16707 vdd.n1386 vdd.n1385 185
R16708 vdd.n1411 vdd.n1388 185
R16709 vdd.n1410 vdd.n1389 185
R16710 vdd.n1409 vdd.n1390 185
R16711 vdd.n1392 vdd.n1391 185
R16712 vdd.n1405 vdd.n1394 185
R16713 vdd.n1404 vdd.n1395 185
R16714 vdd.n1403 vdd.n1396 185
R16715 vdd.n1400 vdd.n1304 185
R16716 vdd.n1498 vdd.n1304 185
R16717 vdd.n2199 vdd.n2198 185
R16718 vdd.n2203 vdd.n1149 185
R16719 vdd.n2079 vdd.n1148 185
R16720 vdd.n2082 vdd.n2081 185
R16721 vdd.n2084 vdd.n2083 185
R16722 vdd.n2087 vdd.n2086 185
R16723 vdd.n2089 vdd.n2088 185
R16724 vdd.n2091 vdd.n2077 185
R16725 vdd.n2093 vdd.n2092 185
R16726 vdd.n2094 vdd.n2071 185
R16727 vdd.n2096 vdd.n2095 185
R16728 vdd.n2098 vdd.n2069 185
R16729 vdd.n2100 vdd.n2099 185
R16730 vdd.n2101 vdd.n2064 185
R16731 vdd.n2103 vdd.n2102 185
R16732 vdd.n2105 vdd.n2062 185
R16733 vdd.n2107 vdd.n2106 185
R16734 vdd.n2108 vdd.n2058 185
R16735 vdd.n2110 vdd.n2109 185
R16736 vdd.n2112 vdd.n2055 185
R16737 vdd.n2114 vdd.n2113 185
R16738 vdd.n2056 vdd.n2049 185
R16739 vdd.n2118 vdd.n2053 185
R16740 vdd.n2119 vdd.n2045 185
R16741 vdd.n2121 vdd.n2120 185
R16742 vdd.n2123 vdd.n2043 185
R16743 vdd.n2125 vdd.n2124 185
R16744 vdd.n2126 vdd.n2038 185
R16745 vdd.n2128 vdd.n2127 185
R16746 vdd.n2130 vdd.n2036 185
R16747 vdd.n2132 vdd.n2131 185
R16748 vdd.n2133 vdd.n2031 185
R16749 vdd.n2135 vdd.n2134 185
R16750 vdd.n2137 vdd.n2029 185
R16751 vdd.n2139 vdd.n2138 185
R16752 vdd.n2140 vdd.n2024 185
R16753 vdd.n2142 vdd.n2141 185
R16754 vdd.n2144 vdd.n2022 185
R16755 vdd.n2146 vdd.n2145 185
R16756 vdd.n2147 vdd.n2018 185
R16757 vdd.n2149 vdd.n2148 185
R16758 vdd.n2151 vdd.n2015 185
R16759 vdd.n2153 vdd.n2152 185
R16760 vdd.n2016 vdd.n2009 185
R16761 vdd.n2157 vdd.n2013 185
R16762 vdd.n2158 vdd.n2005 185
R16763 vdd.n2160 vdd.n2159 185
R16764 vdd.n2162 vdd.n2003 185
R16765 vdd.n2164 vdd.n2163 185
R16766 vdd.n2165 vdd.n1998 185
R16767 vdd.n2167 vdd.n2166 185
R16768 vdd.n2169 vdd.n1996 185
R16769 vdd.n2171 vdd.n2170 185
R16770 vdd.n2172 vdd.n1991 185
R16771 vdd.n2174 vdd.n2173 185
R16772 vdd.n2176 vdd.n1990 185
R16773 vdd.n2177 vdd.n1987 185
R16774 vdd.n2180 vdd.n2179 185
R16775 vdd.n1989 vdd.n1985 185
R16776 vdd.n2184 vdd.n1983 185
R16777 vdd.n2186 vdd.n2185 185
R16778 vdd.n2188 vdd.n1981 185
R16779 vdd.n2190 vdd.n2189 185
R16780 vdd.n2191 vdd.n1155 185
R16781 vdd.n2197 vdd.n1152 185
R16782 vdd.n2197 vdd.n2196 185
R16783 vdd.n1163 vdd.n1151 185
R16784 vdd.n1974 vdd.n1151 185
R16785 vdd.n1973 vdd.n1972 185
R16786 vdd.n1975 vdd.n1973 185
R16787 vdd.n1162 vdd.n1161 185
R16788 vdd.n1161 vdd.n1160 185
R16789 vdd.n1966 vdd.n1965 185
R16790 vdd.n1965 vdd.n1964 185
R16791 vdd.n1166 vdd.n1165 185
R16792 vdd.n1955 vdd.n1166 185
R16793 vdd.n1954 vdd.n1953 185
R16794 vdd.n1956 vdd.n1954 185
R16795 vdd.n1173 vdd.n1172 185
R16796 vdd.n1178 vdd.n1172 185
R16797 vdd.n1949 vdd.n1948 185
R16798 vdd.n1948 vdd.n1947 185
R16799 vdd.n1176 vdd.n1175 185
R16800 vdd.n1177 vdd.n1176 185
R16801 vdd.n1938 vdd.n1937 185
R16802 vdd.n1939 vdd.n1938 185
R16803 vdd.n1186 vdd.n1185 185
R16804 vdd.n1185 vdd.n1184 185
R16805 vdd.n1933 vdd.n1932 185
R16806 vdd.n1932 vdd.n1931 185
R16807 vdd.n1189 vdd.n1188 185
R16808 vdd.n1922 vdd.n1189 185
R16809 vdd.n1921 vdd.n1920 185
R16810 vdd.n1923 vdd.n1921 185
R16811 vdd.n1196 vdd.n1195 185
R16812 vdd.n1200 vdd.n1195 185
R16813 vdd.n1916 vdd.n1915 185
R16814 vdd.n1915 vdd.n1914 185
R16815 vdd.n1199 vdd.n1198 185
R16816 vdd.n1905 vdd.n1199 185
R16817 vdd.n1904 vdd.n1903 185
R16818 vdd.n1906 vdd.n1904 185
R16819 vdd.n1208 vdd.n1207 185
R16820 vdd.n1207 vdd.n1206 185
R16821 vdd.n1899 vdd.n1898 185
R16822 vdd.n1898 vdd.n1897 185
R16823 vdd.n1211 vdd.n1210 185
R16824 vdd.n1212 vdd.n1211 185
R16825 vdd.n1581 vdd.n1580 185
R16826 vdd.n1582 vdd.n1581 185
R16827 vdd.n1219 vdd.n1218 185
R16828 vdd.n1223 vdd.n1218 185
R16829 vdd.n1576 vdd.n1575 185
R16830 vdd.n1575 vdd.n1574 185
R16831 vdd.n1222 vdd.n1221 185
R16832 vdd.n1565 vdd.n1222 185
R16833 vdd.n1564 vdd.n1563 185
R16834 vdd.n1566 vdd.n1564 185
R16835 vdd.n1230 vdd.n1229 185
R16836 vdd.n1235 vdd.n1229 185
R16837 vdd.n1559 vdd.n1558 185
R16838 vdd.n1558 vdd.n1557 185
R16839 vdd.n1233 vdd.n1232 185
R16840 vdd.n1234 vdd.n1233 185
R16841 vdd.n1548 vdd.n1547 185
R16842 vdd.n1549 vdd.n1548 185
R16843 vdd.n1243 vdd.n1242 185
R16844 vdd.n1242 vdd.n1241 185
R16845 vdd.n1543 vdd.n1542 185
R16846 vdd.n1542 vdd.n1541 185
R16847 vdd.n1246 vdd.n1245 185
R16848 vdd.n1532 vdd.n1246 185
R16849 vdd.n1531 vdd.n1530 185
R16850 vdd.n1533 vdd.n1531 185
R16851 vdd.n1253 vdd.n1252 185
R16852 vdd.n1257 vdd.n1252 185
R16853 vdd.n1526 vdd.n1525 185
R16854 vdd.n1525 vdd.n1524 185
R16855 vdd.n1256 vdd.n1255 185
R16856 vdd.n1515 vdd.n1256 185
R16857 vdd.n1514 vdd.n1513 185
R16858 vdd.n1516 vdd.n1514 185
R16859 vdd.n1265 vdd.n1264 185
R16860 vdd.n1264 vdd.n1263 185
R16861 vdd.n1509 vdd.n1508 185
R16862 vdd.n1508 vdd.n1507 185
R16863 vdd.n1268 vdd.n1267 185
R16864 vdd.n1305 vdd.n1268 185
R16865 vdd.n987 vdd.n985 185
R16866 vdd.n2654 vdd.n985 185
R16867 vdd.n2576 vdd.n1005 185
R16868 vdd.n1005 vdd.n992 185
R16869 vdd.n2578 vdd.n2577 185
R16870 vdd.n2579 vdd.n2578 185
R16871 vdd.n2575 vdd.n1004 185
R16872 vdd.n2334 vdd.n1004 185
R16873 vdd.n2574 vdd.n2573 185
R16874 vdd.n2573 vdd.n2572 185
R16875 vdd.n1007 vdd.n1006 185
R16876 vdd.n1008 vdd.n1007 185
R16877 vdd.n2563 vdd.n2562 185
R16878 vdd.n2564 vdd.n2563 185
R16879 vdd.n2561 vdd.n1018 185
R16880 vdd.n1018 vdd.n1015 185
R16881 vdd.n2560 vdd.n2559 185
R16882 vdd.n2559 vdd.n2558 185
R16883 vdd.n1020 vdd.n1019 185
R16884 vdd.n2346 vdd.n1020 185
R16885 vdd.n2551 vdd.n2550 185
R16886 vdd.n2552 vdd.n2551 185
R16887 vdd.n2549 vdd.n1028 185
R16888 vdd.n1033 vdd.n1028 185
R16889 vdd.n2548 vdd.n2547 185
R16890 vdd.n2547 vdd.n2546 185
R16891 vdd.n1030 vdd.n1029 185
R16892 vdd.n1039 vdd.n1030 185
R16893 vdd.n2539 vdd.n2538 185
R16894 vdd.n2540 vdd.n2539 185
R16895 vdd.n2537 vdd.n1040 185
R16896 vdd.n2358 vdd.n1040 185
R16897 vdd.n2536 vdd.n2535 185
R16898 vdd.n2535 vdd.n2534 185
R16899 vdd.n1042 vdd.n1041 185
R16900 vdd.n1043 vdd.n1042 185
R16901 vdd.n2527 vdd.n2526 185
R16902 vdd.n2528 vdd.n2527 185
R16903 vdd.n2525 vdd.n1052 185
R16904 vdd.n1052 vdd.n1049 185
R16905 vdd.n2524 vdd.n2523 185
R16906 vdd.n2523 vdd.n2522 185
R16907 vdd.n1054 vdd.n1053 185
R16908 vdd.n1063 vdd.n1054 185
R16909 vdd.n2514 vdd.n2513 185
R16910 vdd.n2515 vdd.n2514 185
R16911 vdd.n2512 vdd.n1064 185
R16912 vdd.n1070 vdd.n1064 185
R16913 vdd.n2511 vdd.n2510 185
R16914 vdd.n2510 vdd.n2509 185
R16915 vdd.n1066 vdd.n1065 185
R16916 vdd.n1067 vdd.n1066 185
R16917 vdd.n2502 vdd.n2501 185
R16918 vdd.n2503 vdd.n2502 185
R16919 vdd.n2500 vdd.n1077 185
R16920 vdd.n1077 vdd.n1074 185
R16921 vdd.n2499 vdd.n2498 185
R16922 vdd.n2498 vdd.n2497 185
R16923 vdd.n1079 vdd.n1078 185
R16924 vdd.n1080 vdd.n1079 185
R16925 vdd.n2490 vdd.n2489 185
R16926 vdd.n2491 vdd.n2490 185
R16927 vdd.n2488 vdd.n1089 185
R16928 vdd.n1089 vdd.n1086 185
R16929 vdd.n2487 vdd.n2486 185
R16930 vdd.n2486 vdd.n2485 185
R16931 vdd.n1091 vdd.n1090 185
R16932 vdd.n1092 vdd.n1091 185
R16933 vdd.n2478 vdd.n2477 185
R16934 vdd.n2479 vdd.n2478 185
R16935 vdd.n2476 vdd.n1101 185
R16936 vdd.n1101 vdd.n1098 185
R16937 vdd.n2475 vdd.n2474 185
R16938 vdd.n2474 vdd.n2473 185
R16939 vdd.n1103 vdd.n1102 185
R16940 vdd.n1104 vdd.n1103 185
R16941 vdd.n2466 vdd.n2465 185
R16942 vdd.n2467 vdd.n2466 185
R16943 vdd.n2464 vdd.n1113 185
R16944 vdd.n2463 vdd.n2462 185
R16945 vdd.n2460 vdd.n1114 185
R16946 vdd.n2460 vdd.n1110 185
R16947 vdd.n2459 vdd.n2458 185
R16948 vdd.n2457 vdd.n2456 185
R16949 vdd.n2455 vdd.n1116 185
R16950 vdd.n2453 vdd.n2452 185
R16951 vdd.n2451 vdd.n1117 185
R16952 vdd.n2450 vdd.n2449 185
R16953 vdd.n2447 vdd.n1118 185
R16954 vdd.n2445 vdd.n2444 185
R16955 vdd.n2443 vdd.n1119 185
R16956 vdd.n2442 vdd.n2441 185
R16957 vdd.n2439 vdd.n1120 185
R16958 vdd.n2437 vdd.n2436 185
R16959 vdd.n2435 vdd.n1121 185
R16960 vdd.n2434 vdd.n2433 185
R16961 vdd.n2431 vdd.n1122 185
R16962 vdd.n2429 vdd.n2428 185
R16963 vdd.n2427 vdd.n1123 185
R16964 vdd.n2426 vdd.n2425 185
R16965 vdd.n2423 vdd.n1124 185
R16966 vdd.n2421 vdd.n2420 185
R16967 vdd.n2419 vdd.n1125 185
R16968 vdd.n2418 vdd.n2417 185
R16969 vdd.n2415 vdd.n1126 185
R16970 vdd.n2413 vdd.n2412 185
R16971 vdd.n2411 vdd.n1127 185
R16972 vdd.n2410 vdd.n2409 185
R16973 vdd.n2407 vdd.n1128 185
R16974 vdd.n2405 vdd.n2404 185
R16975 vdd.n2403 vdd.n1129 185
R16976 vdd.n2401 vdd.n2400 185
R16977 vdd.n2398 vdd.n1132 185
R16978 vdd.n2396 vdd.n2395 185
R16979 vdd.n2657 vdd.n2656 185
R16980 vdd.n2659 vdd.n2658 185
R16981 vdd.n2661 vdd.n2660 185
R16982 vdd.n2664 vdd.n2663 185
R16983 vdd.n2666 vdd.n2665 185
R16984 vdd.n2668 vdd.n2667 185
R16985 vdd.n2670 vdd.n2669 185
R16986 vdd.n2672 vdd.n2671 185
R16987 vdd.n2674 vdd.n2673 185
R16988 vdd.n2676 vdd.n2675 185
R16989 vdd.n2678 vdd.n2677 185
R16990 vdd.n2680 vdd.n2679 185
R16991 vdd.n2682 vdd.n2681 185
R16992 vdd.n2684 vdd.n2683 185
R16993 vdd.n2686 vdd.n2685 185
R16994 vdd.n2688 vdd.n2687 185
R16995 vdd.n2690 vdd.n2689 185
R16996 vdd.n2692 vdd.n2691 185
R16997 vdd.n2694 vdd.n2693 185
R16998 vdd.n2696 vdd.n2695 185
R16999 vdd.n2698 vdd.n2697 185
R17000 vdd.n2700 vdd.n2699 185
R17001 vdd.n2702 vdd.n2701 185
R17002 vdd.n2704 vdd.n2703 185
R17003 vdd.n2706 vdd.n2705 185
R17004 vdd.n2708 vdd.n2707 185
R17005 vdd.n2710 vdd.n2709 185
R17006 vdd.n2712 vdd.n2711 185
R17007 vdd.n2714 vdd.n2713 185
R17008 vdd.n2716 vdd.n2715 185
R17009 vdd.n2718 vdd.n2717 185
R17010 vdd.n2720 vdd.n2719 185
R17011 vdd.n2722 vdd.n2721 185
R17012 vdd.n2723 vdd.n986 185
R17013 vdd.n2725 vdd.n2724 185
R17014 vdd.n2726 vdd.n2725 185
R17015 vdd.n2655 vdd.n990 185
R17016 vdd.n2655 vdd.n2654 185
R17017 vdd.n2332 vdd.n991 185
R17018 vdd.n992 vdd.n991 185
R17019 vdd.n2333 vdd.n1002 185
R17020 vdd.n2579 vdd.n1002 185
R17021 vdd.n2336 vdd.n2335 185
R17022 vdd.n2335 vdd.n2334 185
R17023 vdd.n2337 vdd.n1009 185
R17024 vdd.n2572 vdd.n1009 185
R17025 vdd.n2339 vdd.n2338 185
R17026 vdd.n2338 vdd.n1008 185
R17027 vdd.n2340 vdd.n1016 185
R17028 vdd.n2564 vdd.n1016 185
R17029 vdd.n2342 vdd.n2341 185
R17030 vdd.n2341 vdd.n1015 185
R17031 vdd.n2343 vdd.n1021 185
R17032 vdd.n2558 vdd.n1021 185
R17033 vdd.n2345 vdd.n2344 185
R17034 vdd.n2346 vdd.n2345 185
R17035 vdd.n2331 vdd.n1026 185
R17036 vdd.n2552 vdd.n1026 185
R17037 vdd.n2330 vdd.n2329 185
R17038 vdd.n2329 vdd.n1033 185
R17039 vdd.n2328 vdd.n1031 185
R17040 vdd.n2546 vdd.n1031 185
R17041 vdd.n2327 vdd.n2326 185
R17042 vdd.n2326 vdd.n1039 185
R17043 vdd.n1133 vdd.n1037 185
R17044 vdd.n2540 vdd.n1037 185
R17045 vdd.n2360 vdd.n2359 185
R17046 vdd.n2359 vdd.n2358 185
R17047 vdd.n2361 vdd.n1044 185
R17048 vdd.n2534 vdd.n1044 185
R17049 vdd.n2363 vdd.n2362 185
R17050 vdd.n2362 vdd.n1043 185
R17051 vdd.n2364 vdd.n1050 185
R17052 vdd.n2528 vdd.n1050 185
R17053 vdd.n2366 vdd.n2365 185
R17054 vdd.n2365 vdd.n1049 185
R17055 vdd.n2367 vdd.n1055 185
R17056 vdd.n2522 vdd.n1055 185
R17057 vdd.n2369 vdd.n2368 185
R17058 vdd.n2368 vdd.n1063 185
R17059 vdd.n2370 vdd.n1061 185
R17060 vdd.n2515 vdd.n1061 185
R17061 vdd.n2372 vdd.n2371 185
R17062 vdd.n2371 vdd.n1070 185
R17063 vdd.n2373 vdd.n1068 185
R17064 vdd.n2509 vdd.n1068 185
R17065 vdd.n2375 vdd.n2374 185
R17066 vdd.n2374 vdd.n1067 185
R17067 vdd.n2376 vdd.n1075 185
R17068 vdd.n2503 vdd.n1075 185
R17069 vdd.n2378 vdd.n2377 185
R17070 vdd.n2377 vdd.n1074 185
R17071 vdd.n2379 vdd.n1081 185
R17072 vdd.n2497 vdd.n1081 185
R17073 vdd.n2381 vdd.n2380 185
R17074 vdd.n2380 vdd.n1080 185
R17075 vdd.n2382 vdd.n1087 185
R17076 vdd.n2491 vdd.n1087 185
R17077 vdd.n2384 vdd.n2383 185
R17078 vdd.n2383 vdd.n1086 185
R17079 vdd.n2385 vdd.n1093 185
R17080 vdd.n2485 vdd.n1093 185
R17081 vdd.n2387 vdd.n2386 185
R17082 vdd.n2386 vdd.n1092 185
R17083 vdd.n2388 vdd.n1099 185
R17084 vdd.n2479 vdd.n1099 185
R17085 vdd.n2390 vdd.n2389 185
R17086 vdd.n2389 vdd.n1098 185
R17087 vdd.n2391 vdd.n1105 185
R17088 vdd.n2473 vdd.n1105 185
R17089 vdd.n2393 vdd.n2392 185
R17090 vdd.n2392 vdd.n1104 185
R17091 vdd.n2394 vdd.n1111 185
R17092 vdd.n2467 vdd.n1111 185
R17093 vdd.n3539 vdd.n3538 185
R17094 vdd.n3538 vdd.n3537 185
R17095 vdd.n3540 vdd.n387 185
R17096 vdd.n387 vdd.n386 185
R17097 vdd.n3542 vdd.n3541 185
R17098 vdd.n3543 vdd.n3542 185
R17099 vdd.n382 vdd.n381 185
R17100 vdd.n3544 vdd.n382 185
R17101 vdd.n3547 vdd.n3546 185
R17102 vdd.n3546 vdd.n3545 185
R17103 vdd.n3548 vdd.n376 185
R17104 vdd.n376 vdd.n375 185
R17105 vdd.n3550 vdd.n3549 185
R17106 vdd.n3551 vdd.n3550 185
R17107 vdd.n371 vdd.n370 185
R17108 vdd.n3552 vdd.n371 185
R17109 vdd.n3555 vdd.n3554 185
R17110 vdd.n3554 vdd.n3553 185
R17111 vdd.n3556 vdd.n365 185
R17112 vdd.n3513 vdd.n365 185
R17113 vdd.n3558 vdd.n3557 185
R17114 vdd.n3559 vdd.n3558 185
R17115 vdd.n360 vdd.n359 185
R17116 vdd.n3560 vdd.n360 185
R17117 vdd.n3563 vdd.n3562 185
R17118 vdd.n3562 vdd.n3561 185
R17119 vdd.n3564 vdd.n354 185
R17120 vdd.n361 vdd.n354 185
R17121 vdd.n3566 vdd.n3565 185
R17122 vdd.n3567 vdd.n3566 185
R17123 vdd.n350 vdd.n349 185
R17124 vdd.n3568 vdd.n350 185
R17125 vdd.n3571 vdd.n3570 185
R17126 vdd.n3570 vdd.n3569 185
R17127 vdd.n3572 vdd.n345 185
R17128 vdd.n345 vdd.n344 185
R17129 vdd.n3574 vdd.n3573 185
R17130 vdd.n3575 vdd.n3574 185
R17131 vdd.n339 vdd.n337 185
R17132 vdd.n3576 vdd.n339 185
R17133 vdd.n3579 vdd.n3578 185
R17134 vdd.n3578 vdd.n3577 185
R17135 vdd.n338 vdd.n336 185
R17136 vdd.n340 vdd.n338 185
R17137 vdd.n3489 vdd.n3488 185
R17138 vdd.n3490 vdd.n3489 185
R17139 vdd.n635 vdd.n634 185
R17140 vdd.n634 vdd.n633 185
R17141 vdd.n3484 vdd.n3483 185
R17142 vdd.n3483 vdd.n3482 185
R17143 vdd.n638 vdd.n637 185
R17144 vdd.n644 vdd.n638 185
R17145 vdd.n3470 vdd.n3469 185
R17146 vdd.n3471 vdd.n3470 185
R17147 vdd.n646 vdd.n645 185
R17148 vdd.n3462 vdd.n645 185
R17149 vdd.n3465 vdd.n3464 185
R17150 vdd.n3464 vdd.n3463 185
R17151 vdd.n649 vdd.n648 185
R17152 vdd.n656 vdd.n649 185
R17153 vdd.n3453 vdd.n3452 185
R17154 vdd.n3454 vdd.n3453 185
R17155 vdd.n658 vdd.n657 185
R17156 vdd.n657 vdd.n655 185
R17157 vdd.n3448 vdd.n3447 185
R17158 vdd.n3447 vdd.n3446 185
R17159 vdd.n661 vdd.n660 185
R17160 vdd.n662 vdd.n661 185
R17161 vdd.n3437 vdd.n3436 185
R17162 vdd.n3438 vdd.n3437 185
R17163 vdd.n669 vdd.n668 185
R17164 vdd.n3429 vdd.n668 185
R17165 vdd.n3432 vdd.n3431 185
R17166 vdd.n3431 vdd.n3430 185
R17167 vdd.n672 vdd.n671 185
R17168 vdd.n679 vdd.n672 185
R17169 vdd.n3420 vdd.n3419 185
R17170 vdd.n3421 vdd.n3420 185
R17171 vdd.n681 vdd.n680 185
R17172 vdd.n680 vdd.n678 185
R17173 vdd.n3415 vdd.n3414 185
R17174 vdd.n3414 vdd.n3413 185
R17175 vdd.n684 vdd.n683 185
R17176 vdd.n723 vdd.n684 185
R17177 vdd.n3403 vdd.n3402 185
R17178 vdd.n3401 vdd.n725 185
R17179 vdd.n3400 vdd.n724 185
R17180 vdd.n3405 vdd.n724 185
R17181 vdd.n729 vdd.n728 185
R17182 vdd.n733 vdd.n732 185
R17183 vdd.n3396 vdd.n734 185
R17184 vdd.n3395 vdd.n3394 185
R17185 vdd.n3393 vdd.n3392 185
R17186 vdd.n3391 vdd.n3390 185
R17187 vdd.n3389 vdd.n3388 185
R17188 vdd.n3387 vdd.n3386 185
R17189 vdd.n3385 vdd.n3384 185
R17190 vdd.n3383 vdd.n3382 185
R17191 vdd.n3381 vdd.n3380 185
R17192 vdd.n3379 vdd.n3378 185
R17193 vdd.n3377 vdd.n3376 185
R17194 vdd.n3375 vdd.n3374 185
R17195 vdd.n3373 vdd.n3372 185
R17196 vdd.n3371 vdd.n3370 185
R17197 vdd.n3369 vdd.n3368 185
R17198 vdd.n3360 vdd.n747 185
R17199 vdd.n3362 vdd.n3361 185
R17200 vdd.n3359 vdd.n3358 185
R17201 vdd.n3357 vdd.n3356 185
R17202 vdd.n3355 vdd.n3354 185
R17203 vdd.n3353 vdd.n3352 185
R17204 vdd.n3351 vdd.n3350 185
R17205 vdd.n3349 vdd.n3348 185
R17206 vdd.n3347 vdd.n3346 185
R17207 vdd.n3345 vdd.n3344 185
R17208 vdd.n3343 vdd.n3342 185
R17209 vdd.n3341 vdd.n3340 185
R17210 vdd.n3339 vdd.n3338 185
R17211 vdd.n3337 vdd.n3336 185
R17212 vdd.n3335 vdd.n3334 185
R17213 vdd.n3333 vdd.n3332 185
R17214 vdd.n3331 vdd.n3330 185
R17215 vdd.n3329 vdd.n3328 185
R17216 vdd.n3327 vdd.n3326 185
R17217 vdd.n3325 vdd.n3324 185
R17218 vdd.n3323 vdd.n3322 185
R17219 vdd.n3321 vdd.n3320 185
R17220 vdd.n3314 vdd.n767 185
R17221 vdd.n3316 vdd.n3315 185
R17222 vdd.n3313 vdd.n3312 185
R17223 vdd.n3311 vdd.n3310 185
R17224 vdd.n3309 vdd.n3308 185
R17225 vdd.n3307 vdd.n3306 185
R17226 vdd.n3305 vdd.n3304 185
R17227 vdd.n3303 vdd.n3302 185
R17228 vdd.n3301 vdd.n3300 185
R17229 vdd.n3299 vdd.n3298 185
R17230 vdd.n3297 vdd.n3296 185
R17231 vdd.n3295 vdd.n3294 185
R17232 vdd.n3293 vdd.n3292 185
R17233 vdd.n3291 vdd.n3290 185
R17234 vdd.n3289 vdd.n3288 185
R17235 vdd.n3287 vdd.n3286 185
R17236 vdd.n3285 vdd.n3284 185
R17237 vdd.n3283 vdd.n3282 185
R17238 vdd.n3281 vdd.n3280 185
R17239 vdd.n3279 vdd.n3278 185
R17240 vdd.n3277 vdd.n691 185
R17241 vdd.n3407 vdd.n3406 185
R17242 vdd.n3406 vdd.n3405 185
R17243 vdd.n3534 vdd.n3533 185
R17244 vdd.n618 vdd.n425 185
R17245 vdd.n617 vdd.n616 185
R17246 vdd.n615 vdd.n614 185
R17247 vdd.n613 vdd.n430 185
R17248 vdd.n609 vdd.n608 185
R17249 vdd.n607 vdd.n606 185
R17250 vdd.n605 vdd.n604 185
R17251 vdd.n603 vdd.n432 185
R17252 vdd.n599 vdd.n598 185
R17253 vdd.n597 vdd.n596 185
R17254 vdd.n595 vdd.n594 185
R17255 vdd.n593 vdd.n434 185
R17256 vdd.n589 vdd.n588 185
R17257 vdd.n587 vdd.n586 185
R17258 vdd.n585 vdd.n584 185
R17259 vdd.n583 vdd.n436 185
R17260 vdd.n579 vdd.n578 185
R17261 vdd.n577 vdd.n576 185
R17262 vdd.n575 vdd.n574 185
R17263 vdd.n573 vdd.n438 185
R17264 vdd.n569 vdd.n568 185
R17265 vdd.n567 vdd.n566 185
R17266 vdd.n565 vdd.n564 185
R17267 vdd.n563 vdd.n442 185
R17268 vdd.n559 vdd.n558 185
R17269 vdd.n557 vdd.n556 185
R17270 vdd.n555 vdd.n554 185
R17271 vdd.n553 vdd.n444 185
R17272 vdd.n549 vdd.n548 185
R17273 vdd.n547 vdd.n546 185
R17274 vdd.n545 vdd.n544 185
R17275 vdd.n543 vdd.n446 185
R17276 vdd.n539 vdd.n538 185
R17277 vdd.n537 vdd.n536 185
R17278 vdd.n535 vdd.n534 185
R17279 vdd.n533 vdd.n448 185
R17280 vdd.n529 vdd.n528 185
R17281 vdd.n527 vdd.n526 185
R17282 vdd.n525 vdd.n524 185
R17283 vdd.n523 vdd.n450 185
R17284 vdd.n519 vdd.n518 185
R17285 vdd.n517 vdd.n516 185
R17286 vdd.n515 vdd.n514 185
R17287 vdd.n513 vdd.n454 185
R17288 vdd.n509 vdd.n508 185
R17289 vdd.n507 vdd.n506 185
R17290 vdd.n505 vdd.n504 185
R17291 vdd.n503 vdd.n456 185
R17292 vdd.n499 vdd.n498 185
R17293 vdd.n497 vdd.n496 185
R17294 vdd.n495 vdd.n494 185
R17295 vdd.n493 vdd.n458 185
R17296 vdd.n489 vdd.n488 185
R17297 vdd.n487 vdd.n486 185
R17298 vdd.n485 vdd.n484 185
R17299 vdd.n483 vdd.n460 185
R17300 vdd.n479 vdd.n478 185
R17301 vdd.n477 vdd.n476 185
R17302 vdd.n475 vdd.n474 185
R17303 vdd.n473 vdd.n462 185
R17304 vdd.n469 vdd.n468 185
R17305 vdd.n467 vdd.n466 185
R17306 vdd.n465 vdd.n392 185
R17307 vdd.n3530 vdd.n393 185
R17308 vdd.n3537 vdd.n393 185
R17309 vdd.n3529 vdd.n3528 185
R17310 vdd.n3528 vdd.n386 185
R17311 vdd.n3527 vdd.n385 185
R17312 vdd.n3543 vdd.n385 185
R17313 vdd.n621 vdd.n384 185
R17314 vdd.n3544 vdd.n384 185
R17315 vdd.n3523 vdd.n383 185
R17316 vdd.n3545 vdd.n383 185
R17317 vdd.n3522 vdd.n3521 185
R17318 vdd.n3521 vdd.n375 185
R17319 vdd.n3520 vdd.n374 185
R17320 vdd.n3551 vdd.n374 185
R17321 vdd.n623 vdd.n373 185
R17322 vdd.n3552 vdd.n373 185
R17323 vdd.n3516 vdd.n372 185
R17324 vdd.n3553 vdd.n372 185
R17325 vdd.n3515 vdd.n3514 185
R17326 vdd.n3514 vdd.n3513 185
R17327 vdd.n3512 vdd.n364 185
R17328 vdd.n3559 vdd.n364 185
R17329 vdd.n625 vdd.n363 185
R17330 vdd.n3560 vdd.n363 185
R17331 vdd.n3508 vdd.n362 185
R17332 vdd.n3561 vdd.n362 185
R17333 vdd.n3507 vdd.n3506 185
R17334 vdd.n3506 vdd.n361 185
R17335 vdd.n3505 vdd.n353 185
R17336 vdd.n3567 vdd.n353 185
R17337 vdd.n627 vdd.n352 185
R17338 vdd.n3568 vdd.n352 185
R17339 vdd.n3501 vdd.n351 185
R17340 vdd.n3569 vdd.n351 185
R17341 vdd.n3500 vdd.n3499 185
R17342 vdd.n3499 vdd.n344 185
R17343 vdd.n3498 vdd.n343 185
R17344 vdd.n3575 vdd.n343 185
R17345 vdd.n629 vdd.n342 185
R17346 vdd.n3576 vdd.n342 185
R17347 vdd.n3494 vdd.n341 185
R17348 vdd.n3577 vdd.n341 185
R17349 vdd.n3493 vdd.n3492 185
R17350 vdd.n3492 vdd.n340 185
R17351 vdd.n3491 vdd.n631 185
R17352 vdd.n3491 vdd.n3490 185
R17353 vdd.n3479 vdd.n632 185
R17354 vdd.n633 vdd.n632 185
R17355 vdd.n3481 vdd.n3480 185
R17356 vdd.n3482 vdd.n3481 185
R17357 vdd.n640 vdd.n639 185
R17358 vdd.n644 vdd.n639 185
R17359 vdd.n3473 vdd.n3472 185
R17360 vdd.n3472 vdd.n3471 185
R17361 vdd.n643 vdd.n642 185
R17362 vdd.n3462 vdd.n643 185
R17363 vdd.n3461 vdd.n3460 185
R17364 vdd.n3463 vdd.n3461 185
R17365 vdd.n651 vdd.n650 185
R17366 vdd.n656 vdd.n650 185
R17367 vdd.n3456 vdd.n3455 185
R17368 vdd.n3455 vdd.n3454 185
R17369 vdd.n654 vdd.n653 185
R17370 vdd.n655 vdd.n654 185
R17371 vdd.n3445 vdd.n3444 185
R17372 vdd.n3446 vdd.n3445 185
R17373 vdd.n664 vdd.n663 185
R17374 vdd.n663 vdd.n662 185
R17375 vdd.n3440 vdd.n3439 185
R17376 vdd.n3439 vdd.n3438 185
R17377 vdd.n667 vdd.n666 185
R17378 vdd.n3429 vdd.n667 185
R17379 vdd.n3428 vdd.n3427 185
R17380 vdd.n3430 vdd.n3428 185
R17381 vdd.n674 vdd.n673 185
R17382 vdd.n679 vdd.n673 185
R17383 vdd.n3423 vdd.n3422 185
R17384 vdd.n3422 vdd.n3421 185
R17385 vdd.n677 vdd.n676 185
R17386 vdd.n678 vdd.n677 185
R17387 vdd.n3412 vdd.n3411 185
R17388 vdd.n3413 vdd.n3412 185
R17389 vdd.n686 vdd.n685 185
R17390 vdd.n723 vdd.n685 185
R17391 vdd.n3014 vdd.n947 185
R17392 vdd.n3013 vdd.n3012 185
R17393 vdd.n949 vdd.n948 185
R17394 vdd.n3010 vdd.n949 185
R17395 vdd.n2833 vdd.n2832 185
R17396 vdd.n2835 vdd.n2834 185
R17397 vdd.n2837 vdd.n2836 185
R17398 vdd.n2839 vdd.n2838 185
R17399 vdd.n2841 vdd.n2840 185
R17400 vdd.n2843 vdd.n2842 185
R17401 vdd.n2845 vdd.n2844 185
R17402 vdd.n2847 vdd.n2846 185
R17403 vdd.n2849 vdd.n2848 185
R17404 vdd.n2851 vdd.n2850 185
R17405 vdd.n2853 vdd.n2852 185
R17406 vdd.n2855 vdd.n2854 185
R17407 vdd.n2857 vdd.n2856 185
R17408 vdd.n2859 vdd.n2858 185
R17409 vdd.n2861 vdd.n2860 185
R17410 vdd.n2863 vdd.n2862 185
R17411 vdd.n2865 vdd.n2864 185
R17412 vdd.n2867 vdd.n2866 185
R17413 vdd.n2869 vdd.n2868 185
R17414 vdd.n2871 vdd.n2870 185
R17415 vdd.n2873 vdd.n2872 185
R17416 vdd.n2875 vdd.n2874 185
R17417 vdd.n2877 vdd.n2876 185
R17418 vdd.n2879 vdd.n2878 185
R17419 vdd.n2881 vdd.n2880 185
R17420 vdd.n2883 vdd.n2882 185
R17421 vdd.n2885 vdd.n2884 185
R17422 vdd.n2887 vdd.n2886 185
R17423 vdd.n2889 vdd.n2888 185
R17424 vdd.n2892 vdd.n2891 185
R17425 vdd.n2894 vdd.n2893 185
R17426 vdd.n2896 vdd.n2895 185
R17427 vdd.n3177 vdd.n3176 185
R17428 vdd.n3179 vdd.n834 185
R17429 vdd.n3181 vdd.n3180 185
R17430 vdd.n3183 vdd.n831 185
R17431 vdd.n3185 vdd.n3184 185
R17432 vdd.n3187 vdd.n829 185
R17433 vdd.n3189 vdd.n3188 185
R17434 vdd.n3190 vdd.n828 185
R17435 vdd.n3192 vdd.n3191 185
R17436 vdd.n3194 vdd.n826 185
R17437 vdd.n3196 vdd.n3195 185
R17438 vdd.n3197 vdd.n825 185
R17439 vdd.n3199 vdd.n3198 185
R17440 vdd.n3201 vdd.n823 185
R17441 vdd.n3203 vdd.n3202 185
R17442 vdd.n3204 vdd.n822 185
R17443 vdd.n3206 vdd.n3205 185
R17444 vdd.n3208 vdd.n731 185
R17445 vdd.n3210 vdd.n3209 185
R17446 vdd.n3212 vdd.n820 185
R17447 vdd.n3214 vdd.n3213 185
R17448 vdd.n3215 vdd.n819 185
R17449 vdd.n3217 vdd.n3216 185
R17450 vdd.n3219 vdd.n817 185
R17451 vdd.n3221 vdd.n3220 185
R17452 vdd.n3222 vdd.n816 185
R17453 vdd.n3224 vdd.n3223 185
R17454 vdd.n3226 vdd.n814 185
R17455 vdd.n3228 vdd.n3227 185
R17456 vdd.n3229 vdd.n813 185
R17457 vdd.n3231 vdd.n3230 185
R17458 vdd.n3233 vdd.n812 185
R17459 vdd.n3234 vdd.n811 185
R17460 vdd.n3237 vdd.n3236 185
R17461 vdd.n3238 vdd.n809 185
R17462 vdd.n809 vdd.n692 185
R17463 vdd.n3175 vdd.n806 185
R17464 vdd.n3241 vdd.n806 185
R17465 vdd.n3174 vdd.n3173 185
R17466 vdd.n3173 vdd.n805 185
R17467 vdd.n3172 vdd.n836 185
R17468 vdd.n3172 vdd.n3171 185
R17469 vdd.n2946 vdd.n837 185
R17470 vdd.n846 vdd.n837 185
R17471 vdd.n2947 vdd.n844 185
R17472 vdd.n3165 vdd.n844 185
R17473 vdd.n2949 vdd.n2948 185
R17474 vdd.n2948 vdd.n843 185
R17475 vdd.n2950 vdd.n852 185
R17476 vdd.n3114 vdd.n852 185
R17477 vdd.n2952 vdd.n2951 185
R17478 vdd.n2951 vdd.n851 185
R17479 vdd.n2953 vdd.n857 185
R17480 vdd.n3108 vdd.n857 185
R17481 vdd.n2955 vdd.n2954 185
R17482 vdd.n2954 vdd.n864 185
R17483 vdd.n2956 vdd.n862 185
R17484 vdd.n3102 vdd.n862 185
R17485 vdd.n2958 vdd.n2957 185
R17486 vdd.n2957 vdd.n870 185
R17487 vdd.n2959 vdd.n868 185
R17488 vdd.n3096 vdd.n868 185
R17489 vdd.n2961 vdd.n2960 185
R17490 vdd.n2960 vdd.n877 185
R17491 vdd.n2962 vdd.n875 185
R17492 vdd.n3090 vdd.n875 185
R17493 vdd.n2964 vdd.n2963 185
R17494 vdd.n2963 vdd.n874 185
R17495 vdd.n2965 vdd.n882 185
R17496 vdd.n3084 vdd.n882 185
R17497 vdd.n2967 vdd.n2966 185
R17498 vdd.n2966 vdd.n881 185
R17499 vdd.n2968 vdd.n889 185
R17500 vdd.n3077 vdd.n889 185
R17501 vdd.n2970 vdd.n2969 185
R17502 vdd.n2969 vdd.n888 185
R17503 vdd.n2971 vdd.n894 185
R17504 vdd.n3071 vdd.n894 185
R17505 vdd.n2973 vdd.n2972 185
R17506 vdd.n2972 vdd.n901 185
R17507 vdd.n2974 vdd.n899 185
R17508 vdd.n3065 vdd.n899 185
R17509 vdd.n2976 vdd.n2975 185
R17510 vdd.n2977 vdd.n2976 185
R17511 vdd.n2945 vdd.n906 185
R17512 vdd.n3059 vdd.n906 185
R17513 vdd.n2944 vdd.n2943 185
R17514 vdd.n2943 vdd.n905 185
R17515 vdd.n2942 vdd.n912 185
R17516 vdd.n3053 vdd.n912 185
R17517 vdd.n2941 vdd.n2940 185
R17518 vdd.n2940 vdd.n911 185
R17519 vdd.n2901 vdd.n917 185
R17520 vdd.n3047 vdd.n917 185
R17521 vdd.n2991 vdd.n2990 185
R17522 vdd.n2990 vdd.n2989 185
R17523 vdd.n2992 vdd.n922 185
R17524 vdd.n3041 vdd.n922 185
R17525 vdd.n2994 vdd.n2993 185
R17526 vdd.n2993 vdd.n930 185
R17527 vdd.n2995 vdd.n928 185
R17528 vdd.n3035 vdd.n928 185
R17529 vdd.n2997 vdd.n2996 185
R17530 vdd.n2996 vdd.n927 185
R17531 vdd.n2998 vdd.n934 185
R17532 vdd.n3029 vdd.n934 185
R17533 vdd.n3000 vdd.n2999 185
R17534 vdd.n3001 vdd.n3000 185
R17535 vdd.n2900 vdd.n939 185
R17536 vdd.n3023 vdd.n939 185
R17537 vdd.n2899 vdd.n2898 185
R17538 vdd.n2898 vdd.n946 185
R17539 vdd.n2897 vdd.n944 185
R17540 vdd.n3017 vdd.n944 185
R17541 vdd.n3016 vdd.n3015 185
R17542 vdd.n3017 vdd.n3016 185
R17543 vdd.n938 vdd.n937 185
R17544 vdd.n946 vdd.n938 185
R17545 vdd.n3025 vdd.n3024 185
R17546 vdd.n3024 vdd.n3023 185
R17547 vdd.n3026 vdd.n936 185
R17548 vdd.n3001 vdd.n936 185
R17549 vdd.n3028 vdd.n3027 185
R17550 vdd.n3029 vdd.n3028 185
R17551 vdd.n926 vdd.n925 185
R17552 vdd.n927 vdd.n926 185
R17553 vdd.n3037 vdd.n3036 185
R17554 vdd.n3036 vdd.n3035 185
R17555 vdd.n3038 vdd.n924 185
R17556 vdd.n930 vdd.n924 185
R17557 vdd.n3040 vdd.n3039 185
R17558 vdd.n3041 vdd.n3040 185
R17559 vdd.n916 vdd.n915 185
R17560 vdd.n2989 vdd.n916 185
R17561 vdd.n3049 vdd.n3048 185
R17562 vdd.n3048 vdd.n3047 185
R17563 vdd.n3050 vdd.n914 185
R17564 vdd.n914 vdd.n911 185
R17565 vdd.n3052 vdd.n3051 185
R17566 vdd.n3053 vdd.n3052 185
R17567 vdd.n904 vdd.n903 185
R17568 vdd.n905 vdd.n904 185
R17569 vdd.n3061 vdd.n3060 185
R17570 vdd.n3060 vdd.n3059 185
R17571 vdd.n3062 vdd.n902 185
R17572 vdd.n2977 vdd.n902 185
R17573 vdd.n3064 vdd.n3063 185
R17574 vdd.n3065 vdd.n3064 185
R17575 vdd.n893 vdd.n892 185
R17576 vdd.n901 vdd.n893 185
R17577 vdd.n3073 vdd.n3072 185
R17578 vdd.n3072 vdd.n3071 185
R17579 vdd.n3074 vdd.n891 185
R17580 vdd.n891 vdd.n888 185
R17581 vdd.n3076 vdd.n3075 185
R17582 vdd.n3077 vdd.n3076 185
R17583 vdd.n880 vdd.n879 185
R17584 vdd.n881 vdd.n880 185
R17585 vdd.n3086 vdd.n3085 185
R17586 vdd.n3085 vdd.n3084 185
R17587 vdd.n3087 vdd.n878 185
R17588 vdd.n878 vdd.n874 185
R17589 vdd.n3089 vdd.n3088 185
R17590 vdd.n3090 vdd.n3089 185
R17591 vdd.n867 vdd.n866 185
R17592 vdd.n877 vdd.n867 185
R17593 vdd.n3098 vdd.n3097 185
R17594 vdd.n3097 vdd.n3096 185
R17595 vdd.n3099 vdd.n865 185
R17596 vdd.n870 vdd.n865 185
R17597 vdd.n3101 vdd.n3100 185
R17598 vdd.n3102 vdd.n3101 185
R17599 vdd.n856 vdd.n855 185
R17600 vdd.n864 vdd.n856 185
R17601 vdd.n3110 vdd.n3109 185
R17602 vdd.n3109 vdd.n3108 185
R17603 vdd.n3111 vdd.n854 185
R17604 vdd.n854 vdd.n851 185
R17605 vdd.n3113 vdd.n3112 185
R17606 vdd.n3114 vdd.n3113 185
R17607 vdd.n842 vdd.n841 185
R17608 vdd.n843 vdd.n842 185
R17609 vdd.n3167 vdd.n3166 185
R17610 vdd.n3166 vdd.n3165 185
R17611 vdd.n3168 vdd.n840 185
R17612 vdd.n846 vdd.n840 185
R17613 vdd.n3170 vdd.n3169 185
R17614 vdd.n3171 vdd.n3170 185
R17615 vdd.n810 vdd.n808 185
R17616 vdd.n808 vdd.n805 185
R17617 vdd.n3240 vdd.n3239 185
R17618 vdd.n3241 vdd.n3240 185
R17619 vdd.n2653 vdd.n2652 185
R17620 vdd.n2654 vdd.n2653 185
R17621 vdd.n996 vdd.n994 185
R17622 vdd.n994 vdd.n992 185
R17623 vdd.n2568 vdd.n1003 185
R17624 vdd.n2579 vdd.n1003 185
R17625 vdd.n2569 vdd.n1012 185
R17626 vdd.n2334 vdd.n1012 185
R17627 vdd.n2571 vdd.n2570 185
R17628 vdd.n2572 vdd.n2571 185
R17629 vdd.n2567 vdd.n1011 185
R17630 vdd.n1011 vdd.n1008 185
R17631 vdd.n2566 vdd.n2565 185
R17632 vdd.n2565 vdd.n2564 185
R17633 vdd.n1014 vdd.n1013 185
R17634 vdd.n1015 vdd.n1014 185
R17635 vdd.n2557 vdd.n2556 185
R17636 vdd.n2558 vdd.n2557 185
R17637 vdd.n2555 vdd.n1023 185
R17638 vdd.n2346 vdd.n1023 185
R17639 vdd.n2554 vdd.n2553 185
R17640 vdd.n2553 vdd.n2552 185
R17641 vdd.n1025 vdd.n1024 185
R17642 vdd.n1033 vdd.n1025 185
R17643 vdd.n2545 vdd.n2544 185
R17644 vdd.n2546 vdd.n2545 185
R17645 vdd.n2543 vdd.n1034 185
R17646 vdd.n1039 vdd.n1034 185
R17647 vdd.n2542 vdd.n2541 185
R17648 vdd.n2541 vdd.n2540 185
R17649 vdd.n1036 vdd.n1035 185
R17650 vdd.n2358 vdd.n1036 185
R17651 vdd.n2533 vdd.n2532 185
R17652 vdd.n2534 vdd.n2533 185
R17653 vdd.n2531 vdd.n1046 185
R17654 vdd.n1046 vdd.n1043 185
R17655 vdd.n2530 vdd.n2529 185
R17656 vdd.n2529 vdd.n2528 185
R17657 vdd.n1048 vdd.n1047 185
R17658 vdd.n1049 vdd.n1048 185
R17659 vdd.n2521 vdd.n2520 185
R17660 vdd.n2522 vdd.n2521 185
R17661 vdd.n2518 vdd.n1057 185
R17662 vdd.n1063 vdd.n1057 185
R17663 vdd.n2517 vdd.n2516 185
R17664 vdd.n2516 vdd.n2515 185
R17665 vdd.n1060 vdd.n1059 185
R17666 vdd.n1070 vdd.n1060 185
R17667 vdd.n2508 vdd.n2507 185
R17668 vdd.n2509 vdd.n2508 185
R17669 vdd.n2506 vdd.n1071 185
R17670 vdd.n1071 vdd.n1067 185
R17671 vdd.n2505 vdd.n2504 185
R17672 vdd.n2504 vdd.n2503 185
R17673 vdd.n1073 vdd.n1072 185
R17674 vdd.n1074 vdd.n1073 185
R17675 vdd.n2496 vdd.n2495 185
R17676 vdd.n2497 vdd.n2496 185
R17677 vdd.n2494 vdd.n1083 185
R17678 vdd.n1083 vdd.n1080 185
R17679 vdd.n2493 vdd.n2492 185
R17680 vdd.n2492 vdd.n2491 185
R17681 vdd.n1085 vdd.n1084 185
R17682 vdd.n1086 vdd.n1085 185
R17683 vdd.n2484 vdd.n2483 185
R17684 vdd.n2485 vdd.n2484 185
R17685 vdd.n2482 vdd.n1095 185
R17686 vdd.n1095 vdd.n1092 185
R17687 vdd.n2481 vdd.n2480 185
R17688 vdd.n2480 vdd.n2479 185
R17689 vdd.n1097 vdd.n1096 185
R17690 vdd.n1098 vdd.n1097 185
R17691 vdd.n2472 vdd.n2471 185
R17692 vdd.n2473 vdd.n2472 185
R17693 vdd.n2470 vdd.n1107 185
R17694 vdd.n1107 vdd.n1104 185
R17695 vdd.n2469 vdd.n2468 185
R17696 vdd.n2468 vdd.n2467 185
R17697 vdd.n2584 vdd.n967 185
R17698 vdd.n2726 vdd.n967 185
R17699 vdd.n2586 vdd.n2585 185
R17700 vdd.n2588 vdd.n2587 185
R17701 vdd.n2590 vdd.n2589 185
R17702 vdd.n2592 vdd.n2591 185
R17703 vdd.n2594 vdd.n2593 185
R17704 vdd.n2596 vdd.n2595 185
R17705 vdd.n2598 vdd.n2597 185
R17706 vdd.n2600 vdd.n2599 185
R17707 vdd.n2602 vdd.n2601 185
R17708 vdd.n2604 vdd.n2603 185
R17709 vdd.n2606 vdd.n2605 185
R17710 vdd.n2608 vdd.n2607 185
R17711 vdd.n2610 vdd.n2609 185
R17712 vdd.n2612 vdd.n2611 185
R17713 vdd.n2614 vdd.n2613 185
R17714 vdd.n2616 vdd.n2615 185
R17715 vdd.n2618 vdd.n2617 185
R17716 vdd.n2620 vdd.n2619 185
R17717 vdd.n2622 vdd.n2621 185
R17718 vdd.n2624 vdd.n2623 185
R17719 vdd.n2626 vdd.n2625 185
R17720 vdd.n2628 vdd.n2627 185
R17721 vdd.n2630 vdd.n2629 185
R17722 vdd.n2632 vdd.n2631 185
R17723 vdd.n2634 vdd.n2633 185
R17724 vdd.n2636 vdd.n2635 185
R17725 vdd.n2638 vdd.n2637 185
R17726 vdd.n2640 vdd.n2639 185
R17727 vdd.n2642 vdd.n2641 185
R17728 vdd.n2644 vdd.n2643 185
R17729 vdd.n2646 vdd.n2645 185
R17730 vdd.n2648 vdd.n2647 185
R17731 vdd.n2650 vdd.n2649 185
R17732 vdd.n2651 vdd.n995 185
R17733 vdd.n2583 vdd.n993 185
R17734 vdd.n2654 vdd.n993 185
R17735 vdd.n2582 vdd.n2581 185
R17736 vdd.n2581 vdd.n992 185
R17737 vdd.n2580 vdd.n1000 185
R17738 vdd.n2580 vdd.n2579 185
R17739 vdd.n2318 vdd.n1001 185
R17740 vdd.n2334 vdd.n1001 185
R17741 vdd.n2319 vdd.n1010 185
R17742 vdd.n2572 vdd.n1010 185
R17743 vdd.n2321 vdd.n2320 185
R17744 vdd.n2320 vdd.n1008 185
R17745 vdd.n2322 vdd.n1017 185
R17746 vdd.n2564 vdd.n1017 185
R17747 vdd.n2324 vdd.n2323 185
R17748 vdd.n2323 vdd.n1015 185
R17749 vdd.n2325 vdd.n1022 185
R17750 vdd.n2558 vdd.n1022 185
R17751 vdd.n2348 vdd.n2347 185
R17752 vdd.n2347 vdd.n2346 185
R17753 vdd.n2349 vdd.n1027 185
R17754 vdd.n2552 vdd.n1027 185
R17755 vdd.n2351 vdd.n2350 185
R17756 vdd.n2350 vdd.n1033 185
R17757 vdd.n2352 vdd.n1032 185
R17758 vdd.n2546 vdd.n1032 185
R17759 vdd.n2354 vdd.n2353 185
R17760 vdd.n2353 vdd.n1039 185
R17761 vdd.n2355 vdd.n1038 185
R17762 vdd.n2540 vdd.n1038 185
R17763 vdd.n2357 vdd.n2356 185
R17764 vdd.n2358 vdd.n2357 185
R17765 vdd.n2317 vdd.n1045 185
R17766 vdd.n2534 vdd.n1045 185
R17767 vdd.n2316 vdd.n2315 185
R17768 vdd.n2315 vdd.n1043 185
R17769 vdd.n2314 vdd.n1051 185
R17770 vdd.n2528 vdd.n1051 185
R17771 vdd.n2313 vdd.n2312 185
R17772 vdd.n2312 vdd.n1049 185
R17773 vdd.n2311 vdd.n1056 185
R17774 vdd.n2522 vdd.n1056 185
R17775 vdd.n2310 vdd.n2309 185
R17776 vdd.n2309 vdd.n1063 185
R17777 vdd.n2308 vdd.n1062 185
R17778 vdd.n2515 vdd.n1062 185
R17779 vdd.n2307 vdd.n2306 185
R17780 vdd.n2306 vdd.n1070 185
R17781 vdd.n2305 vdd.n1069 185
R17782 vdd.n2509 vdd.n1069 185
R17783 vdd.n2304 vdd.n2303 185
R17784 vdd.n2303 vdd.n1067 185
R17785 vdd.n2302 vdd.n1076 185
R17786 vdd.n2503 vdd.n1076 185
R17787 vdd.n2301 vdd.n2300 185
R17788 vdd.n2300 vdd.n1074 185
R17789 vdd.n2299 vdd.n1082 185
R17790 vdd.n2497 vdd.n1082 185
R17791 vdd.n2298 vdd.n2297 185
R17792 vdd.n2297 vdd.n1080 185
R17793 vdd.n2296 vdd.n1088 185
R17794 vdd.n2491 vdd.n1088 185
R17795 vdd.n2295 vdd.n2294 185
R17796 vdd.n2294 vdd.n1086 185
R17797 vdd.n2293 vdd.n1094 185
R17798 vdd.n2485 vdd.n1094 185
R17799 vdd.n2292 vdd.n2291 185
R17800 vdd.n2291 vdd.n1092 185
R17801 vdd.n2290 vdd.n1100 185
R17802 vdd.n2479 vdd.n1100 185
R17803 vdd.n2289 vdd.n2288 185
R17804 vdd.n2288 vdd.n1098 185
R17805 vdd.n2287 vdd.n1106 185
R17806 vdd.n2473 vdd.n1106 185
R17807 vdd.n2286 vdd.n2285 185
R17808 vdd.n2285 vdd.n1104 185
R17809 vdd.n2284 vdd.n1112 185
R17810 vdd.n2467 vdd.n1112 185
R17811 vdd.n1109 vdd.n1108 185
R17812 vdd.n2216 vdd.n2214 185
R17813 vdd.n2219 vdd.n2218 185
R17814 vdd.n2220 vdd.n2213 185
R17815 vdd.n2222 vdd.n2221 185
R17816 vdd.n2224 vdd.n2212 185
R17817 vdd.n2227 vdd.n2226 185
R17818 vdd.n2228 vdd.n2211 185
R17819 vdd.n2230 vdd.n2229 185
R17820 vdd.n2232 vdd.n2210 185
R17821 vdd.n2235 vdd.n2234 185
R17822 vdd.n2236 vdd.n2209 185
R17823 vdd.n2238 vdd.n2237 185
R17824 vdd.n2240 vdd.n2208 185
R17825 vdd.n2243 vdd.n2242 185
R17826 vdd.n2244 vdd.n2207 185
R17827 vdd.n2246 vdd.n2245 185
R17828 vdd.n2248 vdd.n2206 185
R17829 vdd.n2251 vdd.n2250 185
R17830 vdd.n2252 vdd.n1143 185
R17831 vdd.n2254 vdd.n2253 185
R17832 vdd.n2256 vdd.n1142 185
R17833 vdd.n2259 vdd.n2258 185
R17834 vdd.n2260 vdd.n1141 185
R17835 vdd.n2262 vdd.n2261 185
R17836 vdd.n2264 vdd.n1140 185
R17837 vdd.n2267 vdd.n2266 185
R17838 vdd.n2268 vdd.n1139 185
R17839 vdd.n2270 vdd.n2269 185
R17840 vdd.n2272 vdd.n1138 185
R17841 vdd.n2275 vdd.n2274 185
R17842 vdd.n2276 vdd.n1135 185
R17843 vdd.n2279 vdd.n2278 185
R17844 vdd.n2281 vdd.n1134 185
R17845 vdd.n2283 vdd.n2282 185
R17846 vdd.n2282 vdd.n1110 185
R17847 vdd.n327 vdd.n326 171.744
R17848 vdd.n326 vdd.n325 171.744
R17849 vdd.n325 vdd.n294 171.744
R17850 vdd.n318 vdd.n294 171.744
R17851 vdd.n318 vdd.n317 171.744
R17852 vdd.n317 vdd.n299 171.744
R17853 vdd.n310 vdd.n299 171.744
R17854 vdd.n310 vdd.n309 171.744
R17855 vdd.n309 vdd.n303 171.744
R17856 vdd.n268 vdd.n267 171.744
R17857 vdd.n267 vdd.n266 171.744
R17858 vdd.n266 vdd.n235 171.744
R17859 vdd.n259 vdd.n235 171.744
R17860 vdd.n259 vdd.n258 171.744
R17861 vdd.n258 vdd.n240 171.744
R17862 vdd.n251 vdd.n240 171.744
R17863 vdd.n251 vdd.n250 171.744
R17864 vdd.n250 vdd.n244 171.744
R17865 vdd.n225 vdd.n224 171.744
R17866 vdd.n224 vdd.n223 171.744
R17867 vdd.n223 vdd.n192 171.744
R17868 vdd.n216 vdd.n192 171.744
R17869 vdd.n216 vdd.n215 171.744
R17870 vdd.n215 vdd.n197 171.744
R17871 vdd.n208 vdd.n197 171.744
R17872 vdd.n208 vdd.n207 171.744
R17873 vdd.n207 vdd.n201 171.744
R17874 vdd.n166 vdd.n165 171.744
R17875 vdd.n165 vdd.n164 171.744
R17876 vdd.n164 vdd.n133 171.744
R17877 vdd.n157 vdd.n133 171.744
R17878 vdd.n157 vdd.n156 171.744
R17879 vdd.n156 vdd.n138 171.744
R17880 vdd.n149 vdd.n138 171.744
R17881 vdd.n149 vdd.n148 171.744
R17882 vdd.n148 vdd.n142 171.744
R17883 vdd.n124 vdd.n123 171.744
R17884 vdd.n123 vdd.n122 171.744
R17885 vdd.n122 vdd.n91 171.744
R17886 vdd.n115 vdd.n91 171.744
R17887 vdd.n115 vdd.n114 171.744
R17888 vdd.n114 vdd.n96 171.744
R17889 vdd.n107 vdd.n96 171.744
R17890 vdd.n107 vdd.n106 171.744
R17891 vdd.n106 vdd.n100 171.744
R17892 vdd.n65 vdd.n64 171.744
R17893 vdd.n64 vdd.n63 171.744
R17894 vdd.n63 vdd.n32 171.744
R17895 vdd.n56 vdd.n32 171.744
R17896 vdd.n56 vdd.n55 171.744
R17897 vdd.n55 vdd.n37 171.744
R17898 vdd.n48 vdd.n37 171.744
R17899 vdd.n48 vdd.n47 171.744
R17900 vdd.n47 vdd.n41 171.744
R17901 vdd.n1826 vdd.n1825 171.744
R17902 vdd.n1825 vdd.n1824 171.744
R17903 vdd.n1824 vdd.n1793 171.744
R17904 vdd.n1817 vdd.n1793 171.744
R17905 vdd.n1817 vdd.n1816 171.744
R17906 vdd.n1816 vdd.n1798 171.744
R17907 vdd.n1809 vdd.n1798 171.744
R17908 vdd.n1809 vdd.n1808 171.744
R17909 vdd.n1808 vdd.n1802 171.744
R17910 vdd.n1885 vdd.n1884 171.744
R17911 vdd.n1884 vdd.n1883 171.744
R17912 vdd.n1883 vdd.n1852 171.744
R17913 vdd.n1876 vdd.n1852 171.744
R17914 vdd.n1876 vdd.n1875 171.744
R17915 vdd.n1875 vdd.n1857 171.744
R17916 vdd.n1868 vdd.n1857 171.744
R17917 vdd.n1868 vdd.n1867 171.744
R17918 vdd.n1867 vdd.n1861 171.744
R17919 vdd.n1724 vdd.n1723 171.744
R17920 vdd.n1723 vdd.n1722 171.744
R17921 vdd.n1722 vdd.n1691 171.744
R17922 vdd.n1715 vdd.n1691 171.744
R17923 vdd.n1715 vdd.n1714 171.744
R17924 vdd.n1714 vdd.n1696 171.744
R17925 vdd.n1707 vdd.n1696 171.744
R17926 vdd.n1707 vdd.n1706 171.744
R17927 vdd.n1706 vdd.n1700 171.744
R17928 vdd.n1783 vdd.n1782 171.744
R17929 vdd.n1782 vdd.n1781 171.744
R17930 vdd.n1781 vdd.n1750 171.744
R17931 vdd.n1774 vdd.n1750 171.744
R17932 vdd.n1774 vdd.n1773 171.744
R17933 vdd.n1773 vdd.n1755 171.744
R17934 vdd.n1766 vdd.n1755 171.744
R17935 vdd.n1766 vdd.n1765 171.744
R17936 vdd.n1765 vdd.n1759 171.744
R17937 vdd.n1623 vdd.n1622 171.744
R17938 vdd.n1622 vdd.n1621 171.744
R17939 vdd.n1621 vdd.n1590 171.744
R17940 vdd.n1614 vdd.n1590 171.744
R17941 vdd.n1614 vdd.n1613 171.744
R17942 vdd.n1613 vdd.n1595 171.744
R17943 vdd.n1606 vdd.n1595 171.744
R17944 vdd.n1606 vdd.n1605 171.744
R17945 vdd.n1605 vdd.n1599 171.744
R17946 vdd.n1682 vdd.n1681 171.744
R17947 vdd.n1681 vdd.n1680 171.744
R17948 vdd.n1680 vdd.n1649 171.744
R17949 vdd.n1673 vdd.n1649 171.744
R17950 vdd.n1673 vdd.n1672 171.744
R17951 vdd.n1672 vdd.n1654 171.744
R17952 vdd.n1665 vdd.n1654 171.744
R17953 vdd.n1665 vdd.n1664 171.744
R17954 vdd.n1664 vdd.n1658 171.744
R17955 vdd.n468 vdd.n467 146.341
R17956 vdd.n474 vdd.n473 146.341
R17957 vdd.n478 vdd.n477 146.341
R17958 vdd.n484 vdd.n483 146.341
R17959 vdd.n488 vdd.n487 146.341
R17960 vdd.n494 vdd.n493 146.341
R17961 vdd.n498 vdd.n497 146.341
R17962 vdd.n504 vdd.n503 146.341
R17963 vdd.n508 vdd.n507 146.341
R17964 vdd.n514 vdd.n513 146.341
R17965 vdd.n518 vdd.n517 146.341
R17966 vdd.n524 vdd.n523 146.341
R17967 vdd.n528 vdd.n527 146.341
R17968 vdd.n534 vdd.n533 146.341
R17969 vdd.n538 vdd.n537 146.341
R17970 vdd.n544 vdd.n543 146.341
R17971 vdd.n548 vdd.n547 146.341
R17972 vdd.n554 vdd.n553 146.341
R17973 vdd.n558 vdd.n557 146.341
R17974 vdd.n564 vdd.n563 146.341
R17975 vdd.n568 vdd.n567 146.341
R17976 vdd.n574 vdd.n573 146.341
R17977 vdd.n578 vdd.n577 146.341
R17978 vdd.n584 vdd.n583 146.341
R17979 vdd.n588 vdd.n587 146.341
R17980 vdd.n594 vdd.n593 146.341
R17981 vdd.n598 vdd.n597 146.341
R17982 vdd.n604 vdd.n603 146.341
R17983 vdd.n608 vdd.n607 146.341
R17984 vdd.n614 vdd.n613 146.341
R17985 vdd.n616 vdd.n425 146.341
R17986 vdd.n3412 vdd.n685 146.341
R17987 vdd.n3412 vdd.n677 146.341
R17988 vdd.n3422 vdd.n677 146.341
R17989 vdd.n3422 vdd.n673 146.341
R17990 vdd.n3428 vdd.n673 146.341
R17991 vdd.n3428 vdd.n667 146.341
R17992 vdd.n3439 vdd.n667 146.341
R17993 vdd.n3439 vdd.n663 146.341
R17994 vdd.n3445 vdd.n663 146.341
R17995 vdd.n3445 vdd.n654 146.341
R17996 vdd.n3455 vdd.n654 146.341
R17997 vdd.n3455 vdd.n650 146.341
R17998 vdd.n3461 vdd.n650 146.341
R17999 vdd.n3461 vdd.n643 146.341
R18000 vdd.n3472 vdd.n643 146.341
R18001 vdd.n3472 vdd.n639 146.341
R18002 vdd.n3481 vdd.n639 146.341
R18003 vdd.n3481 vdd.n632 146.341
R18004 vdd.n3491 vdd.n632 146.341
R18005 vdd.n3492 vdd.n3491 146.341
R18006 vdd.n3492 vdd.n341 146.341
R18007 vdd.n342 vdd.n341 146.341
R18008 vdd.n343 vdd.n342 146.341
R18009 vdd.n3499 vdd.n343 146.341
R18010 vdd.n3499 vdd.n351 146.341
R18011 vdd.n352 vdd.n351 146.341
R18012 vdd.n353 vdd.n352 146.341
R18013 vdd.n3506 vdd.n353 146.341
R18014 vdd.n3506 vdd.n362 146.341
R18015 vdd.n363 vdd.n362 146.341
R18016 vdd.n364 vdd.n363 146.341
R18017 vdd.n3514 vdd.n364 146.341
R18018 vdd.n3514 vdd.n372 146.341
R18019 vdd.n373 vdd.n372 146.341
R18020 vdd.n374 vdd.n373 146.341
R18021 vdd.n3521 vdd.n374 146.341
R18022 vdd.n3521 vdd.n383 146.341
R18023 vdd.n384 vdd.n383 146.341
R18024 vdd.n385 vdd.n384 146.341
R18025 vdd.n3528 vdd.n385 146.341
R18026 vdd.n3528 vdd.n393 146.341
R18027 vdd.n725 vdd.n724 146.341
R18028 vdd.n728 vdd.n724 146.341
R18029 vdd.n734 vdd.n733 146.341
R18030 vdd.n3394 vdd.n3393 146.341
R18031 vdd.n3390 vdd.n3389 146.341
R18032 vdd.n3386 vdd.n3385 146.341
R18033 vdd.n3382 vdd.n3381 146.341
R18034 vdd.n3378 vdd.n3377 146.341
R18035 vdd.n3374 vdd.n3373 146.341
R18036 vdd.n3370 vdd.n3369 146.341
R18037 vdd.n3361 vdd.n3360 146.341
R18038 vdd.n3358 vdd.n3357 146.341
R18039 vdd.n3354 vdd.n3353 146.341
R18040 vdd.n3350 vdd.n3349 146.341
R18041 vdd.n3346 vdd.n3345 146.341
R18042 vdd.n3342 vdd.n3341 146.341
R18043 vdd.n3338 vdd.n3337 146.341
R18044 vdd.n3334 vdd.n3333 146.341
R18045 vdd.n3330 vdd.n3329 146.341
R18046 vdd.n3326 vdd.n3325 146.341
R18047 vdd.n3322 vdd.n3321 146.341
R18048 vdd.n3315 vdd.n3314 146.341
R18049 vdd.n3312 vdd.n3311 146.341
R18050 vdd.n3308 vdd.n3307 146.341
R18051 vdd.n3304 vdd.n3303 146.341
R18052 vdd.n3300 vdd.n3299 146.341
R18053 vdd.n3296 vdd.n3295 146.341
R18054 vdd.n3292 vdd.n3291 146.341
R18055 vdd.n3288 vdd.n3287 146.341
R18056 vdd.n3284 vdd.n3283 146.341
R18057 vdd.n3280 vdd.n3279 146.341
R18058 vdd.n3406 vdd.n691 146.341
R18059 vdd.n3414 vdd.n684 146.341
R18060 vdd.n3414 vdd.n680 146.341
R18061 vdd.n3420 vdd.n680 146.341
R18062 vdd.n3420 vdd.n672 146.341
R18063 vdd.n3431 vdd.n672 146.341
R18064 vdd.n3431 vdd.n668 146.341
R18065 vdd.n3437 vdd.n668 146.341
R18066 vdd.n3437 vdd.n661 146.341
R18067 vdd.n3447 vdd.n661 146.341
R18068 vdd.n3447 vdd.n657 146.341
R18069 vdd.n3453 vdd.n657 146.341
R18070 vdd.n3453 vdd.n649 146.341
R18071 vdd.n3464 vdd.n649 146.341
R18072 vdd.n3464 vdd.n645 146.341
R18073 vdd.n3470 vdd.n645 146.341
R18074 vdd.n3470 vdd.n638 146.341
R18075 vdd.n3483 vdd.n638 146.341
R18076 vdd.n3483 vdd.n634 146.341
R18077 vdd.n3489 vdd.n634 146.341
R18078 vdd.n3489 vdd.n338 146.341
R18079 vdd.n3578 vdd.n338 146.341
R18080 vdd.n3578 vdd.n339 146.341
R18081 vdd.n3574 vdd.n339 146.341
R18082 vdd.n3574 vdd.n345 146.341
R18083 vdd.n3570 vdd.n345 146.341
R18084 vdd.n3570 vdd.n350 146.341
R18085 vdd.n3566 vdd.n350 146.341
R18086 vdd.n3566 vdd.n354 146.341
R18087 vdd.n3562 vdd.n354 146.341
R18088 vdd.n3562 vdd.n360 146.341
R18089 vdd.n3558 vdd.n360 146.341
R18090 vdd.n3558 vdd.n365 146.341
R18091 vdd.n3554 vdd.n365 146.341
R18092 vdd.n3554 vdd.n371 146.341
R18093 vdd.n3550 vdd.n371 146.341
R18094 vdd.n3550 vdd.n376 146.341
R18095 vdd.n3546 vdd.n376 146.341
R18096 vdd.n3546 vdd.n382 146.341
R18097 vdd.n3542 vdd.n382 146.341
R18098 vdd.n3542 vdd.n387 146.341
R18099 vdd.n3538 vdd.n387 146.341
R18100 vdd.n2189 vdd.n2188 146.341
R18101 vdd.n2186 vdd.n1983 146.341
R18102 vdd.n2179 vdd.n1989 146.341
R18103 vdd.n2177 vdd.n2176 146.341
R18104 vdd.n2174 vdd.n1991 146.341
R18105 vdd.n2170 vdd.n2169 146.341
R18106 vdd.n2167 vdd.n1998 146.341
R18107 vdd.n2163 vdd.n2162 146.341
R18108 vdd.n2160 vdd.n2005 146.341
R18109 vdd.n2016 vdd.n2013 146.341
R18110 vdd.n2152 vdd.n2151 146.341
R18111 vdd.n2149 vdd.n2018 146.341
R18112 vdd.n2145 vdd.n2144 146.341
R18113 vdd.n2142 vdd.n2024 146.341
R18114 vdd.n2138 vdd.n2137 146.341
R18115 vdd.n2135 vdd.n2031 146.341
R18116 vdd.n2131 vdd.n2130 146.341
R18117 vdd.n2128 vdd.n2038 146.341
R18118 vdd.n2124 vdd.n2123 146.341
R18119 vdd.n2121 vdd.n2045 146.341
R18120 vdd.n2056 vdd.n2053 146.341
R18121 vdd.n2113 vdd.n2112 146.341
R18122 vdd.n2110 vdd.n2058 146.341
R18123 vdd.n2106 vdd.n2105 146.341
R18124 vdd.n2103 vdd.n2064 146.341
R18125 vdd.n2099 vdd.n2098 146.341
R18126 vdd.n2096 vdd.n2071 146.341
R18127 vdd.n2092 vdd.n2091 146.341
R18128 vdd.n2089 vdd.n2086 146.341
R18129 vdd.n2084 vdd.n2081 146.341
R18130 vdd.n2079 vdd.n1149 146.341
R18131 vdd.n1508 vdd.n1268 146.341
R18132 vdd.n1508 vdd.n1264 146.341
R18133 vdd.n1514 vdd.n1264 146.341
R18134 vdd.n1514 vdd.n1256 146.341
R18135 vdd.n1525 vdd.n1256 146.341
R18136 vdd.n1525 vdd.n1252 146.341
R18137 vdd.n1531 vdd.n1252 146.341
R18138 vdd.n1531 vdd.n1246 146.341
R18139 vdd.n1542 vdd.n1246 146.341
R18140 vdd.n1542 vdd.n1242 146.341
R18141 vdd.n1548 vdd.n1242 146.341
R18142 vdd.n1548 vdd.n1233 146.341
R18143 vdd.n1558 vdd.n1233 146.341
R18144 vdd.n1558 vdd.n1229 146.341
R18145 vdd.n1564 vdd.n1229 146.341
R18146 vdd.n1564 vdd.n1222 146.341
R18147 vdd.n1575 vdd.n1222 146.341
R18148 vdd.n1575 vdd.n1218 146.341
R18149 vdd.n1581 vdd.n1218 146.341
R18150 vdd.n1581 vdd.n1211 146.341
R18151 vdd.n1898 vdd.n1211 146.341
R18152 vdd.n1898 vdd.n1207 146.341
R18153 vdd.n1904 vdd.n1207 146.341
R18154 vdd.n1904 vdd.n1199 146.341
R18155 vdd.n1915 vdd.n1199 146.341
R18156 vdd.n1915 vdd.n1195 146.341
R18157 vdd.n1921 vdd.n1195 146.341
R18158 vdd.n1921 vdd.n1189 146.341
R18159 vdd.n1932 vdd.n1189 146.341
R18160 vdd.n1932 vdd.n1185 146.341
R18161 vdd.n1938 vdd.n1185 146.341
R18162 vdd.n1938 vdd.n1176 146.341
R18163 vdd.n1948 vdd.n1176 146.341
R18164 vdd.n1948 vdd.n1172 146.341
R18165 vdd.n1954 vdd.n1172 146.341
R18166 vdd.n1954 vdd.n1166 146.341
R18167 vdd.n1965 vdd.n1166 146.341
R18168 vdd.n1965 vdd.n1161 146.341
R18169 vdd.n1973 vdd.n1161 146.341
R18170 vdd.n1973 vdd.n1151 146.341
R18171 vdd.n2197 vdd.n1151 146.341
R18172 vdd.n1497 vdd.n1273 146.341
R18173 vdd.n1497 vdd.n1306 146.341
R18174 vdd.n1310 vdd.n1309 146.341
R18175 vdd.n1312 vdd.n1311 146.341
R18176 vdd.n1316 vdd.n1315 146.341
R18177 vdd.n1318 vdd.n1317 146.341
R18178 vdd.n1322 vdd.n1321 146.341
R18179 vdd.n1324 vdd.n1323 146.341
R18180 vdd.n1328 vdd.n1327 146.341
R18181 vdd.n1330 vdd.n1329 146.341
R18182 vdd.n1336 vdd.n1335 146.341
R18183 vdd.n1338 vdd.n1337 146.341
R18184 vdd.n1342 vdd.n1341 146.341
R18185 vdd.n1344 vdd.n1343 146.341
R18186 vdd.n1348 vdd.n1347 146.341
R18187 vdd.n1350 vdd.n1349 146.341
R18188 vdd.n1354 vdd.n1353 146.341
R18189 vdd.n1356 vdd.n1355 146.341
R18190 vdd.n1360 vdd.n1359 146.341
R18191 vdd.n1362 vdd.n1361 146.341
R18192 vdd.n1434 vdd.n1365 146.341
R18193 vdd.n1367 vdd.n1366 146.341
R18194 vdd.n1371 vdd.n1370 146.341
R18195 vdd.n1373 vdd.n1372 146.341
R18196 vdd.n1377 vdd.n1376 146.341
R18197 vdd.n1379 vdd.n1378 146.341
R18198 vdd.n1383 vdd.n1382 146.341
R18199 vdd.n1385 vdd.n1384 146.341
R18200 vdd.n1389 vdd.n1388 146.341
R18201 vdd.n1391 vdd.n1390 146.341
R18202 vdd.n1395 vdd.n1394 146.341
R18203 vdd.n1396 vdd.n1304 146.341
R18204 vdd.n1506 vdd.n1269 146.341
R18205 vdd.n1506 vdd.n1262 146.341
R18206 vdd.n1517 vdd.n1262 146.341
R18207 vdd.n1517 vdd.n1258 146.341
R18208 vdd.n1523 vdd.n1258 146.341
R18209 vdd.n1523 vdd.n1251 146.341
R18210 vdd.n1534 vdd.n1251 146.341
R18211 vdd.n1534 vdd.n1247 146.341
R18212 vdd.n1540 vdd.n1247 146.341
R18213 vdd.n1540 vdd.n1240 146.341
R18214 vdd.n1550 vdd.n1240 146.341
R18215 vdd.n1550 vdd.n1236 146.341
R18216 vdd.n1556 vdd.n1236 146.341
R18217 vdd.n1556 vdd.n1228 146.341
R18218 vdd.n1567 vdd.n1228 146.341
R18219 vdd.n1567 vdd.n1224 146.341
R18220 vdd.n1573 vdd.n1224 146.341
R18221 vdd.n1573 vdd.n1217 146.341
R18222 vdd.n1583 vdd.n1217 146.341
R18223 vdd.n1583 vdd.n1213 146.341
R18224 vdd.n1896 vdd.n1213 146.341
R18225 vdd.n1896 vdd.n1205 146.341
R18226 vdd.n1907 vdd.n1205 146.341
R18227 vdd.n1907 vdd.n1201 146.341
R18228 vdd.n1913 vdd.n1201 146.341
R18229 vdd.n1913 vdd.n1194 146.341
R18230 vdd.n1924 vdd.n1194 146.341
R18231 vdd.n1924 vdd.n1190 146.341
R18232 vdd.n1930 vdd.n1190 146.341
R18233 vdd.n1930 vdd.n1183 146.341
R18234 vdd.n1940 vdd.n1183 146.341
R18235 vdd.n1940 vdd.n1179 146.341
R18236 vdd.n1946 vdd.n1179 146.341
R18237 vdd.n1946 vdd.n1171 146.341
R18238 vdd.n1957 vdd.n1171 146.341
R18239 vdd.n1957 vdd.n1167 146.341
R18240 vdd.n1963 vdd.n1167 146.341
R18241 vdd.n1963 vdd.n1159 146.341
R18242 vdd.n1976 vdd.n1159 146.341
R18243 vdd.n1976 vdd.n1154 146.341
R18244 vdd.n2195 vdd.n1154 146.341
R18245 vdd.n1136 vdd.t68 127.284
R18246 vdd.n997 vdd.t105 127.284
R18247 vdd.n1130 vdd.t132 127.284
R18248 vdd.n988 vdd.t128 127.284
R18249 vdd.n885 vdd.t78 127.284
R18250 vdd.n885 vdd.t79 127.284
R18251 vdd.n2761 vdd.t123 127.284
R18252 vdd.n832 vdd.t91 127.284
R18253 vdd.n2830 vdd.t110 127.284
R18254 vdd.n799 vdd.t63 127.284
R18255 vdd.n1058 vdd.t119 127.284
R18256 vdd.n1058 vdd.t120 127.284
R18257 vdd.n22 vdd.n20 117.314
R18258 vdd.n17 vdd.n15 117.314
R18259 vdd.n27 vdd.n26 116.927
R18260 vdd.n24 vdd.n23 116.927
R18261 vdd.n22 vdd.n21 116.927
R18262 vdd.n17 vdd.n16 116.927
R18263 vdd.n19 vdd.n18 116.927
R18264 vdd.n27 vdd.n25 116.927
R18265 vdd.n1137 vdd.t67 111.188
R18266 vdd.n998 vdd.t106 111.188
R18267 vdd.n1131 vdd.t131 111.188
R18268 vdd.n989 vdd.t129 111.188
R18269 vdd.n2762 vdd.t122 111.188
R18270 vdd.n833 vdd.t92 111.188
R18271 vdd.n2831 vdd.t109 111.188
R18272 vdd.n800 vdd.t64 111.188
R18273 vdd.n3016 vdd.n938 99.5127
R18274 vdd.n3024 vdd.n938 99.5127
R18275 vdd.n3024 vdd.n936 99.5127
R18276 vdd.n3028 vdd.n936 99.5127
R18277 vdd.n3028 vdd.n926 99.5127
R18278 vdd.n3036 vdd.n926 99.5127
R18279 vdd.n3036 vdd.n924 99.5127
R18280 vdd.n3040 vdd.n924 99.5127
R18281 vdd.n3040 vdd.n916 99.5127
R18282 vdd.n3048 vdd.n916 99.5127
R18283 vdd.n3048 vdd.n914 99.5127
R18284 vdd.n3052 vdd.n914 99.5127
R18285 vdd.n3052 vdd.n904 99.5127
R18286 vdd.n3060 vdd.n904 99.5127
R18287 vdd.n3060 vdd.n902 99.5127
R18288 vdd.n3064 vdd.n902 99.5127
R18289 vdd.n3064 vdd.n893 99.5127
R18290 vdd.n3072 vdd.n893 99.5127
R18291 vdd.n3072 vdd.n891 99.5127
R18292 vdd.n3076 vdd.n891 99.5127
R18293 vdd.n3076 vdd.n880 99.5127
R18294 vdd.n3085 vdd.n880 99.5127
R18295 vdd.n3085 vdd.n878 99.5127
R18296 vdd.n3089 vdd.n878 99.5127
R18297 vdd.n3089 vdd.n867 99.5127
R18298 vdd.n3097 vdd.n867 99.5127
R18299 vdd.n3097 vdd.n865 99.5127
R18300 vdd.n3101 vdd.n865 99.5127
R18301 vdd.n3101 vdd.n856 99.5127
R18302 vdd.n3109 vdd.n856 99.5127
R18303 vdd.n3109 vdd.n854 99.5127
R18304 vdd.n3113 vdd.n854 99.5127
R18305 vdd.n3113 vdd.n842 99.5127
R18306 vdd.n3166 vdd.n842 99.5127
R18307 vdd.n3166 vdd.n840 99.5127
R18308 vdd.n3170 vdd.n840 99.5127
R18309 vdd.n3170 vdd.n808 99.5127
R18310 vdd.n3240 vdd.n808 99.5127
R18311 vdd.n3236 vdd.n809 99.5127
R18312 vdd.n3234 vdd.n3233 99.5127
R18313 vdd.n3231 vdd.n813 99.5127
R18314 vdd.n3227 vdd.n3226 99.5127
R18315 vdd.n3224 vdd.n816 99.5127
R18316 vdd.n3220 vdd.n3219 99.5127
R18317 vdd.n3217 vdd.n819 99.5127
R18318 vdd.n3213 vdd.n3212 99.5127
R18319 vdd.n3210 vdd.n3208 99.5127
R18320 vdd.n3206 vdd.n822 99.5127
R18321 vdd.n3202 vdd.n3201 99.5127
R18322 vdd.n3199 vdd.n825 99.5127
R18323 vdd.n3195 vdd.n3194 99.5127
R18324 vdd.n3192 vdd.n828 99.5127
R18325 vdd.n3188 vdd.n3187 99.5127
R18326 vdd.n3185 vdd.n831 99.5127
R18327 vdd.n3180 vdd.n3179 99.5127
R18328 vdd.n2898 vdd.n944 99.5127
R18329 vdd.n2898 vdd.n939 99.5127
R18330 vdd.n3000 vdd.n939 99.5127
R18331 vdd.n3000 vdd.n934 99.5127
R18332 vdd.n2996 vdd.n934 99.5127
R18333 vdd.n2996 vdd.n928 99.5127
R18334 vdd.n2993 vdd.n928 99.5127
R18335 vdd.n2993 vdd.n922 99.5127
R18336 vdd.n2990 vdd.n922 99.5127
R18337 vdd.n2990 vdd.n917 99.5127
R18338 vdd.n2940 vdd.n917 99.5127
R18339 vdd.n2940 vdd.n912 99.5127
R18340 vdd.n2943 vdd.n912 99.5127
R18341 vdd.n2943 vdd.n906 99.5127
R18342 vdd.n2976 vdd.n906 99.5127
R18343 vdd.n2976 vdd.n899 99.5127
R18344 vdd.n2972 vdd.n899 99.5127
R18345 vdd.n2972 vdd.n894 99.5127
R18346 vdd.n2969 vdd.n894 99.5127
R18347 vdd.n2969 vdd.n889 99.5127
R18348 vdd.n2966 vdd.n889 99.5127
R18349 vdd.n2966 vdd.n882 99.5127
R18350 vdd.n2963 vdd.n882 99.5127
R18351 vdd.n2963 vdd.n875 99.5127
R18352 vdd.n2960 vdd.n875 99.5127
R18353 vdd.n2960 vdd.n868 99.5127
R18354 vdd.n2957 vdd.n868 99.5127
R18355 vdd.n2957 vdd.n862 99.5127
R18356 vdd.n2954 vdd.n862 99.5127
R18357 vdd.n2954 vdd.n857 99.5127
R18358 vdd.n2951 vdd.n857 99.5127
R18359 vdd.n2951 vdd.n852 99.5127
R18360 vdd.n2948 vdd.n852 99.5127
R18361 vdd.n2948 vdd.n844 99.5127
R18362 vdd.n844 vdd.n837 99.5127
R18363 vdd.n3172 vdd.n837 99.5127
R18364 vdd.n3173 vdd.n3172 99.5127
R18365 vdd.n3173 vdd.n806 99.5127
R18366 vdd.n3012 vdd.n949 99.5127
R18367 vdd.n2832 vdd.n949 99.5127
R18368 vdd.n2836 vdd.n2835 99.5127
R18369 vdd.n2840 vdd.n2839 99.5127
R18370 vdd.n2844 vdd.n2843 99.5127
R18371 vdd.n2848 vdd.n2847 99.5127
R18372 vdd.n2852 vdd.n2851 99.5127
R18373 vdd.n2856 vdd.n2855 99.5127
R18374 vdd.n2860 vdd.n2859 99.5127
R18375 vdd.n2864 vdd.n2863 99.5127
R18376 vdd.n2868 vdd.n2867 99.5127
R18377 vdd.n2872 vdd.n2871 99.5127
R18378 vdd.n2876 vdd.n2875 99.5127
R18379 vdd.n2880 vdd.n2879 99.5127
R18380 vdd.n2884 vdd.n2883 99.5127
R18381 vdd.n2888 vdd.n2887 99.5127
R18382 vdd.n2893 vdd.n2892 99.5127
R18383 vdd.n2725 vdd.n986 99.5127
R18384 vdd.n2721 vdd.n2720 99.5127
R18385 vdd.n2717 vdd.n2716 99.5127
R18386 vdd.n2713 vdd.n2712 99.5127
R18387 vdd.n2709 vdd.n2708 99.5127
R18388 vdd.n2705 vdd.n2704 99.5127
R18389 vdd.n2701 vdd.n2700 99.5127
R18390 vdd.n2697 vdd.n2696 99.5127
R18391 vdd.n2693 vdd.n2692 99.5127
R18392 vdd.n2689 vdd.n2688 99.5127
R18393 vdd.n2685 vdd.n2684 99.5127
R18394 vdd.n2681 vdd.n2680 99.5127
R18395 vdd.n2677 vdd.n2676 99.5127
R18396 vdd.n2673 vdd.n2672 99.5127
R18397 vdd.n2669 vdd.n2668 99.5127
R18398 vdd.n2665 vdd.n2664 99.5127
R18399 vdd.n2660 vdd.n2659 99.5127
R18400 vdd.n2392 vdd.n1111 99.5127
R18401 vdd.n2392 vdd.n1105 99.5127
R18402 vdd.n2389 vdd.n1105 99.5127
R18403 vdd.n2389 vdd.n1099 99.5127
R18404 vdd.n2386 vdd.n1099 99.5127
R18405 vdd.n2386 vdd.n1093 99.5127
R18406 vdd.n2383 vdd.n1093 99.5127
R18407 vdd.n2383 vdd.n1087 99.5127
R18408 vdd.n2380 vdd.n1087 99.5127
R18409 vdd.n2380 vdd.n1081 99.5127
R18410 vdd.n2377 vdd.n1081 99.5127
R18411 vdd.n2377 vdd.n1075 99.5127
R18412 vdd.n2374 vdd.n1075 99.5127
R18413 vdd.n2374 vdd.n1068 99.5127
R18414 vdd.n2371 vdd.n1068 99.5127
R18415 vdd.n2371 vdd.n1061 99.5127
R18416 vdd.n2368 vdd.n1061 99.5127
R18417 vdd.n2368 vdd.n1055 99.5127
R18418 vdd.n2365 vdd.n1055 99.5127
R18419 vdd.n2365 vdd.n1050 99.5127
R18420 vdd.n2362 vdd.n1050 99.5127
R18421 vdd.n2362 vdd.n1044 99.5127
R18422 vdd.n2359 vdd.n1044 99.5127
R18423 vdd.n2359 vdd.n1037 99.5127
R18424 vdd.n2326 vdd.n1037 99.5127
R18425 vdd.n2326 vdd.n1031 99.5127
R18426 vdd.n2329 vdd.n1031 99.5127
R18427 vdd.n2329 vdd.n1026 99.5127
R18428 vdd.n2345 vdd.n1026 99.5127
R18429 vdd.n2345 vdd.n1021 99.5127
R18430 vdd.n2341 vdd.n1021 99.5127
R18431 vdd.n2341 vdd.n1016 99.5127
R18432 vdd.n2338 vdd.n1016 99.5127
R18433 vdd.n2338 vdd.n1009 99.5127
R18434 vdd.n2335 vdd.n1009 99.5127
R18435 vdd.n2335 vdd.n1002 99.5127
R18436 vdd.n1002 vdd.n991 99.5127
R18437 vdd.n2655 vdd.n991 99.5127
R18438 vdd.n2462 vdd.n2460 99.5127
R18439 vdd.n2460 vdd.n2459 99.5127
R18440 vdd.n2456 vdd.n2455 99.5127
R18441 vdd.n2453 vdd.n1117 99.5127
R18442 vdd.n2449 vdd.n2447 99.5127
R18443 vdd.n2445 vdd.n1119 99.5127
R18444 vdd.n2441 vdd.n2439 99.5127
R18445 vdd.n2437 vdd.n1121 99.5127
R18446 vdd.n2433 vdd.n2431 99.5127
R18447 vdd.n2429 vdd.n1123 99.5127
R18448 vdd.n2425 vdd.n2423 99.5127
R18449 vdd.n2421 vdd.n1125 99.5127
R18450 vdd.n2417 vdd.n2415 99.5127
R18451 vdd.n2413 vdd.n1127 99.5127
R18452 vdd.n2409 vdd.n2407 99.5127
R18453 vdd.n2405 vdd.n1129 99.5127
R18454 vdd.n2400 vdd.n2398 99.5127
R18455 vdd.n2466 vdd.n1103 99.5127
R18456 vdd.n2474 vdd.n1103 99.5127
R18457 vdd.n2474 vdd.n1101 99.5127
R18458 vdd.n2478 vdd.n1101 99.5127
R18459 vdd.n2478 vdd.n1091 99.5127
R18460 vdd.n2486 vdd.n1091 99.5127
R18461 vdd.n2486 vdd.n1089 99.5127
R18462 vdd.n2490 vdd.n1089 99.5127
R18463 vdd.n2490 vdd.n1079 99.5127
R18464 vdd.n2498 vdd.n1079 99.5127
R18465 vdd.n2498 vdd.n1077 99.5127
R18466 vdd.n2502 vdd.n1077 99.5127
R18467 vdd.n2502 vdd.n1066 99.5127
R18468 vdd.n2510 vdd.n1066 99.5127
R18469 vdd.n2510 vdd.n1064 99.5127
R18470 vdd.n2514 vdd.n1064 99.5127
R18471 vdd.n2514 vdd.n1054 99.5127
R18472 vdd.n2523 vdd.n1054 99.5127
R18473 vdd.n2523 vdd.n1052 99.5127
R18474 vdd.n2527 vdd.n1052 99.5127
R18475 vdd.n2527 vdd.n1042 99.5127
R18476 vdd.n2535 vdd.n1042 99.5127
R18477 vdd.n2535 vdd.n1040 99.5127
R18478 vdd.n2539 vdd.n1040 99.5127
R18479 vdd.n2539 vdd.n1030 99.5127
R18480 vdd.n2547 vdd.n1030 99.5127
R18481 vdd.n2547 vdd.n1028 99.5127
R18482 vdd.n2551 vdd.n1028 99.5127
R18483 vdd.n2551 vdd.n1020 99.5127
R18484 vdd.n2559 vdd.n1020 99.5127
R18485 vdd.n2559 vdd.n1018 99.5127
R18486 vdd.n2563 vdd.n1018 99.5127
R18487 vdd.n2563 vdd.n1007 99.5127
R18488 vdd.n2573 vdd.n1007 99.5127
R18489 vdd.n2573 vdd.n1004 99.5127
R18490 vdd.n2578 vdd.n1004 99.5127
R18491 vdd.n2578 vdd.n1005 99.5127
R18492 vdd.n1005 vdd.n985 99.5127
R18493 vdd.n3156 vdd.n3155 99.5127
R18494 vdd.n3153 vdd.n3119 99.5127
R18495 vdd.n3149 vdd.n3148 99.5127
R18496 vdd.n3146 vdd.n3122 99.5127
R18497 vdd.n3142 vdd.n3141 99.5127
R18498 vdd.n3139 vdd.n3125 99.5127
R18499 vdd.n3135 vdd.n3134 99.5127
R18500 vdd.n3132 vdd.n3129 99.5127
R18501 vdd.n3273 vdd.n787 99.5127
R18502 vdd.n3271 vdd.n3270 99.5127
R18503 vdd.n3268 vdd.n789 99.5127
R18504 vdd.n3264 vdd.n3263 99.5127
R18505 vdd.n3261 vdd.n792 99.5127
R18506 vdd.n3257 vdd.n3256 99.5127
R18507 vdd.n3254 vdd.n795 99.5127
R18508 vdd.n3250 vdd.n3249 99.5127
R18509 vdd.n3247 vdd.n798 99.5127
R18510 vdd.n3005 vdd.n945 99.5127
R18511 vdd.n3005 vdd.n940 99.5127
R18512 vdd.n3002 vdd.n940 99.5127
R18513 vdd.n3002 vdd.n935 99.5127
R18514 vdd.n2902 vdd.n935 99.5127
R18515 vdd.n2902 vdd.n929 99.5127
R18516 vdd.n2905 vdd.n929 99.5127
R18517 vdd.n2905 vdd.n923 99.5127
R18518 vdd.n2988 vdd.n923 99.5127
R18519 vdd.n2988 vdd.n918 99.5127
R18520 vdd.n2984 vdd.n918 99.5127
R18521 vdd.n2984 vdd.n913 99.5127
R18522 vdd.n2981 vdd.n913 99.5127
R18523 vdd.n2981 vdd.n907 99.5127
R18524 vdd.n2978 vdd.n907 99.5127
R18525 vdd.n2978 vdd.n900 99.5127
R18526 vdd.n2937 vdd.n900 99.5127
R18527 vdd.n2937 vdd.n895 99.5127
R18528 vdd.n2934 vdd.n895 99.5127
R18529 vdd.n2934 vdd.n890 99.5127
R18530 vdd.n2931 vdd.n890 99.5127
R18531 vdd.n2931 vdd.n883 99.5127
R18532 vdd.n2928 vdd.n883 99.5127
R18533 vdd.n2928 vdd.n876 99.5127
R18534 vdd.n2925 vdd.n876 99.5127
R18535 vdd.n2925 vdd.n869 99.5127
R18536 vdd.n2922 vdd.n869 99.5127
R18537 vdd.n2922 vdd.n863 99.5127
R18538 vdd.n2919 vdd.n863 99.5127
R18539 vdd.n2919 vdd.n858 99.5127
R18540 vdd.n2916 vdd.n858 99.5127
R18541 vdd.n2916 vdd.n853 99.5127
R18542 vdd.n2913 vdd.n853 99.5127
R18543 vdd.n2913 vdd.n845 99.5127
R18544 vdd.n2910 vdd.n845 99.5127
R18545 vdd.n2910 vdd.n838 99.5127
R18546 vdd.n838 vdd.n804 99.5127
R18547 vdd.n3242 vdd.n804 99.5127
R18548 vdd.n2766 vdd.n2765 99.5127
R18549 vdd.n2770 vdd.n2769 99.5127
R18550 vdd.n2774 vdd.n2773 99.5127
R18551 vdd.n2778 vdd.n2777 99.5127
R18552 vdd.n2782 vdd.n2781 99.5127
R18553 vdd.n2786 vdd.n2785 99.5127
R18554 vdd.n2790 vdd.n2789 99.5127
R18555 vdd.n2794 vdd.n2793 99.5127
R18556 vdd.n2798 vdd.n2797 99.5127
R18557 vdd.n2802 vdd.n2801 99.5127
R18558 vdd.n2806 vdd.n2805 99.5127
R18559 vdd.n2810 vdd.n2809 99.5127
R18560 vdd.n2814 vdd.n2813 99.5127
R18561 vdd.n2818 vdd.n2817 99.5127
R18562 vdd.n2822 vdd.n2821 99.5127
R18563 vdd.n2826 vdd.n2825 99.5127
R18564 vdd.n3009 vdd.n2760 99.5127
R18565 vdd.n3018 vdd.n941 99.5127
R18566 vdd.n3022 vdd.n941 99.5127
R18567 vdd.n3022 vdd.n933 99.5127
R18568 vdd.n3030 vdd.n933 99.5127
R18569 vdd.n3030 vdd.n931 99.5127
R18570 vdd.n3034 vdd.n931 99.5127
R18571 vdd.n3034 vdd.n921 99.5127
R18572 vdd.n3042 vdd.n921 99.5127
R18573 vdd.n3042 vdd.n919 99.5127
R18574 vdd.n3046 vdd.n919 99.5127
R18575 vdd.n3046 vdd.n910 99.5127
R18576 vdd.n3054 vdd.n910 99.5127
R18577 vdd.n3054 vdd.n908 99.5127
R18578 vdd.n3058 vdd.n908 99.5127
R18579 vdd.n3058 vdd.n898 99.5127
R18580 vdd.n3066 vdd.n898 99.5127
R18581 vdd.n3066 vdd.n896 99.5127
R18582 vdd.n3070 vdd.n896 99.5127
R18583 vdd.n3070 vdd.n887 99.5127
R18584 vdd.n3078 vdd.n887 99.5127
R18585 vdd.n3078 vdd.n884 99.5127
R18586 vdd.n3083 vdd.n884 99.5127
R18587 vdd.n3083 vdd.n873 99.5127
R18588 vdd.n3091 vdd.n873 99.5127
R18589 vdd.n3091 vdd.n871 99.5127
R18590 vdd.n3095 vdd.n871 99.5127
R18591 vdd.n3095 vdd.n861 99.5127
R18592 vdd.n3103 vdd.n861 99.5127
R18593 vdd.n3103 vdd.n859 99.5127
R18594 vdd.n3107 vdd.n859 99.5127
R18595 vdd.n3107 vdd.n850 99.5127
R18596 vdd.n3115 vdd.n850 99.5127
R18597 vdd.n3115 vdd.n847 99.5127
R18598 vdd.n3164 vdd.n847 99.5127
R18599 vdd.n3164 vdd.n848 99.5127
R18600 vdd.n848 vdd.n839 99.5127
R18601 vdd.n3159 vdd.n839 99.5127
R18602 vdd.n3159 vdd.n807 99.5127
R18603 vdd.n2649 vdd.n2648 99.5127
R18604 vdd.n2645 vdd.n2644 99.5127
R18605 vdd.n2641 vdd.n2640 99.5127
R18606 vdd.n2637 vdd.n2636 99.5127
R18607 vdd.n2633 vdd.n2632 99.5127
R18608 vdd.n2629 vdd.n2628 99.5127
R18609 vdd.n2625 vdd.n2624 99.5127
R18610 vdd.n2621 vdd.n2620 99.5127
R18611 vdd.n2617 vdd.n2616 99.5127
R18612 vdd.n2613 vdd.n2612 99.5127
R18613 vdd.n2609 vdd.n2608 99.5127
R18614 vdd.n2605 vdd.n2604 99.5127
R18615 vdd.n2601 vdd.n2600 99.5127
R18616 vdd.n2597 vdd.n2596 99.5127
R18617 vdd.n2593 vdd.n2592 99.5127
R18618 vdd.n2589 vdd.n2588 99.5127
R18619 vdd.n2585 vdd.n967 99.5127
R18620 vdd.n2285 vdd.n1112 99.5127
R18621 vdd.n2285 vdd.n1106 99.5127
R18622 vdd.n2288 vdd.n1106 99.5127
R18623 vdd.n2288 vdd.n1100 99.5127
R18624 vdd.n2291 vdd.n1100 99.5127
R18625 vdd.n2291 vdd.n1094 99.5127
R18626 vdd.n2294 vdd.n1094 99.5127
R18627 vdd.n2294 vdd.n1088 99.5127
R18628 vdd.n2297 vdd.n1088 99.5127
R18629 vdd.n2297 vdd.n1082 99.5127
R18630 vdd.n2300 vdd.n1082 99.5127
R18631 vdd.n2300 vdd.n1076 99.5127
R18632 vdd.n2303 vdd.n1076 99.5127
R18633 vdd.n2303 vdd.n1069 99.5127
R18634 vdd.n2306 vdd.n1069 99.5127
R18635 vdd.n2306 vdd.n1062 99.5127
R18636 vdd.n2309 vdd.n1062 99.5127
R18637 vdd.n2309 vdd.n1056 99.5127
R18638 vdd.n2312 vdd.n1056 99.5127
R18639 vdd.n2312 vdd.n1051 99.5127
R18640 vdd.n2315 vdd.n1051 99.5127
R18641 vdd.n2315 vdd.n1045 99.5127
R18642 vdd.n2357 vdd.n1045 99.5127
R18643 vdd.n2357 vdd.n1038 99.5127
R18644 vdd.n2353 vdd.n1038 99.5127
R18645 vdd.n2353 vdd.n1032 99.5127
R18646 vdd.n2350 vdd.n1032 99.5127
R18647 vdd.n2350 vdd.n1027 99.5127
R18648 vdd.n2347 vdd.n1027 99.5127
R18649 vdd.n2347 vdd.n1022 99.5127
R18650 vdd.n2323 vdd.n1022 99.5127
R18651 vdd.n2323 vdd.n1017 99.5127
R18652 vdd.n2320 vdd.n1017 99.5127
R18653 vdd.n2320 vdd.n1010 99.5127
R18654 vdd.n1010 vdd.n1001 99.5127
R18655 vdd.n2580 vdd.n1001 99.5127
R18656 vdd.n2581 vdd.n2580 99.5127
R18657 vdd.n2581 vdd.n993 99.5127
R18658 vdd.n2218 vdd.n2216 99.5127
R18659 vdd.n2222 vdd.n2213 99.5127
R18660 vdd.n2226 vdd.n2224 99.5127
R18661 vdd.n2230 vdd.n2211 99.5127
R18662 vdd.n2234 vdd.n2232 99.5127
R18663 vdd.n2238 vdd.n2209 99.5127
R18664 vdd.n2242 vdd.n2240 99.5127
R18665 vdd.n2246 vdd.n2207 99.5127
R18666 vdd.n2250 vdd.n2248 99.5127
R18667 vdd.n2254 vdd.n1143 99.5127
R18668 vdd.n2258 vdd.n2256 99.5127
R18669 vdd.n2262 vdd.n1141 99.5127
R18670 vdd.n2266 vdd.n2264 99.5127
R18671 vdd.n2270 vdd.n1139 99.5127
R18672 vdd.n2274 vdd.n2272 99.5127
R18673 vdd.n2279 vdd.n1135 99.5127
R18674 vdd.n2282 vdd.n2281 99.5127
R18675 vdd.n2468 vdd.n1107 99.5127
R18676 vdd.n2472 vdd.n1107 99.5127
R18677 vdd.n2472 vdd.n1097 99.5127
R18678 vdd.n2480 vdd.n1097 99.5127
R18679 vdd.n2480 vdd.n1095 99.5127
R18680 vdd.n2484 vdd.n1095 99.5127
R18681 vdd.n2484 vdd.n1085 99.5127
R18682 vdd.n2492 vdd.n1085 99.5127
R18683 vdd.n2492 vdd.n1083 99.5127
R18684 vdd.n2496 vdd.n1083 99.5127
R18685 vdd.n2496 vdd.n1073 99.5127
R18686 vdd.n2504 vdd.n1073 99.5127
R18687 vdd.n2504 vdd.n1071 99.5127
R18688 vdd.n2508 vdd.n1071 99.5127
R18689 vdd.n2508 vdd.n1060 99.5127
R18690 vdd.n2516 vdd.n1060 99.5127
R18691 vdd.n2516 vdd.n1057 99.5127
R18692 vdd.n2521 vdd.n1057 99.5127
R18693 vdd.n2521 vdd.n1048 99.5127
R18694 vdd.n2529 vdd.n1048 99.5127
R18695 vdd.n2529 vdd.n1046 99.5127
R18696 vdd.n2533 vdd.n1046 99.5127
R18697 vdd.n2533 vdd.n1036 99.5127
R18698 vdd.n2541 vdd.n1036 99.5127
R18699 vdd.n2541 vdd.n1034 99.5127
R18700 vdd.n2545 vdd.n1034 99.5127
R18701 vdd.n2545 vdd.n1025 99.5127
R18702 vdd.n2553 vdd.n1025 99.5127
R18703 vdd.n2553 vdd.n1023 99.5127
R18704 vdd.n2557 vdd.n1023 99.5127
R18705 vdd.n2557 vdd.n1014 99.5127
R18706 vdd.n2565 vdd.n1014 99.5127
R18707 vdd.n2565 vdd.n1011 99.5127
R18708 vdd.n2571 vdd.n1011 99.5127
R18709 vdd.n2571 vdd.n1012 99.5127
R18710 vdd.n1012 vdd.n1003 99.5127
R18711 vdd.n1003 vdd.n994 99.5127
R18712 vdd.n2653 vdd.n994 99.5127
R18713 vdd.n9 vdd.n7 98.9633
R18714 vdd.n2 vdd.n0 98.9633
R18715 vdd.n9 vdd.n8 98.6055
R18716 vdd.n11 vdd.n10 98.6055
R18717 vdd.n13 vdd.n12 98.6055
R18718 vdd.n6 vdd.n5 98.6055
R18719 vdd.n4 vdd.n3 98.6055
R18720 vdd.n2 vdd.n1 98.6055
R18721 vdd.t172 vdd.n303 85.8723
R18722 vdd.t213 vdd.n244 85.8723
R18723 vdd.t152 vdd.n201 85.8723
R18724 vdd.t193 vdd.n142 85.8723
R18725 vdd.t236 vdd.n100 85.8723
R18726 vdd.t262 vdd.n41 85.8723
R18727 vdd.t292 vdd.n1802 85.8723
R18728 vdd.t241 vdd.n1861 85.8723
R18729 vdd.t280 vdd.n1700 85.8723
R18730 vdd.t229 vdd.n1759 85.8723
R18731 vdd.t233 vdd.n1599 85.8723
R18732 vdd.t238 vdd.n1658 85.8723
R18733 vdd.n3080 vdd.n885 78.546
R18734 vdd.n2519 vdd.n1058 78.546
R18735 vdd.n290 vdd.n289 75.1835
R18736 vdd.n288 vdd.n287 75.1835
R18737 vdd.n286 vdd.n285 75.1835
R18738 vdd.n284 vdd.n283 75.1835
R18739 vdd.n282 vdd.n281 75.1835
R18740 vdd.n280 vdd.n279 75.1835
R18741 vdd.n278 vdd.n277 75.1835
R18742 vdd.n276 vdd.n275 75.1835
R18743 vdd.n274 vdd.n273 75.1835
R18744 vdd.n188 vdd.n187 75.1835
R18745 vdd.n186 vdd.n185 75.1835
R18746 vdd.n184 vdd.n183 75.1835
R18747 vdd.n182 vdd.n181 75.1835
R18748 vdd.n180 vdd.n179 75.1835
R18749 vdd.n178 vdd.n177 75.1835
R18750 vdd.n176 vdd.n175 75.1835
R18751 vdd.n174 vdd.n173 75.1835
R18752 vdd.n172 vdd.n171 75.1835
R18753 vdd.n87 vdd.n86 75.1835
R18754 vdd.n85 vdd.n84 75.1835
R18755 vdd.n83 vdd.n82 75.1835
R18756 vdd.n81 vdd.n80 75.1835
R18757 vdd.n79 vdd.n78 75.1835
R18758 vdd.n77 vdd.n76 75.1835
R18759 vdd.n75 vdd.n74 75.1835
R18760 vdd.n73 vdd.n72 75.1835
R18761 vdd.n71 vdd.n70 75.1835
R18762 vdd.n1832 vdd.n1831 75.1835
R18763 vdd.n1834 vdd.n1833 75.1835
R18764 vdd.n1836 vdd.n1835 75.1835
R18765 vdd.n1838 vdd.n1837 75.1835
R18766 vdd.n1840 vdd.n1839 75.1835
R18767 vdd.n1842 vdd.n1841 75.1835
R18768 vdd.n1844 vdd.n1843 75.1835
R18769 vdd.n1846 vdd.n1845 75.1835
R18770 vdd.n1848 vdd.n1847 75.1835
R18771 vdd.n1730 vdd.n1729 75.1835
R18772 vdd.n1732 vdd.n1731 75.1835
R18773 vdd.n1734 vdd.n1733 75.1835
R18774 vdd.n1736 vdd.n1735 75.1835
R18775 vdd.n1738 vdd.n1737 75.1835
R18776 vdd.n1740 vdd.n1739 75.1835
R18777 vdd.n1742 vdd.n1741 75.1835
R18778 vdd.n1744 vdd.n1743 75.1835
R18779 vdd.n1746 vdd.n1745 75.1835
R18780 vdd.n1629 vdd.n1628 75.1835
R18781 vdd.n1631 vdd.n1630 75.1835
R18782 vdd.n1633 vdd.n1632 75.1835
R18783 vdd.n1635 vdd.n1634 75.1835
R18784 vdd.n1637 vdd.n1636 75.1835
R18785 vdd.n1639 vdd.n1638 75.1835
R18786 vdd.n1641 vdd.n1640 75.1835
R18787 vdd.n1643 vdd.n1642 75.1835
R18788 vdd.n1645 vdd.n1644 75.1835
R18789 vdd.n3010 vdd.n2743 72.8958
R18790 vdd.n3010 vdd.n2744 72.8958
R18791 vdd.n3010 vdd.n2745 72.8958
R18792 vdd.n3010 vdd.n2746 72.8958
R18793 vdd.n3010 vdd.n2747 72.8958
R18794 vdd.n3010 vdd.n2748 72.8958
R18795 vdd.n3010 vdd.n2749 72.8958
R18796 vdd.n3010 vdd.n2750 72.8958
R18797 vdd.n3010 vdd.n2751 72.8958
R18798 vdd.n3010 vdd.n2752 72.8958
R18799 vdd.n3010 vdd.n2753 72.8958
R18800 vdd.n3010 vdd.n2754 72.8958
R18801 vdd.n3010 vdd.n2755 72.8958
R18802 vdd.n3010 vdd.n2756 72.8958
R18803 vdd.n3010 vdd.n2757 72.8958
R18804 vdd.n3010 vdd.n2758 72.8958
R18805 vdd.n3010 vdd.n2759 72.8958
R18806 vdd.n803 vdd.n692 72.8958
R18807 vdd.n3248 vdd.n692 72.8958
R18808 vdd.n797 vdd.n692 72.8958
R18809 vdd.n3255 vdd.n692 72.8958
R18810 vdd.n794 vdd.n692 72.8958
R18811 vdd.n3262 vdd.n692 72.8958
R18812 vdd.n791 vdd.n692 72.8958
R18813 vdd.n3269 vdd.n692 72.8958
R18814 vdd.n3272 vdd.n692 72.8958
R18815 vdd.n3128 vdd.n692 72.8958
R18816 vdd.n3133 vdd.n692 72.8958
R18817 vdd.n3127 vdd.n692 72.8958
R18818 vdd.n3140 vdd.n692 72.8958
R18819 vdd.n3124 vdd.n692 72.8958
R18820 vdd.n3147 vdd.n692 72.8958
R18821 vdd.n3121 vdd.n692 72.8958
R18822 vdd.n3154 vdd.n692 72.8958
R18823 vdd.n2461 vdd.n1110 72.8958
R18824 vdd.n1115 vdd.n1110 72.8958
R18825 vdd.n2454 vdd.n1110 72.8958
R18826 vdd.n2448 vdd.n1110 72.8958
R18827 vdd.n2446 vdd.n1110 72.8958
R18828 vdd.n2440 vdd.n1110 72.8958
R18829 vdd.n2438 vdd.n1110 72.8958
R18830 vdd.n2432 vdd.n1110 72.8958
R18831 vdd.n2430 vdd.n1110 72.8958
R18832 vdd.n2424 vdd.n1110 72.8958
R18833 vdd.n2422 vdd.n1110 72.8958
R18834 vdd.n2416 vdd.n1110 72.8958
R18835 vdd.n2414 vdd.n1110 72.8958
R18836 vdd.n2408 vdd.n1110 72.8958
R18837 vdd.n2406 vdd.n1110 72.8958
R18838 vdd.n2399 vdd.n1110 72.8958
R18839 vdd.n2397 vdd.n1110 72.8958
R18840 vdd.n2726 vdd.n968 72.8958
R18841 vdd.n2726 vdd.n969 72.8958
R18842 vdd.n2726 vdd.n970 72.8958
R18843 vdd.n2726 vdd.n971 72.8958
R18844 vdd.n2726 vdd.n972 72.8958
R18845 vdd.n2726 vdd.n973 72.8958
R18846 vdd.n2726 vdd.n974 72.8958
R18847 vdd.n2726 vdd.n975 72.8958
R18848 vdd.n2726 vdd.n976 72.8958
R18849 vdd.n2726 vdd.n977 72.8958
R18850 vdd.n2726 vdd.n978 72.8958
R18851 vdd.n2726 vdd.n979 72.8958
R18852 vdd.n2726 vdd.n980 72.8958
R18853 vdd.n2726 vdd.n981 72.8958
R18854 vdd.n2726 vdd.n982 72.8958
R18855 vdd.n2726 vdd.n983 72.8958
R18856 vdd.n2726 vdd.n984 72.8958
R18857 vdd.n3011 vdd.n3010 72.8958
R18858 vdd.n3010 vdd.n2727 72.8958
R18859 vdd.n3010 vdd.n2728 72.8958
R18860 vdd.n3010 vdd.n2729 72.8958
R18861 vdd.n3010 vdd.n2730 72.8958
R18862 vdd.n3010 vdd.n2731 72.8958
R18863 vdd.n3010 vdd.n2732 72.8958
R18864 vdd.n3010 vdd.n2733 72.8958
R18865 vdd.n3010 vdd.n2734 72.8958
R18866 vdd.n3010 vdd.n2735 72.8958
R18867 vdd.n3010 vdd.n2736 72.8958
R18868 vdd.n3010 vdd.n2737 72.8958
R18869 vdd.n3010 vdd.n2738 72.8958
R18870 vdd.n3010 vdd.n2739 72.8958
R18871 vdd.n3010 vdd.n2740 72.8958
R18872 vdd.n3010 vdd.n2741 72.8958
R18873 vdd.n3010 vdd.n2742 72.8958
R18874 vdd.n3178 vdd.n692 72.8958
R18875 vdd.n835 vdd.n692 72.8958
R18876 vdd.n3186 vdd.n692 72.8958
R18877 vdd.n830 vdd.n692 72.8958
R18878 vdd.n3193 vdd.n692 72.8958
R18879 vdd.n827 vdd.n692 72.8958
R18880 vdd.n3200 vdd.n692 72.8958
R18881 vdd.n824 vdd.n692 72.8958
R18882 vdd.n3207 vdd.n692 72.8958
R18883 vdd.n3211 vdd.n692 72.8958
R18884 vdd.n821 vdd.n692 72.8958
R18885 vdd.n3218 vdd.n692 72.8958
R18886 vdd.n818 vdd.n692 72.8958
R18887 vdd.n3225 vdd.n692 72.8958
R18888 vdd.n815 vdd.n692 72.8958
R18889 vdd.n3232 vdd.n692 72.8958
R18890 vdd.n3235 vdd.n692 72.8958
R18891 vdd.n2726 vdd.n966 72.8958
R18892 vdd.n2726 vdd.n965 72.8958
R18893 vdd.n2726 vdd.n964 72.8958
R18894 vdd.n2726 vdd.n963 72.8958
R18895 vdd.n2726 vdd.n962 72.8958
R18896 vdd.n2726 vdd.n961 72.8958
R18897 vdd.n2726 vdd.n960 72.8958
R18898 vdd.n2726 vdd.n959 72.8958
R18899 vdd.n2726 vdd.n958 72.8958
R18900 vdd.n2726 vdd.n957 72.8958
R18901 vdd.n2726 vdd.n956 72.8958
R18902 vdd.n2726 vdd.n955 72.8958
R18903 vdd.n2726 vdd.n954 72.8958
R18904 vdd.n2726 vdd.n953 72.8958
R18905 vdd.n2726 vdd.n952 72.8958
R18906 vdd.n2726 vdd.n951 72.8958
R18907 vdd.n2726 vdd.n950 72.8958
R18908 vdd.n2215 vdd.n1110 72.8958
R18909 vdd.n2217 vdd.n1110 72.8958
R18910 vdd.n2223 vdd.n1110 72.8958
R18911 vdd.n2225 vdd.n1110 72.8958
R18912 vdd.n2231 vdd.n1110 72.8958
R18913 vdd.n2233 vdd.n1110 72.8958
R18914 vdd.n2239 vdd.n1110 72.8958
R18915 vdd.n2241 vdd.n1110 72.8958
R18916 vdd.n2247 vdd.n1110 72.8958
R18917 vdd.n2249 vdd.n1110 72.8958
R18918 vdd.n2255 vdd.n1110 72.8958
R18919 vdd.n2257 vdd.n1110 72.8958
R18920 vdd.n2263 vdd.n1110 72.8958
R18921 vdd.n2265 vdd.n1110 72.8958
R18922 vdd.n2271 vdd.n1110 72.8958
R18923 vdd.n2273 vdd.n1110 72.8958
R18924 vdd.n2280 vdd.n1110 72.8958
R18925 vdd.n1499 vdd.n1498 66.2847
R18926 vdd.n1498 vdd.n1274 66.2847
R18927 vdd.n1498 vdd.n1275 66.2847
R18928 vdd.n1498 vdd.n1276 66.2847
R18929 vdd.n1498 vdd.n1277 66.2847
R18930 vdd.n1498 vdd.n1278 66.2847
R18931 vdd.n1498 vdd.n1279 66.2847
R18932 vdd.n1498 vdd.n1280 66.2847
R18933 vdd.n1498 vdd.n1281 66.2847
R18934 vdd.n1498 vdd.n1282 66.2847
R18935 vdd.n1498 vdd.n1283 66.2847
R18936 vdd.n1498 vdd.n1284 66.2847
R18937 vdd.n1498 vdd.n1285 66.2847
R18938 vdd.n1498 vdd.n1286 66.2847
R18939 vdd.n1498 vdd.n1287 66.2847
R18940 vdd.n1498 vdd.n1288 66.2847
R18941 vdd.n1498 vdd.n1289 66.2847
R18942 vdd.n1498 vdd.n1290 66.2847
R18943 vdd.n1498 vdd.n1291 66.2847
R18944 vdd.n1498 vdd.n1292 66.2847
R18945 vdd.n1498 vdd.n1293 66.2847
R18946 vdd.n1498 vdd.n1294 66.2847
R18947 vdd.n1498 vdd.n1295 66.2847
R18948 vdd.n1498 vdd.n1296 66.2847
R18949 vdd.n1498 vdd.n1297 66.2847
R18950 vdd.n1498 vdd.n1298 66.2847
R18951 vdd.n1498 vdd.n1299 66.2847
R18952 vdd.n1498 vdd.n1300 66.2847
R18953 vdd.n1498 vdd.n1301 66.2847
R18954 vdd.n1498 vdd.n1302 66.2847
R18955 vdd.n1498 vdd.n1303 66.2847
R18956 vdd.n1153 vdd.n1150 66.2847
R18957 vdd.n2080 vdd.n1153 66.2847
R18958 vdd.n2085 vdd.n1153 66.2847
R18959 vdd.n2090 vdd.n1153 66.2847
R18960 vdd.n2078 vdd.n1153 66.2847
R18961 vdd.n2097 vdd.n1153 66.2847
R18962 vdd.n2070 vdd.n1153 66.2847
R18963 vdd.n2104 vdd.n1153 66.2847
R18964 vdd.n2063 vdd.n1153 66.2847
R18965 vdd.n2111 vdd.n1153 66.2847
R18966 vdd.n2057 vdd.n1153 66.2847
R18967 vdd.n2052 vdd.n1153 66.2847
R18968 vdd.n2122 vdd.n1153 66.2847
R18969 vdd.n2044 vdd.n1153 66.2847
R18970 vdd.n2129 vdd.n1153 66.2847
R18971 vdd.n2037 vdd.n1153 66.2847
R18972 vdd.n2136 vdd.n1153 66.2847
R18973 vdd.n2030 vdd.n1153 66.2847
R18974 vdd.n2143 vdd.n1153 66.2847
R18975 vdd.n2023 vdd.n1153 66.2847
R18976 vdd.n2150 vdd.n1153 66.2847
R18977 vdd.n2017 vdd.n1153 66.2847
R18978 vdd.n2012 vdd.n1153 66.2847
R18979 vdd.n2161 vdd.n1153 66.2847
R18980 vdd.n2004 vdd.n1153 66.2847
R18981 vdd.n2168 vdd.n1153 66.2847
R18982 vdd.n1997 vdd.n1153 66.2847
R18983 vdd.n2175 vdd.n1153 66.2847
R18984 vdd.n2178 vdd.n1153 66.2847
R18985 vdd.n1988 vdd.n1153 66.2847
R18986 vdd.n2187 vdd.n1153 66.2847
R18987 vdd.n1982 vdd.n1153 66.2847
R18988 vdd.n3405 vdd.n3404 66.2847
R18989 vdd.n3405 vdd.n693 66.2847
R18990 vdd.n3405 vdd.n694 66.2847
R18991 vdd.n3405 vdd.n695 66.2847
R18992 vdd.n3405 vdd.n696 66.2847
R18993 vdd.n3405 vdd.n697 66.2847
R18994 vdd.n3405 vdd.n698 66.2847
R18995 vdd.n3405 vdd.n699 66.2847
R18996 vdd.n3405 vdd.n700 66.2847
R18997 vdd.n3405 vdd.n701 66.2847
R18998 vdd.n3405 vdd.n702 66.2847
R18999 vdd.n3405 vdd.n703 66.2847
R19000 vdd.n3405 vdd.n704 66.2847
R19001 vdd.n3405 vdd.n705 66.2847
R19002 vdd.n3405 vdd.n706 66.2847
R19003 vdd.n3405 vdd.n707 66.2847
R19004 vdd.n3405 vdd.n708 66.2847
R19005 vdd.n3405 vdd.n709 66.2847
R19006 vdd.n3405 vdd.n710 66.2847
R19007 vdd.n3405 vdd.n711 66.2847
R19008 vdd.n3405 vdd.n712 66.2847
R19009 vdd.n3405 vdd.n713 66.2847
R19010 vdd.n3405 vdd.n714 66.2847
R19011 vdd.n3405 vdd.n715 66.2847
R19012 vdd.n3405 vdd.n716 66.2847
R19013 vdd.n3405 vdd.n717 66.2847
R19014 vdd.n3405 vdd.n718 66.2847
R19015 vdd.n3405 vdd.n719 66.2847
R19016 vdd.n3405 vdd.n720 66.2847
R19017 vdd.n3405 vdd.n721 66.2847
R19018 vdd.n3405 vdd.n722 66.2847
R19019 vdd.n3536 vdd.n3535 66.2847
R19020 vdd.n3536 vdd.n424 66.2847
R19021 vdd.n3536 vdd.n423 66.2847
R19022 vdd.n3536 vdd.n422 66.2847
R19023 vdd.n3536 vdd.n421 66.2847
R19024 vdd.n3536 vdd.n420 66.2847
R19025 vdd.n3536 vdd.n419 66.2847
R19026 vdd.n3536 vdd.n418 66.2847
R19027 vdd.n3536 vdd.n417 66.2847
R19028 vdd.n3536 vdd.n416 66.2847
R19029 vdd.n3536 vdd.n415 66.2847
R19030 vdd.n3536 vdd.n414 66.2847
R19031 vdd.n3536 vdd.n413 66.2847
R19032 vdd.n3536 vdd.n412 66.2847
R19033 vdd.n3536 vdd.n411 66.2847
R19034 vdd.n3536 vdd.n410 66.2847
R19035 vdd.n3536 vdd.n409 66.2847
R19036 vdd.n3536 vdd.n408 66.2847
R19037 vdd.n3536 vdd.n407 66.2847
R19038 vdd.n3536 vdd.n406 66.2847
R19039 vdd.n3536 vdd.n405 66.2847
R19040 vdd.n3536 vdd.n404 66.2847
R19041 vdd.n3536 vdd.n403 66.2847
R19042 vdd.n3536 vdd.n402 66.2847
R19043 vdd.n3536 vdd.n401 66.2847
R19044 vdd.n3536 vdd.n400 66.2847
R19045 vdd.n3536 vdd.n399 66.2847
R19046 vdd.n3536 vdd.n398 66.2847
R19047 vdd.n3536 vdd.n397 66.2847
R19048 vdd.n3536 vdd.n396 66.2847
R19049 vdd.n3536 vdd.n395 66.2847
R19050 vdd.n3536 vdd.n394 66.2847
R19051 vdd.n467 vdd.n394 52.4337
R19052 vdd.n473 vdd.n395 52.4337
R19053 vdd.n477 vdd.n396 52.4337
R19054 vdd.n483 vdd.n397 52.4337
R19055 vdd.n487 vdd.n398 52.4337
R19056 vdd.n493 vdd.n399 52.4337
R19057 vdd.n497 vdd.n400 52.4337
R19058 vdd.n503 vdd.n401 52.4337
R19059 vdd.n507 vdd.n402 52.4337
R19060 vdd.n513 vdd.n403 52.4337
R19061 vdd.n517 vdd.n404 52.4337
R19062 vdd.n523 vdd.n405 52.4337
R19063 vdd.n527 vdd.n406 52.4337
R19064 vdd.n533 vdd.n407 52.4337
R19065 vdd.n537 vdd.n408 52.4337
R19066 vdd.n543 vdd.n409 52.4337
R19067 vdd.n547 vdd.n410 52.4337
R19068 vdd.n553 vdd.n411 52.4337
R19069 vdd.n557 vdd.n412 52.4337
R19070 vdd.n563 vdd.n413 52.4337
R19071 vdd.n567 vdd.n414 52.4337
R19072 vdd.n573 vdd.n415 52.4337
R19073 vdd.n577 vdd.n416 52.4337
R19074 vdd.n583 vdd.n417 52.4337
R19075 vdd.n587 vdd.n418 52.4337
R19076 vdd.n593 vdd.n419 52.4337
R19077 vdd.n597 vdd.n420 52.4337
R19078 vdd.n603 vdd.n421 52.4337
R19079 vdd.n607 vdd.n422 52.4337
R19080 vdd.n613 vdd.n423 52.4337
R19081 vdd.n616 vdd.n424 52.4337
R19082 vdd.n3535 vdd.n3534 52.4337
R19083 vdd.n3404 vdd.n3403 52.4337
R19084 vdd.n728 vdd.n693 52.4337
R19085 vdd.n734 vdd.n694 52.4337
R19086 vdd.n3393 vdd.n695 52.4337
R19087 vdd.n3389 vdd.n696 52.4337
R19088 vdd.n3385 vdd.n697 52.4337
R19089 vdd.n3381 vdd.n698 52.4337
R19090 vdd.n3377 vdd.n699 52.4337
R19091 vdd.n3373 vdd.n700 52.4337
R19092 vdd.n3369 vdd.n701 52.4337
R19093 vdd.n3361 vdd.n702 52.4337
R19094 vdd.n3357 vdd.n703 52.4337
R19095 vdd.n3353 vdd.n704 52.4337
R19096 vdd.n3349 vdd.n705 52.4337
R19097 vdd.n3345 vdd.n706 52.4337
R19098 vdd.n3341 vdd.n707 52.4337
R19099 vdd.n3337 vdd.n708 52.4337
R19100 vdd.n3333 vdd.n709 52.4337
R19101 vdd.n3329 vdd.n710 52.4337
R19102 vdd.n3325 vdd.n711 52.4337
R19103 vdd.n3321 vdd.n712 52.4337
R19104 vdd.n3315 vdd.n713 52.4337
R19105 vdd.n3311 vdd.n714 52.4337
R19106 vdd.n3307 vdd.n715 52.4337
R19107 vdd.n3303 vdd.n716 52.4337
R19108 vdd.n3299 vdd.n717 52.4337
R19109 vdd.n3295 vdd.n718 52.4337
R19110 vdd.n3291 vdd.n719 52.4337
R19111 vdd.n3287 vdd.n720 52.4337
R19112 vdd.n3283 vdd.n721 52.4337
R19113 vdd.n3279 vdd.n722 52.4337
R19114 vdd.n2189 vdd.n1982 52.4337
R19115 vdd.n2187 vdd.n2186 52.4337
R19116 vdd.n1989 vdd.n1988 52.4337
R19117 vdd.n2178 vdd.n2177 52.4337
R19118 vdd.n2175 vdd.n2174 52.4337
R19119 vdd.n2170 vdd.n1997 52.4337
R19120 vdd.n2168 vdd.n2167 52.4337
R19121 vdd.n2163 vdd.n2004 52.4337
R19122 vdd.n2161 vdd.n2160 52.4337
R19123 vdd.n2013 vdd.n2012 52.4337
R19124 vdd.n2152 vdd.n2017 52.4337
R19125 vdd.n2150 vdd.n2149 52.4337
R19126 vdd.n2145 vdd.n2023 52.4337
R19127 vdd.n2143 vdd.n2142 52.4337
R19128 vdd.n2138 vdd.n2030 52.4337
R19129 vdd.n2136 vdd.n2135 52.4337
R19130 vdd.n2131 vdd.n2037 52.4337
R19131 vdd.n2129 vdd.n2128 52.4337
R19132 vdd.n2124 vdd.n2044 52.4337
R19133 vdd.n2122 vdd.n2121 52.4337
R19134 vdd.n2053 vdd.n2052 52.4337
R19135 vdd.n2113 vdd.n2057 52.4337
R19136 vdd.n2111 vdd.n2110 52.4337
R19137 vdd.n2106 vdd.n2063 52.4337
R19138 vdd.n2104 vdd.n2103 52.4337
R19139 vdd.n2099 vdd.n2070 52.4337
R19140 vdd.n2097 vdd.n2096 52.4337
R19141 vdd.n2092 vdd.n2078 52.4337
R19142 vdd.n2090 vdd.n2089 52.4337
R19143 vdd.n2085 vdd.n2084 52.4337
R19144 vdd.n2080 vdd.n2079 52.4337
R19145 vdd.n2198 vdd.n1150 52.4337
R19146 vdd.n1500 vdd.n1499 52.4337
R19147 vdd.n1306 vdd.n1274 52.4337
R19148 vdd.n1310 vdd.n1275 52.4337
R19149 vdd.n1312 vdd.n1276 52.4337
R19150 vdd.n1316 vdd.n1277 52.4337
R19151 vdd.n1318 vdd.n1278 52.4337
R19152 vdd.n1322 vdd.n1279 52.4337
R19153 vdd.n1324 vdd.n1280 52.4337
R19154 vdd.n1328 vdd.n1281 52.4337
R19155 vdd.n1330 vdd.n1282 52.4337
R19156 vdd.n1336 vdd.n1283 52.4337
R19157 vdd.n1338 vdd.n1284 52.4337
R19158 vdd.n1342 vdd.n1285 52.4337
R19159 vdd.n1344 vdd.n1286 52.4337
R19160 vdd.n1348 vdd.n1287 52.4337
R19161 vdd.n1350 vdd.n1288 52.4337
R19162 vdd.n1354 vdd.n1289 52.4337
R19163 vdd.n1356 vdd.n1290 52.4337
R19164 vdd.n1360 vdd.n1291 52.4337
R19165 vdd.n1362 vdd.n1292 52.4337
R19166 vdd.n1434 vdd.n1293 52.4337
R19167 vdd.n1367 vdd.n1294 52.4337
R19168 vdd.n1371 vdd.n1295 52.4337
R19169 vdd.n1373 vdd.n1296 52.4337
R19170 vdd.n1377 vdd.n1297 52.4337
R19171 vdd.n1379 vdd.n1298 52.4337
R19172 vdd.n1383 vdd.n1299 52.4337
R19173 vdd.n1385 vdd.n1300 52.4337
R19174 vdd.n1389 vdd.n1301 52.4337
R19175 vdd.n1391 vdd.n1302 52.4337
R19176 vdd.n1395 vdd.n1303 52.4337
R19177 vdd.n1499 vdd.n1273 52.4337
R19178 vdd.n1309 vdd.n1274 52.4337
R19179 vdd.n1311 vdd.n1275 52.4337
R19180 vdd.n1315 vdd.n1276 52.4337
R19181 vdd.n1317 vdd.n1277 52.4337
R19182 vdd.n1321 vdd.n1278 52.4337
R19183 vdd.n1323 vdd.n1279 52.4337
R19184 vdd.n1327 vdd.n1280 52.4337
R19185 vdd.n1329 vdd.n1281 52.4337
R19186 vdd.n1335 vdd.n1282 52.4337
R19187 vdd.n1337 vdd.n1283 52.4337
R19188 vdd.n1341 vdd.n1284 52.4337
R19189 vdd.n1343 vdd.n1285 52.4337
R19190 vdd.n1347 vdd.n1286 52.4337
R19191 vdd.n1349 vdd.n1287 52.4337
R19192 vdd.n1353 vdd.n1288 52.4337
R19193 vdd.n1355 vdd.n1289 52.4337
R19194 vdd.n1359 vdd.n1290 52.4337
R19195 vdd.n1361 vdd.n1291 52.4337
R19196 vdd.n1365 vdd.n1292 52.4337
R19197 vdd.n1366 vdd.n1293 52.4337
R19198 vdd.n1370 vdd.n1294 52.4337
R19199 vdd.n1372 vdd.n1295 52.4337
R19200 vdd.n1376 vdd.n1296 52.4337
R19201 vdd.n1378 vdd.n1297 52.4337
R19202 vdd.n1382 vdd.n1298 52.4337
R19203 vdd.n1384 vdd.n1299 52.4337
R19204 vdd.n1388 vdd.n1300 52.4337
R19205 vdd.n1390 vdd.n1301 52.4337
R19206 vdd.n1394 vdd.n1302 52.4337
R19207 vdd.n1396 vdd.n1303 52.4337
R19208 vdd.n1150 vdd.n1149 52.4337
R19209 vdd.n2081 vdd.n2080 52.4337
R19210 vdd.n2086 vdd.n2085 52.4337
R19211 vdd.n2091 vdd.n2090 52.4337
R19212 vdd.n2078 vdd.n2071 52.4337
R19213 vdd.n2098 vdd.n2097 52.4337
R19214 vdd.n2070 vdd.n2064 52.4337
R19215 vdd.n2105 vdd.n2104 52.4337
R19216 vdd.n2063 vdd.n2058 52.4337
R19217 vdd.n2112 vdd.n2111 52.4337
R19218 vdd.n2057 vdd.n2056 52.4337
R19219 vdd.n2052 vdd.n2045 52.4337
R19220 vdd.n2123 vdd.n2122 52.4337
R19221 vdd.n2044 vdd.n2038 52.4337
R19222 vdd.n2130 vdd.n2129 52.4337
R19223 vdd.n2037 vdd.n2031 52.4337
R19224 vdd.n2137 vdd.n2136 52.4337
R19225 vdd.n2030 vdd.n2024 52.4337
R19226 vdd.n2144 vdd.n2143 52.4337
R19227 vdd.n2023 vdd.n2018 52.4337
R19228 vdd.n2151 vdd.n2150 52.4337
R19229 vdd.n2017 vdd.n2016 52.4337
R19230 vdd.n2012 vdd.n2005 52.4337
R19231 vdd.n2162 vdd.n2161 52.4337
R19232 vdd.n2004 vdd.n1998 52.4337
R19233 vdd.n2169 vdd.n2168 52.4337
R19234 vdd.n1997 vdd.n1991 52.4337
R19235 vdd.n2176 vdd.n2175 52.4337
R19236 vdd.n2179 vdd.n2178 52.4337
R19237 vdd.n1988 vdd.n1983 52.4337
R19238 vdd.n2188 vdd.n2187 52.4337
R19239 vdd.n1982 vdd.n1155 52.4337
R19240 vdd.n3404 vdd.n725 52.4337
R19241 vdd.n733 vdd.n693 52.4337
R19242 vdd.n3394 vdd.n694 52.4337
R19243 vdd.n3390 vdd.n695 52.4337
R19244 vdd.n3386 vdd.n696 52.4337
R19245 vdd.n3382 vdd.n697 52.4337
R19246 vdd.n3378 vdd.n698 52.4337
R19247 vdd.n3374 vdd.n699 52.4337
R19248 vdd.n3370 vdd.n700 52.4337
R19249 vdd.n3360 vdd.n701 52.4337
R19250 vdd.n3358 vdd.n702 52.4337
R19251 vdd.n3354 vdd.n703 52.4337
R19252 vdd.n3350 vdd.n704 52.4337
R19253 vdd.n3346 vdd.n705 52.4337
R19254 vdd.n3342 vdd.n706 52.4337
R19255 vdd.n3338 vdd.n707 52.4337
R19256 vdd.n3334 vdd.n708 52.4337
R19257 vdd.n3330 vdd.n709 52.4337
R19258 vdd.n3326 vdd.n710 52.4337
R19259 vdd.n3322 vdd.n711 52.4337
R19260 vdd.n3314 vdd.n712 52.4337
R19261 vdd.n3312 vdd.n713 52.4337
R19262 vdd.n3308 vdd.n714 52.4337
R19263 vdd.n3304 vdd.n715 52.4337
R19264 vdd.n3300 vdd.n716 52.4337
R19265 vdd.n3296 vdd.n717 52.4337
R19266 vdd.n3292 vdd.n718 52.4337
R19267 vdd.n3288 vdd.n719 52.4337
R19268 vdd.n3284 vdd.n720 52.4337
R19269 vdd.n3280 vdd.n721 52.4337
R19270 vdd.n722 vdd.n691 52.4337
R19271 vdd.n3535 vdd.n425 52.4337
R19272 vdd.n614 vdd.n424 52.4337
R19273 vdd.n608 vdd.n423 52.4337
R19274 vdd.n604 vdd.n422 52.4337
R19275 vdd.n598 vdd.n421 52.4337
R19276 vdd.n594 vdd.n420 52.4337
R19277 vdd.n588 vdd.n419 52.4337
R19278 vdd.n584 vdd.n418 52.4337
R19279 vdd.n578 vdd.n417 52.4337
R19280 vdd.n574 vdd.n416 52.4337
R19281 vdd.n568 vdd.n415 52.4337
R19282 vdd.n564 vdd.n414 52.4337
R19283 vdd.n558 vdd.n413 52.4337
R19284 vdd.n554 vdd.n412 52.4337
R19285 vdd.n548 vdd.n411 52.4337
R19286 vdd.n544 vdd.n410 52.4337
R19287 vdd.n538 vdd.n409 52.4337
R19288 vdd.n534 vdd.n408 52.4337
R19289 vdd.n528 vdd.n407 52.4337
R19290 vdd.n524 vdd.n406 52.4337
R19291 vdd.n518 vdd.n405 52.4337
R19292 vdd.n514 vdd.n404 52.4337
R19293 vdd.n508 vdd.n403 52.4337
R19294 vdd.n504 vdd.n402 52.4337
R19295 vdd.n498 vdd.n401 52.4337
R19296 vdd.n494 vdd.n400 52.4337
R19297 vdd.n488 vdd.n399 52.4337
R19298 vdd.n484 vdd.n398 52.4337
R19299 vdd.n478 vdd.n397 52.4337
R19300 vdd.n474 vdd.n396 52.4337
R19301 vdd.n468 vdd.n395 52.4337
R19302 vdd.n394 vdd.n392 52.4337
R19303 vdd.t298 vdd.t43 51.4683
R19304 vdd.n274 vdd.n272 42.0461
R19305 vdd.n172 vdd.n170 42.0461
R19306 vdd.n71 vdd.n69 42.0461
R19307 vdd.n1832 vdd.n1830 42.0461
R19308 vdd.n1730 vdd.n1728 42.0461
R19309 vdd.n1629 vdd.n1627 42.0461
R19310 vdd.n332 vdd.n331 41.6884
R19311 vdd.n230 vdd.n229 41.6884
R19312 vdd.n129 vdd.n128 41.6884
R19313 vdd.n1890 vdd.n1889 41.6884
R19314 vdd.n1788 vdd.n1787 41.6884
R19315 vdd.n1687 vdd.n1686 41.6884
R19316 vdd.n1399 vdd.n1398 41.1157
R19317 vdd.n1437 vdd.n1436 41.1157
R19318 vdd.n1333 vdd.n1332 41.1157
R19319 vdd.n428 vdd.n427 41.1157
R19320 vdd.n566 vdd.n441 41.1157
R19321 vdd.n454 vdd.n453 41.1157
R19322 vdd.n3235 vdd.n3234 39.2114
R19323 vdd.n3232 vdd.n3231 39.2114
R19324 vdd.n3227 vdd.n815 39.2114
R19325 vdd.n3225 vdd.n3224 39.2114
R19326 vdd.n3220 vdd.n818 39.2114
R19327 vdd.n3218 vdd.n3217 39.2114
R19328 vdd.n3213 vdd.n821 39.2114
R19329 vdd.n3211 vdd.n3210 39.2114
R19330 vdd.n3207 vdd.n3206 39.2114
R19331 vdd.n3202 vdd.n824 39.2114
R19332 vdd.n3200 vdd.n3199 39.2114
R19333 vdd.n3195 vdd.n827 39.2114
R19334 vdd.n3193 vdd.n3192 39.2114
R19335 vdd.n3188 vdd.n830 39.2114
R19336 vdd.n3186 vdd.n3185 39.2114
R19337 vdd.n3180 vdd.n835 39.2114
R19338 vdd.n3178 vdd.n3177 39.2114
R19339 vdd.n3011 vdd.n947 39.2114
R19340 vdd.n2832 vdd.n2727 39.2114
R19341 vdd.n2836 vdd.n2728 39.2114
R19342 vdd.n2840 vdd.n2729 39.2114
R19343 vdd.n2844 vdd.n2730 39.2114
R19344 vdd.n2848 vdd.n2731 39.2114
R19345 vdd.n2852 vdd.n2732 39.2114
R19346 vdd.n2856 vdd.n2733 39.2114
R19347 vdd.n2860 vdd.n2734 39.2114
R19348 vdd.n2864 vdd.n2735 39.2114
R19349 vdd.n2868 vdd.n2736 39.2114
R19350 vdd.n2872 vdd.n2737 39.2114
R19351 vdd.n2876 vdd.n2738 39.2114
R19352 vdd.n2880 vdd.n2739 39.2114
R19353 vdd.n2884 vdd.n2740 39.2114
R19354 vdd.n2888 vdd.n2741 39.2114
R19355 vdd.n2893 vdd.n2742 39.2114
R19356 vdd.n2721 vdd.n984 39.2114
R19357 vdd.n2717 vdd.n983 39.2114
R19358 vdd.n2713 vdd.n982 39.2114
R19359 vdd.n2709 vdd.n981 39.2114
R19360 vdd.n2705 vdd.n980 39.2114
R19361 vdd.n2701 vdd.n979 39.2114
R19362 vdd.n2697 vdd.n978 39.2114
R19363 vdd.n2693 vdd.n977 39.2114
R19364 vdd.n2689 vdd.n976 39.2114
R19365 vdd.n2685 vdd.n975 39.2114
R19366 vdd.n2681 vdd.n974 39.2114
R19367 vdd.n2677 vdd.n973 39.2114
R19368 vdd.n2673 vdd.n972 39.2114
R19369 vdd.n2669 vdd.n971 39.2114
R19370 vdd.n2665 vdd.n970 39.2114
R19371 vdd.n2660 vdd.n969 39.2114
R19372 vdd.n2656 vdd.n968 39.2114
R19373 vdd.n2461 vdd.n1113 39.2114
R19374 vdd.n2459 vdd.n1115 39.2114
R19375 vdd.n2455 vdd.n2454 39.2114
R19376 vdd.n2448 vdd.n1117 39.2114
R19377 vdd.n2447 vdd.n2446 39.2114
R19378 vdd.n2440 vdd.n1119 39.2114
R19379 vdd.n2439 vdd.n2438 39.2114
R19380 vdd.n2432 vdd.n1121 39.2114
R19381 vdd.n2431 vdd.n2430 39.2114
R19382 vdd.n2424 vdd.n1123 39.2114
R19383 vdd.n2423 vdd.n2422 39.2114
R19384 vdd.n2416 vdd.n1125 39.2114
R19385 vdd.n2415 vdd.n2414 39.2114
R19386 vdd.n2408 vdd.n1127 39.2114
R19387 vdd.n2407 vdd.n2406 39.2114
R19388 vdd.n2399 vdd.n1129 39.2114
R19389 vdd.n2398 vdd.n2397 39.2114
R19390 vdd.n3154 vdd.n3153 39.2114
R19391 vdd.n3149 vdd.n3121 39.2114
R19392 vdd.n3147 vdd.n3146 39.2114
R19393 vdd.n3142 vdd.n3124 39.2114
R19394 vdd.n3140 vdd.n3139 39.2114
R19395 vdd.n3135 vdd.n3127 39.2114
R19396 vdd.n3133 vdd.n3132 39.2114
R19397 vdd.n3128 vdd.n787 39.2114
R19398 vdd.n3272 vdd.n3271 39.2114
R19399 vdd.n3269 vdd.n3268 39.2114
R19400 vdd.n3264 vdd.n791 39.2114
R19401 vdd.n3262 vdd.n3261 39.2114
R19402 vdd.n3257 vdd.n794 39.2114
R19403 vdd.n3255 vdd.n3254 39.2114
R19404 vdd.n3250 vdd.n797 39.2114
R19405 vdd.n3248 vdd.n3247 39.2114
R19406 vdd.n3243 vdd.n803 39.2114
R19407 vdd.n2743 vdd.n943 39.2114
R19408 vdd.n2766 vdd.n2744 39.2114
R19409 vdd.n2770 vdd.n2745 39.2114
R19410 vdd.n2774 vdd.n2746 39.2114
R19411 vdd.n2778 vdd.n2747 39.2114
R19412 vdd.n2782 vdd.n2748 39.2114
R19413 vdd.n2786 vdd.n2749 39.2114
R19414 vdd.n2790 vdd.n2750 39.2114
R19415 vdd.n2794 vdd.n2751 39.2114
R19416 vdd.n2798 vdd.n2752 39.2114
R19417 vdd.n2802 vdd.n2753 39.2114
R19418 vdd.n2806 vdd.n2754 39.2114
R19419 vdd.n2810 vdd.n2755 39.2114
R19420 vdd.n2814 vdd.n2756 39.2114
R19421 vdd.n2818 vdd.n2757 39.2114
R19422 vdd.n2822 vdd.n2758 39.2114
R19423 vdd.n2826 vdd.n2759 39.2114
R19424 vdd.n2765 vdd.n2743 39.2114
R19425 vdd.n2769 vdd.n2744 39.2114
R19426 vdd.n2773 vdd.n2745 39.2114
R19427 vdd.n2777 vdd.n2746 39.2114
R19428 vdd.n2781 vdd.n2747 39.2114
R19429 vdd.n2785 vdd.n2748 39.2114
R19430 vdd.n2789 vdd.n2749 39.2114
R19431 vdd.n2793 vdd.n2750 39.2114
R19432 vdd.n2797 vdd.n2751 39.2114
R19433 vdd.n2801 vdd.n2752 39.2114
R19434 vdd.n2805 vdd.n2753 39.2114
R19435 vdd.n2809 vdd.n2754 39.2114
R19436 vdd.n2813 vdd.n2755 39.2114
R19437 vdd.n2817 vdd.n2756 39.2114
R19438 vdd.n2821 vdd.n2757 39.2114
R19439 vdd.n2825 vdd.n2758 39.2114
R19440 vdd.n2760 vdd.n2759 39.2114
R19441 vdd.n803 vdd.n798 39.2114
R19442 vdd.n3249 vdd.n3248 39.2114
R19443 vdd.n797 vdd.n795 39.2114
R19444 vdd.n3256 vdd.n3255 39.2114
R19445 vdd.n794 vdd.n792 39.2114
R19446 vdd.n3263 vdd.n3262 39.2114
R19447 vdd.n791 vdd.n789 39.2114
R19448 vdd.n3270 vdd.n3269 39.2114
R19449 vdd.n3273 vdd.n3272 39.2114
R19450 vdd.n3129 vdd.n3128 39.2114
R19451 vdd.n3134 vdd.n3133 39.2114
R19452 vdd.n3127 vdd.n3125 39.2114
R19453 vdd.n3141 vdd.n3140 39.2114
R19454 vdd.n3124 vdd.n3122 39.2114
R19455 vdd.n3148 vdd.n3147 39.2114
R19456 vdd.n3121 vdd.n3119 39.2114
R19457 vdd.n3155 vdd.n3154 39.2114
R19458 vdd.n2462 vdd.n2461 39.2114
R19459 vdd.n2456 vdd.n1115 39.2114
R19460 vdd.n2454 vdd.n2453 39.2114
R19461 vdd.n2449 vdd.n2448 39.2114
R19462 vdd.n2446 vdd.n2445 39.2114
R19463 vdd.n2441 vdd.n2440 39.2114
R19464 vdd.n2438 vdd.n2437 39.2114
R19465 vdd.n2433 vdd.n2432 39.2114
R19466 vdd.n2430 vdd.n2429 39.2114
R19467 vdd.n2425 vdd.n2424 39.2114
R19468 vdd.n2422 vdd.n2421 39.2114
R19469 vdd.n2417 vdd.n2416 39.2114
R19470 vdd.n2414 vdd.n2413 39.2114
R19471 vdd.n2409 vdd.n2408 39.2114
R19472 vdd.n2406 vdd.n2405 39.2114
R19473 vdd.n2400 vdd.n2399 39.2114
R19474 vdd.n2397 vdd.n2396 39.2114
R19475 vdd.n2659 vdd.n968 39.2114
R19476 vdd.n2664 vdd.n969 39.2114
R19477 vdd.n2668 vdd.n970 39.2114
R19478 vdd.n2672 vdd.n971 39.2114
R19479 vdd.n2676 vdd.n972 39.2114
R19480 vdd.n2680 vdd.n973 39.2114
R19481 vdd.n2684 vdd.n974 39.2114
R19482 vdd.n2688 vdd.n975 39.2114
R19483 vdd.n2692 vdd.n976 39.2114
R19484 vdd.n2696 vdd.n977 39.2114
R19485 vdd.n2700 vdd.n978 39.2114
R19486 vdd.n2704 vdd.n979 39.2114
R19487 vdd.n2708 vdd.n980 39.2114
R19488 vdd.n2712 vdd.n981 39.2114
R19489 vdd.n2716 vdd.n982 39.2114
R19490 vdd.n2720 vdd.n983 39.2114
R19491 vdd.n986 vdd.n984 39.2114
R19492 vdd.n3012 vdd.n3011 39.2114
R19493 vdd.n2835 vdd.n2727 39.2114
R19494 vdd.n2839 vdd.n2728 39.2114
R19495 vdd.n2843 vdd.n2729 39.2114
R19496 vdd.n2847 vdd.n2730 39.2114
R19497 vdd.n2851 vdd.n2731 39.2114
R19498 vdd.n2855 vdd.n2732 39.2114
R19499 vdd.n2859 vdd.n2733 39.2114
R19500 vdd.n2863 vdd.n2734 39.2114
R19501 vdd.n2867 vdd.n2735 39.2114
R19502 vdd.n2871 vdd.n2736 39.2114
R19503 vdd.n2875 vdd.n2737 39.2114
R19504 vdd.n2879 vdd.n2738 39.2114
R19505 vdd.n2883 vdd.n2739 39.2114
R19506 vdd.n2887 vdd.n2740 39.2114
R19507 vdd.n2892 vdd.n2741 39.2114
R19508 vdd.n2895 vdd.n2742 39.2114
R19509 vdd.n3179 vdd.n3178 39.2114
R19510 vdd.n835 vdd.n831 39.2114
R19511 vdd.n3187 vdd.n3186 39.2114
R19512 vdd.n830 vdd.n828 39.2114
R19513 vdd.n3194 vdd.n3193 39.2114
R19514 vdd.n827 vdd.n825 39.2114
R19515 vdd.n3201 vdd.n3200 39.2114
R19516 vdd.n824 vdd.n822 39.2114
R19517 vdd.n3208 vdd.n3207 39.2114
R19518 vdd.n3212 vdd.n3211 39.2114
R19519 vdd.n821 vdd.n819 39.2114
R19520 vdd.n3219 vdd.n3218 39.2114
R19521 vdd.n818 vdd.n816 39.2114
R19522 vdd.n3226 vdd.n3225 39.2114
R19523 vdd.n815 vdd.n813 39.2114
R19524 vdd.n3233 vdd.n3232 39.2114
R19525 vdd.n3236 vdd.n3235 39.2114
R19526 vdd.n995 vdd.n950 39.2114
R19527 vdd.n2648 vdd.n951 39.2114
R19528 vdd.n2644 vdd.n952 39.2114
R19529 vdd.n2640 vdd.n953 39.2114
R19530 vdd.n2636 vdd.n954 39.2114
R19531 vdd.n2632 vdd.n955 39.2114
R19532 vdd.n2628 vdd.n956 39.2114
R19533 vdd.n2624 vdd.n957 39.2114
R19534 vdd.n2620 vdd.n958 39.2114
R19535 vdd.n2616 vdd.n959 39.2114
R19536 vdd.n2612 vdd.n960 39.2114
R19537 vdd.n2608 vdd.n961 39.2114
R19538 vdd.n2604 vdd.n962 39.2114
R19539 vdd.n2600 vdd.n963 39.2114
R19540 vdd.n2596 vdd.n964 39.2114
R19541 vdd.n2592 vdd.n965 39.2114
R19542 vdd.n2588 vdd.n966 39.2114
R19543 vdd.n2215 vdd.n1109 39.2114
R19544 vdd.n2218 vdd.n2217 39.2114
R19545 vdd.n2223 vdd.n2222 39.2114
R19546 vdd.n2226 vdd.n2225 39.2114
R19547 vdd.n2231 vdd.n2230 39.2114
R19548 vdd.n2234 vdd.n2233 39.2114
R19549 vdd.n2239 vdd.n2238 39.2114
R19550 vdd.n2242 vdd.n2241 39.2114
R19551 vdd.n2247 vdd.n2246 39.2114
R19552 vdd.n2250 vdd.n2249 39.2114
R19553 vdd.n2255 vdd.n2254 39.2114
R19554 vdd.n2258 vdd.n2257 39.2114
R19555 vdd.n2263 vdd.n2262 39.2114
R19556 vdd.n2266 vdd.n2265 39.2114
R19557 vdd.n2271 vdd.n2270 39.2114
R19558 vdd.n2274 vdd.n2273 39.2114
R19559 vdd.n2280 vdd.n2279 39.2114
R19560 vdd.n2585 vdd.n966 39.2114
R19561 vdd.n2589 vdd.n965 39.2114
R19562 vdd.n2593 vdd.n964 39.2114
R19563 vdd.n2597 vdd.n963 39.2114
R19564 vdd.n2601 vdd.n962 39.2114
R19565 vdd.n2605 vdd.n961 39.2114
R19566 vdd.n2609 vdd.n960 39.2114
R19567 vdd.n2613 vdd.n959 39.2114
R19568 vdd.n2617 vdd.n958 39.2114
R19569 vdd.n2621 vdd.n957 39.2114
R19570 vdd.n2625 vdd.n956 39.2114
R19571 vdd.n2629 vdd.n955 39.2114
R19572 vdd.n2633 vdd.n954 39.2114
R19573 vdd.n2637 vdd.n953 39.2114
R19574 vdd.n2641 vdd.n952 39.2114
R19575 vdd.n2645 vdd.n951 39.2114
R19576 vdd.n2649 vdd.n950 39.2114
R19577 vdd.n2216 vdd.n2215 39.2114
R19578 vdd.n2217 vdd.n2213 39.2114
R19579 vdd.n2224 vdd.n2223 39.2114
R19580 vdd.n2225 vdd.n2211 39.2114
R19581 vdd.n2232 vdd.n2231 39.2114
R19582 vdd.n2233 vdd.n2209 39.2114
R19583 vdd.n2240 vdd.n2239 39.2114
R19584 vdd.n2241 vdd.n2207 39.2114
R19585 vdd.n2248 vdd.n2247 39.2114
R19586 vdd.n2249 vdd.n1143 39.2114
R19587 vdd.n2256 vdd.n2255 39.2114
R19588 vdd.n2257 vdd.n1141 39.2114
R19589 vdd.n2264 vdd.n2263 39.2114
R19590 vdd.n2265 vdd.n1139 39.2114
R19591 vdd.n2272 vdd.n2271 39.2114
R19592 vdd.n2273 vdd.n1135 39.2114
R19593 vdd.n2281 vdd.n2280 39.2114
R19594 vdd.n2202 vdd.n2201 37.2369
R19595 vdd.n2118 vdd.n2051 37.2369
R19596 vdd.n2157 vdd.n2011 37.2369
R19597 vdd.n3320 vdd.n769 37.2369
R19598 vdd.n3368 vdd.n3367 37.2369
R19599 vdd.n690 vdd.n689 37.2369
R19600 vdd.n2277 vdd.n1137 30.449
R19601 vdd.n999 vdd.n998 30.449
R19602 vdd.n2402 vdd.n1131 30.449
R19603 vdd.n2662 vdd.n989 30.449
R19604 vdd.n2763 vdd.n2762 30.449
R19605 vdd.n3182 vdd.n833 30.449
R19606 vdd.n2890 vdd.n2831 30.449
R19607 vdd.n801 vdd.n800 30.449
R19608 vdd.n2465 vdd.n2464 30.4395
R19609 vdd.n2724 vdd.n987 30.4395
R19610 vdd.n2657 vdd.n990 30.4395
R19611 vdd.n2395 vdd.n2394 30.4395
R19612 vdd.n2897 vdd.n2896 30.4395
R19613 vdd.n3176 vdd.n3175 30.4395
R19614 vdd.n3015 vdd.n3014 30.4395
R19615 vdd.n3239 vdd.n3238 30.4395
R19616 vdd.n3158 vdd.n3157 30.4395
R19617 vdd.n3244 vdd.n802 30.4395
R19618 vdd.n3008 vdd.n3007 30.4395
R19619 vdd.n3019 vdd.n942 30.4395
R19620 vdd.n2469 vdd.n1108 30.4395
R19621 vdd.n2652 vdd.n2651 30.4395
R19622 vdd.n2584 vdd.n2583 30.4395
R19623 vdd.n2284 vdd.n2283 30.4395
R19624 vdd.n1498 vdd.n1305 22.2201
R19625 vdd.n2196 vdd.n1153 22.2201
R19626 vdd.n3405 vdd.n723 22.2201
R19627 vdd.n3537 vdd.n3536 22.2201
R19628 vdd.n1509 vdd.n1267 19.3944
R19629 vdd.n1509 vdd.n1265 19.3944
R19630 vdd.n1513 vdd.n1265 19.3944
R19631 vdd.n1513 vdd.n1255 19.3944
R19632 vdd.n1526 vdd.n1255 19.3944
R19633 vdd.n1526 vdd.n1253 19.3944
R19634 vdd.n1530 vdd.n1253 19.3944
R19635 vdd.n1530 vdd.n1245 19.3944
R19636 vdd.n1543 vdd.n1245 19.3944
R19637 vdd.n1543 vdd.n1243 19.3944
R19638 vdd.n1547 vdd.n1243 19.3944
R19639 vdd.n1547 vdd.n1232 19.3944
R19640 vdd.n1559 vdd.n1232 19.3944
R19641 vdd.n1559 vdd.n1230 19.3944
R19642 vdd.n1563 vdd.n1230 19.3944
R19643 vdd.n1563 vdd.n1221 19.3944
R19644 vdd.n1576 vdd.n1221 19.3944
R19645 vdd.n1576 vdd.n1219 19.3944
R19646 vdd.n1580 vdd.n1219 19.3944
R19647 vdd.n1580 vdd.n1210 19.3944
R19648 vdd.n1899 vdd.n1210 19.3944
R19649 vdd.n1899 vdd.n1208 19.3944
R19650 vdd.n1903 vdd.n1208 19.3944
R19651 vdd.n1903 vdd.n1198 19.3944
R19652 vdd.n1916 vdd.n1198 19.3944
R19653 vdd.n1916 vdd.n1196 19.3944
R19654 vdd.n1920 vdd.n1196 19.3944
R19655 vdd.n1920 vdd.n1188 19.3944
R19656 vdd.n1933 vdd.n1188 19.3944
R19657 vdd.n1933 vdd.n1186 19.3944
R19658 vdd.n1937 vdd.n1186 19.3944
R19659 vdd.n1937 vdd.n1175 19.3944
R19660 vdd.n1949 vdd.n1175 19.3944
R19661 vdd.n1949 vdd.n1173 19.3944
R19662 vdd.n1953 vdd.n1173 19.3944
R19663 vdd.n1953 vdd.n1165 19.3944
R19664 vdd.n1966 vdd.n1165 19.3944
R19665 vdd.n1966 vdd.n1162 19.3944
R19666 vdd.n1972 vdd.n1162 19.3944
R19667 vdd.n1972 vdd.n1163 19.3944
R19668 vdd.n1163 vdd.n1152 19.3944
R19669 vdd.n1433 vdd.n1368 19.3944
R19670 vdd.n1429 vdd.n1368 19.3944
R19671 vdd.n1429 vdd.n1428 19.3944
R19672 vdd.n1428 vdd.n1427 19.3944
R19673 vdd.n1427 vdd.n1374 19.3944
R19674 vdd.n1423 vdd.n1374 19.3944
R19675 vdd.n1423 vdd.n1422 19.3944
R19676 vdd.n1422 vdd.n1421 19.3944
R19677 vdd.n1421 vdd.n1380 19.3944
R19678 vdd.n1417 vdd.n1380 19.3944
R19679 vdd.n1417 vdd.n1416 19.3944
R19680 vdd.n1416 vdd.n1415 19.3944
R19681 vdd.n1415 vdd.n1386 19.3944
R19682 vdd.n1411 vdd.n1386 19.3944
R19683 vdd.n1411 vdd.n1410 19.3944
R19684 vdd.n1410 vdd.n1409 19.3944
R19685 vdd.n1409 vdd.n1392 19.3944
R19686 vdd.n1405 vdd.n1392 19.3944
R19687 vdd.n1405 vdd.n1404 19.3944
R19688 vdd.n1404 vdd.n1403 19.3944
R19689 vdd.n1468 vdd.n1467 19.3944
R19690 vdd.n1467 vdd.n1466 19.3944
R19691 vdd.n1466 vdd.n1339 19.3944
R19692 vdd.n1462 vdd.n1339 19.3944
R19693 vdd.n1462 vdd.n1461 19.3944
R19694 vdd.n1461 vdd.n1460 19.3944
R19695 vdd.n1460 vdd.n1345 19.3944
R19696 vdd.n1456 vdd.n1345 19.3944
R19697 vdd.n1456 vdd.n1455 19.3944
R19698 vdd.n1455 vdd.n1454 19.3944
R19699 vdd.n1454 vdd.n1351 19.3944
R19700 vdd.n1450 vdd.n1351 19.3944
R19701 vdd.n1450 vdd.n1449 19.3944
R19702 vdd.n1449 vdd.n1448 19.3944
R19703 vdd.n1448 vdd.n1357 19.3944
R19704 vdd.n1444 vdd.n1357 19.3944
R19705 vdd.n1444 vdd.n1443 19.3944
R19706 vdd.n1443 vdd.n1442 19.3944
R19707 vdd.n1442 vdd.n1363 19.3944
R19708 vdd.n1438 vdd.n1363 19.3944
R19709 vdd.n1501 vdd.n1272 19.3944
R19710 vdd.n1496 vdd.n1272 19.3944
R19711 vdd.n1496 vdd.n1307 19.3944
R19712 vdd.n1492 vdd.n1307 19.3944
R19713 vdd.n1492 vdd.n1491 19.3944
R19714 vdd.n1491 vdd.n1490 19.3944
R19715 vdd.n1490 vdd.n1313 19.3944
R19716 vdd.n1486 vdd.n1313 19.3944
R19717 vdd.n1486 vdd.n1485 19.3944
R19718 vdd.n1485 vdd.n1484 19.3944
R19719 vdd.n1484 vdd.n1319 19.3944
R19720 vdd.n1480 vdd.n1319 19.3944
R19721 vdd.n1480 vdd.n1479 19.3944
R19722 vdd.n1479 vdd.n1478 19.3944
R19723 vdd.n1478 vdd.n1325 19.3944
R19724 vdd.n1474 vdd.n1325 19.3944
R19725 vdd.n1474 vdd.n1473 19.3944
R19726 vdd.n1473 vdd.n1472 19.3944
R19727 vdd.n2114 vdd.n2049 19.3944
R19728 vdd.n2114 vdd.n2055 19.3944
R19729 vdd.n2109 vdd.n2055 19.3944
R19730 vdd.n2109 vdd.n2108 19.3944
R19731 vdd.n2108 vdd.n2107 19.3944
R19732 vdd.n2107 vdd.n2062 19.3944
R19733 vdd.n2102 vdd.n2062 19.3944
R19734 vdd.n2102 vdd.n2101 19.3944
R19735 vdd.n2101 vdd.n2100 19.3944
R19736 vdd.n2100 vdd.n2069 19.3944
R19737 vdd.n2095 vdd.n2069 19.3944
R19738 vdd.n2095 vdd.n2094 19.3944
R19739 vdd.n2094 vdd.n2093 19.3944
R19740 vdd.n2093 vdd.n2077 19.3944
R19741 vdd.n2088 vdd.n2077 19.3944
R19742 vdd.n2088 vdd.n2087 19.3944
R19743 vdd.n2083 vdd.n2082 19.3944
R19744 vdd.n2203 vdd.n1148 19.3944
R19745 vdd.n2153 vdd.n2009 19.3944
R19746 vdd.n2153 vdd.n2015 19.3944
R19747 vdd.n2148 vdd.n2015 19.3944
R19748 vdd.n2148 vdd.n2147 19.3944
R19749 vdd.n2147 vdd.n2146 19.3944
R19750 vdd.n2146 vdd.n2022 19.3944
R19751 vdd.n2141 vdd.n2022 19.3944
R19752 vdd.n2141 vdd.n2140 19.3944
R19753 vdd.n2140 vdd.n2139 19.3944
R19754 vdd.n2139 vdd.n2029 19.3944
R19755 vdd.n2134 vdd.n2029 19.3944
R19756 vdd.n2134 vdd.n2133 19.3944
R19757 vdd.n2133 vdd.n2132 19.3944
R19758 vdd.n2132 vdd.n2036 19.3944
R19759 vdd.n2127 vdd.n2036 19.3944
R19760 vdd.n2127 vdd.n2126 19.3944
R19761 vdd.n2126 vdd.n2125 19.3944
R19762 vdd.n2125 vdd.n2043 19.3944
R19763 vdd.n2120 vdd.n2043 19.3944
R19764 vdd.n2120 vdd.n2119 19.3944
R19765 vdd.n2191 vdd.n2190 19.3944
R19766 vdd.n2190 vdd.n1981 19.3944
R19767 vdd.n2185 vdd.n2184 19.3944
R19768 vdd.n2180 vdd.n1985 19.3944
R19769 vdd.n2180 vdd.n1987 19.3944
R19770 vdd.n1990 vdd.n1987 19.3944
R19771 vdd.n2173 vdd.n1990 19.3944
R19772 vdd.n2173 vdd.n2172 19.3944
R19773 vdd.n2172 vdd.n2171 19.3944
R19774 vdd.n2171 vdd.n1996 19.3944
R19775 vdd.n2166 vdd.n1996 19.3944
R19776 vdd.n2166 vdd.n2165 19.3944
R19777 vdd.n2165 vdd.n2164 19.3944
R19778 vdd.n2164 vdd.n2003 19.3944
R19779 vdd.n2159 vdd.n2003 19.3944
R19780 vdd.n2159 vdd.n2158 19.3944
R19781 vdd.n1505 vdd.n1270 19.3944
R19782 vdd.n1505 vdd.n1261 19.3944
R19783 vdd.n1518 vdd.n1261 19.3944
R19784 vdd.n1518 vdd.n1259 19.3944
R19785 vdd.n1522 vdd.n1259 19.3944
R19786 vdd.n1522 vdd.n1250 19.3944
R19787 vdd.n1535 vdd.n1250 19.3944
R19788 vdd.n1535 vdd.n1248 19.3944
R19789 vdd.n1539 vdd.n1248 19.3944
R19790 vdd.n1539 vdd.n1239 19.3944
R19791 vdd.n1551 vdd.n1239 19.3944
R19792 vdd.n1551 vdd.n1237 19.3944
R19793 vdd.n1555 vdd.n1237 19.3944
R19794 vdd.n1555 vdd.n1227 19.3944
R19795 vdd.n1568 vdd.n1227 19.3944
R19796 vdd.n1568 vdd.n1225 19.3944
R19797 vdd.n1572 vdd.n1225 19.3944
R19798 vdd.n1572 vdd.n1216 19.3944
R19799 vdd.n1584 vdd.n1216 19.3944
R19800 vdd.n1584 vdd.n1214 19.3944
R19801 vdd.n1895 vdd.n1214 19.3944
R19802 vdd.n1895 vdd.n1204 19.3944
R19803 vdd.n1908 vdd.n1204 19.3944
R19804 vdd.n1908 vdd.n1202 19.3944
R19805 vdd.n1912 vdd.n1202 19.3944
R19806 vdd.n1912 vdd.n1193 19.3944
R19807 vdd.n1925 vdd.n1193 19.3944
R19808 vdd.n1925 vdd.n1191 19.3944
R19809 vdd.n1929 vdd.n1191 19.3944
R19810 vdd.n1929 vdd.n1182 19.3944
R19811 vdd.n1941 vdd.n1182 19.3944
R19812 vdd.n1941 vdd.n1180 19.3944
R19813 vdd.n1945 vdd.n1180 19.3944
R19814 vdd.n1945 vdd.n1170 19.3944
R19815 vdd.n1958 vdd.n1170 19.3944
R19816 vdd.n1958 vdd.n1168 19.3944
R19817 vdd.n1962 vdd.n1168 19.3944
R19818 vdd.n1962 vdd.n1158 19.3944
R19819 vdd.n1977 vdd.n1158 19.3944
R19820 vdd.n1977 vdd.n1156 19.3944
R19821 vdd.n2194 vdd.n1156 19.3944
R19822 vdd.n3411 vdd.n686 19.3944
R19823 vdd.n3411 vdd.n676 19.3944
R19824 vdd.n3423 vdd.n676 19.3944
R19825 vdd.n3423 vdd.n674 19.3944
R19826 vdd.n3427 vdd.n674 19.3944
R19827 vdd.n3427 vdd.n666 19.3944
R19828 vdd.n3440 vdd.n666 19.3944
R19829 vdd.n3440 vdd.n664 19.3944
R19830 vdd.n3444 vdd.n664 19.3944
R19831 vdd.n3444 vdd.n653 19.3944
R19832 vdd.n3456 vdd.n653 19.3944
R19833 vdd.n3456 vdd.n651 19.3944
R19834 vdd.n3460 vdd.n651 19.3944
R19835 vdd.n3460 vdd.n642 19.3944
R19836 vdd.n3473 vdd.n642 19.3944
R19837 vdd.n3473 vdd.n640 19.3944
R19838 vdd.n3480 vdd.n640 19.3944
R19839 vdd.n3480 vdd.n3479 19.3944
R19840 vdd.n3479 vdd.n631 19.3944
R19841 vdd.n3493 vdd.n631 19.3944
R19842 vdd.n3494 vdd.n3493 19.3944
R19843 vdd.n3494 vdd.n629 19.3944
R19844 vdd.n3498 vdd.n629 19.3944
R19845 vdd.n3500 vdd.n3498 19.3944
R19846 vdd.n3501 vdd.n3500 19.3944
R19847 vdd.n3501 vdd.n627 19.3944
R19848 vdd.n3505 vdd.n627 19.3944
R19849 vdd.n3507 vdd.n3505 19.3944
R19850 vdd.n3508 vdd.n3507 19.3944
R19851 vdd.n3508 vdd.n625 19.3944
R19852 vdd.n3512 vdd.n625 19.3944
R19853 vdd.n3515 vdd.n3512 19.3944
R19854 vdd.n3516 vdd.n3515 19.3944
R19855 vdd.n3516 vdd.n623 19.3944
R19856 vdd.n3520 vdd.n623 19.3944
R19857 vdd.n3522 vdd.n3520 19.3944
R19858 vdd.n3523 vdd.n3522 19.3944
R19859 vdd.n3523 vdd.n621 19.3944
R19860 vdd.n3527 vdd.n621 19.3944
R19861 vdd.n3529 vdd.n3527 19.3944
R19862 vdd.n3530 vdd.n3529 19.3944
R19863 vdd.n569 vdd.n438 19.3944
R19864 vdd.n575 vdd.n438 19.3944
R19865 vdd.n576 vdd.n575 19.3944
R19866 vdd.n579 vdd.n576 19.3944
R19867 vdd.n579 vdd.n436 19.3944
R19868 vdd.n585 vdd.n436 19.3944
R19869 vdd.n586 vdd.n585 19.3944
R19870 vdd.n589 vdd.n586 19.3944
R19871 vdd.n589 vdd.n434 19.3944
R19872 vdd.n595 vdd.n434 19.3944
R19873 vdd.n596 vdd.n595 19.3944
R19874 vdd.n599 vdd.n596 19.3944
R19875 vdd.n599 vdd.n432 19.3944
R19876 vdd.n605 vdd.n432 19.3944
R19877 vdd.n606 vdd.n605 19.3944
R19878 vdd.n609 vdd.n606 19.3944
R19879 vdd.n609 vdd.n430 19.3944
R19880 vdd.n615 vdd.n430 19.3944
R19881 vdd.n617 vdd.n615 19.3944
R19882 vdd.n618 vdd.n617 19.3944
R19883 vdd.n516 vdd.n515 19.3944
R19884 vdd.n519 vdd.n516 19.3944
R19885 vdd.n519 vdd.n450 19.3944
R19886 vdd.n525 vdd.n450 19.3944
R19887 vdd.n526 vdd.n525 19.3944
R19888 vdd.n529 vdd.n526 19.3944
R19889 vdd.n529 vdd.n448 19.3944
R19890 vdd.n535 vdd.n448 19.3944
R19891 vdd.n536 vdd.n535 19.3944
R19892 vdd.n539 vdd.n536 19.3944
R19893 vdd.n539 vdd.n446 19.3944
R19894 vdd.n545 vdd.n446 19.3944
R19895 vdd.n546 vdd.n545 19.3944
R19896 vdd.n549 vdd.n546 19.3944
R19897 vdd.n549 vdd.n444 19.3944
R19898 vdd.n555 vdd.n444 19.3944
R19899 vdd.n556 vdd.n555 19.3944
R19900 vdd.n559 vdd.n556 19.3944
R19901 vdd.n559 vdd.n442 19.3944
R19902 vdd.n565 vdd.n442 19.3944
R19903 vdd.n466 vdd.n465 19.3944
R19904 vdd.n469 vdd.n466 19.3944
R19905 vdd.n469 vdd.n462 19.3944
R19906 vdd.n475 vdd.n462 19.3944
R19907 vdd.n476 vdd.n475 19.3944
R19908 vdd.n479 vdd.n476 19.3944
R19909 vdd.n479 vdd.n460 19.3944
R19910 vdd.n485 vdd.n460 19.3944
R19911 vdd.n486 vdd.n485 19.3944
R19912 vdd.n489 vdd.n486 19.3944
R19913 vdd.n489 vdd.n458 19.3944
R19914 vdd.n495 vdd.n458 19.3944
R19915 vdd.n496 vdd.n495 19.3944
R19916 vdd.n499 vdd.n496 19.3944
R19917 vdd.n499 vdd.n456 19.3944
R19918 vdd.n505 vdd.n456 19.3944
R19919 vdd.n506 vdd.n505 19.3944
R19920 vdd.n509 vdd.n506 19.3944
R19921 vdd.n3415 vdd.n683 19.3944
R19922 vdd.n3415 vdd.n681 19.3944
R19923 vdd.n3419 vdd.n681 19.3944
R19924 vdd.n3419 vdd.n671 19.3944
R19925 vdd.n3432 vdd.n671 19.3944
R19926 vdd.n3432 vdd.n669 19.3944
R19927 vdd.n3436 vdd.n669 19.3944
R19928 vdd.n3436 vdd.n660 19.3944
R19929 vdd.n3448 vdd.n660 19.3944
R19930 vdd.n3448 vdd.n658 19.3944
R19931 vdd.n3452 vdd.n658 19.3944
R19932 vdd.n3452 vdd.n648 19.3944
R19933 vdd.n3465 vdd.n648 19.3944
R19934 vdd.n3465 vdd.n646 19.3944
R19935 vdd.n3469 vdd.n646 19.3944
R19936 vdd.n3469 vdd.n637 19.3944
R19937 vdd.n3484 vdd.n637 19.3944
R19938 vdd.n3484 vdd.n635 19.3944
R19939 vdd.n3488 vdd.n635 19.3944
R19940 vdd.n3488 vdd.n336 19.3944
R19941 vdd.n3579 vdd.n336 19.3944
R19942 vdd.n3579 vdd.n337 19.3944
R19943 vdd.n3573 vdd.n337 19.3944
R19944 vdd.n3573 vdd.n3572 19.3944
R19945 vdd.n3572 vdd.n3571 19.3944
R19946 vdd.n3571 vdd.n349 19.3944
R19947 vdd.n3565 vdd.n349 19.3944
R19948 vdd.n3565 vdd.n3564 19.3944
R19949 vdd.n3564 vdd.n3563 19.3944
R19950 vdd.n3563 vdd.n359 19.3944
R19951 vdd.n3557 vdd.n359 19.3944
R19952 vdd.n3557 vdd.n3556 19.3944
R19953 vdd.n3556 vdd.n3555 19.3944
R19954 vdd.n3555 vdd.n370 19.3944
R19955 vdd.n3549 vdd.n370 19.3944
R19956 vdd.n3549 vdd.n3548 19.3944
R19957 vdd.n3548 vdd.n3547 19.3944
R19958 vdd.n3547 vdd.n381 19.3944
R19959 vdd.n3541 vdd.n381 19.3944
R19960 vdd.n3541 vdd.n3540 19.3944
R19961 vdd.n3540 vdd.n3539 19.3944
R19962 vdd.n3362 vdd.n747 19.3944
R19963 vdd.n3362 vdd.n3359 19.3944
R19964 vdd.n3359 vdd.n3356 19.3944
R19965 vdd.n3356 vdd.n3355 19.3944
R19966 vdd.n3355 vdd.n3352 19.3944
R19967 vdd.n3352 vdd.n3351 19.3944
R19968 vdd.n3351 vdd.n3348 19.3944
R19969 vdd.n3348 vdd.n3347 19.3944
R19970 vdd.n3347 vdd.n3344 19.3944
R19971 vdd.n3344 vdd.n3343 19.3944
R19972 vdd.n3343 vdd.n3340 19.3944
R19973 vdd.n3340 vdd.n3339 19.3944
R19974 vdd.n3339 vdd.n3336 19.3944
R19975 vdd.n3336 vdd.n3335 19.3944
R19976 vdd.n3335 vdd.n3332 19.3944
R19977 vdd.n3332 vdd.n3331 19.3944
R19978 vdd.n3331 vdd.n3328 19.3944
R19979 vdd.n3328 vdd.n3327 19.3944
R19980 vdd.n3327 vdd.n3324 19.3944
R19981 vdd.n3324 vdd.n3323 19.3944
R19982 vdd.n3402 vdd.n3401 19.3944
R19983 vdd.n3401 vdd.n3400 19.3944
R19984 vdd.n732 vdd.n729 19.3944
R19985 vdd.n3396 vdd.n3395 19.3944
R19986 vdd.n3395 vdd.n3392 19.3944
R19987 vdd.n3392 vdd.n3391 19.3944
R19988 vdd.n3391 vdd.n3388 19.3944
R19989 vdd.n3388 vdd.n3387 19.3944
R19990 vdd.n3387 vdd.n3384 19.3944
R19991 vdd.n3384 vdd.n3383 19.3944
R19992 vdd.n3383 vdd.n3380 19.3944
R19993 vdd.n3380 vdd.n3379 19.3944
R19994 vdd.n3379 vdd.n3376 19.3944
R19995 vdd.n3376 vdd.n3375 19.3944
R19996 vdd.n3375 vdd.n3372 19.3944
R19997 vdd.n3372 vdd.n3371 19.3944
R19998 vdd.n3316 vdd.n767 19.3944
R19999 vdd.n3316 vdd.n3313 19.3944
R20000 vdd.n3313 vdd.n3310 19.3944
R20001 vdd.n3310 vdd.n3309 19.3944
R20002 vdd.n3309 vdd.n3306 19.3944
R20003 vdd.n3306 vdd.n3305 19.3944
R20004 vdd.n3305 vdd.n3302 19.3944
R20005 vdd.n3302 vdd.n3301 19.3944
R20006 vdd.n3301 vdd.n3298 19.3944
R20007 vdd.n3298 vdd.n3297 19.3944
R20008 vdd.n3297 vdd.n3294 19.3944
R20009 vdd.n3294 vdd.n3293 19.3944
R20010 vdd.n3293 vdd.n3290 19.3944
R20011 vdd.n3290 vdd.n3289 19.3944
R20012 vdd.n3289 vdd.n3286 19.3944
R20013 vdd.n3286 vdd.n3285 19.3944
R20014 vdd.n3282 vdd.n3281 19.3944
R20015 vdd.n3278 vdd.n3277 19.3944
R20016 vdd.n1437 vdd.n1433 19.0066
R20017 vdd.n2118 vdd.n2049 19.0066
R20018 vdd.n569 vdd.n566 19.0066
R20019 vdd.n3320 vdd.n767 19.0066
R20020 vdd.n1137 vdd.n1136 16.0975
R20021 vdd.n998 vdd.n997 16.0975
R20022 vdd.n1398 vdd.n1397 16.0975
R20023 vdd.n1436 vdd.n1435 16.0975
R20024 vdd.n1332 vdd.n1331 16.0975
R20025 vdd.n2201 vdd.n2200 16.0975
R20026 vdd.n2051 vdd.n2050 16.0975
R20027 vdd.n2011 vdd.n2010 16.0975
R20028 vdd.n1131 vdd.n1130 16.0975
R20029 vdd.n989 vdd.n988 16.0975
R20030 vdd.n2762 vdd.n2761 16.0975
R20031 vdd.n427 vdd.n426 16.0975
R20032 vdd.n441 vdd.n440 16.0975
R20033 vdd.n453 vdd.n452 16.0975
R20034 vdd.n769 vdd.n768 16.0975
R20035 vdd.n3367 vdd.n3366 16.0975
R20036 vdd.n833 vdd.n832 16.0975
R20037 vdd.n2831 vdd.n2830 16.0975
R20038 vdd.n689 vdd.n688 16.0975
R20039 vdd.n800 vdd.n799 16.0975
R20040 vdd.t43 vdd.n2726 15.4182
R20041 vdd.n3010 vdd.t298 15.4182
R20042 vdd.n28 vdd.n27 14.6905
R20043 vdd.n2467 vdd.n1110 13.6043
R20044 vdd.n3241 vdd.n692 13.6043
R20045 vdd.n328 vdd.n293 13.1884
R20046 vdd.n269 vdd.n234 13.1884
R20047 vdd.n226 vdd.n191 13.1884
R20048 vdd.n167 vdd.n132 13.1884
R20049 vdd.n125 vdd.n90 13.1884
R20050 vdd.n66 vdd.n31 13.1884
R20051 vdd.n1827 vdd.n1792 13.1884
R20052 vdd.n1886 vdd.n1851 13.1884
R20053 vdd.n1725 vdd.n1690 13.1884
R20054 vdd.n1784 vdd.n1749 13.1884
R20055 vdd.n1624 vdd.n1589 13.1884
R20056 vdd.n1683 vdd.n1648 13.1884
R20057 vdd.n1468 vdd.n1333 12.9944
R20058 vdd.n1472 vdd.n1333 12.9944
R20059 vdd.n2157 vdd.n2009 12.9944
R20060 vdd.n2158 vdd.n2157 12.9944
R20061 vdd.n515 vdd.n454 12.9944
R20062 vdd.n509 vdd.n454 12.9944
R20063 vdd.n3368 vdd.n747 12.9944
R20064 vdd.n3371 vdd.n3368 12.9944
R20065 vdd.n329 vdd.n291 12.8005
R20066 vdd.n324 vdd.n295 12.8005
R20067 vdd.n270 vdd.n232 12.8005
R20068 vdd.n265 vdd.n236 12.8005
R20069 vdd.n227 vdd.n189 12.8005
R20070 vdd.n222 vdd.n193 12.8005
R20071 vdd.n168 vdd.n130 12.8005
R20072 vdd.n163 vdd.n134 12.8005
R20073 vdd.n126 vdd.n88 12.8005
R20074 vdd.n121 vdd.n92 12.8005
R20075 vdd.n67 vdd.n29 12.8005
R20076 vdd.n62 vdd.n33 12.8005
R20077 vdd.n1828 vdd.n1790 12.8005
R20078 vdd.n1823 vdd.n1794 12.8005
R20079 vdd.n1887 vdd.n1849 12.8005
R20080 vdd.n1882 vdd.n1853 12.8005
R20081 vdd.n1726 vdd.n1688 12.8005
R20082 vdd.n1721 vdd.n1692 12.8005
R20083 vdd.n1785 vdd.n1747 12.8005
R20084 vdd.n1780 vdd.n1751 12.8005
R20085 vdd.n1625 vdd.n1587 12.8005
R20086 vdd.n1620 vdd.n1591 12.8005
R20087 vdd.n1684 vdd.n1646 12.8005
R20088 vdd.n1679 vdd.n1650 12.8005
R20089 vdd.n323 vdd.n296 12.0247
R20090 vdd.n264 vdd.n237 12.0247
R20091 vdd.n221 vdd.n194 12.0247
R20092 vdd.n162 vdd.n135 12.0247
R20093 vdd.n120 vdd.n93 12.0247
R20094 vdd.n61 vdd.n34 12.0247
R20095 vdd.n1822 vdd.n1795 12.0247
R20096 vdd.n1881 vdd.n1854 12.0247
R20097 vdd.n1720 vdd.n1693 12.0247
R20098 vdd.n1779 vdd.n1752 12.0247
R20099 vdd.n1619 vdd.n1592 12.0247
R20100 vdd.n1678 vdd.n1651 12.0247
R20101 vdd.n1507 vdd.n1263 11.337
R20102 vdd.n1516 vdd.n1263 11.337
R20103 vdd.n1516 vdd.n1515 11.337
R20104 vdd.n1524 vdd.n1257 11.337
R20105 vdd.n1533 vdd.n1532 11.337
R20106 vdd.n1549 vdd.n1241 11.337
R20107 vdd.n1557 vdd.n1234 11.337
R20108 vdd.n1566 vdd.n1565 11.337
R20109 vdd.n1574 vdd.n1223 11.337
R20110 vdd.n1897 vdd.n1212 11.337
R20111 vdd.n1906 vdd.n1206 11.337
R20112 vdd.n1914 vdd.n1200 11.337
R20113 vdd.n1923 vdd.n1922 11.337
R20114 vdd.n1939 vdd.n1184 11.337
R20115 vdd.n1947 vdd.n1177 11.337
R20116 vdd.n1956 vdd.n1955 11.337
R20117 vdd.n1964 vdd.n1160 11.337
R20118 vdd.n1975 vdd.n1160 11.337
R20119 vdd.n1975 vdd.n1974 11.337
R20120 vdd.n3413 vdd.n678 11.337
R20121 vdd.n3421 vdd.n678 11.337
R20122 vdd.n3421 vdd.n679 11.337
R20123 vdd.n3430 vdd.n3429 11.337
R20124 vdd.n3446 vdd.n662 11.337
R20125 vdd.n3454 vdd.n655 11.337
R20126 vdd.n3463 vdd.n3462 11.337
R20127 vdd.n3471 vdd.n644 11.337
R20128 vdd.n3490 vdd.n633 11.337
R20129 vdd.n3577 vdd.n340 11.337
R20130 vdd.n3575 vdd.n344 11.337
R20131 vdd.n3569 vdd.n3568 11.337
R20132 vdd.n3561 vdd.n361 11.337
R20133 vdd.n3560 vdd.n3559 11.337
R20134 vdd.n3553 vdd.n3552 11.337
R20135 vdd.n3551 vdd.n375 11.337
R20136 vdd.n3545 vdd.n3544 11.337
R20137 vdd.n3544 vdd.n3543 11.337
R20138 vdd.n3543 vdd.n386 11.337
R20139 vdd.n320 vdd.n319 11.249
R20140 vdd.n261 vdd.n260 11.249
R20141 vdd.n218 vdd.n217 11.249
R20142 vdd.n159 vdd.n158 11.249
R20143 vdd.n117 vdd.n116 11.249
R20144 vdd.n58 vdd.n57 11.249
R20145 vdd.n1819 vdd.n1818 11.249
R20146 vdd.n1878 vdd.n1877 11.249
R20147 vdd.n1717 vdd.n1716 11.249
R20148 vdd.n1776 vdd.n1775 11.249
R20149 vdd.n1616 vdd.n1615 11.249
R20150 vdd.n1675 vdd.n1674 11.249
R20151 vdd.n1305 vdd.t100 11.2237
R20152 vdd.n3537 vdd.t70 11.2237
R20153 vdd.t196 vdd.n1178 10.7702
R20154 vdd.n3438 vdd.t179 10.7702
R20155 vdd.n305 vdd.n304 10.7238
R20156 vdd.n246 vdd.n245 10.7238
R20157 vdd.n203 vdd.n202 10.7238
R20158 vdd.n144 vdd.n143 10.7238
R20159 vdd.n102 vdd.n101 10.7238
R20160 vdd.n43 vdd.n42 10.7238
R20161 vdd.n1804 vdd.n1803 10.7238
R20162 vdd.n1863 vdd.n1862 10.7238
R20163 vdd.n1702 vdd.n1701 10.7238
R20164 vdd.n1761 vdd.n1760 10.7238
R20165 vdd.n1601 vdd.n1600 10.7238
R20166 vdd.n1660 vdd.n1659 10.7238
R20167 vdd.n2465 vdd.n1102 10.6151
R20168 vdd.n2475 vdd.n1102 10.6151
R20169 vdd.n2476 vdd.n2475 10.6151
R20170 vdd.n2477 vdd.n2476 10.6151
R20171 vdd.n2477 vdd.n1090 10.6151
R20172 vdd.n2487 vdd.n1090 10.6151
R20173 vdd.n2488 vdd.n2487 10.6151
R20174 vdd.n2489 vdd.n2488 10.6151
R20175 vdd.n2489 vdd.n1078 10.6151
R20176 vdd.n2499 vdd.n1078 10.6151
R20177 vdd.n2500 vdd.n2499 10.6151
R20178 vdd.n2501 vdd.n2500 10.6151
R20179 vdd.n2501 vdd.n1065 10.6151
R20180 vdd.n2511 vdd.n1065 10.6151
R20181 vdd.n2512 vdd.n2511 10.6151
R20182 vdd.n2513 vdd.n2512 10.6151
R20183 vdd.n2513 vdd.n1053 10.6151
R20184 vdd.n2524 vdd.n1053 10.6151
R20185 vdd.n2525 vdd.n2524 10.6151
R20186 vdd.n2526 vdd.n2525 10.6151
R20187 vdd.n2526 vdd.n1041 10.6151
R20188 vdd.n2536 vdd.n1041 10.6151
R20189 vdd.n2537 vdd.n2536 10.6151
R20190 vdd.n2538 vdd.n2537 10.6151
R20191 vdd.n2538 vdd.n1029 10.6151
R20192 vdd.n2548 vdd.n1029 10.6151
R20193 vdd.n2549 vdd.n2548 10.6151
R20194 vdd.n2550 vdd.n2549 10.6151
R20195 vdd.n2550 vdd.n1019 10.6151
R20196 vdd.n2560 vdd.n1019 10.6151
R20197 vdd.n2561 vdd.n2560 10.6151
R20198 vdd.n2562 vdd.n2561 10.6151
R20199 vdd.n2562 vdd.n1006 10.6151
R20200 vdd.n2574 vdd.n1006 10.6151
R20201 vdd.n2575 vdd.n2574 10.6151
R20202 vdd.n2577 vdd.n2575 10.6151
R20203 vdd.n2577 vdd.n2576 10.6151
R20204 vdd.n2576 vdd.n987 10.6151
R20205 vdd.n2724 vdd.n2723 10.6151
R20206 vdd.n2723 vdd.n2722 10.6151
R20207 vdd.n2722 vdd.n2719 10.6151
R20208 vdd.n2719 vdd.n2718 10.6151
R20209 vdd.n2718 vdd.n2715 10.6151
R20210 vdd.n2715 vdd.n2714 10.6151
R20211 vdd.n2714 vdd.n2711 10.6151
R20212 vdd.n2711 vdd.n2710 10.6151
R20213 vdd.n2710 vdd.n2707 10.6151
R20214 vdd.n2707 vdd.n2706 10.6151
R20215 vdd.n2706 vdd.n2703 10.6151
R20216 vdd.n2703 vdd.n2702 10.6151
R20217 vdd.n2702 vdd.n2699 10.6151
R20218 vdd.n2699 vdd.n2698 10.6151
R20219 vdd.n2698 vdd.n2695 10.6151
R20220 vdd.n2695 vdd.n2694 10.6151
R20221 vdd.n2694 vdd.n2691 10.6151
R20222 vdd.n2691 vdd.n2690 10.6151
R20223 vdd.n2690 vdd.n2687 10.6151
R20224 vdd.n2687 vdd.n2686 10.6151
R20225 vdd.n2686 vdd.n2683 10.6151
R20226 vdd.n2683 vdd.n2682 10.6151
R20227 vdd.n2682 vdd.n2679 10.6151
R20228 vdd.n2679 vdd.n2678 10.6151
R20229 vdd.n2678 vdd.n2675 10.6151
R20230 vdd.n2675 vdd.n2674 10.6151
R20231 vdd.n2674 vdd.n2671 10.6151
R20232 vdd.n2671 vdd.n2670 10.6151
R20233 vdd.n2670 vdd.n2667 10.6151
R20234 vdd.n2667 vdd.n2666 10.6151
R20235 vdd.n2666 vdd.n2663 10.6151
R20236 vdd.n2661 vdd.n2658 10.6151
R20237 vdd.n2658 vdd.n2657 10.6151
R20238 vdd.n2394 vdd.n2393 10.6151
R20239 vdd.n2393 vdd.n2391 10.6151
R20240 vdd.n2391 vdd.n2390 10.6151
R20241 vdd.n2390 vdd.n2388 10.6151
R20242 vdd.n2388 vdd.n2387 10.6151
R20243 vdd.n2387 vdd.n2385 10.6151
R20244 vdd.n2385 vdd.n2384 10.6151
R20245 vdd.n2384 vdd.n2382 10.6151
R20246 vdd.n2382 vdd.n2381 10.6151
R20247 vdd.n2381 vdd.n2379 10.6151
R20248 vdd.n2379 vdd.n2378 10.6151
R20249 vdd.n2378 vdd.n2376 10.6151
R20250 vdd.n2376 vdd.n2375 10.6151
R20251 vdd.n2375 vdd.n2373 10.6151
R20252 vdd.n2373 vdd.n2372 10.6151
R20253 vdd.n2372 vdd.n2370 10.6151
R20254 vdd.n2370 vdd.n2369 10.6151
R20255 vdd.n2369 vdd.n2367 10.6151
R20256 vdd.n2367 vdd.n2366 10.6151
R20257 vdd.n2366 vdd.n2364 10.6151
R20258 vdd.n2364 vdd.n2363 10.6151
R20259 vdd.n2363 vdd.n2361 10.6151
R20260 vdd.n2361 vdd.n2360 10.6151
R20261 vdd.n2360 vdd.n1133 10.6151
R20262 vdd.n2327 vdd.n1133 10.6151
R20263 vdd.n2328 vdd.n2327 10.6151
R20264 vdd.n2330 vdd.n2328 10.6151
R20265 vdd.n2331 vdd.n2330 10.6151
R20266 vdd.n2344 vdd.n2331 10.6151
R20267 vdd.n2344 vdd.n2343 10.6151
R20268 vdd.n2343 vdd.n2342 10.6151
R20269 vdd.n2342 vdd.n2340 10.6151
R20270 vdd.n2340 vdd.n2339 10.6151
R20271 vdd.n2339 vdd.n2337 10.6151
R20272 vdd.n2337 vdd.n2336 10.6151
R20273 vdd.n2336 vdd.n2333 10.6151
R20274 vdd.n2333 vdd.n2332 10.6151
R20275 vdd.n2332 vdd.n990 10.6151
R20276 vdd.n2464 vdd.n2463 10.6151
R20277 vdd.n2463 vdd.n1114 10.6151
R20278 vdd.n2458 vdd.n1114 10.6151
R20279 vdd.n2458 vdd.n2457 10.6151
R20280 vdd.n2457 vdd.n1116 10.6151
R20281 vdd.n2452 vdd.n1116 10.6151
R20282 vdd.n2452 vdd.n2451 10.6151
R20283 vdd.n2451 vdd.n2450 10.6151
R20284 vdd.n2450 vdd.n1118 10.6151
R20285 vdd.n2444 vdd.n1118 10.6151
R20286 vdd.n2444 vdd.n2443 10.6151
R20287 vdd.n2443 vdd.n2442 10.6151
R20288 vdd.n2442 vdd.n1120 10.6151
R20289 vdd.n2436 vdd.n1120 10.6151
R20290 vdd.n2436 vdd.n2435 10.6151
R20291 vdd.n2435 vdd.n2434 10.6151
R20292 vdd.n2434 vdd.n1122 10.6151
R20293 vdd.n2428 vdd.n1122 10.6151
R20294 vdd.n2428 vdd.n2427 10.6151
R20295 vdd.n2427 vdd.n2426 10.6151
R20296 vdd.n2426 vdd.n1124 10.6151
R20297 vdd.n2420 vdd.n1124 10.6151
R20298 vdd.n2420 vdd.n2419 10.6151
R20299 vdd.n2419 vdd.n2418 10.6151
R20300 vdd.n2418 vdd.n1126 10.6151
R20301 vdd.n2412 vdd.n1126 10.6151
R20302 vdd.n2412 vdd.n2411 10.6151
R20303 vdd.n2411 vdd.n2410 10.6151
R20304 vdd.n2410 vdd.n1128 10.6151
R20305 vdd.n2404 vdd.n1128 10.6151
R20306 vdd.n2404 vdd.n2403 10.6151
R20307 vdd.n2401 vdd.n1132 10.6151
R20308 vdd.n2395 vdd.n1132 10.6151
R20309 vdd.n2899 vdd.n2897 10.6151
R20310 vdd.n2900 vdd.n2899 10.6151
R20311 vdd.n2999 vdd.n2900 10.6151
R20312 vdd.n2999 vdd.n2998 10.6151
R20313 vdd.n2998 vdd.n2997 10.6151
R20314 vdd.n2997 vdd.n2995 10.6151
R20315 vdd.n2995 vdd.n2994 10.6151
R20316 vdd.n2994 vdd.n2992 10.6151
R20317 vdd.n2992 vdd.n2991 10.6151
R20318 vdd.n2991 vdd.n2901 10.6151
R20319 vdd.n2941 vdd.n2901 10.6151
R20320 vdd.n2942 vdd.n2941 10.6151
R20321 vdd.n2944 vdd.n2942 10.6151
R20322 vdd.n2945 vdd.n2944 10.6151
R20323 vdd.n2975 vdd.n2945 10.6151
R20324 vdd.n2975 vdd.n2974 10.6151
R20325 vdd.n2974 vdd.n2973 10.6151
R20326 vdd.n2973 vdd.n2971 10.6151
R20327 vdd.n2971 vdd.n2970 10.6151
R20328 vdd.n2970 vdd.n2968 10.6151
R20329 vdd.n2968 vdd.n2967 10.6151
R20330 vdd.n2967 vdd.n2965 10.6151
R20331 vdd.n2965 vdd.n2964 10.6151
R20332 vdd.n2964 vdd.n2962 10.6151
R20333 vdd.n2962 vdd.n2961 10.6151
R20334 vdd.n2961 vdd.n2959 10.6151
R20335 vdd.n2959 vdd.n2958 10.6151
R20336 vdd.n2958 vdd.n2956 10.6151
R20337 vdd.n2956 vdd.n2955 10.6151
R20338 vdd.n2955 vdd.n2953 10.6151
R20339 vdd.n2953 vdd.n2952 10.6151
R20340 vdd.n2952 vdd.n2950 10.6151
R20341 vdd.n2950 vdd.n2949 10.6151
R20342 vdd.n2949 vdd.n2947 10.6151
R20343 vdd.n2947 vdd.n2946 10.6151
R20344 vdd.n2946 vdd.n836 10.6151
R20345 vdd.n3174 vdd.n836 10.6151
R20346 vdd.n3175 vdd.n3174 10.6151
R20347 vdd.n3014 vdd.n3013 10.6151
R20348 vdd.n3013 vdd.n948 10.6151
R20349 vdd.n2833 vdd.n948 10.6151
R20350 vdd.n2834 vdd.n2833 10.6151
R20351 vdd.n2837 vdd.n2834 10.6151
R20352 vdd.n2838 vdd.n2837 10.6151
R20353 vdd.n2841 vdd.n2838 10.6151
R20354 vdd.n2842 vdd.n2841 10.6151
R20355 vdd.n2845 vdd.n2842 10.6151
R20356 vdd.n2846 vdd.n2845 10.6151
R20357 vdd.n2849 vdd.n2846 10.6151
R20358 vdd.n2850 vdd.n2849 10.6151
R20359 vdd.n2853 vdd.n2850 10.6151
R20360 vdd.n2854 vdd.n2853 10.6151
R20361 vdd.n2857 vdd.n2854 10.6151
R20362 vdd.n2858 vdd.n2857 10.6151
R20363 vdd.n2861 vdd.n2858 10.6151
R20364 vdd.n2862 vdd.n2861 10.6151
R20365 vdd.n2865 vdd.n2862 10.6151
R20366 vdd.n2866 vdd.n2865 10.6151
R20367 vdd.n2869 vdd.n2866 10.6151
R20368 vdd.n2870 vdd.n2869 10.6151
R20369 vdd.n2873 vdd.n2870 10.6151
R20370 vdd.n2874 vdd.n2873 10.6151
R20371 vdd.n2877 vdd.n2874 10.6151
R20372 vdd.n2878 vdd.n2877 10.6151
R20373 vdd.n2881 vdd.n2878 10.6151
R20374 vdd.n2882 vdd.n2881 10.6151
R20375 vdd.n2885 vdd.n2882 10.6151
R20376 vdd.n2886 vdd.n2885 10.6151
R20377 vdd.n2889 vdd.n2886 10.6151
R20378 vdd.n2894 vdd.n2891 10.6151
R20379 vdd.n2896 vdd.n2894 10.6151
R20380 vdd.n3015 vdd.n937 10.6151
R20381 vdd.n3025 vdd.n937 10.6151
R20382 vdd.n3026 vdd.n3025 10.6151
R20383 vdd.n3027 vdd.n3026 10.6151
R20384 vdd.n3027 vdd.n925 10.6151
R20385 vdd.n3037 vdd.n925 10.6151
R20386 vdd.n3038 vdd.n3037 10.6151
R20387 vdd.n3039 vdd.n3038 10.6151
R20388 vdd.n3039 vdd.n915 10.6151
R20389 vdd.n3049 vdd.n915 10.6151
R20390 vdd.n3050 vdd.n3049 10.6151
R20391 vdd.n3051 vdd.n3050 10.6151
R20392 vdd.n3051 vdd.n903 10.6151
R20393 vdd.n3061 vdd.n903 10.6151
R20394 vdd.n3062 vdd.n3061 10.6151
R20395 vdd.n3063 vdd.n3062 10.6151
R20396 vdd.n3063 vdd.n892 10.6151
R20397 vdd.n3073 vdd.n892 10.6151
R20398 vdd.n3074 vdd.n3073 10.6151
R20399 vdd.n3075 vdd.n3074 10.6151
R20400 vdd.n3075 vdd.n879 10.6151
R20401 vdd.n3086 vdd.n879 10.6151
R20402 vdd.n3087 vdd.n3086 10.6151
R20403 vdd.n3088 vdd.n3087 10.6151
R20404 vdd.n3088 vdd.n866 10.6151
R20405 vdd.n3098 vdd.n866 10.6151
R20406 vdd.n3099 vdd.n3098 10.6151
R20407 vdd.n3100 vdd.n3099 10.6151
R20408 vdd.n3100 vdd.n855 10.6151
R20409 vdd.n3110 vdd.n855 10.6151
R20410 vdd.n3111 vdd.n3110 10.6151
R20411 vdd.n3112 vdd.n3111 10.6151
R20412 vdd.n3112 vdd.n841 10.6151
R20413 vdd.n3167 vdd.n841 10.6151
R20414 vdd.n3168 vdd.n3167 10.6151
R20415 vdd.n3169 vdd.n3168 10.6151
R20416 vdd.n3169 vdd.n810 10.6151
R20417 vdd.n3239 vdd.n810 10.6151
R20418 vdd.n3238 vdd.n3237 10.6151
R20419 vdd.n3237 vdd.n811 10.6151
R20420 vdd.n812 vdd.n811 10.6151
R20421 vdd.n3230 vdd.n812 10.6151
R20422 vdd.n3230 vdd.n3229 10.6151
R20423 vdd.n3229 vdd.n3228 10.6151
R20424 vdd.n3228 vdd.n814 10.6151
R20425 vdd.n3223 vdd.n814 10.6151
R20426 vdd.n3223 vdd.n3222 10.6151
R20427 vdd.n3222 vdd.n3221 10.6151
R20428 vdd.n3221 vdd.n817 10.6151
R20429 vdd.n3216 vdd.n817 10.6151
R20430 vdd.n3216 vdd.n3215 10.6151
R20431 vdd.n3215 vdd.n3214 10.6151
R20432 vdd.n3214 vdd.n820 10.6151
R20433 vdd.n3209 vdd.n820 10.6151
R20434 vdd.n3209 vdd.n731 10.6151
R20435 vdd.n3205 vdd.n731 10.6151
R20436 vdd.n3205 vdd.n3204 10.6151
R20437 vdd.n3204 vdd.n3203 10.6151
R20438 vdd.n3203 vdd.n823 10.6151
R20439 vdd.n3198 vdd.n823 10.6151
R20440 vdd.n3198 vdd.n3197 10.6151
R20441 vdd.n3197 vdd.n3196 10.6151
R20442 vdd.n3196 vdd.n826 10.6151
R20443 vdd.n3191 vdd.n826 10.6151
R20444 vdd.n3191 vdd.n3190 10.6151
R20445 vdd.n3190 vdd.n3189 10.6151
R20446 vdd.n3189 vdd.n829 10.6151
R20447 vdd.n3184 vdd.n829 10.6151
R20448 vdd.n3184 vdd.n3183 10.6151
R20449 vdd.n3181 vdd.n834 10.6151
R20450 vdd.n3176 vdd.n834 10.6151
R20451 vdd.n3157 vdd.n3118 10.6151
R20452 vdd.n3152 vdd.n3118 10.6151
R20453 vdd.n3152 vdd.n3151 10.6151
R20454 vdd.n3151 vdd.n3150 10.6151
R20455 vdd.n3150 vdd.n3120 10.6151
R20456 vdd.n3145 vdd.n3120 10.6151
R20457 vdd.n3145 vdd.n3144 10.6151
R20458 vdd.n3144 vdd.n3143 10.6151
R20459 vdd.n3143 vdd.n3123 10.6151
R20460 vdd.n3138 vdd.n3123 10.6151
R20461 vdd.n3138 vdd.n3137 10.6151
R20462 vdd.n3137 vdd.n3136 10.6151
R20463 vdd.n3136 vdd.n3126 10.6151
R20464 vdd.n3131 vdd.n3126 10.6151
R20465 vdd.n3131 vdd.n3130 10.6151
R20466 vdd.n3130 vdd.n785 10.6151
R20467 vdd.n3274 vdd.n785 10.6151
R20468 vdd.n3274 vdd.n786 10.6151
R20469 vdd.n788 vdd.n786 10.6151
R20470 vdd.n3267 vdd.n788 10.6151
R20471 vdd.n3267 vdd.n3266 10.6151
R20472 vdd.n3266 vdd.n3265 10.6151
R20473 vdd.n3265 vdd.n790 10.6151
R20474 vdd.n3260 vdd.n790 10.6151
R20475 vdd.n3260 vdd.n3259 10.6151
R20476 vdd.n3259 vdd.n3258 10.6151
R20477 vdd.n3258 vdd.n793 10.6151
R20478 vdd.n3253 vdd.n793 10.6151
R20479 vdd.n3253 vdd.n3252 10.6151
R20480 vdd.n3252 vdd.n3251 10.6151
R20481 vdd.n3251 vdd.n796 10.6151
R20482 vdd.n3246 vdd.n3245 10.6151
R20483 vdd.n3245 vdd.n3244 10.6151
R20484 vdd.n3007 vdd.n3006 10.6151
R20485 vdd.n3006 vdd.n3004 10.6151
R20486 vdd.n3004 vdd.n3003 10.6151
R20487 vdd.n3003 vdd.n2829 10.6151
R20488 vdd.n2903 vdd.n2829 10.6151
R20489 vdd.n2904 vdd.n2903 10.6151
R20490 vdd.n2906 vdd.n2904 10.6151
R20491 vdd.n2907 vdd.n2906 10.6151
R20492 vdd.n2987 vdd.n2907 10.6151
R20493 vdd.n2987 vdd.n2986 10.6151
R20494 vdd.n2986 vdd.n2985 10.6151
R20495 vdd.n2985 vdd.n2983 10.6151
R20496 vdd.n2983 vdd.n2982 10.6151
R20497 vdd.n2982 vdd.n2980 10.6151
R20498 vdd.n2980 vdd.n2979 10.6151
R20499 vdd.n2979 vdd.n2939 10.6151
R20500 vdd.n2939 vdd.n2938 10.6151
R20501 vdd.n2938 vdd.n2936 10.6151
R20502 vdd.n2936 vdd.n2935 10.6151
R20503 vdd.n2935 vdd.n2933 10.6151
R20504 vdd.n2933 vdd.n2932 10.6151
R20505 vdd.n2932 vdd.n2930 10.6151
R20506 vdd.n2930 vdd.n2929 10.6151
R20507 vdd.n2929 vdd.n2927 10.6151
R20508 vdd.n2927 vdd.n2926 10.6151
R20509 vdd.n2926 vdd.n2924 10.6151
R20510 vdd.n2924 vdd.n2923 10.6151
R20511 vdd.n2923 vdd.n2921 10.6151
R20512 vdd.n2921 vdd.n2920 10.6151
R20513 vdd.n2920 vdd.n2918 10.6151
R20514 vdd.n2918 vdd.n2917 10.6151
R20515 vdd.n2917 vdd.n2915 10.6151
R20516 vdd.n2915 vdd.n2914 10.6151
R20517 vdd.n2914 vdd.n2912 10.6151
R20518 vdd.n2912 vdd.n2911 10.6151
R20519 vdd.n2911 vdd.n2909 10.6151
R20520 vdd.n2909 vdd.n2908 10.6151
R20521 vdd.n2908 vdd.n802 10.6151
R20522 vdd.n2764 vdd.n942 10.6151
R20523 vdd.n2767 vdd.n2764 10.6151
R20524 vdd.n2768 vdd.n2767 10.6151
R20525 vdd.n2771 vdd.n2768 10.6151
R20526 vdd.n2772 vdd.n2771 10.6151
R20527 vdd.n2775 vdd.n2772 10.6151
R20528 vdd.n2776 vdd.n2775 10.6151
R20529 vdd.n2779 vdd.n2776 10.6151
R20530 vdd.n2780 vdd.n2779 10.6151
R20531 vdd.n2783 vdd.n2780 10.6151
R20532 vdd.n2784 vdd.n2783 10.6151
R20533 vdd.n2787 vdd.n2784 10.6151
R20534 vdd.n2788 vdd.n2787 10.6151
R20535 vdd.n2791 vdd.n2788 10.6151
R20536 vdd.n2792 vdd.n2791 10.6151
R20537 vdd.n2795 vdd.n2792 10.6151
R20538 vdd.n2796 vdd.n2795 10.6151
R20539 vdd.n2799 vdd.n2796 10.6151
R20540 vdd.n2800 vdd.n2799 10.6151
R20541 vdd.n2803 vdd.n2800 10.6151
R20542 vdd.n2804 vdd.n2803 10.6151
R20543 vdd.n2807 vdd.n2804 10.6151
R20544 vdd.n2808 vdd.n2807 10.6151
R20545 vdd.n2811 vdd.n2808 10.6151
R20546 vdd.n2812 vdd.n2811 10.6151
R20547 vdd.n2815 vdd.n2812 10.6151
R20548 vdd.n2816 vdd.n2815 10.6151
R20549 vdd.n2819 vdd.n2816 10.6151
R20550 vdd.n2820 vdd.n2819 10.6151
R20551 vdd.n2823 vdd.n2820 10.6151
R20552 vdd.n2824 vdd.n2823 10.6151
R20553 vdd.n2828 vdd.n2827 10.6151
R20554 vdd.n3008 vdd.n2828 10.6151
R20555 vdd.n3020 vdd.n3019 10.6151
R20556 vdd.n3021 vdd.n3020 10.6151
R20557 vdd.n3021 vdd.n932 10.6151
R20558 vdd.n3031 vdd.n932 10.6151
R20559 vdd.n3032 vdd.n3031 10.6151
R20560 vdd.n3033 vdd.n3032 10.6151
R20561 vdd.n3033 vdd.n920 10.6151
R20562 vdd.n3043 vdd.n920 10.6151
R20563 vdd.n3044 vdd.n3043 10.6151
R20564 vdd.n3045 vdd.n3044 10.6151
R20565 vdd.n3045 vdd.n909 10.6151
R20566 vdd.n3055 vdd.n909 10.6151
R20567 vdd.n3056 vdd.n3055 10.6151
R20568 vdd.n3057 vdd.n3056 10.6151
R20569 vdd.n3057 vdd.n897 10.6151
R20570 vdd.n3067 vdd.n897 10.6151
R20571 vdd.n3068 vdd.n3067 10.6151
R20572 vdd.n3069 vdd.n3068 10.6151
R20573 vdd.n3069 vdd.n886 10.6151
R20574 vdd.n3079 vdd.n886 10.6151
R20575 vdd.n3082 vdd.n3081 10.6151
R20576 vdd.n3082 vdd.n872 10.6151
R20577 vdd.n3092 vdd.n872 10.6151
R20578 vdd.n3093 vdd.n3092 10.6151
R20579 vdd.n3094 vdd.n3093 10.6151
R20580 vdd.n3094 vdd.n860 10.6151
R20581 vdd.n3104 vdd.n860 10.6151
R20582 vdd.n3105 vdd.n3104 10.6151
R20583 vdd.n3106 vdd.n3105 10.6151
R20584 vdd.n3106 vdd.n849 10.6151
R20585 vdd.n3116 vdd.n849 10.6151
R20586 vdd.n3117 vdd.n3116 10.6151
R20587 vdd.n3163 vdd.n3117 10.6151
R20588 vdd.n3163 vdd.n3162 10.6151
R20589 vdd.n3162 vdd.n3161 10.6151
R20590 vdd.n3161 vdd.n3160 10.6151
R20591 vdd.n3160 vdd.n3158 10.6151
R20592 vdd.n2470 vdd.n2469 10.6151
R20593 vdd.n2471 vdd.n2470 10.6151
R20594 vdd.n2471 vdd.n1096 10.6151
R20595 vdd.n2481 vdd.n1096 10.6151
R20596 vdd.n2482 vdd.n2481 10.6151
R20597 vdd.n2483 vdd.n2482 10.6151
R20598 vdd.n2483 vdd.n1084 10.6151
R20599 vdd.n2493 vdd.n1084 10.6151
R20600 vdd.n2494 vdd.n2493 10.6151
R20601 vdd.n2495 vdd.n2494 10.6151
R20602 vdd.n2495 vdd.n1072 10.6151
R20603 vdd.n2505 vdd.n1072 10.6151
R20604 vdd.n2506 vdd.n2505 10.6151
R20605 vdd.n2507 vdd.n2506 10.6151
R20606 vdd.n2507 vdd.n1059 10.6151
R20607 vdd.n2517 vdd.n1059 10.6151
R20608 vdd.n2518 vdd.n2517 10.6151
R20609 vdd.n2520 vdd.n1047 10.6151
R20610 vdd.n2530 vdd.n1047 10.6151
R20611 vdd.n2531 vdd.n2530 10.6151
R20612 vdd.n2532 vdd.n2531 10.6151
R20613 vdd.n2532 vdd.n1035 10.6151
R20614 vdd.n2542 vdd.n1035 10.6151
R20615 vdd.n2543 vdd.n2542 10.6151
R20616 vdd.n2544 vdd.n2543 10.6151
R20617 vdd.n2544 vdd.n1024 10.6151
R20618 vdd.n2554 vdd.n1024 10.6151
R20619 vdd.n2555 vdd.n2554 10.6151
R20620 vdd.n2556 vdd.n2555 10.6151
R20621 vdd.n2556 vdd.n1013 10.6151
R20622 vdd.n2566 vdd.n1013 10.6151
R20623 vdd.n2567 vdd.n2566 10.6151
R20624 vdd.n2570 vdd.n2567 10.6151
R20625 vdd.n2570 vdd.n2569 10.6151
R20626 vdd.n2569 vdd.n2568 10.6151
R20627 vdd.n2568 vdd.n996 10.6151
R20628 vdd.n2652 vdd.n996 10.6151
R20629 vdd.n2651 vdd.n2650 10.6151
R20630 vdd.n2650 vdd.n2647 10.6151
R20631 vdd.n2647 vdd.n2646 10.6151
R20632 vdd.n2646 vdd.n2643 10.6151
R20633 vdd.n2643 vdd.n2642 10.6151
R20634 vdd.n2642 vdd.n2639 10.6151
R20635 vdd.n2639 vdd.n2638 10.6151
R20636 vdd.n2638 vdd.n2635 10.6151
R20637 vdd.n2635 vdd.n2634 10.6151
R20638 vdd.n2634 vdd.n2631 10.6151
R20639 vdd.n2631 vdd.n2630 10.6151
R20640 vdd.n2630 vdd.n2627 10.6151
R20641 vdd.n2627 vdd.n2626 10.6151
R20642 vdd.n2626 vdd.n2623 10.6151
R20643 vdd.n2623 vdd.n2622 10.6151
R20644 vdd.n2622 vdd.n2619 10.6151
R20645 vdd.n2619 vdd.n2618 10.6151
R20646 vdd.n2618 vdd.n2615 10.6151
R20647 vdd.n2615 vdd.n2614 10.6151
R20648 vdd.n2614 vdd.n2611 10.6151
R20649 vdd.n2611 vdd.n2610 10.6151
R20650 vdd.n2610 vdd.n2607 10.6151
R20651 vdd.n2607 vdd.n2606 10.6151
R20652 vdd.n2606 vdd.n2603 10.6151
R20653 vdd.n2603 vdd.n2602 10.6151
R20654 vdd.n2602 vdd.n2599 10.6151
R20655 vdd.n2599 vdd.n2598 10.6151
R20656 vdd.n2598 vdd.n2595 10.6151
R20657 vdd.n2595 vdd.n2594 10.6151
R20658 vdd.n2594 vdd.n2591 10.6151
R20659 vdd.n2591 vdd.n2590 10.6151
R20660 vdd.n2587 vdd.n2586 10.6151
R20661 vdd.n2586 vdd.n2584 10.6151
R20662 vdd.n2286 vdd.n2284 10.6151
R20663 vdd.n2287 vdd.n2286 10.6151
R20664 vdd.n2289 vdd.n2287 10.6151
R20665 vdd.n2290 vdd.n2289 10.6151
R20666 vdd.n2292 vdd.n2290 10.6151
R20667 vdd.n2293 vdd.n2292 10.6151
R20668 vdd.n2295 vdd.n2293 10.6151
R20669 vdd.n2296 vdd.n2295 10.6151
R20670 vdd.n2298 vdd.n2296 10.6151
R20671 vdd.n2299 vdd.n2298 10.6151
R20672 vdd.n2301 vdd.n2299 10.6151
R20673 vdd.n2302 vdd.n2301 10.6151
R20674 vdd.n2304 vdd.n2302 10.6151
R20675 vdd.n2305 vdd.n2304 10.6151
R20676 vdd.n2307 vdd.n2305 10.6151
R20677 vdd.n2308 vdd.n2307 10.6151
R20678 vdd.n2310 vdd.n2308 10.6151
R20679 vdd.n2311 vdd.n2310 10.6151
R20680 vdd.n2313 vdd.n2311 10.6151
R20681 vdd.n2314 vdd.n2313 10.6151
R20682 vdd.n2316 vdd.n2314 10.6151
R20683 vdd.n2317 vdd.n2316 10.6151
R20684 vdd.n2356 vdd.n2317 10.6151
R20685 vdd.n2356 vdd.n2355 10.6151
R20686 vdd.n2355 vdd.n2354 10.6151
R20687 vdd.n2354 vdd.n2352 10.6151
R20688 vdd.n2352 vdd.n2351 10.6151
R20689 vdd.n2351 vdd.n2349 10.6151
R20690 vdd.n2349 vdd.n2348 10.6151
R20691 vdd.n2348 vdd.n2325 10.6151
R20692 vdd.n2325 vdd.n2324 10.6151
R20693 vdd.n2324 vdd.n2322 10.6151
R20694 vdd.n2322 vdd.n2321 10.6151
R20695 vdd.n2321 vdd.n2319 10.6151
R20696 vdd.n2319 vdd.n2318 10.6151
R20697 vdd.n2318 vdd.n1000 10.6151
R20698 vdd.n2582 vdd.n1000 10.6151
R20699 vdd.n2583 vdd.n2582 10.6151
R20700 vdd.n2214 vdd.n1108 10.6151
R20701 vdd.n2219 vdd.n2214 10.6151
R20702 vdd.n2220 vdd.n2219 10.6151
R20703 vdd.n2221 vdd.n2220 10.6151
R20704 vdd.n2221 vdd.n2212 10.6151
R20705 vdd.n2227 vdd.n2212 10.6151
R20706 vdd.n2228 vdd.n2227 10.6151
R20707 vdd.n2229 vdd.n2228 10.6151
R20708 vdd.n2229 vdd.n2210 10.6151
R20709 vdd.n2235 vdd.n2210 10.6151
R20710 vdd.n2236 vdd.n2235 10.6151
R20711 vdd.n2237 vdd.n2236 10.6151
R20712 vdd.n2237 vdd.n2208 10.6151
R20713 vdd.n2243 vdd.n2208 10.6151
R20714 vdd.n2244 vdd.n2243 10.6151
R20715 vdd.n2245 vdd.n2244 10.6151
R20716 vdd.n2245 vdd.n2206 10.6151
R20717 vdd.n2251 vdd.n2206 10.6151
R20718 vdd.n2252 vdd.n2251 10.6151
R20719 vdd.n2253 vdd.n2252 10.6151
R20720 vdd.n2253 vdd.n1142 10.6151
R20721 vdd.n2259 vdd.n1142 10.6151
R20722 vdd.n2260 vdd.n2259 10.6151
R20723 vdd.n2261 vdd.n2260 10.6151
R20724 vdd.n2261 vdd.n1140 10.6151
R20725 vdd.n2267 vdd.n1140 10.6151
R20726 vdd.n2268 vdd.n2267 10.6151
R20727 vdd.n2269 vdd.n2268 10.6151
R20728 vdd.n2269 vdd.n1138 10.6151
R20729 vdd.n2275 vdd.n1138 10.6151
R20730 vdd.n2276 vdd.n2275 10.6151
R20731 vdd.n2278 vdd.n1134 10.6151
R20732 vdd.n2283 vdd.n1134 10.6151
R20733 vdd.n1931 vdd.t226 10.5435
R20734 vdd.n656 vdd.t184 10.5435
R20735 vdd.n316 vdd.n298 10.4732
R20736 vdd.n257 vdd.n239 10.4732
R20737 vdd.n214 vdd.n196 10.4732
R20738 vdd.n155 vdd.n137 10.4732
R20739 vdd.n113 vdd.n95 10.4732
R20740 vdd.n54 vdd.n36 10.4732
R20741 vdd.n1815 vdd.n1797 10.4732
R20742 vdd.n1874 vdd.n1856 10.4732
R20743 vdd.n1713 vdd.n1695 10.4732
R20744 vdd.n1772 vdd.n1754 10.4732
R20745 vdd.n1612 vdd.n1594 10.4732
R20746 vdd.n1671 vdd.n1653 10.4732
R20747 vdd.t168 vdd.n1905 10.3167
R20748 vdd.n3482 vdd.t248 10.3167
R20749 vdd.n2654 vdd.t296 10.2034
R20750 vdd.n3017 vdd.t53 10.2034
R20751 vdd.n1582 vdd.t139 10.09
R20752 vdd.n3576 vdd.t202 10.09
R20753 vdd.n2182 vdd.n1122 9.88581
R20754 vdd.n3398 vdd.n731 9.88581
R20755 vdd.n3275 vdd.n3274 9.88581
R20756 vdd.n2206 vdd.n2205 9.88581
R20757 vdd.t133 vdd.n1235 9.86327
R20758 vdd.n3567 vdd.t252 9.86327
R20759 vdd.n315 vdd.n300 9.69747
R20760 vdd.n256 vdd.n241 9.69747
R20761 vdd.n213 vdd.n198 9.69747
R20762 vdd.n154 vdd.n139 9.69747
R20763 vdd.n112 vdd.n97 9.69747
R20764 vdd.n53 vdd.n38 9.69747
R20765 vdd.n1814 vdd.n1799 9.69747
R20766 vdd.n1873 vdd.n1858 9.69747
R20767 vdd.n1712 vdd.n1697 9.69747
R20768 vdd.n1771 vdd.n1756 9.69747
R20769 vdd.n1611 vdd.n1596 9.69747
R20770 vdd.n1670 vdd.n1655 9.69747
R20771 vdd.n1541 vdd.t214 9.63654
R20772 vdd.n3513 vdd.t211 9.63654
R20773 vdd.n331 vdd.n330 9.45567
R20774 vdd.n272 vdd.n271 9.45567
R20775 vdd.n229 vdd.n228 9.45567
R20776 vdd.n170 vdd.n169 9.45567
R20777 vdd.n128 vdd.n127 9.45567
R20778 vdd.n69 vdd.n68 9.45567
R20779 vdd.n1830 vdd.n1829 9.45567
R20780 vdd.n1889 vdd.n1888 9.45567
R20781 vdd.n1728 vdd.n1727 9.45567
R20782 vdd.n1787 vdd.n1786 9.45567
R20783 vdd.n1627 vdd.n1626 9.45567
R20784 vdd.n1686 vdd.n1685 9.45567
R20785 vdd.n1515 vdd.t228 9.40981
R20786 vdd.n3545 vdd.t151 9.40981
R20787 vdd.n2155 vdd.n2009 9.3005
R20788 vdd.n2154 vdd.n2153 9.3005
R20789 vdd.n2015 vdd.n2014 9.3005
R20790 vdd.n2148 vdd.n2019 9.3005
R20791 vdd.n2147 vdd.n2020 9.3005
R20792 vdd.n2146 vdd.n2021 9.3005
R20793 vdd.n2025 vdd.n2022 9.3005
R20794 vdd.n2141 vdd.n2026 9.3005
R20795 vdd.n2140 vdd.n2027 9.3005
R20796 vdd.n2139 vdd.n2028 9.3005
R20797 vdd.n2032 vdd.n2029 9.3005
R20798 vdd.n2134 vdd.n2033 9.3005
R20799 vdd.n2133 vdd.n2034 9.3005
R20800 vdd.n2132 vdd.n2035 9.3005
R20801 vdd.n2039 vdd.n2036 9.3005
R20802 vdd.n2127 vdd.n2040 9.3005
R20803 vdd.n2126 vdd.n2041 9.3005
R20804 vdd.n2125 vdd.n2042 9.3005
R20805 vdd.n2046 vdd.n2043 9.3005
R20806 vdd.n2120 vdd.n2047 9.3005
R20807 vdd.n2119 vdd.n2048 9.3005
R20808 vdd.n2118 vdd.n2117 9.3005
R20809 vdd.n2116 vdd.n2049 9.3005
R20810 vdd.n2115 vdd.n2114 9.3005
R20811 vdd.n2055 vdd.n2054 9.3005
R20812 vdd.n2109 vdd.n2059 9.3005
R20813 vdd.n2108 vdd.n2060 9.3005
R20814 vdd.n2107 vdd.n2061 9.3005
R20815 vdd.n2065 vdd.n2062 9.3005
R20816 vdd.n2102 vdd.n2066 9.3005
R20817 vdd.n2101 vdd.n2067 9.3005
R20818 vdd.n2100 vdd.n2068 9.3005
R20819 vdd.n2072 vdd.n2069 9.3005
R20820 vdd.n2095 vdd.n2073 9.3005
R20821 vdd.n2094 vdd.n2074 9.3005
R20822 vdd.n2093 vdd.n2075 9.3005
R20823 vdd.n2077 vdd.n2076 9.3005
R20824 vdd.n2088 vdd.n1144 9.3005
R20825 vdd.n2157 vdd.n2156 9.3005
R20826 vdd.n2181 vdd.n2180 9.3005
R20827 vdd.n1987 vdd.n1986 9.3005
R20828 vdd.n1992 vdd.n1990 9.3005
R20829 vdd.n2173 vdd.n1993 9.3005
R20830 vdd.n2172 vdd.n1994 9.3005
R20831 vdd.n2171 vdd.n1995 9.3005
R20832 vdd.n1999 vdd.n1996 9.3005
R20833 vdd.n2166 vdd.n2000 9.3005
R20834 vdd.n2165 vdd.n2001 9.3005
R20835 vdd.n2164 vdd.n2002 9.3005
R20836 vdd.n2006 vdd.n2003 9.3005
R20837 vdd.n2159 vdd.n2007 9.3005
R20838 vdd.n2158 vdd.n2008 9.3005
R20839 vdd.n2190 vdd.n1980 9.3005
R20840 vdd.n2192 vdd.n2191 9.3005
R20841 vdd.n1895 vdd.n1894 9.3005
R20842 vdd.n1204 vdd.n1203 9.3005
R20843 vdd.n1909 vdd.n1908 9.3005
R20844 vdd.n1910 vdd.n1202 9.3005
R20845 vdd.n1912 vdd.n1911 9.3005
R20846 vdd.n1193 vdd.n1192 9.3005
R20847 vdd.n1926 vdd.n1925 9.3005
R20848 vdd.n1927 vdd.n1191 9.3005
R20849 vdd.n1929 vdd.n1928 9.3005
R20850 vdd.n1182 vdd.n1181 9.3005
R20851 vdd.n1942 vdd.n1941 9.3005
R20852 vdd.n1943 vdd.n1180 9.3005
R20853 vdd.n1945 vdd.n1944 9.3005
R20854 vdd.n1170 vdd.n1169 9.3005
R20855 vdd.n1959 vdd.n1958 9.3005
R20856 vdd.n1960 vdd.n1168 9.3005
R20857 vdd.n1962 vdd.n1961 9.3005
R20858 vdd.n1158 vdd.n1157 9.3005
R20859 vdd.n1978 vdd.n1977 9.3005
R20860 vdd.n1979 vdd.n1156 9.3005
R20861 vdd.n2194 vdd.n2193 9.3005
R20862 vdd.n307 vdd.n306 9.3005
R20863 vdd.n302 vdd.n301 9.3005
R20864 vdd.n313 vdd.n312 9.3005
R20865 vdd.n315 vdd.n314 9.3005
R20866 vdd.n298 vdd.n297 9.3005
R20867 vdd.n321 vdd.n320 9.3005
R20868 vdd.n323 vdd.n322 9.3005
R20869 vdd.n295 vdd.n292 9.3005
R20870 vdd.n330 vdd.n329 9.3005
R20871 vdd.n248 vdd.n247 9.3005
R20872 vdd.n243 vdd.n242 9.3005
R20873 vdd.n254 vdd.n253 9.3005
R20874 vdd.n256 vdd.n255 9.3005
R20875 vdd.n239 vdd.n238 9.3005
R20876 vdd.n262 vdd.n261 9.3005
R20877 vdd.n264 vdd.n263 9.3005
R20878 vdd.n236 vdd.n233 9.3005
R20879 vdd.n271 vdd.n270 9.3005
R20880 vdd.n205 vdd.n204 9.3005
R20881 vdd.n200 vdd.n199 9.3005
R20882 vdd.n211 vdd.n210 9.3005
R20883 vdd.n213 vdd.n212 9.3005
R20884 vdd.n196 vdd.n195 9.3005
R20885 vdd.n219 vdd.n218 9.3005
R20886 vdd.n221 vdd.n220 9.3005
R20887 vdd.n193 vdd.n190 9.3005
R20888 vdd.n228 vdd.n227 9.3005
R20889 vdd.n146 vdd.n145 9.3005
R20890 vdd.n141 vdd.n140 9.3005
R20891 vdd.n152 vdd.n151 9.3005
R20892 vdd.n154 vdd.n153 9.3005
R20893 vdd.n137 vdd.n136 9.3005
R20894 vdd.n160 vdd.n159 9.3005
R20895 vdd.n162 vdd.n161 9.3005
R20896 vdd.n134 vdd.n131 9.3005
R20897 vdd.n169 vdd.n168 9.3005
R20898 vdd.n104 vdd.n103 9.3005
R20899 vdd.n99 vdd.n98 9.3005
R20900 vdd.n110 vdd.n109 9.3005
R20901 vdd.n112 vdd.n111 9.3005
R20902 vdd.n95 vdd.n94 9.3005
R20903 vdd.n118 vdd.n117 9.3005
R20904 vdd.n120 vdd.n119 9.3005
R20905 vdd.n92 vdd.n89 9.3005
R20906 vdd.n127 vdd.n126 9.3005
R20907 vdd.n45 vdd.n44 9.3005
R20908 vdd.n40 vdd.n39 9.3005
R20909 vdd.n51 vdd.n50 9.3005
R20910 vdd.n53 vdd.n52 9.3005
R20911 vdd.n36 vdd.n35 9.3005
R20912 vdd.n59 vdd.n58 9.3005
R20913 vdd.n61 vdd.n60 9.3005
R20914 vdd.n33 vdd.n30 9.3005
R20915 vdd.n68 vdd.n67 9.3005
R20916 vdd.n3320 vdd.n3319 9.3005
R20917 vdd.n3323 vdd.n766 9.3005
R20918 vdd.n3324 vdd.n765 9.3005
R20919 vdd.n3327 vdd.n764 9.3005
R20920 vdd.n3328 vdd.n763 9.3005
R20921 vdd.n3331 vdd.n762 9.3005
R20922 vdd.n3332 vdd.n761 9.3005
R20923 vdd.n3335 vdd.n760 9.3005
R20924 vdd.n3336 vdd.n759 9.3005
R20925 vdd.n3339 vdd.n758 9.3005
R20926 vdd.n3340 vdd.n757 9.3005
R20927 vdd.n3343 vdd.n756 9.3005
R20928 vdd.n3344 vdd.n755 9.3005
R20929 vdd.n3347 vdd.n754 9.3005
R20930 vdd.n3348 vdd.n753 9.3005
R20931 vdd.n3351 vdd.n752 9.3005
R20932 vdd.n3352 vdd.n751 9.3005
R20933 vdd.n3355 vdd.n750 9.3005
R20934 vdd.n3356 vdd.n749 9.3005
R20935 vdd.n3359 vdd.n748 9.3005
R20936 vdd.n3363 vdd.n3362 9.3005
R20937 vdd.n3364 vdd.n747 9.3005
R20938 vdd.n3368 vdd.n3365 9.3005
R20939 vdd.n3371 vdd.n746 9.3005
R20940 vdd.n3372 vdd.n745 9.3005
R20941 vdd.n3375 vdd.n744 9.3005
R20942 vdd.n3376 vdd.n743 9.3005
R20943 vdd.n3379 vdd.n742 9.3005
R20944 vdd.n3380 vdd.n741 9.3005
R20945 vdd.n3383 vdd.n740 9.3005
R20946 vdd.n3384 vdd.n739 9.3005
R20947 vdd.n3387 vdd.n738 9.3005
R20948 vdd.n3388 vdd.n737 9.3005
R20949 vdd.n3391 vdd.n736 9.3005
R20950 vdd.n3392 vdd.n735 9.3005
R20951 vdd.n3395 vdd.n730 9.3005
R20952 vdd.n3401 vdd.n727 9.3005
R20953 vdd.n3402 vdd.n726 9.3005
R20954 vdd.n3416 vdd.n3415 9.3005
R20955 vdd.n3417 vdd.n681 9.3005
R20956 vdd.n3419 vdd.n3418 9.3005
R20957 vdd.n671 vdd.n670 9.3005
R20958 vdd.n3433 vdd.n3432 9.3005
R20959 vdd.n3434 vdd.n669 9.3005
R20960 vdd.n3436 vdd.n3435 9.3005
R20961 vdd.n660 vdd.n659 9.3005
R20962 vdd.n3449 vdd.n3448 9.3005
R20963 vdd.n3450 vdd.n658 9.3005
R20964 vdd.n3452 vdd.n3451 9.3005
R20965 vdd.n648 vdd.n647 9.3005
R20966 vdd.n3466 vdd.n3465 9.3005
R20967 vdd.n3467 vdd.n646 9.3005
R20968 vdd.n3469 vdd.n3468 9.3005
R20969 vdd.n637 vdd.n636 9.3005
R20970 vdd.n3485 vdd.n3484 9.3005
R20971 vdd.n3486 vdd.n635 9.3005
R20972 vdd.n3488 vdd.n3487 9.3005
R20973 vdd.n336 vdd.n334 9.3005
R20974 vdd.n683 vdd.n682 9.3005
R20975 vdd.n3580 vdd.n3579 9.3005
R20976 vdd.n337 vdd.n335 9.3005
R20977 vdd.n3573 vdd.n346 9.3005
R20978 vdd.n3572 vdd.n347 9.3005
R20979 vdd.n3571 vdd.n348 9.3005
R20980 vdd.n355 vdd.n349 9.3005
R20981 vdd.n3565 vdd.n356 9.3005
R20982 vdd.n3564 vdd.n357 9.3005
R20983 vdd.n3563 vdd.n358 9.3005
R20984 vdd.n366 vdd.n359 9.3005
R20985 vdd.n3557 vdd.n367 9.3005
R20986 vdd.n3556 vdd.n368 9.3005
R20987 vdd.n3555 vdd.n369 9.3005
R20988 vdd.n377 vdd.n370 9.3005
R20989 vdd.n3549 vdd.n378 9.3005
R20990 vdd.n3548 vdd.n379 9.3005
R20991 vdd.n3547 vdd.n380 9.3005
R20992 vdd.n388 vdd.n381 9.3005
R20993 vdd.n3541 vdd.n389 9.3005
R20994 vdd.n3540 vdd.n390 9.3005
R20995 vdd.n3539 vdd.n391 9.3005
R20996 vdd.n466 vdd.n463 9.3005
R20997 vdd.n470 vdd.n469 9.3005
R20998 vdd.n471 vdd.n462 9.3005
R20999 vdd.n475 vdd.n472 9.3005
R21000 vdd.n476 vdd.n461 9.3005
R21001 vdd.n480 vdd.n479 9.3005
R21002 vdd.n481 vdd.n460 9.3005
R21003 vdd.n485 vdd.n482 9.3005
R21004 vdd.n486 vdd.n459 9.3005
R21005 vdd.n490 vdd.n489 9.3005
R21006 vdd.n491 vdd.n458 9.3005
R21007 vdd.n495 vdd.n492 9.3005
R21008 vdd.n496 vdd.n457 9.3005
R21009 vdd.n500 vdd.n499 9.3005
R21010 vdd.n501 vdd.n456 9.3005
R21011 vdd.n505 vdd.n502 9.3005
R21012 vdd.n506 vdd.n455 9.3005
R21013 vdd.n510 vdd.n509 9.3005
R21014 vdd.n511 vdd.n454 9.3005
R21015 vdd.n515 vdd.n512 9.3005
R21016 vdd.n516 vdd.n451 9.3005
R21017 vdd.n520 vdd.n519 9.3005
R21018 vdd.n521 vdd.n450 9.3005
R21019 vdd.n525 vdd.n522 9.3005
R21020 vdd.n526 vdd.n449 9.3005
R21021 vdd.n530 vdd.n529 9.3005
R21022 vdd.n531 vdd.n448 9.3005
R21023 vdd.n535 vdd.n532 9.3005
R21024 vdd.n536 vdd.n447 9.3005
R21025 vdd.n540 vdd.n539 9.3005
R21026 vdd.n541 vdd.n446 9.3005
R21027 vdd.n545 vdd.n542 9.3005
R21028 vdd.n546 vdd.n445 9.3005
R21029 vdd.n550 vdd.n549 9.3005
R21030 vdd.n551 vdd.n444 9.3005
R21031 vdd.n555 vdd.n552 9.3005
R21032 vdd.n556 vdd.n443 9.3005
R21033 vdd.n560 vdd.n559 9.3005
R21034 vdd.n561 vdd.n442 9.3005
R21035 vdd.n565 vdd.n562 9.3005
R21036 vdd.n566 vdd.n439 9.3005
R21037 vdd.n570 vdd.n569 9.3005
R21038 vdd.n571 vdd.n438 9.3005
R21039 vdd.n575 vdd.n572 9.3005
R21040 vdd.n576 vdd.n437 9.3005
R21041 vdd.n580 vdd.n579 9.3005
R21042 vdd.n581 vdd.n436 9.3005
R21043 vdd.n585 vdd.n582 9.3005
R21044 vdd.n586 vdd.n435 9.3005
R21045 vdd.n590 vdd.n589 9.3005
R21046 vdd.n591 vdd.n434 9.3005
R21047 vdd.n595 vdd.n592 9.3005
R21048 vdd.n596 vdd.n433 9.3005
R21049 vdd.n600 vdd.n599 9.3005
R21050 vdd.n601 vdd.n432 9.3005
R21051 vdd.n605 vdd.n602 9.3005
R21052 vdd.n606 vdd.n431 9.3005
R21053 vdd.n610 vdd.n609 9.3005
R21054 vdd.n611 vdd.n430 9.3005
R21055 vdd.n615 vdd.n612 9.3005
R21056 vdd.n617 vdd.n429 9.3005
R21057 vdd.n619 vdd.n618 9.3005
R21058 vdd.n3533 vdd.n3532 9.3005
R21059 vdd.n465 vdd.n464 9.3005
R21060 vdd.n3411 vdd.n3410 9.3005
R21061 vdd.n676 vdd.n675 9.3005
R21062 vdd.n3424 vdd.n3423 9.3005
R21063 vdd.n3425 vdd.n674 9.3005
R21064 vdd.n3427 vdd.n3426 9.3005
R21065 vdd.n666 vdd.n665 9.3005
R21066 vdd.n3441 vdd.n3440 9.3005
R21067 vdd.n3442 vdd.n664 9.3005
R21068 vdd.n3444 vdd.n3443 9.3005
R21069 vdd.n653 vdd.n652 9.3005
R21070 vdd.n3457 vdd.n3456 9.3005
R21071 vdd.n3458 vdd.n651 9.3005
R21072 vdd.n3460 vdd.n3459 9.3005
R21073 vdd.n642 vdd.n641 9.3005
R21074 vdd.n3474 vdd.n3473 9.3005
R21075 vdd.n3475 vdd.n640 9.3005
R21076 vdd.n3480 vdd.n3476 9.3005
R21077 vdd.n3479 vdd.n3478 9.3005
R21078 vdd.n3477 vdd.n631 9.3005
R21079 vdd.n3493 vdd.n630 9.3005
R21080 vdd.n3495 vdd.n3494 9.3005
R21081 vdd.n3496 vdd.n629 9.3005
R21082 vdd.n3498 vdd.n3497 9.3005
R21083 vdd.n3500 vdd.n628 9.3005
R21084 vdd.n3502 vdd.n3501 9.3005
R21085 vdd.n3503 vdd.n627 9.3005
R21086 vdd.n3505 vdd.n3504 9.3005
R21087 vdd.n3507 vdd.n626 9.3005
R21088 vdd.n3509 vdd.n3508 9.3005
R21089 vdd.n3510 vdd.n625 9.3005
R21090 vdd.n3512 vdd.n3511 9.3005
R21091 vdd.n3515 vdd.n624 9.3005
R21092 vdd.n3517 vdd.n3516 9.3005
R21093 vdd.n3518 vdd.n623 9.3005
R21094 vdd.n3520 vdd.n3519 9.3005
R21095 vdd.n3522 vdd.n622 9.3005
R21096 vdd.n3524 vdd.n3523 9.3005
R21097 vdd.n3525 vdd.n621 9.3005
R21098 vdd.n3527 vdd.n3526 9.3005
R21099 vdd.n3529 vdd.n620 9.3005
R21100 vdd.n3531 vdd.n3530 9.3005
R21101 vdd.n3409 vdd.n686 9.3005
R21102 vdd.n3408 vdd.n3407 9.3005
R21103 vdd.n3277 vdd.n687 9.3005
R21104 vdd.n3286 vdd.n783 9.3005
R21105 vdd.n3289 vdd.n782 9.3005
R21106 vdd.n3290 vdd.n781 9.3005
R21107 vdd.n3293 vdd.n780 9.3005
R21108 vdd.n3294 vdd.n779 9.3005
R21109 vdd.n3297 vdd.n778 9.3005
R21110 vdd.n3298 vdd.n777 9.3005
R21111 vdd.n3301 vdd.n776 9.3005
R21112 vdd.n3302 vdd.n775 9.3005
R21113 vdd.n3305 vdd.n774 9.3005
R21114 vdd.n3306 vdd.n773 9.3005
R21115 vdd.n3309 vdd.n772 9.3005
R21116 vdd.n3310 vdd.n771 9.3005
R21117 vdd.n3313 vdd.n770 9.3005
R21118 vdd.n3317 vdd.n3316 9.3005
R21119 vdd.n3318 vdd.n767 9.3005
R21120 vdd.n2204 vdd.n2203 9.3005
R21121 vdd.n2199 vdd.n1147 9.3005
R21122 vdd.n1510 vdd.n1509 9.3005
R21123 vdd.n1511 vdd.n1265 9.3005
R21124 vdd.n1513 vdd.n1512 9.3005
R21125 vdd.n1255 vdd.n1254 9.3005
R21126 vdd.n1527 vdd.n1526 9.3005
R21127 vdd.n1528 vdd.n1253 9.3005
R21128 vdd.n1530 vdd.n1529 9.3005
R21129 vdd.n1245 vdd.n1244 9.3005
R21130 vdd.n1544 vdd.n1543 9.3005
R21131 vdd.n1545 vdd.n1243 9.3005
R21132 vdd.n1547 vdd.n1546 9.3005
R21133 vdd.n1232 vdd.n1231 9.3005
R21134 vdd.n1560 vdd.n1559 9.3005
R21135 vdd.n1561 vdd.n1230 9.3005
R21136 vdd.n1563 vdd.n1562 9.3005
R21137 vdd.n1221 vdd.n1220 9.3005
R21138 vdd.n1577 vdd.n1576 9.3005
R21139 vdd.n1578 vdd.n1219 9.3005
R21140 vdd.n1580 vdd.n1579 9.3005
R21141 vdd.n1210 vdd.n1209 9.3005
R21142 vdd.n1900 vdd.n1899 9.3005
R21143 vdd.n1901 vdd.n1208 9.3005
R21144 vdd.n1903 vdd.n1902 9.3005
R21145 vdd.n1198 vdd.n1197 9.3005
R21146 vdd.n1917 vdd.n1916 9.3005
R21147 vdd.n1918 vdd.n1196 9.3005
R21148 vdd.n1920 vdd.n1919 9.3005
R21149 vdd.n1188 vdd.n1187 9.3005
R21150 vdd.n1934 vdd.n1933 9.3005
R21151 vdd.n1935 vdd.n1186 9.3005
R21152 vdd.n1937 vdd.n1936 9.3005
R21153 vdd.n1175 vdd.n1174 9.3005
R21154 vdd.n1950 vdd.n1949 9.3005
R21155 vdd.n1951 vdd.n1173 9.3005
R21156 vdd.n1953 vdd.n1952 9.3005
R21157 vdd.n1165 vdd.n1164 9.3005
R21158 vdd.n1967 vdd.n1966 9.3005
R21159 vdd.n1968 vdd.n1162 9.3005
R21160 vdd.n1972 vdd.n1971 9.3005
R21161 vdd.n1970 vdd.n1163 9.3005
R21162 vdd.n1969 vdd.n1152 9.3005
R21163 vdd.n1267 vdd.n1266 9.3005
R21164 vdd.n1403 vdd.n1402 9.3005
R21165 vdd.n1404 vdd.n1393 9.3005
R21166 vdd.n1406 vdd.n1405 9.3005
R21167 vdd.n1407 vdd.n1392 9.3005
R21168 vdd.n1409 vdd.n1408 9.3005
R21169 vdd.n1410 vdd.n1387 9.3005
R21170 vdd.n1412 vdd.n1411 9.3005
R21171 vdd.n1413 vdd.n1386 9.3005
R21172 vdd.n1415 vdd.n1414 9.3005
R21173 vdd.n1416 vdd.n1381 9.3005
R21174 vdd.n1418 vdd.n1417 9.3005
R21175 vdd.n1419 vdd.n1380 9.3005
R21176 vdd.n1421 vdd.n1420 9.3005
R21177 vdd.n1422 vdd.n1375 9.3005
R21178 vdd.n1424 vdd.n1423 9.3005
R21179 vdd.n1425 vdd.n1374 9.3005
R21180 vdd.n1427 vdd.n1426 9.3005
R21181 vdd.n1428 vdd.n1369 9.3005
R21182 vdd.n1430 vdd.n1429 9.3005
R21183 vdd.n1431 vdd.n1368 9.3005
R21184 vdd.n1433 vdd.n1432 9.3005
R21185 vdd.n1437 vdd.n1364 9.3005
R21186 vdd.n1439 vdd.n1438 9.3005
R21187 vdd.n1440 vdd.n1363 9.3005
R21188 vdd.n1442 vdd.n1441 9.3005
R21189 vdd.n1443 vdd.n1358 9.3005
R21190 vdd.n1445 vdd.n1444 9.3005
R21191 vdd.n1446 vdd.n1357 9.3005
R21192 vdd.n1448 vdd.n1447 9.3005
R21193 vdd.n1449 vdd.n1352 9.3005
R21194 vdd.n1451 vdd.n1450 9.3005
R21195 vdd.n1452 vdd.n1351 9.3005
R21196 vdd.n1454 vdd.n1453 9.3005
R21197 vdd.n1455 vdd.n1346 9.3005
R21198 vdd.n1457 vdd.n1456 9.3005
R21199 vdd.n1458 vdd.n1345 9.3005
R21200 vdd.n1460 vdd.n1459 9.3005
R21201 vdd.n1461 vdd.n1340 9.3005
R21202 vdd.n1463 vdd.n1462 9.3005
R21203 vdd.n1464 vdd.n1339 9.3005
R21204 vdd.n1466 vdd.n1465 9.3005
R21205 vdd.n1467 vdd.n1334 9.3005
R21206 vdd.n1469 vdd.n1468 9.3005
R21207 vdd.n1470 vdd.n1333 9.3005
R21208 vdd.n1472 vdd.n1471 9.3005
R21209 vdd.n1473 vdd.n1326 9.3005
R21210 vdd.n1475 vdd.n1474 9.3005
R21211 vdd.n1476 vdd.n1325 9.3005
R21212 vdd.n1478 vdd.n1477 9.3005
R21213 vdd.n1479 vdd.n1320 9.3005
R21214 vdd.n1481 vdd.n1480 9.3005
R21215 vdd.n1482 vdd.n1319 9.3005
R21216 vdd.n1484 vdd.n1483 9.3005
R21217 vdd.n1485 vdd.n1314 9.3005
R21218 vdd.n1487 vdd.n1486 9.3005
R21219 vdd.n1488 vdd.n1313 9.3005
R21220 vdd.n1490 vdd.n1489 9.3005
R21221 vdd.n1491 vdd.n1308 9.3005
R21222 vdd.n1493 vdd.n1492 9.3005
R21223 vdd.n1494 vdd.n1307 9.3005
R21224 vdd.n1496 vdd.n1495 9.3005
R21225 vdd.n1272 vdd.n1271 9.3005
R21226 vdd.n1502 vdd.n1501 9.3005
R21227 vdd.n1401 vdd.n1400 9.3005
R21228 vdd.n1505 vdd.n1504 9.3005
R21229 vdd.n1261 vdd.n1260 9.3005
R21230 vdd.n1519 vdd.n1518 9.3005
R21231 vdd.n1520 vdd.n1259 9.3005
R21232 vdd.n1522 vdd.n1521 9.3005
R21233 vdd.n1250 vdd.n1249 9.3005
R21234 vdd.n1536 vdd.n1535 9.3005
R21235 vdd.n1537 vdd.n1248 9.3005
R21236 vdd.n1539 vdd.n1538 9.3005
R21237 vdd.n1239 vdd.n1238 9.3005
R21238 vdd.n1552 vdd.n1551 9.3005
R21239 vdd.n1553 vdd.n1237 9.3005
R21240 vdd.n1555 vdd.n1554 9.3005
R21241 vdd.n1227 vdd.n1226 9.3005
R21242 vdd.n1569 vdd.n1568 9.3005
R21243 vdd.n1570 vdd.n1225 9.3005
R21244 vdd.n1572 vdd.n1571 9.3005
R21245 vdd.n1216 vdd.n1215 9.3005
R21246 vdd.n1585 vdd.n1584 9.3005
R21247 vdd.n1586 vdd.n1214 9.3005
R21248 vdd.n1503 vdd.n1270 9.3005
R21249 vdd.n1806 vdd.n1805 9.3005
R21250 vdd.n1801 vdd.n1800 9.3005
R21251 vdd.n1812 vdd.n1811 9.3005
R21252 vdd.n1814 vdd.n1813 9.3005
R21253 vdd.n1797 vdd.n1796 9.3005
R21254 vdd.n1820 vdd.n1819 9.3005
R21255 vdd.n1822 vdd.n1821 9.3005
R21256 vdd.n1794 vdd.n1791 9.3005
R21257 vdd.n1829 vdd.n1828 9.3005
R21258 vdd.n1865 vdd.n1864 9.3005
R21259 vdd.n1860 vdd.n1859 9.3005
R21260 vdd.n1871 vdd.n1870 9.3005
R21261 vdd.n1873 vdd.n1872 9.3005
R21262 vdd.n1856 vdd.n1855 9.3005
R21263 vdd.n1879 vdd.n1878 9.3005
R21264 vdd.n1881 vdd.n1880 9.3005
R21265 vdd.n1853 vdd.n1850 9.3005
R21266 vdd.n1888 vdd.n1887 9.3005
R21267 vdd.n1704 vdd.n1703 9.3005
R21268 vdd.n1699 vdd.n1698 9.3005
R21269 vdd.n1710 vdd.n1709 9.3005
R21270 vdd.n1712 vdd.n1711 9.3005
R21271 vdd.n1695 vdd.n1694 9.3005
R21272 vdd.n1718 vdd.n1717 9.3005
R21273 vdd.n1720 vdd.n1719 9.3005
R21274 vdd.n1692 vdd.n1689 9.3005
R21275 vdd.n1727 vdd.n1726 9.3005
R21276 vdd.n1763 vdd.n1762 9.3005
R21277 vdd.n1758 vdd.n1757 9.3005
R21278 vdd.n1769 vdd.n1768 9.3005
R21279 vdd.n1771 vdd.n1770 9.3005
R21280 vdd.n1754 vdd.n1753 9.3005
R21281 vdd.n1777 vdd.n1776 9.3005
R21282 vdd.n1779 vdd.n1778 9.3005
R21283 vdd.n1751 vdd.n1748 9.3005
R21284 vdd.n1786 vdd.n1785 9.3005
R21285 vdd.n1603 vdd.n1602 9.3005
R21286 vdd.n1598 vdd.n1597 9.3005
R21287 vdd.n1609 vdd.n1608 9.3005
R21288 vdd.n1611 vdd.n1610 9.3005
R21289 vdd.n1594 vdd.n1593 9.3005
R21290 vdd.n1617 vdd.n1616 9.3005
R21291 vdd.n1619 vdd.n1618 9.3005
R21292 vdd.n1591 vdd.n1588 9.3005
R21293 vdd.n1626 vdd.n1625 9.3005
R21294 vdd.n1662 vdd.n1661 9.3005
R21295 vdd.n1657 vdd.n1656 9.3005
R21296 vdd.n1668 vdd.n1667 9.3005
R21297 vdd.n1670 vdd.n1669 9.3005
R21298 vdd.n1653 vdd.n1652 9.3005
R21299 vdd.n1676 vdd.n1675 9.3005
R21300 vdd.n1678 vdd.n1677 9.3005
R21301 vdd.n1650 vdd.n1647 9.3005
R21302 vdd.n1685 vdd.n1684 9.3005
R21303 vdd.n1541 vdd.t245 9.18308
R21304 vdd.n3513 vdd.t181 9.18308
R21305 vdd.n1235 vdd.t224 8.95635
R21306 vdd.n2196 vdd.t84 8.95635
R21307 vdd.n723 vdd.t58 8.95635
R21308 vdd.t190 vdd.n3567 8.95635
R21309 vdd.n312 vdd.n311 8.92171
R21310 vdd.n253 vdd.n252 8.92171
R21311 vdd.n210 vdd.n209 8.92171
R21312 vdd.n151 vdd.n150 8.92171
R21313 vdd.n109 vdd.n108 8.92171
R21314 vdd.n50 vdd.n49 8.92171
R21315 vdd.n1811 vdd.n1810 8.92171
R21316 vdd.n1870 vdd.n1869 8.92171
R21317 vdd.n1709 vdd.n1708 8.92171
R21318 vdd.n1768 vdd.n1767 8.92171
R21319 vdd.n1608 vdd.n1607 8.92171
R21320 vdd.n1667 vdd.n1666 8.92171
R21321 vdd.n231 vdd.n129 8.81535
R21322 vdd.n1789 vdd.n1687 8.81535
R21323 vdd.n1582 vdd.t135 8.72962
R21324 vdd.t217 vdd.n3576 8.72962
R21325 vdd.n1905 vdd.t143 8.50289
R21326 vdd.n3482 vdd.t160 8.50289
R21327 vdd.n28 vdd.n14 8.42249
R21328 vdd.n1931 vdd.t173 8.27616
R21329 vdd.t219 vdd.n656 8.27616
R21330 vdd.n3582 vdd.n3581 8.16225
R21331 vdd.n1893 vdd.n1892 8.16225
R21332 vdd.n308 vdd.n302 8.14595
R21333 vdd.n249 vdd.n243 8.14595
R21334 vdd.n206 vdd.n200 8.14595
R21335 vdd.n147 vdd.n141 8.14595
R21336 vdd.n105 vdd.n99 8.14595
R21337 vdd.n46 vdd.n40 8.14595
R21338 vdd.n1807 vdd.n1801 8.14595
R21339 vdd.n1866 vdd.n1860 8.14595
R21340 vdd.n1705 vdd.n1699 8.14595
R21341 vdd.n1764 vdd.n1758 8.14595
R21342 vdd.n1604 vdd.n1598 8.14595
R21343 vdd.n1663 vdd.n1657 8.14595
R21344 vdd.n1178 vdd.t145 8.04943
R21345 vdd.n3438 vdd.t141 8.04943
R21346 vdd.n2467 vdd.n1104 7.70933
R21347 vdd.n2473 vdd.n1104 7.70933
R21348 vdd.n2479 vdd.n1098 7.70933
R21349 vdd.n2479 vdd.n1092 7.70933
R21350 vdd.n2485 vdd.n1092 7.70933
R21351 vdd.n2485 vdd.n1086 7.70933
R21352 vdd.n2491 vdd.n1086 7.70933
R21353 vdd.n2497 vdd.n1080 7.70933
R21354 vdd.n2503 vdd.n1074 7.70933
R21355 vdd.n2509 vdd.n1067 7.70933
R21356 vdd.n2509 vdd.n1070 7.70933
R21357 vdd.n2515 vdd.n1063 7.70933
R21358 vdd.n2522 vdd.n1049 7.70933
R21359 vdd.n2528 vdd.n1049 7.70933
R21360 vdd.n2534 vdd.n1043 7.70933
R21361 vdd.n2540 vdd.n1039 7.70933
R21362 vdd.n2546 vdd.n1033 7.70933
R21363 vdd.n2564 vdd.n1015 7.70933
R21364 vdd.n2564 vdd.n1008 7.70933
R21365 vdd.n2572 vdd.n1008 7.70933
R21366 vdd.n2654 vdd.n992 7.70933
R21367 vdd.n3017 vdd.n946 7.70933
R21368 vdd.n3029 vdd.n927 7.70933
R21369 vdd.n3035 vdd.n927 7.70933
R21370 vdd.n3035 vdd.n930 7.70933
R21371 vdd.n3053 vdd.n911 7.70933
R21372 vdd.n3059 vdd.n905 7.70933
R21373 vdd.n3065 vdd.n901 7.70933
R21374 vdd.n3071 vdd.n888 7.70933
R21375 vdd.n3077 vdd.n888 7.70933
R21376 vdd.n3084 vdd.n881 7.70933
R21377 vdd.n3090 vdd.n874 7.70933
R21378 vdd.n3090 vdd.n877 7.70933
R21379 vdd.n3096 vdd.n870 7.70933
R21380 vdd.n3102 vdd.n864 7.70933
R21381 vdd.n3108 vdd.n851 7.70933
R21382 vdd.n3114 vdd.n851 7.70933
R21383 vdd.n3114 vdd.n843 7.70933
R21384 vdd.n3165 vdd.n843 7.70933
R21385 vdd.n3165 vdd.n846 7.70933
R21386 vdd.n3171 vdd.n805 7.70933
R21387 vdd.n3241 vdd.n805 7.70933
R21388 vdd.t18 vdd.n1080 7.59597
R21389 vdd.n2346 vdd.t293 7.59597
R21390 vdd.n2989 vdd.t11 7.59597
R21391 vdd.n864 vdd.t55 7.59597
R21392 vdd.n307 vdd.n304 7.3702
R21393 vdd.n248 vdd.n245 7.3702
R21394 vdd.n205 vdd.n202 7.3702
R21395 vdd.n146 vdd.n143 7.3702
R21396 vdd.n104 vdd.n101 7.3702
R21397 vdd.n45 vdd.n42 7.3702
R21398 vdd.n1806 vdd.n1803 7.3702
R21399 vdd.n1865 vdd.n1862 7.3702
R21400 vdd.n1704 vdd.n1701 7.3702
R21401 vdd.n1763 vdd.n1760 7.3702
R21402 vdd.n1603 vdd.n1600 7.3702
R21403 vdd.n1662 vdd.n1659 7.3702
R21404 vdd.n1964 vdd.t232 7.1425
R21405 vdd.n679 vdd.t192 7.1425
R21406 vdd.n1438 vdd.n1437 6.98232
R21407 vdd.n2119 vdd.n2118 6.98232
R21408 vdd.n566 vdd.n565 6.98232
R21409 vdd.n3323 vdd.n3320 6.98232
R21410 vdd.t158 vdd.n1177 6.91577
R21411 vdd.n2503 vdd.t17 6.91577
R21412 vdd.n3096 vdd.t56 6.91577
R21413 vdd.n3446 vdd.t155 6.91577
R21414 vdd.n3081 vdd.n3080 6.86879
R21415 vdd.n2519 vdd.n2518 6.86879
R21416 vdd.n2579 vdd.t294 6.80241
R21417 vdd.n3023 vdd.t51 6.80241
R21418 vdd.n1923 vdd.t230 6.68904
R21419 vdd.n3462 vdd.t153 6.68904
R21420 vdd.t170 vdd.n1206 6.46231
R21421 vdd.n3490 vdd.t147 6.46231
R21422 vdd.n3582 vdd.n333 6.38151
R21423 vdd.n1892 vdd.n1891 6.38151
R21424 vdd.n2346 vdd.t12 6.34895
R21425 vdd.n2989 vdd.t0 6.34895
R21426 vdd.n1574 vdd.t198 6.23558
R21427 vdd.t137 vdd.n344 6.23558
R21428 vdd.t186 vdd.n1234 6.00885
R21429 vdd.t45 vdd.n1043 6.00885
R21430 vdd.n901 vdd.t39 6.00885
R21431 vdd.n3561 vdd.t149 6.00885
R21432 vdd.n308 vdd.n307 5.81868
R21433 vdd.n249 vdd.n248 5.81868
R21434 vdd.n206 vdd.n205 5.81868
R21435 vdd.n147 vdd.n146 5.81868
R21436 vdd.n105 vdd.n104 5.81868
R21437 vdd.n46 vdd.n45 5.81868
R21438 vdd.n1807 vdd.n1806 5.81868
R21439 vdd.n1866 vdd.n1865 5.81868
R21440 vdd.n1705 vdd.n1704 5.81868
R21441 vdd.n1764 vdd.n1763 5.81868
R21442 vdd.n1604 vdd.n1603 5.81868
R21443 vdd.n1663 vdd.n1662 5.81868
R21444 vdd.n1533 vdd.t175 5.78212
R21445 vdd.n3552 vdd.t272 5.78212
R21446 vdd.n2662 vdd.n2661 5.77611
R21447 vdd.n2402 vdd.n2401 5.77611
R21448 vdd.n2891 vdd.n2890 5.77611
R21449 vdd.n3182 vdd.n3181 5.77611
R21450 vdd.n3246 vdd.n801 5.77611
R21451 vdd.n2827 vdd.n2763 5.77611
R21452 vdd.n2587 vdd.n999 5.77611
R21453 vdd.n2278 vdd.n2277 5.77611
R21454 vdd.n1400 vdd.n1399 5.62474
R21455 vdd.n2202 vdd.n2199 5.62474
R21456 vdd.n3533 vdd.n428 5.62474
R21457 vdd.n3407 vdd.n690 5.62474
R21458 vdd.n1257 vdd.t175 5.55539
R21459 vdd.t272 vdd.n3551 5.55539
R21460 vdd.n2540 vdd.t2 5.44203
R21461 vdd.n3059 vdd.t302 5.44203
R21462 vdd.n1549 vdd.t186 5.32866
R21463 vdd.t149 vdd.n3560 5.32866
R21464 vdd.n1565 vdd.t198 5.10193
R21465 vdd.n2515 vdd.t4 5.10193
R21466 vdd.n2534 vdd.t16 5.10193
R21467 vdd.n3065 vdd.t5 5.10193
R21468 vdd.n3084 vdd.t7 5.10193
R21469 vdd.n3569 vdd.t137 5.10193
R21470 vdd.n311 vdd.n302 5.04292
R21471 vdd.n252 vdd.n243 5.04292
R21472 vdd.n209 vdd.n200 5.04292
R21473 vdd.n150 vdd.n141 5.04292
R21474 vdd.n108 vdd.n99 5.04292
R21475 vdd.n49 vdd.n40 5.04292
R21476 vdd.n1810 vdd.n1801 5.04292
R21477 vdd.n1869 vdd.n1860 5.04292
R21478 vdd.n1708 vdd.n1699 5.04292
R21479 vdd.n1767 vdd.n1758 5.04292
R21480 vdd.n1607 vdd.n1598 5.04292
R21481 vdd.n1666 vdd.n1657 5.04292
R21482 vdd.n1063 vdd.t118 4.98857
R21483 vdd.t77 vdd.n881 4.98857
R21484 vdd.n1897 vdd.t170 4.8752
R21485 vdd.t66 vdd.n1098 4.8752
R21486 vdd.t8 vdd.t49 4.8752
R21487 vdd.n2334 vdd.t104 4.8752
R21488 vdd.n3001 vdd.t108 4.8752
R21489 vdd.t14 vdd.t19 4.8752
R21490 vdd.n846 vdd.t62 4.8752
R21491 vdd.t147 vdd.n340 4.8752
R21492 vdd.n2663 vdd.n2662 4.83952
R21493 vdd.n2403 vdd.n2402 4.83952
R21494 vdd.n2890 vdd.n2889 4.83952
R21495 vdd.n3183 vdd.n3182 4.83952
R21496 vdd.n801 vdd.n796 4.83952
R21497 vdd.n2824 vdd.n2763 4.83952
R21498 vdd.n2590 vdd.n999 4.83952
R21499 vdd.n2277 vdd.n2276 4.83952
R21500 vdd.n2558 vdd.t37 4.76184
R21501 vdd.n3041 vdd.t47 4.76184
R21502 vdd.n2087 vdd.n1145 4.74817
R21503 vdd.n2082 vdd.n1146 4.74817
R21504 vdd.n1984 vdd.n1981 4.74817
R21505 vdd.n2183 vdd.n1985 4.74817
R21506 vdd.n2185 vdd.n1984 4.74817
R21507 vdd.n2184 vdd.n2183 4.74817
R21508 vdd.n3400 vdd.n3399 4.74817
R21509 vdd.n3397 vdd.n3396 4.74817
R21510 vdd.n3397 vdd.n732 4.74817
R21511 vdd.n3399 vdd.n729 4.74817
R21512 vdd.n3282 vdd.n784 4.74817
R21513 vdd.n3278 vdd.n3276 4.74817
R21514 vdd.n3281 vdd.n3276 4.74817
R21515 vdd.n3285 vdd.n784 4.74817
R21516 vdd.n2083 vdd.n1145 4.74817
R21517 vdd.n1148 vdd.n1146 4.74817
R21518 vdd.n333 vdd.n332 4.7074
R21519 vdd.n231 vdd.n230 4.7074
R21520 vdd.n1891 vdd.n1890 4.7074
R21521 vdd.n1789 vdd.n1788 4.7074
R21522 vdd.n1200 vdd.t230 4.64847
R21523 vdd.n3471 vdd.t153 4.64847
R21524 vdd.n1939 vdd.t158 4.42174
R21525 vdd.t155 vdd.n655 4.42174
R21526 vdd.n2334 vdd.t300 4.30838
R21527 vdd.n3001 vdd.t40 4.30838
R21528 vdd.n312 vdd.n300 4.26717
R21529 vdd.n253 vdd.n241 4.26717
R21530 vdd.n210 vdd.n198 4.26717
R21531 vdd.n151 vdd.n139 4.26717
R21532 vdd.n109 vdd.n97 4.26717
R21533 vdd.n50 vdd.n38 4.26717
R21534 vdd.n1811 vdd.n1799 4.26717
R21535 vdd.n1870 vdd.n1858 4.26717
R21536 vdd.n1709 vdd.n1697 4.26717
R21537 vdd.n1768 vdd.n1756 4.26717
R21538 vdd.n1608 vdd.n1596 4.26717
R21539 vdd.n1667 vdd.n1655 4.26717
R21540 vdd.n1955 vdd.t232 4.19501
R21541 vdd.t10 vdd.n1074 4.19501
R21542 vdd.n1033 vdd.t42 4.19501
R21543 vdd.t9 vdd.n911 4.19501
R21544 vdd.n870 vdd.t6 4.19501
R21545 vdd.n3430 vdd.t192 4.19501
R21546 vdd.n333 vdd.n231 4.10845
R21547 vdd.n1891 vdd.n1789 4.10845
R21548 vdd.n289 vdd.t243 4.06363
R21549 vdd.n289 vdd.t284 4.06363
R21550 vdd.n287 vdd.t150 4.06363
R21551 vdd.n287 vdd.t207 4.06363
R21552 vdd.n285 vdd.t210 4.06363
R21553 vdd.n285 vdd.t263 4.06363
R21554 vdd.n283 vdd.t265 4.06363
R21555 vdd.n283 vdd.t138 4.06363
R21556 vdd.n281 vdd.t167 4.06363
R21557 vdd.n281 vdd.t237 4.06363
R21558 vdd.n279 vdd.t266 4.06363
R21559 vdd.n279 vdd.t281 4.06363
R21560 vdd.n277 vdd.t285 4.06363
R21561 vdd.n277 vdd.t177 4.06363
R21562 vdd.n275 vdd.t208 4.06363
R21563 vdd.n275 vdd.t283 4.06363
R21564 vdd.n273 vdd.t289 4.06363
R21565 vdd.n273 vdd.t206 4.06363
R21566 vdd.n187 vdd.t235 4.06363
R21567 vdd.n187 vdd.t273 4.06363
R21568 vdd.n185 vdd.t290 4.06363
R21569 vdd.n185 vdd.t182 4.06363
R21570 vdd.n183 vdd.t191 4.06363
R21571 vdd.n183 vdd.t253 4.06363
R21572 vdd.n181 vdd.t254 4.06363
R21573 vdd.n181 vdd.t282 4.06363
R21574 vdd.n179 vdd.t148 4.06363
R21575 vdd.n179 vdd.t218 4.06363
R21576 vdd.n177 vdd.t257 4.06363
R21577 vdd.n177 vdd.t267 4.06363
R21578 vdd.n175 vdd.t275 4.06363
R21579 vdd.n175 vdd.t154 4.06363
R21580 vdd.n173 vdd.t183 4.06363
R21581 vdd.n173 vdd.t274 4.06363
R21582 vdd.n171 vdd.t277 4.06363
R21583 vdd.n171 vdd.t180 4.06363
R21584 vdd.n86 vdd.t212 4.06363
R21585 vdd.n86 vdd.t286 4.06363
R21586 vdd.n84 vdd.t188 4.06363
R21587 vdd.n84 vdd.t270 4.06363
R21588 vdd.n82 vdd.t223 4.06363
R21589 vdd.n82 vdd.t255 4.06363
R21590 vdd.n80 vdd.t203 4.06363
R21591 vdd.n80 vdd.t278 4.06363
R21592 vdd.n78 vdd.t166 4.06363
R21593 vdd.n78 vdd.t264 4.06363
R21594 vdd.n76 vdd.t161 4.06363
R21595 vdd.n76 vdd.t249 4.06363
R21596 vdd.n74 vdd.t185 4.06363
R21597 vdd.n74 vdd.t268 4.06363
R21598 vdd.n72 vdd.t156 4.06363
R21599 vdd.n72 vdd.t220 4.06363
R21600 vdd.n70 vdd.t142 4.06363
R21601 vdd.n70 vdd.t194 4.06363
R21602 vdd.n1831 vdd.t258 4.06363
R21603 vdd.n1831 vdd.t205 4.06363
R21604 vdd.n1833 vdd.t200 4.06363
R21605 vdd.n1833 vdd.t260 4.06363
R21606 vdd.n1835 vdd.t242 4.06363
R21607 vdd.n1835 vdd.t240 4.06363
R21608 vdd.n1837 vdd.t195 4.06363
R21609 vdd.n1837 vdd.t165 4.06363
R21610 vdd.n1839 vdd.t163 4.06363
R21611 vdd.n1839 vdd.t239 4.06363
R21612 vdd.n1841 vdd.t216 4.06363
R21613 vdd.n1841 vdd.t164 4.06363
R21614 vdd.n1843 vdd.t157 4.06363
R21615 vdd.n1843 vdd.t261 4.06363
R21616 vdd.n1845 vdd.t259 4.06363
R21617 vdd.n1845 vdd.t209 4.06363
R21618 vdd.n1847 vdd.t201 4.06363
R21619 vdd.n1847 vdd.t288 4.06363
R21620 vdd.n1729 vdd.t244 4.06363
R21621 vdd.n1729 vdd.t178 4.06363
R21622 vdd.n1731 vdd.t174 4.06363
R21623 vdd.n1731 vdd.t247 4.06363
R21624 vdd.n1733 vdd.t231 4.06363
R21625 vdd.n1733 vdd.t227 4.06363
R21626 vdd.n1735 vdd.t169 4.06363
R21627 vdd.n1735 vdd.t144 4.06363
R21628 vdd.n1737 vdd.t136 4.06363
R21629 vdd.n1737 vdd.t222 4.06363
R21630 vdd.n1739 vdd.t199 4.06363
R21631 vdd.n1739 vdd.t140 4.06363
R21632 vdd.n1741 vdd.t134 4.06363
R21633 vdd.n1741 vdd.t251 4.06363
R21634 vdd.n1743 vdd.t246 4.06363
R21635 vdd.n1743 vdd.t189 4.06363
R21636 vdd.n1745 vdd.t176 4.06363
R21637 vdd.n1745 vdd.t276 4.06363
R21638 vdd.n1628 vdd.t197 4.06363
R21639 vdd.n1628 vdd.t146 4.06363
R21640 vdd.n1630 vdd.t221 4.06363
R21641 vdd.n1630 vdd.t159 4.06363
R21642 vdd.n1632 vdd.t269 4.06363
R21643 vdd.n1632 vdd.t291 4.06363
R21644 vdd.n1634 vdd.t250 4.06363
R21645 vdd.n1634 vdd.t162 4.06363
R21646 vdd.n1636 vdd.t234 4.06363
R21647 vdd.n1636 vdd.t171 4.06363
R21648 vdd.n1638 vdd.t279 4.06363
R21649 vdd.n1638 vdd.t204 4.06363
R21650 vdd.n1640 vdd.t256 4.06363
R21651 vdd.n1640 vdd.t225 4.06363
R21652 vdd.n1642 vdd.t271 4.06363
R21653 vdd.n1642 vdd.t187 4.06363
R21654 vdd.n1644 vdd.t287 4.06363
R21655 vdd.n1644 vdd.t215 4.06363
R21656 vdd.n26 vdd.t34 3.9605
R21657 vdd.n26 vdd.t30 3.9605
R21658 vdd.n23 vdd.t36 3.9605
R21659 vdd.n23 vdd.t33 3.9605
R21660 vdd.n21 vdd.t27 3.9605
R21661 vdd.n21 vdd.t31 3.9605
R21662 vdd.n20 vdd.t22 3.9605
R21663 vdd.n20 vdd.t23 3.9605
R21664 vdd.n15 vdd.t21 3.9605
R21665 vdd.n15 vdd.t24 3.9605
R21666 vdd.n16 vdd.t25 3.9605
R21667 vdd.n16 vdd.t32 3.9605
R21668 vdd.n18 vdd.t28 3.9605
R21669 vdd.n18 vdd.t35 3.9605
R21670 vdd.n25 vdd.t29 3.9605
R21671 vdd.n25 vdd.t26 3.9605
R21672 vdd.n3080 vdd.n3079 3.74684
R21673 vdd.n2520 vdd.n2519 3.74684
R21674 vdd.n7 vdd.t15 3.61217
R21675 vdd.n7 vdd.t303 3.61217
R21676 vdd.n8 vdd.t48 3.61217
R21677 vdd.n8 vdd.t1 3.61217
R21678 vdd.n10 vdd.t52 3.61217
R21679 vdd.n10 vdd.t41 3.61217
R21680 vdd.n12 vdd.t299 3.61217
R21681 vdd.n12 vdd.t54 3.61217
R21682 vdd.n5 vdd.t297 3.61217
R21683 vdd.n5 vdd.t44 3.61217
R21684 vdd.n3 vdd.t301 3.61217
R21685 vdd.n3 vdd.t295 3.61217
R21686 vdd.n1 vdd.t13 3.61217
R21687 vdd.n1 vdd.t38 3.61217
R21688 vdd.n0 vdd.t3 3.61217
R21689 vdd.n0 vdd.t50 3.61217
R21690 vdd.n2497 vdd.t10 3.51482
R21691 vdd.n2552 vdd.t42 3.51482
R21692 vdd.n3047 vdd.t9 3.51482
R21693 vdd.n3102 vdd.t6 3.51482
R21694 vdd.n316 vdd.n315 3.49141
R21695 vdd.n257 vdd.n256 3.49141
R21696 vdd.n214 vdd.n213 3.49141
R21697 vdd.n155 vdd.n154 3.49141
R21698 vdd.n113 vdd.n112 3.49141
R21699 vdd.n54 vdd.n53 3.49141
R21700 vdd.n1815 vdd.n1814 3.49141
R21701 vdd.n1874 vdd.n1873 3.49141
R21702 vdd.n1713 vdd.n1712 3.49141
R21703 vdd.n1772 vdd.n1771 3.49141
R21704 vdd.n1612 vdd.n1611 3.49141
R21705 vdd.n1671 vdd.n1670 3.49141
R21706 vdd.n2572 vdd.t300 3.40145
R21707 vdd.n2726 vdd.t296 3.40145
R21708 vdd.n3010 vdd.t53 3.40145
R21709 vdd.n3029 vdd.t40 3.40145
R21710 vdd.n1956 vdd.t145 3.28809
R21711 vdd.n3429 vdd.t141 3.28809
R21712 vdd.t173 vdd.n1184 3.06136
R21713 vdd.n3454 vdd.t219 3.06136
R21714 vdd.t37 vdd.n1015 2.94799
R21715 vdd.n930 vdd.t47 2.94799
R21716 vdd.n1914 vdd.t143 2.83463
R21717 vdd.n2473 vdd.t66 2.83463
R21718 vdd.n2579 vdd.t104 2.83463
R21719 vdd.n3023 vdd.t108 2.83463
R21720 vdd.n3171 vdd.t62 2.83463
R21721 vdd.n644 vdd.t160 2.83463
R21722 vdd.n319 vdd.n298 2.71565
R21723 vdd.n260 vdd.n239 2.71565
R21724 vdd.n217 vdd.n196 2.71565
R21725 vdd.n158 vdd.n137 2.71565
R21726 vdd.n116 vdd.n95 2.71565
R21727 vdd.n57 vdd.n36 2.71565
R21728 vdd.n1818 vdd.n1797 2.71565
R21729 vdd.n1877 vdd.n1856 2.71565
R21730 vdd.n1716 vdd.n1695 2.71565
R21731 vdd.n1775 vdd.n1754 2.71565
R21732 vdd.n1615 vdd.n1594 2.71565
R21733 vdd.n1674 vdd.n1653 2.71565
R21734 vdd.t135 vdd.n1212 2.6079
R21735 vdd.n1070 vdd.t4 2.6079
R21736 vdd.n2358 vdd.t16 2.6079
R21737 vdd.n2977 vdd.t5 2.6079
R21738 vdd.t7 vdd.n874 2.6079
R21739 vdd.n3577 vdd.t217 2.6079
R21740 vdd.n306 vdd.n305 2.4129
R21741 vdd.n247 vdd.n246 2.4129
R21742 vdd.n204 vdd.n203 2.4129
R21743 vdd.n145 vdd.n144 2.4129
R21744 vdd.n103 vdd.n102 2.4129
R21745 vdd.n44 vdd.n43 2.4129
R21746 vdd.n1805 vdd.n1804 2.4129
R21747 vdd.n1864 vdd.n1863 2.4129
R21748 vdd.n1703 vdd.n1702 2.4129
R21749 vdd.n1762 vdd.n1761 2.4129
R21750 vdd.n1602 vdd.n1601 2.4129
R21751 vdd.n1661 vdd.n1660 2.4129
R21752 vdd.n1566 vdd.t224 2.38117
R21753 vdd.n1974 vdd.t84 2.38117
R21754 vdd.n3413 vdd.t58 2.38117
R21755 vdd.n3568 vdd.t190 2.38117
R21756 vdd.n2182 vdd.n1984 2.27742
R21757 vdd.n2183 vdd.n2182 2.27742
R21758 vdd.n3398 vdd.n3397 2.27742
R21759 vdd.n3399 vdd.n3398 2.27742
R21760 vdd.n3276 vdd.n3275 2.27742
R21761 vdd.n3275 vdd.n784 2.27742
R21762 vdd.n2205 vdd.n1145 2.27742
R21763 vdd.n2205 vdd.n1146 2.27742
R21764 vdd.n2358 vdd.t2 2.2678
R21765 vdd.n2977 vdd.t302 2.2678
R21766 vdd.t245 vdd.n1241 2.15444
R21767 vdd.n3559 vdd.t181 2.15444
R21768 vdd.n2546 vdd.t49 2.04107
R21769 vdd.n3053 vdd.t14 2.04107
R21770 vdd.n320 vdd.n296 1.93989
R21771 vdd.n261 vdd.n237 1.93989
R21772 vdd.n218 vdd.n194 1.93989
R21773 vdd.n159 vdd.n135 1.93989
R21774 vdd.n117 vdd.n93 1.93989
R21775 vdd.n58 vdd.n34 1.93989
R21776 vdd.n1819 vdd.n1795 1.93989
R21777 vdd.n1878 vdd.n1854 1.93989
R21778 vdd.n1717 vdd.n1693 1.93989
R21779 vdd.n1776 vdd.n1752 1.93989
R21780 vdd.n1616 vdd.n1592 1.93989
R21781 vdd.n1675 vdd.n1651 1.93989
R21782 vdd.n1524 vdd.t228 1.92771
R21783 vdd.t151 vdd.n375 1.92771
R21784 vdd.n1532 vdd.t214 1.70098
R21785 vdd.n2522 vdd.t46 1.70098
R21786 vdd.n2528 vdd.t45 1.70098
R21787 vdd.n3071 vdd.t39 1.70098
R21788 vdd.n3077 vdd.t20 1.70098
R21789 vdd.n3553 vdd.t211 1.70098
R21790 vdd.n1557 vdd.t133 1.47425
R21791 vdd.n361 vdd.t252 1.47425
R21792 vdd.n2552 vdd.t12 1.36088
R21793 vdd.n3047 vdd.t0 1.36088
R21794 vdd.n1223 vdd.t139 1.24752
R21795 vdd.t202 vdd.n3575 1.24752
R21796 vdd.n331 vdd.n291 1.16414
R21797 vdd.n324 vdd.n323 1.16414
R21798 vdd.n272 vdd.n232 1.16414
R21799 vdd.n265 vdd.n264 1.16414
R21800 vdd.n229 vdd.n189 1.16414
R21801 vdd.n222 vdd.n221 1.16414
R21802 vdd.n170 vdd.n130 1.16414
R21803 vdd.n163 vdd.n162 1.16414
R21804 vdd.n128 vdd.n88 1.16414
R21805 vdd.n121 vdd.n120 1.16414
R21806 vdd.n69 vdd.n29 1.16414
R21807 vdd.n62 vdd.n61 1.16414
R21808 vdd.n1830 vdd.n1790 1.16414
R21809 vdd.n1823 vdd.n1822 1.16414
R21810 vdd.n1889 vdd.n1849 1.16414
R21811 vdd.n1882 vdd.n1881 1.16414
R21812 vdd.n1728 vdd.n1688 1.16414
R21813 vdd.n1721 vdd.n1720 1.16414
R21814 vdd.n1787 vdd.n1747 1.16414
R21815 vdd.n1780 vdd.n1779 1.16414
R21816 vdd.n1627 vdd.n1587 1.16414
R21817 vdd.n1620 vdd.n1619 1.16414
R21818 vdd.n1686 vdd.n1646 1.16414
R21819 vdd.n1679 vdd.n1678 1.16414
R21820 vdd.n1892 vdd.n28 1.11236
R21821 vdd vdd.n3582 1.10453
R21822 vdd.n1906 vdd.t168 1.02079
R21823 vdd.t118 vdd.t46 1.02079
R21824 vdd.t20 vdd.t77 1.02079
R21825 vdd.t248 vdd.n633 1.02079
R21826 vdd.n1403 vdd.n1399 0.970197
R21827 vdd.n2203 vdd.n2202 0.970197
R21828 vdd.n618 vdd.n428 0.970197
R21829 vdd.n3277 vdd.n690 0.970197
R21830 vdd.t294 vdd.n992 0.907421
R21831 vdd.n946 vdd.t51 0.907421
R21832 vdd.n1922 vdd.t226 0.794056
R21833 vdd.t17 vdd.n1067 0.794056
R21834 vdd.n1039 vdd.t8 0.794056
R21835 vdd.t19 vdd.n905 0.794056
R21836 vdd.n877 vdd.t56 0.794056
R21837 vdd.n3463 vdd.t184 0.794056
R21838 vdd.n1947 vdd.t196 0.567326
R21839 vdd.t179 vdd.n662 0.567326
R21840 vdd.n2193 vdd.n2192 0.530988
R21841 vdd.n726 vdd.n682 0.530988
R21842 vdd.n464 vdd.n391 0.530988
R21843 vdd.n3532 vdd.n3531 0.530988
R21844 vdd.n3409 vdd.n3408 0.530988
R21845 vdd.n1969 vdd.n1147 0.530988
R21846 vdd.n1401 vdd.n1266 0.530988
R21847 vdd.n1503 vdd.n1502 0.530988
R21848 vdd.n4 vdd.n2 0.459552
R21849 vdd.n11 vdd.n9 0.459552
R21850 vdd.n329 vdd.n328 0.388379
R21851 vdd.n295 vdd.n293 0.388379
R21852 vdd.n270 vdd.n269 0.388379
R21853 vdd.n236 vdd.n234 0.388379
R21854 vdd.n227 vdd.n226 0.388379
R21855 vdd.n193 vdd.n191 0.388379
R21856 vdd.n168 vdd.n167 0.388379
R21857 vdd.n134 vdd.n132 0.388379
R21858 vdd.n126 vdd.n125 0.388379
R21859 vdd.n92 vdd.n90 0.388379
R21860 vdd.n67 vdd.n66 0.388379
R21861 vdd.n33 vdd.n31 0.388379
R21862 vdd.n1828 vdd.n1827 0.388379
R21863 vdd.n1794 vdd.n1792 0.388379
R21864 vdd.n1887 vdd.n1886 0.388379
R21865 vdd.n1853 vdd.n1851 0.388379
R21866 vdd.n1726 vdd.n1725 0.388379
R21867 vdd.n1692 vdd.n1690 0.388379
R21868 vdd.n1785 vdd.n1784 0.388379
R21869 vdd.n1751 vdd.n1749 0.388379
R21870 vdd.n1625 vdd.n1624 0.388379
R21871 vdd.n1591 vdd.n1589 0.388379
R21872 vdd.n1684 vdd.n1683 0.388379
R21873 vdd.n1650 vdd.n1648 0.388379
R21874 vdd.n19 vdd.n17 0.387128
R21875 vdd.n24 vdd.n22 0.387128
R21876 vdd.n6 vdd.n4 0.358259
R21877 vdd.n13 vdd.n11 0.358259
R21878 vdd.n276 vdd.n274 0.358259
R21879 vdd.n278 vdd.n276 0.358259
R21880 vdd.n280 vdd.n278 0.358259
R21881 vdd.n282 vdd.n280 0.358259
R21882 vdd.n284 vdd.n282 0.358259
R21883 vdd.n286 vdd.n284 0.358259
R21884 vdd.n288 vdd.n286 0.358259
R21885 vdd.n290 vdd.n288 0.358259
R21886 vdd.n332 vdd.n290 0.358259
R21887 vdd.n174 vdd.n172 0.358259
R21888 vdd.n176 vdd.n174 0.358259
R21889 vdd.n178 vdd.n176 0.358259
R21890 vdd.n180 vdd.n178 0.358259
R21891 vdd.n182 vdd.n180 0.358259
R21892 vdd.n184 vdd.n182 0.358259
R21893 vdd.n186 vdd.n184 0.358259
R21894 vdd.n188 vdd.n186 0.358259
R21895 vdd.n230 vdd.n188 0.358259
R21896 vdd.n73 vdd.n71 0.358259
R21897 vdd.n75 vdd.n73 0.358259
R21898 vdd.n77 vdd.n75 0.358259
R21899 vdd.n79 vdd.n77 0.358259
R21900 vdd.n81 vdd.n79 0.358259
R21901 vdd.n83 vdd.n81 0.358259
R21902 vdd.n85 vdd.n83 0.358259
R21903 vdd.n87 vdd.n85 0.358259
R21904 vdd.n129 vdd.n87 0.358259
R21905 vdd.n1890 vdd.n1848 0.358259
R21906 vdd.n1848 vdd.n1846 0.358259
R21907 vdd.n1846 vdd.n1844 0.358259
R21908 vdd.n1844 vdd.n1842 0.358259
R21909 vdd.n1842 vdd.n1840 0.358259
R21910 vdd.n1840 vdd.n1838 0.358259
R21911 vdd.n1838 vdd.n1836 0.358259
R21912 vdd.n1836 vdd.n1834 0.358259
R21913 vdd.n1834 vdd.n1832 0.358259
R21914 vdd.n1788 vdd.n1746 0.358259
R21915 vdd.n1746 vdd.n1744 0.358259
R21916 vdd.n1744 vdd.n1742 0.358259
R21917 vdd.n1742 vdd.n1740 0.358259
R21918 vdd.n1740 vdd.n1738 0.358259
R21919 vdd.n1738 vdd.n1736 0.358259
R21920 vdd.n1736 vdd.n1734 0.358259
R21921 vdd.n1734 vdd.n1732 0.358259
R21922 vdd.n1732 vdd.n1730 0.358259
R21923 vdd.n1687 vdd.n1645 0.358259
R21924 vdd.n1645 vdd.n1643 0.358259
R21925 vdd.n1643 vdd.n1641 0.358259
R21926 vdd.n1641 vdd.n1639 0.358259
R21927 vdd.n1639 vdd.n1637 0.358259
R21928 vdd.n1637 vdd.n1635 0.358259
R21929 vdd.n1635 vdd.n1633 0.358259
R21930 vdd.n1633 vdd.n1631 0.358259
R21931 vdd.n1631 vdd.n1629 0.358259
R21932 vdd.n14 vdd.n6 0.334552
R21933 vdd.n14 vdd.n13 0.334552
R21934 vdd.n27 vdd.n19 0.21707
R21935 vdd.n27 vdd.n24 0.21707
R21936 vdd.n330 vdd.n292 0.155672
R21937 vdd.n322 vdd.n292 0.155672
R21938 vdd.n322 vdd.n321 0.155672
R21939 vdd.n321 vdd.n297 0.155672
R21940 vdd.n314 vdd.n297 0.155672
R21941 vdd.n314 vdd.n313 0.155672
R21942 vdd.n313 vdd.n301 0.155672
R21943 vdd.n306 vdd.n301 0.155672
R21944 vdd.n271 vdd.n233 0.155672
R21945 vdd.n263 vdd.n233 0.155672
R21946 vdd.n263 vdd.n262 0.155672
R21947 vdd.n262 vdd.n238 0.155672
R21948 vdd.n255 vdd.n238 0.155672
R21949 vdd.n255 vdd.n254 0.155672
R21950 vdd.n254 vdd.n242 0.155672
R21951 vdd.n247 vdd.n242 0.155672
R21952 vdd.n228 vdd.n190 0.155672
R21953 vdd.n220 vdd.n190 0.155672
R21954 vdd.n220 vdd.n219 0.155672
R21955 vdd.n219 vdd.n195 0.155672
R21956 vdd.n212 vdd.n195 0.155672
R21957 vdd.n212 vdd.n211 0.155672
R21958 vdd.n211 vdd.n199 0.155672
R21959 vdd.n204 vdd.n199 0.155672
R21960 vdd.n169 vdd.n131 0.155672
R21961 vdd.n161 vdd.n131 0.155672
R21962 vdd.n161 vdd.n160 0.155672
R21963 vdd.n160 vdd.n136 0.155672
R21964 vdd.n153 vdd.n136 0.155672
R21965 vdd.n153 vdd.n152 0.155672
R21966 vdd.n152 vdd.n140 0.155672
R21967 vdd.n145 vdd.n140 0.155672
R21968 vdd.n127 vdd.n89 0.155672
R21969 vdd.n119 vdd.n89 0.155672
R21970 vdd.n119 vdd.n118 0.155672
R21971 vdd.n118 vdd.n94 0.155672
R21972 vdd.n111 vdd.n94 0.155672
R21973 vdd.n111 vdd.n110 0.155672
R21974 vdd.n110 vdd.n98 0.155672
R21975 vdd.n103 vdd.n98 0.155672
R21976 vdd.n68 vdd.n30 0.155672
R21977 vdd.n60 vdd.n30 0.155672
R21978 vdd.n60 vdd.n59 0.155672
R21979 vdd.n59 vdd.n35 0.155672
R21980 vdd.n52 vdd.n35 0.155672
R21981 vdd.n52 vdd.n51 0.155672
R21982 vdd.n51 vdd.n39 0.155672
R21983 vdd.n44 vdd.n39 0.155672
R21984 vdd.n1829 vdd.n1791 0.155672
R21985 vdd.n1821 vdd.n1791 0.155672
R21986 vdd.n1821 vdd.n1820 0.155672
R21987 vdd.n1820 vdd.n1796 0.155672
R21988 vdd.n1813 vdd.n1796 0.155672
R21989 vdd.n1813 vdd.n1812 0.155672
R21990 vdd.n1812 vdd.n1800 0.155672
R21991 vdd.n1805 vdd.n1800 0.155672
R21992 vdd.n1888 vdd.n1850 0.155672
R21993 vdd.n1880 vdd.n1850 0.155672
R21994 vdd.n1880 vdd.n1879 0.155672
R21995 vdd.n1879 vdd.n1855 0.155672
R21996 vdd.n1872 vdd.n1855 0.155672
R21997 vdd.n1872 vdd.n1871 0.155672
R21998 vdd.n1871 vdd.n1859 0.155672
R21999 vdd.n1864 vdd.n1859 0.155672
R22000 vdd.n1727 vdd.n1689 0.155672
R22001 vdd.n1719 vdd.n1689 0.155672
R22002 vdd.n1719 vdd.n1718 0.155672
R22003 vdd.n1718 vdd.n1694 0.155672
R22004 vdd.n1711 vdd.n1694 0.155672
R22005 vdd.n1711 vdd.n1710 0.155672
R22006 vdd.n1710 vdd.n1698 0.155672
R22007 vdd.n1703 vdd.n1698 0.155672
R22008 vdd.n1786 vdd.n1748 0.155672
R22009 vdd.n1778 vdd.n1748 0.155672
R22010 vdd.n1778 vdd.n1777 0.155672
R22011 vdd.n1777 vdd.n1753 0.155672
R22012 vdd.n1770 vdd.n1753 0.155672
R22013 vdd.n1770 vdd.n1769 0.155672
R22014 vdd.n1769 vdd.n1757 0.155672
R22015 vdd.n1762 vdd.n1757 0.155672
R22016 vdd.n1626 vdd.n1588 0.155672
R22017 vdd.n1618 vdd.n1588 0.155672
R22018 vdd.n1618 vdd.n1617 0.155672
R22019 vdd.n1617 vdd.n1593 0.155672
R22020 vdd.n1610 vdd.n1593 0.155672
R22021 vdd.n1610 vdd.n1609 0.155672
R22022 vdd.n1609 vdd.n1597 0.155672
R22023 vdd.n1602 vdd.n1597 0.155672
R22024 vdd.n1685 vdd.n1647 0.155672
R22025 vdd.n1677 vdd.n1647 0.155672
R22026 vdd.n1677 vdd.n1676 0.155672
R22027 vdd.n1676 vdd.n1652 0.155672
R22028 vdd.n1669 vdd.n1652 0.155672
R22029 vdd.n1669 vdd.n1668 0.155672
R22030 vdd.n1668 vdd.n1656 0.155672
R22031 vdd.n1661 vdd.n1656 0.155672
R22032 vdd.n2181 vdd.n1986 0.152939
R22033 vdd.n1992 vdd.n1986 0.152939
R22034 vdd.n1993 vdd.n1992 0.152939
R22035 vdd.n1994 vdd.n1993 0.152939
R22036 vdd.n1995 vdd.n1994 0.152939
R22037 vdd.n1999 vdd.n1995 0.152939
R22038 vdd.n2000 vdd.n1999 0.152939
R22039 vdd.n2001 vdd.n2000 0.152939
R22040 vdd.n2002 vdd.n2001 0.152939
R22041 vdd.n2006 vdd.n2002 0.152939
R22042 vdd.n2007 vdd.n2006 0.152939
R22043 vdd.n2008 vdd.n2007 0.152939
R22044 vdd.n2156 vdd.n2008 0.152939
R22045 vdd.n2156 vdd.n2155 0.152939
R22046 vdd.n2155 vdd.n2154 0.152939
R22047 vdd.n2154 vdd.n2014 0.152939
R22048 vdd.n2019 vdd.n2014 0.152939
R22049 vdd.n2020 vdd.n2019 0.152939
R22050 vdd.n2021 vdd.n2020 0.152939
R22051 vdd.n2025 vdd.n2021 0.152939
R22052 vdd.n2026 vdd.n2025 0.152939
R22053 vdd.n2027 vdd.n2026 0.152939
R22054 vdd.n2028 vdd.n2027 0.152939
R22055 vdd.n2032 vdd.n2028 0.152939
R22056 vdd.n2033 vdd.n2032 0.152939
R22057 vdd.n2034 vdd.n2033 0.152939
R22058 vdd.n2035 vdd.n2034 0.152939
R22059 vdd.n2039 vdd.n2035 0.152939
R22060 vdd.n2040 vdd.n2039 0.152939
R22061 vdd.n2041 vdd.n2040 0.152939
R22062 vdd.n2042 vdd.n2041 0.152939
R22063 vdd.n2046 vdd.n2042 0.152939
R22064 vdd.n2047 vdd.n2046 0.152939
R22065 vdd.n2048 vdd.n2047 0.152939
R22066 vdd.n2117 vdd.n2048 0.152939
R22067 vdd.n2117 vdd.n2116 0.152939
R22068 vdd.n2116 vdd.n2115 0.152939
R22069 vdd.n2115 vdd.n2054 0.152939
R22070 vdd.n2059 vdd.n2054 0.152939
R22071 vdd.n2060 vdd.n2059 0.152939
R22072 vdd.n2061 vdd.n2060 0.152939
R22073 vdd.n2065 vdd.n2061 0.152939
R22074 vdd.n2066 vdd.n2065 0.152939
R22075 vdd.n2067 vdd.n2066 0.152939
R22076 vdd.n2068 vdd.n2067 0.152939
R22077 vdd.n2072 vdd.n2068 0.152939
R22078 vdd.n2073 vdd.n2072 0.152939
R22079 vdd.n2074 vdd.n2073 0.152939
R22080 vdd.n2075 vdd.n2074 0.152939
R22081 vdd.n2076 vdd.n2075 0.152939
R22082 vdd.n2076 vdd.n1144 0.152939
R22083 vdd.n2192 vdd.n1980 0.152939
R22084 vdd.n1894 vdd.n1203 0.152939
R22085 vdd.n1909 vdd.n1203 0.152939
R22086 vdd.n1910 vdd.n1909 0.152939
R22087 vdd.n1911 vdd.n1910 0.152939
R22088 vdd.n1911 vdd.n1192 0.152939
R22089 vdd.n1926 vdd.n1192 0.152939
R22090 vdd.n1927 vdd.n1926 0.152939
R22091 vdd.n1928 vdd.n1927 0.152939
R22092 vdd.n1928 vdd.n1181 0.152939
R22093 vdd.n1942 vdd.n1181 0.152939
R22094 vdd.n1943 vdd.n1942 0.152939
R22095 vdd.n1944 vdd.n1943 0.152939
R22096 vdd.n1944 vdd.n1169 0.152939
R22097 vdd.n1959 vdd.n1169 0.152939
R22098 vdd.n1960 vdd.n1959 0.152939
R22099 vdd.n1961 vdd.n1960 0.152939
R22100 vdd.n1961 vdd.n1157 0.152939
R22101 vdd.n1978 vdd.n1157 0.152939
R22102 vdd.n1979 vdd.n1978 0.152939
R22103 vdd.n2193 vdd.n1979 0.152939
R22104 vdd.n735 vdd.n730 0.152939
R22105 vdd.n736 vdd.n735 0.152939
R22106 vdd.n737 vdd.n736 0.152939
R22107 vdd.n738 vdd.n737 0.152939
R22108 vdd.n739 vdd.n738 0.152939
R22109 vdd.n740 vdd.n739 0.152939
R22110 vdd.n741 vdd.n740 0.152939
R22111 vdd.n742 vdd.n741 0.152939
R22112 vdd.n743 vdd.n742 0.152939
R22113 vdd.n744 vdd.n743 0.152939
R22114 vdd.n745 vdd.n744 0.152939
R22115 vdd.n746 vdd.n745 0.152939
R22116 vdd.n3365 vdd.n746 0.152939
R22117 vdd.n3365 vdd.n3364 0.152939
R22118 vdd.n3364 vdd.n3363 0.152939
R22119 vdd.n3363 vdd.n748 0.152939
R22120 vdd.n749 vdd.n748 0.152939
R22121 vdd.n750 vdd.n749 0.152939
R22122 vdd.n751 vdd.n750 0.152939
R22123 vdd.n752 vdd.n751 0.152939
R22124 vdd.n753 vdd.n752 0.152939
R22125 vdd.n754 vdd.n753 0.152939
R22126 vdd.n755 vdd.n754 0.152939
R22127 vdd.n756 vdd.n755 0.152939
R22128 vdd.n757 vdd.n756 0.152939
R22129 vdd.n758 vdd.n757 0.152939
R22130 vdd.n759 vdd.n758 0.152939
R22131 vdd.n760 vdd.n759 0.152939
R22132 vdd.n761 vdd.n760 0.152939
R22133 vdd.n762 vdd.n761 0.152939
R22134 vdd.n763 vdd.n762 0.152939
R22135 vdd.n764 vdd.n763 0.152939
R22136 vdd.n765 vdd.n764 0.152939
R22137 vdd.n766 vdd.n765 0.152939
R22138 vdd.n3319 vdd.n766 0.152939
R22139 vdd.n3319 vdd.n3318 0.152939
R22140 vdd.n3318 vdd.n3317 0.152939
R22141 vdd.n3317 vdd.n770 0.152939
R22142 vdd.n771 vdd.n770 0.152939
R22143 vdd.n772 vdd.n771 0.152939
R22144 vdd.n773 vdd.n772 0.152939
R22145 vdd.n774 vdd.n773 0.152939
R22146 vdd.n775 vdd.n774 0.152939
R22147 vdd.n776 vdd.n775 0.152939
R22148 vdd.n777 vdd.n776 0.152939
R22149 vdd.n778 vdd.n777 0.152939
R22150 vdd.n779 vdd.n778 0.152939
R22151 vdd.n780 vdd.n779 0.152939
R22152 vdd.n781 vdd.n780 0.152939
R22153 vdd.n782 vdd.n781 0.152939
R22154 vdd.n783 vdd.n782 0.152939
R22155 vdd.n727 vdd.n726 0.152939
R22156 vdd.n3416 vdd.n682 0.152939
R22157 vdd.n3417 vdd.n3416 0.152939
R22158 vdd.n3418 vdd.n3417 0.152939
R22159 vdd.n3418 vdd.n670 0.152939
R22160 vdd.n3433 vdd.n670 0.152939
R22161 vdd.n3434 vdd.n3433 0.152939
R22162 vdd.n3435 vdd.n3434 0.152939
R22163 vdd.n3435 vdd.n659 0.152939
R22164 vdd.n3449 vdd.n659 0.152939
R22165 vdd.n3450 vdd.n3449 0.152939
R22166 vdd.n3451 vdd.n3450 0.152939
R22167 vdd.n3451 vdd.n647 0.152939
R22168 vdd.n3466 vdd.n647 0.152939
R22169 vdd.n3467 vdd.n3466 0.152939
R22170 vdd.n3468 vdd.n3467 0.152939
R22171 vdd.n3468 vdd.n636 0.152939
R22172 vdd.n3485 vdd.n636 0.152939
R22173 vdd.n3486 vdd.n3485 0.152939
R22174 vdd.n3487 vdd.n3486 0.152939
R22175 vdd.n3487 vdd.n334 0.152939
R22176 vdd.n3580 vdd.n335 0.152939
R22177 vdd.n346 vdd.n335 0.152939
R22178 vdd.n347 vdd.n346 0.152939
R22179 vdd.n348 vdd.n347 0.152939
R22180 vdd.n355 vdd.n348 0.152939
R22181 vdd.n356 vdd.n355 0.152939
R22182 vdd.n357 vdd.n356 0.152939
R22183 vdd.n358 vdd.n357 0.152939
R22184 vdd.n366 vdd.n358 0.152939
R22185 vdd.n367 vdd.n366 0.152939
R22186 vdd.n368 vdd.n367 0.152939
R22187 vdd.n369 vdd.n368 0.152939
R22188 vdd.n377 vdd.n369 0.152939
R22189 vdd.n378 vdd.n377 0.152939
R22190 vdd.n379 vdd.n378 0.152939
R22191 vdd.n380 vdd.n379 0.152939
R22192 vdd.n388 vdd.n380 0.152939
R22193 vdd.n389 vdd.n388 0.152939
R22194 vdd.n390 vdd.n389 0.152939
R22195 vdd.n391 vdd.n390 0.152939
R22196 vdd.n464 vdd.n463 0.152939
R22197 vdd.n470 vdd.n463 0.152939
R22198 vdd.n471 vdd.n470 0.152939
R22199 vdd.n472 vdd.n471 0.152939
R22200 vdd.n472 vdd.n461 0.152939
R22201 vdd.n480 vdd.n461 0.152939
R22202 vdd.n481 vdd.n480 0.152939
R22203 vdd.n482 vdd.n481 0.152939
R22204 vdd.n482 vdd.n459 0.152939
R22205 vdd.n490 vdd.n459 0.152939
R22206 vdd.n491 vdd.n490 0.152939
R22207 vdd.n492 vdd.n491 0.152939
R22208 vdd.n492 vdd.n457 0.152939
R22209 vdd.n500 vdd.n457 0.152939
R22210 vdd.n501 vdd.n500 0.152939
R22211 vdd.n502 vdd.n501 0.152939
R22212 vdd.n502 vdd.n455 0.152939
R22213 vdd.n510 vdd.n455 0.152939
R22214 vdd.n511 vdd.n510 0.152939
R22215 vdd.n512 vdd.n511 0.152939
R22216 vdd.n512 vdd.n451 0.152939
R22217 vdd.n520 vdd.n451 0.152939
R22218 vdd.n521 vdd.n520 0.152939
R22219 vdd.n522 vdd.n521 0.152939
R22220 vdd.n522 vdd.n449 0.152939
R22221 vdd.n530 vdd.n449 0.152939
R22222 vdd.n531 vdd.n530 0.152939
R22223 vdd.n532 vdd.n531 0.152939
R22224 vdd.n532 vdd.n447 0.152939
R22225 vdd.n540 vdd.n447 0.152939
R22226 vdd.n541 vdd.n540 0.152939
R22227 vdd.n542 vdd.n541 0.152939
R22228 vdd.n542 vdd.n445 0.152939
R22229 vdd.n550 vdd.n445 0.152939
R22230 vdd.n551 vdd.n550 0.152939
R22231 vdd.n552 vdd.n551 0.152939
R22232 vdd.n552 vdd.n443 0.152939
R22233 vdd.n560 vdd.n443 0.152939
R22234 vdd.n561 vdd.n560 0.152939
R22235 vdd.n562 vdd.n561 0.152939
R22236 vdd.n562 vdd.n439 0.152939
R22237 vdd.n570 vdd.n439 0.152939
R22238 vdd.n571 vdd.n570 0.152939
R22239 vdd.n572 vdd.n571 0.152939
R22240 vdd.n572 vdd.n437 0.152939
R22241 vdd.n580 vdd.n437 0.152939
R22242 vdd.n581 vdd.n580 0.152939
R22243 vdd.n582 vdd.n581 0.152939
R22244 vdd.n582 vdd.n435 0.152939
R22245 vdd.n590 vdd.n435 0.152939
R22246 vdd.n591 vdd.n590 0.152939
R22247 vdd.n592 vdd.n591 0.152939
R22248 vdd.n592 vdd.n433 0.152939
R22249 vdd.n600 vdd.n433 0.152939
R22250 vdd.n601 vdd.n600 0.152939
R22251 vdd.n602 vdd.n601 0.152939
R22252 vdd.n602 vdd.n431 0.152939
R22253 vdd.n610 vdd.n431 0.152939
R22254 vdd.n611 vdd.n610 0.152939
R22255 vdd.n612 vdd.n611 0.152939
R22256 vdd.n612 vdd.n429 0.152939
R22257 vdd.n619 vdd.n429 0.152939
R22258 vdd.n3532 vdd.n619 0.152939
R22259 vdd.n3410 vdd.n3409 0.152939
R22260 vdd.n3410 vdd.n675 0.152939
R22261 vdd.n3424 vdd.n675 0.152939
R22262 vdd.n3425 vdd.n3424 0.152939
R22263 vdd.n3426 vdd.n3425 0.152939
R22264 vdd.n3426 vdd.n665 0.152939
R22265 vdd.n3441 vdd.n665 0.152939
R22266 vdd.n3442 vdd.n3441 0.152939
R22267 vdd.n3443 vdd.n3442 0.152939
R22268 vdd.n3443 vdd.n652 0.152939
R22269 vdd.n3457 vdd.n652 0.152939
R22270 vdd.n3458 vdd.n3457 0.152939
R22271 vdd.n3459 vdd.n3458 0.152939
R22272 vdd.n3459 vdd.n641 0.152939
R22273 vdd.n3474 vdd.n641 0.152939
R22274 vdd.n3475 vdd.n3474 0.152939
R22275 vdd.n3476 vdd.n3475 0.152939
R22276 vdd.n3478 vdd.n3476 0.152939
R22277 vdd.n3478 vdd.n3477 0.152939
R22278 vdd.n3477 vdd.n630 0.152939
R22279 vdd.n3495 vdd.n630 0.152939
R22280 vdd.n3496 vdd.n3495 0.152939
R22281 vdd.n3497 vdd.n3496 0.152939
R22282 vdd.n3497 vdd.n628 0.152939
R22283 vdd.n3502 vdd.n628 0.152939
R22284 vdd.n3503 vdd.n3502 0.152939
R22285 vdd.n3504 vdd.n3503 0.152939
R22286 vdd.n3504 vdd.n626 0.152939
R22287 vdd.n3509 vdd.n626 0.152939
R22288 vdd.n3510 vdd.n3509 0.152939
R22289 vdd.n3511 vdd.n3510 0.152939
R22290 vdd.n3511 vdd.n624 0.152939
R22291 vdd.n3517 vdd.n624 0.152939
R22292 vdd.n3518 vdd.n3517 0.152939
R22293 vdd.n3519 vdd.n3518 0.152939
R22294 vdd.n3519 vdd.n622 0.152939
R22295 vdd.n3524 vdd.n622 0.152939
R22296 vdd.n3525 vdd.n3524 0.152939
R22297 vdd.n3526 vdd.n3525 0.152939
R22298 vdd.n3526 vdd.n620 0.152939
R22299 vdd.n3531 vdd.n620 0.152939
R22300 vdd.n3408 vdd.n687 0.152939
R22301 vdd.n2204 vdd.n1147 0.152939
R22302 vdd.n1510 vdd.n1266 0.152939
R22303 vdd.n1511 vdd.n1510 0.152939
R22304 vdd.n1512 vdd.n1511 0.152939
R22305 vdd.n1512 vdd.n1254 0.152939
R22306 vdd.n1527 vdd.n1254 0.152939
R22307 vdd.n1528 vdd.n1527 0.152939
R22308 vdd.n1529 vdd.n1528 0.152939
R22309 vdd.n1529 vdd.n1244 0.152939
R22310 vdd.n1544 vdd.n1244 0.152939
R22311 vdd.n1545 vdd.n1544 0.152939
R22312 vdd.n1546 vdd.n1545 0.152939
R22313 vdd.n1546 vdd.n1231 0.152939
R22314 vdd.n1560 vdd.n1231 0.152939
R22315 vdd.n1561 vdd.n1560 0.152939
R22316 vdd.n1562 vdd.n1561 0.152939
R22317 vdd.n1562 vdd.n1220 0.152939
R22318 vdd.n1577 vdd.n1220 0.152939
R22319 vdd.n1578 vdd.n1577 0.152939
R22320 vdd.n1579 vdd.n1578 0.152939
R22321 vdd.n1579 vdd.n1209 0.152939
R22322 vdd.n1900 vdd.n1209 0.152939
R22323 vdd.n1901 vdd.n1900 0.152939
R22324 vdd.n1902 vdd.n1901 0.152939
R22325 vdd.n1902 vdd.n1197 0.152939
R22326 vdd.n1917 vdd.n1197 0.152939
R22327 vdd.n1918 vdd.n1917 0.152939
R22328 vdd.n1919 vdd.n1918 0.152939
R22329 vdd.n1919 vdd.n1187 0.152939
R22330 vdd.n1934 vdd.n1187 0.152939
R22331 vdd.n1935 vdd.n1934 0.152939
R22332 vdd.n1936 vdd.n1935 0.152939
R22333 vdd.n1936 vdd.n1174 0.152939
R22334 vdd.n1950 vdd.n1174 0.152939
R22335 vdd.n1951 vdd.n1950 0.152939
R22336 vdd.n1952 vdd.n1951 0.152939
R22337 vdd.n1952 vdd.n1164 0.152939
R22338 vdd.n1967 vdd.n1164 0.152939
R22339 vdd.n1968 vdd.n1967 0.152939
R22340 vdd.n1971 vdd.n1968 0.152939
R22341 vdd.n1971 vdd.n1970 0.152939
R22342 vdd.n1970 vdd.n1969 0.152939
R22343 vdd.n1502 vdd.n1271 0.152939
R22344 vdd.n1495 vdd.n1271 0.152939
R22345 vdd.n1495 vdd.n1494 0.152939
R22346 vdd.n1494 vdd.n1493 0.152939
R22347 vdd.n1493 vdd.n1308 0.152939
R22348 vdd.n1489 vdd.n1308 0.152939
R22349 vdd.n1489 vdd.n1488 0.152939
R22350 vdd.n1488 vdd.n1487 0.152939
R22351 vdd.n1487 vdd.n1314 0.152939
R22352 vdd.n1483 vdd.n1314 0.152939
R22353 vdd.n1483 vdd.n1482 0.152939
R22354 vdd.n1482 vdd.n1481 0.152939
R22355 vdd.n1481 vdd.n1320 0.152939
R22356 vdd.n1477 vdd.n1320 0.152939
R22357 vdd.n1477 vdd.n1476 0.152939
R22358 vdd.n1476 vdd.n1475 0.152939
R22359 vdd.n1475 vdd.n1326 0.152939
R22360 vdd.n1471 vdd.n1326 0.152939
R22361 vdd.n1471 vdd.n1470 0.152939
R22362 vdd.n1470 vdd.n1469 0.152939
R22363 vdd.n1469 vdd.n1334 0.152939
R22364 vdd.n1465 vdd.n1334 0.152939
R22365 vdd.n1465 vdd.n1464 0.152939
R22366 vdd.n1464 vdd.n1463 0.152939
R22367 vdd.n1463 vdd.n1340 0.152939
R22368 vdd.n1459 vdd.n1340 0.152939
R22369 vdd.n1459 vdd.n1458 0.152939
R22370 vdd.n1458 vdd.n1457 0.152939
R22371 vdd.n1457 vdd.n1346 0.152939
R22372 vdd.n1453 vdd.n1346 0.152939
R22373 vdd.n1453 vdd.n1452 0.152939
R22374 vdd.n1452 vdd.n1451 0.152939
R22375 vdd.n1451 vdd.n1352 0.152939
R22376 vdd.n1447 vdd.n1352 0.152939
R22377 vdd.n1447 vdd.n1446 0.152939
R22378 vdd.n1446 vdd.n1445 0.152939
R22379 vdd.n1445 vdd.n1358 0.152939
R22380 vdd.n1441 vdd.n1358 0.152939
R22381 vdd.n1441 vdd.n1440 0.152939
R22382 vdd.n1440 vdd.n1439 0.152939
R22383 vdd.n1439 vdd.n1364 0.152939
R22384 vdd.n1432 vdd.n1364 0.152939
R22385 vdd.n1432 vdd.n1431 0.152939
R22386 vdd.n1431 vdd.n1430 0.152939
R22387 vdd.n1430 vdd.n1369 0.152939
R22388 vdd.n1426 vdd.n1369 0.152939
R22389 vdd.n1426 vdd.n1425 0.152939
R22390 vdd.n1425 vdd.n1424 0.152939
R22391 vdd.n1424 vdd.n1375 0.152939
R22392 vdd.n1420 vdd.n1375 0.152939
R22393 vdd.n1420 vdd.n1419 0.152939
R22394 vdd.n1419 vdd.n1418 0.152939
R22395 vdd.n1418 vdd.n1381 0.152939
R22396 vdd.n1414 vdd.n1381 0.152939
R22397 vdd.n1414 vdd.n1413 0.152939
R22398 vdd.n1413 vdd.n1412 0.152939
R22399 vdd.n1412 vdd.n1387 0.152939
R22400 vdd.n1408 vdd.n1387 0.152939
R22401 vdd.n1408 vdd.n1407 0.152939
R22402 vdd.n1407 vdd.n1406 0.152939
R22403 vdd.n1406 vdd.n1393 0.152939
R22404 vdd.n1402 vdd.n1393 0.152939
R22405 vdd.n1402 vdd.n1401 0.152939
R22406 vdd.n1504 vdd.n1503 0.152939
R22407 vdd.n1504 vdd.n1260 0.152939
R22408 vdd.n1519 vdd.n1260 0.152939
R22409 vdd.n1520 vdd.n1519 0.152939
R22410 vdd.n1521 vdd.n1520 0.152939
R22411 vdd.n1521 vdd.n1249 0.152939
R22412 vdd.n1536 vdd.n1249 0.152939
R22413 vdd.n1537 vdd.n1536 0.152939
R22414 vdd.n1538 vdd.n1537 0.152939
R22415 vdd.n1538 vdd.n1238 0.152939
R22416 vdd.n1552 vdd.n1238 0.152939
R22417 vdd.n1553 vdd.n1552 0.152939
R22418 vdd.n1554 vdd.n1553 0.152939
R22419 vdd.n1554 vdd.n1226 0.152939
R22420 vdd.n1569 vdd.n1226 0.152939
R22421 vdd.n1570 vdd.n1569 0.152939
R22422 vdd.n1571 vdd.n1570 0.152939
R22423 vdd.n1571 vdd.n1215 0.152939
R22424 vdd.n1585 vdd.n1215 0.152939
R22425 vdd.n1586 vdd.n1585 0.152939
R22426 vdd.n1507 vdd.t100 0.113865
R22427 vdd.n2491 vdd.t18 0.113865
R22428 vdd.n2558 vdd.t293 0.113865
R22429 vdd.n3041 vdd.t11 0.113865
R22430 vdd.n3108 vdd.t55 0.113865
R22431 vdd.t70 vdd.n386 0.113865
R22432 vdd.n2182 vdd.n1980 0.110256
R22433 vdd.n3398 vdd.n727 0.110256
R22434 vdd.n3275 vdd.n687 0.110256
R22435 vdd.n2205 vdd.n2204 0.110256
R22436 vdd.n1894 vdd.n1893 0.0695946
R22437 vdd.n3581 vdd.n334 0.0695946
R22438 vdd.n3581 vdd.n3580 0.0695946
R22439 vdd.n1893 vdd.n1586 0.0695946
R22440 vdd.n2182 vdd.n2181 0.0431829
R22441 vdd.n2205 vdd.n1144 0.0431829
R22442 vdd.n3398 vdd.n730 0.0431829
R22443 vdd.n3275 vdd.n783 0.0431829
R22444 vdd vdd.n28 0.00833333
R22445 a_n2650_13878.n88 a_n2650_13878.t98 512.366
R22446 a_n2650_13878.n87 a_n2650_13878.t77 512.366
R22447 a_n2650_13878.n80 a_n2650_13878.t82 512.366
R22448 a_n2650_13878.n86 a_n2650_13878.t71 512.366
R22449 a_n2650_13878.n85 a_n2650_13878.t87 512.366
R22450 a_n2650_13878.n81 a_n2650_13878.t95 512.366
R22451 a_n2650_13878.n84 a_n2650_13878.t96 512.366
R22452 a_n2650_13878.n83 a_n2650_13878.t66 512.366
R22453 a_n2650_13878.n82 a_n2650_13878.t79 512.366
R22454 a_n2650_13878.n70 a_n2650_13878.t42 533.335
R22455 a_n2650_13878.n106 a_n2650_13878.t44 512.366
R22456 a_n2650_13878.n105 a_n2650_13878.t12 512.366
R22457 a_n2650_13878.n77 a_n2650_13878.t28 512.366
R22458 a_n2650_13878.n104 a_n2650_13878.t36 512.366
R22459 a_n2650_13878.n103 a_n2650_13878.t38 512.366
R22460 a_n2650_13878.n78 a_n2650_13878.t16 512.366
R22461 a_n2650_13878.n102 a_n2650_13878.t26 512.366
R22462 a_n2650_13878.n101 a_n2650_13878.t46 512.366
R22463 a_n2650_13878.n79 a_n2650_13878.t40 512.366
R22464 a_n2650_13878.n133 a_n2650_13878.t30 512.366
R22465 a_n2650_13878.n134 a_n2650_13878.t34 512.366
R22466 a_n2650_13878.n74 a_n2650_13878.t32 512.366
R22467 a_n2650_13878.n135 a_n2650_13878.t22 512.366
R22468 a_n2650_13878.n136 a_n2650_13878.t14 512.366
R22469 a_n2650_13878.n137 a_n2650_13878.t8 512.366
R22470 a_n2650_13878.n138 a_n2650_13878.t24 512.366
R22471 a_n2650_13878.n73 a_n2650_13878.t18 512.366
R22472 a_n2650_13878.n139 a_n2650_13878.t10 512.366
R22473 a_n2650_13878.n126 a_n2650_13878.t70 512.366
R22474 a_n2650_13878.n127 a_n2650_13878.t93 512.366
R22475 a_n2650_13878.n76 a_n2650_13878.t94 512.366
R22476 a_n2650_13878.n128 a_n2650_13878.t68 512.366
R22477 a_n2650_13878.n129 a_n2650_13878.t90 512.366
R22478 a_n2650_13878.n130 a_n2650_13878.t91 512.366
R22479 a_n2650_13878.n131 a_n2650_13878.t65 512.366
R22480 a_n2650_13878.n75 a_n2650_13878.t76 512.366
R22481 a_n2650_13878.n132 a_n2650_13878.t86 512.366
R22482 a_n2650_13878.n118 a_n2650_13878.t84 512.366
R22483 a_n2650_13878.n117 a_n2650_13878.t74 512.366
R22484 a_n2650_13878.n116 a_n2650_13878.t64 512.366
R22485 a_n2650_13878.n120 a_n2650_13878.t92 512.366
R22486 a_n2650_13878.n119 a_n2650_13878.t81 512.366
R22487 a_n2650_13878.n115 a_n2650_13878.t80 512.366
R22488 a_n2650_13878.n122 a_n2650_13878.t88 512.366
R22489 a_n2650_13878.n121 a_n2650_13878.t72 512.366
R22490 a_n2650_13878.n114 a_n2650_13878.t73 512.366
R22491 a_n2650_13878.n124 a_n2650_13878.t75 512.366
R22492 a_n2650_13878.n123 a_n2650_13878.t85 512.366
R22493 a_n2650_13878.n113 a_n2650_13878.t99 512.366
R22494 a_n2650_13878.n1 a_n2650_13878.n69 70.1674
R22495 a_n2650_13878.n70 a_n2650_13878.n79 20.9683
R22496 a_n2650_13878.n16 a_n2650_13878.n47 70.1674
R22497 a_n2650_13878.n20 a_n2650_13878.n40 70.1674
R22498 a_n2650_13878.n132 a_n2650_13878.n40 20.9683
R22499 a_n2650_13878.n39 a_n2650_13878.n20 74.73
R22500 a_n2650_13878.n39 a_n2650_13878.n75 11.843
R22501 a_n2650_13878.n19 a_n2650_13878.n38 80.4688
R22502 a_n2650_13878.n131 a_n2650_13878.n38 0.365327
R22503 a_n2650_13878.n37 a_n2650_13878.n19 75.0448
R22504 a_n2650_13878.n21 a_n2650_13878.n36 70.1674
R22505 a_n2650_13878.n128 a_n2650_13878.n36 20.9683
R22506 a_n2650_13878.n35 a_n2650_13878.n21 70.3058
R22507 a_n2650_13878.n35 a_n2650_13878.n76 20.6913
R22508 a_n2650_13878.n22 a_n2650_13878.n34 75.3623
R22509 a_n2650_13878.n127 a_n2650_13878.n34 10.5784
R22510 a_n2650_13878.n126 a_n2650_13878.n22 161.3
R22511 a_n2650_13878.n139 a_n2650_13878.n47 20.9683
R22512 a_n2650_13878.n46 a_n2650_13878.n16 74.73
R22513 a_n2650_13878.n46 a_n2650_13878.n73 11.843
R22514 a_n2650_13878.n15 a_n2650_13878.n45 80.4688
R22515 a_n2650_13878.n138 a_n2650_13878.n45 0.365327
R22516 a_n2650_13878.n44 a_n2650_13878.n15 75.0448
R22517 a_n2650_13878.n17 a_n2650_13878.n43 70.1674
R22518 a_n2650_13878.n135 a_n2650_13878.n43 20.9683
R22519 a_n2650_13878.n42 a_n2650_13878.n17 70.3058
R22520 a_n2650_13878.n42 a_n2650_13878.n74 20.6913
R22521 a_n2650_13878.n18 a_n2650_13878.n41 75.3623
R22522 a_n2650_13878.n134 a_n2650_13878.n41 10.5784
R22523 a_n2650_13878.n133 a_n2650_13878.n18 161.3
R22524 a_n2650_13878.n7 a_n2650_13878.n56 70.1674
R22525 a_n2650_13878.n9 a_n2650_13878.n53 70.1674
R22526 a_n2650_13878.n11 a_n2650_13878.n51 70.1674
R22527 a_n2650_13878.n13 a_n2650_13878.n49 70.1674
R22528 a_n2650_13878.n49 a_n2650_13878.n113 20.9683
R22529 a_n2650_13878.n48 a_n2650_13878.n14 75.0448
R22530 a_n2650_13878.n123 a_n2650_13878.n48 11.2134
R22531 a_n2650_13878.n14 a_n2650_13878.n124 161.3
R22532 a_n2650_13878.n51 a_n2650_13878.n114 20.9683
R22533 a_n2650_13878.n50 a_n2650_13878.n12 75.0448
R22534 a_n2650_13878.n121 a_n2650_13878.n50 11.2134
R22535 a_n2650_13878.n12 a_n2650_13878.n122 161.3
R22536 a_n2650_13878.n53 a_n2650_13878.n115 20.9683
R22537 a_n2650_13878.n52 a_n2650_13878.n10 75.0448
R22538 a_n2650_13878.n119 a_n2650_13878.n52 11.2134
R22539 a_n2650_13878.n10 a_n2650_13878.n120 161.3
R22540 a_n2650_13878.n56 a_n2650_13878.n116 20.9683
R22541 a_n2650_13878.n54 a_n2650_13878.n8 75.0448
R22542 a_n2650_13878.n117 a_n2650_13878.n54 11.2134
R22543 a_n2650_13878.n8 a_n2650_13878.n118 161.3
R22544 a_n2650_13878.n62 a_n2650_13878.n33 74.73
R22545 a_n2650_13878.n101 a_n2650_13878.n62 11.843
R22546 a_n2650_13878.n61 a_n2650_13878.n5 80.4688
R22547 a_n2650_13878.n61 a_n2650_13878.n102 0.365327
R22548 a_n2650_13878.n5 a_n2650_13878.n60 75.0448
R22549 a_n2650_13878.n59 a_n2650_13878.n4 70.1674
R22550 a_n2650_13878.n104 a_n2650_13878.n59 20.9683
R22551 a_n2650_13878.n4 a_n2650_13878.n58 70.3058
R22552 a_n2650_13878.n58 a_n2650_13878.n77 20.6913
R22553 a_n2650_13878.n57 a_n2650_13878.n6 75.3623
R22554 a_n2650_13878.n105 a_n2650_13878.n57 10.5784
R22555 a_n2650_13878.n6 a_n2650_13878.n106 161.3
R22556 a_n2650_13878.n33 a_n2650_13878.n70 70.1674
R22557 a_n2650_13878.n69 a_n2650_13878.n82 20.9683
R22558 a_n2650_13878.n68 a_n2650_13878.n1 74.73
R22559 a_n2650_13878.n83 a_n2650_13878.n68 11.843
R22560 a_n2650_13878.n67 a_n2650_13878.n0 80.4688
R22561 a_n2650_13878.n67 a_n2650_13878.n84 0.365327
R22562 a_n2650_13878.n0 a_n2650_13878.n66 75.0448
R22563 a_n2650_13878.n65 a_n2650_13878.n2 70.1674
R22564 a_n2650_13878.n86 a_n2650_13878.n65 20.9683
R22565 a_n2650_13878.n2 a_n2650_13878.n64 70.3058
R22566 a_n2650_13878.n64 a_n2650_13878.n80 20.6913
R22567 a_n2650_13878.n63 a_n2650_13878.n3 75.3623
R22568 a_n2650_13878.n87 a_n2650_13878.n63 10.5784
R22569 a_n2650_13878.n3 a_n2650_13878.n88 161.3
R22570 a_n2650_13878.n31 a_n2650_13878.n98 81.2902
R22571 a_n2650_13878.n32 a_n2650_13878.n92 81.2902
R22572 a_n2650_13878.n23 a_n2650_13878.n89 81.2902
R22573 a_n2650_13878.n31 a_n2650_13878.n99 80.9324
R22574 a_n2650_13878.n25 a_n2650_13878.n100 80.9324
R22575 a_n2650_13878.n25 a_n2650_13878.n97 80.9324
R22576 a_n2650_13878.n25 a_n2650_13878.n96 80.9324
R22577 a_n2650_13878.n24 a_n2650_13878.n95 80.9324
R22578 a_n2650_13878.n32 a_n2650_13878.n93 80.9324
R22579 a_n2650_13878.n23 a_n2650_13878.n94 80.9324
R22580 a_n2650_13878.n23 a_n2650_13878.n91 80.9324
R22581 a_n2650_13878.n23 a_n2650_13878.n90 80.9324
R22582 a_n2650_13878.n29 a_n2650_13878.t31 74.6477
R22583 a_n2650_13878.n26 a_n2650_13878.t43 74.6477
R22584 a_n2650_13878.n111 a_n2650_13878.t45 74.2899
R22585 a_n2650_13878.n28 a_n2650_13878.t21 74.2897
R22586 a_n2650_13878.n28 a_n2650_13878.n141 70.6783
R22587 a_n2650_13878.n30 a_n2650_13878.n72 70.6783
R22588 a_n2650_13878.n29 a_n2650_13878.n71 70.6783
R22589 a_n2650_13878.n26 a_n2650_13878.n107 70.6783
R22590 a_n2650_13878.n26 a_n2650_13878.n108 70.6783
R22591 a_n2650_13878.n27 a_n2650_13878.n109 70.6783
R22592 a_n2650_13878.n27 a_n2650_13878.n110 70.6783
R22593 a_n2650_13878.n142 a_n2650_13878.n30 70.6782
R22594 a_n2650_13878.n88 a_n2650_13878.n87 48.2005
R22595 a_n2650_13878.n65 a_n2650_13878.n85 20.9683
R22596 a_n2650_13878.n84 a_n2650_13878.n81 48.2005
R22597 a_n2650_13878.t69 a_n2650_13878.n69 533.335
R22598 a_n2650_13878.n106 a_n2650_13878.n105 48.2005
R22599 a_n2650_13878.n59 a_n2650_13878.n103 20.9683
R22600 a_n2650_13878.n102 a_n2650_13878.n78 48.2005
R22601 a_n2650_13878.n134 a_n2650_13878.n133 48.2005
R22602 a_n2650_13878.n136 a_n2650_13878.n43 20.9683
R22603 a_n2650_13878.n138 a_n2650_13878.n137 48.2005
R22604 a_n2650_13878.t20 a_n2650_13878.n47 533.335
R22605 a_n2650_13878.n127 a_n2650_13878.n126 48.2005
R22606 a_n2650_13878.n129 a_n2650_13878.n36 20.9683
R22607 a_n2650_13878.n131 a_n2650_13878.n130 48.2005
R22608 a_n2650_13878.t67 a_n2650_13878.n40 533.335
R22609 a_n2650_13878.n118 a_n2650_13878.n117 48.2005
R22610 a_n2650_13878.t89 a_n2650_13878.n56 533.335
R22611 a_n2650_13878.n120 a_n2650_13878.n119 48.2005
R22612 a_n2650_13878.t97 a_n2650_13878.n53 533.335
R22613 a_n2650_13878.n122 a_n2650_13878.n121 48.2005
R22614 a_n2650_13878.t83 a_n2650_13878.n51 533.335
R22615 a_n2650_13878.n124 a_n2650_13878.n123 48.2005
R22616 a_n2650_13878.t78 a_n2650_13878.n49 533.335
R22617 a_n2650_13878.n86 a_n2650_13878.n64 21.4216
R22618 a_n2650_13878.n104 a_n2650_13878.n58 21.4216
R22619 a_n2650_13878.n135 a_n2650_13878.n42 21.4216
R22620 a_n2650_13878.n128 a_n2650_13878.n35 21.4216
R22621 a_n2650_13878.n24 a_n2650_13878.n23 31.7747
R22622 a_n2650_13878.n68 a_n2650_13878.n82 34.4824
R22623 a_n2650_13878.n62 a_n2650_13878.n79 34.4824
R22624 a_n2650_13878.n139 a_n2650_13878.n46 34.4824
R22625 a_n2650_13878.n132 a_n2650_13878.n39 34.4824
R22626 a_n2650_13878.n85 a_n2650_13878.n66 35.3134
R22627 a_n2650_13878.n66 a_n2650_13878.n81 11.2134
R22628 a_n2650_13878.n103 a_n2650_13878.n60 35.3134
R22629 a_n2650_13878.n60 a_n2650_13878.n78 11.2134
R22630 a_n2650_13878.n136 a_n2650_13878.n44 35.3134
R22631 a_n2650_13878.n137 a_n2650_13878.n44 11.2134
R22632 a_n2650_13878.n129 a_n2650_13878.n37 35.3134
R22633 a_n2650_13878.n130 a_n2650_13878.n37 11.2134
R22634 a_n2650_13878.n54 a_n2650_13878.n116 35.3134
R22635 a_n2650_13878.n52 a_n2650_13878.n115 35.3134
R22636 a_n2650_13878.n50 a_n2650_13878.n114 35.3134
R22637 a_n2650_13878.n48 a_n2650_13878.n113 35.3134
R22638 a_n2650_13878.n33 a_n2650_13878.n25 23.891
R22639 a_n2650_13878.n63 a_n2650_13878.n80 36.139
R22640 a_n2650_13878.n57 a_n2650_13878.n77 36.139
R22641 a_n2650_13878.n74 a_n2650_13878.n41 36.139
R22642 a_n2650_13878.n76 a_n2650_13878.n34 36.139
R22643 a_n2650_13878.n22 a_n2650_13878.n125 13.3641
R22644 a_n2650_13878.n1 a_n2650_13878.n55 13.1596
R22645 a_n2650_13878.n112 a_n2650_13878.n6 11.8547
R22646 a_n2650_13878.n28 a_n2650_13878.n140 10.2167
R22647 a_n2650_13878.n7 a_n2650_13878.n55 9.99103
R22648 a_n2650_13878.n125 a_n2650_13878.n14 9.99103
R22649 a_n2650_13878.n140 a_n2650_13878.n16 8.01944
R22650 a_n2650_13878.n112 a_n2650_13878.n111 6.37334
R22651 a_n2650_13878.n140 a_n2650_13878.n55 5.3452
R22652 a_n2650_13878.n18 a_n2650_13878.n20 4.07247
R22653 a_n2650_13878.n33 a_n2650_13878.n3 4.06674
R22654 a_n2650_13878.n141 a_n2650_13878.t19 3.61217
R22655 a_n2650_13878.n141 a_n2650_13878.t11 3.61217
R22656 a_n2650_13878.n72 a_n2650_13878.t23 3.61217
R22657 a_n2650_13878.n72 a_n2650_13878.t15 3.61217
R22658 a_n2650_13878.n71 a_n2650_13878.t35 3.61217
R22659 a_n2650_13878.n71 a_n2650_13878.t33 3.61217
R22660 a_n2650_13878.n107 a_n2650_13878.t47 3.61217
R22661 a_n2650_13878.n107 a_n2650_13878.t41 3.61217
R22662 a_n2650_13878.n108 a_n2650_13878.t17 3.61217
R22663 a_n2650_13878.n108 a_n2650_13878.t27 3.61217
R22664 a_n2650_13878.n109 a_n2650_13878.t37 3.61217
R22665 a_n2650_13878.n109 a_n2650_13878.t39 3.61217
R22666 a_n2650_13878.n110 a_n2650_13878.t13 3.61217
R22667 a_n2650_13878.n110 a_n2650_13878.t29 3.61217
R22668 a_n2650_13878.t9 a_n2650_13878.n142 3.61217
R22669 a_n2650_13878.n142 a_n2650_13878.t25 3.61217
R22670 a_n2650_13878.n98 a_n2650_13878.t55 2.82907
R22671 a_n2650_13878.n98 a_n2650_13878.t59 2.82907
R22672 a_n2650_13878.n99 a_n2650_13878.t3 2.82907
R22673 a_n2650_13878.n99 a_n2650_13878.t52 2.82907
R22674 a_n2650_13878.n100 a_n2650_13878.t1 2.82907
R22675 a_n2650_13878.n100 a_n2650_13878.t4 2.82907
R22676 a_n2650_13878.n97 a_n2650_13878.t58 2.82907
R22677 a_n2650_13878.n97 a_n2650_13878.t54 2.82907
R22678 a_n2650_13878.n96 a_n2650_13878.t49 2.82907
R22679 a_n2650_13878.n96 a_n2650_13878.t63 2.82907
R22680 a_n2650_13878.n95 a_n2650_13878.t2 2.82907
R22681 a_n2650_13878.n95 a_n2650_13878.t6 2.82907
R22682 a_n2650_13878.n92 a_n2650_13878.t60 2.82907
R22683 a_n2650_13878.n92 a_n2650_13878.t48 2.82907
R22684 a_n2650_13878.n93 a_n2650_13878.t51 2.82907
R22685 a_n2650_13878.n93 a_n2650_13878.t61 2.82907
R22686 a_n2650_13878.n94 a_n2650_13878.t5 2.82907
R22687 a_n2650_13878.n94 a_n2650_13878.t57 2.82907
R22688 a_n2650_13878.n91 a_n2650_13878.t56 2.82907
R22689 a_n2650_13878.n91 a_n2650_13878.t7 2.82907
R22690 a_n2650_13878.n90 a_n2650_13878.t50 2.82907
R22691 a_n2650_13878.n90 a_n2650_13878.t53 2.82907
R22692 a_n2650_13878.n89 a_n2650_13878.t0 2.82907
R22693 a_n2650_13878.n89 a_n2650_13878.t62 2.82907
R22694 a_n2650_13878.n125 a_n2650_13878.n112 1.30542
R22695 a_n2650_13878.n11 a_n2650_13878.n10 1.04595
R22696 a_n2650_13878.n67 a_n2650_13878.n83 47.835
R22697 a_n2650_13878.n61 a_n2650_13878.n101 47.835
R22698 a_n2650_13878.n73 a_n2650_13878.n45 47.835
R22699 a_n2650_13878.n75 a_n2650_13878.n38 47.835
R22700 a_n2650_13878.n20 a_n2650_13878.n19 1.13686
R22701 a_n2650_13878.n16 a_n2650_13878.n15 1.13686
R22702 a_n2650_13878.n1 a_n2650_13878.n0 1.13686
R22703 a_n2650_13878.n33 a_n2650_13878.n5 1.10471
R22704 a_n2650_13878.n23 a_n2650_13878.n32 1.07378
R22705 a_n2650_13878.n21 a_n2650_13878.n22 0.758076
R22706 a_n2650_13878.n19 a_n2650_13878.n21 0.758076
R22707 a_n2650_13878.n17 a_n2650_13878.n18 0.758076
R22708 a_n2650_13878.n15 a_n2650_13878.n17 0.758076
R22709 a_n2650_13878.n14 a_n2650_13878.n13 0.758076
R22710 a_n2650_13878.n12 a_n2650_13878.n11 0.758076
R22711 a_n2650_13878.n10 a_n2650_13878.n9 0.758076
R22712 a_n2650_13878.n8 a_n2650_13878.n7 0.758076
R22713 a_n2650_13878.n6 a_n2650_13878.n4 0.758076
R22714 a_n2650_13878.n5 a_n2650_13878.n4 0.758076
R22715 a_n2650_13878.n3 a_n2650_13878.n2 0.758076
R22716 a_n2650_13878.n0 a_n2650_13878.n2 0.758076
R22717 a_n2650_13878.n25 a_n2650_13878.n31 0.716017
R22718 a_n2650_13878.n30 a_n2650_13878.n28 0.716017
R22719 a_n2650_13878.n30 a_n2650_13878.n29 0.716017
R22720 a_n2650_13878.n27 a_n2650_13878.n26 0.716017
R22721 a_n2650_13878.n111 a_n2650_13878.n27 0.716017
R22722 a_n2650_13878.n25 a_n2650_13878.n24 0.716017
R22723 a_n2650_13878.n13 a_n2650_13878.n12 0.67853
R22724 a_n2650_13878.n9 a_n2650_13878.n8 0.67853
R22725 a_n2472_13878.n25 a_n2472_13878.n24 98.9632
R22726 a_n2472_13878.n2 a_n2472_13878.n0 98.7517
R22727 a_n2472_13878.n20 a_n2472_13878.n19 98.6055
R22728 a_n2472_13878.n22 a_n2472_13878.n21 98.6055
R22729 a_n2472_13878.n24 a_n2472_13878.n23 98.6055
R22730 a_n2472_13878.n8 a_n2472_13878.n7 98.6055
R22731 a_n2472_13878.n6 a_n2472_13878.n5 98.6055
R22732 a_n2472_13878.n4 a_n2472_13878.n3 98.6055
R22733 a_n2472_13878.n2 a_n2472_13878.n1 98.6055
R22734 a_n2472_13878.n18 a_n2472_13878.n17 98.6054
R22735 a_n2472_13878.n10 a_n2472_13878.t21 74.6477
R22736 a_n2472_13878.n15 a_n2472_13878.t22 74.2899
R22737 a_n2472_13878.n12 a_n2472_13878.t23 74.2899
R22738 a_n2472_13878.n11 a_n2472_13878.t20 74.2899
R22739 a_n2472_13878.n14 a_n2472_13878.n13 70.6783
R22740 a_n2472_13878.n10 a_n2472_13878.n9 70.6783
R22741 a_n2472_13878.n16 a_n2472_13878.n8 15.0004
R22742 a_n2472_13878.n18 a_n2472_13878.n16 12.2917
R22743 a_n2472_13878.n16 a_n2472_13878.n15 7.67184
R22744 a_n2472_13878.n17 a_n2472_13878.t16 3.61217
R22745 a_n2472_13878.n17 a_n2472_13878.t5 3.61217
R22746 a_n2472_13878.n19 a_n2472_13878.t8 3.61217
R22747 a_n2472_13878.n19 a_n2472_13878.t9 3.61217
R22748 a_n2472_13878.n21 a_n2472_13878.t17 3.61217
R22749 a_n2472_13878.n21 a_n2472_13878.t18 3.61217
R22750 a_n2472_13878.n23 a_n2472_13878.t0 3.61217
R22751 a_n2472_13878.n23 a_n2472_13878.t10 3.61217
R22752 a_n2472_13878.n13 a_n2472_13878.t26 3.61217
R22753 a_n2472_13878.n13 a_n2472_13878.t27 3.61217
R22754 a_n2472_13878.n9 a_n2472_13878.t24 3.61217
R22755 a_n2472_13878.n9 a_n2472_13878.t25 3.61217
R22756 a_n2472_13878.n7 a_n2472_13878.t11 3.61217
R22757 a_n2472_13878.n7 a_n2472_13878.t1 3.61217
R22758 a_n2472_13878.n5 a_n2472_13878.t14 3.61217
R22759 a_n2472_13878.n5 a_n2472_13878.t3 3.61217
R22760 a_n2472_13878.n3 a_n2472_13878.t2 3.61217
R22761 a_n2472_13878.n3 a_n2472_13878.t4 3.61217
R22762 a_n2472_13878.n1 a_n2472_13878.t12 3.61217
R22763 a_n2472_13878.n1 a_n2472_13878.t6 3.61217
R22764 a_n2472_13878.n0 a_n2472_13878.t15 3.61217
R22765 a_n2472_13878.n0 a_n2472_13878.t7 3.61217
R22766 a_n2472_13878.n25 a_n2472_13878.t13 3.61217
R22767 a_n2472_13878.t19 a_n2472_13878.n25 3.61217
R22768 a_n2472_13878.n11 a_n2472_13878.n10 0.358259
R22769 a_n2472_13878.n14 a_n2472_13878.n12 0.358259
R22770 a_n2472_13878.n15 a_n2472_13878.n14 0.358259
R22771 a_n2472_13878.n24 a_n2472_13878.n22 0.358259
R22772 a_n2472_13878.n22 a_n2472_13878.n20 0.358259
R22773 a_n2472_13878.n20 a_n2472_13878.n18 0.358259
R22774 a_n2472_13878.n4 a_n2472_13878.n2 0.146627
R22775 a_n2472_13878.n6 a_n2472_13878.n4 0.146627
R22776 a_n2472_13878.n8 a_n2472_13878.n6 0.146627
R22777 a_n2472_13878.n12 a_n2472_13878.n11 0.101793
R22778 a_n2650_8322.n10 a_n2650_8322.t3 74.6477
R22779 a_n2650_8322.n1 a_n2650_8322.t23 74.6477
R22780 a_n2650_8322.n24 a_n2650_8322.t25 74.6474
R22781 a_n2650_8322.n18 a_n2650_8322.t22 74.2899
R22782 a_n2650_8322.n11 a_n2650_8322.t1 74.2899
R22783 a_n2650_8322.n12 a_n2650_8322.t4 74.2899
R22784 a_n2650_8322.n15 a_n2650_8322.t5 74.2899
R22785 a_n2650_8322.n8 a_n2650_8322.t8 74.2899
R22786 a_n2650_8322.n24 a_n2650_8322.n23 70.6783
R22787 a_n2650_8322.n22 a_n2650_8322.n21 70.6783
R22788 a_n2650_8322.n20 a_n2650_8322.n19 70.6783
R22789 a_n2650_8322.n10 a_n2650_8322.n9 70.6783
R22790 a_n2650_8322.n14 a_n2650_8322.n13 70.6783
R22791 a_n2650_8322.n1 a_n2650_8322.n0 70.6783
R22792 a_n2650_8322.n3 a_n2650_8322.n2 70.6783
R22793 a_n2650_8322.n5 a_n2650_8322.n4 70.6783
R22794 a_n2650_8322.n7 a_n2650_8322.n6 70.6783
R22795 a_n2650_8322.n26 a_n2650_8322.n25 70.6782
R22796 a_n2650_8322.n16 a_n2650_8322.n8 24.1867
R22797 a_n2650_8322.n17 a_n2650_8322.t29 9.75584
R22798 a_n2650_8322.n16 a_n2650_8322.n15 7.67184
R22799 a_n2650_8322.n18 a_n2650_8322.n17 6.55222
R22800 a_n2650_8322.n17 a_n2650_8322.n16 5.3452
R22801 a_n2650_8322.n23 a_n2650_8322.t20 3.61217
R22802 a_n2650_8322.n23 a_n2650_8322.t16 3.61217
R22803 a_n2650_8322.n21 a_n2650_8322.t24 3.61217
R22804 a_n2650_8322.n21 a_n2650_8322.t14 3.61217
R22805 a_n2650_8322.n19 a_n2650_8322.t12 3.61217
R22806 a_n2650_8322.n19 a_n2650_8322.t11 3.61217
R22807 a_n2650_8322.n9 a_n2650_8322.t7 3.61217
R22808 a_n2650_8322.n9 a_n2650_8322.t6 3.61217
R22809 a_n2650_8322.n13 a_n2650_8322.t2 3.61217
R22810 a_n2650_8322.n13 a_n2650_8322.t0 3.61217
R22811 a_n2650_8322.n0 a_n2650_8322.t26 3.61217
R22812 a_n2650_8322.n0 a_n2650_8322.t18 3.61217
R22813 a_n2650_8322.n2 a_n2650_8322.t10 3.61217
R22814 a_n2650_8322.n2 a_n2650_8322.t9 3.61217
R22815 a_n2650_8322.n4 a_n2650_8322.t21 3.61217
R22816 a_n2650_8322.n4 a_n2650_8322.t15 3.61217
R22817 a_n2650_8322.n6 a_n2650_8322.t19 3.61217
R22818 a_n2650_8322.n6 a_n2650_8322.t17 3.61217
R22819 a_n2650_8322.n26 a_n2650_8322.t13 3.61217
R22820 a_n2650_8322.t27 a_n2650_8322.n26 3.61217
R22821 a_n2650_8322.n15 a_n2650_8322.n14 0.358259
R22822 a_n2650_8322.n14 a_n2650_8322.n12 0.358259
R22823 a_n2650_8322.n11 a_n2650_8322.n10 0.358259
R22824 a_n2650_8322.n8 a_n2650_8322.n7 0.358259
R22825 a_n2650_8322.n7 a_n2650_8322.n5 0.358259
R22826 a_n2650_8322.n5 a_n2650_8322.n3 0.358259
R22827 a_n2650_8322.n3 a_n2650_8322.n1 0.358259
R22828 a_n2650_8322.n20 a_n2650_8322.n18 0.358259
R22829 a_n2650_8322.n22 a_n2650_8322.n20 0.358259
R22830 a_n2650_8322.n25 a_n2650_8322.n22 0.358259
R22831 a_n2650_8322.n25 a_n2650_8322.n24 0.358259
R22832 a_n2650_8322.n12 a_n2650_8322.n11 0.101793
R22833 a_n2650_8322.t32 a_n2650_8322.t30 0.0788333
R22834 a_n2650_8322.t28 a_n2650_8322.t33 0.0788333
R22835 a_n2650_8322.t29 a_n2650_8322.t31 0.0788333
R22836 a_n2650_8322.t28 a_n2650_8322.t32 0.0318333
R22837 a_n2650_8322.t29 a_n2650_8322.t33 0.0318333
R22838 a_n2650_8322.t30 a_n2650_8322.t33 0.0318333
R22839 a_n2650_8322.t31 a_n2650_8322.t28 0.0318333
R22840 output.n41 output.n15 289.615
R22841 output.n72 output.n46 289.615
R22842 output.n104 output.n78 289.615
R22843 output.n136 output.n110 289.615
R22844 output.n77 output.n45 197.26
R22845 output.n77 output.n76 196.298
R22846 output.n109 output.n108 196.298
R22847 output.n141 output.n140 196.298
R22848 output.n42 output.n41 185
R22849 output.n40 output.n39 185
R22850 output.n19 output.n18 185
R22851 output.n34 output.n33 185
R22852 output.n32 output.n31 185
R22853 output.n23 output.n22 185
R22854 output.n26 output.n25 185
R22855 output.n73 output.n72 185
R22856 output.n71 output.n70 185
R22857 output.n50 output.n49 185
R22858 output.n65 output.n64 185
R22859 output.n63 output.n62 185
R22860 output.n54 output.n53 185
R22861 output.n57 output.n56 185
R22862 output.n105 output.n104 185
R22863 output.n103 output.n102 185
R22864 output.n82 output.n81 185
R22865 output.n97 output.n96 185
R22866 output.n95 output.n94 185
R22867 output.n86 output.n85 185
R22868 output.n89 output.n88 185
R22869 output.n137 output.n136 185
R22870 output.n135 output.n134 185
R22871 output.n114 output.n113 185
R22872 output.n129 output.n128 185
R22873 output.n127 output.n126 185
R22874 output.n118 output.n117 185
R22875 output.n121 output.n120 185
R22876 output.t0 output.n24 147.661
R22877 output.t18 output.n55 147.661
R22878 output.t1 output.n87 147.661
R22879 output.t19 output.n119 147.661
R22880 output.n41 output.n40 104.615
R22881 output.n40 output.n18 104.615
R22882 output.n33 output.n18 104.615
R22883 output.n33 output.n32 104.615
R22884 output.n32 output.n22 104.615
R22885 output.n25 output.n22 104.615
R22886 output.n72 output.n71 104.615
R22887 output.n71 output.n49 104.615
R22888 output.n64 output.n49 104.615
R22889 output.n64 output.n63 104.615
R22890 output.n63 output.n53 104.615
R22891 output.n56 output.n53 104.615
R22892 output.n104 output.n103 104.615
R22893 output.n103 output.n81 104.615
R22894 output.n96 output.n81 104.615
R22895 output.n96 output.n95 104.615
R22896 output.n95 output.n85 104.615
R22897 output.n88 output.n85 104.615
R22898 output.n136 output.n135 104.615
R22899 output.n135 output.n113 104.615
R22900 output.n128 output.n113 104.615
R22901 output.n128 output.n127 104.615
R22902 output.n127 output.n117 104.615
R22903 output.n120 output.n117 104.615
R22904 output.n1 output.t13 77.056
R22905 output.n14 output.t15 76.6694
R22906 output.n1 output.n0 72.7095
R22907 output.n3 output.n2 72.7095
R22908 output.n5 output.n4 72.7095
R22909 output.n7 output.n6 72.7095
R22910 output.n9 output.n8 72.7095
R22911 output.n11 output.n10 72.7095
R22912 output.n13 output.n12 72.7095
R22913 output.n25 output.t0 52.3082
R22914 output.n56 output.t18 52.3082
R22915 output.n88 output.t1 52.3082
R22916 output.n120 output.t19 52.3082
R22917 output.n26 output.n24 15.6674
R22918 output.n57 output.n55 15.6674
R22919 output.n89 output.n87 15.6674
R22920 output.n121 output.n119 15.6674
R22921 output.n27 output.n23 12.8005
R22922 output.n58 output.n54 12.8005
R22923 output.n90 output.n86 12.8005
R22924 output.n122 output.n118 12.8005
R22925 output.n31 output.n30 12.0247
R22926 output.n62 output.n61 12.0247
R22927 output.n94 output.n93 12.0247
R22928 output.n126 output.n125 12.0247
R22929 output.n34 output.n21 11.249
R22930 output.n65 output.n52 11.249
R22931 output.n97 output.n84 11.249
R22932 output.n129 output.n116 11.249
R22933 output.n35 output.n19 10.4732
R22934 output.n66 output.n50 10.4732
R22935 output.n98 output.n82 10.4732
R22936 output.n130 output.n114 10.4732
R22937 output.n39 output.n38 9.69747
R22938 output.n70 output.n69 9.69747
R22939 output.n102 output.n101 9.69747
R22940 output.n134 output.n133 9.69747
R22941 output.n45 output.n44 9.45567
R22942 output.n76 output.n75 9.45567
R22943 output.n108 output.n107 9.45567
R22944 output.n140 output.n139 9.45567
R22945 output.n44 output.n43 9.3005
R22946 output.n17 output.n16 9.3005
R22947 output.n38 output.n37 9.3005
R22948 output.n36 output.n35 9.3005
R22949 output.n21 output.n20 9.3005
R22950 output.n30 output.n29 9.3005
R22951 output.n28 output.n27 9.3005
R22952 output.n75 output.n74 9.3005
R22953 output.n48 output.n47 9.3005
R22954 output.n69 output.n68 9.3005
R22955 output.n67 output.n66 9.3005
R22956 output.n52 output.n51 9.3005
R22957 output.n61 output.n60 9.3005
R22958 output.n59 output.n58 9.3005
R22959 output.n107 output.n106 9.3005
R22960 output.n80 output.n79 9.3005
R22961 output.n101 output.n100 9.3005
R22962 output.n99 output.n98 9.3005
R22963 output.n84 output.n83 9.3005
R22964 output.n93 output.n92 9.3005
R22965 output.n91 output.n90 9.3005
R22966 output.n139 output.n138 9.3005
R22967 output.n112 output.n111 9.3005
R22968 output.n133 output.n132 9.3005
R22969 output.n131 output.n130 9.3005
R22970 output.n116 output.n115 9.3005
R22971 output.n125 output.n124 9.3005
R22972 output.n123 output.n122 9.3005
R22973 output.n42 output.n17 8.92171
R22974 output.n73 output.n48 8.92171
R22975 output.n105 output.n80 8.92171
R22976 output.n137 output.n112 8.92171
R22977 output output.n141 8.15037
R22978 output.n43 output.n15 8.14595
R22979 output.n74 output.n46 8.14595
R22980 output.n106 output.n78 8.14595
R22981 output.n138 output.n110 8.14595
R22982 output.n45 output.n15 5.81868
R22983 output.n76 output.n46 5.81868
R22984 output.n108 output.n78 5.81868
R22985 output.n140 output.n110 5.81868
R22986 output.n43 output.n42 5.04292
R22987 output.n74 output.n73 5.04292
R22988 output.n106 output.n105 5.04292
R22989 output.n138 output.n137 5.04292
R22990 output.n28 output.n24 4.38594
R22991 output.n59 output.n55 4.38594
R22992 output.n91 output.n87 4.38594
R22993 output.n123 output.n119 4.38594
R22994 output.n39 output.n17 4.26717
R22995 output.n70 output.n48 4.26717
R22996 output.n102 output.n80 4.26717
R22997 output.n134 output.n112 4.26717
R22998 output.n0 output.t3 3.9605
R22999 output.n0 output.t8 3.9605
R23000 output.n2 output.t12 3.9605
R23001 output.n2 output.t4 3.9605
R23002 output.n4 output.t6 3.9605
R23003 output.n4 output.t5 3.9605
R23004 output.n6 output.t11 3.9605
R23005 output.n6 output.t14 3.9605
R23006 output.n8 output.t16 3.9605
R23007 output.n8 output.t9 3.9605
R23008 output.n10 output.t10 3.9605
R23009 output.n10 output.t17 3.9605
R23010 output.n12 output.t2 3.9605
R23011 output.n12 output.t7 3.9605
R23012 output.n38 output.n19 3.49141
R23013 output.n69 output.n50 3.49141
R23014 output.n101 output.n82 3.49141
R23015 output.n133 output.n114 3.49141
R23016 output.n35 output.n34 2.71565
R23017 output.n66 output.n65 2.71565
R23018 output.n98 output.n97 2.71565
R23019 output.n130 output.n129 2.71565
R23020 output.n31 output.n21 1.93989
R23021 output.n62 output.n52 1.93989
R23022 output.n94 output.n84 1.93989
R23023 output.n126 output.n116 1.93989
R23024 output.n30 output.n23 1.16414
R23025 output.n61 output.n54 1.16414
R23026 output.n93 output.n86 1.16414
R23027 output.n125 output.n118 1.16414
R23028 output.n141 output.n109 0.962709
R23029 output.n109 output.n77 0.962709
R23030 output.n27 output.n26 0.388379
R23031 output.n58 output.n57 0.388379
R23032 output.n90 output.n89 0.388379
R23033 output.n122 output.n121 0.388379
R23034 output.n14 output.n13 0.387128
R23035 output.n13 output.n11 0.387128
R23036 output.n11 output.n9 0.387128
R23037 output.n9 output.n7 0.387128
R23038 output.n7 output.n5 0.387128
R23039 output.n5 output.n3 0.387128
R23040 output.n3 output.n1 0.387128
R23041 output.n44 output.n16 0.155672
R23042 output.n37 output.n16 0.155672
R23043 output.n37 output.n36 0.155672
R23044 output.n36 output.n20 0.155672
R23045 output.n29 output.n20 0.155672
R23046 output.n29 output.n28 0.155672
R23047 output.n75 output.n47 0.155672
R23048 output.n68 output.n47 0.155672
R23049 output.n68 output.n67 0.155672
R23050 output.n67 output.n51 0.155672
R23051 output.n60 output.n51 0.155672
R23052 output.n60 output.n59 0.155672
R23053 output.n107 output.n79 0.155672
R23054 output.n100 output.n79 0.155672
R23055 output.n100 output.n99 0.155672
R23056 output.n99 output.n83 0.155672
R23057 output.n92 output.n83 0.155672
R23058 output.n92 output.n91 0.155672
R23059 output.n139 output.n111 0.155672
R23060 output.n132 output.n111 0.155672
R23061 output.n132 output.n131 0.155672
R23062 output.n131 output.n115 0.155672
R23063 output.n124 output.n115 0.155672
R23064 output.n124 output.n123 0.155672
R23065 output output.n14 0.126227
R23066 plus.n43 plus.t25 442.325
R23067 plus.n11 plus.t12 442.325
R23068 plus.n42 plus.t5 415.966
R23069 plus.n41 plus.t20 415.966
R23070 plus.n47 plus.t26 415.966
R23071 plus.n39 plus.t11 415.966
R23072 plus.n52 plus.t6 415.966
R23073 plus.n54 plus.t10 415.966
R23074 plus.n37 plus.t19 415.966
R23075 plus.n59 plus.t8 415.966
R23076 plus.n35 plus.t16 415.966
R23077 plus.n64 plus.t28 415.966
R23078 plus.n66 plus.t21 415.966
R23079 plus.n32 plus.t23 415.966
R23080 plus.n30 plus.t13 415.966
R23081 plus.n29 plus.t27 415.966
R23082 plus.n3 plus.t22 415.966
R23083 plus.n23 plus.t7 415.966
R23084 plus.n22 plus.t18 415.966
R23085 plus.n6 plus.t14 415.966
R23086 plus.n17 plus.t24 415.966
R23087 plus.n15 plus.t17 415.966
R23088 plus.n9 plus.t9 415.966
R23089 plus.n10 plus.t15 415.966
R23090 plus.n70 plus.t3 243.97
R23091 plus.n70 plus.n69 223.454
R23092 plus.n72 plus.n71 223.454
R23093 plus.n67 plus.n66 161.3
R23094 plus.n65 plus.n34 161.3
R23095 plus.n64 plus.n63 161.3
R23096 plus.n62 plus.n35 161.3
R23097 plus.n61 plus.n60 161.3
R23098 plus.n59 plus.n36 161.3
R23099 plus.n58 plus.n57 161.3
R23100 plus.n56 plus.n37 161.3
R23101 plus.n55 plus.n54 161.3
R23102 plus.n53 plus.n38 161.3
R23103 plus.n52 plus.n51 161.3
R23104 plus.n50 plus.n39 161.3
R23105 plus.n49 plus.n48 161.3
R23106 plus.n47 plus.n40 161.3
R23107 plus.n46 plus.n45 161.3
R23108 plus.n44 plus.n41 161.3
R23109 plus.n12 plus.n9 161.3
R23110 plus.n14 plus.n13 161.3
R23111 plus.n15 plus.n8 161.3
R23112 plus.n16 plus.n7 161.3
R23113 plus.n18 plus.n17 161.3
R23114 plus.n19 plus.n6 161.3
R23115 plus.n21 plus.n20 161.3
R23116 plus.n22 plus.n5 161.3
R23117 plus.n23 plus.n4 161.3
R23118 plus.n25 plus.n24 161.3
R23119 plus.n26 plus.n3 161.3
R23120 plus.n28 plus.n27 161.3
R23121 plus.n29 plus.n2 161.3
R23122 plus.n30 plus.n1 161.3
R23123 plus.n31 plus.n0 161.3
R23124 plus.n33 plus.n32 161.3
R23125 plus.n42 plus.n41 48.2005
R23126 plus.n52 plus.n39 48.2005
R23127 plus.n54 plus.n37 48.2005
R23128 plus.n64 plus.n35 48.2005
R23129 plus.n30 plus.n29 48.2005
R23130 plus.n23 plus.n22 48.2005
R23131 plus.n17 plus.n6 48.2005
R23132 plus.n10 plus.n9 48.2005
R23133 plus.n48 plus.n47 47.4702
R23134 plus.n59 plus.n58 47.4702
R23135 plus.n24 plus.n3 47.4702
R23136 plus.n16 plus.n15 47.4702
R23137 plus.n66 plus.n65 46.0096
R23138 plus.n32 plus.n31 46.0096
R23139 plus.n44 plus.n43 45.0871
R23140 plus.n12 plus.n11 45.0871
R23141 plus.n68 plus.n67 31.0554
R23142 plus.n47 plus.n46 25.5611
R23143 plus.n60 plus.n59 25.5611
R23144 plus.n28 plus.n3 25.5611
R23145 plus.n15 plus.n14 25.5611
R23146 plus.n53 plus.n52 24.1005
R23147 plus.n54 plus.n53 24.1005
R23148 plus.n22 plus.n21 24.1005
R23149 plus.n21 plus.n6 24.1005
R23150 plus.n46 plus.n41 22.6399
R23151 plus.n60 plus.n35 22.6399
R23152 plus.n29 plus.n28 22.6399
R23153 plus.n14 plus.n9 22.6399
R23154 plus.n69 plus.t4 19.8005
R23155 plus.n69 plus.t1 19.8005
R23156 plus.n71 plus.t0 19.8005
R23157 plus.n71 plus.t2 19.8005
R23158 plus plus.n73 14.4109
R23159 plus.n43 plus.n42 14.1472
R23160 plus.n11 plus.n10 14.1472
R23161 plus.n68 plus.n33 11.7259
R23162 plus.n73 plus.n72 5.40567
R23163 plus.n65 plus.n64 2.19141
R23164 plus.n31 plus.n30 2.19141
R23165 plus.n73 plus.n68 1.188
R23166 plus.n48 plus.n39 0.730803
R23167 plus.n58 plus.n37 0.730803
R23168 plus.n24 plus.n23 0.730803
R23169 plus.n17 plus.n16 0.730803
R23170 plus.n72 plus.n70 0.716017
R23171 plus.n45 plus.n44 0.189894
R23172 plus.n45 plus.n40 0.189894
R23173 plus.n49 plus.n40 0.189894
R23174 plus.n50 plus.n49 0.189894
R23175 plus.n51 plus.n50 0.189894
R23176 plus.n51 plus.n38 0.189894
R23177 plus.n55 plus.n38 0.189894
R23178 plus.n56 plus.n55 0.189894
R23179 plus.n57 plus.n56 0.189894
R23180 plus.n57 plus.n36 0.189894
R23181 plus.n61 plus.n36 0.189894
R23182 plus.n62 plus.n61 0.189894
R23183 plus.n63 plus.n62 0.189894
R23184 plus.n63 plus.n34 0.189894
R23185 plus.n67 plus.n34 0.189894
R23186 plus.n33 plus.n0 0.189894
R23187 plus.n1 plus.n0 0.189894
R23188 plus.n2 plus.n1 0.189894
R23189 plus.n27 plus.n2 0.189894
R23190 plus.n27 plus.n26 0.189894
R23191 plus.n26 plus.n25 0.189894
R23192 plus.n25 plus.n4 0.189894
R23193 plus.n5 plus.n4 0.189894
R23194 plus.n20 plus.n5 0.189894
R23195 plus.n20 plus.n19 0.189894
R23196 plus.n19 plus.n18 0.189894
R23197 plus.n18 plus.n7 0.189894
R23198 plus.n8 plus.n7 0.189894
R23199 plus.n13 plus.n8 0.189894
R23200 plus.n13 plus.n12 0.189894
R23201 a_n2903_n3924.n14 a_n2903_n3924.t49 214.994
R23202 a_n2903_n3924.n1 a_n2903_n3924.t34 214.493
R23203 a_n2903_n3924.n15 a_n2903_n3924.t46 214.321
R23204 a_n2903_n3924.n16 a_n2903_n3924.t44 214.321
R23205 a_n2903_n3924.n17 a_n2903_n3924.t48 214.321
R23206 a_n2903_n3924.n18 a_n2903_n3924.t45 214.321
R23207 a_n2903_n3924.n19 a_n2903_n3924.t4 214.321
R23208 a_n2903_n3924.n14 a_n2903_n3924.t9 214.321
R23209 a_n2903_n3924.n0 a_n2903_n3924.t13 55.8337
R23210 a_n2903_n3924.n2 a_n2903_n3924.t51 55.8337
R23211 a_n2903_n3924.n13 a_n2903_n3924.t2 55.8337
R23212 a_n2903_n3924.n47 a_n2903_n3924.t17 55.8335
R23213 a_n2903_n3924.n45 a_n2903_n3924.t35 55.8335
R23214 a_n2903_n3924.n34 a_n2903_n3924.t0 55.8335
R23215 a_n2903_n3924.n33 a_n2903_n3924.t26 55.8335
R23216 a_n2903_n3924.n22 a_n2903_n3924.t15 55.8335
R23217 a_n2903_n3924.n49 a_n2903_n3924.n48 53.0052
R23218 a_n2903_n3924.n51 a_n2903_n3924.n50 53.0052
R23219 a_n2903_n3924.n53 a_n2903_n3924.n52 53.0052
R23220 a_n2903_n3924.n55 a_n2903_n3924.n54 53.0052
R23221 a_n2903_n3924.n4 a_n2903_n3924.n3 53.0052
R23222 a_n2903_n3924.n6 a_n2903_n3924.n5 53.0052
R23223 a_n2903_n3924.n8 a_n2903_n3924.n7 53.0052
R23224 a_n2903_n3924.n10 a_n2903_n3924.n9 53.0052
R23225 a_n2903_n3924.n12 a_n2903_n3924.n11 53.0052
R23226 a_n2903_n3924.n44 a_n2903_n3924.n43 53.0051
R23227 a_n2903_n3924.n42 a_n2903_n3924.n41 53.0051
R23228 a_n2903_n3924.n40 a_n2903_n3924.n39 53.0051
R23229 a_n2903_n3924.n38 a_n2903_n3924.n37 53.0051
R23230 a_n2903_n3924.n36 a_n2903_n3924.n35 53.0051
R23231 a_n2903_n3924.n32 a_n2903_n3924.n31 53.0051
R23232 a_n2903_n3924.n30 a_n2903_n3924.n29 53.0051
R23233 a_n2903_n3924.n28 a_n2903_n3924.n27 53.0051
R23234 a_n2903_n3924.n26 a_n2903_n3924.n25 53.0051
R23235 a_n2903_n3924.n24 a_n2903_n3924.n23 53.0051
R23236 a_n2903_n3924.n57 a_n2903_n3924.n56 53.0051
R23237 a_n2903_n3924.n21 a_n2903_n3924.n13 12.1555
R23238 a_n2903_n3924.n47 a_n2903_n3924.n46 12.1555
R23239 a_n2903_n3924.n22 a_n2903_n3924.n21 5.07593
R23240 a_n2903_n3924.n46 a_n2903_n3924.n45 5.07593
R23241 a_n2903_n3924.n48 a_n2903_n3924.t22 2.82907
R23242 a_n2903_n3924.n48 a_n2903_n3924.t10 2.82907
R23243 a_n2903_n3924.n50 a_n2903_n3924.t19 2.82907
R23244 a_n2903_n3924.n50 a_n2903_n3924.t30 2.82907
R23245 a_n2903_n3924.n52 a_n2903_n3924.t32 2.82907
R23246 a_n2903_n3924.n52 a_n2903_n3924.t28 2.82907
R23247 a_n2903_n3924.n54 a_n2903_n3924.t12 2.82907
R23248 a_n2903_n3924.n54 a_n2903_n3924.t27 2.82907
R23249 a_n2903_n3924.n3 a_n2903_n3924.t39 2.82907
R23250 a_n2903_n3924.n3 a_n2903_n3924.t42 2.82907
R23251 a_n2903_n3924.n5 a_n2903_n3924.t5 2.82907
R23252 a_n2903_n3924.n5 a_n2903_n3924.t3 2.82907
R23253 a_n2903_n3924.n7 a_n2903_n3924.t41 2.82907
R23254 a_n2903_n3924.n7 a_n2903_n3924.t1 2.82907
R23255 a_n2903_n3924.n9 a_n2903_n3924.t55 2.82907
R23256 a_n2903_n3924.n9 a_n2903_n3924.t50 2.82907
R23257 a_n2903_n3924.n11 a_n2903_n3924.t7 2.82907
R23258 a_n2903_n3924.n11 a_n2903_n3924.t36 2.82907
R23259 a_n2903_n3924.n43 a_n2903_n3924.t53 2.82907
R23260 a_n2903_n3924.n43 a_n2903_n3924.t52 2.82907
R23261 a_n2903_n3924.n41 a_n2903_n3924.t47 2.82907
R23262 a_n2903_n3924.n41 a_n2903_n3924.t38 2.82907
R23263 a_n2903_n3924.n39 a_n2903_n3924.t8 2.82907
R23264 a_n2903_n3924.n39 a_n2903_n3924.t6 2.82907
R23265 a_n2903_n3924.n37 a_n2903_n3924.t40 2.82907
R23266 a_n2903_n3924.n37 a_n2903_n3924.t43 2.82907
R23267 a_n2903_n3924.n35 a_n2903_n3924.t54 2.82907
R23268 a_n2903_n3924.n35 a_n2903_n3924.t37 2.82907
R23269 a_n2903_n3924.n31 a_n2903_n3924.t29 2.82907
R23270 a_n2903_n3924.n31 a_n2903_n3924.t23 2.82907
R23271 a_n2903_n3924.n29 a_n2903_n3924.t14 2.82907
R23272 a_n2903_n3924.n29 a_n2903_n3924.t21 2.82907
R23273 a_n2903_n3924.n27 a_n2903_n3924.t20 2.82907
R23274 a_n2903_n3924.n27 a_n2903_n3924.t24 2.82907
R23275 a_n2903_n3924.n25 a_n2903_n3924.t16 2.82907
R23276 a_n2903_n3924.n25 a_n2903_n3924.t31 2.82907
R23277 a_n2903_n3924.n23 a_n2903_n3924.t25 2.82907
R23278 a_n2903_n3924.n23 a_n2903_n3924.t11 2.82907
R23279 a_n2903_n3924.t33 a_n2903_n3924.n57 2.82907
R23280 a_n2903_n3924.n57 a_n2903_n3924.t18 2.82907
R23281 a_n2903_n3924.n46 a_n2903_n3924.n1 1.95694
R23282 a_n2903_n3924.n21 a_n2903_n3924.n20 1.95694
R23283 a_n2903_n3924.n19 a_n2903_n3924.n18 0.672012
R23284 a_n2903_n3924.n18 a_n2903_n3924.n17 0.672012
R23285 a_n2903_n3924.n17 a_n2903_n3924.n16 0.672012
R23286 a_n2903_n3924.n16 a_n2903_n3924.n15 0.672012
R23287 a_n2903_n3924.n20 a_n2903_n3924.n19 0.643669
R23288 a_n2903_n3924.n15 a_n2903_n3924.n1 0.501227
R23289 a_n2903_n3924.n24 a_n2903_n3924.n22 0.358259
R23290 a_n2903_n3924.n26 a_n2903_n3924.n24 0.358259
R23291 a_n2903_n3924.n28 a_n2903_n3924.n26 0.358259
R23292 a_n2903_n3924.n30 a_n2903_n3924.n28 0.358259
R23293 a_n2903_n3924.n32 a_n2903_n3924.n30 0.358259
R23294 a_n2903_n3924.n33 a_n2903_n3924.n32 0.358259
R23295 a_n2903_n3924.n36 a_n2903_n3924.n34 0.358259
R23296 a_n2903_n3924.n38 a_n2903_n3924.n36 0.358259
R23297 a_n2903_n3924.n40 a_n2903_n3924.n38 0.358259
R23298 a_n2903_n3924.n42 a_n2903_n3924.n40 0.358259
R23299 a_n2903_n3924.n44 a_n2903_n3924.n42 0.358259
R23300 a_n2903_n3924.n45 a_n2903_n3924.n44 0.358259
R23301 a_n2903_n3924.n13 a_n2903_n3924.n12 0.358259
R23302 a_n2903_n3924.n12 a_n2903_n3924.n10 0.358259
R23303 a_n2903_n3924.n10 a_n2903_n3924.n8 0.358259
R23304 a_n2903_n3924.n8 a_n2903_n3924.n6 0.358259
R23305 a_n2903_n3924.n6 a_n2903_n3924.n4 0.358259
R23306 a_n2903_n3924.n4 a_n2903_n3924.n2 0.358259
R23307 a_n2903_n3924.n56 a_n2903_n3924.n0 0.358259
R23308 a_n2903_n3924.n56 a_n2903_n3924.n55 0.358259
R23309 a_n2903_n3924.n55 a_n2903_n3924.n53 0.358259
R23310 a_n2903_n3924.n53 a_n2903_n3924.n51 0.358259
R23311 a_n2903_n3924.n51 a_n2903_n3924.n49 0.358259
R23312 a_n2903_n3924.n49 a_n2903_n3924.n47 0.358259
R23313 a_n2903_n3924.n34 a_n2903_n3924.n33 0.235414
R23314 a_n2903_n3924.n2 a_n2903_n3924.n0 0.235414
R23315 a_n2903_n3924.n20 a_n2903_n3924.n14 0.028843
R23316 minus.n45 minus.t26 442.325
R23317 minus.n9 minus.t12 442.325
R23318 minus.n66 minus.t16 415.966
R23319 minus.n64 minus.t28 415.966
R23320 minus.n63 minus.t21 415.966
R23321 minus.n37 minus.t14 415.966
R23322 minus.n57 minus.t23 415.966
R23323 minus.n56 minus.t11 415.966
R23324 minus.n40 minus.t5 415.966
R23325 minus.n51 minus.t17 415.966
R23326 minus.n49 minus.t10 415.966
R23327 minus.n43 minus.t25 415.966
R23328 minus.n44 minus.t7 415.966
R23329 minus.n8 minus.t18 415.966
R23330 minus.n7 minus.t8 415.966
R23331 minus.n13 minus.t13 415.966
R23332 minus.n5 minus.t24 415.966
R23333 minus.n18 minus.t19 415.966
R23334 minus.n20 minus.t22 415.966
R23335 minus.n3 minus.t6 415.966
R23336 minus.n25 minus.t20 415.966
R23337 minus.n1 minus.t27 415.966
R23338 minus.n30 minus.t15 415.966
R23339 minus.n32 minus.t9 415.966
R23340 minus.n72 minus.t3 243.255
R23341 minus.n71 minus.n69 224.169
R23342 minus.n71 minus.n70 223.454
R23343 minus.n46 minus.n43 161.3
R23344 minus.n48 minus.n47 161.3
R23345 minus.n49 minus.n42 161.3
R23346 minus.n50 minus.n41 161.3
R23347 minus.n52 minus.n51 161.3
R23348 minus.n53 minus.n40 161.3
R23349 minus.n55 minus.n54 161.3
R23350 minus.n56 minus.n39 161.3
R23351 minus.n57 minus.n38 161.3
R23352 minus.n59 minus.n58 161.3
R23353 minus.n60 minus.n37 161.3
R23354 minus.n62 minus.n61 161.3
R23355 minus.n63 minus.n36 161.3
R23356 minus.n64 minus.n35 161.3
R23357 minus.n65 minus.n34 161.3
R23358 minus.n67 minus.n66 161.3
R23359 minus.n33 minus.n32 161.3
R23360 minus.n31 minus.n0 161.3
R23361 minus.n30 minus.n29 161.3
R23362 minus.n28 minus.n1 161.3
R23363 minus.n27 minus.n26 161.3
R23364 minus.n25 minus.n2 161.3
R23365 minus.n24 minus.n23 161.3
R23366 minus.n22 minus.n3 161.3
R23367 minus.n21 minus.n20 161.3
R23368 minus.n19 minus.n4 161.3
R23369 minus.n18 minus.n17 161.3
R23370 minus.n16 minus.n5 161.3
R23371 minus.n15 minus.n14 161.3
R23372 minus.n13 minus.n6 161.3
R23373 minus.n12 minus.n11 161.3
R23374 minus.n10 minus.n7 161.3
R23375 minus.n64 minus.n63 48.2005
R23376 minus.n57 minus.n56 48.2005
R23377 minus.n51 minus.n40 48.2005
R23378 minus.n44 minus.n43 48.2005
R23379 minus.n8 minus.n7 48.2005
R23380 minus.n18 minus.n5 48.2005
R23381 minus.n20 minus.n3 48.2005
R23382 minus.n30 minus.n1 48.2005
R23383 minus.n58 minus.n37 47.4702
R23384 minus.n50 minus.n49 47.4702
R23385 minus.n14 minus.n13 47.4702
R23386 minus.n25 minus.n24 47.4702
R23387 minus.n66 minus.n65 46.0096
R23388 minus.n32 minus.n31 46.0096
R23389 minus.n10 minus.n9 45.0871
R23390 minus.n46 minus.n45 45.0871
R23391 minus.n68 minus.n67 31.2713
R23392 minus.n62 minus.n37 25.5611
R23393 minus.n49 minus.n48 25.5611
R23394 minus.n13 minus.n12 25.5611
R23395 minus.n26 minus.n25 25.5611
R23396 minus.n56 minus.n55 24.1005
R23397 minus.n55 minus.n40 24.1005
R23398 minus.n19 minus.n18 24.1005
R23399 minus.n20 minus.n19 24.1005
R23400 minus.n63 minus.n62 22.6399
R23401 minus.n48 minus.n43 22.6399
R23402 minus.n12 minus.n7 22.6399
R23403 minus.n26 minus.n1 22.6399
R23404 minus.n70 minus.t2 19.8005
R23405 minus.n70 minus.t0 19.8005
R23406 minus.n69 minus.t1 19.8005
R23407 minus.n69 minus.t4 19.8005
R23408 minus.n45 minus.n44 14.1472
R23409 minus.n9 minus.n8 14.1472
R23410 minus.n68 minus.n33 11.9418
R23411 minus minus.n73 11.5737
R23412 minus.n73 minus.n72 4.80222
R23413 minus.n65 minus.n64 2.19141
R23414 minus.n31 minus.n30 2.19141
R23415 minus.n73 minus.n68 0.972091
R23416 minus.n58 minus.n57 0.730803
R23417 minus.n51 minus.n50 0.730803
R23418 minus.n14 minus.n5 0.730803
R23419 minus.n24 minus.n3 0.730803
R23420 minus.n72 minus.n71 0.716017
R23421 minus.n67 minus.n34 0.189894
R23422 minus.n35 minus.n34 0.189894
R23423 minus.n36 minus.n35 0.189894
R23424 minus.n61 minus.n36 0.189894
R23425 minus.n61 minus.n60 0.189894
R23426 minus.n60 minus.n59 0.189894
R23427 minus.n59 minus.n38 0.189894
R23428 minus.n39 minus.n38 0.189894
R23429 minus.n54 minus.n39 0.189894
R23430 minus.n54 minus.n53 0.189894
R23431 minus.n53 minus.n52 0.189894
R23432 minus.n52 minus.n41 0.189894
R23433 minus.n42 minus.n41 0.189894
R23434 minus.n47 minus.n42 0.189894
R23435 minus.n47 minus.n46 0.189894
R23436 minus.n11 minus.n10 0.189894
R23437 minus.n11 minus.n6 0.189894
R23438 minus.n15 minus.n6 0.189894
R23439 minus.n16 minus.n15 0.189894
R23440 minus.n17 minus.n16 0.189894
R23441 minus.n17 minus.n4 0.189894
R23442 minus.n21 minus.n4 0.189894
R23443 minus.n22 minus.n21 0.189894
R23444 minus.n23 minus.n22 0.189894
R23445 minus.n23 minus.n2 0.189894
R23446 minus.n27 minus.n2 0.189894
R23447 minus.n28 minus.n27 0.189894
R23448 minus.n29 minus.n28 0.189894
R23449 minus.n29 minus.n0 0.189894
R23450 minus.n33 minus.n0 0.189894
R23451 outputibias.n27 outputibias.n1 289.615
R23452 outputibias.n58 outputibias.n32 289.615
R23453 outputibias.n90 outputibias.n64 289.615
R23454 outputibias.n122 outputibias.n96 289.615
R23455 outputibias.n28 outputibias.n27 185
R23456 outputibias.n26 outputibias.n25 185
R23457 outputibias.n5 outputibias.n4 185
R23458 outputibias.n20 outputibias.n19 185
R23459 outputibias.n18 outputibias.n17 185
R23460 outputibias.n9 outputibias.n8 185
R23461 outputibias.n12 outputibias.n11 185
R23462 outputibias.n59 outputibias.n58 185
R23463 outputibias.n57 outputibias.n56 185
R23464 outputibias.n36 outputibias.n35 185
R23465 outputibias.n51 outputibias.n50 185
R23466 outputibias.n49 outputibias.n48 185
R23467 outputibias.n40 outputibias.n39 185
R23468 outputibias.n43 outputibias.n42 185
R23469 outputibias.n91 outputibias.n90 185
R23470 outputibias.n89 outputibias.n88 185
R23471 outputibias.n68 outputibias.n67 185
R23472 outputibias.n83 outputibias.n82 185
R23473 outputibias.n81 outputibias.n80 185
R23474 outputibias.n72 outputibias.n71 185
R23475 outputibias.n75 outputibias.n74 185
R23476 outputibias.n123 outputibias.n122 185
R23477 outputibias.n121 outputibias.n120 185
R23478 outputibias.n100 outputibias.n99 185
R23479 outputibias.n115 outputibias.n114 185
R23480 outputibias.n113 outputibias.n112 185
R23481 outputibias.n104 outputibias.n103 185
R23482 outputibias.n107 outputibias.n106 185
R23483 outputibias.n0 outputibias.t8 178.945
R23484 outputibias.n133 outputibias.t9 177.018
R23485 outputibias.n132 outputibias.t10 177.018
R23486 outputibias.n0 outputibias.t11 177.018
R23487 outputibias.t7 outputibias.n10 147.661
R23488 outputibias.t5 outputibias.n41 147.661
R23489 outputibias.t1 outputibias.n73 147.661
R23490 outputibias.t3 outputibias.n105 147.661
R23491 outputibias.n128 outputibias.t6 132.363
R23492 outputibias.n128 outputibias.t4 130.436
R23493 outputibias.n129 outputibias.t0 130.436
R23494 outputibias.n130 outputibias.t2 130.436
R23495 outputibias.n27 outputibias.n26 104.615
R23496 outputibias.n26 outputibias.n4 104.615
R23497 outputibias.n19 outputibias.n4 104.615
R23498 outputibias.n19 outputibias.n18 104.615
R23499 outputibias.n18 outputibias.n8 104.615
R23500 outputibias.n11 outputibias.n8 104.615
R23501 outputibias.n58 outputibias.n57 104.615
R23502 outputibias.n57 outputibias.n35 104.615
R23503 outputibias.n50 outputibias.n35 104.615
R23504 outputibias.n50 outputibias.n49 104.615
R23505 outputibias.n49 outputibias.n39 104.615
R23506 outputibias.n42 outputibias.n39 104.615
R23507 outputibias.n90 outputibias.n89 104.615
R23508 outputibias.n89 outputibias.n67 104.615
R23509 outputibias.n82 outputibias.n67 104.615
R23510 outputibias.n82 outputibias.n81 104.615
R23511 outputibias.n81 outputibias.n71 104.615
R23512 outputibias.n74 outputibias.n71 104.615
R23513 outputibias.n122 outputibias.n121 104.615
R23514 outputibias.n121 outputibias.n99 104.615
R23515 outputibias.n114 outputibias.n99 104.615
R23516 outputibias.n114 outputibias.n113 104.615
R23517 outputibias.n113 outputibias.n103 104.615
R23518 outputibias.n106 outputibias.n103 104.615
R23519 outputibias.n63 outputibias.n31 95.6354
R23520 outputibias.n63 outputibias.n62 94.6732
R23521 outputibias.n95 outputibias.n94 94.6732
R23522 outputibias.n127 outputibias.n126 94.6732
R23523 outputibias.n11 outputibias.t7 52.3082
R23524 outputibias.n42 outputibias.t5 52.3082
R23525 outputibias.n74 outputibias.t1 52.3082
R23526 outputibias.n106 outputibias.t3 52.3082
R23527 outputibias.n12 outputibias.n10 15.6674
R23528 outputibias.n43 outputibias.n41 15.6674
R23529 outputibias.n75 outputibias.n73 15.6674
R23530 outputibias.n107 outputibias.n105 15.6674
R23531 outputibias.n13 outputibias.n9 12.8005
R23532 outputibias.n44 outputibias.n40 12.8005
R23533 outputibias.n76 outputibias.n72 12.8005
R23534 outputibias.n108 outputibias.n104 12.8005
R23535 outputibias.n17 outputibias.n16 12.0247
R23536 outputibias.n48 outputibias.n47 12.0247
R23537 outputibias.n80 outputibias.n79 12.0247
R23538 outputibias.n112 outputibias.n111 12.0247
R23539 outputibias.n20 outputibias.n7 11.249
R23540 outputibias.n51 outputibias.n38 11.249
R23541 outputibias.n83 outputibias.n70 11.249
R23542 outputibias.n115 outputibias.n102 11.249
R23543 outputibias.n21 outputibias.n5 10.4732
R23544 outputibias.n52 outputibias.n36 10.4732
R23545 outputibias.n84 outputibias.n68 10.4732
R23546 outputibias.n116 outputibias.n100 10.4732
R23547 outputibias.n25 outputibias.n24 9.69747
R23548 outputibias.n56 outputibias.n55 9.69747
R23549 outputibias.n88 outputibias.n87 9.69747
R23550 outputibias.n120 outputibias.n119 9.69747
R23551 outputibias.n31 outputibias.n30 9.45567
R23552 outputibias.n62 outputibias.n61 9.45567
R23553 outputibias.n94 outputibias.n93 9.45567
R23554 outputibias.n126 outputibias.n125 9.45567
R23555 outputibias.n30 outputibias.n29 9.3005
R23556 outputibias.n3 outputibias.n2 9.3005
R23557 outputibias.n24 outputibias.n23 9.3005
R23558 outputibias.n22 outputibias.n21 9.3005
R23559 outputibias.n7 outputibias.n6 9.3005
R23560 outputibias.n16 outputibias.n15 9.3005
R23561 outputibias.n14 outputibias.n13 9.3005
R23562 outputibias.n61 outputibias.n60 9.3005
R23563 outputibias.n34 outputibias.n33 9.3005
R23564 outputibias.n55 outputibias.n54 9.3005
R23565 outputibias.n53 outputibias.n52 9.3005
R23566 outputibias.n38 outputibias.n37 9.3005
R23567 outputibias.n47 outputibias.n46 9.3005
R23568 outputibias.n45 outputibias.n44 9.3005
R23569 outputibias.n93 outputibias.n92 9.3005
R23570 outputibias.n66 outputibias.n65 9.3005
R23571 outputibias.n87 outputibias.n86 9.3005
R23572 outputibias.n85 outputibias.n84 9.3005
R23573 outputibias.n70 outputibias.n69 9.3005
R23574 outputibias.n79 outputibias.n78 9.3005
R23575 outputibias.n77 outputibias.n76 9.3005
R23576 outputibias.n125 outputibias.n124 9.3005
R23577 outputibias.n98 outputibias.n97 9.3005
R23578 outputibias.n119 outputibias.n118 9.3005
R23579 outputibias.n117 outputibias.n116 9.3005
R23580 outputibias.n102 outputibias.n101 9.3005
R23581 outputibias.n111 outputibias.n110 9.3005
R23582 outputibias.n109 outputibias.n108 9.3005
R23583 outputibias.n28 outputibias.n3 8.92171
R23584 outputibias.n59 outputibias.n34 8.92171
R23585 outputibias.n91 outputibias.n66 8.92171
R23586 outputibias.n123 outputibias.n98 8.92171
R23587 outputibias.n29 outputibias.n1 8.14595
R23588 outputibias.n60 outputibias.n32 8.14595
R23589 outputibias.n92 outputibias.n64 8.14595
R23590 outputibias.n124 outputibias.n96 8.14595
R23591 outputibias.n31 outputibias.n1 5.81868
R23592 outputibias.n62 outputibias.n32 5.81868
R23593 outputibias.n94 outputibias.n64 5.81868
R23594 outputibias.n126 outputibias.n96 5.81868
R23595 outputibias.n131 outputibias.n130 5.20947
R23596 outputibias.n29 outputibias.n28 5.04292
R23597 outputibias.n60 outputibias.n59 5.04292
R23598 outputibias.n92 outputibias.n91 5.04292
R23599 outputibias.n124 outputibias.n123 5.04292
R23600 outputibias.n131 outputibias.n127 4.42209
R23601 outputibias.n14 outputibias.n10 4.38594
R23602 outputibias.n45 outputibias.n41 4.38594
R23603 outputibias.n77 outputibias.n73 4.38594
R23604 outputibias.n109 outputibias.n105 4.38594
R23605 outputibias.n132 outputibias.n131 4.28454
R23606 outputibias.n25 outputibias.n3 4.26717
R23607 outputibias.n56 outputibias.n34 4.26717
R23608 outputibias.n88 outputibias.n66 4.26717
R23609 outputibias.n120 outputibias.n98 4.26717
R23610 outputibias.n24 outputibias.n5 3.49141
R23611 outputibias.n55 outputibias.n36 3.49141
R23612 outputibias.n87 outputibias.n68 3.49141
R23613 outputibias.n119 outputibias.n100 3.49141
R23614 outputibias.n21 outputibias.n20 2.71565
R23615 outputibias.n52 outputibias.n51 2.71565
R23616 outputibias.n84 outputibias.n83 2.71565
R23617 outputibias.n116 outputibias.n115 2.71565
R23618 outputibias.n17 outputibias.n7 1.93989
R23619 outputibias.n48 outputibias.n38 1.93989
R23620 outputibias.n80 outputibias.n70 1.93989
R23621 outputibias.n112 outputibias.n102 1.93989
R23622 outputibias.n130 outputibias.n129 1.9266
R23623 outputibias.n129 outputibias.n128 1.9266
R23624 outputibias.n133 outputibias.n132 1.92658
R23625 outputibias.n134 outputibias.n133 1.29913
R23626 outputibias.n16 outputibias.n9 1.16414
R23627 outputibias.n47 outputibias.n40 1.16414
R23628 outputibias.n79 outputibias.n72 1.16414
R23629 outputibias.n111 outputibias.n104 1.16414
R23630 outputibias.n127 outputibias.n95 0.962709
R23631 outputibias.n95 outputibias.n63 0.962709
R23632 outputibias.n13 outputibias.n12 0.388379
R23633 outputibias.n44 outputibias.n43 0.388379
R23634 outputibias.n76 outputibias.n75 0.388379
R23635 outputibias.n108 outputibias.n107 0.388379
R23636 outputibias.n134 outputibias.n0 0.337251
R23637 outputibias outputibias.n134 0.302375
R23638 outputibias.n30 outputibias.n2 0.155672
R23639 outputibias.n23 outputibias.n2 0.155672
R23640 outputibias.n23 outputibias.n22 0.155672
R23641 outputibias.n22 outputibias.n6 0.155672
R23642 outputibias.n15 outputibias.n6 0.155672
R23643 outputibias.n15 outputibias.n14 0.155672
R23644 outputibias.n61 outputibias.n33 0.155672
R23645 outputibias.n54 outputibias.n33 0.155672
R23646 outputibias.n54 outputibias.n53 0.155672
R23647 outputibias.n53 outputibias.n37 0.155672
R23648 outputibias.n46 outputibias.n37 0.155672
R23649 outputibias.n46 outputibias.n45 0.155672
R23650 outputibias.n93 outputibias.n65 0.155672
R23651 outputibias.n86 outputibias.n65 0.155672
R23652 outputibias.n86 outputibias.n85 0.155672
R23653 outputibias.n85 outputibias.n69 0.155672
R23654 outputibias.n78 outputibias.n69 0.155672
R23655 outputibias.n78 outputibias.n77 0.155672
R23656 outputibias.n125 outputibias.n97 0.155672
R23657 outputibias.n118 outputibias.n97 0.155672
R23658 outputibias.n118 outputibias.n117 0.155672
R23659 outputibias.n117 outputibias.n101 0.155672
R23660 outputibias.n110 outputibias.n101 0.155672
R23661 outputibias.n110 outputibias.n109 0.155672
R23662 diffpairibias.n0 diffpairibias.t18 436.822
R23663 diffpairibias.n21 diffpairibias.t19 435.479
R23664 diffpairibias.n20 diffpairibias.t16 435.479
R23665 diffpairibias.n19 diffpairibias.t17 435.479
R23666 diffpairibias.n18 diffpairibias.t21 435.479
R23667 diffpairibias.n0 diffpairibias.t22 435.479
R23668 diffpairibias.n1 diffpairibias.t20 435.479
R23669 diffpairibias.n2 diffpairibias.t23 435.479
R23670 diffpairibias.n10 diffpairibias.t0 377.536
R23671 diffpairibias.n10 diffpairibias.t8 376.193
R23672 diffpairibias.n11 diffpairibias.t10 376.193
R23673 diffpairibias.n12 diffpairibias.t6 376.193
R23674 diffpairibias.n13 diffpairibias.t2 376.193
R23675 diffpairibias.n14 diffpairibias.t12 376.193
R23676 diffpairibias.n15 diffpairibias.t4 376.193
R23677 diffpairibias.n16 diffpairibias.t14 376.193
R23678 diffpairibias.n3 diffpairibias.t1 113.368
R23679 diffpairibias.n3 diffpairibias.t9 112.698
R23680 diffpairibias.n4 diffpairibias.t11 112.698
R23681 diffpairibias.n5 diffpairibias.t7 112.698
R23682 diffpairibias.n6 diffpairibias.t3 112.698
R23683 diffpairibias.n7 diffpairibias.t13 112.698
R23684 diffpairibias.n8 diffpairibias.t5 112.698
R23685 diffpairibias.n9 diffpairibias.t15 112.698
R23686 diffpairibias.n17 diffpairibias.n16 4.77242
R23687 diffpairibias.n17 diffpairibias.n9 4.30807
R23688 diffpairibias.n18 diffpairibias.n17 4.13945
R23689 diffpairibias.n16 diffpairibias.n15 1.34352
R23690 diffpairibias.n15 diffpairibias.n14 1.34352
R23691 diffpairibias.n14 diffpairibias.n13 1.34352
R23692 diffpairibias.n13 diffpairibias.n12 1.34352
R23693 diffpairibias.n12 diffpairibias.n11 1.34352
R23694 diffpairibias.n11 diffpairibias.n10 1.34352
R23695 diffpairibias.n2 diffpairibias.n1 1.34352
R23696 diffpairibias.n1 diffpairibias.n0 1.34352
R23697 diffpairibias.n19 diffpairibias.n18 1.34352
R23698 diffpairibias.n20 diffpairibias.n19 1.34352
R23699 diffpairibias.n21 diffpairibias.n20 1.34352
R23700 diffpairibias.n22 diffpairibias.n21 0.862419
R23701 diffpairibias diffpairibias.n22 0.684875
R23702 diffpairibias.n9 diffpairibias.n8 0.672012
R23703 diffpairibias.n8 diffpairibias.n7 0.672012
R23704 diffpairibias.n7 diffpairibias.n6 0.672012
R23705 diffpairibias.n6 diffpairibias.n5 0.672012
R23706 diffpairibias.n5 diffpairibias.n4 0.672012
R23707 diffpairibias.n4 diffpairibias.n3 0.672012
R23708 diffpairibias.n22 diffpairibias.n2 0.190907
C0 minus commonsourceibias 0.322616f
C1 plus commonsourceibias 0.276969f
C2 output outputibias 2.34152f
C3 vdd output 7.23429f
C4 CSoutput output 6.13571f
C5 CSoutput outputibias 0.032386f
C6 vdd CSoutput 0.141661p
C7 minus diffpairibias 2.98e-19
C8 commonsourceibias output 0.006808f
C9 CSoutput minus 2.78935f
C10 vdd plus 0.096545f
C11 commonsourceibias outputibias 0.003832f
C12 plus diffpairibias 2.75e-19
C13 vdd commonsourceibias 0.004218f
C14 CSoutput plus 0.854749f
C15 commonsourceibias diffpairibias 0.052851f
C16 CSoutput commonsourceibias 36.982002f
C17 minus plus 9.1398f
C18 diffpairibias gnd 48.968437f
C19 outputibias gnd 32.465668f
C20 output gnd 15.47879f
C21 commonsourceibias gnd 0.150131p
C22 plus gnd 33.224503f
C23 minus gnd 27.5984f
C24 CSoutput gnd 0.100649p
C25 vdd gnd 0.508603p
C26 diffpairibias.t18 gnd 0.087401f
C27 diffpairibias.t22 gnd 0.087239f
C28 diffpairibias.n0 gnd 0.102784f
C29 diffpairibias.t20 gnd 0.087239f
C30 diffpairibias.n1 gnd 0.050171f
C31 diffpairibias.t23 gnd 0.087239f
C32 diffpairibias.n2 gnd 0.039841f
C33 diffpairibias.t1 gnd 0.083757f
C34 diffpairibias.t9 gnd 0.083392f
C35 diffpairibias.n3 gnd 0.131682f
C36 diffpairibias.t11 gnd 0.083392f
C37 diffpairibias.n4 gnd 0.07027f
C38 diffpairibias.t7 gnd 0.083392f
C39 diffpairibias.n5 gnd 0.07027f
C40 diffpairibias.t3 gnd 0.083392f
C41 diffpairibias.n6 gnd 0.07027f
C42 diffpairibias.t13 gnd 0.083392f
C43 diffpairibias.n7 gnd 0.07027f
C44 diffpairibias.t5 gnd 0.083392f
C45 diffpairibias.n8 gnd 0.07027f
C46 diffpairibias.t15 gnd 0.083392f
C47 diffpairibias.n9 gnd 0.099771f
C48 diffpairibias.t0 gnd 0.08427f
C49 diffpairibias.t8 gnd 0.084123f
C50 diffpairibias.n10 gnd 0.091784f
C51 diffpairibias.t10 gnd 0.084123f
C52 diffpairibias.n11 gnd 0.050681f
C53 diffpairibias.t6 gnd 0.084123f
C54 diffpairibias.n12 gnd 0.050681f
C55 diffpairibias.t2 gnd 0.084123f
C56 diffpairibias.n13 gnd 0.050681f
C57 diffpairibias.t12 gnd 0.084123f
C58 diffpairibias.n14 gnd 0.050681f
C59 diffpairibias.t4 gnd 0.084123f
C60 diffpairibias.n15 gnd 0.050681f
C61 diffpairibias.t14 gnd 0.084123f
C62 diffpairibias.n16 gnd 0.059977f
C63 diffpairibias.n17 gnd 0.226448f
C64 diffpairibias.t21 gnd 0.087239f
C65 diffpairibias.n18 gnd 0.050181f
C66 diffpairibias.t17 gnd 0.087239f
C67 diffpairibias.n19 gnd 0.050171f
C68 diffpairibias.t16 gnd 0.087239f
C69 diffpairibias.n20 gnd 0.050171f
C70 diffpairibias.t19 gnd 0.087239f
C71 diffpairibias.n21 gnd 0.045859f
C72 diffpairibias.n22 gnd 0.046268f
C73 outputibias.t11 gnd 0.11477f
C74 outputibias.t8 gnd 0.115567f
C75 outputibias.n0 gnd 0.130108f
C76 outputibias.n1 gnd 0.001372f
C77 outputibias.n2 gnd 9.76e-19
C78 outputibias.n3 gnd 5.24e-19
C79 outputibias.n4 gnd 0.001239f
C80 outputibias.n5 gnd 5.55e-19
C81 outputibias.n6 gnd 9.76e-19
C82 outputibias.n7 gnd 5.24e-19
C83 outputibias.n8 gnd 0.001239f
C84 outputibias.n9 gnd 5.55e-19
C85 outputibias.n10 gnd 0.004176f
C86 outputibias.t7 gnd 0.00202f
C87 outputibias.n11 gnd 9.3e-19
C88 outputibias.n12 gnd 7.32e-19
C89 outputibias.n13 gnd 5.24e-19
C90 outputibias.n14 gnd 0.02322f
C91 outputibias.n15 gnd 9.76e-19
C92 outputibias.n16 gnd 5.24e-19
C93 outputibias.n17 gnd 5.55e-19
C94 outputibias.n18 gnd 0.001239f
C95 outputibias.n19 gnd 0.001239f
C96 outputibias.n20 gnd 5.55e-19
C97 outputibias.n21 gnd 5.24e-19
C98 outputibias.n22 gnd 9.76e-19
C99 outputibias.n23 gnd 9.76e-19
C100 outputibias.n24 gnd 5.24e-19
C101 outputibias.n25 gnd 5.55e-19
C102 outputibias.n26 gnd 0.001239f
C103 outputibias.n27 gnd 0.002683f
C104 outputibias.n28 gnd 5.55e-19
C105 outputibias.n29 gnd 5.24e-19
C106 outputibias.n30 gnd 0.002256f
C107 outputibias.n31 gnd 0.005781f
C108 outputibias.n32 gnd 0.001372f
C109 outputibias.n33 gnd 9.76e-19
C110 outputibias.n34 gnd 5.24e-19
C111 outputibias.n35 gnd 0.001239f
C112 outputibias.n36 gnd 5.55e-19
C113 outputibias.n37 gnd 9.76e-19
C114 outputibias.n38 gnd 5.24e-19
C115 outputibias.n39 gnd 0.001239f
C116 outputibias.n40 gnd 5.55e-19
C117 outputibias.n41 gnd 0.004176f
C118 outputibias.t5 gnd 0.00202f
C119 outputibias.n42 gnd 9.3e-19
C120 outputibias.n43 gnd 7.32e-19
C121 outputibias.n44 gnd 5.24e-19
C122 outputibias.n45 gnd 0.02322f
C123 outputibias.n46 gnd 9.76e-19
C124 outputibias.n47 gnd 5.24e-19
C125 outputibias.n48 gnd 5.55e-19
C126 outputibias.n49 gnd 0.001239f
C127 outputibias.n50 gnd 0.001239f
C128 outputibias.n51 gnd 5.55e-19
C129 outputibias.n52 gnd 5.24e-19
C130 outputibias.n53 gnd 9.76e-19
C131 outputibias.n54 gnd 9.76e-19
C132 outputibias.n55 gnd 5.24e-19
C133 outputibias.n56 gnd 5.55e-19
C134 outputibias.n57 gnd 0.001239f
C135 outputibias.n58 gnd 0.002683f
C136 outputibias.n59 gnd 5.55e-19
C137 outputibias.n60 gnd 5.24e-19
C138 outputibias.n61 gnd 0.002256f
C139 outputibias.n62 gnd 0.005197f
C140 outputibias.n63 gnd 0.121892f
C141 outputibias.n64 gnd 0.001372f
C142 outputibias.n65 gnd 9.76e-19
C143 outputibias.n66 gnd 5.24e-19
C144 outputibias.n67 gnd 0.001239f
C145 outputibias.n68 gnd 5.55e-19
C146 outputibias.n69 gnd 9.76e-19
C147 outputibias.n70 gnd 5.24e-19
C148 outputibias.n71 gnd 0.001239f
C149 outputibias.n72 gnd 5.55e-19
C150 outputibias.n73 gnd 0.004176f
C151 outputibias.t1 gnd 0.00202f
C152 outputibias.n74 gnd 9.3e-19
C153 outputibias.n75 gnd 7.32e-19
C154 outputibias.n76 gnd 5.24e-19
C155 outputibias.n77 gnd 0.02322f
C156 outputibias.n78 gnd 9.76e-19
C157 outputibias.n79 gnd 5.24e-19
C158 outputibias.n80 gnd 5.55e-19
C159 outputibias.n81 gnd 0.001239f
C160 outputibias.n82 gnd 0.001239f
C161 outputibias.n83 gnd 5.55e-19
C162 outputibias.n84 gnd 5.24e-19
C163 outputibias.n85 gnd 9.76e-19
C164 outputibias.n86 gnd 9.76e-19
C165 outputibias.n87 gnd 5.24e-19
C166 outputibias.n88 gnd 5.55e-19
C167 outputibias.n89 gnd 0.001239f
C168 outputibias.n90 gnd 0.002683f
C169 outputibias.n91 gnd 5.55e-19
C170 outputibias.n92 gnd 5.24e-19
C171 outputibias.n93 gnd 0.002256f
C172 outputibias.n94 gnd 0.005197f
C173 outputibias.n95 gnd 0.064513f
C174 outputibias.n96 gnd 0.001372f
C175 outputibias.n97 gnd 9.76e-19
C176 outputibias.n98 gnd 5.24e-19
C177 outputibias.n99 gnd 0.001239f
C178 outputibias.n100 gnd 5.55e-19
C179 outputibias.n101 gnd 9.76e-19
C180 outputibias.n102 gnd 5.24e-19
C181 outputibias.n103 gnd 0.001239f
C182 outputibias.n104 gnd 5.55e-19
C183 outputibias.n105 gnd 0.004176f
C184 outputibias.t3 gnd 0.00202f
C185 outputibias.n106 gnd 9.3e-19
C186 outputibias.n107 gnd 7.32e-19
C187 outputibias.n108 gnd 5.24e-19
C188 outputibias.n109 gnd 0.02322f
C189 outputibias.n110 gnd 9.76e-19
C190 outputibias.n111 gnd 5.24e-19
C191 outputibias.n112 gnd 5.55e-19
C192 outputibias.n113 gnd 0.001239f
C193 outputibias.n114 gnd 0.001239f
C194 outputibias.n115 gnd 5.55e-19
C195 outputibias.n116 gnd 5.24e-19
C196 outputibias.n117 gnd 9.76e-19
C197 outputibias.n118 gnd 9.76e-19
C198 outputibias.n119 gnd 5.24e-19
C199 outputibias.n120 gnd 5.55e-19
C200 outputibias.n121 gnd 0.001239f
C201 outputibias.n122 gnd 0.002683f
C202 outputibias.n123 gnd 5.55e-19
C203 outputibias.n124 gnd 5.24e-19
C204 outputibias.n125 gnd 0.002256f
C205 outputibias.n126 gnd 0.005197f
C206 outputibias.n127 gnd 0.084814f
C207 outputibias.t2 gnd 0.108319f
C208 outputibias.t0 gnd 0.108319f
C209 outputibias.t4 gnd 0.108319f
C210 outputibias.t6 gnd 0.109238f
C211 outputibias.n128 gnd 0.134674f
C212 outputibias.n129 gnd 0.07244f
C213 outputibias.n130 gnd 0.079818f
C214 outputibias.n131 gnd 0.164901f
C215 outputibias.t10 gnd 0.11477f
C216 outputibias.n132 gnd 0.067481f
C217 outputibias.t9 gnd 0.11477f
C218 outputibias.n133 gnd 0.065115f
C219 outputibias.n134 gnd 0.029159f
C220 minus.n0 gnd 0.032888f
C221 minus.t27 gnd 0.332265f
C222 minus.n1 gnd 0.153313f
C223 minus.n2 gnd 0.032888f
C224 minus.t6 gnd 0.332265f
C225 minus.n3 gnd 0.150271f
C226 minus.n4 gnd 0.032888f
C227 minus.t24 gnd 0.332265f
C228 minus.n5 gnd 0.150271f
C229 minus.n6 gnd 0.032888f
C230 minus.t8 gnd 0.332265f
C231 minus.n7 gnd 0.153313f
C232 minus.t12 gnd 0.341211f
C233 minus.t18 gnd 0.332265f
C234 minus.n8 gnd 0.157204f
C235 minus.n9 gnd 0.142301f
C236 minus.n10 gnd 0.133539f
C237 minus.n11 gnd 0.032888f
C238 minus.n12 gnd 0.007463f
C239 minus.t13 gnd 0.332265f
C240 minus.n13 gnd 0.153617f
C241 minus.n14 gnd 0.007463f
C242 minus.n15 gnd 0.032888f
C243 minus.n16 gnd 0.032888f
C244 minus.n17 gnd 0.032888f
C245 minus.t19 gnd 0.332265f
C246 minus.n18 gnd 0.153515f
C247 minus.n19 gnd 0.007463f
C248 minus.t22 gnd 0.332265f
C249 minus.n20 gnd 0.153515f
C250 minus.n21 gnd 0.032888f
C251 minus.n22 gnd 0.032888f
C252 minus.n23 gnd 0.032888f
C253 minus.n24 gnd 0.007463f
C254 minus.t20 gnd 0.332265f
C255 minus.n25 gnd 0.153617f
C256 minus.n26 gnd 0.007463f
C257 minus.n27 gnd 0.032888f
C258 minus.n28 gnd 0.032888f
C259 minus.n29 gnd 0.032888f
C260 minus.t15 gnd 0.332265f
C261 minus.n30 gnd 0.150474f
C262 minus.n31 gnd 0.007463f
C263 minus.t9 gnd 0.332265f
C264 minus.n32 gnd 0.149866f
C265 minus.n33 gnd 0.369096f
C266 minus.n34 gnd 0.032888f
C267 minus.t16 gnd 0.332265f
C268 minus.t28 gnd 0.332265f
C269 minus.n35 gnd 0.032888f
C270 minus.t21 gnd 0.332265f
C271 minus.n36 gnd 0.032888f
C272 minus.t14 gnd 0.332265f
C273 minus.n37 gnd 0.153617f
C274 minus.n38 gnd 0.032888f
C275 minus.t23 gnd 0.332265f
C276 minus.t11 gnd 0.332265f
C277 minus.n39 gnd 0.032888f
C278 minus.t5 gnd 0.332265f
C279 minus.n40 gnd 0.153515f
C280 minus.n41 gnd 0.032888f
C281 minus.t17 gnd 0.332265f
C282 minus.t10 gnd 0.332265f
C283 minus.n42 gnd 0.032888f
C284 minus.t25 gnd 0.332265f
C285 minus.n43 gnd 0.153313f
C286 minus.t26 gnd 0.341211f
C287 minus.t7 gnd 0.332265f
C288 minus.n44 gnd 0.157204f
C289 minus.n45 gnd 0.142301f
C290 minus.n46 gnd 0.133539f
C291 minus.n47 gnd 0.032888f
C292 minus.n48 gnd 0.007463f
C293 minus.n49 gnd 0.153617f
C294 minus.n50 gnd 0.007463f
C295 minus.n51 gnd 0.150271f
C296 minus.n52 gnd 0.032888f
C297 minus.n53 gnd 0.032888f
C298 minus.n54 gnd 0.032888f
C299 minus.n55 gnd 0.007463f
C300 minus.n56 gnd 0.153515f
C301 minus.n57 gnd 0.150271f
C302 minus.n58 gnd 0.007463f
C303 minus.n59 gnd 0.032888f
C304 minus.n60 gnd 0.032888f
C305 minus.n61 gnd 0.032888f
C306 minus.n62 gnd 0.007463f
C307 minus.n63 gnd 0.153313f
C308 minus.n64 gnd 0.150474f
C309 minus.n65 gnd 0.007463f
C310 minus.n66 gnd 0.149866f
C311 minus.n67 gnd 0.998001f
C312 minus.n68 gnd 1.51388f
C313 minus.t1 gnd 0.010139f
C314 minus.t4 gnd 0.010139f
C315 minus.n69 gnd 0.033338f
C316 minus.t2 gnd 0.010139f
C317 minus.t0 gnd 0.010139f
C318 minus.n70 gnd 0.032881f
C319 minus.n71 gnd 0.280622f
C320 minus.t3 gnd 0.056429f
C321 minus.n72 gnd 0.153133f
C322 minus.n73 gnd 2.08976f
C323 a_n2903_n3924.t18 gnd 0.108618f
C324 a_n2903_n3924.t13 gnd 1.12888f
C325 a_n2903_n3924.n0 gnd 0.383133f
C326 a_n2903_n3924.t34 gnd 1.40337f
C327 a_n2903_n3924.n1 gnd 1.48426f
C328 a_n2903_n3924.t51 gnd 1.12888f
C329 a_n2903_n3924.n2 gnd 0.383133f
C330 a_n2903_n3924.t39 gnd 0.108618f
C331 a_n2903_n3924.t42 gnd 0.108618f
C332 a_n2903_n3924.n3 gnd 0.887099f
C333 a_n2903_n3924.n4 gnd 0.359777f
C334 a_n2903_n3924.t5 gnd 0.108618f
C335 a_n2903_n3924.t3 gnd 0.108618f
C336 a_n2903_n3924.n5 gnd 0.887099f
C337 a_n2903_n3924.n6 gnd 0.359777f
C338 a_n2903_n3924.t41 gnd 0.108618f
C339 a_n2903_n3924.t1 gnd 0.108618f
C340 a_n2903_n3924.n7 gnd 0.887099f
C341 a_n2903_n3924.n8 gnd 0.359777f
C342 a_n2903_n3924.t55 gnd 0.108618f
C343 a_n2903_n3924.t50 gnd 0.108618f
C344 a_n2903_n3924.n9 gnd 0.887099f
C345 a_n2903_n3924.n10 gnd 0.359777f
C346 a_n2903_n3924.t7 gnd 0.108618f
C347 a_n2903_n3924.t36 gnd 0.108618f
C348 a_n2903_n3924.n11 gnd 0.887099f
C349 a_n2903_n3924.n12 gnd 0.359777f
C350 a_n2903_n3924.t2 gnd 1.12888f
C351 a_n2903_n3924.n13 gnd 0.974186f
C352 a_n2903_n3924.t49 gnd 1.40461f
C353 a_n2903_n3924.t9 gnd 1.40261f
C354 a_n2903_n3924.n14 gnd 1.26893f
C355 a_n2903_n3924.t46 gnd 1.40261f
C356 a_n2903_n3924.n15 gnd 0.892855f
C357 a_n2903_n3924.t44 gnd 1.40261f
C358 a_n2903_n3924.n16 gnd 0.987884f
C359 a_n2903_n3924.t48 gnd 1.40261f
C360 a_n2903_n3924.n17 gnd 0.987884f
C361 a_n2903_n3924.t45 gnd 1.40261f
C362 a_n2903_n3924.n18 gnd 0.987884f
C363 a_n2903_n3924.t4 gnd 1.40261f
C364 a_n2903_n3924.n19 gnd 0.972113f
C365 a_n2903_n3924.n20 gnd 0.533935f
C366 a_n2903_n3924.n21 gnd 1.01395f
C367 a_n2903_n3924.t15 gnd 1.12888f
C368 a_n2903_n3924.n22 gnd 0.619233f
C369 a_n2903_n3924.t25 gnd 0.108618f
C370 a_n2903_n3924.t11 gnd 0.108618f
C371 a_n2903_n3924.n23 gnd 0.887098f
C372 a_n2903_n3924.n24 gnd 0.359779f
C373 a_n2903_n3924.t16 gnd 0.108618f
C374 a_n2903_n3924.t31 gnd 0.108618f
C375 a_n2903_n3924.n25 gnd 0.887098f
C376 a_n2903_n3924.n26 gnd 0.359779f
C377 a_n2903_n3924.t20 gnd 0.108618f
C378 a_n2903_n3924.t24 gnd 0.108618f
C379 a_n2903_n3924.n27 gnd 0.887098f
C380 a_n2903_n3924.n28 gnd 0.359779f
C381 a_n2903_n3924.t14 gnd 0.108618f
C382 a_n2903_n3924.t21 gnd 0.108618f
C383 a_n2903_n3924.n29 gnd 0.887098f
C384 a_n2903_n3924.n30 gnd 0.359779f
C385 a_n2903_n3924.t29 gnd 0.108618f
C386 a_n2903_n3924.t23 gnd 0.108618f
C387 a_n2903_n3924.n31 gnd 0.887098f
C388 a_n2903_n3924.n32 gnd 0.359779f
C389 a_n2903_n3924.t26 gnd 1.12888f
C390 a_n2903_n3924.n33 gnd 0.383138f
C391 a_n2903_n3924.t0 gnd 1.12888f
C392 a_n2903_n3924.n34 gnd 0.383138f
C393 a_n2903_n3924.t54 gnd 0.108618f
C394 a_n2903_n3924.t37 gnd 0.108618f
C395 a_n2903_n3924.n35 gnd 0.887098f
C396 a_n2903_n3924.n36 gnd 0.359779f
C397 a_n2903_n3924.t40 gnd 0.108618f
C398 a_n2903_n3924.t43 gnd 0.108618f
C399 a_n2903_n3924.n37 gnd 0.887098f
C400 a_n2903_n3924.n38 gnd 0.359779f
C401 a_n2903_n3924.t8 gnd 0.108618f
C402 a_n2903_n3924.t6 gnd 0.108618f
C403 a_n2903_n3924.n39 gnd 0.887098f
C404 a_n2903_n3924.n40 gnd 0.359779f
C405 a_n2903_n3924.t47 gnd 0.108618f
C406 a_n2903_n3924.t38 gnd 0.108618f
C407 a_n2903_n3924.n41 gnd 0.887098f
C408 a_n2903_n3924.n42 gnd 0.359779f
C409 a_n2903_n3924.t53 gnd 0.108618f
C410 a_n2903_n3924.t52 gnd 0.108618f
C411 a_n2903_n3924.n43 gnd 0.887098f
C412 a_n2903_n3924.n44 gnd 0.359779f
C413 a_n2903_n3924.t35 gnd 1.12888f
C414 a_n2903_n3924.n45 gnd 0.619233f
C415 a_n2903_n3924.n46 gnd 1.01395f
C416 a_n2903_n3924.t17 gnd 1.12888f
C417 a_n2903_n3924.n47 gnd 0.97419f
C418 a_n2903_n3924.t22 gnd 0.108618f
C419 a_n2903_n3924.t10 gnd 0.108618f
C420 a_n2903_n3924.n48 gnd 0.887099f
C421 a_n2903_n3924.n49 gnd 0.359777f
C422 a_n2903_n3924.t19 gnd 0.108618f
C423 a_n2903_n3924.t30 gnd 0.108618f
C424 a_n2903_n3924.n50 gnd 0.887099f
C425 a_n2903_n3924.n51 gnd 0.359777f
C426 a_n2903_n3924.t32 gnd 0.108618f
C427 a_n2903_n3924.t28 gnd 0.108618f
C428 a_n2903_n3924.n52 gnd 0.887099f
C429 a_n2903_n3924.n53 gnd 0.359777f
C430 a_n2903_n3924.t12 gnd 0.108618f
C431 a_n2903_n3924.t27 gnd 0.108618f
C432 a_n2903_n3924.n54 gnd 0.887099f
C433 a_n2903_n3924.n55 gnd 0.359777f
C434 a_n2903_n3924.n56 gnd 0.359776f
C435 a_n2903_n3924.n57 gnd 0.887101f
C436 a_n2903_n3924.t33 gnd 0.108618f
C437 plus.n0 gnd 0.023857f
C438 plus.t23 gnd 0.241028f
C439 plus.n1 gnd 0.023857f
C440 plus.t13 gnd 0.241028f
C441 plus.n2 gnd 0.023857f
C442 plus.t27 gnd 0.241028f
C443 plus.t22 gnd 0.241028f
C444 plus.n3 gnd 0.111435f
C445 plus.n4 gnd 0.023857f
C446 plus.t7 gnd 0.241028f
C447 plus.n5 gnd 0.023857f
C448 plus.t18 gnd 0.241028f
C449 plus.t14 gnd 0.241028f
C450 plus.n6 gnd 0.111361f
C451 plus.n7 gnd 0.023857f
C452 plus.t24 gnd 0.241028f
C453 plus.n8 gnd 0.023857f
C454 plus.t17 gnd 0.241028f
C455 plus.t9 gnd 0.241028f
C456 plus.n9 gnd 0.111214f
C457 plus.t12 gnd 0.247518f
C458 plus.t15 gnd 0.241028f
C459 plus.n10 gnd 0.114037f
C460 plus.n11 gnd 0.103227f
C461 plus.n12 gnd 0.096871f
C462 plus.n13 gnd 0.023857f
C463 plus.n14 gnd 0.005414f
C464 plus.n15 gnd 0.111435f
C465 plus.n16 gnd 0.005414f
C466 plus.n17 gnd 0.109008f
C467 plus.n18 gnd 0.023857f
C468 plus.n19 gnd 0.023857f
C469 plus.n20 gnd 0.023857f
C470 plus.n21 gnd 0.005414f
C471 plus.n22 gnd 0.111361f
C472 plus.n23 gnd 0.109008f
C473 plus.n24 gnd 0.005414f
C474 plus.n25 gnd 0.023857f
C475 plus.n26 gnd 0.023857f
C476 plus.n27 gnd 0.023857f
C477 plus.n28 gnd 0.005414f
C478 plus.n29 gnd 0.111214f
C479 plus.n30 gnd 0.109155f
C480 plus.n31 gnd 0.005414f
C481 plus.n32 gnd 0.108714f
C482 plus.n33 gnd 0.261581f
C483 plus.n34 gnd 0.023857f
C484 plus.t16 gnd 0.241028f
C485 plus.n35 gnd 0.111214f
C486 plus.t28 gnd 0.241028f
C487 plus.n36 gnd 0.023857f
C488 plus.t19 gnd 0.241028f
C489 plus.n37 gnd 0.109008f
C490 plus.n38 gnd 0.023857f
C491 plus.t11 gnd 0.241028f
C492 plus.n39 gnd 0.109008f
C493 plus.t6 gnd 0.241028f
C494 plus.n40 gnd 0.023857f
C495 plus.t20 gnd 0.241028f
C496 plus.n41 gnd 0.111214f
C497 plus.t25 gnd 0.247518f
C498 plus.t5 gnd 0.241028f
C499 plus.n42 gnd 0.114037f
C500 plus.n43 gnd 0.103227f
C501 plus.n44 gnd 0.096871f
C502 plus.n45 gnd 0.023857f
C503 plus.n46 gnd 0.005414f
C504 plus.t26 gnd 0.241028f
C505 plus.n47 gnd 0.111435f
C506 plus.n48 gnd 0.005414f
C507 plus.n49 gnd 0.023857f
C508 plus.n50 gnd 0.023857f
C509 plus.n51 gnd 0.023857f
C510 plus.n52 gnd 0.111361f
C511 plus.n53 gnd 0.005414f
C512 plus.t10 gnd 0.241028f
C513 plus.n54 gnd 0.111361f
C514 plus.n55 gnd 0.023857f
C515 plus.n56 gnd 0.023857f
C516 plus.n57 gnd 0.023857f
C517 plus.n58 gnd 0.005414f
C518 plus.t8 gnd 0.241028f
C519 plus.n59 gnd 0.111435f
C520 plus.n60 gnd 0.005414f
C521 plus.n61 gnd 0.023857f
C522 plus.n62 gnd 0.023857f
C523 plus.n63 gnd 0.023857f
C524 plus.n64 gnd 0.109155f
C525 plus.n65 gnd 0.005414f
C526 plus.t21 gnd 0.241028f
C527 plus.n66 gnd 0.108714f
C528 plus.n67 gnd 0.714366f
C529 plus.n68 gnd 1.08878f
C530 plus.t3 gnd 0.041185f
C531 plus.t4 gnd 0.007355f
C532 plus.t1 gnd 0.007355f
C533 plus.n69 gnd 0.023852f
C534 plus.n70 gnd 0.185165f
C535 plus.t0 gnd 0.007355f
C536 plus.t2 gnd 0.007355f
C537 plus.n71 gnd 0.023852f
C538 plus.n72 gnd 0.138989f
C539 plus.n73 gnd 2.67147f
C540 output.t13 gnd 0.464308f
C541 output.t3 gnd 0.044422f
C542 output.t8 gnd 0.044422f
C543 output.n0 gnd 0.364624f
C544 output.n1 gnd 0.614102f
C545 output.t12 gnd 0.044422f
C546 output.t4 gnd 0.044422f
C547 output.n2 gnd 0.364624f
C548 output.n3 gnd 0.350265f
C549 output.t6 gnd 0.044422f
C550 output.t5 gnd 0.044422f
C551 output.n4 gnd 0.364624f
C552 output.n5 gnd 0.350265f
C553 output.t11 gnd 0.044422f
C554 output.t14 gnd 0.044422f
C555 output.n6 gnd 0.364624f
C556 output.n7 gnd 0.350265f
C557 output.t16 gnd 0.044422f
C558 output.t9 gnd 0.044422f
C559 output.n8 gnd 0.364624f
C560 output.n9 gnd 0.350265f
C561 output.t10 gnd 0.044422f
C562 output.t17 gnd 0.044422f
C563 output.n10 gnd 0.364624f
C564 output.n11 gnd 0.350265f
C565 output.t2 gnd 0.044422f
C566 output.t7 gnd 0.044422f
C567 output.n12 gnd 0.364624f
C568 output.n13 gnd 0.350265f
C569 output.t15 gnd 0.462979f
C570 output.n14 gnd 0.28994f
C571 output.n15 gnd 0.015803f
C572 output.n16 gnd 0.011243f
C573 output.n17 gnd 0.006041f
C574 output.n18 gnd 0.01428f
C575 output.n19 gnd 0.006397f
C576 output.n20 gnd 0.011243f
C577 output.n21 gnd 0.006041f
C578 output.n22 gnd 0.01428f
C579 output.n23 gnd 0.006397f
C580 output.n24 gnd 0.048111f
C581 output.t0 gnd 0.023274f
C582 output.n25 gnd 0.01071f
C583 output.n26 gnd 0.008435f
C584 output.n27 gnd 0.006041f
C585 output.n28 gnd 0.267512f
C586 output.n29 gnd 0.011243f
C587 output.n30 gnd 0.006041f
C588 output.n31 gnd 0.006397f
C589 output.n32 gnd 0.01428f
C590 output.n33 gnd 0.01428f
C591 output.n34 gnd 0.006397f
C592 output.n35 gnd 0.006041f
C593 output.n36 gnd 0.011243f
C594 output.n37 gnd 0.011243f
C595 output.n38 gnd 0.006041f
C596 output.n39 gnd 0.006397f
C597 output.n40 gnd 0.01428f
C598 output.n41 gnd 0.030913f
C599 output.n42 gnd 0.006397f
C600 output.n43 gnd 0.006041f
C601 output.n44 gnd 0.025987f
C602 output.n45 gnd 0.097665f
C603 output.n46 gnd 0.015803f
C604 output.n47 gnd 0.011243f
C605 output.n48 gnd 0.006041f
C606 output.n49 gnd 0.01428f
C607 output.n50 gnd 0.006397f
C608 output.n51 gnd 0.011243f
C609 output.n52 gnd 0.006041f
C610 output.n53 gnd 0.01428f
C611 output.n54 gnd 0.006397f
C612 output.n55 gnd 0.048111f
C613 output.t18 gnd 0.023274f
C614 output.n56 gnd 0.01071f
C615 output.n57 gnd 0.008435f
C616 output.n58 gnd 0.006041f
C617 output.n59 gnd 0.267512f
C618 output.n60 gnd 0.011243f
C619 output.n61 gnd 0.006041f
C620 output.n62 gnd 0.006397f
C621 output.n63 gnd 0.01428f
C622 output.n64 gnd 0.01428f
C623 output.n65 gnd 0.006397f
C624 output.n66 gnd 0.006041f
C625 output.n67 gnd 0.011243f
C626 output.n68 gnd 0.011243f
C627 output.n69 gnd 0.006041f
C628 output.n70 gnd 0.006397f
C629 output.n71 gnd 0.01428f
C630 output.n72 gnd 0.030913f
C631 output.n73 gnd 0.006397f
C632 output.n74 gnd 0.006041f
C633 output.n75 gnd 0.025987f
C634 output.n76 gnd 0.09306f
C635 output.n77 gnd 1.65264f
C636 output.n78 gnd 0.015803f
C637 output.n79 gnd 0.011243f
C638 output.n80 gnd 0.006041f
C639 output.n81 gnd 0.01428f
C640 output.n82 gnd 0.006397f
C641 output.n83 gnd 0.011243f
C642 output.n84 gnd 0.006041f
C643 output.n85 gnd 0.01428f
C644 output.n86 gnd 0.006397f
C645 output.n87 gnd 0.048111f
C646 output.t1 gnd 0.023274f
C647 output.n88 gnd 0.01071f
C648 output.n89 gnd 0.008435f
C649 output.n90 gnd 0.006041f
C650 output.n91 gnd 0.267512f
C651 output.n92 gnd 0.011243f
C652 output.n93 gnd 0.006041f
C653 output.n94 gnd 0.006397f
C654 output.n95 gnd 0.01428f
C655 output.n96 gnd 0.01428f
C656 output.n97 gnd 0.006397f
C657 output.n98 gnd 0.006041f
C658 output.n99 gnd 0.011243f
C659 output.n100 gnd 0.011243f
C660 output.n101 gnd 0.006041f
C661 output.n102 gnd 0.006397f
C662 output.n103 gnd 0.01428f
C663 output.n104 gnd 0.030913f
C664 output.n105 gnd 0.006397f
C665 output.n106 gnd 0.006041f
C666 output.n107 gnd 0.025987f
C667 output.n108 gnd 0.09306f
C668 output.n109 gnd 0.713089f
C669 output.n110 gnd 0.015803f
C670 output.n111 gnd 0.011243f
C671 output.n112 gnd 0.006041f
C672 output.n113 gnd 0.01428f
C673 output.n114 gnd 0.006397f
C674 output.n115 gnd 0.011243f
C675 output.n116 gnd 0.006041f
C676 output.n117 gnd 0.01428f
C677 output.n118 gnd 0.006397f
C678 output.n119 gnd 0.048111f
C679 output.t19 gnd 0.023274f
C680 output.n120 gnd 0.01071f
C681 output.n121 gnd 0.008435f
C682 output.n122 gnd 0.006041f
C683 output.n123 gnd 0.267512f
C684 output.n124 gnd 0.011243f
C685 output.n125 gnd 0.006041f
C686 output.n126 gnd 0.006397f
C687 output.n127 gnd 0.01428f
C688 output.n128 gnd 0.01428f
C689 output.n129 gnd 0.006397f
C690 output.n130 gnd 0.006041f
C691 output.n131 gnd 0.011243f
C692 output.n132 gnd 0.011243f
C693 output.n133 gnd 0.006041f
C694 output.n134 gnd 0.006397f
C695 output.n135 gnd 0.01428f
C696 output.n136 gnd 0.030913f
C697 output.n137 gnd 0.006397f
C698 output.n138 gnd 0.006041f
C699 output.n139 gnd 0.025987f
C700 output.n140 gnd 0.09306f
C701 output.n141 gnd 1.67353f
C702 a_n2650_8322.t13 gnd 0.098003f
C703 a_n2650_8322.t33 gnd 20.3315f
C704 a_n2650_8322.t30 gnd 20.189f
C705 a_n2650_8322.t32 gnd 20.189f
C706 a_n2650_8322.t28 gnd 20.3315f
C707 a_n2650_8322.t31 gnd 20.189f
C708 a_n2650_8322.t29 gnd 28.6388f
C709 a_n2650_8322.t23 gnd 0.917645f
C710 a_n2650_8322.t26 gnd 0.098003f
C711 a_n2650_8322.t18 gnd 0.098003f
C712 a_n2650_8322.n0 gnd 0.690329f
C713 a_n2650_8322.n1 gnd 0.771341f
C714 a_n2650_8322.t10 gnd 0.098003f
C715 a_n2650_8322.t9 gnd 0.098003f
C716 a_n2650_8322.n2 gnd 0.690329f
C717 a_n2650_8322.n3 gnd 0.391909f
C718 a_n2650_8322.t21 gnd 0.098003f
C719 a_n2650_8322.t15 gnd 0.098003f
C720 a_n2650_8322.n4 gnd 0.690329f
C721 a_n2650_8322.n5 gnd 0.391909f
C722 a_n2650_8322.t19 gnd 0.098003f
C723 a_n2650_8322.t17 gnd 0.098003f
C724 a_n2650_8322.n6 gnd 0.690329f
C725 a_n2650_8322.n7 gnd 0.391909f
C726 a_n2650_8322.t8 gnd 0.915818f
C727 a_n2650_8322.n8 gnd 1.70901f
C728 a_n2650_8322.t3 gnd 0.917645f
C729 a_n2650_8322.t7 gnd 0.098003f
C730 a_n2650_8322.t6 gnd 0.098003f
C731 a_n2650_8322.n9 gnd 0.690329f
C732 a_n2650_8322.n10 gnd 0.771341f
C733 a_n2650_8322.t1 gnd 0.915818f
C734 a_n2650_8322.n11 gnd 0.38815f
C735 a_n2650_8322.t4 gnd 0.915818f
C736 a_n2650_8322.n12 gnd 0.38815f
C737 a_n2650_8322.t2 gnd 0.098003f
C738 a_n2650_8322.t0 gnd 0.098003f
C739 a_n2650_8322.n13 gnd 0.690329f
C740 a_n2650_8322.n14 gnd 0.391909f
C741 a_n2650_8322.t5 gnd 0.915818f
C742 a_n2650_8322.n15 gnd 1.27346f
C743 a_n2650_8322.n16 gnd 2.08071f
C744 a_n2650_8322.n17 gnd 3.34289f
C745 a_n2650_8322.t22 gnd 0.915818f
C746 a_n2650_8322.n18 gnd 0.996146f
C747 a_n2650_8322.t12 gnd 0.098003f
C748 a_n2650_8322.t11 gnd 0.098003f
C749 a_n2650_8322.n19 gnd 0.690329f
C750 a_n2650_8322.n20 gnd 0.391909f
C751 a_n2650_8322.t24 gnd 0.098003f
C752 a_n2650_8322.t14 gnd 0.098003f
C753 a_n2650_8322.n21 gnd 0.690329f
C754 a_n2650_8322.n22 gnd 0.391909f
C755 a_n2650_8322.t25 gnd 0.917643f
C756 a_n2650_8322.t20 gnd 0.098003f
C757 a_n2650_8322.t16 gnd 0.098003f
C758 a_n2650_8322.n23 gnd 0.690329f
C759 a_n2650_8322.n24 gnd 0.771343f
C760 a_n2650_8322.n25 gnd 0.391907f
C761 a_n2650_8322.n26 gnd 0.690331f
C762 a_n2650_8322.t27 gnd 0.098003f
C763 a_n2472_13878.t13 gnd 0.187752f
C764 a_n2472_13878.t15 gnd 0.187752f
C765 a_n2472_13878.t7 gnd 0.187752f
C766 a_n2472_13878.n0 gnd 1.47995f
C767 a_n2472_13878.t12 gnd 0.187752f
C768 a_n2472_13878.t6 gnd 0.187752f
C769 a_n2472_13878.n1 gnd 1.47838f
C770 a_n2472_13878.n2 gnd 2.06575f
C771 a_n2472_13878.t2 gnd 0.187752f
C772 a_n2472_13878.t4 gnd 0.187752f
C773 a_n2472_13878.n3 gnd 1.47838f
C774 a_n2472_13878.n4 gnd 1.00763f
C775 a_n2472_13878.t14 gnd 0.187752f
C776 a_n2472_13878.t3 gnd 0.187752f
C777 a_n2472_13878.n5 gnd 1.47838f
C778 a_n2472_13878.n6 gnd 1.00763f
C779 a_n2472_13878.t11 gnd 0.187752f
C780 a_n2472_13878.t1 gnd 0.187752f
C781 a_n2472_13878.n7 gnd 1.47838f
C782 a_n2472_13878.n8 gnd 4.40971f
C783 a_n2472_13878.t21 gnd 1.75801f
C784 a_n2472_13878.t24 gnd 0.187752f
C785 a_n2472_13878.t25 gnd 0.187752f
C786 a_n2472_13878.n9 gnd 1.32252f
C787 a_n2472_13878.n10 gnd 1.47772f
C788 a_n2472_13878.t20 gnd 1.75451f
C789 a_n2472_13878.n11 gnd 0.743612f
C790 a_n2472_13878.t23 gnd 1.75451f
C791 a_n2472_13878.n12 gnd 0.743612f
C792 a_n2472_13878.t26 gnd 0.187752f
C793 a_n2472_13878.t27 gnd 0.187752f
C794 a_n2472_13878.n13 gnd 1.32252f
C795 a_n2472_13878.n14 gnd 0.750813f
C796 a_n2472_13878.t22 gnd 1.75451f
C797 a_n2472_13878.n15 gnd 2.43968f
C798 a_n2472_13878.n16 gnd 3.23176f
C799 a_n2472_13878.t16 gnd 0.187752f
C800 a_n2472_13878.t5 gnd 0.187752f
C801 a_n2472_13878.n17 gnd 1.47838f
C802 a_n2472_13878.n18 gnd 2.22265f
C803 a_n2472_13878.t8 gnd 0.187752f
C804 a_n2472_13878.t9 gnd 0.187752f
C805 a_n2472_13878.n19 gnd 1.47838f
C806 a_n2472_13878.n20 gnd 0.655033f
C807 a_n2472_13878.t17 gnd 0.187752f
C808 a_n2472_13878.t18 gnd 0.187752f
C809 a_n2472_13878.n21 gnd 1.47838f
C810 a_n2472_13878.n22 gnd 0.655033f
C811 a_n2472_13878.t0 gnd 0.187752f
C812 a_n2472_13878.t10 gnd 0.187752f
C813 a_n2472_13878.n23 gnd 1.47838f
C814 a_n2472_13878.n24 gnd 1.32888f
C815 a_n2472_13878.n25 gnd 1.48083f
C816 a_n2472_13878.t19 gnd 0.187752f
C817 a_n2650_13878.n0 gnd 0.21772f
C818 a_n2650_13878.n1 gnd 0.942749f
C819 a_n2650_13878.n2 gnd 0.21772f
C820 a_n2650_13878.n3 gnd 0.506761f
C821 a_n2650_13878.n4 gnd 0.21772f
C822 a_n2650_13878.n5 gnd 0.21772f
C823 a_n2650_13878.n6 gnd 0.809668f
C824 a_n2650_13878.n7 gnd 0.809584f
C825 a_n2650_13878.n8 gnd 0.20658f
C826 a_n2650_13878.n9 gnd 0.15215f
C827 a_n2650_13878.n10 gnd 0.239132f
C828 a_n2650_13878.n11 gnd 0.184702f
C829 a_n2650_13878.n12 gnd 0.20658f
C830 a_n2650_13878.n13 gnd 0.15215f
C831 a_n2650_13878.n14 gnd 0.864014f
C832 a_n2650_13878.n15 gnd 0.21772f
C833 a_n2650_13878.n16 gnd 0.702566f
C834 a_n2650_13878.n17 gnd 0.21772f
C835 a_n2650_13878.n18 gnd 0.507263f
C836 a_n2650_13878.n19 gnd 0.21772f
C837 a_n2650_13878.n20 gnd 0.561693f
C838 a_n2650_13878.n21 gnd 0.21772f
C839 a_n2650_13878.n22 gnd 0.901302f
C840 a_n2650_13878.n23 gnd 3.52187f
C841 a_n2650_13878.n24 gnd 2.68251f
C842 a_n2650_13878.n25 gnd 3.77855f
C843 a_n2650_13878.n26 gnd 1.79246f
C844 a_n2650_13878.n27 gnd 1.20779f
C845 a_n2650_13878.n28 gnd 2.25634f
C846 a_n2650_13878.n29 gnd 1.18856f
C847 a_n2650_13878.n30 gnd 1.20779f
C848 a_n2650_13878.n31 gnd 0.732993f
C849 a_n2650_13878.n32 gnd 0.732995f
C850 a_n2650_13878.n33 gnd 3.25198f
C851 a_n2650_13878.n34 gnd 0.008736f
C852 a_n2650_13878.n35 gnd 4.21e-19
C853 a_n2650_13878.n37 gnd 0.008429f
C854 a_n2650_13878.n38 gnd 0.012257f
C855 a_n2650_13878.n39 gnd 0.008109f
C856 a_n2650_13878.n40 gnd 0.287607f
C857 a_n2650_13878.n41 gnd 0.008736f
C858 a_n2650_13878.n42 gnd 4.21e-19
C859 a_n2650_13878.n44 gnd 0.008429f
C860 a_n2650_13878.n45 gnd 0.012257f
C861 a_n2650_13878.n46 gnd 0.008109f
C862 a_n2650_13878.n47 gnd 0.287607f
C863 a_n2650_13878.n48 gnd 0.008429f
C864 a_n2650_13878.n49 gnd 0.287607f
C865 a_n2650_13878.n50 gnd 0.008429f
C866 a_n2650_13878.n51 gnd 0.287607f
C867 a_n2650_13878.n52 gnd 0.008429f
C868 a_n2650_13878.n53 gnd 0.287607f
C869 a_n2650_13878.n54 gnd 0.008429f
C870 a_n2650_13878.n55 gnd 1.58548f
C871 a_n2650_13878.n56 gnd 0.287607f
C872 a_n2650_13878.n57 gnd 0.008736f
C873 a_n2650_13878.n58 gnd 4.21e-19
C874 a_n2650_13878.n60 gnd 0.008429f
C875 a_n2650_13878.n61 gnd 0.012257f
C876 a_n2650_13878.n62 gnd 0.008109f
C877 a_n2650_13878.n63 gnd 0.008736f
C878 a_n2650_13878.n64 gnd 4.21e-19
C879 a_n2650_13878.n66 gnd 0.008429f
C880 a_n2650_13878.n67 gnd 0.012257f
C881 a_n2650_13878.n68 gnd 0.008109f
C882 a_n2650_13878.n69 gnd 0.287607f
C883 a_n2650_13878.n70 gnd 0.287607f
C884 a_n2650_13878.t25 gnd 0.151013f
C885 a_n2650_13878.t31 gnd 1.41401f
C886 a_n2650_13878.t35 gnd 0.151013f
C887 a_n2650_13878.t33 gnd 0.151013f
C888 a_n2650_13878.n71 gnd 1.06373f
C889 a_n2650_13878.t23 gnd 0.151013f
C890 a_n2650_13878.t15 gnd 0.151013f
C891 a_n2650_13878.n72 gnd 1.06373f
C892 a_n2650_13878.t18 gnd 0.702438f
C893 a_n2650_13878.n73 gnd 0.305176f
C894 a_n2650_13878.t8 gnd 0.702438f
C895 a_n2650_13878.t32 gnd 0.702438f
C896 a_n2650_13878.n74 gnd 0.308697f
C897 a_n2650_13878.t30 gnd 0.702438f
C898 a_n2650_13878.t76 gnd 0.702438f
C899 a_n2650_13878.n75 gnd 0.305176f
C900 a_n2650_13878.t91 gnd 0.702438f
C901 a_n2650_13878.t94 gnd 0.702438f
C902 a_n2650_13878.n76 gnd 0.308697f
C903 a_n2650_13878.t70 gnd 0.702438f
C904 a_n2650_13878.t44 gnd 0.702438f
C905 a_n2650_13878.t12 gnd 0.702438f
C906 a_n2650_13878.t28 gnd 0.702438f
C907 a_n2650_13878.n77 gnd 0.308697f
C908 a_n2650_13878.t36 gnd 0.702438f
C909 a_n2650_13878.t38 gnd 0.702438f
C910 a_n2650_13878.t16 gnd 0.702438f
C911 a_n2650_13878.n78 gnd 0.304914f
C912 a_n2650_13878.t26 gnd 0.702438f
C913 a_n2650_13878.t46 gnd 0.702438f
C914 a_n2650_13878.t40 gnd 0.702438f
C915 a_n2650_13878.n79 gnd 0.308821f
C916 a_n2650_13878.t98 gnd 0.702438f
C917 a_n2650_13878.t77 gnd 0.702438f
C918 a_n2650_13878.t82 gnd 0.702438f
C919 a_n2650_13878.n80 gnd 0.308697f
C920 a_n2650_13878.t71 gnd 0.702438f
C921 a_n2650_13878.t87 gnd 0.702438f
C922 a_n2650_13878.t95 gnd 0.702438f
C923 a_n2650_13878.n81 gnd 0.304914f
C924 a_n2650_13878.t96 gnd 0.702438f
C925 a_n2650_13878.t66 gnd 0.702438f
C926 a_n2650_13878.t79 gnd 0.702438f
C927 a_n2650_13878.n82 gnd 0.308821f
C928 a_n2650_13878.t69 gnd 0.714208f
C929 a_n2650_13878.n83 gnd 0.305176f
C930 a_n2650_13878.n84 gnd 0.299545f
C931 a_n2650_13878.n85 gnd 0.308836f
C932 a_n2650_13878.n86 gnd 0.311475f
C933 a_n2650_13878.n87 gnd 0.304579f
C934 a_n2650_13878.n88 gnd 0.299377f
C935 a_n2650_13878.t42 gnd 0.714208f
C936 a_n2650_13878.t0 gnd 0.117454f
C937 a_n2650_13878.t62 gnd 0.117454f
C938 a_n2650_13878.n89 gnd 1.03952f
C939 a_n2650_13878.t50 gnd 0.117454f
C940 a_n2650_13878.t53 gnd 0.117454f
C941 a_n2650_13878.n90 gnd 1.03787f
C942 a_n2650_13878.t56 gnd 0.117454f
C943 a_n2650_13878.t7 gnd 0.117454f
C944 a_n2650_13878.n91 gnd 1.03787f
C945 a_n2650_13878.t60 gnd 0.117454f
C946 a_n2650_13878.t48 gnd 0.117454f
C947 a_n2650_13878.n92 gnd 1.03952f
C948 a_n2650_13878.t51 gnd 0.117454f
C949 a_n2650_13878.t61 gnd 0.117454f
C950 a_n2650_13878.n93 gnd 1.03787f
C951 a_n2650_13878.t5 gnd 0.117454f
C952 a_n2650_13878.t57 gnd 0.117454f
C953 a_n2650_13878.n94 gnd 1.03787f
C954 a_n2650_13878.t2 gnd 0.117454f
C955 a_n2650_13878.t6 gnd 0.117454f
C956 a_n2650_13878.n95 gnd 1.03787f
C957 a_n2650_13878.t49 gnd 0.117454f
C958 a_n2650_13878.t63 gnd 0.117454f
C959 a_n2650_13878.n96 gnd 1.03787f
C960 a_n2650_13878.t58 gnd 0.117454f
C961 a_n2650_13878.t54 gnd 0.117454f
C962 a_n2650_13878.n97 gnd 1.03787f
C963 a_n2650_13878.t55 gnd 0.117454f
C964 a_n2650_13878.t59 gnd 0.117454f
C965 a_n2650_13878.n98 gnd 1.03952f
C966 a_n2650_13878.t3 gnd 0.117454f
C967 a_n2650_13878.t52 gnd 0.117454f
C968 a_n2650_13878.n99 gnd 1.03787f
C969 a_n2650_13878.t1 gnd 0.117454f
C970 a_n2650_13878.t4 gnd 0.117454f
C971 a_n2650_13878.n100 gnd 1.03787f
C972 a_n2650_13878.n101 gnd 0.305176f
C973 a_n2650_13878.n102 gnd 0.299545f
C974 a_n2650_13878.n103 gnd 0.308836f
C975 a_n2650_13878.n104 gnd 0.311475f
C976 a_n2650_13878.n105 gnd 0.304579f
C977 a_n2650_13878.n106 gnd 0.299377f
C978 a_n2650_13878.t43 gnd 1.41401f
C979 a_n2650_13878.t47 gnd 0.151013f
C980 a_n2650_13878.t41 gnd 0.151013f
C981 a_n2650_13878.n107 gnd 1.06373f
C982 a_n2650_13878.t17 gnd 0.151013f
C983 a_n2650_13878.t27 gnd 0.151013f
C984 a_n2650_13878.n108 gnd 1.06373f
C985 a_n2650_13878.t37 gnd 0.151013f
C986 a_n2650_13878.t39 gnd 0.151013f
C987 a_n2650_13878.n109 gnd 1.06373f
C988 a_n2650_13878.t13 gnd 0.151013f
C989 a_n2650_13878.t29 gnd 0.151013f
C990 a_n2650_13878.n110 gnd 1.06373f
C991 a_n2650_13878.t45 gnd 1.41119f
C992 a_n2650_13878.n111 gnd 1.45813f
C993 a_n2650_13878.n112 gnd 0.949282f
C994 a_n2650_13878.t75 gnd 0.702438f
C995 a_n2650_13878.t85 gnd 0.702438f
C996 a_n2650_13878.t99 gnd 0.702438f
C997 a_n2650_13878.n113 gnd 0.308836f
C998 a_n2650_13878.t88 gnd 0.702438f
C999 a_n2650_13878.t72 gnd 0.702438f
C1000 a_n2650_13878.t73 gnd 0.702438f
C1001 a_n2650_13878.n114 gnd 0.308836f
C1002 a_n2650_13878.t92 gnd 0.702438f
C1003 a_n2650_13878.t81 gnd 0.702438f
C1004 a_n2650_13878.t80 gnd 0.702438f
C1005 a_n2650_13878.n115 gnd 0.308836f
C1006 a_n2650_13878.t84 gnd 0.702438f
C1007 a_n2650_13878.t74 gnd 0.702438f
C1008 a_n2650_13878.t64 gnd 0.702438f
C1009 a_n2650_13878.n116 gnd 0.308836f
C1010 a_n2650_13878.t89 gnd 0.714208f
C1011 a_n2650_13878.n117 gnd 0.304914f
C1012 a_n2650_13878.n118 gnd 0.299377f
C1013 a_n2650_13878.t97 gnd 0.714208f
C1014 a_n2650_13878.n119 gnd 0.304914f
C1015 a_n2650_13878.n120 gnd 0.299377f
C1016 a_n2650_13878.t83 gnd 0.714208f
C1017 a_n2650_13878.n121 gnd 0.304914f
C1018 a_n2650_13878.n122 gnd 0.299377f
C1019 a_n2650_13878.t78 gnd 0.714208f
C1020 a_n2650_13878.n123 gnd 0.304914f
C1021 a_n2650_13878.n124 gnd 0.299377f
C1022 a_n2650_13878.n125 gnd 1.25084f
C1023 a_n2650_13878.n126 gnd 0.299377f
C1024 a_n2650_13878.t93 gnd 0.702438f
C1025 a_n2650_13878.n127 gnd 0.304579f
C1026 a_n2650_13878.t68 gnd 0.702438f
C1027 a_n2650_13878.n128 gnd 0.311475f
C1028 a_n2650_13878.t90 gnd 0.702438f
C1029 a_n2650_13878.n129 gnd 0.308836f
C1030 a_n2650_13878.n130 gnd 0.304914f
C1031 a_n2650_13878.t65 gnd 0.702438f
C1032 a_n2650_13878.n131 gnd 0.299545f
C1033 a_n2650_13878.t86 gnd 0.702438f
C1034 a_n2650_13878.n132 gnd 0.308821f
C1035 a_n2650_13878.t67 gnd 0.714208f
C1036 a_n2650_13878.n133 gnd 0.299377f
C1037 a_n2650_13878.t34 gnd 0.702438f
C1038 a_n2650_13878.n134 gnd 0.304579f
C1039 a_n2650_13878.t22 gnd 0.702438f
C1040 a_n2650_13878.n135 gnd 0.311475f
C1041 a_n2650_13878.t14 gnd 0.702438f
C1042 a_n2650_13878.n136 gnd 0.308836f
C1043 a_n2650_13878.n137 gnd 0.304914f
C1044 a_n2650_13878.t24 gnd 0.702438f
C1045 a_n2650_13878.n138 gnd 0.299545f
C1046 a_n2650_13878.t10 gnd 0.702438f
C1047 a_n2650_13878.n139 gnd 0.308821f
C1048 a_n2650_13878.t20 gnd 0.714208f
C1049 a_n2650_13878.n140 gnd 1.28381f
C1050 a_n2650_13878.t21 gnd 1.41119f
C1051 a_n2650_13878.t19 gnd 0.151013f
C1052 a_n2650_13878.t11 gnd 0.151013f
C1053 a_n2650_13878.n141 gnd 1.06373f
C1054 a_n2650_13878.n142 gnd 1.06374f
C1055 a_n2650_13878.t9 gnd 0.151013f
C1056 vdd.t3 gnd 0.038016f
C1057 vdd.t50 gnd 0.038016f
C1058 vdd.n0 gnd 0.299836f
C1059 vdd.t13 gnd 0.038016f
C1060 vdd.t38 gnd 0.038016f
C1061 vdd.n1 gnd 0.299341f
C1062 vdd.n2 gnd 0.27605f
C1063 vdd.t301 gnd 0.038016f
C1064 vdd.t295 gnd 0.038016f
C1065 vdd.n3 gnd 0.299341f
C1066 vdd.n4 gnd 0.139609f
C1067 vdd.t297 gnd 0.038016f
C1068 vdd.t44 gnd 0.038016f
C1069 vdd.n5 gnd 0.299341f
C1070 vdd.n6 gnd 0.130997f
C1071 vdd.t15 gnd 0.038016f
C1072 vdd.t303 gnd 0.038016f
C1073 vdd.n7 gnd 0.299836f
C1074 vdd.t48 gnd 0.038016f
C1075 vdd.t1 gnd 0.038016f
C1076 vdd.n8 gnd 0.299341f
C1077 vdd.n9 gnd 0.27605f
C1078 vdd.t52 gnd 0.038016f
C1079 vdd.t41 gnd 0.038016f
C1080 vdd.n10 gnd 0.299341f
C1081 vdd.n11 gnd 0.139609f
C1082 vdd.t299 gnd 0.038016f
C1083 vdd.t54 gnd 0.038016f
C1084 vdd.n12 gnd 0.299341f
C1085 vdd.n13 gnd 0.130997f
C1086 vdd.n14 gnd 0.092612f
C1087 vdd.t21 gnd 0.02112f
C1088 vdd.t24 gnd 0.02112f
C1089 vdd.n15 gnd 0.194399f
C1090 vdd.t25 gnd 0.02112f
C1091 vdd.t32 gnd 0.02112f
C1092 vdd.n16 gnd 0.19383f
C1093 vdd.n17 gnd 0.337325f
C1094 vdd.t28 gnd 0.02112f
C1095 vdd.t35 gnd 0.02112f
C1096 vdd.n18 gnd 0.19383f
C1097 vdd.n19 gnd 0.139556f
C1098 vdd.t22 gnd 0.02112f
C1099 vdd.t23 gnd 0.02112f
C1100 vdd.n20 gnd 0.194399f
C1101 vdd.t27 gnd 0.02112f
C1102 vdd.t31 gnd 0.02112f
C1103 vdd.n21 gnd 0.19383f
C1104 vdd.n22 gnd 0.337325f
C1105 vdd.t36 gnd 0.02112f
C1106 vdd.t33 gnd 0.02112f
C1107 vdd.n23 gnd 0.19383f
C1108 vdd.n24 gnd 0.139556f
C1109 vdd.t29 gnd 0.02112f
C1110 vdd.t26 gnd 0.02112f
C1111 vdd.n25 gnd 0.19383f
C1112 vdd.t34 gnd 0.02112f
C1113 vdd.t30 gnd 0.02112f
C1114 vdd.n26 gnd 0.19383f
C1115 vdd.n27 gnd 22.3309f
C1116 vdd.n28 gnd 8.566401f
C1117 vdd.n29 gnd 0.00576f
C1118 vdd.n30 gnd 0.005345f
C1119 vdd.n31 gnd 0.002957f
C1120 vdd.n32 gnd 0.006789f
C1121 vdd.n33 gnd 0.002872f
C1122 vdd.n34 gnd 0.003041f
C1123 vdd.n35 gnd 0.005345f
C1124 vdd.n36 gnd 0.002872f
C1125 vdd.n37 gnd 0.006789f
C1126 vdd.n38 gnd 0.003041f
C1127 vdd.n39 gnd 0.005345f
C1128 vdd.n40 gnd 0.002872f
C1129 vdd.n41 gnd 0.005092f
C1130 vdd.n42 gnd 0.005107f
C1131 vdd.t262 gnd 0.014586f
C1132 vdd.n43 gnd 0.032453f
C1133 vdd.n44 gnd 0.168893f
C1134 vdd.n45 gnd 0.002872f
C1135 vdd.n46 gnd 0.003041f
C1136 vdd.n47 gnd 0.006789f
C1137 vdd.n48 gnd 0.006789f
C1138 vdd.n49 gnd 0.003041f
C1139 vdd.n50 gnd 0.002872f
C1140 vdd.n51 gnd 0.005345f
C1141 vdd.n52 gnd 0.005345f
C1142 vdd.n53 gnd 0.002872f
C1143 vdd.n54 gnd 0.003041f
C1144 vdd.n55 gnd 0.006789f
C1145 vdd.n56 gnd 0.006789f
C1146 vdd.n57 gnd 0.003041f
C1147 vdd.n58 gnd 0.002872f
C1148 vdd.n59 gnd 0.005345f
C1149 vdd.n60 gnd 0.005345f
C1150 vdd.n61 gnd 0.002872f
C1151 vdd.n62 gnd 0.003041f
C1152 vdd.n63 gnd 0.006789f
C1153 vdd.n64 gnd 0.006789f
C1154 vdd.n65 gnd 0.016051f
C1155 vdd.n66 gnd 0.002957f
C1156 vdd.n67 gnd 0.002872f
C1157 vdd.n68 gnd 0.013816f
C1158 vdd.n69 gnd 0.009645f
C1159 vdd.t142 gnd 0.033792f
C1160 vdd.t194 gnd 0.033792f
C1161 vdd.n70 gnd 0.23224f
C1162 vdd.n71 gnd 0.182621f
C1163 vdd.t156 gnd 0.033792f
C1164 vdd.t220 gnd 0.033792f
C1165 vdd.n72 gnd 0.23224f
C1166 vdd.n73 gnd 0.147374f
C1167 vdd.t185 gnd 0.033792f
C1168 vdd.t268 gnd 0.033792f
C1169 vdd.n74 gnd 0.23224f
C1170 vdd.n75 gnd 0.147374f
C1171 vdd.t161 gnd 0.033792f
C1172 vdd.t249 gnd 0.033792f
C1173 vdd.n76 gnd 0.23224f
C1174 vdd.n77 gnd 0.147374f
C1175 vdd.t166 gnd 0.033792f
C1176 vdd.t264 gnd 0.033792f
C1177 vdd.n78 gnd 0.23224f
C1178 vdd.n79 gnd 0.147374f
C1179 vdd.t203 gnd 0.033792f
C1180 vdd.t278 gnd 0.033792f
C1181 vdd.n80 gnd 0.23224f
C1182 vdd.n81 gnd 0.147374f
C1183 vdd.t223 gnd 0.033792f
C1184 vdd.t255 gnd 0.033792f
C1185 vdd.n82 gnd 0.23224f
C1186 vdd.n83 gnd 0.147374f
C1187 vdd.t188 gnd 0.033792f
C1188 vdd.t270 gnd 0.033792f
C1189 vdd.n84 gnd 0.23224f
C1190 vdd.n85 gnd 0.147374f
C1191 vdd.t212 gnd 0.033792f
C1192 vdd.t286 gnd 0.033792f
C1193 vdd.n86 gnd 0.23224f
C1194 vdd.n87 gnd 0.147374f
C1195 vdd.n88 gnd 0.00576f
C1196 vdd.n89 gnd 0.005345f
C1197 vdd.n90 gnd 0.002957f
C1198 vdd.n91 gnd 0.006789f
C1199 vdd.n92 gnd 0.002872f
C1200 vdd.n93 gnd 0.003041f
C1201 vdd.n94 gnd 0.005345f
C1202 vdd.n95 gnd 0.002872f
C1203 vdd.n96 gnd 0.006789f
C1204 vdd.n97 gnd 0.003041f
C1205 vdd.n98 gnd 0.005345f
C1206 vdd.n99 gnd 0.002872f
C1207 vdd.n100 gnd 0.005092f
C1208 vdd.n101 gnd 0.005107f
C1209 vdd.t236 gnd 0.014586f
C1210 vdd.n102 gnd 0.032453f
C1211 vdd.n103 gnd 0.168893f
C1212 vdd.n104 gnd 0.002872f
C1213 vdd.n105 gnd 0.003041f
C1214 vdd.n106 gnd 0.006789f
C1215 vdd.n107 gnd 0.006789f
C1216 vdd.n108 gnd 0.003041f
C1217 vdd.n109 gnd 0.002872f
C1218 vdd.n110 gnd 0.005345f
C1219 vdd.n111 gnd 0.005345f
C1220 vdd.n112 gnd 0.002872f
C1221 vdd.n113 gnd 0.003041f
C1222 vdd.n114 gnd 0.006789f
C1223 vdd.n115 gnd 0.006789f
C1224 vdd.n116 gnd 0.003041f
C1225 vdd.n117 gnd 0.002872f
C1226 vdd.n118 gnd 0.005345f
C1227 vdd.n119 gnd 0.005345f
C1228 vdd.n120 gnd 0.002872f
C1229 vdd.n121 gnd 0.003041f
C1230 vdd.n122 gnd 0.006789f
C1231 vdd.n123 gnd 0.006789f
C1232 vdd.n124 gnd 0.016051f
C1233 vdd.n125 gnd 0.002957f
C1234 vdd.n126 gnd 0.002872f
C1235 vdd.n127 gnd 0.013816f
C1236 vdd.n128 gnd 0.009343f
C1237 vdd.n129 gnd 0.109647f
C1238 vdd.n130 gnd 0.00576f
C1239 vdd.n131 gnd 0.005345f
C1240 vdd.n132 gnd 0.002957f
C1241 vdd.n133 gnd 0.006789f
C1242 vdd.n134 gnd 0.002872f
C1243 vdd.n135 gnd 0.003041f
C1244 vdd.n136 gnd 0.005345f
C1245 vdd.n137 gnd 0.002872f
C1246 vdd.n138 gnd 0.006789f
C1247 vdd.n139 gnd 0.003041f
C1248 vdd.n140 gnd 0.005345f
C1249 vdd.n141 gnd 0.002872f
C1250 vdd.n142 gnd 0.005092f
C1251 vdd.n143 gnd 0.005107f
C1252 vdd.t193 gnd 0.014586f
C1253 vdd.n144 gnd 0.032453f
C1254 vdd.n145 gnd 0.168893f
C1255 vdd.n146 gnd 0.002872f
C1256 vdd.n147 gnd 0.003041f
C1257 vdd.n148 gnd 0.006789f
C1258 vdd.n149 gnd 0.006789f
C1259 vdd.n150 gnd 0.003041f
C1260 vdd.n151 gnd 0.002872f
C1261 vdd.n152 gnd 0.005345f
C1262 vdd.n153 gnd 0.005345f
C1263 vdd.n154 gnd 0.002872f
C1264 vdd.n155 gnd 0.003041f
C1265 vdd.n156 gnd 0.006789f
C1266 vdd.n157 gnd 0.006789f
C1267 vdd.n158 gnd 0.003041f
C1268 vdd.n159 gnd 0.002872f
C1269 vdd.n160 gnd 0.005345f
C1270 vdd.n161 gnd 0.005345f
C1271 vdd.n162 gnd 0.002872f
C1272 vdd.n163 gnd 0.003041f
C1273 vdd.n164 gnd 0.006789f
C1274 vdd.n165 gnd 0.006789f
C1275 vdd.n166 gnd 0.016051f
C1276 vdd.n167 gnd 0.002957f
C1277 vdd.n168 gnd 0.002872f
C1278 vdd.n169 gnd 0.013816f
C1279 vdd.n170 gnd 0.009645f
C1280 vdd.t277 gnd 0.033792f
C1281 vdd.t180 gnd 0.033792f
C1282 vdd.n171 gnd 0.23224f
C1283 vdd.n172 gnd 0.182621f
C1284 vdd.t183 gnd 0.033792f
C1285 vdd.t274 gnd 0.033792f
C1286 vdd.n173 gnd 0.23224f
C1287 vdd.n174 gnd 0.147374f
C1288 vdd.t275 gnd 0.033792f
C1289 vdd.t154 gnd 0.033792f
C1290 vdd.n175 gnd 0.23224f
C1291 vdd.n176 gnd 0.147374f
C1292 vdd.t257 gnd 0.033792f
C1293 vdd.t267 gnd 0.033792f
C1294 vdd.n177 gnd 0.23224f
C1295 vdd.n178 gnd 0.147374f
C1296 vdd.t148 gnd 0.033792f
C1297 vdd.t218 gnd 0.033792f
C1298 vdd.n179 gnd 0.23224f
C1299 vdd.n180 gnd 0.147374f
C1300 vdd.t254 gnd 0.033792f
C1301 vdd.t282 gnd 0.033792f
C1302 vdd.n181 gnd 0.23224f
C1303 vdd.n182 gnd 0.147374f
C1304 vdd.t191 gnd 0.033792f
C1305 vdd.t253 gnd 0.033792f
C1306 vdd.n183 gnd 0.23224f
C1307 vdd.n184 gnd 0.147374f
C1308 vdd.t290 gnd 0.033792f
C1309 vdd.t182 gnd 0.033792f
C1310 vdd.n185 gnd 0.23224f
C1311 vdd.n186 gnd 0.147374f
C1312 vdd.t235 gnd 0.033792f
C1313 vdd.t273 gnd 0.033792f
C1314 vdd.n187 gnd 0.23224f
C1315 vdd.n188 gnd 0.147374f
C1316 vdd.n189 gnd 0.00576f
C1317 vdd.n190 gnd 0.005345f
C1318 vdd.n191 gnd 0.002957f
C1319 vdd.n192 gnd 0.006789f
C1320 vdd.n193 gnd 0.002872f
C1321 vdd.n194 gnd 0.003041f
C1322 vdd.n195 gnd 0.005345f
C1323 vdd.n196 gnd 0.002872f
C1324 vdd.n197 gnd 0.006789f
C1325 vdd.n198 gnd 0.003041f
C1326 vdd.n199 gnd 0.005345f
C1327 vdd.n200 gnd 0.002872f
C1328 vdd.n201 gnd 0.005092f
C1329 vdd.n202 gnd 0.005107f
C1330 vdd.t152 gnd 0.014586f
C1331 vdd.n203 gnd 0.032453f
C1332 vdd.n204 gnd 0.168893f
C1333 vdd.n205 gnd 0.002872f
C1334 vdd.n206 gnd 0.003041f
C1335 vdd.n207 gnd 0.006789f
C1336 vdd.n208 gnd 0.006789f
C1337 vdd.n209 gnd 0.003041f
C1338 vdd.n210 gnd 0.002872f
C1339 vdd.n211 gnd 0.005345f
C1340 vdd.n212 gnd 0.005345f
C1341 vdd.n213 gnd 0.002872f
C1342 vdd.n214 gnd 0.003041f
C1343 vdd.n215 gnd 0.006789f
C1344 vdd.n216 gnd 0.006789f
C1345 vdd.n217 gnd 0.003041f
C1346 vdd.n218 gnd 0.002872f
C1347 vdd.n219 gnd 0.005345f
C1348 vdd.n220 gnd 0.005345f
C1349 vdd.n221 gnd 0.002872f
C1350 vdd.n222 gnd 0.003041f
C1351 vdd.n223 gnd 0.006789f
C1352 vdd.n224 gnd 0.006789f
C1353 vdd.n225 gnd 0.016051f
C1354 vdd.n226 gnd 0.002957f
C1355 vdd.n227 gnd 0.002872f
C1356 vdd.n228 gnd 0.013816f
C1357 vdd.n229 gnd 0.009343f
C1358 vdd.n230 gnd 0.065229f
C1359 vdd.n231 gnd 0.235038f
C1360 vdd.n232 gnd 0.00576f
C1361 vdd.n233 gnd 0.005345f
C1362 vdd.n234 gnd 0.002957f
C1363 vdd.n235 gnd 0.006789f
C1364 vdd.n236 gnd 0.002872f
C1365 vdd.n237 gnd 0.003041f
C1366 vdd.n238 gnd 0.005345f
C1367 vdd.n239 gnd 0.002872f
C1368 vdd.n240 gnd 0.006789f
C1369 vdd.n241 gnd 0.003041f
C1370 vdd.n242 gnd 0.005345f
C1371 vdd.n243 gnd 0.002872f
C1372 vdd.n244 gnd 0.005092f
C1373 vdd.n245 gnd 0.005107f
C1374 vdd.t213 gnd 0.014586f
C1375 vdd.n246 gnd 0.032453f
C1376 vdd.n247 gnd 0.168893f
C1377 vdd.n248 gnd 0.002872f
C1378 vdd.n249 gnd 0.003041f
C1379 vdd.n250 gnd 0.006789f
C1380 vdd.n251 gnd 0.006789f
C1381 vdd.n252 gnd 0.003041f
C1382 vdd.n253 gnd 0.002872f
C1383 vdd.n254 gnd 0.005345f
C1384 vdd.n255 gnd 0.005345f
C1385 vdd.n256 gnd 0.002872f
C1386 vdd.n257 gnd 0.003041f
C1387 vdd.n258 gnd 0.006789f
C1388 vdd.n259 gnd 0.006789f
C1389 vdd.n260 gnd 0.003041f
C1390 vdd.n261 gnd 0.002872f
C1391 vdd.n262 gnd 0.005345f
C1392 vdd.n263 gnd 0.005345f
C1393 vdd.n264 gnd 0.002872f
C1394 vdd.n265 gnd 0.003041f
C1395 vdd.n266 gnd 0.006789f
C1396 vdd.n267 gnd 0.006789f
C1397 vdd.n268 gnd 0.016051f
C1398 vdd.n269 gnd 0.002957f
C1399 vdd.n270 gnd 0.002872f
C1400 vdd.n271 gnd 0.013816f
C1401 vdd.n272 gnd 0.009645f
C1402 vdd.t289 gnd 0.033792f
C1403 vdd.t206 gnd 0.033792f
C1404 vdd.n273 gnd 0.23224f
C1405 vdd.n274 gnd 0.182621f
C1406 vdd.t208 gnd 0.033792f
C1407 vdd.t283 gnd 0.033792f
C1408 vdd.n275 gnd 0.23224f
C1409 vdd.n276 gnd 0.147374f
C1410 vdd.t285 gnd 0.033792f
C1411 vdd.t177 gnd 0.033792f
C1412 vdd.n277 gnd 0.23224f
C1413 vdd.n278 gnd 0.147374f
C1414 vdd.t266 gnd 0.033792f
C1415 vdd.t281 gnd 0.033792f
C1416 vdd.n279 gnd 0.23224f
C1417 vdd.n280 gnd 0.147374f
C1418 vdd.t167 gnd 0.033792f
C1419 vdd.t237 gnd 0.033792f
C1420 vdd.n281 gnd 0.23224f
C1421 vdd.n282 gnd 0.147374f
C1422 vdd.t265 gnd 0.033792f
C1423 vdd.t138 gnd 0.033792f
C1424 vdd.n283 gnd 0.23224f
C1425 vdd.n284 gnd 0.147374f
C1426 vdd.t210 gnd 0.033792f
C1427 vdd.t263 gnd 0.033792f
C1428 vdd.n285 gnd 0.23224f
C1429 vdd.n286 gnd 0.147374f
C1430 vdd.t150 gnd 0.033792f
C1431 vdd.t207 gnd 0.033792f
C1432 vdd.n287 gnd 0.23224f
C1433 vdd.n288 gnd 0.147374f
C1434 vdd.t243 gnd 0.033792f
C1435 vdd.t284 gnd 0.033792f
C1436 vdd.n289 gnd 0.23224f
C1437 vdd.n290 gnd 0.147374f
C1438 vdd.n291 gnd 0.00576f
C1439 vdd.n292 gnd 0.005345f
C1440 vdd.n293 gnd 0.002957f
C1441 vdd.n294 gnd 0.006789f
C1442 vdd.n295 gnd 0.002872f
C1443 vdd.n296 gnd 0.003041f
C1444 vdd.n297 gnd 0.005345f
C1445 vdd.n298 gnd 0.002872f
C1446 vdd.n299 gnd 0.006789f
C1447 vdd.n300 gnd 0.003041f
C1448 vdd.n301 gnd 0.005345f
C1449 vdd.n302 gnd 0.002872f
C1450 vdd.n303 gnd 0.005092f
C1451 vdd.n304 gnd 0.005107f
C1452 vdd.t172 gnd 0.014586f
C1453 vdd.n305 gnd 0.032453f
C1454 vdd.n306 gnd 0.168893f
C1455 vdd.n307 gnd 0.002872f
C1456 vdd.n308 gnd 0.003041f
C1457 vdd.n309 gnd 0.006789f
C1458 vdd.n310 gnd 0.006789f
C1459 vdd.n311 gnd 0.003041f
C1460 vdd.n312 gnd 0.002872f
C1461 vdd.n313 gnd 0.005345f
C1462 vdd.n314 gnd 0.005345f
C1463 vdd.n315 gnd 0.002872f
C1464 vdd.n316 gnd 0.003041f
C1465 vdd.n317 gnd 0.006789f
C1466 vdd.n318 gnd 0.006789f
C1467 vdd.n319 gnd 0.003041f
C1468 vdd.n320 gnd 0.002872f
C1469 vdd.n321 gnd 0.005345f
C1470 vdd.n322 gnd 0.005345f
C1471 vdd.n323 gnd 0.002872f
C1472 vdd.n324 gnd 0.003041f
C1473 vdd.n325 gnd 0.006789f
C1474 vdd.n326 gnd 0.006789f
C1475 vdd.n327 gnd 0.016051f
C1476 vdd.n328 gnd 0.002957f
C1477 vdd.n329 gnd 0.002872f
C1478 vdd.n330 gnd 0.013816f
C1479 vdd.n331 gnd 0.009343f
C1480 vdd.n332 gnd 0.065229f
C1481 vdd.n333 gnd 0.269067f
C1482 vdd.n334 gnd 0.008067f
C1483 vdd.n335 gnd 0.010496f
C1484 vdd.n336 gnd 0.008448f
C1485 vdd.n337 gnd 0.008448f
C1486 vdd.n338 gnd 0.010496f
C1487 vdd.n339 gnd 0.010496f
C1488 vdd.n340 gnd 0.766932f
C1489 vdd.n341 gnd 0.010496f
C1490 vdd.n342 gnd 0.010496f
C1491 vdd.n343 gnd 0.010496f
C1492 vdd.n344 gnd 0.83129f
C1493 vdd.n345 gnd 0.010496f
C1494 vdd.n346 gnd 0.010496f
C1495 vdd.n347 gnd 0.010496f
C1496 vdd.n348 gnd 0.010496f
C1497 vdd.n349 gnd 0.008448f
C1498 vdd.n350 gnd 0.010496f
C1499 vdd.t137 gnd 0.536316f
C1500 vdd.n351 gnd 0.010496f
C1501 vdd.n352 gnd 0.010496f
C1502 vdd.n353 gnd 0.010496f
C1503 vdd.t252 gnd 0.536316f
C1504 vdd.n354 gnd 0.010496f
C1505 vdd.n355 gnd 0.010496f
C1506 vdd.n356 gnd 0.010496f
C1507 vdd.n357 gnd 0.010496f
C1508 vdd.n358 gnd 0.010496f
C1509 vdd.n359 gnd 0.008448f
C1510 vdd.n360 gnd 0.010496f
C1511 vdd.n361 gnd 0.606037f
C1512 vdd.n362 gnd 0.010496f
C1513 vdd.n363 gnd 0.010496f
C1514 vdd.n364 gnd 0.010496f
C1515 vdd.t181 gnd 0.536316f
C1516 vdd.n365 gnd 0.010496f
C1517 vdd.n366 gnd 0.010496f
C1518 vdd.n367 gnd 0.010496f
C1519 vdd.n368 gnd 0.010496f
C1520 vdd.n369 gnd 0.010496f
C1521 vdd.n370 gnd 0.008448f
C1522 vdd.n371 gnd 0.010496f
C1523 vdd.t211 gnd 0.536316f
C1524 vdd.n372 gnd 0.010496f
C1525 vdd.n373 gnd 0.010496f
C1526 vdd.n374 gnd 0.010496f
C1527 vdd.n375 gnd 0.62749f
C1528 vdd.n376 gnd 0.010496f
C1529 vdd.n377 gnd 0.010496f
C1530 vdd.n378 gnd 0.010496f
C1531 vdd.n379 gnd 0.010496f
C1532 vdd.n380 gnd 0.010496f
C1533 vdd.n381 gnd 0.008448f
C1534 vdd.n382 gnd 0.010496f
C1535 vdd.t151 gnd 0.536316f
C1536 vdd.n383 gnd 0.010496f
C1537 vdd.n384 gnd 0.010496f
C1538 vdd.n385 gnd 0.010496f
C1539 vdd.n386 gnd 0.541679f
C1540 vdd.n387 gnd 0.010496f
C1541 vdd.n388 gnd 0.010496f
C1542 vdd.n389 gnd 0.010496f
C1543 vdd.n390 gnd 0.010496f
C1544 vdd.n391 gnd 0.02539f
C1545 vdd.n392 gnd 0.025935f
C1546 vdd.t70 gnd 0.536316f
C1547 vdd.n393 gnd 0.02539f
C1548 vdd.n425 gnd 0.010496f
C1549 vdd.t98 gnd 0.129127f
C1550 vdd.t97 gnd 0.138001f
C1551 vdd.t96 gnd 0.168639f
C1552 vdd.n426 gnd 0.216171f
C1553 vdd.n427 gnd 0.182467f
C1554 vdd.n428 gnd 0.013855f
C1555 vdd.n429 gnd 0.010496f
C1556 vdd.n430 gnd 0.008448f
C1557 vdd.n431 gnd 0.010496f
C1558 vdd.n432 gnd 0.008448f
C1559 vdd.n433 gnd 0.010496f
C1560 vdd.n434 gnd 0.008448f
C1561 vdd.n435 gnd 0.010496f
C1562 vdd.n436 gnd 0.008448f
C1563 vdd.n437 gnd 0.010496f
C1564 vdd.n438 gnd 0.008448f
C1565 vdd.n439 gnd 0.010496f
C1566 vdd.t72 gnd 0.129127f
C1567 vdd.t71 gnd 0.138001f
C1568 vdd.t69 gnd 0.168639f
C1569 vdd.n440 gnd 0.216171f
C1570 vdd.n441 gnd 0.182467f
C1571 vdd.n442 gnd 0.008448f
C1572 vdd.n443 gnd 0.010496f
C1573 vdd.n444 gnd 0.008448f
C1574 vdd.n445 gnd 0.010496f
C1575 vdd.n446 gnd 0.008448f
C1576 vdd.n447 gnd 0.010496f
C1577 vdd.n448 gnd 0.008448f
C1578 vdd.n449 gnd 0.010496f
C1579 vdd.n450 gnd 0.008448f
C1580 vdd.n451 gnd 0.010496f
C1581 vdd.t89 gnd 0.129127f
C1582 vdd.t88 gnd 0.138001f
C1583 vdd.t87 gnd 0.168639f
C1584 vdd.n452 gnd 0.216171f
C1585 vdd.n453 gnd 0.182467f
C1586 vdd.n454 gnd 0.018079f
C1587 vdd.n455 gnd 0.010496f
C1588 vdd.n456 gnd 0.008448f
C1589 vdd.n457 gnd 0.010496f
C1590 vdd.n458 gnd 0.008448f
C1591 vdd.n459 gnd 0.010496f
C1592 vdd.n460 gnd 0.008448f
C1593 vdd.n461 gnd 0.010496f
C1594 vdd.n462 gnd 0.008448f
C1595 vdd.n463 gnd 0.010496f
C1596 vdd.n464 gnd 0.025935f
C1597 vdd.n465 gnd 0.007012f
C1598 vdd.n466 gnd 0.008448f
C1599 vdd.n467 gnd 0.010496f
C1600 vdd.n468 gnd 0.010496f
C1601 vdd.n469 gnd 0.008448f
C1602 vdd.n470 gnd 0.010496f
C1603 vdd.n471 gnd 0.010496f
C1604 vdd.n472 gnd 0.010496f
C1605 vdd.n473 gnd 0.010496f
C1606 vdd.n474 gnd 0.010496f
C1607 vdd.n475 gnd 0.008448f
C1608 vdd.n476 gnd 0.008448f
C1609 vdd.n477 gnd 0.010496f
C1610 vdd.n478 gnd 0.010496f
C1611 vdd.n479 gnd 0.008448f
C1612 vdd.n480 gnd 0.010496f
C1613 vdd.n481 gnd 0.010496f
C1614 vdd.n482 gnd 0.010496f
C1615 vdd.n483 gnd 0.010496f
C1616 vdd.n484 gnd 0.010496f
C1617 vdd.n485 gnd 0.008448f
C1618 vdd.n486 gnd 0.008448f
C1619 vdd.n487 gnd 0.010496f
C1620 vdd.n488 gnd 0.010496f
C1621 vdd.n489 gnd 0.008448f
C1622 vdd.n490 gnd 0.010496f
C1623 vdd.n491 gnd 0.010496f
C1624 vdd.n492 gnd 0.010496f
C1625 vdd.n493 gnd 0.010496f
C1626 vdd.n494 gnd 0.010496f
C1627 vdd.n495 gnd 0.008448f
C1628 vdd.n496 gnd 0.008448f
C1629 vdd.n497 gnd 0.010496f
C1630 vdd.n498 gnd 0.010496f
C1631 vdd.n499 gnd 0.008448f
C1632 vdd.n500 gnd 0.010496f
C1633 vdd.n501 gnd 0.010496f
C1634 vdd.n502 gnd 0.010496f
C1635 vdd.n503 gnd 0.010496f
C1636 vdd.n504 gnd 0.010496f
C1637 vdd.n505 gnd 0.008448f
C1638 vdd.n506 gnd 0.008448f
C1639 vdd.n507 gnd 0.010496f
C1640 vdd.n508 gnd 0.010496f
C1641 vdd.n509 gnd 0.007054f
C1642 vdd.n510 gnd 0.010496f
C1643 vdd.n511 gnd 0.010496f
C1644 vdd.n512 gnd 0.010496f
C1645 vdd.n513 gnd 0.010496f
C1646 vdd.n514 gnd 0.010496f
C1647 vdd.n515 gnd 0.007054f
C1648 vdd.n516 gnd 0.008448f
C1649 vdd.n517 gnd 0.010496f
C1650 vdd.n518 gnd 0.010496f
C1651 vdd.n519 gnd 0.008448f
C1652 vdd.n520 gnd 0.010496f
C1653 vdd.n521 gnd 0.010496f
C1654 vdd.n522 gnd 0.010496f
C1655 vdd.n523 gnd 0.010496f
C1656 vdd.n524 gnd 0.010496f
C1657 vdd.n525 gnd 0.008448f
C1658 vdd.n526 gnd 0.008448f
C1659 vdd.n527 gnd 0.010496f
C1660 vdd.n528 gnd 0.010496f
C1661 vdd.n529 gnd 0.008448f
C1662 vdd.n530 gnd 0.010496f
C1663 vdd.n531 gnd 0.010496f
C1664 vdd.n532 gnd 0.010496f
C1665 vdd.n533 gnd 0.010496f
C1666 vdd.n534 gnd 0.010496f
C1667 vdd.n535 gnd 0.008448f
C1668 vdd.n536 gnd 0.008448f
C1669 vdd.n537 gnd 0.010496f
C1670 vdd.n538 gnd 0.010496f
C1671 vdd.n539 gnd 0.008448f
C1672 vdd.n540 gnd 0.010496f
C1673 vdd.n541 gnd 0.010496f
C1674 vdd.n542 gnd 0.010496f
C1675 vdd.n543 gnd 0.010496f
C1676 vdd.n544 gnd 0.010496f
C1677 vdd.n545 gnd 0.008448f
C1678 vdd.n546 gnd 0.008448f
C1679 vdd.n547 gnd 0.010496f
C1680 vdd.n548 gnd 0.010496f
C1681 vdd.n549 gnd 0.008448f
C1682 vdd.n550 gnd 0.010496f
C1683 vdd.n551 gnd 0.010496f
C1684 vdd.n552 gnd 0.010496f
C1685 vdd.n553 gnd 0.010496f
C1686 vdd.n554 gnd 0.010496f
C1687 vdd.n555 gnd 0.008448f
C1688 vdd.n556 gnd 0.008448f
C1689 vdd.n557 gnd 0.010496f
C1690 vdd.n558 gnd 0.010496f
C1691 vdd.n559 gnd 0.008448f
C1692 vdd.n560 gnd 0.010496f
C1693 vdd.n561 gnd 0.010496f
C1694 vdd.n562 gnd 0.010496f
C1695 vdd.n563 gnd 0.010496f
C1696 vdd.n564 gnd 0.010496f
C1697 vdd.n565 gnd 0.005745f
C1698 vdd.n566 gnd 0.018079f
C1699 vdd.n567 gnd 0.010496f
C1700 vdd.n568 gnd 0.010496f
C1701 vdd.n569 gnd 0.008363f
C1702 vdd.n570 gnd 0.010496f
C1703 vdd.n571 gnd 0.010496f
C1704 vdd.n572 gnd 0.010496f
C1705 vdd.n573 gnd 0.010496f
C1706 vdd.n574 gnd 0.010496f
C1707 vdd.n575 gnd 0.008448f
C1708 vdd.n576 gnd 0.008448f
C1709 vdd.n577 gnd 0.010496f
C1710 vdd.n578 gnd 0.010496f
C1711 vdd.n579 gnd 0.008448f
C1712 vdd.n580 gnd 0.010496f
C1713 vdd.n581 gnd 0.010496f
C1714 vdd.n582 gnd 0.010496f
C1715 vdd.n583 gnd 0.010496f
C1716 vdd.n584 gnd 0.010496f
C1717 vdd.n585 gnd 0.008448f
C1718 vdd.n586 gnd 0.008448f
C1719 vdd.n587 gnd 0.010496f
C1720 vdd.n588 gnd 0.010496f
C1721 vdd.n589 gnd 0.008448f
C1722 vdd.n590 gnd 0.010496f
C1723 vdd.n591 gnd 0.010496f
C1724 vdd.n592 gnd 0.010496f
C1725 vdd.n593 gnd 0.010496f
C1726 vdd.n594 gnd 0.010496f
C1727 vdd.n595 gnd 0.008448f
C1728 vdd.n596 gnd 0.008448f
C1729 vdd.n597 gnd 0.010496f
C1730 vdd.n598 gnd 0.010496f
C1731 vdd.n599 gnd 0.008448f
C1732 vdd.n600 gnd 0.010496f
C1733 vdd.n601 gnd 0.010496f
C1734 vdd.n602 gnd 0.010496f
C1735 vdd.n603 gnd 0.010496f
C1736 vdd.n604 gnd 0.010496f
C1737 vdd.n605 gnd 0.008448f
C1738 vdd.n606 gnd 0.008448f
C1739 vdd.n607 gnd 0.010496f
C1740 vdd.n608 gnd 0.010496f
C1741 vdd.n609 gnd 0.008448f
C1742 vdd.n610 gnd 0.010496f
C1743 vdd.n611 gnd 0.010496f
C1744 vdd.n612 gnd 0.010496f
C1745 vdd.n613 gnd 0.010496f
C1746 vdd.n614 gnd 0.010496f
C1747 vdd.n615 gnd 0.008448f
C1748 vdd.n616 gnd 0.010496f
C1749 vdd.n617 gnd 0.008448f
C1750 vdd.n618 gnd 0.004435f
C1751 vdd.n619 gnd 0.010496f
C1752 vdd.n620 gnd 0.010496f
C1753 vdd.n621 gnd 0.008448f
C1754 vdd.n622 gnd 0.010496f
C1755 vdd.n623 gnd 0.008448f
C1756 vdd.n624 gnd 0.010496f
C1757 vdd.n625 gnd 0.008448f
C1758 vdd.n626 gnd 0.010496f
C1759 vdd.n627 gnd 0.008448f
C1760 vdd.n628 gnd 0.010496f
C1761 vdd.n629 gnd 0.008448f
C1762 vdd.n630 gnd 0.010496f
C1763 vdd.n631 gnd 0.008448f
C1764 vdd.n632 gnd 0.010496f
C1765 vdd.n633 gnd 0.584585f
C1766 vdd.t147 gnd 0.536316f
C1767 vdd.n634 gnd 0.010496f
C1768 vdd.n635 gnd 0.008448f
C1769 vdd.n636 gnd 0.010496f
C1770 vdd.n637 gnd 0.008448f
C1771 vdd.n638 gnd 0.010496f
C1772 vdd.t160 gnd 0.536316f
C1773 vdd.n639 gnd 0.010496f
C1774 vdd.n640 gnd 0.008448f
C1775 vdd.n641 gnd 0.010496f
C1776 vdd.n642 gnd 0.008448f
C1777 vdd.n643 gnd 0.010496f
C1778 vdd.t153 gnd 0.536316f
C1779 vdd.n644 gnd 0.670395f
C1780 vdd.n645 gnd 0.010496f
C1781 vdd.n646 gnd 0.008448f
C1782 vdd.n647 gnd 0.010496f
C1783 vdd.n648 gnd 0.008448f
C1784 vdd.n649 gnd 0.010496f
C1785 vdd.t184 gnd 0.536316f
C1786 vdd.n650 gnd 0.010496f
C1787 vdd.n651 gnd 0.008448f
C1788 vdd.n652 gnd 0.010496f
C1789 vdd.n653 gnd 0.008448f
C1790 vdd.n654 gnd 0.010496f
C1791 vdd.n655 gnd 0.745479f
C1792 vdd.n656 gnd 0.890285f
C1793 vdd.t219 gnd 0.536316f
C1794 vdd.n657 gnd 0.010496f
C1795 vdd.n658 gnd 0.008448f
C1796 vdd.n659 gnd 0.010496f
C1797 vdd.n660 gnd 0.008448f
C1798 vdd.n661 gnd 0.010496f
C1799 vdd.n662 gnd 0.563132f
C1800 vdd.n663 gnd 0.010496f
C1801 vdd.n664 gnd 0.008448f
C1802 vdd.n665 gnd 0.010496f
C1803 vdd.n666 gnd 0.008448f
C1804 vdd.n667 gnd 0.010496f
C1805 vdd.t141 gnd 0.536316f
C1806 vdd.t179 gnd 0.536316f
C1807 vdd.n668 gnd 0.010496f
C1808 vdd.n669 gnd 0.008448f
C1809 vdd.n670 gnd 0.010496f
C1810 vdd.n671 gnd 0.008448f
C1811 vdd.n672 gnd 0.010496f
C1812 vdd.t192 gnd 0.536316f
C1813 vdd.n673 gnd 0.010496f
C1814 vdd.n674 gnd 0.008448f
C1815 vdd.n675 gnd 0.010496f
C1816 vdd.n676 gnd 0.008448f
C1817 vdd.n677 gnd 0.010496f
C1818 vdd.n678 gnd 1.07263f
C1819 vdd.n679 gnd 0.874195f
C1820 vdd.n680 gnd 0.010496f
C1821 vdd.n681 gnd 0.008448f
C1822 vdd.n682 gnd 0.02539f
C1823 vdd.n683 gnd 0.007012f
C1824 vdd.n684 gnd 0.02539f
C1825 vdd.t58 gnd 0.536316f
C1826 vdd.n685 gnd 0.02539f
C1827 vdd.n686 gnd 0.007012f
C1828 vdd.n687 gnd 0.009026f
C1829 vdd.t81 gnd 0.129127f
C1830 vdd.t82 gnd 0.138001f
C1831 vdd.t80 gnd 0.168639f
C1832 vdd.n688 gnd 0.216171f
C1833 vdd.n689 gnd 0.181623f
C1834 vdd.n690 gnd 0.01301f
C1835 vdd.n691 gnd 0.010496f
C1836 vdd.n692 gnd 10.9087f
C1837 vdd.n723 gnd 1.47487f
C1838 vdd.n724 gnd 0.010496f
C1839 vdd.n725 gnd 0.010496f
C1840 vdd.n726 gnd 0.025935f
C1841 vdd.n727 gnd 0.009026f
C1842 vdd.n728 gnd 0.010496f
C1843 vdd.n729 gnd 0.008448f
C1844 vdd.n730 gnd 0.006717f
C1845 vdd.n731 gnd 0.033502f
C1846 vdd.n732 gnd 0.008448f
C1847 vdd.n733 gnd 0.010496f
C1848 vdd.n734 gnd 0.010496f
C1849 vdd.n735 gnd 0.010496f
C1850 vdd.n736 gnd 0.010496f
C1851 vdd.n737 gnd 0.010496f
C1852 vdd.n738 gnd 0.010496f
C1853 vdd.n739 gnd 0.010496f
C1854 vdd.n740 gnd 0.010496f
C1855 vdd.n741 gnd 0.010496f
C1856 vdd.n742 gnd 0.010496f
C1857 vdd.n743 gnd 0.010496f
C1858 vdd.n744 gnd 0.010496f
C1859 vdd.n745 gnd 0.010496f
C1860 vdd.n746 gnd 0.010496f
C1861 vdd.n747 gnd 0.007054f
C1862 vdd.n748 gnd 0.010496f
C1863 vdd.n749 gnd 0.010496f
C1864 vdd.n750 gnd 0.010496f
C1865 vdd.n751 gnd 0.010496f
C1866 vdd.n752 gnd 0.010496f
C1867 vdd.n753 gnd 0.010496f
C1868 vdd.n754 gnd 0.010496f
C1869 vdd.n755 gnd 0.010496f
C1870 vdd.n756 gnd 0.010496f
C1871 vdd.n757 gnd 0.010496f
C1872 vdd.n758 gnd 0.010496f
C1873 vdd.n759 gnd 0.010496f
C1874 vdd.n760 gnd 0.010496f
C1875 vdd.n761 gnd 0.010496f
C1876 vdd.n762 gnd 0.010496f
C1877 vdd.n763 gnd 0.010496f
C1878 vdd.n764 gnd 0.010496f
C1879 vdd.n765 gnd 0.010496f
C1880 vdd.n766 gnd 0.010496f
C1881 vdd.n767 gnd 0.008363f
C1882 vdd.t59 gnd 0.129127f
C1883 vdd.t60 gnd 0.138001f
C1884 vdd.t57 gnd 0.168639f
C1885 vdd.n768 gnd 0.216171f
C1886 vdd.n769 gnd 0.181623f
C1887 vdd.n770 gnd 0.010496f
C1888 vdd.n771 gnd 0.010496f
C1889 vdd.n772 gnd 0.010496f
C1890 vdd.n773 gnd 0.010496f
C1891 vdd.n774 gnd 0.010496f
C1892 vdd.n775 gnd 0.010496f
C1893 vdd.n776 gnd 0.010496f
C1894 vdd.n777 gnd 0.010496f
C1895 vdd.n778 gnd 0.010496f
C1896 vdd.n779 gnd 0.010496f
C1897 vdd.n780 gnd 0.010496f
C1898 vdd.n781 gnd 0.010496f
C1899 vdd.n782 gnd 0.010496f
C1900 vdd.n783 gnd 0.006717f
C1901 vdd.n785 gnd 0.007137f
C1902 vdd.n786 gnd 0.007137f
C1903 vdd.n787 gnd 0.007137f
C1904 vdd.n788 gnd 0.007137f
C1905 vdd.n789 gnd 0.007137f
C1906 vdd.n790 gnd 0.007137f
C1907 vdd.n792 gnd 0.007137f
C1908 vdd.n793 gnd 0.007137f
C1909 vdd.n795 gnd 0.007137f
C1910 vdd.n796 gnd 0.005195f
C1911 vdd.n798 gnd 0.007137f
C1912 vdd.t64 gnd 0.288414f
C1913 vdd.t63 gnd 0.295228f
C1914 vdd.t61 gnd 0.188288f
C1915 vdd.n799 gnd 0.101759f
C1916 vdd.n800 gnd 0.057721f
C1917 vdd.n801 gnd 0.0102f
C1918 vdd.n802 gnd 0.016362f
C1919 vdd.n804 gnd 0.007137f
C1920 vdd.n805 gnd 0.72939f
C1921 vdd.n806 gnd 0.015457f
C1922 vdd.n807 gnd 0.015457f
C1923 vdd.n808 gnd 0.007137f
C1924 vdd.n809 gnd 0.01645f
C1925 vdd.n810 gnd 0.007137f
C1926 vdd.n811 gnd 0.007137f
C1927 vdd.n812 gnd 0.007137f
C1928 vdd.n813 gnd 0.007137f
C1929 vdd.n814 gnd 0.007137f
C1930 vdd.n816 gnd 0.007137f
C1931 vdd.n817 gnd 0.007137f
C1932 vdd.n819 gnd 0.007137f
C1933 vdd.n820 gnd 0.007137f
C1934 vdd.n822 gnd 0.007137f
C1935 vdd.n823 gnd 0.007137f
C1936 vdd.n825 gnd 0.007137f
C1937 vdd.n826 gnd 0.007137f
C1938 vdd.n828 gnd 0.007137f
C1939 vdd.n829 gnd 0.007137f
C1940 vdd.n831 gnd 0.007137f
C1941 vdd.t92 gnd 0.288414f
C1942 vdd.t91 gnd 0.295228f
C1943 vdd.t90 gnd 0.188288f
C1944 vdd.n832 gnd 0.101759f
C1945 vdd.n833 gnd 0.057721f
C1946 vdd.n834 gnd 0.007137f
C1947 vdd.n836 gnd 0.007137f
C1948 vdd.n837 gnd 0.007137f
C1949 vdd.t62 gnd 0.364695f
C1950 vdd.n838 gnd 0.007137f
C1951 vdd.n839 gnd 0.007137f
C1952 vdd.n840 gnd 0.007137f
C1953 vdd.n841 gnd 0.007137f
C1954 vdd.n842 gnd 0.007137f
C1955 vdd.n843 gnd 0.72939f
C1956 vdd.n844 gnd 0.007137f
C1957 vdd.n845 gnd 0.007137f
C1958 vdd.n846 gnd 0.595311f
C1959 vdd.n847 gnd 0.007137f
C1960 vdd.n848 gnd 0.007137f
C1961 vdd.n849 gnd 0.007137f
C1962 vdd.n850 gnd 0.007137f
C1963 vdd.n851 gnd 0.72939f
C1964 vdd.n852 gnd 0.007137f
C1965 vdd.n853 gnd 0.007137f
C1966 vdd.n854 gnd 0.007137f
C1967 vdd.n855 gnd 0.007137f
C1968 vdd.n856 gnd 0.007137f
C1969 vdd.t55 gnd 0.364695f
C1970 vdd.n857 gnd 0.007137f
C1971 vdd.n858 gnd 0.007137f
C1972 vdd.n859 gnd 0.007137f
C1973 vdd.n860 gnd 0.007137f
C1974 vdd.n861 gnd 0.007137f
C1975 vdd.t6 gnd 0.364695f
C1976 vdd.n862 gnd 0.007137f
C1977 vdd.n863 gnd 0.007137f
C1978 vdd.n864 gnd 0.724027f
C1979 vdd.n865 gnd 0.007137f
C1980 vdd.n866 gnd 0.007137f
C1981 vdd.n867 gnd 0.007137f
C1982 vdd.t56 gnd 0.364695f
C1983 vdd.n868 gnd 0.007137f
C1984 vdd.n869 gnd 0.007137f
C1985 vdd.n870 gnd 0.563132f
C1986 vdd.n871 gnd 0.007137f
C1987 vdd.n872 gnd 0.007137f
C1988 vdd.n873 gnd 0.007137f
C1989 vdd.n874 gnd 0.488048f
C1990 vdd.n875 gnd 0.007137f
C1991 vdd.n876 gnd 0.007137f
C1992 vdd.n877 gnd 0.402237f
C1993 vdd.n878 gnd 0.007137f
C1994 vdd.n879 gnd 0.007137f
C1995 vdd.n880 gnd 0.007137f
C1996 vdd.n881 gnd 0.600674f
C1997 vdd.n882 gnd 0.007137f
C1998 vdd.n883 gnd 0.007137f
C1999 vdd.t7 gnd 0.364695f
C2000 vdd.n884 gnd 0.007137f
C2001 vdd.t78 gnd 0.295228f
C2002 vdd.t76 gnd 0.188288f
C2003 vdd.t79 gnd 0.295228f
C2004 vdd.n885 gnd 0.16593f
C2005 vdd.n886 gnd 0.007137f
C2006 vdd.n887 gnd 0.007137f
C2007 vdd.n888 gnd 0.72939f
C2008 vdd.n889 gnd 0.007137f
C2009 vdd.n890 gnd 0.007137f
C2010 vdd.t77 gnd 0.284248f
C2011 vdd.t20 gnd 0.128716f
C2012 vdd.n891 gnd 0.007137f
C2013 vdd.n892 gnd 0.007137f
C2014 vdd.n893 gnd 0.007137f
C2015 vdd.t39 gnd 0.364695f
C2016 vdd.n894 gnd 0.007137f
C2017 vdd.n895 gnd 0.007137f
C2018 vdd.n896 gnd 0.007137f
C2019 vdd.n897 gnd 0.007137f
C2020 vdd.n898 gnd 0.007137f
C2021 vdd.t5 gnd 0.364695f
C2022 vdd.n899 gnd 0.007137f
C2023 vdd.n900 gnd 0.007137f
C2024 vdd.n901 gnd 0.648942f
C2025 vdd.n902 gnd 0.007137f
C2026 vdd.n903 gnd 0.007137f
C2027 vdd.n904 gnd 0.007137f
C2028 vdd.n905 gnd 0.402237f
C2029 vdd.n906 gnd 0.007137f
C2030 vdd.n907 gnd 0.007137f
C2031 vdd.t302 gnd 0.364695f
C2032 vdd.n908 gnd 0.007137f
C2033 vdd.n909 gnd 0.007137f
C2034 vdd.n910 gnd 0.007137f
C2035 vdd.n911 gnd 0.563132f
C2036 vdd.n912 gnd 0.007137f
C2037 vdd.n913 gnd 0.007137f
C2038 vdd.t19 gnd 0.268158f
C2039 vdd.t14 gnd 0.327153f
C2040 vdd.n914 gnd 0.007137f
C2041 vdd.n915 gnd 0.007137f
C2042 vdd.n916 gnd 0.007137f
C2043 vdd.t0 gnd 0.364695f
C2044 vdd.n917 gnd 0.007137f
C2045 vdd.n918 gnd 0.007137f
C2046 vdd.t9 gnd 0.364695f
C2047 vdd.n919 gnd 0.007137f
C2048 vdd.n920 gnd 0.007137f
C2049 vdd.n921 gnd 0.007137f
C2050 vdd.t47 gnd 0.364695f
C2051 vdd.n922 gnd 0.007137f
C2052 vdd.n923 gnd 0.007137f
C2053 vdd.t11 gnd 0.364695f
C2054 vdd.n924 gnd 0.007137f
C2055 vdd.n925 gnd 0.007137f
C2056 vdd.n926 gnd 0.007137f
C2057 vdd.n927 gnd 0.72939f
C2058 vdd.n928 gnd 0.007137f
C2059 vdd.n929 gnd 0.007137f
C2060 vdd.n930 gnd 0.504137f
C2061 vdd.n931 gnd 0.007137f
C2062 vdd.n932 gnd 0.007137f
C2063 vdd.n933 gnd 0.007137f
C2064 vdd.t40 gnd 0.364695f
C2065 vdd.n934 gnd 0.007137f
C2066 vdd.n935 gnd 0.007137f
C2067 vdd.n936 gnd 0.007137f
C2068 vdd.n937 gnd 0.007137f
C2069 vdd.n938 gnd 0.007137f
C2070 vdd.t51 gnd 0.364695f
C2071 vdd.n939 gnd 0.007137f
C2072 vdd.n940 gnd 0.007137f
C2073 vdd.t108 gnd 0.364695f
C2074 vdd.n941 gnd 0.007137f
C2075 vdd.n942 gnd 0.01645f
C2076 vdd.n943 gnd 0.01645f
C2077 vdd.t53 gnd 0.643579f
C2078 vdd.n944 gnd 0.015457f
C2079 vdd.n945 gnd 0.015457f
C2080 vdd.n946 gnd 0.4076f
C2081 vdd.n947 gnd 0.01645f
C2082 vdd.n948 gnd 0.007137f
C2083 vdd.n949 gnd 0.007137f
C2084 vdd.t296 gnd 0.643579f
C2085 vdd.n967 gnd 0.01645f
C2086 vdd.n985 gnd 0.015457f
C2087 vdd.n986 gnd 0.007137f
C2088 vdd.n987 gnd 0.015457f
C2089 vdd.t129 gnd 0.288414f
C2090 vdd.t128 gnd 0.295228f
C2091 vdd.t127 gnd 0.188288f
C2092 vdd.n988 gnd 0.101759f
C2093 vdd.n989 gnd 0.057721f
C2094 vdd.n990 gnd 0.016362f
C2095 vdd.n991 gnd 0.007137f
C2096 vdd.n992 gnd 0.4076f
C2097 vdd.n993 gnd 0.015457f
C2098 vdd.n994 gnd 0.007137f
C2099 vdd.n995 gnd 0.01645f
C2100 vdd.n996 gnd 0.007137f
C2101 vdd.t106 gnd 0.288414f
C2102 vdd.t105 gnd 0.295228f
C2103 vdd.t103 gnd 0.188288f
C2104 vdd.n997 gnd 0.101759f
C2105 vdd.n998 gnd 0.057721f
C2106 vdd.n999 gnd 0.0102f
C2107 vdd.n1000 gnd 0.007137f
C2108 vdd.n1001 gnd 0.007137f
C2109 vdd.t104 gnd 0.364695f
C2110 vdd.n1002 gnd 0.007137f
C2111 vdd.t294 gnd 0.364695f
C2112 vdd.n1003 gnd 0.007137f
C2113 vdd.n1004 gnd 0.007137f
C2114 vdd.n1005 gnd 0.007137f
C2115 vdd.n1006 gnd 0.007137f
C2116 vdd.n1007 gnd 0.007137f
C2117 vdd.n1008 gnd 0.72939f
C2118 vdd.n1009 gnd 0.007137f
C2119 vdd.n1010 gnd 0.007137f
C2120 vdd.t300 gnd 0.364695f
C2121 vdd.n1011 gnd 0.007137f
C2122 vdd.n1012 gnd 0.007137f
C2123 vdd.n1013 gnd 0.007137f
C2124 vdd.n1014 gnd 0.007137f
C2125 vdd.n1015 gnd 0.504137f
C2126 vdd.n1016 gnd 0.007137f
C2127 vdd.n1017 gnd 0.007137f
C2128 vdd.n1018 gnd 0.007137f
C2129 vdd.n1019 gnd 0.007137f
C2130 vdd.n1020 gnd 0.007137f
C2131 vdd.t293 gnd 0.364695f
C2132 vdd.n1021 gnd 0.007137f
C2133 vdd.n1022 gnd 0.007137f
C2134 vdd.t37 gnd 0.364695f
C2135 vdd.n1023 gnd 0.007137f
C2136 vdd.n1024 gnd 0.007137f
C2137 vdd.n1025 gnd 0.007137f
C2138 vdd.t42 gnd 0.364695f
C2139 vdd.n1026 gnd 0.007137f
C2140 vdd.n1027 gnd 0.007137f
C2141 vdd.t12 gnd 0.364695f
C2142 vdd.n1028 gnd 0.007137f
C2143 vdd.n1029 gnd 0.007137f
C2144 vdd.n1030 gnd 0.007137f
C2145 vdd.t49 gnd 0.327153f
C2146 vdd.n1031 gnd 0.007137f
C2147 vdd.n1032 gnd 0.007137f
C2148 vdd.n1033 gnd 0.563132f
C2149 vdd.n1034 gnd 0.007137f
C2150 vdd.n1035 gnd 0.007137f
C2151 vdd.n1036 gnd 0.007137f
C2152 vdd.t2 gnd 0.364695f
C2153 vdd.n1037 gnd 0.007137f
C2154 vdd.n1038 gnd 0.007137f
C2155 vdd.t8 gnd 0.268158f
C2156 vdd.n1039 gnd 0.402237f
C2157 vdd.n1040 gnd 0.007137f
C2158 vdd.n1041 gnd 0.007137f
C2159 vdd.n1042 gnd 0.007137f
C2160 vdd.n1043 gnd 0.648942f
C2161 vdd.n1044 gnd 0.007137f
C2162 vdd.n1045 gnd 0.007137f
C2163 vdd.t16 gnd 0.364695f
C2164 vdd.n1046 gnd 0.007137f
C2165 vdd.n1047 gnd 0.007137f
C2166 vdd.n1048 gnd 0.007137f
C2167 vdd.n1049 gnd 0.72939f
C2168 vdd.n1050 gnd 0.007137f
C2169 vdd.n1051 gnd 0.007137f
C2170 vdd.t45 gnd 0.364695f
C2171 vdd.n1052 gnd 0.007137f
C2172 vdd.n1053 gnd 0.007137f
C2173 vdd.n1054 gnd 0.007137f
C2174 vdd.t46 gnd 0.128716f
C2175 vdd.n1055 gnd 0.007137f
C2176 vdd.n1056 gnd 0.007137f
C2177 vdd.n1057 gnd 0.007137f
C2178 vdd.t119 gnd 0.295228f
C2179 vdd.t117 gnd 0.188288f
C2180 vdd.t120 gnd 0.295228f
C2181 vdd.n1058 gnd 0.16593f
C2182 vdd.n1059 gnd 0.007137f
C2183 vdd.n1060 gnd 0.007137f
C2184 vdd.t4 gnd 0.364695f
C2185 vdd.n1061 gnd 0.007137f
C2186 vdd.n1062 gnd 0.007137f
C2187 vdd.t118 gnd 0.284248f
C2188 vdd.n1063 gnd 0.600674f
C2189 vdd.n1064 gnd 0.007137f
C2190 vdd.n1065 gnd 0.007137f
C2191 vdd.n1066 gnd 0.007137f
C2192 vdd.n1067 gnd 0.402237f
C2193 vdd.n1068 gnd 0.007137f
C2194 vdd.n1069 gnd 0.007137f
C2195 vdd.n1070 gnd 0.488048f
C2196 vdd.n1071 gnd 0.007137f
C2197 vdd.n1072 gnd 0.007137f
C2198 vdd.n1073 gnd 0.007137f
C2199 vdd.n1074 gnd 0.563132f
C2200 vdd.n1075 gnd 0.007137f
C2201 vdd.n1076 gnd 0.007137f
C2202 vdd.t17 gnd 0.364695f
C2203 vdd.n1077 gnd 0.007137f
C2204 vdd.n1078 gnd 0.007137f
C2205 vdd.n1079 gnd 0.007137f
C2206 vdd.n1080 gnd 0.724027f
C2207 vdd.n1081 gnd 0.007137f
C2208 vdd.n1082 gnd 0.007137f
C2209 vdd.t10 gnd 0.364695f
C2210 vdd.n1083 gnd 0.007137f
C2211 vdd.n1084 gnd 0.007137f
C2212 vdd.n1085 gnd 0.007137f
C2213 vdd.n1086 gnd 0.72939f
C2214 vdd.n1087 gnd 0.007137f
C2215 vdd.n1088 gnd 0.007137f
C2216 vdd.t18 gnd 0.364695f
C2217 vdd.n1089 gnd 0.007137f
C2218 vdd.n1090 gnd 0.007137f
C2219 vdd.n1091 gnd 0.007137f
C2220 vdd.n1092 gnd 0.72939f
C2221 vdd.n1093 gnd 0.007137f
C2222 vdd.n1094 gnd 0.007137f
C2223 vdd.n1095 gnd 0.007137f
C2224 vdd.n1096 gnd 0.007137f
C2225 vdd.n1097 gnd 0.007137f
C2226 vdd.n1098 gnd 0.595311f
C2227 vdd.n1099 gnd 0.007137f
C2228 vdd.n1100 gnd 0.007137f
C2229 vdd.n1101 gnd 0.007137f
C2230 vdd.n1102 gnd 0.007137f
C2231 vdd.n1103 gnd 0.007137f
C2232 vdd.n1104 gnd 0.72939f
C2233 vdd.n1105 gnd 0.007137f
C2234 vdd.n1106 gnd 0.007137f
C2235 vdd.t66 gnd 0.364695f
C2236 vdd.n1107 gnd 0.007137f
C2237 vdd.n1108 gnd 0.01645f
C2238 vdd.n1109 gnd 0.01645f
C2239 vdd.n1110 gnd 10.9087f
C2240 vdd.n1111 gnd 0.015457f
C2241 vdd.n1112 gnd 0.015457f
C2242 vdd.n1113 gnd 0.01645f
C2243 vdd.n1114 gnd 0.007137f
C2244 vdd.n1116 gnd 0.007137f
C2245 vdd.n1117 gnd 0.007137f
C2246 vdd.n1118 gnd 0.007137f
C2247 vdd.n1119 gnd 0.007137f
C2248 vdd.n1120 gnd 0.007137f
C2249 vdd.n1121 gnd 0.007137f
C2250 vdd.n1122 gnd 0.037553f
C2251 vdd.n1123 gnd 0.007137f
C2252 vdd.n1124 gnd 0.007137f
C2253 vdd.n1125 gnd 0.007137f
C2254 vdd.n1126 gnd 0.007137f
C2255 vdd.n1127 gnd 0.007137f
C2256 vdd.n1128 gnd 0.007137f
C2257 vdd.n1129 gnd 0.007137f
C2258 vdd.t131 gnd 0.288414f
C2259 vdd.t132 gnd 0.295228f
C2260 vdd.t130 gnd 0.188288f
C2261 vdd.n1130 gnd 0.101759f
C2262 vdd.n1131 gnd 0.057721f
C2263 vdd.n1132 gnd 0.007137f
C2264 vdd.n1133 gnd 0.007137f
C2265 vdd.n1134 gnd 0.007137f
C2266 vdd.n1135 gnd 0.007137f
C2267 vdd.t67 gnd 0.288414f
C2268 vdd.t68 gnd 0.295228f
C2269 vdd.t65 gnd 0.188288f
C2270 vdd.n1136 gnd 0.101759f
C2271 vdd.n1137 gnd 0.057721f
C2272 vdd.n1138 gnd 0.007137f
C2273 vdd.n1139 gnd 0.007137f
C2274 vdd.n1140 gnd 0.007137f
C2275 vdd.n1141 gnd 0.007137f
C2276 vdd.n1142 gnd 0.007137f
C2277 vdd.n1143 gnd 0.007137f
C2278 vdd.n1144 gnd 0.006717f
C2279 vdd.n1147 gnd 0.025935f
C2280 vdd.n1148 gnd 0.008448f
C2281 vdd.n1149 gnd 0.010496f
C2282 vdd.n1151 gnd 0.010496f
C2283 vdd.n1152 gnd 0.007012f
C2284 vdd.t84 gnd 0.536316f
C2285 vdd.n1153 gnd 11.3163f
C2286 vdd.n1154 gnd 0.010496f
C2287 vdd.n1155 gnd 0.025935f
C2288 vdd.n1156 gnd 0.008448f
C2289 vdd.n1157 gnd 0.010496f
C2290 vdd.n1158 gnd 0.008448f
C2291 vdd.n1159 gnd 0.010496f
C2292 vdd.n1160 gnd 1.07263f
C2293 vdd.n1161 gnd 0.010496f
C2294 vdd.n1162 gnd 0.008448f
C2295 vdd.n1163 gnd 0.008448f
C2296 vdd.n1164 gnd 0.010496f
C2297 vdd.n1165 gnd 0.008448f
C2298 vdd.n1166 gnd 0.010496f
C2299 vdd.t232 gnd 0.536316f
C2300 vdd.n1167 gnd 0.010496f
C2301 vdd.n1168 gnd 0.008448f
C2302 vdd.n1169 gnd 0.010496f
C2303 vdd.n1170 gnd 0.008448f
C2304 vdd.n1171 gnd 0.010496f
C2305 vdd.t145 gnd 0.536316f
C2306 vdd.n1172 gnd 0.010496f
C2307 vdd.n1173 gnd 0.008448f
C2308 vdd.n1174 gnd 0.010496f
C2309 vdd.n1175 gnd 0.008448f
C2310 vdd.n1176 gnd 0.010496f
C2311 vdd.n1177 gnd 0.863469f
C2312 vdd.n1178 gnd 0.890285f
C2313 vdd.t196 gnd 0.536316f
C2314 vdd.n1179 gnd 0.010496f
C2315 vdd.n1180 gnd 0.008448f
C2316 vdd.n1181 gnd 0.010496f
C2317 vdd.n1182 gnd 0.008448f
C2318 vdd.n1183 gnd 0.010496f
C2319 vdd.n1184 gnd 0.681121f
C2320 vdd.n1185 gnd 0.010496f
C2321 vdd.n1186 gnd 0.008448f
C2322 vdd.n1187 gnd 0.010496f
C2323 vdd.n1188 gnd 0.008448f
C2324 vdd.n1189 gnd 0.010496f
C2325 vdd.t226 gnd 0.536316f
C2326 vdd.t173 gnd 0.536316f
C2327 vdd.n1190 gnd 0.010496f
C2328 vdd.n1191 gnd 0.008448f
C2329 vdd.n1192 gnd 0.010496f
C2330 vdd.n1193 gnd 0.008448f
C2331 vdd.n1194 gnd 0.010496f
C2332 vdd.t230 gnd 0.536316f
C2333 vdd.n1195 gnd 0.010496f
C2334 vdd.n1196 gnd 0.008448f
C2335 vdd.n1197 gnd 0.010496f
C2336 vdd.n1198 gnd 0.008448f
C2337 vdd.n1199 gnd 0.010496f
C2338 vdd.t143 gnd 0.536316f
C2339 vdd.n1200 gnd 0.756206f
C2340 vdd.n1201 gnd 0.010496f
C2341 vdd.n1202 gnd 0.008448f
C2342 vdd.n1203 gnd 0.010496f
C2343 vdd.n1204 gnd 0.008448f
C2344 vdd.n1205 gnd 0.010496f
C2345 vdd.n1206 gnd 0.842016f
C2346 vdd.n1207 gnd 0.010496f
C2347 vdd.n1208 gnd 0.008448f
C2348 vdd.n1209 gnd 0.010496f
C2349 vdd.n1210 gnd 0.008448f
C2350 vdd.n1211 gnd 0.010496f
C2351 vdd.n1212 gnd 0.659669f
C2352 vdd.t170 gnd 0.536316f
C2353 vdd.n1213 gnd 0.010496f
C2354 vdd.n1214 gnd 0.008448f
C2355 vdd.n1215 gnd 0.010496f
C2356 vdd.n1216 gnd 0.008448f
C2357 vdd.n1217 gnd 0.010496f
C2358 vdd.t139 gnd 0.536316f
C2359 vdd.n1218 gnd 0.010496f
C2360 vdd.n1219 gnd 0.008448f
C2361 vdd.n1220 gnd 0.010496f
C2362 vdd.n1221 gnd 0.008448f
C2363 vdd.n1222 gnd 0.010496f
C2364 vdd.t198 gnd 0.536316f
C2365 vdd.n1223 gnd 0.595311f
C2366 vdd.n1224 gnd 0.010496f
C2367 vdd.n1225 gnd 0.008448f
C2368 vdd.n1226 gnd 0.010496f
C2369 vdd.n1227 gnd 0.008448f
C2370 vdd.n1228 gnd 0.010496f
C2371 vdd.t224 gnd 0.536316f
C2372 vdd.n1229 gnd 0.010496f
C2373 vdd.n1230 gnd 0.008448f
C2374 vdd.n1231 gnd 0.010496f
C2375 vdd.n1232 gnd 0.008448f
C2376 vdd.n1233 gnd 0.010496f
C2377 vdd.n1234 gnd 0.820564f
C2378 vdd.n1235 gnd 0.890285f
C2379 vdd.t133 gnd 0.536316f
C2380 vdd.n1236 gnd 0.010496f
C2381 vdd.n1237 gnd 0.008448f
C2382 vdd.n1238 gnd 0.010496f
C2383 vdd.n1239 gnd 0.008448f
C2384 vdd.n1240 gnd 0.010496f
C2385 vdd.n1241 gnd 0.638216f
C2386 vdd.n1242 gnd 0.010496f
C2387 vdd.n1243 gnd 0.008448f
C2388 vdd.n1244 gnd 0.010496f
C2389 vdd.n1245 gnd 0.008448f
C2390 vdd.n1246 gnd 0.010496f
C2391 vdd.t214 gnd 0.536316f
C2392 vdd.t245 gnd 0.536316f
C2393 vdd.n1247 gnd 0.010496f
C2394 vdd.n1248 gnd 0.008448f
C2395 vdd.n1249 gnd 0.010496f
C2396 vdd.n1250 gnd 0.008448f
C2397 vdd.n1251 gnd 0.010496f
C2398 vdd.t175 gnd 0.536316f
C2399 vdd.n1252 gnd 0.010496f
C2400 vdd.n1253 gnd 0.008448f
C2401 vdd.n1254 gnd 0.010496f
C2402 vdd.n1255 gnd 0.008448f
C2403 vdd.n1256 gnd 0.010496f
C2404 vdd.t228 gnd 0.536316f
C2405 vdd.n1257 gnd 0.799111f
C2406 vdd.n1258 gnd 0.010496f
C2407 vdd.n1259 gnd 0.008448f
C2408 vdd.n1260 gnd 0.010496f
C2409 vdd.n1261 gnd 0.008448f
C2410 vdd.n1262 gnd 0.010496f
C2411 vdd.n1263 gnd 1.07263f
C2412 vdd.n1264 gnd 0.010496f
C2413 vdd.n1265 gnd 0.008448f
C2414 vdd.n1266 gnd 0.02539f
C2415 vdd.n1267 gnd 0.007012f
C2416 vdd.n1268 gnd 0.02539f
C2417 vdd.t100 gnd 0.536316f
C2418 vdd.n1269 gnd 0.02539f
C2419 vdd.n1270 gnd 0.007012f
C2420 vdd.n1271 gnd 0.010496f
C2421 vdd.n1272 gnd 0.008448f
C2422 vdd.n1273 gnd 0.010496f
C2423 vdd.n1304 gnd 0.025935f
C2424 vdd.n1305 gnd 1.58213f
C2425 vdd.n1306 gnd 0.010496f
C2426 vdd.n1307 gnd 0.008448f
C2427 vdd.n1308 gnd 0.010496f
C2428 vdd.n1309 gnd 0.010496f
C2429 vdd.n1310 gnd 0.010496f
C2430 vdd.n1311 gnd 0.010496f
C2431 vdd.n1312 gnd 0.010496f
C2432 vdd.n1313 gnd 0.008448f
C2433 vdd.n1314 gnd 0.010496f
C2434 vdd.n1315 gnd 0.010496f
C2435 vdd.n1316 gnd 0.010496f
C2436 vdd.n1317 gnd 0.010496f
C2437 vdd.n1318 gnd 0.010496f
C2438 vdd.n1319 gnd 0.008448f
C2439 vdd.n1320 gnd 0.010496f
C2440 vdd.n1321 gnd 0.010496f
C2441 vdd.n1322 gnd 0.010496f
C2442 vdd.n1323 gnd 0.010496f
C2443 vdd.n1324 gnd 0.010496f
C2444 vdd.n1325 gnd 0.008448f
C2445 vdd.n1326 gnd 0.010496f
C2446 vdd.n1327 gnd 0.010496f
C2447 vdd.n1328 gnd 0.010496f
C2448 vdd.n1329 gnd 0.010496f
C2449 vdd.n1330 gnd 0.010496f
C2450 vdd.t125 gnd 0.129127f
C2451 vdd.t126 gnd 0.138001f
C2452 vdd.t124 gnd 0.168639f
C2453 vdd.n1331 gnd 0.216171f
C2454 vdd.n1332 gnd 0.182467f
C2455 vdd.n1333 gnd 0.018079f
C2456 vdd.n1334 gnd 0.010496f
C2457 vdd.n1335 gnd 0.010496f
C2458 vdd.n1336 gnd 0.010496f
C2459 vdd.n1337 gnd 0.010496f
C2460 vdd.n1338 gnd 0.010496f
C2461 vdd.n1339 gnd 0.008448f
C2462 vdd.n1340 gnd 0.010496f
C2463 vdd.n1341 gnd 0.010496f
C2464 vdd.n1342 gnd 0.010496f
C2465 vdd.n1343 gnd 0.010496f
C2466 vdd.n1344 gnd 0.010496f
C2467 vdd.n1345 gnd 0.008448f
C2468 vdd.n1346 gnd 0.010496f
C2469 vdd.n1347 gnd 0.010496f
C2470 vdd.n1348 gnd 0.010496f
C2471 vdd.n1349 gnd 0.010496f
C2472 vdd.n1350 gnd 0.010496f
C2473 vdd.n1351 gnd 0.008448f
C2474 vdd.n1352 gnd 0.010496f
C2475 vdd.n1353 gnd 0.010496f
C2476 vdd.n1354 gnd 0.010496f
C2477 vdd.n1355 gnd 0.010496f
C2478 vdd.n1356 gnd 0.010496f
C2479 vdd.n1357 gnd 0.008448f
C2480 vdd.n1358 gnd 0.010496f
C2481 vdd.n1359 gnd 0.010496f
C2482 vdd.n1360 gnd 0.010496f
C2483 vdd.n1361 gnd 0.010496f
C2484 vdd.n1362 gnd 0.010496f
C2485 vdd.n1363 gnd 0.008448f
C2486 vdd.n1364 gnd 0.010496f
C2487 vdd.n1365 gnd 0.010496f
C2488 vdd.n1366 gnd 0.010496f
C2489 vdd.n1367 gnd 0.010496f
C2490 vdd.n1368 gnd 0.008448f
C2491 vdd.n1369 gnd 0.010496f
C2492 vdd.n1370 gnd 0.010496f
C2493 vdd.n1371 gnd 0.010496f
C2494 vdd.n1372 gnd 0.010496f
C2495 vdd.n1373 gnd 0.010496f
C2496 vdd.n1374 gnd 0.008448f
C2497 vdd.n1375 gnd 0.010496f
C2498 vdd.n1376 gnd 0.010496f
C2499 vdd.n1377 gnd 0.010496f
C2500 vdd.n1378 gnd 0.010496f
C2501 vdd.n1379 gnd 0.010496f
C2502 vdd.n1380 gnd 0.008448f
C2503 vdd.n1381 gnd 0.010496f
C2504 vdd.n1382 gnd 0.010496f
C2505 vdd.n1383 gnd 0.010496f
C2506 vdd.n1384 gnd 0.010496f
C2507 vdd.n1385 gnd 0.010496f
C2508 vdd.n1386 gnd 0.008448f
C2509 vdd.n1387 gnd 0.010496f
C2510 vdd.n1388 gnd 0.010496f
C2511 vdd.n1389 gnd 0.010496f
C2512 vdd.n1390 gnd 0.010496f
C2513 vdd.n1391 gnd 0.010496f
C2514 vdd.n1392 gnd 0.008448f
C2515 vdd.n1393 gnd 0.010496f
C2516 vdd.n1394 gnd 0.010496f
C2517 vdd.n1395 gnd 0.010496f
C2518 vdd.n1396 gnd 0.010496f
C2519 vdd.t101 gnd 0.129127f
C2520 vdd.t102 gnd 0.138001f
C2521 vdd.t99 gnd 0.168639f
C2522 vdd.n1397 gnd 0.216171f
C2523 vdd.n1398 gnd 0.182467f
C2524 vdd.n1399 gnd 0.013855f
C2525 vdd.n1400 gnd 0.004013f
C2526 vdd.n1401 gnd 0.025935f
C2527 vdd.n1402 gnd 0.010496f
C2528 vdd.n1403 gnd 0.004435f
C2529 vdd.n1404 gnd 0.008448f
C2530 vdd.n1405 gnd 0.008448f
C2531 vdd.n1406 gnd 0.010496f
C2532 vdd.n1407 gnd 0.010496f
C2533 vdd.n1408 gnd 0.010496f
C2534 vdd.n1409 gnd 0.008448f
C2535 vdd.n1410 gnd 0.008448f
C2536 vdd.n1411 gnd 0.008448f
C2537 vdd.n1412 gnd 0.010496f
C2538 vdd.n1413 gnd 0.010496f
C2539 vdd.n1414 gnd 0.010496f
C2540 vdd.n1415 gnd 0.008448f
C2541 vdd.n1416 gnd 0.008448f
C2542 vdd.n1417 gnd 0.008448f
C2543 vdd.n1418 gnd 0.010496f
C2544 vdd.n1419 gnd 0.010496f
C2545 vdd.n1420 gnd 0.010496f
C2546 vdd.n1421 gnd 0.008448f
C2547 vdd.n1422 gnd 0.008448f
C2548 vdd.n1423 gnd 0.008448f
C2549 vdd.n1424 gnd 0.010496f
C2550 vdd.n1425 gnd 0.010496f
C2551 vdd.n1426 gnd 0.010496f
C2552 vdd.n1427 gnd 0.008448f
C2553 vdd.n1428 gnd 0.008448f
C2554 vdd.n1429 gnd 0.008448f
C2555 vdd.n1430 gnd 0.010496f
C2556 vdd.n1431 gnd 0.010496f
C2557 vdd.n1432 gnd 0.010496f
C2558 vdd.n1433 gnd 0.008363f
C2559 vdd.n1434 gnd 0.010496f
C2560 vdd.t112 gnd 0.129127f
C2561 vdd.t113 gnd 0.138001f
C2562 vdd.t111 gnd 0.168639f
C2563 vdd.n1435 gnd 0.216171f
C2564 vdd.n1436 gnd 0.182467f
C2565 vdd.n1437 gnd 0.018079f
C2566 vdd.n1438 gnd 0.005745f
C2567 vdd.n1439 gnd 0.010496f
C2568 vdd.n1440 gnd 0.010496f
C2569 vdd.n1441 gnd 0.010496f
C2570 vdd.n1442 gnd 0.008448f
C2571 vdd.n1443 gnd 0.008448f
C2572 vdd.n1444 gnd 0.008448f
C2573 vdd.n1445 gnd 0.010496f
C2574 vdd.n1446 gnd 0.010496f
C2575 vdd.n1447 gnd 0.010496f
C2576 vdd.n1448 gnd 0.008448f
C2577 vdd.n1449 gnd 0.008448f
C2578 vdd.n1450 gnd 0.008448f
C2579 vdd.n1451 gnd 0.010496f
C2580 vdd.n1452 gnd 0.010496f
C2581 vdd.n1453 gnd 0.010496f
C2582 vdd.n1454 gnd 0.008448f
C2583 vdd.n1455 gnd 0.008448f
C2584 vdd.n1456 gnd 0.008448f
C2585 vdd.n1457 gnd 0.010496f
C2586 vdd.n1458 gnd 0.010496f
C2587 vdd.n1459 gnd 0.010496f
C2588 vdd.n1460 gnd 0.008448f
C2589 vdd.n1461 gnd 0.008448f
C2590 vdd.n1462 gnd 0.008448f
C2591 vdd.n1463 gnd 0.010496f
C2592 vdd.n1464 gnd 0.010496f
C2593 vdd.n1465 gnd 0.010496f
C2594 vdd.n1466 gnd 0.008448f
C2595 vdd.n1467 gnd 0.008448f
C2596 vdd.n1468 gnd 0.007054f
C2597 vdd.n1469 gnd 0.010496f
C2598 vdd.n1470 gnd 0.010496f
C2599 vdd.n1471 gnd 0.010496f
C2600 vdd.n1472 gnd 0.007054f
C2601 vdd.n1473 gnd 0.008448f
C2602 vdd.n1474 gnd 0.008448f
C2603 vdd.n1475 gnd 0.010496f
C2604 vdd.n1476 gnd 0.010496f
C2605 vdd.n1477 gnd 0.010496f
C2606 vdd.n1478 gnd 0.008448f
C2607 vdd.n1479 gnd 0.008448f
C2608 vdd.n1480 gnd 0.008448f
C2609 vdd.n1481 gnd 0.010496f
C2610 vdd.n1482 gnd 0.010496f
C2611 vdd.n1483 gnd 0.010496f
C2612 vdd.n1484 gnd 0.008448f
C2613 vdd.n1485 gnd 0.008448f
C2614 vdd.n1486 gnd 0.008448f
C2615 vdd.n1487 gnd 0.010496f
C2616 vdd.n1488 gnd 0.010496f
C2617 vdd.n1489 gnd 0.010496f
C2618 vdd.n1490 gnd 0.008448f
C2619 vdd.n1491 gnd 0.008448f
C2620 vdd.n1492 gnd 0.008448f
C2621 vdd.n1493 gnd 0.010496f
C2622 vdd.n1494 gnd 0.010496f
C2623 vdd.n1495 gnd 0.010496f
C2624 vdd.n1496 gnd 0.008448f
C2625 vdd.n1497 gnd 0.010496f
C2626 vdd.n1498 gnd 2.54214f
C2627 vdd.n1500 gnd 0.025935f
C2628 vdd.n1501 gnd 0.007012f
C2629 vdd.n1502 gnd 0.025935f
C2630 vdd.n1503 gnd 0.02539f
C2631 vdd.n1504 gnd 0.010496f
C2632 vdd.n1505 gnd 0.008448f
C2633 vdd.n1506 gnd 0.010496f
C2634 vdd.n1507 gnd 0.541679f
C2635 vdd.n1508 gnd 0.010496f
C2636 vdd.n1509 gnd 0.008448f
C2637 vdd.n1510 gnd 0.010496f
C2638 vdd.n1511 gnd 0.010496f
C2639 vdd.n1512 gnd 0.010496f
C2640 vdd.n1513 gnd 0.008448f
C2641 vdd.n1514 gnd 0.010496f
C2642 vdd.n1515 gnd 0.981458f
C2643 vdd.n1516 gnd 1.07263f
C2644 vdd.n1517 gnd 0.010496f
C2645 vdd.n1518 gnd 0.008448f
C2646 vdd.n1519 gnd 0.010496f
C2647 vdd.n1520 gnd 0.010496f
C2648 vdd.n1521 gnd 0.010496f
C2649 vdd.n1522 gnd 0.008448f
C2650 vdd.n1523 gnd 0.010496f
C2651 vdd.n1524 gnd 0.62749f
C2652 vdd.n1525 gnd 0.010496f
C2653 vdd.n1526 gnd 0.008448f
C2654 vdd.n1527 gnd 0.010496f
C2655 vdd.n1528 gnd 0.010496f
C2656 vdd.n1529 gnd 0.010496f
C2657 vdd.n1530 gnd 0.008448f
C2658 vdd.n1531 gnd 0.010496f
C2659 vdd.n1532 gnd 0.616763f
C2660 vdd.n1533 gnd 0.809837f
C2661 vdd.n1534 gnd 0.010496f
C2662 vdd.n1535 gnd 0.008448f
C2663 vdd.n1536 gnd 0.010496f
C2664 vdd.n1537 gnd 0.010496f
C2665 vdd.n1538 gnd 0.010496f
C2666 vdd.n1539 gnd 0.008448f
C2667 vdd.n1540 gnd 0.010496f
C2668 vdd.n1541 gnd 0.890285f
C2669 vdd.n1542 gnd 0.010496f
C2670 vdd.n1543 gnd 0.008448f
C2671 vdd.n1544 gnd 0.010496f
C2672 vdd.n1545 gnd 0.010496f
C2673 vdd.n1546 gnd 0.010496f
C2674 vdd.n1547 gnd 0.008448f
C2675 vdd.n1548 gnd 0.010496f
C2676 vdd.t186 gnd 0.536316f
C2677 vdd.n1549 gnd 0.788385f
C2678 vdd.n1550 gnd 0.010496f
C2679 vdd.n1551 gnd 0.008448f
C2680 vdd.n1552 gnd 0.010496f
C2681 vdd.n1553 gnd 0.010496f
C2682 vdd.n1554 gnd 0.010496f
C2683 vdd.n1555 gnd 0.008448f
C2684 vdd.n1556 gnd 0.010496f
C2685 vdd.n1557 gnd 0.606037f
C2686 vdd.n1558 gnd 0.010496f
C2687 vdd.n1559 gnd 0.008448f
C2688 vdd.n1560 gnd 0.010496f
C2689 vdd.n1561 gnd 0.010496f
C2690 vdd.n1562 gnd 0.010496f
C2691 vdd.n1563 gnd 0.008448f
C2692 vdd.n1564 gnd 0.010496f
C2693 vdd.n1565 gnd 0.777658f
C2694 vdd.n1566 gnd 0.648942f
C2695 vdd.n1567 gnd 0.010496f
C2696 vdd.n1568 gnd 0.008448f
C2697 vdd.n1569 gnd 0.010496f
C2698 vdd.n1570 gnd 0.010496f
C2699 vdd.n1571 gnd 0.010496f
C2700 vdd.n1572 gnd 0.008448f
C2701 vdd.n1573 gnd 0.010496f
C2702 vdd.n1574 gnd 0.83129f
C2703 vdd.n1575 gnd 0.010496f
C2704 vdd.n1576 gnd 0.008448f
C2705 vdd.n1577 gnd 0.010496f
C2706 vdd.n1578 gnd 0.010496f
C2707 vdd.n1579 gnd 0.010496f
C2708 vdd.n1580 gnd 0.008448f
C2709 vdd.n1581 gnd 0.010496f
C2710 vdd.t135 gnd 0.536316f
C2711 vdd.n1582 gnd 0.890285f
C2712 vdd.n1583 gnd 0.010496f
C2713 vdd.n1584 gnd 0.008448f
C2714 vdd.n1585 gnd 0.010496f
C2715 vdd.n1586 gnd 0.008067f
C2716 vdd.n1587 gnd 0.00576f
C2717 vdd.n1588 gnd 0.005345f
C2718 vdd.n1589 gnd 0.002957f
C2719 vdd.n1590 gnd 0.006789f
C2720 vdd.n1591 gnd 0.002872f
C2721 vdd.n1592 gnd 0.003041f
C2722 vdd.n1593 gnd 0.005345f
C2723 vdd.n1594 gnd 0.002872f
C2724 vdd.n1595 gnd 0.006789f
C2725 vdd.n1596 gnd 0.003041f
C2726 vdd.n1597 gnd 0.005345f
C2727 vdd.n1598 gnd 0.002872f
C2728 vdd.n1599 gnd 0.005092f
C2729 vdd.n1600 gnd 0.005107f
C2730 vdd.t233 gnd 0.014586f
C2731 vdd.n1601 gnd 0.032453f
C2732 vdd.n1602 gnd 0.168893f
C2733 vdd.n1603 gnd 0.002872f
C2734 vdd.n1604 gnd 0.003041f
C2735 vdd.n1605 gnd 0.006789f
C2736 vdd.n1606 gnd 0.006789f
C2737 vdd.n1607 gnd 0.003041f
C2738 vdd.n1608 gnd 0.002872f
C2739 vdd.n1609 gnd 0.005345f
C2740 vdd.n1610 gnd 0.005345f
C2741 vdd.n1611 gnd 0.002872f
C2742 vdd.n1612 gnd 0.003041f
C2743 vdd.n1613 gnd 0.006789f
C2744 vdd.n1614 gnd 0.006789f
C2745 vdd.n1615 gnd 0.003041f
C2746 vdd.n1616 gnd 0.002872f
C2747 vdd.n1617 gnd 0.005345f
C2748 vdd.n1618 gnd 0.005345f
C2749 vdd.n1619 gnd 0.002872f
C2750 vdd.n1620 gnd 0.003041f
C2751 vdd.n1621 gnd 0.006789f
C2752 vdd.n1622 gnd 0.006789f
C2753 vdd.n1623 gnd 0.016051f
C2754 vdd.n1624 gnd 0.002957f
C2755 vdd.n1625 gnd 0.002872f
C2756 vdd.n1626 gnd 0.013816f
C2757 vdd.n1627 gnd 0.009645f
C2758 vdd.t197 gnd 0.033792f
C2759 vdd.t146 gnd 0.033792f
C2760 vdd.n1628 gnd 0.23224f
C2761 vdd.n1629 gnd 0.182621f
C2762 vdd.t221 gnd 0.033792f
C2763 vdd.t159 gnd 0.033792f
C2764 vdd.n1630 gnd 0.23224f
C2765 vdd.n1631 gnd 0.147374f
C2766 vdd.t269 gnd 0.033792f
C2767 vdd.t291 gnd 0.033792f
C2768 vdd.n1632 gnd 0.23224f
C2769 vdd.n1633 gnd 0.147374f
C2770 vdd.t250 gnd 0.033792f
C2771 vdd.t162 gnd 0.033792f
C2772 vdd.n1634 gnd 0.23224f
C2773 vdd.n1635 gnd 0.147374f
C2774 vdd.t234 gnd 0.033792f
C2775 vdd.t171 gnd 0.033792f
C2776 vdd.n1636 gnd 0.23224f
C2777 vdd.n1637 gnd 0.147374f
C2778 vdd.t279 gnd 0.033792f
C2779 vdd.t204 gnd 0.033792f
C2780 vdd.n1638 gnd 0.23224f
C2781 vdd.n1639 gnd 0.147374f
C2782 vdd.t256 gnd 0.033792f
C2783 vdd.t225 gnd 0.033792f
C2784 vdd.n1640 gnd 0.23224f
C2785 vdd.n1641 gnd 0.147374f
C2786 vdd.t271 gnd 0.033792f
C2787 vdd.t187 gnd 0.033792f
C2788 vdd.n1642 gnd 0.23224f
C2789 vdd.n1643 gnd 0.147374f
C2790 vdd.t287 gnd 0.033792f
C2791 vdd.t215 gnd 0.033792f
C2792 vdd.n1644 gnd 0.23224f
C2793 vdd.n1645 gnd 0.147374f
C2794 vdd.n1646 gnd 0.00576f
C2795 vdd.n1647 gnd 0.005345f
C2796 vdd.n1648 gnd 0.002957f
C2797 vdd.n1649 gnd 0.006789f
C2798 vdd.n1650 gnd 0.002872f
C2799 vdd.n1651 gnd 0.003041f
C2800 vdd.n1652 gnd 0.005345f
C2801 vdd.n1653 gnd 0.002872f
C2802 vdd.n1654 gnd 0.006789f
C2803 vdd.n1655 gnd 0.003041f
C2804 vdd.n1656 gnd 0.005345f
C2805 vdd.n1657 gnd 0.002872f
C2806 vdd.n1658 gnd 0.005092f
C2807 vdd.n1659 gnd 0.005107f
C2808 vdd.t238 gnd 0.014586f
C2809 vdd.n1660 gnd 0.032453f
C2810 vdd.n1661 gnd 0.168893f
C2811 vdd.n1662 gnd 0.002872f
C2812 vdd.n1663 gnd 0.003041f
C2813 vdd.n1664 gnd 0.006789f
C2814 vdd.n1665 gnd 0.006789f
C2815 vdd.n1666 gnd 0.003041f
C2816 vdd.n1667 gnd 0.002872f
C2817 vdd.n1668 gnd 0.005345f
C2818 vdd.n1669 gnd 0.005345f
C2819 vdd.n1670 gnd 0.002872f
C2820 vdd.n1671 gnd 0.003041f
C2821 vdd.n1672 gnd 0.006789f
C2822 vdd.n1673 gnd 0.006789f
C2823 vdd.n1674 gnd 0.003041f
C2824 vdd.n1675 gnd 0.002872f
C2825 vdd.n1676 gnd 0.005345f
C2826 vdd.n1677 gnd 0.005345f
C2827 vdd.n1678 gnd 0.002872f
C2828 vdd.n1679 gnd 0.003041f
C2829 vdd.n1680 gnd 0.006789f
C2830 vdd.n1681 gnd 0.006789f
C2831 vdd.n1682 gnd 0.016051f
C2832 vdd.n1683 gnd 0.002957f
C2833 vdd.n1684 gnd 0.002872f
C2834 vdd.n1685 gnd 0.013816f
C2835 vdd.n1686 gnd 0.009343f
C2836 vdd.n1687 gnd 0.109647f
C2837 vdd.n1688 gnd 0.00576f
C2838 vdd.n1689 gnd 0.005345f
C2839 vdd.n1690 gnd 0.002957f
C2840 vdd.n1691 gnd 0.006789f
C2841 vdd.n1692 gnd 0.002872f
C2842 vdd.n1693 gnd 0.003041f
C2843 vdd.n1694 gnd 0.005345f
C2844 vdd.n1695 gnd 0.002872f
C2845 vdd.n1696 gnd 0.006789f
C2846 vdd.n1697 gnd 0.003041f
C2847 vdd.n1698 gnd 0.005345f
C2848 vdd.n1699 gnd 0.002872f
C2849 vdd.n1700 gnd 0.005092f
C2850 vdd.n1701 gnd 0.005107f
C2851 vdd.t280 gnd 0.014586f
C2852 vdd.n1702 gnd 0.032453f
C2853 vdd.n1703 gnd 0.168893f
C2854 vdd.n1704 gnd 0.002872f
C2855 vdd.n1705 gnd 0.003041f
C2856 vdd.n1706 gnd 0.006789f
C2857 vdd.n1707 gnd 0.006789f
C2858 vdd.n1708 gnd 0.003041f
C2859 vdd.n1709 gnd 0.002872f
C2860 vdd.n1710 gnd 0.005345f
C2861 vdd.n1711 gnd 0.005345f
C2862 vdd.n1712 gnd 0.002872f
C2863 vdd.n1713 gnd 0.003041f
C2864 vdd.n1714 gnd 0.006789f
C2865 vdd.n1715 gnd 0.006789f
C2866 vdd.n1716 gnd 0.003041f
C2867 vdd.n1717 gnd 0.002872f
C2868 vdd.n1718 gnd 0.005345f
C2869 vdd.n1719 gnd 0.005345f
C2870 vdd.n1720 gnd 0.002872f
C2871 vdd.n1721 gnd 0.003041f
C2872 vdd.n1722 gnd 0.006789f
C2873 vdd.n1723 gnd 0.006789f
C2874 vdd.n1724 gnd 0.016051f
C2875 vdd.n1725 gnd 0.002957f
C2876 vdd.n1726 gnd 0.002872f
C2877 vdd.n1727 gnd 0.013816f
C2878 vdd.n1728 gnd 0.009645f
C2879 vdd.t244 gnd 0.033792f
C2880 vdd.t178 gnd 0.033792f
C2881 vdd.n1729 gnd 0.23224f
C2882 vdd.n1730 gnd 0.182621f
C2883 vdd.t174 gnd 0.033792f
C2884 vdd.t247 gnd 0.033792f
C2885 vdd.n1731 gnd 0.23224f
C2886 vdd.n1732 gnd 0.147374f
C2887 vdd.t231 gnd 0.033792f
C2888 vdd.t227 gnd 0.033792f
C2889 vdd.n1733 gnd 0.23224f
C2890 vdd.n1734 gnd 0.147374f
C2891 vdd.t169 gnd 0.033792f
C2892 vdd.t144 gnd 0.033792f
C2893 vdd.n1735 gnd 0.23224f
C2894 vdd.n1736 gnd 0.147374f
C2895 vdd.t136 gnd 0.033792f
C2896 vdd.t222 gnd 0.033792f
C2897 vdd.n1737 gnd 0.23224f
C2898 vdd.n1738 gnd 0.147374f
C2899 vdd.t199 gnd 0.033792f
C2900 vdd.t140 gnd 0.033792f
C2901 vdd.n1739 gnd 0.23224f
C2902 vdd.n1740 gnd 0.147374f
C2903 vdd.t134 gnd 0.033792f
C2904 vdd.t251 gnd 0.033792f
C2905 vdd.n1741 gnd 0.23224f
C2906 vdd.n1742 gnd 0.147374f
C2907 vdd.t246 gnd 0.033792f
C2908 vdd.t189 gnd 0.033792f
C2909 vdd.n1743 gnd 0.23224f
C2910 vdd.n1744 gnd 0.147374f
C2911 vdd.t176 gnd 0.033792f
C2912 vdd.t276 gnd 0.033792f
C2913 vdd.n1745 gnd 0.23224f
C2914 vdd.n1746 gnd 0.147374f
C2915 vdd.n1747 gnd 0.00576f
C2916 vdd.n1748 gnd 0.005345f
C2917 vdd.n1749 gnd 0.002957f
C2918 vdd.n1750 gnd 0.006789f
C2919 vdd.n1751 gnd 0.002872f
C2920 vdd.n1752 gnd 0.003041f
C2921 vdd.n1753 gnd 0.005345f
C2922 vdd.n1754 gnd 0.002872f
C2923 vdd.n1755 gnd 0.006789f
C2924 vdd.n1756 gnd 0.003041f
C2925 vdd.n1757 gnd 0.005345f
C2926 vdd.n1758 gnd 0.002872f
C2927 vdd.n1759 gnd 0.005092f
C2928 vdd.n1760 gnd 0.005107f
C2929 vdd.t229 gnd 0.014586f
C2930 vdd.n1761 gnd 0.032453f
C2931 vdd.n1762 gnd 0.168893f
C2932 vdd.n1763 gnd 0.002872f
C2933 vdd.n1764 gnd 0.003041f
C2934 vdd.n1765 gnd 0.006789f
C2935 vdd.n1766 gnd 0.006789f
C2936 vdd.n1767 gnd 0.003041f
C2937 vdd.n1768 gnd 0.002872f
C2938 vdd.n1769 gnd 0.005345f
C2939 vdd.n1770 gnd 0.005345f
C2940 vdd.n1771 gnd 0.002872f
C2941 vdd.n1772 gnd 0.003041f
C2942 vdd.n1773 gnd 0.006789f
C2943 vdd.n1774 gnd 0.006789f
C2944 vdd.n1775 gnd 0.003041f
C2945 vdd.n1776 gnd 0.002872f
C2946 vdd.n1777 gnd 0.005345f
C2947 vdd.n1778 gnd 0.005345f
C2948 vdd.n1779 gnd 0.002872f
C2949 vdd.n1780 gnd 0.003041f
C2950 vdd.n1781 gnd 0.006789f
C2951 vdd.n1782 gnd 0.006789f
C2952 vdd.n1783 gnd 0.016051f
C2953 vdd.n1784 gnd 0.002957f
C2954 vdd.n1785 gnd 0.002872f
C2955 vdd.n1786 gnd 0.013816f
C2956 vdd.n1787 gnd 0.009343f
C2957 vdd.n1788 gnd 0.065229f
C2958 vdd.n1789 gnd 0.235038f
C2959 vdd.n1790 gnd 0.00576f
C2960 vdd.n1791 gnd 0.005345f
C2961 vdd.n1792 gnd 0.002957f
C2962 vdd.n1793 gnd 0.006789f
C2963 vdd.n1794 gnd 0.002872f
C2964 vdd.n1795 gnd 0.003041f
C2965 vdd.n1796 gnd 0.005345f
C2966 vdd.n1797 gnd 0.002872f
C2967 vdd.n1798 gnd 0.006789f
C2968 vdd.n1799 gnd 0.003041f
C2969 vdd.n1800 gnd 0.005345f
C2970 vdd.n1801 gnd 0.002872f
C2971 vdd.n1802 gnd 0.005092f
C2972 vdd.n1803 gnd 0.005107f
C2973 vdd.t292 gnd 0.014586f
C2974 vdd.n1804 gnd 0.032453f
C2975 vdd.n1805 gnd 0.168893f
C2976 vdd.n1806 gnd 0.002872f
C2977 vdd.n1807 gnd 0.003041f
C2978 vdd.n1808 gnd 0.006789f
C2979 vdd.n1809 gnd 0.006789f
C2980 vdd.n1810 gnd 0.003041f
C2981 vdd.n1811 gnd 0.002872f
C2982 vdd.n1812 gnd 0.005345f
C2983 vdd.n1813 gnd 0.005345f
C2984 vdd.n1814 gnd 0.002872f
C2985 vdd.n1815 gnd 0.003041f
C2986 vdd.n1816 gnd 0.006789f
C2987 vdd.n1817 gnd 0.006789f
C2988 vdd.n1818 gnd 0.003041f
C2989 vdd.n1819 gnd 0.002872f
C2990 vdd.n1820 gnd 0.005345f
C2991 vdd.n1821 gnd 0.005345f
C2992 vdd.n1822 gnd 0.002872f
C2993 vdd.n1823 gnd 0.003041f
C2994 vdd.n1824 gnd 0.006789f
C2995 vdd.n1825 gnd 0.006789f
C2996 vdd.n1826 gnd 0.016051f
C2997 vdd.n1827 gnd 0.002957f
C2998 vdd.n1828 gnd 0.002872f
C2999 vdd.n1829 gnd 0.013816f
C3000 vdd.n1830 gnd 0.009645f
C3001 vdd.t258 gnd 0.033792f
C3002 vdd.t205 gnd 0.033792f
C3003 vdd.n1831 gnd 0.23224f
C3004 vdd.n1832 gnd 0.182621f
C3005 vdd.t200 gnd 0.033792f
C3006 vdd.t260 gnd 0.033792f
C3007 vdd.n1833 gnd 0.23224f
C3008 vdd.n1834 gnd 0.147374f
C3009 vdd.t242 gnd 0.033792f
C3010 vdd.t240 gnd 0.033792f
C3011 vdd.n1835 gnd 0.23224f
C3012 vdd.n1836 gnd 0.147374f
C3013 vdd.t195 gnd 0.033792f
C3014 vdd.t165 gnd 0.033792f
C3015 vdd.n1837 gnd 0.23224f
C3016 vdd.n1838 gnd 0.147374f
C3017 vdd.t163 gnd 0.033792f
C3018 vdd.t239 gnd 0.033792f
C3019 vdd.n1839 gnd 0.23224f
C3020 vdd.n1840 gnd 0.147374f
C3021 vdd.t216 gnd 0.033792f
C3022 vdd.t164 gnd 0.033792f
C3023 vdd.n1841 gnd 0.23224f
C3024 vdd.n1842 gnd 0.147374f
C3025 vdd.t157 gnd 0.033792f
C3026 vdd.t261 gnd 0.033792f
C3027 vdd.n1843 gnd 0.23224f
C3028 vdd.n1844 gnd 0.147374f
C3029 vdd.t259 gnd 0.033792f
C3030 vdd.t209 gnd 0.033792f
C3031 vdd.n1845 gnd 0.23224f
C3032 vdd.n1846 gnd 0.147374f
C3033 vdd.t201 gnd 0.033792f
C3034 vdd.t288 gnd 0.033792f
C3035 vdd.n1847 gnd 0.23224f
C3036 vdd.n1848 gnd 0.147374f
C3037 vdd.n1849 gnd 0.00576f
C3038 vdd.n1850 gnd 0.005345f
C3039 vdd.n1851 gnd 0.002957f
C3040 vdd.n1852 gnd 0.006789f
C3041 vdd.n1853 gnd 0.002872f
C3042 vdd.n1854 gnd 0.003041f
C3043 vdd.n1855 gnd 0.005345f
C3044 vdd.n1856 gnd 0.002872f
C3045 vdd.n1857 gnd 0.006789f
C3046 vdd.n1858 gnd 0.003041f
C3047 vdd.n1859 gnd 0.005345f
C3048 vdd.n1860 gnd 0.002872f
C3049 vdd.n1861 gnd 0.005092f
C3050 vdd.n1862 gnd 0.005107f
C3051 vdd.t241 gnd 0.014586f
C3052 vdd.n1863 gnd 0.032453f
C3053 vdd.n1864 gnd 0.168893f
C3054 vdd.n1865 gnd 0.002872f
C3055 vdd.n1866 gnd 0.003041f
C3056 vdd.n1867 gnd 0.006789f
C3057 vdd.n1868 gnd 0.006789f
C3058 vdd.n1869 gnd 0.003041f
C3059 vdd.n1870 gnd 0.002872f
C3060 vdd.n1871 gnd 0.005345f
C3061 vdd.n1872 gnd 0.005345f
C3062 vdd.n1873 gnd 0.002872f
C3063 vdd.n1874 gnd 0.003041f
C3064 vdd.n1875 gnd 0.006789f
C3065 vdd.n1876 gnd 0.006789f
C3066 vdd.n1877 gnd 0.003041f
C3067 vdd.n1878 gnd 0.002872f
C3068 vdd.n1879 gnd 0.005345f
C3069 vdd.n1880 gnd 0.005345f
C3070 vdd.n1881 gnd 0.002872f
C3071 vdd.n1882 gnd 0.003041f
C3072 vdd.n1883 gnd 0.006789f
C3073 vdd.n1884 gnd 0.006789f
C3074 vdd.n1885 gnd 0.016051f
C3075 vdd.n1886 gnd 0.002957f
C3076 vdd.n1887 gnd 0.002872f
C3077 vdd.n1888 gnd 0.013816f
C3078 vdd.n1889 gnd 0.009343f
C3079 vdd.n1890 gnd 0.065229f
C3080 vdd.n1891 gnd 0.269067f
C3081 vdd.n1892 gnd 2.94957f
C3082 vdd.n1893 gnd 0.619089f
C3083 vdd.n1894 gnd 0.008067f
C3084 vdd.n1895 gnd 0.008448f
C3085 vdd.n1896 gnd 0.010496f
C3086 vdd.n1897 gnd 0.766932f
C3087 vdd.n1898 gnd 0.010496f
C3088 vdd.n1899 gnd 0.008448f
C3089 vdd.n1900 gnd 0.010496f
C3090 vdd.n1901 gnd 0.010496f
C3091 vdd.n1902 gnd 0.010496f
C3092 vdd.n1903 gnd 0.008448f
C3093 vdd.n1904 gnd 0.010496f
C3094 vdd.n1905 gnd 0.890285f
C3095 vdd.t168 gnd 0.536316f
C3096 vdd.n1906 gnd 0.584585f
C3097 vdd.n1907 gnd 0.010496f
C3098 vdd.n1908 gnd 0.008448f
C3099 vdd.n1909 gnd 0.010496f
C3100 vdd.n1910 gnd 0.010496f
C3101 vdd.n1911 gnd 0.010496f
C3102 vdd.n1912 gnd 0.008448f
C3103 vdd.n1913 gnd 0.010496f
C3104 vdd.n1914 gnd 0.670395f
C3105 vdd.n1915 gnd 0.010496f
C3106 vdd.n1916 gnd 0.008448f
C3107 vdd.n1917 gnd 0.010496f
C3108 vdd.n1918 gnd 0.010496f
C3109 vdd.n1919 gnd 0.010496f
C3110 vdd.n1920 gnd 0.008448f
C3111 vdd.n1921 gnd 0.010496f
C3112 vdd.n1922 gnd 0.573858f
C3113 vdd.n1923 gnd 0.852743f
C3114 vdd.n1924 gnd 0.010496f
C3115 vdd.n1925 gnd 0.008448f
C3116 vdd.n1926 gnd 0.010496f
C3117 vdd.n1927 gnd 0.010496f
C3118 vdd.n1928 gnd 0.010496f
C3119 vdd.n1929 gnd 0.008448f
C3120 vdd.n1930 gnd 0.010496f
C3121 vdd.n1931 gnd 0.890285f
C3122 vdd.n1932 gnd 0.010496f
C3123 vdd.n1933 gnd 0.008448f
C3124 vdd.n1934 gnd 0.010496f
C3125 vdd.n1935 gnd 0.010496f
C3126 vdd.n1936 gnd 0.010496f
C3127 vdd.n1937 gnd 0.008448f
C3128 vdd.n1938 gnd 0.010496f
C3129 vdd.t158 gnd 0.536316f
C3130 vdd.n1939 gnd 0.745479f
C3131 vdd.n1940 gnd 0.010496f
C3132 vdd.n1941 gnd 0.008448f
C3133 vdd.n1942 gnd 0.010496f
C3134 vdd.n1943 gnd 0.010496f
C3135 vdd.n1944 gnd 0.010496f
C3136 vdd.n1945 gnd 0.008448f
C3137 vdd.n1946 gnd 0.010496f
C3138 vdd.n1947 gnd 0.563132f
C3139 vdd.n1948 gnd 0.010496f
C3140 vdd.n1949 gnd 0.008448f
C3141 vdd.n1950 gnd 0.010496f
C3142 vdd.n1951 gnd 0.010496f
C3143 vdd.n1952 gnd 0.010496f
C3144 vdd.n1953 gnd 0.008448f
C3145 vdd.n1954 gnd 0.010496f
C3146 vdd.n1955 gnd 0.734753f
C3147 vdd.n1956 gnd 0.691848f
C3148 vdd.n1957 gnd 0.010496f
C3149 vdd.n1958 gnd 0.008448f
C3150 vdd.n1959 gnd 0.010496f
C3151 vdd.n1960 gnd 0.010496f
C3152 vdd.n1961 gnd 0.010496f
C3153 vdd.n1962 gnd 0.008448f
C3154 vdd.n1963 gnd 0.010496f
C3155 vdd.n1964 gnd 0.874195f
C3156 vdd.n1965 gnd 0.010496f
C3157 vdd.n1966 gnd 0.008448f
C3158 vdd.n1967 gnd 0.010496f
C3159 vdd.n1968 gnd 0.010496f
C3160 vdd.n1969 gnd 0.02539f
C3161 vdd.n1970 gnd 0.010496f
C3162 vdd.n1971 gnd 0.010496f
C3163 vdd.n1972 gnd 0.008448f
C3164 vdd.n1973 gnd 0.010496f
C3165 vdd.n1974 gnd 0.648942f
C3166 vdd.n1975 gnd 1.07263f
C3167 vdd.n1976 gnd 0.010496f
C3168 vdd.n1977 gnd 0.008448f
C3169 vdd.n1978 gnd 0.010496f
C3170 vdd.n1979 gnd 0.010496f
C3171 vdd.n1980 gnd 0.009026f
C3172 vdd.n1981 gnd 0.008448f
C3173 vdd.n1983 gnd 0.010496f
C3174 vdd.n1985 gnd 0.008448f
C3175 vdd.n1986 gnd 0.010496f
C3176 vdd.n1987 gnd 0.008448f
C3177 vdd.n1989 gnd 0.010496f
C3178 vdd.n1990 gnd 0.008448f
C3179 vdd.n1991 gnd 0.010496f
C3180 vdd.n1992 gnd 0.010496f
C3181 vdd.n1993 gnd 0.010496f
C3182 vdd.n1994 gnd 0.010496f
C3183 vdd.n1995 gnd 0.010496f
C3184 vdd.n1996 gnd 0.008448f
C3185 vdd.n1998 gnd 0.010496f
C3186 vdd.n1999 gnd 0.010496f
C3187 vdd.n2000 gnd 0.010496f
C3188 vdd.n2001 gnd 0.010496f
C3189 vdd.n2002 gnd 0.010496f
C3190 vdd.n2003 gnd 0.008448f
C3191 vdd.n2005 gnd 0.010496f
C3192 vdd.n2006 gnd 0.010496f
C3193 vdd.n2007 gnd 0.010496f
C3194 vdd.n2008 gnd 0.010496f
C3195 vdd.n2009 gnd 0.007054f
C3196 vdd.t116 gnd 0.129127f
C3197 vdd.t115 gnd 0.138001f
C3198 vdd.t114 gnd 0.168639f
C3199 vdd.n2010 gnd 0.216171f
C3200 vdd.n2011 gnd 0.181623f
C3201 vdd.n2013 gnd 0.010496f
C3202 vdd.n2014 gnd 0.010496f
C3203 vdd.n2015 gnd 0.008448f
C3204 vdd.n2016 gnd 0.010496f
C3205 vdd.n2018 gnd 0.010496f
C3206 vdd.n2019 gnd 0.010496f
C3207 vdd.n2020 gnd 0.010496f
C3208 vdd.n2021 gnd 0.010496f
C3209 vdd.n2022 gnd 0.008448f
C3210 vdd.n2024 gnd 0.010496f
C3211 vdd.n2025 gnd 0.010496f
C3212 vdd.n2026 gnd 0.010496f
C3213 vdd.n2027 gnd 0.010496f
C3214 vdd.n2028 gnd 0.010496f
C3215 vdd.n2029 gnd 0.008448f
C3216 vdd.n2031 gnd 0.010496f
C3217 vdd.n2032 gnd 0.010496f
C3218 vdd.n2033 gnd 0.010496f
C3219 vdd.n2034 gnd 0.010496f
C3220 vdd.n2035 gnd 0.010496f
C3221 vdd.n2036 gnd 0.008448f
C3222 vdd.n2038 gnd 0.010496f
C3223 vdd.n2039 gnd 0.010496f
C3224 vdd.n2040 gnd 0.010496f
C3225 vdd.n2041 gnd 0.010496f
C3226 vdd.n2042 gnd 0.010496f
C3227 vdd.n2043 gnd 0.008448f
C3228 vdd.n2045 gnd 0.010496f
C3229 vdd.n2046 gnd 0.010496f
C3230 vdd.n2047 gnd 0.010496f
C3231 vdd.n2048 gnd 0.010496f
C3232 vdd.n2049 gnd 0.008363f
C3233 vdd.t95 gnd 0.129127f
C3234 vdd.t94 gnd 0.138001f
C3235 vdd.t93 gnd 0.168639f
C3236 vdd.n2050 gnd 0.216171f
C3237 vdd.n2051 gnd 0.181623f
C3238 vdd.n2053 gnd 0.010496f
C3239 vdd.n2054 gnd 0.010496f
C3240 vdd.n2055 gnd 0.008448f
C3241 vdd.n2056 gnd 0.010496f
C3242 vdd.n2058 gnd 0.010496f
C3243 vdd.n2059 gnd 0.010496f
C3244 vdd.n2060 gnd 0.010496f
C3245 vdd.n2061 gnd 0.010496f
C3246 vdd.n2062 gnd 0.008448f
C3247 vdd.n2064 gnd 0.010496f
C3248 vdd.n2065 gnd 0.010496f
C3249 vdd.n2066 gnd 0.010496f
C3250 vdd.n2067 gnd 0.010496f
C3251 vdd.n2068 gnd 0.010496f
C3252 vdd.n2069 gnd 0.008448f
C3253 vdd.n2071 gnd 0.010496f
C3254 vdd.n2072 gnd 0.010496f
C3255 vdd.n2073 gnd 0.010496f
C3256 vdd.n2074 gnd 0.010496f
C3257 vdd.n2075 gnd 0.010496f
C3258 vdd.n2076 gnd 0.010496f
C3259 vdd.n2077 gnd 0.008448f
C3260 vdd.n2079 gnd 0.010496f
C3261 vdd.n2081 gnd 0.010496f
C3262 vdd.n2082 gnd 0.008448f
C3263 vdd.n2083 gnd 0.008448f
C3264 vdd.n2084 gnd 0.010496f
C3265 vdd.n2086 gnd 0.010496f
C3266 vdd.n2087 gnd 0.008448f
C3267 vdd.n2088 gnd 0.008448f
C3268 vdd.n2089 gnd 0.010496f
C3269 vdd.n2091 gnd 0.010496f
C3270 vdd.n2092 gnd 0.010496f
C3271 vdd.n2093 gnd 0.008448f
C3272 vdd.n2094 gnd 0.008448f
C3273 vdd.n2095 gnd 0.008448f
C3274 vdd.n2096 gnd 0.010496f
C3275 vdd.n2098 gnd 0.010496f
C3276 vdd.n2099 gnd 0.010496f
C3277 vdd.n2100 gnd 0.008448f
C3278 vdd.n2101 gnd 0.008448f
C3279 vdd.n2102 gnd 0.008448f
C3280 vdd.n2103 gnd 0.010496f
C3281 vdd.n2105 gnd 0.010496f
C3282 vdd.n2106 gnd 0.010496f
C3283 vdd.n2107 gnd 0.008448f
C3284 vdd.n2108 gnd 0.008448f
C3285 vdd.n2109 gnd 0.008448f
C3286 vdd.n2110 gnd 0.010496f
C3287 vdd.n2112 gnd 0.010496f
C3288 vdd.n2113 gnd 0.010496f
C3289 vdd.n2114 gnd 0.008448f
C3290 vdd.n2115 gnd 0.010496f
C3291 vdd.n2116 gnd 0.010496f
C3292 vdd.n2117 gnd 0.010496f
C3293 vdd.n2118 gnd 0.017234f
C3294 vdd.n2119 gnd 0.005745f
C3295 vdd.n2120 gnd 0.008448f
C3296 vdd.n2121 gnd 0.010496f
C3297 vdd.n2123 gnd 0.010496f
C3298 vdd.n2124 gnd 0.010496f
C3299 vdd.n2125 gnd 0.008448f
C3300 vdd.n2126 gnd 0.008448f
C3301 vdd.n2127 gnd 0.008448f
C3302 vdd.n2128 gnd 0.010496f
C3303 vdd.n2130 gnd 0.010496f
C3304 vdd.n2131 gnd 0.010496f
C3305 vdd.n2132 gnd 0.008448f
C3306 vdd.n2133 gnd 0.008448f
C3307 vdd.n2134 gnd 0.008448f
C3308 vdd.n2135 gnd 0.010496f
C3309 vdd.n2137 gnd 0.010496f
C3310 vdd.n2138 gnd 0.010496f
C3311 vdd.n2139 gnd 0.008448f
C3312 vdd.n2140 gnd 0.008448f
C3313 vdd.n2141 gnd 0.008448f
C3314 vdd.n2142 gnd 0.010496f
C3315 vdd.n2144 gnd 0.010496f
C3316 vdd.n2145 gnd 0.010496f
C3317 vdd.n2146 gnd 0.008448f
C3318 vdd.n2147 gnd 0.008448f
C3319 vdd.n2148 gnd 0.008448f
C3320 vdd.n2149 gnd 0.010496f
C3321 vdd.n2151 gnd 0.010496f
C3322 vdd.n2152 gnd 0.010496f
C3323 vdd.n2153 gnd 0.008448f
C3324 vdd.n2154 gnd 0.010496f
C3325 vdd.n2155 gnd 0.010496f
C3326 vdd.n2156 gnd 0.010496f
C3327 vdd.n2157 gnd 0.017234f
C3328 vdd.n2158 gnd 0.007054f
C3329 vdd.n2159 gnd 0.008448f
C3330 vdd.n2160 gnd 0.010496f
C3331 vdd.n2162 gnd 0.010496f
C3332 vdd.n2163 gnd 0.010496f
C3333 vdd.n2164 gnd 0.008448f
C3334 vdd.n2165 gnd 0.008448f
C3335 vdd.n2166 gnd 0.008448f
C3336 vdd.n2167 gnd 0.010496f
C3337 vdd.n2169 gnd 0.010496f
C3338 vdd.n2170 gnd 0.010496f
C3339 vdd.n2171 gnd 0.008448f
C3340 vdd.n2172 gnd 0.008448f
C3341 vdd.n2173 gnd 0.008448f
C3342 vdd.n2174 gnd 0.010496f
C3343 vdd.n2176 gnd 0.010496f
C3344 vdd.n2177 gnd 0.010496f
C3345 vdd.n2179 gnd 0.010496f
C3346 vdd.n2180 gnd 0.008448f
C3347 vdd.n2181 gnd 0.006717f
C3348 vdd.n2182 gnd 0.954793f
C3349 vdd.n2184 gnd 0.008448f
C3350 vdd.n2185 gnd 0.008448f
C3351 vdd.n2186 gnd 0.010496f
C3352 vdd.n2188 gnd 0.010496f
C3353 vdd.n2189 gnd 0.010496f
C3354 vdd.n2190 gnd 0.008448f
C3355 vdd.n2191 gnd 0.007012f
C3356 vdd.n2192 gnd 0.025935f
C3357 vdd.n2193 gnd 0.02539f
C3358 vdd.n2194 gnd 0.007012f
C3359 vdd.n2195 gnd 0.02539f
C3360 vdd.n2196 gnd 1.47487f
C3361 vdd.n2197 gnd 0.02539f
C3362 vdd.n2198 gnd 0.025935f
C3363 vdd.n2199 gnd 0.004013f
C3364 vdd.t86 gnd 0.129127f
C3365 vdd.t85 gnd 0.138001f
C3366 vdd.t83 gnd 0.168639f
C3367 vdd.n2200 gnd 0.216171f
C3368 vdd.n2201 gnd 0.181623f
C3369 vdd.n2202 gnd 0.01301f
C3370 vdd.n2203 gnd 0.004435f
C3371 vdd.n2204 gnd 0.009026f
C3372 vdd.n2205 gnd 0.954793f
C3373 vdd.n2206 gnd 0.037553f
C3374 vdd.n2207 gnd 0.007137f
C3375 vdd.n2208 gnd 0.007137f
C3376 vdd.n2209 gnd 0.007137f
C3377 vdd.n2210 gnd 0.007137f
C3378 vdd.n2211 gnd 0.007137f
C3379 vdd.n2212 gnd 0.007137f
C3380 vdd.n2213 gnd 0.007137f
C3381 vdd.n2214 gnd 0.007137f
C3382 vdd.n2216 gnd 0.007137f
C3383 vdd.n2218 gnd 0.007137f
C3384 vdd.n2219 gnd 0.007137f
C3385 vdd.n2220 gnd 0.007137f
C3386 vdd.n2221 gnd 0.007137f
C3387 vdd.n2222 gnd 0.007137f
C3388 vdd.n2224 gnd 0.007137f
C3389 vdd.n2226 gnd 0.007137f
C3390 vdd.n2227 gnd 0.007137f
C3391 vdd.n2228 gnd 0.007137f
C3392 vdd.n2229 gnd 0.007137f
C3393 vdd.n2230 gnd 0.007137f
C3394 vdd.n2232 gnd 0.007137f
C3395 vdd.n2234 gnd 0.007137f
C3396 vdd.n2235 gnd 0.007137f
C3397 vdd.n2236 gnd 0.007137f
C3398 vdd.n2237 gnd 0.007137f
C3399 vdd.n2238 gnd 0.007137f
C3400 vdd.n2240 gnd 0.007137f
C3401 vdd.n2242 gnd 0.007137f
C3402 vdd.n2243 gnd 0.007137f
C3403 vdd.n2244 gnd 0.007137f
C3404 vdd.n2245 gnd 0.007137f
C3405 vdd.n2246 gnd 0.007137f
C3406 vdd.n2248 gnd 0.007137f
C3407 vdd.n2250 gnd 0.007137f
C3408 vdd.n2251 gnd 0.007137f
C3409 vdd.n2252 gnd 0.007137f
C3410 vdd.n2253 gnd 0.007137f
C3411 vdd.n2254 gnd 0.007137f
C3412 vdd.n2256 gnd 0.007137f
C3413 vdd.n2258 gnd 0.007137f
C3414 vdd.n2259 gnd 0.007137f
C3415 vdd.n2260 gnd 0.007137f
C3416 vdd.n2261 gnd 0.007137f
C3417 vdd.n2262 gnd 0.007137f
C3418 vdd.n2264 gnd 0.007137f
C3419 vdd.n2266 gnd 0.007137f
C3420 vdd.n2267 gnd 0.007137f
C3421 vdd.n2268 gnd 0.007137f
C3422 vdd.n2269 gnd 0.007137f
C3423 vdd.n2270 gnd 0.007137f
C3424 vdd.n2272 gnd 0.007137f
C3425 vdd.n2274 gnd 0.007137f
C3426 vdd.n2275 gnd 0.007137f
C3427 vdd.n2276 gnd 0.005195f
C3428 vdd.n2277 gnd 0.0102f
C3429 vdd.n2278 gnd 0.00551f
C3430 vdd.n2279 gnd 0.007137f
C3431 vdd.n2281 gnd 0.007137f
C3432 vdd.n2282 gnd 0.01645f
C3433 vdd.n2283 gnd 0.01645f
C3434 vdd.n2284 gnd 0.015457f
C3435 vdd.n2285 gnd 0.007137f
C3436 vdd.n2286 gnd 0.007137f
C3437 vdd.n2287 gnd 0.007137f
C3438 vdd.n2288 gnd 0.007137f
C3439 vdd.n2289 gnd 0.007137f
C3440 vdd.n2290 gnd 0.007137f
C3441 vdd.n2291 gnd 0.007137f
C3442 vdd.n2292 gnd 0.007137f
C3443 vdd.n2293 gnd 0.007137f
C3444 vdd.n2294 gnd 0.007137f
C3445 vdd.n2295 gnd 0.007137f
C3446 vdd.n2296 gnd 0.007137f
C3447 vdd.n2297 gnd 0.007137f
C3448 vdd.n2298 gnd 0.007137f
C3449 vdd.n2299 gnd 0.007137f
C3450 vdd.n2300 gnd 0.007137f
C3451 vdd.n2301 gnd 0.007137f
C3452 vdd.n2302 gnd 0.007137f
C3453 vdd.n2303 gnd 0.007137f
C3454 vdd.n2304 gnd 0.007137f
C3455 vdd.n2305 gnd 0.007137f
C3456 vdd.n2306 gnd 0.007137f
C3457 vdd.n2307 gnd 0.007137f
C3458 vdd.n2308 gnd 0.007137f
C3459 vdd.n2309 gnd 0.007137f
C3460 vdd.n2310 gnd 0.007137f
C3461 vdd.n2311 gnd 0.007137f
C3462 vdd.n2312 gnd 0.007137f
C3463 vdd.n2313 gnd 0.007137f
C3464 vdd.n2314 gnd 0.007137f
C3465 vdd.n2315 gnd 0.007137f
C3466 vdd.n2316 gnd 0.007137f
C3467 vdd.n2317 gnd 0.007137f
C3468 vdd.n2318 gnd 0.007137f
C3469 vdd.n2319 gnd 0.007137f
C3470 vdd.n2320 gnd 0.007137f
C3471 vdd.n2321 gnd 0.007137f
C3472 vdd.n2322 gnd 0.007137f
C3473 vdd.n2323 gnd 0.007137f
C3474 vdd.n2324 gnd 0.007137f
C3475 vdd.n2325 gnd 0.007137f
C3476 vdd.n2326 gnd 0.007137f
C3477 vdd.n2327 gnd 0.007137f
C3478 vdd.n2328 gnd 0.007137f
C3479 vdd.n2329 gnd 0.007137f
C3480 vdd.n2330 gnd 0.007137f
C3481 vdd.n2331 gnd 0.007137f
C3482 vdd.n2332 gnd 0.007137f
C3483 vdd.n2333 gnd 0.007137f
C3484 vdd.n2334 gnd 0.434416f
C3485 vdd.n2335 gnd 0.007137f
C3486 vdd.n2336 gnd 0.007137f
C3487 vdd.n2337 gnd 0.007137f
C3488 vdd.n2338 gnd 0.007137f
C3489 vdd.n2339 gnd 0.007137f
C3490 vdd.n2340 gnd 0.007137f
C3491 vdd.n2341 gnd 0.007137f
C3492 vdd.n2342 gnd 0.007137f
C3493 vdd.n2343 gnd 0.007137f
C3494 vdd.n2344 gnd 0.007137f
C3495 vdd.n2345 gnd 0.007137f
C3496 vdd.n2346 gnd 0.659669f
C3497 vdd.n2347 gnd 0.007137f
C3498 vdd.n2348 gnd 0.007137f
C3499 vdd.n2349 gnd 0.007137f
C3500 vdd.n2350 gnd 0.007137f
C3501 vdd.n2351 gnd 0.007137f
C3502 vdd.n2352 gnd 0.007137f
C3503 vdd.n2353 gnd 0.007137f
C3504 vdd.n2354 gnd 0.007137f
C3505 vdd.n2355 gnd 0.007137f
C3506 vdd.n2356 gnd 0.007137f
C3507 vdd.n2357 gnd 0.007137f
C3508 vdd.n2358 gnd 0.230616f
C3509 vdd.n2359 gnd 0.007137f
C3510 vdd.n2360 gnd 0.007137f
C3511 vdd.n2361 gnd 0.007137f
C3512 vdd.n2362 gnd 0.007137f
C3513 vdd.n2363 gnd 0.007137f
C3514 vdd.n2364 gnd 0.007137f
C3515 vdd.n2365 gnd 0.007137f
C3516 vdd.n2366 gnd 0.007137f
C3517 vdd.n2367 gnd 0.007137f
C3518 vdd.n2368 gnd 0.007137f
C3519 vdd.n2369 gnd 0.007137f
C3520 vdd.n2370 gnd 0.007137f
C3521 vdd.n2371 gnd 0.007137f
C3522 vdd.n2372 gnd 0.007137f
C3523 vdd.n2373 gnd 0.007137f
C3524 vdd.n2374 gnd 0.007137f
C3525 vdd.n2375 gnd 0.007137f
C3526 vdd.n2376 gnd 0.007137f
C3527 vdd.n2377 gnd 0.007137f
C3528 vdd.n2378 gnd 0.007137f
C3529 vdd.n2379 gnd 0.007137f
C3530 vdd.n2380 gnd 0.007137f
C3531 vdd.n2381 gnd 0.007137f
C3532 vdd.n2382 gnd 0.007137f
C3533 vdd.n2383 gnd 0.007137f
C3534 vdd.n2384 gnd 0.007137f
C3535 vdd.n2385 gnd 0.007137f
C3536 vdd.n2386 gnd 0.007137f
C3537 vdd.n2387 gnd 0.007137f
C3538 vdd.n2388 gnd 0.007137f
C3539 vdd.n2389 gnd 0.007137f
C3540 vdd.n2390 gnd 0.007137f
C3541 vdd.n2391 gnd 0.007137f
C3542 vdd.n2392 gnd 0.007137f
C3543 vdd.n2393 gnd 0.007137f
C3544 vdd.n2394 gnd 0.015457f
C3545 vdd.n2395 gnd 0.01645f
C3546 vdd.n2396 gnd 0.01645f
C3547 vdd.n2398 gnd 0.007137f
C3548 vdd.n2400 gnd 0.007137f
C3549 vdd.n2401 gnd 0.00551f
C3550 vdd.n2402 gnd 0.0102f
C3551 vdd.n2403 gnd 0.005195f
C3552 vdd.n2404 gnd 0.007137f
C3553 vdd.n2405 gnd 0.007137f
C3554 vdd.n2407 gnd 0.007137f
C3555 vdd.n2409 gnd 0.007137f
C3556 vdd.n2410 gnd 0.007137f
C3557 vdd.n2411 gnd 0.007137f
C3558 vdd.n2412 gnd 0.007137f
C3559 vdd.n2413 gnd 0.007137f
C3560 vdd.n2415 gnd 0.007137f
C3561 vdd.n2417 gnd 0.007137f
C3562 vdd.n2418 gnd 0.007137f
C3563 vdd.n2419 gnd 0.007137f
C3564 vdd.n2420 gnd 0.007137f
C3565 vdd.n2421 gnd 0.007137f
C3566 vdd.n2423 gnd 0.007137f
C3567 vdd.n2425 gnd 0.007137f
C3568 vdd.n2426 gnd 0.007137f
C3569 vdd.n2427 gnd 0.007137f
C3570 vdd.n2428 gnd 0.007137f
C3571 vdd.n2429 gnd 0.007137f
C3572 vdd.n2431 gnd 0.007137f
C3573 vdd.n2433 gnd 0.007137f
C3574 vdd.n2434 gnd 0.007137f
C3575 vdd.n2435 gnd 0.007137f
C3576 vdd.n2436 gnd 0.007137f
C3577 vdd.n2437 gnd 0.007137f
C3578 vdd.n2439 gnd 0.007137f
C3579 vdd.n2441 gnd 0.007137f
C3580 vdd.n2442 gnd 0.007137f
C3581 vdd.n2443 gnd 0.007137f
C3582 vdd.n2444 gnd 0.007137f
C3583 vdd.n2445 gnd 0.007137f
C3584 vdd.n2447 gnd 0.007137f
C3585 vdd.n2449 gnd 0.007137f
C3586 vdd.n2450 gnd 0.007137f
C3587 vdd.n2451 gnd 0.007137f
C3588 vdd.n2452 gnd 0.007137f
C3589 vdd.n2453 gnd 0.007137f
C3590 vdd.n2455 gnd 0.007137f
C3591 vdd.n2456 gnd 0.007137f
C3592 vdd.n2457 gnd 0.007137f
C3593 vdd.n2458 gnd 0.007137f
C3594 vdd.n2459 gnd 0.007137f
C3595 vdd.n2460 gnd 0.007137f
C3596 vdd.n2462 gnd 0.007137f
C3597 vdd.n2463 gnd 0.007137f
C3598 vdd.n2464 gnd 0.01645f
C3599 vdd.n2465 gnd 0.015457f
C3600 vdd.n2466 gnd 0.015457f
C3601 vdd.n2467 gnd 1.00827f
C3602 vdd.n2468 gnd 0.015457f
C3603 vdd.n2469 gnd 0.015457f
C3604 vdd.n2470 gnd 0.007137f
C3605 vdd.n2471 gnd 0.007137f
C3606 vdd.n2472 gnd 0.007137f
C3607 vdd.n2473 gnd 0.498774f
C3608 vdd.n2474 gnd 0.007137f
C3609 vdd.n2475 gnd 0.007137f
C3610 vdd.n2476 gnd 0.007137f
C3611 vdd.n2477 gnd 0.007137f
C3612 vdd.n2478 gnd 0.007137f
C3613 vdd.n2479 gnd 0.72939f
C3614 vdd.n2480 gnd 0.007137f
C3615 vdd.n2481 gnd 0.007137f
C3616 vdd.n2482 gnd 0.007137f
C3617 vdd.n2483 gnd 0.007137f
C3618 vdd.n2484 gnd 0.007137f
C3619 vdd.n2485 gnd 0.72939f
C3620 vdd.n2486 gnd 0.007137f
C3621 vdd.n2487 gnd 0.007137f
C3622 vdd.n2488 gnd 0.007137f
C3623 vdd.n2489 gnd 0.007137f
C3624 vdd.n2490 gnd 0.007137f
C3625 vdd.n2491 gnd 0.370058f
C3626 vdd.n2492 gnd 0.007137f
C3627 vdd.n2493 gnd 0.007137f
C3628 vdd.n2494 gnd 0.007137f
C3629 vdd.n2495 gnd 0.007137f
C3630 vdd.n2496 gnd 0.007137f
C3631 vdd.n2497 gnd 0.530953f
C3632 vdd.n2498 gnd 0.007137f
C3633 vdd.n2499 gnd 0.007137f
C3634 vdd.n2500 gnd 0.007137f
C3635 vdd.n2501 gnd 0.007137f
C3636 vdd.n2502 gnd 0.007137f
C3637 vdd.n2503 gnd 0.691848f
C3638 vdd.n2504 gnd 0.007137f
C3639 vdd.n2505 gnd 0.007137f
C3640 vdd.n2506 gnd 0.007137f
C3641 vdd.n2507 gnd 0.007137f
C3642 vdd.n2508 gnd 0.007137f
C3643 vdd.n2509 gnd 0.72939f
C3644 vdd.n2510 gnd 0.007137f
C3645 vdd.n2511 gnd 0.007137f
C3646 vdd.n2512 gnd 0.007137f
C3647 vdd.n2513 gnd 0.007137f
C3648 vdd.n2514 gnd 0.007137f
C3649 vdd.n2515 gnd 0.606037f
C3650 vdd.n2516 gnd 0.007137f
C3651 vdd.n2517 gnd 0.007137f
C3652 vdd.n2518 gnd 0.005878f
C3653 vdd.n2519 gnd 0.020676f
C3654 vdd.n2520 gnd 0.004828f
C3655 vdd.n2521 gnd 0.007137f
C3656 vdd.n2522 gnd 0.445142f
C3657 vdd.n2523 gnd 0.007137f
C3658 vdd.n2524 gnd 0.007137f
C3659 vdd.n2525 gnd 0.007137f
C3660 vdd.n2526 gnd 0.007137f
C3661 vdd.n2527 gnd 0.007137f
C3662 vdd.n2528 gnd 0.445142f
C3663 vdd.n2529 gnd 0.007137f
C3664 vdd.n2530 gnd 0.007137f
C3665 vdd.n2531 gnd 0.007137f
C3666 vdd.n2532 gnd 0.007137f
C3667 vdd.n2533 gnd 0.007137f
C3668 vdd.n2534 gnd 0.606037f
C3669 vdd.n2535 gnd 0.007137f
C3670 vdd.n2536 gnd 0.007137f
C3671 vdd.n2537 gnd 0.007137f
C3672 vdd.n2538 gnd 0.007137f
C3673 vdd.n2539 gnd 0.007137f
C3674 vdd.n2540 gnd 0.622127f
C3675 vdd.n2541 gnd 0.007137f
C3676 vdd.n2542 gnd 0.007137f
C3677 vdd.n2543 gnd 0.007137f
C3678 vdd.n2544 gnd 0.007137f
C3679 vdd.n2545 gnd 0.007137f
C3680 vdd.n2546 gnd 0.461232f
C3681 vdd.n2547 gnd 0.007137f
C3682 vdd.n2548 gnd 0.007137f
C3683 vdd.n2549 gnd 0.007137f
C3684 vdd.n2550 gnd 0.007137f
C3685 vdd.n2551 gnd 0.007137f
C3686 vdd.n2552 gnd 0.230616f
C3687 vdd.n2553 gnd 0.007137f
C3688 vdd.n2554 gnd 0.007137f
C3689 vdd.n2555 gnd 0.007137f
C3690 vdd.n2556 gnd 0.007137f
C3691 vdd.n2557 gnd 0.007137f
C3692 vdd.n2558 gnd 0.230616f
C3693 vdd.n2559 gnd 0.007137f
C3694 vdd.n2560 gnd 0.007137f
C3695 vdd.n2561 gnd 0.007137f
C3696 vdd.n2562 gnd 0.007137f
C3697 vdd.n2563 gnd 0.007137f
C3698 vdd.n2564 gnd 0.72939f
C3699 vdd.n2565 gnd 0.007137f
C3700 vdd.n2566 gnd 0.007137f
C3701 vdd.n2567 gnd 0.007137f
C3702 vdd.n2568 gnd 0.007137f
C3703 vdd.n2569 gnd 0.007137f
C3704 vdd.n2570 gnd 0.007137f
C3705 vdd.n2571 gnd 0.007137f
C3706 vdd.n2572 gnd 0.52559f
C3707 vdd.n2573 gnd 0.007137f
C3708 vdd.n2574 gnd 0.007137f
C3709 vdd.n2575 gnd 0.007137f
C3710 vdd.n2576 gnd 0.007137f
C3711 vdd.n2577 gnd 0.007137f
C3712 vdd.n2578 gnd 0.007137f
C3713 vdd.n2579 gnd 0.455869f
C3714 vdd.n2580 gnd 0.007137f
C3715 vdd.n2581 gnd 0.007137f
C3716 vdd.n2582 gnd 0.007137f
C3717 vdd.n2583 gnd 0.016362f
C3718 vdd.n2584 gnd 0.015545f
C3719 vdd.n2585 gnd 0.007137f
C3720 vdd.n2586 gnd 0.007137f
C3721 vdd.n2587 gnd 0.00551f
C3722 vdd.n2588 gnd 0.007137f
C3723 vdd.n2589 gnd 0.007137f
C3724 vdd.n2590 gnd 0.005195f
C3725 vdd.n2591 gnd 0.007137f
C3726 vdd.n2592 gnd 0.007137f
C3727 vdd.n2593 gnd 0.007137f
C3728 vdd.n2594 gnd 0.007137f
C3729 vdd.n2595 gnd 0.007137f
C3730 vdd.n2596 gnd 0.007137f
C3731 vdd.n2597 gnd 0.007137f
C3732 vdd.n2598 gnd 0.007137f
C3733 vdd.n2599 gnd 0.007137f
C3734 vdd.n2600 gnd 0.007137f
C3735 vdd.n2601 gnd 0.007137f
C3736 vdd.n2602 gnd 0.007137f
C3737 vdd.n2603 gnd 0.007137f
C3738 vdd.n2604 gnd 0.007137f
C3739 vdd.n2605 gnd 0.007137f
C3740 vdd.n2606 gnd 0.007137f
C3741 vdd.n2607 gnd 0.007137f
C3742 vdd.n2608 gnd 0.007137f
C3743 vdd.n2609 gnd 0.007137f
C3744 vdd.n2610 gnd 0.007137f
C3745 vdd.n2611 gnd 0.007137f
C3746 vdd.n2612 gnd 0.007137f
C3747 vdd.n2613 gnd 0.007137f
C3748 vdd.n2614 gnd 0.007137f
C3749 vdd.n2615 gnd 0.007137f
C3750 vdd.n2616 gnd 0.007137f
C3751 vdd.n2617 gnd 0.007137f
C3752 vdd.n2618 gnd 0.007137f
C3753 vdd.n2619 gnd 0.007137f
C3754 vdd.n2620 gnd 0.007137f
C3755 vdd.n2621 gnd 0.007137f
C3756 vdd.n2622 gnd 0.007137f
C3757 vdd.n2623 gnd 0.007137f
C3758 vdd.n2624 gnd 0.007137f
C3759 vdd.n2625 gnd 0.007137f
C3760 vdd.n2626 gnd 0.007137f
C3761 vdd.n2627 gnd 0.007137f
C3762 vdd.n2628 gnd 0.007137f
C3763 vdd.n2629 gnd 0.007137f
C3764 vdd.n2630 gnd 0.007137f
C3765 vdd.n2631 gnd 0.007137f
C3766 vdd.n2632 gnd 0.007137f
C3767 vdd.n2633 gnd 0.007137f
C3768 vdd.n2634 gnd 0.007137f
C3769 vdd.n2635 gnd 0.007137f
C3770 vdd.n2636 gnd 0.007137f
C3771 vdd.n2637 gnd 0.007137f
C3772 vdd.n2638 gnd 0.007137f
C3773 vdd.n2639 gnd 0.007137f
C3774 vdd.n2640 gnd 0.007137f
C3775 vdd.n2641 gnd 0.007137f
C3776 vdd.n2642 gnd 0.007137f
C3777 vdd.n2643 gnd 0.007137f
C3778 vdd.n2644 gnd 0.007137f
C3779 vdd.n2645 gnd 0.007137f
C3780 vdd.n2646 gnd 0.007137f
C3781 vdd.n2647 gnd 0.007137f
C3782 vdd.n2648 gnd 0.007137f
C3783 vdd.n2649 gnd 0.007137f
C3784 vdd.n2650 gnd 0.007137f
C3785 vdd.n2651 gnd 0.01645f
C3786 vdd.n2652 gnd 0.015457f
C3787 vdd.n2653 gnd 0.015457f
C3788 vdd.n2654 gnd 0.847379f
C3789 vdd.n2655 gnd 0.015457f
C3790 vdd.n2656 gnd 0.01645f
C3791 vdd.n2657 gnd 0.015545f
C3792 vdd.n2658 gnd 0.007137f
C3793 vdd.n2659 gnd 0.007137f
C3794 vdd.n2660 gnd 0.007137f
C3795 vdd.n2661 gnd 0.00551f
C3796 vdd.n2662 gnd 0.0102f
C3797 vdd.n2663 gnd 0.005195f
C3798 vdd.n2664 gnd 0.007137f
C3799 vdd.n2665 gnd 0.007137f
C3800 vdd.n2666 gnd 0.007137f
C3801 vdd.n2667 gnd 0.007137f
C3802 vdd.n2668 gnd 0.007137f
C3803 vdd.n2669 gnd 0.007137f
C3804 vdd.n2670 gnd 0.007137f
C3805 vdd.n2671 gnd 0.007137f
C3806 vdd.n2672 gnd 0.007137f
C3807 vdd.n2673 gnd 0.007137f
C3808 vdd.n2674 gnd 0.007137f
C3809 vdd.n2675 gnd 0.007137f
C3810 vdd.n2676 gnd 0.007137f
C3811 vdd.n2677 gnd 0.007137f
C3812 vdd.n2678 gnd 0.007137f
C3813 vdd.n2679 gnd 0.007137f
C3814 vdd.n2680 gnd 0.007137f
C3815 vdd.n2681 gnd 0.007137f
C3816 vdd.n2682 gnd 0.007137f
C3817 vdd.n2683 gnd 0.007137f
C3818 vdd.n2684 gnd 0.007137f
C3819 vdd.n2685 gnd 0.007137f
C3820 vdd.n2686 gnd 0.007137f
C3821 vdd.n2687 gnd 0.007137f
C3822 vdd.n2688 gnd 0.007137f
C3823 vdd.n2689 gnd 0.007137f
C3824 vdd.n2690 gnd 0.007137f
C3825 vdd.n2691 gnd 0.007137f
C3826 vdd.n2692 gnd 0.007137f
C3827 vdd.n2693 gnd 0.007137f
C3828 vdd.n2694 gnd 0.007137f
C3829 vdd.n2695 gnd 0.007137f
C3830 vdd.n2696 gnd 0.007137f
C3831 vdd.n2697 gnd 0.007137f
C3832 vdd.n2698 gnd 0.007137f
C3833 vdd.n2699 gnd 0.007137f
C3834 vdd.n2700 gnd 0.007137f
C3835 vdd.n2701 gnd 0.007137f
C3836 vdd.n2702 gnd 0.007137f
C3837 vdd.n2703 gnd 0.007137f
C3838 vdd.n2704 gnd 0.007137f
C3839 vdd.n2705 gnd 0.007137f
C3840 vdd.n2706 gnd 0.007137f
C3841 vdd.n2707 gnd 0.007137f
C3842 vdd.n2708 gnd 0.007137f
C3843 vdd.n2709 gnd 0.007137f
C3844 vdd.n2710 gnd 0.007137f
C3845 vdd.n2711 gnd 0.007137f
C3846 vdd.n2712 gnd 0.007137f
C3847 vdd.n2713 gnd 0.007137f
C3848 vdd.n2714 gnd 0.007137f
C3849 vdd.n2715 gnd 0.007137f
C3850 vdd.n2716 gnd 0.007137f
C3851 vdd.n2717 gnd 0.007137f
C3852 vdd.n2718 gnd 0.007137f
C3853 vdd.n2719 gnd 0.007137f
C3854 vdd.n2720 gnd 0.007137f
C3855 vdd.n2721 gnd 0.007137f
C3856 vdd.n2722 gnd 0.007137f
C3857 vdd.n2723 gnd 0.007137f
C3858 vdd.n2724 gnd 0.01645f
C3859 vdd.n2725 gnd 0.01645f
C3860 vdd.n2726 gnd 0.890285f
C3861 vdd.t43 gnd 3.16426f
C3862 vdd.t298 gnd 3.16426f
C3863 vdd.n2760 gnd 0.007137f
C3864 vdd.t122 gnd 0.288414f
C3865 vdd.t123 gnd 0.295228f
C3866 vdd.t121 gnd 0.188288f
C3867 vdd.n2761 gnd 0.101759f
C3868 vdd.n2762 gnd 0.057721f
C3869 vdd.n2763 gnd 0.0102f
C3870 vdd.n2764 gnd 0.007137f
C3871 vdd.n2765 gnd 0.007137f
C3872 vdd.n2766 gnd 0.007137f
C3873 vdd.n2767 gnd 0.007137f
C3874 vdd.n2768 gnd 0.007137f
C3875 vdd.n2769 gnd 0.007137f
C3876 vdd.n2770 gnd 0.007137f
C3877 vdd.n2771 gnd 0.007137f
C3878 vdd.n2772 gnd 0.007137f
C3879 vdd.n2773 gnd 0.007137f
C3880 vdd.n2774 gnd 0.007137f
C3881 vdd.n2775 gnd 0.007137f
C3882 vdd.n2776 gnd 0.007137f
C3883 vdd.n2777 gnd 0.007137f
C3884 vdd.n2778 gnd 0.007137f
C3885 vdd.n2779 gnd 0.007137f
C3886 vdd.n2780 gnd 0.007137f
C3887 vdd.n2781 gnd 0.007137f
C3888 vdd.n2782 gnd 0.007137f
C3889 vdd.n2783 gnd 0.007137f
C3890 vdd.n2784 gnd 0.007137f
C3891 vdd.n2785 gnd 0.007137f
C3892 vdd.n2786 gnd 0.007137f
C3893 vdd.n2787 gnd 0.007137f
C3894 vdd.n2788 gnd 0.007137f
C3895 vdd.n2789 gnd 0.007137f
C3896 vdd.n2790 gnd 0.007137f
C3897 vdd.n2791 gnd 0.007137f
C3898 vdd.n2792 gnd 0.007137f
C3899 vdd.n2793 gnd 0.007137f
C3900 vdd.n2794 gnd 0.007137f
C3901 vdd.n2795 gnd 0.007137f
C3902 vdd.n2796 gnd 0.007137f
C3903 vdd.n2797 gnd 0.007137f
C3904 vdd.n2798 gnd 0.007137f
C3905 vdd.n2799 gnd 0.007137f
C3906 vdd.n2800 gnd 0.007137f
C3907 vdd.n2801 gnd 0.007137f
C3908 vdd.n2802 gnd 0.007137f
C3909 vdd.n2803 gnd 0.007137f
C3910 vdd.n2804 gnd 0.007137f
C3911 vdd.n2805 gnd 0.007137f
C3912 vdd.n2806 gnd 0.007137f
C3913 vdd.n2807 gnd 0.007137f
C3914 vdd.n2808 gnd 0.007137f
C3915 vdd.n2809 gnd 0.007137f
C3916 vdd.n2810 gnd 0.007137f
C3917 vdd.n2811 gnd 0.007137f
C3918 vdd.n2812 gnd 0.007137f
C3919 vdd.n2813 gnd 0.007137f
C3920 vdd.n2814 gnd 0.007137f
C3921 vdd.n2815 gnd 0.007137f
C3922 vdd.n2816 gnd 0.007137f
C3923 vdd.n2817 gnd 0.007137f
C3924 vdd.n2818 gnd 0.007137f
C3925 vdd.n2819 gnd 0.007137f
C3926 vdd.n2820 gnd 0.007137f
C3927 vdd.n2821 gnd 0.007137f
C3928 vdd.n2822 gnd 0.007137f
C3929 vdd.n2823 gnd 0.007137f
C3930 vdd.n2824 gnd 0.005195f
C3931 vdd.n2825 gnd 0.007137f
C3932 vdd.n2826 gnd 0.007137f
C3933 vdd.n2827 gnd 0.00551f
C3934 vdd.n2828 gnd 0.007137f
C3935 vdd.n2829 gnd 0.007137f
C3936 vdd.t109 gnd 0.288414f
C3937 vdd.t110 gnd 0.295228f
C3938 vdd.t107 gnd 0.188288f
C3939 vdd.n2830 gnd 0.101759f
C3940 vdd.n2831 gnd 0.057721f
C3941 vdd.n2832 gnd 0.007137f
C3942 vdd.n2833 gnd 0.007137f
C3943 vdd.n2834 gnd 0.007137f
C3944 vdd.n2835 gnd 0.007137f
C3945 vdd.n2836 gnd 0.007137f
C3946 vdd.n2837 gnd 0.007137f
C3947 vdd.n2838 gnd 0.007137f
C3948 vdd.n2839 gnd 0.007137f
C3949 vdd.n2840 gnd 0.007137f
C3950 vdd.n2841 gnd 0.007137f
C3951 vdd.n2842 gnd 0.007137f
C3952 vdd.n2843 gnd 0.007137f
C3953 vdd.n2844 gnd 0.007137f
C3954 vdd.n2845 gnd 0.007137f
C3955 vdd.n2846 gnd 0.007137f
C3956 vdd.n2847 gnd 0.007137f
C3957 vdd.n2848 gnd 0.007137f
C3958 vdd.n2849 gnd 0.007137f
C3959 vdd.n2850 gnd 0.007137f
C3960 vdd.n2851 gnd 0.007137f
C3961 vdd.n2852 gnd 0.007137f
C3962 vdd.n2853 gnd 0.007137f
C3963 vdd.n2854 gnd 0.007137f
C3964 vdd.n2855 gnd 0.007137f
C3965 vdd.n2856 gnd 0.007137f
C3966 vdd.n2857 gnd 0.007137f
C3967 vdd.n2858 gnd 0.007137f
C3968 vdd.n2859 gnd 0.007137f
C3969 vdd.n2860 gnd 0.007137f
C3970 vdd.n2861 gnd 0.007137f
C3971 vdd.n2862 gnd 0.007137f
C3972 vdd.n2863 gnd 0.007137f
C3973 vdd.n2864 gnd 0.007137f
C3974 vdd.n2865 gnd 0.007137f
C3975 vdd.n2866 gnd 0.007137f
C3976 vdd.n2867 gnd 0.007137f
C3977 vdd.n2868 gnd 0.007137f
C3978 vdd.n2869 gnd 0.007137f
C3979 vdd.n2870 gnd 0.007137f
C3980 vdd.n2871 gnd 0.007137f
C3981 vdd.n2872 gnd 0.007137f
C3982 vdd.n2873 gnd 0.007137f
C3983 vdd.n2874 gnd 0.007137f
C3984 vdd.n2875 gnd 0.007137f
C3985 vdd.n2876 gnd 0.007137f
C3986 vdd.n2877 gnd 0.007137f
C3987 vdd.n2878 gnd 0.007137f
C3988 vdd.n2879 gnd 0.007137f
C3989 vdd.n2880 gnd 0.007137f
C3990 vdd.n2881 gnd 0.007137f
C3991 vdd.n2882 gnd 0.007137f
C3992 vdd.n2883 gnd 0.007137f
C3993 vdd.n2884 gnd 0.007137f
C3994 vdd.n2885 gnd 0.007137f
C3995 vdd.n2886 gnd 0.007137f
C3996 vdd.n2887 gnd 0.007137f
C3997 vdd.n2888 gnd 0.007137f
C3998 vdd.n2889 gnd 0.005195f
C3999 vdd.n2890 gnd 0.0102f
C4000 vdd.n2891 gnd 0.00551f
C4001 vdd.n2892 gnd 0.007137f
C4002 vdd.n2893 gnd 0.007137f
C4003 vdd.n2894 gnd 0.007137f
C4004 vdd.n2895 gnd 0.01645f
C4005 vdd.n2896 gnd 0.01645f
C4006 vdd.n2897 gnd 0.015457f
C4007 vdd.n2898 gnd 0.007137f
C4008 vdd.n2899 gnd 0.007137f
C4009 vdd.n2900 gnd 0.007137f
C4010 vdd.n2901 gnd 0.007137f
C4011 vdd.n2902 gnd 0.007137f
C4012 vdd.n2903 gnd 0.007137f
C4013 vdd.n2904 gnd 0.007137f
C4014 vdd.n2905 gnd 0.007137f
C4015 vdd.n2906 gnd 0.007137f
C4016 vdd.n2907 gnd 0.007137f
C4017 vdd.n2908 gnd 0.007137f
C4018 vdd.n2909 gnd 0.007137f
C4019 vdd.n2910 gnd 0.007137f
C4020 vdd.n2911 gnd 0.007137f
C4021 vdd.n2912 gnd 0.007137f
C4022 vdd.n2913 gnd 0.007137f
C4023 vdd.n2914 gnd 0.007137f
C4024 vdd.n2915 gnd 0.007137f
C4025 vdd.n2916 gnd 0.007137f
C4026 vdd.n2917 gnd 0.007137f
C4027 vdd.n2918 gnd 0.007137f
C4028 vdd.n2919 gnd 0.007137f
C4029 vdd.n2920 gnd 0.007137f
C4030 vdd.n2921 gnd 0.007137f
C4031 vdd.n2922 gnd 0.007137f
C4032 vdd.n2923 gnd 0.007137f
C4033 vdd.n2924 gnd 0.007137f
C4034 vdd.n2925 gnd 0.007137f
C4035 vdd.n2926 gnd 0.007137f
C4036 vdd.n2927 gnd 0.007137f
C4037 vdd.n2928 gnd 0.007137f
C4038 vdd.n2929 gnd 0.007137f
C4039 vdd.n2930 gnd 0.007137f
C4040 vdd.n2931 gnd 0.007137f
C4041 vdd.n2932 gnd 0.007137f
C4042 vdd.n2933 gnd 0.007137f
C4043 vdd.n2934 gnd 0.007137f
C4044 vdd.n2935 gnd 0.007137f
C4045 vdd.n2936 gnd 0.007137f
C4046 vdd.n2937 gnd 0.007137f
C4047 vdd.n2938 gnd 0.007137f
C4048 vdd.n2939 gnd 0.007137f
C4049 vdd.n2940 gnd 0.007137f
C4050 vdd.n2941 gnd 0.007137f
C4051 vdd.n2942 gnd 0.007137f
C4052 vdd.n2943 gnd 0.007137f
C4053 vdd.n2944 gnd 0.007137f
C4054 vdd.n2945 gnd 0.007137f
C4055 vdd.n2946 gnd 0.007137f
C4056 vdd.n2947 gnd 0.007137f
C4057 vdd.n2948 gnd 0.007137f
C4058 vdd.n2949 gnd 0.007137f
C4059 vdd.n2950 gnd 0.007137f
C4060 vdd.n2951 gnd 0.007137f
C4061 vdd.n2952 gnd 0.007137f
C4062 vdd.n2953 gnd 0.007137f
C4063 vdd.n2954 gnd 0.007137f
C4064 vdd.n2955 gnd 0.007137f
C4065 vdd.n2956 gnd 0.007137f
C4066 vdd.n2957 gnd 0.007137f
C4067 vdd.n2958 gnd 0.007137f
C4068 vdd.n2959 gnd 0.007137f
C4069 vdd.n2960 gnd 0.007137f
C4070 vdd.n2961 gnd 0.007137f
C4071 vdd.n2962 gnd 0.007137f
C4072 vdd.n2963 gnd 0.007137f
C4073 vdd.n2964 gnd 0.007137f
C4074 vdd.n2965 gnd 0.007137f
C4075 vdd.n2966 gnd 0.007137f
C4076 vdd.n2967 gnd 0.007137f
C4077 vdd.n2968 gnd 0.007137f
C4078 vdd.n2969 gnd 0.007137f
C4079 vdd.n2970 gnd 0.007137f
C4080 vdd.n2971 gnd 0.007137f
C4081 vdd.n2972 gnd 0.007137f
C4082 vdd.n2973 gnd 0.007137f
C4083 vdd.n2974 gnd 0.007137f
C4084 vdd.n2975 gnd 0.007137f
C4085 vdd.n2976 gnd 0.007137f
C4086 vdd.n2977 gnd 0.230616f
C4087 vdd.n2978 gnd 0.007137f
C4088 vdd.n2979 gnd 0.007137f
C4089 vdd.n2980 gnd 0.007137f
C4090 vdd.n2981 gnd 0.007137f
C4091 vdd.n2982 gnd 0.007137f
C4092 vdd.n2983 gnd 0.007137f
C4093 vdd.n2984 gnd 0.007137f
C4094 vdd.n2985 gnd 0.007137f
C4095 vdd.n2986 gnd 0.007137f
C4096 vdd.n2987 gnd 0.007137f
C4097 vdd.n2988 gnd 0.007137f
C4098 vdd.n2989 gnd 0.659669f
C4099 vdd.n2990 gnd 0.007137f
C4100 vdd.n2991 gnd 0.007137f
C4101 vdd.n2992 gnd 0.007137f
C4102 vdd.n2993 gnd 0.007137f
C4103 vdd.n2994 gnd 0.007137f
C4104 vdd.n2995 gnd 0.007137f
C4105 vdd.n2996 gnd 0.007137f
C4106 vdd.n2997 gnd 0.007137f
C4107 vdd.n2998 gnd 0.007137f
C4108 vdd.n2999 gnd 0.007137f
C4109 vdd.n3000 gnd 0.007137f
C4110 vdd.n3001 gnd 0.434416f
C4111 vdd.n3002 gnd 0.007137f
C4112 vdd.n3003 gnd 0.007137f
C4113 vdd.n3004 gnd 0.007137f
C4114 vdd.n3005 gnd 0.007137f
C4115 vdd.n3006 gnd 0.007137f
C4116 vdd.n3007 gnd 0.015457f
C4117 vdd.n3008 gnd 0.01645f
C4118 vdd.n3009 gnd 0.01645f
C4119 vdd.n3010 gnd 0.890285f
C4120 vdd.n3012 gnd 0.007137f
C4121 vdd.n3013 gnd 0.007137f
C4122 vdd.n3014 gnd 0.01645f
C4123 vdd.n3015 gnd 0.015457f
C4124 vdd.n3016 gnd 0.015457f
C4125 vdd.n3017 gnd 0.847379f
C4126 vdd.n3018 gnd 0.015457f
C4127 vdd.n3019 gnd 0.015457f
C4128 vdd.n3020 gnd 0.007137f
C4129 vdd.n3021 gnd 0.007137f
C4130 vdd.n3022 gnd 0.007137f
C4131 vdd.n3023 gnd 0.455869f
C4132 vdd.n3024 gnd 0.007137f
C4133 vdd.n3025 gnd 0.007137f
C4134 vdd.n3026 gnd 0.007137f
C4135 vdd.n3027 gnd 0.007137f
C4136 vdd.n3028 gnd 0.007137f
C4137 vdd.n3029 gnd 0.52559f
C4138 vdd.n3030 gnd 0.007137f
C4139 vdd.n3031 gnd 0.007137f
C4140 vdd.n3032 gnd 0.007137f
C4141 vdd.n3033 gnd 0.007137f
C4142 vdd.n3034 gnd 0.007137f
C4143 vdd.n3035 gnd 0.72939f
C4144 vdd.n3036 gnd 0.007137f
C4145 vdd.n3037 gnd 0.007137f
C4146 vdd.n3038 gnd 0.007137f
C4147 vdd.n3039 gnd 0.007137f
C4148 vdd.n3040 gnd 0.007137f
C4149 vdd.n3041 gnd 0.230616f
C4150 vdd.n3042 gnd 0.007137f
C4151 vdd.n3043 gnd 0.007137f
C4152 vdd.n3044 gnd 0.007137f
C4153 vdd.n3045 gnd 0.007137f
C4154 vdd.n3046 gnd 0.007137f
C4155 vdd.n3047 gnd 0.230616f
C4156 vdd.n3048 gnd 0.007137f
C4157 vdd.n3049 gnd 0.007137f
C4158 vdd.n3050 gnd 0.007137f
C4159 vdd.n3051 gnd 0.007137f
C4160 vdd.n3052 gnd 0.007137f
C4161 vdd.n3053 gnd 0.461232f
C4162 vdd.n3054 gnd 0.007137f
C4163 vdd.n3055 gnd 0.007137f
C4164 vdd.n3056 gnd 0.007137f
C4165 vdd.n3057 gnd 0.007137f
C4166 vdd.n3058 gnd 0.007137f
C4167 vdd.n3059 gnd 0.622127f
C4168 vdd.n3060 gnd 0.007137f
C4169 vdd.n3061 gnd 0.007137f
C4170 vdd.n3062 gnd 0.007137f
C4171 vdd.n3063 gnd 0.007137f
C4172 vdd.n3064 gnd 0.007137f
C4173 vdd.n3065 gnd 0.606037f
C4174 vdd.n3066 gnd 0.007137f
C4175 vdd.n3067 gnd 0.007137f
C4176 vdd.n3068 gnd 0.007137f
C4177 vdd.n3069 gnd 0.007137f
C4178 vdd.n3070 gnd 0.007137f
C4179 vdd.n3071 gnd 0.445142f
C4180 vdd.n3072 gnd 0.007137f
C4181 vdd.n3073 gnd 0.007137f
C4182 vdd.n3074 gnd 0.007137f
C4183 vdd.n3075 gnd 0.007137f
C4184 vdd.n3076 gnd 0.007137f
C4185 vdd.n3077 gnd 0.445142f
C4186 vdd.n3078 gnd 0.007137f
C4187 vdd.n3079 gnd 0.004828f
C4188 vdd.n3080 gnd 0.020676f
C4189 vdd.n3081 gnd 0.005878f
C4190 vdd.n3082 gnd 0.007137f
C4191 vdd.n3083 gnd 0.007137f
C4192 vdd.n3084 gnd 0.606037f
C4193 vdd.n3085 gnd 0.007137f
C4194 vdd.n3086 gnd 0.007137f
C4195 vdd.n3087 gnd 0.007137f
C4196 vdd.n3088 gnd 0.007137f
C4197 vdd.n3089 gnd 0.007137f
C4198 vdd.n3090 gnd 0.72939f
C4199 vdd.n3091 gnd 0.007137f
C4200 vdd.n3092 gnd 0.007137f
C4201 vdd.n3093 gnd 0.007137f
C4202 vdd.n3094 gnd 0.007137f
C4203 vdd.n3095 gnd 0.007137f
C4204 vdd.n3096 gnd 0.691848f
C4205 vdd.n3097 gnd 0.007137f
C4206 vdd.n3098 gnd 0.007137f
C4207 vdd.n3099 gnd 0.007137f
C4208 vdd.n3100 gnd 0.007137f
C4209 vdd.n3101 gnd 0.007137f
C4210 vdd.n3102 gnd 0.530953f
C4211 vdd.n3103 gnd 0.007137f
C4212 vdd.n3104 gnd 0.007137f
C4213 vdd.n3105 gnd 0.007137f
C4214 vdd.n3106 gnd 0.007137f
C4215 vdd.n3107 gnd 0.007137f
C4216 vdd.n3108 gnd 0.370058f
C4217 vdd.n3109 gnd 0.007137f
C4218 vdd.n3110 gnd 0.007137f
C4219 vdd.n3111 gnd 0.007137f
C4220 vdd.n3112 gnd 0.007137f
C4221 vdd.n3113 gnd 0.007137f
C4222 vdd.n3114 gnd 0.72939f
C4223 vdd.n3115 gnd 0.007137f
C4224 vdd.n3116 gnd 0.007137f
C4225 vdd.n3117 gnd 0.007137f
C4226 vdd.n3118 gnd 0.007137f
C4227 vdd.n3119 gnd 0.007137f
C4228 vdd.n3120 gnd 0.007137f
C4229 vdd.n3122 gnd 0.007137f
C4230 vdd.n3123 gnd 0.007137f
C4231 vdd.n3125 gnd 0.007137f
C4232 vdd.n3126 gnd 0.007137f
C4233 vdd.n3129 gnd 0.007137f
C4234 vdd.n3130 gnd 0.007137f
C4235 vdd.n3131 gnd 0.007137f
C4236 vdd.n3132 gnd 0.007137f
C4237 vdd.n3134 gnd 0.007137f
C4238 vdd.n3135 gnd 0.007137f
C4239 vdd.n3136 gnd 0.007137f
C4240 vdd.n3137 gnd 0.007137f
C4241 vdd.n3138 gnd 0.007137f
C4242 vdd.n3139 gnd 0.007137f
C4243 vdd.n3141 gnd 0.007137f
C4244 vdd.n3142 gnd 0.007137f
C4245 vdd.n3143 gnd 0.007137f
C4246 vdd.n3144 gnd 0.007137f
C4247 vdd.n3145 gnd 0.007137f
C4248 vdd.n3146 gnd 0.007137f
C4249 vdd.n3148 gnd 0.007137f
C4250 vdd.n3149 gnd 0.007137f
C4251 vdd.n3150 gnd 0.007137f
C4252 vdd.n3151 gnd 0.007137f
C4253 vdd.n3152 gnd 0.007137f
C4254 vdd.n3153 gnd 0.007137f
C4255 vdd.n3155 gnd 0.007137f
C4256 vdd.n3156 gnd 0.01645f
C4257 vdd.n3157 gnd 0.01645f
C4258 vdd.n3158 gnd 0.015457f
C4259 vdd.n3159 gnd 0.007137f
C4260 vdd.n3160 gnd 0.007137f
C4261 vdd.n3161 gnd 0.007137f
C4262 vdd.n3162 gnd 0.007137f
C4263 vdd.n3163 gnd 0.007137f
C4264 vdd.n3164 gnd 0.007137f
C4265 vdd.n3165 gnd 0.72939f
C4266 vdd.n3166 gnd 0.007137f
C4267 vdd.n3167 gnd 0.007137f
C4268 vdd.n3168 gnd 0.007137f
C4269 vdd.n3169 gnd 0.007137f
C4270 vdd.n3170 gnd 0.007137f
C4271 vdd.n3171 gnd 0.498774f
C4272 vdd.n3172 gnd 0.007137f
C4273 vdd.n3173 gnd 0.007137f
C4274 vdd.n3174 gnd 0.007137f
C4275 vdd.n3175 gnd 0.016362f
C4276 vdd.n3176 gnd 0.015545f
C4277 vdd.n3177 gnd 0.01645f
C4278 vdd.n3179 gnd 0.007137f
C4279 vdd.n3180 gnd 0.007137f
C4280 vdd.n3181 gnd 0.00551f
C4281 vdd.n3182 gnd 0.0102f
C4282 vdd.n3183 gnd 0.005195f
C4283 vdd.n3184 gnd 0.007137f
C4284 vdd.n3185 gnd 0.007137f
C4285 vdd.n3187 gnd 0.007137f
C4286 vdd.n3188 gnd 0.007137f
C4287 vdd.n3189 gnd 0.007137f
C4288 vdd.n3190 gnd 0.007137f
C4289 vdd.n3191 gnd 0.007137f
C4290 vdd.n3192 gnd 0.007137f
C4291 vdd.n3194 gnd 0.007137f
C4292 vdd.n3195 gnd 0.007137f
C4293 vdd.n3196 gnd 0.007137f
C4294 vdd.n3197 gnd 0.007137f
C4295 vdd.n3198 gnd 0.007137f
C4296 vdd.n3199 gnd 0.007137f
C4297 vdd.n3201 gnd 0.007137f
C4298 vdd.n3202 gnd 0.007137f
C4299 vdd.n3203 gnd 0.007137f
C4300 vdd.n3204 gnd 0.007137f
C4301 vdd.n3205 gnd 0.007137f
C4302 vdd.n3206 gnd 0.007137f
C4303 vdd.n3208 gnd 0.007137f
C4304 vdd.n3209 gnd 0.007137f
C4305 vdd.n3210 gnd 0.007137f
C4306 vdd.n3212 gnd 0.007137f
C4307 vdd.n3213 gnd 0.007137f
C4308 vdd.n3214 gnd 0.007137f
C4309 vdd.n3215 gnd 0.007137f
C4310 vdd.n3216 gnd 0.007137f
C4311 vdd.n3217 gnd 0.007137f
C4312 vdd.n3219 gnd 0.007137f
C4313 vdd.n3220 gnd 0.007137f
C4314 vdd.n3221 gnd 0.007137f
C4315 vdd.n3222 gnd 0.007137f
C4316 vdd.n3223 gnd 0.007137f
C4317 vdd.n3224 gnd 0.007137f
C4318 vdd.n3226 gnd 0.007137f
C4319 vdd.n3227 gnd 0.007137f
C4320 vdd.n3228 gnd 0.007137f
C4321 vdd.n3229 gnd 0.007137f
C4322 vdd.n3230 gnd 0.007137f
C4323 vdd.n3231 gnd 0.007137f
C4324 vdd.n3233 gnd 0.007137f
C4325 vdd.n3234 gnd 0.007137f
C4326 vdd.n3236 gnd 0.007137f
C4327 vdd.n3237 gnd 0.007137f
C4328 vdd.n3238 gnd 0.01645f
C4329 vdd.n3239 gnd 0.015457f
C4330 vdd.n3240 gnd 0.015457f
C4331 vdd.n3241 gnd 1.00827f
C4332 vdd.n3242 gnd 0.015457f
C4333 vdd.n3243 gnd 0.01645f
C4334 vdd.n3244 gnd 0.015545f
C4335 vdd.n3245 gnd 0.007137f
C4336 vdd.n3246 gnd 0.00551f
C4337 vdd.n3247 gnd 0.007137f
C4338 vdd.n3249 gnd 0.007137f
C4339 vdd.n3250 gnd 0.007137f
C4340 vdd.n3251 gnd 0.007137f
C4341 vdd.n3252 gnd 0.007137f
C4342 vdd.n3253 gnd 0.007137f
C4343 vdd.n3254 gnd 0.007137f
C4344 vdd.n3256 gnd 0.007137f
C4345 vdd.n3257 gnd 0.007137f
C4346 vdd.n3258 gnd 0.007137f
C4347 vdd.n3259 gnd 0.007137f
C4348 vdd.n3260 gnd 0.007137f
C4349 vdd.n3261 gnd 0.007137f
C4350 vdd.n3263 gnd 0.007137f
C4351 vdd.n3264 gnd 0.007137f
C4352 vdd.n3265 gnd 0.007137f
C4353 vdd.n3266 gnd 0.007137f
C4354 vdd.n3267 gnd 0.007137f
C4355 vdd.n3268 gnd 0.007137f
C4356 vdd.n3270 gnd 0.007137f
C4357 vdd.n3271 gnd 0.007137f
C4358 vdd.n3273 gnd 0.007137f
C4359 vdd.n3274 gnd 0.033502f
C4360 vdd.n3275 gnd 0.958844f
C4361 vdd.n3277 gnd 0.004435f
C4362 vdd.n3278 gnd 0.008448f
C4363 vdd.n3279 gnd 0.010496f
C4364 vdd.n3280 gnd 0.010496f
C4365 vdd.n3281 gnd 0.008448f
C4366 vdd.n3282 gnd 0.008448f
C4367 vdd.n3283 gnd 0.010496f
C4368 vdd.n3284 gnd 0.010496f
C4369 vdd.n3285 gnd 0.008448f
C4370 vdd.n3286 gnd 0.008448f
C4371 vdd.n3287 gnd 0.010496f
C4372 vdd.n3288 gnd 0.010496f
C4373 vdd.n3289 gnd 0.008448f
C4374 vdd.n3290 gnd 0.008448f
C4375 vdd.n3291 gnd 0.010496f
C4376 vdd.n3292 gnd 0.010496f
C4377 vdd.n3293 gnd 0.008448f
C4378 vdd.n3294 gnd 0.008448f
C4379 vdd.n3295 gnd 0.010496f
C4380 vdd.n3296 gnd 0.010496f
C4381 vdd.n3297 gnd 0.008448f
C4382 vdd.n3298 gnd 0.008448f
C4383 vdd.n3299 gnd 0.010496f
C4384 vdd.n3300 gnd 0.010496f
C4385 vdd.n3301 gnd 0.008448f
C4386 vdd.n3302 gnd 0.008448f
C4387 vdd.n3303 gnd 0.010496f
C4388 vdd.n3304 gnd 0.010496f
C4389 vdd.n3305 gnd 0.008448f
C4390 vdd.n3306 gnd 0.008448f
C4391 vdd.n3307 gnd 0.010496f
C4392 vdd.n3308 gnd 0.010496f
C4393 vdd.n3309 gnd 0.008448f
C4394 vdd.n3310 gnd 0.008448f
C4395 vdd.n3311 gnd 0.010496f
C4396 vdd.n3312 gnd 0.010496f
C4397 vdd.n3313 gnd 0.008448f
C4398 vdd.n3314 gnd 0.010496f
C4399 vdd.n3315 gnd 0.010496f
C4400 vdd.n3316 gnd 0.008448f
C4401 vdd.n3317 gnd 0.010496f
C4402 vdd.n3318 gnd 0.010496f
C4403 vdd.n3319 gnd 0.010496f
C4404 vdd.n3320 gnd 0.017234f
C4405 vdd.n3321 gnd 0.010496f
C4406 vdd.n3322 gnd 0.010496f
C4407 vdd.n3323 gnd 0.005745f
C4408 vdd.n3324 gnd 0.008448f
C4409 vdd.n3325 gnd 0.010496f
C4410 vdd.n3326 gnd 0.010496f
C4411 vdd.n3327 gnd 0.008448f
C4412 vdd.n3328 gnd 0.008448f
C4413 vdd.n3329 gnd 0.010496f
C4414 vdd.n3330 gnd 0.010496f
C4415 vdd.n3331 gnd 0.008448f
C4416 vdd.n3332 gnd 0.008448f
C4417 vdd.n3333 gnd 0.010496f
C4418 vdd.n3334 gnd 0.010496f
C4419 vdd.n3335 gnd 0.008448f
C4420 vdd.n3336 gnd 0.008448f
C4421 vdd.n3337 gnd 0.010496f
C4422 vdd.n3338 gnd 0.010496f
C4423 vdd.n3339 gnd 0.008448f
C4424 vdd.n3340 gnd 0.008448f
C4425 vdd.n3341 gnd 0.010496f
C4426 vdd.n3342 gnd 0.010496f
C4427 vdd.n3343 gnd 0.008448f
C4428 vdd.n3344 gnd 0.008448f
C4429 vdd.n3345 gnd 0.010496f
C4430 vdd.n3346 gnd 0.010496f
C4431 vdd.n3347 gnd 0.008448f
C4432 vdd.n3348 gnd 0.008448f
C4433 vdd.n3349 gnd 0.010496f
C4434 vdd.n3350 gnd 0.010496f
C4435 vdd.n3351 gnd 0.008448f
C4436 vdd.n3352 gnd 0.008448f
C4437 vdd.n3353 gnd 0.010496f
C4438 vdd.n3354 gnd 0.010496f
C4439 vdd.n3355 gnd 0.008448f
C4440 vdd.n3356 gnd 0.008448f
C4441 vdd.n3357 gnd 0.010496f
C4442 vdd.n3358 gnd 0.010496f
C4443 vdd.n3359 gnd 0.008448f
C4444 vdd.n3360 gnd 0.010496f
C4445 vdd.n3361 gnd 0.010496f
C4446 vdd.n3362 gnd 0.008448f
C4447 vdd.n3363 gnd 0.010496f
C4448 vdd.n3364 gnd 0.010496f
C4449 vdd.n3365 gnd 0.010496f
C4450 vdd.t74 gnd 0.129127f
C4451 vdd.t75 gnd 0.138001f
C4452 vdd.t73 gnd 0.168639f
C4453 vdd.n3366 gnd 0.216171f
C4454 vdd.n3367 gnd 0.181623f
C4455 vdd.n3368 gnd 0.017234f
C4456 vdd.n3369 gnd 0.010496f
C4457 vdd.n3370 gnd 0.010496f
C4458 vdd.n3371 gnd 0.007054f
C4459 vdd.n3372 gnd 0.008448f
C4460 vdd.n3373 gnd 0.010496f
C4461 vdd.n3374 gnd 0.010496f
C4462 vdd.n3375 gnd 0.008448f
C4463 vdd.n3376 gnd 0.008448f
C4464 vdd.n3377 gnd 0.010496f
C4465 vdd.n3378 gnd 0.010496f
C4466 vdd.n3379 gnd 0.008448f
C4467 vdd.n3380 gnd 0.008448f
C4468 vdd.n3381 gnd 0.010496f
C4469 vdd.n3382 gnd 0.010496f
C4470 vdd.n3383 gnd 0.008448f
C4471 vdd.n3384 gnd 0.008448f
C4472 vdd.n3385 gnd 0.010496f
C4473 vdd.n3386 gnd 0.010496f
C4474 vdd.n3387 gnd 0.008448f
C4475 vdd.n3388 gnd 0.008448f
C4476 vdd.n3389 gnd 0.010496f
C4477 vdd.n3390 gnd 0.010496f
C4478 vdd.n3391 gnd 0.008448f
C4479 vdd.n3392 gnd 0.008448f
C4480 vdd.n3393 gnd 0.010496f
C4481 vdd.n3394 gnd 0.010496f
C4482 vdd.n3395 gnd 0.008448f
C4483 vdd.n3396 gnd 0.008448f
C4484 vdd.n3398 gnd 0.958844f
C4485 vdd.n3400 gnd 0.008448f
C4486 vdd.n3401 gnd 0.008448f
C4487 vdd.n3402 gnd 0.007012f
C4488 vdd.n3403 gnd 0.025935f
C4489 vdd.n3405 gnd 11.3163f
C4490 vdd.n3406 gnd 0.025935f
C4491 vdd.n3407 gnd 0.004013f
C4492 vdd.n3408 gnd 0.025935f
C4493 vdd.n3409 gnd 0.02539f
C4494 vdd.n3410 gnd 0.010496f
C4495 vdd.n3411 gnd 0.008448f
C4496 vdd.n3412 gnd 0.010496f
C4497 vdd.n3413 gnd 0.648942f
C4498 vdd.n3414 gnd 0.010496f
C4499 vdd.n3415 gnd 0.008448f
C4500 vdd.n3416 gnd 0.010496f
C4501 vdd.n3417 gnd 0.010496f
C4502 vdd.n3418 gnd 0.010496f
C4503 vdd.n3419 gnd 0.008448f
C4504 vdd.n3420 gnd 0.010496f
C4505 vdd.n3421 gnd 1.07263f
C4506 vdd.n3422 gnd 0.010496f
C4507 vdd.n3423 gnd 0.008448f
C4508 vdd.n3424 gnd 0.010496f
C4509 vdd.n3425 gnd 0.010496f
C4510 vdd.n3426 gnd 0.010496f
C4511 vdd.n3427 gnd 0.008448f
C4512 vdd.n3428 gnd 0.010496f
C4513 vdd.n3429 gnd 0.691848f
C4514 vdd.n3430 gnd 0.734753f
C4515 vdd.n3431 gnd 0.010496f
C4516 vdd.n3432 gnd 0.008448f
C4517 vdd.n3433 gnd 0.010496f
C4518 vdd.n3434 gnd 0.010496f
C4519 vdd.n3435 gnd 0.010496f
C4520 vdd.n3436 gnd 0.008448f
C4521 vdd.n3437 gnd 0.010496f
C4522 vdd.n3438 gnd 0.890285f
C4523 vdd.n3439 gnd 0.010496f
C4524 vdd.n3440 gnd 0.008448f
C4525 vdd.n3441 gnd 0.010496f
C4526 vdd.n3442 gnd 0.010496f
C4527 vdd.n3443 gnd 0.010496f
C4528 vdd.n3444 gnd 0.008448f
C4529 vdd.n3445 gnd 0.010496f
C4530 vdd.t155 gnd 0.536316f
C4531 vdd.n3446 gnd 0.863469f
C4532 vdd.n3447 gnd 0.010496f
C4533 vdd.n3448 gnd 0.008448f
C4534 vdd.n3449 gnd 0.010496f
C4535 vdd.n3450 gnd 0.010496f
C4536 vdd.n3451 gnd 0.010496f
C4537 vdd.n3452 gnd 0.008448f
C4538 vdd.n3453 gnd 0.010496f
C4539 vdd.n3454 gnd 0.681121f
C4540 vdd.n3455 gnd 0.010496f
C4541 vdd.n3456 gnd 0.008448f
C4542 vdd.n3457 gnd 0.010496f
C4543 vdd.n3458 gnd 0.010496f
C4544 vdd.n3459 gnd 0.010496f
C4545 vdd.n3460 gnd 0.008448f
C4546 vdd.n3461 gnd 0.010496f
C4547 vdd.n3462 gnd 0.852743f
C4548 vdd.n3463 gnd 0.573858f
C4549 vdd.n3464 gnd 0.010496f
C4550 vdd.n3465 gnd 0.008448f
C4551 vdd.n3466 gnd 0.010496f
C4552 vdd.n3467 gnd 0.010496f
C4553 vdd.n3468 gnd 0.010496f
C4554 vdd.n3469 gnd 0.008448f
C4555 vdd.n3470 gnd 0.010496f
C4556 vdd.n3471 gnd 0.756206f
C4557 vdd.n3472 gnd 0.010496f
C4558 vdd.n3473 gnd 0.008448f
C4559 vdd.n3474 gnd 0.010496f
C4560 vdd.n3475 gnd 0.010496f
C4561 vdd.n3476 gnd 0.010496f
C4562 vdd.n3477 gnd 0.010496f
C4563 vdd.n3478 gnd 0.010496f
C4564 vdd.n3479 gnd 0.008448f
C4565 vdd.n3480 gnd 0.008448f
C4566 vdd.n3481 gnd 0.010496f
C4567 vdd.t248 gnd 0.536316f
C4568 vdd.n3482 gnd 0.890285f
C4569 vdd.n3483 gnd 0.010496f
C4570 vdd.n3484 gnd 0.008448f
C4571 vdd.n3485 gnd 0.010496f
C4572 vdd.n3486 gnd 0.010496f
C4573 vdd.n3487 gnd 0.010496f
C4574 vdd.n3488 gnd 0.008448f
C4575 vdd.n3489 gnd 0.010496f
C4576 vdd.n3490 gnd 0.842016f
C4577 vdd.n3491 gnd 0.010496f
C4578 vdd.n3492 gnd 0.010496f
C4579 vdd.n3493 gnd 0.008448f
C4580 vdd.n3494 gnd 0.008448f
C4581 vdd.n3495 gnd 0.010496f
C4582 vdd.n3496 gnd 0.010496f
C4583 vdd.n3497 gnd 0.010496f
C4584 vdd.n3498 gnd 0.008448f
C4585 vdd.n3499 gnd 0.010496f
C4586 vdd.n3500 gnd 0.008448f
C4587 vdd.n3501 gnd 0.008448f
C4588 vdd.n3502 gnd 0.010496f
C4589 vdd.n3503 gnd 0.010496f
C4590 vdd.n3504 gnd 0.010496f
C4591 vdd.n3505 gnd 0.008448f
C4592 vdd.n3506 gnd 0.010496f
C4593 vdd.n3507 gnd 0.008448f
C4594 vdd.n3508 gnd 0.008448f
C4595 vdd.n3509 gnd 0.010496f
C4596 vdd.n3510 gnd 0.010496f
C4597 vdd.n3511 gnd 0.010496f
C4598 vdd.n3512 gnd 0.008448f
C4599 vdd.n3513 gnd 0.890285f
C4600 vdd.n3514 gnd 0.010496f
C4601 vdd.n3515 gnd 0.008448f
C4602 vdd.n3516 gnd 0.008448f
C4603 vdd.n3517 gnd 0.010496f
C4604 vdd.n3518 gnd 0.010496f
C4605 vdd.n3519 gnd 0.010496f
C4606 vdd.n3520 gnd 0.008448f
C4607 vdd.n3521 gnd 0.010496f
C4608 vdd.n3522 gnd 0.008448f
C4609 vdd.n3523 gnd 0.008448f
C4610 vdd.n3524 gnd 0.010496f
C4611 vdd.n3525 gnd 0.010496f
C4612 vdd.n3526 gnd 0.010496f
C4613 vdd.n3527 gnd 0.008448f
C4614 vdd.n3528 gnd 0.010496f
C4615 vdd.n3529 gnd 0.008448f
C4616 vdd.n3530 gnd 0.007012f
C4617 vdd.n3531 gnd 0.02539f
C4618 vdd.n3532 gnd 0.025935f
C4619 vdd.n3533 gnd 0.004013f
C4620 vdd.n3534 gnd 0.025935f
C4621 vdd.n3536 gnd 2.54214f
C4622 vdd.n3537 gnd 1.58213f
C4623 vdd.n3538 gnd 0.02539f
C4624 vdd.n3539 gnd 0.007012f
C4625 vdd.n3540 gnd 0.008448f
C4626 vdd.n3541 gnd 0.008448f
C4627 vdd.n3542 gnd 0.010496f
C4628 vdd.n3543 gnd 1.07263f
C4629 vdd.n3544 gnd 1.07263f
C4630 vdd.n3545 gnd 0.981458f
C4631 vdd.n3546 gnd 0.010496f
C4632 vdd.n3547 gnd 0.008448f
C4633 vdd.n3548 gnd 0.008448f
C4634 vdd.n3549 gnd 0.008448f
C4635 vdd.n3550 gnd 0.010496f
C4636 vdd.n3551 gnd 0.799111f
C4637 vdd.t272 gnd 0.536316f
C4638 vdd.n3552 gnd 0.809837f
C4639 vdd.n3553 gnd 0.616763f
C4640 vdd.n3554 gnd 0.010496f
C4641 vdd.n3555 gnd 0.008448f
C4642 vdd.n3556 gnd 0.008448f
C4643 vdd.n3557 gnd 0.008448f
C4644 vdd.n3558 gnd 0.010496f
C4645 vdd.n3559 gnd 0.638216f
C4646 vdd.n3560 gnd 0.788385f
C4647 vdd.t149 gnd 0.536316f
C4648 vdd.n3561 gnd 0.820564f
C4649 vdd.n3562 gnd 0.010496f
C4650 vdd.n3563 gnd 0.008448f
C4651 vdd.n3564 gnd 0.008448f
C4652 vdd.n3565 gnd 0.008448f
C4653 vdd.n3566 gnd 0.010496f
C4654 vdd.n3567 gnd 0.890285f
C4655 vdd.t190 gnd 0.536316f
C4656 vdd.n3568 gnd 0.648942f
C4657 vdd.n3569 gnd 0.777658f
C4658 vdd.n3570 gnd 0.010496f
C4659 vdd.n3571 gnd 0.008448f
C4660 vdd.n3572 gnd 0.008448f
C4661 vdd.n3573 gnd 0.008448f
C4662 vdd.n3574 gnd 0.010496f
C4663 vdd.n3575 gnd 0.595311f
C4664 vdd.t202 gnd 0.536316f
C4665 vdd.n3576 gnd 0.890285f
C4666 vdd.t217 gnd 0.536316f
C4667 vdd.n3577 gnd 0.659669f
C4668 vdd.n3578 gnd 0.010496f
C4669 vdd.n3579 gnd 0.008448f
C4670 vdd.n3580 gnd 0.008067f
C4671 vdd.n3581 gnd 0.619088f
C4672 vdd.n3582 gnd 2.93817f
C4673 a_n8964_8799.n0 gnd 0.211341f
C4674 a_n8964_8799.n1 gnd 0.290199f
C4675 a_n8964_8799.n2 gnd 0.211341f
C4676 a_n8964_8799.n3 gnd 0.211341f
C4677 a_n8964_8799.n4 gnd 0.211341f
C4678 a_n8964_8799.n5 gnd 0.211341f
C4679 a_n8964_8799.n6 gnd 0.211341f
C4680 a_n8964_8799.n7 gnd 0.219756f
C4681 a_n8964_8799.n8 gnd 0.211341f
C4682 a_n8964_8799.n9 gnd 0.290199f
C4683 a_n8964_8799.n10 gnd 0.211341f
C4684 a_n8964_8799.n11 gnd 0.211341f
C4685 a_n8964_8799.n12 gnd 0.211341f
C4686 a_n8964_8799.n13 gnd 0.211341f
C4687 a_n8964_8799.n14 gnd 0.211341f
C4688 a_n8964_8799.n15 gnd 0.219756f
C4689 a_n8964_8799.n16 gnd 0.211341f
C4690 a_n8964_8799.n17 gnd 0.458068f
C4691 a_n8964_8799.n18 gnd 0.211341f
C4692 a_n8964_8799.n19 gnd 0.211341f
C4693 a_n8964_8799.n20 gnd 0.211341f
C4694 a_n8964_8799.n21 gnd 0.211341f
C4695 a_n8964_8799.n22 gnd 0.211341f
C4696 a_n8964_8799.n23 gnd 0.219756f
C4697 a_n8964_8799.n24 gnd 0.211341f
C4698 a_n8964_8799.n25 gnd 0.325427f
C4699 a_n8964_8799.n26 gnd 0.211341f
C4700 a_n8964_8799.n27 gnd 0.211341f
C4701 a_n8964_8799.n28 gnd 0.211341f
C4702 a_n8964_8799.n29 gnd 0.211341f
C4703 a_n8964_8799.n30 gnd 0.211341f
C4704 a_n8964_8799.n31 gnd 0.184528f
C4705 a_n8964_8799.n32 gnd 0.211341f
C4706 a_n8964_8799.n33 gnd 0.325427f
C4707 a_n8964_8799.n34 gnd 0.211341f
C4708 a_n8964_8799.n35 gnd 0.211341f
C4709 a_n8964_8799.n36 gnd 0.211341f
C4710 a_n8964_8799.n37 gnd 0.211341f
C4711 a_n8964_8799.n38 gnd 0.211341f
C4712 a_n8964_8799.n39 gnd 0.184528f
C4713 a_n8964_8799.n40 gnd 0.211341f
C4714 a_n8964_8799.n41 gnd 0.325427f
C4715 a_n8964_8799.n42 gnd 0.211341f
C4716 a_n8964_8799.n43 gnd 0.211341f
C4717 a_n8964_8799.n44 gnd 0.211341f
C4718 a_n8964_8799.n45 gnd 0.211341f
C4719 a_n8964_8799.n46 gnd 0.211341f
C4720 a_n8964_8799.n47 gnd 0.352398f
C4721 a_n8964_8799.n48 gnd 3.4684f
C4722 a_n8964_8799.n49 gnd 1.7685f
C4723 a_n8964_8799.n50 gnd 3.009f
C4724 a_n8964_8799.n51 gnd 1.54896f
C4725 a_n8964_8799.n52 gnd 2.82598f
C4726 a_n8964_8799.n53 gnd 4.00249f
C4727 a_n8964_8799.n54 gnd 1.54896f
C4728 a_n8964_8799.n55 gnd 0.71152f
C4729 a_n8964_8799.n56 gnd 0.254435f
C4730 a_n8964_8799.n57 gnd 0.00372f
C4731 a_n8964_8799.n58 gnd 0.009805f
C4732 a_n8964_8799.n59 gnd 0.010713f
C4733 a_n8964_8799.n60 gnd 0.005661f
C4734 a_n8964_8799.n62 gnd 0.00475f
C4735 a_n8964_8799.n63 gnd 0.010273f
C4736 a_n8964_8799.n64 gnd 0.010273f
C4737 a_n8964_8799.n65 gnd 0.00475f
C4738 a_n8964_8799.n67 gnd 0.005661f
C4739 a_n8964_8799.n68 gnd 0.010713f
C4740 a_n8964_8799.n69 gnd 0.009805f
C4741 a_n8964_8799.n70 gnd 0.00372f
C4742 a_n8964_8799.n71 gnd 0.254435f
C4743 a_n8964_8799.n72 gnd 0.00372f
C4744 a_n8964_8799.n73 gnd 0.009805f
C4745 a_n8964_8799.n74 gnd 0.010713f
C4746 a_n8964_8799.n75 gnd 0.005661f
C4747 a_n8964_8799.n77 gnd 0.00475f
C4748 a_n8964_8799.n78 gnd 0.010273f
C4749 a_n8964_8799.n79 gnd 0.010273f
C4750 a_n8964_8799.n80 gnd 0.00475f
C4751 a_n8964_8799.n82 gnd 0.005661f
C4752 a_n8964_8799.n83 gnd 0.010713f
C4753 a_n8964_8799.n84 gnd 0.009805f
C4754 a_n8964_8799.n85 gnd 0.00372f
C4755 a_n8964_8799.n86 gnd 0.254435f
C4756 a_n8964_8799.n87 gnd 0.00372f
C4757 a_n8964_8799.n88 gnd 0.009805f
C4758 a_n8964_8799.n89 gnd 0.010713f
C4759 a_n8964_8799.n90 gnd 0.005661f
C4760 a_n8964_8799.n92 gnd 0.00475f
C4761 a_n8964_8799.n93 gnd 0.010273f
C4762 a_n8964_8799.n94 gnd 0.010273f
C4763 a_n8964_8799.n95 gnd 0.00475f
C4764 a_n8964_8799.n97 gnd 0.005661f
C4765 a_n8964_8799.n98 gnd 0.010713f
C4766 a_n8964_8799.n99 gnd 0.009805f
C4767 a_n8964_8799.n100 gnd 0.00372f
C4768 a_n8964_8799.n101 gnd 0.00372f
C4769 a_n8964_8799.n102 gnd 0.009805f
C4770 a_n8964_8799.n103 gnd 0.010713f
C4771 a_n8964_8799.n104 gnd 0.005661f
C4772 a_n8964_8799.n106 gnd 0.00475f
C4773 a_n8964_8799.n107 gnd 0.010273f
C4774 a_n8964_8799.n108 gnd 0.010273f
C4775 a_n8964_8799.n109 gnd 0.00475f
C4776 a_n8964_8799.n111 gnd 0.005661f
C4777 a_n8964_8799.n112 gnd 0.010713f
C4778 a_n8964_8799.n113 gnd 0.009805f
C4779 a_n8964_8799.n114 gnd 0.00372f
C4780 a_n8964_8799.n115 gnd 0.254435f
C4781 a_n8964_8799.n116 gnd 0.00372f
C4782 a_n8964_8799.n117 gnd 0.009805f
C4783 a_n8964_8799.n118 gnd 0.010713f
C4784 a_n8964_8799.n119 gnd 0.005661f
C4785 a_n8964_8799.n121 gnd 0.00475f
C4786 a_n8964_8799.n122 gnd 0.010273f
C4787 a_n8964_8799.n123 gnd 0.010273f
C4788 a_n8964_8799.n124 gnd 0.00475f
C4789 a_n8964_8799.n126 gnd 0.005661f
C4790 a_n8964_8799.n127 gnd 0.010713f
C4791 a_n8964_8799.n128 gnd 0.009805f
C4792 a_n8964_8799.n129 gnd 0.00372f
C4793 a_n8964_8799.n130 gnd 0.254435f
C4794 a_n8964_8799.n131 gnd 0.00372f
C4795 a_n8964_8799.n132 gnd 0.009805f
C4796 a_n8964_8799.n133 gnd 0.010713f
C4797 a_n8964_8799.n134 gnd 0.005661f
C4798 a_n8964_8799.n136 gnd 0.00475f
C4799 a_n8964_8799.n137 gnd 0.010273f
C4800 a_n8964_8799.n138 gnd 0.010273f
C4801 a_n8964_8799.n139 gnd 0.00475f
C4802 a_n8964_8799.n141 gnd 0.005661f
C4803 a_n8964_8799.n142 gnd 0.010713f
C4804 a_n8964_8799.n143 gnd 0.009805f
C4805 a_n8964_8799.n144 gnd 0.00372f
C4806 a_n8964_8799.n145 gnd 0.254435f
C4807 a_n8964_8799.t17 gnd 0.146589f
C4808 a_n8964_8799.t8 gnd 0.146589f
C4809 a_n8964_8799.t7 gnd 0.146589f
C4810 a_n8964_8799.n146 gnd 1.15617f
C4811 a_n8964_8799.t29 gnd 0.146589f
C4812 a_n8964_8799.t21 gnd 0.146589f
C4813 a_n8964_8799.n147 gnd 1.15426f
C4814 a_n8964_8799.t28 gnd 0.146589f
C4815 a_n8964_8799.t24 gnd 0.146589f
C4816 a_n8964_8799.n148 gnd 1.15426f
C4817 a_n8964_8799.t26 gnd 0.146589f
C4818 a_n8964_8799.t36 gnd 0.146589f
C4819 a_n8964_8799.n149 gnd 1.15426f
C4820 a_n8964_8799.t25 gnd 0.146589f
C4821 a_n8964_8799.t41 gnd 0.146589f
C4822 a_n8964_8799.n150 gnd 1.15426f
C4823 a_n8964_8799.t14 gnd 0.114013f
C4824 a_n8964_8799.t30 gnd 0.114013f
C4825 a_n8964_8799.n151 gnd 1.00907f
C4826 a_n8964_8799.t15 gnd 0.114013f
C4827 a_n8964_8799.t0 gnd 0.114013f
C4828 a_n8964_8799.n152 gnd 1.00746f
C4829 a_n8964_8799.t12 gnd 0.114013f
C4830 a_n8964_8799.t38 gnd 0.114013f
C4831 a_n8964_8799.n153 gnd 1.00746f
C4832 a_n8964_8799.t2 gnd 0.114013f
C4833 a_n8964_8799.t31 gnd 0.114013f
C4834 a_n8964_8799.n154 gnd 1.00907f
C4835 a_n8964_8799.t9 gnd 0.114013f
C4836 a_n8964_8799.t3 gnd 0.114013f
C4837 a_n8964_8799.n155 gnd 1.00746f
C4838 a_n8964_8799.t18 gnd 0.114013f
C4839 a_n8964_8799.t5 gnd 0.114013f
C4840 a_n8964_8799.n156 gnd 1.00746f
C4841 a_n8964_8799.t32 gnd 0.114013f
C4842 a_n8964_8799.t11 gnd 0.114013f
C4843 a_n8964_8799.n157 gnd 1.00907f
C4844 a_n8964_8799.t19 gnd 0.114013f
C4845 a_n8964_8799.t1 gnd 0.114013f
C4846 a_n8964_8799.n158 gnd 1.00746f
C4847 a_n8964_8799.t16 gnd 0.114013f
C4848 a_n8964_8799.t10 gnd 0.114013f
C4849 a_n8964_8799.n159 gnd 1.00746f
C4850 a_n8964_8799.t43 gnd 0.114013f
C4851 a_n8964_8799.t39 gnd 0.114013f
C4852 a_n8964_8799.n160 gnd 1.00746f
C4853 a_n8964_8799.t33 gnd 0.114013f
C4854 a_n8964_8799.t13 gnd 0.114013f
C4855 a_n8964_8799.n161 gnd 1.00746f
C4856 a_n8964_8799.t4 gnd 0.114013f
C4857 a_n8964_8799.t22 gnd 0.114013f
C4858 a_n8964_8799.n162 gnd 1.00746f
C4859 a_n8964_8799.t77 gnd 0.607824f
C4860 a_n8964_8799.n163 gnd 0.27365f
C4861 a_n8964_8799.t122 gnd 0.607824f
C4862 a_n8964_8799.t145 gnd 0.607824f
C4863 a_n8964_8799.n164 gnd 0.275611f
C4864 a_n8964_8799.t90 gnd 0.607824f
C4865 a_n8964_8799.t93 gnd 0.607824f
C4866 a_n8964_8799.n165 gnd 0.268697f
C4867 a_n8964_8799.t146 gnd 0.607824f
C4868 a_n8964_8799.t151 gnd 0.607824f
C4869 a_n8964_8799.n166 gnd 0.272742f
C4870 a_n8964_8799.t76 gnd 0.607824f
C4871 a_n8964_8799.t121 gnd 0.607824f
C4872 a_n8964_8799.t91 gnd 0.619328f
C4873 a_n8964_8799.n167 gnd 0.254804f
C4874 a_n8964_8799.n168 gnd 0.275989f
C4875 a_n8964_8799.t48 gnd 0.607824f
C4876 a_n8964_8799.n169 gnd 0.27365f
C4877 a_n8964_8799.n170 gnd 0.269348f
C4878 a_n8964_8799.t114 gnd 0.607824f
C4879 a_n8964_8799.n171 gnd 0.268045f
C4880 a_n8964_8799.t74 gnd 0.607824f
C4881 a_n8964_8799.n172 gnd 0.275351f
C4882 a_n8964_8799.t109 gnd 0.607824f
C4883 a_n8964_8799.n173 gnd 0.275611f
C4884 a_n8964_8799.n174 gnd 0.273182f
C4885 a_n8964_8799.t147 gnd 0.607824f
C4886 a_n8964_8799.n175 gnd 0.268697f
C4887 a_n8964_8799.t125 gnd 0.607824f
C4888 a_n8964_8799.n176 gnd 0.273182f
C4889 a_n8964_8799.n177 gnd 0.275351f
C4890 a_n8964_8799.t92 gnd 0.607824f
C4891 a_n8964_8799.n178 gnd 0.272742f
C4892 a_n8964_8799.n179 gnd 0.268045f
C4893 a_n8964_8799.t75 gnd 0.607824f
C4894 a_n8964_8799.n180 gnd 0.269348f
C4895 a_n8964_8799.t118 gnd 0.607824f
C4896 a_n8964_8799.n181 gnd 0.275989f
C4897 a_n8964_8799.t44 gnd 0.619318f
C4898 a_n8964_8799.t88 gnd 0.607824f
C4899 a_n8964_8799.n182 gnd 0.27365f
C4900 a_n8964_8799.t139 gnd 0.607824f
C4901 a_n8964_8799.t158 gnd 0.607824f
C4902 a_n8964_8799.n183 gnd 0.275611f
C4903 a_n8964_8799.t100 gnd 0.607824f
C4904 a_n8964_8799.t105 gnd 0.607824f
C4905 a_n8964_8799.n184 gnd 0.268697f
C4906 a_n8964_8799.t160 gnd 0.607824f
C4907 a_n8964_8799.t163 gnd 0.607824f
C4908 a_n8964_8799.n185 gnd 0.272742f
C4909 a_n8964_8799.t87 gnd 0.607824f
C4910 a_n8964_8799.t138 gnd 0.607824f
C4911 a_n8964_8799.t101 gnd 0.619328f
C4912 a_n8964_8799.n186 gnd 0.254804f
C4913 a_n8964_8799.n187 gnd 0.275989f
C4914 a_n8964_8799.t60 gnd 0.607824f
C4915 a_n8964_8799.n188 gnd 0.27365f
C4916 a_n8964_8799.n189 gnd 0.269348f
C4917 a_n8964_8799.t129 gnd 0.607824f
C4918 a_n8964_8799.n190 gnd 0.268045f
C4919 a_n8964_8799.t83 gnd 0.607824f
C4920 a_n8964_8799.n191 gnd 0.275351f
C4921 a_n8964_8799.t123 gnd 0.607824f
C4922 a_n8964_8799.n192 gnd 0.275611f
C4923 a_n8964_8799.n193 gnd 0.273182f
C4924 a_n8964_8799.t162 gnd 0.607824f
C4925 a_n8964_8799.n194 gnd 0.268697f
C4926 a_n8964_8799.t142 gnd 0.607824f
C4927 a_n8964_8799.n195 gnd 0.273182f
C4928 a_n8964_8799.n196 gnd 0.275351f
C4929 a_n8964_8799.t102 gnd 0.607824f
C4930 a_n8964_8799.n197 gnd 0.272742f
C4931 a_n8964_8799.n198 gnd 0.268045f
C4932 a_n8964_8799.t86 gnd 0.607824f
C4933 a_n8964_8799.n199 gnd 0.269348f
C4934 a_n8964_8799.t136 gnd 0.607824f
C4935 a_n8964_8799.n200 gnd 0.275989f
C4936 a_n8964_8799.t56 gnd 0.619318f
C4937 a_n8964_8799.n201 gnd 0.913779f
C4938 a_n8964_8799.t124 gnd 0.607824f
C4939 a_n8964_8799.n202 gnd 0.27365f
C4940 a_n8964_8799.t106 gnd 0.607824f
C4941 a_n8964_8799.t148 gnd 0.607824f
C4942 a_n8964_8799.n203 gnd 0.275611f
C4943 a_n8964_8799.t66 gnd 0.607824f
C4944 a_n8964_8799.t141 gnd 0.607824f
C4945 a_n8964_8799.n204 gnd 0.268697f
C4946 a_n8964_8799.t119 gnd 0.607824f
C4947 a_n8964_8799.t79 gnd 0.607824f
C4948 a_n8964_8799.n205 gnd 0.272742f
C4949 a_n8964_8799.t64 gnd 0.607824f
C4950 a_n8964_8799.t49 gnd 0.607824f
C4951 a_n8964_8799.t94 gnd 0.619328f
C4952 a_n8964_8799.n206 gnd 0.254804f
C4953 a_n8964_8799.n207 gnd 0.275989f
C4954 a_n8964_8799.t110 gnd 0.607824f
C4955 a_n8964_8799.n208 gnd 0.27365f
C4956 a_n8964_8799.n209 gnd 0.269348f
C4957 a_n8964_8799.t131 gnd 0.607824f
C4958 a_n8964_8799.n210 gnd 0.268045f
C4959 a_n8964_8799.t103 gnd 0.607824f
C4960 a_n8964_8799.n211 gnd 0.275351f
C4961 a_n8964_8799.t57 gnd 0.607824f
C4962 a_n8964_8799.n212 gnd 0.275611f
C4963 a_n8964_8799.n213 gnd 0.273182f
C4964 a_n8964_8799.t98 gnd 0.607824f
C4965 a_n8964_8799.n214 gnd 0.268697f
C4966 a_n8964_8799.t84 gnd 0.607824f
C4967 a_n8964_8799.n215 gnd 0.273182f
C4968 a_n8964_8799.n216 gnd 0.275351f
C4969 a_n8964_8799.t45 gnd 0.607824f
C4970 a_n8964_8799.n217 gnd 0.272742f
C4971 a_n8964_8799.n218 gnd 0.268045f
C4972 a_n8964_8799.t150 gnd 0.607824f
C4973 a_n8964_8799.n219 gnd 0.269348f
C4974 a_n8964_8799.t157 gnd 0.607824f
C4975 a_n8964_8799.n220 gnd 0.275989f
C4976 a_n8964_8799.t99 gnd 0.619318f
C4977 a_n8964_8799.n221 gnd 1.7332f
C4978 a_n8964_8799.t111 gnd 0.619318f
C4979 a_n8964_8799.t47 gnd 0.607824f
C4980 a_n8964_8799.t117 gnd 0.607824f
C4981 a_n8964_8799.n222 gnd 0.27365f
C4982 a_n8964_8799.t115 gnd 0.607824f
C4983 a_n8964_8799.t53 gnd 0.607824f
C4984 a_n8964_8799.t51 gnd 0.607824f
C4985 a_n8964_8799.n223 gnd 0.272742f
C4986 a_n8964_8799.t137 gnd 0.607824f
C4987 a_n8964_8799.t69 gnd 0.607824f
C4988 a_n8964_8799.t55 gnd 0.607824f
C4989 a_n8964_8799.n224 gnd 0.273182f
C4990 a_n8964_8799.t143 gnd 0.607824f
C4991 a_n8964_8799.t95 gnd 0.607824f
C4992 a_n8964_8799.t70 gnd 0.607824f
C4993 a_n8964_8799.n225 gnd 0.273182f
C4994 a_n8964_8799.t161 gnd 0.607824f
C4995 a_n8964_8799.t113 gnd 0.607824f
C4996 a_n8964_8799.t72 gnd 0.607824f
C4997 a_n8964_8799.n226 gnd 0.272742f
C4998 a_n8964_8799.t155 gnd 0.607824f
C4999 a_n8964_8799.t116 gnd 0.607824f
C5000 a_n8964_8799.t89 gnd 0.607824f
C5001 a_n8964_8799.n227 gnd 0.27365f
C5002 a_n8964_8799.t140 gnd 0.619328f
C5003 a_n8964_8799.n228 gnd 0.254804f
C5004 a_n8964_8799.t52 gnd 0.607824f
C5005 a_n8964_8799.n229 gnd 0.275989f
C5006 a_n8964_8799.n230 gnd 0.269348f
C5007 a_n8964_8799.n231 gnd 0.268045f
C5008 a_n8964_8799.n232 gnd 0.275351f
C5009 a_n8964_8799.n233 gnd 0.275611f
C5010 a_n8964_8799.n234 gnd 0.268697f
C5011 a_n8964_8799.n235 gnd 0.268697f
C5012 a_n8964_8799.n236 gnd 0.275611f
C5013 a_n8964_8799.n237 gnd 0.275351f
C5014 a_n8964_8799.n238 gnd 0.268045f
C5015 a_n8964_8799.n239 gnd 0.269348f
C5016 a_n8964_8799.n240 gnd 0.275989f
C5017 a_n8964_8799.t127 gnd 0.619318f
C5018 a_n8964_8799.t59 gnd 0.607824f
C5019 a_n8964_8799.t135 gnd 0.607824f
C5020 a_n8964_8799.n241 gnd 0.27365f
C5021 a_n8964_8799.t133 gnd 0.607824f
C5022 a_n8964_8799.t62 gnd 0.607824f
C5023 a_n8964_8799.t61 gnd 0.607824f
C5024 a_n8964_8799.n242 gnd 0.272742f
C5025 a_n8964_8799.t153 gnd 0.607824f
C5026 a_n8964_8799.t78 gnd 0.607824f
C5027 a_n8964_8799.t68 gnd 0.607824f
C5028 a_n8964_8799.n243 gnd 0.273182f
C5029 a_n8964_8799.t156 gnd 0.607824f
C5030 a_n8964_8799.t108 gnd 0.607824f
C5031 a_n8964_8799.t81 gnd 0.607824f
C5032 a_n8964_8799.n244 gnd 0.273182f
C5033 a_n8964_8799.t54 gnd 0.607824f
C5034 a_n8964_8799.t128 gnd 0.607824f
C5035 a_n8964_8799.t82 gnd 0.607824f
C5036 a_n8964_8799.n245 gnd 0.272742f
C5037 a_n8964_8799.t46 gnd 0.607824f
C5038 a_n8964_8799.t134 gnd 0.607824f
C5039 a_n8964_8799.t97 gnd 0.607824f
C5040 a_n8964_8799.n246 gnd 0.27365f
C5041 a_n8964_8799.t154 gnd 0.619328f
C5042 a_n8964_8799.n247 gnd 0.254804f
C5043 a_n8964_8799.t63 gnd 0.607824f
C5044 a_n8964_8799.n248 gnd 0.275989f
C5045 a_n8964_8799.n249 gnd 0.269348f
C5046 a_n8964_8799.n250 gnd 0.268045f
C5047 a_n8964_8799.n251 gnd 0.275351f
C5048 a_n8964_8799.n252 gnd 0.275611f
C5049 a_n8964_8799.n253 gnd 0.268697f
C5050 a_n8964_8799.n254 gnd 0.268697f
C5051 a_n8964_8799.n255 gnd 0.275611f
C5052 a_n8964_8799.n256 gnd 0.275351f
C5053 a_n8964_8799.n257 gnd 0.268045f
C5054 a_n8964_8799.n258 gnd 0.269348f
C5055 a_n8964_8799.n259 gnd 0.275989f
C5056 a_n8964_8799.n260 gnd 0.913779f
C5057 a_n8964_8799.t73 gnd 0.619318f
C5058 a_n8964_8799.t159 gnd 0.607824f
C5059 a_n8964_8799.t126 gnd 0.607824f
C5060 a_n8964_8799.n261 gnd 0.27365f
C5061 a_n8964_8799.t152 gnd 0.607824f
C5062 a_n8964_8799.t107 gnd 0.607824f
C5063 a_n8964_8799.t132 gnd 0.607824f
C5064 a_n8964_8799.n262 gnd 0.272742f
C5065 a_n8964_8799.t67 gnd 0.607824f
C5066 a_n8964_8799.t149 gnd 0.607824f
C5067 a_n8964_8799.t85 gnd 0.607824f
C5068 a_n8964_8799.n263 gnd 0.273182f
C5069 a_n8964_8799.t144 gnd 0.607824f
C5070 a_n8964_8799.t71 gnd 0.607824f
C5071 a_n8964_8799.t120 gnd 0.607824f
C5072 a_n8964_8799.n264 gnd 0.273182f
C5073 a_n8964_8799.t58 gnd 0.607824f
C5074 a_n8964_8799.t104 gnd 0.607824f
C5075 a_n8964_8799.t80 gnd 0.607824f
C5076 a_n8964_8799.n265 gnd 0.272742f
C5077 a_n8964_8799.t130 gnd 0.607824f
C5078 a_n8964_8799.t65 gnd 0.607824f
C5079 a_n8964_8799.t112 gnd 0.607824f
C5080 a_n8964_8799.n266 gnd 0.27365f
C5081 a_n8964_8799.t96 gnd 0.619328f
C5082 a_n8964_8799.n267 gnd 0.254804f
C5083 a_n8964_8799.t50 gnd 0.607824f
C5084 a_n8964_8799.n268 gnd 0.275989f
C5085 a_n8964_8799.n269 gnd 0.269348f
C5086 a_n8964_8799.n270 gnd 0.268045f
C5087 a_n8964_8799.n271 gnd 0.275351f
C5088 a_n8964_8799.n272 gnd 0.275611f
C5089 a_n8964_8799.n273 gnd 0.268697f
C5090 a_n8964_8799.n274 gnd 0.268697f
C5091 a_n8964_8799.n275 gnd 0.275611f
C5092 a_n8964_8799.n276 gnd 0.275351f
C5093 a_n8964_8799.n277 gnd 0.268045f
C5094 a_n8964_8799.n278 gnd 0.269348f
C5095 a_n8964_8799.n279 gnd 0.275989f
C5096 a_n8964_8799.n280 gnd 1.33295f
C5097 a_n8964_8799.n281 gnd 15.9505f
C5098 a_n8964_8799.n282 gnd 4.44839f
C5099 a_n8964_8799.n283 gnd 7.10849f
C5100 a_n8964_8799.t20 gnd 0.146589f
C5101 a_n8964_8799.t42 gnd 0.146589f
C5102 a_n8964_8799.n284 gnd 1.15426f
C5103 a_n8964_8799.t23 gnd 0.146589f
C5104 a_n8964_8799.t40 gnd 0.146589f
C5105 a_n8964_8799.n285 gnd 1.15426f
C5106 a_n8964_8799.t34 gnd 0.146589f
C5107 a_n8964_8799.t35 gnd 0.146589f
C5108 a_n8964_8799.n286 gnd 1.15426f
C5109 a_n8964_8799.t27 gnd 0.146589f
C5110 a_n8964_8799.t37 gnd 0.146589f
C5111 a_n8964_8799.n287 gnd 1.15616f
C5112 a_n8964_8799.n288 gnd 1.15426f
C5113 a_n8964_8799.t6 gnd 0.146589f
C5114 CSoutput.n0 gnd 0.048592f
C5115 CSoutput.t198 gnd 0.321424f
C5116 CSoutput.n1 gnd 0.145139f
C5117 CSoutput.n2 gnd 0.048592f
C5118 CSoutput.t204 gnd 0.321424f
C5119 CSoutput.n3 gnd 0.038513f
C5120 CSoutput.n4 gnd 0.048592f
C5121 CSoutput.t192 gnd 0.321424f
C5122 CSoutput.n5 gnd 0.03321f
C5123 CSoutput.n6 gnd 0.048592f
C5124 CSoutput.t201 gnd 0.321424f
C5125 CSoutput.t200 gnd 0.321424f
C5126 CSoutput.n7 gnd 0.143557f
C5127 CSoutput.n8 gnd 0.048592f
C5128 CSoutput.t189 gnd 0.321424f
C5129 CSoutput.n9 gnd 0.031664f
C5130 CSoutput.n10 gnd 0.048592f
C5131 CSoutput.t195 gnd 0.321424f
C5132 CSoutput.t197 gnd 0.321424f
C5133 CSoutput.n11 gnd 0.143557f
C5134 CSoutput.n12 gnd 0.048592f
C5135 CSoutput.t187 gnd 0.321424f
C5136 CSoutput.n13 gnd 0.03321f
C5137 CSoutput.n14 gnd 0.048592f
C5138 CSoutput.t185 gnd 0.321424f
C5139 CSoutput.t196 gnd 0.321424f
C5140 CSoutput.n15 gnd 0.143557f
C5141 CSoutput.n16 gnd 0.048592f
C5142 CSoutput.t199 gnd 0.321424f
C5143 CSoutput.n17 gnd 0.03547f
C5144 CSoutput.t188 gnd 0.38411f
C5145 CSoutput.t205 gnd 0.321424f
C5146 CSoutput.n18 gnd 0.183267f
C5147 CSoutput.n19 gnd 0.177832f
C5148 CSoutput.n20 gnd 0.206306f
C5149 CSoutput.n21 gnd 0.048592f
C5150 CSoutput.n22 gnd 0.040555f
C5151 CSoutput.n23 gnd 0.143557f
C5152 CSoutput.n24 gnd 0.039094f
C5153 CSoutput.n25 gnd 0.038513f
C5154 CSoutput.n26 gnd 0.048592f
C5155 CSoutput.n27 gnd 0.048592f
C5156 CSoutput.n28 gnd 0.040243f
C5157 CSoutput.n29 gnd 0.034168f
C5158 CSoutput.n30 gnd 0.146753f
C5159 CSoutput.n31 gnd 0.034638f
C5160 CSoutput.n32 gnd 0.048592f
C5161 CSoutput.n33 gnd 0.048592f
C5162 CSoutput.n34 gnd 0.048592f
C5163 CSoutput.n35 gnd 0.039815f
C5164 CSoutput.n36 gnd 0.143557f
C5165 CSoutput.n37 gnd 0.038077f
C5166 CSoutput.n38 gnd 0.03953f
C5167 CSoutput.n39 gnd 0.048592f
C5168 CSoutput.n40 gnd 0.048592f
C5169 CSoutput.n41 gnd 0.040547f
C5170 CSoutput.n42 gnd 0.03706f
C5171 CSoutput.n43 gnd 0.143557f
C5172 CSoutput.n44 gnd 0.038f
C5173 CSoutput.n45 gnd 0.048592f
C5174 CSoutput.n46 gnd 0.048592f
C5175 CSoutput.n47 gnd 0.048592f
C5176 CSoutput.n48 gnd 0.038f
C5177 CSoutput.n49 gnd 0.143557f
C5178 CSoutput.n50 gnd 0.03706f
C5179 CSoutput.n51 gnd 0.040547f
C5180 CSoutput.n52 gnd 0.048592f
C5181 CSoutput.n53 gnd 0.048592f
C5182 CSoutput.n54 gnd 0.03953f
C5183 CSoutput.n55 gnd 0.038077f
C5184 CSoutput.n56 gnd 0.143557f
C5185 CSoutput.n57 gnd 0.039815f
C5186 CSoutput.n58 gnd 0.048592f
C5187 CSoutput.n59 gnd 0.048592f
C5188 CSoutput.n60 gnd 0.048592f
C5189 CSoutput.n61 gnd 0.034638f
C5190 CSoutput.n62 gnd 0.146753f
C5191 CSoutput.n63 gnd 0.034168f
C5192 CSoutput.t202 gnd 0.321424f
C5193 CSoutput.n64 gnd 0.143557f
C5194 CSoutput.n65 gnd 0.040243f
C5195 CSoutput.n66 gnd 0.048592f
C5196 CSoutput.n67 gnd 0.048592f
C5197 CSoutput.n68 gnd 0.048592f
C5198 CSoutput.n69 gnd 0.039094f
C5199 CSoutput.n70 gnd 0.143557f
C5200 CSoutput.n71 gnd 0.040555f
C5201 CSoutput.n72 gnd 0.03547f
C5202 CSoutput.n73 gnd 0.048592f
C5203 CSoutput.n74 gnd 0.048592f
C5204 CSoutput.n75 gnd 0.036785f
C5205 CSoutput.n76 gnd 0.021847f
C5206 CSoutput.t190 gnd 0.361143f
C5207 CSoutput.n77 gnd 0.179401f
C5208 CSoutput.n78 gnd 0.767641f
C5209 CSoutput.t15 gnd 0.060611f
C5210 CSoutput.t55 gnd 0.060611f
C5211 CSoutput.n79 gnd 0.469273f
C5212 CSoutput.t170 gnd 0.060611f
C5213 CSoutput.t28 gnd 0.060611f
C5214 CSoutput.n80 gnd 0.468436f
C5215 CSoutput.n81 gnd 0.475462f
C5216 CSoutput.t9 gnd 0.060611f
C5217 CSoutput.t70 gnd 0.060611f
C5218 CSoutput.n82 gnd 0.468436f
C5219 CSoutput.n83 gnd 0.234288f
C5220 CSoutput.t47 gnd 0.060611f
C5221 CSoutput.t62 gnd 0.060611f
C5222 CSoutput.n84 gnd 0.468436f
C5223 CSoutput.n85 gnd 0.234288f
C5224 CSoutput.t90 gnd 0.060611f
C5225 CSoutput.t165 gnd 0.060611f
C5226 CSoutput.n86 gnd 0.468436f
C5227 CSoutput.n87 gnd 0.234288f
C5228 CSoutput.t89 gnd 0.060611f
C5229 CSoutput.t183 gnd 0.060611f
C5230 CSoutput.n88 gnd 0.468436f
C5231 CSoutput.n89 gnd 0.234288f
C5232 CSoutput.t60 gnd 0.060611f
C5233 CSoutput.t12 gnd 0.060611f
C5234 CSoutput.n90 gnd 0.468436f
C5235 CSoutput.n91 gnd 0.234288f
C5236 CSoutput.t82 gnd 0.060611f
C5237 CSoutput.t32 gnd 0.060611f
C5238 CSoutput.n92 gnd 0.468436f
C5239 CSoutput.n93 gnd 0.234288f
C5240 CSoutput.t180 gnd 0.060611f
C5241 CSoutput.t35 gnd 0.060611f
C5242 CSoutput.n94 gnd 0.468436f
C5243 CSoutput.n95 gnd 0.234288f
C5244 CSoutput.t3 gnd 0.060611f
C5245 CSoutput.t49 gnd 0.060611f
C5246 CSoutput.n96 gnd 0.468436f
C5247 CSoutput.n97 gnd 0.42963f
C5248 CSoutput.t0 gnd 0.060611f
C5249 CSoutput.t36 gnd 0.060611f
C5250 CSoutput.n98 gnd 0.469273f
C5251 CSoutput.t175 gnd 0.060611f
C5252 CSoutput.t177 gnd 0.060611f
C5253 CSoutput.n99 gnd 0.468436f
C5254 CSoutput.n100 gnd 0.475462f
C5255 CSoutput.t37 gnd 0.060611f
C5256 CSoutput.t75 gnd 0.060611f
C5257 CSoutput.n101 gnd 0.468436f
C5258 CSoutput.n102 gnd 0.234288f
C5259 CSoutput.t41 gnd 0.060611f
C5260 CSoutput.t85 gnd 0.060611f
C5261 CSoutput.n103 gnd 0.468436f
C5262 CSoutput.n104 gnd 0.234288f
C5263 CSoutput.t176 gnd 0.060611f
C5264 CSoutput.t22 gnd 0.060611f
C5265 CSoutput.n105 gnd 0.468436f
C5266 CSoutput.n106 gnd 0.234288f
C5267 CSoutput.t18 gnd 0.060611f
C5268 CSoutput.t65 gnd 0.060611f
C5269 CSoutput.n107 gnd 0.468436f
C5270 CSoutput.n108 gnd 0.234288f
C5271 CSoutput.t30 gnd 0.060611f
C5272 CSoutput.t31 gnd 0.060611f
C5273 CSoutput.n109 gnd 0.468436f
C5274 CSoutput.n110 gnd 0.234288f
C5275 CSoutput.t51 gnd 0.060611f
C5276 CSoutput.t63 gnd 0.060611f
C5277 CSoutput.n111 gnd 0.468436f
C5278 CSoutput.n112 gnd 0.234288f
C5279 CSoutput.t64 gnd 0.060611f
C5280 CSoutput.t83 gnd 0.060611f
C5281 CSoutput.n113 gnd 0.468436f
C5282 CSoutput.n114 gnd 0.234288f
C5283 CSoutput.t67 gnd 0.060611f
C5284 CSoutput.t76 gnd 0.060611f
C5285 CSoutput.n115 gnd 0.468436f
C5286 CSoutput.n116 gnd 0.349382f
C5287 CSoutput.n117 gnd 0.440569f
C5288 CSoutput.t38 gnd 0.060611f
C5289 CSoutput.t71 gnd 0.060611f
C5290 CSoutput.n118 gnd 0.469273f
C5291 CSoutput.t6 gnd 0.060611f
C5292 CSoutput.t21 gnd 0.060611f
C5293 CSoutput.n119 gnd 0.468436f
C5294 CSoutput.n120 gnd 0.475462f
C5295 CSoutput.t182 gnd 0.060611f
C5296 CSoutput.t168 gnd 0.060611f
C5297 CSoutput.n121 gnd 0.468436f
C5298 CSoutput.n122 gnd 0.234288f
C5299 CSoutput.t25 gnd 0.060611f
C5300 CSoutput.t57 gnd 0.060611f
C5301 CSoutput.n123 gnd 0.468436f
C5302 CSoutput.n124 gnd 0.234288f
C5303 CSoutput.t19 gnd 0.060611f
C5304 CSoutput.t163 gnd 0.060611f
C5305 CSoutput.n125 gnd 0.468436f
C5306 CSoutput.n126 gnd 0.234288f
C5307 CSoutput.t39 gnd 0.060611f
C5308 CSoutput.t53 gnd 0.060611f
C5309 CSoutput.n127 gnd 0.468436f
C5310 CSoutput.n128 gnd 0.234288f
C5311 CSoutput.t5 gnd 0.060611f
C5312 CSoutput.t20 gnd 0.060611f
C5313 CSoutput.n129 gnd 0.468436f
C5314 CSoutput.n130 gnd 0.234288f
C5315 CSoutput.t96 gnd 0.060611f
C5316 CSoutput.t14 gnd 0.060611f
C5317 CSoutput.n131 gnd 0.468436f
C5318 CSoutput.n132 gnd 0.234288f
C5319 CSoutput.t174 gnd 0.060611f
C5320 CSoutput.t10 gnd 0.060611f
C5321 CSoutput.n133 gnd 0.468436f
C5322 CSoutput.n134 gnd 0.234288f
C5323 CSoutput.t69 gnd 0.060611f
C5324 CSoutput.t48 gnd 0.060611f
C5325 CSoutput.n135 gnd 0.468436f
C5326 CSoutput.n136 gnd 0.349382f
C5327 CSoutput.n137 gnd 0.492443f
C5328 CSoutput.n138 gnd 9.227429f
C5329 CSoutput.n140 gnd 0.859579f
C5330 CSoutput.n141 gnd 0.644684f
C5331 CSoutput.n142 gnd 0.859579f
C5332 CSoutput.n143 gnd 0.859579f
C5333 CSoutput.n144 gnd 2.31425f
C5334 CSoutput.n145 gnd 0.859579f
C5335 CSoutput.n146 gnd 0.859579f
C5336 CSoutput.t193 gnd 1.07447f
C5337 CSoutput.n147 gnd 0.859579f
C5338 CSoutput.n148 gnd 0.859579f
C5339 CSoutput.n152 gnd 0.859579f
C5340 CSoutput.n156 gnd 0.859579f
C5341 CSoutput.n157 gnd 0.859579f
C5342 CSoutput.n159 gnd 0.859579f
C5343 CSoutput.n164 gnd 0.859579f
C5344 CSoutput.n166 gnd 0.859579f
C5345 CSoutput.n167 gnd 0.859579f
C5346 CSoutput.n169 gnd 0.859579f
C5347 CSoutput.n170 gnd 0.859579f
C5348 CSoutput.n172 gnd 0.859579f
C5349 CSoutput.t186 gnd 14.363501f
C5350 CSoutput.n174 gnd 0.859579f
C5351 CSoutput.n175 gnd 0.644684f
C5352 CSoutput.n176 gnd 0.859579f
C5353 CSoutput.n177 gnd 0.859579f
C5354 CSoutput.n178 gnd 2.31425f
C5355 CSoutput.n179 gnd 0.859579f
C5356 CSoutput.n180 gnd 0.859579f
C5357 CSoutput.t203 gnd 1.07447f
C5358 CSoutput.n181 gnd 0.859579f
C5359 CSoutput.n182 gnd 0.859579f
C5360 CSoutput.n186 gnd 0.859579f
C5361 CSoutput.n190 gnd 0.859579f
C5362 CSoutput.n191 gnd 0.859579f
C5363 CSoutput.n193 gnd 0.859579f
C5364 CSoutput.n198 gnd 0.859579f
C5365 CSoutput.n200 gnd 0.859579f
C5366 CSoutput.n201 gnd 0.859579f
C5367 CSoutput.n203 gnd 0.859579f
C5368 CSoutput.n204 gnd 0.859579f
C5369 CSoutput.n206 gnd 0.859579f
C5370 CSoutput.n207 gnd 0.644684f
C5371 CSoutput.n209 gnd 0.859579f
C5372 CSoutput.n210 gnd 0.644684f
C5373 CSoutput.n211 gnd 0.859579f
C5374 CSoutput.n212 gnd 0.859579f
C5375 CSoutput.n213 gnd 2.31425f
C5376 CSoutput.n214 gnd 0.859579f
C5377 CSoutput.n215 gnd 0.859579f
C5378 CSoutput.t184 gnd 1.07447f
C5379 CSoutput.n216 gnd 0.859579f
C5380 CSoutput.n217 gnd 2.31425f
C5381 CSoutput.n219 gnd 0.859579f
C5382 CSoutput.n220 gnd 0.859579f
C5383 CSoutput.n222 gnd 0.859579f
C5384 CSoutput.n223 gnd 0.859579f
C5385 CSoutput.t194 gnd 14.1294f
C5386 CSoutput.t191 gnd 14.363501f
C5387 CSoutput.n229 gnd 2.69663f
C5388 CSoutput.n230 gnd 10.9851f
C5389 CSoutput.n231 gnd 11.4447f
C5390 CSoutput.n236 gnd 2.92117f
C5391 CSoutput.n242 gnd 0.859579f
C5392 CSoutput.n244 gnd 0.859579f
C5393 CSoutput.n246 gnd 0.859579f
C5394 CSoutput.n248 gnd 0.859579f
C5395 CSoutput.n250 gnd 0.859579f
C5396 CSoutput.n256 gnd 0.859579f
C5397 CSoutput.n263 gnd 1.577f
C5398 CSoutput.n264 gnd 1.577f
C5399 CSoutput.n265 gnd 0.859579f
C5400 CSoutput.n266 gnd 0.859579f
C5401 CSoutput.n268 gnd 0.644684f
C5402 CSoutput.n269 gnd 0.552114f
C5403 CSoutput.n271 gnd 0.644684f
C5404 CSoutput.n272 gnd 0.552114f
C5405 CSoutput.n273 gnd 0.644684f
C5406 CSoutput.n275 gnd 0.859579f
C5407 CSoutput.n277 gnd 2.31425f
C5408 CSoutput.n278 gnd 2.69663f
C5409 CSoutput.n279 gnd 10.1034f
C5410 CSoutput.n281 gnd 0.644684f
C5411 CSoutput.n282 gnd 1.65881f
C5412 CSoutput.n283 gnd 0.644684f
C5413 CSoutput.n285 gnd 0.859579f
C5414 CSoutput.n287 gnd 2.31425f
C5415 CSoutput.n288 gnd 5.04081f
C5416 CSoutput.t45 gnd 0.060611f
C5417 CSoutput.t77 gnd 0.060611f
C5418 CSoutput.n289 gnd 0.469273f
C5419 CSoutput.t16 gnd 0.060611f
C5420 CSoutput.t81 gnd 0.060611f
C5421 CSoutput.n290 gnd 0.468436f
C5422 CSoutput.n291 gnd 0.475462f
C5423 CSoutput.t178 gnd 0.060611f
C5424 CSoutput.t23 gnd 0.060611f
C5425 CSoutput.n292 gnd 0.468436f
C5426 CSoutput.n293 gnd 0.234288f
C5427 CSoutput.t46 gnd 0.060611f
C5428 CSoutput.t86 gnd 0.060611f
C5429 CSoutput.n294 gnd 0.468436f
C5430 CSoutput.n295 gnd 0.234288f
C5431 CSoutput.t61 gnd 0.060611f
C5432 CSoutput.t92 gnd 0.060611f
C5433 CSoutput.n296 gnd 0.468436f
C5434 CSoutput.n297 gnd 0.234288f
C5435 CSoutput.t52 gnd 0.060611f
C5436 CSoutput.t50 gnd 0.060611f
C5437 CSoutput.n298 gnd 0.468436f
C5438 CSoutput.n299 gnd 0.234288f
C5439 CSoutput.t93 gnd 0.060611f
C5440 CSoutput.t68 gnd 0.060611f
C5441 CSoutput.n300 gnd 0.468436f
C5442 CSoutput.n301 gnd 0.234288f
C5443 CSoutput.t11 gnd 0.060611f
C5444 CSoutput.t24 gnd 0.060611f
C5445 CSoutput.n302 gnd 0.468436f
C5446 CSoutput.n303 gnd 0.234288f
C5447 CSoutput.t91 gnd 0.060611f
C5448 CSoutput.t80 gnd 0.060611f
C5449 CSoutput.n304 gnd 0.468436f
C5450 CSoutput.n305 gnd 0.234288f
C5451 CSoutput.t29 gnd 0.060611f
C5452 CSoutput.t79 gnd 0.060611f
C5453 CSoutput.n306 gnd 0.468436f
C5454 CSoutput.n307 gnd 0.42963f
C5455 CSoutput.t27 gnd 0.060611f
C5456 CSoutput.t164 gnd 0.060611f
C5457 CSoutput.n308 gnd 0.469273f
C5458 CSoutput.t173 gnd 0.060611f
C5459 CSoutput.t88 gnd 0.060611f
C5460 CSoutput.n309 gnd 0.468436f
C5461 CSoutput.n310 gnd 0.475462f
C5462 CSoutput.t74 gnd 0.060611f
C5463 CSoutput.t2 gnd 0.060611f
C5464 CSoutput.n311 gnd 0.468436f
C5465 CSoutput.n312 gnd 0.234288f
C5466 CSoutput.t34 gnd 0.060611f
C5467 CSoutput.t171 gnd 0.060611f
C5468 CSoutput.n313 gnd 0.468436f
C5469 CSoutput.n314 gnd 0.234288f
C5470 CSoutput.t54 gnd 0.060611f
C5471 CSoutput.t73 gnd 0.060611f
C5472 CSoutput.n315 gnd 0.468436f
C5473 CSoutput.n316 gnd 0.234288f
C5474 CSoutput.t44 gnd 0.060611f
C5475 CSoutput.t56 gnd 0.060611f
C5476 CSoutput.n317 gnd 0.468436f
C5477 CSoutput.n318 gnd 0.234288f
C5478 CSoutput.t17 gnd 0.060611f
C5479 CSoutput.t13 gnd 0.060611f
C5480 CSoutput.n319 gnd 0.468436f
C5481 CSoutput.n320 gnd 0.234288f
C5482 CSoutput.t94 gnd 0.060611f
C5483 CSoutput.t42 gnd 0.060611f
C5484 CSoutput.n321 gnd 0.468436f
C5485 CSoutput.n322 gnd 0.234288f
C5486 CSoutput.t8 gnd 0.060611f
C5487 CSoutput.t172 gnd 0.060611f
C5488 CSoutput.n323 gnd 0.468436f
C5489 CSoutput.n324 gnd 0.234288f
C5490 CSoutput.t1 gnd 0.060611f
C5491 CSoutput.t66 gnd 0.060611f
C5492 CSoutput.n325 gnd 0.468436f
C5493 CSoutput.n326 gnd 0.349382f
C5494 CSoutput.n327 gnd 0.440569f
C5495 CSoutput.t78 gnd 0.060611f
C5496 CSoutput.t40 gnd 0.060611f
C5497 CSoutput.n328 gnd 0.469273f
C5498 CSoutput.t33 gnd 0.060611f
C5499 CSoutput.t87 gnd 0.060611f
C5500 CSoutput.n329 gnd 0.468436f
C5501 CSoutput.n330 gnd 0.475462f
C5502 CSoutput.t167 gnd 0.060611f
C5503 CSoutput.t169 gnd 0.060611f
C5504 CSoutput.n331 gnd 0.468436f
C5505 CSoutput.n332 gnd 0.234288f
C5506 CSoutput.t4 gnd 0.060611f
C5507 CSoutput.t72 gnd 0.060611f
C5508 CSoutput.n333 gnd 0.468436f
C5509 CSoutput.n334 gnd 0.234288f
C5510 CSoutput.t166 gnd 0.060611f
C5511 CSoutput.t181 gnd 0.060611f
C5512 CSoutput.n335 gnd 0.468436f
C5513 CSoutput.n336 gnd 0.234288f
C5514 CSoutput.t84 gnd 0.060611f
C5515 CSoutput.t7 gnd 0.060611f
C5516 CSoutput.n337 gnd 0.468436f
C5517 CSoutput.n338 gnd 0.234288f
C5518 CSoutput.t43 gnd 0.060611f
C5519 CSoutput.t95 gnd 0.060611f
C5520 CSoutput.n339 gnd 0.468436f
C5521 CSoutput.n340 gnd 0.234288f
C5522 CSoutput.t97 gnd 0.060611f
C5523 CSoutput.t59 gnd 0.060611f
C5524 CSoutput.n341 gnd 0.468436f
C5525 CSoutput.n342 gnd 0.234288f
C5526 CSoutput.t98 gnd 0.060611f
C5527 CSoutput.t179 gnd 0.060611f
C5528 CSoutput.n343 gnd 0.468436f
C5529 CSoutput.n344 gnd 0.234288f
C5530 CSoutput.t58 gnd 0.060611f
C5531 CSoutput.t26 gnd 0.060611f
C5532 CSoutput.n345 gnd 0.468435f
C5533 CSoutput.n346 gnd 0.349384f
C5534 CSoutput.n347 gnd 0.492443f
C5535 CSoutput.n348 gnd 13.177999f
C5536 CSoutput.t134 gnd 0.053035f
C5537 CSoutput.t144 gnd 0.053035f
C5538 CSoutput.n349 gnd 0.470204f
C5539 CSoutput.t102 gnd 0.053035f
C5540 CSoutput.t104 gnd 0.053035f
C5541 CSoutput.n350 gnd 0.468635f
C5542 CSoutput.n351 gnd 0.436681f
C5543 CSoutput.t118 gnd 0.053035f
C5544 CSoutput.t126 gnd 0.053035f
C5545 CSoutput.n352 gnd 0.468635f
C5546 CSoutput.n353 gnd 0.215263f
C5547 CSoutput.t160 gnd 0.053035f
C5548 CSoutput.t135 gnd 0.053035f
C5549 CSoutput.n354 gnd 0.468635f
C5550 CSoutput.n355 gnd 0.215263f
C5551 CSoutput.t108 gnd 0.053035f
C5552 CSoutput.t116 gnd 0.053035f
C5553 CSoutput.n356 gnd 0.468635f
C5554 CSoutput.n357 gnd 0.215263f
C5555 CSoutput.t110 gnd 0.053035f
C5556 CSoutput.t152 gnd 0.053035f
C5557 CSoutput.n358 gnd 0.468635f
C5558 CSoutput.n359 gnd 0.215263f
C5559 CSoutput.t131 gnd 0.053035f
C5560 CSoutput.t142 gnd 0.053035f
C5561 CSoutput.n360 gnd 0.468635f
C5562 CSoutput.n361 gnd 0.215263f
C5563 CSoutput.t99 gnd 0.053035f
C5564 CSoutput.t107 gnd 0.053035f
C5565 CSoutput.n362 gnd 0.468635f
C5566 CSoutput.n363 gnd 0.396988f
C5567 CSoutput.t153 gnd 0.053035f
C5568 CSoutput.t132 gnd 0.053035f
C5569 CSoutput.n364 gnd 0.470204f
C5570 CSoutput.t161 gnd 0.053035f
C5571 CSoutput.t151 gnd 0.053035f
C5572 CSoutput.n365 gnd 0.468635f
C5573 CSoutput.n366 gnd 0.436681f
C5574 CSoutput.t109 gnd 0.053035f
C5575 CSoutput.t117 gnd 0.053035f
C5576 CSoutput.n367 gnd 0.468635f
C5577 CSoutput.n368 gnd 0.215263f
C5578 CSoutput.t150 gnd 0.053035f
C5579 CSoutput.t154 gnd 0.053035f
C5580 CSoutput.n369 gnd 0.468635f
C5581 CSoutput.n370 gnd 0.215263f
C5582 CSoutput.t158 gnd 0.053035f
C5583 CSoutput.t138 gnd 0.053035f
C5584 CSoutput.n371 gnd 0.468635f
C5585 CSoutput.n372 gnd 0.215263f
C5586 CSoutput.t100 gnd 0.053035f
C5587 CSoutput.t103 gnd 0.053035f
C5588 CSoutput.n373 gnd 0.468635f
C5589 CSoutput.n374 gnd 0.215263f
C5590 CSoutput.t113 gnd 0.053035f
C5591 CSoutput.t130 gnd 0.053035f
C5592 CSoutput.n375 gnd 0.468635f
C5593 CSoutput.n376 gnd 0.215263f
C5594 CSoutput.t159 gnd 0.053035f
C5595 CSoutput.t157 gnd 0.053035f
C5596 CSoutput.n377 gnd 0.468635f
C5597 CSoutput.n378 gnd 0.326815f
C5598 CSoutput.n379 gnd 0.607248f
C5599 CSoutput.n380 gnd 13.284401f
C5600 CSoutput.t149 gnd 0.053035f
C5601 CSoutput.t140 gnd 0.053035f
C5602 CSoutput.n381 gnd 0.470204f
C5603 CSoutput.t112 gnd 0.053035f
C5604 CSoutput.t106 gnd 0.053035f
C5605 CSoutput.n382 gnd 0.468635f
C5606 CSoutput.n383 gnd 0.436681f
C5607 CSoutput.t162 gnd 0.053035f
C5608 CSoutput.t125 gnd 0.053035f
C5609 CSoutput.n384 gnd 0.468635f
C5610 CSoutput.n385 gnd 0.215263f
C5611 CSoutput.t141 gnd 0.053035f
C5612 CSoutput.t146 gnd 0.053035f
C5613 CSoutput.n386 gnd 0.468635f
C5614 CSoutput.n387 gnd 0.215263f
C5615 CSoutput.t123 gnd 0.053035f
C5616 CSoutput.t114 gnd 0.053035f
C5617 CSoutput.n388 gnd 0.468635f
C5618 CSoutput.n389 gnd 0.215263f
C5619 CSoutput.t120 gnd 0.053035f
C5620 CSoutput.t156 gnd 0.053035f
C5621 CSoutput.n390 gnd 0.468635f
C5622 CSoutput.n391 gnd 0.215263f
C5623 CSoutput.t147 gnd 0.053035f
C5624 CSoutput.t129 gnd 0.053035f
C5625 CSoutput.n392 gnd 0.468635f
C5626 CSoutput.n393 gnd 0.215263f
C5627 CSoutput.t145 gnd 0.053035f
C5628 CSoutput.t137 gnd 0.053035f
C5629 CSoutput.n394 gnd 0.468635f
C5630 CSoutput.n395 gnd 0.396988f
C5631 CSoutput.t139 gnd 0.053035f
C5632 CSoutput.t121 gnd 0.053035f
C5633 CSoutput.n396 gnd 0.470204f
C5634 CSoutput.t101 gnd 0.053035f
C5635 CSoutput.t148 gnd 0.053035f
C5636 CSoutput.n397 gnd 0.468635f
C5637 CSoutput.n398 gnd 0.436681f
C5638 CSoutput.t124 gnd 0.053035f
C5639 CSoutput.t115 gnd 0.053035f
C5640 CSoutput.n399 gnd 0.468635f
C5641 CSoutput.n400 gnd 0.215263f
C5642 CSoutput.t122 gnd 0.053035f
C5643 CSoutput.t127 gnd 0.053035f
C5644 CSoutput.n401 gnd 0.468635f
C5645 CSoutput.n402 gnd 0.215263f
C5646 CSoutput.t143 gnd 0.053035f
C5647 CSoutput.t136 gnd 0.053035f
C5648 CSoutput.n403 gnd 0.468635f
C5649 CSoutput.n404 gnd 0.215263f
C5650 CSoutput.t111 gnd 0.053035f
C5651 CSoutput.t105 gnd 0.053035f
C5652 CSoutput.n405 gnd 0.468635f
C5653 CSoutput.n406 gnd 0.215263f
C5654 CSoutput.t128 gnd 0.053035f
C5655 CSoutput.t119 gnd 0.053035f
C5656 CSoutput.n407 gnd 0.468635f
C5657 CSoutput.n408 gnd 0.215263f
C5658 CSoutput.t133 gnd 0.053035f
C5659 CSoutput.t155 gnd 0.053035f
C5660 CSoutput.n409 gnd 0.468635f
C5661 CSoutput.n410 gnd 0.326815f
C5662 CSoutput.n411 gnd 0.607248f
C5663 CSoutput.n412 gnd 7.80511f
C5664 CSoutput.n413 gnd 15.498599f
C5665 commonsourceibias.n0 gnd 0.010545f
C5666 commonsourceibias.t94 gnd 0.159685f
C5667 commonsourceibias.t109 gnd 0.147652f
C5668 commonsourceibias.n1 gnd 0.006423f
C5669 commonsourceibias.n2 gnd 0.007903f
C5670 commonsourceibias.t72 gnd 0.147652f
C5671 commonsourceibias.n3 gnd 0.008017f
C5672 commonsourceibias.n4 gnd 0.007903f
C5673 commonsourceibias.t70 gnd 0.147652f
C5674 commonsourceibias.n5 gnd 0.058913f
C5675 commonsourceibias.t102 gnd 0.147652f
C5676 commonsourceibias.n6 gnd 0.006393f
C5677 commonsourceibias.n7 gnd 0.007903f
C5678 commonsourceibias.t118 gnd 0.147652f
C5679 commonsourceibias.n8 gnd 0.00763f
C5680 commonsourceibias.n9 gnd 0.007903f
C5681 commonsourceibias.t66 gnd 0.147652f
C5682 commonsourceibias.n10 gnd 0.058913f
C5683 commonsourceibias.t93 gnd 0.147652f
C5684 commonsourceibias.n11 gnd 0.006383f
C5685 commonsourceibias.n12 gnd 0.010545f
C5686 commonsourceibias.t54 gnd 0.159685f
C5687 commonsourceibias.t24 gnd 0.147652f
C5688 commonsourceibias.n13 gnd 0.006423f
C5689 commonsourceibias.n14 gnd 0.007903f
C5690 commonsourceibias.t14 gnd 0.147652f
C5691 commonsourceibias.n15 gnd 0.008017f
C5692 commonsourceibias.n16 gnd 0.007903f
C5693 commonsourceibias.t52 gnd 0.147652f
C5694 commonsourceibias.n17 gnd 0.058913f
C5695 commonsourceibias.t20 gnd 0.147652f
C5696 commonsourceibias.n18 gnd 0.006393f
C5697 commonsourceibias.n19 gnd 0.007903f
C5698 commonsourceibias.t58 gnd 0.147652f
C5699 commonsourceibias.n20 gnd 0.00763f
C5700 commonsourceibias.n21 gnd 0.007903f
C5701 commonsourceibias.t60 gnd 0.147652f
C5702 commonsourceibias.n22 gnd 0.058913f
C5703 commonsourceibias.t16 gnd 0.147652f
C5704 commonsourceibias.n23 gnd 0.006383f
C5705 commonsourceibias.n24 gnd 0.007903f
C5706 commonsourceibias.t56 gnd 0.147652f
C5707 commonsourceibias.t38 gnd 0.147652f
C5708 commonsourceibias.n25 gnd 0.058913f
C5709 commonsourceibias.n26 gnd 0.007903f
C5710 commonsourceibias.t6 gnd 0.147652f
C5711 commonsourceibias.n27 gnd 0.058913f
C5712 commonsourceibias.n28 gnd 0.007903f
C5713 commonsourceibias.t62 gnd 0.147652f
C5714 commonsourceibias.n29 gnd 0.058913f
C5715 commonsourceibias.n30 gnd 0.007903f
C5716 commonsourceibias.t32 gnd 0.147652f
C5717 commonsourceibias.n31 gnd 0.008983f
C5718 commonsourceibias.n32 gnd 0.007903f
C5719 commonsourceibias.t0 gnd 0.147652f
C5720 commonsourceibias.n33 gnd 0.010623f
C5721 commonsourceibias.t10 gnd 0.164481f
C5722 commonsourceibias.t26 gnd 0.147652f
C5723 commonsourceibias.n34 gnd 0.065644f
C5724 commonsourceibias.n35 gnd 0.070328f
C5725 commonsourceibias.n36 gnd 0.033639f
C5726 commonsourceibias.n37 gnd 0.007903f
C5727 commonsourceibias.n38 gnd 0.006423f
C5728 commonsourceibias.n39 gnd 0.01089f
C5729 commonsourceibias.n40 gnd 0.058913f
C5730 commonsourceibias.n41 gnd 0.010937f
C5731 commonsourceibias.n42 gnd 0.007903f
C5732 commonsourceibias.n43 gnd 0.007903f
C5733 commonsourceibias.n44 gnd 0.007903f
C5734 commonsourceibias.n45 gnd 0.008017f
C5735 commonsourceibias.n46 gnd 0.058913f
C5736 commonsourceibias.n47 gnd 0.009741f
C5737 commonsourceibias.n48 gnd 0.010776f
C5738 commonsourceibias.n49 gnd 0.007903f
C5739 commonsourceibias.n50 gnd 0.007903f
C5740 commonsourceibias.n51 gnd 0.010705f
C5741 commonsourceibias.n52 gnd 0.006393f
C5742 commonsourceibias.n53 gnd 0.010838f
C5743 commonsourceibias.n54 gnd 0.007903f
C5744 commonsourceibias.n55 gnd 0.007903f
C5745 commonsourceibias.n56 gnd 0.010904f
C5746 commonsourceibias.n57 gnd 0.009403f
C5747 commonsourceibias.n58 gnd 0.00763f
C5748 commonsourceibias.n59 gnd 0.007903f
C5749 commonsourceibias.n60 gnd 0.007903f
C5750 commonsourceibias.n61 gnd 0.009667f
C5751 commonsourceibias.n62 gnd 0.01085f
C5752 commonsourceibias.n63 gnd 0.058913f
C5753 commonsourceibias.n64 gnd 0.010777f
C5754 commonsourceibias.n65 gnd 0.007903f
C5755 commonsourceibias.n66 gnd 0.007903f
C5756 commonsourceibias.n67 gnd 0.007903f
C5757 commonsourceibias.n68 gnd 0.010777f
C5758 commonsourceibias.n69 gnd 0.058913f
C5759 commonsourceibias.n70 gnd 0.01085f
C5760 commonsourceibias.n71 gnd 0.009667f
C5761 commonsourceibias.n72 gnd 0.007903f
C5762 commonsourceibias.n73 gnd 0.007903f
C5763 commonsourceibias.n74 gnd 0.007903f
C5764 commonsourceibias.n75 gnd 0.009403f
C5765 commonsourceibias.n76 gnd 0.010904f
C5766 commonsourceibias.n77 gnd 0.058913f
C5767 commonsourceibias.n78 gnd 0.010838f
C5768 commonsourceibias.n79 gnd 0.007903f
C5769 commonsourceibias.n80 gnd 0.007903f
C5770 commonsourceibias.n81 gnd 0.007903f
C5771 commonsourceibias.n82 gnd 0.010705f
C5772 commonsourceibias.n83 gnd 0.058913f
C5773 commonsourceibias.n84 gnd 0.010776f
C5774 commonsourceibias.n85 gnd 0.009741f
C5775 commonsourceibias.n86 gnd 0.007903f
C5776 commonsourceibias.n87 gnd 0.007903f
C5777 commonsourceibias.n88 gnd 0.007903f
C5778 commonsourceibias.n89 gnd 0.008983f
C5779 commonsourceibias.n90 gnd 0.010937f
C5780 commonsourceibias.n91 gnd 0.058913f
C5781 commonsourceibias.n92 gnd 0.01089f
C5782 commonsourceibias.n93 gnd 0.007903f
C5783 commonsourceibias.n94 gnd 0.007903f
C5784 commonsourceibias.n95 gnd 0.007903f
C5785 commonsourceibias.n96 gnd 0.010623f
C5786 commonsourceibias.n97 gnd 0.058913f
C5787 commonsourceibias.n98 gnd 0.010649f
C5788 commonsourceibias.n99 gnd 0.071041f
C5789 commonsourceibias.n100 gnd 0.079434f
C5790 commonsourceibias.t55 gnd 0.017054f
C5791 commonsourceibias.t25 gnd 0.017054f
C5792 commonsourceibias.n101 gnd 0.150693f
C5793 commonsourceibias.n102 gnd 0.130533f
C5794 commonsourceibias.t15 gnd 0.017054f
C5795 commonsourceibias.t53 gnd 0.017054f
C5796 commonsourceibias.n103 gnd 0.150693f
C5797 commonsourceibias.n104 gnd 0.069219f
C5798 commonsourceibias.t21 gnd 0.017054f
C5799 commonsourceibias.t59 gnd 0.017054f
C5800 commonsourceibias.n105 gnd 0.150693f
C5801 commonsourceibias.n106 gnd 0.069219f
C5802 commonsourceibias.t61 gnd 0.017054f
C5803 commonsourceibias.t17 gnd 0.017054f
C5804 commonsourceibias.n107 gnd 0.150693f
C5805 commonsourceibias.n108 gnd 0.057829f
C5806 commonsourceibias.t27 gnd 0.017054f
C5807 commonsourceibias.t11 gnd 0.017054f
C5808 commonsourceibias.n109 gnd 0.151197f
C5809 commonsourceibias.t33 gnd 0.017054f
C5810 commonsourceibias.t1 gnd 0.017054f
C5811 commonsourceibias.n110 gnd 0.150693f
C5812 commonsourceibias.n111 gnd 0.140418f
C5813 commonsourceibias.t7 gnd 0.017054f
C5814 commonsourceibias.t63 gnd 0.017054f
C5815 commonsourceibias.n112 gnd 0.150693f
C5816 commonsourceibias.n113 gnd 0.069219f
C5817 commonsourceibias.t57 gnd 0.017054f
C5818 commonsourceibias.t39 gnd 0.017054f
C5819 commonsourceibias.n114 gnd 0.150693f
C5820 commonsourceibias.n115 gnd 0.057829f
C5821 commonsourceibias.n116 gnd 0.070025f
C5822 commonsourceibias.n117 gnd 0.007903f
C5823 commonsourceibias.t88 gnd 0.147652f
C5824 commonsourceibias.t105 gnd 0.147652f
C5825 commonsourceibias.n118 gnd 0.058913f
C5826 commonsourceibias.n119 gnd 0.007903f
C5827 commonsourceibias.t86 gnd 0.147652f
C5828 commonsourceibias.n120 gnd 0.058913f
C5829 commonsourceibias.n121 gnd 0.007903f
C5830 commonsourceibias.t82 gnd 0.147652f
C5831 commonsourceibias.n122 gnd 0.058913f
C5832 commonsourceibias.n123 gnd 0.007903f
C5833 commonsourceibias.t97 gnd 0.147652f
C5834 commonsourceibias.n124 gnd 0.008983f
C5835 commonsourceibias.n125 gnd 0.007903f
C5836 commonsourceibias.t111 gnd 0.147652f
C5837 commonsourceibias.n126 gnd 0.010623f
C5838 commonsourceibias.t89 gnd 0.164481f
C5839 commonsourceibias.t75 gnd 0.147652f
C5840 commonsourceibias.n127 gnd 0.065644f
C5841 commonsourceibias.n128 gnd 0.070328f
C5842 commonsourceibias.n129 gnd 0.033639f
C5843 commonsourceibias.n130 gnd 0.007903f
C5844 commonsourceibias.n131 gnd 0.006423f
C5845 commonsourceibias.n132 gnd 0.01089f
C5846 commonsourceibias.n133 gnd 0.058913f
C5847 commonsourceibias.n134 gnd 0.010937f
C5848 commonsourceibias.n135 gnd 0.007903f
C5849 commonsourceibias.n136 gnd 0.007903f
C5850 commonsourceibias.n137 gnd 0.007903f
C5851 commonsourceibias.n138 gnd 0.008017f
C5852 commonsourceibias.n139 gnd 0.058913f
C5853 commonsourceibias.n140 gnd 0.009741f
C5854 commonsourceibias.n141 gnd 0.010776f
C5855 commonsourceibias.n142 gnd 0.007903f
C5856 commonsourceibias.n143 gnd 0.007903f
C5857 commonsourceibias.n144 gnd 0.010705f
C5858 commonsourceibias.n145 gnd 0.006393f
C5859 commonsourceibias.n146 gnd 0.010838f
C5860 commonsourceibias.n147 gnd 0.007903f
C5861 commonsourceibias.n148 gnd 0.007903f
C5862 commonsourceibias.n149 gnd 0.010904f
C5863 commonsourceibias.n150 gnd 0.009403f
C5864 commonsourceibias.n151 gnd 0.00763f
C5865 commonsourceibias.n152 gnd 0.007903f
C5866 commonsourceibias.n153 gnd 0.007903f
C5867 commonsourceibias.n154 gnd 0.009667f
C5868 commonsourceibias.n155 gnd 0.01085f
C5869 commonsourceibias.n156 gnd 0.058913f
C5870 commonsourceibias.n157 gnd 0.010777f
C5871 commonsourceibias.n158 gnd 0.007865f
C5872 commonsourceibias.n159 gnd 0.057129f
C5873 commonsourceibias.n160 gnd 0.007865f
C5874 commonsourceibias.n161 gnd 0.010777f
C5875 commonsourceibias.n162 gnd 0.058913f
C5876 commonsourceibias.n163 gnd 0.01085f
C5877 commonsourceibias.n164 gnd 0.009667f
C5878 commonsourceibias.n165 gnd 0.007903f
C5879 commonsourceibias.n166 gnd 0.007903f
C5880 commonsourceibias.n167 gnd 0.007903f
C5881 commonsourceibias.n168 gnd 0.009403f
C5882 commonsourceibias.n169 gnd 0.010904f
C5883 commonsourceibias.n170 gnd 0.058913f
C5884 commonsourceibias.n171 gnd 0.010838f
C5885 commonsourceibias.n172 gnd 0.007903f
C5886 commonsourceibias.n173 gnd 0.007903f
C5887 commonsourceibias.n174 gnd 0.007903f
C5888 commonsourceibias.n175 gnd 0.010705f
C5889 commonsourceibias.n176 gnd 0.058913f
C5890 commonsourceibias.n177 gnd 0.010776f
C5891 commonsourceibias.n178 gnd 0.009741f
C5892 commonsourceibias.n179 gnd 0.007903f
C5893 commonsourceibias.n180 gnd 0.007903f
C5894 commonsourceibias.n181 gnd 0.007903f
C5895 commonsourceibias.n182 gnd 0.008983f
C5896 commonsourceibias.n183 gnd 0.010937f
C5897 commonsourceibias.n184 gnd 0.058913f
C5898 commonsourceibias.n185 gnd 0.01089f
C5899 commonsourceibias.n186 gnd 0.007903f
C5900 commonsourceibias.n187 gnd 0.007903f
C5901 commonsourceibias.n188 gnd 0.007903f
C5902 commonsourceibias.n189 gnd 0.010623f
C5903 commonsourceibias.n190 gnd 0.058913f
C5904 commonsourceibias.n191 gnd 0.010649f
C5905 commonsourceibias.n192 gnd 0.071041f
C5906 commonsourceibias.n193 gnd 0.046914f
C5907 commonsourceibias.n194 gnd 0.010545f
C5908 commonsourceibias.t96 gnd 0.147652f
C5909 commonsourceibias.n195 gnd 0.006423f
C5910 commonsourceibias.n196 gnd 0.007903f
C5911 commonsourceibias.t65 gnd 0.147652f
C5912 commonsourceibias.n197 gnd 0.008017f
C5913 commonsourceibias.n198 gnd 0.007903f
C5914 commonsourceibias.t127 gnd 0.147652f
C5915 commonsourceibias.n199 gnd 0.058913f
C5916 commonsourceibias.t87 gnd 0.147652f
C5917 commonsourceibias.n200 gnd 0.006393f
C5918 commonsourceibias.n201 gnd 0.007903f
C5919 commonsourceibias.t104 gnd 0.147652f
C5920 commonsourceibias.n202 gnd 0.00763f
C5921 commonsourceibias.n203 gnd 0.007903f
C5922 commonsourceibias.t122 gnd 0.147652f
C5923 commonsourceibias.n204 gnd 0.058913f
C5924 commonsourceibias.t80 gnd 0.147652f
C5925 commonsourceibias.n205 gnd 0.006383f
C5926 commonsourceibias.n206 gnd 0.007903f
C5927 commonsourceibias.t76 gnd 0.147652f
C5928 commonsourceibias.t90 gnd 0.147652f
C5929 commonsourceibias.n207 gnd 0.058913f
C5930 commonsourceibias.n208 gnd 0.007903f
C5931 commonsourceibias.t74 gnd 0.147652f
C5932 commonsourceibias.n209 gnd 0.058913f
C5933 commonsourceibias.n210 gnd 0.007903f
C5934 commonsourceibias.t71 gnd 0.147652f
C5935 commonsourceibias.n211 gnd 0.058913f
C5936 commonsourceibias.n212 gnd 0.007903f
C5937 commonsourceibias.t83 gnd 0.147652f
C5938 commonsourceibias.n213 gnd 0.008983f
C5939 commonsourceibias.n214 gnd 0.007903f
C5940 commonsourceibias.t98 gnd 0.147652f
C5941 commonsourceibias.n215 gnd 0.010623f
C5942 commonsourceibias.t77 gnd 0.164481f
C5943 commonsourceibias.t67 gnd 0.147652f
C5944 commonsourceibias.n216 gnd 0.065644f
C5945 commonsourceibias.n217 gnd 0.070328f
C5946 commonsourceibias.n218 gnd 0.033639f
C5947 commonsourceibias.n219 gnd 0.007903f
C5948 commonsourceibias.n220 gnd 0.006423f
C5949 commonsourceibias.n221 gnd 0.01089f
C5950 commonsourceibias.n222 gnd 0.058913f
C5951 commonsourceibias.n223 gnd 0.010937f
C5952 commonsourceibias.n224 gnd 0.007903f
C5953 commonsourceibias.n225 gnd 0.007903f
C5954 commonsourceibias.n226 gnd 0.007903f
C5955 commonsourceibias.n227 gnd 0.008017f
C5956 commonsourceibias.n228 gnd 0.058913f
C5957 commonsourceibias.n229 gnd 0.009741f
C5958 commonsourceibias.n230 gnd 0.010776f
C5959 commonsourceibias.n231 gnd 0.007903f
C5960 commonsourceibias.n232 gnd 0.007903f
C5961 commonsourceibias.n233 gnd 0.010705f
C5962 commonsourceibias.n234 gnd 0.006393f
C5963 commonsourceibias.n235 gnd 0.010838f
C5964 commonsourceibias.n236 gnd 0.007903f
C5965 commonsourceibias.n237 gnd 0.007903f
C5966 commonsourceibias.n238 gnd 0.010904f
C5967 commonsourceibias.n239 gnd 0.009403f
C5968 commonsourceibias.n240 gnd 0.00763f
C5969 commonsourceibias.n241 gnd 0.007903f
C5970 commonsourceibias.n242 gnd 0.007903f
C5971 commonsourceibias.n243 gnd 0.009667f
C5972 commonsourceibias.n244 gnd 0.01085f
C5973 commonsourceibias.n245 gnd 0.058913f
C5974 commonsourceibias.n246 gnd 0.010777f
C5975 commonsourceibias.n247 gnd 0.007903f
C5976 commonsourceibias.n248 gnd 0.007903f
C5977 commonsourceibias.n249 gnd 0.007903f
C5978 commonsourceibias.n250 gnd 0.010777f
C5979 commonsourceibias.n251 gnd 0.058913f
C5980 commonsourceibias.n252 gnd 0.01085f
C5981 commonsourceibias.n253 gnd 0.009667f
C5982 commonsourceibias.n254 gnd 0.007903f
C5983 commonsourceibias.n255 gnd 0.007903f
C5984 commonsourceibias.n256 gnd 0.007903f
C5985 commonsourceibias.n257 gnd 0.009403f
C5986 commonsourceibias.n258 gnd 0.010904f
C5987 commonsourceibias.n259 gnd 0.058913f
C5988 commonsourceibias.n260 gnd 0.010838f
C5989 commonsourceibias.n261 gnd 0.007903f
C5990 commonsourceibias.n262 gnd 0.007903f
C5991 commonsourceibias.n263 gnd 0.007903f
C5992 commonsourceibias.n264 gnd 0.010705f
C5993 commonsourceibias.n265 gnd 0.058913f
C5994 commonsourceibias.n266 gnd 0.010776f
C5995 commonsourceibias.n267 gnd 0.009741f
C5996 commonsourceibias.n268 gnd 0.007903f
C5997 commonsourceibias.n269 gnd 0.007903f
C5998 commonsourceibias.n270 gnd 0.007903f
C5999 commonsourceibias.n271 gnd 0.008983f
C6000 commonsourceibias.n272 gnd 0.010937f
C6001 commonsourceibias.n273 gnd 0.058913f
C6002 commonsourceibias.n274 gnd 0.01089f
C6003 commonsourceibias.n275 gnd 0.007903f
C6004 commonsourceibias.n276 gnd 0.007903f
C6005 commonsourceibias.n277 gnd 0.007903f
C6006 commonsourceibias.n278 gnd 0.010623f
C6007 commonsourceibias.n279 gnd 0.058913f
C6008 commonsourceibias.n280 gnd 0.010649f
C6009 commonsourceibias.t81 gnd 0.159685f
C6010 commonsourceibias.n281 gnd 0.071041f
C6011 commonsourceibias.n282 gnd 0.02535f
C6012 commonsourceibias.n283 gnd 0.398385f
C6013 commonsourceibias.n284 gnd 0.010545f
C6014 commonsourceibias.t113 gnd 0.159685f
C6015 commonsourceibias.t123 gnd 0.147652f
C6016 commonsourceibias.n285 gnd 0.006423f
C6017 commonsourceibias.n286 gnd 0.007903f
C6018 commonsourceibias.t68 gnd 0.147652f
C6019 commonsourceibias.n287 gnd 0.008017f
C6020 commonsourceibias.n288 gnd 0.007903f
C6021 commonsourceibias.t119 gnd 0.147652f
C6022 commonsourceibias.n289 gnd 0.006393f
C6023 commonsourceibias.n290 gnd 0.007903f
C6024 commonsourceibias.t64 gnd 0.147652f
C6025 commonsourceibias.n291 gnd 0.00763f
C6026 commonsourceibias.n292 gnd 0.007903f
C6027 commonsourceibias.t112 gnd 0.147652f
C6028 commonsourceibias.n293 gnd 0.006383f
C6029 commonsourceibias.n294 gnd 0.007903f
C6030 commonsourceibias.t107 gnd 0.147652f
C6031 commonsourceibias.t121 gnd 0.147652f
C6032 commonsourceibias.n295 gnd 0.058913f
C6033 commonsourceibias.n296 gnd 0.007903f
C6034 commonsourceibias.t78 gnd 0.147652f
C6035 commonsourceibias.n297 gnd 0.058913f
C6036 commonsourceibias.n298 gnd 0.007903f
C6037 commonsourceibias.t101 gnd 0.147652f
C6038 commonsourceibias.n299 gnd 0.058913f
C6039 commonsourceibias.n300 gnd 0.007903f
C6040 commonsourceibias.t115 gnd 0.147652f
C6041 commonsourceibias.n301 gnd 0.008983f
C6042 commonsourceibias.n302 gnd 0.007903f
C6043 commonsourceibias.t125 gnd 0.147652f
C6044 commonsourceibias.n303 gnd 0.010623f
C6045 commonsourceibias.t108 gnd 0.164481f
C6046 commonsourceibias.t91 gnd 0.147652f
C6047 commonsourceibias.n304 gnd 0.065644f
C6048 commonsourceibias.n305 gnd 0.070328f
C6049 commonsourceibias.n306 gnd 0.033639f
C6050 commonsourceibias.n307 gnd 0.007903f
C6051 commonsourceibias.n308 gnd 0.006423f
C6052 commonsourceibias.n309 gnd 0.01089f
C6053 commonsourceibias.n310 gnd 0.058913f
C6054 commonsourceibias.n311 gnd 0.010937f
C6055 commonsourceibias.n312 gnd 0.007903f
C6056 commonsourceibias.n313 gnd 0.007903f
C6057 commonsourceibias.n314 gnd 0.007903f
C6058 commonsourceibias.n315 gnd 0.008017f
C6059 commonsourceibias.n316 gnd 0.058913f
C6060 commonsourceibias.n317 gnd 0.009741f
C6061 commonsourceibias.n318 gnd 0.010776f
C6062 commonsourceibias.n319 gnd 0.007903f
C6063 commonsourceibias.n320 gnd 0.007903f
C6064 commonsourceibias.n321 gnd 0.010705f
C6065 commonsourceibias.n322 gnd 0.006393f
C6066 commonsourceibias.n323 gnd 0.010838f
C6067 commonsourceibias.n324 gnd 0.007903f
C6068 commonsourceibias.n325 gnd 0.007903f
C6069 commonsourceibias.n326 gnd 0.010904f
C6070 commonsourceibias.n327 gnd 0.009403f
C6071 commonsourceibias.n328 gnd 0.00763f
C6072 commonsourceibias.n329 gnd 0.007903f
C6073 commonsourceibias.n330 gnd 0.007903f
C6074 commonsourceibias.n331 gnd 0.009667f
C6075 commonsourceibias.n332 gnd 0.01085f
C6076 commonsourceibias.n333 gnd 0.058913f
C6077 commonsourceibias.n334 gnd 0.010777f
C6078 commonsourceibias.n335 gnd 0.007865f
C6079 commonsourceibias.t5 gnd 0.017054f
C6080 commonsourceibias.t29 gnd 0.017054f
C6081 commonsourceibias.n336 gnd 0.151197f
C6082 commonsourceibias.t35 gnd 0.017054f
C6083 commonsourceibias.t13 gnd 0.017054f
C6084 commonsourceibias.n337 gnd 0.150693f
C6085 commonsourceibias.n338 gnd 0.140418f
C6086 commonsourceibias.t31 gnd 0.017054f
C6087 commonsourceibias.t37 gnd 0.017054f
C6088 commonsourceibias.n339 gnd 0.150693f
C6089 commonsourceibias.n340 gnd 0.069219f
C6090 commonsourceibias.t19 gnd 0.017054f
C6091 commonsourceibias.t47 gnd 0.017054f
C6092 commonsourceibias.n341 gnd 0.150693f
C6093 commonsourceibias.n342 gnd 0.057829f
C6094 commonsourceibias.n343 gnd 0.010545f
C6095 commonsourceibias.t22 gnd 0.147652f
C6096 commonsourceibias.n344 gnd 0.006423f
C6097 commonsourceibias.n345 gnd 0.007903f
C6098 commonsourceibias.t2 gnd 0.147652f
C6099 commonsourceibias.n346 gnd 0.008017f
C6100 commonsourceibias.n347 gnd 0.007903f
C6101 commonsourceibias.t50 gnd 0.147652f
C6102 commonsourceibias.n348 gnd 0.006393f
C6103 commonsourceibias.n349 gnd 0.007903f
C6104 commonsourceibias.t48 gnd 0.147652f
C6105 commonsourceibias.n350 gnd 0.00763f
C6106 commonsourceibias.n351 gnd 0.007903f
C6107 commonsourceibias.t8 gnd 0.147652f
C6108 commonsourceibias.n352 gnd 0.006383f
C6109 commonsourceibias.n353 gnd 0.007903f
C6110 commonsourceibias.t46 gnd 0.147652f
C6111 commonsourceibias.t18 gnd 0.147652f
C6112 commonsourceibias.n354 gnd 0.058913f
C6113 commonsourceibias.n355 gnd 0.007903f
C6114 commonsourceibias.t36 gnd 0.147652f
C6115 commonsourceibias.n356 gnd 0.058913f
C6116 commonsourceibias.n357 gnd 0.007903f
C6117 commonsourceibias.t30 gnd 0.147652f
C6118 commonsourceibias.n358 gnd 0.058913f
C6119 commonsourceibias.n359 gnd 0.007903f
C6120 commonsourceibias.t12 gnd 0.147652f
C6121 commonsourceibias.n360 gnd 0.008983f
C6122 commonsourceibias.n361 gnd 0.007903f
C6123 commonsourceibias.t34 gnd 0.147652f
C6124 commonsourceibias.n362 gnd 0.010623f
C6125 commonsourceibias.t4 gnd 0.164481f
C6126 commonsourceibias.t28 gnd 0.147652f
C6127 commonsourceibias.n363 gnd 0.065644f
C6128 commonsourceibias.n364 gnd 0.070328f
C6129 commonsourceibias.n365 gnd 0.033639f
C6130 commonsourceibias.n366 gnd 0.007903f
C6131 commonsourceibias.n367 gnd 0.006423f
C6132 commonsourceibias.n368 gnd 0.01089f
C6133 commonsourceibias.n369 gnd 0.058913f
C6134 commonsourceibias.n370 gnd 0.010937f
C6135 commonsourceibias.n371 gnd 0.007903f
C6136 commonsourceibias.n372 gnd 0.007903f
C6137 commonsourceibias.n373 gnd 0.007903f
C6138 commonsourceibias.n374 gnd 0.008017f
C6139 commonsourceibias.n375 gnd 0.058913f
C6140 commonsourceibias.n376 gnd 0.009741f
C6141 commonsourceibias.n377 gnd 0.010776f
C6142 commonsourceibias.n378 gnd 0.007903f
C6143 commonsourceibias.n379 gnd 0.007903f
C6144 commonsourceibias.n380 gnd 0.010705f
C6145 commonsourceibias.n381 gnd 0.006393f
C6146 commonsourceibias.n382 gnd 0.010838f
C6147 commonsourceibias.n383 gnd 0.007903f
C6148 commonsourceibias.n384 gnd 0.007903f
C6149 commonsourceibias.n385 gnd 0.010904f
C6150 commonsourceibias.n386 gnd 0.009403f
C6151 commonsourceibias.n387 gnd 0.00763f
C6152 commonsourceibias.n388 gnd 0.007903f
C6153 commonsourceibias.n389 gnd 0.007903f
C6154 commonsourceibias.n390 gnd 0.009667f
C6155 commonsourceibias.n391 gnd 0.01085f
C6156 commonsourceibias.n392 gnd 0.058913f
C6157 commonsourceibias.n393 gnd 0.010777f
C6158 commonsourceibias.n394 gnd 0.007903f
C6159 commonsourceibias.n395 gnd 0.007903f
C6160 commonsourceibias.n396 gnd 0.007903f
C6161 commonsourceibias.n397 gnd 0.010777f
C6162 commonsourceibias.n398 gnd 0.058913f
C6163 commonsourceibias.n399 gnd 0.01085f
C6164 commonsourceibias.t40 gnd 0.147652f
C6165 commonsourceibias.n400 gnd 0.058913f
C6166 commonsourceibias.n401 gnd 0.009667f
C6167 commonsourceibias.n402 gnd 0.007903f
C6168 commonsourceibias.n403 gnd 0.007903f
C6169 commonsourceibias.n404 gnd 0.007903f
C6170 commonsourceibias.n405 gnd 0.009403f
C6171 commonsourceibias.n406 gnd 0.010904f
C6172 commonsourceibias.n407 gnd 0.058913f
C6173 commonsourceibias.n408 gnd 0.010838f
C6174 commonsourceibias.n409 gnd 0.007903f
C6175 commonsourceibias.n410 gnd 0.007903f
C6176 commonsourceibias.n411 gnd 0.007903f
C6177 commonsourceibias.n412 gnd 0.010705f
C6178 commonsourceibias.n413 gnd 0.058913f
C6179 commonsourceibias.n414 gnd 0.010776f
C6180 commonsourceibias.t42 gnd 0.147652f
C6181 commonsourceibias.n415 gnd 0.058913f
C6182 commonsourceibias.n416 gnd 0.009741f
C6183 commonsourceibias.n417 gnd 0.007903f
C6184 commonsourceibias.n418 gnd 0.007903f
C6185 commonsourceibias.n419 gnd 0.007903f
C6186 commonsourceibias.n420 gnd 0.008983f
C6187 commonsourceibias.n421 gnd 0.010937f
C6188 commonsourceibias.n422 gnd 0.058913f
C6189 commonsourceibias.n423 gnd 0.01089f
C6190 commonsourceibias.n424 gnd 0.007903f
C6191 commonsourceibias.n425 gnd 0.007903f
C6192 commonsourceibias.n426 gnd 0.007903f
C6193 commonsourceibias.n427 gnd 0.010623f
C6194 commonsourceibias.n428 gnd 0.058913f
C6195 commonsourceibias.n429 gnd 0.010649f
C6196 commonsourceibias.t44 gnd 0.159685f
C6197 commonsourceibias.n430 gnd 0.071041f
C6198 commonsourceibias.n431 gnd 0.079434f
C6199 commonsourceibias.t23 gnd 0.017054f
C6200 commonsourceibias.t45 gnd 0.017054f
C6201 commonsourceibias.n432 gnd 0.150693f
C6202 commonsourceibias.n433 gnd 0.130533f
C6203 commonsourceibias.t43 gnd 0.017054f
C6204 commonsourceibias.t3 gnd 0.017054f
C6205 commonsourceibias.n434 gnd 0.150693f
C6206 commonsourceibias.n435 gnd 0.069219f
C6207 commonsourceibias.t49 gnd 0.017054f
C6208 commonsourceibias.t51 gnd 0.017054f
C6209 commonsourceibias.n436 gnd 0.150693f
C6210 commonsourceibias.n437 gnd 0.069219f
C6211 commonsourceibias.t9 gnd 0.017054f
C6212 commonsourceibias.t41 gnd 0.017054f
C6213 commonsourceibias.n438 gnd 0.150693f
C6214 commonsourceibias.n439 gnd 0.057829f
C6215 commonsourceibias.n440 gnd 0.070025f
C6216 commonsourceibias.n441 gnd 0.057129f
C6217 commonsourceibias.n442 gnd 0.007865f
C6218 commonsourceibias.n443 gnd 0.010777f
C6219 commonsourceibias.n444 gnd 0.058913f
C6220 commonsourceibias.n445 gnd 0.01085f
C6221 commonsourceibias.t126 gnd 0.147652f
C6222 commonsourceibias.n446 gnd 0.058913f
C6223 commonsourceibias.n447 gnd 0.009667f
C6224 commonsourceibias.n448 gnd 0.007903f
C6225 commonsourceibias.n449 gnd 0.007903f
C6226 commonsourceibias.n450 gnd 0.007903f
C6227 commonsourceibias.n451 gnd 0.009403f
C6228 commonsourceibias.n452 gnd 0.010904f
C6229 commonsourceibias.n453 gnd 0.058913f
C6230 commonsourceibias.n454 gnd 0.010838f
C6231 commonsourceibias.n455 gnd 0.007903f
C6232 commonsourceibias.n456 gnd 0.007903f
C6233 commonsourceibias.n457 gnd 0.007903f
C6234 commonsourceibias.n458 gnd 0.010705f
C6235 commonsourceibias.n459 gnd 0.058913f
C6236 commonsourceibias.n460 gnd 0.010776f
C6237 commonsourceibias.t84 gnd 0.147652f
C6238 commonsourceibias.n461 gnd 0.058913f
C6239 commonsourceibias.n462 gnd 0.009741f
C6240 commonsourceibias.n463 gnd 0.007903f
C6241 commonsourceibias.n464 gnd 0.007903f
C6242 commonsourceibias.n465 gnd 0.007903f
C6243 commonsourceibias.n466 gnd 0.008983f
C6244 commonsourceibias.n467 gnd 0.010937f
C6245 commonsourceibias.n468 gnd 0.058913f
C6246 commonsourceibias.n469 gnd 0.01089f
C6247 commonsourceibias.n470 gnd 0.007903f
C6248 commonsourceibias.n471 gnd 0.007903f
C6249 commonsourceibias.n472 gnd 0.007903f
C6250 commonsourceibias.n473 gnd 0.010623f
C6251 commonsourceibias.n474 gnd 0.058913f
C6252 commonsourceibias.n475 gnd 0.010649f
C6253 commonsourceibias.n476 gnd 0.071041f
C6254 commonsourceibias.n477 gnd 0.046914f
C6255 commonsourceibias.n478 gnd 0.010545f
C6256 commonsourceibias.t114 gnd 0.147652f
C6257 commonsourceibias.n479 gnd 0.006423f
C6258 commonsourceibias.n480 gnd 0.007903f
C6259 commonsourceibias.t124 gnd 0.147652f
C6260 commonsourceibias.n481 gnd 0.008017f
C6261 commonsourceibias.n482 gnd 0.007903f
C6262 commonsourceibias.t106 gnd 0.147652f
C6263 commonsourceibias.n483 gnd 0.006393f
C6264 commonsourceibias.n484 gnd 0.007903f
C6265 commonsourceibias.t120 gnd 0.147652f
C6266 commonsourceibias.n485 gnd 0.00763f
C6267 commonsourceibias.n486 gnd 0.007903f
C6268 commonsourceibias.t99 gnd 0.147652f
C6269 commonsourceibias.n487 gnd 0.006383f
C6270 commonsourceibias.n488 gnd 0.007903f
C6271 commonsourceibias.t92 gnd 0.147652f
C6272 commonsourceibias.t110 gnd 0.147652f
C6273 commonsourceibias.n489 gnd 0.058913f
C6274 commonsourceibias.n490 gnd 0.007903f
C6275 commonsourceibias.t69 gnd 0.147652f
C6276 commonsourceibias.n491 gnd 0.058913f
C6277 commonsourceibias.n492 gnd 0.007903f
C6278 commonsourceibias.t85 gnd 0.147652f
C6279 commonsourceibias.n493 gnd 0.058913f
C6280 commonsourceibias.n494 gnd 0.007903f
C6281 commonsourceibias.t103 gnd 0.147652f
C6282 commonsourceibias.n495 gnd 0.008983f
C6283 commonsourceibias.n496 gnd 0.007903f
C6284 commonsourceibias.t116 gnd 0.147652f
C6285 commonsourceibias.n497 gnd 0.010623f
C6286 commonsourceibias.t95 gnd 0.164481f
C6287 commonsourceibias.t79 gnd 0.147652f
C6288 commonsourceibias.n498 gnd 0.065644f
C6289 commonsourceibias.n499 gnd 0.070328f
C6290 commonsourceibias.n500 gnd 0.033639f
C6291 commonsourceibias.n501 gnd 0.007903f
C6292 commonsourceibias.n502 gnd 0.006423f
C6293 commonsourceibias.n503 gnd 0.01089f
C6294 commonsourceibias.n504 gnd 0.058913f
C6295 commonsourceibias.n505 gnd 0.010937f
C6296 commonsourceibias.n506 gnd 0.007903f
C6297 commonsourceibias.n507 gnd 0.007903f
C6298 commonsourceibias.n508 gnd 0.007903f
C6299 commonsourceibias.n509 gnd 0.008017f
C6300 commonsourceibias.n510 gnd 0.058913f
C6301 commonsourceibias.n511 gnd 0.009741f
C6302 commonsourceibias.n512 gnd 0.010776f
C6303 commonsourceibias.n513 gnd 0.007903f
C6304 commonsourceibias.n514 gnd 0.007903f
C6305 commonsourceibias.n515 gnd 0.010705f
C6306 commonsourceibias.n516 gnd 0.006393f
C6307 commonsourceibias.n517 gnd 0.010838f
C6308 commonsourceibias.n518 gnd 0.007903f
C6309 commonsourceibias.n519 gnd 0.007903f
C6310 commonsourceibias.n520 gnd 0.010904f
C6311 commonsourceibias.n521 gnd 0.009403f
C6312 commonsourceibias.n522 gnd 0.00763f
C6313 commonsourceibias.n523 gnd 0.007903f
C6314 commonsourceibias.n524 gnd 0.007903f
C6315 commonsourceibias.n525 gnd 0.009667f
C6316 commonsourceibias.n526 gnd 0.01085f
C6317 commonsourceibias.n527 gnd 0.058913f
C6318 commonsourceibias.n528 gnd 0.010777f
C6319 commonsourceibias.n529 gnd 0.007903f
C6320 commonsourceibias.n530 gnd 0.007903f
C6321 commonsourceibias.n531 gnd 0.007903f
C6322 commonsourceibias.n532 gnd 0.010777f
C6323 commonsourceibias.n533 gnd 0.058913f
C6324 commonsourceibias.n534 gnd 0.01085f
C6325 commonsourceibias.t117 gnd 0.147652f
C6326 commonsourceibias.n535 gnd 0.058913f
C6327 commonsourceibias.n536 gnd 0.009667f
C6328 commonsourceibias.n537 gnd 0.007903f
C6329 commonsourceibias.n538 gnd 0.007903f
C6330 commonsourceibias.n539 gnd 0.007903f
C6331 commonsourceibias.n540 gnd 0.009403f
C6332 commonsourceibias.n541 gnd 0.010904f
C6333 commonsourceibias.n542 gnd 0.058913f
C6334 commonsourceibias.n543 gnd 0.010838f
C6335 commonsourceibias.n544 gnd 0.007903f
C6336 commonsourceibias.n545 gnd 0.007903f
C6337 commonsourceibias.n546 gnd 0.007903f
C6338 commonsourceibias.n547 gnd 0.010705f
C6339 commonsourceibias.n548 gnd 0.058913f
C6340 commonsourceibias.n549 gnd 0.010776f
C6341 commonsourceibias.t73 gnd 0.147652f
C6342 commonsourceibias.n550 gnd 0.058913f
C6343 commonsourceibias.n551 gnd 0.009741f
C6344 commonsourceibias.n552 gnd 0.007903f
C6345 commonsourceibias.n553 gnd 0.007903f
C6346 commonsourceibias.n554 gnd 0.007903f
C6347 commonsourceibias.n555 gnd 0.008983f
C6348 commonsourceibias.n556 gnd 0.010937f
C6349 commonsourceibias.n557 gnd 0.058913f
C6350 commonsourceibias.n558 gnd 0.01089f
C6351 commonsourceibias.n559 gnd 0.007903f
C6352 commonsourceibias.n560 gnd 0.007903f
C6353 commonsourceibias.n561 gnd 0.007903f
C6354 commonsourceibias.n562 gnd 0.010623f
C6355 commonsourceibias.n563 gnd 0.058913f
C6356 commonsourceibias.n564 gnd 0.010649f
C6357 commonsourceibias.t100 gnd 0.159685f
C6358 commonsourceibias.n565 gnd 0.071041f
C6359 commonsourceibias.n566 gnd 0.02535f
C6360 commonsourceibias.n567 gnd 0.218509f
C6361 commonsourceibias.n568 gnd 4.2686f
.ends

