* NGSPICE file created from diffpair.ext - technology: sky130A

.subckt diffpair minus drain_right drain_left source plus
X0 source.t47 plus.t0 drain_left.t21 a_n4174_n2688# sky130_fd_pr__nfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=1
X1 source.t22 minus.t0 drain_right.t23 a_n4174_n2688# sky130_fd_pr__nfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=1
X2 drain_right.t22 minus.t1 source.t6 a_n4174_n2688# sky130_fd_pr__nfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=1
X3 source.t8 minus.t2 drain_right.t21 a_n4174_n2688# sky130_fd_pr__nfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=1
X4 source.t46 plus.t1 drain_left.t23 a_n4174_n2688# sky130_fd_pr__nfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=1
X5 drain_left.t9 plus.t2 source.t45 a_n4174_n2688# sky130_fd_pr__nfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=1
X6 source.t1 minus.t3 drain_right.t20 a_n4174_n2688# sky130_fd_pr__nfet_01v8 ad=3.51 pd=18.78 as=1.485 ps=9.33 w=9 l=1
X7 source.t2 minus.t4 drain_right.t19 a_n4174_n2688# sky130_fd_pr__nfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=1
X8 drain_left.t1 plus.t3 source.t44 a_n4174_n2688# sky130_fd_pr__nfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=1
X9 drain_right.t18 minus.t5 source.t15 a_n4174_n2688# sky130_fd_pr__nfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=1
X10 source.t11 minus.t6 drain_right.t17 a_n4174_n2688# sky130_fd_pr__nfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=1
X11 drain_left.t7 plus.t4 source.t43 a_n4174_n2688# sky130_fd_pr__nfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=1
X12 drain_left.t18 plus.t5 source.t42 a_n4174_n2688# sky130_fd_pr__nfet_01v8 ad=1.485 pd=9.33 as=3.51 ps=18.78 w=9 l=1
X13 source.t41 plus.t6 drain_left.t16 a_n4174_n2688# sky130_fd_pr__nfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=1
X14 a_n4174_n2688# a_n4174_n2688# a_n4174_n2688# a_n4174_n2688# sky130_fd_pr__nfet_01v8 ad=3.51 pd=18.78 as=28.08 ps=150.24 w=9 l=1
X15 drain_right.t16 minus.t7 source.t9 a_n4174_n2688# sky130_fd_pr__nfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=1
X16 source.t4 minus.t8 drain_right.t15 a_n4174_n2688# sky130_fd_pr__nfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=1
X17 source.t40 plus.t7 drain_left.t4 a_n4174_n2688# sky130_fd_pr__nfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=1
X18 source.t39 plus.t8 drain_left.t20 a_n4174_n2688# sky130_fd_pr__nfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=1
X19 drain_left.t17 plus.t9 source.t38 a_n4174_n2688# sky130_fd_pr__nfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=1
X20 source.t37 plus.t10 drain_left.t6 a_n4174_n2688# sky130_fd_pr__nfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=1
X21 drain_left.t3 plus.t11 source.t36 a_n4174_n2688# sky130_fd_pr__nfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=1
X22 drain_right.t14 minus.t9 source.t16 a_n4174_n2688# sky130_fd_pr__nfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=1
X23 drain_left.t2 plus.t12 source.t35 a_n4174_n2688# sky130_fd_pr__nfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=1
X24 drain_left.t19 plus.t13 source.t34 a_n4174_n2688# sky130_fd_pr__nfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=1
X25 source.t33 plus.t14 drain_left.t11 a_n4174_n2688# sky130_fd_pr__nfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=1
X26 source.t32 plus.t15 drain_left.t12 a_n4174_n2688# sky130_fd_pr__nfet_01v8 ad=3.51 pd=18.78 as=1.485 ps=9.33 w=9 l=1
X27 drain_right.t13 minus.t10 source.t7 a_n4174_n2688# sky130_fd_pr__nfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=1
X28 drain_left.t10 plus.t16 source.t31 a_n4174_n2688# sky130_fd_pr__nfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=1
X29 drain_right.t12 minus.t11 source.t14 a_n4174_n2688# sky130_fd_pr__nfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=1
X30 source.t3 minus.t12 drain_right.t11 a_n4174_n2688# sky130_fd_pr__nfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=1
X31 source.t30 plus.t17 drain_left.t5 a_n4174_n2688# sky130_fd_pr__nfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=1
X32 source.t29 plus.t18 drain_left.t14 a_n4174_n2688# sky130_fd_pr__nfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=1
X33 source.t28 plus.t19 drain_left.t15 a_n4174_n2688# sky130_fd_pr__nfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=1
X34 drain_right.t10 minus.t13 source.t10 a_n4174_n2688# sky130_fd_pr__nfet_01v8 ad=1.485 pd=9.33 as=3.51 ps=18.78 w=9 l=1
X35 drain_right.t9 minus.t14 source.t13 a_n4174_n2688# sky130_fd_pr__nfet_01v8 ad=1.485 pd=9.33 as=3.51 ps=18.78 w=9 l=1
X36 drain_left.t13 plus.t20 source.t27 a_n4174_n2688# sky130_fd_pr__nfet_01v8 ad=1.485 pd=9.33 as=3.51 ps=18.78 w=9 l=1
X37 drain_right.t8 minus.t15 source.t18 a_n4174_n2688# sky130_fd_pr__nfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=1
X38 drain_right.t7 minus.t16 source.t0 a_n4174_n2688# sky130_fd_pr__nfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=1
X39 a_n4174_n2688# a_n4174_n2688# a_n4174_n2688# a_n4174_n2688# sky130_fd_pr__nfet_01v8 ad=3.51 pd=18.78 as=0 ps=0 w=9 l=1
X40 source.t5 minus.t17 drain_right.t6 a_n4174_n2688# sky130_fd_pr__nfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=1
X41 source.t17 minus.t18 drain_right.t5 a_n4174_n2688# sky130_fd_pr__nfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=1
X42 source.t12 minus.t19 drain_right.t4 a_n4174_n2688# sky130_fd_pr__nfet_01v8 ad=3.51 pd=18.78 as=1.485 ps=9.33 w=9 l=1
X43 source.t21 minus.t20 drain_right.t3 a_n4174_n2688# sky130_fd_pr__nfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=1
X44 source.t20 minus.t21 drain_right.t2 a_n4174_n2688# sky130_fd_pr__nfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=1
X45 drain_right.t1 minus.t22 source.t19 a_n4174_n2688# sky130_fd_pr__nfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=1
X46 a_n4174_n2688# a_n4174_n2688# a_n4174_n2688# a_n4174_n2688# sky130_fd_pr__nfet_01v8 ad=3.51 pd=18.78 as=0 ps=0 w=9 l=1
X47 source.t26 plus.t21 drain_left.t22 a_n4174_n2688# sky130_fd_pr__nfet_01v8 ad=3.51 pd=18.78 as=1.485 ps=9.33 w=9 l=1
X48 drain_right.t0 minus.t23 source.t23 a_n4174_n2688# sky130_fd_pr__nfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=1
X49 drain_left.t8 plus.t22 source.t25 a_n4174_n2688# sky130_fd_pr__nfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=1
X50 drain_left.t0 plus.t23 source.t24 a_n4174_n2688# sky130_fd_pr__nfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=1
X51 a_n4174_n2688# a_n4174_n2688# a_n4174_n2688# a_n4174_n2688# sky130_fd_pr__nfet_01v8 ad=3.51 pd=18.78 as=0 ps=0 w=9 l=1
R0 plus.n15 plus.t21 278.204
R1 plus.n79 plus.t20 278.204
R2 plus.n61 plus.t5 256.183
R3 plus.n124 plus.t15 256.183
R4 plus.n1 plus.t8 216.9
R5 plus.n54 plus.t13 216.9
R6 plus.n48 plus.t6 216.9
R7 plus.n41 plus.t9 216.9
R8 plus.n39 plus.t14 216.9
R9 plus.n33 plus.t4 216.9
R10 plus.n9 plus.t10 216.9
R11 plus.n11 plus.t3 216.9
R12 plus.n13 plus.t0 216.9
R13 plus.n16 plus.t2 216.9
R14 plus.n64 plus.t23 216.9
R15 plus.n117 plus.t7 216.9
R16 plus.n111 plus.t12 216.9
R17 plus.n70 plus.t1 216.9
R18 plus.n103 plus.t16 216.9
R19 plus.n97 plus.t19 216.9
R20 plus.n73 plus.t11 216.9
R21 plus.n75 plus.t17 216.9
R22 plus.n77 plus.t22 216.9
R23 plus.n80 plus.t18 216.9
R24 plus.n17 plus.n14 161.3
R25 plus.n19 plus.n18 161.3
R26 plus.n21 plus.n20 161.3
R27 plus.n22 plus.n12 161.3
R28 plus.n24 plus.n23 161.3
R29 plus.n26 plus.n25 161.3
R30 plus.n27 plus.n10 161.3
R31 plus.n29 plus.n28 161.3
R32 plus.n31 plus.n30 161.3
R33 plus.n32 plus.n8 161.3
R34 plus.n35 plus.n34 161.3
R35 plus.n36 plus.n7 161.3
R36 plus.n38 plus.n37 161.3
R37 plus.n40 plus.n6 161.3
R38 plus.n43 plus.n42 161.3
R39 plus.n44 plus.n5 161.3
R40 plus.n46 plus.n45 161.3
R41 plus.n47 plus.n4 161.3
R42 plus.n50 plus.n49 161.3
R43 plus.n51 plus.n3 161.3
R44 plus.n53 plus.n52 161.3
R45 plus.n55 plus.n2 161.3
R46 plus.n57 plus.n56 161.3
R47 plus.n59 plus.n58 161.3
R48 plus.n60 plus.n0 161.3
R49 plus.n81 plus.n78 161.3
R50 plus.n83 plus.n82 161.3
R51 plus.n85 plus.n84 161.3
R52 plus.n86 plus.n76 161.3
R53 plus.n88 plus.n87 161.3
R54 plus.n90 plus.n89 161.3
R55 plus.n91 plus.n74 161.3
R56 plus.n93 plus.n92 161.3
R57 plus.n95 plus.n94 161.3
R58 plus.n96 plus.n72 161.3
R59 plus.n99 plus.n98 161.3
R60 plus.n100 plus.n71 161.3
R61 plus.n102 plus.n101 161.3
R62 plus.n104 plus.n69 161.3
R63 plus.n106 plus.n105 161.3
R64 plus.n107 plus.n68 161.3
R65 plus.n109 plus.n108 161.3
R66 plus.n110 plus.n67 161.3
R67 plus.n113 plus.n112 161.3
R68 plus.n114 plus.n66 161.3
R69 plus.n116 plus.n115 161.3
R70 plus.n118 plus.n65 161.3
R71 plus.n120 plus.n119 161.3
R72 plus.n122 plus.n121 161.3
R73 plus.n123 plus.n63 161.3
R74 plus.n62 plus.n61 80.6037
R75 plus.n125 plus.n124 80.6037
R76 plus.n56 plus.n55 56.5617
R77 plus.n42 plus.n40 56.5617
R78 plus.n32 plus.n31 56.5617
R79 plus.n18 plus.n17 56.5617
R80 plus.n119 plus.n118 56.5617
R81 plus.n105 plus.n104 56.5617
R82 plus.n96 plus.n95 56.5617
R83 plus.n82 plus.n81 56.5617
R84 plus.n47 plus.n46 56.0773
R85 plus.n27 plus.n26 56.0773
R86 plus.n110 plus.n109 56.0773
R87 plus.n91 plus.n90 56.0773
R88 plus.n61 plus.n60 46.0096
R89 plus.n124 plus.n123 46.0096
R90 plus.n49 plus.n3 41.5458
R91 plus.n23 plus.n22 41.5458
R92 plus.n112 plus.n66 41.5458
R93 plus.n87 plus.n86 41.5458
R94 plus.n38 plus.n7 40.577
R95 plus.n34 plus.n7 40.577
R96 plus.n102 plus.n71 40.577
R97 plus.n98 plus.n71 40.577
R98 plus.n53 plus.n3 39.6083
R99 plus.n22 plus.n21 39.6083
R100 plus.n116 plus.n66 39.6083
R101 plus.n86 plus.n85 39.6083
R102 plus plus.n125 37.9881
R103 plus.n16 plus.n15 33.0515
R104 plus.n80 plus.n79 33.0515
R105 plus.n15 plus.n14 28.5514
R106 plus.n79 plus.n78 28.5514
R107 plus.n60 plus.n59 26.0455
R108 plus.n123 plus.n122 26.0455
R109 plus.n46 plus.n5 25.0767
R110 plus.n28 plus.n27 25.0767
R111 plus.n109 plus.n68 25.0767
R112 plus.n92 plus.n91 25.0767
R113 plus.n42 plus.n41 24.3464
R114 plus.n31 plus.n9 24.3464
R115 plus.n105 plus.n70 24.3464
R116 plus.n95 plus.n73 24.3464
R117 plus.n56 plus.n1 23.8546
R118 plus.n17 plus.n16 23.8546
R119 plus.n119 plus.n64 23.8546
R120 plus.n81 plus.n80 23.8546
R121 plus.n55 plus.n54 16.9689
R122 plus.n18 plus.n13 16.9689
R123 plus.n118 plus.n117 16.9689
R124 plus.n82 plus.n77 16.9689
R125 plus.n40 plus.n39 16.477
R126 plus.n33 plus.n32 16.477
R127 plus.n104 plus.n103 16.477
R128 plus.n97 plus.n96 16.477
R129 plus.n48 plus.n47 15.9852
R130 plus.n26 plus.n11 15.9852
R131 plus.n111 plus.n110 15.9852
R132 plus.n90 plus.n75 15.9852
R133 plus plus.n62 11.3191
R134 plus.n49 plus.n48 8.60764
R135 plus.n23 plus.n11 8.60764
R136 plus.n112 plus.n111 8.60764
R137 plus.n87 plus.n75 8.60764
R138 plus.n39 plus.n38 8.11581
R139 plus.n34 plus.n33 8.11581
R140 plus.n103 plus.n102 8.11581
R141 plus.n98 plus.n97 8.11581
R142 plus.n54 plus.n53 7.62397
R143 plus.n21 plus.n13 7.62397
R144 plus.n117 plus.n116 7.62397
R145 plus.n85 plus.n77 7.62397
R146 plus.n59 plus.n1 0.738255
R147 plus.n122 plus.n64 0.738255
R148 plus.n62 plus.n0 0.285035
R149 plus.n125 plus.n63 0.285035
R150 plus.n41 plus.n5 0.246418
R151 plus.n28 plus.n9 0.246418
R152 plus.n70 plus.n68 0.246418
R153 plus.n92 plus.n73 0.246418
R154 plus.n19 plus.n14 0.189894
R155 plus.n20 plus.n19 0.189894
R156 plus.n20 plus.n12 0.189894
R157 plus.n24 plus.n12 0.189894
R158 plus.n25 plus.n24 0.189894
R159 plus.n25 plus.n10 0.189894
R160 plus.n29 plus.n10 0.189894
R161 plus.n30 plus.n29 0.189894
R162 plus.n30 plus.n8 0.189894
R163 plus.n35 plus.n8 0.189894
R164 plus.n36 plus.n35 0.189894
R165 plus.n37 plus.n36 0.189894
R166 plus.n37 plus.n6 0.189894
R167 plus.n43 plus.n6 0.189894
R168 plus.n44 plus.n43 0.189894
R169 plus.n45 plus.n44 0.189894
R170 plus.n45 plus.n4 0.189894
R171 plus.n50 plus.n4 0.189894
R172 plus.n51 plus.n50 0.189894
R173 plus.n52 plus.n51 0.189894
R174 plus.n52 plus.n2 0.189894
R175 plus.n57 plus.n2 0.189894
R176 plus.n58 plus.n57 0.189894
R177 plus.n58 plus.n0 0.189894
R178 plus.n121 plus.n63 0.189894
R179 plus.n121 plus.n120 0.189894
R180 plus.n120 plus.n65 0.189894
R181 plus.n115 plus.n65 0.189894
R182 plus.n115 plus.n114 0.189894
R183 plus.n114 plus.n113 0.189894
R184 plus.n113 plus.n67 0.189894
R185 plus.n108 plus.n67 0.189894
R186 plus.n108 plus.n107 0.189894
R187 plus.n107 plus.n106 0.189894
R188 plus.n106 plus.n69 0.189894
R189 plus.n101 plus.n69 0.189894
R190 plus.n101 plus.n100 0.189894
R191 plus.n100 plus.n99 0.189894
R192 plus.n99 plus.n72 0.189894
R193 plus.n94 plus.n72 0.189894
R194 plus.n94 plus.n93 0.189894
R195 plus.n93 plus.n74 0.189894
R196 plus.n89 plus.n74 0.189894
R197 plus.n89 plus.n88 0.189894
R198 plus.n88 plus.n76 0.189894
R199 plus.n84 plus.n76 0.189894
R200 plus.n84 plus.n83 0.189894
R201 plus.n83 plus.n78 0.189894
R202 drain_left.n13 drain_left.n11 66.6841
R203 drain_left.n7 drain_left.n5 66.6839
R204 drain_left.n2 drain_left.n0 66.6839
R205 drain_left.n19 drain_left.n18 65.5376
R206 drain_left.n17 drain_left.n16 65.5376
R207 drain_left.n15 drain_left.n14 65.5376
R208 drain_left.n13 drain_left.n12 65.5376
R209 drain_left.n21 drain_left.n20 65.5374
R210 drain_left.n7 drain_left.n6 65.5373
R211 drain_left.n9 drain_left.n8 65.5373
R212 drain_left.n4 drain_left.n3 65.5373
R213 drain_left.n2 drain_left.n1 65.5373
R214 drain_left drain_left.n10 35.9866
R215 drain_left drain_left.n21 6.79977
R216 drain_left.n5 drain_left.t14 2.2005
R217 drain_left.n5 drain_left.t13 2.2005
R218 drain_left.n6 drain_left.t5 2.2005
R219 drain_left.n6 drain_left.t8 2.2005
R220 drain_left.n8 drain_left.t15 2.2005
R221 drain_left.n8 drain_left.t3 2.2005
R222 drain_left.n3 drain_left.t23 2.2005
R223 drain_left.n3 drain_left.t10 2.2005
R224 drain_left.n1 drain_left.t4 2.2005
R225 drain_left.n1 drain_left.t2 2.2005
R226 drain_left.n0 drain_left.t12 2.2005
R227 drain_left.n0 drain_left.t0 2.2005
R228 drain_left.n20 drain_left.t20 2.2005
R229 drain_left.n20 drain_left.t18 2.2005
R230 drain_left.n18 drain_left.t16 2.2005
R231 drain_left.n18 drain_left.t19 2.2005
R232 drain_left.n16 drain_left.t11 2.2005
R233 drain_left.n16 drain_left.t17 2.2005
R234 drain_left.n14 drain_left.t6 2.2005
R235 drain_left.n14 drain_left.t7 2.2005
R236 drain_left.n12 drain_left.t21 2.2005
R237 drain_left.n12 drain_left.t1 2.2005
R238 drain_left.n11 drain_left.t22 2.2005
R239 drain_left.n11 drain_left.t9 2.2005
R240 drain_left.n9 drain_left.n7 1.14705
R241 drain_left.n4 drain_left.n2 1.14705
R242 drain_left.n15 drain_left.n13 1.14705
R243 drain_left.n17 drain_left.n15 1.14705
R244 drain_left.n19 drain_left.n17 1.14705
R245 drain_left.n21 drain_left.n19 1.14705
R246 drain_left.n10 drain_left.n9 0.51843
R247 drain_left.n10 drain_left.n4 0.51843
R248 source.n11 source.t26 51.0588
R249 source.n12 source.t10 51.0588
R250 source.n23 source.t1 51.0588
R251 source.n47 source.t13 51.0586
R252 source.n36 source.t12 51.0586
R253 source.n35 source.t27 51.0586
R254 source.n24 source.t32 51.0586
R255 source.n0 source.t42 51.0586
R256 source.n2 source.n1 48.8588
R257 source.n4 source.n3 48.8588
R258 source.n6 source.n5 48.8588
R259 source.n8 source.n7 48.8588
R260 source.n10 source.n9 48.8588
R261 source.n14 source.n13 48.8588
R262 source.n16 source.n15 48.8588
R263 source.n18 source.n17 48.8588
R264 source.n20 source.n19 48.8588
R265 source.n22 source.n21 48.8588
R266 source.n46 source.n45 48.8586
R267 source.n44 source.n43 48.8586
R268 source.n42 source.n41 48.8586
R269 source.n40 source.n39 48.8586
R270 source.n38 source.n37 48.8586
R271 source.n34 source.n33 48.8586
R272 source.n32 source.n31 48.8586
R273 source.n30 source.n29 48.8586
R274 source.n28 source.n27 48.8586
R275 source.n26 source.n25 48.8586
R276 source.n24 source.n23 20.1616
R277 source.n48 source.n0 14.3253
R278 source.n48 source.n47 5.83671
R279 source.n45 source.t14 2.2005
R280 source.n45 source.t2 2.2005
R281 source.n43 source.t16 2.2005
R282 source.n43 source.t20 2.2005
R283 source.n41 source.t19 2.2005
R284 source.n41 source.t5 2.2005
R285 source.n39 source.t23 2.2005
R286 source.n39 source.t3 2.2005
R287 source.n37 source.t0 2.2005
R288 source.n37 source.t8 2.2005
R289 source.n33 source.t25 2.2005
R290 source.n33 source.t29 2.2005
R291 source.n31 source.t36 2.2005
R292 source.n31 source.t30 2.2005
R293 source.n29 source.t31 2.2005
R294 source.n29 source.t28 2.2005
R295 source.n27 source.t35 2.2005
R296 source.n27 source.t46 2.2005
R297 source.n25 source.t24 2.2005
R298 source.n25 source.t40 2.2005
R299 source.n1 source.t34 2.2005
R300 source.n1 source.t39 2.2005
R301 source.n3 source.t38 2.2005
R302 source.n3 source.t41 2.2005
R303 source.n5 source.t43 2.2005
R304 source.n5 source.t33 2.2005
R305 source.n7 source.t44 2.2005
R306 source.n7 source.t37 2.2005
R307 source.n9 source.t45 2.2005
R308 source.n9 source.t47 2.2005
R309 source.n13 source.t18 2.2005
R310 source.n13 source.t17 2.2005
R311 source.n15 source.t15 2.2005
R312 source.n15 source.t21 2.2005
R313 source.n17 source.t9 2.2005
R314 source.n17 source.t22 2.2005
R315 source.n19 source.t6 2.2005
R316 source.n19 source.t11 2.2005
R317 source.n21 source.t7 2.2005
R318 source.n21 source.t4 2.2005
R319 source.n23 source.n22 1.14705
R320 source.n22 source.n20 1.14705
R321 source.n20 source.n18 1.14705
R322 source.n18 source.n16 1.14705
R323 source.n16 source.n14 1.14705
R324 source.n14 source.n12 1.14705
R325 source.n11 source.n10 1.14705
R326 source.n10 source.n8 1.14705
R327 source.n8 source.n6 1.14705
R328 source.n6 source.n4 1.14705
R329 source.n4 source.n2 1.14705
R330 source.n2 source.n0 1.14705
R331 source.n26 source.n24 1.14705
R332 source.n28 source.n26 1.14705
R333 source.n30 source.n28 1.14705
R334 source.n32 source.n30 1.14705
R335 source.n34 source.n32 1.14705
R336 source.n35 source.n34 1.14705
R337 source.n38 source.n36 1.14705
R338 source.n40 source.n38 1.14705
R339 source.n42 source.n40 1.14705
R340 source.n44 source.n42 1.14705
R341 source.n46 source.n44 1.14705
R342 source.n47 source.n46 1.14705
R343 source.n12 source.n11 0.470328
R344 source.n36 source.n35 0.470328
R345 source source.n48 0.188
R346 minus.n16 minus.t13 278.204
R347 minus.n78 minus.t19 278.204
R348 minus.n61 minus.t3 256.183
R349 minus.n124 minus.t14 256.183
R350 minus.n17 minus.t18 216.9
R351 minus.n14 minus.t15 216.9
R352 minus.n12 minus.t20 216.9
R353 minus.n10 minus.t5 216.9
R354 minus.n34 minus.t0 216.9
R355 minus.n40 minus.t7 216.9
R356 minus.n7 minus.t6 216.9
R357 minus.n48 minus.t1 216.9
R358 minus.n54 minus.t8 216.9
R359 minus.n1 minus.t10 216.9
R360 minus.n79 minus.t16 216.9
R361 minus.n76 minus.t2 216.9
R362 minus.n74 minus.t23 216.9
R363 minus.n72 minus.t12 216.9
R364 minus.n96 minus.t22 216.9
R365 minus.n102 minus.t17 216.9
R366 minus.n104 minus.t9 216.9
R367 minus.n111 minus.t21 216.9
R368 minus.n117 minus.t11 216.9
R369 minus.n64 minus.t4 216.9
R370 minus.n60 minus.n0 161.3
R371 minus.n59 minus.n58 161.3
R372 minus.n57 minus.n56 161.3
R373 minus.n55 minus.n2 161.3
R374 minus.n53 minus.n52 161.3
R375 minus.n51 minus.n3 161.3
R376 minus.n50 minus.n49 161.3
R377 minus.n47 minus.n4 161.3
R378 minus.n46 minus.n45 161.3
R379 minus.n44 minus.n5 161.3
R380 minus.n43 minus.n42 161.3
R381 minus.n41 minus.n6 161.3
R382 minus.n39 minus.n38 161.3
R383 minus.n37 minus.n8 161.3
R384 minus.n36 minus.n35 161.3
R385 minus.n33 minus.n9 161.3
R386 minus.n32 minus.n31 161.3
R387 minus.n30 minus.n29 161.3
R388 minus.n28 minus.n11 161.3
R389 minus.n27 minus.n26 161.3
R390 minus.n25 minus.n24 161.3
R391 minus.n23 minus.n13 161.3
R392 minus.n22 minus.n21 161.3
R393 minus.n20 minus.n19 161.3
R394 minus.n18 minus.n15 161.3
R395 minus.n123 minus.n63 161.3
R396 minus.n122 minus.n121 161.3
R397 minus.n120 minus.n119 161.3
R398 minus.n118 minus.n65 161.3
R399 minus.n116 minus.n115 161.3
R400 minus.n114 minus.n66 161.3
R401 minus.n113 minus.n112 161.3
R402 minus.n110 minus.n67 161.3
R403 minus.n109 minus.n108 161.3
R404 minus.n107 minus.n68 161.3
R405 minus.n106 minus.n105 161.3
R406 minus.n103 minus.n69 161.3
R407 minus.n101 minus.n100 161.3
R408 minus.n99 minus.n70 161.3
R409 minus.n98 minus.n97 161.3
R410 minus.n95 minus.n71 161.3
R411 minus.n94 minus.n93 161.3
R412 minus.n92 minus.n91 161.3
R413 minus.n90 minus.n73 161.3
R414 minus.n89 minus.n88 161.3
R415 minus.n87 minus.n86 161.3
R416 minus.n85 minus.n75 161.3
R417 minus.n84 minus.n83 161.3
R418 minus.n82 minus.n81 161.3
R419 minus.n80 minus.n77 161.3
R420 minus.n62 minus.n61 80.6037
R421 minus.n125 minus.n124 80.6037
R422 minus.n19 minus.n18 56.5617
R423 minus.n33 minus.n32 56.5617
R424 minus.n42 minus.n41 56.5617
R425 minus.n56 minus.n55 56.5617
R426 minus.n81 minus.n80 56.5617
R427 minus.n95 minus.n94 56.5617
R428 minus.n105 minus.n103 56.5617
R429 minus.n119 minus.n118 56.5617
R430 minus.n28 minus.n27 56.0773
R431 minus.n47 minus.n46 56.0773
R432 minus.n90 minus.n89 56.0773
R433 minus.n110 minus.n109 56.0773
R434 minus.n61 minus.n60 46.0096
R435 minus.n124 minus.n123 46.0096
R436 minus.n126 minus.n62 42.9706
R437 minus.n24 minus.n23 41.5458
R438 minus.n49 minus.n3 41.5458
R439 minus.n86 minus.n85 41.5458
R440 minus.n112 minus.n66 41.5458
R441 minus.n35 minus.n8 40.577
R442 minus.n39 minus.n8 40.577
R443 minus.n97 minus.n70 40.577
R444 minus.n101 minus.n70 40.577
R445 minus.n23 minus.n22 39.6083
R446 minus.n53 minus.n3 39.6083
R447 minus.n85 minus.n84 39.6083
R448 minus.n116 minus.n66 39.6083
R449 minus.n17 minus.n16 33.0515
R450 minus.n79 minus.n78 33.0515
R451 minus.n16 minus.n15 28.5514
R452 minus.n78 minus.n77 28.5514
R453 minus.n60 minus.n59 26.0455
R454 minus.n123 minus.n122 26.0455
R455 minus.n29 minus.n28 25.0767
R456 minus.n46 minus.n5 25.0767
R457 minus.n91 minus.n90 25.0767
R458 minus.n109 minus.n68 25.0767
R459 minus.n32 minus.n10 24.3464
R460 minus.n42 minus.n7 24.3464
R461 minus.n94 minus.n72 24.3464
R462 minus.n105 minus.n104 24.3464
R463 minus.n18 minus.n17 23.8546
R464 minus.n56 minus.n1 23.8546
R465 minus.n80 minus.n79 23.8546
R466 minus.n119 minus.n64 23.8546
R467 minus.n19 minus.n14 16.9689
R468 minus.n55 minus.n54 16.9689
R469 minus.n81 minus.n76 16.9689
R470 minus.n118 minus.n117 16.9689
R471 minus.n34 minus.n33 16.477
R472 minus.n41 minus.n40 16.477
R473 minus.n96 minus.n95 16.477
R474 minus.n103 minus.n102 16.477
R475 minus.n27 minus.n12 15.9852
R476 minus.n48 minus.n47 15.9852
R477 minus.n89 minus.n74 15.9852
R478 minus.n111 minus.n110 15.9852
R479 minus.n24 minus.n12 8.60764
R480 minus.n49 minus.n48 8.60764
R481 minus.n86 minus.n74 8.60764
R482 minus.n112 minus.n111 8.60764
R483 minus.n35 minus.n34 8.11581
R484 minus.n40 minus.n39 8.11581
R485 minus.n97 minus.n96 8.11581
R486 minus.n102 minus.n101 8.11581
R487 minus.n22 minus.n14 7.62397
R488 minus.n54 minus.n53 7.62397
R489 minus.n84 minus.n76 7.62397
R490 minus.n117 minus.n116 7.62397
R491 minus.n126 minus.n125 6.81155
R492 minus.n59 minus.n1 0.738255
R493 minus.n122 minus.n64 0.738255
R494 minus.n62 minus.n0 0.285035
R495 minus.n125 minus.n63 0.285035
R496 minus.n29 minus.n10 0.246418
R497 minus.n7 minus.n5 0.246418
R498 minus.n91 minus.n72 0.246418
R499 minus.n104 minus.n68 0.246418
R500 minus.n58 minus.n0 0.189894
R501 minus.n58 minus.n57 0.189894
R502 minus.n57 minus.n2 0.189894
R503 minus.n52 minus.n2 0.189894
R504 minus.n52 minus.n51 0.189894
R505 minus.n51 minus.n50 0.189894
R506 minus.n50 minus.n4 0.189894
R507 minus.n45 minus.n4 0.189894
R508 minus.n45 minus.n44 0.189894
R509 minus.n44 minus.n43 0.189894
R510 minus.n43 minus.n6 0.189894
R511 minus.n38 minus.n6 0.189894
R512 minus.n38 minus.n37 0.189894
R513 minus.n37 minus.n36 0.189894
R514 minus.n36 minus.n9 0.189894
R515 minus.n31 minus.n9 0.189894
R516 minus.n31 minus.n30 0.189894
R517 minus.n30 minus.n11 0.189894
R518 minus.n26 minus.n11 0.189894
R519 minus.n26 minus.n25 0.189894
R520 minus.n25 minus.n13 0.189894
R521 minus.n21 minus.n13 0.189894
R522 minus.n21 minus.n20 0.189894
R523 minus.n20 minus.n15 0.189894
R524 minus.n82 minus.n77 0.189894
R525 minus.n83 minus.n82 0.189894
R526 minus.n83 minus.n75 0.189894
R527 minus.n87 minus.n75 0.189894
R528 minus.n88 minus.n87 0.189894
R529 minus.n88 minus.n73 0.189894
R530 minus.n92 minus.n73 0.189894
R531 minus.n93 minus.n92 0.189894
R532 minus.n93 minus.n71 0.189894
R533 minus.n98 minus.n71 0.189894
R534 minus.n99 minus.n98 0.189894
R535 minus.n100 minus.n99 0.189894
R536 minus.n100 minus.n69 0.189894
R537 minus.n106 minus.n69 0.189894
R538 minus.n107 minus.n106 0.189894
R539 minus.n108 minus.n107 0.189894
R540 minus.n108 minus.n67 0.189894
R541 minus.n113 minus.n67 0.189894
R542 minus.n114 minus.n113 0.189894
R543 minus.n115 minus.n114 0.189894
R544 minus.n115 minus.n65 0.189894
R545 minus.n120 minus.n65 0.189894
R546 minus.n121 minus.n120 0.189894
R547 minus.n121 minus.n63 0.189894
R548 minus minus.n126 0.188
R549 drain_right.n13 drain_right.n11 66.684
R550 drain_right.n7 drain_right.n5 66.6839
R551 drain_right.n2 drain_right.n0 66.6839
R552 drain_right.n13 drain_right.n12 65.5376
R553 drain_right.n15 drain_right.n14 65.5376
R554 drain_right.n17 drain_right.n16 65.5376
R555 drain_right.n19 drain_right.n18 65.5376
R556 drain_right.n21 drain_right.n20 65.5376
R557 drain_right.n7 drain_right.n6 65.5373
R558 drain_right.n9 drain_right.n8 65.5373
R559 drain_right.n4 drain_right.n3 65.5373
R560 drain_right.n2 drain_right.n1 65.5373
R561 drain_right drain_right.n10 35.4334
R562 drain_right drain_right.n21 6.79977
R563 drain_right.n5 drain_right.t19 2.2005
R564 drain_right.n5 drain_right.t9 2.2005
R565 drain_right.n6 drain_right.t2 2.2005
R566 drain_right.n6 drain_right.t12 2.2005
R567 drain_right.n8 drain_right.t6 2.2005
R568 drain_right.n8 drain_right.t14 2.2005
R569 drain_right.n3 drain_right.t11 2.2005
R570 drain_right.n3 drain_right.t1 2.2005
R571 drain_right.n1 drain_right.t21 2.2005
R572 drain_right.n1 drain_right.t0 2.2005
R573 drain_right.n0 drain_right.t4 2.2005
R574 drain_right.n0 drain_right.t7 2.2005
R575 drain_right.n11 drain_right.t5 2.2005
R576 drain_right.n11 drain_right.t10 2.2005
R577 drain_right.n12 drain_right.t3 2.2005
R578 drain_right.n12 drain_right.t8 2.2005
R579 drain_right.n14 drain_right.t23 2.2005
R580 drain_right.n14 drain_right.t18 2.2005
R581 drain_right.n16 drain_right.t17 2.2005
R582 drain_right.n16 drain_right.t16 2.2005
R583 drain_right.n18 drain_right.t15 2.2005
R584 drain_right.n18 drain_right.t22 2.2005
R585 drain_right.n20 drain_right.t20 2.2005
R586 drain_right.n20 drain_right.t13 2.2005
R587 drain_right.n9 drain_right.n7 1.14705
R588 drain_right.n4 drain_right.n2 1.14705
R589 drain_right.n21 drain_right.n19 1.14705
R590 drain_right.n19 drain_right.n17 1.14705
R591 drain_right.n17 drain_right.n15 1.14705
R592 drain_right.n15 drain_right.n13 1.14705
R593 drain_right.n10 drain_right.n9 0.51843
R594 drain_right.n10 drain_right.n4 0.51843
C0 minus source 14.400201f
C1 plus source 14.4142f
C2 plus minus 7.80076f
C3 drain_right drain_left 2.34071f
C4 drain_left source 19.2095f
C5 drain_left minus 0.176388f
C6 plus drain_left 14.0894f
C7 drain_right source 19.2138f
C8 drain_right minus 13.6678f
C9 plus drain_right 0.582226f
C10 drain_right a_n4174_n2688# 8.271871f
C11 drain_left a_n4174_n2688# 8.8429f
C12 source a_n4174_n2688# 8.344078f
C13 minus a_n4174_n2688# 16.914732f
C14 plus a_n4174_n2688# 18.57304f
C15 drain_right.t4 a_n4174_n2688# 0.19501f
C16 drain_right.t7 a_n4174_n2688# 0.19501f
C17 drain_right.n0 a_n4174_n2688# 1.71314f
C18 drain_right.t21 a_n4174_n2688# 0.19501f
C19 drain_right.t0 a_n4174_n2688# 0.19501f
C20 drain_right.n1 a_n4174_n2688# 1.70569f
C21 drain_right.n2 a_n4174_n2688# 0.848064f
C22 drain_right.t11 a_n4174_n2688# 0.19501f
C23 drain_right.t1 a_n4174_n2688# 0.19501f
C24 drain_right.n3 a_n4174_n2688# 1.70569f
C25 drain_right.n4 a_n4174_n2688# 0.367922f
C26 drain_right.t19 a_n4174_n2688# 0.19501f
C27 drain_right.t9 a_n4174_n2688# 0.19501f
C28 drain_right.n5 a_n4174_n2688# 1.71314f
C29 drain_right.t2 a_n4174_n2688# 0.19501f
C30 drain_right.t12 a_n4174_n2688# 0.19501f
C31 drain_right.n6 a_n4174_n2688# 1.70569f
C32 drain_right.n7 a_n4174_n2688# 0.848064f
C33 drain_right.t6 a_n4174_n2688# 0.19501f
C34 drain_right.t14 a_n4174_n2688# 0.19501f
C35 drain_right.n8 a_n4174_n2688# 1.70569f
C36 drain_right.n9 a_n4174_n2688# 0.367922f
C37 drain_right.n10 a_n4174_n2688# 1.80677f
C38 drain_right.t5 a_n4174_n2688# 0.19501f
C39 drain_right.t10 a_n4174_n2688# 0.19501f
C40 drain_right.n11 a_n4174_n2688# 1.71314f
C41 drain_right.t3 a_n4174_n2688# 0.19501f
C42 drain_right.t8 a_n4174_n2688# 0.19501f
C43 drain_right.n12 a_n4174_n2688# 1.70569f
C44 drain_right.n13 a_n4174_n2688# 0.848065f
C45 drain_right.t23 a_n4174_n2688# 0.19501f
C46 drain_right.t18 a_n4174_n2688# 0.19501f
C47 drain_right.n14 a_n4174_n2688# 1.70569f
C48 drain_right.n15 a_n4174_n2688# 0.422232f
C49 drain_right.t17 a_n4174_n2688# 0.19501f
C50 drain_right.t16 a_n4174_n2688# 0.19501f
C51 drain_right.n16 a_n4174_n2688# 1.70569f
C52 drain_right.n17 a_n4174_n2688# 0.422232f
C53 drain_right.t15 a_n4174_n2688# 0.19501f
C54 drain_right.t22 a_n4174_n2688# 0.19501f
C55 drain_right.n18 a_n4174_n2688# 1.70569f
C56 drain_right.n19 a_n4174_n2688# 0.422232f
C57 drain_right.t20 a_n4174_n2688# 0.19501f
C58 drain_right.t13 a_n4174_n2688# 0.19501f
C59 drain_right.n20 a_n4174_n2688# 1.70569f
C60 drain_right.n21 a_n4174_n2688# 0.674531f
C61 minus.n0 a_n4174_n2688# 0.045577f
C62 minus.t10 a_n4174_n2688# 0.829579f
C63 minus.n1 a_n4174_n2688# 0.318431f
C64 minus.n2 a_n4174_n2688# 0.034156f
C65 minus.t8 a_n4174_n2688# 0.829579f
C66 minus.n3 a_n4174_n2688# 0.02763f
C67 minus.n4 a_n4174_n2688# 0.034156f
C68 minus.t1 a_n4174_n2688# 0.829579f
C69 minus.n5 a_n4174_n2688# 0.032975f
C70 minus.n6 a_n4174_n2688# 0.034156f
C71 minus.t6 a_n4174_n2688# 0.829579f
C72 minus.n7 a_n4174_n2688# 0.318431f
C73 minus.t7 a_n4174_n2688# 0.829579f
C74 minus.n8 a_n4174_n2688# 0.027586f
C75 minus.n9 a_n4174_n2688# 0.034156f
C76 minus.t0 a_n4174_n2688# 0.829579f
C77 minus.t5 a_n4174_n2688# 0.829579f
C78 minus.n10 a_n4174_n2688# 0.318431f
C79 minus.n11 a_n4174_n2688# 0.034156f
C80 minus.t20 a_n4174_n2688# 0.829579f
C81 minus.n12 a_n4174_n2688# 0.318431f
C82 minus.n13 a_n4174_n2688# 0.034156f
C83 minus.t15 a_n4174_n2688# 0.829579f
C84 minus.n14 a_n4174_n2688# 0.318431f
C85 minus.n15 a_n4174_n2688# 0.171949f
C86 minus.t18 a_n4174_n2688# 0.829579f
C87 minus.t13 a_n4174_n2688# 0.911374f
C88 minus.n16 a_n4174_n2688# 0.359428f
C89 minus.n17 a_n4174_n2688# 0.369716f
C90 minus.n18 a_n4174_n2688# 0.042098f
C91 minus.n19 a_n4174_n2688# 0.046572f
C92 minus.n20 a_n4174_n2688# 0.034156f
C93 minus.n21 a_n4174_n2688# 0.034156f
C94 minus.n22 a_n4174_n2688# 0.046268f
C95 minus.n23 a_n4174_n2688# 0.02763f
C96 minus.n24 a_n4174_n2688# 0.046842f
C97 minus.n25 a_n4174_n2688# 0.034156f
C98 minus.n26 a_n4174_n2688# 0.034156f
C99 minus.n27 a_n4174_n2688# 0.047128f
C100 minus.n28 a_n4174_n2688# 0.040638f
C101 minus.n29 a_n4174_n2688# 0.032975f
C102 minus.n30 a_n4174_n2688# 0.034156f
C103 minus.n31 a_n4174_n2688# 0.034156f
C104 minus.n32 a_n4174_n2688# 0.041778f
C105 minus.n33 a_n4174_n2688# 0.046892f
C106 minus.n34 a_n4174_n2688# 0.318431f
C107 minus.n35 a_n4174_n2688# 0.046577f
C108 minus.n36 a_n4174_n2688# 0.034156f
C109 minus.n37 a_n4174_n2688# 0.034156f
C110 minus.n38 a_n4174_n2688# 0.034156f
C111 minus.n39 a_n4174_n2688# 0.046577f
C112 minus.n40 a_n4174_n2688# 0.318431f
C113 minus.n41 a_n4174_n2688# 0.046892f
C114 minus.n42 a_n4174_n2688# 0.041778f
C115 minus.n43 a_n4174_n2688# 0.034156f
C116 minus.n44 a_n4174_n2688# 0.034156f
C117 minus.n45 a_n4174_n2688# 0.034156f
C118 minus.n46 a_n4174_n2688# 0.040638f
C119 minus.n47 a_n4174_n2688# 0.047128f
C120 minus.n48 a_n4174_n2688# 0.318431f
C121 minus.n49 a_n4174_n2688# 0.046842f
C122 minus.n50 a_n4174_n2688# 0.034156f
C123 minus.n51 a_n4174_n2688# 0.034156f
C124 minus.n52 a_n4174_n2688# 0.034156f
C125 minus.n53 a_n4174_n2688# 0.046268f
C126 minus.n54 a_n4174_n2688# 0.318431f
C127 minus.n55 a_n4174_n2688# 0.046572f
C128 minus.n56 a_n4174_n2688# 0.042098f
C129 minus.n57 a_n4174_n2688# 0.034156f
C130 minus.n58 a_n4174_n2688# 0.034156f
C131 minus.n59 a_n4174_n2688# 0.034648f
C132 minus.n60 a_n4174_n2688# 0.035819f
C133 minus.t3 a_n4174_n2688# 0.881587f
C134 minus.n61 a_n4174_n2688# 0.368465f
C135 minus.n62 a_n4174_n2688# 1.5832f
C136 minus.n63 a_n4174_n2688# 0.045577f
C137 minus.t4 a_n4174_n2688# 0.829579f
C138 minus.n64 a_n4174_n2688# 0.318431f
C139 minus.n65 a_n4174_n2688# 0.034156f
C140 minus.t11 a_n4174_n2688# 0.829579f
C141 minus.n66 a_n4174_n2688# 0.02763f
C142 minus.n67 a_n4174_n2688# 0.034156f
C143 minus.t21 a_n4174_n2688# 0.829579f
C144 minus.n68 a_n4174_n2688# 0.032975f
C145 minus.n69 a_n4174_n2688# 0.034156f
C146 minus.t17 a_n4174_n2688# 0.829579f
C147 minus.n70 a_n4174_n2688# 0.027586f
C148 minus.n71 a_n4174_n2688# 0.034156f
C149 minus.t22 a_n4174_n2688# 0.829579f
C150 minus.t12 a_n4174_n2688# 0.829579f
C151 minus.n72 a_n4174_n2688# 0.318431f
C152 minus.n73 a_n4174_n2688# 0.034156f
C153 minus.t23 a_n4174_n2688# 0.829579f
C154 minus.n74 a_n4174_n2688# 0.318431f
C155 minus.n75 a_n4174_n2688# 0.034156f
C156 minus.t2 a_n4174_n2688# 0.829579f
C157 minus.n76 a_n4174_n2688# 0.318431f
C158 minus.n77 a_n4174_n2688# 0.171949f
C159 minus.t16 a_n4174_n2688# 0.829579f
C160 minus.t19 a_n4174_n2688# 0.911374f
C161 minus.n78 a_n4174_n2688# 0.359428f
C162 minus.n79 a_n4174_n2688# 0.369716f
C163 minus.n80 a_n4174_n2688# 0.042098f
C164 minus.n81 a_n4174_n2688# 0.046572f
C165 minus.n82 a_n4174_n2688# 0.034156f
C166 minus.n83 a_n4174_n2688# 0.034156f
C167 minus.n84 a_n4174_n2688# 0.046268f
C168 minus.n85 a_n4174_n2688# 0.02763f
C169 minus.n86 a_n4174_n2688# 0.046842f
C170 minus.n87 a_n4174_n2688# 0.034156f
C171 minus.n88 a_n4174_n2688# 0.034156f
C172 minus.n89 a_n4174_n2688# 0.047128f
C173 minus.n90 a_n4174_n2688# 0.040638f
C174 minus.n91 a_n4174_n2688# 0.032975f
C175 minus.n92 a_n4174_n2688# 0.034156f
C176 minus.n93 a_n4174_n2688# 0.034156f
C177 minus.n94 a_n4174_n2688# 0.041778f
C178 minus.n95 a_n4174_n2688# 0.046892f
C179 minus.n96 a_n4174_n2688# 0.318431f
C180 minus.n97 a_n4174_n2688# 0.046577f
C181 minus.n98 a_n4174_n2688# 0.034156f
C182 minus.n99 a_n4174_n2688# 0.034156f
C183 minus.n100 a_n4174_n2688# 0.034156f
C184 minus.n101 a_n4174_n2688# 0.046577f
C185 minus.n102 a_n4174_n2688# 0.318431f
C186 minus.n103 a_n4174_n2688# 0.046892f
C187 minus.t9 a_n4174_n2688# 0.829579f
C188 minus.n104 a_n4174_n2688# 0.318431f
C189 minus.n105 a_n4174_n2688# 0.041778f
C190 minus.n106 a_n4174_n2688# 0.034156f
C191 minus.n107 a_n4174_n2688# 0.034156f
C192 minus.n108 a_n4174_n2688# 0.034156f
C193 minus.n109 a_n4174_n2688# 0.040638f
C194 minus.n110 a_n4174_n2688# 0.047128f
C195 minus.n111 a_n4174_n2688# 0.318431f
C196 minus.n112 a_n4174_n2688# 0.046842f
C197 minus.n113 a_n4174_n2688# 0.034156f
C198 minus.n114 a_n4174_n2688# 0.034156f
C199 minus.n115 a_n4174_n2688# 0.034156f
C200 minus.n116 a_n4174_n2688# 0.046268f
C201 minus.n117 a_n4174_n2688# 0.318431f
C202 minus.n118 a_n4174_n2688# 0.046572f
C203 minus.n119 a_n4174_n2688# 0.042098f
C204 minus.n120 a_n4174_n2688# 0.034156f
C205 minus.n121 a_n4174_n2688# 0.034156f
C206 minus.n122 a_n4174_n2688# 0.034648f
C207 minus.n123 a_n4174_n2688# 0.035819f
C208 minus.t14 a_n4174_n2688# 0.881587f
C209 minus.n124 a_n4174_n2688# 0.368465f
C210 minus.n125 a_n4174_n2688# 0.259918f
C211 minus.n126 a_n4174_n2688# 1.86604f
C212 source.t42 a_n4174_n2688# 1.86195f
C213 source.n0 a_n4174_n2688# 1.15042f
C214 source.t34 a_n4174_n2688# 0.17461f
C215 source.t39 a_n4174_n2688# 0.17461f
C216 source.n1 a_n4174_n2688# 1.46172f
C217 source.n2 a_n4174_n2688# 0.410228f
C218 source.t38 a_n4174_n2688# 0.17461f
C219 source.t41 a_n4174_n2688# 0.17461f
C220 source.n3 a_n4174_n2688# 1.46172f
C221 source.n4 a_n4174_n2688# 0.410228f
C222 source.t43 a_n4174_n2688# 0.17461f
C223 source.t33 a_n4174_n2688# 0.17461f
C224 source.n5 a_n4174_n2688# 1.46172f
C225 source.n6 a_n4174_n2688# 0.410228f
C226 source.t44 a_n4174_n2688# 0.17461f
C227 source.t37 a_n4174_n2688# 0.17461f
C228 source.n7 a_n4174_n2688# 1.46172f
C229 source.n8 a_n4174_n2688# 0.410228f
C230 source.t45 a_n4174_n2688# 0.17461f
C231 source.t47 a_n4174_n2688# 0.17461f
C232 source.n9 a_n4174_n2688# 1.46172f
C233 source.n10 a_n4174_n2688# 0.410228f
C234 source.t26 a_n4174_n2688# 1.86195f
C235 source.n11 a_n4174_n2688# 0.432671f
C236 source.t10 a_n4174_n2688# 1.86195f
C237 source.n12 a_n4174_n2688# 0.432671f
C238 source.t18 a_n4174_n2688# 0.17461f
C239 source.t17 a_n4174_n2688# 0.17461f
C240 source.n13 a_n4174_n2688# 1.46172f
C241 source.n14 a_n4174_n2688# 0.410228f
C242 source.t15 a_n4174_n2688# 0.17461f
C243 source.t21 a_n4174_n2688# 0.17461f
C244 source.n15 a_n4174_n2688# 1.46172f
C245 source.n16 a_n4174_n2688# 0.410228f
C246 source.t9 a_n4174_n2688# 0.17461f
C247 source.t22 a_n4174_n2688# 0.17461f
C248 source.n17 a_n4174_n2688# 1.46172f
C249 source.n18 a_n4174_n2688# 0.410228f
C250 source.t6 a_n4174_n2688# 0.17461f
C251 source.t11 a_n4174_n2688# 0.17461f
C252 source.n19 a_n4174_n2688# 1.46172f
C253 source.n20 a_n4174_n2688# 0.410228f
C254 source.t7 a_n4174_n2688# 0.17461f
C255 source.t4 a_n4174_n2688# 0.17461f
C256 source.n21 a_n4174_n2688# 1.46172f
C257 source.n22 a_n4174_n2688# 0.410228f
C258 source.t1 a_n4174_n2688# 1.86195f
C259 source.n23 a_n4174_n2688# 1.52287f
C260 source.t32 a_n4174_n2688# 1.86195f
C261 source.n24 a_n4174_n2688# 1.52288f
C262 source.t24 a_n4174_n2688# 0.17461f
C263 source.t40 a_n4174_n2688# 0.17461f
C264 source.n25 a_n4174_n2688# 1.46172f
C265 source.n26 a_n4174_n2688# 0.410232f
C266 source.t35 a_n4174_n2688# 0.17461f
C267 source.t46 a_n4174_n2688# 0.17461f
C268 source.n27 a_n4174_n2688# 1.46172f
C269 source.n28 a_n4174_n2688# 0.410232f
C270 source.t31 a_n4174_n2688# 0.17461f
C271 source.t28 a_n4174_n2688# 0.17461f
C272 source.n29 a_n4174_n2688# 1.46172f
C273 source.n30 a_n4174_n2688# 0.410232f
C274 source.t36 a_n4174_n2688# 0.17461f
C275 source.t30 a_n4174_n2688# 0.17461f
C276 source.n31 a_n4174_n2688# 1.46172f
C277 source.n32 a_n4174_n2688# 0.410232f
C278 source.t25 a_n4174_n2688# 0.17461f
C279 source.t29 a_n4174_n2688# 0.17461f
C280 source.n33 a_n4174_n2688# 1.46172f
C281 source.n34 a_n4174_n2688# 0.410232f
C282 source.t27 a_n4174_n2688# 1.86195f
C283 source.n35 a_n4174_n2688# 0.432675f
C284 source.t12 a_n4174_n2688# 1.86195f
C285 source.n36 a_n4174_n2688# 0.432675f
C286 source.t0 a_n4174_n2688# 0.17461f
C287 source.t8 a_n4174_n2688# 0.17461f
C288 source.n37 a_n4174_n2688# 1.46172f
C289 source.n38 a_n4174_n2688# 0.410232f
C290 source.t23 a_n4174_n2688# 0.17461f
C291 source.t3 a_n4174_n2688# 0.17461f
C292 source.n39 a_n4174_n2688# 1.46172f
C293 source.n40 a_n4174_n2688# 0.410232f
C294 source.t19 a_n4174_n2688# 0.17461f
C295 source.t5 a_n4174_n2688# 0.17461f
C296 source.n41 a_n4174_n2688# 1.46172f
C297 source.n42 a_n4174_n2688# 0.410232f
C298 source.t16 a_n4174_n2688# 0.17461f
C299 source.t20 a_n4174_n2688# 0.17461f
C300 source.n43 a_n4174_n2688# 1.46172f
C301 source.n44 a_n4174_n2688# 0.410232f
C302 source.t14 a_n4174_n2688# 0.17461f
C303 source.t2 a_n4174_n2688# 0.17461f
C304 source.n45 a_n4174_n2688# 1.46172f
C305 source.n46 a_n4174_n2688# 0.410232f
C306 source.t13 a_n4174_n2688# 1.86195f
C307 source.n47 a_n4174_n2688# 0.608685f
C308 source.n48 a_n4174_n2688# 1.30411f
C309 drain_left.t12 a_n4174_n2688# 0.196627f
C310 drain_left.t0 a_n4174_n2688# 0.196627f
C311 drain_left.n0 a_n4174_n2688# 1.72734f
C312 drain_left.t4 a_n4174_n2688# 0.196627f
C313 drain_left.t2 a_n4174_n2688# 0.196627f
C314 drain_left.n1 a_n4174_n2688# 1.71983f
C315 drain_left.n2 a_n4174_n2688# 0.855096f
C316 drain_left.t23 a_n4174_n2688# 0.196627f
C317 drain_left.t10 a_n4174_n2688# 0.196627f
C318 drain_left.n3 a_n4174_n2688# 1.71983f
C319 drain_left.n4 a_n4174_n2688# 0.370973f
C320 drain_left.t14 a_n4174_n2688# 0.196627f
C321 drain_left.t13 a_n4174_n2688# 0.196627f
C322 drain_left.n5 a_n4174_n2688# 1.72734f
C323 drain_left.t5 a_n4174_n2688# 0.196627f
C324 drain_left.t8 a_n4174_n2688# 0.196627f
C325 drain_left.n6 a_n4174_n2688# 1.71983f
C326 drain_left.n7 a_n4174_n2688# 0.855096f
C327 drain_left.t15 a_n4174_n2688# 0.196627f
C328 drain_left.t3 a_n4174_n2688# 0.196627f
C329 drain_left.n8 a_n4174_n2688# 1.71983f
C330 drain_left.n9 a_n4174_n2688# 0.370973f
C331 drain_left.n10 a_n4174_n2688# 1.87677f
C332 drain_left.t22 a_n4174_n2688# 0.196627f
C333 drain_left.t9 a_n4174_n2688# 0.196627f
C334 drain_left.n11 a_n4174_n2688# 1.72735f
C335 drain_left.t21 a_n4174_n2688# 0.196627f
C336 drain_left.t1 a_n4174_n2688# 0.196627f
C337 drain_left.n12 a_n4174_n2688# 1.71984f
C338 drain_left.n13 a_n4174_n2688# 0.855089f
C339 drain_left.t6 a_n4174_n2688# 0.196627f
C340 drain_left.t7 a_n4174_n2688# 0.196627f
C341 drain_left.n14 a_n4174_n2688# 1.71984f
C342 drain_left.n15 a_n4174_n2688# 0.425732f
C343 drain_left.t11 a_n4174_n2688# 0.196627f
C344 drain_left.t17 a_n4174_n2688# 0.196627f
C345 drain_left.n16 a_n4174_n2688# 1.71984f
C346 drain_left.n17 a_n4174_n2688# 0.425732f
C347 drain_left.t16 a_n4174_n2688# 0.196627f
C348 drain_left.t19 a_n4174_n2688# 0.196627f
C349 drain_left.n18 a_n4174_n2688# 1.71984f
C350 drain_left.n19 a_n4174_n2688# 0.425732f
C351 drain_left.t20 a_n4174_n2688# 0.196627f
C352 drain_left.t18 a_n4174_n2688# 0.196627f
C353 drain_left.n20 a_n4174_n2688# 1.71983f
C354 drain_left.n21 a_n4174_n2688# 0.680131f
C355 plus.n0 a_n4174_n2688# 0.046173f
C356 plus.t5 a_n4174_n2688# 0.893128f
C357 plus.t8 a_n4174_n2688# 0.840439f
C358 plus.n1 a_n4174_n2688# 0.322599f
C359 plus.n2 a_n4174_n2688# 0.034603f
C360 plus.t13 a_n4174_n2688# 0.840439f
C361 plus.n3 a_n4174_n2688# 0.027992f
C362 plus.n4 a_n4174_n2688# 0.034603f
C363 plus.t6 a_n4174_n2688# 0.840439f
C364 plus.n5 a_n4174_n2688# 0.033406f
C365 plus.n6 a_n4174_n2688# 0.034603f
C366 plus.t14 a_n4174_n2688# 0.840439f
C367 plus.n7 a_n4174_n2688# 0.027948f
C368 plus.n8 a_n4174_n2688# 0.034603f
C369 plus.t4 a_n4174_n2688# 0.840439f
C370 plus.t10 a_n4174_n2688# 0.840439f
C371 plus.n9 a_n4174_n2688# 0.322599f
C372 plus.n10 a_n4174_n2688# 0.034603f
C373 plus.t3 a_n4174_n2688# 0.840439f
C374 plus.n11 a_n4174_n2688# 0.322599f
C375 plus.n12 a_n4174_n2688# 0.034603f
C376 plus.t0 a_n4174_n2688# 0.840439f
C377 plus.n13 a_n4174_n2688# 0.322599f
C378 plus.n14 a_n4174_n2688# 0.174201f
C379 plus.t2 a_n4174_n2688# 0.840439f
C380 plus.t21 a_n4174_n2688# 0.923305f
C381 plus.n15 a_n4174_n2688# 0.364133f
C382 plus.n16 a_n4174_n2688# 0.374556f
C383 plus.n17 a_n4174_n2688# 0.042649f
C384 plus.n18 a_n4174_n2688# 0.047182f
C385 plus.n19 a_n4174_n2688# 0.034603f
C386 plus.n20 a_n4174_n2688# 0.034603f
C387 plus.n21 a_n4174_n2688# 0.046874f
C388 plus.n22 a_n4174_n2688# 0.027992f
C389 plus.n23 a_n4174_n2688# 0.047455f
C390 plus.n24 a_n4174_n2688# 0.034603f
C391 plus.n25 a_n4174_n2688# 0.034603f
C392 plus.n26 a_n4174_n2688# 0.047745f
C393 plus.n27 a_n4174_n2688# 0.04117f
C394 plus.n28 a_n4174_n2688# 0.033406f
C395 plus.n29 a_n4174_n2688# 0.034603f
C396 plus.n30 a_n4174_n2688# 0.034603f
C397 plus.n31 a_n4174_n2688# 0.042325f
C398 plus.n32 a_n4174_n2688# 0.047506f
C399 plus.n33 a_n4174_n2688# 0.322599f
C400 plus.n34 a_n4174_n2688# 0.047187f
C401 plus.n35 a_n4174_n2688# 0.034603f
C402 plus.n36 a_n4174_n2688# 0.034603f
C403 plus.n37 a_n4174_n2688# 0.034603f
C404 plus.n38 a_n4174_n2688# 0.047187f
C405 plus.n39 a_n4174_n2688# 0.322599f
C406 plus.n40 a_n4174_n2688# 0.047506f
C407 plus.t9 a_n4174_n2688# 0.840439f
C408 plus.n41 a_n4174_n2688# 0.322599f
C409 plus.n42 a_n4174_n2688# 0.042325f
C410 plus.n43 a_n4174_n2688# 0.034603f
C411 plus.n44 a_n4174_n2688# 0.034603f
C412 plus.n45 a_n4174_n2688# 0.034603f
C413 plus.n46 a_n4174_n2688# 0.04117f
C414 plus.n47 a_n4174_n2688# 0.047745f
C415 plus.n48 a_n4174_n2688# 0.322599f
C416 plus.n49 a_n4174_n2688# 0.047455f
C417 plus.n50 a_n4174_n2688# 0.034603f
C418 plus.n51 a_n4174_n2688# 0.034603f
C419 plus.n52 a_n4174_n2688# 0.034603f
C420 plus.n53 a_n4174_n2688# 0.046874f
C421 plus.n54 a_n4174_n2688# 0.322599f
C422 plus.n55 a_n4174_n2688# 0.047182f
C423 plus.n56 a_n4174_n2688# 0.042649f
C424 plus.n57 a_n4174_n2688# 0.034603f
C425 plus.n58 a_n4174_n2688# 0.034603f
C426 plus.n59 a_n4174_n2688# 0.035102f
C427 plus.n60 a_n4174_n2688# 0.036288f
C428 plus.n61 a_n4174_n2688# 0.373289f
C429 plus.n62 a_n4174_n2688# 0.377978f
C430 plus.n63 a_n4174_n2688# 0.046173f
C431 plus.t15 a_n4174_n2688# 0.893128f
C432 plus.t23 a_n4174_n2688# 0.840439f
C433 plus.n64 a_n4174_n2688# 0.322599f
C434 plus.n65 a_n4174_n2688# 0.034603f
C435 plus.t7 a_n4174_n2688# 0.840439f
C436 plus.n66 a_n4174_n2688# 0.027992f
C437 plus.n67 a_n4174_n2688# 0.034603f
C438 plus.t12 a_n4174_n2688# 0.840439f
C439 plus.n68 a_n4174_n2688# 0.033406f
C440 plus.n69 a_n4174_n2688# 0.034603f
C441 plus.t1 a_n4174_n2688# 0.840439f
C442 plus.n70 a_n4174_n2688# 0.322599f
C443 plus.t16 a_n4174_n2688# 0.840439f
C444 plus.n71 a_n4174_n2688# 0.027948f
C445 plus.n72 a_n4174_n2688# 0.034603f
C446 plus.t19 a_n4174_n2688# 0.840439f
C447 plus.t11 a_n4174_n2688# 0.840439f
C448 plus.n73 a_n4174_n2688# 0.322599f
C449 plus.n74 a_n4174_n2688# 0.034603f
C450 plus.t17 a_n4174_n2688# 0.840439f
C451 plus.n75 a_n4174_n2688# 0.322599f
C452 plus.n76 a_n4174_n2688# 0.034603f
C453 plus.t22 a_n4174_n2688# 0.840439f
C454 plus.n77 a_n4174_n2688# 0.322599f
C455 plus.n78 a_n4174_n2688# 0.174201f
C456 plus.t18 a_n4174_n2688# 0.840439f
C457 plus.t20 a_n4174_n2688# 0.923305f
C458 plus.n79 a_n4174_n2688# 0.364133f
C459 plus.n80 a_n4174_n2688# 0.374556f
C460 plus.n81 a_n4174_n2688# 0.042649f
C461 plus.n82 a_n4174_n2688# 0.047182f
C462 plus.n83 a_n4174_n2688# 0.034603f
C463 plus.n84 a_n4174_n2688# 0.034603f
C464 plus.n85 a_n4174_n2688# 0.046874f
C465 plus.n86 a_n4174_n2688# 0.027992f
C466 plus.n87 a_n4174_n2688# 0.047455f
C467 plus.n88 a_n4174_n2688# 0.034603f
C468 plus.n89 a_n4174_n2688# 0.034603f
C469 plus.n90 a_n4174_n2688# 0.047745f
C470 plus.n91 a_n4174_n2688# 0.04117f
C471 plus.n92 a_n4174_n2688# 0.033406f
C472 plus.n93 a_n4174_n2688# 0.034603f
C473 plus.n94 a_n4174_n2688# 0.034603f
C474 plus.n95 a_n4174_n2688# 0.042325f
C475 plus.n96 a_n4174_n2688# 0.047506f
C476 plus.n97 a_n4174_n2688# 0.322599f
C477 plus.n98 a_n4174_n2688# 0.047187f
C478 plus.n99 a_n4174_n2688# 0.034603f
C479 plus.n100 a_n4174_n2688# 0.034603f
C480 plus.n101 a_n4174_n2688# 0.034603f
C481 plus.n102 a_n4174_n2688# 0.047187f
C482 plus.n103 a_n4174_n2688# 0.322599f
C483 plus.n104 a_n4174_n2688# 0.047506f
C484 plus.n105 a_n4174_n2688# 0.042325f
C485 plus.n106 a_n4174_n2688# 0.034603f
C486 plus.n107 a_n4174_n2688# 0.034603f
C487 plus.n108 a_n4174_n2688# 0.034603f
C488 plus.n109 a_n4174_n2688# 0.04117f
C489 plus.n110 a_n4174_n2688# 0.047745f
C490 plus.n111 a_n4174_n2688# 0.322599f
C491 plus.n112 a_n4174_n2688# 0.047455f
C492 plus.n113 a_n4174_n2688# 0.034603f
C493 plus.n114 a_n4174_n2688# 0.034603f
C494 plus.n115 a_n4174_n2688# 0.034603f
C495 plus.n116 a_n4174_n2688# 0.046874f
C496 plus.n117 a_n4174_n2688# 0.322599f
C497 plus.n118 a_n4174_n2688# 0.047182f
C498 plus.n119 a_n4174_n2688# 0.042649f
C499 plus.n120 a_n4174_n2688# 0.034603f
C500 plus.n121 a_n4174_n2688# 0.034603f
C501 plus.n122 a_n4174_n2688# 0.035102f
C502 plus.n123 a_n4174_n2688# 0.036288f
C503 plus.n124 a_n4174_n2688# 0.373289f
C504 plus.n125 a_n4174_n2688# 1.42684f
.ends

