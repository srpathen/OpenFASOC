* NGSPICE file created from diffpair.ext - technology: sky130A

.subckt diffpair minus drain_right drain_left source plus
X0 a_n2874_n2688# a_n2874_n2688# a_n2874_n2688# a_n2874_n2688# sky130_fd_pr__nfet_01v8 ad=3.51 pd=18.78 as=28.08 ps=150.24 w=9 l=0.5
X1 drain_right.t23 minus.t0 source.t26 a_n2874_n2688# sky130_fd_pr__nfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X2 source.t30 minus.t1 drain_right.t22 a_n2874_n2688# sky130_fd_pr__nfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X3 drain_left.t23 plus.t0 source.t1 a_n2874_n2688# sky130_fd_pr__nfet_01v8 ad=1.485 pd=9.33 as=3.51 ps=18.78 w=9 l=0.5
X4 source.t5 plus.t1 drain_left.t22 a_n2874_n2688# sky130_fd_pr__nfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X5 drain_left.t21 plus.t2 source.t35 a_n2874_n2688# sky130_fd_pr__nfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X6 drain_left.t20 plus.t3 source.t37 a_n2874_n2688# sky130_fd_pr__nfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X7 source.t23 minus.t2 drain_right.t21 a_n2874_n2688# sky130_fd_pr__nfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X8 source.t42 plus.t4 drain_left.t19 a_n2874_n2688# sky130_fd_pr__nfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X9 drain_right.t20 minus.t3 source.t22 a_n2874_n2688# sky130_fd_pr__nfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X10 a_n2874_n2688# a_n2874_n2688# a_n2874_n2688# a_n2874_n2688# sky130_fd_pr__nfet_01v8 ad=3.51 pd=18.78 as=0 ps=0 w=9 l=0.5
X11 source.t43 plus.t5 drain_left.t18 a_n2874_n2688# sky130_fd_pr__nfet_01v8 ad=3.51 pd=18.78 as=1.485 ps=9.33 w=9 l=0.5
X12 source.t20 minus.t4 drain_right.t19 a_n2874_n2688# sky130_fd_pr__nfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X13 drain_left.t17 plus.t6 source.t46 a_n2874_n2688# sky130_fd_pr__nfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X14 source.t47 plus.t7 drain_left.t16 a_n2874_n2688# sky130_fd_pr__nfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X15 drain_right.t18 minus.t5 source.t32 a_n2874_n2688# sky130_fd_pr__nfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X16 source.t3 plus.t8 drain_left.t15 a_n2874_n2688# sky130_fd_pr__nfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X17 drain_right.t17 minus.t6 source.t24 a_n2874_n2688# sky130_fd_pr__nfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X18 drain_right.t16 minus.t7 source.t18 a_n2874_n2688# sky130_fd_pr__nfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X19 source.t34 minus.t8 drain_right.t15 a_n2874_n2688# sky130_fd_pr__nfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X20 source.t19 minus.t9 drain_right.t14 a_n2874_n2688# sky130_fd_pr__nfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X21 drain_left.t14 plus.t9 source.t0 a_n2874_n2688# sky130_fd_pr__nfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X22 source.t27 minus.t10 drain_right.t13 a_n2874_n2688# sky130_fd_pr__nfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X23 drain_right.t12 minus.t11 source.t31 a_n2874_n2688# sky130_fd_pr__nfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X24 source.t2 plus.t10 drain_left.t13 a_n2874_n2688# sky130_fd_pr__nfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X25 source.t25 minus.t12 drain_right.t11 a_n2874_n2688# sky130_fd_pr__nfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X26 source.t21 minus.t13 drain_right.t10 a_n2874_n2688# sky130_fd_pr__nfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X27 a_n2874_n2688# a_n2874_n2688# a_n2874_n2688# a_n2874_n2688# sky130_fd_pr__nfet_01v8 ad=3.51 pd=18.78 as=0 ps=0 w=9 l=0.5
X28 drain_right.t9 minus.t14 source.t33 a_n2874_n2688# sky130_fd_pr__nfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X29 source.t41 plus.t11 drain_left.t12 a_n2874_n2688# sky130_fd_pr__nfet_01v8 ad=3.51 pd=18.78 as=1.485 ps=9.33 w=9 l=0.5
X30 drain_left.t11 plus.t12 source.t38 a_n2874_n2688# sky130_fd_pr__nfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X31 drain_right.t8 minus.t15 source.t14 a_n2874_n2688# sky130_fd_pr__nfet_01v8 ad=1.485 pd=9.33 as=3.51 ps=18.78 w=9 l=0.5
X32 drain_right.t7 minus.t16 source.t17 a_n2874_n2688# sky130_fd_pr__nfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X33 a_n2874_n2688# a_n2874_n2688# a_n2874_n2688# a_n2874_n2688# sky130_fd_pr__nfet_01v8 ad=3.51 pd=18.78 as=0 ps=0 w=9 l=0.5
X34 drain_left.t10 plus.t13 source.t9 a_n2874_n2688# sky130_fd_pr__nfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X35 drain_right.t6 minus.t17 source.t15 a_n2874_n2688# sky130_fd_pr__nfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X36 drain_left.t9 plus.t14 source.t36 a_n2874_n2688# sky130_fd_pr__nfet_01v8 ad=1.485 pd=9.33 as=3.51 ps=18.78 w=9 l=0.5
X37 source.t39 plus.t15 drain_left.t8 a_n2874_n2688# sky130_fd_pr__nfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X38 source.t12 minus.t18 drain_right.t5 a_n2874_n2688# sky130_fd_pr__nfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X39 source.t6 plus.t16 drain_left.t7 a_n2874_n2688# sky130_fd_pr__nfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X40 source.t28 minus.t19 drain_right.t4 a_n2874_n2688# sky130_fd_pr__nfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X41 source.t8 plus.t17 drain_left.t6 a_n2874_n2688# sky130_fd_pr__nfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X42 drain_right.t3 minus.t20 source.t11 a_n2874_n2688# sky130_fd_pr__nfet_01v8 ad=1.485 pd=9.33 as=3.51 ps=18.78 w=9 l=0.5
X43 source.t45 plus.t18 drain_left.t5 a_n2874_n2688# sky130_fd_pr__nfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X44 drain_left.t4 plus.t19 source.t44 a_n2874_n2688# sky130_fd_pr__nfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X45 source.t29 minus.t21 drain_right.t2 a_n2874_n2688# sky130_fd_pr__nfet_01v8 ad=3.51 pd=18.78 as=1.485 ps=9.33 w=9 l=0.5
X46 drain_left.t3 plus.t20 source.t10 a_n2874_n2688# sky130_fd_pr__nfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X47 source.t7 plus.t21 drain_left.t2 a_n2874_n2688# sky130_fd_pr__nfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X48 drain_right.t1 minus.t22 source.t16 a_n2874_n2688# sky130_fd_pr__nfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X49 source.t13 minus.t23 drain_right.t0 a_n2874_n2688# sky130_fd_pr__nfet_01v8 ad=3.51 pd=18.78 as=1.485 ps=9.33 w=9 l=0.5
X50 drain_left.t1 plus.t22 source.t4 a_n2874_n2688# sky130_fd_pr__nfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X51 drain_left.t0 plus.t23 source.t40 a_n2874_n2688# sky130_fd_pr__nfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
R0 minus.n9 minus.t15 538.725
R1 minus.n43 minus.t23 538.725
R2 minus.n8 minus.t2 512.366
R3 minus.n7 minus.t7 512.366
R4 minus.n13 minus.t18 512.366
R5 minus.n5 minus.t5 512.366
R6 minus.n18 minus.t12 512.366
R7 minus.n20 minus.t0 512.366
R8 minus.n3 minus.t13 512.366
R9 minus.n25 minus.t17 512.366
R10 minus.n1 minus.t4 512.366
R11 minus.n30 minus.t16 512.366
R12 minus.n32 minus.t21 512.366
R13 minus.n42 minus.t22 512.366
R14 minus.n41 minus.t9 512.366
R15 minus.n47 minus.t6 512.366
R16 minus.n39 minus.t1 512.366
R17 minus.n52 minus.t11 512.366
R18 minus.n54 minus.t10 512.366
R19 minus.n37 minus.t3 512.366
R20 minus.n59 minus.t19 512.366
R21 minus.n35 minus.t14 512.366
R22 minus.n64 minus.t8 512.366
R23 minus.n66 minus.t20 512.366
R24 minus.n33 minus.n32 161.3
R25 minus.n31 minus.n0 161.3
R26 minus.n30 minus.n29 161.3
R27 minus.n28 minus.n1 161.3
R28 minus.n27 minus.n26 161.3
R29 minus.n25 minus.n2 161.3
R30 minus.n24 minus.n23 161.3
R31 minus.n22 minus.n3 161.3
R32 minus.n21 minus.n20 161.3
R33 minus.n19 minus.n4 161.3
R34 minus.n18 minus.n17 161.3
R35 minus.n16 minus.n5 161.3
R36 minus.n15 minus.n14 161.3
R37 minus.n13 minus.n6 161.3
R38 minus.n12 minus.n11 161.3
R39 minus.n10 minus.n7 161.3
R40 minus.n67 minus.n66 161.3
R41 minus.n65 minus.n34 161.3
R42 minus.n64 minus.n63 161.3
R43 minus.n62 minus.n35 161.3
R44 minus.n61 minus.n60 161.3
R45 minus.n59 minus.n36 161.3
R46 minus.n58 minus.n57 161.3
R47 minus.n56 minus.n37 161.3
R48 minus.n55 minus.n54 161.3
R49 minus.n53 minus.n38 161.3
R50 minus.n52 minus.n51 161.3
R51 minus.n50 minus.n39 161.3
R52 minus.n49 minus.n48 161.3
R53 minus.n47 minus.n40 161.3
R54 minus.n46 minus.n45 161.3
R55 minus.n44 minus.n41 161.3
R56 minus.n8 minus.n7 48.2005
R57 minus.n18 minus.n5 48.2005
R58 minus.n20 minus.n3 48.2005
R59 minus.n30 minus.n1 48.2005
R60 minus.n42 minus.n41 48.2005
R61 minus.n52 minus.n39 48.2005
R62 minus.n54 minus.n37 48.2005
R63 minus.n64 minus.n35 48.2005
R64 minus.n14 minus.n13 47.4702
R65 minus.n25 minus.n24 47.4702
R66 minus.n48 minus.n47 47.4702
R67 minus.n59 minus.n58 47.4702
R68 minus.n32 minus.n31 46.0096
R69 minus.n66 minus.n65 46.0096
R70 minus.n10 minus.n9 45.0871
R71 minus.n44 minus.n43 45.0871
R72 minus.n68 minus.n33 37.7619
R73 minus.n13 minus.n12 25.5611
R74 minus.n26 minus.n25 25.5611
R75 minus.n47 minus.n46 25.5611
R76 minus.n60 minus.n59 25.5611
R77 minus.n20 minus.n19 24.1005
R78 minus.n19 minus.n18 24.1005
R79 minus.n53 minus.n52 24.1005
R80 minus.n54 minus.n53 24.1005
R81 minus.n12 minus.n7 22.6399
R82 minus.n26 minus.n1 22.6399
R83 minus.n46 minus.n41 22.6399
R84 minus.n60 minus.n35 22.6399
R85 minus.n9 minus.n8 14.1472
R86 minus.n43 minus.n42 14.1472
R87 minus.n68 minus.n67 6.52702
R88 minus.n31 minus.n30 2.19141
R89 minus.n65 minus.n64 2.19141
R90 minus.n14 minus.n5 0.730803
R91 minus.n24 minus.n3 0.730803
R92 minus.n48 minus.n39 0.730803
R93 minus.n58 minus.n37 0.730803
R94 minus.n33 minus.n0 0.189894
R95 minus.n29 minus.n0 0.189894
R96 minus.n29 minus.n28 0.189894
R97 minus.n28 minus.n27 0.189894
R98 minus.n27 minus.n2 0.189894
R99 minus.n23 minus.n2 0.189894
R100 minus.n23 minus.n22 0.189894
R101 minus.n22 minus.n21 0.189894
R102 minus.n21 minus.n4 0.189894
R103 minus.n17 minus.n4 0.189894
R104 minus.n17 minus.n16 0.189894
R105 minus.n16 minus.n15 0.189894
R106 minus.n15 minus.n6 0.189894
R107 minus.n11 minus.n6 0.189894
R108 minus.n11 minus.n10 0.189894
R109 minus.n45 minus.n44 0.189894
R110 minus.n45 minus.n40 0.189894
R111 minus.n49 minus.n40 0.189894
R112 minus.n50 minus.n49 0.189894
R113 minus.n51 minus.n50 0.189894
R114 minus.n51 minus.n38 0.189894
R115 minus.n55 minus.n38 0.189894
R116 minus.n56 minus.n55 0.189894
R117 minus.n57 minus.n56 0.189894
R118 minus.n57 minus.n36 0.189894
R119 minus.n61 minus.n36 0.189894
R120 minus.n62 minus.n61 0.189894
R121 minus.n63 minus.n62 0.189894
R122 minus.n63 minus.n34 0.189894
R123 minus.n67 minus.n34 0.189894
R124 minus minus.n68 0.188
R125 source.n11 source.t43 51.0588
R126 source.n12 source.t14 51.0588
R127 source.n23 source.t29 51.0588
R128 source.n47 source.t11 51.0586
R129 source.n36 source.t13 51.0586
R130 source.n35 source.t36 51.0586
R131 source.n24 source.t41 51.0586
R132 source.n0 source.t1 51.0586
R133 source.n2 source.n1 48.8588
R134 source.n4 source.n3 48.8588
R135 source.n6 source.n5 48.8588
R136 source.n8 source.n7 48.8588
R137 source.n10 source.n9 48.8588
R138 source.n14 source.n13 48.8588
R139 source.n16 source.n15 48.8588
R140 source.n18 source.n17 48.8588
R141 source.n20 source.n19 48.8588
R142 source.n22 source.n21 48.8588
R143 source.n46 source.n45 48.8586
R144 source.n44 source.n43 48.8586
R145 source.n42 source.n41 48.8586
R146 source.n40 source.n39 48.8586
R147 source.n38 source.n37 48.8586
R148 source.n34 source.n33 48.8586
R149 source.n32 source.n31 48.8586
R150 source.n30 source.n29 48.8586
R151 source.n28 source.n27 48.8586
R152 source.n26 source.n25 48.8586
R153 source.n24 source.n23 19.7305
R154 source.n48 source.n0 14.1098
R155 source.n48 source.n47 5.62119
R156 source.n45 source.t33 2.2005
R157 source.n45 source.t34 2.2005
R158 source.n43 source.t22 2.2005
R159 source.n43 source.t28 2.2005
R160 source.n41 source.t31 2.2005
R161 source.n41 source.t27 2.2005
R162 source.n39 source.t24 2.2005
R163 source.n39 source.t30 2.2005
R164 source.n37 source.t16 2.2005
R165 source.n37 source.t19 2.2005
R166 source.n33 source.t37 2.2005
R167 source.n33 source.t39 2.2005
R168 source.n31 source.t44 2.2005
R169 source.n31 source.t45 2.2005
R170 source.n29 source.t35 2.2005
R171 source.n29 source.t3 2.2005
R172 source.n27 source.t46 2.2005
R173 source.n27 source.t6 2.2005
R174 source.n25 source.t4 2.2005
R175 source.n25 source.t47 2.2005
R176 source.n1 source.t38 2.2005
R177 source.n1 source.t5 2.2005
R178 source.n3 source.t10 2.2005
R179 source.n3 source.t42 2.2005
R180 source.n5 source.t40 2.2005
R181 source.n5 source.t2 2.2005
R182 source.n7 source.t0 2.2005
R183 source.n7 source.t8 2.2005
R184 source.n9 source.t9 2.2005
R185 source.n9 source.t7 2.2005
R186 source.n13 source.t18 2.2005
R187 source.n13 source.t23 2.2005
R188 source.n15 source.t32 2.2005
R189 source.n15 source.t12 2.2005
R190 source.n17 source.t26 2.2005
R191 source.n17 source.t25 2.2005
R192 source.n19 source.t15 2.2005
R193 source.n19 source.t21 2.2005
R194 source.n21 source.t17 2.2005
R195 source.n21 source.t20 2.2005
R196 source.n23 source.n22 0.716017
R197 source.n22 source.n20 0.716017
R198 source.n20 source.n18 0.716017
R199 source.n18 source.n16 0.716017
R200 source.n16 source.n14 0.716017
R201 source.n14 source.n12 0.716017
R202 source.n11 source.n10 0.716017
R203 source.n10 source.n8 0.716017
R204 source.n8 source.n6 0.716017
R205 source.n6 source.n4 0.716017
R206 source.n4 source.n2 0.716017
R207 source.n2 source.n0 0.716017
R208 source.n26 source.n24 0.716017
R209 source.n28 source.n26 0.716017
R210 source.n30 source.n28 0.716017
R211 source.n32 source.n30 0.716017
R212 source.n34 source.n32 0.716017
R213 source.n35 source.n34 0.716017
R214 source.n38 source.n36 0.716017
R215 source.n40 source.n38 0.716017
R216 source.n42 source.n40 0.716017
R217 source.n44 source.n42 0.716017
R218 source.n46 source.n44 0.716017
R219 source.n47 source.n46 0.716017
R220 source.n12 source.n11 0.470328
R221 source.n36 source.n35 0.470328
R222 source source.n48 0.188
R223 drain_right.n13 drain_right.n11 66.2529
R224 drain_right.n7 drain_right.n5 66.2529
R225 drain_right.n2 drain_right.n0 66.2529
R226 drain_right.n13 drain_right.n12 65.5376
R227 drain_right.n15 drain_right.n14 65.5376
R228 drain_right.n17 drain_right.n16 65.5376
R229 drain_right.n19 drain_right.n18 65.5376
R230 drain_right.n21 drain_right.n20 65.5376
R231 drain_right.n7 drain_right.n6 65.5373
R232 drain_right.n9 drain_right.n8 65.5373
R233 drain_right.n4 drain_right.n3 65.5373
R234 drain_right.n2 drain_right.n1 65.5373
R235 drain_right drain_right.n10 31.3385
R236 drain_right drain_right.n21 6.36873
R237 drain_right.n5 drain_right.t15 2.2005
R238 drain_right.n5 drain_right.t3 2.2005
R239 drain_right.n6 drain_right.t4 2.2005
R240 drain_right.n6 drain_right.t9 2.2005
R241 drain_right.n8 drain_right.t13 2.2005
R242 drain_right.n8 drain_right.t20 2.2005
R243 drain_right.n3 drain_right.t22 2.2005
R244 drain_right.n3 drain_right.t12 2.2005
R245 drain_right.n1 drain_right.t14 2.2005
R246 drain_right.n1 drain_right.t17 2.2005
R247 drain_right.n0 drain_right.t0 2.2005
R248 drain_right.n0 drain_right.t1 2.2005
R249 drain_right.n11 drain_right.t21 2.2005
R250 drain_right.n11 drain_right.t8 2.2005
R251 drain_right.n12 drain_right.t5 2.2005
R252 drain_right.n12 drain_right.t16 2.2005
R253 drain_right.n14 drain_right.t11 2.2005
R254 drain_right.n14 drain_right.t18 2.2005
R255 drain_right.n16 drain_right.t10 2.2005
R256 drain_right.n16 drain_right.t23 2.2005
R257 drain_right.n18 drain_right.t19 2.2005
R258 drain_right.n18 drain_right.t6 2.2005
R259 drain_right.n20 drain_right.t2 2.2005
R260 drain_right.n20 drain_right.t7 2.2005
R261 drain_right.n9 drain_right.n7 0.716017
R262 drain_right.n4 drain_right.n2 0.716017
R263 drain_right.n21 drain_right.n19 0.716017
R264 drain_right.n19 drain_right.n17 0.716017
R265 drain_right.n17 drain_right.n15 0.716017
R266 drain_right.n15 drain_right.n13 0.716017
R267 drain_right.n10 drain_right.n9 0.302913
R268 drain_right.n10 drain_right.n4 0.302913
R269 plus.n11 plus.t5 538.725
R270 plus.n45 plus.t14 538.725
R271 plus.n32 plus.t0 512.366
R272 plus.n30 plus.t1 512.366
R273 plus.n29 plus.t12 512.366
R274 plus.n3 plus.t4 512.366
R275 plus.n23 plus.t20 512.366
R276 plus.n22 plus.t10 512.366
R277 plus.n6 plus.t23 512.366
R278 plus.n17 plus.t17 512.366
R279 plus.n15 plus.t9 512.366
R280 plus.n9 plus.t21 512.366
R281 plus.n10 plus.t13 512.366
R282 plus.n66 plus.t11 512.366
R283 plus.n64 plus.t22 512.366
R284 plus.n63 plus.t7 512.366
R285 plus.n37 plus.t6 512.366
R286 plus.n57 plus.t16 512.366
R287 plus.n56 plus.t2 512.366
R288 plus.n40 plus.t8 512.366
R289 plus.n51 plus.t19 512.366
R290 plus.n49 plus.t18 512.366
R291 plus.n43 plus.t3 512.366
R292 plus.n44 plus.t15 512.366
R293 plus.n12 plus.n9 161.3
R294 plus.n14 plus.n13 161.3
R295 plus.n15 plus.n8 161.3
R296 plus.n16 plus.n7 161.3
R297 plus.n18 plus.n17 161.3
R298 plus.n19 plus.n6 161.3
R299 plus.n21 plus.n20 161.3
R300 plus.n22 plus.n5 161.3
R301 plus.n23 plus.n4 161.3
R302 plus.n25 plus.n24 161.3
R303 plus.n26 plus.n3 161.3
R304 plus.n28 plus.n27 161.3
R305 plus.n29 plus.n2 161.3
R306 plus.n30 plus.n1 161.3
R307 plus.n31 plus.n0 161.3
R308 plus.n33 plus.n32 161.3
R309 plus.n46 plus.n43 161.3
R310 plus.n48 plus.n47 161.3
R311 plus.n49 plus.n42 161.3
R312 plus.n50 plus.n41 161.3
R313 plus.n52 plus.n51 161.3
R314 plus.n53 plus.n40 161.3
R315 plus.n55 plus.n54 161.3
R316 plus.n56 plus.n39 161.3
R317 plus.n57 plus.n38 161.3
R318 plus.n59 plus.n58 161.3
R319 plus.n60 plus.n37 161.3
R320 plus.n62 plus.n61 161.3
R321 plus.n63 plus.n36 161.3
R322 plus.n64 plus.n35 161.3
R323 plus.n65 plus.n34 161.3
R324 plus.n67 plus.n66 161.3
R325 plus.n30 plus.n29 48.2005
R326 plus.n23 plus.n22 48.2005
R327 plus.n17 plus.n6 48.2005
R328 plus.n10 plus.n9 48.2005
R329 plus.n64 plus.n63 48.2005
R330 plus.n57 plus.n56 48.2005
R331 plus.n51 plus.n40 48.2005
R332 plus.n44 plus.n43 48.2005
R333 plus.n24 plus.n3 47.4702
R334 plus.n16 plus.n15 47.4702
R335 plus.n58 plus.n37 47.4702
R336 plus.n50 plus.n49 47.4702
R337 plus.n32 plus.n31 46.0096
R338 plus.n66 plus.n65 46.0096
R339 plus.n12 plus.n11 45.0871
R340 plus.n46 plus.n45 45.0871
R341 plus plus.n67 32.7793
R342 plus.n28 plus.n3 25.5611
R343 plus.n15 plus.n14 25.5611
R344 plus.n62 plus.n37 25.5611
R345 plus.n49 plus.n48 25.5611
R346 plus.n21 plus.n6 24.1005
R347 plus.n22 plus.n21 24.1005
R348 plus.n56 plus.n55 24.1005
R349 plus.n55 plus.n40 24.1005
R350 plus.n29 plus.n28 22.6399
R351 plus.n14 plus.n9 22.6399
R352 plus.n63 plus.n62 22.6399
R353 plus.n48 plus.n43 22.6399
R354 plus.n11 plus.n10 14.1472
R355 plus.n45 plus.n44 14.1472
R356 plus plus.n33 11.0346
R357 plus.n31 plus.n30 2.19141
R358 plus.n65 plus.n64 2.19141
R359 plus.n24 plus.n23 0.730803
R360 plus.n17 plus.n16 0.730803
R361 plus.n58 plus.n57 0.730803
R362 plus.n51 plus.n50 0.730803
R363 plus.n13 plus.n12 0.189894
R364 plus.n13 plus.n8 0.189894
R365 plus.n8 plus.n7 0.189894
R366 plus.n18 plus.n7 0.189894
R367 plus.n19 plus.n18 0.189894
R368 plus.n20 plus.n19 0.189894
R369 plus.n20 plus.n5 0.189894
R370 plus.n5 plus.n4 0.189894
R371 plus.n25 plus.n4 0.189894
R372 plus.n26 plus.n25 0.189894
R373 plus.n27 plus.n26 0.189894
R374 plus.n27 plus.n2 0.189894
R375 plus.n2 plus.n1 0.189894
R376 plus.n1 plus.n0 0.189894
R377 plus.n33 plus.n0 0.189894
R378 plus.n67 plus.n34 0.189894
R379 plus.n35 plus.n34 0.189894
R380 plus.n36 plus.n35 0.189894
R381 plus.n61 plus.n36 0.189894
R382 plus.n61 plus.n60 0.189894
R383 plus.n60 plus.n59 0.189894
R384 plus.n59 plus.n38 0.189894
R385 plus.n39 plus.n38 0.189894
R386 plus.n54 plus.n39 0.189894
R387 plus.n54 plus.n53 0.189894
R388 plus.n53 plus.n52 0.189894
R389 plus.n52 plus.n41 0.189894
R390 plus.n42 plus.n41 0.189894
R391 plus.n47 plus.n42 0.189894
R392 plus.n47 plus.n46 0.189894
R393 drain_left.n13 drain_left.n11 66.2531
R394 drain_left.n7 drain_left.n5 66.2529
R395 drain_left.n2 drain_left.n0 66.2529
R396 drain_left.n19 drain_left.n18 65.5376
R397 drain_left.n17 drain_left.n16 65.5376
R398 drain_left.n15 drain_left.n14 65.5376
R399 drain_left.n13 drain_left.n12 65.5376
R400 drain_left.n21 drain_left.n20 65.5374
R401 drain_left.n7 drain_left.n6 65.5373
R402 drain_left.n9 drain_left.n8 65.5373
R403 drain_left.n4 drain_left.n3 65.5373
R404 drain_left.n2 drain_left.n1 65.5373
R405 drain_left drain_left.n10 31.8918
R406 drain_left drain_left.n21 6.36873
R407 drain_left.n5 drain_left.t8 2.2005
R408 drain_left.n5 drain_left.t9 2.2005
R409 drain_left.n6 drain_left.t5 2.2005
R410 drain_left.n6 drain_left.t20 2.2005
R411 drain_left.n8 drain_left.t15 2.2005
R412 drain_left.n8 drain_left.t4 2.2005
R413 drain_left.n3 drain_left.t7 2.2005
R414 drain_left.n3 drain_left.t21 2.2005
R415 drain_left.n1 drain_left.t16 2.2005
R416 drain_left.n1 drain_left.t17 2.2005
R417 drain_left.n0 drain_left.t12 2.2005
R418 drain_left.n0 drain_left.t1 2.2005
R419 drain_left.n20 drain_left.t22 2.2005
R420 drain_left.n20 drain_left.t23 2.2005
R421 drain_left.n18 drain_left.t19 2.2005
R422 drain_left.n18 drain_left.t11 2.2005
R423 drain_left.n16 drain_left.t13 2.2005
R424 drain_left.n16 drain_left.t3 2.2005
R425 drain_left.n14 drain_left.t6 2.2005
R426 drain_left.n14 drain_left.t0 2.2005
R427 drain_left.n12 drain_left.t2 2.2005
R428 drain_left.n12 drain_left.t14 2.2005
R429 drain_left.n11 drain_left.t18 2.2005
R430 drain_left.n11 drain_left.t10 2.2005
R431 drain_left.n9 drain_left.n7 0.716017
R432 drain_left.n4 drain_left.n2 0.716017
R433 drain_left.n15 drain_left.n13 0.716017
R434 drain_left.n17 drain_left.n15 0.716017
R435 drain_left.n19 drain_left.n17 0.716017
R436 drain_left.n21 drain_left.n19 0.716017
R437 drain_left.n10 drain_left.n9 0.302913
R438 drain_left.n10 drain_left.n4 0.302913
C0 drain_left drain_right 1.55979f
C1 minus drain_right 9.2836f
C2 source drain_right 26.5441f
C3 plus drain_left 9.56992f
C4 minus plus 6.18598f
C5 plus source 9.471821f
C6 minus drain_left 0.173624f
C7 source drain_left 26.542599f
C8 minus source 9.45778f
C9 plus drain_right 0.443411f
C10 drain_right a_n2874_n2688# 6.93073f
C11 drain_left a_n2874_n2688# 7.34347f
C12 source a_n2874_n2688# 7.63688f
C13 minus a_n2874_n2688# 11.318554f
C14 plus a_n2874_n2688# 13.126781f
C15 drain_left.t12 a_n2874_n2688# 0.209323f
C16 drain_left.t1 a_n2874_n2688# 0.209323f
C17 drain_left.n0 a_n2874_n2688# 1.83502f
C18 drain_left.t16 a_n2874_n2688# 0.209323f
C19 drain_left.t17 a_n2874_n2688# 0.209323f
C20 drain_left.n1 a_n2874_n2688# 1.83088f
C21 drain_left.n2 a_n2874_n2688# 0.750653f
C22 drain_left.t7 a_n2874_n2688# 0.209323f
C23 drain_left.t21 a_n2874_n2688# 0.209323f
C24 drain_left.n3 a_n2874_n2688# 1.83088f
C25 drain_left.n4 a_n2874_n2688# 0.334548f
C26 drain_left.t8 a_n2874_n2688# 0.209323f
C27 drain_left.t9 a_n2874_n2688# 0.209323f
C28 drain_left.n5 a_n2874_n2688# 1.83502f
C29 drain_left.t5 a_n2874_n2688# 0.209323f
C30 drain_left.t20 a_n2874_n2688# 0.209323f
C31 drain_left.n6 a_n2874_n2688# 1.83088f
C32 drain_left.n7 a_n2874_n2688# 0.750653f
C33 drain_left.t15 a_n2874_n2688# 0.209323f
C34 drain_left.t4 a_n2874_n2688# 0.209323f
C35 drain_left.n8 a_n2874_n2688# 1.83088f
C36 drain_left.n9 a_n2874_n2688# 0.334548f
C37 drain_left.n10 a_n2874_n2688# 1.56935f
C38 drain_left.t18 a_n2874_n2688# 0.209323f
C39 drain_left.t10 a_n2874_n2688# 0.209323f
C40 drain_left.n11 a_n2874_n2688# 1.83502f
C41 drain_left.t2 a_n2874_n2688# 0.209323f
C42 drain_left.t14 a_n2874_n2688# 0.209323f
C43 drain_left.n12 a_n2874_n2688# 1.83088f
C44 drain_left.n13 a_n2874_n2688# 0.750646f
C45 drain_left.t6 a_n2874_n2688# 0.209323f
C46 drain_left.t0 a_n2874_n2688# 0.209323f
C47 drain_left.n14 a_n2874_n2688# 1.83088f
C48 drain_left.n15 a_n2874_n2688# 0.371465f
C49 drain_left.t13 a_n2874_n2688# 0.209323f
C50 drain_left.t3 a_n2874_n2688# 0.209323f
C51 drain_left.n16 a_n2874_n2688# 1.83088f
C52 drain_left.n17 a_n2874_n2688# 0.371465f
C53 drain_left.t19 a_n2874_n2688# 0.209323f
C54 drain_left.t11 a_n2874_n2688# 0.209323f
C55 drain_left.n18 a_n2874_n2688# 1.83088f
C56 drain_left.n19 a_n2874_n2688# 0.371465f
C57 drain_left.t22 a_n2874_n2688# 0.209323f
C58 drain_left.t23 a_n2874_n2688# 0.209323f
C59 drain_left.n20 a_n2874_n2688# 1.83087f
C60 drain_left.n21 a_n2874_n2688# 0.624336f
C61 plus.n0 a_n2874_n2688# 0.044314f
C62 plus.t0 a_n2874_n2688# 0.571887f
C63 plus.t1 a_n2874_n2688# 0.571887f
C64 plus.n1 a_n2874_n2688# 0.044314f
C65 plus.t12 a_n2874_n2688# 0.571887f
C66 plus.n2 a_n2874_n2688# 0.044314f
C67 plus.t4 a_n2874_n2688# 0.571887f
C68 plus.n3 a_n2874_n2688# 0.248381f
C69 plus.n4 a_n2874_n2688# 0.044314f
C70 plus.t20 a_n2874_n2688# 0.571887f
C71 plus.t10 a_n2874_n2688# 0.571887f
C72 plus.n5 a_n2874_n2688# 0.044314f
C73 plus.t23 a_n2874_n2688# 0.571887f
C74 plus.n6 a_n2874_n2688# 0.248245f
C75 plus.n7 a_n2874_n2688# 0.044314f
C76 plus.t17 a_n2874_n2688# 0.571887f
C77 plus.t9 a_n2874_n2688# 0.571887f
C78 plus.n8 a_n2874_n2688# 0.044314f
C79 plus.t21 a_n2874_n2688# 0.571887f
C80 plus.n9 a_n2874_n2688# 0.247971f
C81 plus.t13 a_n2874_n2688# 0.571887f
C82 plus.n10 a_n2874_n2688# 0.253215f
C83 plus.t5 a_n2874_n2688# 0.583809f
C84 plus.n11 a_n2874_n2688# 0.233266f
C85 plus.n12 a_n2874_n2688# 0.179933f
C86 plus.n13 a_n2874_n2688# 0.044314f
C87 plus.n14 a_n2874_n2688# 0.010056f
C88 plus.n15 a_n2874_n2688# 0.248381f
C89 plus.n16 a_n2874_n2688# 0.010056f
C90 plus.n17 a_n2874_n2688# 0.243873f
C91 plus.n18 a_n2874_n2688# 0.044314f
C92 plus.n19 a_n2874_n2688# 0.044314f
C93 plus.n20 a_n2874_n2688# 0.044314f
C94 plus.n21 a_n2874_n2688# 0.010056f
C95 plus.n22 a_n2874_n2688# 0.248245f
C96 plus.n23 a_n2874_n2688# 0.243873f
C97 plus.n24 a_n2874_n2688# 0.010056f
C98 plus.n25 a_n2874_n2688# 0.044314f
C99 plus.n26 a_n2874_n2688# 0.044314f
C100 plus.n27 a_n2874_n2688# 0.044314f
C101 plus.n28 a_n2874_n2688# 0.010056f
C102 plus.n29 a_n2874_n2688# 0.247971f
C103 plus.n30 a_n2874_n2688# 0.244146f
C104 plus.n31 a_n2874_n2688# 0.010056f
C105 plus.n32 a_n2874_n2688# 0.243327f
C106 plus.n33 a_n2874_n2688# 0.438196f
C107 plus.n34 a_n2874_n2688# 0.044314f
C108 plus.t11 a_n2874_n2688# 0.571887f
C109 plus.n35 a_n2874_n2688# 0.044314f
C110 plus.t22 a_n2874_n2688# 0.571887f
C111 plus.n36 a_n2874_n2688# 0.044314f
C112 plus.t7 a_n2874_n2688# 0.571887f
C113 plus.t6 a_n2874_n2688# 0.571887f
C114 plus.n37 a_n2874_n2688# 0.248381f
C115 plus.n38 a_n2874_n2688# 0.044314f
C116 plus.t16 a_n2874_n2688# 0.571887f
C117 plus.n39 a_n2874_n2688# 0.044314f
C118 plus.t2 a_n2874_n2688# 0.571887f
C119 plus.t8 a_n2874_n2688# 0.571887f
C120 plus.n40 a_n2874_n2688# 0.248245f
C121 plus.n41 a_n2874_n2688# 0.044314f
C122 plus.t19 a_n2874_n2688# 0.571887f
C123 plus.n42 a_n2874_n2688# 0.044314f
C124 plus.t18 a_n2874_n2688# 0.571887f
C125 plus.t3 a_n2874_n2688# 0.571887f
C126 plus.n43 a_n2874_n2688# 0.247971f
C127 plus.t14 a_n2874_n2688# 0.583809f
C128 plus.t15 a_n2874_n2688# 0.571887f
C129 plus.n44 a_n2874_n2688# 0.253215f
C130 plus.n45 a_n2874_n2688# 0.233266f
C131 plus.n46 a_n2874_n2688# 0.179933f
C132 plus.n47 a_n2874_n2688# 0.044314f
C133 plus.n48 a_n2874_n2688# 0.010056f
C134 plus.n49 a_n2874_n2688# 0.248381f
C135 plus.n50 a_n2874_n2688# 0.010056f
C136 plus.n51 a_n2874_n2688# 0.243873f
C137 plus.n52 a_n2874_n2688# 0.044314f
C138 plus.n53 a_n2874_n2688# 0.044314f
C139 plus.n54 a_n2874_n2688# 0.044314f
C140 plus.n55 a_n2874_n2688# 0.010056f
C141 plus.n56 a_n2874_n2688# 0.248245f
C142 plus.n57 a_n2874_n2688# 0.243873f
C143 plus.n58 a_n2874_n2688# 0.010056f
C144 plus.n59 a_n2874_n2688# 0.044314f
C145 plus.n60 a_n2874_n2688# 0.044314f
C146 plus.n61 a_n2874_n2688# 0.044314f
C147 plus.n62 a_n2874_n2688# 0.010056f
C148 plus.n63 a_n2874_n2688# 0.247971f
C149 plus.n64 a_n2874_n2688# 0.244146f
C150 plus.n65 a_n2874_n2688# 0.010056f
C151 plus.n66 a_n2874_n2688# 0.243327f
C152 plus.n67 a_n2874_n2688# 1.46929f
C153 drain_right.t0 a_n2874_n2688# 0.208248f
C154 drain_right.t1 a_n2874_n2688# 0.208248f
C155 drain_right.n0 a_n2874_n2688# 1.82559f
C156 drain_right.t14 a_n2874_n2688# 0.208248f
C157 drain_right.t17 a_n2874_n2688# 0.208248f
C158 drain_right.n1 a_n2874_n2688# 1.82147f
C159 drain_right.n2 a_n2874_n2688# 0.746796f
C160 drain_right.t22 a_n2874_n2688# 0.208248f
C161 drain_right.t12 a_n2874_n2688# 0.208248f
C162 drain_right.n3 a_n2874_n2688# 1.82147f
C163 drain_right.n4 a_n2874_n2688# 0.332829f
C164 drain_right.t15 a_n2874_n2688# 0.208248f
C165 drain_right.t3 a_n2874_n2688# 0.208248f
C166 drain_right.n5 a_n2874_n2688# 1.82559f
C167 drain_right.t4 a_n2874_n2688# 0.208248f
C168 drain_right.t9 a_n2874_n2688# 0.208248f
C169 drain_right.n6 a_n2874_n2688# 1.82147f
C170 drain_right.n7 a_n2874_n2688# 0.746796f
C171 drain_right.t13 a_n2874_n2688# 0.208248f
C172 drain_right.t20 a_n2874_n2688# 0.208248f
C173 drain_right.n8 a_n2874_n2688# 1.82147f
C174 drain_right.n9 a_n2874_n2688# 0.332829f
C175 drain_right.n10 a_n2874_n2688# 1.50202f
C176 drain_right.t21 a_n2874_n2688# 0.208248f
C177 drain_right.t8 a_n2874_n2688# 0.208248f
C178 drain_right.n11 a_n2874_n2688# 1.82559f
C179 drain_right.t5 a_n2874_n2688# 0.208248f
C180 drain_right.t16 a_n2874_n2688# 0.208248f
C181 drain_right.n12 a_n2874_n2688# 1.82148f
C182 drain_right.n13 a_n2874_n2688# 0.746797f
C183 drain_right.t11 a_n2874_n2688# 0.208248f
C184 drain_right.t18 a_n2874_n2688# 0.208248f
C185 drain_right.n14 a_n2874_n2688# 1.82148f
C186 drain_right.n15 a_n2874_n2688# 0.369557f
C187 drain_right.t10 a_n2874_n2688# 0.208248f
C188 drain_right.t23 a_n2874_n2688# 0.208248f
C189 drain_right.n16 a_n2874_n2688# 1.82148f
C190 drain_right.n17 a_n2874_n2688# 0.369557f
C191 drain_right.t19 a_n2874_n2688# 0.208248f
C192 drain_right.t6 a_n2874_n2688# 0.208248f
C193 drain_right.n18 a_n2874_n2688# 1.82148f
C194 drain_right.n19 a_n2874_n2688# 0.369557f
C195 drain_right.t2 a_n2874_n2688# 0.208248f
C196 drain_right.t7 a_n2874_n2688# 0.208248f
C197 drain_right.n20 a_n2874_n2688# 1.82148f
C198 drain_right.n21 a_n2874_n2688# 0.621121f
C199 source.t1 a_n2874_n2688# 2.04901f
C200 source.n0 a_n2874_n2688# 1.20335f
C201 source.t38 a_n2874_n2688# 0.192152f
C202 source.t5 a_n2874_n2688# 0.192152f
C203 source.n1 a_n2874_n2688# 1.60857f
C204 source.n2 a_n2874_n2688# 0.376392f
C205 source.t10 a_n2874_n2688# 0.192152f
C206 source.t42 a_n2874_n2688# 0.192152f
C207 source.n3 a_n2874_n2688# 1.60857f
C208 source.n4 a_n2874_n2688# 0.376392f
C209 source.t40 a_n2874_n2688# 0.192152f
C210 source.t2 a_n2874_n2688# 0.192152f
C211 source.n5 a_n2874_n2688# 1.60857f
C212 source.n6 a_n2874_n2688# 0.376392f
C213 source.t0 a_n2874_n2688# 0.192152f
C214 source.t8 a_n2874_n2688# 0.192152f
C215 source.n7 a_n2874_n2688# 1.60857f
C216 source.n8 a_n2874_n2688# 0.376392f
C217 source.t9 a_n2874_n2688# 0.192152f
C218 source.t7 a_n2874_n2688# 0.192152f
C219 source.n9 a_n2874_n2688# 1.60857f
C220 source.n10 a_n2874_n2688# 0.376392f
C221 source.t43 a_n2874_n2688# 2.04902f
C222 source.n11 a_n2874_n2688# 0.438614f
C223 source.t14 a_n2874_n2688# 2.04902f
C224 source.n12 a_n2874_n2688# 0.438614f
C225 source.t18 a_n2874_n2688# 0.192152f
C226 source.t23 a_n2874_n2688# 0.192152f
C227 source.n13 a_n2874_n2688# 1.60857f
C228 source.n14 a_n2874_n2688# 0.376392f
C229 source.t32 a_n2874_n2688# 0.192152f
C230 source.t12 a_n2874_n2688# 0.192152f
C231 source.n15 a_n2874_n2688# 1.60857f
C232 source.n16 a_n2874_n2688# 0.376392f
C233 source.t26 a_n2874_n2688# 0.192152f
C234 source.t25 a_n2874_n2688# 0.192152f
C235 source.n17 a_n2874_n2688# 1.60857f
C236 source.n18 a_n2874_n2688# 0.376392f
C237 source.t15 a_n2874_n2688# 0.192152f
C238 source.t21 a_n2874_n2688# 0.192152f
C239 source.n19 a_n2874_n2688# 1.60857f
C240 source.n20 a_n2874_n2688# 0.376392f
C241 source.t17 a_n2874_n2688# 0.192152f
C242 source.t20 a_n2874_n2688# 0.192152f
C243 source.n21 a_n2874_n2688# 1.60857f
C244 source.n22 a_n2874_n2688# 0.376392f
C245 source.t29 a_n2874_n2688# 2.04902f
C246 source.n23 a_n2874_n2688# 1.60082f
C247 source.t41 a_n2874_n2688# 2.04901f
C248 source.n24 a_n2874_n2688# 1.60082f
C249 source.t4 a_n2874_n2688# 0.192152f
C250 source.t47 a_n2874_n2688# 0.192152f
C251 source.n25 a_n2874_n2688# 1.60857f
C252 source.n26 a_n2874_n2688# 0.376397f
C253 source.t46 a_n2874_n2688# 0.192152f
C254 source.t6 a_n2874_n2688# 0.192152f
C255 source.n27 a_n2874_n2688# 1.60857f
C256 source.n28 a_n2874_n2688# 0.376397f
C257 source.t35 a_n2874_n2688# 0.192152f
C258 source.t3 a_n2874_n2688# 0.192152f
C259 source.n29 a_n2874_n2688# 1.60857f
C260 source.n30 a_n2874_n2688# 0.376397f
C261 source.t44 a_n2874_n2688# 0.192152f
C262 source.t45 a_n2874_n2688# 0.192152f
C263 source.n31 a_n2874_n2688# 1.60857f
C264 source.n32 a_n2874_n2688# 0.376397f
C265 source.t37 a_n2874_n2688# 0.192152f
C266 source.t39 a_n2874_n2688# 0.192152f
C267 source.n33 a_n2874_n2688# 1.60857f
C268 source.n34 a_n2874_n2688# 0.376397f
C269 source.t36 a_n2874_n2688# 2.04901f
C270 source.n35 a_n2874_n2688# 0.438619f
C271 source.t13 a_n2874_n2688# 2.04901f
C272 source.n36 a_n2874_n2688# 0.438619f
C273 source.t16 a_n2874_n2688# 0.192152f
C274 source.t19 a_n2874_n2688# 0.192152f
C275 source.n37 a_n2874_n2688# 1.60857f
C276 source.n38 a_n2874_n2688# 0.376397f
C277 source.t24 a_n2874_n2688# 0.192152f
C278 source.t30 a_n2874_n2688# 0.192152f
C279 source.n39 a_n2874_n2688# 1.60857f
C280 source.n40 a_n2874_n2688# 0.376397f
C281 source.t31 a_n2874_n2688# 0.192152f
C282 source.t27 a_n2874_n2688# 0.192152f
C283 source.n41 a_n2874_n2688# 1.60857f
C284 source.n42 a_n2874_n2688# 0.376397f
C285 source.t22 a_n2874_n2688# 0.192152f
C286 source.t28 a_n2874_n2688# 0.192152f
C287 source.n43 a_n2874_n2688# 1.60857f
C288 source.n44 a_n2874_n2688# 0.376397f
C289 source.t33 a_n2874_n2688# 0.192152f
C290 source.t34 a_n2874_n2688# 0.192152f
C291 source.n45 a_n2874_n2688# 1.60857f
C292 source.n46 a_n2874_n2688# 0.376397f
C293 source.t11 a_n2874_n2688# 2.04901f
C294 source.n47 a_n2874_n2688# 0.603063f
C295 source.n48 a_n2874_n2688# 1.41445f
C296 minus.n0 a_n2874_n2688# 0.043634f
C297 minus.t4 a_n2874_n2688# 0.563111f
C298 minus.n1 a_n2874_n2688# 0.244166f
C299 minus.t16 a_n2874_n2688# 0.563111f
C300 minus.n2 a_n2874_n2688# 0.043634f
C301 minus.t13 a_n2874_n2688# 0.563111f
C302 minus.n3 a_n2874_n2688# 0.240131f
C303 minus.n4 a_n2874_n2688# 0.043634f
C304 minus.t5 a_n2874_n2688# 0.563111f
C305 minus.n5 a_n2874_n2688# 0.240131f
C306 minus.t12 a_n2874_n2688# 0.563111f
C307 minus.n6 a_n2874_n2688# 0.043634f
C308 minus.t7 a_n2874_n2688# 0.563111f
C309 minus.n7 a_n2874_n2688# 0.244166f
C310 minus.t15 a_n2874_n2688# 0.57485f
C311 minus.t2 a_n2874_n2688# 0.563111f
C312 minus.n8 a_n2874_n2688# 0.249329f
C313 minus.n9 a_n2874_n2688# 0.229687f
C314 minus.n10 a_n2874_n2688# 0.177172f
C315 minus.n11 a_n2874_n2688# 0.043634f
C316 minus.n12 a_n2874_n2688# 0.009901f
C317 minus.t18 a_n2874_n2688# 0.563111f
C318 minus.n13 a_n2874_n2688# 0.24457f
C319 minus.n14 a_n2874_n2688# 0.009901f
C320 minus.n15 a_n2874_n2688# 0.043634f
C321 minus.n16 a_n2874_n2688# 0.043634f
C322 minus.n17 a_n2874_n2688# 0.043634f
C323 minus.n18 a_n2874_n2688# 0.244435f
C324 minus.n19 a_n2874_n2688# 0.009901f
C325 minus.t0 a_n2874_n2688# 0.563111f
C326 minus.n20 a_n2874_n2688# 0.244435f
C327 minus.n21 a_n2874_n2688# 0.043634f
C328 minus.n22 a_n2874_n2688# 0.043634f
C329 minus.n23 a_n2874_n2688# 0.043634f
C330 minus.n24 a_n2874_n2688# 0.009901f
C331 minus.t17 a_n2874_n2688# 0.563111f
C332 minus.n25 a_n2874_n2688# 0.24457f
C333 minus.n26 a_n2874_n2688# 0.009901f
C334 minus.n27 a_n2874_n2688# 0.043634f
C335 minus.n28 a_n2874_n2688# 0.043634f
C336 minus.n29 a_n2874_n2688# 0.043634f
C337 minus.n30 a_n2874_n2688# 0.2404f
C338 minus.n31 a_n2874_n2688# 0.009901f
C339 minus.t21 a_n2874_n2688# 0.563111f
C340 minus.n32 a_n2874_n2688# 0.239593f
C341 minus.n33 a_n2874_n2688# 1.64768f
C342 minus.n34 a_n2874_n2688# 0.043634f
C343 minus.t14 a_n2874_n2688# 0.563111f
C344 minus.n35 a_n2874_n2688# 0.244166f
C345 minus.n36 a_n2874_n2688# 0.043634f
C346 minus.t3 a_n2874_n2688# 0.563111f
C347 minus.n37 a_n2874_n2688# 0.240131f
C348 minus.n38 a_n2874_n2688# 0.043634f
C349 minus.t1 a_n2874_n2688# 0.563111f
C350 minus.n39 a_n2874_n2688# 0.240131f
C351 minus.n40 a_n2874_n2688# 0.043634f
C352 minus.t9 a_n2874_n2688# 0.563111f
C353 minus.n41 a_n2874_n2688# 0.244166f
C354 minus.t23 a_n2874_n2688# 0.57485f
C355 minus.t22 a_n2874_n2688# 0.563111f
C356 minus.n42 a_n2874_n2688# 0.249329f
C357 minus.n43 a_n2874_n2688# 0.229687f
C358 minus.n44 a_n2874_n2688# 0.177172f
C359 minus.n45 a_n2874_n2688# 0.043634f
C360 minus.n46 a_n2874_n2688# 0.009901f
C361 minus.t6 a_n2874_n2688# 0.563111f
C362 minus.n47 a_n2874_n2688# 0.24457f
C363 minus.n48 a_n2874_n2688# 0.009901f
C364 minus.n49 a_n2874_n2688# 0.043634f
C365 minus.n50 a_n2874_n2688# 0.043634f
C366 minus.n51 a_n2874_n2688# 0.043634f
C367 minus.t11 a_n2874_n2688# 0.563111f
C368 minus.n52 a_n2874_n2688# 0.244435f
C369 minus.n53 a_n2874_n2688# 0.009901f
C370 minus.t10 a_n2874_n2688# 0.563111f
C371 minus.n54 a_n2874_n2688# 0.244435f
C372 minus.n55 a_n2874_n2688# 0.043634f
C373 minus.n56 a_n2874_n2688# 0.043634f
C374 minus.n57 a_n2874_n2688# 0.043634f
C375 minus.n58 a_n2874_n2688# 0.009901f
C376 minus.t19 a_n2874_n2688# 0.563111f
C377 minus.n59 a_n2874_n2688# 0.24457f
C378 minus.n60 a_n2874_n2688# 0.009901f
C379 minus.n61 a_n2874_n2688# 0.043634f
C380 minus.n62 a_n2874_n2688# 0.043634f
C381 minus.n63 a_n2874_n2688# 0.043634f
C382 minus.t8 a_n2874_n2688# 0.563111f
C383 minus.n64 a_n2874_n2688# 0.2404f
C384 minus.n65 a_n2874_n2688# 0.009901f
C385 minus.t20 a_n2874_n2688# 0.563111f
C386 minus.n66 a_n2874_n2688# 0.239593f
C387 minus.n67 a_n2874_n2688# 0.28804f
C388 minus.n68 a_n2874_n2688# 1.99135f
.ends

