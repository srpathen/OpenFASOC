* NGSPICE file created from opamp233.ext - technology: sky130A

.subckt opamp233 gnd CSoutput output vdd plus minus commonsourceibias outputibias
+ diffpairibias
X0 CSoutput.t158 a_n6972_8799.t40 vdd.t233 vdd.t199 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X1 a_n6972_8799.t3 plus.t5 a_n2903_n3924.t41 gnd.t53 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.7
X2 a_n2140_13878.t15 a_n2408_n452.t24 a_n2408_n452.t25 vdd.t2 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X3 CSoutput.t39 commonsourceibias.t80 gnd.t142 gnd.t141 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X4 a_n2140_13878.t23 a_n2408_n452.t56 vdd.t235 vdd.t234 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X5 gnd.t401 gnd.t399 gnd.t400 gnd.t349 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=0 ps=0 w=7 l=0.7
X6 vdd.t232 a_n6972_8799.t41 CSoutput.t157 vdd.t140 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X7 vdd.t106 vdd.t104 vdd.t105 vdd.t48 sky130_fd_pr__pfet_01v8 ad=3.12 pd=16.78 as=0 ps=0 w=8 l=0.5
X8 gnd.t146 commonsourceibias.t81 CSoutput.t41 gnd.t103 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X9 gnd.t398 gnd.t396 minus.t4 gnd.t397 sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.5
X10 CSoutput.t47 commonsourceibias.t82 gnd.t159 gnd.t20 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X11 CSoutput.t165 commonsourceibias.t83 gnd.t239 gnd.t184 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X12 CSoutput.t156 a_n6972_8799.t42 vdd.t231 vdd.t146 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X13 a_n2903_n3924.t40 plus.t6 a_n6972_8799.t28 gnd.t54 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.7
X14 gnd.t33 commonsourceibias.t84 CSoutput.t15 gnd.t32 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X15 CSoutput.t192 a_n2318_8322.t27 sky130_fd_pr__cap_mim_m3_1 l=12 w=12
X16 a_n2903_n3924.t17 minus.t5 a_n2408_n452.t44 gnd.t100 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.7
X17 a_n2318_8322.t23 a_n2408_n452.t57 a_n6972_8799.t39 vdd.t107 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X18 vdd.t4 CSoutput.t193 output.t15 gnd.t133 sky130_fd_pr__nfet_01v8 ad=0.825 pd=5.33 as=0.825 ps=5.33 w=5 l=1
X19 CSoutput.t155 a_n6972_8799.t43 vdd.t230 vdd.t174 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X20 CSoutput.t26 commonsourceibias.t85 gnd.t68 gnd.t67 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X21 gnd.t195 commonsourceibias.t86 CSoutput.t66 gnd.t172 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X22 CSoutput.t60 commonsourceibias.t87 gnd.t182 gnd.t165 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X23 gnd.t227 commonsourceibias.t88 CSoutput.t86 gnd.t60 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=1.155 ps=7.33 w=7 l=1
X24 vdd.t229 a_n6972_8799.t44 CSoutput.t154 vdd.t194 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X25 CSoutput.t74 commonsourceibias.t89 gnd.t204 gnd.t165 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X26 CSoutput.t14 commonsourceibias.t90 gnd.t31 gnd.t0 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X27 gnd.t5 commonsourceibias.t91 CSoutput.t2 gnd.t4 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X28 a_n2408_n452.t47 minus.t6 a_n2903_n3924.t45 gnd.t111 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.7
X29 gnd.t395 gnd.t392 gnd.t394 gnd.t393 sky130_fd_pr__nfet_01v8 ad=2.34 pd=12.78 as=0 ps=0 w=6 l=2
X30 gnd.t391 gnd.t389 gnd.t390 gnd.t308 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=0 ps=0 w=7 l=1
X31 commonsourceibias.t79 commonsourceibias.t78 gnd.t257 gnd.t67 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X32 CSoutput.t73 commonsourceibias.t92 gnd.t203 gnd.t184 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X33 gnd.t388 gnd.t386 gnd.t387 gnd.t297 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=0 ps=0 w=7 l=1
X34 a_n6972_8799.t17 a_n2408_n452.t58 a_n2318_8322.t22 vdd.t16 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=3.51 ps=18.78 w=9 l=0.5
X35 vdd.t228 a_n6972_8799.t45 CSoutput.t153 vdd.t206 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X36 a_n2408_n452.t52 minus.t7 a_n2903_n3924.t51 gnd.t110 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.7
X37 CSoutput.t152 a_n6972_8799.t46 vdd.t227 vdd.t176 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X38 a_n6972_8799.t18 a_n2408_n452.t59 a_n2318_8322.t21 vdd.t21 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=3.51 ps=18.78 w=9 l=0.5
X39 CSoutput.t178 commonsourceibias.t93 gnd.t256 gnd.t141 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X40 gnd.t278 commonsourceibias.t94 CSoutput.t189 gnd.t58 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X41 gnd.t385 gnd.t383 gnd.t384 gnd.t312 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=0 ps=0 w=7 l=1
X42 CSoutput.t59 commonsourceibias.t95 gnd.t181 gnd.t74 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X43 CSoutput.t72 commonsourceibias.t96 gnd.t202 gnd.t24 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X44 a_n2903_n3924.t47 minus.t8 a_n2408_n452.t49 gnd.t109 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=1.155 ps=7.33 w=7 l=0.7
X45 vdd.t103 vdd.t101 vdd.t102 vdd.t32 sky130_fd_pr__pfet_01v8 ad=3.51 pd=18.78 as=0 ps=0 w=9 l=0.5
X46 CSoutput.t177 commonsourceibias.t97 gnd.t255 gnd.t139 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X47 CSoutput.t151 a_n6972_8799.t47 vdd.t226 vdd.t199 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X48 CSoutput.t150 a_n6972_8799.t48 vdd.t225 vdd.t168 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=3.12 ps=16.78 w=8 l=0.5
X49 a_n2903_n3924.t48 diffpairibias.t16 gnd.t169 gnd.t168 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=2.73 ps=14.78 w=7 l=1
X50 gnd.t277 commonsourceibias.t98 CSoutput.t188 gnd.t51 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=1.155 ps=7.33 w=7 l=1
X51 gnd.t180 commonsourceibias.t99 CSoutput.t58 gnd.t105 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X52 vdd.t100 vdd.t98 vdd.t99 vdd.t48 sky130_fd_pr__pfet_01v8 ad=3.12 pd=16.78 as=0 ps=0 w=8 l=0.5
X53 CSoutput.t176 commonsourceibias.t100 gnd.t254 gnd.t43 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X54 CSoutput.t182 commonsourceibias.t101 gnd.t268 gnd.t2 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=2.73 ps=14.78 w=7 l=1
X55 gnd.t70 commonsourceibias.t76 commonsourceibias.t77 gnd.t69 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X56 CSoutput.t38 commonsourceibias.t102 gnd.t140 gnd.t139 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X57 CSoutput.t149 a_n6972_8799.t49 vdd.t224 vdd.t146 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X58 gnd.t158 commonsourceibias.t103 CSoutput.t46 gnd.t22 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X59 a_n2903_n3924.t39 plus.t7 a_n6972_8799.t12 gnd.t117 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.7
X60 a_n2140_13878.t14 a_n2408_n452.t10 a_n2408_n452.t11 vdd.t20 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X61 CSoutput.t164 commonsourceibias.t104 gnd.t238 gnd.t137 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X62 CSoutput.t13 commonsourceibias.t105 gnd.t30 gnd.t29 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X63 gnd.t66 commonsourceibias.t106 CSoutput.t25 gnd.t22 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X64 vdd.t5 CSoutput.t194 output.t14 gnd.t132 sky130_fd_pr__nfet_01v8 ad=0.825 pd=5.33 as=0.825 ps=5.33 w=5 l=1
X65 a_n6972_8799.t13 plus.t8 a_n2903_n3924.t38 gnd.t116 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=2.73 ps=14.78 w=7 l=0.7
X66 a_n2408_n452.t21 a_n2408_n452.t20 a_n2140_13878.t13 vdd.t0 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X67 CSoutput.t65 commonsourceibias.t107 gnd.t194 gnd.t39 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X68 gnd.t179 commonsourceibias.t108 CSoutput.t57 gnd.t103 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X69 CSoutput.t195 a_n2318_8322.t26 sky130_fd_pr__cap_mim_m3_1 l=12 w=12
X70 a_n6972_8799.t11 plus.t9 a_n2903_n3924.t37 gnd.t115 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.7
X71 CSoutput.t148 a_n6972_8799.t50 vdd.t223 vdd.t174 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X72 vdd.t97 vdd.t95 vdd.t96 vdd.t78 sky130_fd_pr__pfet_01v8 ad=3.51 pd=18.78 as=0 ps=0 w=9 l=0.5
X73 gnd.t183 commonsourceibias.t74 commonsourceibias.t75 gnd.t14 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X74 CSoutput.t85 commonsourceibias.t109 gnd.t226 gnd.t165 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X75 vdd.t222 a_n6972_8799.t51 CSoutput.t147 vdd.t194 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X76 gnd.t382 gnd.t380 gnd.t381 gnd.t312 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=0 ps=0 w=7 l=1
X77 CSoutput.t71 commonsourceibias.t110 gnd.t201 gnd.t29 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X78 diffpairibias.t15 diffpairibias.t14 gnd.t151 gnd.t150 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=2.73 ps=14.78 w=7 l=1
X79 a_n2903_n3924.t36 plus.t10 a_n6972_8799.t38 gnd.t91 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.7
X80 gnd.t28 commonsourceibias.t111 CSoutput.t12 gnd.t27 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X81 a_n2408_n452.t40 minus.t9 a_n2903_n3924.t11 gnd.t86 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.7
X82 CSoutput.t1 commonsourceibias.t112 gnd.t3 gnd.t2 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=2.73 ps=14.78 w=7 l=1
X83 CSoutput.t70 commonsourceibias.t113 gnd.t200 gnd.t45 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X84 gnd.t237 commonsourceibias.t114 CSoutput.t163 gnd.t101 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X85 a_n6972_8799.t5 a_n2408_n452.t60 a_n2318_8322.t20 vdd.t18 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X86 gnd.t65 commonsourceibias.t115 CSoutput.t24 gnd.t35 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X87 CSoutput.t146 a_n6972_8799.t52 vdd.t221 vdd.t196 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X88 gnd.t193 commonsourceibias.t116 CSoutput.t64 gnd.t10 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X89 gnd.t379 gnd.t377 plus.t2 gnd.t378 sky130_fd_pr__nfet_01v8 ad=0.39 pd=2.78 as=0.165 ps=1.33 w=1 l=0.5
X90 vdd.t220 a_n6972_8799.t53 CSoutput.t145 vdd.t152 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X91 CSoutput.t84 commonsourceibias.t117 gnd.t225 gnd.t45 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X92 diffpairibias.t13 diffpairibias.t12 gnd.t229 gnd.t228 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=2.73 ps=14.78 w=7 l=1
X93 CSoutput.t144 a_n6972_8799.t54 vdd.t219 vdd.t159 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=3.12 ps=16.78 w=8 l=0.5
X94 gnd.t258 commonsourceibias.t72 commonsourceibias.t73 gnd.t12 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X95 gnd.t253 commonsourceibias.t118 CSoutput.t175 gnd.t4 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X96 CSoutput.t187 commonsourceibias.t119 gnd.t276 gnd.t39 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X97 gnd.t178 commonsourceibias.t120 CSoutput.t56 gnd.t12 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X98 CSoutput.t69 commonsourceibias.t121 gnd.t199 gnd.t0 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X99 CSoutput.t11 commonsourceibias.t122 gnd.t26 gnd.t18 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X100 vdd.t218 a_n6972_8799.t55 CSoutput.t143 vdd.t144 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X101 CSoutput.t48 commonsourceibias.t123 gnd.t162 gnd.t16 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X102 CSoutput.t142 a_n6972_8799.t56 vdd.t217 vdd.t208 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X103 gnd.t252 commonsourceibias.t124 CSoutput.t174 gnd.t58 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X104 CSoutput.t141 a_n6972_8799.t57 vdd.t216 vdd.t168 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=3.12 ps=16.78 w=8 l=0.5
X105 CSoutput.t140 a_n6972_8799.t58 vdd.t212 vdd.t208 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X106 gnd.t406 commonsourceibias.t70 commonsourceibias.t71 gnd.t196 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X107 gnd.t205 commonsourceibias.t68 commonsourceibias.t69 gnd.t51 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=1.155 ps=7.33 w=7 l=1
X108 gnd.t376 gnd.t374 gnd.t375 gnd.t304 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=0 ps=0 w=7 l=0.7
X109 CSoutput.t181 commonsourceibias.t125 gnd.t267 gnd.t43 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X110 vdd.t122 CSoutput.t196 output.t13 gnd.t131 sky130_fd_pr__nfet_01v8 ad=0.825 pd=5.33 as=0.825 ps=5.33 w=5 l=1
X111 gnd.t363 gnd.t361 plus.t4 gnd.t362 sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.5
X112 output.t12 CSoutput.t197 vdd.t123 gnd.t130 sky130_fd_pr__nfet_01v8 ad=0.825 pd=5.33 as=0.825 ps=5.33 w=5 l=1
X113 CSoutput.t37 commonsourceibias.t126 gnd.t138 gnd.t137 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X114 a_n2903_n3924.t35 plus.t11 a_n6972_8799.t10 gnd.t114 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.7
X115 gnd.t157 commonsourceibias.t127 CSoutput.t45 gnd.t12 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X116 a_n2903_n3924.t12 diffpairibias.t17 gnd.t88 gnd.t87 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=2.73 ps=14.78 w=7 l=1
X117 CSoutput.t198 a_n2318_8322.t24 sky130_fd_pr__cap_mim_m3_1 l=12 w=12
X118 gnd.t373 gnd.t371 gnd.t372 gnd.t293 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=0 ps=0 w=7 l=1
X119 a_n2408_n452.t3 a_n2408_n452.t2 a_n2140_13878.t12 vdd.t107 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X120 vdd.t215 a_n6972_8799.t59 CSoutput.t139 vdd.t178 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X121 vdd.t214 a_n6972_8799.t60 CSoutput.t138 vdd.t206 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X122 gnd.t236 commonsourceibias.t128 CSoutput.t162 gnd.t105 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X123 gnd.t370 gnd.t367 gnd.t369 gnd.t368 sky130_fd_pr__nfet_01v8 ad=1.95 pd=10.78 as=0 ps=0 w=5 l=1
X124 a_n6972_8799.t6 a_n2408_n452.t61 a_n2318_8322.t19 vdd.t19 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X125 a_n2408_n452.t19 a_n2408_n452.t18 a_n2140_13878.t11 vdd.t10 sky130_fd_pr__pfet_01v8 ad=3.51 pd=18.78 as=1.485 ps=9.33 w=9 l=0.5
X126 gnd.t366 gnd.t364 gnd.t365 gnd.t293 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=0 ps=0 w=7 l=1
X127 gnd.t233 commonsourceibias.t129 CSoutput.t160 gnd.t27 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X128 CSoutput.t10 commonsourceibias.t130 gnd.t25 gnd.t24 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X129 commonsourceibias.t67 commonsourceibias.t66 gnd.t216 gnd.t137 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X130 vdd.t213 a_n6972_8799.t61 CSoutput.t137 vdd.t156 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X131 CSoutput.t136 a_n6972_8799.t62 vdd.t211 vdd.t181 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X132 gnd.t64 commonsourceibias.t131 CSoutput.t23 gnd.t63 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X133 a_n2408_n452.t38 minus.t10 a_n2903_n3924.t8 gnd.t79 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.7
X134 gnd.t192 commonsourceibias.t132 CSoutput.t63 gnd.t47 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X135 vdd.t94 vdd.t92 vdd.t93 vdd.t44 sky130_fd_pr__pfet_01v8 ad=3.12 pd=16.78 as=0 ps=0 w=8 l=0.5
X136 vdd.t91 vdd.t89 vdd.t90 vdd.t82 sky130_fd_pr__pfet_01v8 ad=3.51 pd=18.78 as=0 ps=0 w=9 l=0.5
X137 gnd.t206 commonsourceibias.t64 commonsourceibias.t65 gnd.t172 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X138 gnd.t177 commonsourceibias.t133 CSoutput.t55 gnd.t69 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X139 CSoutput.t135 a_n6972_8799.t63 vdd.t210 vdd.t159 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=3.12 ps=16.78 w=8 l=0.5
X140 vdd.t88 vdd.t85 vdd.t87 vdd.t86 sky130_fd_pr__pfet_01v8 ad=3.51 pd=18.78 as=0 ps=0 w=9 l=0.5
X141 a_n2903_n3924.t0 minus.t11 a_n2408_n452.t0 gnd.t6 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.7
X142 gnd.t360 gnd.t358 gnd.t359 gnd.t297 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=0 ps=0 w=7 l=1
X143 vdd.t109 a_n2408_n452.t62 a_n2318_8322.t7 vdd.t108 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X144 a_n2408_n452.t9 a_n2408_n452.t8 a_n2140_13878.t10 vdd.t6 sky130_fd_pr__pfet_01v8 ad=3.51 pd=18.78 as=1.485 ps=9.33 w=9 l=0.5
X145 CSoutput.t83 commonsourceibias.t134 gnd.t224 gnd.t189 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=2.73 ps=14.78 w=7 l=1
X146 a_n2318_8322.t6 a_n2408_n452.t63 vdd.t111 vdd.t110 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X147 gnd.t198 commonsourceibias.t135 CSoutput.t68 gnd.t4 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X148 a_n2903_n3924.t52 diffpairibias.t18 gnd.t262 gnd.t261 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=2.73 ps=14.78 w=7 l=1
X149 output.t11 CSoutput.t199 vdd.t124 gnd.t129 sky130_fd_pr__nfet_01v8 ad=0.825 pd=5.33 as=0.825 ps=5.33 w=5 l=1
X150 CSoutput.t134 a_n6972_8799.t64 vdd.t209 vdd.t208 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X151 vdd.t125 CSoutput.t200 output.t10 gnd.t128 sky130_fd_pr__nfet_01v8 ad=0.825 pd=5.33 as=0.825 ps=5.33 w=5 l=1
X152 gnd.t23 commonsourceibias.t136 CSoutput.t9 gnd.t22 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X153 gnd.t217 commonsourceibias.t62 commonsourceibias.t63 gnd.t101 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X154 CSoutput.t0 commonsourceibias.t137 gnd.t1 gnd.t0 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X155 gnd.t197 commonsourceibias.t138 CSoutput.t67 gnd.t196 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X156 CSoutput.t36 commonsourceibias.t139 gnd.t136 gnd.t135 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X157 CSoutput.t161 commonsourceibias.t140 gnd.t235 gnd.t189 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=2.73 ps=14.78 w=7 l=1
X158 CSoutput.t159 commonsourceibias.t141 gnd.t232 gnd.t141 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X159 a_n2903_n3924.t1 minus.t12 a_n2408_n452.t1 gnd.t7 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.7
X160 a_n2903_n3924.t53 minus.t13 a_n2408_n452.t53 gnd.t108 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=1.155 ps=7.33 w=7 l=0.7
X161 vdd.t26 a_n2408_n452.t64 a_n2140_13878.t22 vdd.t25 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X162 a_n2408_n452.t43 minus.t14 a_n2903_n3924.t16 gnd.t99 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.7
X163 a_n2903_n3924.t34 plus.t12 a_n6972_8799.t27 gnd.t78 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.7
X164 a_n2903_n3924.t33 plus.t13 a_n6972_8799.t26 gnd.t77 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.7
X165 vdd.t84 vdd.t81 vdd.t83 vdd.t82 sky130_fd_pr__pfet_01v8 ad=3.51 pd=18.78 as=0 ps=0 w=9 l=0.5
X166 vdd.t126 CSoutput.t201 output.t9 gnd.t127 sky130_fd_pr__nfet_01v8 ad=0.825 pd=5.33 as=0.825 ps=5.33 w=5 l=1
X167 a_n2408_n452.t39 minus.t15 a_n2903_n3924.t10 gnd.t85 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.7
X168 gnd.t357 gnd.t355 gnd.t356 gnd.t293 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=0 ps=0 w=7 l=1
X169 vdd.t207 a_n6972_8799.t65 CSoutput.t133 vdd.t206 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X170 gnd.t354 gnd.t352 plus.t3 gnd.t353 sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.39 ps=2.78 w=1 l=0.5
X171 a_n6972_8799.t25 plus.t14 a_n2903_n3924.t32 gnd.t113 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.7
X172 a_n6972_8799.t0 plus.t15 a_n2903_n3924.t31 gnd.t112 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=2.73 ps=14.78 w=7 l=0.7
X173 vdd.t80 vdd.t77 vdd.t79 vdd.t78 sky130_fd_pr__pfet_01v8 ad=3.51 pd=18.78 as=0 ps=0 w=9 l=0.5
X174 a_n2318_8322.t5 a_n2408_n452.t65 vdd.t28 vdd.t27 sky130_fd_pr__pfet_01v8 ad=3.51 pd=18.78 as=1.485 ps=9.33 w=9 l=0.5
X175 a_n6972_8799.t32 a_n2408_n452.t66 a_n2318_8322.t18 vdd.t3 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X176 diffpairibias.t11 diffpairibias.t10 gnd.t403 gnd.t402 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=2.73 ps=14.78 w=7 l=1
X177 a_n2408_n452.t51 minus.t16 a_n2903_n3924.t50 gnd.t107 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.7
X178 a_n2408_n452.t5 a_n2408_n452.t4 a_n2140_13878.t9 vdd.t15 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X179 vdd.t205 a_n6972_8799.t66 CSoutput.t132 vdd.t156 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X180 CSoutput.t22 commonsourceibias.t142 gnd.t62 gnd.t20 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X181 a_n6972_8799.t33 a_n2408_n452.t67 a_n2318_8322.t17 vdd.t2 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X182 CSoutput.t131 a_n6972_8799.t67 vdd.t204 vdd.t181 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X183 commonsourceibias.t61 commonsourceibias.t60 gnd.t185 gnd.t184 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X184 output.t8 CSoutput.t202 vdd.t127 gnd.t126 sky130_fd_pr__nfet_01v8 ad=0.825 pd=5.33 as=0.825 ps=5.33 w=5 l=1
X185 gnd.t191 commonsourceibias.t143 CSoutput.t62 gnd.t103 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X186 a_n2140_13878.t8 a_n2408_n452.t32 a_n2408_n452.t33 vdd.t19 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X187 gnd.t57 commonsourceibias.t58 commonsourceibias.t59 gnd.t32 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X188 vdd.t76 vdd.t74 vdd.t75 vdd.t44 sky130_fd_pr__pfet_01v8 ad=3.12 pd=16.78 as=0 ps=0 w=8 l=0.5
X189 a_n2903_n3924.t14 minus.t17 a_n2408_n452.t42 gnd.t92 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.7
X190 CSoutput.t82 commonsourceibias.t144 gnd.t223 gnd.t24 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X191 CSoutput.t130 a_n6972_8799.t68 vdd.t203 vdd.t196 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X192 output.t7 CSoutput.t203 vdd.t128 gnd.t125 sky130_fd_pr__nfet_01v8 ad=0.825 pd=5.33 as=0.825 ps=5.33 w=5 l=1
X193 gnd.t351 gnd.t348 gnd.t350 gnd.t349 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=0 ps=0 w=7 l=0.7
X194 CSoutput.t17 commonsourceibias.t145 gnd.t41 gnd.t29 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X195 vdd.t117 a_n2408_n452.t68 a_n2318_8322.t4 vdd.t116 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=3.51 ps=18.78 w=9 l=0.5
X196 a_n2140_13878.t7 a_n2408_n452.t26 a_n2408_n452.t27 vdd.t16 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=3.51 ps=18.78 w=9 l=0.5
X197 vdd.t202 a_n6972_8799.t69 CSoutput.t129 vdd.t140 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X198 gnd.t266 commonsourceibias.t146 CSoutput.t180 gnd.t47 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X199 gnd.t97 commonsourceibias.t147 CSoutput.t33 gnd.t32 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X200 a_n2408_n452.t29 a_n2408_n452.t28 a_n2140_13878.t6 vdd.t17 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X201 gnd.t245 commonsourceibias.t148 CSoutput.t167 gnd.t35 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X202 gnd.t214 commonsourceibias.t149 CSoutput.t79 gnd.t58 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X203 commonsourceibias.t57 commonsourceibias.t56 gnd.t34 gnd.t0 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X204 gnd.t83 commonsourceibias.t150 CSoutput.t30 gnd.t32 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X205 gnd.t347 gnd.t345 gnd.t346 gnd.t308 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=0 ps=0 w=7 l=1
X206 minus.t3 gnd.t342 gnd.t344 gnd.t343 sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.5
X207 gnd.t405 commonsourceibias.t151 CSoutput.t191 gnd.t60 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=1.155 ps=7.33 w=7 l=1
X208 a_n2903_n3924.t30 plus.t16 a_n6972_8799.t24 gnd.t100 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.7
X209 CSoutput.t28 commonsourceibias.t152 gnd.t75 gnd.t74 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X210 a_n2903_n3924.t15 diffpairibias.t19 gnd.t94 gnd.t93 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=2.73 ps=14.78 w=7 l=1
X211 gnd.t341 gnd.t338 gnd.t340 gnd.t339 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=0 ps=0 w=7 l=1
X212 a_n2903_n3924.t42 diffpairibias.t20 gnd.t149 gnd.t148 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=2.73 ps=14.78 w=7 l=1
X213 commonsourceibias.t55 commonsourceibias.t54 gnd.t241 gnd.t141 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X214 vdd.t201 a_n6972_8799.t70 CSoutput.t128 vdd.t166 sky130_fd_pr__pfet_01v8 ad=3.12 pd=16.78 as=1.32 ps=8.33 w=8 l=0.5
X215 a_n6972_8799.t8 plus.t17 a_n2903_n3924.t29 gnd.t111 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.7
X216 gnd.t337 gnd.t335 gnd.t336 gnd.t312 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=0 ps=0 w=7 l=1
X217 CSoutput.t8 commonsourceibias.t153 gnd.t21 gnd.t20 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X218 CSoutput.t7 commonsourceibias.t154 gnd.t19 gnd.t18 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X219 commonsourceibias.t53 commonsourceibias.t52 gnd.t160 gnd.t43 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X220 gnd.t334 gnd.t331 gnd.t333 gnd.t332 sky130_fd_pr__nfet_01v8 ad=1.95 pd=10.78 as=0 ps=0 w=5 l=1
X221 output.t18 outputibias.t8 gnd.t219 gnd.t218 sky130_fd_pr__nfet_01v8 ad=2.34 pd=12.78 as=2.34 ps=12.78 w=6 l=2
X222 CSoutput.t19 commonsourceibias.t155 gnd.t44 gnd.t43 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X223 CSoutput.t127 a_n6972_8799.t71 vdd.t200 vdd.t199 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X224 commonsourceibias.t51 commonsourceibias.t50 gnd.t269 gnd.t139 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X225 CSoutput.t126 a_n6972_8799.t72 vdd.t198 vdd.t185 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X226 CSoutput.t40 commonsourceibias.t156 gnd.t145 gnd.t16 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X227 outputibias.t7 outputibias.t6 gnd.t243 gnd.t242 sky130_fd_pr__nfet_01v8 ad=2.34 pd=12.78 as=2.34 ps=12.78 w=6 l=2
X228 gnd.t259 commonsourceibias.t48 commonsourceibias.t49 gnd.t22 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X229 vdd.t129 CSoutput.t204 output.t6 gnd.t124 sky130_fd_pr__nfet_01v8 ad=0.825 pd=5.33 as=0.825 ps=5.33 w=5 l=1
X230 diffpairibias.t9 diffpairibias.t8 gnd.t72 gnd.t71 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=2.73 ps=14.78 w=7 l=1
X231 a_n2140_13878.t21 a_n2408_n452.t69 vdd.t119 vdd.t118 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X232 output.t17 outputibias.t9 gnd.t208 gnd.t207 sky130_fd_pr__nfet_01v8 ad=2.34 pd=12.78 as=2.34 ps=12.78 w=6 l=2
X233 vdd.t8 a_n2408_n452.t70 a_n2140_13878.t20 vdd.t7 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X234 CSoutput.t44 commonsourceibias.t157 gnd.t156 gnd.t74 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X235 CSoutput.t166 commonsourceibias.t158 gnd.t240 gnd.t143 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X236 CSoutput.t125 a_n6972_8799.t73 vdd.t197 vdd.t196 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X237 CSoutput.t6 commonsourceibias.t159 gnd.t17 gnd.t16 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X238 gnd.t104 commonsourceibias.t46 commonsourceibias.t47 gnd.t103 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X239 vdd.t141 a_n6972_8799.t74 CSoutput.t124 vdd.t140 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X240 outputibias.t5 outputibias.t4 gnd.t271 gnd.t270 sky130_fd_pr__nfet_01v8 ad=2.34 pd=12.78 as=2.34 ps=12.78 w=6 l=2
X241 commonsourceibias.t45 commonsourceibias.t44 gnd.t166 gnd.t165 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X242 gnd.t212 commonsourceibias.t160 CSoutput.t78 gnd.t47 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X243 plus.t1 gnd.t328 gnd.t330 gnd.t329 sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.5
X244 a_n2140_13878.t5 a_n2408_n452.t16 a_n2408_n452.t17 vdd.t18 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X245 gnd.t76 commonsourceibias.t42 commonsourceibias.t43 gnd.t27 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X246 a_n2903_n3924.t46 minus.t18 a_n2408_n452.t48 gnd.t117 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.7
X247 gnd.t404 commonsourceibias.t161 CSoutput.t190 gnd.t37 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X248 commonsourceibias.t41 commonsourceibias.t40 gnd.t84 gnd.t2 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=2.73 ps=14.78 w=7 l=1
X249 a_n2408_n452.t46 minus.t19 a_n2903_n3924.t44 gnd.t116 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=2.73 ps=14.78 w=7 l=0.7
X250 gnd.t98 commonsourceibias.t38 commonsourceibias.t39 gnd.t10 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X251 a_n2318_8322.t16 a_n2408_n452.t71 a_n6972_8799.t4 vdd.t9 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X252 CSoutput.t16 commonsourceibias.t162 gnd.t40 gnd.t39 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X253 CSoutput.t123 a_n6972_8799.t75 vdd.t143 vdd.t142 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X254 diffpairibias.t7 diffpairibias.t6 gnd.t153 gnd.t152 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=2.73 ps=14.78 w=7 l=1
X255 vdd.t195 a_n6972_8799.t76 CSoutput.t122 vdd.t194 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X256 commonsourceibias.t37 commonsourceibias.t36 gnd.t46 gnd.t45 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X257 a_n2408_n452.t50 minus.t20 a_n2903_n3924.t49 gnd.t115 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.7
X258 a_n2408_n452.t34 minus.t21 a_n2903_n3924.t3 gnd.t53 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.7
X259 gnd.t327 gnd.t325 gnd.t326 gnd.t308 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=0 ps=0 w=7 l=1
X260 vdd.t12 a_n2408_n452.t72 a_n2318_8322.t3 vdd.t11 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=3.51 ps=18.78 w=9 l=0.5
X261 vdd.t193 a_n6972_8799.t77 CSoutput.t121 vdd.t166 sky130_fd_pr__pfet_01v8 ad=3.12 pd=16.78 as=1.32 ps=8.33 w=8 l=0.5
X262 a_n2903_n3924.t13 minus.t22 a_n2408_n452.t41 gnd.t91 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.7
X263 a_n6972_8799.t1 plus.t18 a_n2903_n3924.t28 gnd.t86 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.7
X264 gnd.t251 commonsourceibias.t163 CSoutput.t173 gnd.t37 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X265 a_n2903_n3924.t4 minus.t23 a_n2408_n452.t35 gnd.t54 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.7
X266 gnd.t59 commonsourceibias.t34 commonsourceibias.t35 gnd.t58 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X267 CSoutput.t186 commonsourceibias.t164 gnd.t275 gnd.t135 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X268 a_n2140_13878.t19 a_n2408_n452.t73 vdd.t14 vdd.t13 sky130_fd_pr__pfet_01v8 ad=3.51 pd=18.78 as=1.485 ps=9.33 w=9 l=0.5
X269 output.t5 CSoutput.t205 vdd.t130 gnd.t123 sky130_fd_pr__nfet_01v8 ad=0.825 pd=5.33 as=0.825 ps=5.33 w=5 l=1
X270 vdd.t192 a_n6972_8799.t78 CSoutput.t120 vdd.t178 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X271 CSoutput.t119 a_n6972_8799.t79 vdd.t191 vdd.t185 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X272 CSoutput.t118 a_n6972_8799.t80 vdd.t190 vdd.t176 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X273 gnd.t324 gnd.t322 minus.t2 gnd.t323 sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.39 ps=2.78 w=1 l=0.5
X274 gnd.t176 commonsourceibias.t165 CSoutput.t54 gnd.t101 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X275 gnd.t321 gnd.t318 gnd.t320 gnd.t319 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=0 ps=0 w=7 l=1
X276 a_n2903_n3924.t2 diffpairibias.t21 gnd.t50 gnd.t49 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=2.73 ps=14.78 w=7 l=1
X277 a_n2318_8322.t15 a_n2408_n452.t74 a_n6972_8799.t36 vdd.t15 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X278 vdd.t121 a_n2408_n452.t75 a_n2318_8322.t2 vdd.t120 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X279 CSoutput.t206 a_n2318_8322.t25 sky130_fd_pr__cap_mim_m3_1 l=12 w=12
X280 CSoutput.t117 a_n6972_8799.t81 vdd.t186 vdd.t185 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X281 gnd.t106 commonsourceibias.t32 commonsourceibias.t33 gnd.t105 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X282 vdd.t73 vdd.t71 vdd.t72 vdd.t52 sky130_fd_pr__pfet_01v8 ad=3.12 pd=16.78 as=0 ps=0 w=8 l=0.5
X283 vdd.t189 a_n6972_8799.t82 CSoutput.t116 vdd.t138 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X284 outputibias.t3 outputibias.t2 gnd.t90 gnd.t89 sky130_fd_pr__nfet_01v8 ad=2.34 pd=12.78 as=2.34 ps=12.78 w=6 l=2
X285 CSoutput.t115 a_n6972_8799.t83 vdd.t188 vdd.t154 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X286 vdd.t187 a_n6972_8799.t84 CSoutput.t114 vdd.t171 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X287 vdd.t184 a_n6972_8799.t85 CSoutput.t113 vdd.t150 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X288 a_n6972_8799.t7 plus.t19 a_n2903_n3924.t27 gnd.t110 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.7
X289 output.t19 outputibias.t10 gnd.t280 gnd.t279 sky130_fd_pr__nfet_01v8 ad=2.34 pd=12.78 as=2.34 ps=12.78 w=6 l=2
X290 vdd.t70 vdd.t68 vdd.t69 vdd.t40 sky130_fd_pr__pfet_01v8 ad=3.12 pd=16.78 as=0 ps=0 w=8 l=0.5
X291 gnd.t188 commonsourceibias.t30 commonsourceibias.t31 gnd.t63 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X292 vdd.t67 vdd.t64 vdd.t66 vdd.t65 sky130_fd_pr__pfet_01v8 ad=3.51 pd=18.78 as=0 ps=0 w=9 l=0.5
X293 CSoutput.t172 commonsourceibias.t166 gnd.t250 gnd.t67 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X294 a_n2903_n3924.t26 plus.t20 a_n6972_8799.t2 gnd.t109 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=1.155 ps=7.33 w=7 l=0.7
X295 gnd.t317 gnd.t315 gnd.t316 gnd.t297 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=0 ps=0 w=7 l=1
X296 vdd.t131 CSoutput.t207 output.t4 gnd.t122 sky130_fd_pr__nfet_01v8 ad=0.825 pd=5.33 as=0.825 ps=5.33 w=5 l=1
X297 CSoutput.t185 commonsourceibias.t167 gnd.t274 gnd.t139 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X298 CSoutput.t112 a_n6972_8799.t86 vdd.t183 vdd.t142 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X299 a_n2140_13878.t4 a_n2408_n452.t14 a_n2408_n452.t15 vdd.t1 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X300 a_n2318_8322.t14 a_n2408_n452.t76 a_n6972_8799.t34 vdd.t0 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X301 diffpairibias.t5 diffpairibias.t4 gnd.t264 gnd.t263 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=2.73 ps=14.78 w=7 l=1
X302 CSoutput.t208 a_n2318_8322.t25 sky130_fd_pr__cap_mim_m3_1 l=12 w=12
X303 gnd.t314 gnd.t311 gnd.t313 gnd.t312 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=0 ps=0 w=7 l=1
X304 CSoutput.t111 a_n6972_8799.t87 vdd.t182 vdd.t181 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X305 gnd.t281 commonsourceibias.t28 commonsourceibias.t29 gnd.t4 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X306 output.t3 CSoutput.t209 vdd.t132 gnd.t121 sky130_fd_pr__nfet_01v8 ad=0.825 pd=5.33 as=0.825 ps=5.33 w=5 l=1
X307 vdd.t180 a_n6972_8799.t88 CSoutput.t110 vdd.t171 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X308 CSoutput.t53 commonsourceibias.t168 gnd.t175 gnd.t45 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X309 commonsourceibias.t27 commonsourceibias.t26 gnd.t260 gnd.t189 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=2.73 ps=14.78 w=7 l=1
X310 vdd.t179 a_n6972_8799.t89 CSoutput.t109 vdd.t178 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X311 a_n2318_8322.t1 a_n2408_n452.t77 vdd.t113 vdd.t112 sky130_fd_pr__pfet_01v8 ad=3.51 pd=18.78 as=1.485 ps=9.33 w=9 l=0.5
X312 CSoutput.t108 a_n6972_8799.t90 vdd.t177 vdd.t176 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X313 vdd.t63 vdd.t61 vdd.t62 vdd.t36 sky130_fd_pr__pfet_01v8 ad=3.51 pd=18.78 as=0 ps=0 w=9 l=0.5
X314 gnd.t155 commonsourceibias.t169 CSoutput.t43 gnd.t69 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X315 vdd.t23 a_n2408_n452.t78 a_n2140_13878.t18 vdd.t22 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=3.51 ps=18.78 w=9 l=0.5
X316 plus.t0 gnd.t289 gnd.t291 gnd.t290 sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.5
X317 CSoutput.t107 a_n6972_8799.t91 vdd.t175 vdd.t174 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X318 vdd.t60 vdd.t58 vdd.t59 vdd.t52 sky130_fd_pr__pfet_01v8 ad=3.12 pd=16.78 as=0 ps=0 w=8 l=0.5
X319 CSoutput.t106 a_n6972_8799.t92 vdd.t173 vdd.t154 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X320 a_n2903_n3924.t25 plus.t21 a_n6972_8799.t14 gnd.t108 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=1.155 ps=7.33 w=7 l=0.7
X321 vdd.t172 a_n6972_8799.t93 CSoutput.t105 vdd.t171 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X322 vdd.t170 a_n6972_8799.t94 CSoutput.t104 vdd.t150 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X323 gnd.t249 commonsourceibias.t170 CSoutput.t171 gnd.t10 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X324 gnd.t15 commonsourceibias.t171 CSoutput.t5 gnd.t14 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X325 vdd.t57 vdd.t55 vdd.t56 vdd.t40 sky130_fd_pr__pfet_01v8 ad=3.12 pd=16.78 as=0 ps=0 w=8 l=0.5
X326 output.t2 CSoutput.t210 vdd.t133 gnd.t120 sky130_fd_pr__nfet_01v8 ad=0.825 pd=5.33 as=0.825 ps=5.33 w=5 l=1
X327 a_n2903_n3924.t7 minus.t24 a_n2408_n452.t37 gnd.t78 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.7
X328 a_n2318_8322.t13 a_n2408_n452.t79 a_n6972_8799.t19 vdd.t24 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X329 commonsourceibias.t25 commonsourceibias.t24 gnd.t234 gnd.t20 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X330 CSoutput.t103 a_n6972_8799.t95 vdd.t169 vdd.t168 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=3.12 ps=16.78 w=8 l=0.5
X331 a_n6972_8799.t31 a_n2408_n452.t80 a_n2318_8322.t12 vdd.t1 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X332 a_n6972_8799.t16 plus.t22 a_n2903_n3924.t24 gnd.t85 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.7
X333 vdd.t167 a_n6972_8799.t96 CSoutput.t102 vdd.t166 sky130_fd_pr__pfet_01v8 ad=3.12 pd=16.78 as=1.32 ps=8.33 w=8 l=0.5
X334 a_n2140_13878.t17 a_n2408_n452.t81 vdd.t30 vdd.t29 sky130_fd_pr__pfet_01v8 ad=3.51 pd=18.78 as=1.485 ps=9.33 w=9 l=0.5
X335 gnd.t174 commonsourceibias.t172 CSoutput.t52 gnd.t63 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X336 vdd.t165 a_n6972_8799.t97 CSoutput.t101 vdd.t152 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X337 a_n2408_n452.t55 minus.t25 a_n2903_n3924.t55 gnd.t113 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.7
X338 CSoutput.t100 a_n6972_8799.t98 vdd.t164 vdd.t142 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X339 commonsourceibias.t23 commonsourceibias.t22 gnd.t407 gnd.t24 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X340 output.t1 CSoutput.t211 vdd.t134 gnd.t119 sky130_fd_pr__nfet_01v8 ad=1.95 pd=10.78 as=0.825 ps=5.33 w=5 l=1
X341 gnd.t310 gnd.t307 gnd.t309 gnd.t308 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=0 ps=0 w=7 l=1
X342 gnd.t42 commonsourceibias.t173 CSoutput.t18 gnd.t35 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X343 vdd.t54 vdd.t51 vdd.t53 vdd.t52 sky130_fd_pr__pfet_01v8 ad=3.12 pd=16.78 as=0 ps=0 w=8 l=0.5
X344 a_n2318_8322.t11 a_n2408_n452.t82 a_n6972_8799.t29 vdd.t6 sky130_fd_pr__pfet_01v8 ad=3.51 pd=18.78 as=1.485 ps=9.33 w=9 l=0.5
X345 commonsourceibias.t21 commonsourceibias.t20 gnd.t213 gnd.t29 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X346 a_n6972_8799.t15 plus.t23 a_n2903_n3924.t23 gnd.t107 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.7
X347 gnd.t306 gnd.t303 gnd.t305 gnd.t304 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=0 ps=0 w=7 l=0.7
X348 gnd.t302 gnd.t300 minus.t1 gnd.t301 sky130_fd_pr__nfet_01v8 ad=0.39 pd=2.78 as=0.165 ps=1.33 w=1 l=0.5
X349 gnd.t13 commonsourceibias.t174 CSoutput.t4 gnd.t12 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X350 vdd.t50 vdd.t47 vdd.t49 vdd.t48 sky130_fd_pr__pfet_01v8 ad=3.12 pd=16.78 as=0 ps=0 w=8 l=0.5
X351 CSoutput.t77 commonsourceibias.t175 gnd.t211 gnd.t135 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X352 a_n2903_n3924.t54 minus.t26 a_n2408_n452.t54 gnd.t114 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.7
X353 gnd.t36 commonsourceibias.t18 commonsourceibias.t19 gnd.t35 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X354 a_n2140_13878.t3 a_n2408_n452.t22 a_n2408_n452.t23 vdd.t3 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X355 outputibias.t1 outputibias.t0 gnd.t187 gnd.t186 sky130_fd_pr__nfet_01v8 ad=2.34 pd=12.78 as=2.34 ps=12.78 w=6 l=2
X356 vdd.t163 a_n6972_8799.t99 CSoutput.t99 vdd.t148 sky130_fd_pr__pfet_01v8 ad=3.12 pd=16.78 as=1.32 ps=8.33 w=8 l=0.5
X357 a_n2903_n3924.t22 plus.t24 a_n6972_8799.t22 gnd.t92 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.7
X358 gnd.t244 commonsourceibias.t16 commonsourceibias.t17 gnd.t60 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=1.155 ps=7.33 w=7 l=1
X359 vdd.t46 vdd.t43 vdd.t45 vdd.t44 sky130_fd_pr__pfet_01v8 ad=3.12 pd=16.78 as=0 ps=0 w=8 l=0.5
X360 vdd.t42 vdd.t39 vdd.t41 vdd.t40 sky130_fd_pr__pfet_01v8 ad=3.12 pd=16.78 as=0 ps=0 w=8 l=0.5
X361 commonsourceibias.t15 commonsourceibias.t14 gnd.t161 gnd.t74 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X362 gnd.t299 gnd.t296 gnd.t298 gnd.t297 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=0 ps=0 w=7 l=1
X363 gnd.t265 commonsourceibias.t176 CSoutput.t179 gnd.t196 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X364 gnd.t96 commonsourceibias.t177 CSoutput.t32 gnd.t51 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=1.155 ps=7.33 w=7 l=1
X365 a_n2903_n3924.t5 diffpairibias.t22 gnd.t56 gnd.t55 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=2.73 ps=14.78 w=7 l=1
X366 gnd.t134 commonsourceibias.t178 CSoutput.t35 gnd.t105 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X367 vdd.t162 a_n6972_8799.t100 CSoutput.t98 vdd.t144 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X368 CSoutput.t42 commonsourceibias.t179 gnd.t154 gnd.t18 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X369 gnd.t82 commonsourceibias.t180 CSoutput.t29 gnd.t69 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X370 CSoutput.t27 commonsourceibias.t181 gnd.t73 gnd.t67 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X371 a_n2408_n452.t7 a_n2408_n452.t6 a_n2140_13878.t2 vdd.t24 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X372 gnd.t295 gnd.t292 gnd.t294 gnd.t293 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=0 ps=0 w=7 l=1
X373 a_n6972_8799.t30 a_n2408_n452.t83 a_n2318_8322.t10 vdd.t20 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X374 vdd.t135 CSoutput.t212 output.t0 gnd.t118 sky130_fd_pr__nfet_01v8 ad=0.825 pd=5.33 as=1.95 ps=10.78 w=5 l=1
X375 vdd.t161 a_n6972_8799.t101 CSoutput.t97 vdd.t148 sky130_fd_pr__pfet_01v8 ad=3.12 pd=16.78 as=1.32 ps=8.33 w=8 l=0.5
X376 CSoutput.t96 a_n6972_8799.t102 vdd.t160 vdd.t159 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=3.12 ps=16.78 w=8 l=0.5
X377 a_n6972_8799.t21 plus.t25 a_n2903_n3924.t21 gnd.t79 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.7
X378 vdd.t158 a_n6972_8799.t103 CSoutput.t95 vdd.t138 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X379 CSoutput.t76 commonsourceibias.t182 gnd.t210 gnd.t143 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X380 gnd.t61 commonsourceibias.t183 CSoutput.t21 gnd.t60 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=1.155 ps=7.33 w=7 l=1
X381 commonsourceibias.t13 commonsourceibias.t12 gnd.t147 gnd.t18 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X382 CSoutput.t61 commonsourceibias.t184 gnd.t190 gnd.t189 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=2.73 ps=14.78 w=7 l=1
X383 gnd.t288 gnd.t285 gnd.t287 gnd.t286 sky130_fd_pr__nfet_01v8 ad=2.34 pd=12.78 as=0 ps=0 w=6 l=2
X384 diffpairibias.t3 diffpairibias.t2 gnd.t9 gnd.t8 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=2.73 ps=14.78 w=7 l=1
X385 vdd.t157 a_n6972_8799.t104 CSoutput.t94 vdd.t156 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X386 CSoutput.t93 a_n6972_8799.t105 vdd.t155 vdd.t154 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X387 a_n2318_8322.t9 a_n2408_n452.t84 a_n6972_8799.t35 vdd.t17 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X388 CSoutput.t81 commonsourceibias.t185 gnd.t222 gnd.t137 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X389 gnd.t248 commonsourceibias.t186 CSoutput.t170 gnd.t37 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X390 a_n2903_n3924.t20 plus.t26 a_n6972_8799.t9 gnd.t6 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.7
X391 vdd.t153 a_n6972_8799.t106 CSoutput.t92 vdd.t152 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X392 diffpairibias.t1 diffpairibias.t0 gnd.t231 gnd.t230 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=2.73 ps=14.78 w=7 l=1
X393 gnd.t273 commonsourceibias.t187 CSoutput.t184 gnd.t196 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X394 CSoutput.t213 a_n2318_8322.t24 sky130_fd_pr__cap_mim_m3_1 l=12 w=12
X395 commonsourceibias.t11 commonsourceibias.t10 gnd.t144 gnd.t143 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X396 gnd.t173 commonsourceibias.t188 CSoutput.t51 gnd.t172 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X397 a_n2903_n3924.t19 plus.t27 a_n6972_8799.t20 gnd.t7 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.7
X398 commonsourceibias.t9 commonsourceibias.t8 gnd.t167 gnd.t16 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X399 CSoutput.t31 commonsourceibias.t189 gnd.t95 gnd.t2 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=2.73 ps=14.78 w=7 l=1
X400 vdd.t38 vdd.t35 vdd.t37 vdd.t36 sky130_fd_pr__pfet_01v8 ad=3.51 pd=18.78 as=0 ps=0 w=9 l=0.5
X401 vdd.t115 a_n2408_n452.t85 a_n2140_13878.t16 vdd.t114 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=3.51 ps=18.78 w=9 l=0.5
X402 a_n6972_8799.t23 plus.t28 a_n2903_n3924.t18 gnd.t99 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.7
X403 gnd.t48 commonsourceibias.t6 commonsourceibias.t7 gnd.t47 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X404 vdd.t34 vdd.t31 vdd.t33 vdd.t32 sky130_fd_pr__pfet_01v8 ad=3.51 pd=18.78 as=0 ps=0 w=9 l=0.5
X405 a_n2903_n3924.t6 minus.t27 a_n2408_n452.t36 gnd.t77 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.7
X406 vdd.t151 a_n6972_8799.t107 CSoutput.t91 vdd.t150 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X407 vdd.t149 a_n6972_8799.t108 CSoutput.t90 vdd.t148 sky130_fd_pr__pfet_01v8 ad=3.12 pd=16.78 as=1.32 ps=8.33 w=8 l=0.5
X408 gnd.t38 commonsourceibias.t4 commonsourceibias.t5 gnd.t37 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X409 CSoutput.t89 a_n6972_8799.t109 vdd.t147 vdd.t146 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X410 gnd.t102 commonsourceibias.t190 CSoutput.t34 gnd.t101 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X411 a_n2408_n452.t45 minus.t28 a_n2903_n3924.t43 gnd.t112 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=2.73 ps=14.78 w=7 l=0.7
X412 commonsourceibias.t3 commonsourceibias.t2 gnd.t220 gnd.t39 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X413 gnd.t52 commonsourceibias.t191 CSoutput.t20 gnd.t51 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=1.155 ps=7.33 w=7 l=1
X414 gnd.t247 commonsourceibias.t192 CSoutput.t169 gnd.t172 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X415 gnd.t11 commonsourceibias.t193 CSoutput.t3 gnd.t10 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X416 a_n2318_8322.t8 a_n2408_n452.t86 a_n6972_8799.t37 vdd.t10 sky130_fd_pr__pfet_01v8 ad=3.51 pd=18.78 as=1.485 ps=9.33 w=9 l=0.5
X417 vdd.t145 a_n6972_8799.t110 CSoutput.t88 vdd.t144 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X418 output.t16 outputibias.t11 gnd.t164 gnd.t163 sky130_fd_pr__nfet_01v8 ad=2.34 pd=12.78 as=2.34 ps=12.78 w=6 l=2
X419 gnd.t171 commonsourceibias.t194 CSoutput.t50 gnd.t14 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X420 a_n2318_8322.t0 a_n2408_n452.t87 vdd.t137 vdd.t136 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X421 gnd.t215 commonsourceibias.t195 CSoutput.t80 gnd.t63 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X422 a_n2140_13878.t1 a_n2408_n452.t12 a_n2408_n452.t13 vdd.t21 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=3.51 ps=18.78 w=9 l=0.5
X423 gnd.t209 commonsourceibias.t196 CSoutput.t75 gnd.t14 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X424 CSoutput.t168 commonsourceibias.t197 gnd.t246 gnd.t143 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X425 vdd.t139 a_n6972_8799.t111 CSoutput.t87 vdd.t138 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X426 commonsourceibias.t1 commonsourceibias.t0 gnd.t221 gnd.t135 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X427 CSoutput.t183 commonsourceibias.t198 gnd.t272 gnd.t184 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X428 minus.t0 gnd.t282 gnd.t284 gnd.t283 sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.5
X429 a_n2903_n3924.t9 diffpairibias.t23 gnd.t81 gnd.t80 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=2.73 ps=14.78 w=7 l=1
X430 a_n2408_n452.t31 a_n2408_n452.t30 a_n2140_13878.t0 vdd.t9 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X431 gnd.t170 commonsourceibias.t199 CSoutput.t49 gnd.t27 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
R0 a_n6972_8799.n141 a_n6972_8799.t54 490.524
R1 a_n6972_8799.n152 a_n6972_8799.t63 490.524
R2 a_n6972_8799.n164 a_n6972_8799.t102 490.524
R3 a_n6972_8799.n107 a_n6972_8799.t99 490.524
R4 a_n6972_8799.n118 a_n6972_8799.t108 490.524
R5 a_n6972_8799.n130 a_n6972_8799.t101 490.524
R6 a_n6972_8799.n30 a_n6972_8799.t70 484.3
R7 a_n6972_8799.n147 a_n6972_8799.t58 464.166
R8 a_n6972_8799.n146 a_n6972_8799.t103 464.166
R9 a_n6972_8799.n137 a_n6972_8799.t80 464.166
R10 a_n6972_8799.n145 a_n6972_8799.t78 464.166
R11 a_n6972_8799.n144 a_n6972_8799.t42 464.166
R12 a_n6972_8799.n138 a_n6972_8799.t84 464.166
R13 a_n6972_8799.n143 a_n6972_8799.t83 464.166
R14 a_n6972_8799.n142 a_n6972_8799.t44 464.166
R15 a_n6972_8799.n139 a_n6972_8799.t43 464.166
R16 a_n6972_8799.n140 a_n6972_8799.t97 464.166
R17 a_n6972_8799.n39 a_n6972_8799.t77 484.3
R18 a_n6972_8799.n158 a_n6972_8799.t64 464.166
R19 a_n6972_8799.n157 a_n6972_8799.t111 464.166
R20 a_n6972_8799.n148 a_n6972_8799.t90 464.166
R21 a_n6972_8799.n156 a_n6972_8799.t89 464.166
R22 a_n6972_8799.n155 a_n6972_8799.t49 464.166
R23 a_n6972_8799.n149 a_n6972_8799.t93 464.166
R24 a_n6972_8799.n154 a_n6972_8799.t92 464.166
R25 a_n6972_8799.n153 a_n6972_8799.t51 464.166
R26 a_n6972_8799.n150 a_n6972_8799.t50 464.166
R27 a_n6972_8799.n151 a_n6972_8799.t106 464.166
R28 a_n6972_8799.n48 a_n6972_8799.t96 484.3
R29 a_n6972_8799.n170 a_n6972_8799.t56 464.166
R30 a_n6972_8799.n169 a_n6972_8799.t82 464.166
R31 a_n6972_8799.n160 a_n6972_8799.t46 464.166
R32 a_n6972_8799.n168 a_n6972_8799.t59 464.166
R33 a_n6972_8799.n167 a_n6972_8799.t109 464.166
R34 a_n6972_8799.n161 a_n6972_8799.t88 464.166
R35 a_n6972_8799.n166 a_n6972_8799.t105 464.166
R36 a_n6972_8799.n165 a_n6972_8799.t76 464.166
R37 a_n6972_8799.n162 a_n6972_8799.t91 464.166
R38 a_n6972_8799.n163 a_n6972_8799.t53 464.166
R39 a_n6972_8799.n106 a_n6972_8799.t68 464.166
R40 a_n6972_8799.n105 a_n6972_8799.t69 464.166
R41 a_n6972_8799.n108 a_n6972_8799.t86 464.166
R42 a_n6972_8799.n104 a_n6972_8799.t61 464.166
R43 a_n6972_8799.n109 a_n6972_8799.t62 464.166
R44 a_n6972_8799.n110 a_n6972_8799.t85 464.166
R45 a_n6972_8799.n103 a_n6972_8799.t40 464.166
R46 a_n6972_8799.n111 a_n6972_8799.t60 464.166
R47 a_n6972_8799.n102 a_n6972_8799.t72 464.166
R48 a_n6972_8799.n112 a_n6972_8799.t100 464.166
R49 a_n6972_8799.n117 a_n6972_8799.t73 464.166
R50 a_n6972_8799.n116 a_n6972_8799.t74 464.166
R51 a_n6972_8799.n119 a_n6972_8799.t98 464.166
R52 a_n6972_8799.n115 a_n6972_8799.t66 464.166
R53 a_n6972_8799.n120 a_n6972_8799.t67 464.166
R54 a_n6972_8799.n121 a_n6972_8799.t94 464.166
R55 a_n6972_8799.n114 a_n6972_8799.t47 464.166
R56 a_n6972_8799.n122 a_n6972_8799.t65 464.166
R57 a_n6972_8799.n113 a_n6972_8799.t79 464.166
R58 a_n6972_8799.n123 a_n6972_8799.t110 464.166
R59 a_n6972_8799.n129 a_n6972_8799.t52 464.166
R60 a_n6972_8799.n128 a_n6972_8799.t41 464.166
R61 a_n6972_8799.n131 a_n6972_8799.t75 464.166
R62 a_n6972_8799.n127 a_n6972_8799.t104 464.166
R63 a_n6972_8799.n132 a_n6972_8799.t87 464.166
R64 a_n6972_8799.n133 a_n6972_8799.t107 464.166
R65 a_n6972_8799.n126 a_n6972_8799.t71 464.166
R66 a_n6972_8799.n134 a_n6972_8799.t45 464.166
R67 a_n6972_8799.n125 a_n6972_8799.t81 464.166
R68 a_n6972_8799.n135 a_n6972_8799.t55 464.166
R69 a_n6972_8799.n38 a_n6972_8799.n37 75.3623
R70 a_n6972_8799.n36 a_n6972_8799.n24 70.3058
R71 a_n6972_8799.n24 a_n6972_8799.n35 70.1674
R72 a_n6972_8799.n35 a_n6972_8799.n138 20.9683
R73 a_n6972_8799.n34 a_n6972_8799.n25 75.0448
R74 a_n6972_8799.n144 a_n6972_8799.n34 11.2134
R75 a_n6972_8799.n33 a_n6972_8799.n25 80.4688
R76 a_n6972_8799.n27 a_n6972_8799.n32 74.73
R77 a_n6972_8799.n31 a_n6972_8799.n27 70.1674
R78 a_n6972_8799.n147 a_n6972_8799.n31 20.9683
R79 a_n6972_8799.n26 a_n6972_8799.n30 70.5844
R80 a_n6972_8799.n47 a_n6972_8799.n46 75.3623
R81 a_n6972_8799.n45 a_n6972_8799.n20 70.3058
R82 a_n6972_8799.n20 a_n6972_8799.n44 70.1674
R83 a_n6972_8799.n44 a_n6972_8799.n149 20.9683
R84 a_n6972_8799.n43 a_n6972_8799.n21 75.0448
R85 a_n6972_8799.n155 a_n6972_8799.n43 11.2134
R86 a_n6972_8799.n42 a_n6972_8799.n21 80.4688
R87 a_n6972_8799.n23 a_n6972_8799.n41 74.73
R88 a_n6972_8799.n40 a_n6972_8799.n23 70.1674
R89 a_n6972_8799.n158 a_n6972_8799.n40 20.9683
R90 a_n6972_8799.n22 a_n6972_8799.n39 70.5844
R91 a_n6972_8799.n56 a_n6972_8799.n55 75.3623
R92 a_n6972_8799.n54 a_n6972_8799.n16 70.3058
R93 a_n6972_8799.n16 a_n6972_8799.n53 70.1674
R94 a_n6972_8799.n53 a_n6972_8799.n161 20.9683
R95 a_n6972_8799.n52 a_n6972_8799.n17 75.0448
R96 a_n6972_8799.n167 a_n6972_8799.n52 11.2134
R97 a_n6972_8799.n51 a_n6972_8799.n17 80.4688
R98 a_n6972_8799.n19 a_n6972_8799.n50 74.73
R99 a_n6972_8799.n49 a_n6972_8799.n19 70.1674
R100 a_n6972_8799.n170 a_n6972_8799.n49 20.9683
R101 a_n6972_8799.n18 a_n6972_8799.n48 70.5844
R102 a_n6972_8799.n12 a_n6972_8799.n65 70.5844
R103 a_n6972_8799.n64 a_n6972_8799.n13 70.1674
R104 a_n6972_8799.n64 a_n6972_8799.n102 20.9683
R105 a_n6972_8799.n13 a_n6972_8799.n63 74.73
R106 a_n6972_8799.n111 a_n6972_8799.n63 11.843
R107 a_n6972_8799.n62 a_n6972_8799.n14 80.4688
R108 a_n6972_8799.n62 a_n6972_8799.n103 0.365327
R109 a_n6972_8799.n14 a_n6972_8799.n61 75.0448
R110 a_n6972_8799.n60 a_n6972_8799.n15 70.1674
R111 a_n6972_8799.n60 a_n6972_8799.n104 20.9683
R112 a_n6972_8799.n15 a_n6972_8799.n59 70.3058
R113 a_n6972_8799.n108 a_n6972_8799.n59 20.6913
R114 a_n6972_8799.n58 a_n6972_8799.n57 75.3623
R115 a_n6972_8799.n8 a_n6972_8799.n74 70.5844
R116 a_n6972_8799.n73 a_n6972_8799.n9 70.1674
R117 a_n6972_8799.n73 a_n6972_8799.n113 20.9683
R118 a_n6972_8799.n9 a_n6972_8799.n72 74.73
R119 a_n6972_8799.n122 a_n6972_8799.n72 11.843
R120 a_n6972_8799.n71 a_n6972_8799.n10 80.4688
R121 a_n6972_8799.n71 a_n6972_8799.n114 0.365327
R122 a_n6972_8799.n10 a_n6972_8799.n70 75.0448
R123 a_n6972_8799.n69 a_n6972_8799.n11 70.1674
R124 a_n6972_8799.n69 a_n6972_8799.n115 20.9683
R125 a_n6972_8799.n11 a_n6972_8799.n68 70.3058
R126 a_n6972_8799.n119 a_n6972_8799.n68 20.6913
R127 a_n6972_8799.n67 a_n6972_8799.n66 75.3623
R128 a_n6972_8799.n4 a_n6972_8799.n83 70.5844
R129 a_n6972_8799.n82 a_n6972_8799.n5 70.1674
R130 a_n6972_8799.n82 a_n6972_8799.n125 20.9683
R131 a_n6972_8799.n5 a_n6972_8799.n81 74.73
R132 a_n6972_8799.n134 a_n6972_8799.n81 11.843
R133 a_n6972_8799.n80 a_n6972_8799.n6 80.4688
R134 a_n6972_8799.n80 a_n6972_8799.n126 0.365327
R135 a_n6972_8799.n6 a_n6972_8799.n79 75.0448
R136 a_n6972_8799.n78 a_n6972_8799.n7 70.1674
R137 a_n6972_8799.n78 a_n6972_8799.n127 20.9683
R138 a_n6972_8799.n7 a_n6972_8799.n77 70.3058
R139 a_n6972_8799.n131 a_n6972_8799.n77 20.6913
R140 a_n6972_8799.n76 a_n6972_8799.n75 75.3623
R141 a_n6972_8799.n177 a_n6972_8799.n84 98.9633
R142 a_n6972_8799.n28 a_n6972_8799.n85 98.9631
R143 a_n6972_8799.n29 a_n6972_8799.n175 98.6055
R144 a_n6972_8799.n29 a_n6972_8799.n176 98.6055
R145 a_n6972_8799.n28 a_n6972_8799.n86 98.6055
R146 a_n6972_8799.n28 a_n6972_8799.n87 98.6055
R147 a_n6972_8799.n89 a_n6972_8799.n88 98.6055
R148 a_n6972_8799.n178 a_n6972_8799.n177 98.6054
R149 a_n6972_8799.n1 a_n6972_8799.n90 81.3764
R150 a_n6972_8799.n3 a_n6972_8799.n96 81.3764
R151 a_n6972_8799.n0 a_n6972_8799.n93 81.3764
R152 a_n6972_8799.n2 a_n6972_8799.n99 80.9324
R153 a_n6972_8799.n2 a_n6972_8799.n100 80.9324
R154 a_n6972_8799.n1 a_n6972_8799.n101 80.9324
R155 a_n6972_8799.n1 a_n6972_8799.n92 80.9324
R156 a_n6972_8799.n1 a_n6972_8799.n91 80.9324
R157 a_n6972_8799.n3 a_n6972_8799.n97 80.9324
R158 a_n6972_8799.n0 a_n6972_8799.n98 80.9324
R159 a_n6972_8799.n0 a_n6972_8799.n95 80.9324
R160 a_n6972_8799.n0 a_n6972_8799.n94 80.9324
R161 a_n6972_8799.n31 a_n6972_8799.n146 20.9683
R162 a_n6972_8799.n145 a_n6972_8799.n144 48.2005
R163 a_n6972_8799.n143 a_n6972_8799.n35 20.9683
R164 a_n6972_8799.n140 a_n6972_8799.n139 48.2005
R165 a_n6972_8799.n40 a_n6972_8799.n157 20.9683
R166 a_n6972_8799.n156 a_n6972_8799.n155 48.2005
R167 a_n6972_8799.n154 a_n6972_8799.n44 20.9683
R168 a_n6972_8799.n151 a_n6972_8799.n150 48.2005
R169 a_n6972_8799.n49 a_n6972_8799.n169 20.9683
R170 a_n6972_8799.n168 a_n6972_8799.n167 48.2005
R171 a_n6972_8799.n166 a_n6972_8799.n53 20.9683
R172 a_n6972_8799.n163 a_n6972_8799.n162 48.2005
R173 a_n6972_8799.n106 a_n6972_8799.n105 48.2005
R174 a_n6972_8799.n109 a_n6972_8799.n60 20.9683
R175 a_n6972_8799.n110 a_n6972_8799.n103 48.2005
R176 a_n6972_8799.n112 a_n6972_8799.n64 20.9683
R177 a_n6972_8799.n117 a_n6972_8799.n116 48.2005
R178 a_n6972_8799.n120 a_n6972_8799.n69 20.9683
R179 a_n6972_8799.n121 a_n6972_8799.n114 48.2005
R180 a_n6972_8799.n123 a_n6972_8799.n73 20.9683
R181 a_n6972_8799.n129 a_n6972_8799.n128 48.2005
R182 a_n6972_8799.n132 a_n6972_8799.n78 20.9683
R183 a_n6972_8799.n133 a_n6972_8799.n126 48.2005
R184 a_n6972_8799.n135 a_n6972_8799.n82 20.9683
R185 a_n6972_8799.n33 a_n6972_8799.n137 47.835
R186 a_n6972_8799.n36 a_n6972_8799.n142 20.6913
R187 a_n6972_8799.n42 a_n6972_8799.n148 47.835
R188 a_n6972_8799.n45 a_n6972_8799.n153 20.6913
R189 a_n6972_8799.n51 a_n6972_8799.n160 47.835
R190 a_n6972_8799.n54 a_n6972_8799.n165 20.6913
R191 a_n6972_8799.n104 a_n6972_8799.n59 21.4216
R192 a_n6972_8799.n115 a_n6972_8799.n68 21.4216
R193 a_n6972_8799.n127 a_n6972_8799.n77 21.4216
R194 a_n6972_8799.t48 a_n6972_8799.n65 484.3
R195 a_n6972_8799.t57 a_n6972_8799.n74 484.3
R196 a_n6972_8799.t95 a_n6972_8799.n83 484.3
R197 a_n6972_8799.n58 a_n6972_8799.n107 45.0871
R198 a_n6972_8799.n67 a_n6972_8799.n118 45.0871
R199 a_n6972_8799.n76 a_n6972_8799.n130 45.0871
R200 a_n6972_8799.n38 a_n6972_8799.n141 45.0871
R201 a_n6972_8799.n47 a_n6972_8799.n152 45.0871
R202 a_n6972_8799.n56 a_n6972_8799.n164 45.0871
R203 a_n6972_8799.n2 a_n6972_8799.n0 33.4185
R204 a_n6972_8799.n174 a_n6972_8799.n89 32.0088
R205 a_n6972_8799.n32 a_n6972_8799.n137 11.843
R206 a_n6972_8799.n142 a_n6972_8799.n37 36.139
R207 a_n6972_8799.n41 a_n6972_8799.n148 11.843
R208 a_n6972_8799.n153 a_n6972_8799.n46 36.139
R209 a_n6972_8799.n50 a_n6972_8799.n160 11.843
R210 a_n6972_8799.n165 a_n6972_8799.n55 36.139
R211 a_n6972_8799.n108 a_n6972_8799.n57 36.139
R212 a_n6972_8799.n102 a_n6972_8799.n63 34.4824
R213 a_n6972_8799.n119 a_n6972_8799.n66 36.139
R214 a_n6972_8799.n113 a_n6972_8799.n72 34.4824
R215 a_n6972_8799.n131 a_n6972_8799.n75 36.139
R216 a_n6972_8799.n125 a_n6972_8799.n81 34.4824
R217 a_n6972_8799.n34 a_n6972_8799.n138 35.3134
R218 a_n6972_8799.n43 a_n6972_8799.n149 35.3134
R219 a_n6972_8799.n52 a_n6972_8799.n161 35.3134
R220 a_n6972_8799.n61 a_n6972_8799.n109 35.3134
R221 a_n6972_8799.n110 a_n6972_8799.n61 11.2134
R222 a_n6972_8799.n70 a_n6972_8799.n120 35.3134
R223 a_n6972_8799.n121 a_n6972_8799.n70 11.2134
R224 a_n6972_8799.n79 a_n6972_8799.n132 35.3134
R225 a_n6972_8799.n133 a_n6972_8799.n79 11.2134
R226 a_n6972_8799.n146 a_n6972_8799.n32 34.4824
R227 a_n6972_8799.n37 a_n6972_8799.n139 10.5784
R228 a_n6972_8799.n157 a_n6972_8799.n41 34.4824
R229 a_n6972_8799.n46 a_n6972_8799.n150 10.5784
R230 a_n6972_8799.n169 a_n6972_8799.n50 34.4824
R231 a_n6972_8799.n55 a_n6972_8799.n162 10.5784
R232 a_n6972_8799.n57 a_n6972_8799.n105 10.5784
R233 a_n6972_8799.n66 a_n6972_8799.n116 10.5784
R234 a_n6972_8799.n75 a_n6972_8799.n128 10.5784
R235 a_n6972_8799.n29 a_n6972_8799.n174 18.5874
R236 a_n6972_8799.n141 a_n6972_8799.n140 14.1472
R237 a_n6972_8799.n152 a_n6972_8799.n151 14.1472
R238 a_n6972_8799.n164 a_n6972_8799.n163 14.1472
R239 a_n6972_8799.n107 a_n6972_8799.n106 14.1472
R240 a_n6972_8799.n118 a_n6972_8799.n117 14.1472
R241 a_n6972_8799.n130 a_n6972_8799.n129 14.1472
R242 a_n6972_8799.n173 a_n6972_8799.n1 12.3339
R243 a_n6972_8799.n174 a_n6972_8799.n173 11.4887
R244 a_n6972_8799.n159 a_n6972_8799.n26 9.01755
R245 a_n6972_8799.n124 a_n6972_8799.n12 9.01755
R246 a_n6972_8799.n172 a_n6972_8799.n136 7.00615
R247 a_n6972_8799.n172 a_n6972_8799.n171 6.58471
R248 a_n6972_8799.n159 a_n6972_8799.n22 4.90959
R249 a_n6972_8799.n171 a_n6972_8799.n18 4.90959
R250 a_n6972_8799.n124 a_n6972_8799.n8 4.90959
R251 a_n6972_8799.n136 a_n6972_8799.n4 4.90959
R252 a_n6972_8799.n171 a_n6972_8799.n159 4.10845
R253 a_n6972_8799.n136 a_n6972_8799.n124 4.10845
R254 a_n6972_8799.n175 a_n6972_8799.t35 3.61217
R255 a_n6972_8799.n175 a_n6972_8799.t17 3.61217
R256 a_n6972_8799.n176 a_n6972_8799.t34 3.61217
R257 a_n6972_8799.n176 a_n6972_8799.t30 3.61217
R258 a_n6972_8799.n84 a_n6972_8799.t37 3.61217
R259 a_n6972_8799.n84 a_n6972_8799.t33 3.61217
R260 a_n6972_8799.n85 a_n6972_8799.t36 3.61217
R261 a_n6972_8799.n85 a_n6972_8799.t18 3.61217
R262 a_n6972_8799.n86 a_n6972_8799.t39 3.61217
R263 a_n6972_8799.n86 a_n6972_8799.t32 3.61217
R264 a_n6972_8799.n87 a_n6972_8799.t19 3.61217
R265 a_n6972_8799.n87 a_n6972_8799.t31 3.61217
R266 a_n6972_8799.n88 a_n6972_8799.t29 3.61217
R267 a_n6972_8799.n88 a_n6972_8799.t5 3.61217
R268 a_n6972_8799.t4 a_n6972_8799.n178 3.61217
R269 a_n6972_8799.n178 a_n6972_8799.t6 3.61217
R270 a_n6972_8799.n173 a_n6972_8799.n172 3.4105
R271 a_n6972_8799.n99 a_n6972_8799.t38 2.82907
R272 a_n6972_8799.n99 a_n6972_8799.t13 2.82907
R273 a_n6972_8799.n100 a_n6972_8799.t27 2.82907
R274 a_n6972_8799.n100 a_n6972_8799.t23 2.82907
R275 a_n6972_8799.n101 a_n6972_8799.t12 2.82907
R276 a_n6972_8799.n101 a_n6972_8799.t25 2.82907
R277 a_n6972_8799.n92 a_n6972_8799.t20 2.82907
R278 a_n6972_8799.n92 a_n6972_8799.t11 2.82907
R279 a_n6972_8799.n91 a_n6972_8799.t9 2.82907
R280 a_n6972_8799.n91 a_n6972_8799.t21 2.82907
R281 a_n6972_8799.n90 a_n6972_8799.t2 2.82907
R282 a_n6972_8799.n90 a_n6972_8799.t7 2.82907
R283 a_n6972_8799.n96 a_n6972_8799.t26 2.82907
R284 a_n6972_8799.n96 a_n6972_8799.t0 2.82907
R285 a_n6972_8799.n97 a_n6972_8799.t22 2.82907
R286 a_n6972_8799.n97 a_n6972_8799.t1 2.82907
R287 a_n6972_8799.n98 a_n6972_8799.t28 2.82907
R288 a_n6972_8799.n98 a_n6972_8799.t15 2.82907
R289 a_n6972_8799.n95 a_n6972_8799.t10 2.82907
R290 a_n6972_8799.n95 a_n6972_8799.t3 2.82907
R291 a_n6972_8799.n94 a_n6972_8799.t24 2.82907
R292 a_n6972_8799.n94 a_n6972_8799.t8 2.82907
R293 a_n6972_8799.n93 a_n6972_8799.t14 2.82907
R294 a_n6972_8799.n93 a_n6972_8799.t16 2.82907
R295 a_n6972_8799.n30 a_n6972_8799.n147 22.3251
R296 a_n6972_8799.n39 a_n6972_8799.n158 22.3251
R297 a_n6972_8799.n48 a_n6972_8799.n170 22.3251
R298 a_n6972_8799.n65 a_n6972_8799.n112 22.3251
R299 a_n6972_8799.n74 a_n6972_8799.n123 22.3251
R300 a_n6972_8799.n83 a_n6972_8799.n135 22.3251
R301 a_n6972_8799.n33 a_n6972_8799.n145 0.365327
R302 a_n6972_8799.n143 a_n6972_8799.n36 21.4216
R303 a_n6972_8799.n42 a_n6972_8799.n156 0.365327
R304 a_n6972_8799.n154 a_n6972_8799.n45 21.4216
R305 a_n6972_8799.n51 a_n6972_8799.n168 0.365327
R306 a_n6972_8799.n166 a_n6972_8799.n54 21.4216
R307 a_n6972_8799.n111 a_n6972_8799.n62 47.835
R308 a_n6972_8799.n122 a_n6972_8799.n71 47.835
R309 a_n6972_8799.n134 a_n6972_8799.n80 47.835
R310 a_n6972_8799.n1 a_n6972_8799.n2 1.77636
R311 a_n6972_8799.n0 a_n6972_8799.n3 1.3324
R312 a_n6972_8799.n27 a_n6972_8799.n25 0.758076
R313 a_n6972_8799.n25 a_n6972_8799.n24 0.758076
R314 a_n6972_8799.n38 a_n6972_8799.n24 0.758076
R315 a_n6972_8799.n23 a_n6972_8799.n21 0.758076
R316 a_n6972_8799.n21 a_n6972_8799.n20 0.758076
R317 a_n6972_8799.n47 a_n6972_8799.n20 0.758076
R318 a_n6972_8799.n19 a_n6972_8799.n17 0.758076
R319 a_n6972_8799.n17 a_n6972_8799.n16 0.758076
R320 a_n6972_8799.n56 a_n6972_8799.n16 0.758076
R321 a_n6972_8799.n15 a_n6972_8799.n14 0.758076
R322 a_n6972_8799.n14 a_n6972_8799.n13 0.758076
R323 a_n6972_8799.n13 a_n6972_8799.n12 0.758076
R324 a_n6972_8799.n11 a_n6972_8799.n10 0.758076
R325 a_n6972_8799.n10 a_n6972_8799.n9 0.758076
R326 a_n6972_8799.n9 a_n6972_8799.n8 0.758076
R327 a_n6972_8799.n7 a_n6972_8799.n6 0.758076
R328 a_n6972_8799.n6 a_n6972_8799.n5 0.758076
R329 a_n6972_8799.n5 a_n6972_8799.n4 0.758076
R330 a_n6972_8799.n177 a_n6972_8799.n29 0.716017
R331 a_n6972_8799.n89 a_n6972_8799.n28 0.716017
R332 a_n6972_8799.n76 a_n6972_8799.n7 0.568682
R333 a_n6972_8799.n67 a_n6972_8799.n11 0.568682
R334 a_n6972_8799.n58 a_n6972_8799.n15 0.568682
R335 a_n6972_8799.n19 a_n6972_8799.n18 0.568682
R336 a_n6972_8799.n23 a_n6972_8799.n22 0.568682
R337 a_n6972_8799.n27 a_n6972_8799.n26 0.568682
R338 vdd.n303 vdd.n267 756.745
R339 vdd.n252 vdd.n216 756.745
R340 vdd.n209 vdd.n173 756.745
R341 vdd.n158 vdd.n122 756.745
R342 vdd.n116 vdd.n80 756.745
R343 vdd.n65 vdd.n29 756.745
R344 vdd.n1860 vdd.n1824 756.745
R345 vdd.n1911 vdd.n1875 756.745
R346 vdd.n1766 vdd.n1730 756.745
R347 vdd.n1817 vdd.n1781 756.745
R348 vdd.n1673 vdd.n1637 756.745
R349 vdd.n1724 vdd.n1688 756.745
R350 vdd.n1081 vdd.t35 640.208
R351 vdd.n809 vdd.t77 640.208
R352 vdd.n1101 vdd.t61 640.208
R353 vdd.n800 vdd.t95 640.208
R354 vdd.n700 vdd.t64 640.208
R355 vdd.n2416 vdd.t89 640.208
R356 vdd.n661 vdd.t101 640.208
R357 vdd.n2413 vdd.t81 640.208
R358 vdd.n625 vdd.t31 640.208
R359 vdd.n871 vdd.t85 640.208
R360 vdd.n1472 vdd.t51 592.009
R361 vdd.n1509 vdd.t58 592.009
R362 vdd.n1383 vdd.t71 592.009
R363 vdd.n1981 vdd.t43 592.009
R364 vdd.n1018 vdd.t74 592.009
R365 vdd.n978 vdd.t92 592.009
R366 vdd.n3113 vdd.t47 592.009
R367 vdd.n427 vdd.t98 592.009
R368 vdd.n387 vdd.t104 592.009
R369 vdd.n580 vdd.t55 592.009
R370 vdd.n543 vdd.t68 592.009
R371 vdd.n2900 vdd.t39 592.009
R372 vdd.n304 vdd.n303 585
R373 vdd.n302 vdd.n269 585
R374 vdd.n301 vdd.n300 585
R375 vdd.n272 vdd.n270 585
R376 vdd.n295 vdd.n294 585
R377 vdd.n293 vdd.n292 585
R378 vdd.n276 vdd.n275 585
R379 vdd.n287 vdd.n286 585
R380 vdd.n285 vdd.n284 585
R381 vdd.n280 vdd.n279 585
R382 vdd.n253 vdd.n252 585
R383 vdd.n251 vdd.n218 585
R384 vdd.n250 vdd.n249 585
R385 vdd.n221 vdd.n219 585
R386 vdd.n244 vdd.n243 585
R387 vdd.n242 vdd.n241 585
R388 vdd.n225 vdd.n224 585
R389 vdd.n236 vdd.n235 585
R390 vdd.n234 vdd.n233 585
R391 vdd.n229 vdd.n228 585
R392 vdd.n210 vdd.n209 585
R393 vdd.n208 vdd.n175 585
R394 vdd.n207 vdd.n206 585
R395 vdd.n178 vdd.n176 585
R396 vdd.n201 vdd.n200 585
R397 vdd.n199 vdd.n198 585
R398 vdd.n182 vdd.n181 585
R399 vdd.n193 vdd.n192 585
R400 vdd.n191 vdd.n190 585
R401 vdd.n186 vdd.n185 585
R402 vdd.n159 vdd.n158 585
R403 vdd.n157 vdd.n124 585
R404 vdd.n156 vdd.n155 585
R405 vdd.n127 vdd.n125 585
R406 vdd.n150 vdd.n149 585
R407 vdd.n148 vdd.n147 585
R408 vdd.n131 vdd.n130 585
R409 vdd.n142 vdd.n141 585
R410 vdd.n140 vdd.n139 585
R411 vdd.n135 vdd.n134 585
R412 vdd.n117 vdd.n116 585
R413 vdd.n115 vdd.n82 585
R414 vdd.n114 vdd.n113 585
R415 vdd.n85 vdd.n83 585
R416 vdd.n108 vdd.n107 585
R417 vdd.n106 vdd.n105 585
R418 vdd.n89 vdd.n88 585
R419 vdd.n100 vdd.n99 585
R420 vdd.n98 vdd.n97 585
R421 vdd.n93 vdd.n92 585
R422 vdd.n66 vdd.n65 585
R423 vdd.n64 vdd.n31 585
R424 vdd.n63 vdd.n62 585
R425 vdd.n34 vdd.n32 585
R426 vdd.n57 vdd.n56 585
R427 vdd.n55 vdd.n54 585
R428 vdd.n38 vdd.n37 585
R429 vdd.n49 vdd.n48 585
R430 vdd.n47 vdd.n46 585
R431 vdd.n42 vdd.n41 585
R432 vdd.n1861 vdd.n1860 585
R433 vdd.n1859 vdd.n1826 585
R434 vdd.n1858 vdd.n1857 585
R435 vdd.n1829 vdd.n1827 585
R436 vdd.n1852 vdd.n1851 585
R437 vdd.n1850 vdd.n1849 585
R438 vdd.n1833 vdd.n1832 585
R439 vdd.n1844 vdd.n1843 585
R440 vdd.n1842 vdd.n1841 585
R441 vdd.n1837 vdd.n1836 585
R442 vdd.n1912 vdd.n1911 585
R443 vdd.n1910 vdd.n1877 585
R444 vdd.n1909 vdd.n1908 585
R445 vdd.n1880 vdd.n1878 585
R446 vdd.n1903 vdd.n1902 585
R447 vdd.n1901 vdd.n1900 585
R448 vdd.n1884 vdd.n1883 585
R449 vdd.n1895 vdd.n1894 585
R450 vdd.n1893 vdd.n1892 585
R451 vdd.n1888 vdd.n1887 585
R452 vdd.n1767 vdd.n1766 585
R453 vdd.n1765 vdd.n1732 585
R454 vdd.n1764 vdd.n1763 585
R455 vdd.n1735 vdd.n1733 585
R456 vdd.n1758 vdd.n1757 585
R457 vdd.n1756 vdd.n1755 585
R458 vdd.n1739 vdd.n1738 585
R459 vdd.n1750 vdd.n1749 585
R460 vdd.n1748 vdd.n1747 585
R461 vdd.n1743 vdd.n1742 585
R462 vdd.n1818 vdd.n1817 585
R463 vdd.n1816 vdd.n1783 585
R464 vdd.n1815 vdd.n1814 585
R465 vdd.n1786 vdd.n1784 585
R466 vdd.n1809 vdd.n1808 585
R467 vdd.n1807 vdd.n1806 585
R468 vdd.n1790 vdd.n1789 585
R469 vdd.n1801 vdd.n1800 585
R470 vdd.n1799 vdd.n1798 585
R471 vdd.n1794 vdd.n1793 585
R472 vdd.n1674 vdd.n1673 585
R473 vdd.n1672 vdd.n1639 585
R474 vdd.n1671 vdd.n1670 585
R475 vdd.n1642 vdd.n1640 585
R476 vdd.n1665 vdd.n1664 585
R477 vdd.n1663 vdd.n1662 585
R478 vdd.n1646 vdd.n1645 585
R479 vdd.n1657 vdd.n1656 585
R480 vdd.n1655 vdd.n1654 585
R481 vdd.n1650 vdd.n1649 585
R482 vdd.n1725 vdd.n1724 585
R483 vdd.n1723 vdd.n1690 585
R484 vdd.n1722 vdd.n1721 585
R485 vdd.n1693 vdd.n1691 585
R486 vdd.n1716 vdd.n1715 585
R487 vdd.n1714 vdd.n1713 585
R488 vdd.n1697 vdd.n1696 585
R489 vdd.n1708 vdd.n1707 585
R490 vdd.n1706 vdd.n1705 585
R491 vdd.n1701 vdd.n1700 585
R492 vdd.n3229 vdd.n352 488.781
R493 vdd.n3111 vdd.n350 488.781
R494 vdd.n3033 vdd.n515 488.781
R495 vdd.n3031 vdd.n517 488.781
R496 vdd.n1976 vdd.n1265 488.781
R497 vdd.n1979 vdd.n1978 488.781
R498 vdd.n1578 vdd.n1343 488.781
R499 vdd.n1576 vdd.n1346 488.781
R500 vdd.n281 vdd.t219 329.043
R501 vdd.n230 vdd.t201 329.043
R502 vdd.n187 vdd.t210 329.043
R503 vdd.n136 vdd.t193 329.043
R504 vdd.n94 vdd.t160 329.043
R505 vdd.n43 vdd.t167 329.043
R506 vdd.n1838 vdd.t225 329.043
R507 vdd.n1889 vdd.t163 329.043
R508 vdd.n1744 vdd.t216 329.043
R509 vdd.n1795 vdd.t149 329.043
R510 vdd.n1651 vdd.t169 329.043
R511 vdd.n1702 vdd.t161 329.043
R512 vdd.n1472 vdd.t54 319.788
R513 vdd.n1509 vdd.t60 319.788
R514 vdd.n1383 vdd.t73 319.788
R515 vdd.n1981 vdd.t45 319.788
R516 vdd.n1018 vdd.t75 319.788
R517 vdd.n978 vdd.t93 319.788
R518 vdd.n3113 vdd.t49 319.788
R519 vdd.n427 vdd.t99 319.788
R520 vdd.n387 vdd.t105 319.788
R521 vdd.n580 vdd.t57 319.788
R522 vdd.n543 vdd.t70 319.788
R523 vdd.n2900 vdd.t42 319.788
R524 vdd.n1473 vdd.t53 303.69
R525 vdd.n1510 vdd.t59 303.69
R526 vdd.n1384 vdd.t72 303.69
R527 vdd.n1982 vdd.t46 303.69
R528 vdd.n1019 vdd.t76 303.69
R529 vdd.n979 vdd.t94 303.69
R530 vdd.n3114 vdd.t50 303.69
R531 vdd.n428 vdd.t100 303.69
R532 vdd.n388 vdd.t106 303.69
R533 vdd.n581 vdd.t56 303.69
R534 vdd.n544 vdd.t69 303.69
R535 vdd.n2901 vdd.t41 303.69
R536 vdd.n2648 vdd.n755 291.221
R537 vdd.n2862 vdd.n635 291.221
R538 vdd.n2799 vdd.n632 291.221
R539 vdd.n2580 vdd.n2579 291.221
R540 vdd.n2376 vdd.n797 291.221
R541 vdd.n2307 vdd.n2306 291.221
R542 vdd.n1137 vdd.n1136 291.221
R543 vdd.n2127 vdd.n903 291.221
R544 vdd.n2778 vdd.n633 291.221
R545 vdd.n2865 vdd.n2864 291.221
R546 vdd.n2484 vdd.n2410 291.221
R547 vdd.n2652 vdd.n759 291.221
R548 vdd.n2304 vdd.n807 291.221
R549 vdd.n805 vdd.n779 291.221
R550 vdd.n1215 vdd.n944 291.221
R551 vdd.n2131 vdd.n908 291.221
R552 vdd.n2780 vdd.n633 185
R553 vdd.n2863 vdd.n633 185
R554 vdd.n2782 vdd.n2781 185
R555 vdd.n2781 vdd.n631 185
R556 vdd.n2783 vdd.n667 185
R557 vdd.n2793 vdd.n667 185
R558 vdd.n2784 vdd.n676 185
R559 vdd.n676 vdd.n674 185
R560 vdd.n2786 vdd.n2785 185
R561 vdd.n2787 vdd.n2786 185
R562 vdd.n2739 vdd.n675 185
R563 vdd.n675 vdd.n671 185
R564 vdd.n2738 vdd.n2737 185
R565 vdd.n2737 vdd.n2736 185
R566 vdd.n678 vdd.n677 185
R567 vdd.n679 vdd.n678 185
R568 vdd.n2729 vdd.n2728 185
R569 vdd.n2730 vdd.n2729 185
R570 vdd.n2727 vdd.n688 185
R571 vdd.n688 vdd.n685 185
R572 vdd.n2726 vdd.n2725 185
R573 vdd.n2725 vdd.n2724 185
R574 vdd.n690 vdd.n689 185
R575 vdd.n698 vdd.n690 185
R576 vdd.n2717 vdd.n2716 185
R577 vdd.n2718 vdd.n2717 185
R578 vdd.n2714 vdd.n699 185
R579 vdd.n706 vdd.n699 185
R580 vdd.n2713 vdd.n2712 185
R581 vdd.n2712 vdd.n2711 185
R582 vdd.n702 vdd.n701 185
R583 vdd.n703 vdd.n702 185
R584 vdd.n2704 vdd.n2703 185
R585 vdd.n2705 vdd.n2704 185
R586 vdd.n2702 vdd.n713 185
R587 vdd.n713 vdd.n710 185
R588 vdd.n2701 vdd.n2700 185
R589 vdd.n2700 vdd.n2699 185
R590 vdd.n715 vdd.n714 185
R591 vdd.n723 vdd.n715 185
R592 vdd.n2692 vdd.n2691 185
R593 vdd.n2693 vdd.n2692 185
R594 vdd.n2690 vdd.n724 185
R595 vdd.n729 vdd.n724 185
R596 vdd.n2689 vdd.n2688 185
R597 vdd.n2688 vdd.n2687 185
R598 vdd.n726 vdd.n725 185
R599 vdd.n2559 vdd.n726 185
R600 vdd.n2680 vdd.n2679 185
R601 vdd.n2681 vdd.n2680 185
R602 vdd.n2678 vdd.n736 185
R603 vdd.n736 vdd.n733 185
R604 vdd.n2677 vdd.n2676 185
R605 vdd.n2676 vdd.n2675 185
R606 vdd.n738 vdd.n737 185
R607 vdd.n739 vdd.n738 185
R608 vdd.n2668 vdd.n2667 185
R609 vdd.n2669 vdd.n2668 185
R610 vdd.n2666 vdd.n748 185
R611 vdd.n748 vdd.n745 185
R612 vdd.n2665 vdd.n2664 185
R613 vdd.n2664 vdd.n2663 185
R614 vdd.n750 vdd.n749 185
R615 vdd.n2574 vdd.n750 185
R616 vdd.n2656 vdd.n2655 185
R617 vdd.n2657 vdd.n2656 185
R618 vdd.n2654 vdd.n759 185
R619 vdd.n759 vdd.n756 185
R620 vdd.n2653 vdd.n2652 185
R621 vdd.n761 vdd.n760 185
R622 vdd.n2420 vdd.n2419 185
R623 vdd.n2422 vdd.n2421 185
R624 vdd.n2424 vdd.n2423 185
R625 vdd.n2426 vdd.n2425 185
R626 vdd.n2428 vdd.n2427 185
R627 vdd.n2430 vdd.n2429 185
R628 vdd.n2432 vdd.n2431 185
R629 vdd.n2434 vdd.n2433 185
R630 vdd.n2436 vdd.n2435 185
R631 vdd.n2438 vdd.n2437 185
R632 vdd.n2440 vdd.n2439 185
R633 vdd.n2442 vdd.n2441 185
R634 vdd.n2444 vdd.n2443 185
R635 vdd.n2446 vdd.n2445 185
R636 vdd.n2448 vdd.n2447 185
R637 vdd.n2450 vdd.n2449 185
R638 vdd.n2452 vdd.n2451 185
R639 vdd.n2454 vdd.n2453 185
R640 vdd.n2456 vdd.n2455 185
R641 vdd.n2458 vdd.n2457 185
R642 vdd.n2460 vdd.n2459 185
R643 vdd.n2462 vdd.n2461 185
R644 vdd.n2464 vdd.n2463 185
R645 vdd.n2466 vdd.n2465 185
R646 vdd.n2468 vdd.n2467 185
R647 vdd.n2470 vdd.n2469 185
R648 vdd.n2472 vdd.n2471 185
R649 vdd.n2474 vdd.n2473 185
R650 vdd.n2476 vdd.n2475 185
R651 vdd.n2478 vdd.n2477 185
R652 vdd.n2480 vdd.n2479 185
R653 vdd.n2482 vdd.n2481 185
R654 vdd.n2483 vdd.n2410 185
R655 vdd.n2650 vdd.n2410 185
R656 vdd.n2866 vdd.n2865 185
R657 vdd.n2867 vdd.n624 185
R658 vdd.n2869 vdd.n2868 185
R659 vdd.n2871 vdd.n622 185
R660 vdd.n2873 vdd.n2872 185
R661 vdd.n2874 vdd.n621 185
R662 vdd.n2876 vdd.n2875 185
R663 vdd.n2878 vdd.n619 185
R664 vdd.n2880 vdd.n2879 185
R665 vdd.n2881 vdd.n618 185
R666 vdd.n2883 vdd.n2882 185
R667 vdd.n2885 vdd.n616 185
R668 vdd.n2887 vdd.n2886 185
R669 vdd.n2888 vdd.n615 185
R670 vdd.n2890 vdd.n2889 185
R671 vdd.n2892 vdd.n614 185
R672 vdd.n2893 vdd.n611 185
R673 vdd.n2896 vdd.n2895 185
R674 vdd.n612 vdd.n610 185
R675 vdd.n2752 vdd.n2751 185
R676 vdd.n2754 vdd.n2753 185
R677 vdd.n2756 vdd.n2748 185
R678 vdd.n2758 vdd.n2757 185
R679 vdd.n2759 vdd.n2747 185
R680 vdd.n2761 vdd.n2760 185
R681 vdd.n2763 vdd.n2745 185
R682 vdd.n2765 vdd.n2764 185
R683 vdd.n2766 vdd.n2744 185
R684 vdd.n2768 vdd.n2767 185
R685 vdd.n2770 vdd.n2742 185
R686 vdd.n2772 vdd.n2771 185
R687 vdd.n2773 vdd.n2741 185
R688 vdd.n2775 vdd.n2774 185
R689 vdd.n2777 vdd.n2740 185
R690 vdd.n2779 vdd.n2778 185
R691 vdd.n2778 vdd.n613 185
R692 vdd.n2864 vdd.n628 185
R693 vdd.n2864 vdd.n2863 185
R694 vdd.n2487 vdd.n630 185
R695 vdd.n631 vdd.n630 185
R696 vdd.n2488 vdd.n666 185
R697 vdd.n2793 vdd.n666 185
R698 vdd.n2490 vdd.n2489 185
R699 vdd.n2489 vdd.n674 185
R700 vdd.n2491 vdd.n673 185
R701 vdd.n2787 vdd.n673 185
R702 vdd.n2493 vdd.n2492 185
R703 vdd.n2492 vdd.n671 185
R704 vdd.n2494 vdd.n681 185
R705 vdd.n2736 vdd.n681 185
R706 vdd.n2496 vdd.n2495 185
R707 vdd.n2495 vdd.n679 185
R708 vdd.n2497 vdd.n687 185
R709 vdd.n2730 vdd.n687 185
R710 vdd.n2499 vdd.n2498 185
R711 vdd.n2498 vdd.n685 185
R712 vdd.n2500 vdd.n692 185
R713 vdd.n2724 vdd.n692 185
R714 vdd.n2502 vdd.n2501 185
R715 vdd.n2501 vdd.n698 185
R716 vdd.n2503 vdd.n697 185
R717 vdd.n2718 vdd.n697 185
R718 vdd.n2505 vdd.n2504 185
R719 vdd.n2504 vdd.n706 185
R720 vdd.n2506 vdd.n705 185
R721 vdd.n2711 vdd.n705 185
R722 vdd.n2508 vdd.n2507 185
R723 vdd.n2507 vdd.n703 185
R724 vdd.n2509 vdd.n712 185
R725 vdd.n2705 vdd.n712 185
R726 vdd.n2511 vdd.n2510 185
R727 vdd.n2510 vdd.n710 185
R728 vdd.n2512 vdd.n717 185
R729 vdd.n2699 vdd.n717 185
R730 vdd.n2514 vdd.n2513 185
R731 vdd.n2513 vdd.n723 185
R732 vdd.n2515 vdd.n722 185
R733 vdd.n2693 vdd.n722 185
R734 vdd.n2517 vdd.n2516 185
R735 vdd.n2516 vdd.n729 185
R736 vdd.n2518 vdd.n728 185
R737 vdd.n2687 vdd.n728 185
R738 vdd.n2561 vdd.n2560 185
R739 vdd.n2560 vdd.n2559 185
R740 vdd.n2562 vdd.n735 185
R741 vdd.n2681 vdd.n735 185
R742 vdd.n2564 vdd.n2563 185
R743 vdd.n2563 vdd.n733 185
R744 vdd.n2565 vdd.n741 185
R745 vdd.n2675 vdd.n741 185
R746 vdd.n2567 vdd.n2566 185
R747 vdd.n2566 vdd.n739 185
R748 vdd.n2568 vdd.n747 185
R749 vdd.n2669 vdd.n747 185
R750 vdd.n2570 vdd.n2569 185
R751 vdd.n2569 vdd.n745 185
R752 vdd.n2571 vdd.n752 185
R753 vdd.n2663 vdd.n752 185
R754 vdd.n2573 vdd.n2572 185
R755 vdd.n2574 vdd.n2573 185
R756 vdd.n2486 vdd.n758 185
R757 vdd.n2657 vdd.n758 185
R758 vdd.n2485 vdd.n2484 185
R759 vdd.n2484 vdd.n756 185
R760 vdd.n1976 vdd.n1975 185
R761 vdd.n1977 vdd.n1976 185
R762 vdd.n1266 vdd.n1264 185
R763 vdd.n1968 vdd.n1264 185
R764 vdd.n1971 vdd.n1970 185
R765 vdd.n1970 vdd.n1969 185
R766 vdd.n1269 vdd.n1268 185
R767 vdd.n1270 vdd.n1269 185
R768 vdd.n1957 vdd.n1956 185
R769 vdd.n1958 vdd.n1957 185
R770 vdd.n1278 vdd.n1277 185
R771 vdd.n1949 vdd.n1277 185
R772 vdd.n1952 vdd.n1951 185
R773 vdd.n1951 vdd.n1950 185
R774 vdd.n1281 vdd.n1280 185
R775 vdd.n1287 vdd.n1281 185
R776 vdd.n1940 vdd.n1939 185
R777 vdd.n1941 vdd.n1940 185
R778 vdd.n1289 vdd.n1288 185
R779 vdd.n1932 vdd.n1288 185
R780 vdd.n1935 vdd.n1934 185
R781 vdd.n1934 vdd.n1933 185
R782 vdd.n1292 vdd.n1291 185
R783 vdd.n1293 vdd.n1292 185
R784 vdd.n1923 vdd.n1922 185
R785 vdd.n1924 vdd.n1923 185
R786 vdd.n1301 vdd.n1300 185
R787 vdd.n1300 vdd.n1299 185
R788 vdd.n1636 vdd.n1635 185
R789 vdd.n1635 vdd.n1634 185
R790 vdd.n1304 vdd.n1303 185
R791 vdd.n1310 vdd.n1304 185
R792 vdd.n1625 vdd.n1624 185
R793 vdd.n1626 vdd.n1625 185
R794 vdd.n1312 vdd.n1311 185
R795 vdd.n1617 vdd.n1311 185
R796 vdd.n1620 vdd.n1619 185
R797 vdd.n1619 vdd.n1618 185
R798 vdd.n1315 vdd.n1314 185
R799 vdd.n1322 vdd.n1315 185
R800 vdd.n1608 vdd.n1607 185
R801 vdd.n1609 vdd.n1608 185
R802 vdd.n1324 vdd.n1323 185
R803 vdd.n1323 vdd.n1321 185
R804 vdd.n1603 vdd.n1602 185
R805 vdd.n1602 vdd.n1601 185
R806 vdd.n1327 vdd.n1326 185
R807 vdd.n1328 vdd.n1327 185
R808 vdd.n1592 vdd.n1591 185
R809 vdd.n1593 vdd.n1592 185
R810 vdd.n1336 vdd.n1335 185
R811 vdd.n1335 vdd.n1334 185
R812 vdd.n1587 vdd.n1586 185
R813 vdd.n1586 vdd.n1585 185
R814 vdd.n1339 vdd.n1338 185
R815 vdd.n1345 vdd.n1339 185
R816 vdd.n1576 vdd.n1575 185
R817 vdd.n1577 vdd.n1576 185
R818 vdd.n1572 vdd.n1346 185
R819 vdd.n1571 vdd.n1349 185
R820 vdd.n1570 vdd.n1350 185
R821 vdd.n1350 vdd.n1344 185
R822 vdd.n1353 vdd.n1351 185
R823 vdd.n1566 vdd.n1355 185
R824 vdd.n1565 vdd.n1356 185
R825 vdd.n1564 vdd.n1358 185
R826 vdd.n1361 vdd.n1359 185
R827 vdd.n1560 vdd.n1363 185
R828 vdd.n1559 vdd.n1364 185
R829 vdd.n1558 vdd.n1366 185
R830 vdd.n1369 vdd.n1367 185
R831 vdd.n1554 vdd.n1371 185
R832 vdd.n1553 vdd.n1372 185
R833 vdd.n1552 vdd.n1374 185
R834 vdd.n1377 vdd.n1375 185
R835 vdd.n1548 vdd.n1379 185
R836 vdd.n1547 vdd.n1380 185
R837 vdd.n1546 vdd.n1382 185
R838 vdd.n1387 vdd.n1385 185
R839 vdd.n1542 vdd.n1389 185
R840 vdd.n1541 vdd.n1390 185
R841 vdd.n1540 vdd.n1392 185
R842 vdd.n1395 vdd.n1393 185
R843 vdd.n1536 vdd.n1397 185
R844 vdd.n1535 vdd.n1398 185
R845 vdd.n1534 vdd.n1400 185
R846 vdd.n1403 vdd.n1401 185
R847 vdd.n1530 vdd.n1405 185
R848 vdd.n1529 vdd.n1406 185
R849 vdd.n1528 vdd.n1408 185
R850 vdd.n1411 vdd.n1409 185
R851 vdd.n1524 vdd.n1413 185
R852 vdd.n1523 vdd.n1414 185
R853 vdd.n1522 vdd.n1416 185
R854 vdd.n1419 vdd.n1417 185
R855 vdd.n1518 vdd.n1421 185
R856 vdd.n1517 vdd.n1422 185
R857 vdd.n1516 vdd.n1424 185
R858 vdd.n1427 vdd.n1425 185
R859 vdd.n1512 vdd.n1429 185
R860 vdd.n1511 vdd.n1508 185
R861 vdd.n1506 vdd.n1430 185
R862 vdd.n1505 vdd.n1504 185
R863 vdd.n1435 vdd.n1432 185
R864 vdd.n1500 vdd.n1436 185
R865 vdd.n1499 vdd.n1438 185
R866 vdd.n1498 vdd.n1439 185
R867 vdd.n1443 vdd.n1440 185
R868 vdd.n1494 vdd.n1444 185
R869 vdd.n1493 vdd.n1446 185
R870 vdd.n1492 vdd.n1447 185
R871 vdd.n1451 vdd.n1448 185
R872 vdd.n1488 vdd.n1452 185
R873 vdd.n1487 vdd.n1454 185
R874 vdd.n1486 vdd.n1455 185
R875 vdd.n1459 vdd.n1456 185
R876 vdd.n1482 vdd.n1460 185
R877 vdd.n1481 vdd.n1462 185
R878 vdd.n1480 vdd.n1463 185
R879 vdd.n1467 vdd.n1464 185
R880 vdd.n1476 vdd.n1468 185
R881 vdd.n1475 vdd.n1470 185
R882 vdd.n1471 vdd.n1343 185
R883 vdd.n1344 vdd.n1343 185
R884 vdd.n1980 vdd.n1979 185
R885 vdd.n1984 vdd.n1260 185
R886 vdd.n1259 vdd.n1253 185
R887 vdd.n1257 vdd.n1256 185
R888 vdd.n1255 vdd.n1049 185
R889 vdd.n1988 vdd.n1046 185
R890 vdd.n1990 vdd.n1989 185
R891 vdd.n1992 vdd.n1044 185
R892 vdd.n1994 vdd.n1993 185
R893 vdd.n1995 vdd.n1039 185
R894 vdd.n1997 vdd.n1996 185
R895 vdd.n1999 vdd.n1037 185
R896 vdd.n2001 vdd.n2000 185
R897 vdd.n2002 vdd.n1032 185
R898 vdd.n2004 vdd.n2003 185
R899 vdd.n2006 vdd.n1030 185
R900 vdd.n2008 vdd.n2007 185
R901 vdd.n2009 vdd.n1026 185
R902 vdd.n2011 vdd.n2010 185
R903 vdd.n2013 vdd.n1023 185
R904 vdd.n2015 vdd.n2014 185
R905 vdd.n1024 vdd.n1017 185
R906 vdd.n2019 vdd.n1021 185
R907 vdd.n2020 vdd.n1013 185
R908 vdd.n2022 vdd.n2021 185
R909 vdd.n2024 vdd.n1011 185
R910 vdd.n2026 vdd.n2025 185
R911 vdd.n2027 vdd.n1006 185
R912 vdd.n2029 vdd.n2028 185
R913 vdd.n2031 vdd.n1004 185
R914 vdd.n2033 vdd.n2032 185
R915 vdd.n2034 vdd.n999 185
R916 vdd.n2036 vdd.n2035 185
R917 vdd.n2038 vdd.n997 185
R918 vdd.n2040 vdd.n2039 185
R919 vdd.n2041 vdd.n992 185
R920 vdd.n2043 vdd.n2042 185
R921 vdd.n2045 vdd.n990 185
R922 vdd.n2047 vdd.n2046 185
R923 vdd.n2048 vdd.n986 185
R924 vdd.n2050 vdd.n2049 185
R925 vdd.n2052 vdd.n983 185
R926 vdd.n2054 vdd.n2053 185
R927 vdd.n984 vdd.n977 185
R928 vdd.n2058 vdd.n981 185
R929 vdd.n2059 vdd.n973 185
R930 vdd.n2061 vdd.n2060 185
R931 vdd.n2063 vdd.n971 185
R932 vdd.n2065 vdd.n2064 185
R933 vdd.n2066 vdd.n966 185
R934 vdd.n2068 vdd.n2067 185
R935 vdd.n2070 vdd.n964 185
R936 vdd.n2072 vdd.n2071 185
R937 vdd.n2073 vdd.n959 185
R938 vdd.n2075 vdd.n2074 185
R939 vdd.n2077 vdd.n957 185
R940 vdd.n2079 vdd.n2078 185
R941 vdd.n2080 vdd.n955 185
R942 vdd.n2082 vdd.n2081 185
R943 vdd.n2085 vdd.n2084 185
R944 vdd.n2087 vdd.n2086 185
R945 vdd.n2089 vdd.n953 185
R946 vdd.n2091 vdd.n2090 185
R947 vdd.n1265 vdd.n952 185
R948 vdd.n1978 vdd.n1263 185
R949 vdd.n1978 vdd.n1977 185
R950 vdd.n1273 vdd.n1262 185
R951 vdd.n1968 vdd.n1262 185
R952 vdd.n1967 vdd.n1966 185
R953 vdd.n1969 vdd.n1967 185
R954 vdd.n1272 vdd.n1271 185
R955 vdd.n1271 vdd.n1270 185
R956 vdd.n1960 vdd.n1959 185
R957 vdd.n1959 vdd.n1958 185
R958 vdd.n1276 vdd.n1275 185
R959 vdd.n1949 vdd.n1276 185
R960 vdd.n1948 vdd.n1947 185
R961 vdd.n1950 vdd.n1948 185
R962 vdd.n1283 vdd.n1282 185
R963 vdd.n1287 vdd.n1282 185
R964 vdd.n1943 vdd.n1942 185
R965 vdd.n1942 vdd.n1941 185
R966 vdd.n1286 vdd.n1285 185
R967 vdd.n1932 vdd.n1286 185
R968 vdd.n1931 vdd.n1930 185
R969 vdd.n1933 vdd.n1931 185
R970 vdd.n1295 vdd.n1294 185
R971 vdd.n1294 vdd.n1293 185
R972 vdd.n1926 vdd.n1925 185
R973 vdd.n1925 vdd.n1924 185
R974 vdd.n1298 vdd.n1297 185
R975 vdd.n1299 vdd.n1298 185
R976 vdd.n1633 vdd.n1632 185
R977 vdd.n1634 vdd.n1633 185
R978 vdd.n1306 vdd.n1305 185
R979 vdd.n1310 vdd.n1305 185
R980 vdd.n1628 vdd.n1627 185
R981 vdd.n1627 vdd.n1626 185
R982 vdd.n1309 vdd.n1308 185
R983 vdd.n1617 vdd.n1309 185
R984 vdd.n1616 vdd.n1615 185
R985 vdd.n1618 vdd.n1616 185
R986 vdd.n1317 vdd.n1316 185
R987 vdd.n1322 vdd.n1316 185
R988 vdd.n1611 vdd.n1610 185
R989 vdd.n1610 vdd.n1609 185
R990 vdd.n1320 vdd.n1319 185
R991 vdd.n1321 vdd.n1320 185
R992 vdd.n1600 vdd.n1599 185
R993 vdd.n1601 vdd.n1600 185
R994 vdd.n1330 vdd.n1329 185
R995 vdd.n1329 vdd.n1328 185
R996 vdd.n1595 vdd.n1594 185
R997 vdd.n1594 vdd.n1593 185
R998 vdd.n1333 vdd.n1332 185
R999 vdd.n1334 vdd.n1333 185
R1000 vdd.n1584 vdd.n1583 185
R1001 vdd.n1585 vdd.n1584 185
R1002 vdd.n1341 vdd.n1340 185
R1003 vdd.n1345 vdd.n1340 185
R1004 vdd.n1579 vdd.n1578 185
R1005 vdd.n1578 vdd.n1577 185
R1006 vdd.n799 vdd.n797 185
R1007 vdd.n2305 vdd.n797 185
R1008 vdd.n2227 vdd.n817 185
R1009 vdd.n817 vdd.n804 185
R1010 vdd.n2229 vdd.n2228 185
R1011 vdd.n2230 vdd.n2229 185
R1012 vdd.n2226 vdd.n816 185
R1013 vdd.n1166 vdd.n816 185
R1014 vdd.n2225 vdd.n2224 185
R1015 vdd.n2224 vdd.n2223 185
R1016 vdd.n819 vdd.n818 185
R1017 vdd.n820 vdd.n819 185
R1018 vdd.n2214 vdd.n2213 185
R1019 vdd.n2215 vdd.n2214 185
R1020 vdd.n2212 vdd.n830 185
R1021 vdd.n830 vdd.n827 185
R1022 vdd.n2211 vdd.n2210 185
R1023 vdd.n2210 vdd.n2209 185
R1024 vdd.n832 vdd.n831 185
R1025 vdd.n833 vdd.n832 185
R1026 vdd.n2202 vdd.n2201 185
R1027 vdd.n2203 vdd.n2202 185
R1028 vdd.n2200 vdd.n841 185
R1029 vdd.n846 vdd.n841 185
R1030 vdd.n2199 vdd.n2198 185
R1031 vdd.n2198 vdd.n2197 185
R1032 vdd.n843 vdd.n842 185
R1033 vdd.n852 vdd.n843 185
R1034 vdd.n2190 vdd.n2189 185
R1035 vdd.n2191 vdd.n2190 185
R1036 vdd.n2188 vdd.n853 185
R1037 vdd.n1187 vdd.n853 185
R1038 vdd.n2187 vdd.n2186 185
R1039 vdd.n2186 vdd.n2185 185
R1040 vdd.n855 vdd.n854 185
R1041 vdd.n856 vdd.n855 185
R1042 vdd.n2178 vdd.n2177 185
R1043 vdd.n2179 vdd.n2178 185
R1044 vdd.n2176 vdd.n865 185
R1045 vdd.n865 vdd.n862 185
R1046 vdd.n2175 vdd.n2174 185
R1047 vdd.n2174 vdd.n2173 185
R1048 vdd.n867 vdd.n866 185
R1049 vdd.n876 vdd.n867 185
R1050 vdd.n2165 vdd.n2164 185
R1051 vdd.n2166 vdd.n2165 185
R1052 vdd.n2163 vdd.n877 185
R1053 vdd.n883 vdd.n877 185
R1054 vdd.n2162 vdd.n2161 185
R1055 vdd.n2161 vdd.n2160 185
R1056 vdd.n879 vdd.n878 185
R1057 vdd.n880 vdd.n879 185
R1058 vdd.n2153 vdd.n2152 185
R1059 vdd.n2154 vdd.n2153 185
R1060 vdd.n2151 vdd.n890 185
R1061 vdd.n890 vdd.n887 185
R1062 vdd.n2150 vdd.n2149 185
R1063 vdd.n2149 vdd.n2148 185
R1064 vdd.n892 vdd.n891 185
R1065 vdd.n893 vdd.n892 185
R1066 vdd.n2141 vdd.n2140 185
R1067 vdd.n2142 vdd.n2141 185
R1068 vdd.n2139 vdd.n901 185
R1069 vdd.n907 vdd.n901 185
R1070 vdd.n2138 vdd.n2137 185
R1071 vdd.n2137 vdd.n2136 185
R1072 vdd.n903 vdd.n902 185
R1073 vdd.n904 vdd.n903 185
R1074 vdd.n2127 vdd.n2126 185
R1075 vdd.n2125 vdd.n946 185
R1076 vdd.n2124 vdd.n945 185
R1077 vdd.n2129 vdd.n945 185
R1078 vdd.n2123 vdd.n2122 185
R1079 vdd.n2121 vdd.n2120 185
R1080 vdd.n2119 vdd.n2118 185
R1081 vdd.n2117 vdd.n2116 185
R1082 vdd.n2115 vdd.n2114 185
R1083 vdd.n2113 vdd.n2112 185
R1084 vdd.n2111 vdd.n2110 185
R1085 vdd.n2109 vdd.n2108 185
R1086 vdd.n2107 vdd.n2106 185
R1087 vdd.n2105 vdd.n2104 185
R1088 vdd.n2103 vdd.n2102 185
R1089 vdd.n2101 vdd.n2100 185
R1090 vdd.n2099 vdd.n2098 185
R1091 vdd.n2097 vdd.n2096 185
R1092 vdd.n2095 vdd.n2094 185
R1093 vdd.n1103 vdd.n947 185
R1094 vdd.n1105 vdd.n1104 185
R1095 vdd.n1107 vdd.n1106 185
R1096 vdd.n1109 vdd.n1108 185
R1097 vdd.n1111 vdd.n1110 185
R1098 vdd.n1113 vdd.n1112 185
R1099 vdd.n1115 vdd.n1114 185
R1100 vdd.n1117 vdd.n1116 185
R1101 vdd.n1119 vdd.n1118 185
R1102 vdd.n1121 vdd.n1120 185
R1103 vdd.n1123 vdd.n1122 185
R1104 vdd.n1125 vdd.n1124 185
R1105 vdd.n1127 vdd.n1126 185
R1106 vdd.n1129 vdd.n1128 185
R1107 vdd.n1132 vdd.n1131 185
R1108 vdd.n1134 vdd.n1133 185
R1109 vdd.n1136 vdd.n1135 185
R1110 vdd.n2308 vdd.n2307 185
R1111 vdd.n2310 vdd.n2309 185
R1112 vdd.n2312 vdd.n2311 185
R1113 vdd.n2315 vdd.n2314 185
R1114 vdd.n2317 vdd.n2316 185
R1115 vdd.n2319 vdd.n2318 185
R1116 vdd.n2321 vdd.n2320 185
R1117 vdd.n2323 vdd.n2322 185
R1118 vdd.n2325 vdd.n2324 185
R1119 vdd.n2327 vdd.n2326 185
R1120 vdd.n2329 vdd.n2328 185
R1121 vdd.n2331 vdd.n2330 185
R1122 vdd.n2333 vdd.n2332 185
R1123 vdd.n2335 vdd.n2334 185
R1124 vdd.n2337 vdd.n2336 185
R1125 vdd.n2339 vdd.n2338 185
R1126 vdd.n2341 vdd.n2340 185
R1127 vdd.n2343 vdd.n2342 185
R1128 vdd.n2345 vdd.n2344 185
R1129 vdd.n2347 vdd.n2346 185
R1130 vdd.n2349 vdd.n2348 185
R1131 vdd.n2351 vdd.n2350 185
R1132 vdd.n2353 vdd.n2352 185
R1133 vdd.n2355 vdd.n2354 185
R1134 vdd.n2357 vdd.n2356 185
R1135 vdd.n2359 vdd.n2358 185
R1136 vdd.n2361 vdd.n2360 185
R1137 vdd.n2363 vdd.n2362 185
R1138 vdd.n2365 vdd.n2364 185
R1139 vdd.n2367 vdd.n2366 185
R1140 vdd.n2369 vdd.n2368 185
R1141 vdd.n2371 vdd.n2370 185
R1142 vdd.n2373 vdd.n2372 185
R1143 vdd.n2374 vdd.n798 185
R1144 vdd.n2376 vdd.n2375 185
R1145 vdd.n2377 vdd.n2376 185
R1146 vdd.n2306 vdd.n802 185
R1147 vdd.n2306 vdd.n2305 185
R1148 vdd.n1164 vdd.n803 185
R1149 vdd.n804 vdd.n803 185
R1150 vdd.n1165 vdd.n814 185
R1151 vdd.n2230 vdd.n814 185
R1152 vdd.n1168 vdd.n1167 185
R1153 vdd.n1167 vdd.n1166 185
R1154 vdd.n1169 vdd.n821 185
R1155 vdd.n2223 vdd.n821 185
R1156 vdd.n1171 vdd.n1170 185
R1157 vdd.n1170 vdd.n820 185
R1158 vdd.n1172 vdd.n828 185
R1159 vdd.n2215 vdd.n828 185
R1160 vdd.n1174 vdd.n1173 185
R1161 vdd.n1173 vdd.n827 185
R1162 vdd.n1175 vdd.n834 185
R1163 vdd.n2209 vdd.n834 185
R1164 vdd.n1177 vdd.n1176 185
R1165 vdd.n1176 vdd.n833 185
R1166 vdd.n1178 vdd.n839 185
R1167 vdd.n2203 vdd.n839 185
R1168 vdd.n1180 vdd.n1179 185
R1169 vdd.n1179 vdd.n846 185
R1170 vdd.n1181 vdd.n844 185
R1171 vdd.n2197 vdd.n844 185
R1172 vdd.n1183 vdd.n1182 185
R1173 vdd.n1182 vdd.n852 185
R1174 vdd.n1184 vdd.n850 185
R1175 vdd.n2191 vdd.n850 185
R1176 vdd.n1186 vdd.n1185 185
R1177 vdd.n1187 vdd.n1186 185
R1178 vdd.n1163 vdd.n857 185
R1179 vdd.n2185 vdd.n857 185
R1180 vdd.n1162 vdd.n1161 185
R1181 vdd.n1161 vdd.n856 185
R1182 vdd.n1160 vdd.n863 185
R1183 vdd.n2179 vdd.n863 185
R1184 vdd.n1159 vdd.n1158 185
R1185 vdd.n1158 vdd.n862 185
R1186 vdd.n1157 vdd.n868 185
R1187 vdd.n2173 vdd.n868 185
R1188 vdd.n1156 vdd.n1155 185
R1189 vdd.n1155 vdd.n876 185
R1190 vdd.n1154 vdd.n874 185
R1191 vdd.n2166 vdd.n874 185
R1192 vdd.n1153 vdd.n1152 185
R1193 vdd.n1152 vdd.n883 185
R1194 vdd.n1151 vdd.n881 185
R1195 vdd.n2160 vdd.n881 185
R1196 vdd.n1150 vdd.n1149 185
R1197 vdd.n1149 vdd.n880 185
R1198 vdd.n1148 vdd.n888 185
R1199 vdd.n2154 vdd.n888 185
R1200 vdd.n1147 vdd.n1146 185
R1201 vdd.n1146 vdd.n887 185
R1202 vdd.n1145 vdd.n894 185
R1203 vdd.n2148 vdd.n894 185
R1204 vdd.n1144 vdd.n1143 185
R1205 vdd.n1143 vdd.n893 185
R1206 vdd.n1142 vdd.n899 185
R1207 vdd.n2142 vdd.n899 185
R1208 vdd.n1141 vdd.n1140 185
R1209 vdd.n1140 vdd.n907 185
R1210 vdd.n1139 vdd.n905 185
R1211 vdd.n2136 vdd.n905 185
R1212 vdd.n1138 vdd.n1137 185
R1213 vdd.n1137 vdd.n904 185
R1214 vdd.n3229 vdd.n3228 185
R1215 vdd.n3230 vdd.n3229 185
R1216 vdd.n347 vdd.n346 185
R1217 vdd.n3231 vdd.n347 185
R1218 vdd.n3234 vdd.n3233 185
R1219 vdd.n3233 vdd.n3232 185
R1220 vdd.n3235 vdd.n341 185
R1221 vdd.n341 vdd.n340 185
R1222 vdd.n3237 vdd.n3236 185
R1223 vdd.n3238 vdd.n3237 185
R1224 vdd.n336 vdd.n335 185
R1225 vdd.n3239 vdd.n336 185
R1226 vdd.n3242 vdd.n3241 185
R1227 vdd.n3241 vdd.n3240 185
R1228 vdd.n3243 vdd.n330 185
R1229 vdd.n330 vdd.n329 185
R1230 vdd.n3245 vdd.n3244 185
R1231 vdd.n3246 vdd.n3245 185
R1232 vdd.n324 vdd.n323 185
R1233 vdd.n3247 vdd.n324 185
R1234 vdd.n3250 vdd.n3249 185
R1235 vdd.n3249 vdd.n3248 185
R1236 vdd.n3251 vdd.n319 185
R1237 vdd.n325 vdd.n319 185
R1238 vdd.n3253 vdd.n3252 185
R1239 vdd.n3254 vdd.n3253 185
R1240 vdd.n315 vdd.n313 185
R1241 vdd.n3255 vdd.n315 185
R1242 vdd.n3258 vdd.n3257 185
R1243 vdd.n3257 vdd.n3256 185
R1244 vdd.n314 vdd.n312 185
R1245 vdd.n481 vdd.n314 185
R1246 vdd.n3080 vdd.n3079 185
R1247 vdd.n3081 vdd.n3080 185
R1248 vdd.n483 vdd.n482 185
R1249 vdd.n3072 vdd.n482 185
R1250 vdd.n3075 vdd.n3074 185
R1251 vdd.n3074 vdd.n3073 185
R1252 vdd.n486 vdd.n485 185
R1253 vdd.n493 vdd.n486 185
R1254 vdd.n3063 vdd.n3062 185
R1255 vdd.n3064 vdd.n3063 185
R1256 vdd.n495 vdd.n494 185
R1257 vdd.n494 vdd.n492 185
R1258 vdd.n3058 vdd.n3057 185
R1259 vdd.n3057 vdd.n3056 185
R1260 vdd.n498 vdd.n497 185
R1261 vdd.n499 vdd.n498 185
R1262 vdd.n3047 vdd.n3046 185
R1263 vdd.n3048 vdd.n3047 185
R1264 vdd.n507 vdd.n506 185
R1265 vdd.n506 vdd.n505 185
R1266 vdd.n3042 vdd.n3041 185
R1267 vdd.n3041 vdd.n3040 185
R1268 vdd.n510 vdd.n509 185
R1269 vdd.n511 vdd.n510 185
R1270 vdd.n3031 vdd.n3030 185
R1271 vdd.n3032 vdd.n3031 185
R1272 vdd.n3027 vdd.n517 185
R1273 vdd.n3026 vdd.n3025 185
R1274 vdd.n3023 vdd.n519 185
R1275 vdd.n3023 vdd.n516 185
R1276 vdd.n3022 vdd.n3021 185
R1277 vdd.n3020 vdd.n3019 185
R1278 vdd.n3018 vdd.n3017 185
R1279 vdd.n3016 vdd.n3015 185
R1280 vdd.n3014 vdd.n525 185
R1281 vdd.n3012 vdd.n3011 185
R1282 vdd.n3010 vdd.n526 185
R1283 vdd.n3009 vdd.n3008 185
R1284 vdd.n3006 vdd.n531 185
R1285 vdd.n3004 vdd.n3003 185
R1286 vdd.n3002 vdd.n532 185
R1287 vdd.n3001 vdd.n3000 185
R1288 vdd.n2998 vdd.n537 185
R1289 vdd.n2996 vdd.n2995 185
R1290 vdd.n2994 vdd.n538 185
R1291 vdd.n2993 vdd.n2992 185
R1292 vdd.n2990 vdd.n545 185
R1293 vdd.n2988 vdd.n2987 185
R1294 vdd.n2986 vdd.n546 185
R1295 vdd.n2985 vdd.n2984 185
R1296 vdd.n2982 vdd.n551 185
R1297 vdd.n2980 vdd.n2979 185
R1298 vdd.n2978 vdd.n552 185
R1299 vdd.n2977 vdd.n2976 185
R1300 vdd.n2974 vdd.n557 185
R1301 vdd.n2972 vdd.n2971 185
R1302 vdd.n2970 vdd.n558 185
R1303 vdd.n2969 vdd.n2968 185
R1304 vdd.n2966 vdd.n563 185
R1305 vdd.n2964 vdd.n2963 185
R1306 vdd.n2962 vdd.n564 185
R1307 vdd.n2961 vdd.n2960 185
R1308 vdd.n2958 vdd.n569 185
R1309 vdd.n2956 vdd.n2955 185
R1310 vdd.n2954 vdd.n570 185
R1311 vdd.n2953 vdd.n2952 185
R1312 vdd.n2950 vdd.n575 185
R1313 vdd.n2948 vdd.n2947 185
R1314 vdd.n2946 vdd.n576 185
R1315 vdd.n585 vdd.n579 185
R1316 vdd.n2942 vdd.n2941 185
R1317 vdd.n2939 vdd.n583 185
R1318 vdd.n2938 vdd.n2937 185
R1319 vdd.n2936 vdd.n2935 185
R1320 vdd.n2934 vdd.n589 185
R1321 vdd.n2932 vdd.n2931 185
R1322 vdd.n2930 vdd.n590 185
R1323 vdd.n2929 vdd.n2928 185
R1324 vdd.n2926 vdd.n595 185
R1325 vdd.n2924 vdd.n2923 185
R1326 vdd.n2922 vdd.n596 185
R1327 vdd.n2921 vdd.n2920 185
R1328 vdd.n2918 vdd.n601 185
R1329 vdd.n2916 vdd.n2915 185
R1330 vdd.n2914 vdd.n602 185
R1331 vdd.n2913 vdd.n2912 185
R1332 vdd.n2910 vdd.n2909 185
R1333 vdd.n2908 vdd.n2907 185
R1334 vdd.n2906 vdd.n2905 185
R1335 vdd.n2904 vdd.n2903 185
R1336 vdd.n2899 vdd.n515 185
R1337 vdd.n516 vdd.n515 185
R1338 vdd.n3112 vdd.n3111 185
R1339 vdd.n3116 vdd.n462 185
R1340 vdd.n3118 vdd.n3117 185
R1341 vdd.n3120 vdd.n460 185
R1342 vdd.n3122 vdd.n3121 185
R1343 vdd.n3123 vdd.n455 185
R1344 vdd.n3125 vdd.n3124 185
R1345 vdd.n3127 vdd.n453 185
R1346 vdd.n3129 vdd.n3128 185
R1347 vdd.n3130 vdd.n448 185
R1348 vdd.n3132 vdd.n3131 185
R1349 vdd.n3134 vdd.n446 185
R1350 vdd.n3136 vdd.n3135 185
R1351 vdd.n3137 vdd.n441 185
R1352 vdd.n3139 vdd.n3138 185
R1353 vdd.n3141 vdd.n439 185
R1354 vdd.n3143 vdd.n3142 185
R1355 vdd.n3144 vdd.n435 185
R1356 vdd.n3146 vdd.n3145 185
R1357 vdd.n3148 vdd.n432 185
R1358 vdd.n3150 vdd.n3149 185
R1359 vdd.n433 vdd.n426 185
R1360 vdd.n3154 vdd.n430 185
R1361 vdd.n3155 vdd.n422 185
R1362 vdd.n3157 vdd.n3156 185
R1363 vdd.n3159 vdd.n420 185
R1364 vdd.n3161 vdd.n3160 185
R1365 vdd.n3162 vdd.n415 185
R1366 vdd.n3164 vdd.n3163 185
R1367 vdd.n3166 vdd.n413 185
R1368 vdd.n3168 vdd.n3167 185
R1369 vdd.n3169 vdd.n408 185
R1370 vdd.n3171 vdd.n3170 185
R1371 vdd.n3173 vdd.n406 185
R1372 vdd.n3175 vdd.n3174 185
R1373 vdd.n3176 vdd.n401 185
R1374 vdd.n3178 vdd.n3177 185
R1375 vdd.n3180 vdd.n399 185
R1376 vdd.n3182 vdd.n3181 185
R1377 vdd.n3183 vdd.n395 185
R1378 vdd.n3185 vdd.n3184 185
R1379 vdd.n3187 vdd.n392 185
R1380 vdd.n3189 vdd.n3188 185
R1381 vdd.n393 vdd.n386 185
R1382 vdd.n3193 vdd.n390 185
R1383 vdd.n3194 vdd.n382 185
R1384 vdd.n3196 vdd.n3195 185
R1385 vdd.n3198 vdd.n380 185
R1386 vdd.n3200 vdd.n3199 185
R1387 vdd.n3201 vdd.n375 185
R1388 vdd.n3203 vdd.n3202 185
R1389 vdd.n3205 vdd.n373 185
R1390 vdd.n3207 vdd.n3206 185
R1391 vdd.n3208 vdd.n368 185
R1392 vdd.n3210 vdd.n3209 185
R1393 vdd.n3212 vdd.n366 185
R1394 vdd.n3214 vdd.n3213 185
R1395 vdd.n3215 vdd.n360 185
R1396 vdd.n3217 vdd.n3216 185
R1397 vdd.n3219 vdd.n359 185
R1398 vdd.n3220 vdd.n358 185
R1399 vdd.n3223 vdd.n3222 185
R1400 vdd.n3224 vdd.n356 185
R1401 vdd.n3225 vdd.n352 185
R1402 vdd.n3107 vdd.n350 185
R1403 vdd.n3230 vdd.n350 185
R1404 vdd.n3106 vdd.n349 185
R1405 vdd.n3231 vdd.n349 185
R1406 vdd.n3105 vdd.n348 185
R1407 vdd.n3232 vdd.n348 185
R1408 vdd.n468 vdd.n467 185
R1409 vdd.n467 vdd.n340 185
R1410 vdd.n3101 vdd.n339 185
R1411 vdd.n3238 vdd.n339 185
R1412 vdd.n3100 vdd.n338 185
R1413 vdd.n3239 vdd.n338 185
R1414 vdd.n3099 vdd.n337 185
R1415 vdd.n3240 vdd.n337 185
R1416 vdd.n471 vdd.n470 185
R1417 vdd.n470 vdd.n329 185
R1418 vdd.n3095 vdd.n328 185
R1419 vdd.n3246 vdd.n328 185
R1420 vdd.n3094 vdd.n327 185
R1421 vdd.n3247 vdd.n327 185
R1422 vdd.n3093 vdd.n326 185
R1423 vdd.n3248 vdd.n326 185
R1424 vdd.n474 vdd.n473 185
R1425 vdd.n473 vdd.n325 185
R1426 vdd.n3089 vdd.n318 185
R1427 vdd.n3254 vdd.n318 185
R1428 vdd.n3088 vdd.n317 185
R1429 vdd.n3255 vdd.n317 185
R1430 vdd.n3087 vdd.n316 185
R1431 vdd.n3256 vdd.n316 185
R1432 vdd.n480 vdd.n476 185
R1433 vdd.n481 vdd.n480 185
R1434 vdd.n3083 vdd.n3082 185
R1435 vdd.n3082 vdd.n3081 185
R1436 vdd.n479 vdd.n478 185
R1437 vdd.n3072 vdd.n479 185
R1438 vdd.n3071 vdd.n3070 185
R1439 vdd.n3073 vdd.n3071 185
R1440 vdd.n488 vdd.n487 185
R1441 vdd.n493 vdd.n487 185
R1442 vdd.n3066 vdd.n3065 185
R1443 vdd.n3065 vdd.n3064 185
R1444 vdd.n491 vdd.n490 185
R1445 vdd.n492 vdd.n491 185
R1446 vdd.n3055 vdd.n3054 185
R1447 vdd.n3056 vdd.n3055 185
R1448 vdd.n501 vdd.n500 185
R1449 vdd.n500 vdd.n499 185
R1450 vdd.n3050 vdd.n3049 185
R1451 vdd.n3049 vdd.n3048 185
R1452 vdd.n504 vdd.n503 185
R1453 vdd.n505 vdd.n504 185
R1454 vdd.n3039 vdd.n3038 185
R1455 vdd.n3040 vdd.n3039 185
R1456 vdd.n513 vdd.n512 185
R1457 vdd.n512 vdd.n511 185
R1458 vdd.n3034 vdd.n3033 185
R1459 vdd.n3033 vdd.n3032 185
R1460 vdd.n2648 vdd.n2647 185
R1461 vdd.n2646 vdd.n2412 185
R1462 vdd.n2645 vdd.n2411 185
R1463 vdd.n2650 vdd.n2411 185
R1464 vdd.n2644 vdd.n2643 185
R1465 vdd.n2642 vdd.n2641 185
R1466 vdd.n2640 vdd.n2639 185
R1467 vdd.n2638 vdd.n2637 185
R1468 vdd.n2636 vdd.n2635 185
R1469 vdd.n2634 vdd.n2633 185
R1470 vdd.n2632 vdd.n2631 185
R1471 vdd.n2630 vdd.n2629 185
R1472 vdd.n2628 vdd.n2627 185
R1473 vdd.n2626 vdd.n2625 185
R1474 vdd.n2624 vdd.n2623 185
R1475 vdd.n2622 vdd.n2621 185
R1476 vdd.n2620 vdd.n2619 185
R1477 vdd.n2618 vdd.n2617 185
R1478 vdd.n2616 vdd.n2615 185
R1479 vdd.n2614 vdd.n2613 185
R1480 vdd.n2612 vdd.n2611 185
R1481 vdd.n2610 vdd.n2609 185
R1482 vdd.n2608 vdd.n2607 185
R1483 vdd.n2606 vdd.n2605 185
R1484 vdd.n2604 vdd.n2603 185
R1485 vdd.n2602 vdd.n2601 185
R1486 vdd.n2600 vdd.n2599 185
R1487 vdd.n2598 vdd.n2597 185
R1488 vdd.n2596 vdd.n2595 185
R1489 vdd.n2594 vdd.n2593 185
R1490 vdd.n2592 vdd.n2591 185
R1491 vdd.n2590 vdd.n2589 185
R1492 vdd.n2588 vdd.n2587 185
R1493 vdd.n2585 vdd.n2584 185
R1494 vdd.n2583 vdd.n2582 185
R1495 vdd.n2581 vdd.n2580 185
R1496 vdd.n2800 vdd.n2799 185
R1497 vdd.n2801 vdd.n660 185
R1498 vdd.n2803 vdd.n2802 185
R1499 vdd.n2805 vdd.n658 185
R1500 vdd.n2807 vdd.n2806 185
R1501 vdd.n2808 vdd.n657 185
R1502 vdd.n2810 vdd.n2809 185
R1503 vdd.n2812 vdd.n655 185
R1504 vdd.n2814 vdd.n2813 185
R1505 vdd.n2815 vdd.n654 185
R1506 vdd.n2817 vdd.n2816 185
R1507 vdd.n2819 vdd.n652 185
R1508 vdd.n2821 vdd.n2820 185
R1509 vdd.n2822 vdd.n651 185
R1510 vdd.n2824 vdd.n2823 185
R1511 vdd.n2826 vdd.n649 185
R1512 vdd.n2828 vdd.n2827 185
R1513 vdd.n2830 vdd.n648 185
R1514 vdd.n2832 vdd.n2831 185
R1515 vdd.n2834 vdd.n646 185
R1516 vdd.n2836 vdd.n2835 185
R1517 vdd.n2837 vdd.n645 185
R1518 vdd.n2839 vdd.n2838 185
R1519 vdd.n2841 vdd.n643 185
R1520 vdd.n2843 vdd.n2842 185
R1521 vdd.n2844 vdd.n642 185
R1522 vdd.n2846 vdd.n2845 185
R1523 vdd.n2848 vdd.n640 185
R1524 vdd.n2850 vdd.n2849 185
R1525 vdd.n2851 vdd.n639 185
R1526 vdd.n2853 vdd.n2852 185
R1527 vdd.n2855 vdd.n638 185
R1528 vdd.n2856 vdd.n637 185
R1529 vdd.n2859 vdd.n2858 185
R1530 vdd.n2860 vdd.n635 185
R1531 vdd.n635 vdd.n613 185
R1532 vdd.n2797 vdd.n632 185
R1533 vdd.n2863 vdd.n632 185
R1534 vdd.n2796 vdd.n2795 185
R1535 vdd.n2795 vdd.n631 185
R1536 vdd.n2794 vdd.n664 185
R1537 vdd.n2794 vdd.n2793 185
R1538 vdd.n2528 vdd.n665 185
R1539 vdd.n674 vdd.n665 185
R1540 vdd.n2529 vdd.n672 185
R1541 vdd.n2787 vdd.n672 185
R1542 vdd.n2531 vdd.n2530 185
R1543 vdd.n2530 vdd.n671 185
R1544 vdd.n2532 vdd.n680 185
R1545 vdd.n2736 vdd.n680 185
R1546 vdd.n2534 vdd.n2533 185
R1547 vdd.n2533 vdd.n679 185
R1548 vdd.n2535 vdd.n686 185
R1549 vdd.n2730 vdd.n686 185
R1550 vdd.n2537 vdd.n2536 185
R1551 vdd.n2536 vdd.n685 185
R1552 vdd.n2538 vdd.n691 185
R1553 vdd.n2724 vdd.n691 185
R1554 vdd.n2540 vdd.n2539 185
R1555 vdd.n2539 vdd.n698 185
R1556 vdd.n2541 vdd.n696 185
R1557 vdd.n2718 vdd.n696 185
R1558 vdd.n2543 vdd.n2542 185
R1559 vdd.n2542 vdd.n706 185
R1560 vdd.n2544 vdd.n704 185
R1561 vdd.n2711 vdd.n704 185
R1562 vdd.n2546 vdd.n2545 185
R1563 vdd.n2545 vdd.n703 185
R1564 vdd.n2547 vdd.n711 185
R1565 vdd.n2705 vdd.n711 185
R1566 vdd.n2549 vdd.n2548 185
R1567 vdd.n2548 vdd.n710 185
R1568 vdd.n2550 vdd.n716 185
R1569 vdd.n2699 vdd.n716 185
R1570 vdd.n2552 vdd.n2551 185
R1571 vdd.n2551 vdd.n723 185
R1572 vdd.n2553 vdd.n721 185
R1573 vdd.n2693 vdd.n721 185
R1574 vdd.n2555 vdd.n2554 185
R1575 vdd.n2554 vdd.n729 185
R1576 vdd.n2556 vdd.n727 185
R1577 vdd.n2687 vdd.n727 185
R1578 vdd.n2558 vdd.n2557 185
R1579 vdd.n2559 vdd.n2558 185
R1580 vdd.n2527 vdd.n734 185
R1581 vdd.n2681 vdd.n734 185
R1582 vdd.n2526 vdd.n2525 185
R1583 vdd.n2525 vdd.n733 185
R1584 vdd.n2524 vdd.n740 185
R1585 vdd.n2675 vdd.n740 185
R1586 vdd.n2523 vdd.n2522 185
R1587 vdd.n2522 vdd.n739 185
R1588 vdd.n2521 vdd.n746 185
R1589 vdd.n2669 vdd.n746 185
R1590 vdd.n2520 vdd.n2519 185
R1591 vdd.n2519 vdd.n745 185
R1592 vdd.n2415 vdd.n751 185
R1593 vdd.n2663 vdd.n751 185
R1594 vdd.n2576 vdd.n2575 185
R1595 vdd.n2575 vdd.n2574 185
R1596 vdd.n2577 vdd.n757 185
R1597 vdd.n2657 vdd.n757 185
R1598 vdd.n2579 vdd.n2578 185
R1599 vdd.n2579 vdd.n756 185
R1600 vdd.n755 vdd.n754 185
R1601 vdd.n756 vdd.n755 185
R1602 vdd.n2659 vdd.n2658 185
R1603 vdd.n2658 vdd.n2657 185
R1604 vdd.n2660 vdd.n753 185
R1605 vdd.n2574 vdd.n753 185
R1606 vdd.n2662 vdd.n2661 185
R1607 vdd.n2663 vdd.n2662 185
R1608 vdd.n744 vdd.n743 185
R1609 vdd.n745 vdd.n744 185
R1610 vdd.n2671 vdd.n2670 185
R1611 vdd.n2670 vdd.n2669 185
R1612 vdd.n2672 vdd.n742 185
R1613 vdd.n742 vdd.n739 185
R1614 vdd.n2674 vdd.n2673 185
R1615 vdd.n2675 vdd.n2674 185
R1616 vdd.n732 vdd.n731 185
R1617 vdd.n733 vdd.n732 185
R1618 vdd.n2683 vdd.n2682 185
R1619 vdd.n2682 vdd.n2681 185
R1620 vdd.n2684 vdd.n730 185
R1621 vdd.n2559 vdd.n730 185
R1622 vdd.n2686 vdd.n2685 185
R1623 vdd.n2687 vdd.n2686 185
R1624 vdd.n720 vdd.n719 185
R1625 vdd.n729 vdd.n720 185
R1626 vdd.n2695 vdd.n2694 185
R1627 vdd.n2694 vdd.n2693 185
R1628 vdd.n2696 vdd.n718 185
R1629 vdd.n723 vdd.n718 185
R1630 vdd.n2698 vdd.n2697 185
R1631 vdd.n2699 vdd.n2698 185
R1632 vdd.n709 vdd.n708 185
R1633 vdd.n710 vdd.n709 185
R1634 vdd.n2707 vdd.n2706 185
R1635 vdd.n2706 vdd.n2705 185
R1636 vdd.n2708 vdd.n707 185
R1637 vdd.n707 vdd.n703 185
R1638 vdd.n2710 vdd.n2709 185
R1639 vdd.n2711 vdd.n2710 185
R1640 vdd.n695 vdd.n694 185
R1641 vdd.n706 vdd.n695 185
R1642 vdd.n2720 vdd.n2719 185
R1643 vdd.n2719 vdd.n2718 185
R1644 vdd.n2721 vdd.n693 185
R1645 vdd.n698 vdd.n693 185
R1646 vdd.n2723 vdd.n2722 185
R1647 vdd.n2724 vdd.n2723 185
R1648 vdd.n684 vdd.n683 185
R1649 vdd.n685 vdd.n684 185
R1650 vdd.n2732 vdd.n2731 185
R1651 vdd.n2731 vdd.n2730 185
R1652 vdd.n2733 vdd.n682 185
R1653 vdd.n682 vdd.n679 185
R1654 vdd.n2735 vdd.n2734 185
R1655 vdd.n2736 vdd.n2735 185
R1656 vdd.n670 vdd.n669 185
R1657 vdd.n671 vdd.n670 185
R1658 vdd.n2789 vdd.n2788 185
R1659 vdd.n2788 vdd.n2787 185
R1660 vdd.n2790 vdd.n668 185
R1661 vdd.n674 vdd.n668 185
R1662 vdd.n2792 vdd.n2791 185
R1663 vdd.n2793 vdd.n2792 185
R1664 vdd.n636 vdd.n634 185
R1665 vdd.n634 vdd.n631 185
R1666 vdd.n2862 vdd.n2861 185
R1667 vdd.n2863 vdd.n2862 185
R1668 vdd.n2304 vdd.n2303 185
R1669 vdd.n2305 vdd.n2304 185
R1670 vdd.n808 vdd.n806 185
R1671 vdd.n806 vdd.n804 185
R1672 vdd.n2219 vdd.n815 185
R1673 vdd.n2230 vdd.n815 185
R1674 vdd.n2220 vdd.n824 185
R1675 vdd.n1166 vdd.n824 185
R1676 vdd.n2222 vdd.n2221 185
R1677 vdd.n2223 vdd.n2222 185
R1678 vdd.n2218 vdd.n823 185
R1679 vdd.n823 vdd.n820 185
R1680 vdd.n2217 vdd.n2216 185
R1681 vdd.n2216 vdd.n2215 185
R1682 vdd.n826 vdd.n825 185
R1683 vdd.n827 vdd.n826 185
R1684 vdd.n2208 vdd.n2207 185
R1685 vdd.n2209 vdd.n2208 185
R1686 vdd.n2206 vdd.n836 185
R1687 vdd.n836 vdd.n833 185
R1688 vdd.n2205 vdd.n2204 185
R1689 vdd.n2204 vdd.n2203 185
R1690 vdd.n838 vdd.n837 185
R1691 vdd.n846 vdd.n838 185
R1692 vdd.n2196 vdd.n2195 185
R1693 vdd.n2197 vdd.n2196 185
R1694 vdd.n2194 vdd.n847 185
R1695 vdd.n852 vdd.n847 185
R1696 vdd.n2193 vdd.n2192 185
R1697 vdd.n2192 vdd.n2191 185
R1698 vdd.n849 vdd.n848 185
R1699 vdd.n1187 vdd.n849 185
R1700 vdd.n2184 vdd.n2183 185
R1701 vdd.n2185 vdd.n2184 185
R1702 vdd.n2182 vdd.n859 185
R1703 vdd.n859 vdd.n856 185
R1704 vdd.n2181 vdd.n2180 185
R1705 vdd.n2180 vdd.n2179 185
R1706 vdd.n861 vdd.n860 185
R1707 vdd.n862 vdd.n861 185
R1708 vdd.n2172 vdd.n2171 185
R1709 vdd.n2173 vdd.n2172 185
R1710 vdd.n2169 vdd.n870 185
R1711 vdd.n876 vdd.n870 185
R1712 vdd.n2168 vdd.n2167 185
R1713 vdd.n2167 vdd.n2166 185
R1714 vdd.n873 vdd.n872 185
R1715 vdd.n883 vdd.n873 185
R1716 vdd.n2159 vdd.n2158 185
R1717 vdd.n2160 vdd.n2159 185
R1718 vdd.n2157 vdd.n884 185
R1719 vdd.n884 vdd.n880 185
R1720 vdd.n2156 vdd.n2155 185
R1721 vdd.n2155 vdd.n2154 185
R1722 vdd.n886 vdd.n885 185
R1723 vdd.n887 vdd.n886 185
R1724 vdd.n2147 vdd.n2146 185
R1725 vdd.n2148 vdd.n2147 185
R1726 vdd.n2145 vdd.n896 185
R1727 vdd.n896 vdd.n893 185
R1728 vdd.n2144 vdd.n2143 185
R1729 vdd.n2143 vdd.n2142 185
R1730 vdd.n898 vdd.n897 185
R1731 vdd.n907 vdd.n898 185
R1732 vdd.n2135 vdd.n2134 185
R1733 vdd.n2136 vdd.n2135 185
R1734 vdd.n2133 vdd.n908 185
R1735 vdd.n908 vdd.n904 185
R1736 vdd.n2235 vdd.n779 185
R1737 vdd.n2377 vdd.n779 185
R1738 vdd.n2237 vdd.n2236 185
R1739 vdd.n2239 vdd.n2238 185
R1740 vdd.n2241 vdd.n2240 185
R1741 vdd.n2243 vdd.n2242 185
R1742 vdd.n2245 vdd.n2244 185
R1743 vdd.n2247 vdd.n2246 185
R1744 vdd.n2249 vdd.n2248 185
R1745 vdd.n2251 vdd.n2250 185
R1746 vdd.n2253 vdd.n2252 185
R1747 vdd.n2255 vdd.n2254 185
R1748 vdd.n2257 vdd.n2256 185
R1749 vdd.n2259 vdd.n2258 185
R1750 vdd.n2261 vdd.n2260 185
R1751 vdd.n2263 vdd.n2262 185
R1752 vdd.n2265 vdd.n2264 185
R1753 vdd.n2267 vdd.n2266 185
R1754 vdd.n2269 vdd.n2268 185
R1755 vdd.n2271 vdd.n2270 185
R1756 vdd.n2273 vdd.n2272 185
R1757 vdd.n2275 vdd.n2274 185
R1758 vdd.n2277 vdd.n2276 185
R1759 vdd.n2279 vdd.n2278 185
R1760 vdd.n2281 vdd.n2280 185
R1761 vdd.n2283 vdd.n2282 185
R1762 vdd.n2285 vdd.n2284 185
R1763 vdd.n2287 vdd.n2286 185
R1764 vdd.n2289 vdd.n2288 185
R1765 vdd.n2291 vdd.n2290 185
R1766 vdd.n2293 vdd.n2292 185
R1767 vdd.n2295 vdd.n2294 185
R1768 vdd.n2297 vdd.n2296 185
R1769 vdd.n2299 vdd.n2298 185
R1770 vdd.n2301 vdd.n2300 185
R1771 vdd.n2302 vdd.n807 185
R1772 vdd.n2234 vdd.n805 185
R1773 vdd.n2305 vdd.n805 185
R1774 vdd.n2233 vdd.n2232 185
R1775 vdd.n2232 vdd.n804 185
R1776 vdd.n2231 vdd.n812 185
R1777 vdd.n2231 vdd.n2230 185
R1778 vdd.n1084 vdd.n813 185
R1779 vdd.n1166 vdd.n813 185
R1780 vdd.n1085 vdd.n822 185
R1781 vdd.n2223 vdd.n822 185
R1782 vdd.n1087 vdd.n1086 185
R1783 vdd.n1086 vdd.n820 185
R1784 vdd.n1088 vdd.n829 185
R1785 vdd.n2215 vdd.n829 185
R1786 vdd.n1090 vdd.n1089 185
R1787 vdd.n1089 vdd.n827 185
R1788 vdd.n1091 vdd.n835 185
R1789 vdd.n2209 vdd.n835 185
R1790 vdd.n1093 vdd.n1092 185
R1791 vdd.n1092 vdd.n833 185
R1792 vdd.n1094 vdd.n840 185
R1793 vdd.n2203 vdd.n840 185
R1794 vdd.n1096 vdd.n1095 185
R1795 vdd.n1095 vdd.n846 185
R1796 vdd.n1097 vdd.n845 185
R1797 vdd.n2197 vdd.n845 185
R1798 vdd.n1099 vdd.n1098 185
R1799 vdd.n1098 vdd.n852 185
R1800 vdd.n1100 vdd.n851 185
R1801 vdd.n2191 vdd.n851 185
R1802 vdd.n1189 vdd.n1188 185
R1803 vdd.n1188 vdd.n1187 185
R1804 vdd.n1190 vdd.n858 185
R1805 vdd.n2185 vdd.n858 185
R1806 vdd.n1192 vdd.n1191 185
R1807 vdd.n1191 vdd.n856 185
R1808 vdd.n1193 vdd.n864 185
R1809 vdd.n2179 vdd.n864 185
R1810 vdd.n1195 vdd.n1194 185
R1811 vdd.n1194 vdd.n862 185
R1812 vdd.n1196 vdd.n869 185
R1813 vdd.n2173 vdd.n869 185
R1814 vdd.n1198 vdd.n1197 185
R1815 vdd.n1197 vdd.n876 185
R1816 vdd.n1199 vdd.n875 185
R1817 vdd.n2166 vdd.n875 185
R1818 vdd.n1201 vdd.n1200 185
R1819 vdd.n1200 vdd.n883 185
R1820 vdd.n1202 vdd.n882 185
R1821 vdd.n2160 vdd.n882 185
R1822 vdd.n1204 vdd.n1203 185
R1823 vdd.n1203 vdd.n880 185
R1824 vdd.n1205 vdd.n889 185
R1825 vdd.n2154 vdd.n889 185
R1826 vdd.n1207 vdd.n1206 185
R1827 vdd.n1206 vdd.n887 185
R1828 vdd.n1208 vdd.n895 185
R1829 vdd.n2148 vdd.n895 185
R1830 vdd.n1210 vdd.n1209 185
R1831 vdd.n1209 vdd.n893 185
R1832 vdd.n1211 vdd.n900 185
R1833 vdd.n2142 vdd.n900 185
R1834 vdd.n1213 vdd.n1212 185
R1835 vdd.n1212 vdd.n907 185
R1836 vdd.n1214 vdd.n906 185
R1837 vdd.n2136 vdd.n906 185
R1838 vdd.n1216 vdd.n1215 185
R1839 vdd.n1215 vdd.n904 185
R1840 vdd.n2132 vdd.n2131 185
R1841 vdd.n910 vdd.n909 185
R1842 vdd.n1051 vdd.n1050 185
R1843 vdd.n1053 vdd.n1052 185
R1844 vdd.n1055 vdd.n1054 185
R1845 vdd.n1057 vdd.n1056 185
R1846 vdd.n1059 vdd.n1058 185
R1847 vdd.n1061 vdd.n1060 185
R1848 vdd.n1063 vdd.n1062 185
R1849 vdd.n1065 vdd.n1064 185
R1850 vdd.n1067 vdd.n1066 185
R1851 vdd.n1069 vdd.n1068 185
R1852 vdd.n1071 vdd.n1070 185
R1853 vdd.n1073 vdd.n1072 185
R1854 vdd.n1075 vdd.n1074 185
R1855 vdd.n1077 vdd.n1076 185
R1856 vdd.n1079 vdd.n1078 185
R1857 vdd.n1250 vdd.n1080 185
R1858 vdd.n1249 vdd.n1248 185
R1859 vdd.n1247 vdd.n1246 185
R1860 vdd.n1245 vdd.n1244 185
R1861 vdd.n1243 vdd.n1242 185
R1862 vdd.n1241 vdd.n1240 185
R1863 vdd.n1239 vdd.n1238 185
R1864 vdd.n1237 vdd.n1236 185
R1865 vdd.n1235 vdd.n1234 185
R1866 vdd.n1233 vdd.n1232 185
R1867 vdd.n1231 vdd.n1230 185
R1868 vdd.n1229 vdd.n1228 185
R1869 vdd.n1227 vdd.n1226 185
R1870 vdd.n1225 vdd.n1224 185
R1871 vdd.n1223 vdd.n1222 185
R1872 vdd.n1221 vdd.n1220 185
R1873 vdd.n1219 vdd.n1218 185
R1874 vdd.n1217 vdd.n944 185
R1875 vdd.n2129 vdd.n944 185
R1876 vdd.n2129 vdd.n911 179.345
R1877 vdd.n613 vdd.n516 179.345
R1878 vdd.n303 vdd.n302 171.744
R1879 vdd.n302 vdd.n301 171.744
R1880 vdd.n301 vdd.n270 171.744
R1881 vdd.n294 vdd.n270 171.744
R1882 vdd.n294 vdd.n293 171.744
R1883 vdd.n293 vdd.n275 171.744
R1884 vdd.n286 vdd.n275 171.744
R1885 vdd.n286 vdd.n285 171.744
R1886 vdd.n285 vdd.n279 171.744
R1887 vdd.n252 vdd.n251 171.744
R1888 vdd.n251 vdd.n250 171.744
R1889 vdd.n250 vdd.n219 171.744
R1890 vdd.n243 vdd.n219 171.744
R1891 vdd.n243 vdd.n242 171.744
R1892 vdd.n242 vdd.n224 171.744
R1893 vdd.n235 vdd.n224 171.744
R1894 vdd.n235 vdd.n234 171.744
R1895 vdd.n234 vdd.n228 171.744
R1896 vdd.n209 vdd.n208 171.744
R1897 vdd.n208 vdd.n207 171.744
R1898 vdd.n207 vdd.n176 171.744
R1899 vdd.n200 vdd.n176 171.744
R1900 vdd.n200 vdd.n199 171.744
R1901 vdd.n199 vdd.n181 171.744
R1902 vdd.n192 vdd.n181 171.744
R1903 vdd.n192 vdd.n191 171.744
R1904 vdd.n191 vdd.n185 171.744
R1905 vdd.n158 vdd.n157 171.744
R1906 vdd.n157 vdd.n156 171.744
R1907 vdd.n156 vdd.n125 171.744
R1908 vdd.n149 vdd.n125 171.744
R1909 vdd.n149 vdd.n148 171.744
R1910 vdd.n148 vdd.n130 171.744
R1911 vdd.n141 vdd.n130 171.744
R1912 vdd.n141 vdd.n140 171.744
R1913 vdd.n140 vdd.n134 171.744
R1914 vdd.n116 vdd.n115 171.744
R1915 vdd.n115 vdd.n114 171.744
R1916 vdd.n114 vdd.n83 171.744
R1917 vdd.n107 vdd.n83 171.744
R1918 vdd.n107 vdd.n106 171.744
R1919 vdd.n106 vdd.n88 171.744
R1920 vdd.n99 vdd.n88 171.744
R1921 vdd.n99 vdd.n98 171.744
R1922 vdd.n98 vdd.n92 171.744
R1923 vdd.n65 vdd.n64 171.744
R1924 vdd.n64 vdd.n63 171.744
R1925 vdd.n63 vdd.n32 171.744
R1926 vdd.n56 vdd.n32 171.744
R1927 vdd.n56 vdd.n55 171.744
R1928 vdd.n55 vdd.n37 171.744
R1929 vdd.n48 vdd.n37 171.744
R1930 vdd.n48 vdd.n47 171.744
R1931 vdd.n47 vdd.n41 171.744
R1932 vdd.n1860 vdd.n1859 171.744
R1933 vdd.n1859 vdd.n1858 171.744
R1934 vdd.n1858 vdd.n1827 171.744
R1935 vdd.n1851 vdd.n1827 171.744
R1936 vdd.n1851 vdd.n1850 171.744
R1937 vdd.n1850 vdd.n1832 171.744
R1938 vdd.n1843 vdd.n1832 171.744
R1939 vdd.n1843 vdd.n1842 171.744
R1940 vdd.n1842 vdd.n1836 171.744
R1941 vdd.n1911 vdd.n1910 171.744
R1942 vdd.n1910 vdd.n1909 171.744
R1943 vdd.n1909 vdd.n1878 171.744
R1944 vdd.n1902 vdd.n1878 171.744
R1945 vdd.n1902 vdd.n1901 171.744
R1946 vdd.n1901 vdd.n1883 171.744
R1947 vdd.n1894 vdd.n1883 171.744
R1948 vdd.n1894 vdd.n1893 171.744
R1949 vdd.n1893 vdd.n1887 171.744
R1950 vdd.n1766 vdd.n1765 171.744
R1951 vdd.n1765 vdd.n1764 171.744
R1952 vdd.n1764 vdd.n1733 171.744
R1953 vdd.n1757 vdd.n1733 171.744
R1954 vdd.n1757 vdd.n1756 171.744
R1955 vdd.n1756 vdd.n1738 171.744
R1956 vdd.n1749 vdd.n1738 171.744
R1957 vdd.n1749 vdd.n1748 171.744
R1958 vdd.n1748 vdd.n1742 171.744
R1959 vdd.n1817 vdd.n1816 171.744
R1960 vdd.n1816 vdd.n1815 171.744
R1961 vdd.n1815 vdd.n1784 171.744
R1962 vdd.n1808 vdd.n1784 171.744
R1963 vdd.n1808 vdd.n1807 171.744
R1964 vdd.n1807 vdd.n1789 171.744
R1965 vdd.n1800 vdd.n1789 171.744
R1966 vdd.n1800 vdd.n1799 171.744
R1967 vdd.n1799 vdd.n1793 171.744
R1968 vdd.n1673 vdd.n1672 171.744
R1969 vdd.n1672 vdd.n1671 171.744
R1970 vdd.n1671 vdd.n1640 171.744
R1971 vdd.n1664 vdd.n1640 171.744
R1972 vdd.n1664 vdd.n1663 171.744
R1973 vdd.n1663 vdd.n1645 171.744
R1974 vdd.n1656 vdd.n1645 171.744
R1975 vdd.n1656 vdd.n1655 171.744
R1976 vdd.n1655 vdd.n1649 171.744
R1977 vdd.n1724 vdd.n1723 171.744
R1978 vdd.n1723 vdd.n1722 171.744
R1979 vdd.n1722 vdd.n1691 171.744
R1980 vdd.n1715 vdd.n1691 171.744
R1981 vdd.n1715 vdd.n1714 171.744
R1982 vdd.n1714 vdd.n1696 171.744
R1983 vdd.n1707 vdd.n1696 171.744
R1984 vdd.n1707 vdd.n1706 171.744
R1985 vdd.n1706 vdd.n1700 171.744
R1986 vdd.n3222 vdd.n356 146.341
R1987 vdd.n3220 vdd.n3219 146.341
R1988 vdd.n3217 vdd.n360 146.341
R1989 vdd.n3213 vdd.n3212 146.341
R1990 vdd.n3210 vdd.n368 146.341
R1991 vdd.n3206 vdd.n3205 146.341
R1992 vdd.n3203 vdd.n375 146.341
R1993 vdd.n3199 vdd.n3198 146.341
R1994 vdd.n3196 vdd.n382 146.341
R1995 vdd.n393 vdd.n390 146.341
R1996 vdd.n3188 vdd.n3187 146.341
R1997 vdd.n3185 vdd.n395 146.341
R1998 vdd.n3181 vdd.n3180 146.341
R1999 vdd.n3178 vdd.n401 146.341
R2000 vdd.n3174 vdd.n3173 146.341
R2001 vdd.n3171 vdd.n408 146.341
R2002 vdd.n3167 vdd.n3166 146.341
R2003 vdd.n3164 vdd.n415 146.341
R2004 vdd.n3160 vdd.n3159 146.341
R2005 vdd.n3157 vdd.n422 146.341
R2006 vdd.n433 vdd.n430 146.341
R2007 vdd.n3149 vdd.n3148 146.341
R2008 vdd.n3146 vdd.n435 146.341
R2009 vdd.n3142 vdd.n3141 146.341
R2010 vdd.n3139 vdd.n441 146.341
R2011 vdd.n3135 vdd.n3134 146.341
R2012 vdd.n3132 vdd.n448 146.341
R2013 vdd.n3128 vdd.n3127 146.341
R2014 vdd.n3125 vdd.n455 146.341
R2015 vdd.n3121 vdd.n3120 146.341
R2016 vdd.n3118 vdd.n462 146.341
R2017 vdd.n3033 vdd.n512 146.341
R2018 vdd.n3039 vdd.n512 146.341
R2019 vdd.n3039 vdd.n504 146.341
R2020 vdd.n3049 vdd.n504 146.341
R2021 vdd.n3049 vdd.n500 146.341
R2022 vdd.n3055 vdd.n500 146.341
R2023 vdd.n3055 vdd.n491 146.341
R2024 vdd.n3065 vdd.n491 146.341
R2025 vdd.n3065 vdd.n487 146.341
R2026 vdd.n3071 vdd.n487 146.341
R2027 vdd.n3071 vdd.n479 146.341
R2028 vdd.n3082 vdd.n479 146.341
R2029 vdd.n3082 vdd.n480 146.341
R2030 vdd.n480 vdd.n316 146.341
R2031 vdd.n317 vdd.n316 146.341
R2032 vdd.n318 vdd.n317 146.341
R2033 vdd.n473 vdd.n318 146.341
R2034 vdd.n473 vdd.n326 146.341
R2035 vdd.n327 vdd.n326 146.341
R2036 vdd.n328 vdd.n327 146.341
R2037 vdd.n470 vdd.n328 146.341
R2038 vdd.n470 vdd.n337 146.341
R2039 vdd.n338 vdd.n337 146.341
R2040 vdd.n339 vdd.n338 146.341
R2041 vdd.n467 vdd.n339 146.341
R2042 vdd.n467 vdd.n348 146.341
R2043 vdd.n349 vdd.n348 146.341
R2044 vdd.n350 vdd.n349 146.341
R2045 vdd.n3025 vdd.n3023 146.341
R2046 vdd.n3023 vdd.n3022 146.341
R2047 vdd.n3019 vdd.n3018 146.341
R2048 vdd.n3015 vdd.n3014 146.341
R2049 vdd.n3012 vdd.n526 146.341
R2050 vdd.n3008 vdd.n3006 146.341
R2051 vdd.n3004 vdd.n532 146.341
R2052 vdd.n3000 vdd.n2998 146.341
R2053 vdd.n2996 vdd.n538 146.341
R2054 vdd.n2992 vdd.n2990 146.341
R2055 vdd.n2988 vdd.n546 146.341
R2056 vdd.n2984 vdd.n2982 146.341
R2057 vdd.n2980 vdd.n552 146.341
R2058 vdd.n2976 vdd.n2974 146.341
R2059 vdd.n2972 vdd.n558 146.341
R2060 vdd.n2968 vdd.n2966 146.341
R2061 vdd.n2964 vdd.n564 146.341
R2062 vdd.n2960 vdd.n2958 146.341
R2063 vdd.n2956 vdd.n570 146.341
R2064 vdd.n2952 vdd.n2950 146.341
R2065 vdd.n2948 vdd.n576 146.341
R2066 vdd.n2941 vdd.n585 146.341
R2067 vdd.n2939 vdd.n2938 146.341
R2068 vdd.n2935 vdd.n2934 146.341
R2069 vdd.n2932 vdd.n590 146.341
R2070 vdd.n2928 vdd.n2926 146.341
R2071 vdd.n2924 vdd.n596 146.341
R2072 vdd.n2920 vdd.n2918 146.341
R2073 vdd.n2916 vdd.n602 146.341
R2074 vdd.n2912 vdd.n2910 146.341
R2075 vdd.n2907 vdd.n2906 146.341
R2076 vdd.n2903 vdd.n515 146.341
R2077 vdd.n3031 vdd.n510 146.341
R2078 vdd.n3041 vdd.n510 146.341
R2079 vdd.n3041 vdd.n506 146.341
R2080 vdd.n3047 vdd.n506 146.341
R2081 vdd.n3047 vdd.n498 146.341
R2082 vdd.n3057 vdd.n498 146.341
R2083 vdd.n3057 vdd.n494 146.341
R2084 vdd.n3063 vdd.n494 146.341
R2085 vdd.n3063 vdd.n486 146.341
R2086 vdd.n3074 vdd.n486 146.341
R2087 vdd.n3074 vdd.n482 146.341
R2088 vdd.n3080 vdd.n482 146.341
R2089 vdd.n3080 vdd.n314 146.341
R2090 vdd.n3257 vdd.n314 146.341
R2091 vdd.n3257 vdd.n315 146.341
R2092 vdd.n3253 vdd.n315 146.341
R2093 vdd.n3253 vdd.n319 146.341
R2094 vdd.n3249 vdd.n319 146.341
R2095 vdd.n3249 vdd.n324 146.341
R2096 vdd.n3245 vdd.n324 146.341
R2097 vdd.n3245 vdd.n330 146.341
R2098 vdd.n3241 vdd.n330 146.341
R2099 vdd.n3241 vdd.n336 146.341
R2100 vdd.n3237 vdd.n336 146.341
R2101 vdd.n3237 vdd.n341 146.341
R2102 vdd.n3233 vdd.n341 146.341
R2103 vdd.n3233 vdd.n347 146.341
R2104 vdd.n3229 vdd.n347 146.341
R2105 vdd.n2090 vdd.n2089 146.341
R2106 vdd.n2087 vdd.n2084 146.341
R2107 vdd.n2082 vdd.n955 146.341
R2108 vdd.n2078 vdd.n2077 146.341
R2109 vdd.n2075 vdd.n959 146.341
R2110 vdd.n2071 vdd.n2070 146.341
R2111 vdd.n2068 vdd.n966 146.341
R2112 vdd.n2064 vdd.n2063 146.341
R2113 vdd.n2061 vdd.n973 146.341
R2114 vdd.n984 vdd.n981 146.341
R2115 vdd.n2053 vdd.n2052 146.341
R2116 vdd.n2050 vdd.n986 146.341
R2117 vdd.n2046 vdd.n2045 146.341
R2118 vdd.n2043 vdd.n992 146.341
R2119 vdd.n2039 vdd.n2038 146.341
R2120 vdd.n2036 vdd.n999 146.341
R2121 vdd.n2032 vdd.n2031 146.341
R2122 vdd.n2029 vdd.n1006 146.341
R2123 vdd.n2025 vdd.n2024 146.341
R2124 vdd.n2022 vdd.n1013 146.341
R2125 vdd.n1024 vdd.n1021 146.341
R2126 vdd.n2014 vdd.n2013 146.341
R2127 vdd.n2011 vdd.n1026 146.341
R2128 vdd.n2007 vdd.n2006 146.341
R2129 vdd.n2004 vdd.n1032 146.341
R2130 vdd.n2000 vdd.n1999 146.341
R2131 vdd.n1997 vdd.n1039 146.341
R2132 vdd.n1993 vdd.n1992 146.341
R2133 vdd.n1990 vdd.n1046 146.341
R2134 vdd.n1257 vdd.n1255 146.341
R2135 vdd.n1260 vdd.n1259 146.341
R2136 vdd.n1578 vdd.n1340 146.341
R2137 vdd.n1584 vdd.n1340 146.341
R2138 vdd.n1584 vdd.n1333 146.341
R2139 vdd.n1594 vdd.n1333 146.341
R2140 vdd.n1594 vdd.n1329 146.341
R2141 vdd.n1600 vdd.n1329 146.341
R2142 vdd.n1600 vdd.n1320 146.341
R2143 vdd.n1610 vdd.n1320 146.341
R2144 vdd.n1610 vdd.n1316 146.341
R2145 vdd.n1616 vdd.n1316 146.341
R2146 vdd.n1616 vdd.n1309 146.341
R2147 vdd.n1627 vdd.n1309 146.341
R2148 vdd.n1627 vdd.n1305 146.341
R2149 vdd.n1633 vdd.n1305 146.341
R2150 vdd.n1633 vdd.n1298 146.341
R2151 vdd.n1925 vdd.n1298 146.341
R2152 vdd.n1925 vdd.n1294 146.341
R2153 vdd.n1931 vdd.n1294 146.341
R2154 vdd.n1931 vdd.n1286 146.341
R2155 vdd.n1942 vdd.n1286 146.341
R2156 vdd.n1942 vdd.n1282 146.341
R2157 vdd.n1948 vdd.n1282 146.341
R2158 vdd.n1948 vdd.n1276 146.341
R2159 vdd.n1959 vdd.n1276 146.341
R2160 vdd.n1959 vdd.n1271 146.341
R2161 vdd.n1967 vdd.n1271 146.341
R2162 vdd.n1967 vdd.n1262 146.341
R2163 vdd.n1978 vdd.n1262 146.341
R2164 vdd.n1350 vdd.n1349 146.341
R2165 vdd.n1353 vdd.n1350 146.341
R2166 vdd.n1356 vdd.n1355 146.341
R2167 vdd.n1361 vdd.n1358 146.341
R2168 vdd.n1364 vdd.n1363 146.341
R2169 vdd.n1369 vdd.n1366 146.341
R2170 vdd.n1372 vdd.n1371 146.341
R2171 vdd.n1377 vdd.n1374 146.341
R2172 vdd.n1380 vdd.n1379 146.341
R2173 vdd.n1387 vdd.n1382 146.341
R2174 vdd.n1390 vdd.n1389 146.341
R2175 vdd.n1395 vdd.n1392 146.341
R2176 vdd.n1398 vdd.n1397 146.341
R2177 vdd.n1403 vdd.n1400 146.341
R2178 vdd.n1406 vdd.n1405 146.341
R2179 vdd.n1411 vdd.n1408 146.341
R2180 vdd.n1414 vdd.n1413 146.341
R2181 vdd.n1419 vdd.n1416 146.341
R2182 vdd.n1422 vdd.n1421 146.341
R2183 vdd.n1427 vdd.n1424 146.341
R2184 vdd.n1508 vdd.n1429 146.341
R2185 vdd.n1506 vdd.n1505 146.341
R2186 vdd.n1436 vdd.n1435 146.341
R2187 vdd.n1439 vdd.n1438 146.341
R2188 vdd.n1444 vdd.n1443 146.341
R2189 vdd.n1447 vdd.n1446 146.341
R2190 vdd.n1452 vdd.n1451 146.341
R2191 vdd.n1455 vdd.n1454 146.341
R2192 vdd.n1460 vdd.n1459 146.341
R2193 vdd.n1463 vdd.n1462 146.341
R2194 vdd.n1468 vdd.n1467 146.341
R2195 vdd.n1470 vdd.n1343 146.341
R2196 vdd.n1576 vdd.n1339 146.341
R2197 vdd.n1586 vdd.n1339 146.341
R2198 vdd.n1586 vdd.n1335 146.341
R2199 vdd.n1592 vdd.n1335 146.341
R2200 vdd.n1592 vdd.n1327 146.341
R2201 vdd.n1602 vdd.n1327 146.341
R2202 vdd.n1602 vdd.n1323 146.341
R2203 vdd.n1608 vdd.n1323 146.341
R2204 vdd.n1608 vdd.n1315 146.341
R2205 vdd.n1619 vdd.n1315 146.341
R2206 vdd.n1619 vdd.n1311 146.341
R2207 vdd.n1625 vdd.n1311 146.341
R2208 vdd.n1625 vdd.n1304 146.341
R2209 vdd.n1635 vdd.n1304 146.341
R2210 vdd.n1635 vdd.n1300 146.341
R2211 vdd.n1923 vdd.n1300 146.341
R2212 vdd.n1923 vdd.n1292 146.341
R2213 vdd.n1934 vdd.n1292 146.341
R2214 vdd.n1934 vdd.n1288 146.341
R2215 vdd.n1940 vdd.n1288 146.341
R2216 vdd.n1940 vdd.n1281 146.341
R2217 vdd.n1951 vdd.n1281 146.341
R2218 vdd.n1951 vdd.n1277 146.341
R2219 vdd.n1957 vdd.n1277 146.341
R2220 vdd.n1957 vdd.n1269 146.341
R2221 vdd.n1970 vdd.n1269 146.341
R2222 vdd.n1970 vdd.n1264 146.341
R2223 vdd.n1976 vdd.n1264 146.341
R2224 vdd.n1081 vdd.t38 127.284
R2225 vdd.n809 vdd.t79 127.284
R2226 vdd.n1101 vdd.t63 127.284
R2227 vdd.n800 vdd.t96 127.284
R2228 vdd.n700 vdd.t66 127.284
R2229 vdd.n700 vdd.t67 127.284
R2230 vdd.n2416 vdd.t91 127.284
R2231 vdd.n661 vdd.t102 127.284
R2232 vdd.n2413 vdd.t84 127.284
R2233 vdd.n625 vdd.t33 127.284
R2234 vdd.n871 vdd.t87 127.284
R2235 vdd.n871 vdd.t88 127.284
R2236 vdd.n22 vdd.n20 117.314
R2237 vdd.n17 vdd.n15 117.314
R2238 vdd.n27 vdd.n26 116.927
R2239 vdd.n24 vdd.n23 116.927
R2240 vdd.n22 vdd.n21 116.927
R2241 vdd.n17 vdd.n16 116.927
R2242 vdd.n19 vdd.n18 116.927
R2243 vdd.n27 vdd.n25 116.927
R2244 vdd.n1082 vdd.t37 111.188
R2245 vdd.n810 vdd.t80 111.188
R2246 vdd.n1102 vdd.t62 111.188
R2247 vdd.n801 vdd.t97 111.188
R2248 vdd.n2417 vdd.t90 111.188
R2249 vdd.n662 vdd.t103 111.188
R2250 vdd.n2414 vdd.t83 111.188
R2251 vdd.n626 vdd.t34 111.188
R2252 vdd.n2658 vdd.n755 99.5127
R2253 vdd.n2658 vdd.n753 99.5127
R2254 vdd.n2662 vdd.n753 99.5127
R2255 vdd.n2662 vdd.n744 99.5127
R2256 vdd.n2670 vdd.n744 99.5127
R2257 vdd.n2670 vdd.n742 99.5127
R2258 vdd.n2674 vdd.n742 99.5127
R2259 vdd.n2674 vdd.n732 99.5127
R2260 vdd.n2682 vdd.n732 99.5127
R2261 vdd.n2682 vdd.n730 99.5127
R2262 vdd.n2686 vdd.n730 99.5127
R2263 vdd.n2686 vdd.n720 99.5127
R2264 vdd.n2694 vdd.n720 99.5127
R2265 vdd.n2694 vdd.n718 99.5127
R2266 vdd.n2698 vdd.n718 99.5127
R2267 vdd.n2698 vdd.n709 99.5127
R2268 vdd.n2706 vdd.n709 99.5127
R2269 vdd.n2706 vdd.n707 99.5127
R2270 vdd.n2710 vdd.n707 99.5127
R2271 vdd.n2710 vdd.n695 99.5127
R2272 vdd.n2719 vdd.n695 99.5127
R2273 vdd.n2719 vdd.n693 99.5127
R2274 vdd.n2723 vdd.n693 99.5127
R2275 vdd.n2723 vdd.n684 99.5127
R2276 vdd.n2731 vdd.n684 99.5127
R2277 vdd.n2731 vdd.n682 99.5127
R2278 vdd.n2735 vdd.n682 99.5127
R2279 vdd.n2735 vdd.n670 99.5127
R2280 vdd.n2788 vdd.n670 99.5127
R2281 vdd.n2788 vdd.n668 99.5127
R2282 vdd.n2792 vdd.n668 99.5127
R2283 vdd.n2792 vdd.n634 99.5127
R2284 vdd.n2862 vdd.n634 99.5127
R2285 vdd.n2858 vdd.n635 99.5127
R2286 vdd.n2856 vdd.n2855 99.5127
R2287 vdd.n2853 vdd.n639 99.5127
R2288 vdd.n2849 vdd.n2848 99.5127
R2289 vdd.n2846 vdd.n642 99.5127
R2290 vdd.n2842 vdd.n2841 99.5127
R2291 vdd.n2839 vdd.n645 99.5127
R2292 vdd.n2835 vdd.n2834 99.5127
R2293 vdd.n2832 vdd.n648 99.5127
R2294 vdd.n2827 vdd.n2826 99.5127
R2295 vdd.n2824 vdd.n651 99.5127
R2296 vdd.n2820 vdd.n2819 99.5127
R2297 vdd.n2817 vdd.n654 99.5127
R2298 vdd.n2813 vdd.n2812 99.5127
R2299 vdd.n2810 vdd.n657 99.5127
R2300 vdd.n2806 vdd.n2805 99.5127
R2301 vdd.n2803 vdd.n660 99.5127
R2302 vdd.n2579 vdd.n757 99.5127
R2303 vdd.n2575 vdd.n757 99.5127
R2304 vdd.n2575 vdd.n751 99.5127
R2305 vdd.n2519 vdd.n751 99.5127
R2306 vdd.n2519 vdd.n746 99.5127
R2307 vdd.n2522 vdd.n746 99.5127
R2308 vdd.n2522 vdd.n740 99.5127
R2309 vdd.n2525 vdd.n740 99.5127
R2310 vdd.n2525 vdd.n734 99.5127
R2311 vdd.n2558 vdd.n734 99.5127
R2312 vdd.n2558 vdd.n727 99.5127
R2313 vdd.n2554 vdd.n727 99.5127
R2314 vdd.n2554 vdd.n721 99.5127
R2315 vdd.n2551 vdd.n721 99.5127
R2316 vdd.n2551 vdd.n716 99.5127
R2317 vdd.n2548 vdd.n716 99.5127
R2318 vdd.n2548 vdd.n711 99.5127
R2319 vdd.n2545 vdd.n711 99.5127
R2320 vdd.n2545 vdd.n704 99.5127
R2321 vdd.n2542 vdd.n704 99.5127
R2322 vdd.n2542 vdd.n696 99.5127
R2323 vdd.n2539 vdd.n696 99.5127
R2324 vdd.n2539 vdd.n691 99.5127
R2325 vdd.n2536 vdd.n691 99.5127
R2326 vdd.n2536 vdd.n686 99.5127
R2327 vdd.n2533 vdd.n686 99.5127
R2328 vdd.n2533 vdd.n680 99.5127
R2329 vdd.n2530 vdd.n680 99.5127
R2330 vdd.n2530 vdd.n672 99.5127
R2331 vdd.n672 vdd.n665 99.5127
R2332 vdd.n2794 vdd.n665 99.5127
R2333 vdd.n2795 vdd.n2794 99.5127
R2334 vdd.n2795 vdd.n632 99.5127
R2335 vdd.n2412 vdd.n2411 99.5127
R2336 vdd.n2643 vdd.n2411 99.5127
R2337 vdd.n2641 vdd.n2640 99.5127
R2338 vdd.n2637 vdd.n2636 99.5127
R2339 vdd.n2633 vdd.n2632 99.5127
R2340 vdd.n2629 vdd.n2628 99.5127
R2341 vdd.n2625 vdd.n2624 99.5127
R2342 vdd.n2621 vdd.n2620 99.5127
R2343 vdd.n2617 vdd.n2616 99.5127
R2344 vdd.n2613 vdd.n2612 99.5127
R2345 vdd.n2609 vdd.n2608 99.5127
R2346 vdd.n2605 vdd.n2604 99.5127
R2347 vdd.n2601 vdd.n2600 99.5127
R2348 vdd.n2597 vdd.n2596 99.5127
R2349 vdd.n2593 vdd.n2592 99.5127
R2350 vdd.n2589 vdd.n2588 99.5127
R2351 vdd.n2584 vdd.n2583 99.5127
R2352 vdd.n2376 vdd.n798 99.5127
R2353 vdd.n2372 vdd.n2371 99.5127
R2354 vdd.n2368 vdd.n2367 99.5127
R2355 vdd.n2364 vdd.n2363 99.5127
R2356 vdd.n2360 vdd.n2359 99.5127
R2357 vdd.n2356 vdd.n2355 99.5127
R2358 vdd.n2352 vdd.n2351 99.5127
R2359 vdd.n2348 vdd.n2347 99.5127
R2360 vdd.n2344 vdd.n2343 99.5127
R2361 vdd.n2340 vdd.n2339 99.5127
R2362 vdd.n2336 vdd.n2335 99.5127
R2363 vdd.n2332 vdd.n2331 99.5127
R2364 vdd.n2328 vdd.n2327 99.5127
R2365 vdd.n2324 vdd.n2323 99.5127
R2366 vdd.n2320 vdd.n2319 99.5127
R2367 vdd.n2316 vdd.n2315 99.5127
R2368 vdd.n2311 vdd.n2310 99.5127
R2369 vdd.n1137 vdd.n905 99.5127
R2370 vdd.n1140 vdd.n905 99.5127
R2371 vdd.n1140 vdd.n899 99.5127
R2372 vdd.n1143 vdd.n899 99.5127
R2373 vdd.n1143 vdd.n894 99.5127
R2374 vdd.n1146 vdd.n894 99.5127
R2375 vdd.n1146 vdd.n888 99.5127
R2376 vdd.n1149 vdd.n888 99.5127
R2377 vdd.n1149 vdd.n881 99.5127
R2378 vdd.n1152 vdd.n881 99.5127
R2379 vdd.n1152 vdd.n874 99.5127
R2380 vdd.n1155 vdd.n874 99.5127
R2381 vdd.n1155 vdd.n868 99.5127
R2382 vdd.n1158 vdd.n868 99.5127
R2383 vdd.n1158 vdd.n863 99.5127
R2384 vdd.n1161 vdd.n863 99.5127
R2385 vdd.n1161 vdd.n857 99.5127
R2386 vdd.n1186 vdd.n857 99.5127
R2387 vdd.n1186 vdd.n850 99.5127
R2388 vdd.n1182 vdd.n850 99.5127
R2389 vdd.n1182 vdd.n844 99.5127
R2390 vdd.n1179 vdd.n844 99.5127
R2391 vdd.n1179 vdd.n839 99.5127
R2392 vdd.n1176 vdd.n839 99.5127
R2393 vdd.n1176 vdd.n834 99.5127
R2394 vdd.n1173 vdd.n834 99.5127
R2395 vdd.n1173 vdd.n828 99.5127
R2396 vdd.n1170 vdd.n828 99.5127
R2397 vdd.n1170 vdd.n821 99.5127
R2398 vdd.n1167 vdd.n821 99.5127
R2399 vdd.n1167 vdd.n814 99.5127
R2400 vdd.n814 vdd.n803 99.5127
R2401 vdd.n2306 vdd.n803 99.5127
R2402 vdd.n946 vdd.n945 99.5127
R2403 vdd.n2122 vdd.n945 99.5127
R2404 vdd.n2120 vdd.n2119 99.5127
R2405 vdd.n2116 vdd.n2115 99.5127
R2406 vdd.n2112 vdd.n2111 99.5127
R2407 vdd.n2108 vdd.n2107 99.5127
R2408 vdd.n2104 vdd.n2103 99.5127
R2409 vdd.n2100 vdd.n2099 99.5127
R2410 vdd.n2096 vdd.n2095 99.5127
R2411 vdd.n1104 vdd.n1103 99.5127
R2412 vdd.n1108 vdd.n1107 99.5127
R2413 vdd.n1112 vdd.n1111 99.5127
R2414 vdd.n1116 vdd.n1115 99.5127
R2415 vdd.n1120 vdd.n1119 99.5127
R2416 vdd.n1124 vdd.n1123 99.5127
R2417 vdd.n1128 vdd.n1127 99.5127
R2418 vdd.n1133 vdd.n1132 99.5127
R2419 vdd.n2137 vdd.n903 99.5127
R2420 vdd.n2137 vdd.n901 99.5127
R2421 vdd.n2141 vdd.n901 99.5127
R2422 vdd.n2141 vdd.n892 99.5127
R2423 vdd.n2149 vdd.n892 99.5127
R2424 vdd.n2149 vdd.n890 99.5127
R2425 vdd.n2153 vdd.n890 99.5127
R2426 vdd.n2153 vdd.n879 99.5127
R2427 vdd.n2161 vdd.n879 99.5127
R2428 vdd.n2161 vdd.n877 99.5127
R2429 vdd.n2165 vdd.n877 99.5127
R2430 vdd.n2165 vdd.n867 99.5127
R2431 vdd.n2174 vdd.n867 99.5127
R2432 vdd.n2174 vdd.n865 99.5127
R2433 vdd.n2178 vdd.n865 99.5127
R2434 vdd.n2178 vdd.n855 99.5127
R2435 vdd.n2186 vdd.n855 99.5127
R2436 vdd.n2186 vdd.n853 99.5127
R2437 vdd.n2190 vdd.n853 99.5127
R2438 vdd.n2190 vdd.n843 99.5127
R2439 vdd.n2198 vdd.n843 99.5127
R2440 vdd.n2198 vdd.n841 99.5127
R2441 vdd.n2202 vdd.n841 99.5127
R2442 vdd.n2202 vdd.n832 99.5127
R2443 vdd.n2210 vdd.n832 99.5127
R2444 vdd.n2210 vdd.n830 99.5127
R2445 vdd.n2214 vdd.n830 99.5127
R2446 vdd.n2214 vdd.n819 99.5127
R2447 vdd.n2224 vdd.n819 99.5127
R2448 vdd.n2224 vdd.n816 99.5127
R2449 vdd.n2229 vdd.n816 99.5127
R2450 vdd.n2229 vdd.n817 99.5127
R2451 vdd.n817 vdd.n797 99.5127
R2452 vdd.n2778 vdd.n2777 99.5127
R2453 vdd.n2775 vdd.n2741 99.5127
R2454 vdd.n2771 vdd.n2770 99.5127
R2455 vdd.n2768 vdd.n2744 99.5127
R2456 vdd.n2764 vdd.n2763 99.5127
R2457 vdd.n2761 vdd.n2747 99.5127
R2458 vdd.n2757 vdd.n2756 99.5127
R2459 vdd.n2754 vdd.n2751 99.5127
R2460 vdd.n2895 vdd.n612 99.5127
R2461 vdd.n2893 vdd.n2892 99.5127
R2462 vdd.n2890 vdd.n615 99.5127
R2463 vdd.n2886 vdd.n2885 99.5127
R2464 vdd.n2883 vdd.n618 99.5127
R2465 vdd.n2879 vdd.n2878 99.5127
R2466 vdd.n2876 vdd.n621 99.5127
R2467 vdd.n2872 vdd.n2871 99.5127
R2468 vdd.n2869 vdd.n624 99.5127
R2469 vdd.n2484 vdd.n758 99.5127
R2470 vdd.n2573 vdd.n758 99.5127
R2471 vdd.n2573 vdd.n752 99.5127
R2472 vdd.n2569 vdd.n752 99.5127
R2473 vdd.n2569 vdd.n747 99.5127
R2474 vdd.n2566 vdd.n747 99.5127
R2475 vdd.n2566 vdd.n741 99.5127
R2476 vdd.n2563 vdd.n741 99.5127
R2477 vdd.n2563 vdd.n735 99.5127
R2478 vdd.n2560 vdd.n735 99.5127
R2479 vdd.n2560 vdd.n728 99.5127
R2480 vdd.n2516 vdd.n728 99.5127
R2481 vdd.n2516 vdd.n722 99.5127
R2482 vdd.n2513 vdd.n722 99.5127
R2483 vdd.n2513 vdd.n717 99.5127
R2484 vdd.n2510 vdd.n717 99.5127
R2485 vdd.n2510 vdd.n712 99.5127
R2486 vdd.n2507 vdd.n712 99.5127
R2487 vdd.n2507 vdd.n705 99.5127
R2488 vdd.n2504 vdd.n705 99.5127
R2489 vdd.n2504 vdd.n697 99.5127
R2490 vdd.n2501 vdd.n697 99.5127
R2491 vdd.n2501 vdd.n692 99.5127
R2492 vdd.n2498 vdd.n692 99.5127
R2493 vdd.n2498 vdd.n687 99.5127
R2494 vdd.n2495 vdd.n687 99.5127
R2495 vdd.n2495 vdd.n681 99.5127
R2496 vdd.n2492 vdd.n681 99.5127
R2497 vdd.n2492 vdd.n673 99.5127
R2498 vdd.n2489 vdd.n673 99.5127
R2499 vdd.n2489 vdd.n666 99.5127
R2500 vdd.n666 vdd.n630 99.5127
R2501 vdd.n2864 vdd.n630 99.5127
R2502 vdd.n2419 vdd.n761 99.5127
R2503 vdd.n2423 vdd.n2422 99.5127
R2504 vdd.n2427 vdd.n2426 99.5127
R2505 vdd.n2431 vdd.n2430 99.5127
R2506 vdd.n2435 vdd.n2434 99.5127
R2507 vdd.n2439 vdd.n2438 99.5127
R2508 vdd.n2443 vdd.n2442 99.5127
R2509 vdd.n2447 vdd.n2446 99.5127
R2510 vdd.n2451 vdd.n2450 99.5127
R2511 vdd.n2455 vdd.n2454 99.5127
R2512 vdd.n2459 vdd.n2458 99.5127
R2513 vdd.n2463 vdd.n2462 99.5127
R2514 vdd.n2467 vdd.n2466 99.5127
R2515 vdd.n2471 vdd.n2470 99.5127
R2516 vdd.n2475 vdd.n2474 99.5127
R2517 vdd.n2479 vdd.n2478 99.5127
R2518 vdd.n2481 vdd.n2410 99.5127
R2519 vdd.n2656 vdd.n759 99.5127
R2520 vdd.n2656 vdd.n750 99.5127
R2521 vdd.n2664 vdd.n750 99.5127
R2522 vdd.n2664 vdd.n748 99.5127
R2523 vdd.n2668 vdd.n748 99.5127
R2524 vdd.n2668 vdd.n738 99.5127
R2525 vdd.n2676 vdd.n738 99.5127
R2526 vdd.n2676 vdd.n736 99.5127
R2527 vdd.n2680 vdd.n736 99.5127
R2528 vdd.n2680 vdd.n726 99.5127
R2529 vdd.n2688 vdd.n726 99.5127
R2530 vdd.n2688 vdd.n724 99.5127
R2531 vdd.n2692 vdd.n724 99.5127
R2532 vdd.n2692 vdd.n715 99.5127
R2533 vdd.n2700 vdd.n715 99.5127
R2534 vdd.n2700 vdd.n713 99.5127
R2535 vdd.n2704 vdd.n713 99.5127
R2536 vdd.n2704 vdd.n702 99.5127
R2537 vdd.n2712 vdd.n702 99.5127
R2538 vdd.n2712 vdd.n699 99.5127
R2539 vdd.n2717 vdd.n699 99.5127
R2540 vdd.n2717 vdd.n690 99.5127
R2541 vdd.n2725 vdd.n690 99.5127
R2542 vdd.n2725 vdd.n688 99.5127
R2543 vdd.n2729 vdd.n688 99.5127
R2544 vdd.n2729 vdd.n678 99.5127
R2545 vdd.n2737 vdd.n678 99.5127
R2546 vdd.n2737 vdd.n675 99.5127
R2547 vdd.n2786 vdd.n675 99.5127
R2548 vdd.n2786 vdd.n676 99.5127
R2549 vdd.n676 vdd.n667 99.5127
R2550 vdd.n2781 vdd.n667 99.5127
R2551 vdd.n2781 vdd.n633 99.5127
R2552 vdd.n2300 vdd.n2299 99.5127
R2553 vdd.n2296 vdd.n2295 99.5127
R2554 vdd.n2292 vdd.n2291 99.5127
R2555 vdd.n2288 vdd.n2287 99.5127
R2556 vdd.n2284 vdd.n2283 99.5127
R2557 vdd.n2280 vdd.n2279 99.5127
R2558 vdd.n2276 vdd.n2275 99.5127
R2559 vdd.n2272 vdd.n2271 99.5127
R2560 vdd.n2268 vdd.n2267 99.5127
R2561 vdd.n2264 vdd.n2263 99.5127
R2562 vdd.n2260 vdd.n2259 99.5127
R2563 vdd.n2256 vdd.n2255 99.5127
R2564 vdd.n2252 vdd.n2251 99.5127
R2565 vdd.n2248 vdd.n2247 99.5127
R2566 vdd.n2244 vdd.n2243 99.5127
R2567 vdd.n2240 vdd.n2239 99.5127
R2568 vdd.n2236 vdd.n779 99.5127
R2569 vdd.n1215 vdd.n906 99.5127
R2570 vdd.n1212 vdd.n906 99.5127
R2571 vdd.n1212 vdd.n900 99.5127
R2572 vdd.n1209 vdd.n900 99.5127
R2573 vdd.n1209 vdd.n895 99.5127
R2574 vdd.n1206 vdd.n895 99.5127
R2575 vdd.n1206 vdd.n889 99.5127
R2576 vdd.n1203 vdd.n889 99.5127
R2577 vdd.n1203 vdd.n882 99.5127
R2578 vdd.n1200 vdd.n882 99.5127
R2579 vdd.n1200 vdd.n875 99.5127
R2580 vdd.n1197 vdd.n875 99.5127
R2581 vdd.n1197 vdd.n869 99.5127
R2582 vdd.n1194 vdd.n869 99.5127
R2583 vdd.n1194 vdd.n864 99.5127
R2584 vdd.n1191 vdd.n864 99.5127
R2585 vdd.n1191 vdd.n858 99.5127
R2586 vdd.n1188 vdd.n858 99.5127
R2587 vdd.n1188 vdd.n851 99.5127
R2588 vdd.n1098 vdd.n851 99.5127
R2589 vdd.n1098 vdd.n845 99.5127
R2590 vdd.n1095 vdd.n845 99.5127
R2591 vdd.n1095 vdd.n840 99.5127
R2592 vdd.n1092 vdd.n840 99.5127
R2593 vdd.n1092 vdd.n835 99.5127
R2594 vdd.n1089 vdd.n835 99.5127
R2595 vdd.n1089 vdd.n829 99.5127
R2596 vdd.n1086 vdd.n829 99.5127
R2597 vdd.n1086 vdd.n822 99.5127
R2598 vdd.n822 vdd.n813 99.5127
R2599 vdd.n2231 vdd.n813 99.5127
R2600 vdd.n2232 vdd.n2231 99.5127
R2601 vdd.n2232 vdd.n805 99.5127
R2602 vdd.n1050 vdd.n910 99.5127
R2603 vdd.n1054 vdd.n1053 99.5127
R2604 vdd.n1058 vdd.n1057 99.5127
R2605 vdd.n1062 vdd.n1061 99.5127
R2606 vdd.n1066 vdd.n1065 99.5127
R2607 vdd.n1070 vdd.n1069 99.5127
R2608 vdd.n1074 vdd.n1073 99.5127
R2609 vdd.n1078 vdd.n1077 99.5127
R2610 vdd.n1248 vdd.n1080 99.5127
R2611 vdd.n1246 vdd.n1245 99.5127
R2612 vdd.n1242 vdd.n1241 99.5127
R2613 vdd.n1238 vdd.n1237 99.5127
R2614 vdd.n1234 vdd.n1233 99.5127
R2615 vdd.n1230 vdd.n1229 99.5127
R2616 vdd.n1226 vdd.n1225 99.5127
R2617 vdd.n1222 vdd.n1221 99.5127
R2618 vdd.n1218 vdd.n944 99.5127
R2619 vdd.n2135 vdd.n908 99.5127
R2620 vdd.n2135 vdd.n898 99.5127
R2621 vdd.n2143 vdd.n898 99.5127
R2622 vdd.n2143 vdd.n896 99.5127
R2623 vdd.n2147 vdd.n896 99.5127
R2624 vdd.n2147 vdd.n886 99.5127
R2625 vdd.n2155 vdd.n886 99.5127
R2626 vdd.n2155 vdd.n884 99.5127
R2627 vdd.n2159 vdd.n884 99.5127
R2628 vdd.n2159 vdd.n873 99.5127
R2629 vdd.n2167 vdd.n873 99.5127
R2630 vdd.n2167 vdd.n870 99.5127
R2631 vdd.n2172 vdd.n870 99.5127
R2632 vdd.n2172 vdd.n861 99.5127
R2633 vdd.n2180 vdd.n861 99.5127
R2634 vdd.n2180 vdd.n859 99.5127
R2635 vdd.n2184 vdd.n859 99.5127
R2636 vdd.n2184 vdd.n849 99.5127
R2637 vdd.n2192 vdd.n849 99.5127
R2638 vdd.n2192 vdd.n847 99.5127
R2639 vdd.n2196 vdd.n847 99.5127
R2640 vdd.n2196 vdd.n838 99.5127
R2641 vdd.n2204 vdd.n838 99.5127
R2642 vdd.n2204 vdd.n836 99.5127
R2643 vdd.n2208 vdd.n836 99.5127
R2644 vdd.n2208 vdd.n826 99.5127
R2645 vdd.n2216 vdd.n826 99.5127
R2646 vdd.n2216 vdd.n823 99.5127
R2647 vdd.n2222 vdd.n823 99.5127
R2648 vdd.n2222 vdd.n824 99.5127
R2649 vdd.n824 vdd.n815 99.5127
R2650 vdd.n815 vdd.n806 99.5127
R2651 vdd.n2304 vdd.n806 99.5127
R2652 vdd.n9 vdd.n7 98.9633
R2653 vdd.n2 vdd.n0 98.9633
R2654 vdd.n9 vdd.n8 98.6055
R2655 vdd.n11 vdd.n10 98.6055
R2656 vdd.n13 vdd.n12 98.6055
R2657 vdd.n6 vdd.n5 98.6055
R2658 vdd.n4 vdd.n3 98.6055
R2659 vdd.n2 vdd.n1 98.6055
R2660 vdd.t219 vdd.n279 85.8723
R2661 vdd.t201 vdd.n228 85.8723
R2662 vdd.t210 vdd.n185 85.8723
R2663 vdd.t193 vdd.n134 85.8723
R2664 vdd.t160 vdd.n92 85.8723
R2665 vdd.t167 vdd.n41 85.8723
R2666 vdd.t225 vdd.n1836 85.8723
R2667 vdd.t163 vdd.n1887 85.8723
R2668 vdd.t216 vdd.n1742 85.8723
R2669 vdd.t149 vdd.n1793 85.8723
R2670 vdd.t169 vdd.n1649 85.8723
R2671 vdd.t161 vdd.n1700 85.8723
R2672 vdd.n2715 vdd.n700 78.546
R2673 vdd.n2170 vdd.n871 78.546
R2674 vdd.n266 vdd.n265 75.1835
R2675 vdd.n264 vdd.n263 75.1835
R2676 vdd.n262 vdd.n261 75.1835
R2677 vdd.n260 vdd.n259 75.1835
R2678 vdd.n258 vdd.n257 75.1835
R2679 vdd.n172 vdd.n171 75.1835
R2680 vdd.n170 vdd.n169 75.1835
R2681 vdd.n168 vdd.n167 75.1835
R2682 vdd.n166 vdd.n165 75.1835
R2683 vdd.n164 vdd.n163 75.1835
R2684 vdd.n79 vdd.n78 75.1835
R2685 vdd.n77 vdd.n76 75.1835
R2686 vdd.n75 vdd.n74 75.1835
R2687 vdd.n73 vdd.n72 75.1835
R2688 vdd.n71 vdd.n70 75.1835
R2689 vdd.n1866 vdd.n1865 75.1835
R2690 vdd.n1868 vdd.n1867 75.1835
R2691 vdd.n1870 vdd.n1869 75.1835
R2692 vdd.n1872 vdd.n1871 75.1835
R2693 vdd.n1874 vdd.n1873 75.1835
R2694 vdd.n1772 vdd.n1771 75.1835
R2695 vdd.n1774 vdd.n1773 75.1835
R2696 vdd.n1776 vdd.n1775 75.1835
R2697 vdd.n1778 vdd.n1777 75.1835
R2698 vdd.n1780 vdd.n1779 75.1835
R2699 vdd.n1679 vdd.n1678 75.1835
R2700 vdd.n1681 vdd.n1680 75.1835
R2701 vdd.n1683 vdd.n1682 75.1835
R2702 vdd.n1685 vdd.n1684 75.1835
R2703 vdd.n1687 vdd.n1686 75.1835
R2704 vdd.n2651 vdd.n2650 72.8958
R2705 vdd.n2650 vdd.n2394 72.8958
R2706 vdd.n2650 vdd.n2395 72.8958
R2707 vdd.n2650 vdd.n2396 72.8958
R2708 vdd.n2650 vdd.n2397 72.8958
R2709 vdd.n2650 vdd.n2398 72.8958
R2710 vdd.n2650 vdd.n2399 72.8958
R2711 vdd.n2650 vdd.n2400 72.8958
R2712 vdd.n2650 vdd.n2401 72.8958
R2713 vdd.n2650 vdd.n2402 72.8958
R2714 vdd.n2650 vdd.n2403 72.8958
R2715 vdd.n2650 vdd.n2404 72.8958
R2716 vdd.n2650 vdd.n2405 72.8958
R2717 vdd.n2650 vdd.n2406 72.8958
R2718 vdd.n2650 vdd.n2407 72.8958
R2719 vdd.n2650 vdd.n2408 72.8958
R2720 vdd.n2650 vdd.n2409 72.8958
R2721 vdd.n629 vdd.n613 72.8958
R2722 vdd.n2870 vdd.n613 72.8958
R2723 vdd.n623 vdd.n613 72.8958
R2724 vdd.n2877 vdd.n613 72.8958
R2725 vdd.n620 vdd.n613 72.8958
R2726 vdd.n2884 vdd.n613 72.8958
R2727 vdd.n617 vdd.n613 72.8958
R2728 vdd.n2891 vdd.n613 72.8958
R2729 vdd.n2894 vdd.n613 72.8958
R2730 vdd.n2750 vdd.n613 72.8958
R2731 vdd.n2755 vdd.n613 72.8958
R2732 vdd.n2749 vdd.n613 72.8958
R2733 vdd.n2762 vdd.n613 72.8958
R2734 vdd.n2746 vdd.n613 72.8958
R2735 vdd.n2769 vdd.n613 72.8958
R2736 vdd.n2743 vdd.n613 72.8958
R2737 vdd.n2776 vdd.n613 72.8958
R2738 vdd.n2129 vdd.n2128 72.8958
R2739 vdd.n2129 vdd.n912 72.8958
R2740 vdd.n2129 vdd.n913 72.8958
R2741 vdd.n2129 vdd.n914 72.8958
R2742 vdd.n2129 vdd.n915 72.8958
R2743 vdd.n2129 vdd.n916 72.8958
R2744 vdd.n2129 vdd.n917 72.8958
R2745 vdd.n2129 vdd.n918 72.8958
R2746 vdd.n2129 vdd.n919 72.8958
R2747 vdd.n2129 vdd.n920 72.8958
R2748 vdd.n2129 vdd.n921 72.8958
R2749 vdd.n2129 vdd.n922 72.8958
R2750 vdd.n2129 vdd.n923 72.8958
R2751 vdd.n2129 vdd.n924 72.8958
R2752 vdd.n2129 vdd.n925 72.8958
R2753 vdd.n2129 vdd.n926 72.8958
R2754 vdd.n2129 vdd.n927 72.8958
R2755 vdd.n2377 vdd.n780 72.8958
R2756 vdd.n2377 vdd.n781 72.8958
R2757 vdd.n2377 vdd.n782 72.8958
R2758 vdd.n2377 vdd.n783 72.8958
R2759 vdd.n2377 vdd.n784 72.8958
R2760 vdd.n2377 vdd.n785 72.8958
R2761 vdd.n2377 vdd.n786 72.8958
R2762 vdd.n2377 vdd.n787 72.8958
R2763 vdd.n2377 vdd.n788 72.8958
R2764 vdd.n2377 vdd.n789 72.8958
R2765 vdd.n2377 vdd.n790 72.8958
R2766 vdd.n2377 vdd.n791 72.8958
R2767 vdd.n2377 vdd.n792 72.8958
R2768 vdd.n2377 vdd.n793 72.8958
R2769 vdd.n2377 vdd.n794 72.8958
R2770 vdd.n2377 vdd.n795 72.8958
R2771 vdd.n2377 vdd.n796 72.8958
R2772 vdd.n2650 vdd.n2649 72.8958
R2773 vdd.n2650 vdd.n2378 72.8958
R2774 vdd.n2650 vdd.n2379 72.8958
R2775 vdd.n2650 vdd.n2380 72.8958
R2776 vdd.n2650 vdd.n2381 72.8958
R2777 vdd.n2650 vdd.n2382 72.8958
R2778 vdd.n2650 vdd.n2383 72.8958
R2779 vdd.n2650 vdd.n2384 72.8958
R2780 vdd.n2650 vdd.n2385 72.8958
R2781 vdd.n2650 vdd.n2386 72.8958
R2782 vdd.n2650 vdd.n2387 72.8958
R2783 vdd.n2650 vdd.n2388 72.8958
R2784 vdd.n2650 vdd.n2389 72.8958
R2785 vdd.n2650 vdd.n2390 72.8958
R2786 vdd.n2650 vdd.n2391 72.8958
R2787 vdd.n2650 vdd.n2392 72.8958
R2788 vdd.n2650 vdd.n2393 72.8958
R2789 vdd.n2798 vdd.n613 72.8958
R2790 vdd.n2804 vdd.n613 72.8958
R2791 vdd.n659 vdd.n613 72.8958
R2792 vdd.n2811 vdd.n613 72.8958
R2793 vdd.n656 vdd.n613 72.8958
R2794 vdd.n2818 vdd.n613 72.8958
R2795 vdd.n653 vdd.n613 72.8958
R2796 vdd.n2825 vdd.n613 72.8958
R2797 vdd.n650 vdd.n613 72.8958
R2798 vdd.n2833 vdd.n613 72.8958
R2799 vdd.n647 vdd.n613 72.8958
R2800 vdd.n2840 vdd.n613 72.8958
R2801 vdd.n644 vdd.n613 72.8958
R2802 vdd.n2847 vdd.n613 72.8958
R2803 vdd.n641 vdd.n613 72.8958
R2804 vdd.n2854 vdd.n613 72.8958
R2805 vdd.n2857 vdd.n613 72.8958
R2806 vdd.n2377 vdd.n778 72.8958
R2807 vdd.n2377 vdd.n777 72.8958
R2808 vdd.n2377 vdd.n776 72.8958
R2809 vdd.n2377 vdd.n775 72.8958
R2810 vdd.n2377 vdd.n774 72.8958
R2811 vdd.n2377 vdd.n773 72.8958
R2812 vdd.n2377 vdd.n772 72.8958
R2813 vdd.n2377 vdd.n771 72.8958
R2814 vdd.n2377 vdd.n770 72.8958
R2815 vdd.n2377 vdd.n769 72.8958
R2816 vdd.n2377 vdd.n768 72.8958
R2817 vdd.n2377 vdd.n767 72.8958
R2818 vdd.n2377 vdd.n766 72.8958
R2819 vdd.n2377 vdd.n765 72.8958
R2820 vdd.n2377 vdd.n764 72.8958
R2821 vdd.n2377 vdd.n763 72.8958
R2822 vdd.n2377 vdd.n762 72.8958
R2823 vdd.n2130 vdd.n2129 72.8958
R2824 vdd.n2129 vdd.n928 72.8958
R2825 vdd.n2129 vdd.n929 72.8958
R2826 vdd.n2129 vdd.n930 72.8958
R2827 vdd.n2129 vdd.n931 72.8958
R2828 vdd.n2129 vdd.n932 72.8958
R2829 vdd.n2129 vdd.n933 72.8958
R2830 vdd.n2129 vdd.n934 72.8958
R2831 vdd.n2129 vdd.n935 72.8958
R2832 vdd.n2129 vdd.n936 72.8958
R2833 vdd.n2129 vdd.n937 72.8958
R2834 vdd.n2129 vdd.n938 72.8958
R2835 vdd.n2129 vdd.n939 72.8958
R2836 vdd.n2129 vdd.n940 72.8958
R2837 vdd.n2129 vdd.n941 72.8958
R2838 vdd.n2129 vdd.n942 72.8958
R2839 vdd.n2129 vdd.n943 72.8958
R2840 vdd.n1348 vdd.n1344 66.2847
R2841 vdd.n1354 vdd.n1344 66.2847
R2842 vdd.n1357 vdd.n1344 66.2847
R2843 vdd.n1362 vdd.n1344 66.2847
R2844 vdd.n1365 vdd.n1344 66.2847
R2845 vdd.n1370 vdd.n1344 66.2847
R2846 vdd.n1373 vdd.n1344 66.2847
R2847 vdd.n1378 vdd.n1344 66.2847
R2848 vdd.n1381 vdd.n1344 66.2847
R2849 vdd.n1388 vdd.n1344 66.2847
R2850 vdd.n1391 vdd.n1344 66.2847
R2851 vdd.n1396 vdd.n1344 66.2847
R2852 vdd.n1399 vdd.n1344 66.2847
R2853 vdd.n1404 vdd.n1344 66.2847
R2854 vdd.n1407 vdd.n1344 66.2847
R2855 vdd.n1412 vdd.n1344 66.2847
R2856 vdd.n1415 vdd.n1344 66.2847
R2857 vdd.n1420 vdd.n1344 66.2847
R2858 vdd.n1423 vdd.n1344 66.2847
R2859 vdd.n1428 vdd.n1344 66.2847
R2860 vdd.n1507 vdd.n1344 66.2847
R2861 vdd.n1431 vdd.n1344 66.2847
R2862 vdd.n1437 vdd.n1344 66.2847
R2863 vdd.n1442 vdd.n1344 66.2847
R2864 vdd.n1445 vdd.n1344 66.2847
R2865 vdd.n1450 vdd.n1344 66.2847
R2866 vdd.n1453 vdd.n1344 66.2847
R2867 vdd.n1458 vdd.n1344 66.2847
R2868 vdd.n1461 vdd.n1344 66.2847
R2869 vdd.n1466 vdd.n1344 66.2847
R2870 vdd.n1469 vdd.n1344 66.2847
R2871 vdd.n1261 vdd.n911 66.2847
R2872 vdd.n1258 vdd.n911 66.2847
R2873 vdd.n1254 vdd.n911 66.2847
R2874 vdd.n1991 vdd.n911 66.2847
R2875 vdd.n1045 vdd.n911 66.2847
R2876 vdd.n1998 vdd.n911 66.2847
R2877 vdd.n1038 vdd.n911 66.2847
R2878 vdd.n2005 vdd.n911 66.2847
R2879 vdd.n1031 vdd.n911 66.2847
R2880 vdd.n2012 vdd.n911 66.2847
R2881 vdd.n1025 vdd.n911 66.2847
R2882 vdd.n1020 vdd.n911 66.2847
R2883 vdd.n2023 vdd.n911 66.2847
R2884 vdd.n1012 vdd.n911 66.2847
R2885 vdd.n2030 vdd.n911 66.2847
R2886 vdd.n1005 vdd.n911 66.2847
R2887 vdd.n2037 vdd.n911 66.2847
R2888 vdd.n998 vdd.n911 66.2847
R2889 vdd.n2044 vdd.n911 66.2847
R2890 vdd.n991 vdd.n911 66.2847
R2891 vdd.n2051 vdd.n911 66.2847
R2892 vdd.n985 vdd.n911 66.2847
R2893 vdd.n980 vdd.n911 66.2847
R2894 vdd.n2062 vdd.n911 66.2847
R2895 vdd.n972 vdd.n911 66.2847
R2896 vdd.n2069 vdd.n911 66.2847
R2897 vdd.n965 vdd.n911 66.2847
R2898 vdd.n2076 vdd.n911 66.2847
R2899 vdd.n958 vdd.n911 66.2847
R2900 vdd.n2083 vdd.n911 66.2847
R2901 vdd.n2088 vdd.n911 66.2847
R2902 vdd.n954 vdd.n911 66.2847
R2903 vdd.n3024 vdd.n516 66.2847
R2904 vdd.n520 vdd.n516 66.2847
R2905 vdd.n523 vdd.n516 66.2847
R2906 vdd.n3013 vdd.n516 66.2847
R2907 vdd.n3007 vdd.n516 66.2847
R2908 vdd.n3005 vdd.n516 66.2847
R2909 vdd.n2999 vdd.n516 66.2847
R2910 vdd.n2997 vdd.n516 66.2847
R2911 vdd.n2991 vdd.n516 66.2847
R2912 vdd.n2989 vdd.n516 66.2847
R2913 vdd.n2983 vdd.n516 66.2847
R2914 vdd.n2981 vdd.n516 66.2847
R2915 vdd.n2975 vdd.n516 66.2847
R2916 vdd.n2973 vdd.n516 66.2847
R2917 vdd.n2967 vdd.n516 66.2847
R2918 vdd.n2965 vdd.n516 66.2847
R2919 vdd.n2959 vdd.n516 66.2847
R2920 vdd.n2957 vdd.n516 66.2847
R2921 vdd.n2951 vdd.n516 66.2847
R2922 vdd.n2949 vdd.n516 66.2847
R2923 vdd.n584 vdd.n516 66.2847
R2924 vdd.n2940 vdd.n516 66.2847
R2925 vdd.n586 vdd.n516 66.2847
R2926 vdd.n2933 vdd.n516 66.2847
R2927 vdd.n2927 vdd.n516 66.2847
R2928 vdd.n2925 vdd.n516 66.2847
R2929 vdd.n2919 vdd.n516 66.2847
R2930 vdd.n2917 vdd.n516 66.2847
R2931 vdd.n2911 vdd.n516 66.2847
R2932 vdd.n607 vdd.n516 66.2847
R2933 vdd.n609 vdd.n516 66.2847
R2934 vdd.n3110 vdd.n351 66.2847
R2935 vdd.n3119 vdd.n351 66.2847
R2936 vdd.n461 vdd.n351 66.2847
R2937 vdd.n3126 vdd.n351 66.2847
R2938 vdd.n454 vdd.n351 66.2847
R2939 vdd.n3133 vdd.n351 66.2847
R2940 vdd.n447 vdd.n351 66.2847
R2941 vdd.n3140 vdd.n351 66.2847
R2942 vdd.n440 vdd.n351 66.2847
R2943 vdd.n3147 vdd.n351 66.2847
R2944 vdd.n434 vdd.n351 66.2847
R2945 vdd.n429 vdd.n351 66.2847
R2946 vdd.n3158 vdd.n351 66.2847
R2947 vdd.n421 vdd.n351 66.2847
R2948 vdd.n3165 vdd.n351 66.2847
R2949 vdd.n414 vdd.n351 66.2847
R2950 vdd.n3172 vdd.n351 66.2847
R2951 vdd.n407 vdd.n351 66.2847
R2952 vdd.n3179 vdd.n351 66.2847
R2953 vdd.n400 vdd.n351 66.2847
R2954 vdd.n3186 vdd.n351 66.2847
R2955 vdd.n394 vdd.n351 66.2847
R2956 vdd.n389 vdd.n351 66.2847
R2957 vdd.n3197 vdd.n351 66.2847
R2958 vdd.n381 vdd.n351 66.2847
R2959 vdd.n3204 vdd.n351 66.2847
R2960 vdd.n374 vdd.n351 66.2847
R2961 vdd.n3211 vdd.n351 66.2847
R2962 vdd.n367 vdd.n351 66.2847
R2963 vdd.n3218 vdd.n351 66.2847
R2964 vdd.n3221 vdd.n351 66.2847
R2965 vdd.n355 vdd.n351 66.2847
R2966 vdd.n356 vdd.n355 52.4337
R2967 vdd.n3221 vdd.n3220 52.4337
R2968 vdd.n3218 vdd.n3217 52.4337
R2969 vdd.n3213 vdd.n367 52.4337
R2970 vdd.n3211 vdd.n3210 52.4337
R2971 vdd.n3206 vdd.n374 52.4337
R2972 vdd.n3204 vdd.n3203 52.4337
R2973 vdd.n3199 vdd.n381 52.4337
R2974 vdd.n3197 vdd.n3196 52.4337
R2975 vdd.n390 vdd.n389 52.4337
R2976 vdd.n3188 vdd.n394 52.4337
R2977 vdd.n3186 vdd.n3185 52.4337
R2978 vdd.n3181 vdd.n400 52.4337
R2979 vdd.n3179 vdd.n3178 52.4337
R2980 vdd.n3174 vdd.n407 52.4337
R2981 vdd.n3172 vdd.n3171 52.4337
R2982 vdd.n3167 vdd.n414 52.4337
R2983 vdd.n3165 vdd.n3164 52.4337
R2984 vdd.n3160 vdd.n421 52.4337
R2985 vdd.n3158 vdd.n3157 52.4337
R2986 vdd.n430 vdd.n429 52.4337
R2987 vdd.n3149 vdd.n434 52.4337
R2988 vdd.n3147 vdd.n3146 52.4337
R2989 vdd.n3142 vdd.n440 52.4337
R2990 vdd.n3140 vdd.n3139 52.4337
R2991 vdd.n3135 vdd.n447 52.4337
R2992 vdd.n3133 vdd.n3132 52.4337
R2993 vdd.n3128 vdd.n454 52.4337
R2994 vdd.n3126 vdd.n3125 52.4337
R2995 vdd.n3121 vdd.n461 52.4337
R2996 vdd.n3119 vdd.n3118 52.4337
R2997 vdd.n3111 vdd.n3110 52.4337
R2998 vdd.n3024 vdd.n517 52.4337
R2999 vdd.n3022 vdd.n520 52.4337
R3000 vdd.n3018 vdd.n523 52.4337
R3001 vdd.n3014 vdd.n3013 52.4337
R3002 vdd.n3007 vdd.n526 52.4337
R3003 vdd.n3006 vdd.n3005 52.4337
R3004 vdd.n2999 vdd.n532 52.4337
R3005 vdd.n2998 vdd.n2997 52.4337
R3006 vdd.n2991 vdd.n538 52.4337
R3007 vdd.n2990 vdd.n2989 52.4337
R3008 vdd.n2983 vdd.n546 52.4337
R3009 vdd.n2982 vdd.n2981 52.4337
R3010 vdd.n2975 vdd.n552 52.4337
R3011 vdd.n2974 vdd.n2973 52.4337
R3012 vdd.n2967 vdd.n558 52.4337
R3013 vdd.n2966 vdd.n2965 52.4337
R3014 vdd.n2959 vdd.n564 52.4337
R3015 vdd.n2958 vdd.n2957 52.4337
R3016 vdd.n2951 vdd.n570 52.4337
R3017 vdd.n2950 vdd.n2949 52.4337
R3018 vdd.n584 vdd.n576 52.4337
R3019 vdd.n2941 vdd.n2940 52.4337
R3020 vdd.n2938 vdd.n586 52.4337
R3021 vdd.n2934 vdd.n2933 52.4337
R3022 vdd.n2927 vdd.n590 52.4337
R3023 vdd.n2926 vdd.n2925 52.4337
R3024 vdd.n2919 vdd.n596 52.4337
R3025 vdd.n2918 vdd.n2917 52.4337
R3026 vdd.n2911 vdd.n602 52.4337
R3027 vdd.n2910 vdd.n607 52.4337
R3028 vdd.n2906 vdd.n609 52.4337
R3029 vdd.n2090 vdd.n954 52.4337
R3030 vdd.n2088 vdd.n2087 52.4337
R3031 vdd.n2083 vdd.n2082 52.4337
R3032 vdd.n2078 vdd.n958 52.4337
R3033 vdd.n2076 vdd.n2075 52.4337
R3034 vdd.n2071 vdd.n965 52.4337
R3035 vdd.n2069 vdd.n2068 52.4337
R3036 vdd.n2064 vdd.n972 52.4337
R3037 vdd.n2062 vdd.n2061 52.4337
R3038 vdd.n981 vdd.n980 52.4337
R3039 vdd.n2053 vdd.n985 52.4337
R3040 vdd.n2051 vdd.n2050 52.4337
R3041 vdd.n2046 vdd.n991 52.4337
R3042 vdd.n2044 vdd.n2043 52.4337
R3043 vdd.n2039 vdd.n998 52.4337
R3044 vdd.n2037 vdd.n2036 52.4337
R3045 vdd.n2032 vdd.n1005 52.4337
R3046 vdd.n2030 vdd.n2029 52.4337
R3047 vdd.n2025 vdd.n1012 52.4337
R3048 vdd.n2023 vdd.n2022 52.4337
R3049 vdd.n1021 vdd.n1020 52.4337
R3050 vdd.n2014 vdd.n1025 52.4337
R3051 vdd.n2012 vdd.n2011 52.4337
R3052 vdd.n2007 vdd.n1031 52.4337
R3053 vdd.n2005 vdd.n2004 52.4337
R3054 vdd.n2000 vdd.n1038 52.4337
R3055 vdd.n1998 vdd.n1997 52.4337
R3056 vdd.n1993 vdd.n1045 52.4337
R3057 vdd.n1991 vdd.n1990 52.4337
R3058 vdd.n1255 vdd.n1254 52.4337
R3059 vdd.n1259 vdd.n1258 52.4337
R3060 vdd.n1979 vdd.n1261 52.4337
R3061 vdd.n1348 vdd.n1346 52.4337
R3062 vdd.n1354 vdd.n1353 52.4337
R3063 vdd.n1357 vdd.n1356 52.4337
R3064 vdd.n1362 vdd.n1361 52.4337
R3065 vdd.n1365 vdd.n1364 52.4337
R3066 vdd.n1370 vdd.n1369 52.4337
R3067 vdd.n1373 vdd.n1372 52.4337
R3068 vdd.n1378 vdd.n1377 52.4337
R3069 vdd.n1381 vdd.n1380 52.4337
R3070 vdd.n1388 vdd.n1387 52.4337
R3071 vdd.n1391 vdd.n1390 52.4337
R3072 vdd.n1396 vdd.n1395 52.4337
R3073 vdd.n1399 vdd.n1398 52.4337
R3074 vdd.n1404 vdd.n1403 52.4337
R3075 vdd.n1407 vdd.n1406 52.4337
R3076 vdd.n1412 vdd.n1411 52.4337
R3077 vdd.n1415 vdd.n1414 52.4337
R3078 vdd.n1420 vdd.n1419 52.4337
R3079 vdd.n1423 vdd.n1422 52.4337
R3080 vdd.n1428 vdd.n1427 52.4337
R3081 vdd.n1508 vdd.n1507 52.4337
R3082 vdd.n1505 vdd.n1431 52.4337
R3083 vdd.n1437 vdd.n1436 52.4337
R3084 vdd.n1442 vdd.n1439 52.4337
R3085 vdd.n1445 vdd.n1444 52.4337
R3086 vdd.n1450 vdd.n1447 52.4337
R3087 vdd.n1453 vdd.n1452 52.4337
R3088 vdd.n1458 vdd.n1455 52.4337
R3089 vdd.n1461 vdd.n1460 52.4337
R3090 vdd.n1466 vdd.n1463 52.4337
R3091 vdd.n1469 vdd.n1468 52.4337
R3092 vdd.n1349 vdd.n1348 52.4337
R3093 vdd.n1355 vdd.n1354 52.4337
R3094 vdd.n1358 vdd.n1357 52.4337
R3095 vdd.n1363 vdd.n1362 52.4337
R3096 vdd.n1366 vdd.n1365 52.4337
R3097 vdd.n1371 vdd.n1370 52.4337
R3098 vdd.n1374 vdd.n1373 52.4337
R3099 vdd.n1379 vdd.n1378 52.4337
R3100 vdd.n1382 vdd.n1381 52.4337
R3101 vdd.n1389 vdd.n1388 52.4337
R3102 vdd.n1392 vdd.n1391 52.4337
R3103 vdd.n1397 vdd.n1396 52.4337
R3104 vdd.n1400 vdd.n1399 52.4337
R3105 vdd.n1405 vdd.n1404 52.4337
R3106 vdd.n1408 vdd.n1407 52.4337
R3107 vdd.n1413 vdd.n1412 52.4337
R3108 vdd.n1416 vdd.n1415 52.4337
R3109 vdd.n1421 vdd.n1420 52.4337
R3110 vdd.n1424 vdd.n1423 52.4337
R3111 vdd.n1429 vdd.n1428 52.4337
R3112 vdd.n1507 vdd.n1506 52.4337
R3113 vdd.n1435 vdd.n1431 52.4337
R3114 vdd.n1438 vdd.n1437 52.4337
R3115 vdd.n1443 vdd.n1442 52.4337
R3116 vdd.n1446 vdd.n1445 52.4337
R3117 vdd.n1451 vdd.n1450 52.4337
R3118 vdd.n1454 vdd.n1453 52.4337
R3119 vdd.n1459 vdd.n1458 52.4337
R3120 vdd.n1462 vdd.n1461 52.4337
R3121 vdd.n1467 vdd.n1466 52.4337
R3122 vdd.n1470 vdd.n1469 52.4337
R3123 vdd.n1261 vdd.n1260 52.4337
R3124 vdd.n1258 vdd.n1257 52.4337
R3125 vdd.n1254 vdd.n1046 52.4337
R3126 vdd.n1992 vdd.n1991 52.4337
R3127 vdd.n1045 vdd.n1039 52.4337
R3128 vdd.n1999 vdd.n1998 52.4337
R3129 vdd.n1038 vdd.n1032 52.4337
R3130 vdd.n2006 vdd.n2005 52.4337
R3131 vdd.n1031 vdd.n1026 52.4337
R3132 vdd.n2013 vdd.n2012 52.4337
R3133 vdd.n1025 vdd.n1024 52.4337
R3134 vdd.n1020 vdd.n1013 52.4337
R3135 vdd.n2024 vdd.n2023 52.4337
R3136 vdd.n1012 vdd.n1006 52.4337
R3137 vdd.n2031 vdd.n2030 52.4337
R3138 vdd.n1005 vdd.n999 52.4337
R3139 vdd.n2038 vdd.n2037 52.4337
R3140 vdd.n998 vdd.n992 52.4337
R3141 vdd.n2045 vdd.n2044 52.4337
R3142 vdd.n991 vdd.n986 52.4337
R3143 vdd.n2052 vdd.n2051 52.4337
R3144 vdd.n985 vdd.n984 52.4337
R3145 vdd.n980 vdd.n973 52.4337
R3146 vdd.n2063 vdd.n2062 52.4337
R3147 vdd.n972 vdd.n966 52.4337
R3148 vdd.n2070 vdd.n2069 52.4337
R3149 vdd.n965 vdd.n959 52.4337
R3150 vdd.n2077 vdd.n2076 52.4337
R3151 vdd.n958 vdd.n955 52.4337
R3152 vdd.n2084 vdd.n2083 52.4337
R3153 vdd.n2089 vdd.n2088 52.4337
R3154 vdd.n1265 vdd.n954 52.4337
R3155 vdd.n3025 vdd.n3024 52.4337
R3156 vdd.n3019 vdd.n520 52.4337
R3157 vdd.n3015 vdd.n523 52.4337
R3158 vdd.n3013 vdd.n3012 52.4337
R3159 vdd.n3008 vdd.n3007 52.4337
R3160 vdd.n3005 vdd.n3004 52.4337
R3161 vdd.n3000 vdd.n2999 52.4337
R3162 vdd.n2997 vdd.n2996 52.4337
R3163 vdd.n2992 vdd.n2991 52.4337
R3164 vdd.n2989 vdd.n2988 52.4337
R3165 vdd.n2984 vdd.n2983 52.4337
R3166 vdd.n2981 vdd.n2980 52.4337
R3167 vdd.n2976 vdd.n2975 52.4337
R3168 vdd.n2973 vdd.n2972 52.4337
R3169 vdd.n2968 vdd.n2967 52.4337
R3170 vdd.n2965 vdd.n2964 52.4337
R3171 vdd.n2960 vdd.n2959 52.4337
R3172 vdd.n2957 vdd.n2956 52.4337
R3173 vdd.n2952 vdd.n2951 52.4337
R3174 vdd.n2949 vdd.n2948 52.4337
R3175 vdd.n585 vdd.n584 52.4337
R3176 vdd.n2940 vdd.n2939 52.4337
R3177 vdd.n2935 vdd.n586 52.4337
R3178 vdd.n2933 vdd.n2932 52.4337
R3179 vdd.n2928 vdd.n2927 52.4337
R3180 vdd.n2925 vdd.n2924 52.4337
R3181 vdd.n2920 vdd.n2919 52.4337
R3182 vdd.n2917 vdd.n2916 52.4337
R3183 vdd.n2912 vdd.n2911 52.4337
R3184 vdd.n2907 vdd.n607 52.4337
R3185 vdd.n2903 vdd.n609 52.4337
R3186 vdd.n3110 vdd.n462 52.4337
R3187 vdd.n3120 vdd.n3119 52.4337
R3188 vdd.n461 vdd.n455 52.4337
R3189 vdd.n3127 vdd.n3126 52.4337
R3190 vdd.n454 vdd.n448 52.4337
R3191 vdd.n3134 vdd.n3133 52.4337
R3192 vdd.n447 vdd.n441 52.4337
R3193 vdd.n3141 vdd.n3140 52.4337
R3194 vdd.n440 vdd.n435 52.4337
R3195 vdd.n3148 vdd.n3147 52.4337
R3196 vdd.n434 vdd.n433 52.4337
R3197 vdd.n429 vdd.n422 52.4337
R3198 vdd.n3159 vdd.n3158 52.4337
R3199 vdd.n421 vdd.n415 52.4337
R3200 vdd.n3166 vdd.n3165 52.4337
R3201 vdd.n414 vdd.n408 52.4337
R3202 vdd.n3173 vdd.n3172 52.4337
R3203 vdd.n407 vdd.n401 52.4337
R3204 vdd.n3180 vdd.n3179 52.4337
R3205 vdd.n400 vdd.n395 52.4337
R3206 vdd.n3187 vdd.n3186 52.4337
R3207 vdd.n394 vdd.n393 52.4337
R3208 vdd.n389 vdd.n382 52.4337
R3209 vdd.n3198 vdd.n3197 52.4337
R3210 vdd.n381 vdd.n375 52.4337
R3211 vdd.n3205 vdd.n3204 52.4337
R3212 vdd.n374 vdd.n368 52.4337
R3213 vdd.n3212 vdd.n3211 52.4337
R3214 vdd.n367 vdd.n360 52.4337
R3215 vdd.n3219 vdd.n3218 52.4337
R3216 vdd.n3222 vdd.n3221 52.4337
R3217 vdd.n355 vdd.n352 52.4337
R3218 vdd.t29 vdd.t11 51.4683
R3219 vdd.n258 vdd.n256 42.0461
R3220 vdd.n164 vdd.n162 42.0461
R3221 vdd.n71 vdd.n69 42.0461
R3222 vdd.n1866 vdd.n1864 42.0461
R3223 vdd.n1772 vdd.n1770 42.0461
R3224 vdd.n1679 vdd.n1677 42.0461
R3225 vdd.n308 vdd.n307 41.6884
R3226 vdd.n214 vdd.n213 41.6884
R3227 vdd.n121 vdd.n120 41.6884
R3228 vdd.n1916 vdd.n1915 41.6884
R3229 vdd.n1822 vdd.n1821 41.6884
R3230 vdd.n1729 vdd.n1728 41.6884
R3231 vdd.n1474 vdd.n1473 41.1157
R3232 vdd.n1511 vdd.n1510 41.1157
R3233 vdd.n1385 vdd.n1384 41.1157
R3234 vdd.n3115 vdd.n3114 41.1157
R3235 vdd.n3154 vdd.n428 41.1157
R3236 vdd.n3193 vdd.n388 41.1157
R3237 vdd.n2857 vdd.n2856 39.2114
R3238 vdd.n2854 vdd.n2853 39.2114
R3239 vdd.n2849 vdd.n641 39.2114
R3240 vdd.n2847 vdd.n2846 39.2114
R3241 vdd.n2842 vdd.n644 39.2114
R3242 vdd.n2840 vdd.n2839 39.2114
R3243 vdd.n2835 vdd.n647 39.2114
R3244 vdd.n2833 vdd.n2832 39.2114
R3245 vdd.n2827 vdd.n650 39.2114
R3246 vdd.n2825 vdd.n2824 39.2114
R3247 vdd.n2820 vdd.n653 39.2114
R3248 vdd.n2818 vdd.n2817 39.2114
R3249 vdd.n2813 vdd.n656 39.2114
R3250 vdd.n2811 vdd.n2810 39.2114
R3251 vdd.n2806 vdd.n659 39.2114
R3252 vdd.n2804 vdd.n2803 39.2114
R3253 vdd.n2799 vdd.n2798 39.2114
R3254 vdd.n2649 vdd.n2648 39.2114
R3255 vdd.n2643 vdd.n2378 39.2114
R3256 vdd.n2640 vdd.n2379 39.2114
R3257 vdd.n2636 vdd.n2380 39.2114
R3258 vdd.n2632 vdd.n2381 39.2114
R3259 vdd.n2628 vdd.n2382 39.2114
R3260 vdd.n2624 vdd.n2383 39.2114
R3261 vdd.n2620 vdd.n2384 39.2114
R3262 vdd.n2616 vdd.n2385 39.2114
R3263 vdd.n2612 vdd.n2386 39.2114
R3264 vdd.n2608 vdd.n2387 39.2114
R3265 vdd.n2604 vdd.n2388 39.2114
R3266 vdd.n2600 vdd.n2389 39.2114
R3267 vdd.n2596 vdd.n2390 39.2114
R3268 vdd.n2592 vdd.n2391 39.2114
R3269 vdd.n2588 vdd.n2392 39.2114
R3270 vdd.n2583 vdd.n2393 39.2114
R3271 vdd.n2372 vdd.n796 39.2114
R3272 vdd.n2368 vdd.n795 39.2114
R3273 vdd.n2364 vdd.n794 39.2114
R3274 vdd.n2360 vdd.n793 39.2114
R3275 vdd.n2356 vdd.n792 39.2114
R3276 vdd.n2352 vdd.n791 39.2114
R3277 vdd.n2348 vdd.n790 39.2114
R3278 vdd.n2344 vdd.n789 39.2114
R3279 vdd.n2340 vdd.n788 39.2114
R3280 vdd.n2336 vdd.n787 39.2114
R3281 vdd.n2332 vdd.n786 39.2114
R3282 vdd.n2328 vdd.n785 39.2114
R3283 vdd.n2324 vdd.n784 39.2114
R3284 vdd.n2320 vdd.n783 39.2114
R3285 vdd.n2316 vdd.n782 39.2114
R3286 vdd.n2311 vdd.n781 39.2114
R3287 vdd.n2307 vdd.n780 39.2114
R3288 vdd.n2128 vdd.n2127 39.2114
R3289 vdd.n2122 vdd.n912 39.2114
R3290 vdd.n2119 vdd.n913 39.2114
R3291 vdd.n2115 vdd.n914 39.2114
R3292 vdd.n2111 vdd.n915 39.2114
R3293 vdd.n2107 vdd.n916 39.2114
R3294 vdd.n2103 vdd.n917 39.2114
R3295 vdd.n2099 vdd.n918 39.2114
R3296 vdd.n2095 vdd.n919 39.2114
R3297 vdd.n1104 vdd.n920 39.2114
R3298 vdd.n1108 vdd.n921 39.2114
R3299 vdd.n1112 vdd.n922 39.2114
R3300 vdd.n1116 vdd.n923 39.2114
R3301 vdd.n1120 vdd.n924 39.2114
R3302 vdd.n1124 vdd.n925 39.2114
R3303 vdd.n1128 vdd.n926 39.2114
R3304 vdd.n1133 vdd.n927 39.2114
R3305 vdd.n2776 vdd.n2775 39.2114
R3306 vdd.n2771 vdd.n2743 39.2114
R3307 vdd.n2769 vdd.n2768 39.2114
R3308 vdd.n2764 vdd.n2746 39.2114
R3309 vdd.n2762 vdd.n2761 39.2114
R3310 vdd.n2757 vdd.n2749 39.2114
R3311 vdd.n2755 vdd.n2754 39.2114
R3312 vdd.n2750 vdd.n612 39.2114
R3313 vdd.n2894 vdd.n2893 39.2114
R3314 vdd.n2891 vdd.n2890 39.2114
R3315 vdd.n2886 vdd.n617 39.2114
R3316 vdd.n2884 vdd.n2883 39.2114
R3317 vdd.n2879 vdd.n620 39.2114
R3318 vdd.n2877 vdd.n2876 39.2114
R3319 vdd.n2872 vdd.n623 39.2114
R3320 vdd.n2870 vdd.n2869 39.2114
R3321 vdd.n2865 vdd.n629 39.2114
R3322 vdd.n2652 vdd.n2651 39.2114
R3323 vdd.n2419 vdd.n2394 39.2114
R3324 vdd.n2423 vdd.n2395 39.2114
R3325 vdd.n2427 vdd.n2396 39.2114
R3326 vdd.n2431 vdd.n2397 39.2114
R3327 vdd.n2435 vdd.n2398 39.2114
R3328 vdd.n2439 vdd.n2399 39.2114
R3329 vdd.n2443 vdd.n2400 39.2114
R3330 vdd.n2447 vdd.n2401 39.2114
R3331 vdd.n2451 vdd.n2402 39.2114
R3332 vdd.n2455 vdd.n2403 39.2114
R3333 vdd.n2459 vdd.n2404 39.2114
R3334 vdd.n2463 vdd.n2405 39.2114
R3335 vdd.n2467 vdd.n2406 39.2114
R3336 vdd.n2471 vdd.n2407 39.2114
R3337 vdd.n2475 vdd.n2408 39.2114
R3338 vdd.n2479 vdd.n2409 39.2114
R3339 vdd.n2651 vdd.n761 39.2114
R3340 vdd.n2422 vdd.n2394 39.2114
R3341 vdd.n2426 vdd.n2395 39.2114
R3342 vdd.n2430 vdd.n2396 39.2114
R3343 vdd.n2434 vdd.n2397 39.2114
R3344 vdd.n2438 vdd.n2398 39.2114
R3345 vdd.n2442 vdd.n2399 39.2114
R3346 vdd.n2446 vdd.n2400 39.2114
R3347 vdd.n2450 vdd.n2401 39.2114
R3348 vdd.n2454 vdd.n2402 39.2114
R3349 vdd.n2458 vdd.n2403 39.2114
R3350 vdd.n2462 vdd.n2404 39.2114
R3351 vdd.n2466 vdd.n2405 39.2114
R3352 vdd.n2470 vdd.n2406 39.2114
R3353 vdd.n2474 vdd.n2407 39.2114
R3354 vdd.n2478 vdd.n2408 39.2114
R3355 vdd.n2481 vdd.n2409 39.2114
R3356 vdd.n629 vdd.n624 39.2114
R3357 vdd.n2871 vdd.n2870 39.2114
R3358 vdd.n623 vdd.n621 39.2114
R3359 vdd.n2878 vdd.n2877 39.2114
R3360 vdd.n620 vdd.n618 39.2114
R3361 vdd.n2885 vdd.n2884 39.2114
R3362 vdd.n617 vdd.n615 39.2114
R3363 vdd.n2892 vdd.n2891 39.2114
R3364 vdd.n2895 vdd.n2894 39.2114
R3365 vdd.n2751 vdd.n2750 39.2114
R3366 vdd.n2756 vdd.n2755 39.2114
R3367 vdd.n2749 vdd.n2747 39.2114
R3368 vdd.n2763 vdd.n2762 39.2114
R3369 vdd.n2746 vdd.n2744 39.2114
R3370 vdd.n2770 vdd.n2769 39.2114
R3371 vdd.n2743 vdd.n2741 39.2114
R3372 vdd.n2777 vdd.n2776 39.2114
R3373 vdd.n2128 vdd.n946 39.2114
R3374 vdd.n2120 vdd.n912 39.2114
R3375 vdd.n2116 vdd.n913 39.2114
R3376 vdd.n2112 vdd.n914 39.2114
R3377 vdd.n2108 vdd.n915 39.2114
R3378 vdd.n2104 vdd.n916 39.2114
R3379 vdd.n2100 vdd.n917 39.2114
R3380 vdd.n2096 vdd.n918 39.2114
R3381 vdd.n1103 vdd.n919 39.2114
R3382 vdd.n1107 vdd.n920 39.2114
R3383 vdd.n1111 vdd.n921 39.2114
R3384 vdd.n1115 vdd.n922 39.2114
R3385 vdd.n1119 vdd.n923 39.2114
R3386 vdd.n1123 vdd.n924 39.2114
R3387 vdd.n1127 vdd.n925 39.2114
R3388 vdd.n1132 vdd.n926 39.2114
R3389 vdd.n1136 vdd.n927 39.2114
R3390 vdd.n2310 vdd.n780 39.2114
R3391 vdd.n2315 vdd.n781 39.2114
R3392 vdd.n2319 vdd.n782 39.2114
R3393 vdd.n2323 vdd.n783 39.2114
R3394 vdd.n2327 vdd.n784 39.2114
R3395 vdd.n2331 vdd.n785 39.2114
R3396 vdd.n2335 vdd.n786 39.2114
R3397 vdd.n2339 vdd.n787 39.2114
R3398 vdd.n2343 vdd.n788 39.2114
R3399 vdd.n2347 vdd.n789 39.2114
R3400 vdd.n2351 vdd.n790 39.2114
R3401 vdd.n2355 vdd.n791 39.2114
R3402 vdd.n2359 vdd.n792 39.2114
R3403 vdd.n2363 vdd.n793 39.2114
R3404 vdd.n2367 vdd.n794 39.2114
R3405 vdd.n2371 vdd.n795 39.2114
R3406 vdd.n798 vdd.n796 39.2114
R3407 vdd.n2649 vdd.n2412 39.2114
R3408 vdd.n2641 vdd.n2378 39.2114
R3409 vdd.n2637 vdd.n2379 39.2114
R3410 vdd.n2633 vdd.n2380 39.2114
R3411 vdd.n2629 vdd.n2381 39.2114
R3412 vdd.n2625 vdd.n2382 39.2114
R3413 vdd.n2621 vdd.n2383 39.2114
R3414 vdd.n2617 vdd.n2384 39.2114
R3415 vdd.n2613 vdd.n2385 39.2114
R3416 vdd.n2609 vdd.n2386 39.2114
R3417 vdd.n2605 vdd.n2387 39.2114
R3418 vdd.n2601 vdd.n2388 39.2114
R3419 vdd.n2597 vdd.n2389 39.2114
R3420 vdd.n2593 vdd.n2390 39.2114
R3421 vdd.n2589 vdd.n2391 39.2114
R3422 vdd.n2584 vdd.n2392 39.2114
R3423 vdd.n2580 vdd.n2393 39.2114
R3424 vdd.n2798 vdd.n660 39.2114
R3425 vdd.n2805 vdd.n2804 39.2114
R3426 vdd.n659 vdd.n657 39.2114
R3427 vdd.n2812 vdd.n2811 39.2114
R3428 vdd.n656 vdd.n654 39.2114
R3429 vdd.n2819 vdd.n2818 39.2114
R3430 vdd.n653 vdd.n651 39.2114
R3431 vdd.n2826 vdd.n2825 39.2114
R3432 vdd.n650 vdd.n648 39.2114
R3433 vdd.n2834 vdd.n2833 39.2114
R3434 vdd.n647 vdd.n645 39.2114
R3435 vdd.n2841 vdd.n2840 39.2114
R3436 vdd.n644 vdd.n642 39.2114
R3437 vdd.n2848 vdd.n2847 39.2114
R3438 vdd.n641 vdd.n639 39.2114
R3439 vdd.n2855 vdd.n2854 39.2114
R3440 vdd.n2858 vdd.n2857 39.2114
R3441 vdd.n807 vdd.n762 39.2114
R3442 vdd.n2299 vdd.n763 39.2114
R3443 vdd.n2295 vdd.n764 39.2114
R3444 vdd.n2291 vdd.n765 39.2114
R3445 vdd.n2287 vdd.n766 39.2114
R3446 vdd.n2283 vdd.n767 39.2114
R3447 vdd.n2279 vdd.n768 39.2114
R3448 vdd.n2275 vdd.n769 39.2114
R3449 vdd.n2271 vdd.n770 39.2114
R3450 vdd.n2267 vdd.n771 39.2114
R3451 vdd.n2263 vdd.n772 39.2114
R3452 vdd.n2259 vdd.n773 39.2114
R3453 vdd.n2255 vdd.n774 39.2114
R3454 vdd.n2251 vdd.n775 39.2114
R3455 vdd.n2247 vdd.n776 39.2114
R3456 vdd.n2243 vdd.n777 39.2114
R3457 vdd.n2239 vdd.n778 39.2114
R3458 vdd.n2131 vdd.n2130 39.2114
R3459 vdd.n1050 vdd.n928 39.2114
R3460 vdd.n1054 vdd.n929 39.2114
R3461 vdd.n1058 vdd.n930 39.2114
R3462 vdd.n1062 vdd.n931 39.2114
R3463 vdd.n1066 vdd.n932 39.2114
R3464 vdd.n1070 vdd.n933 39.2114
R3465 vdd.n1074 vdd.n934 39.2114
R3466 vdd.n1078 vdd.n935 39.2114
R3467 vdd.n1248 vdd.n936 39.2114
R3468 vdd.n1245 vdd.n937 39.2114
R3469 vdd.n1241 vdd.n938 39.2114
R3470 vdd.n1237 vdd.n939 39.2114
R3471 vdd.n1233 vdd.n940 39.2114
R3472 vdd.n1229 vdd.n941 39.2114
R3473 vdd.n1225 vdd.n942 39.2114
R3474 vdd.n1221 vdd.n943 39.2114
R3475 vdd.n2236 vdd.n778 39.2114
R3476 vdd.n2240 vdd.n777 39.2114
R3477 vdd.n2244 vdd.n776 39.2114
R3478 vdd.n2248 vdd.n775 39.2114
R3479 vdd.n2252 vdd.n774 39.2114
R3480 vdd.n2256 vdd.n773 39.2114
R3481 vdd.n2260 vdd.n772 39.2114
R3482 vdd.n2264 vdd.n771 39.2114
R3483 vdd.n2268 vdd.n770 39.2114
R3484 vdd.n2272 vdd.n769 39.2114
R3485 vdd.n2276 vdd.n768 39.2114
R3486 vdd.n2280 vdd.n767 39.2114
R3487 vdd.n2284 vdd.n766 39.2114
R3488 vdd.n2288 vdd.n765 39.2114
R3489 vdd.n2292 vdd.n764 39.2114
R3490 vdd.n2296 vdd.n763 39.2114
R3491 vdd.n2300 vdd.n762 39.2114
R3492 vdd.n2130 vdd.n910 39.2114
R3493 vdd.n1053 vdd.n928 39.2114
R3494 vdd.n1057 vdd.n929 39.2114
R3495 vdd.n1061 vdd.n930 39.2114
R3496 vdd.n1065 vdd.n931 39.2114
R3497 vdd.n1069 vdd.n932 39.2114
R3498 vdd.n1073 vdd.n933 39.2114
R3499 vdd.n1077 vdd.n934 39.2114
R3500 vdd.n1080 vdd.n935 39.2114
R3501 vdd.n1246 vdd.n936 39.2114
R3502 vdd.n1242 vdd.n937 39.2114
R3503 vdd.n1238 vdd.n938 39.2114
R3504 vdd.n1234 vdd.n939 39.2114
R3505 vdd.n1230 vdd.n940 39.2114
R3506 vdd.n1226 vdd.n941 39.2114
R3507 vdd.n1222 vdd.n942 39.2114
R3508 vdd.n1218 vdd.n943 39.2114
R3509 vdd.n1983 vdd.n1982 37.2369
R3510 vdd.n2019 vdd.n1019 37.2369
R3511 vdd.n2058 vdd.n979 37.2369
R3512 vdd.n2946 vdd.n581 37.2369
R3513 vdd.n545 vdd.n544 37.2369
R3514 vdd.n2902 vdd.n2901 37.2369
R3515 vdd.n2126 vdd.n902 31.0639
R3516 vdd.n2375 vdd.n799 31.0639
R3517 vdd.n2308 vdd.n802 31.0639
R3518 vdd.n1138 vdd.n1135 31.0639
R3519 vdd.n2581 vdd.n2578 31.0639
R3520 vdd.n2800 vdd.n2797 31.0639
R3521 vdd.n2647 vdd.n754 31.0639
R3522 vdd.n2861 vdd.n2860 31.0639
R3523 vdd.n2780 vdd.n2779 31.0639
R3524 vdd.n2866 vdd.n628 31.0639
R3525 vdd.n2485 vdd.n2483 31.0639
R3526 vdd.n2654 vdd.n2653 31.0639
R3527 vdd.n2133 vdd.n2132 31.0639
R3528 vdd.n2303 vdd.n2302 31.0639
R3529 vdd.n2235 vdd.n2234 31.0639
R3530 vdd.n1217 vdd.n1216 31.0639
R3531 vdd.n1083 vdd.n1082 30.449
R3532 vdd.n811 vdd.n810 30.449
R3533 vdd.n1130 vdd.n1102 30.449
R3534 vdd.n2313 vdd.n801 30.449
R3535 vdd.n2418 vdd.n2417 30.449
R3536 vdd.n663 vdd.n662 30.449
R3537 vdd.n2586 vdd.n2414 30.449
R3538 vdd.n627 vdd.n626 30.449
R3539 vdd.n1577 vdd.n1344 20.633
R3540 vdd.n1977 vdd.n911 20.633
R3541 vdd.n3032 vdd.n516 20.633
R3542 vdd.n3230 vdd.n351 20.633
R3543 vdd.n1579 vdd.n1341 19.3944
R3544 vdd.n1583 vdd.n1341 19.3944
R3545 vdd.n1583 vdd.n1332 19.3944
R3546 vdd.n1595 vdd.n1332 19.3944
R3547 vdd.n1595 vdd.n1330 19.3944
R3548 vdd.n1599 vdd.n1330 19.3944
R3549 vdd.n1599 vdd.n1319 19.3944
R3550 vdd.n1611 vdd.n1319 19.3944
R3551 vdd.n1611 vdd.n1317 19.3944
R3552 vdd.n1615 vdd.n1317 19.3944
R3553 vdd.n1615 vdd.n1308 19.3944
R3554 vdd.n1628 vdd.n1308 19.3944
R3555 vdd.n1628 vdd.n1306 19.3944
R3556 vdd.n1632 vdd.n1306 19.3944
R3557 vdd.n1632 vdd.n1297 19.3944
R3558 vdd.n1926 vdd.n1297 19.3944
R3559 vdd.n1926 vdd.n1295 19.3944
R3560 vdd.n1930 vdd.n1295 19.3944
R3561 vdd.n1930 vdd.n1285 19.3944
R3562 vdd.n1943 vdd.n1285 19.3944
R3563 vdd.n1943 vdd.n1283 19.3944
R3564 vdd.n1947 vdd.n1283 19.3944
R3565 vdd.n1947 vdd.n1275 19.3944
R3566 vdd.n1960 vdd.n1275 19.3944
R3567 vdd.n1960 vdd.n1272 19.3944
R3568 vdd.n1966 vdd.n1272 19.3944
R3569 vdd.n1966 vdd.n1273 19.3944
R3570 vdd.n1273 vdd.n1263 19.3944
R3571 vdd.n1504 vdd.n1430 19.3944
R3572 vdd.n1504 vdd.n1432 19.3944
R3573 vdd.n1500 vdd.n1432 19.3944
R3574 vdd.n1500 vdd.n1499 19.3944
R3575 vdd.n1499 vdd.n1498 19.3944
R3576 vdd.n1498 vdd.n1440 19.3944
R3577 vdd.n1494 vdd.n1440 19.3944
R3578 vdd.n1494 vdd.n1493 19.3944
R3579 vdd.n1493 vdd.n1492 19.3944
R3580 vdd.n1492 vdd.n1448 19.3944
R3581 vdd.n1488 vdd.n1448 19.3944
R3582 vdd.n1488 vdd.n1487 19.3944
R3583 vdd.n1487 vdd.n1486 19.3944
R3584 vdd.n1486 vdd.n1456 19.3944
R3585 vdd.n1482 vdd.n1456 19.3944
R3586 vdd.n1482 vdd.n1481 19.3944
R3587 vdd.n1481 vdd.n1480 19.3944
R3588 vdd.n1480 vdd.n1464 19.3944
R3589 vdd.n1476 vdd.n1464 19.3944
R3590 vdd.n1476 vdd.n1475 19.3944
R3591 vdd.n1542 vdd.n1541 19.3944
R3592 vdd.n1541 vdd.n1540 19.3944
R3593 vdd.n1540 vdd.n1393 19.3944
R3594 vdd.n1536 vdd.n1393 19.3944
R3595 vdd.n1536 vdd.n1535 19.3944
R3596 vdd.n1535 vdd.n1534 19.3944
R3597 vdd.n1534 vdd.n1401 19.3944
R3598 vdd.n1530 vdd.n1401 19.3944
R3599 vdd.n1530 vdd.n1529 19.3944
R3600 vdd.n1529 vdd.n1528 19.3944
R3601 vdd.n1528 vdd.n1409 19.3944
R3602 vdd.n1524 vdd.n1409 19.3944
R3603 vdd.n1524 vdd.n1523 19.3944
R3604 vdd.n1523 vdd.n1522 19.3944
R3605 vdd.n1522 vdd.n1417 19.3944
R3606 vdd.n1518 vdd.n1417 19.3944
R3607 vdd.n1518 vdd.n1517 19.3944
R3608 vdd.n1517 vdd.n1516 19.3944
R3609 vdd.n1516 vdd.n1425 19.3944
R3610 vdd.n1512 vdd.n1425 19.3944
R3611 vdd.n1572 vdd.n1571 19.3944
R3612 vdd.n1571 vdd.n1570 19.3944
R3613 vdd.n1570 vdd.n1351 19.3944
R3614 vdd.n1566 vdd.n1351 19.3944
R3615 vdd.n1566 vdd.n1565 19.3944
R3616 vdd.n1565 vdd.n1564 19.3944
R3617 vdd.n1564 vdd.n1359 19.3944
R3618 vdd.n1560 vdd.n1359 19.3944
R3619 vdd.n1560 vdd.n1559 19.3944
R3620 vdd.n1559 vdd.n1558 19.3944
R3621 vdd.n1558 vdd.n1367 19.3944
R3622 vdd.n1554 vdd.n1367 19.3944
R3623 vdd.n1554 vdd.n1553 19.3944
R3624 vdd.n1553 vdd.n1552 19.3944
R3625 vdd.n1552 vdd.n1375 19.3944
R3626 vdd.n1548 vdd.n1375 19.3944
R3627 vdd.n1548 vdd.n1547 19.3944
R3628 vdd.n1547 vdd.n1546 19.3944
R3629 vdd.n2015 vdd.n1017 19.3944
R3630 vdd.n2015 vdd.n1023 19.3944
R3631 vdd.n2010 vdd.n1023 19.3944
R3632 vdd.n2010 vdd.n2009 19.3944
R3633 vdd.n2009 vdd.n2008 19.3944
R3634 vdd.n2008 vdd.n1030 19.3944
R3635 vdd.n2003 vdd.n1030 19.3944
R3636 vdd.n2003 vdd.n2002 19.3944
R3637 vdd.n2002 vdd.n2001 19.3944
R3638 vdd.n2001 vdd.n1037 19.3944
R3639 vdd.n1996 vdd.n1037 19.3944
R3640 vdd.n1996 vdd.n1995 19.3944
R3641 vdd.n1995 vdd.n1994 19.3944
R3642 vdd.n1994 vdd.n1044 19.3944
R3643 vdd.n1989 vdd.n1044 19.3944
R3644 vdd.n1989 vdd.n1988 19.3944
R3645 vdd.n1256 vdd.n1049 19.3944
R3646 vdd.n1984 vdd.n1253 19.3944
R3647 vdd.n2054 vdd.n977 19.3944
R3648 vdd.n2054 vdd.n983 19.3944
R3649 vdd.n2049 vdd.n983 19.3944
R3650 vdd.n2049 vdd.n2048 19.3944
R3651 vdd.n2048 vdd.n2047 19.3944
R3652 vdd.n2047 vdd.n990 19.3944
R3653 vdd.n2042 vdd.n990 19.3944
R3654 vdd.n2042 vdd.n2041 19.3944
R3655 vdd.n2041 vdd.n2040 19.3944
R3656 vdd.n2040 vdd.n997 19.3944
R3657 vdd.n2035 vdd.n997 19.3944
R3658 vdd.n2035 vdd.n2034 19.3944
R3659 vdd.n2034 vdd.n2033 19.3944
R3660 vdd.n2033 vdd.n1004 19.3944
R3661 vdd.n2028 vdd.n1004 19.3944
R3662 vdd.n2028 vdd.n2027 19.3944
R3663 vdd.n2027 vdd.n2026 19.3944
R3664 vdd.n2026 vdd.n1011 19.3944
R3665 vdd.n2021 vdd.n1011 19.3944
R3666 vdd.n2021 vdd.n2020 19.3944
R3667 vdd.n2091 vdd.n952 19.3944
R3668 vdd.n2091 vdd.n953 19.3944
R3669 vdd.n2086 vdd.n2085 19.3944
R3670 vdd.n2081 vdd.n2080 19.3944
R3671 vdd.n2080 vdd.n2079 19.3944
R3672 vdd.n2079 vdd.n957 19.3944
R3673 vdd.n2074 vdd.n957 19.3944
R3674 vdd.n2074 vdd.n2073 19.3944
R3675 vdd.n2073 vdd.n2072 19.3944
R3676 vdd.n2072 vdd.n964 19.3944
R3677 vdd.n2067 vdd.n964 19.3944
R3678 vdd.n2067 vdd.n2066 19.3944
R3679 vdd.n2066 vdd.n2065 19.3944
R3680 vdd.n2065 vdd.n971 19.3944
R3681 vdd.n2060 vdd.n971 19.3944
R3682 vdd.n2060 vdd.n2059 19.3944
R3683 vdd.n1575 vdd.n1338 19.3944
R3684 vdd.n1587 vdd.n1338 19.3944
R3685 vdd.n1587 vdd.n1336 19.3944
R3686 vdd.n1591 vdd.n1336 19.3944
R3687 vdd.n1591 vdd.n1326 19.3944
R3688 vdd.n1603 vdd.n1326 19.3944
R3689 vdd.n1603 vdd.n1324 19.3944
R3690 vdd.n1607 vdd.n1324 19.3944
R3691 vdd.n1607 vdd.n1314 19.3944
R3692 vdd.n1620 vdd.n1314 19.3944
R3693 vdd.n1620 vdd.n1312 19.3944
R3694 vdd.n1624 vdd.n1312 19.3944
R3695 vdd.n1624 vdd.n1303 19.3944
R3696 vdd.n1636 vdd.n1303 19.3944
R3697 vdd.n1636 vdd.n1301 19.3944
R3698 vdd.n1922 vdd.n1301 19.3944
R3699 vdd.n1922 vdd.n1291 19.3944
R3700 vdd.n1935 vdd.n1291 19.3944
R3701 vdd.n1935 vdd.n1289 19.3944
R3702 vdd.n1939 vdd.n1289 19.3944
R3703 vdd.n1939 vdd.n1280 19.3944
R3704 vdd.n1952 vdd.n1280 19.3944
R3705 vdd.n1952 vdd.n1278 19.3944
R3706 vdd.n1956 vdd.n1278 19.3944
R3707 vdd.n1956 vdd.n1268 19.3944
R3708 vdd.n1971 vdd.n1268 19.3944
R3709 vdd.n1971 vdd.n1266 19.3944
R3710 vdd.n1975 vdd.n1266 19.3944
R3711 vdd.n3034 vdd.n513 19.3944
R3712 vdd.n3038 vdd.n513 19.3944
R3713 vdd.n3038 vdd.n503 19.3944
R3714 vdd.n3050 vdd.n503 19.3944
R3715 vdd.n3050 vdd.n501 19.3944
R3716 vdd.n3054 vdd.n501 19.3944
R3717 vdd.n3054 vdd.n490 19.3944
R3718 vdd.n3066 vdd.n490 19.3944
R3719 vdd.n3066 vdd.n488 19.3944
R3720 vdd.n3070 vdd.n488 19.3944
R3721 vdd.n3070 vdd.n478 19.3944
R3722 vdd.n3083 vdd.n478 19.3944
R3723 vdd.n3083 vdd.n476 19.3944
R3724 vdd.n3087 vdd.n476 19.3944
R3725 vdd.n3088 vdd.n3087 19.3944
R3726 vdd.n3089 vdd.n3088 19.3944
R3727 vdd.n3089 vdd.n474 19.3944
R3728 vdd.n3093 vdd.n474 19.3944
R3729 vdd.n3094 vdd.n3093 19.3944
R3730 vdd.n3095 vdd.n3094 19.3944
R3731 vdd.n3095 vdd.n471 19.3944
R3732 vdd.n3099 vdd.n471 19.3944
R3733 vdd.n3100 vdd.n3099 19.3944
R3734 vdd.n3101 vdd.n3100 19.3944
R3735 vdd.n3101 vdd.n468 19.3944
R3736 vdd.n3105 vdd.n468 19.3944
R3737 vdd.n3106 vdd.n3105 19.3944
R3738 vdd.n3107 vdd.n3106 19.3944
R3739 vdd.n3150 vdd.n426 19.3944
R3740 vdd.n3150 vdd.n432 19.3944
R3741 vdd.n3145 vdd.n432 19.3944
R3742 vdd.n3145 vdd.n3144 19.3944
R3743 vdd.n3144 vdd.n3143 19.3944
R3744 vdd.n3143 vdd.n439 19.3944
R3745 vdd.n3138 vdd.n439 19.3944
R3746 vdd.n3138 vdd.n3137 19.3944
R3747 vdd.n3137 vdd.n3136 19.3944
R3748 vdd.n3136 vdd.n446 19.3944
R3749 vdd.n3131 vdd.n446 19.3944
R3750 vdd.n3131 vdd.n3130 19.3944
R3751 vdd.n3130 vdd.n3129 19.3944
R3752 vdd.n3129 vdd.n453 19.3944
R3753 vdd.n3124 vdd.n453 19.3944
R3754 vdd.n3124 vdd.n3123 19.3944
R3755 vdd.n3123 vdd.n3122 19.3944
R3756 vdd.n3122 vdd.n460 19.3944
R3757 vdd.n3117 vdd.n460 19.3944
R3758 vdd.n3117 vdd.n3116 19.3944
R3759 vdd.n3189 vdd.n386 19.3944
R3760 vdd.n3189 vdd.n392 19.3944
R3761 vdd.n3184 vdd.n392 19.3944
R3762 vdd.n3184 vdd.n3183 19.3944
R3763 vdd.n3183 vdd.n3182 19.3944
R3764 vdd.n3182 vdd.n399 19.3944
R3765 vdd.n3177 vdd.n399 19.3944
R3766 vdd.n3177 vdd.n3176 19.3944
R3767 vdd.n3176 vdd.n3175 19.3944
R3768 vdd.n3175 vdd.n406 19.3944
R3769 vdd.n3170 vdd.n406 19.3944
R3770 vdd.n3170 vdd.n3169 19.3944
R3771 vdd.n3169 vdd.n3168 19.3944
R3772 vdd.n3168 vdd.n413 19.3944
R3773 vdd.n3163 vdd.n413 19.3944
R3774 vdd.n3163 vdd.n3162 19.3944
R3775 vdd.n3162 vdd.n3161 19.3944
R3776 vdd.n3161 vdd.n420 19.3944
R3777 vdd.n3156 vdd.n420 19.3944
R3778 vdd.n3156 vdd.n3155 19.3944
R3779 vdd.n3225 vdd.n3224 19.3944
R3780 vdd.n3224 vdd.n3223 19.3944
R3781 vdd.n3223 vdd.n358 19.3944
R3782 vdd.n359 vdd.n358 19.3944
R3783 vdd.n3216 vdd.n359 19.3944
R3784 vdd.n3216 vdd.n3215 19.3944
R3785 vdd.n3215 vdd.n3214 19.3944
R3786 vdd.n3214 vdd.n366 19.3944
R3787 vdd.n3209 vdd.n366 19.3944
R3788 vdd.n3209 vdd.n3208 19.3944
R3789 vdd.n3208 vdd.n3207 19.3944
R3790 vdd.n3207 vdd.n373 19.3944
R3791 vdd.n3202 vdd.n373 19.3944
R3792 vdd.n3202 vdd.n3201 19.3944
R3793 vdd.n3201 vdd.n3200 19.3944
R3794 vdd.n3200 vdd.n380 19.3944
R3795 vdd.n3195 vdd.n380 19.3944
R3796 vdd.n3195 vdd.n3194 19.3944
R3797 vdd.n3030 vdd.n509 19.3944
R3798 vdd.n3042 vdd.n509 19.3944
R3799 vdd.n3042 vdd.n507 19.3944
R3800 vdd.n3046 vdd.n507 19.3944
R3801 vdd.n3046 vdd.n497 19.3944
R3802 vdd.n3058 vdd.n497 19.3944
R3803 vdd.n3058 vdd.n495 19.3944
R3804 vdd.n3062 vdd.n495 19.3944
R3805 vdd.n3062 vdd.n485 19.3944
R3806 vdd.n3075 vdd.n485 19.3944
R3807 vdd.n3075 vdd.n483 19.3944
R3808 vdd.n3079 vdd.n483 19.3944
R3809 vdd.n3079 vdd.n312 19.3944
R3810 vdd.n3258 vdd.n312 19.3944
R3811 vdd.n3258 vdd.n313 19.3944
R3812 vdd.n3252 vdd.n313 19.3944
R3813 vdd.n3252 vdd.n3251 19.3944
R3814 vdd.n3251 vdd.n3250 19.3944
R3815 vdd.n3250 vdd.n323 19.3944
R3816 vdd.n3244 vdd.n323 19.3944
R3817 vdd.n3244 vdd.n3243 19.3944
R3818 vdd.n3243 vdd.n3242 19.3944
R3819 vdd.n3242 vdd.n335 19.3944
R3820 vdd.n3236 vdd.n335 19.3944
R3821 vdd.n3236 vdd.n3235 19.3944
R3822 vdd.n3235 vdd.n3234 19.3944
R3823 vdd.n3234 vdd.n346 19.3944
R3824 vdd.n3228 vdd.n346 19.3944
R3825 vdd.n2987 vdd.n2986 19.3944
R3826 vdd.n2986 vdd.n2985 19.3944
R3827 vdd.n2985 vdd.n551 19.3944
R3828 vdd.n2979 vdd.n551 19.3944
R3829 vdd.n2979 vdd.n2978 19.3944
R3830 vdd.n2978 vdd.n2977 19.3944
R3831 vdd.n2977 vdd.n557 19.3944
R3832 vdd.n2971 vdd.n557 19.3944
R3833 vdd.n2971 vdd.n2970 19.3944
R3834 vdd.n2970 vdd.n2969 19.3944
R3835 vdd.n2969 vdd.n563 19.3944
R3836 vdd.n2963 vdd.n563 19.3944
R3837 vdd.n2963 vdd.n2962 19.3944
R3838 vdd.n2962 vdd.n2961 19.3944
R3839 vdd.n2961 vdd.n569 19.3944
R3840 vdd.n2955 vdd.n569 19.3944
R3841 vdd.n2955 vdd.n2954 19.3944
R3842 vdd.n2954 vdd.n2953 19.3944
R3843 vdd.n2953 vdd.n575 19.3944
R3844 vdd.n2947 vdd.n575 19.3944
R3845 vdd.n3027 vdd.n3026 19.3944
R3846 vdd.n3026 vdd.n519 19.3944
R3847 vdd.n3021 vdd.n3020 19.3944
R3848 vdd.n3017 vdd.n3016 19.3944
R3849 vdd.n3016 vdd.n525 19.3944
R3850 vdd.n3011 vdd.n525 19.3944
R3851 vdd.n3011 vdd.n3010 19.3944
R3852 vdd.n3010 vdd.n3009 19.3944
R3853 vdd.n3009 vdd.n531 19.3944
R3854 vdd.n3003 vdd.n531 19.3944
R3855 vdd.n3003 vdd.n3002 19.3944
R3856 vdd.n3002 vdd.n3001 19.3944
R3857 vdd.n3001 vdd.n537 19.3944
R3858 vdd.n2995 vdd.n537 19.3944
R3859 vdd.n2995 vdd.n2994 19.3944
R3860 vdd.n2994 vdd.n2993 19.3944
R3861 vdd.n2942 vdd.n579 19.3944
R3862 vdd.n2942 vdd.n583 19.3944
R3863 vdd.n2937 vdd.n583 19.3944
R3864 vdd.n2937 vdd.n2936 19.3944
R3865 vdd.n2936 vdd.n589 19.3944
R3866 vdd.n2931 vdd.n589 19.3944
R3867 vdd.n2931 vdd.n2930 19.3944
R3868 vdd.n2930 vdd.n2929 19.3944
R3869 vdd.n2929 vdd.n595 19.3944
R3870 vdd.n2923 vdd.n595 19.3944
R3871 vdd.n2923 vdd.n2922 19.3944
R3872 vdd.n2922 vdd.n2921 19.3944
R3873 vdd.n2921 vdd.n601 19.3944
R3874 vdd.n2915 vdd.n601 19.3944
R3875 vdd.n2915 vdd.n2914 19.3944
R3876 vdd.n2914 vdd.n2913 19.3944
R3877 vdd.n2909 vdd.n2908 19.3944
R3878 vdd.n2905 vdd.n2904 19.3944
R3879 vdd.n1511 vdd.n1430 19.0066
R3880 vdd.n2019 vdd.n1017 19.0066
R3881 vdd.n3154 vdd.n426 19.0066
R3882 vdd.n2946 vdd.n579 19.0066
R3883 vdd.n1082 vdd.n1081 16.0975
R3884 vdd.n810 vdd.n809 16.0975
R3885 vdd.n1473 vdd.n1472 16.0975
R3886 vdd.n1510 vdd.n1509 16.0975
R3887 vdd.n1384 vdd.n1383 16.0975
R3888 vdd.n1982 vdd.n1981 16.0975
R3889 vdd.n1019 vdd.n1018 16.0975
R3890 vdd.n979 vdd.n978 16.0975
R3891 vdd.n1102 vdd.n1101 16.0975
R3892 vdd.n801 vdd.n800 16.0975
R3893 vdd.n2417 vdd.n2416 16.0975
R3894 vdd.n3114 vdd.n3113 16.0975
R3895 vdd.n428 vdd.n427 16.0975
R3896 vdd.n388 vdd.n387 16.0975
R3897 vdd.n581 vdd.n580 16.0975
R3898 vdd.n544 vdd.n543 16.0975
R3899 vdd.n662 vdd.n661 16.0975
R3900 vdd.n2414 vdd.n2413 16.0975
R3901 vdd.n2901 vdd.n2900 16.0975
R3902 vdd.n626 vdd.n625 16.0975
R3903 vdd.t11 vdd.n2377 15.4182
R3904 vdd.n2650 vdd.t29 15.4182
R3905 vdd.n28 vdd.n27 14.7341
R3906 vdd.n2129 vdd.n904 14.0578
R3907 vdd.n2863 vdd.n613 14.0578
R3908 vdd.n304 vdd.n269 13.1884
R3909 vdd.n253 vdd.n218 13.1884
R3910 vdd.n210 vdd.n175 13.1884
R3911 vdd.n159 vdd.n124 13.1884
R3912 vdd.n117 vdd.n82 13.1884
R3913 vdd.n66 vdd.n31 13.1884
R3914 vdd.n1861 vdd.n1826 13.1884
R3915 vdd.n1912 vdd.n1877 13.1884
R3916 vdd.n1767 vdd.n1732 13.1884
R3917 vdd.n1818 vdd.n1783 13.1884
R3918 vdd.n1674 vdd.n1639 13.1884
R3919 vdd.n1725 vdd.n1690 13.1884
R3920 vdd.n1542 vdd.n1385 12.9944
R3921 vdd.n1546 vdd.n1385 12.9944
R3922 vdd.n2058 vdd.n977 12.9944
R3923 vdd.n2059 vdd.n2058 12.9944
R3924 vdd.n3193 vdd.n386 12.9944
R3925 vdd.n3194 vdd.n3193 12.9944
R3926 vdd.n2987 vdd.n545 12.9944
R3927 vdd.n2993 vdd.n545 12.9944
R3928 vdd.n305 vdd.n267 12.8005
R3929 vdd.n300 vdd.n271 12.8005
R3930 vdd.n254 vdd.n216 12.8005
R3931 vdd.n249 vdd.n220 12.8005
R3932 vdd.n211 vdd.n173 12.8005
R3933 vdd.n206 vdd.n177 12.8005
R3934 vdd.n160 vdd.n122 12.8005
R3935 vdd.n155 vdd.n126 12.8005
R3936 vdd.n118 vdd.n80 12.8005
R3937 vdd.n113 vdd.n84 12.8005
R3938 vdd.n67 vdd.n29 12.8005
R3939 vdd.n62 vdd.n33 12.8005
R3940 vdd.n1862 vdd.n1824 12.8005
R3941 vdd.n1857 vdd.n1828 12.8005
R3942 vdd.n1913 vdd.n1875 12.8005
R3943 vdd.n1908 vdd.n1879 12.8005
R3944 vdd.n1768 vdd.n1730 12.8005
R3945 vdd.n1763 vdd.n1734 12.8005
R3946 vdd.n1819 vdd.n1781 12.8005
R3947 vdd.n1814 vdd.n1785 12.8005
R3948 vdd.n1675 vdd.n1637 12.8005
R3949 vdd.n1670 vdd.n1641 12.8005
R3950 vdd.n1726 vdd.n1688 12.8005
R3951 vdd.n1721 vdd.n1692 12.8005
R3952 vdd.n299 vdd.n272 12.0247
R3953 vdd.n248 vdd.n221 12.0247
R3954 vdd.n205 vdd.n178 12.0247
R3955 vdd.n154 vdd.n127 12.0247
R3956 vdd.n112 vdd.n85 12.0247
R3957 vdd.n61 vdd.n34 12.0247
R3958 vdd.n1856 vdd.n1829 12.0247
R3959 vdd.n1907 vdd.n1880 12.0247
R3960 vdd.n1762 vdd.n1735 12.0247
R3961 vdd.n1813 vdd.n1786 12.0247
R3962 vdd.n1669 vdd.n1642 12.0247
R3963 vdd.n1720 vdd.n1693 12.0247
R3964 vdd.n1577 vdd.n1345 11.337
R3965 vdd.n1585 vdd.n1334 11.337
R3966 vdd.n1593 vdd.n1334 11.337
R3967 vdd.n1601 vdd.n1328 11.337
R3968 vdd.n1609 vdd.n1321 11.337
R3969 vdd.n1618 vdd.n1617 11.337
R3970 vdd.n1626 vdd.n1310 11.337
R3971 vdd.n1924 vdd.n1299 11.337
R3972 vdd.n1933 vdd.n1293 11.337
R3973 vdd.n1941 vdd.n1287 11.337
R3974 vdd.n1950 vdd.n1949 11.337
R3975 vdd.n1958 vdd.n1270 11.337
R3976 vdd.n1969 vdd.n1270 11.337
R3977 vdd.n1969 vdd.n1968 11.337
R3978 vdd.n3040 vdd.n511 11.337
R3979 vdd.n3040 vdd.n505 11.337
R3980 vdd.n3048 vdd.n505 11.337
R3981 vdd.n3056 vdd.n499 11.337
R3982 vdd.n3064 vdd.n492 11.337
R3983 vdd.n3073 vdd.n3072 11.337
R3984 vdd.n3081 vdd.n481 11.337
R3985 vdd.n3255 vdd.n3254 11.337
R3986 vdd.n3248 vdd.n325 11.337
R3987 vdd.n3246 vdd.n329 11.337
R3988 vdd.n3240 vdd.n3239 11.337
R3989 vdd.n3238 vdd.n340 11.337
R3990 vdd.n3232 vdd.n340 11.337
R3991 vdd.n3231 vdd.n3230 11.337
R3992 vdd.n296 vdd.n295 11.249
R3993 vdd.n245 vdd.n244 11.249
R3994 vdd.n202 vdd.n201 11.249
R3995 vdd.n151 vdd.n150 11.249
R3996 vdd.n109 vdd.n108 11.249
R3997 vdd.n58 vdd.n57 11.249
R3998 vdd.n1853 vdd.n1852 11.249
R3999 vdd.n1904 vdd.n1903 11.249
R4000 vdd.n1759 vdd.n1758 11.249
R4001 vdd.n1810 vdd.n1809 11.249
R4002 vdd.n1666 vdd.n1665 11.249
R4003 vdd.n1717 vdd.n1716 11.249
R4004 vdd.n1593 vdd.t148 10.9969
R4005 vdd.t159 vdd.n3238 10.9969
R4006 vdd.n1322 vdd.t142 10.7702
R4007 vdd.t194 vdd.n3247 10.7702
R4008 vdd.n281 vdd.n280 10.7238
R4009 vdd.n230 vdd.n229 10.7238
R4010 vdd.n187 vdd.n186 10.7238
R4011 vdd.n136 vdd.n135 10.7238
R4012 vdd.n94 vdd.n93 10.7238
R4013 vdd.n43 vdd.n42 10.7238
R4014 vdd.n1838 vdd.n1837 10.7238
R4015 vdd.n1889 vdd.n1888 10.7238
R4016 vdd.n1744 vdd.n1743 10.7238
R4017 vdd.n1795 vdd.n1794 10.7238
R4018 vdd.n1651 vdd.n1650 10.7238
R4019 vdd.n1702 vdd.n1701 10.7238
R4020 vdd.n2305 vdd.t110 10.6568
R4021 vdd.t7 vdd.n756 10.6568
R4022 vdd.n2138 vdd.n902 10.6151
R4023 vdd.n2139 vdd.n2138 10.6151
R4024 vdd.n2140 vdd.n2139 10.6151
R4025 vdd.n2140 vdd.n891 10.6151
R4026 vdd.n2150 vdd.n891 10.6151
R4027 vdd.n2151 vdd.n2150 10.6151
R4028 vdd.n2152 vdd.n2151 10.6151
R4029 vdd.n2152 vdd.n878 10.6151
R4030 vdd.n2162 vdd.n878 10.6151
R4031 vdd.n2163 vdd.n2162 10.6151
R4032 vdd.n2164 vdd.n2163 10.6151
R4033 vdd.n2164 vdd.n866 10.6151
R4034 vdd.n2175 vdd.n866 10.6151
R4035 vdd.n2176 vdd.n2175 10.6151
R4036 vdd.n2177 vdd.n2176 10.6151
R4037 vdd.n2177 vdd.n854 10.6151
R4038 vdd.n2187 vdd.n854 10.6151
R4039 vdd.n2188 vdd.n2187 10.6151
R4040 vdd.n2189 vdd.n2188 10.6151
R4041 vdd.n2189 vdd.n842 10.6151
R4042 vdd.n2199 vdd.n842 10.6151
R4043 vdd.n2200 vdd.n2199 10.6151
R4044 vdd.n2201 vdd.n2200 10.6151
R4045 vdd.n2201 vdd.n831 10.6151
R4046 vdd.n2211 vdd.n831 10.6151
R4047 vdd.n2212 vdd.n2211 10.6151
R4048 vdd.n2213 vdd.n2212 10.6151
R4049 vdd.n2213 vdd.n818 10.6151
R4050 vdd.n2225 vdd.n818 10.6151
R4051 vdd.n2226 vdd.n2225 10.6151
R4052 vdd.n2228 vdd.n2226 10.6151
R4053 vdd.n2228 vdd.n2227 10.6151
R4054 vdd.n2227 vdd.n799 10.6151
R4055 vdd.n2375 vdd.n2374 10.6151
R4056 vdd.n2374 vdd.n2373 10.6151
R4057 vdd.n2373 vdd.n2370 10.6151
R4058 vdd.n2370 vdd.n2369 10.6151
R4059 vdd.n2369 vdd.n2366 10.6151
R4060 vdd.n2366 vdd.n2365 10.6151
R4061 vdd.n2365 vdd.n2362 10.6151
R4062 vdd.n2362 vdd.n2361 10.6151
R4063 vdd.n2361 vdd.n2358 10.6151
R4064 vdd.n2358 vdd.n2357 10.6151
R4065 vdd.n2357 vdd.n2354 10.6151
R4066 vdd.n2354 vdd.n2353 10.6151
R4067 vdd.n2353 vdd.n2350 10.6151
R4068 vdd.n2350 vdd.n2349 10.6151
R4069 vdd.n2349 vdd.n2346 10.6151
R4070 vdd.n2346 vdd.n2345 10.6151
R4071 vdd.n2345 vdd.n2342 10.6151
R4072 vdd.n2342 vdd.n2341 10.6151
R4073 vdd.n2341 vdd.n2338 10.6151
R4074 vdd.n2338 vdd.n2337 10.6151
R4075 vdd.n2337 vdd.n2334 10.6151
R4076 vdd.n2334 vdd.n2333 10.6151
R4077 vdd.n2333 vdd.n2330 10.6151
R4078 vdd.n2330 vdd.n2329 10.6151
R4079 vdd.n2329 vdd.n2326 10.6151
R4080 vdd.n2326 vdd.n2325 10.6151
R4081 vdd.n2325 vdd.n2322 10.6151
R4082 vdd.n2322 vdd.n2321 10.6151
R4083 vdd.n2321 vdd.n2318 10.6151
R4084 vdd.n2318 vdd.n2317 10.6151
R4085 vdd.n2317 vdd.n2314 10.6151
R4086 vdd.n2312 vdd.n2309 10.6151
R4087 vdd.n2309 vdd.n2308 10.6151
R4088 vdd.n1139 vdd.n1138 10.6151
R4089 vdd.n1141 vdd.n1139 10.6151
R4090 vdd.n1142 vdd.n1141 10.6151
R4091 vdd.n1144 vdd.n1142 10.6151
R4092 vdd.n1145 vdd.n1144 10.6151
R4093 vdd.n1147 vdd.n1145 10.6151
R4094 vdd.n1148 vdd.n1147 10.6151
R4095 vdd.n1150 vdd.n1148 10.6151
R4096 vdd.n1151 vdd.n1150 10.6151
R4097 vdd.n1153 vdd.n1151 10.6151
R4098 vdd.n1154 vdd.n1153 10.6151
R4099 vdd.n1156 vdd.n1154 10.6151
R4100 vdd.n1157 vdd.n1156 10.6151
R4101 vdd.n1159 vdd.n1157 10.6151
R4102 vdd.n1160 vdd.n1159 10.6151
R4103 vdd.n1162 vdd.n1160 10.6151
R4104 vdd.n1163 vdd.n1162 10.6151
R4105 vdd.n1185 vdd.n1163 10.6151
R4106 vdd.n1185 vdd.n1184 10.6151
R4107 vdd.n1184 vdd.n1183 10.6151
R4108 vdd.n1183 vdd.n1181 10.6151
R4109 vdd.n1181 vdd.n1180 10.6151
R4110 vdd.n1180 vdd.n1178 10.6151
R4111 vdd.n1178 vdd.n1177 10.6151
R4112 vdd.n1177 vdd.n1175 10.6151
R4113 vdd.n1175 vdd.n1174 10.6151
R4114 vdd.n1174 vdd.n1172 10.6151
R4115 vdd.n1172 vdd.n1171 10.6151
R4116 vdd.n1171 vdd.n1169 10.6151
R4117 vdd.n1169 vdd.n1168 10.6151
R4118 vdd.n1168 vdd.n1165 10.6151
R4119 vdd.n1165 vdd.n1164 10.6151
R4120 vdd.n1164 vdd.n802 10.6151
R4121 vdd.n2126 vdd.n2125 10.6151
R4122 vdd.n2125 vdd.n2124 10.6151
R4123 vdd.n2124 vdd.n2123 10.6151
R4124 vdd.n2123 vdd.n2121 10.6151
R4125 vdd.n2121 vdd.n2118 10.6151
R4126 vdd.n2118 vdd.n2117 10.6151
R4127 vdd.n2117 vdd.n2114 10.6151
R4128 vdd.n2114 vdd.n2113 10.6151
R4129 vdd.n2113 vdd.n2110 10.6151
R4130 vdd.n2110 vdd.n2109 10.6151
R4131 vdd.n2109 vdd.n2106 10.6151
R4132 vdd.n2106 vdd.n2105 10.6151
R4133 vdd.n2105 vdd.n2102 10.6151
R4134 vdd.n2102 vdd.n2101 10.6151
R4135 vdd.n2101 vdd.n2098 10.6151
R4136 vdd.n2098 vdd.n2097 10.6151
R4137 vdd.n2097 vdd.n2094 10.6151
R4138 vdd.n2094 vdd.n947 10.6151
R4139 vdd.n1105 vdd.n947 10.6151
R4140 vdd.n1106 vdd.n1105 10.6151
R4141 vdd.n1109 vdd.n1106 10.6151
R4142 vdd.n1110 vdd.n1109 10.6151
R4143 vdd.n1113 vdd.n1110 10.6151
R4144 vdd.n1114 vdd.n1113 10.6151
R4145 vdd.n1117 vdd.n1114 10.6151
R4146 vdd.n1118 vdd.n1117 10.6151
R4147 vdd.n1121 vdd.n1118 10.6151
R4148 vdd.n1122 vdd.n1121 10.6151
R4149 vdd.n1125 vdd.n1122 10.6151
R4150 vdd.n1126 vdd.n1125 10.6151
R4151 vdd.n1129 vdd.n1126 10.6151
R4152 vdd.n1134 vdd.n1131 10.6151
R4153 vdd.n1135 vdd.n1134 10.6151
R4154 vdd.n2578 vdd.n2577 10.6151
R4155 vdd.n2577 vdd.n2576 10.6151
R4156 vdd.n2576 vdd.n2415 10.6151
R4157 vdd.n2520 vdd.n2415 10.6151
R4158 vdd.n2521 vdd.n2520 10.6151
R4159 vdd.n2523 vdd.n2521 10.6151
R4160 vdd.n2524 vdd.n2523 10.6151
R4161 vdd.n2526 vdd.n2524 10.6151
R4162 vdd.n2527 vdd.n2526 10.6151
R4163 vdd.n2557 vdd.n2527 10.6151
R4164 vdd.n2557 vdd.n2556 10.6151
R4165 vdd.n2556 vdd.n2555 10.6151
R4166 vdd.n2555 vdd.n2553 10.6151
R4167 vdd.n2553 vdd.n2552 10.6151
R4168 vdd.n2552 vdd.n2550 10.6151
R4169 vdd.n2550 vdd.n2549 10.6151
R4170 vdd.n2549 vdd.n2547 10.6151
R4171 vdd.n2547 vdd.n2546 10.6151
R4172 vdd.n2546 vdd.n2544 10.6151
R4173 vdd.n2544 vdd.n2543 10.6151
R4174 vdd.n2543 vdd.n2541 10.6151
R4175 vdd.n2541 vdd.n2540 10.6151
R4176 vdd.n2540 vdd.n2538 10.6151
R4177 vdd.n2538 vdd.n2537 10.6151
R4178 vdd.n2537 vdd.n2535 10.6151
R4179 vdd.n2535 vdd.n2534 10.6151
R4180 vdd.n2534 vdd.n2532 10.6151
R4181 vdd.n2532 vdd.n2531 10.6151
R4182 vdd.n2531 vdd.n2529 10.6151
R4183 vdd.n2529 vdd.n2528 10.6151
R4184 vdd.n2528 vdd.n664 10.6151
R4185 vdd.n2796 vdd.n664 10.6151
R4186 vdd.n2797 vdd.n2796 10.6151
R4187 vdd.n2647 vdd.n2646 10.6151
R4188 vdd.n2646 vdd.n2645 10.6151
R4189 vdd.n2645 vdd.n2644 10.6151
R4190 vdd.n2644 vdd.n2642 10.6151
R4191 vdd.n2642 vdd.n2639 10.6151
R4192 vdd.n2639 vdd.n2638 10.6151
R4193 vdd.n2638 vdd.n2635 10.6151
R4194 vdd.n2635 vdd.n2634 10.6151
R4195 vdd.n2634 vdd.n2631 10.6151
R4196 vdd.n2631 vdd.n2630 10.6151
R4197 vdd.n2630 vdd.n2627 10.6151
R4198 vdd.n2627 vdd.n2626 10.6151
R4199 vdd.n2626 vdd.n2623 10.6151
R4200 vdd.n2623 vdd.n2622 10.6151
R4201 vdd.n2622 vdd.n2619 10.6151
R4202 vdd.n2619 vdd.n2618 10.6151
R4203 vdd.n2618 vdd.n2615 10.6151
R4204 vdd.n2615 vdd.n2614 10.6151
R4205 vdd.n2614 vdd.n2611 10.6151
R4206 vdd.n2611 vdd.n2610 10.6151
R4207 vdd.n2610 vdd.n2607 10.6151
R4208 vdd.n2607 vdd.n2606 10.6151
R4209 vdd.n2606 vdd.n2603 10.6151
R4210 vdd.n2603 vdd.n2602 10.6151
R4211 vdd.n2602 vdd.n2599 10.6151
R4212 vdd.n2599 vdd.n2598 10.6151
R4213 vdd.n2598 vdd.n2595 10.6151
R4214 vdd.n2595 vdd.n2594 10.6151
R4215 vdd.n2594 vdd.n2591 10.6151
R4216 vdd.n2591 vdd.n2590 10.6151
R4217 vdd.n2590 vdd.n2587 10.6151
R4218 vdd.n2585 vdd.n2582 10.6151
R4219 vdd.n2582 vdd.n2581 10.6151
R4220 vdd.n2659 vdd.n754 10.6151
R4221 vdd.n2660 vdd.n2659 10.6151
R4222 vdd.n2661 vdd.n2660 10.6151
R4223 vdd.n2661 vdd.n743 10.6151
R4224 vdd.n2671 vdd.n743 10.6151
R4225 vdd.n2672 vdd.n2671 10.6151
R4226 vdd.n2673 vdd.n2672 10.6151
R4227 vdd.n2673 vdd.n731 10.6151
R4228 vdd.n2683 vdd.n731 10.6151
R4229 vdd.n2684 vdd.n2683 10.6151
R4230 vdd.n2685 vdd.n2684 10.6151
R4231 vdd.n2685 vdd.n719 10.6151
R4232 vdd.n2695 vdd.n719 10.6151
R4233 vdd.n2696 vdd.n2695 10.6151
R4234 vdd.n2697 vdd.n2696 10.6151
R4235 vdd.n2697 vdd.n708 10.6151
R4236 vdd.n2707 vdd.n708 10.6151
R4237 vdd.n2708 vdd.n2707 10.6151
R4238 vdd.n2709 vdd.n2708 10.6151
R4239 vdd.n2709 vdd.n694 10.6151
R4240 vdd.n2720 vdd.n694 10.6151
R4241 vdd.n2721 vdd.n2720 10.6151
R4242 vdd.n2722 vdd.n2721 10.6151
R4243 vdd.n2722 vdd.n683 10.6151
R4244 vdd.n2732 vdd.n683 10.6151
R4245 vdd.n2733 vdd.n2732 10.6151
R4246 vdd.n2734 vdd.n2733 10.6151
R4247 vdd.n2734 vdd.n669 10.6151
R4248 vdd.n2789 vdd.n669 10.6151
R4249 vdd.n2790 vdd.n2789 10.6151
R4250 vdd.n2791 vdd.n2790 10.6151
R4251 vdd.n2791 vdd.n636 10.6151
R4252 vdd.n2861 vdd.n636 10.6151
R4253 vdd.n2860 vdd.n2859 10.6151
R4254 vdd.n2859 vdd.n637 10.6151
R4255 vdd.n638 vdd.n637 10.6151
R4256 vdd.n2852 vdd.n638 10.6151
R4257 vdd.n2852 vdd.n2851 10.6151
R4258 vdd.n2851 vdd.n2850 10.6151
R4259 vdd.n2850 vdd.n640 10.6151
R4260 vdd.n2845 vdd.n640 10.6151
R4261 vdd.n2845 vdd.n2844 10.6151
R4262 vdd.n2844 vdd.n2843 10.6151
R4263 vdd.n2843 vdd.n643 10.6151
R4264 vdd.n2838 vdd.n643 10.6151
R4265 vdd.n2838 vdd.n2837 10.6151
R4266 vdd.n2837 vdd.n2836 10.6151
R4267 vdd.n2836 vdd.n646 10.6151
R4268 vdd.n2831 vdd.n646 10.6151
R4269 vdd.n2831 vdd.n2830 10.6151
R4270 vdd.n2830 vdd.n2828 10.6151
R4271 vdd.n2828 vdd.n649 10.6151
R4272 vdd.n2823 vdd.n649 10.6151
R4273 vdd.n2823 vdd.n2822 10.6151
R4274 vdd.n2822 vdd.n2821 10.6151
R4275 vdd.n2821 vdd.n652 10.6151
R4276 vdd.n2816 vdd.n652 10.6151
R4277 vdd.n2816 vdd.n2815 10.6151
R4278 vdd.n2815 vdd.n2814 10.6151
R4279 vdd.n2814 vdd.n655 10.6151
R4280 vdd.n2809 vdd.n655 10.6151
R4281 vdd.n2809 vdd.n2808 10.6151
R4282 vdd.n2808 vdd.n2807 10.6151
R4283 vdd.n2807 vdd.n658 10.6151
R4284 vdd.n2802 vdd.n2801 10.6151
R4285 vdd.n2801 vdd.n2800 10.6151
R4286 vdd.n2779 vdd.n2740 10.6151
R4287 vdd.n2774 vdd.n2740 10.6151
R4288 vdd.n2774 vdd.n2773 10.6151
R4289 vdd.n2773 vdd.n2772 10.6151
R4290 vdd.n2772 vdd.n2742 10.6151
R4291 vdd.n2767 vdd.n2742 10.6151
R4292 vdd.n2767 vdd.n2766 10.6151
R4293 vdd.n2766 vdd.n2765 10.6151
R4294 vdd.n2765 vdd.n2745 10.6151
R4295 vdd.n2760 vdd.n2745 10.6151
R4296 vdd.n2760 vdd.n2759 10.6151
R4297 vdd.n2759 vdd.n2758 10.6151
R4298 vdd.n2758 vdd.n2748 10.6151
R4299 vdd.n2753 vdd.n2748 10.6151
R4300 vdd.n2753 vdd.n2752 10.6151
R4301 vdd.n2752 vdd.n610 10.6151
R4302 vdd.n2896 vdd.n610 10.6151
R4303 vdd.n2896 vdd.n611 10.6151
R4304 vdd.n614 vdd.n611 10.6151
R4305 vdd.n2889 vdd.n614 10.6151
R4306 vdd.n2889 vdd.n2888 10.6151
R4307 vdd.n2888 vdd.n2887 10.6151
R4308 vdd.n2887 vdd.n616 10.6151
R4309 vdd.n2882 vdd.n616 10.6151
R4310 vdd.n2882 vdd.n2881 10.6151
R4311 vdd.n2881 vdd.n2880 10.6151
R4312 vdd.n2880 vdd.n619 10.6151
R4313 vdd.n2875 vdd.n619 10.6151
R4314 vdd.n2875 vdd.n2874 10.6151
R4315 vdd.n2874 vdd.n2873 10.6151
R4316 vdd.n2873 vdd.n622 10.6151
R4317 vdd.n2868 vdd.n2867 10.6151
R4318 vdd.n2867 vdd.n2866 10.6151
R4319 vdd.n2486 vdd.n2485 10.6151
R4320 vdd.n2572 vdd.n2486 10.6151
R4321 vdd.n2572 vdd.n2571 10.6151
R4322 vdd.n2571 vdd.n2570 10.6151
R4323 vdd.n2570 vdd.n2568 10.6151
R4324 vdd.n2568 vdd.n2567 10.6151
R4325 vdd.n2567 vdd.n2565 10.6151
R4326 vdd.n2565 vdd.n2564 10.6151
R4327 vdd.n2564 vdd.n2562 10.6151
R4328 vdd.n2562 vdd.n2561 10.6151
R4329 vdd.n2561 vdd.n2518 10.6151
R4330 vdd.n2518 vdd.n2517 10.6151
R4331 vdd.n2517 vdd.n2515 10.6151
R4332 vdd.n2515 vdd.n2514 10.6151
R4333 vdd.n2514 vdd.n2512 10.6151
R4334 vdd.n2512 vdd.n2511 10.6151
R4335 vdd.n2511 vdd.n2509 10.6151
R4336 vdd.n2509 vdd.n2508 10.6151
R4337 vdd.n2508 vdd.n2506 10.6151
R4338 vdd.n2506 vdd.n2505 10.6151
R4339 vdd.n2505 vdd.n2503 10.6151
R4340 vdd.n2503 vdd.n2502 10.6151
R4341 vdd.n2502 vdd.n2500 10.6151
R4342 vdd.n2500 vdd.n2499 10.6151
R4343 vdd.n2499 vdd.n2497 10.6151
R4344 vdd.n2497 vdd.n2496 10.6151
R4345 vdd.n2496 vdd.n2494 10.6151
R4346 vdd.n2494 vdd.n2493 10.6151
R4347 vdd.n2493 vdd.n2491 10.6151
R4348 vdd.n2491 vdd.n2490 10.6151
R4349 vdd.n2490 vdd.n2488 10.6151
R4350 vdd.n2488 vdd.n2487 10.6151
R4351 vdd.n2487 vdd.n628 10.6151
R4352 vdd.n2653 vdd.n760 10.6151
R4353 vdd.n2420 vdd.n760 10.6151
R4354 vdd.n2421 vdd.n2420 10.6151
R4355 vdd.n2424 vdd.n2421 10.6151
R4356 vdd.n2425 vdd.n2424 10.6151
R4357 vdd.n2428 vdd.n2425 10.6151
R4358 vdd.n2429 vdd.n2428 10.6151
R4359 vdd.n2432 vdd.n2429 10.6151
R4360 vdd.n2433 vdd.n2432 10.6151
R4361 vdd.n2436 vdd.n2433 10.6151
R4362 vdd.n2437 vdd.n2436 10.6151
R4363 vdd.n2440 vdd.n2437 10.6151
R4364 vdd.n2441 vdd.n2440 10.6151
R4365 vdd.n2444 vdd.n2441 10.6151
R4366 vdd.n2445 vdd.n2444 10.6151
R4367 vdd.n2448 vdd.n2445 10.6151
R4368 vdd.n2449 vdd.n2448 10.6151
R4369 vdd.n2452 vdd.n2449 10.6151
R4370 vdd.n2453 vdd.n2452 10.6151
R4371 vdd.n2456 vdd.n2453 10.6151
R4372 vdd.n2457 vdd.n2456 10.6151
R4373 vdd.n2460 vdd.n2457 10.6151
R4374 vdd.n2461 vdd.n2460 10.6151
R4375 vdd.n2464 vdd.n2461 10.6151
R4376 vdd.n2465 vdd.n2464 10.6151
R4377 vdd.n2468 vdd.n2465 10.6151
R4378 vdd.n2469 vdd.n2468 10.6151
R4379 vdd.n2472 vdd.n2469 10.6151
R4380 vdd.n2473 vdd.n2472 10.6151
R4381 vdd.n2476 vdd.n2473 10.6151
R4382 vdd.n2477 vdd.n2476 10.6151
R4383 vdd.n2482 vdd.n2480 10.6151
R4384 vdd.n2483 vdd.n2482 10.6151
R4385 vdd.n2655 vdd.n2654 10.6151
R4386 vdd.n2655 vdd.n749 10.6151
R4387 vdd.n2665 vdd.n749 10.6151
R4388 vdd.n2666 vdd.n2665 10.6151
R4389 vdd.n2667 vdd.n2666 10.6151
R4390 vdd.n2667 vdd.n737 10.6151
R4391 vdd.n2677 vdd.n737 10.6151
R4392 vdd.n2678 vdd.n2677 10.6151
R4393 vdd.n2679 vdd.n2678 10.6151
R4394 vdd.n2679 vdd.n725 10.6151
R4395 vdd.n2689 vdd.n725 10.6151
R4396 vdd.n2690 vdd.n2689 10.6151
R4397 vdd.n2691 vdd.n2690 10.6151
R4398 vdd.n2691 vdd.n714 10.6151
R4399 vdd.n2701 vdd.n714 10.6151
R4400 vdd.n2702 vdd.n2701 10.6151
R4401 vdd.n2703 vdd.n2702 10.6151
R4402 vdd.n2703 vdd.n701 10.6151
R4403 vdd.n2713 vdd.n701 10.6151
R4404 vdd.n2714 vdd.n2713 10.6151
R4405 vdd.n2716 vdd.n689 10.6151
R4406 vdd.n2726 vdd.n689 10.6151
R4407 vdd.n2727 vdd.n2726 10.6151
R4408 vdd.n2728 vdd.n2727 10.6151
R4409 vdd.n2728 vdd.n677 10.6151
R4410 vdd.n2738 vdd.n677 10.6151
R4411 vdd.n2739 vdd.n2738 10.6151
R4412 vdd.n2785 vdd.n2739 10.6151
R4413 vdd.n2785 vdd.n2784 10.6151
R4414 vdd.n2784 vdd.n2783 10.6151
R4415 vdd.n2783 vdd.n2782 10.6151
R4416 vdd.n2782 vdd.n2780 10.6151
R4417 vdd.n2134 vdd.n2133 10.6151
R4418 vdd.n2134 vdd.n897 10.6151
R4419 vdd.n2144 vdd.n897 10.6151
R4420 vdd.n2145 vdd.n2144 10.6151
R4421 vdd.n2146 vdd.n2145 10.6151
R4422 vdd.n2146 vdd.n885 10.6151
R4423 vdd.n2156 vdd.n885 10.6151
R4424 vdd.n2157 vdd.n2156 10.6151
R4425 vdd.n2158 vdd.n2157 10.6151
R4426 vdd.n2158 vdd.n872 10.6151
R4427 vdd.n2168 vdd.n872 10.6151
R4428 vdd.n2169 vdd.n2168 10.6151
R4429 vdd.n2171 vdd.n860 10.6151
R4430 vdd.n2181 vdd.n860 10.6151
R4431 vdd.n2182 vdd.n2181 10.6151
R4432 vdd.n2183 vdd.n2182 10.6151
R4433 vdd.n2183 vdd.n848 10.6151
R4434 vdd.n2193 vdd.n848 10.6151
R4435 vdd.n2194 vdd.n2193 10.6151
R4436 vdd.n2195 vdd.n2194 10.6151
R4437 vdd.n2195 vdd.n837 10.6151
R4438 vdd.n2205 vdd.n837 10.6151
R4439 vdd.n2206 vdd.n2205 10.6151
R4440 vdd.n2207 vdd.n2206 10.6151
R4441 vdd.n2207 vdd.n825 10.6151
R4442 vdd.n2217 vdd.n825 10.6151
R4443 vdd.n2218 vdd.n2217 10.6151
R4444 vdd.n2221 vdd.n2218 10.6151
R4445 vdd.n2221 vdd.n2220 10.6151
R4446 vdd.n2220 vdd.n2219 10.6151
R4447 vdd.n2219 vdd.n808 10.6151
R4448 vdd.n2303 vdd.n808 10.6151
R4449 vdd.n2302 vdd.n2301 10.6151
R4450 vdd.n2301 vdd.n2298 10.6151
R4451 vdd.n2298 vdd.n2297 10.6151
R4452 vdd.n2297 vdd.n2294 10.6151
R4453 vdd.n2294 vdd.n2293 10.6151
R4454 vdd.n2293 vdd.n2290 10.6151
R4455 vdd.n2290 vdd.n2289 10.6151
R4456 vdd.n2289 vdd.n2286 10.6151
R4457 vdd.n2286 vdd.n2285 10.6151
R4458 vdd.n2285 vdd.n2282 10.6151
R4459 vdd.n2282 vdd.n2281 10.6151
R4460 vdd.n2281 vdd.n2278 10.6151
R4461 vdd.n2278 vdd.n2277 10.6151
R4462 vdd.n2277 vdd.n2274 10.6151
R4463 vdd.n2274 vdd.n2273 10.6151
R4464 vdd.n2273 vdd.n2270 10.6151
R4465 vdd.n2270 vdd.n2269 10.6151
R4466 vdd.n2269 vdd.n2266 10.6151
R4467 vdd.n2266 vdd.n2265 10.6151
R4468 vdd.n2265 vdd.n2262 10.6151
R4469 vdd.n2262 vdd.n2261 10.6151
R4470 vdd.n2261 vdd.n2258 10.6151
R4471 vdd.n2258 vdd.n2257 10.6151
R4472 vdd.n2257 vdd.n2254 10.6151
R4473 vdd.n2254 vdd.n2253 10.6151
R4474 vdd.n2253 vdd.n2250 10.6151
R4475 vdd.n2250 vdd.n2249 10.6151
R4476 vdd.n2249 vdd.n2246 10.6151
R4477 vdd.n2246 vdd.n2245 10.6151
R4478 vdd.n2245 vdd.n2242 10.6151
R4479 vdd.n2242 vdd.n2241 10.6151
R4480 vdd.n2238 vdd.n2237 10.6151
R4481 vdd.n2237 vdd.n2235 10.6151
R4482 vdd.n1216 vdd.n1214 10.6151
R4483 vdd.n1214 vdd.n1213 10.6151
R4484 vdd.n1213 vdd.n1211 10.6151
R4485 vdd.n1211 vdd.n1210 10.6151
R4486 vdd.n1210 vdd.n1208 10.6151
R4487 vdd.n1208 vdd.n1207 10.6151
R4488 vdd.n1207 vdd.n1205 10.6151
R4489 vdd.n1205 vdd.n1204 10.6151
R4490 vdd.n1204 vdd.n1202 10.6151
R4491 vdd.n1202 vdd.n1201 10.6151
R4492 vdd.n1201 vdd.n1199 10.6151
R4493 vdd.n1199 vdd.n1198 10.6151
R4494 vdd.n1198 vdd.n1196 10.6151
R4495 vdd.n1196 vdd.n1195 10.6151
R4496 vdd.n1195 vdd.n1193 10.6151
R4497 vdd.n1193 vdd.n1192 10.6151
R4498 vdd.n1192 vdd.n1190 10.6151
R4499 vdd.n1190 vdd.n1189 10.6151
R4500 vdd.n1189 vdd.n1100 10.6151
R4501 vdd.n1100 vdd.n1099 10.6151
R4502 vdd.n1099 vdd.n1097 10.6151
R4503 vdd.n1097 vdd.n1096 10.6151
R4504 vdd.n1096 vdd.n1094 10.6151
R4505 vdd.n1094 vdd.n1093 10.6151
R4506 vdd.n1093 vdd.n1091 10.6151
R4507 vdd.n1091 vdd.n1090 10.6151
R4508 vdd.n1090 vdd.n1088 10.6151
R4509 vdd.n1088 vdd.n1087 10.6151
R4510 vdd.n1087 vdd.n1085 10.6151
R4511 vdd.n1085 vdd.n1084 10.6151
R4512 vdd.n1084 vdd.n812 10.6151
R4513 vdd.n2233 vdd.n812 10.6151
R4514 vdd.n2234 vdd.n2233 10.6151
R4515 vdd.n2132 vdd.n909 10.6151
R4516 vdd.n1051 vdd.n909 10.6151
R4517 vdd.n1052 vdd.n1051 10.6151
R4518 vdd.n1055 vdd.n1052 10.6151
R4519 vdd.n1056 vdd.n1055 10.6151
R4520 vdd.n1059 vdd.n1056 10.6151
R4521 vdd.n1060 vdd.n1059 10.6151
R4522 vdd.n1063 vdd.n1060 10.6151
R4523 vdd.n1064 vdd.n1063 10.6151
R4524 vdd.n1067 vdd.n1064 10.6151
R4525 vdd.n1068 vdd.n1067 10.6151
R4526 vdd.n1071 vdd.n1068 10.6151
R4527 vdd.n1072 vdd.n1071 10.6151
R4528 vdd.n1075 vdd.n1072 10.6151
R4529 vdd.n1076 vdd.n1075 10.6151
R4530 vdd.n1079 vdd.n1076 10.6151
R4531 vdd.n1250 vdd.n1079 10.6151
R4532 vdd.n1250 vdd.n1249 10.6151
R4533 vdd.n1249 vdd.n1247 10.6151
R4534 vdd.n1247 vdd.n1244 10.6151
R4535 vdd.n1244 vdd.n1243 10.6151
R4536 vdd.n1243 vdd.n1240 10.6151
R4537 vdd.n1240 vdd.n1239 10.6151
R4538 vdd.n1239 vdd.n1236 10.6151
R4539 vdd.n1236 vdd.n1235 10.6151
R4540 vdd.n1235 vdd.n1232 10.6151
R4541 vdd.n1232 vdd.n1231 10.6151
R4542 vdd.n1231 vdd.n1228 10.6151
R4543 vdd.n1228 vdd.n1227 10.6151
R4544 vdd.n1227 vdd.n1224 10.6151
R4545 vdd.n1224 vdd.n1223 10.6151
R4546 vdd.n1220 vdd.n1219 10.6151
R4547 vdd.n1219 vdd.n1217 10.6151
R4548 vdd.n1634 vdd.t150 10.5435
R4549 vdd.n1977 vdd.t44 10.5435
R4550 vdd.n3032 vdd.t40 10.5435
R4551 vdd.n3256 vdd.t146 10.5435
R4552 vdd.n292 vdd.n274 10.4732
R4553 vdd.n241 vdd.n223 10.4732
R4554 vdd.n198 vdd.n180 10.4732
R4555 vdd.n147 vdd.n129 10.4732
R4556 vdd.n105 vdd.n87 10.4732
R4557 vdd.n54 vdd.n36 10.4732
R4558 vdd.n1849 vdd.n1831 10.4732
R4559 vdd.n1900 vdd.n1882 10.4732
R4560 vdd.n1755 vdd.n1737 10.4732
R4561 vdd.n1806 vdd.n1788 10.4732
R4562 vdd.n1662 vdd.n1644 10.4732
R4563 vdd.n1713 vdd.n1695 10.4732
R4564 vdd.n1932 vdd.t185 10.3167
R4565 vdd.t138 vdd.n493 10.3167
R4566 vdd.n1585 vdd.t52 9.86327
R4567 vdd.n3232 vdd.t48 9.86327
R4568 vdd.n2094 vdd.n2093 9.78206
R4569 vdd.n2830 vdd.n2829 9.78206
R4570 vdd.n2897 vdd.n2896 9.78206
R4571 vdd.n1986 vdd.n1250 9.78206
R4572 vdd.n291 vdd.n276 9.69747
R4573 vdd.n240 vdd.n225 9.69747
R4574 vdd.n197 vdd.n182 9.69747
R4575 vdd.n146 vdd.n131 9.69747
R4576 vdd.n104 vdd.n89 9.69747
R4577 vdd.n53 vdd.n38 9.69747
R4578 vdd.n1848 vdd.n1833 9.69747
R4579 vdd.n1899 vdd.n1884 9.69747
R4580 vdd.n1754 vdd.n1739 9.69747
R4581 vdd.n1805 vdd.n1790 9.69747
R4582 vdd.n1661 vdd.n1646 9.69747
R4583 vdd.n1712 vdd.n1697 9.69747
R4584 vdd.n307 vdd.n306 9.45567
R4585 vdd.n256 vdd.n255 9.45567
R4586 vdd.n213 vdd.n212 9.45567
R4587 vdd.n162 vdd.n161 9.45567
R4588 vdd.n120 vdd.n119 9.45567
R4589 vdd.n69 vdd.n68 9.45567
R4590 vdd.n1864 vdd.n1863 9.45567
R4591 vdd.n1915 vdd.n1914 9.45567
R4592 vdd.n1770 vdd.n1769 9.45567
R4593 vdd.n1821 vdd.n1820 9.45567
R4594 vdd.n1677 vdd.n1676 9.45567
R4595 vdd.n1728 vdd.n1727 9.45567
R4596 vdd.n2056 vdd.n977 9.3005
R4597 vdd.n2055 vdd.n2054 9.3005
R4598 vdd.n983 vdd.n982 9.3005
R4599 vdd.n2049 vdd.n987 9.3005
R4600 vdd.n2048 vdd.n988 9.3005
R4601 vdd.n2047 vdd.n989 9.3005
R4602 vdd.n993 vdd.n990 9.3005
R4603 vdd.n2042 vdd.n994 9.3005
R4604 vdd.n2041 vdd.n995 9.3005
R4605 vdd.n2040 vdd.n996 9.3005
R4606 vdd.n1000 vdd.n997 9.3005
R4607 vdd.n2035 vdd.n1001 9.3005
R4608 vdd.n2034 vdd.n1002 9.3005
R4609 vdd.n2033 vdd.n1003 9.3005
R4610 vdd.n1007 vdd.n1004 9.3005
R4611 vdd.n2028 vdd.n1008 9.3005
R4612 vdd.n2027 vdd.n1009 9.3005
R4613 vdd.n2026 vdd.n1010 9.3005
R4614 vdd.n1014 vdd.n1011 9.3005
R4615 vdd.n2021 vdd.n1015 9.3005
R4616 vdd.n2020 vdd.n1016 9.3005
R4617 vdd.n2019 vdd.n2018 9.3005
R4618 vdd.n2017 vdd.n1017 9.3005
R4619 vdd.n2016 vdd.n2015 9.3005
R4620 vdd.n1023 vdd.n1022 9.3005
R4621 vdd.n2010 vdd.n1027 9.3005
R4622 vdd.n2009 vdd.n1028 9.3005
R4623 vdd.n2008 vdd.n1029 9.3005
R4624 vdd.n1033 vdd.n1030 9.3005
R4625 vdd.n2003 vdd.n1034 9.3005
R4626 vdd.n2002 vdd.n1035 9.3005
R4627 vdd.n2001 vdd.n1036 9.3005
R4628 vdd.n1040 vdd.n1037 9.3005
R4629 vdd.n1996 vdd.n1041 9.3005
R4630 vdd.n1995 vdd.n1042 9.3005
R4631 vdd.n1994 vdd.n1043 9.3005
R4632 vdd.n1047 vdd.n1044 9.3005
R4633 vdd.n1989 vdd.n1048 9.3005
R4634 vdd.n2058 vdd.n2057 9.3005
R4635 vdd.n2080 vdd.n948 9.3005
R4636 vdd.n2079 vdd.n956 9.3005
R4637 vdd.n960 vdd.n957 9.3005
R4638 vdd.n2074 vdd.n961 9.3005
R4639 vdd.n2073 vdd.n962 9.3005
R4640 vdd.n2072 vdd.n963 9.3005
R4641 vdd.n967 vdd.n964 9.3005
R4642 vdd.n2067 vdd.n968 9.3005
R4643 vdd.n2066 vdd.n969 9.3005
R4644 vdd.n2065 vdd.n970 9.3005
R4645 vdd.n974 vdd.n971 9.3005
R4646 vdd.n2060 vdd.n975 9.3005
R4647 vdd.n2059 vdd.n976 9.3005
R4648 vdd.n2092 vdd.n2091 9.3005
R4649 vdd.n952 vdd.n951 9.3005
R4650 vdd.n1920 vdd.n1301 9.3005
R4651 vdd.n1922 vdd.n1921 9.3005
R4652 vdd.n1291 vdd.n1290 9.3005
R4653 vdd.n1936 vdd.n1935 9.3005
R4654 vdd.n1937 vdd.n1289 9.3005
R4655 vdd.n1939 vdd.n1938 9.3005
R4656 vdd.n1280 vdd.n1279 9.3005
R4657 vdd.n1953 vdd.n1952 9.3005
R4658 vdd.n1954 vdd.n1278 9.3005
R4659 vdd.n1956 vdd.n1955 9.3005
R4660 vdd.n1268 vdd.n1267 9.3005
R4661 vdd.n1972 vdd.n1971 9.3005
R4662 vdd.n1973 vdd.n1266 9.3005
R4663 vdd.n1975 vdd.n1974 9.3005
R4664 vdd.n283 vdd.n282 9.3005
R4665 vdd.n278 vdd.n277 9.3005
R4666 vdd.n289 vdd.n288 9.3005
R4667 vdd.n291 vdd.n290 9.3005
R4668 vdd.n274 vdd.n273 9.3005
R4669 vdd.n297 vdd.n296 9.3005
R4670 vdd.n299 vdd.n298 9.3005
R4671 vdd.n271 vdd.n268 9.3005
R4672 vdd.n306 vdd.n305 9.3005
R4673 vdd.n232 vdd.n231 9.3005
R4674 vdd.n227 vdd.n226 9.3005
R4675 vdd.n238 vdd.n237 9.3005
R4676 vdd.n240 vdd.n239 9.3005
R4677 vdd.n223 vdd.n222 9.3005
R4678 vdd.n246 vdd.n245 9.3005
R4679 vdd.n248 vdd.n247 9.3005
R4680 vdd.n220 vdd.n217 9.3005
R4681 vdd.n255 vdd.n254 9.3005
R4682 vdd.n189 vdd.n188 9.3005
R4683 vdd.n184 vdd.n183 9.3005
R4684 vdd.n195 vdd.n194 9.3005
R4685 vdd.n197 vdd.n196 9.3005
R4686 vdd.n180 vdd.n179 9.3005
R4687 vdd.n203 vdd.n202 9.3005
R4688 vdd.n205 vdd.n204 9.3005
R4689 vdd.n177 vdd.n174 9.3005
R4690 vdd.n212 vdd.n211 9.3005
R4691 vdd.n138 vdd.n137 9.3005
R4692 vdd.n133 vdd.n132 9.3005
R4693 vdd.n144 vdd.n143 9.3005
R4694 vdd.n146 vdd.n145 9.3005
R4695 vdd.n129 vdd.n128 9.3005
R4696 vdd.n152 vdd.n151 9.3005
R4697 vdd.n154 vdd.n153 9.3005
R4698 vdd.n126 vdd.n123 9.3005
R4699 vdd.n161 vdd.n160 9.3005
R4700 vdd.n96 vdd.n95 9.3005
R4701 vdd.n91 vdd.n90 9.3005
R4702 vdd.n102 vdd.n101 9.3005
R4703 vdd.n104 vdd.n103 9.3005
R4704 vdd.n87 vdd.n86 9.3005
R4705 vdd.n110 vdd.n109 9.3005
R4706 vdd.n112 vdd.n111 9.3005
R4707 vdd.n84 vdd.n81 9.3005
R4708 vdd.n119 vdd.n118 9.3005
R4709 vdd.n45 vdd.n44 9.3005
R4710 vdd.n40 vdd.n39 9.3005
R4711 vdd.n51 vdd.n50 9.3005
R4712 vdd.n53 vdd.n52 9.3005
R4713 vdd.n36 vdd.n35 9.3005
R4714 vdd.n59 vdd.n58 9.3005
R4715 vdd.n61 vdd.n60 9.3005
R4716 vdd.n33 vdd.n30 9.3005
R4717 vdd.n68 vdd.n67 9.3005
R4718 vdd.n2946 vdd.n2945 9.3005
R4719 vdd.n2947 vdd.n578 9.3005
R4720 vdd.n577 vdd.n575 9.3005
R4721 vdd.n2953 vdd.n574 9.3005
R4722 vdd.n2954 vdd.n573 9.3005
R4723 vdd.n2955 vdd.n572 9.3005
R4724 vdd.n571 vdd.n569 9.3005
R4725 vdd.n2961 vdd.n568 9.3005
R4726 vdd.n2962 vdd.n567 9.3005
R4727 vdd.n2963 vdd.n566 9.3005
R4728 vdd.n565 vdd.n563 9.3005
R4729 vdd.n2969 vdd.n562 9.3005
R4730 vdd.n2970 vdd.n561 9.3005
R4731 vdd.n2971 vdd.n560 9.3005
R4732 vdd.n559 vdd.n557 9.3005
R4733 vdd.n2977 vdd.n556 9.3005
R4734 vdd.n2978 vdd.n555 9.3005
R4735 vdd.n2979 vdd.n554 9.3005
R4736 vdd.n553 vdd.n551 9.3005
R4737 vdd.n2985 vdd.n550 9.3005
R4738 vdd.n2986 vdd.n549 9.3005
R4739 vdd.n2987 vdd.n548 9.3005
R4740 vdd.n547 vdd.n545 9.3005
R4741 vdd.n2993 vdd.n542 9.3005
R4742 vdd.n2994 vdd.n541 9.3005
R4743 vdd.n2995 vdd.n540 9.3005
R4744 vdd.n539 vdd.n537 9.3005
R4745 vdd.n3001 vdd.n536 9.3005
R4746 vdd.n3002 vdd.n535 9.3005
R4747 vdd.n3003 vdd.n534 9.3005
R4748 vdd.n533 vdd.n531 9.3005
R4749 vdd.n3009 vdd.n530 9.3005
R4750 vdd.n3010 vdd.n529 9.3005
R4751 vdd.n3011 vdd.n528 9.3005
R4752 vdd.n527 vdd.n525 9.3005
R4753 vdd.n3016 vdd.n524 9.3005
R4754 vdd.n3026 vdd.n518 9.3005
R4755 vdd.n3028 vdd.n3027 9.3005
R4756 vdd.n509 vdd.n508 9.3005
R4757 vdd.n3043 vdd.n3042 9.3005
R4758 vdd.n3044 vdd.n507 9.3005
R4759 vdd.n3046 vdd.n3045 9.3005
R4760 vdd.n497 vdd.n496 9.3005
R4761 vdd.n3059 vdd.n3058 9.3005
R4762 vdd.n3060 vdd.n495 9.3005
R4763 vdd.n3062 vdd.n3061 9.3005
R4764 vdd.n485 vdd.n484 9.3005
R4765 vdd.n3076 vdd.n3075 9.3005
R4766 vdd.n3077 vdd.n483 9.3005
R4767 vdd.n3079 vdd.n3078 9.3005
R4768 vdd.n312 vdd.n310 9.3005
R4769 vdd.n3030 vdd.n3029 9.3005
R4770 vdd.n3259 vdd.n3258 9.3005
R4771 vdd.n313 vdd.n311 9.3005
R4772 vdd.n3252 vdd.n320 9.3005
R4773 vdd.n3251 vdd.n321 9.3005
R4774 vdd.n3250 vdd.n322 9.3005
R4775 vdd.n331 vdd.n323 9.3005
R4776 vdd.n3244 vdd.n332 9.3005
R4777 vdd.n3243 vdd.n333 9.3005
R4778 vdd.n3242 vdd.n334 9.3005
R4779 vdd.n342 vdd.n335 9.3005
R4780 vdd.n3236 vdd.n343 9.3005
R4781 vdd.n3235 vdd.n344 9.3005
R4782 vdd.n3234 vdd.n345 9.3005
R4783 vdd.n353 vdd.n346 9.3005
R4784 vdd.n3228 vdd.n3227 9.3005
R4785 vdd.n3224 vdd.n354 9.3005
R4786 vdd.n3223 vdd.n357 9.3005
R4787 vdd.n361 vdd.n358 9.3005
R4788 vdd.n362 vdd.n359 9.3005
R4789 vdd.n3216 vdd.n363 9.3005
R4790 vdd.n3215 vdd.n364 9.3005
R4791 vdd.n3214 vdd.n365 9.3005
R4792 vdd.n369 vdd.n366 9.3005
R4793 vdd.n3209 vdd.n370 9.3005
R4794 vdd.n3208 vdd.n371 9.3005
R4795 vdd.n3207 vdd.n372 9.3005
R4796 vdd.n376 vdd.n373 9.3005
R4797 vdd.n3202 vdd.n377 9.3005
R4798 vdd.n3201 vdd.n378 9.3005
R4799 vdd.n3200 vdd.n379 9.3005
R4800 vdd.n383 vdd.n380 9.3005
R4801 vdd.n3195 vdd.n384 9.3005
R4802 vdd.n3194 vdd.n385 9.3005
R4803 vdd.n3193 vdd.n3192 9.3005
R4804 vdd.n3191 vdd.n386 9.3005
R4805 vdd.n3190 vdd.n3189 9.3005
R4806 vdd.n392 vdd.n391 9.3005
R4807 vdd.n3184 vdd.n396 9.3005
R4808 vdd.n3183 vdd.n397 9.3005
R4809 vdd.n3182 vdd.n398 9.3005
R4810 vdd.n402 vdd.n399 9.3005
R4811 vdd.n3177 vdd.n403 9.3005
R4812 vdd.n3176 vdd.n404 9.3005
R4813 vdd.n3175 vdd.n405 9.3005
R4814 vdd.n409 vdd.n406 9.3005
R4815 vdd.n3170 vdd.n410 9.3005
R4816 vdd.n3169 vdd.n411 9.3005
R4817 vdd.n3168 vdd.n412 9.3005
R4818 vdd.n416 vdd.n413 9.3005
R4819 vdd.n3163 vdd.n417 9.3005
R4820 vdd.n3162 vdd.n418 9.3005
R4821 vdd.n3161 vdd.n419 9.3005
R4822 vdd.n423 vdd.n420 9.3005
R4823 vdd.n3156 vdd.n424 9.3005
R4824 vdd.n3155 vdd.n425 9.3005
R4825 vdd.n3154 vdd.n3153 9.3005
R4826 vdd.n3152 vdd.n426 9.3005
R4827 vdd.n3151 vdd.n3150 9.3005
R4828 vdd.n432 vdd.n431 9.3005
R4829 vdd.n3145 vdd.n436 9.3005
R4830 vdd.n3144 vdd.n437 9.3005
R4831 vdd.n3143 vdd.n438 9.3005
R4832 vdd.n442 vdd.n439 9.3005
R4833 vdd.n3138 vdd.n443 9.3005
R4834 vdd.n3137 vdd.n444 9.3005
R4835 vdd.n3136 vdd.n445 9.3005
R4836 vdd.n449 vdd.n446 9.3005
R4837 vdd.n3131 vdd.n450 9.3005
R4838 vdd.n3130 vdd.n451 9.3005
R4839 vdd.n3129 vdd.n452 9.3005
R4840 vdd.n456 vdd.n453 9.3005
R4841 vdd.n3124 vdd.n457 9.3005
R4842 vdd.n3123 vdd.n458 9.3005
R4843 vdd.n3122 vdd.n459 9.3005
R4844 vdd.n463 vdd.n460 9.3005
R4845 vdd.n3117 vdd.n464 9.3005
R4846 vdd.n3116 vdd.n465 9.3005
R4847 vdd.n3112 vdd.n3109 9.3005
R4848 vdd.n3226 vdd.n3225 9.3005
R4849 vdd.n3036 vdd.n513 9.3005
R4850 vdd.n3038 vdd.n3037 9.3005
R4851 vdd.n503 vdd.n502 9.3005
R4852 vdd.n3051 vdd.n3050 9.3005
R4853 vdd.n3052 vdd.n501 9.3005
R4854 vdd.n3054 vdd.n3053 9.3005
R4855 vdd.n490 vdd.n489 9.3005
R4856 vdd.n3067 vdd.n3066 9.3005
R4857 vdd.n3068 vdd.n488 9.3005
R4858 vdd.n3070 vdd.n3069 9.3005
R4859 vdd.n478 vdd.n477 9.3005
R4860 vdd.n3084 vdd.n3083 9.3005
R4861 vdd.n3085 vdd.n476 9.3005
R4862 vdd.n3087 vdd.n3086 9.3005
R4863 vdd.n3088 vdd.n475 9.3005
R4864 vdd.n3090 vdd.n3089 9.3005
R4865 vdd.n3091 vdd.n474 9.3005
R4866 vdd.n3093 vdd.n3092 9.3005
R4867 vdd.n3094 vdd.n472 9.3005
R4868 vdd.n3096 vdd.n3095 9.3005
R4869 vdd.n3097 vdd.n471 9.3005
R4870 vdd.n3099 vdd.n3098 9.3005
R4871 vdd.n3100 vdd.n469 9.3005
R4872 vdd.n3102 vdd.n3101 9.3005
R4873 vdd.n3103 vdd.n468 9.3005
R4874 vdd.n3105 vdd.n3104 9.3005
R4875 vdd.n3106 vdd.n466 9.3005
R4876 vdd.n3108 vdd.n3107 9.3005
R4877 vdd.n3035 vdd.n3034 9.3005
R4878 vdd.n2899 vdd.n514 9.3005
R4879 vdd.n2904 vdd.n2898 9.3005
R4880 vdd.n2914 vdd.n605 9.3005
R4881 vdd.n2915 vdd.n604 9.3005
R4882 vdd.n603 vdd.n601 9.3005
R4883 vdd.n2921 vdd.n600 9.3005
R4884 vdd.n2922 vdd.n599 9.3005
R4885 vdd.n2923 vdd.n598 9.3005
R4886 vdd.n597 vdd.n595 9.3005
R4887 vdd.n2929 vdd.n594 9.3005
R4888 vdd.n2930 vdd.n593 9.3005
R4889 vdd.n2931 vdd.n592 9.3005
R4890 vdd.n591 vdd.n589 9.3005
R4891 vdd.n2936 vdd.n588 9.3005
R4892 vdd.n2937 vdd.n587 9.3005
R4893 vdd.n583 vdd.n582 9.3005
R4894 vdd.n2943 vdd.n2942 9.3005
R4895 vdd.n2944 vdd.n579 9.3005
R4896 vdd.n1985 vdd.n1984 9.3005
R4897 vdd.n1980 vdd.n1252 9.3005
R4898 vdd.n1581 vdd.n1341 9.3005
R4899 vdd.n1583 vdd.n1582 9.3005
R4900 vdd.n1332 vdd.n1331 9.3005
R4901 vdd.n1596 vdd.n1595 9.3005
R4902 vdd.n1597 vdd.n1330 9.3005
R4903 vdd.n1599 vdd.n1598 9.3005
R4904 vdd.n1319 vdd.n1318 9.3005
R4905 vdd.n1612 vdd.n1611 9.3005
R4906 vdd.n1613 vdd.n1317 9.3005
R4907 vdd.n1615 vdd.n1614 9.3005
R4908 vdd.n1308 vdd.n1307 9.3005
R4909 vdd.n1629 vdd.n1628 9.3005
R4910 vdd.n1630 vdd.n1306 9.3005
R4911 vdd.n1632 vdd.n1631 9.3005
R4912 vdd.n1297 vdd.n1296 9.3005
R4913 vdd.n1927 vdd.n1926 9.3005
R4914 vdd.n1928 vdd.n1295 9.3005
R4915 vdd.n1930 vdd.n1929 9.3005
R4916 vdd.n1285 vdd.n1284 9.3005
R4917 vdd.n1944 vdd.n1943 9.3005
R4918 vdd.n1945 vdd.n1283 9.3005
R4919 vdd.n1947 vdd.n1946 9.3005
R4920 vdd.n1275 vdd.n1274 9.3005
R4921 vdd.n1961 vdd.n1960 9.3005
R4922 vdd.n1962 vdd.n1272 9.3005
R4923 vdd.n1966 vdd.n1965 9.3005
R4924 vdd.n1964 vdd.n1273 9.3005
R4925 vdd.n1963 vdd.n1263 9.3005
R4926 vdd.n1580 vdd.n1579 9.3005
R4927 vdd.n1475 vdd.n1465 9.3005
R4928 vdd.n1477 vdd.n1476 9.3005
R4929 vdd.n1478 vdd.n1464 9.3005
R4930 vdd.n1480 vdd.n1479 9.3005
R4931 vdd.n1481 vdd.n1457 9.3005
R4932 vdd.n1483 vdd.n1482 9.3005
R4933 vdd.n1484 vdd.n1456 9.3005
R4934 vdd.n1486 vdd.n1485 9.3005
R4935 vdd.n1487 vdd.n1449 9.3005
R4936 vdd.n1489 vdd.n1488 9.3005
R4937 vdd.n1490 vdd.n1448 9.3005
R4938 vdd.n1492 vdd.n1491 9.3005
R4939 vdd.n1493 vdd.n1441 9.3005
R4940 vdd.n1495 vdd.n1494 9.3005
R4941 vdd.n1496 vdd.n1440 9.3005
R4942 vdd.n1498 vdd.n1497 9.3005
R4943 vdd.n1499 vdd.n1434 9.3005
R4944 vdd.n1501 vdd.n1500 9.3005
R4945 vdd.n1502 vdd.n1432 9.3005
R4946 vdd.n1504 vdd.n1503 9.3005
R4947 vdd.n1433 vdd.n1430 9.3005
R4948 vdd.n1511 vdd.n1426 9.3005
R4949 vdd.n1513 vdd.n1512 9.3005
R4950 vdd.n1514 vdd.n1425 9.3005
R4951 vdd.n1516 vdd.n1515 9.3005
R4952 vdd.n1517 vdd.n1418 9.3005
R4953 vdd.n1519 vdd.n1518 9.3005
R4954 vdd.n1520 vdd.n1417 9.3005
R4955 vdd.n1522 vdd.n1521 9.3005
R4956 vdd.n1523 vdd.n1410 9.3005
R4957 vdd.n1525 vdd.n1524 9.3005
R4958 vdd.n1526 vdd.n1409 9.3005
R4959 vdd.n1528 vdd.n1527 9.3005
R4960 vdd.n1529 vdd.n1402 9.3005
R4961 vdd.n1531 vdd.n1530 9.3005
R4962 vdd.n1532 vdd.n1401 9.3005
R4963 vdd.n1534 vdd.n1533 9.3005
R4964 vdd.n1535 vdd.n1394 9.3005
R4965 vdd.n1537 vdd.n1536 9.3005
R4966 vdd.n1538 vdd.n1393 9.3005
R4967 vdd.n1540 vdd.n1539 9.3005
R4968 vdd.n1541 vdd.n1386 9.3005
R4969 vdd.n1543 vdd.n1542 9.3005
R4970 vdd.n1544 vdd.n1385 9.3005
R4971 vdd.n1546 vdd.n1545 9.3005
R4972 vdd.n1547 vdd.n1376 9.3005
R4973 vdd.n1549 vdd.n1548 9.3005
R4974 vdd.n1550 vdd.n1375 9.3005
R4975 vdd.n1552 vdd.n1551 9.3005
R4976 vdd.n1553 vdd.n1368 9.3005
R4977 vdd.n1555 vdd.n1554 9.3005
R4978 vdd.n1556 vdd.n1367 9.3005
R4979 vdd.n1558 vdd.n1557 9.3005
R4980 vdd.n1559 vdd.n1360 9.3005
R4981 vdd.n1561 vdd.n1560 9.3005
R4982 vdd.n1562 vdd.n1359 9.3005
R4983 vdd.n1564 vdd.n1563 9.3005
R4984 vdd.n1565 vdd.n1352 9.3005
R4985 vdd.n1567 vdd.n1566 9.3005
R4986 vdd.n1568 vdd.n1351 9.3005
R4987 vdd.n1570 vdd.n1569 9.3005
R4988 vdd.n1571 vdd.n1347 9.3005
R4989 vdd.n1573 vdd.n1572 9.3005
R4990 vdd.n1471 vdd.n1342 9.3005
R4991 vdd.n1338 vdd.n1337 9.3005
R4992 vdd.n1588 vdd.n1587 9.3005
R4993 vdd.n1589 vdd.n1336 9.3005
R4994 vdd.n1591 vdd.n1590 9.3005
R4995 vdd.n1326 vdd.n1325 9.3005
R4996 vdd.n1604 vdd.n1603 9.3005
R4997 vdd.n1605 vdd.n1324 9.3005
R4998 vdd.n1607 vdd.n1606 9.3005
R4999 vdd.n1314 vdd.n1313 9.3005
R5000 vdd.n1621 vdd.n1620 9.3005
R5001 vdd.n1622 vdd.n1312 9.3005
R5002 vdd.n1624 vdd.n1623 9.3005
R5003 vdd.n1303 vdd.n1302 9.3005
R5004 vdd.n1575 vdd.n1574 9.3005
R5005 vdd.n1919 vdd.n1636 9.3005
R5006 vdd.n1840 vdd.n1839 9.3005
R5007 vdd.n1835 vdd.n1834 9.3005
R5008 vdd.n1846 vdd.n1845 9.3005
R5009 vdd.n1848 vdd.n1847 9.3005
R5010 vdd.n1831 vdd.n1830 9.3005
R5011 vdd.n1854 vdd.n1853 9.3005
R5012 vdd.n1856 vdd.n1855 9.3005
R5013 vdd.n1828 vdd.n1825 9.3005
R5014 vdd.n1863 vdd.n1862 9.3005
R5015 vdd.n1891 vdd.n1890 9.3005
R5016 vdd.n1886 vdd.n1885 9.3005
R5017 vdd.n1897 vdd.n1896 9.3005
R5018 vdd.n1899 vdd.n1898 9.3005
R5019 vdd.n1882 vdd.n1881 9.3005
R5020 vdd.n1905 vdd.n1904 9.3005
R5021 vdd.n1907 vdd.n1906 9.3005
R5022 vdd.n1879 vdd.n1876 9.3005
R5023 vdd.n1914 vdd.n1913 9.3005
R5024 vdd.n1746 vdd.n1745 9.3005
R5025 vdd.n1741 vdd.n1740 9.3005
R5026 vdd.n1752 vdd.n1751 9.3005
R5027 vdd.n1754 vdd.n1753 9.3005
R5028 vdd.n1737 vdd.n1736 9.3005
R5029 vdd.n1760 vdd.n1759 9.3005
R5030 vdd.n1762 vdd.n1761 9.3005
R5031 vdd.n1734 vdd.n1731 9.3005
R5032 vdd.n1769 vdd.n1768 9.3005
R5033 vdd.n1797 vdd.n1796 9.3005
R5034 vdd.n1792 vdd.n1791 9.3005
R5035 vdd.n1803 vdd.n1802 9.3005
R5036 vdd.n1805 vdd.n1804 9.3005
R5037 vdd.n1788 vdd.n1787 9.3005
R5038 vdd.n1811 vdd.n1810 9.3005
R5039 vdd.n1813 vdd.n1812 9.3005
R5040 vdd.n1785 vdd.n1782 9.3005
R5041 vdd.n1820 vdd.n1819 9.3005
R5042 vdd.n1653 vdd.n1652 9.3005
R5043 vdd.n1648 vdd.n1647 9.3005
R5044 vdd.n1659 vdd.n1658 9.3005
R5045 vdd.n1661 vdd.n1660 9.3005
R5046 vdd.n1644 vdd.n1643 9.3005
R5047 vdd.n1667 vdd.n1666 9.3005
R5048 vdd.n1669 vdd.n1668 9.3005
R5049 vdd.n1641 vdd.n1638 9.3005
R5050 vdd.n1676 vdd.n1675 9.3005
R5051 vdd.n1704 vdd.n1703 9.3005
R5052 vdd.n1699 vdd.n1698 9.3005
R5053 vdd.n1710 vdd.n1709 9.3005
R5054 vdd.n1712 vdd.n1711 9.3005
R5055 vdd.n1695 vdd.n1694 9.3005
R5056 vdd.n1718 vdd.n1717 9.3005
R5057 vdd.n1720 vdd.n1719 9.3005
R5058 vdd.n1692 vdd.n1689 9.3005
R5059 vdd.n1727 vdd.n1726 9.3005
R5060 vdd.n288 vdd.n287 8.92171
R5061 vdd.n237 vdd.n236 8.92171
R5062 vdd.n194 vdd.n193 8.92171
R5063 vdd.n143 vdd.n142 8.92171
R5064 vdd.n101 vdd.n100 8.92171
R5065 vdd.n50 vdd.n49 8.92171
R5066 vdd.n1845 vdd.n1844 8.92171
R5067 vdd.n1896 vdd.n1895 8.92171
R5068 vdd.n1751 vdd.n1750 8.92171
R5069 vdd.n1802 vdd.n1801 8.92171
R5070 vdd.n1658 vdd.n1657 8.92171
R5071 vdd.n1709 vdd.n1708 8.92171
R5072 vdd.n215 vdd.n121 8.81535
R5073 vdd.n1823 vdd.n1729 8.81535
R5074 vdd.n1958 vdd.t168 8.72962
R5075 vdd.n3048 vdd.t166 8.72962
R5076 vdd.t206 vdd.n1932 8.50289
R5077 vdd.n493 vdd.t176 8.50289
R5078 vdd.n28 vdd.n14 8.42249
R5079 vdd.n1634 vdd.t181 8.27616
R5080 vdd.n3256 vdd.t171 8.27616
R5081 vdd.n3260 vdd.n3259 8.16225
R5082 vdd.n1919 vdd.n1918 8.16225
R5083 vdd.n284 vdd.n278 8.14595
R5084 vdd.n233 vdd.n227 8.14595
R5085 vdd.n190 vdd.n184 8.14595
R5086 vdd.n139 vdd.n133 8.14595
R5087 vdd.n97 vdd.n91 8.14595
R5088 vdd.n46 vdd.n40 8.14595
R5089 vdd.n1841 vdd.n1835 8.14595
R5090 vdd.n1892 vdd.n1886 8.14595
R5091 vdd.n1747 vdd.n1741 8.14595
R5092 vdd.n1798 vdd.n1792 8.14595
R5093 vdd.n1654 vdd.n1648 8.14595
R5094 vdd.n1705 vdd.n1699 8.14595
R5095 vdd.t140 vdd.n1322 8.04943
R5096 vdd.n3247 vdd.t174 8.04943
R5097 vdd.n2136 vdd.n904 7.70933
R5098 vdd.n2136 vdd.n907 7.70933
R5099 vdd.n2142 vdd.n893 7.70933
R5100 vdd.n2148 vdd.n893 7.70933
R5101 vdd.n2148 vdd.n887 7.70933
R5102 vdd.n2154 vdd.n887 7.70933
R5103 vdd.n2160 vdd.n880 7.70933
R5104 vdd.n2160 vdd.n883 7.70933
R5105 vdd.n2166 vdd.n876 7.70933
R5106 vdd.n2173 vdd.n862 7.70933
R5107 vdd.n2179 vdd.n862 7.70933
R5108 vdd.n2185 vdd.n856 7.70933
R5109 vdd.n2191 vdd.n852 7.70933
R5110 vdd.n2197 vdd.n846 7.70933
R5111 vdd.n2209 vdd.n833 7.70933
R5112 vdd.n2215 vdd.n827 7.70933
R5113 vdd.n2215 vdd.n820 7.70933
R5114 vdd.n2223 vdd.n820 7.70933
R5115 vdd.n2305 vdd.n804 7.70933
R5116 vdd.n2657 vdd.n756 7.70933
R5117 vdd.n2669 vdd.n745 7.70933
R5118 vdd.n2669 vdd.n739 7.70933
R5119 vdd.n2675 vdd.n739 7.70933
R5120 vdd.n2681 vdd.n733 7.70933
R5121 vdd.n2687 vdd.n729 7.70933
R5122 vdd.n2693 vdd.n723 7.70933
R5123 vdd.n2705 vdd.n710 7.70933
R5124 vdd.n2711 vdd.n703 7.70933
R5125 vdd.n2711 vdd.n706 7.70933
R5126 vdd.n2718 vdd.n698 7.70933
R5127 vdd.n2724 vdd.n685 7.70933
R5128 vdd.n2730 vdd.n685 7.70933
R5129 vdd.n2736 vdd.n679 7.70933
R5130 vdd.n2736 vdd.n671 7.70933
R5131 vdd.n2787 vdd.n671 7.70933
R5132 vdd.n2787 vdd.n674 7.70933
R5133 vdd.n2793 vdd.n631 7.70933
R5134 vdd.n2863 vdd.n631 7.70933
R5135 vdd.n2716 vdd.n2715 7.49318
R5136 vdd.n2170 vdd.n2169 7.49318
R5137 vdd.n283 vdd.n280 7.3702
R5138 vdd.n232 vdd.n229 7.3702
R5139 vdd.n189 vdd.n186 7.3702
R5140 vdd.n138 vdd.n135 7.3702
R5141 vdd.n96 vdd.n93 7.3702
R5142 vdd.n45 vdd.n42 7.3702
R5143 vdd.n1840 vdd.n1837 7.3702
R5144 vdd.n1891 vdd.n1888 7.3702
R5145 vdd.n1746 vdd.n1743 7.3702
R5146 vdd.n1797 vdd.n1794 7.3702
R5147 vdd.n1653 vdd.n1650 7.3702
R5148 vdd.n1704 vdd.n1701 7.3702
R5149 vdd.n2154 vdd.t6 7.36923
R5150 vdd.t16 vdd.n679 7.36923
R5151 vdd.n2230 vdd.t108 7.25587
R5152 vdd.n2574 vdd.t118 7.25587
R5153 vdd.n1601 vdd.t196 7.1425
R5154 vdd.n3240 vdd.t152 7.1425
R5155 vdd.n1512 vdd.n1511 6.98232
R5156 vdd.n2020 vdd.n2019 6.98232
R5157 vdd.n3155 vdd.n3154 6.98232
R5158 vdd.n2947 vdd.n2946 6.98232
R5159 vdd.n1617 vdd.t156 6.91577
R5160 vdd.n325 vdd.t154 6.91577
R5161 vdd.n1924 vdd.t199 6.68904
R5162 vdd.n3081 vdd.t178 6.68904
R5163 vdd.n1287 vdd.t144 6.46231
R5164 vdd.t208 vdd.n492 6.46231
R5165 vdd.n3260 vdd.n309 6.27748
R5166 vdd.n1918 vdd.n1917 6.27748
R5167 vdd.t136 vdd.n833 5.89549
R5168 vdd.n2681 vdd.t25 5.89549
R5169 vdd.n284 vdd.n283 5.81868
R5170 vdd.n233 vdd.n232 5.81868
R5171 vdd.n190 vdd.n189 5.81868
R5172 vdd.n139 vdd.n138 5.81868
R5173 vdd.n97 vdd.n96 5.81868
R5174 vdd.n46 vdd.n45 5.81868
R5175 vdd.n1841 vdd.n1840 5.81868
R5176 vdd.n1892 vdd.n1891 5.81868
R5177 vdd.n1747 vdd.n1746 5.81868
R5178 vdd.n1798 vdd.n1797 5.81868
R5179 vdd.n1654 vdd.n1653 5.81868
R5180 vdd.n1705 vdd.n1704 5.81868
R5181 vdd.n2313 vdd.n2312 5.77611
R5182 vdd.n1131 vdd.n1130 5.77611
R5183 vdd.n2586 vdd.n2585 5.77611
R5184 vdd.n2802 vdd.n663 5.77611
R5185 vdd.n2868 vdd.n627 5.77611
R5186 vdd.n2480 vdd.n2418 5.77611
R5187 vdd.n2238 vdd.n811 5.77611
R5188 vdd.n1220 vdd.n1083 5.77611
R5189 vdd.n1474 vdd.n1471 5.62474
R5190 vdd.n1983 vdd.n1980 5.62474
R5191 vdd.n3115 vdd.n3112 5.62474
R5192 vdd.n2902 vdd.n2899 5.62474
R5193 vdd.t1 vdd.n856 5.55539
R5194 vdd.n2185 vdd.t107 5.55539
R5195 vdd.t19 vdd.n710 5.55539
R5196 vdd.n2705 vdd.t0 5.55539
R5197 vdd.n876 vdd.t86 5.44203
R5198 vdd.n2718 vdd.t65 5.44203
R5199 vdd.n2142 vdd.t36 5.32866
R5200 vdd.n1166 vdd.t78 5.32866
R5201 vdd.n2663 vdd.t82 5.32866
R5202 vdd.n674 vdd.t32 5.32866
R5203 vdd.n287 vdd.n278 5.04292
R5204 vdd.n236 vdd.n227 5.04292
R5205 vdd.n193 vdd.n184 5.04292
R5206 vdd.n142 vdd.n133 5.04292
R5207 vdd.n100 vdd.n91 5.04292
R5208 vdd.n49 vdd.n40 5.04292
R5209 vdd.n1844 vdd.n1835 5.04292
R5210 vdd.n1895 vdd.n1886 5.04292
R5211 vdd.n1750 vdd.n1741 5.04292
R5212 vdd.n1801 vdd.n1792 5.04292
R5213 vdd.n1657 vdd.n1648 5.04292
R5214 vdd.n1708 vdd.n1699 5.04292
R5215 vdd.n2191 vdd.t27 4.98857
R5216 vdd.n723 vdd.t22 4.98857
R5217 vdd.n1950 vdd.t144 4.8752
R5218 vdd.t3 vdd.t120 4.8752
R5219 vdd.t21 vdd.t116 4.8752
R5220 vdd.t13 vdd.t10 4.8752
R5221 vdd.t234 vdd.t9 4.8752
R5222 vdd.n3056 vdd.t208 4.8752
R5223 vdd.n2314 vdd.n2313 4.83952
R5224 vdd.n1130 vdd.n1129 4.83952
R5225 vdd.n2587 vdd.n2586 4.83952
R5226 vdd.n663 vdd.n658 4.83952
R5227 vdd.n627 vdd.n622 4.83952
R5228 vdd.n2477 vdd.n2418 4.83952
R5229 vdd.n2241 vdd.n811 4.83952
R5230 vdd.n1223 vdd.n1083 4.83952
R5231 vdd.n1988 vdd.n1987 4.74817
R5232 vdd.n1256 vdd.n1251 4.74817
R5233 vdd.n953 vdd.n950 4.74817
R5234 vdd.n2081 vdd.n949 4.74817
R5235 vdd.n2086 vdd.n950 4.74817
R5236 vdd.n2085 vdd.n949 4.74817
R5237 vdd.n521 vdd.n519 4.74817
R5238 vdd.n3017 vdd.n522 4.74817
R5239 vdd.n3020 vdd.n522 4.74817
R5240 vdd.n3021 vdd.n521 4.74817
R5241 vdd.n2909 vdd.n606 4.74817
R5242 vdd.n2905 vdd.n608 4.74817
R5243 vdd.n2908 vdd.n608 4.74817
R5244 vdd.n2913 vdd.n606 4.74817
R5245 vdd.n1987 vdd.n1049 4.74817
R5246 vdd.n1253 vdd.n1251 4.74817
R5247 vdd.n309 vdd.n308 4.7074
R5248 vdd.n215 vdd.n214 4.7074
R5249 vdd.n1917 vdd.n1916 4.7074
R5250 vdd.n1823 vdd.n1822 4.7074
R5251 vdd.t199 vdd.n1293 4.64847
R5252 vdd.n2166 vdd.t18 4.64847
R5253 vdd.n846 vdd.t15 4.64847
R5254 vdd.n2687 vdd.t2 4.64847
R5255 vdd.n698 vdd.t17 4.64847
R5256 vdd.n3072 vdd.t178 4.64847
R5257 vdd.n1626 vdd.t156 4.42174
R5258 vdd.n3254 vdd.t154 4.42174
R5259 vdd.n288 vdd.n276 4.26717
R5260 vdd.n237 vdd.n225 4.26717
R5261 vdd.n194 vdd.n182 4.26717
R5262 vdd.n143 vdd.n131 4.26717
R5263 vdd.n101 vdd.n89 4.26717
R5264 vdd.n50 vdd.n38 4.26717
R5265 vdd.n1845 vdd.n1833 4.26717
R5266 vdd.n1896 vdd.n1884 4.26717
R5267 vdd.n1751 vdd.n1739 4.26717
R5268 vdd.n1802 vdd.n1790 4.26717
R5269 vdd.n1658 vdd.n1646 4.26717
R5270 vdd.n1709 vdd.n1697 4.26717
R5271 vdd.t196 vdd.n1321 4.19501
R5272 vdd.t152 vdd.n329 4.19501
R5273 vdd.n309 vdd.n215 4.10845
R5274 vdd.n1917 vdd.n1823 4.10845
R5275 vdd.n265 vdd.t230 4.06363
R5276 vdd.n265 vdd.t165 4.06363
R5277 vdd.n263 vdd.t188 4.06363
R5278 vdd.n263 vdd.t229 4.06363
R5279 vdd.n261 vdd.t231 4.06363
R5280 vdd.n261 vdd.t187 4.06363
R5281 vdd.n259 vdd.t190 4.06363
R5282 vdd.n259 vdd.t192 4.06363
R5283 vdd.n257 vdd.t212 4.06363
R5284 vdd.n257 vdd.t158 4.06363
R5285 vdd.n171 vdd.t223 4.06363
R5286 vdd.n171 vdd.t153 4.06363
R5287 vdd.n169 vdd.t173 4.06363
R5288 vdd.n169 vdd.t222 4.06363
R5289 vdd.n167 vdd.t224 4.06363
R5290 vdd.n167 vdd.t172 4.06363
R5291 vdd.n165 vdd.t177 4.06363
R5292 vdd.n165 vdd.t179 4.06363
R5293 vdd.n163 vdd.t209 4.06363
R5294 vdd.n163 vdd.t139 4.06363
R5295 vdd.n78 vdd.t175 4.06363
R5296 vdd.n78 vdd.t220 4.06363
R5297 vdd.n76 vdd.t155 4.06363
R5298 vdd.n76 vdd.t195 4.06363
R5299 vdd.n74 vdd.t147 4.06363
R5300 vdd.n74 vdd.t180 4.06363
R5301 vdd.n72 vdd.t227 4.06363
R5302 vdd.n72 vdd.t215 4.06363
R5303 vdd.n70 vdd.t217 4.06363
R5304 vdd.n70 vdd.t189 4.06363
R5305 vdd.n1865 vdd.t198 4.06363
R5306 vdd.n1865 vdd.t162 4.06363
R5307 vdd.n1867 vdd.t233 4.06363
R5308 vdd.n1867 vdd.t214 4.06363
R5309 vdd.n1869 vdd.t211 4.06363
R5310 vdd.n1869 vdd.t184 4.06363
R5311 vdd.n1871 vdd.t183 4.06363
R5312 vdd.n1871 vdd.t213 4.06363
R5313 vdd.n1873 vdd.t203 4.06363
R5314 vdd.n1873 vdd.t202 4.06363
R5315 vdd.n1771 vdd.t191 4.06363
R5316 vdd.n1771 vdd.t145 4.06363
R5317 vdd.n1773 vdd.t226 4.06363
R5318 vdd.n1773 vdd.t207 4.06363
R5319 vdd.n1775 vdd.t204 4.06363
R5320 vdd.n1775 vdd.t170 4.06363
R5321 vdd.n1777 vdd.t164 4.06363
R5322 vdd.n1777 vdd.t205 4.06363
R5323 vdd.n1779 vdd.t197 4.06363
R5324 vdd.n1779 vdd.t141 4.06363
R5325 vdd.n1678 vdd.t186 4.06363
R5326 vdd.n1678 vdd.t218 4.06363
R5327 vdd.n1680 vdd.t200 4.06363
R5328 vdd.n1680 vdd.t228 4.06363
R5329 vdd.n1682 vdd.t182 4.06363
R5330 vdd.n1682 vdd.t151 4.06363
R5331 vdd.n1684 vdd.t143 4.06363
R5332 vdd.n1684 vdd.t157 4.06363
R5333 vdd.n1686 vdd.t221 4.06363
R5334 vdd.n1686 vdd.t232 4.06363
R5335 vdd.n26 vdd.t130 3.9605
R5336 vdd.n26 vdd.t131 3.9605
R5337 vdd.n23 vdd.t132 3.9605
R5338 vdd.n23 vdd.t129 3.9605
R5339 vdd.n21 vdd.t128 3.9605
R5340 vdd.n21 vdd.t122 3.9605
R5341 vdd.n20 vdd.t134 3.9605
R5342 vdd.n20 vdd.t126 3.9605
R5343 vdd.n15 vdd.t127 3.9605
R5344 vdd.n15 vdd.t135 3.9605
R5345 vdd.n16 vdd.t133 3.9605
R5346 vdd.n16 vdd.t125 3.9605
R5347 vdd.n18 vdd.t123 3.9605
R5348 vdd.n18 vdd.t4 3.9605
R5349 vdd.n25 vdd.t124 3.9605
R5350 vdd.n25 vdd.t5 3.9605
R5351 vdd.n2223 vdd.t112 3.85492
R5352 vdd.n1166 vdd.t112 3.85492
R5353 vdd.n2663 vdd.t114 3.85492
R5354 vdd.t114 vdd.n745 3.85492
R5355 vdd.n7 vdd.t235 3.61217
R5356 vdd.n7 vdd.t23 3.61217
R5357 vdd.n8 vdd.t14 3.61217
R5358 vdd.n8 vdd.t26 3.61217
R5359 vdd.n10 vdd.t119 3.61217
R5360 vdd.n10 vdd.t115 3.61217
R5361 vdd.n12 vdd.t30 3.61217
R5362 vdd.n12 vdd.t8 3.61217
R5363 vdd.n5 vdd.t111 3.61217
R5364 vdd.n5 vdd.t12 3.61217
R5365 vdd.n3 vdd.t113 3.61217
R5366 vdd.n3 vdd.t109 3.61217
R5367 vdd.n1 vdd.t137 3.61217
R5368 vdd.n1 vdd.t117 3.61217
R5369 vdd.n0 vdd.t28 3.61217
R5370 vdd.n0 vdd.t121 3.61217
R5371 vdd.n292 vdd.n291 3.49141
R5372 vdd.n241 vdd.n240 3.49141
R5373 vdd.n198 vdd.n197 3.49141
R5374 vdd.n147 vdd.n146 3.49141
R5375 vdd.n105 vdd.n104 3.49141
R5376 vdd.n54 vdd.n53 3.49141
R5377 vdd.n1849 vdd.n1848 3.49141
R5378 vdd.n1900 vdd.n1899 3.49141
R5379 vdd.n1755 vdd.n1754 3.49141
R5380 vdd.n1806 vdd.n1805 3.49141
R5381 vdd.n1662 vdd.n1661 3.49141
R5382 vdd.n1713 vdd.n1712 3.49141
R5383 vdd.n2377 vdd.t110 3.40145
R5384 vdd.n2650 vdd.t7 3.40145
R5385 vdd.n1609 vdd.t140 3.28809
R5386 vdd.t174 vdd.n3246 3.28809
R5387 vdd.n2715 vdd.n2714 3.12245
R5388 vdd.n2171 vdd.n2170 3.12245
R5389 vdd.n1310 vdd.t181 3.06136
R5390 vdd.n883 vdd.t18 3.06136
R5391 vdd.n2203 vdd.t15 3.06136
R5392 vdd.n2559 vdd.t2 3.06136
R5393 vdd.n2724 vdd.t17 3.06136
R5394 vdd.t171 vdd.n3255 3.06136
R5395 vdd.n1933 vdd.t206 2.83463
R5396 vdd.n3073 vdd.t176 2.83463
R5397 vdd.n1187 vdd.t27 2.72126
R5398 vdd.n2699 vdd.t22 2.72126
R5399 vdd.n295 vdd.n274 2.71565
R5400 vdd.n244 vdd.n223 2.71565
R5401 vdd.n201 vdd.n180 2.71565
R5402 vdd.n150 vdd.n129 2.71565
R5403 vdd.n108 vdd.n87 2.71565
R5404 vdd.n57 vdd.n36 2.71565
R5405 vdd.n1852 vdd.n1831 2.71565
R5406 vdd.n1903 vdd.n1882 2.71565
R5407 vdd.n1758 vdd.n1737 2.71565
R5408 vdd.n1809 vdd.n1788 2.71565
R5409 vdd.n1665 vdd.n1644 2.71565
R5410 vdd.n1716 vdd.n1695 2.71565
R5411 vdd.n1949 vdd.t168 2.6079
R5412 vdd.t166 vdd.n499 2.6079
R5413 vdd.t116 vdd.n827 2.49453
R5414 vdd.n2675 vdd.t13 2.49453
R5415 vdd.n282 vdd.n281 2.4129
R5416 vdd.n231 vdd.n230 2.4129
R5417 vdd.n188 vdd.n187 2.4129
R5418 vdd.n137 vdd.n136 2.4129
R5419 vdd.n95 vdd.n94 2.4129
R5420 vdd.n44 vdd.n43 2.4129
R5421 vdd.n1839 vdd.n1838 2.4129
R5422 vdd.n1890 vdd.n1889 2.4129
R5423 vdd.n1745 vdd.n1744 2.4129
R5424 vdd.n1796 vdd.n1795 2.4129
R5425 vdd.n1652 vdd.n1651 2.4129
R5426 vdd.n1703 vdd.n1702 2.4129
R5427 vdd.n907 vdd.t36 2.38117
R5428 vdd.n2230 vdd.t78 2.38117
R5429 vdd.n2574 vdd.t82 2.38117
R5430 vdd.n2793 vdd.t32 2.38117
R5431 vdd.n2093 vdd.n950 2.27742
R5432 vdd.n2093 vdd.n949 2.27742
R5433 vdd.n2829 vdd.n522 2.27742
R5434 vdd.n2829 vdd.n521 2.27742
R5435 vdd.n2897 vdd.n608 2.27742
R5436 vdd.n2897 vdd.n606 2.27742
R5437 vdd.n1987 vdd.n1986 2.27742
R5438 vdd.n1986 vdd.n1251 2.27742
R5439 vdd.n2179 vdd.t1 2.15444
R5440 vdd.n1187 vdd.t107 2.15444
R5441 vdd.n2699 vdd.t19 2.15444
R5442 vdd.t0 vdd.n703 2.15444
R5443 vdd.n296 vdd.n272 1.93989
R5444 vdd.n245 vdd.n221 1.93989
R5445 vdd.n202 vdd.n178 1.93989
R5446 vdd.n151 vdd.n127 1.93989
R5447 vdd.n109 vdd.n85 1.93989
R5448 vdd.n58 vdd.n34 1.93989
R5449 vdd.n1853 vdd.n1829 1.93989
R5450 vdd.n1904 vdd.n1880 1.93989
R5451 vdd.n1759 vdd.n1735 1.93989
R5452 vdd.n1810 vdd.n1786 1.93989
R5453 vdd.n1666 vdd.n1642 1.93989
R5454 vdd.n1717 vdd.n1693 1.93989
R5455 vdd.n2203 vdd.t136 1.81434
R5456 vdd.n2559 vdd.t25 1.81434
R5457 vdd.n2197 vdd.t120 1.58761
R5458 vdd.n729 vdd.t234 1.58761
R5459 vdd.n1345 vdd.t52 1.47425
R5460 vdd.t48 vdd.n3231 1.47425
R5461 vdd.n2173 vdd.t24 1.24752
R5462 vdd.n852 vdd.t3 1.24752
R5463 vdd.n2693 vdd.t9 1.24752
R5464 vdd.n706 vdd.t20 1.24752
R5465 vdd.n307 vdd.n267 1.16414
R5466 vdd.n300 vdd.n299 1.16414
R5467 vdd.n256 vdd.n216 1.16414
R5468 vdd.n249 vdd.n248 1.16414
R5469 vdd.n213 vdd.n173 1.16414
R5470 vdd.n206 vdd.n205 1.16414
R5471 vdd.n162 vdd.n122 1.16414
R5472 vdd.n155 vdd.n154 1.16414
R5473 vdd.n120 vdd.n80 1.16414
R5474 vdd.n113 vdd.n112 1.16414
R5475 vdd.n69 vdd.n29 1.16414
R5476 vdd.n62 vdd.n61 1.16414
R5477 vdd.n1864 vdd.n1824 1.16414
R5478 vdd.n1857 vdd.n1856 1.16414
R5479 vdd.n1915 vdd.n1875 1.16414
R5480 vdd.n1908 vdd.n1907 1.16414
R5481 vdd.n1770 vdd.n1730 1.16414
R5482 vdd.n1763 vdd.n1762 1.16414
R5483 vdd.n1821 vdd.n1781 1.16414
R5484 vdd.n1814 vdd.n1813 1.16414
R5485 vdd.n1677 vdd.n1637 1.16414
R5486 vdd.n1670 vdd.n1669 1.16414
R5487 vdd.n1728 vdd.n1688 1.16414
R5488 vdd.n1721 vdd.n1720 1.16414
R5489 vdd.n1941 vdd.t185 1.02079
R5490 vdd.t86 vdd.t24 1.02079
R5491 vdd.t20 vdd.t65 1.02079
R5492 vdd.n3064 vdd.t138 1.02079
R5493 vdd.n1475 vdd.n1474 0.970197
R5494 vdd.n1984 vdd.n1983 0.970197
R5495 vdd.n3116 vdd.n3115 0.970197
R5496 vdd.n2904 vdd.n2902 0.970197
R5497 vdd.n1918 vdd.n28 0.90431
R5498 vdd vdd.n3260 0.896477
R5499 vdd.t150 vdd.n1299 0.794056
R5500 vdd.n1968 vdd.t44 0.794056
R5501 vdd.t40 vdd.n511 0.794056
R5502 vdd.n481 vdd.t146 0.794056
R5503 vdd.n1618 vdd.t142 0.567326
R5504 vdd.n3248 vdd.t194 0.567326
R5505 vdd.n1974 vdd.n951 0.509646
R5506 vdd.n3029 vdd.n3028 0.509646
R5507 vdd.n3227 vdd.n3226 0.509646
R5508 vdd.n3109 vdd.n3108 0.509646
R5509 vdd.n3035 vdd.n514 0.509646
R5510 vdd.n1963 vdd.n1252 0.509646
R5511 vdd.n1580 vdd.n1342 0.509646
R5512 vdd.n1574 vdd.n1573 0.509646
R5513 vdd.n4 vdd.n2 0.459552
R5514 vdd.n11 vdd.n9 0.459552
R5515 vdd.t108 vdd.n804 0.453961
R5516 vdd.n2657 vdd.t118 0.453961
R5517 vdd.n305 vdd.n304 0.388379
R5518 vdd.n271 vdd.n269 0.388379
R5519 vdd.n254 vdd.n253 0.388379
R5520 vdd.n220 vdd.n218 0.388379
R5521 vdd.n211 vdd.n210 0.388379
R5522 vdd.n177 vdd.n175 0.388379
R5523 vdd.n160 vdd.n159 0.388379
R5524 vdd.n126 vdd.n124 0.388379
R5525 vdd.n118 vdd.n117 0.388379
R5526 vdd.n84 vdd.n82 0.388379
R5527 vdd.n67 vdd.n66 0.388379
R5528 vdd.n33 vdd.n31 0.388379
R5529 vdd.n1862 vdd.n1861 0.388379
R5530 vdd.n1828 vdd.n1826 0.388379
R5531 vdd.n1913 vdd.n1912 0.388379
R5532 vdd.n1879 vdd.n1877 0.388379
R5533 vdd.n1768 vdd.n1767 0.388379
R5534 vdd.n1734 vdd.n1732 0.388379
R5535 vdd.n1819 vdd.n1818 0.388379
R5536 vdd.n1785 vdd.n1783 0.388379
R5537 vdd.n1675 vdd.n1674 0.388379
R5538 vdd.n1641 vdd.n1639 0.388379
R5539 vdd.n1726 vdd.n1725 0.388379
R5540 vdd.n1692 vdd.n1690 0.388379
R5541 vdd.n19 vdd.n17 0.387128
R5542 vdd.n24 vdd.n22 0.387128
R5543 vdd.n6 vdd.n4 0.358259
R5544 vdd.n13 vdd.n11 0.358259
R5545 vdd.n260 vdd.n258 0.358259
R5546 vdd.n262 vdd.n260 0.358259
R5547 vdd.n264 vdd.n262 0.358259
R5548 vdd.n266 vdd.n264 0.358259
R5549 vdd.n308 vdd.n266 0.358259
R5550 vdd.n166 vdd.n164 0.358259
R5551 vdd.n168 vdd.n166 0.358259
R5552 vdd.n170 vdd.n168 0.358259
R5553 vdd.n172 vdd.n170 0.358259
R5554 vdd.n214 vdd.n172 0.358259
R5555 vdd.n73 vdd.n71 0.358259
R5556 vdd.n75 vdd.n73 0.358259
R5557 vdd.n77 vdd.n75 0.358259
R5558 vdd.n79 vdd.n77 0.358259
R5559 vdd.n121 vdd.n79 0.358259
R5560 vdd.n1916 vdd.n1874 0.358259
R5561 vdd.n1874 vdd.n1872 0.358259
R5562 vdd.n1872 vdd.n1870 0.358259
R5563 vdd.n1870 vdd.n1868 0.358259
R5564 vdd.n1868 vdd.n1866 0.358259
R5565 vdd.n1822 vdd.n1780 0.358259
R5566 vdd.n1780 vdd.n1778 0.358259
R5567 vdd.n1778 vdd.n1776 0.358259
R5568 vdd.n1776 vdd.n1774 0.358259
R5569 vdd.n1774 vdd.n1772 0.358259
R5570 vdd.n1729 vdd.n1687 0.358259
R5571 vdd.n1687 vdd.n1685 0.358259
R5572 vdd.n1685 vdd.n1683 0.358259
R5573 vdd.n1683 vdd.n1681 0.358259
R5574 vdd.n1681 vdd.n1679 0.358259
R5575 vdd.t148 vdd.n1328 0.340595
R5576 vdd.t6 vdd.n880 0.340595
R5577 vdd.n2209 vdd.t21 0.340595
R5578 vdd.t10 vdd.n733 0.340595
R5579 vdd.n2730 vdd.t16 0.340595
R5580 vdd.n3239 vdd.t159 0.340595
R5581 vdd.n14 vdd.n6 0.334552
R5582 vdd.n14 vdd.n13 0.334552
R5583 vdd.n27 vdd.n19 0.21707
R5584 vdd.n27 vdd.n24 0.21707
R5585 vdd.n306 vdd.n268 0.155672
R5586 vdd.n298 vdd.n268 0.155672
R5587 vdd.n298 vdd.n297 0.155672
R5588 vdd.n297 vdd.n273 0.155672
R5589 vdd.n290 vdd.n273 0.155672
R5590 vdd.n290 vdd.n289 0.155672
R5591 vdd.n289 vdd.n277 0.155672
R5592 vdd.n282 vdd.n277 0.155672
R5593 vdd.n255 vdd.n217 0.155672
R5594 vdd.n247 vdd.n217 0.155672
R5595 vdd.n247 vdd.n246 0.155672
R5596 vdd.n246 vdd.n222 0.155672
R5597 vdd.n239 vdd.n222 0.155672
R5598 vdd.n239 vdd.n238 0.155672
R5599 vdd.n238 vdd.n226 0.155672
R5600 vdd.n231 vdd.n226 0.155672
R5601 vdd.n212 vdd.n174 0.155672
R5602 vdd.n204 vdd.n174 0.155672
R5603 vdd.n204 vdd.n203 0.155672
R5604 vdd.n203 vdd.n179 0.155672
R5605 vdd.n196 vdd.n179 0.155672
R5606 vdd.n196 vdd.n195 0.155672
R5607 vdd.n195 vdd.n183 0.155672
R5608 vdd.n188 vdd.n183 0.155672
R5609 vdd.n161 vdd.n123 0.155672
R5610 vdd.n153 vdd.n123 0.155672
R5611 vdd.n153 vdd.n152 0.155672
R5612 vdd.n152 vdd.n128 0.155672
R5613 vdd.n145 vdd.n128 0.155672
R5614 vdd.n145 vdd.n144 0.155672
R5615 vdd.n144 vdd.n132 0.155672
R5616 vdd.n137 vdd.n132 0.155672
R5617 vdd.n119 vdd.n81 0.155672
R5618 vdd.n111 vdd.n81 0.155672
R5619 vdd.n111 vdd.n110 0.155672
R5620 vdd.n110 vdd.n86 0.155672
R5621 vdd.n103 vdd.n86 0.155672
R5622 vdd.n103 vdd.n102 0.155672
R5623 vdd.n102 vdd.n90 0.155672
R5624 vdd.n95 vdd.n90 0.155672
R5625 vdd.n68 vdd.n30 0.155672
R5626 vdd.n60 vdd.n30 0.155672
R5627 vdd.n60 vdd.n59 0.155672
R5628 vdd.n59 vdd.n35 0.155672
R5629 vdd.n52 vdd.n35 0.155672
R5630 vdd.n52 vdd.n51 0.155672
R5631 vdd.n51 vdd.n39 0.155672
R5632 vdd.n44 vdd.n39 0.155672
R5633 vdd.n1863 vdd.n1825 0.155672
R5634 vdd.n1855 vdd.n1825 0.155672
R5635 vdd.n1855 vdd.n1854 0.155672
R5636 vdd.n1854 vdd.n1830 0.155672
R5637 vdd.n1847 vdd.n1830 0.155672
R5638 vdd.n1847 vdd.n1846 0.155672
R5639 vdd.n1846 vdd.n1834 0.155672
R5640 vdd.n1839 vdd.n1834 0.155672
R5641 vdd.n1914 vdd.n1876 0.155672
R5642 vdd.n1906 vdd.n1876 0.155672
R5643 vdd.n1906 vdd.n1905 0.155672
R5644 vdd.n1905 vdd.n1881 0.155672
R5645 vdd.n1898 vdd.n1881 0.155672
R5646 vdd.n1898 vdd.n1897 0.155672
R5647 vdd.n1897 vdd.n1885 0.155672
R5648 vdd.n1890 vdd.n1885 0.155672
R5649 vdd.n1769 vdd.n1731 0.155672
R5650 vdd.n1761 vdd.n1731 0.155672
R5651 vdd.n1761 vdd.n1760 0.155672
R5652 vdd.n1760 vdd.n1736 0.155672
R5653 vdd.n1753 vdd.n1736 0.155672
R5654 vdd.n1753 vdd.n1752 0.155672
R5655 vdd.n1752 vdd.n1740 0.155672
R5656 vdd.n1745 vdd.n1740 0.155672
R5657 vdd.n1820 vdd.n1782 0.155672
R5658 vdd.n1812 vdd.n1782 0.155672
R5659 vdd.n1812 vdd.n1811 0.155672
R5660 vdd.n1811 vdd.n1787 0.155672
R5661 vdd.n1804 vdd.n1787 0.155672
R5662 vdd.n1804 vdd.n1803 0.155672
R5663 vdd.n1803 vdd.n1791 0.155672
R5664 vdd.n1796 vdd.n1791 0.155672
R5665 vdd.n1676 vdd.n1638 0.155672
R5666 vdd.n1668 vdd.n1638 0.155672
R5667 vdd.n1668 vdd.n1667 0.155672
R5668 vdd.n1667 vdd.n1643 0.155672
R5669 vdd.n1660 vdd.n1643 0.155672
R5670 vdd.n1660 vdd.n1659 0.155672
R5671 vdd.n1659 vdd.n1647 0.155672
R5672 vdd.n1652 vdd.n1647 0.155672
R5673 vdd.n1727 vdd.n1689 0.155672
R5674 vdd.n1719 vdd.n1689 0.155672
R5675 vdd.n1719 vdd.n1718 0.155672
R5676 vdd.n1718 vdd.n1694 0.155672
R5677 vdd.n1711 vdd.n1694 0.155672
R5678 vdd.n1711 vdd.n1710 0.155672
R5679 vdd.n1710 vdd.n1698 0.155672
R5680 vdd.n1703 vdd.n1698 0.155672
R5681 vdd.n956 vdd.n948 0.152939
R5682 vdd.n960 vdd.n956 0.152939
R5683 vdd.n961 vdd.n960 0.152939
R5684 vdd.n962 vdd.n961 0.152939
R5685 vdd.n963 vdd.n962 0.152939
R5686 vdd.n967 vdd.n963 0.152939
R5687 vdd.n968 vdd.n967 0.152939
R5688 vdd.n969 vdd.n968 0.152939
R5689 vdd.n970 vdd.n969 0.152939
R5690 vdd.n974 vdd.n970 0.152939
R5691 vdd.n975 vdd.n974 0.152939
R5692 vdd.n976 vdd.n975 0.152939
R5693 vdd.n2057 vdd.n976 0.152939
R5694 vdd.n2057 vdd.n2056 0.152939
R5695 vdd.n2056 vdd.n2055 0.152939
R5696 vdd.n2055 vdd.n982 0.152939
R5697 vdd.n987 vdd.n982 0.152939
R5698 vdd.n988 vdd.n987 0.152939
R5699 vdd.n989 vdd.n988 0.152939
R5700 vdd.n993 vdd.n989 0.152939
R5701 vdd.n994 vdd.n993 0.152939
R5702 vdd.n995 vdd.n994 0.152939
R5703 vdd.n996 vdd.n995 0.152939
R5704 vdd.n1000 vdd.n996 0.152939
R5705 vdd.n1001 vdd.n1000 0.152939
R5706 vdd.n1002 vdd.n1001 0.152939
R5707 vdd.n1003 vdd.n1002 0.152939
R5708 vdd.n1007 vdd.n1003 0.152939
R5709 vdd.n1008 vdd.n1007 0.152939
R5710 vdd.n1009 vdd.n1008 0.152939
R5711 vdd.n1010 vdd.n1009 0.152939
R5712 vdd.n1014 vdd.n1010 0.152939
R5713 vdd.n1015 vdd.n1014 0.152939
R5714 vdd.n1016 vdd.n1015 0.152939
R5715 vdd.n2018 vdd.n1016 0.152939
R5716 vdd.n2018 vdd.n2017 0.152939
R5717 vdd.n2017 vdd.n2016 0.152939
R5718 vdd.n2016 vdd.n1022 0.152939
R5719 vdd.n1027 vdd.n1022 0.152939
R5720 vdd.n1028 vdd.n1027 0.152939
R5721 vdd.n1029 vdd.n1028 0.152939
R5722 vdd.n1033 vdd.n1029 0.152939
R5723 vdd.n1034 vdd.n1033 0.152939
R5724 vdd.n1035 vdd.n1034 0.152939
R5725 vdd.n1036 vdd.n1035 0.152939
R5726 vdd.n1040 vdd.n1036 0.152939
R5727 vdd.n1041 vdd.n1040 0.152939
R5728 vdd.n1042 vdd.n1041 0.152939
R5729 vdd.n1043 vdd.n1042 0.152939
R5730 vdd.n1047 vdd.n1043 0.152939
R5731 vdd.n1048 vdd.n1047 0.152939
R5732 vdd.n2092 vdd.n951 0.152939
R5733 vdd.n1921 vdd.n1920 0.152939
R5734 vdd.n1921 vdd.n1290 0.152939
R5735 vdd.n1936 vdd.n1290 0.152939
R5736 vdd.n1937 vdd.n1936 0.152939
R5737 vdd.n1938 vdd.n1937 0.152939
R5738 vdd.n1938 vdd.n1279 0.152939
R5739 vdd.n1953 vdd.n1279 0.152939
R5740 vdd.n1954 vdd.n1953 0.152939
R5741 vdd.n1955 vdd.n1954 0.152939
R5742 vdd.n1955 vdd.n1267 0.152939
R5743 vdd.n1972 vdd.n1267 0.152939
R5744 vdd.n1973 vdd.n1972 0.152939
R5745 vdd.n1974 vdd.n1973 0.152939
R5746 vdd.n527 vdd.n524 0.152939
R5747 vdd.n528 vdd.n527 0.152939
R5748 vdd.n529 vdd.n528 0.152939
R5749 vdd.n530 vdd.n529 0.152939
R5750 vdd.n533 vdd.n530 0.152939
R5751 vdd.n534 vdd.n533 0.152939
R5752 vdd.n535 vdd.n534 0.152939
R5753 vdd.n536 vdd.n535 0.152939
R5754 vdd.n539 vdd.n536 0.152939
R5755 vdd.n540 vdd.n539 0.152939
R5756 vdd.n541 vdd.n540 0.152939
R5757 vdd.n542 vdd.n541 0.152939
R5758 vdd.n547 vdd.n542 0.152939
R5759 vdd.n548 vdd.n547 0.152939
R5760 vdd.n549 vdd.n548 0.152939
R5761 vdd.n550 vdd.n549 0.152939
R5762 vdd.n553 vdd.n550 0.152939
R5763 vdd.n554 vdd.n553 0.152939
R5764 vdd.n555 vdd.n554 0.152939
R5765 vdd.n556 vdd.n555 0.152939
R5766 vdd.n559 vdd.n556 0.152939
R5767 vdd.n560 vdd.n559 0.152939
R5768 vdd.n561 vdd.n560 0.152939
R5769 vdd.n562 vdd.n561 0.152939
R5770 vdd.n565 vdd.n562 0.152939
R5771 vdd.n566 vdd.n565 0.152939
R5772 vdd.n567 vdd.n566 0.152939
R5773 vdd.n568 vdd.n567 0.152939
R5774 vdd.n571 vdd.n568 0.152939
R5775 vdd.n572 vdd.n571 0.152939
R5776 vdd.n573 vdd.n572 0.152939
R5777 vdd.n574 vdd.n573 0.152939
R5778 vdd.n577 vdd.n574 0.152939
R5779 vdd.n578 vdd.n577 0.152939
R5780 vdd.n2945 vdd.n578 0.152939
R5781 vdd.n2945 vdd.n2944 0.152939
R5782 vdd.n2944 vdd.n2943 0.152939
R5783 vdd.n2943 vdd.n582 0.152939
R5784 vdd.n587 vdd.n582 0.152939
R5785 vdd.n588 vdd.n587 0.152939
R5786 vdd.n591 vdd.n588 0.152939
R5787 vdd.n592 vdd.n591 0.152939
R5788 vdd.n593 vdd.n592 0.152939
R5789 vdd.n594 vdd.n593 0.152939
R5790 vdd.n597 vdd.n594 0.152939
R5791 vdd.n598 vdd.n597 0.152939
R5792 vdd.n599 vdd.n598 0.152939
R5793 vdd.n600 vdd.n599 0.152939
R5794 vdd.n603 vdd.n600 0.152939
R5795 vdd.n604 vdd.n603 0.152939
R5796 vdd.n605 vdd.n604 0.152939
R5797 vdd.n3028 vdd.n518 0.152939
R5798 vdd.n3029 vdd.n508 0.152939
R5799 vdd.n3043 vdd.n508 0.152939
R5800 vdd.n3044 vdd.n3043 0.152939
R5801 vdd.n3045 vdd.n3044 0.152939
R5802 vdd.n3045 vdd.n496 0.152939
R5803 vdd.n3059 vdd.n496 0.152939
R5804 vdd.n3060 vdd.n3059 0.152939
R5805 vdd.n3061 vdd.n3060 0.152939
R5806 vdd.n3061 vdd.n484 0.152939
R5807 vdd.n3076 vdd.n484 0.152939
R5808 vdd.n3077 vdd.n3076 0.152939
R5809 vdd.n3078 vdd.n3077 0.152939
R5810 vdd.n3078 vdd.n310 0.152939
R5811 vdd.n320 vdd.n311 0.152939
R5812 vdd.n321 vdd.n320 0.152939
R5813 vdd.n322 vdd.n321 0.152939
R5814 vdd.n331 vdd.n322 0.152939
R5815 vdd.n332 vdd.n331 0.152939
R5816 vdd.n333 vdd.n332 0.152939
R5817 vdd.n334 vdd.n333 0.152939
R5818 vdd.n342 vdd.n334 0.152939
R5819 vdd.n343 vdd.n342 0.152939
R5820 vdd.n344 vdd.n343 0.152939
R5821 vdd.n345 vdd.n344 0.152939
R5822 vdd.n353 vdd.n345 0.152939
R5823 vdd.n3227 vdd.n353 0.152939
R5824 vdd.n3226 vdd.n354 0.152939
R5825 vdd.n357 vdd.n354 0.152939
R5826 vdd.n361 vdd.n357 0.152939
R5827 vdd.n362 vdd.n361 0.152939
R5828 vdd.n363 vdd.n362 0.152939
R5829 vdd.n364 vdd.n363 0.152939
R5830 vdd.n365 vdd.n364 0.152939
R5831 vdd.n369 vdd.n365 0.152939
R5832 vdd.n370 vdd.n369 0.152939
R5833 vdd.n371 vdd.n370 0.152939
R5834 vdd.n372 vdd.n371 0.152939
R5835 vdd.n376 vdd.n372 0.152939
R5836 vdd.n377 vdd.n376 0.152939
R5837 vdd.n378 vdd.n377 0.152939
R5838 vdd.n379 vdd.n378 0.152939
R5839 vdd.n383 vdd.n379 0.152939
R5840 vdd.n384 vdd.n383 0.152939
R5841 vdd.n385 vdd.n384 0.152939
R5842 vdd.n3192 vdd.n385 0.152939
R5843 vdd.n3192 vdd.n3191 0.152939
R5844 vdd.n3191 vdd.n3190 0.152939
R5845 vdd.n3190 vdd.n391 0.152939
R5846 vdd.n396 vdd.n391 0.152939
R5847 vdd.n397 vdd.n396 0.152939
R5848 vdd.n398 vdd.n397 0.152939
R5849 vdd.n402 vdd.n398 0.152939
R5850 vdd.n403 vdd.n402 0.152939
R5851 vdd.n404 vdd.n403 0.152939
R5852 vdd.n405 vdd.n404 0.152939
R5853 vdd.n409 vdd.n405 0.152939
R5854 vdd.n410 vdd.n409 0.152939
R5855 vdd.n411 vdd.n410 0.152939
R5856 vdd.n412 vdd.n411 0.152939
R5857 vdd.n416 vdd.n412 0.152939
R5858 vdd.n417 vdd.n416 0.152939
R5859 vdd.n418 vdd.n417 0.152939
R5860 vdd.n419 vdd.n418 0.152939
R5861 vdd.n423 vdd.n419 0.152939
R5862 vdd.n424 vdd.n423 0.152939
R5863 vdd.n425 vdd.n424 0.152939
R5864 vdd.n3153 vdd.n425 0.152939
R5865 vdd.n3153 vdd.n3152 0.152939
R5866 vdd.n3152 vdd.n3151 0.152939
R5867 vdd.n3151 vdd.n431 0.152939
R5868 vdd.n436 vdd.n431 0.152939
R5869 vdd.n437 vdd.n436 0.152939
R5870 vdd.n438 vdd.n437 0.152939
R5871 vdd.n442 vdd.n438 0.152939
R5872 vdd.n443 vdd.n442 0.152939
R5873 vdd.n444 vdd.n443 0.152939
R5874 vdd.n445 vdd.n444 0.152939
R5875 vdd.n449 vdd.n445 0.152939
R5876 vdd.n450 vdd.n449 0.152939
R5877 vdd.n451 vdd.n450 0.152939
R5878 vdd.n452 vdd.n451 0.152939
R5879 vdd.n456 vdd.n452 0.152939
R5880 vdd.n457 vdd.n456 0.152939
R5881 vdd.n458 vdd.n457 0.152939
R5882 vdd.n459 vdd.n458 0.152939
R5883 vdd.n463 vdd.n459 0.152939
R5884 vdd.n464 vdd.n463 0.152939
R5885 vdd.n465 vdd.n464 0.152939
R5886 vdd.n3109 vdd.n465 0.152939
R5887 vdd.n3036 vdd.n3035 0.152939
R5888 vdd.n3037 vdd.n3036 0.152939
R5889 vdd.n3037 vdd.n502 0.152939
R5890 vdd.n3051 vdd.n502 0.152939
R5891 vdd.n3052 vdd.n3051 0.152939
R5892 vdd.n3053 vdd.n3052 0.152939
R5893 vdd.n3053 vdd.n489 0.152939
R5894 vdd.n3067 vdd.n489 0.152939
R5895 vdd.n3068 vdd.n3067 0.152939
R5896 vdd.n3069 vdd.n3068 0.152939
R5897 vdd.n3069 vdd.n477 0.152939
R5898 vdd.n3084 vdd.n477 0.152939
R5899 vdd.n3085 vdd.n3084 0.152939
R5900 vdd.n3086 vdd.n3085 0.152939
R5901 vdd.n3086 vdd.n475 0.152939
R5902 vdd.n3090 vdd.n475 0.152939
R5903 vdd.n3091 vdd.n3090 0.152939
R5904 vdd.n3092 vdd.n3091 0.152939
R5905 vdd.n3092 vdd.n472 0.152939
R5906 vdd.n3096 vdd.n472 0.152939
R5907 vdd.n3097 vdd.n3096 0.152939
R5908 vdd.n3098 vdd.n3097 0.152939
R5909 vdd.n3098 vdd.n469 0.152939
R5910 vdd.n3102 vdd.n469 0.152939
R5911 vdd.n3103 vdd.n3102 0.152939
R5912 vdd.n3104 vdd.n3103 0.152939
R5913 vdd.n3104 vdd.n466 0.152939
R5914 vdd.n3108 vdd.n466 0.152939
R5915 vdd.n2898 vdd.n514 0.152939
R5916 vdd.n1985 vdd.n1252 0.152939
R5917 vdd.n1581 vdd.n1580 0.152939
R5918 vdd.n1582 vdd.n1581 0.152939
R5919 vdd.n1582 vdd.n1331 0.152939
R5920 vdd.n1596 vdd.n1331 0.152939
R5921 vdd.n1597 vdd.n1596 0.152939
R5922 vdd.n1598 vdd.n1597 0.152939
R5923 vdd.n1598 vdd.n1318 0.152939
R5924 vdd.n1612 vdd.n1318 0.152939
R5925 vdd.n1613 vdd.n1612 0.152939
R5926 vdd.n1614 vdd.n1613 0.152939
R5927 vdd.n1614 vdd.n1307 0.152939
R5928 vdd.n1629 vdd.n1307 0.152939
R5929 vdd.n1630 vdd.n1629 0.152939
R5930 vdd.n1631 vdd.n1630 0.152939
R5931 vdd.n1631 vdd.n1296 0.152939
R5932 vdd.n1927 vdd.n1296 0.152939
R5933 vdd.n1928 vdd.n1927 0.152939
R5934 vdd.n1929 vdd.n1928 0.152939
R5935 vdd.n1929 vdd.n1284 0.152939
R5936 vdd.n1944 vdd.n1284 0.152939
R5937 vdd.n1945 vdd.n1944 0.152939
R5938 vdd.n1946 vdd.n1945 0.152939
R5939 vdd.n1946 vdd.n1274 0.152939
R5940 vdd.n1961 vdd.n1274 0.152939
R5941 vdd.n1962 vdd.n1961 0.152939
R5942 vdd.n1965 vdd.n1962 0.152939
R5943 vdd.n1965 vdd.n1964 0.152939
R5944 vdd.n1964 vdd.n1963 0.152939
R5945 vdd.n1573 vdd.n1347 0.152939
R5946 vdd.n1569 vdd.n1347 0.152939
R5947 vdd.n1569 vdd.n1568 0.152939
R5948 vdd.n1568 vdd.n1567 0.152939
R5949 vdd.n1567 vdd.n1352 0.152939
R5950 vdd.n1563 vdd.n1352 0.152939
R5951 vdd.n1563 vdd.n1562 0.152939
R5952 vdd.n1562 vdd.n1561 0.152939
R5953 vdd.n1561 vdd.n1360 0.152939
R5954 vdd.n1557 vdd.n1360 0.152939
R5955 vdd.n1557 vdd.n1556 0.152939
R5956 vdd.n1556 vdd.n1555 0.152939
R5957 vdd.n1555 vdd.n1368 0.152939
R5958 vdd.n1551 vdd.n1368 0.152939
R5959 vdd.n1551 vdd.n1550 0.152939
R5960 vdd.n1550 vdd.n1549 0.152939
R5961 vdd.n1549 vdd.n1376 0.152939
R5962 vdd.n1545 vdd.n1376 0.152939
R5963 vdd.n1545 vdd.n1544 0.152939
R5964 vdd.n1544 vdd.n1543 0.152939
R5965 vdd.n1543 vdd.n1386 0.152939
R5966 vdd.n1539 vdd.n1386 0.152939
R5967 vdd.n1539 vdd.n1538 0.152939
R5968 vdd.n1538 vdd.n1537 0.152939
R5969 vdd.n1537 vdd.n1394 0.152939
R5970 vdd.n1533 vdd.n1394 0.152939
R5971 vdd.n1533 vdd.n1532 0.152939
R5972 vdd.n1532 vdd.n1531 0.152939
R5973 vdd.n1531 vdd.n1402 0.152939
R5974 vdd.n1527 vdd.n1402 0.152939
R5975 vdd.n1527 vdd.n1526 0.152939
R5976 vdd.n1526 vdd.n1525 0.152939
R5977 vdd.n1525 vdd.n1410 0.152939
R5978 vdd.n1521 vdd.n1410 0.152939
R5979 vdd.n1521 vdd.n1520 0.152939
R5980 vdd.n1520 vdd.n1519 0.152939
R5981 vdd.n1519 vdd.n1418 0.152939
R5982 vdd.n1515 vdd.n1418 0.152939
R5983 vdd.n1515 vdd.n1514 0.152939
R5984 vdd.n1514 vdd.n1513 0.152939
R5985 vdd.n1513 vdd.n1426 0.152939
R5986 vdd.n1433 vdd.n1426 0.152939
R5987 vdd.n1503 vdd.n1433 0.152939
R5988 vdd.n1503 vdd.n1502 0.152939
R5989 vdd.n1502 vdd.n1501 0.152939
R5990 vdd.n1501 vdd.n1434 0.152939
R5991 vdd.n1497 vdd.n1434 0.152939
R5992 vdd.n1497 vdd.n1496 0.152939
R5993 vdd.n1496 vdd.n1495 0.152939
R5994 vdd.n1495 vdd.n1441 0.152939
R5995 vdd.n1491 vdd.n1441 0.152939
R5996 vdd.n1491 vdd.n1490 0.152939
R5997 vdd.n1490 vdd.n1489 0.152939
R5998 vdd.n1489 vdd.n1449 0.152939
R5999 vdd.n1485 vdd.n1449 0.152939
R6000 vdd.n1485 vdd.n1484 0.152939
R6001 vdd.n1484 vdd.n1483 0.152939
R6002 vdd.n1483 vdd.n1457 0.152939
R6003 vdd.n1479 vdd.n1457 0.152939
R6004 vdd.n1479 vdd.n1478 0.152939
R6005 vdd.n1478 vdd.n1477 0.152939
R6006 vdd.n1477 vdd.n1465 0.152939
R6007 vdd.n1465 vdd.n1342 0.152939
R6008 vdd.n1574 vdd.n1337 0.152939
R6009 vdd.n1588 vdd.n1337 0.152939
R6010 vdd.n1589 vdd.n1588 0.152939
R6011 vdd.n1590 vdd.n1589 0.152939
R6012 vdd.n1590 vdd.n1325 0.152939
R6013 vdd.n1604 vdd.n1325 0.152939
R6014 vdd.n1605 vdd.n1604 0.152939
R6015 vdd.n1606 vdd.n1605 0.152939
R6016 vdd.n1606 vdd.n1313 0.152939
R6017 vdd.n1621 vdd.n1313 0.152939
R6018 vdd.n1622 vdd.n1621 0.152939
R6019 vdd.n1623 vdd.n1622 0.152939
R6020 vdd.n1623 vdd.n1302 0.152939
R6021 vdd.n1920 vdd.n1919 0.145814
R6022 vdd.n3259 vdd.n310 0.145814
R6023 vdd.n3259 vdd.n311 0.145814
R6024 vdd.n1919 vdd.n1302 0.145814
R6025 vdd.n2093 vdd.n2092 0.110256
R6026 vdd.n2829 vdd.n518 0.110256
R6027 vdd.n2898 vdd.n2897 0.110256
R6028 vdd.n1986 vdd.n1985 0.110256
R6029 vdd.n2093 vdd.n948 0.0431829
R6030 vdd.n1986 vdd.n1048 0.0431829
R6031 vdd.n2829 vdd.n524 0.0431829
R6032 vdd.n2897 vdd.n605 0.0431829
R6033 vdd vdd.n28 0.00833333
R6034 CSoutput.n19 CSoutput.t211 184.661
R6035 CSoutput.n78 CSoutput.n77 165.8
R6036 CSoutput.n76 CSoutput.n0 165.8
R6037 CSoutput.n75 CSoutput.n74 165.8
R6038 CSoutput.n73 CSoutput.n72 165.8
R6039 CSoutput.n71 CSoutput.n2 165.8
R6040 CSoutput.n69 CSoutput.n68 165.8
R6041 CSoutput.n67 CSoutput.n3 165.8
R6042 CSoutput.n66 CSoutput.n65 165.8
R6043 CSoutput.n63 CSoutput.n4 165.8
R6044 CSoutput.n61 CSoutput.n60 165.8
R6045 CSoutput.n59 CSoutput.n5 165.8
R6046 CSoutput.n58 CSoutput.n57 165.8
R6047 CSoutput.n55 CSoutput.n6 165.8
R6048 CSoutput.n54 CSoutput.n53 165.8
R6049 CSoutput.n52 CSoutput.n51 165.8
R6050 CSoutput.n50 CSoutput.n8 165.8
R6051 CSoutput.n48 CSoutput.n47 165.8
R6052 CSoutput.n46 CSoutput.n9 165.8
R6053 CSoutput.n45 CSoutput.n44 165.8
R6054 CSoutput.n42 CSoutput.n10 165.8
R6055 CSoutput.n41 CSoutput.n40 165.8
R6056 CSoutput.n39 CSoutput.n38 165.8
R6057 CSoutput.n37 CSoutput.n12 165.8
R6058 CSoutput.n35 CSoutput.n34 165.8
R6059 CSoutput.n33 CSoutput.n13 165.8
R6060 CSoutput.n32 CSoutput.n31 165.8
R6061 CSoutput.n29 CSoutput.n14 165.8
R6062 CSoutput.n28 CSoutput.n27 165.8
R6063 CSoutput.n26 CSoutput.n25 165.8
R6064 CSoutput.n24 CSoutput.n16 165.8
R6065 CSoutput.n22 CSoutput.n21 165.8
R6066 CSoutput.n20 CSoutput.n17 165.8
R6067 CSoutput.n77 CSoutput.t212 162.194
R6068 CSoutput.n18 CSoutput.t201 120.501
R6069 CSoutput.n23 CSoutput.t203 120.501
R6070 CSoutput.n15 CSoutput.t196 120.501
R6071 CSoutput.n30 CSoutput.t209 120.501
R6072 CSoutput.n36 CSoutput.t204 120.501
R6073 CSoutput.n11 CSoutput.t199 120.501
R6074 CSoutput.n43 CSoutput.t194 120.501
R6075 CSoutput.n49 CSoutput.t205 120.501
R6076 CSoutput.n7 CSoutput.t207 120.501
R6077 CSoutput.n56 CSoutput.t197 120.501
R6078 CSoutput.n62 CSoutput.t193 120.501
R6079 CSoutput.n64 CSoutput.t210 120.501
R6080 CSoutput.n70 CSoutput.t200 120.501
R6081 CSoutput.n1 CSoutput.t202 120.501
R6082 CSoutput.n290 CSoutput.n288 103.469
R6083 CSoutput.n278 CSoutput.n276 103.469
R6084 CSoutput.n267 CSoutput.n265 103.469
R6085 CSoutput.n104 CSoutput.n102 103.469
R6086 CSoutput.n92 CSoutput.n90 103.469
R6087 CSoutput.n81 CSoutput.n79 103.469
R6088 CSoutput.n296 CSoutput.n295 103.111
R6089 CSoutput.n294 CSoutput.n293 103.111
R6090 CSoutput.n292 CSoutput.n291 103.111
R6091 CSoutput.n290 CSoutput.n289 103.111
R6092 CSoutput.n286 CSoutput.n285 103.111
R6093 CSoutput.n284 CSoutput.n283 103.111
R6094 CSoutput.n282 CSoutput.n281 103.111
R6095 CSoutput.n280 CSoutput.n279 103.111
R6096 CSoutput.n278 CSoutput.n277 103.111
R6097 CSoutput.n275 CSoutput.n274 103.111
R6098 CSoutput.n273 CSoutput.n272 103.111
R6099 CSoutput.n271 CSoutput.n270 103.111
R6100 CSoutput.n269 CSoutput.n268 103.111
R6101 CSoutput.n267 CSoutput.n266 103.111
R6102 CSoutput.n104 CSoutput.n103 103.111
R6103 CSoutput.n106 CSoutput.n105 103.111
R6104 CSoutput.n108 CSoutput.n107 103.111
R6105 CSoutput.n110 CSoutput.n109 103.111
R6106 CSoutput.n112 CSoutput.n111 103.111
R6107 CSoutput.n92 CSoutput.n91 103.111
R6108 CSoutput.n94 CSoutput.n93 103.111
R6109 CSoutput.n96 CSoutput.n95 103.111
R6110 CSoutput.n98 CSoutput.n97 103.111
R6111 CSoutput.n100 CSoutput.n99 103.111
R6112 CSoutput.n81 CSoutput.n80 103.111
R6113 CSoutput.n83 CSoutput.n82 103.111
R6114 CSoutput.n85 CSoutput.n84 103.111
R6115 CSoutput.n87 CSoutput.n86 103.111
R6116 CSoutput.n89 CSoutput.n88 103.111
R6117 CSoutput.n298 CSoutput.n297 103.111
R6118 CSoutput.n342 CSoutput.n340 81.5057
R6119 CSoutput.n322 CSoutput.n320 81.5057
R6120 CSoutput.n303 CSoutput.n301 81.5057
R6121 CSoutput.n402 CSoutput.n400 81.5057
R6122 CSoutput.n382 CSoutput.n380 81.5057
R6123 CSoutput.n363 CSoutput.n361 81.5057
R6124 CSoutput.n358 CSoutput.n357 80.9324
R6125 CSoutput.n356 CSoutput.n355 80.9324
R6126 CSoutput.n354 CSoutput.n353 80.9324
R6127 CSoutput.n352 CSoutput.n351 80.9324
R6128 CSoutput.n350 CSoutput.n349 80.9324
R6129 CSoutput.n348 CSoutput.n347 80.9324
R6130 CSoutput.n346 CSoutput.n345 80.9324
R6131 CSoutput.n344 CSoutput.n343 80.9324
R6132 CSoutput.n342 CSoutput.n341 80.9324
R6133 CSoutput.n338 CSoutput.n337 80.9324
R6134 CSoutput.n336 CSoutput.n335 80.9324
R6135 CSoutput.n334 CSoutput.n333 80.9324
R6136 CSoutput.n332 CSoutput.n331 80.9324
R6137 CSoutput.n330 CSoutput.n329 80.9324
R6138 CSoutput.n328 CSoutput.n327 80.9324
R6139 CSoutput.n326 CSoutput.n325 80.9324
R6140 CSoutput.n324 CSoutput.n323 80.9324
R6141 CSoutput.n322 CSoutput.n321 80.9324
R6142 CSoutput.n319 CSoutput.n318 80.9324
R6143 CSoutput.n317 CSoutput.n316 80.9324
R6144 CSoutput.n315 CSoutput.n314 80.9324
R6145 CSoutput.n313 CSoutput.n312 80.9324
R6146 CSoutput.n311 CSoutput.n310 80.9324
R6147 CSoutput.n309 CSoutput.n308 80.9324
R6148 CSoutput.n307 CSoutput.n306 80.9324
R6149 CSoutput.n305 CSoutput.n304 80.9324
R6150 CSoutput.n303 CSoutput.n302 80.9324
R6151 CSoutput.n402 CSoutput.n401 80.9324
R6152 CSoutput.n404 CSoutput.n403 80.9324
R6153 CSoutput.n406 CSoutput.n405 80.9324
R6154 CSoutput.n408 CSoutput.n407 80.9324
R6155 CSoutput.n410 CSoutput.n409 80.9324
R6156 CSoutput.n412 CSoutput.n411 80.9324
R6157 CSoutput.n414 CSoutput.n413 80.9324
R6158 CSoutput.n416 CSoutput.n415 80.9324
R6159 CSoutput.n418 CSoutput.n417 80.9324
R6160 CSoutput.n382 CSoutput.n381 80.9324
R6161 CSoutput.n384 CSoutput.n383 80.9324
R6162 CSoutput.n386 CSoutput.n385 80.9324
R6163 CSoutput.n388 CSoutput.n387 80.9324
R6164 CSoutput.n390 CSoutput.n389 80.9324
R6165 CSoutput.n392 CSoutput.n391 80.9324
R6166 CSoutput.n394 CSoutput.n393 80.9324
R6167 CSoutput.n396 CSoutput.n395 80.9324
R6168 CSoutput.n398 CSoutput.n397 80.9324
R6169 CSoutput.n363 CSoutput.n362 80.9324
R6170 CSoutput.n365 CSoutput.n364 80.9324
R6171 CSoutput.n367 CSoutput.n366 80.9324
R6172 CSoutput.n369 CSoutput.n368 80.9324
R6173 CSoutput.n371 CSoutput.n370 80.9324
R6174 CSoutput.n373 CSoutput.n372 80.9324
R6175 CSoutput.n375 CSoutput.n374 80.9324
R6176 CSoutput.n377 CSoutput.n376 80.9324
R6177 CSoutput.n379 CSoutput.n378 80.9324
R6178 CSoutput.n25 CSoutput.n24 48.1486
R6179 CSoutput.n69 CSoutput.n3 48.1486
R6180 CSoutput.n38 CSoutput.n37 48.1486
R6181 CSoutput.n42 CSoutput.n41 48.1486
R6182 CSoutput.n51 CSoutput.n50 48.1486
R6183 CSoutput.n55 CSoutput.n54 48.1486
R6184 CSoutput.n22 CSoutput.n17 46.462
R6185 CSoutput.n72 CSoutput.n71 46.462
R6186 CSoutput.n20 CSoutput.n19 44.9055
R6187 CSoutput.n29 CSoutput.n28 43.7635
R6188 CSoutput.n65 CSoutput.n63 43.7635
R6189 CSoutput.n35 CSoutput.n13 41.7396
R6190 CSoutput.n57 CSoutput.n5 41.7396
R6191 CSoutput.n44 CSoutput.n9 37.0171
R6192 CSoutput.n48 CSoutput.n9 37.0171
R6193 CSoutput.n76 CSoutput.n75 34.9932
R6194 CSoutput.n31 CSoutput.n13 32.2947
R6195 CSoutput.n61 CSoutput.n5 32.2947
R6196 CSoutput.n30 CSoutput.n29 29.6014
R6197 CSoutput.n63 CSoutput.n62 29.6014
R6198 CSoutput.n19 CSoutput.n18 28.4085
R6199 CSoutput.n18 CSoutput.n17 25.1176
R6200 CSoutput.n72 CSoutput.n1 25.1176
R6201 CSoutput.n43 CSoutput.n42 22.0922
R6202 CSoutput.n50 CSoutput.n49 22.0922
R6203 CSoutput.n77 CSoutput.n76 21.8586
R6204 CSoutput.n37 CSoutput.n36 18.9681
R6205 CSoutput.n56 CSoutput.n55 18.9681
R6206 CSoutput.n25 CSoutput.n15 17.6292
R6207 CSoutput.n64 CSoutput.n3 17.6292
R6208 CSoutput.n24 CSoutput.n23 15.844
R6209 CSoutput.n70 CSoutput.n69 15.844
R6210 CSoutput.n38 CSoutput.n11 14.5051
R6211 CSoutput.n54 CSoutput.n7 14.5051
R6212 CSoutput.n421 CSoutput.n78 11.4982
R6213 CSoutput.n41 CSoutput.n11 11.3811
R6214 CSoutput.n51 CSoutput.n7 11.3811
R6215 CSoutput.n23 CSoutput.n22 10.0422
R6216 CSoutput.n71 CSoutput.n70 10.0422
R6217 CSoutput.n287 CSoutput.n275 9.25285
R6218 CSoutput.n101 CSoutput.n89 9.25285
R6219 CSoutput.n360 CSoutput.n300 9.05363
R6220 CSoutput.n339 CSoutput.n319 8.98182
R6221 CSoutput.n399 CSoutput.n379 8.98182
R6222 CSoutput.n28 CSoutput.n15 8.25698
R6223 CSoutput.n65 CSoutput.n64 8.25698
R6224 CSoutput.n300 CSoutput.n299 7.12641
R6225 CSoutput.n114 CSoutput.n113 7.12641
R6226 CSoutput.n36 CSoutput.n35 6.91809
R6227 CSoutput.n57 CSoutput.n56 6.91809
R6228 CSoutput.n360 CSoutput.n359 6.02792
R6229 CSoutput.n420 CSoutput.n419 6.02792
R6230 CSoutput.n421 CSoutput.n114 5.46119
R6231 CSoutput.n359 CSoutput.n358 5.25266
R6232 CSoutput.n339 CSoutput.n338 5.25266
R6233 CSoutput.n419 CSoutput.n418 5.25266
R6234 CSoutput.n399 CSoutput.n398 5.25266
R6235 CSoutput.n299 CSoutput.n298 5.1449
R6236 CSoutput.n287 CSoutput.n286 5.1449
R6237 CSoutput.n113 CSoutput.n112 5.1449
R6238 CSoutput.n101 CSoutput.n100 5.1449
R6239 CSoutput.n205 CSoutput.n158 4.5005
R6240 CSoutput.n174 CSoutput.n158 4.5005
R6241 CSoutput.n169 CSoutput.n153 4.5005
R6242 CSoutput.n169 CSoutput.n155 4.5005
R6243 CSoutput.n169 CSoutput.n152 4.5005
R6244 CSoutput.n169 CSoutput.n156 4.5005
R6245 CSoutput.n169 CSoutput.n151 4.5005
R6246 CSoutput.n169 CSoutput.t213 4.5005
R6247 CSoutput.n169 CSoutput.n150 4.5005
R6248 CSoutput.n169 CSoutput.n157 4.5005
R6249 CSoutput.n169 CSoutput.n158 4.5005
R6250 CSoutput.n167 CSoutput.n153 4.5005
R6251 CSoutput.n167 CSoutput.n155 4.5005
R6252 CSoutput.n167 CSoutput.n152 4.5005
R6253 CSoutput.n167 CSoutput.n156 4.5005
R6254 CSoutput.n167 CSoutput.n151 4.5005
R6255 CSoutput.n167 CSoutput.t213 4.5005
R6256 CSoutput.n167 CSoutput.n150 4.5005
R6257 CSoutput.n167 CSoutput.n157 4.5005
R6258 CSoutput.n167 CSoutput.n158 4.5005
R6259 CSoutput.n166 CSoutput.n153 4.5005
R6260 CSoutput.n166 CSoutput.n155 4.5005
R6261 CSoutput.n166 CSoutput.n152 4.5005
R6262 CSoutput.n166 CSoutput.n156 4.5005
R6263 CSoutput.n166 CSoutput.n151 4.5005
R6264 CSoutput.n166 CSoutput.t213 4.5005
R6265 CSoutput.n166 CSoutput.n150 4.5005
R6266 CSoutput.n166 CSoutput.n157 4.5005
R6267 CSoutput.n166 CSoutput.n158 4.5005
R6268 CSoutput.n251 CSoutput.n153 4.5005
R6269 CSoutput.n251 CSoutput.n155 4.5005
R6270 CSoutput.n251 CSoutput.n152 4.5005
R6271 CSoutput.n251 CSoutput.n156 4.5005
R6272 CSoutput.n251 CSoutput.n151 4.5005
R6273 CSoutput.n251 CSoutput.t213 4.5005
R6274 CSoutput.n251 CSoutput.n150 4.5005
R6275 CSoutput.n251 CSoutput.n157 4.5005
R6276 CSoutput.n251 CSoutput.n158 4.5005
R6277 CSoutput.n249 CSoutput.n153 4.5005
R6278 CSoutput.n249 CSoutput.n155 4.5005
R6279 CSoutput.n249 CSoutput.n152 4.5005
R6280 CSoutput.n249 CSoutput.n156 4.5005
R6281 CSoutput.n249 CSoutput.n151 4.5005
R6282 CSoutput.n249 CSoutput.t213 4.5005
R6283 CSoutput.n249 CSoutput.n150 4.5005
R6284 CSoutput.n249 CSoutput.n157 4.5005
R6285 CSoutput.n247 CSoutput.n153 4.5005
R6286 CSoutput.n247 CSoutput.n155 4.5005
R6287 CSoutput.n247 CSoutput.n152 4.5005
R6288 CSoutput.n247 CSoutput.n156 4.5005
R6289 CSoutput.n247 CSoutput.n151 4.5005
R6290 CSoutput.n247 CSoutput.t213 4.5005
R6291 CSoutput.n247 CSoutput.n150 4.5005
R6292 CSoutput.n247 CSoutput.n157 4.5005
R6293 CSoutput.n177 CSoutput.n153 4.5005
R6294 CSoutput.n177 CSoutput.n155 4.5005
R6295 CSoutput.n177 CSoutput.n152 4.5005
R6296 CSoutput.n177 CSoutput.n156 4.5005
R6297 CSoutput.n177 CSoutput.n151 4.5005
R6298 CSoutput.n177 CSoutput.t213 4.5005
R6299 CSoutput.n177 CSoutput.n150 4.5005
R6300 CSoutput.n177 CSoutput.n157 4.5005
R6301 CSoutput.n177 CSoutput.n158 4.5005
R6302 CSoutput.n176 CSoutput.n153 4.5005
R6303 CSoutput.n176 CSoutput.n155 4.5005
R6304 CSoutput.n176 CSoutput.n152 4.5005
R6305 CSoutput.n176 CSoutput.n156 4.5005
R6306 CSoutput.n176 CSoutput.n151 4.5005
R6307 CSoutput.n176 CSoutput.t213 4.5005
R6308 CSoutput.n176 CSoutput.n150 4.5005
R6309 CSoutput.n176 CSoutput.n157 4.5005
R6310 CSoutput.n176 CSoutput.n158 4.5005
R6311 CSoutput.n180 CSoutput.n153 4.5005
R6312 CSoutput.n180 CSoutput.n155 4.5005
R6313 CSoutput.n180 CSoutput.n152 4.5005
R6314 CSoutput.n180 CSoutput.n156 4.5005
R6315 CSoutput.n180 CSoutput.n151 4.5005
R6316 CSoutput.n180 CSoutput.t213 4.5005
R6317 CSoutput.n180 CSoutput.n150 4.5005
R6318 CSoutput.n180 CSoutput.n157 4.5005
R6319 CSoutput.n180 CSoutput.n158 4.5005
R6320 CSoutput.n179 CSoutput.n153 4.5005
R6321 CSoutput.n179 CSoutput.n155 4.5005
R6322 CSoutput.n179 CSoutput.n152 4.5005
R6323 CSoutput.n179 CSoutput.n156 4.5005
R6324 CSoutput.n179 CSoutput.n151 4.5005
R6325 CSoutput.n179 CSoutput.t213 4.5005
R6326 CSoutput.n179 CSoutput.n150 4.5005
R6327 CSoutput.n179 CSoutput.n157 4.5005
R6328 CSoutput.n179 CSoutput.n158 4.5005
R6329 CSoutput.n162 CSoutput.n153 4.5005
R6330 CSoutput.n162 CSoutput.n155 4.5005
R6331 CSoutput.n162 CSoutput.n152 4.5005
R6332 CSoutput.n162 CSoutput.n156 4.5005
R6333 CSoutput.n162 CSoutput.n151 4.5005
R6334 CSoutput.n162 CSoutput.t213 4.5005
R6335 CSoutput.n162 CSoutput.n150 4.5005
R6336 CSoutput.n162 CSoutput.n157 4.5005
R6337 CSoutput.n162 CSoutput.n158 4.5005
R6338 CSoutput.n254 CSoutput.n153 4.5005
R6339 CSoutput.n254 CSoutput.n155 4.5005
R6340 CSoutput.n254 CSoutput.n152 4.5005
R6341 CSoutput.n254 CSoutput.n156 4.5005
R6342 CSoutput.n254 CSoutput.n151 4.5005
R6343 CSoutput.n254 CSoutput.t213 4.5005
R6344 CSoutput.n254 CSoutput.n150 4.5005
R6345 CSoutput.n254 CSoutput.n157 4.5005
R6346 CSoutput.n254 CSoutput.n158 4.5005
R6347 CSoutput.n241 CSoutput.n212 4.5005
R6348 CSoutput.n241 CSoutput.n218 4.5005
R6349 CSoutput.n199 CSoutput.n188 4.5005
R6350 CSoutput.n199 CSoutput.n190 4.5005
R6351 CSoutput.n199 CSoutput.n187 4.5005
R6352 CSoutput.n199 CSoutput.n191 4.5005
R6353 CSoutput.n199 CSoutput.n186 4.5005
R6354 CSoutput.n199 CSoutput.t208 4.5005
R6355 CSoutput.n199 CSoutput.n185 4.5005
R6356 CSoutput.n199 CSoutput.n192 4.5005
R6357 CSoutput.n241 CSoutput.n199 4.5005
R6358 CSoutput.n220 CSoutput.n188 4.5005
R6359 CSoutput.n220 CSoutput.n190 4.5005
R6360 CSoutput.n220 CSoutput.n187 4.5005
R6361 CSoutput.n220 CSoutput.n191 4.5005
R6362 CSoutput.n220 CSoutput.n186 4.5005
R6363 CSoutput.n220 CSoutput.t208 4.5005
R6364 CSoutput.n220 CSoutput.n185 4.5005
R6365 CSoutput.n220 CSoutput.n192 4.5005
R6366 CSoutput.n241 CSoutput.n220 4.5005
R6367 CSoutput.n198 CSoutput.n188 4.5005
R6368 CSoutput.n198 CSoutput.n190 4.5005
R6369 CSoutput.n198 CSoutput.n187 4.5005
R6370 CSoutput.n198 CSoutput.n191 4.5005
R6371 CSoutput.n198 CSoutput.n186 4.5005
R6372 CSoutput.n198 CSoutput.t208 4.5005
R6373 CSoutput.n198 CSoutput.n185 4.5005
R6374 CSoutput.n198 CSoutput.n192 4.5005
R6375 CSoutput.n241 CSoutput.n198 4.5005
R6376 CSoutput.n222 CSoutput.n188 4.5005
R6377 CSoutput.n222 CSoutput.n190 4.5005
R6378 CSoutput.n222 CSoutput.n187 4.5005
R6379 CSoutput.n222 CSoutput.n191 4.5005
R6380 CSoutput.n222 CSoutput.n186 4.5005
R6381 CSoutput.n222 CSoutput.t208 4.5005
R6382 CSoutput.n222 CSoutput.n185 4.5005
R6383 CSoutput.n222 CSoutput.n192 4.5005
R6384 CSoutput.n241 CSoutput.n222 4.5005
R6385 CSoutput.n188 CSoutput.n183 4.5005
R6386 CSoutput.n190 CSoutput.n183 4.5005
R6387 CSoutput.n187 CSoutput.n183 4.5005
R6388 CSoutput.n191 CSoutput.n183 4.5005
R6389 CSoutput.n186 CSoutput.n183 4.5005
R6390 CSoutput.t208 CSoutput.n183 4.5005
R6391 CSoutput.n185 CSoutput.n183 4.5005
R6392 CSoutput.n192 CSoutput.n183 4.5005
R6393 CSoutput.n244 CSoutput.n188 4.5005
R6394 CSoutput.n244 CSoutput.n190 4.5005
R6395 CSoutput.n244 CSoutput.n187 4.5005
R6396 CSoutput.n244 CSoutput.n191 4.5005
R6397 CSoutput.n244 CSoutput.n186 4.5005
R6398 CSoutput.n244 CSoutput.t208 4.5005
R6399 CSoutput.n244 CSoutput.n185 4.5005
R6400 CSoutput.n244 CSoutput.n192 4.5005
R6401 CSoutput.n242 CSoutput.n188 4.5005
R6402 CSoutput.n242 CSoutput.n190 4.5005
R6403 CSoutput.n242 CSoutput.n187 4.5005
R6404 CSoutput.n242 CSoutput.n191 4.5005
R6405 CSoutput.n242 CSoutput.n186 4.5005
R6406 CSoutput.n242 CSoutput.t208 4.5005
R6407 CSoutput.n242 CSoutput.n185 4.5005
R6408 CSoutput.n242 CSoutput.n192 4.5005
R6409 CSoutput.n242 CSoutput.n241 4.5005
R6410 CSoutput.n224 CSoutput.n188 4.5005
R6411 CSoutput.n224 CSoutput.n190 4.5005
R6412 CSoutput.n224 CSoutput.n187 4.5005
R6413 CSoutput.n224 CSoutput.n191 4.5005
R6414 CSoutput.n224 CSoutput.n186 4.5005
R6415 CSoutput.n224 CSoutput.t208 4.5005
R6416 CSoutput.n224 CSoutput.n185 4.5005
R6417 CSoutput.n224 CSoutput.n192 4.5005
R6418 CSoutput.n241 CSoutput.n224 4.5005
R6419 CSoutput.n196 CSoutput.n188 4.5005
R6420 CSoutput.n196 CSoutput.n190 4.5005
R6421 CSoutput.n196 CSoutput.n187 4.5005
R6422 CSoutput.n196 CSoutput.n191 4.5005
R6423 CSoutput.n196 CSoutput.n186 4.5005
R6424 CSoutput.n196 CSoutput.t208 4.5005
R6425 CSoutput.n196 CSoutput.n185 4.5005
R6426 CSoutput.n196 CSoutput.n192 4.5005
R6427 CSoutput.n241 CSoutput.n196 4.5005
R6428 CSoutput.n226 CSoutput.n188 4.5005
R6429 CSoutput.n226 CSoutput.n190 4.5005
R6430 CSoutput.n226 CSoutput.n187 4.5005
R6431 CSoutput.n226 CSoutput.n191 4.5005
R6432 CSoutput.n226 CSoutput.n186 4.5005
R6433 CSoutput.n226 CSoutput.t208 4.5005
R6434 CSoutput.n226 CSoutput.n185 4.5005
R6435 CSoutput.n226 CSoutput.n192 4.5005
R6436 CSoutput.n241 CSoutput.n226 4.5005
R6437 CSoutput.n195 CSoutput.n188 4.5005
R6438 CSoutput.n195 CSoutput.n190 4.5005
R6439 CSoutput.n195 CSoutput.n187 4.5005
R6440 CSoutput.n195 CSoutput.n191 4.5005
R6441 CSoutput.n195 CSoutput.n186 4.5005
R6442 CSoutput.n195 CSoutput.t208 4.5005
R6443 CSoutput.n195 CSoutput.n185 4.5005
R6444 CSoutput.n195 CSoutput.n192 4.5005
R6445 CSoutput.n241 CSoutput.n195 4.5005
R6446 CSoutput.n240 CSoutput.n188 4.5005
R6447 CSoutput.n240 CSoutput.n190 4.5005
R6448 CSoutput.n240 CSoutput.n187 4.5005
R6449 CSoutput.n240 CSoutput.n191 4.5005
R6450 CSoutput.n240 CSoutput.n186 4.5005
R6451 CSoutput.n240 CSoutput.t208 4.5005
R6452 CSoutput.n240 CSoutput.n185 4.5005
R6453 CSoutput.n240 CSoutput.n192 4.5005
R6454 CSoutput.n241 CSoutput.n240 4.5005
R6455 CSoutput.n239 CSoutput.n124 4.5005
R6456 CSoutput.n140 CSoutput.n124 4.5005
R6457 CSoutput.n135 CSoutput.n119 4.5005
R6458 CSoutput.n135 CSoutput.n121 4.5005
R6459 CSoutput.n135 CSoutput.n118 4.5005
R6460 CSoutput.n135 CSoutput.n122 4.5005
R6461 CSoutput.n135 CSoutput.n117 4.5005
R6462 CSoutput.n135 CSoutput.t206 4.5005
R6463 CSoutput.n135 CSoutput.n116 4.5005
R6464 CSoutput.n135 CSoutput.n123 4.5005
R6465 CSoutput.n135 CSoutput.n124 4.5005
R6466 CSoutput.n133 CSoutput.n119 4.5005
R6467 CSoutput.n133 CSoutput.n121 4.5005
R6468 CSoutput.n133 CSoutput.n118 4.5005
R6469 CSoutput.n133 CSoutput.n122 4.5005
R6470 CSoutput.n133 CSoutput.n117 4.5005
R6471 CSoutput.n133 CSoutput.t206 4.5005
R6472 CSoutput.n133 CSoutput.n116 4.5005
R6473 CSoutput.n133 CSoutput.n123 4.5005
R6474 CSoutput.n133 CSoutput.n124 4.5005
R6475 CSoutput.n132 CSoutput.n119 4.5005
R6476 CSoutput.n132 CSoutput.n121 4.5005
R6477 CSoutput.n132 CSoutput.n118 4.5005
R6478 CSoutput.n132 CSoutput.n122 4.5005
R6479 CSoutput.n132 CSoutput.n117 4.5005
R6480 CSoutput.n132 CSoutput.t206 4.5005
R6481 CSoutput.n132 CSoutput.n116 4.5005
R6482 CSoutput.n132 CSoutput.n123 4.5005
R6483 CSoutput.n132 CSoutput.n124 4.5005
R6484 CSoutput.n261 CSoutput.n119 4.5005
R6485 CSoutput.n261 CSoutput.n121 4.5005
R6486 CSoutput.n261 CSoutput.n118 4.5005
R6487 CSoutput.n261 CSoutput.n122 4.5005
R6488 CSoutput.n261 CSoutput.n117 4.5005
R6489 CSoutput.n261 CSoutput.t206 4.5005
R6490 CSoutput.n261 CSoutput.n116 4.5005
R6491 CSoutput.n261 CSoutput.n123 4.5005
R6492 CSoutput.n261 CSoutput.n124 4.5005
R6493 CSoutput.n259 CSoutput.n119 4.5005
R6494 CSoutput.n259 CSoutput.n121 4.5005
R6495 CSoutput.n259 CSoutput.n118 4.5005
R6496 CSoutput.n259 CSoutput.n122 4.5005
R6497 CSoutput.n259 CSoutput.n117 4.5005
R6498 CSoutput.n259 CSoutput.t206 4.5005
R6499 CSoutput.n259 CSoutput.n116 4.5005
R6500 CSoutput.n259 CSoutput.n123 4.5005
R6501 CSoutput.n257 CSoutput.n119 4.5005
R6502 CSoutput.n257 CSoutput.n121 4.5005
R6503 CSoutput.n257 CSoutput.n118 4.5005
R6504 CSoutput.n257 CSoutput.n122 4.5005
R6505 CSoutput.n257 CSoutput.n117 4.5005
R6506 CSoutput.n257 CSoutput.t206 4.5005
R6507 CSoutput.n257 CSoutput.n116 4.5005
R6508 CSoutput.n257 CSoutput.n123 4.5005
R6509 CSoutput.n143 CSoutput.n119 4.5005
R6510 CSoutput.n143 CSoutput.n121 4.5005
R6511 CSoutput.n143 CSoutput.n118 4.5005
R6512 CSoutput.n143 CSoutput.n122 4.5005
R6513 CSoutput.n143 CSoutput.n117 4.5005
R6514 CSoutput.n143 CSoutput.t206 4.5005
R6515 CSoutput.n143 CSoutput.n116 4.5005
R6516 CSoutput.n143 CSoutput.n123 4.5005
R6517 CSoutput.n143 CSoutput.n124 4.5005
R6518 CSoutput.n142 CSoutput.n119 4.5005
R6519 CSoutput.n142 CSoutput.n121 4.5005
R6520 CSoutput.n142 CSoutput.n118 4.5005
R6521 CSoutput.n142 CSoutput.n122 4.5005
R6522 CSoutput.n142 CSoutput.n117 4.5005
R6523 CSoutput.n142 CSoutput.t206 4.5005
R6524 CSoutput.n142 CSoutput.n116 4.5005
R6525 CSoutput.n142 CSoutput.n123 4.5005
R6526 CSoutput.n142 CSoutput.n124 4.5005
R6527 CSoutput.n146 CSoutput.n119 4.5005
R6528 CSoutput.n146 CSoutput.n121 4.5005
R6529 CSoutput.n146 CSoutput.n118 4.5005
R6530 CSoutput.n146 CSoutput.n122 4.5005
R6531 CSoutput.n146 CSoutput.n117 4.5005
R6532 CSoutput.n146 CSoutput.t206 4.5005
R6533 CSoutput.n146 CSoutput.n116 4.5005
R6534 CSoutput.n146 CSoutput.n123 4.5005
R6535 CSoutput.n146 CSoutput.n124 4.5005
R6536 CSoutput.n145 CSoutput.n119 4.5005
R6537 CSoutput.n145 CSoutput.n121 4.5005
R6538 CSoutput.n145 CSoutput.n118 4.5005
R6539 CSoutput.n145 CSoutput.n122 4.5005
R6540 CSoutput.n145 CSoutput.n117 4.5005
R6541 CSoutput.n145 CSoutput.t206 4.5005
R6542 CSoutput.n145 CSoutput.n116 4.5005
R6543 CSoutput.n145 CSoutput.n123 4.5005
R6544 CSoutput.n145 CSoutput.n124 4.5005
R6545 CSoutput.n128 CSoutput.n119 4.5005
R6546 CSoutput.n128 CSoutput.n121 4.5005
R6547 CSoutput.n128 CSoutput.n118 4.5005
R6548 CSoutput.n128 CSoutput.n122 4.5005
R6549 CSoutput.n128 CSoutput.n117 4.5005
R6550 CSoutput.n128 CSoutput.t206 4.5005
R6551 CSoutput.n128 CSoutput.n116 4.5005
R6552 CSoutput.n128 CSoutput.n123 4.5005
R6553 CSoutput.n128 CSoutput.n124 4.5005
R6554 CSoutput.n264 CSoutput.n119 4.5005
R6555 CSoutput.n264 CSoutput.n121 4.5005
R6556 CSoutput.n264 CSoutput.n118 4.5005
R6557 CSoutput.n264 CSoutput.n122 4.5005
R6558 CSoutput.n264 CSoutput.n117 4.5005
R6559 CSoutput.n264 CSoutput.t206 4.5005
R6560 CSoutput.n264 CSoutput.n116 4.5005
R6561 CSoutput.n264 CSoutput.n123 4.5005
R6562 CSoutput.n264 CSoutput.n124 4.5005
R6563 CSoutput.n299 CSoutput.n287 4.10845
R6564 CSoutput.n113 CSoutput.n101 4.10845
R6565 CSoutput.n297 CSoutput.t101 4.06363
R6566 CSoutput.n297 CSoutput.t144 4.06363
R6567 CSoutput.n295 CSoutput.t154 4.06363
R6568 CSoutput.n295 CSoutput.t155 4.06363
R6569 CSoutput.n293 CSoutput.t114 4.06363
R6570 CSoutput.n293 CSoutput.t115 4.06363
R6571 CSoutput.n291 CSoutput.t120 4.06363
R6572 CSoutput.n291 CSoutput.t156 4.06363
R6573 CSoutput.n289 CSoutput.t95 4.06363
R6574 CSoutput.n289 CSoutput.t118 4.06363
R6575 CSoutput.n288 CSoutput.t128 4.06363
R6576 CSoutput.n288 CSoutput.t140 4.06363
R6577 CSoutput.n285 CSoutput.t92 4.06363
R6578 CSoutput.n285 CSoutput.t135 4.06363
R6579 CSoutput.n283 CSoutput.t147 4.06363
R6580 CSoutput.n283 CSoutput.t148 4.06363
R6581 CSoutput.n281 CSoutput.t105 4.06363
R6582 CSoutput.n281 CSoutput.t106 4.06363
R6583 CSoutput.n279 CSoutput.t109 4.06363
R6584 CSoutput.n279 CSoutput.t149 4.06363
R6585 CSoutput.n277 CSoutput.t87 4.06363
R6586 CSoutput.n277 CSoutput.t108 4.06363
R6587 CSoutput.n276 CSoutput.t121 4.06363
R6588 CSoutput.n276 CSoutput.t134 4.06363
R6589 CSoutput.n274 CSoutput.t145 4.06363
R6590 CSoutput.n274 CSoutput.t96 4.06363
R6591 CSoutput.n272 CSoutput.t122 4.06363
R6592 CSoutput.n272 CSoutput.t107 4.06363
R6593 CSoutput.n270 CSoutput.t110 4.06363
R6594 CSoutput.n270 CSoutput.t93 4.06363
R6595 CSoutput.n268 CSoutput.t139 4.06363
R6596 CSoutput.n268 CSoutput.t89 4.06363
R6597 CSoutput.n266 CSoutput.t116 4.06363
R6598 CSoutput.n266 CSoutput.t152 4.06363
R6599 CSoutput.n265 CSoutput.t102 4.06363
R6600 CSoutput.n265 CSoutput.t142 4.06363
R6601 CSoutput.n102 CSoutput.t98 4.06363
R6602 CSoutput.n102 CSoutput.t150 4.06363
R6603 CSoutput.n103 CSoutput.t138 4.06363
R6604 CSoutput.n103 CSoutput.t126 4.06363
R6605 CSoutput.n105 CSoutput.t113 4.06363
R6606 CSoutput.n105 CSoutput.t158 4.06363
R6607 CSoutput.n107 CSoutput.t137 4.06363
R6608 CSoutput.n107 CSoutput.t136 4.06363
R6609 CSoutput.n109 CSoutput.t129 4.06363
R6610 CSoutput.n109 CSoutput.t112 4.06363
R6611 CSoutput.n111 CSoutput.t99 4.06363
R6612 CSoutput.n111 CSoutput.t130 4.06363
R6613 CSoutput.n90 CSoutput.t88 4.06363
R6614 CSoutput.n90 CSoutput.t141 4.06363
R6615 CSoutput.n91 CSoutput.t133 4.06363
R6616 CSoutput.n91 CSoutput.t119 4.06363
R6617 CSoutput.n93 CSoutput.t104 4.06363
R6618 CSoutput.n93 CSoutput.t151 4.06363
R6619 CSoutput.n95 CSoutput.t132 4.06363
R6620 CSoutput.n95 CSoutput.t131 4.06363
R6621 CSoutput.n97 CSoutput.t124 4.06363
R6622 CSoutput.n97 CSoutput.t100 4.06363
R6623 CSoutput.n99 CSoutput.t90 4.06363
R6624 CSoutput.n99 CSoutput.t125 4.06363
R6625 CSoutput.n79 CSoutput.t143 4.06363
R6626 CSoutput.n79 CSoutput.t103 4.06363
R6627 CSoutput.n80 CSoutput.t153 4.06363
R6628 CSoutput.n80 CSoutput.t117 4.06363
R6629 CSoutput.n82 CSoutput.t91 4.06363
R6630 CSoutput.n82 CSoutput.t127 4.06363
R6631 CSoutput.n84 CSoutput.t94 4.06363
R6632 CSoutput.n84 CSoutput.t111 4.06363
R6633 CSoutput.n86 CSoutput.t157 4.06363
R6634 CSoutput.n86 CSoutput.t123 4.06363
R6635 CSoutput.n88 CSoutput.t97 4.06363
R6636 CSoutput.n88 CSoutput.t146 4.06363
R6637 CSoutput.n44 CSoutput.n43 3.79402
R6638 CSoutput.n49 CSoutput.n48 3.79402
R6639 CSoutput.n359 CSoutput.n339 3.72967
R6640 CSoutput.n419 CSoutput.n399 3.72967
R6641 CSoutput.n421 CSoutput.n420 3.57343
R6642 CSoutput.n420 CSoutput.n360 3.42304
R6643 CSoutput.n357 CSoutput.t30 2.82907
R6644 CSoutput.n357 CSoutput.t61 2.82907
R6645 CSoutput.n355 CSoutput.t49 2.82907
R6646 CSoutput.n355 CSoutput.t19 2.82907
R6647 CSoutput.n353 CSoutput.t54 2.82907
R6648 CSoutput.n353 CSoutput.t77 2.82907
R6649 CSoutput.n351 CSoutput.t184 2.82907
R6650 CSoutput.n351 CSoutput.t72 2.82907
R6651 CSoutput.n349 CSoutput.t52 2.82907
R6652 CSoutput.n349 CSoutput.t53 2.82907
R6653 CSoutput.n347 CSoutput.t18 2.82907
R6654 CSoutput.n347 CSoutput.t39 2.82907
R6655 CSoutput.n345 CSoutput.t79 2.82907
R6656 CSoutput.n345 CSoutput.t76 2.82907
R6657 CSoutput.n343 CSoutput.t50 2.82907
R6658 CSoutput.n343 CSoutput.t71 2.82907
R6659 CSoutput.n341 CSoutput.t173 2.82907
R6660 CSoutput.n341 CSoutput.t44 2.82907
R6661 CSoutput.n340 CSoutput.t21 2.82907
R6662 CSoutput.n340 CSoutput.t73 2.82907
R6663 CSoutput.n337 CSoutput.t33 2.82907
R6664 CSoutput.n337 CSoutput.t83 2.82907
R6665 CSoutput.n335 CSoutput.t160 2.82907
R6666 CSoutput.n335 CSoutput.t181 2.82907
R6667 CSoutput.n333 CSoutput.t163 2.82907
R6668 CSoutput.n333 CSoutput.t36 2.82907
R6669 CSoutput.n331 CSoutput.t67 2.82907
R6670 CSoutput.n331 CSoutput.t10 2.82907
R6671 CSoutput.n329 CSoutput.t80 2.82907
R6672 CSoutput.n329 CSoutput.t70 2.82907
R6673 CSoutput.n327 CSoutput.t24 2.82907
R6674 CSoutput.n327 CSoutput.t159 2.82907
R6675 CSoutput.n325 CSoutput.t189 2.82907
R6676 CSoutput.n325 CSoutput.t168 2.82907
R6677 CSoutput.n323 CSoutput.t75 2.82907
R6678 CSoutput.n323 CSoutput.t13 2.82907
R6679 CSoutput.n321 CSoutput.t170 2.82907
R6680 CSoutput.n321 CSoutput.t59 2.82907
R6681 CSoutput.n320 CSoutput.t86 2.82907
R6682 CSoutput.n320 CSoutput.t183 2.82907
R6683 CSoutput.n318 CSoutput.t15 2.82907
R6684 CSoutput.n318 CSoutput.t161 2.82907
R6685 CSoutput.n316 CSoutput.t12 2.82907
R6686 CSoutput.n316 CSoutput.t176 2.82907
R6687 CSoutput.n314 CSoutput.t34 2.82907
R6688 CSoutput.n314 CSoutput.t186 2.82907
R6689 CSoutput.n312 CSoutput.t179 2.82907
R6690 CSoutput.n312 CSoutput.t82 2.82907
R6691 CSoutput.n310 CSoutput.t23 2.82907
R6692 CSoutput.n310 CSoutput.t84 2.82907
R6693 CSoutput.n308 CSoutput.t167 2.82907
R6694 CSoutput.n308 CSoutput.t178 2.82907
R6695 CSoutput.n306 CSoutput.t174 2.82907
R6696 CSoutput.n306 CSoutput.t166 2.82907
R6697 CSoutput.n304 CSoutput.t5 2.82907
R6698 CSoutput.n304 CSoutput.t17 2.82907
R6699 CSoutput.n302 CSoutput.t190 2.82907
R6700 CSoutput.n302 CSoutput.t28 2.82907
R6701 CSoutput.n301 CSoutput.t191 2.82907
R6702 CSoutput.n301 CSoutput.t165 2.82907
R6703 CSoutput.n400 CSoutput.t55 2.82907
R6704 CSoutput.n400 CSoutput.t182 2.82907
R6705 CSoutput.n401 CSoutput.t171 2.82907
R6706 CSoutput.n401 CSoutput.t8 2.82907
R6707 CSoutput.n403 CSoutput.t62 2.82907
R6708 CSoutput.n403 CSoutput.t11 2.82907
R6709 CSoutput.n405 CSoutput.t58 2.82907
R6710 CSoutput.n405 CSoutput.t0 2.82907
R6711 CSoutput.n407 CSoutput.t45 2.82907
R6712 CSoutput.n407 CSoutput.t60 2.82907
R6713 CSoutput.n409 CSoutput.t169 2.82907
R6714 CSoutput.n409 CSoutput.t185 2.82907
R6715 CSoutput.n411 CSoutput.t9 2.82907
R6716 CSoutput.n411 CSoutput.t65 2.82907
R6717 CSoutput.n413 CSoutput.t2 2.82907
R6718 CSoutput.n413 CSoutput.t27 2.82907
R6719 CSoutput.n415 CSoutput.t180 2.82907
R6720 CSoutput.n415 CSoutput.t37 2.82907
R6721 CSoutput.n417 CSoutput.t20 2.82907
R6722 CSoutput.n417 CSoutput.t40 2.82907
R6723 CSoutput.n380 CSoutput.t29 2.82907
R6724 CSoutput.n380 CSoutput.t31 2.82907
R6725 CSoutput.n381 CSoutput.t3 2.82907
R6726 CSoutput.n381 CSoutput.t47 2.82907
R6727 CSoutput.n383 CSoutput.t41 2.82907
R6728 CSoutput.n383 CSoutput.t42 2.82907
R6729 CSoutput.n385 CSoutput.t35 2.82907
R6730 CSoutput.n385 CSoutput.t69 2.82907
R6731 CSoutput.n387 CSoutput.t56 2.82907
R6732 CSoutput.n387 CSoutput.t74 2.82907
R6733 CSoutput.n389 CSoutput.t66 2.82907
R6734 CSoutput.n389 CSoutput.t177 2.82907
R6735 CSoutput.n391 CSoutput.t25 2.82907
R6736 CSoutput.n391 CSoutput.t187 2.82907
R6737 CSoutput.n393 CSoutput.t175 2.82907
R6738 CSoutput.n393 CSoutput.t26 2.82907
R6739 CSoutput.n395 CSoutput.t63 2.82907
R6740 CSoutput.n395 CSoutput.t164 2.82907
R6741 CSoutput.n397 CSoutput.t188 2.82907
R6742 CSoutput.n397 CSoutput.t48 2.82907
R6743 CSoutput.n361 CSoutput.t43 2.82907
R6744 CSoutput.n361 CSoutput.t1 2.82907
R6745 CSoutput.n362 CSoutput.t64 2.82907
R6746 CSoutput.n362 CSoutput.t22 2.82907
R6747 CSoutput.n364 CSoutput.t57 2.82907
R6748 CSoutput.n364 CSoutput.t7 2.82907
R6749 CSoutput.n366 CSoutput.t162 2.82907
R6750 CSoutput.n366 CSoutput.t14 2.82907
R6751 CSoutput.n368 CSoutput.t4 2.82907
R6752 CSoutput.n368 CSoutput.t85 2.82907
R6753 CSoutput.n370 CSoutput.t51 2.82907
R6754 CSoutput.n370 CSoutput.t38 2.82907
R6755 CSoutput.n372 CSoutput.t46 2.82907
R6756 CSoutput.n372 CSoutput.t16 2.82907
R6757 CSoutput.n374 CSoutput.t68 2.82907
R6758 CSoutput.n374 CSoutput.t172 2.82907
R6759 CSoutput.n376 CSoutput.t78 2.82907
R6760 CSoutput.n376 CSoutput.t81 2.82907
R6761 CSoutput.n378 CSoutput.t32 2.82907
R6762 CSoutput.n378 CSoutput.t6 2.82907
R6763 CSoutput.n75 CSoutput.n1 2.45513
R6764 CSoutput.n300 CSoutput.n114 2.36742
R6765 CSoutput.n205 CSoutput.n203 2.251
R6766 CSoutput.n205 CSoutput.n202 2.251
R6767 CSoutput.n205 CSoutput.n201 2.251
R6768 CSoutput.n205 CSoutput.n200 2.251
R6769 CSoutput.n174 CSoutput.n173 2.251
R6770 CSoutput.n174 CSoutput.n172 2.251
R6771 CSoutput.n174 CSoutput.n171 2.251
R6772 CSoutput.n174 CSoutput.n170 2.251
R6773 CSoutput.n247 CSoutput.n246 2.251
R6774 CSoutput.n212 CSoutput.n210 2.251
R6775 CSoutput.n212 CSoutput.n209 2.251
R6776 CSoutput.n212 CSoutput.n208 2.251
R6777 CSoutput.n230 CSoutput.n212 2.251
R6778 CSoutput.n218 CSoutput.n217 2.251
R6779 CSoutput.n218 CSoutput.n216 2.251
R6780 CSoutput.n218 CSoutput.n215 2.251
R6781 CSoutput.n218 CSoutput.n214 2.251
R6782 CSoutput.n244 CSoutput.n184 2.251
R6783 CSoutput.n239 CSoutput.n237 2.251
R6784 CSoutput.n239 CSoutput.n236 2.251
R6785 CSoutput.n239 CSoutput.n235 2.251
R6786 CSoutput.n239 CSoutput.n234 2.251
R6787 CSoutput.n140 CSoutput.n139 2.251
R6788 CSoutput.n140 CSoutput.n138 2.251
R6789 CSoutput.n140 CSoutput.n137 2.251
R6790 CSoutput.n140 CSoutput.n136 2.251
R6791 CSoutput.n257 CSoutput.n256 2.251
R6792 CSoutput.n174 CSoutput.n154 2.2505
R6793 CSoutput.n169 CSoutput.n154 2.2505
R6794 CSoutput.n167 CSoutput.n154 2.2505
R6795 CSoutput.n166 CSoutput.n154 2.2505
R6796 CSoutput.n251 CSoutput.n154 2.2505
R6797 CSoutput.n249 CSoutput.n154 2.2505
R6798 CSoutput.n247 CSoutput.n154 2.2505
R6799 CSoutput.n177 CSoutput.n154 2.2505
R6800 CSoutput.n176 CSoutput.n154 2.2505
R6801 CSoutput.n180 CSoutput.n154 2.2505
R6802 CSoutput.n179 CSoutput.n154 2.2505
R6803 CSoutput.n162 CSoutput.n154 2.2505
R6804 CSoutput.n254 CSoutput.n154 2.2505
R6805 CSoutput.n254 CSoutput.n253 2.2505
R6806 CSoutput.n218 CSoutput.n189 2.2505
R6807 CSoutput.n199 CSoutput.n189 2.2505
R6808 CSoutput.n220 CSoutput.n189 2.2505
R6809 CSoutput.n198 CSoutput.n189 2.2505
R6810 CSoutput.n222 CSoutput.n189 2.2505
R6811 CSoutput.n189 CSoutput.n183 2.2505
R6812 CSoutput.n244 CSoutput.n189 2.2505
R6813 CSoutput.n242 CSoutput.n189 2.2505
R6814 CSoutput.n224 CSoutput.n189 2.2505
R6815 CSoutput.n196 CSoutput.n189 2.2505
R6816 CSoutput.n226 CSoutput.n189 2.2505
R6817 CSoutput.n195 CSoutput.n189 2.2505
R6818 CSoutput.n240 CSoutput.n189 2.2505
R6819 CSoutput.n240 CSoutput.n193 2.2505
R6820 CSoutput.n140 CSoutput.n120 2.2505
R6821 CSoutput.n135 CSoutput.n120 2.2505
R6822 CSoutput.n133 CSoutput.n120 2.2505
R6823 CSoutput.n132 CSoutput.n120 2.2505
R6824 CSoutput.n261 CSoutput.n120 2.2505
R6825 CSoutput.n259 CSoutput.n120 2.2505
R6826 CSoutput.n257 CSoutput.n120 2.2505
R6827 CSoutput.n143 CSoutput.n120 2.2505
R6828 CSoutput.n142 CSoutput.n120 2.2505
R6829 CSoutput.n146 CSoutput.n120 2.2505
R6830 CSoutput.n145 CSoutput.n120 2.2505
R6831 CSoutput.n128 CSoutput.n120 2.2505
R6832 CSoutput.n264 CSoutput.n120 2.2505
R6833 CSoutput.n264 CSoutput.n263 2.2505
R6834 CSoutput.n182 CSoutput.n175 2.25024
R6835 CSoutput.n182 CSoutput.n168 2.25024
R6836 CSoutput.n250 CSoutput.n182 2.25024
R6837 CSoutput.n182 CSoutput.n178 2.25024
R6838 CSoutput.n182 CSoutput.n181 2.25024
R6839 CSoutput.n182 CSoutput.n149 2.25024
R6840 CSoutput.n232 CSoutput.n229 2.25024
R6841 CSoutput.n232 CSoutput.n228 2.25024
R6842 CSoutput.n232 CSoutput.n227 2.25024
R6843 CSoutput.n232 CSoutput.n194 2.25024
R6844 CSoutput.n232 CSoutput.n231 2.25024
R6845 CSoutput.n233 CSoutput.n232 2.25024
R6846 CSoutput.n148 CSoutput.n141 2.25024
R6847 CSoutput.n148 CSoutput.n134 2.25024
R6848 CSoutput.n260 CSoutput.n148 2.25024
R6849 CSoutput.n148 CSoutput.n144 2.25024
R6850 CSoutput.n148 CSoutput.n147 2.25024
R6851 CSoutput.n148 CSoutput.n115 2.25024
R6852 CSoutput.n249 CSoutput.n159 1.50111
R6853 CSoutput.n197 CSoutput.n183 1.50111
R6854 CSoutput.n259 CSoutput.n125 1.50111
R6855 CSoutput.n205 CSoutput.n204 1.501
R6856 CSoutput.n212 CSoutput.n211 1.501
R6857 CSoutput.n239 CSoutput.n238 1.501
R6858 CSoutput.n253 CSoutput.n164 1.12536
R6859 CSoutput.n253 CSoutput.n165 1.12536
R6860 CSoutput.n253 CSoutput.n252 1.12536
R6861 CSoutput.n213 CSoutput.n193 1.12536
R6862 CSoutput.n219 CSoutput.n193 1.12536
R6863 CSoutput.n221 CSoutput.n193 1.12536
R6864 CSoutput.n263 CSoutput.n130 1.12536
R6865 CSoutput.n263 CSoutput.n131 1.12536
R6866 CSoutput.n263 CSoutput.n262 1.12536
R6867 CSoutput.n253 CSoutput.n160 1.12536
R6868 CSoutput.n253 CSoutput.n161 1.12536
R6869 CSoutput.n253 CSoutput.n163 1.12536
R6870 CSoutput.n243 CSoutput.n193 1.12536
R6871 CSoutput.n223 CSoutput.n193 1.12536
R6872 CSoutput.n225 CSoutput.n193 1.12536
R6873 CSoutput.n263 CSoutput.n126 1.12536
R6874 CSoutput.n263 CSoutput.n127 1.12536
R6875 CSoutput.n263 CSoutput.n129 1.12536
R6876 CSoutput.n31 CSoutput.n30 0.669944
R6877 CSoutput.n62 CSoutput.n61 0.669944
R6878 CSoutput.n344 CSoutput.n342 0.573776
R6879 CSoutput.n346 CSoutput.n344 0.573776
R6880 CSoutput.n348 CSoutput.n346 0.573776
R6881 CSoutput.n350 CSoutput.n348 0.573776
R6882 CSoutput.n352 CSoutput.n350 0.573776
R6883 CSoutput.n354 CSoutput.n352 0.573776
R6884 CSoutput.n356 CSoutput.n354 0.573776
R6885 CSoutput.n358 CSoutput.n356 0.573776
R6886 CSoutput.n324 CSoutput.n322 0.573776
R6887 CSoutput.n326 CSoutput.n324 0.573776
R6888 CSoutput.n328 CSoutput.n326 0.573776
R6889 CSoutput.n330 CSoutput.n328 0.573776
R6890 CSoutput.n332 CSoutput.n330 0.573776
R6891 CSoutput.n334 CSoutput.n332 0.573776
R6892 CSoutput.n336 CSoutput.n334 0.573776
R6893 CSoutput.n338 CSoutput.n336 0.573776
R6894 CSoutput.n305 CSoutput.n303 0.573776
R6895 CSoutput.n307 CSoutput.n305 0.573776
R6896 CSoutput.n309 CSoutput.n307 0.573776
R6897 CSoutput.n311 CSoutput.n309 0.573776
R6898 CSoutput.n313 CSoutput.n311 0.573776
R6899 CSoutput.n315 CSoutput.n313 0.573776
R6900 CSoutput.n317 CSoutput.n315 0.573776
R6901 CSoutput.n319 CSoutput.n317 0.573776
R6902 CSoutput.n418 CSoutput.n416 0.573776
R6903 CSoutput.n416 CSoutput.n414 0.573776
R6904 CSoutput.n414 CSoutput.n412 0.573776
R6905 CSoutput.n412 CSoutput.n410 0.573776
R6906 CSoutput.n410 CSoutput.n408 0.573776
R6907 CSoutput.n408 CSoutput.n406 0.573776
R6908 CSoutput.n406 CSoutput.n404 0.573776
R6909 CSoutput.n404 CSoutput.n402 0.573776
R6910 CSoutput.n398 CSoutput.n396 0.573776
R6911 CSoutput.n396 CSoutput.n394 0.573776
R6912 CSoutput.n394 CSoutput.n392 0.573776
R6913 CSoutput.n392 CSoutput.n390 0.573776
R6914 CSoutput.n390 CSoutput.n388 0.573776
R6915 CSoutput.n388 CSoutput.n386 0.573776
R6916 CSoutput.n386 CSoutput.n384 0.573776
R6917 CSoutput.n384 CSoutput.n382 0.573776
R6918 CSoutput.n379 CSoutput.n377 0.573776
R6919 CSoutput.n377 CSoutput.n375 0.573776
R6920 CSoutput.n375 CSoutput.n373 0.573776
R6921 CSoutput.n373 CSoutput.n371 0.573776
R6922 CSoutput.n371 CSoutput.n369 0.573776
R6923 CSoutput.n369 CSoutput.n367 0.573776
R6924 CSoutput.n367 CSoutput.n365 0.573776
R6925 CSoutput.n365 CSoutput.n363 0.573776
R6926 CSoutput.n421 CSoutput.n264 0.53442
R6927 CSoutput.n292 CSoutput.n290 0.358259
R6928 CSoutput.n294 CSoutput.n292 0.358259
R6929 CSoutput.n296 CSoutput.n294 0.358259
R6930 CSoutput.n298 CSoutput.n296 0.358259
R6931 CSoutput.n280 CSoutput.n278 0.358259
R6932 CSoutput.n282 CSoutput.n280 0.358259
R6933 CSoutput.n284 CSoutput.n282 0.358259
R6934 CSoutput.n286 CSoutput.n284 0.358259
R6935 CSoutput.n269 CSoutput.n267 0.358259
R6936 CSoutput.n271 CSoutput.n269 0.358259
R6937 CSoutput.n273 CSoutput.n271 0.358259
R6938 CSoutput.n275 CSoutput.n273 0.358259
R6939 CSoutput.n112 CSoutput.n110 0.358259
R6940 CSoutput.n110 CSoutput.n108 0.358259
R6941 CSoutput.n108 CSoutput.n106 0.358259
R6942 CSoutput.n106 CSoutput.n104 0.358259
R6943 CSoutput.n100 CSoutput.n98 0.358259
R6944 CSoutput.n98 CSoutput.n96 0.358259
R6945 CSoutput.n96 CSoutput.n94 0.358259
R6946 CSoutput.n94 CSoutput.n92 0.358259
R6947 CSoutput.n89 CSoutput.n87 0.358259
R6948 CSoutput.n87 CSoutput.n85 0.358259
R6949 CSoutput.n85 CSoutput.n83 0.358259
R6950 CSoutput.n83 CSoutput.n81 0.358259
R6951 CSoutput.n21 CSoutput.n20 0.169105
R6952 CSoutput.n21 CSoutput.n16 0.169105
R6953 CSoutput.n26 CSoutput.n16 0.169105
R6954 CSoutput.n27 CSoutput.n26 0.169105
R6955 CSoutput.n27 CSoutput.n14 0.169105
R6956 CSoutput.n32 CSoutput.n14 0.169105
R6957 CSoutput.n33 CSoutput.n32 0.169105
R6958 CSoutput.n34 CSoutput.n33 0.169105
R6959 CSoutput.n34 CSoutput.n12 0.169105
R6960 CSoutput.n39 CSoutput.n12 0.169105
R6961 CSoutput.n40 CSoutput.n39 0.169105
R6962 CSoutput.n40 CSoutput.n10 0.169105
R6963 CSoutput.n45 CSoutput.n10 0.169105
R6964 CSoutput.n46 CSoutput.n45 0.169105
R6965 CSoutput.n47 CSoutput.n46 0.169105
R6966 CSoutput.n47 CSoutput.n8 0.169105
R6967 CSoutput.n52 CSoutput.n8 0.169105
R6968 CSoutput.n53 CSoutput.n52 0.169105
R6969 CSoutput.n53 CSoutput.n6 0.169105
R6970 CSoutput.n58 CSoutput.n6 0.169105
R6971 CSoutput.n59 CSoutput.n58 0.169105
R6972 CSoutput.n60 CSoutput.n59 0.169105
R6973 CSoutput.n60 CSoutput.n4 0.169105
R6974 CSoutput.n66 CSoutput.n4 0.169105
R6975 CSoutput.n67 CSoutput.n66 0.169105
R6976 CSoutput.n68 CSoutput.n67 0.169105
R6977 CSoutput.n68 CSoutput.n2 0.169105
R6978 CSoutput.n73 CSoutput.n2 0.169105
R6979 CSoutput.n74 CSoutput.n73 0.169105
R6980 CSoutput.n74 CSoutput.n0 0.169105
R6981 CSoutput.n78 CSoutput.n0 0.169105
R6982 CSoutput.n207 CSoutput.n206 0.0910737
R6983 CSoutput.n258 CSoutput.n255 0.0723685
R6984 CSoutput.n212 CSoutput.n207 0.0522944
R6985 CSoutput.n255 CSoutput.n254 0.0499135
R6986 CSoutput.n206 CSoutput.n205 0.0499135
R6987 CSoutput.n240 CSoutput.n239 0.0464294
R6988 CSoutput.n248 CSoutput.n245 0.0391444
R6989 CSoutput.n207 CSoutput.t192 0.023435
R6990 CSoutput.n255 CSoutput.t195 0.02262
R6991 CSoutput.n206 CSoutput.t198 0.02262
R6992 CSoutput CSoutput.n421 0.0052
R6993 CSoutput.n177 CSoutput.n160 0.00365111
R6994 CSoutput.n180 CSoutput.n161 0.00365111
R6995 CSoutput.n163 CSoutput.n162 0.00365111
R6996 CSoutput.n205 CSoutput.n164 0.00365111
R6997 CSoutput.n169 CSoutput.n165 0.00365111
R6998 CSoutput.n252 CSoutput.n166 0.00365111
R6999 CSoutput.n243 CSoutput.n242 0.00365111
R7000 CSoutput.n223 CSoutput.n196 0.00365111
R7001 CSoutput.n225 CSoutput.n195 0.00365111
R7002 CSoutput.n213 CSoutput.n212 0.00365111
R7003 CSoutput.n219 CSoutput.n199 0.00365111
R7004 CSoutput.n221 CSoutput.n198 0.00365111
R7005 CSoutput.n143 CSoutput.n126 0.00365111
R7006 CSoutput.n146 CSoutput.n127 0.00365111
R7007 CSoutput.n129 CSoutput.n128 0.00365111
R7008 CSoutput.n239 CSoutput.n130 0.00365111
R7009 CSoutput.n135 CSoutput.n131 0.00365111
R7010 CSoutput.n262 CSoutput.n132 0.00365111
R7011 CSoutput.n174 CSoutput.n164 0.00340054
R7012 CSoutput.n167 CSoutput.n165 0.00340054
R7013 CSoutput.n252 CSoutput.n251 0.00340054
R7014 CSoutput.n247 CSoutput.n160 0.00340054
R7015 CSoutput.n176 CSoutput.n161 0.00340054
R7016 CSoutput.n179 CSoutput.n163 0.00340054
R7017 CSoutput.n218 CSoutput.n213 0.00340054
R7018 CSoutput.n220 CSoutput.n219 0.00340054
R7019 CSoutput.n222 CSoutput.n221 0.00340054
R7020 CSoutput.n244 CSoutput.n243 0.00340054
R7021 CSoutput.n224 CSoutput.n223 0.00340054
R7022 CSoutput.n226 CSoutput.n225 0.00340054
R7023 CSoutput.n140 CSoutput.n130 0.00340054
R7024 CSoutput.n133 CSoutput.n131 0.00340054
R7025 CSoutput.n262 CSoutput.n261 0.00340054
R7026 CSoutput.n257 CSoutput.n126 0.00340054
R7027 CSoutput.n142 CSoutput.n127 0.00340054
R7028 CSoutput.n145 CSoutput.n129 0.00340054
R7029 CSoutput.n175 CSoutput.n169 0.00252698
R7030 CSoutput.n168 CSoutput.n166 0.00252698
R7031 CSoutput.n250 CSoutput.n249 0.00252698
R7032 CSoutput.n178 CSoutput.n176 0.00252698
R7033 CSoutput.n181 CSoutput.n179 0.00252698
R7034 CSoutput.n254 CSoutput.n149 0.00252698
R7035 CSoutput.n175 CSoutput.n174 0.00252698
R7036 CSoutput.n168 CSoutput.n167 0.00252698
R7037 CSoutput.n251 CSoutput.n250 0.00252698
R7038 CSoutput.n178 CSoutput.n177 0.00252698
R7039 CSoutput.n181 CSoutput.n180 0.00252698
R7040 CSoutput.n162 CSoutput.n149 0.00252698
R7041 CSoutput.n229 CSoutput.n199 0.00252698
R7042 CSoutput.n228 CSoutput.n198 0.00252698
R7043 CSoutput.n227 CSoutput.n183 0.00252698
R7044 CSoutput.n224 CSoutput.n194 0.00252698
R7045 CSoutput.n231 CSoutput.n226 0.00252698
R7046 CSoutput.n240 CSoutput.n233 0.00252698
R7047 CSoutput.n229 CSoutput.n218 0.00252698
R7048 CSoutput.n228 CSoutput.n220 0.00252698
R7049 CSoutput.n227 CSoutput.n222 0.00252698
R7050 CSoutput.n242 CSoutput.n194 0.00252698
R7051 CSoutput.n231 CSoutput.n196 0.00252698
R7052 CSoutput.n233 CSoutput.n195 0.00252698
R7053 CSoutput.n141 CSoutput.n135 0.00252698
R7054 CSoutput.n134 CSoutput.n132 0.00252698
R7055 CSoutput.n260 CSoutput.n259 0.00252698
R7056 CSoutput.n144 CSoutput.n142 0.00252698
R7057 CSoutput.n147 CSoutput.n145 0.00252698
R7058 CSoutput.n264 CSoutput.n115 0.00252698
R7059 CSoutput.n141 CSoutput.n140 0.00252698
R7060 CSoutput.n134 CSoutput.n133 0.00252698
R7061 CSoutput.n261 CSoutput.n260 0.00252698
R7062 CSoutput.n144 CSoutput.n143 0.00252698
R7063 CSoutput.n147 CSoutput.n146 0.00252698
R7064 CSoutput.n128 CSoutput.n115 0.00252698
R7065 CSoutput.n249 CSoutput.n248 0.0020275
R7066 CSoutput.n248 CSoutput.n247 0.0020275
R7067 CSoutput.n245 CSoutput.n183 0.0020275
R7068 CSoutput.n245 CSoutput.n244 0.0020275
R7069 CSoutput.n259 CSoutput.n258 0.0020275
R7070 CSoutput.n258 CSoutput.n257 0.0020275
R7071 CSoutput.n159 CSoutput.n158 0.00166668
R7072 CSoutput.n241 CSoutput.n197 0.00166668
R7073 CSoutput.n125 CSoutput.n124 0.00166668
R7074 CSoutput.n263 CSoutput.n125 0.00133328
R7075 CSoutput.n197 CSoutput.n193 0.00133328
R7076 CSoutput.n253 CSoutput.n159 0.00133328
R7077 CSoutput.n256 CSoutput.n148 0.001
R7078 CSoutput.n234 CSoutput.n148 0.001
R7079 CSoutput.n136 CSoutput.n116 0.001
R7080 CSoutput.n235 CSoutput.n116 0.001
R7081 CSoutput.n137 CSoutput.n117 0.001
R7082 CSoutput.n236 CSoutput.n117 0.001
R7083 CSoutput.n138 CSoutput.n118 0.001
R7084 CSoutput.n237 CSoutput.n118 0.001
R7085 CSoutput.n139 CSoutput.n119 0.001
R7086 CSoutput.n238 CSoutput.n119 0.001
R7087 CSoutput.n232 CSoutput.n184 0.001
R7088 CSoutput.n232 CSoutput.n230 0.001
R7089 CSoutput.n214 CSoutput.n185 0.001
R7090 CSoutput.n208 CSoutput.n185 0.001
R7091 CSoutput.n215 CSoutput.n186 0.001
R7092 CSoutput.n209 CSoutput.n186 0.001
R7093 CSoutput.n216 CSoutput.n187 0.001
R7094 CSoutput.n210 CSoutput.n187 0.001
R7095 CSoutput.n217 CSoutput.n188 0.001
R7096 CSoutput.n211 CSoutput.n188 0.001
R7097 CSoutput.n246 CSoutput.n182 0.001
R7098 CSoutput.n200 CSoutput.n182 0.001
R7099 CSoutput.n170 CSoutput.n150 0.001
R7100 CSoutput.n201 CSoutput.n150 0.001
R7101 CSoutput.n171 CSoutput.n151 0.001
R7102 CSoutput.n202 CSoutput.n151 0.001
R7103 CSoutput.n172 CSoutput.n152 0.001
R7104 CSoutput.n203 CSoutput.n152 0.001
R7105 CSoutput.n173 CSoutput.n153 0.001
R7106 CSoutput.n204 CSoutput.n153 0.001
R7107 CSoutput.n204 CSoutput.n154 0.001
R7108 CSoutput.n203 CSoutput.n155 0.001
R7109 CSoutput.n202 CSoutput.n156 0.001
R7110 CSoutput.n201 CSoutput.t213 0.001
R7111 CSoutput.n200 CSoutput.n157 0.001
R7112 CSoutput.n173 CSoutput.n155 0.001
R7113 CSoutput.n172 CSoutput.n156 0.001
R7114 CSoutput.n171 CSoutput.t213 0.001
R7115 CSoutput.n170 CSoutput.n157 0.001
R7116 CSoutput.n246 CSoutput.n158 0.001
R7117 CSoutput.n211 CSoutput.n189 0.001
R7118 CSoutput.n210 CSoutput.n190 0.001
R7119 CSoutput.n209 CSoutput.n191 0.001
R7120 CSoutput.n208 CSoutput.t208 0.001
R7121 CSoutput.n230 CSoutput.n192 0.001
R7122 CSoutput.n217 CSoutput.n190 0.001
R7123 CSoutput.n216 CSoutput.n191 0.001
R7124 CSoutput.n215 CSoutput.t208 0.001
R7125 CSoutput.n214 CSoutput.n192 0.001
R7126 CSoutput.n241 CSoutput.n184 0.001
R7127 CSoutput.n238 CSoutput.n120 0.001
R7128 CSoutput.n237 CSoutput.n121 0.001
R7129 CSoutput.n236 CSoutput.n122 0.001
R7130 CSoutput.n235 CSoutput.t206 0.001
R7131 CSoutput.n234 CSoutput.n123 0.001
R7132 CSoutput.n139 CSoutput.n121 0.001
R7133 CSoutput.n138 CSoutput.n122 0.001
R7134 CSoutput.n137 CSoutput.t206 0.001
R7135 CSoutput.n136 CSoutput.n123 0.001
R7136 CSoutput.n256 CSoutput.n124 0.001
R7137 plus.n53 plus.t20 323.478
R7138 plus.n11 plus.t15 323.478
R7139 plus.n52 plus.t19 297.12
R7140 plus.n56 plus.t26 297.12
R7141 plus.n58 plus.t25 297.12
R7142 plus.n62 plus.t27 297.12
R7143 plus.n64 plus.t9 297.12
R7144 plus.n68 plus.t7 297.12
R7145 plus.n70 plus.t14 297.12
R7146 plus.n74 plus.t12 297.12
R7147 plus.n76 plus.t28 297.12
R7148 plus.n80 plus.t10 297.12
R7149 plus.n82 plus.t8 297.12
R7150 plus.n40 plus.t21 297.12
R7151 plus.n38 plus.t22 297.12
R7152 plus.n2 plus.t16 297.12
R7153 plus.n32 plus.t17 297.12
R7154 plus.n4 plus.t11 297.12
R7155 plus.n26 plus.t5 297.12
R7156 plus.n6 plus.t6 297.12
R7157 plus.n20 plus.t23 297.12
R7158 plus.n8 plus.t24 297.12
R7159 plus.n14 plus.t18 297.12
R7160 plus.n10 plus.t13 297.12
R7161 plus.n86 plus.t3 243.97
R7162 plus.n86 plus.n85 223.454
R7163 plus.n88 plus.n87 223.454
R7164 plus.n83 plus.n82 161.3
R7165 plus.n81 plus.n42 161.3
R7166 plus.n80 plus.n79 161.3
R7167 plus.n78 plus.n43 161.3
R7168 plus.n77 plus.n76 161.3
R7169 plus.n75 plus.n44 161.3
R7170 plus.n74 plus.n73 161.3
R7171 plus.n72 plus.n45 161.3
R7172 plus.n71 plus.n70 161.3
R7173 plus.n69 plus.n46 161.3
R7174 plus.n68 plus.n67 161.3
R7175 plus.n66 plus.n47 161.3
R7176 plus.n65 plus.n64 161.3
R7177 plus.n63 plus.n48 161.3
R7178 plus.n62 plus.n61 161.3
R7179 plus.n60 plus.n49 161.3
R7180 plus.n59 plus.n58 161.3
R7181 plus.n57 plus.n50 161.3
R7182 plus.n56 plus.n55 161.3
R7183 plus.n54 plus.n51 161.3
R7184 plus.n13 plus.n12 161.3
R7185 plus.n14 plus.n9 161.3
R7186 plus.n16 plus.n15 161.3
R7187 plus.n17 plus.n8 161.3
R7188 plus.n19 plus.n18 161.3
R7189 plus.n20 plus.n7 161.3
R7190 plus.n22 plus.n21 161.3
R7191 plus.n23 plus.n6 161.3
R7192 plus.n25 plus.n24 161.3
R7193 plus.n26 plus.n5 161.3
R7194 plus.n28 plus.n27 161.3
R7195 plus.n29 plus.n4 161.3
R7196 plus.n31 plus.n30 161.3
R7197 plus.n32 plus.n3 161.3
R7198 plus.n34 plus.n33 161.3
R7199 plus.n35 plus.n2 161.3
R7200 plus.n37 plus.n36 161.3
R7201 plus.n38 plus.n1 161.3
R7202 plus.n39 plus.n0 161.3
R7203 plus.n41 plus.n40 161.3
R7204 plus.n82 plus.n81 46.0096
R7205 plus.n40 plus.n39 46.0096
R7206 plus.n54 plus.n53 45.0871
R7207 plus.n12 plus.n11 45.0871
R7208 plus.n52 plus.n51 41.6278
R7209 plus.n80 plus.n43 41.6278
R7210 plus.n38 plus.n37 41.6278
R7211 plus.n13 plus.n10 41.6278
R7212 plus.n57 plus.n56 37.246
R7213 plus.n76 plus.n75 37.246
R7214 plus.n33 plus.n2 37.246
R7215 plus.n15 plus.n14 37.246
R7216 plus.n84 plus.n83 33.1766
R7217 plus.n58 plus.n49 32.8641
R7218 plus.n74 plus.n45 32.8641
R7219 plus.n32 plus.n31 32.8641
R7220 plus.n19 plus.n8 32.8641
R7221 plus.n63 plus.n62 28.4823
R7222 plus.n70 plus.n69 28.4823
R7223 plus.n27 plus.n4 28.4823
R7224 plus.n21 plus.n20 28.4823
R7225 plus.n64 plus.n47 24.1005
R7226 plus.n68 plus.n47 24.1005
R7227 plus.n26 plus.n25 24.1005
R7228 plus.n25 plus.n6 24.1005
R7229 plus.n85 plus.t4 19.8005
R7230 plus.n85 plus.t1 19.8005
R7231 plus.n87 plus.t2 19.8005
R7232 plus.n87 plus.t0 19.8005
R7233 plus.n64 plus.n63 19.7187
R7234 plus.n69 plus.n68 19.7187
R7235 plus.n27 plus.n26 19.7187
R7236 plus.n21 plus.n6 19.7187
R7237 plus.n62 plus.n49 15.3369
R7238 plus.n70 plus.n45 15.3369
R7239 plus.n31 plus.n4 15.3369
R7240 plus.n20 plus.n19 15.3369
R7241 plus plus.n89 14.9059
R7242 plus.n53 plus.n52 14.1472
R7243 plus.n11 plus.n10 14.1472
R7244 plus.n84 plus.n41 11.8774
R7245 plus.n58 plus.n57 10.955
R7246 plus.n75 plus.n74 10.955
R7247 plus.n33 plus.n32 10.955
R7248 plus.n15 plus.n8 10.955
R7249 plus.n56 plus.n51 6.57323
R7250 plus.n76 plus.n43 6.57323
R7251 plus.n37 plus.n2 6.57323
R7252 plus.n14 plus.n13 6.57323
R7253 plus.n89 plus.n88 5.40567
R7254 plus.n81 plus.n80 2.19141
R7255 plus.n39 plus.n38 2.19141
R7256 plus.n89 plus.n84 1.188
R7257 plus.n88 plus.n86 0.716017
R7258 plus.n55 plus.n54 0.189894
R7259 plus.n55 plus.n50 0.189894
R7260 plus.n59 plus.n50 0.189894
R7261 plus.n60 plus.n59 0.189894
R7262 plus.n61 plus.n60 0.189894
R7263 plus.n61 plus.n48 0.189894
R7264 plus.n65 plus.n48 0.189894
R7265 plus.n66 plus.n65 0.189894
R7266 plus.n67 plus.n66 0.189894
R7267 plus.n67 plus.n46 0.189894
R7268 plus.n71 plus.n46 0.189894
R7269 plus.n72 plus.n71 0.189894
R7270 plus.n73 plus.n72 0.189894
R7271 plus.n73 plus.n44 0.189894
R7272 plus.n77 plus.n44 0.189894
R7273 plus.n78 plus.n77 0.189894
R7274 plus.n79 plus.n78 0.189894
R7275 plus.n79 plus.n42 0.189894
R7276 plus.n83 plus.n42 0.189894
R7277 plus.n41 plus.n0 0.189894
R7278 plus.n1 plus.n0 0.189894
R7279 plus.n36 plus.n1 0.189894
R7280 plus.n36 plus.n35 0.189894
R7281 plus.n35 plus.n34 0.189894
R7282 plus.n34 plus.n3 0.189894
R7283 plus.n30 plus.n3 0.189894
R7284 plus.n30 plus.n29 0.189894
R7285 plus.n29 plus.n28 0.189894
R7286 plus.n28 plus.n5 0.189894
R7287 plus.n24 plus.n5 0.189894
R7288 plus.n24 plus.n23 0.189894
R7289 plus.n23 plus.n22 0.189894
R7290 plus.n22 plus.n7 0.189894
R7291 plus.n18 plus.n7 0.189894
R7292 plus.n18 plus.n17 0.189894
R7293 plus.n17 plus.n16 0.189894
R7294 plus.n16 plus.n9 0.189894
R7295 plus.n12 plus.n9 0.189894
R7296 a_n2903_n3924.n30 a_n2903_n3924.t2 214.643
R7297 a_n2903_n3924.n37 a_n2903_n3924.t52 214.321
R7298 a_n2903_n3924.n36 a_n2903_n3924.t5 214.321
R7299 a_n2903_n3924.n35 a_n2903_n3924.t42 214.321
R7300 a_n2903_n3924.n34 a_n2903_n3924.t9 214.321
R7301 a_n2903_n3924.n33 a_n2903_n3924.t15 214.321
R7302 a_n2903_n3924.n32 a_n2903_n3924.t48 214.321
R7303 a_n2903_n3924.n31 a_n2903_n3924.t12 214.321
R7304 a_n2903_n3924.n13 a_n2903_n3924.t26 55.8337
R7305 a_n2903_n3924.n14 a_n2903_n3924.t43 55.8337
R7306 a_n2903_n3924.n25 a_n2903_n3924.t53 55.8337
R7307 a_n2903_n3924.n2 a_n2903_n3924.t38 55.8335
R7308 a_n2903_n3924.n39 a_n2903_n3924.t44 55.8335
R7309 a_n2903_n3924.n50 a_n2903_n3924.t47 55.8335
R7310 a_n2903_n3924.n51 a_n2903_n3924.t31 55.8335
R7311 a_n2903_n3924.n28 a_n2903_n3924.t25 55.8335
R7312 a_n2903_n3924.n57 a_n2903_n3924.n56 53.0054
R7313 a_n2903_n3924.n4 a_n2903_n3924.n3 53.0052
R7314 a_n2903_n3924.n6 a_n2903_n3924.n5 53.0052
R7315 a_n2903_n3924.n8 a_n2903_n3924.n7 53.0052
R7316 a_n2903_n3924.n10 a_n2903_n3924.n9 53.0052
R7317 a_n2903_n3924.n12 a_n2903_n3924.n11 53.0052
R7318 a_n2903_n3924.n16 a_n2903_n3924.n15 53.0052
R7319 a_n2903_n3924.n18 a_n2903_n3924.n17 53.0052
R7320 a_n2903_n3924.n20 a_n2903_n3924.n19 53.0052
R7321 a_n2903_n3924.n22 a_n2903_n3924.n21 53.0052
R7322 a_n2903_n3924.n24 a_n2903_n3924.n23 53.0052
R7323 a_n2903_n3924.n41 a_n2903_n3924.n40 53.0051
R7324 a_n2903_n3924.n43 a_n2903_n3924.n42 53.0051
R7325 a_n2903_n3924.n45 a_n2903_n3924.n44 53.0051
R7326 a_n2903_n3924.n47 a_n2903_n3924.n46 53.0051
R7327 a_n2903_n3924.n49 a_n2903_n3924.n48 53.0051
R7328 a_n2903_n3924.n53 a_n2903_n3924.n52 53.0051
R7329 a_n2903_n3924.n55 a_n2903_n3924.n54 53.0051
R7330 a_n2903_n3924.n1 a_n2903_n3924.n0 53.0051
R7331 a_n2903_n3924.n27 a_n2903_n3924.n26 53.0051
R7332 a_n2903_n3924.n29 a_n2903_n3924.n25 12.1986
R7333 a_n2903_n3924.n38 a_n2903_n3924.n2 12.1986
R7334 a_n2903_n3924.n29 a_n2903_n3924.n28 5.11903
R7335 a_n2903_n3924.n39 a_n2903_n3924.n38 5.11903
R7336 a_n2903_n3924.n40 a_n2903_n3924.t16 2.82907
R7337 a_n2903_n3924.n40 a_n2903_n3924.t13 2.82907
R7338 a_n2903_n3924.n42 a_n2903_n3924.t55 2.82907
R7339 a_n2903_n3924.n42 a_n2903_n3924.t7 2.82907
R7340 a_n2903_n3924.n44 a_n2903_n3924.t49 2.82907
R7341 a_n2903_n3924.n44 a_n2903_n3924.t46 2.82907
R7342 a_n2903_n3924.n46 a_n2903_n3924.t8 2.82907
R7343 a_n2903_n3924.n46 a_n2903_n3924.t1 2.82907
R7344 a_n2903_n3924.n48 a_n2903_n3924.t51 2.82907
R7345 a_n2903_n3924.n48 a_n2903_n3924.t0 2.82907
R7346 a_n2903_n3924.n52 a_n2903_n3924.t28 2.82907
R7347 a_n2903_n3924.n52 a_n2903_n3924.t33 2.82907
R7348 a_n2903_n3924.n54 a_n2903_n3924.t23 2.82907
R7349 a_n2903_n3924.n54 a_n2903_n3924.t22 2.82907
R7350 a_n2903_n3924.n0 a_n2903_n3924.t29 2.82907
R7351 a_n2903_n3924.n0 a_n2903_n3924.t35 2.82907
R7352 a_n2903_n3924.n26 a_n2903_n3924.t24 2.82907
R7353 a_n2903_n3924.n26 a_n2903_n3924.t30 2.82907
R7354 a_n2903_n3924.n3 a_n2903_n3924.t18 2.82907
R7355 a_n2903_n3924.n3 a_n2903_n3924.t36 2.82907
R7356 a_n2903_n3924.n5 a_n2903_n3924.t32 2.82907
R7357 a_n2903_n3924.n5 a_n2903_n3924.t34 2.82907
R7358 a_n2903_n3924.n7 a_n2903_n3924.t37 2.82907
R7359 a_n2903_n3924.n7 a_n2903_n3924.t39 2.82907
R7360 a_n2903_n3924.n9 a_n2903_n3924.t21 2.82907
R7361 a_n2903_n3924.n9 a_n2903_n3924.t19 2.82907
R7362 a_n2903_n3924.n11 a_n2903_n3924.t27 2.82907
R7363 a_n2903_n3924.n11 a_n2903_n3924.t20 2.82907
R7364 a_n2903_n3924.n15 a_n2903_n3924.t11 2.82907
R7365 a_n2903_n3924.n15 a_n2903_n3924.t6 2.82907
R7366 a_n2903_n3924.n17 a_n2903_n3924.t50 2.82907
R7367 a_n2903_n3924.n17 a_n2903_n3924.t14 2.82907
R7368 a_n2903_n3924.n19 a_n2903_n3924.t3 2.82907
R7369 a_n2903_n3924.n19 a_n2903_n3924.t4 2.82907
R7370 a_n2903_n3924.n21 a_n2903_n3924.t45 2.82907
R7371 a_n2903_n3924.n21 a_n2903_n3924.t54 2.82907
R7372 a_n2903_n3924.n23 a_n2903_n3924.t10 2.82907
R7373 a_n2903_n3924.n23 a_n2903_n3924.t17 2.82907
R7374 a_n2903_n3924.t41 a_n2903_n3924.n57 2.82907
R7375 a_n2903_n3924.n57 a_n2903_n3924.t40 2.82907
R7376 a_n2903_n3924.n38 a_n2903_n3924.n37 2.16406
R7377 a_n2903_n3924.n30 a_n2903_n3924.n29 1.95694
R7378 a_n2903_n3924.n32 a_n2903_n3924.n31 0.672012
R7379 a_n2903_n3924.n33 a_n2903_n3924.n32 0.672012
R7380 a_n2903_n3924.n34 a_n2903_n3924.n33 0.672012
R7381 a_n2903_n3924.n35 a_n2903_n3924.n34 0.672012
R7382 a_n2903_n3924.n36 a_n2903_n3924.n35 0.672012
R7383 a_n2903_n3924.n37 a_n2903_n3924.n36 0.672012
R7384 a_n2903_n3924.n25 a_n2903_n3924.n24 0.444466
R7385 a_n2903_n3924.n24 a_n2903_n3924.n22 0.444466
R7386 a_n2903_n3924.n22 a_n2903_n3924.n20 0.444466
R7387 a_n2903_n3924.n20 a_n2903_n3924.n18 0.444466
R7388 a_n2903_n3924.n18 a_n2903_n3924.n16 0.444466
R7389 a_n2903_n3924.n16 a_n2903_n3924.n14 0.444466
R7390 a_n2903_n3924.n13 a_n2903_n3924.n12 0.444466
R7391 a_n2903_n3924.n12 a_n2903_n3924.n10 0.444466
R7392 a_n2903_n3924.n10 a_n2903_n3924.n8 0.444466
R7393 a_n2903_n3924.n8 a_n2903_n3924.n6 0.444466
R7394 a_n2903_n3924.n6 a_n2903_n3924.n4 0.444466
R7395 a_n2903_n3924.n4 a_n2903_n3924.n2 0.444466
R7396 a_n2903_n3924.n28 a_n2903_n3924.n27 0.444466
R7397 a_n2903_n3924.n27 a_n2903_n3924.n1 0.444466
R7398 a_n2903_n3924.n56 a_n2903_n3924.n1 0.444466
R7399 a_n2903_n3924.n56 a_n2903_n3924.n55 0.444466
R7400 a_n2903_n3924.n55 a_n2903_n3924.n53 0.444466
R7401 a_n2903_n3924.n53 a_n2903_n3924.n51 0.444466
R7402 a_n2903_n3924.n50 a_n2903_n3924.n49 0.444466
R7403 a_n2903_n3924.n49 a_n2903_n3924.n47 0.444466
R7404 a_n2903_n3924.n47 a_n2903_n3924.n45 0.444466
R7405 a_n2903_n3924.n45 a_n2903_n3924.n43 0.444466
R7406 a_n2903_n3924.n43 a_n2903_n3924.n41 0.444466
R7407 a_n2903_n3924.n41 a_n2903_n3924.n39 0.444466
R7408 a_n2903_n3924.n31 a_n2903_n3924.n30 0.350064
R7409 a_n2903_n3924.n14 a_n2903_n3924.n13 0.235414
R7410 a_n2903_n3924.n51 a_n2903_n3924.n50 0.235414
R7411 gnd.n7135 gnd.n718 978.75
R7412 gnd.n6559 gnd.n5111 939.716
R7413 gnd.n3047 gnd.n3046 771.183
R7414 gnd.n4568 gnd.n1796 771.183
R7415 gnd.n3327 gnd.n2550 771.183
R7416 gnd.n4570 gnd.n1791 771.183
R7417 gnd.n6574 gnd.n1122 766.379
R7418 gnd.n6507 gnd.n1119 766.379
R7419 gnd.n5622 gnd.n5521 766.379
R7420 gnd.n5620 gnd.n5523 766.379
R7421 gnd.n6558 gnd.n5118 756.769
R7422 gnd.n6569 gnd.n6568 756.769
R7423 gnd.n5754 gnd.n5483 756.769
R7424 gnd.n5740 gnd.n5472 756.769
R7425 gnd.n251 gnd.n241 751.963
R7426 gnd.n440 gnd.n439 751.963
R7427 gnd.n1972 gnd.n1860 751.963
R7428 gnd.n4379 gnd.n1974 751.963
R7429 gnd.n1553 gnd.n1541 751.963
R7430 gnd.n3320 gnd.n3319 751.963
R7431 gnd.n2803 gnd.n1185 751.963
R7432 gnd.n2759 gnd.n2758 751.963
R7433 gnd.n6743 gnd.n950 723.135
R7434 gnd.n7134 gnd.n719 723.135
R7435 gnd.n7348 gnd.n7347 723.135
R7436 gnd.n2659 gnd.n2640 723.135
R7437 gnd.n7664 gnd.n245 696.707
R7438 gnd.n7540 gnd.n7539 696.707
R7439 gnd.n4382 gnd.n4381 696.707
R7440 gnd.n4499 gnd.n1906 696.707
R7441 gnd.n4811 gnd.n1546 696.707
R7442 gnd.n3269 gnd.n2581 696.707
R7443 gnd.n4989 gnd.n1258 696.707
R7444 gnd.n5109 gnd.n1189 696.707
R7445 gnd.n6743 gnd.n6742 585
R7446 gnd.n6744 gnd.n6743 585
R7447 gnd.n6741 gnd.n952 585
R7448 gnd.n952 gnd.n951 585
R7449 gnd.n6740 gnd.n6739 585
R7450 gnd.n6739 gnd.n6738 585
R7451 gnd.n957 gnd.n956 585
R7452 gnd.n6737 gnd.n957 585
R7453 gnd.n6735 gnd.n6734 585
R7454 gnd.n6736 gnd.n6735 585
R7455 gnd.n6733 gnd.n959 585
R7456 gnd.n959 gnd.n958 585
R7457 gnd.n6732 gnd.n6731 585
R7458 gnd.n6731 gnd.n6730 585
R7459 gnd.n965 gnd.n964 585
R7460 gnd.n6729 gnd.n965 585
R7461 gnd.n6727 gnd.n6726 585
R7462 gnd.n6728 gnd.n6727 585
R7463 gnd.n6725 gnd.n967 585
R7464 gnd.n967 gnd.n966 585
R7465 gnd.n6724 gnd.n6723 585
R7466 gnd.n6723 gnd.n6722 585
R7467 gnd.n973 gnd.n972 585
R7468 gnd.n6721 gnd.n973 585
R7469 gnd.n6719 gnd.n6718 585
R7470 gnd.n6720 gnd.n6719 585
R7471 gnd.n6717 gnd.n975 585
R7472 gnd.n975 gnd.n974 585
R7473 gnd.n6716 gnd.n6715 585
R7474 gnd.n6715 gnd.n6714 585
R7475 gnd.n981 gnd.n980 585
R7476 gnd.n6713 gnd.n981 585
R7477 gnd.n6711 gnd.n6710 585
R7478 gnd.n6712 gnd.n6711 585
R7479 gnd.n6709 gnd.n983 585
R7480 gnd.n983 gnd.n982 585
R7481 gnd.n6708 gnd.n6707 585
R7482 gnd.n6707 gnd.n6706 585
R7483 gnd.n989 gnd.n988 585
R7484 gnd.n6705 gnd.n989 585
R7485 gnd.n6703 gnd.n6702 585
R7486 gnd.n6704 gnd.n6703 585
R7487 gnd.n6701 gnd.n991 585
R7488 gnd.n991 gnd.n990 585
R7489 gnd.n6700 gnd.n6699 585
R7490 gnd.n6699 gnd.n6698 585
R7491 gnd.n997 gnd.n996 585
R7492 gnd.n6697 gnd.n997 585
R7493 gnd.n6695 gnd.n6694 585
R7494 gnd.n6696 gnd.n6695 585
R7495 gnd.n6693 gnd.n999 585
R7496 gnd.n999 gnd.n998 585
R7497 gnd.n6692 gnd.n6691 585
R7498 gnd.n6691 gnd.n6690 585
R7499 gnd.n1005 gnd.n1004 585
R7500 gnd.n6689 gnd.n1005 585
R7501 gnd.n6687 gnd.n6686 585
R7502 gnd.n6688 gnd.n6687 585
R7503 gnd.n6685 gnd.n1007 585
R7504 gnd.n1007 gnd.n1006 585
R7505 gnd.n6684 gnd.n6683 585
R7506 gnd.n6683 gnd.n6682 585
R7507 gnd.n1013 gnd.n1012 585
R7508 gnd.n6681 gnd.n1013 585
R7509 gnd.n6679 gnd.n6678 585
R7510 gnd.n6680 gnd.n6679 585
R7511 gnd.n6677 gnd.n1015 585
R7512 gnd.n1015 gnd.n1014 585
R7513 gnd.n6676 gnd.n6675 585
R7514 gnd.n6675 gnd.n6674 585
R7515 gnd.n1021 gnd.n1020 585
R7516 gnd.n6673 gnd.n1021 585
R7517 gnd.n6671 gnd.n6670 585
R7518 gnd.n6672 gnd.n6671 585
R7519 gnd.n6669 gnd.n1023 585
R7520 gnd.n1023 gnd.n1022 585
R7521 gnd.n6668 gnd.n6667 585
R7522 gnd.n6667 gnd.n6666 585
R7523 gnd.n1029 gnd.n1028 585
R7524 gnd.n6665 gnd.n1029 585
R7525 gnd.n6663 gnd.n6662 585
R7526 gnd.n6664 gnd.n6663 585
R7527 gnd.n6661 gnd.n1031 585
R7528 gnd.n1031 gnd.n1030 585
R7529 gnd.n6660 gnd.n6659 585
R7530 gnd.n6659 gnd.n6658 585
R7531 gnd.n1037 gnd.n1036 585
R7532 gnd.n6657 gnd.n1037 585
R7533 gnd.n6655 gnd.n6654 585
R7534 gnd.n6656 gnd.n6655 585
R7535 gnd.n6653 gnd.n1039 585
R7536 gnd.n1039 gnd.n1038 585
R7537 gnd.n6652 gnd.n6651 585
R7538 gnd.n6651 gnd.n6650 585
R7539 gnd.n1045 gnd.n1044 585
R7540 gnd.n6649 gnd.n1045 585
R7541 gnd.n6647 gnd.n6646 585
R7542 gnd.n6648 gnd.n6647 585
R7543 gnd.n6645 gnd.n1047 585
R7544 gnd.n1047 gnd.n1046 585
R7545 gnd.n6644 gnd.n6643 585
R7546 gnd.n6643 gnd.n6642 585
R7547 gnd.n1053 gnd.n1052 585
R7548 gnd.n6641 gnd.n1053 585
R7549 gnd.n6639 gnd.n6638 585
R7550 gnd.n6640 gnd.n6639 585
R7551 gnd.n6637 gnd.n1055 585
R7552 gnd.n1055 gnd.n1054 585
R7553 gnd.n6636 gnd.n6635 585
R7554 gnd.n6635 gnd.n6634 585
R7555 gnd.n1061 gnd.n1060 585
R7556 gnd.n6633 gnd.n1061 585
R7557 gnd.n6631 gnd.n6630 585
R7558 gnd.n6632 gnd.n6631 585
R7559 gnd.n6629 gnd.n1063 585
R7560 gnd.n1063 gnd.n1062 585
R7561 gnd.n6628 gnd.n6627 585
R7562 gnd.n6627 gnd.n6626 585
R7563 gnd.n1069 gnd.n1068 585
R7564 gnd.n6625 gnd.n1069 585
R7565 gnd.n6623 gnd.n6622 585
R7566 gnd.n6624 gnd.n6623 585
R7567 gnd.n6621 gnd.n1071 585
R7568 gnd.n1071 gnd.n1070 585
R7569 gnd.n6620 gnd.n6619 585
R7570 gnd.n6619 gnd.n6618 585
R7571 gnd.n1077 gnd.n1076 585
R7572 gnd.n6617 gnd.n1077 585
R7573 gnd.n6615 gnd.n6614 585
R7574 gnd.n6616 gnd.n6615 585
R7575 gnd.n6613 gnd.n1079 585
R7576 gnd.n1079 gnd.n1078 585
R7577 gnd.n6612 gnd.n6611 585
R7578 gnd.n6611 gnd.n6610 585
R7579 gnd.n1085 gnd.n1084 585
R7580 gnd.n6609 gnd.n1085 585
R7581 gnd.n6607 gnd.n6606 585
R7582 gnd.n6608 gnd.n6607 585
R7583 gnd.n6605 gnd.n1087 585
R7584 gnd.n1087 gnd.n1086 585
R7585 gnd.n6604 gnd.n6603 585
R7586 gnd.n6603 gnd.n6602 585
R7587 gnd.n1093 gnd.n1092 585
R7588 gnd.n6601 gnd.n1093 585
R7589 gnd.n6599 gnd.n6598 585
R7590 gnd.n6600 gnd.n6599 585
R7591 gnd.n6597 gnd.n1095 585
R7592 gnd.n1095 gnd.n1094 585
R7593 gnd.n6596 gnd.n6595 585
R7594 gnd.n6595 gnd.n6594 585
R7595 gnd.n1101 gnd.n1100 585
R7596 gnd.n6593 gnd.n1101 585
R7597 gnd.n6591 gnd.n6590 585
R7598 gnd.n6592 gnd.n6591 585
R7599 gnd.n6589 gnd.n1103 585
R7600 gnd.n1103 gnd.n1102 585
R7601 gnd.n6588 gnd.n6587 585
R7602 gnd.n6587 gnd.n6586 585
R7603 gnd.n1109 gnd.n1108 585
R7604 gnd.n6585 gnd.n1109 585
R7605 gnd.n6583 gnd.n6582 585
R7606 gnd.n6584 gnd.n6583 585
R7607 gnd.n6581 gnd.n1111 585
R7608 gnd.n1111 gnd.n1110 585
R7609 gnd.n6580 gnd.n6579 585
R7610 gnd.n6579 gnd.n6578 585
R7611 gnd.n1117 gnd.n1116 585
R7612 gnd.n6577 gnd.n1117 585
R7613 gnd.n950 gnd.n949 585
R7614 gnd.n6745 gnd.n950 585
R7615 gnd.n6748 gnd.n6747 585
R7616 gnd.n6747 gnd.n6746 585
R7617 gnd.n947 gnd.n946 585
R7618 gnd.n946 gnd.n945 585
R7619 gnd.n6753 gnd.n6752 585
R7620 gnd.n6754 gnd.n6753 585
R7621 gnd.n944 gnd.n943 585
R7622 gnd.n6755 gnd.n944 585
R7623 gnd.n6758 gnd.n6757 585
R7624 gnd.n6757 gnd.n6756 585
R7625 gnd.n941 gnd.n940 585
R7626 gnd.n940 gnd.n939 585
R7627 gnd.n6763 gnd.n6762 585
R7628 gnd.n6764 gnd.n6763 585
R7629 gnd.n938 gnd.n937 585
R7630 gnd.n6765 gnd.n938 585
R7631 gnd.n6768 gnd.n6767 585
R7632 gnd.n6767 gnd.n6766 585
R7633 gnd.n935 gnd.n934 585
R7634 gnd.n934 gnd.n933 585
R7635 gnd.n6773 gnd.n6772 585
R7636 gnd.n6774 gnd.n6773 585
R7637 gnd.n932 gnd.n931 585
R7638 gnd.n6775 gnd.n932 585
R7639 gnd.n6778 gnd.n6777 585
R7640 gnd.n6777 gnd.n6776 585
R7641 gnd.n929 gnd.n928 585
R7642 gnd.n928 gnd.n927 585
R7643 gnd.n6783 gnd.n6782 585
R7644 gnd.n6784 gnd.n6783 585
R7645 gnd.n926 gnd.n925 585
R7646 gnd.n6785 gnd.n926 585
R7647 gnd.n6788 gnd.n6787 585
R7648 gnd.n6787 gnd.n6786 585
R7649 gnd.n923 gnd.n922 585
R7650 gnd.n922 gnd.n921 585
R7651 gnd.n6793 gnd.n6792 585
R7652 gnd.n6794 gnd.n6793 585
R7653 gnd.n920 gnd.n919 585
R7654 gnd.n6795 gnd.n920 585
R7655 gnd.n6798 gnd.n6797 585
R7656 gnd.n6797 gnd.n6796 585
R7657 gnd.n917 gnd.n916 585
R7658 gnd.n916 gnd.n915 585
R7659 gnd.n6803 gnd.n6802 585
R7660 gnd.n6804 gnd.n6803 585
R7661 gnd.n914 gnd.n913 585
R7662 gnd.n6805 gnd.n914 585
R7663 gnd.n6808 gnd.n6807 585
R7664 gnd.n6807 gnd.n6806 585
R7665 gnd.n911 gnd.n910 585
R7666 gnd.n910 gnd.n909 585
R7667 gnd.n6813 gnd.n6812 585
R7668 gnd.n6814 gnd.n6813 585
R7669 gnd.n908 gnd.n907 585
R7670 gnd.n6815 gnd.n908 585
R7671 gnd.n6818 gnd.n6817 585
R7672 gnd.n6817 gnd.n6816 585
R7673 gnd.n905 gnd.n904 585
R7674 gnd.n904 gnd.n903 585
R7675 gnd.n6823 gnd.n6822 585
R7676 gnd.n6824 gnd.n6823 585
R7677 gnd.n902 gnd.n901 585
R7678 gnd.n6825 gnd.n902 585
R7679 gnd.n6828 gnd.n6827 585
R7680 gnd.n6827 gnd.n6826 585
R7681 gnd.n899 gnd.n898 585
R7682 gnd.n898 gnd.n897 585
R7683 gnd.n6833 gnd.n6832 585
R7684 gnd.n6834 gnd.n6833 585
R7685 gnd.n896 gnd.n895 585
R7686 gnd.n6835 gnd.n896 585
R7687 gnd.n6838 gnd.n6837 585
R7688 gnd.n6837 gnd.n6836 585
R7689 gnd.n893 gnd.n892 585
R7690 gnd.n892 gnd.n891 585
R7691 gnd.n6843 gnd.n6842 585
R7692 gnd.n6844 gnd.n6843 585
R7693 gnd.n890 gnd.n889 585
R7694 gnd.n6845 gnd.n890 585
R7695 gnd.n6848 gnd.n6847 585
R7696 gnd.n6847 gnd.n6846 585
R7697 gnd.n887 gnd.n886 585
R7698 gnd.n886 gnd.n885 585
R7699 gnd.n6853 gnd.n6852 585
R7700 gnd.n6854 gnd.n6853 585
R7701 gnd.n884 gnd.n883 585
R7702 gnd.n6855 gnd.n884 585
R7703 gnd.n6858 gnd.n6857 585
R7704 gnd.n6857 gnd.n6856 585
R7705 gnd.n881 gnd.n880 585
R7706 gnd.n880 gnd.n879 585
R7707 gnd.n6863 gnd.n6862 585
R7708 gnd.n6864 gnd.n6863 585
R7709 gnd.n878 gnd.n877 585
R7710 gnd.n6865 gnd.n878 585
R7711 gnd.n6868 gnd.n6867 585
R7712 gnd.n6867 gnd.n6866 585
R7713 gnd.n875 gnd.n874 585
R7714 gnd.n874 gnd.n873 585
R7715 gnd.n6873 gnd.n6872 585
R7716 gnd.n6874 gnd.n6873 585
R7717 gnd.n872 gnd.n871 585
R7718 gnd.n6875 gnd.n872 585
R7719 gnd.n6878 gnd.n6877 585
R7720 gnd.n6877 gnd.n6876 585
R7721 gnd.n869 gnd.n868 585
R7722 gnd.n868 gnd.n867 585
R7723 gnd.n6883 gnd.n6882 585
R7724 gnd.n6884 gnd.n6883 585
R7725 gnd.n866 gnd.n865 585
R7726 gnd.n6885 gnd.n866 585
R7727 gnd.n6888 gnd.n6887 585
R7728 gnd.n6887 gnd.n6886 585
R7729 gnd.n863 gnd.n862 585
R7730 gnd.n862 gnd.n861 585
R7731 gnd.n6893 gnd.n6892 585
R7732 gnd.n6894 gnd.n6893 585
R7733 gnd.n860 gnd.n859 585
R7734 gnd.n6895 gnd.n860 585
R7735 gnd.n6898 gnd.n6897 585
R7736 gnd.n6897 gnd.n6896 585
R7737 gnd.n857 gnd.n856 585
R7738 gnd.n856 gnd.n855 585
R7739 gnd.n6903 gnd.n6902 585
R7740 gnd.n6904 gnd.n6903 585
R7741 gnd.n854 gnd.n853 585
R7742 gnd.n6905 gnd.n854 585
R7743 gnd.n6908 gnd.n6907 585
R7744 gnd.n6907 gnd.n6906 585
R7745 gnd.n851 gnd.n850 585
R7746 gnd.n850 gnd.n849 585
R7747 gnd.n6913 gnd.n6912 585
R7748 gnd.n6914 gnd.n6913 585
R7749 gnd.n848 gnd.n847 585
R7750 gnd.n6915 gnd.n848 585
R7751 gnd.n6918 gnd.n6917 585
R7752 gnd.n6917 gnd.n6916 585
R7753 gnd.n845 gnd.n844 585
R7754 gnd.n844 gnd.n843 585
R7755 gnd.n6923 gnd.n6922 585
R7756 gnd.n6924 gnd.n6923 585
R7757 gnd.n842 gnd.n841 585
R7758 gnd.n6925 gnd.n842 585
R7759 gnd.n6928 gnd.n6927 585
R7760 gnd.n6927 gnd.n6926 585
R7761 gnd.n839 gnd.n838 585
R7762 gnd.n838 gnd.n837 585
R7763 gnd.n6933 gnd.n6932 585
R7764 gnd.n6934 gnd.n6933 585
R7765 gnd.n836 gnd.n835 585
R7766 gnd.n6935 gnd.n836 585
R7767 gnd.n6938 gnd.n6937 585
R7768 gnd.n6937 gnd.n6936 585
R7769 gnd.n833 gnd.n832 585
R7770 gnd.n832 gnd.n831 585
R7771 gnd.n6943 gnd.n6942 585
R7772 gnd.n6944 gnd.n6943 585
R7773 gnd.n830 gnd.n829 585
R7774 gnd.n6945 gnd.n830 585
R7775 gnd.n6948 gnd.n6947 585
R7776 gnd.n6947 gnd.n6946 585
R7777 gnd.n827 gnd.n826 585
R7778 gnd.n826 gnd.n825 585
R7779 gnd.n6953 gnd.n6952 585
R7780 gnd.n6954 gnd.n6953 585
R7781 gnd.n824 gnd.n823 585
R7782 gnd.n6955 gnd.n824 585
R7783 gnd.n6958 gnd.n6957 585
R7784 gnd.n6957 gnd.n6956 585
R7785 gnd.n821 gnd.n820 585
R7786 gnd.n820 gnd.n819 585
R7787 gnd.n6963 gnd.n6962 585
R7788 gnd.n6964 gnd.n6963 585
R7789 gnd.n818 gnd.n817 585
R7790 gnd.n6965 gnd.n818 585
R7791 gnd.n6968 gnd.n6967 585
R7792 gnd.n6967 gnd.n6966 585
R7793 gnd.n815 gnd.n814 585
R7794 gnd.n814 gnd.n813 585
R7795 gnd.n6973 gnd.n6972 585
R7796 gnd.n6974 gnd.n6973 585
R7797 gnd.n812 gnd.n811 585
R7798 gnd.n6975 gnd.n812 585
R7799 gnd.n6978 gnd.n6977 585
R7800 gnd.n6977 gnd.n6976 585
R7801 gnd.n809 gnd.n808 585
R7802 gnd.n808 gnd.n807 585
R7803 gnd.n6983 gnd.n6982 585
R7804 gnd.n6984 gnd.n6983 585
R7805 gnd.n806 gnd.n805 585
R7806 gnd.n6985 gnd.n806 585
R7807 gnd.n6988 gnd.n6987 585
R7808 gnd.n6987 gnd.n6986 585
R7809 gnd.n803 gnd.n802 585
R7810 gnd.n802 gnd.n801 585
R7811 gnd.n6993 gnd.n6992 585
R7812 gnd.n6994 gnd.n6993 585
R7813 gnd.n800 gnd.n799 585
R7814 gnd.n6995 gnd.n800 585
R7815 gnd.n6998 gnd.n6997 585
R7816 gnd.n6997 gnd.n6996 585
R7817 gnd.n797 gnd.n796 585
R7818 gnd.n796 gnd.n795 585
R7819 gnd.n7003 gnd.n7002 585
R7820 gnd.n7004 gnd.n7003 585
R7821 gnd.n794 gnd.n793 585
R7822 gnd.n7005 gnd.n794 585
R7823 gnd.n7008 gnd.n7007 585
R7824 gnd.n7007 gnd.n7006 585
R7825 gnd.n791 gnd.n790 585
R7826 gnd.n790 gnd.n789 585
R7827 gnd.n7013 gnd.n7012 585
R7828 gnd.n7014 gnd.n7013 585
R7829 gnd.n788 gnd.n787 585
R7830 gnd.n7015 gnd.n788 585
R7831 gnd.n7018 gnd.n7017 585
R7832 gnd.n7017 gnd.n7016 585
R7833 gnd.n785 gnd.n784 585
R7834 gnd.n784 gnd.n783 585
R7835 gnd.n7023 gnd.n7022 585
R7836 gnd.n7024 gnd.n7023 585
R7837 gnd.n782 gnd.n781 585
R7838 gnd.n7025 gnd.n782 585
R7839 gnd.n7028 gnd.n7027 585
R7840 gnd.n7027 gnd.n7026 585
R7841 gnd.n779 gnd.n778 585
R7842 gnd.n778 gnd.n777 585
R7843 gnd.n7033 gnd.n7032 585
R7844 gnd.n7034 gnd.n7033 585
R7845 gnd.n776 gnd.n775 585
R7846 gnd.n7035 gnd.n776 585
R7847 gnd.n7038 gnd.n7037 585
R7848 gnd.n7037 gnd.n7036 585
R7849 gnd.n773 gnd.n772 585
R7850 gnd.n772 gnd.n771 585
R7851 gnd.n7043 gnd.n7042 585
R7852 gnd.n7044 gnd.n7043 585
R7853 gnd.n770 gnd.n769 585
R7854 gnd.n7045 gnd.n770 585
R7855 gnd.n7048 gnd.n7047 585
R7856 gnd.n7047 gnd.n7046 585
R7857 gnd.n767 gnd.n766 585
R7858 gnd.n766 gnd.n765 585
R7859 gnd.n7053 gnd.n7052 585
R7860 gnd.n7054 gnd.n7053 585
R7861 gnd.n764 gnd.n763 585
R7862 gnd.n7055 gnd.n764 585
R7863 gnd.n7058 gnd.n7057 585
R7864 gnd.n7057 gnd.n7056 585
R7865 gnd.n761 gnd.n760 585
R7866 gnd.n760 gnd.n759 585
R7867 gnd.n7063 gnd.n7062 585
R7868 gnd.n7064 gnd.n7063 585
R7869 gnd.n758 gnd.n757 585
R7870 gnd.n7065 gnd.n758 585
R7871 gnd.n7068 gnd.n7067 585
R7872 gnd.n7067 gnd.n7066 585
R7873 gnd.n755 gnd.n754 585
R7874 gnd.n754 gnd.n753 585
R7875 gnd.n7073 gnd.n7072 585
R7876 gnd.n7074 gnd.n7073 585
R7877 gnd.n752 gnd.n751 585
R7878 gnd.n7075 gnd.n752 585
R7879 gnd.n7078 gnd.n7077 585
R7880 gnd.n7077 gnd.n7076 585
R7881 gnd.n749 gnd.n748 585
R7882 gnd.n748 gnd.n747 585
R7883 gnd.n7083 gnd.n7082 585
R7884 gnd.n7084 gnd.n7083 585
R7885 gnd.n746 gnd.n745 585
R7886 gnd.n7085 gnd.n746 585
R7887 gnd.n7088 gnd.n7087 585
R7888 gnd.n7087 gnd.n7086 585
R7889 gnd.n743 gnd.n742 585
R7890 gnd.n742 gnd.n741 585
R7891 gnd.n7093 gnd.n7092 585
R7892 gnd.n7094 gnd.n7093 585
R7893 gnd.n740 gnd.n739 585
R7894 gnd.n7095 gnd.n740 585
R7895 gnd.n7098 gnd.n7097 585
R7896 gnd.n7097 gnd.n7096 585
R7897 gnd.n737 gnd.n736 585
R7898 gnd.n736 gnd.n735 585
R7899 gnd.n7103 gnd.n7102 585
R7900 gnd.n7104 gnd.n7103 585
R7901 gnd.n734 gnd.n733 585
R7902 gnd.n7105 gnd.n734 585
R7903 gnd.n7108 gnd.n7107 585
R7904 gnd.n7107 gnd.n7106 585
R7905 gnd.n731 gnd.n730 585
R7906 gnd.n730 gnd.n729 585
R7907 gnd.n7113 gnd.n7112 585
R7908 gnd.n7114 gnd.n7113 585
R7909 gnd.n728 gnd.n727 585
R7910 gnd.n7115 gnd.n728 585
R7911 gnd.n7118 gnd.n7117 585
R7912 gnd.n7117 gnd.n7116 585
R7913 gnd.n725 gnd.n724 585
R7914 gnd.n724 gnd.n723 585
R7915 gnd.n7124 gnd.n7123 585
R7916 gnd.n7125 gnd.n7124 585
R7917 gnd.n722 gnd.n721 585
R7918 gnd.n7126 gnd.n722 585
R7919 gnd.n7129 gnd.n7128 585
R7920 gnd.n7128 gnd.n7127 585
R7921 gnd.n7130 gnd.n719 585
R7922 gnd.n719 gnd.n718 585
R7923 gnd.n594 gnd.n593 585
R7924 gnd.n7338 gnd.n593 585
R7925 gnd.n7341 gnd.n7340 585
R7926 gnd.n7340 gnd.n7339 585
R7927 gnd.n597 gnd.n596 585
R7928 gnd.n7336 gnd.n597 585
R7929 gnd.n7334 gnd.n7333 585
R7930 gnd.n7335 gnd.n7334 585
R7931 gnd.n600 gnd.n599 585
R7932 gnd.n599 gnd.n598 585
R7933 gnd.n7329 gnd.n7328 585
R7934 gnd.n7328 gnd.n7327 585
R7935 gnd.n603 gnd.n602 585
R7936 gnd.n7326 gnd.n603 585
R7937 gnd.n7324 gnd.n7323 585
R7938 gnd.n7325 gnd.n7324 585
R7939 gnd.n606 gnd.n605 585
R7940 gnd.n605 gnd.n604 585
R7941 gnd.n7319 gnd.n7318 585
R7942 gnd.n7318 gnd.n7317 585
R7943 gnd.n609 gnd.n608 585
R7944 gnd.n7316 gnd.n609 585
R7945 gnd.n7314 gnd.n7313 585
R7946 gnd.n7315 gnd.n7314 585
R7947 gnd.n612 gnd.n611 585
R7948 gnd.n611 gnd.n610 585
R7949 gnd.n7309 gnd.n7308 585
R7950 gnd.n7308 gnd.n7307 585
R7951 gnd.n615 gnd.n614 585
R7952 gnd.n7306 gnd.n615 585
R7953 gnd.n7304 gnd.n7303 585
R7954 gnd.n7305 gnd.n7304 585
R7955 gnd.n618 gnd.n617 585
R7956 gnd.n617 gnd.n616 585
R7957 gnd.n7299 gnd.n7298 585
R7958 gnd.n7298 gnd.n7297 585
R7959 gnd.n621 gnd.n620 585
R7960 gnd.n7296 gnd.n621 585
R7961 gnd.n7294 gnd.n7293 585
R7962 gnd.n7295 gnd.n7294 585
R7963 gnd.n624 gnd.n623 585
R7964 gnd.n623 gnd.n622 585
R7965 gnd.n7289 gnd.n7288 585
R7966 gnd.n7288 gnd.n7287 585
R7967 gnd.n627 gnd.n626 585
R7968 gnd.n7286 gnd.n627 585
R7969 gnd.n7284 gnd.n7283 585
R7970 gnd.n7285 gnd.n7284 585
R7971 gnd.n630 gnd.n629 585
R7972 gnd.n629 gnd.n628 585
R7973 gnd.n7279 gnd.n7278 585
R7974 gnd.n7278 gnd.n7277 585
R7975 gnd.n633 gnd.n632 585
R7976 gnd.n7276 gnd.n633 585
R7977 gnd.n7274 gnd.n7273 585
R7978 gnd.n7275 gnd.n7274 585
R7979 gnd.n636 gnd.n635 585
R7980 gnd.n635 gnd.n634 585
R7981 gnd.n7269 gnd.n7268 585
R7982 gnd.n7268 gnd.n7267 585
R7983 gnd.n639 gnd.n638 585
R7984 gnd.n7266 gnd.n639 585
R7985 gnd.n7264 gnd.n7263 585
R7986 gnd.n7265 gnd.n7264 585
R7987 gnd.n642 gnd.n641 585
R7988 gnd.n641 gnd.n640 585
R7989 gnd.n7259 gnd.n7258 585
R7990 gnd.n7258 gnd.n7257 585
R7991 gnd.n645 gnd.n644 585
R7992 gnd.n7256 gnd.n645 585
R7993 gnd.n7254 gnd.n7253 585
R7994 gnd.n7255 gnd.n7254 585
R7995 gnd.n648 gnd.n647 585
R7996 gnd.n647 gnd.n646 585
R7997 gnd.n7249 gnd.n7248 585
R7998 gnd.n7248 gnd.n7247 585
R7999 gnd.n651 gnd.n650 585
R8000 gnd.n7246 gnd.n651 585
R8001 gnd.n7244 gnd.n7243 585
R8002 gnd.n7245 gnd.n7244 585
R8003 gnd.n654 gnd.n653 585
R8004 gnd.n653 gnd.n652 585
R8005 gnd.n7239 gnd.n7238 585
R8006 gnd.n7238 gnd.n7237 585
R8007 gnd.n657 gnd.n656 585
R8008 gnd.n7236 gnd.n657 585
R8009 gnd.n7234 gnd.n7233 585
R8010 gnd.n7235 gnd.n7234 585
R8011 gnd.n660 gnd.n659 585
R8012 gnd.n659 gnd.n658 585
R8013 gnd.n7229 gnd.n7228 585
R8014 gnd.n7228 gnd.n7227 585
R8015 gnd.n663 gnd.n662 585
R8016 gnd.n7226 gnd.n663 585
R8017 gnd.n7224 gnd.n7223 585
R8018 gnd.n7225 gnd.n7224 585
R8019 gnd.n666 gnd.n665 585
R8020 gnd.n665 gnd.n664 585
R8021 gnd.n7219 gnd.n7218 585
R8022 gnd.n7218 gnd.n7217 585
R8023 gnd.n669 gnd.n668 585
R8024 gnd.n7216 gnd.n669 585
R8025 gnd.n7214 gnd.n7213 585
R8026 gnd.n7215 gnd.n7214 585
R8027 gnd.n672 gnd.n671 585
R8028 gnd.n671 gnd.n670 585
R8029 gnd.n7209 gnd.n7208 585
R8030 gnd.n7208 gnd.n7207 585
R8031 gnd.n675 gnd.n674 585
R8032 gnd.n7206 gnd.n675 585
R8033 gnd.n7204 gnd.n7203 585
R8034 gnd.n7205 gnd.n7204 585
R8035 gnd.n678 gnd.n677 585
R8036 gnd.n677 gnd.n676 585
R8037 gnd.n7199 gnd.n7198 585
R8038 gnd.n7198 gnd.n7197 585
R8039 gnd.n681 gnd.n680 585
R8040 gnd.n7196 gnd.n681 585
R8041 gnd.n7194 gnd.n7193 585
R8042 gnd.n7195 gnd.n7194 585
R8043 gnd.n684 gnd.n683 585
R8044 gnd.n683 gnd.n682 585
R8045 gnd.n7189 gnd.n7188 585
R8046 gnd.n7188 gnd.n7187 585
R8047 gnd.n687 gnd.n686 585
R8048 gnd.n7186 gnd.n687 585
R8049 gnd.n7184 gnd.n7183 585
R8050 gnd.n7185 gnd.n7184 585
R8051 gnd.n690 gnd.n689 585
R8052 gnd.n689 gnd.n688 585
R8053 gnd.n7179 gnd.n7178 585
R8054 gnd.n7178 gnd.n7177 585
R8055 gnd.n693 gnd.n692 585
R8056 gnd.n7176 gnd.n693 585
R8057 gnd.n7174 gnd.n7173 585
R8058 gnd.n7175 gnd.n7174 585
R8059 gnd.n696 gnd.n695 585
R8060 gnd.n695 gnd.n694 585
R8061 gnd.n7169 gnd.n7168 585
R8062 gnd.n7168 gnd.n7167 585
R8063 gnd.n699 gnd.n698 585
R8064 gnd.n7166 gnd.n699 585
R8065 gnd.n7164 gnd.n7163 585
R8066 gnd.n7165 gnd.n7164 585
R8067 gnd.n702 gnd.n701 585
R8068 gnd.n701 gnd.n700 585
R8069 gnd.n7159 gnd.n7158 585
R8070 gnd.n7158 gnd.n7157 585
R8071 gnd.n705 gnd.n704 585
R8072 gnd.n7156 gnd.n705 585
R8073 gnd.n7154 gnd.n7153 585
R8074 gnd.n7155 gnd.n7154 585
R8075 gnd.n708 gnd.n707 585
R8076 gnd.n707 gnd.n706 585
R8077 gnd.n7149 gnd.n7148 585
R8078 gnd.n7148 gnd.n7147 585
R8079 gnd.n711 gnd.n710 585
R8080 gnd.n7146 gnd.n711 585
R8081 gnd.n7144 gnd.n7143 585
R8082 gnd.n7145 gnd.n7144 585
R8083 gnd.n714 gnd.n713 585
R8084 gnd.n713 gnd.n712 585
R8085 gnd.n7139 gnd.n7138 585
R8086 gnd.n7138 gnd.n7137 585
R8087 gnd.n717 gnd.n716 585
R8088 gnd.n7136 gnd.n717 585
R8089 gnd.n7134 gnd.n7133 585
R8090 gnd.n7135 gnd.n7134 585
R8091 gnd.n1541 gnd.n1540 585
R8092 gnd.n3318 gnd.n1541 585
R8093 gnd.n4820 gnd.n4819 585
R8094 gnd.n4819 gnd.n4818 585
R8095 gnd.n4821 gnd.n1536 585
R8096 gnd.n3278 gnd.n1536 585
R8097 gnd.n4823 gnd.n4822 585
R8098 gnd.n4824 gnd.n4823 585
R8099 gnd.n1520 gnd.n1519 585
R8100 gnd.n3026 gnd.n1520 585
R8101 gnd.n4832 gnd.n4831 585
R8102 gnd.n4831 gnd.n4830 585
R8103 gnd.n4833 gnd.n1515 585
R8104 gnd.n3291 gnd.n1515 585
R8105 gnd.n4835 gnd.n4834 585
R8106 gnd.n4836 gnd.n4835 585
R8107 gnd.n1501 gnd.n1500 585
R8108 gnd.n3019 gnd.n1501 585
R8109 gnd.n4844 gnd.n4843 585
R8110 gnd.n4843 gnd.n4842 585
R8111 gnd.n4845 gnd.n1496 585
R8112 gnd.n3011 gnd.n1496 585
R8113 gnd.n4847 gnd.n4846 585
R8114 gnd.n4848 gnd.n4847 585
R8115 gnd.n1480 gnd.n1479 585
R8116 gnd.n2973 gnd.n1480 585
R8117 gnd.n4856 gnd.n4855 585
R8118 gnd.n4855 gnd.n4854 585
R8119 gnd.n4857 gnd.n1475 585
R8120 gnd.n2964 gnd.n1475 585
R8121 gnd.n4859 gnd.n4858 585
R8122 gnd.n4860 gnd.n4859 585
R8123 gnd.n1461 gnd.n1460 585
R8124 gnd.n2959 gnd.n1461 585
R8125 gnd.n4868 gnd.n4867 585
R8126 gnd.n4867 gnd.n4866 585
R8127 gnd.n4869 gnd.n1456 585
R8128 gnd.n2987 gnd.n1456 585
R8129 gnd.n4871 gnd.n4870 585
R8130 gnd.n4872 gnd.n4871 585
R8131 gnd.n1440 gnd.n1439 585
R8132 gnd.n2952 gnd.n1440 585
R8133 gnd.n4880 gnd.n4879 585
R8134 gnd.n4879 gnd.n4878 585
R8135 gnd.n4881 gnd.n1435 585
R8136 gnd.n2944 gnd.n1435 585
R8137 gnd.n4883 gnd.n4882 585
R8138 gnd.n4884 gnd.n4883 585
R8139 gnd.n1422 gnd.n1421 585
R8140 gnd.n2938 gnd.n1422 585
R8141 gnd.n4892 gnd.n4891 585
R8142 gnd.n4891 gnd.n4890 585
R8143 gnd.n4893 gnd.n1416 585
R8144 gnd.n2930 gnd.n1416 585
R8145 gnd.n4895 gnd.n4894 585
R8146 gnd.n4896 gnd.n4895 585
R8147 gnd.n1417 gnd.n1415 585
R8148 gnd.n2899 gnd.n1415 585
R8149 gnd.n2881 gnd.n2880 585
R8150 gnd.n2880 gnd.n2641 585
R8151 gnd.n2882 gnd.n2650 585
R8152 gnd.n2891 gnd.n2650 585
R8153 gnd.n2884 gnd.n2883 585
R8154 gnd.n2885 gnd.n2884 585
R8155 gnd.n2663 gnd.n2662 585
R8156 gnd.n2869 gnd.n2662 585
R8157 gnd.n2723 gnd.n2722 585
R8158 gnd.n2726 gnd.n2723 585
R8159 gnd.n1395 gnd.n1394 585
R8160 gnd.n1398 gnd.n1395 585
R8161 gnd.n4905 gnd.n4904 585
R8162 gnd.n4904 gnd.n4903 585
R8163 gnd.n4906 gnd.n1390 585
R8164 gnd.n1390 gnd.n1389 585
R8165 gnd.n4908 gnd.n4907 585
R8166 gnd.n4909 gnd.n4908 585
R8167 gnd.n1377 gnd.n1376 585
R8168 gnd.n1386 gnd.n1377 585
R8169 gnd.n4917 gnd.n4916 585
R8170 gnd.n4916 gnd.n4915 585
R8171 gnd.n4918 gnd.n1372 585
R8172 gnd.n1372 gnd.n1371 585
R8173 gnd.n4920 gnd.n4919 585
R8174 gnd.n4921 gnd.n4920 585
R8175 gnd.n1358 gnd.n1357 585
R8176 gnd.n1361 gnd.n1358 585
R8177 gnd.n4929 gnd.n4928 585
R8178 gnd.n4928 gnd.n4927 585
R8179 gnd.n4930 gnd.n1353 585
R8180 gnd.n1353 gnd.n1352 585
R8181 gnd.n4932 gnd.n4931 585
R8182 gnd.n4933 gnd.n4932 585
R8183 gnd.n1339 gnd.n1338 585
R8184 gnd.n1349 gnd.n1339 585
R8185 gnd.n4941 gnd.n4940 585
R8186 gnd.n4940 gnd.n4939 585
R8187 gnd.n4942 gnd.n1334 585
R8188 gnd.n1334 gnd.n1333 585
R8189 gnd.n4944 gnd.n4943 585
R8190 gnd.n4945 gnd.n4944 585
R8191 gnd.n1320 gnd.n1319 585
R8192 gnd.n1323 gnd.n1320 585
R8193 gnd.n4953 gnd.n4952 585
R8194 gnd.n4952 gnd.n4951 585
R8195 gnd.n4954 gnd.n1315 585
R8196 gnd.n1315 gnd.n1314 585
R8197 gnd.n4956 gnd.n4955 585
R8198 gnd.n4957 gnd.n4956 585
R8199 gnd.n1301 gnd.n1300 585
R8200 gnd.n1311 gnd.n1301 585
R8201 gnd.n4965 gnd.n4964 585
R8202 gnd.n4964 gnd.n4963 585
R8203 gnd.n4966 gnd.n1296 585
R8204 gnd.n1296 gnd.n1295 585
R8205 gnd.n4968 gnd.n4967 585
R8206 gnd.n4969 gnd.n4968 585
R8207 gnd.n1282 gnd.n1281 585
R8208 gnd.n1285 gnd.n1282 585
R8209 gnd.n4977 gnd.n4976 585
R8210 gnd.n4976 gnd.n4975 585
R8211 gnd.n4978 gnd.n1275 585
R8212 gnd.n1275 gnd.n1273 585
R8213 gnd.n4980 gnd.n4979 585
R8214 gnd.n4981 gnd.n4980 585
R8215 gnd.n1277 gnd.n1274 585
R8216 gnd.n1274 gnd.n1270 585
R8217 gnd.n1276 gnd.n1261 585
R8218 gnd.n4987 gnd.n1261 585
R8219 gnd.n2758 gnd.n1255 585
R8220 gnd.n2758 gnd.n1186 585
R8221 gnd.n2760 gnd.n2759 585
R8222 gnd.n2762 gnd.n2761 585
R8223 gnd.n2764 gnd.n2763 585
R8224 gnd.n2768 gnd.n2756 585
R8225 gnd.n2770 gnd.n2769 585
R8226 gnd.n2772 gnd.n2771 585
R8227 gnd.n2774 gnd.n2773 585
R8228 gnd.n2778 gnd.n2754 585
R8229 gnd.n2780 gnd.n2779 585
R8230 gnd.n2782 gnd.n2781 585
R8231 gnd.n2784 gnd.n2783 585
R8232 gnd.n2788 gnd.n2752 585
R8233 gnd.n2790 gnd.n2789 585
R8234 gnd.n2792 gnd.n2791 585
R8235 gnd.n2794 gnd.n2793 585
R8236 gnd.n2749 gnd.n2748 585
R8237 gnd.n2798 gnd.n2750 585
R8238 gnd.n2799 gnd.n2745 585
R8239 gnd.n2800 gnd.n1185 585
R8240 gnd.n5111 gnd.n1185 585
R8241 gnd.n3321 gnd.n3320 585
R8242 gnd.n3115 gnd.n2579 585
R8243 gnd.n3127 gnd.n3116 585
R8244 gnd.n3128 gnd.n3114 585
R8245 gnd.n3113 gnd.n3105 585
R8246 gnd.n3135 gnd.n3104 585
R8247 gnd.n3136 gnd.n3103 585
R8248 gnd.n3097 gnd.n3096 585
R8249 gnd.n3143 gnd.n3095 585
R8250 gnd.n3144 gnd.n3094 585
R8251 gnd.n3093 gnd.n3085 585
R8252 gnd.n3151 gnd.n3084 585
R8253 gnd.n3152 gnd.n3083 585
R8254 gnd.n3077 gnd.n3076 585
R8255 gnd.n3159 gnd.n3075 585
R8256 gnd.n3160 gnd.n3074 585
R8257 gnd.n3073 gnd.n3065 585
R8258 gnd.n3167 gnd.n3064 585
R8259 gnd.n3168 gnd.n1553 585
R8260 gnd.n4810 gnd.n1553 585
R8261 gnd.n3319 gnd.n2580 585
R8262 gnd.n3319 gnd.n3318 585
R8263 gnd.n3280 gnd.n1544 585
R8264 gnd.n4818 gnd.n1544 585
R8265 gnd.n3283 gnd.n3279 585
R8266 gnd.n3279 gnd.n3278 585
R8267 gnd.n3284 gnd.n1534 585
R8268 gnd.n4824 gnd.n1534 585
R8269 gnd.n3285 gnd.n2597 585
R8270 gnd.n3026 gnd.n2597 585
R8271 gnd.n2594 gnd.n1523 585
R8272 gnd.n4830 gnd.n1523 585
R8273 gnd.n3290 gnd.n3289 585
R8274 gnd.n3291 gnd.n3290 585
R8275 gnd.n2593 gnd.n1514 585
R8276 gnd.n4836 gnd.n1514 585
R8277 gnd.n3018 gnd.n3017 585
R8278 gnd.n3019 gnd.n3018 585
R8279 gnd.n2600 gnd.n1503 585
R8280 gnd.n4842 gnd.n1503 585
R8281 gnd.n3013 gnd.n3012 585
R8282 gnd.n3012 gnd.n3011 585
R8283 gnd.n2602 gnd.n1494 585
R8284 gnd.n4848 gnd.n1494 585
R8285 gnd.n2975 gnd.n2974 585
R8286 gnd.n2974 gnd.n2973 585
R8287 gnd.n2622 gnd.n1483 585
R8288 gnd.n4854 gnd.n1483 585
R8289 gnd.n2979 gnd.n2621 585
R8290 gnd.n2964 gnd.n2621 585
R8291 gnd.n2980 gnd.n1474 585
R8292 gnd.n4860 gnd.n1474 585
R8293 gnd.n2981 gnd.n2620 585
R8294 gnd.n2959 gnd.n2620 585
R8295 gnd.n2617 gnd.n1463 585
R8296 gnd.n4866 gnd.n1463 585
R8297 gnd.n2986 gnd.n2985 585
R8298 gnd.n2987 gnd.n2986 585
R8299 gnd.n2616 gnd.n1454 585
R8300 gnd.n4872 gnd.n1454 585
R8301 gnd.n2951 gnd.n2950 585
R8302 gnd.n2952 gnd.n2951 585
R8303 gnd.n2625 gnd.n1443 585
R8304 gnd.n4878 gnd.n1443 585
R8305 gnd.n2946 gnd.n2945 585
R8306 gnd.n2945 gnd.n2944 585
R8307 gnd.n2627 gnd.n1434 585
R8308 gnd.n4884 gnd.n1434 585
R8309 gnd.n2937 gnd.n2936 585
R8310 gnd.n2938 gnd.n2937 585
R8311 gnd.n2631 gnd.n1424 585
R8312 gnd.n4890 gnd.n1424 585
R8313 gnd.n2932 gnd.n2931 585
R8314 gnd.n2931 gnd.n2930 585
R8315 gnd.n2633 gnd.n1413 585
R8316 gnd.n4896 gnd.n1413 585
R8317 gnd.n2898 gnd.n2897 585
R8318 gnd.n2899 gnd.n2898 585
R8319 gnd.n2644 gnd.n2643 585
R8320 gnd.n2643 gnd.n2641 585
R8321 gnd.n2893 gnd.n2892 585
R8322 gnd.n2892 gnd.n2891 585
R8323 gnd.n2647 gnd.n2646 585
R8324 gnd.n2885 gnd.n2647 585
R8325 gnd.n2868 gnd.n2867 585
R8326 gnd.n2869 gnd.n2868 585
R8327 gnd.n2728 gnd.n2727 585
R8328 gnd.n2727 gnd.n2726 585
R8329 gnd.n2863 gnd.n2862 585
R8330 gnd.n2862 gnd.n1398 585
R8331 gnd.n2861 gnd.n1397 585
R8332 gnd.n4903 gnd.n1397 585
R8333 gnd.n2860 gnd.n2859 585
R8334 gnd.n2859 gnd.n1389 585
R8335 gnd.n2730 gnd.n1388 585
R8336 gnd.n4909 gnd.n1388 585
R8337 gnd.n2855 gnd.n2854 585
R8338 gnd.n2854 gnd.n1386 585
R8339 gnd.n2853 gnd.n1379 585
R8340 gnd.n4915 gnd.n1379 585
R8341 gnd.n2852 gnd.n2851 585
R8342 gnd.n2851 gnd.n1371 585
R8343 gnd.n2732 gnd.n1370 585
R8344 gnd.n4921 gnd.n1370 585
R8345 gnd.n2847 gnd.n2846 585
R8346 gnd.n2846 gnd.n1361 585
R8347 gnd.n2845 gnd.n1360 585
R8348 gnd.n4927 gnd.n1360 585
R8349 gnd.n2844 gnd.n2843 585
R8350 gnd.n2843 gnd.n1352 585
R8351 gnd.n2734 gnd.n1351 585
R8352 gnd.n4933 gnd.n1351 585
R8353 gnd.n2839 gnd.n2838 585
R8354 gnd.n2838 gnd.n1349 585
R8355 gnd.n2837 gnd.n1341 585
R8356 gnd.n4939 gnd.n1341 585
R8357 gnd.n2836 gnd.n2835 585
R8358 gnd.n2835 gnd.n1333 585
R8359 gnd.n2736 gnd.n1332 585
R8360 gnd.n4945 gnd.n1332 585
R8361 gnd.n2831 gnd.n2830 585
R8362 gnd.n2830 gnd.n1323 585
R8363 gnd.n2829 gnd.n1322 585
R8364 gnd.n4951 gnd.n1322 585
R8365 gnd.n2828 gnd.n2827 585
R8366 gnd.n2827 gnd.n1314 585
R8367 gnd.n2738 gnd.n1313 585
R8368 gnd.n4957 gnd.n1313 585
R8369 gnd.n2823 gnd.n2822 585
R8370 gnd.n2822 gnd.n1311 585
R8371 gnd.n2821 gnd.n1303 585
R8372 gnd.n4963 gnd.n1303 585
R8373 gnd.n2820 gnd.n2819 585
R8374 gnd.n2819 gnd.n1295 585
R8375 gnd.n2740 gnd.n1294 585
R8376 gnd.n4969 gnd.n1294 585
R8377 gnd.n2815 gnd.n2814 585
R8378 gnd.n2814 gnd.n1285 585
R8379 gnd.n2813 gnd.n1284 585
R8380 gnd.n4975 gnd.n1284 585
R8381 gnd.n2812 gnd.n2811 585
R8382 gnd.n2811 gnd.n1273 585
R8383 gnd.n2742 gnd.n1272 585
R8384 gnd.n4981 gnd.n1272 585
R8385 gnd.n2807 gnd.n2806 585
R8386 gnd.n2806 gnd.n1270 585
R8387 gnd.n2805 gnd.n1260 585
R8388 gnd.n4987 gnd.n1260 585
R8389 gnd.n2804 gnd.n2803 585
R8390 gnd.n2803 gnd.n1186 585
R8391 gnd.n6574 gnd.n6573 585
R8392 gnd.n6575 gnd.n6574 585
R8393 gnd.n1123 gnd.n1121 585
R8394 gnd.n6514 gnd.n1121 585
R8395 gnd.n6418 gnd.n5133 585
R8396 gnd.n5133 gnd.n5123 585
R8397 gnd.n6420 gnd.n6419 585
R8398 gnd.n6421 gnd.n6420 585
R8399 gnd.n5134 gnd.n5132 585
R8400 gnd.n5142 gnd.n5132 585
R8401 gnd.n6393 gnd.n5154 585
R8402 gnd.n5154 gnd.n5141 585
R8403 gnd.n6395 gnd.n6394 585
R8404 gnd.n6396 gnd.n6395 585
R8405 gnd.n5155 gnd.n5153 585
R8406 gnd.n5153 gnd.n5149 585
R8407 gnd.n6125 gnd.n6124 585
R8408 gnd.n6124 gnd.n6123 585
R8409 gnd.n5160 gnd.n5159 585
R8410 gnd.n6094 gnd.n5160 585
R8411 gnd.n6114 gnd.n6113 585
R8412 gnd.n6113 gnd.n6112 585
R8413 gnd.n5167 gnd.n5166 585
R8414 gnd.n6100 gnd.n5167 585
R8415 gnd.n6073 gnd.n5187 585
R8416 gnd.n5187 gnd.n5176 585
R8417 gnd.n6075 gnd.n6074 585
R8418 gnd.n6076 gnd.n6075 585
R8419 gnd.n5188 gnd.n5186 585
R8420 gnd.n5196 gnd.n5186 585
R8421 gnd.n6051 gnd.n5207 585
R8422 gnd.n5207 gnd.n5195 585
R8423 gnd.n6053 gnd.n6052 585
R8424 gnd.n6054 gnd.n6053 585
R8425 gnd.n5208 gnd.n5206 585
R8426 gnd.n6035 gnd.n5206 585
R8427 gnd.n6039 gnd.n6038 585
R8428 gnd.n6038 gnd.n6037 585
R8429 gnd.n5213 gnd.n5212 585
R8430 gnd.n6022 gnd.n5213 585
R8431 gnd.n6007 gnd.n5234 585
R8432 gnd.n5234 gnd.n5221 585
R8433 gnd.n6009 gnd.n6008 585
R8434 gnd.n6010 gnd.n6009 585
R8435 gnd.n5235 gnd.n5233 585
R8436 gnd.n5233 gnd.n5229 585
R8437 gnd.n5994 gnd.n5993 585
R8438 gnd.n5993 gnd.n5992 585
R8439 gnd.n5242 gnd.n5241 585
R8440 gnd.n5252 gnd.n5242 585
R8441 gnd.n5983 gnd.n5982 585
R8442 gnd.n5982 gnd.n5981 585
R8443 gnd.n5249 gnd.n5248 585
R8444 gnd.n5969 gnd.n5249 585
R8445 gnd.n5946 gnd.n5350 585
R8446 gnd.n5350 gnd.n5259 585
R8447 gnd.n5948 gnd.n5947 585
R8448 gnd.n5949 gnd.n5948 585
R8449 gnd.n5351 gnd.n5349 585
R8450 gnd.n5359 gnd.n5349 585
R8451 gnd.n5924 gnd.n5371 585
R8452 gnd.n5371 gnd.n5358 585
R8453 gnd.n5926 gnd.n5925 585
R8454 gnd.n5927 gnd.n5926 585
R8455 gnd.n5372 gnd.n5370 585
R8456 gnd.n5370 gnd.n5366 585
R8457 gnd.n5912 gnd.n5911 585
R8458 gnd.n5911 gnd.n5910 585
R8459 gnd.n5377 gnd.n5376 585
R8460 gnd.n5386 gnd.n5377 585
R8461 gnd.n5901 gnd.n5900 585
R8462 gnd.n5900 gnd.n5899 585
R8463 gnd.n5384 gnd.n5383 585
R8464 gnd.n5887 gnd.n5384 585
R8465 gnd.n5859 gnd.n5858 585
R8466 gnd.n5858 gnd.n5393 585
R8467 gnd.n5860 gnd.n5404 585
R8468 gnd.n5851 gnd.n5404 585
R8469 gnd.n5862 gnd.n5861 585
R8470 gnd.n5863 gnd.n5862 585
R8471 gnd.n5405 gnd.n5403 585
R8472 gnd.n5419 gnd.n5403 585
R8473 gnd.n5843 gnd.n5842 585
R8474 gnd.n5842 gnd.n5841 585
R8475 gnd.n5416 gnd.n5415 585
R8476 gnd.n5826 gnd.n5416 585
R8477 gnd.n5813 gnd.n5436 585
R8478 gnd.n5436 gnd.n5426 585
R8479 gnd.n5815 gnd.n5814 585
R8480 gnd.n5816 gnd.n5815 585
R8481 gnd.n5437 gnd.n5435 585
R8482 gnd.n5445 gnd.n5435 585
R8483 gnd.n5789 gnd.n5457 585
R8484 gnd.n5457 gnd.n5444 585
R8485 gnd.n5791 gnd.n5790 585
R8486 gnd.n5792 gnd.n5791 585
R8487 gnd.n5458 gnd.n5456 585
R8488 gnd.n5456 gnd.n5452 585
R8489 gnd.n5777 gnd.n5776 585
R8490 gnd.n5776 gnd.n5775 585
R8491 gnd.n5463 gnd.n5462 585
R8492 gnd.n5467 gnd.n5463 585
R8493 gnd.n5761 gnd.n5760 585
R8494 gnd.n5762 gnd.n5761 585
R8495 gnd.n5478 gnd.n5477 585
R8496 gnd.n5477 gnd.n5473 585
R8497 gnd.n5751 gnd.n5750 585
R8498 gnd.n5752 gnd.n5751 585
R8499 gnd.n5487 gnd.n5486 585
R8500 gnd.n5486 gnd.n5484 585
R8501 gnd.n5745 gnd.n5744 585
R8502 gnd.n5744 gnd.n5743 585
R8503 gnd.n5491 gnd.n5490 585
R8504 gnd.n5499 gnd.n5491 585
R8505 gnd.n5652 gnd.n5651 585
R8506 gnd.n5653 gnd.n5652 585
R8507 gnd.n5501 gnd.n5500 585
R8508 gnd.n5500 gnd.n5498 585
R8509 gnd.n5647 gnd.n5646 585
R8510 gnd.n5646 gnd.n5645 585
R8511 gnd.n5504 gnd.n5503 585
R8512 gnd.n5505 gnd.n5504 585
R8513 gnd.n5636 gnd.n5635 585
R8514 gnd.n5637 gnd.n5636 585
R8515 gnd.n5513 gnd.n5512 585
R8516 gnd.n5512 gnd.n5511 585
R8517 gnd.n5631 gnd.n5630 585
R8518 gnd.n5630 gnd.n5629 585
R8519 gnd.n5516 gnd.n5515 585
R8520 gnd.n5517 gnd.n5516 585
R8521 gnd.n5620 gnd.n5619 585
R8522 gnd.n5621 gnd.n5620 585
R8523 gnd.n5616 gnd.n5523 585
R8524 gnd.n5615 gnd.n5614 585
R8525 gnd.n5612 gnd.n5525 585
R8526 gnd.n5612 gnd.n5522 585
R8527 gnd.n5611 gnd.n5610 585
R8528 gnd.n5609 gnd.n5608 585
R8529 gnd.n5607 gnd.n5530 585
R8530 gnd.n5605 gnd.n5604 585
R8531 gnd.n5603 gnd.n5531 585
R8532 gnd.n5602 gnd.n5601 585
R8533 gnd.n5599 gnd.n5536 585
R8534 gnd.n5597 gnd.n5596 585
R8535 gnd.n5595 gnd.n5537 585
R8536 gnd.n5594 gnd.n5593 585
R8537 gnd.n5591 gnd.n5542 585
R8538 gnd.n5589 gnd.n5588 585
R8539 gnd.n5587 gnd.n5543 585
R8540 gnd.n5586 gnd.n5585 585
R8541 gnd.n5583 gnd.n5548 585
R8542 gnd.n5581 gnd.n5580 585
R8543 gnd.n5579 gnd.n5549 585
R8544 gnd.n5578 gnd.n5577 585
R8545 gnd.n5575 gnd.n5554 585
R8546 gnd.n5573 gnd.n5572 585
R8547 gnd.n5570 gnd.n5555 585
R8548 gnd.n5569 gnd.n5568 585
R8549 gnd.n5566 gnd.n5564 585
R8550 gnd.n5562 gnd.n5521 585
R8551 gnd.n6508 gnd.n6507 585
R8552 gnd.n6506 gnd.n6505 585
R8553 gnd.n6504 gnd.n6503 585
R8554 gnd.n6497 gnd.n6428 585
R8555 gnd.n6499 gnd.n6498 585
R8556 gnd.n6493 gnd.n6492 585
R8557 gnd.n6491 gnd.n6490 585
R8558 gnd.n6484 gnd.n6430 585
R8559 gnd.n6486 gnd.n6485 585
R8560 gnd.n6483 gnd.n6482 585
R8561 gnd.n6481 gnd.n6480 585
R8562 gnd.n6474 gnd.n6432 585
R8563 gnd.n6476 gnd.n6475 585
R8564 gnd.n6473 gnd.n6472 585
R8565 gnd.n6471 gnd.n6470 585
R8566 gnd.n6464 gnd.n6434 585
R8567 gnd.n6466 gnd.n6465 585
R8568 gnd.n6463 gnd.n6462 585
R8569 gnd.n6461 gnd.n6460 585
R8570 gnd.n6454 gnd.n6436 585
R8571 gnd.n6456 gnd.n6455 585
R8572 gnd.n6453 gnd.n6452 585
R8573 gnd.n6451 gnd.n6450 585
R8574 gnd.n6444 gnd.n6438 585
R8575 gnd.n6446 gnd.n6445 585
R8576 gnd.n6443 gnd.n6442 585
R8577 gnd.n6441 gnd.n1122 585
R8578 gnd.n6559 gnd.n1122 585
R8579 gnd.n6511 gnd.n1119 585
R8580 gnd.n6575 gnd.n1119 585
R8581 gnd.n6513 gnd.n6512 585
R8582 gnd.n6514 gnd.n6513 585
R8583 gnd.n5126 gnd.n5125 585
R8584 gnd.n5125 gnd.n5123 585
R8585 gnd.n6423 gnd.n6422 585
R8586 gnd.n6422 gnd.n6421 585
R8587 gnd.n5129 gnd.n5128 585
R8588 gnd.n5142 gnd.n5129 585
R8589 gnd.n6089 gnd.n6088 585
R8590 gnd.n6088 gnd.n5141 585
R8591 gnd.n6090 gnd.n5151 585
R8592 gnd.n6396 gnd.n5151 585
R8593 gnd.n6092 gnd.n6091 585
R8594 gnd.n6091 gnd.n5149 585
R8595 gnd.n6093 gnd.n5162 585
R8596 gnd.n6123 gnd.n5162 585
R8597 gnd.n6096 gnd.n6095 585
R8598 gnd.n6095 gnd.n6094 585
R8599 gnd.n6097 gnd.n5169 585
R8600 gnd.n6112 gnd.n5169 585
R8601 gnd.n6099 gnd.n6098 585
R8602 gnd.n6100 gnd.n6099 585
R8603 gnd.n5180 gnd.n5179 585
R8604 gnd.n5179 gnd.n5176 585
R8605 gnd.n6078 gnd.n6077 585
R8606 gnd.n6077 gnd.n6076 585
R8607 gnd.n5183 gnd.n5182 585
R8608 gnd.n5196 gnd.n5183 585
R8609 gnd.n6031 gnd.n6030 585
R8610 gnd.n6030 gnd.n5195 585
R8611 gnd.n6032 gnd.n5204 585
R8612 gnd.n6054 gnd.n5204 585
R8613 gnd.n6034 gnd.n6033 585
R8614 gnd.n6035 gnd.n6034 585
R8615 gnd.n5217 gnd.n5215 585
R8616 gnd.n6037 gnd.n5215 585
R8617 gnd.n6024 gnd.n6023 585
R8618 gnd.n6023 gnd.n6022 585
R8619 gnd.n5220 gnd.n5219 585
R8620 gnd.n5221 gnd.n5220 585
R8621 gnd.n5960 gnd.n5231 585
R8622 gnd.n6010 gnd.n5231 585
R8623 gnd.n5962 gnd.n5961 585
R8624 gnd.n5961 gnd.n5229 585
R8625 gnd.n5963 gnd.n5244 585
R8626 gnd.n5992 gnd.n5244 585
R8627 gnd.n5965 gnd.n5964 585
R8628 gnd.n5964 gnd.n5252 585
R8629 gnd.n5966 gnd.n5251 585
R8630 gnd.n5981 gnd.n5251 585
R8631 gnd.n5968 gnd.n5967 585
R8632 gnd.n5969 gnd.n5968 585
R8633 gnd.n5263 gnd.n5262 585
R8634 gnd.n5262 gnd.n5259 585
R8635 gnd.n5951 gnd.n5950 585
R8636 gnd.n5950 gnd.n5949 585
R8637 gnd.n5346 gnd.n5345 585
R8638 gnd.n5359 gnd.n5346 585
R8639 gnd.n5872 gnd.n5871 585
R8640 gnd.n5871 gnd.n5358 585
R8641 gnd.n5873 gnd.n5368 585
R8642 gnd.n5927 gnd.n5368 585
R8643 gnd.n5876 gnd.n5875 585
R8644 gnd.n5875 gnd.n5366 585
R8645 gnd.n5877 gnd.n5379 585
R8646 gnd.n5910 gnd.n5379 585
R8647 gnd.n5880 gnd.n5879 585
R8648 gnd.n5879 gnd.n5386 585
R8649 gnd.n5881 gnd.n5385 585
R8650 gnd.n5899 gnd.n5385 585
R8651 gnd.n5884 gnd.n5883 585
R8652 gnd.n5887 gnd.n5884 585
R8653 gnd.n5869 gnd.n5395 585
R8654 gnd.n5395 gnd.n5393 585
R8655 gnd.n5400 gnd.n5396 585
R8656 gnd.n5851 gnd.n5400 585
R8657 gnd.n5865 gnd.n5864 585
R8658 gnd.n5864 gnd.n5863 585
R8659 gnd.n5399 gnd.n5398 585
R8660 gnd.n5419 gnd.n5399 585
R8661 gnd.n5823 gnd.n5418 585
R8662 gnd.n5841 gnd.n5418 585
R8663 gnd.n5825 gnd.n5824 585
R8664 gnd.n5826 gnd.n5825 585
R8665 gnd.n5429 gnd.n5428 585
R8666 gnd.n5428 gnd.n5426 585
R8667 gnd.n5818 gnd.n5817 585
R8668 gnd.n5817 gnd.n5816 585
R8669 gnd.n5432 gnd.n5431 585
R8670 gnd.n5445 gnd.n5432 585
R8671 gnd.n5669 gnd.n5668 585
R8672 gnd.n5668 gnd.n5444 585
R8673 gnd.n5670 gnd.n5454 585
R8674 gnd.n5792 gnd.n5454 585
R8675 gnd.n5672 gnd.n5671 585
R8676 gnd.n5671 gnd.n5452 585
R8677 gnd.n5673 gnd.n5464 585
R8678 gnd.n5775 gnd.n5464 585
R8679 gnd.n5675 gnd.n5674 585
R8680 gnd.n5674 gnd.n5467 585
R8681 gnd.n5676 gnd.n5475 585
R8682 gnd.n5762 gnd.n5475 585
R8683 gnd.n5678 gnd.n5677 585
R8684 gnd.n5677 gnd.n5473 585
R8685 gnd.n5679 gnd.n5485 585
R8686 gnd.n5752 gnd.n5485 585
R8687 gnd.n5680 gnd.n5493 585
R8688 gnd.n5493 gnd.n5484 585
R8689 gnd.n5682 gnd.n5681 585
R8690 gnd.n5743 gnd.n5682 585
R8691 gnd.n5494 gnd.n5492 585
R8692 gnd.n5499 gnd.n5492 585
R8693 gnd.n5655 gnd.n5654 585
R8694 gnd.n5654 gnd.n5653 585
R8695 gnd.n5497 gnd.n5496 585
R8696 gnd.n5498 gnd.n5497 585
R8697 gnd.n5644 gnd.n5643 585
R8698 gnd.n5645 gnd.n5644 585
R8699 gnd.n5507 gnd.n5506 585
R8700 gnd.n5506 gnd.n5505 585
R8701 gnd.n5639 gnd.n5638 585
R8702 gnd.n5638 gnd.n5637 585
R8703 gnd.n5510 gnd.n5509 585
R8704 gnd.n5511 gnd.n5510 585
R8705 gnd.n5628 gnd.n5627 585
R8706 gnd.n5629 gnd.n5628 585
R8707 gnd.n5519 gnd.n5518 585
R8708 gnd.n5518 gnd.n5517 585
R8709 gnd.n5623 gnd.n5622 585
R8710 gnd.n5622 gnd.n5621 585
R8711 gnd.n241 gnd.n240 585
R8712 gnd.n244 gnd.n241 585
R8713 gnd.n7673 gnd.n7672 585
R8714 gnd.n7672 gnd.n7671 585
R8715 gnd.n7674 gnd.n236 585
R8716 gnd.n236 gnd.n235 585
R8717 gnd.n7676 gnd.n7675 585
R8718 gnd.n7677 gnd.n7676 585
R8719 gnd.n221 gnd.n220 585
R8720 gnd.n225 gnd.n221 585
R8721 gnd.n7685 gnd.n7684 585
R8722 gnd.n7684 gnd.n7683 585
R8723 gnd.n7686 gnd.n216 585
R8724 gnd.n222 gnd.n216 585
R8725 gnd.n7688 gnd.n7687 585
R8726 gnd.n7689 gnd.n7688 585
R8727 gnd.n203 gnd.n202 585
R8728 gnd.n206 gnd.n203 585
R8729 gnd.n7697 gnd.n7696 585
R8730 gnd.n7696 gnd.n7695 585
R8731 gnd.n7698 gnd.n198 585
R8732 gnd.n198 gnd.n197 585
R8733 gnd.n7700 gnd.n7699 585
R8734 gnd.n7701 gnd.n7700 585
R8735 gnd.n183 gnd.n182 585
R8736 gnd.n194 gnd.n183 585
R8737 gnd.n7709 gnd.n7708 585
R8738 gnd.n7708 gnd.n7707 585
R8739 gnd.n7710 gnd.n178 585
R8740 gnd.n184 gnd.n178 585
R8741 gnd.n7712 gnd.n7711 585
R8742 gnd.n7713 gnd.n7712 585
R8743 gnd.n165 gnd.n164 585
R8744 gnd.n168 gnd.n165 585
R8745 gnd.n7721 gnd.n7720 585
R8746 gnd.n7720 gnd.n7719 585
R8747 gnd.n7722 gnd.n160 585
R8748 gnd.n160 gnd.n159 585
R8749 gnd.n7724 gnd.n7723 585
R8750 gnd.n7725 gnd.n7724 585
R8751 gnd.n145 gnd.n144 585
R8752 gnd.n156 gnd.n145 585
R8753 gnd.n7733 gnd.n7732 585
R8754 gnd.n7732 gnd.n7731 585
R8755 gnd.n7734 gnd.n140 585
R8756 gnd.n146 gnd.n140 585
R8757 gnd.n7736 gnd.n7735 585
R8758 gnd.n7737 gnd.n7736 585
R8759 gnd.n128 gnd.n127 585
R8760 gnd.n131 gnd.n128 585
R8761 gnd.n7745 gnd.n7744 585
R8762 gnd.n7744 gnd.n7743 585
R8763 gnd.n7746 gnd.n122 585
R8764 gnd.n122 gnd.n120 585
R8765 gnd.n7748 gnd.n7747 585
R8766 gnd.n7749 gnd.n7748 585
R8767 gnd.n123 gnd.n121 585
R8768 gnd.n121 gnd.n117 585
R8769 gnd.n7487 gnd.n7486 585
R8770 gnd.n7486 gnd.n102 585
R8771 gnd.n7485 gnd.n103 585
R8772 gnd.n7757 gnd.n103 585
R8773 gnd.n7484 gnd.n7483 585
R8774 gnd.n7483 gnd.n7482 585
R8775 gnd.n484 gnd.n482 585
R8776 gnd.n485 gnd.n484 585
R8777 gnd.n7475 gnd.n7474 585
R8778 gnd.n7474 gnd.n7473 585
R8779 gnd.n490 gnd.n489 585
R8780 gnd.n7465 gnd.n490 585
R8781 gnd.n7448 gnd.n7447 585
R8782 gnd.n7447 gnd.n7446 585
R8783 gnd.n7449 gnd.n506 585
R8784 gnd.n7457 gnd.n506 585
R8785 gnd.n7451 gnd.n7450 585
R8786 gnd.n7452 gnd.n7451 585
R8787 gnd.n512 gnd.n511 585
R8788 gnd.n7438 gnd.n511 585
R8789 gnd.n7414 gnd.n7413 585
R8790 gnd.n7413 gnd.n7412 585
R8791 gnd.n7415 gnd.n529 585
R8792 gnd.n7430 gnd.n529 585
R8793 gnd.n7416 gnd.n541 585
R8794 gnd.n7406 gnd.n541 585
R8795 gnd.n7418 gnd.n7417 585
R8796 gnd.n7419 gnd.n7418 585
R8797 gnd.n542 gnd.n540 585
R8798 gnd.n7402 gnd.n540 585
R8799 gnd.n7378 gnd.n7377 585
R8800 gnd.n7377 gnd.n7376 585
R8801 gnd.n7379 gnd.n558 585
R8802 gnd.n7393 gnd.n558 585
R8803 gnd.n7380 gnd.n569 585
R8804 gnd.n7370 gnd.n569 585
R8805 gnd.n7382 gnd.n7381 585
R8806 gnd.n7383 gnd.n7382 585
R8807 gnd.n570 gnd.n568 585
R8808 gnd.n2055 gnd.n568 585
R8809 gnd.n2048 gnd.n2047 585
R8810 gnd.n4328 gnd.n2048 585
R8811 gnd.n4338 gnd.n4337 585
R8812 gnd.n4337 gnd.n4336 585
R8813 gnd.n4339 gnd.n2043 585
R8814 gnd.n4316 gnd.n2043 585
R8815 gnd.n4341 gnd.n4340 585
R8816 gnd.n4342 gnd.n4341 585
R8817 gnd.n2028 gnd.n2027 585
R8818 gnd.n4300 gnd.n2028 585
R8819 gnd.n4350 gnd.n4349 585
R8820 gnd.n4349 gnd.n4348 585
R8821 gnd.n4351 gnd.n2023 585
R8822 gnd.n4285 gnd.n2023 585
R8823 gnd.n4353 gnd.n4352 585
R8824 gnd.n4354 gnd.n4353 585
R8825 gnd.n2007 gnd.n2006 585
R8826 gnd.n4277 gnd.n2007 585
R8827 gnd.n4362 gnd.n4361 585
R8828 gnd.n4361 gnd.n4360 585
R8829 gnd.n4363 gnd.n2000 585
R8830 gnd.n4270 gnd.n2000 585
R8831 gnd.n4365 gnd.n4364 585
R8832 gnd.n4366 gnd.n4365 585
R8833 gnd.n2001 gnd.n1999 585
R8834 gnd.n4262 gnd.n1999 585
R8835 gnd.n1983 gnd.n1977 585
R8836 gnd.n4372 gnd.n1983 585
R8837 gnd.n4377 gnd.n1975 585
R8838 gnd.n4238 gnd.n1975 585
R8839 gnd.n4379 gnd.n4378 585
R8840 gnd.n4380 gnd.n4379 585
R8841 gnd.n1974 gnd.n1814 585
R8842 gnd.n4547 gnd.n1815 585
R8843 gnd.n4546 gnd.n1816 585
R8844 gnd.n1891 gnd.n1817 585
R8845 gnd.n4539 gnd.n1823 585
R8846 gnd.n4538 gnd.n1824 585
R8847 gnd.n1894 gnd.n1825 585
R8848 gnd.n4531 gnd.n1831 585
R8849 gnd.n4530 gnd.n1832 585
R8850 gnd.n1896 gnd.n1833 585
R8851 gnd.n4523 gnd.n1839 585
R8852 gnd.n4522 gnd.n1840 585
R8853 gnd.n1899 gnd.n1841 585
R8854 gnd.n4515 gnd.n1847 585
R8855 gnd.n4514 gnd.n1848 585
R8856 gnd.n1901 gnd.n1849 585
R8857 gnd.n4507 gnd.n1857 585
R8858 gnd.n4506 gnd.n4503 585
R8859 gnd.n1860 gnd.n1858 585
R8860 gnd.n4501 gnd.n1860 585
R8861 gnd.n439 gnd.n365 585
R8862 gnd.n446 gnd.n445 585
R8863 gnd.n448 gnd.n447 585
R8864 gnd.n450 gnd.n449 585
R8865 gnd.n452 gnd.n451 585
R8866 gnd.n454 gnd.n453 585
R8867 gnd.n456 gnd.n455 585
R8868 gnd.n458 gnd.n457 585
R8869 gnd.n460 gnd.n459 585
R8870 gnd.n462 gnd.n461 585
R8871 gnd.n464 gnd.n463 585
R8872 gnd.n466 gnd.n465 585
R8873 gnd.n468 gnd.n467 585
R8874 gnd.n470 gnd.n469 585
R8875 gnd.n472 gnd.n471 585
R8876 gnd.n474 gnd.n473 585
R8877 gnd.n476 gnd.n475 585
R8878 gnd.n477 gnd.n349 585
R8879 gnd.n478 gnd.n251 585
R8880 gnd.n7663 gnd.n251 585
R8881 gnd.n441 gnd.n440 585
R8882 gnd.n440 gnd.n244 585
R8883 gnd.n438 gnd.n243 585
R8884 gnd.n7671 gnd.n243 585
R8885 gnd.n437 gnd.n436 585
R8886 gnd.n436 gnd.n235 585
R8887 gnd.n369 gnd.n234 585
R8888 gnd.n7677 gnd.n234 585
R8889 gnd.n432 gnd.n431 585
R8890 gnd.n431 gnd.n225 585
R8891 gnd.n430 gnd.n224 585
R8892 gnd.n7683 gnd.n224 585
R8893 gnd.n429 gnd.n428 585
R8894 gnd.n428 gnd.n222 585
R8895 gnd.n371 gnd.n215 585
R8896 gnd.n7689 gnd.n215 585
R8897 gnd.n424 gnd.n423 585
R8898 gnd.n423 gnd.n206 585
R8899 gnd.n422 gnd.n205 585
R8900 gnd.n7695 gnd.n205 585
R8901 gnd.n421 gnd.n420 585
R8902 gnd.n420 gnd.n197 585
R8903 gnd.n373 gnd.n196 585
R8904 gnd.n7701 gnd.n196 585
R8905 gnd.n416 gnd.n415 585
R8906 gnd.n415 gnd.n194 585
R8907 gnd.n414 gnd.n186 585
R8908 gnd.n7707 gnd.n186 585
R8909 gnd.n413 gnd.n412 585
R8910 gnd.n412 gnd.n184 585
R8911 gnd.n375 gnd.n177 585
R8912 gnd.n7713 gnd.n177 585
R8913 gnd.n408 gnd.n407 585
R8914 gnd.n407 gnd.n168 585
R8915 gnd.n406 gnd.n167 585
R8916 gnd.n7719 gnd.n167 585
R8917 gnd.n405 gnd.n404 585
R8918 gnd.n404 gnd.n159 585
R8919 gnd.n377 gnd.n158 585
R8920 gnd.n7725 gnd.n158 585
R8921 gnd.n400 gnd.n399 585
R8922 gnd.n399 gnd.n156 585
R8923 gnd.n398 gnd.n148 585
R8924 gnd.n7731 gnd.n148 585
R8925 gnd.n397 gnd.n396 585
R8926 gnd.n396 gnd.n146 585
R8927 gnd.n379 gnd.n139 585
R8928 gnd.n7737 gnd.n139 585
R8929 gnd.n392 gnd.n391 585
R8930 gnd.n391 gnd.n131 585
R8931 gnd.n390 gnd.n130 585
R8932 gnd.n7743 gnd.n130 585
R8933 gnd.n389 gnd.n388 585
R8934 gnd.n388 gnd.n120 585
R8935 gnd.n381 gnd.n119 585
R8936 gnd.n7749 gnd.n119 585
R8937 gnd.n384 gnd.n383 585
R8938 gnd.n383 gnd.n117 585
R8939 gnd.n100 gnd.n99 585
R8940 gnd.n102 gnd.n100 585
R8941 gnd.n7759 gnd.n7758 585
R8942 gnd.n7758 gnd.n7757 585
R8943 gnd.n7760 gnd.n98 585
R8944 gnd.n7482 gnd.n98 585
R8945 gnd.n492 gnd.n96 585
R8946 gnd.n492 gnd.n485 585
R8947 gnd.n500 gnd.n493 585
R8948 gnd.n7473 gnd.n493 585
R8949 gnd.n7464 gnd.n7463 585
R8950 gnd.n7465 gnd.n7464 585
R8951 gnd.n499 gnd.n498 585
R8952 gnd.n7446 gnd.n498 585
R8953 gnd.n7459 gnd.n7458 585
R8954 gnd.n7458 gnd.n7457 585
R8955 gnd.n503 gnd.n502 585
R8956 gnd.n7452 gnd.n503 585
R8957 gnd.n7437 gnd.n7436 585
R8958 gnd.n7438 gnd.n7437 585
R8959 gnd.n522 gnd.n521 585
R8960 gnd.n7412 gnd.n521 585
R8961 gnd.n7432 gnd.n7431 585
R8962 gnd.n7431 gnd.n7430 585
R8963 gnd.n525 gnd.n524 585
R8964 gnd.n7406 gnd.n525 585
R8965 gnd.n551 gnd.n538 585
R8966 gnd.n7419 gnd.n538 585
R8967 gnd.n7401 gnd.n7400 585
R8968 gnd.n7402 gnd.n7401 585
R8969 gnd.n550 gnd.n549 585
R8970 gnd.n7376 gnd.n549 585
R8971 gnd.n7395 gnd.n7394 585
R8972 gnd.n7394 gnd.n7393 585
R8973 gnd.n554 gnd.n553 585
R8974 gnd.n7370 gnd.n554 585
R8975 gnd.n4308 gnd.n567 585
R8976 gnd.n7383 gnd.n567 585
R8977 gnd.n4309 gnd.n4306 585
R8978 gnd.n4306 gnd.n2055 585
R8979 gnd.n4310 gnd.n2054 585
R8980 gnd.n4328 gnd.n2054 585
R8981 gnd.n2063 gnd.n2051 585
R8982 gnd.n4336 gnd.n2051 585
R8983 gnd.n4315 gnd.n4314 585
R8984 gnd.n4316 gnd.n4315 585
R8985 gnd.n2062 gnd.n2042 585
R8986 gnd.n4342 gnd.n2042 585
R8987 gnd.n4302 gnd.n4301 585
R8988 gnd.n4301 gnd.n4300 585
R8989 gnd.n2065 gnd.n2031 585
R8990 gnd.n4348 gnd.n2031 585
R8991 gnd.n4284 gnd.n4283 585
R8992 gnd.n4285 gnd.n4284 585
R8993 gnd.n2067 gnd.n2021 585
R8994 gnd.n4354 gnd.n2021 585
R8995 gnd.n4279 gnd.n4278 585
R8996 gnd.n4278 gnd.n4277 585
R8997 gnd.n2069 gnd.n2010 585
R8998 gnd.n4360 gnd.n2010 585
R8999 gnd.n4269 gnd.n4268 585
R9000 gnd.n4270 gnd.n4269 585
R9001 gnd.n2071 gnd.n1997 585
R9002 gnd.n4366 gnd.n1997 585
R9003 gnd.n4264 gnd.n4263 585
R9004 gnd.n4263 gnd.n4262 585
R9005 gnd.n4261 gnd.n1981 585
R9006 gnd.n4372 gnd.n1981 585
R9007 gnd.n4260 gnd.n2074 585
R9008 gnd.n4238 gnd.n2074 585
R9009 gnd.n2073 gnd.n1972 585
R9010 gnd.n4380 gnd.n1972 585
R9011 gnd.n6519 gnd.n5118 585
R9012 gnd.n5118 gnd.n1120 585
R9013 gnd.n6518 gnd.n6517 585
R9014 gnd.n6517 gnd.n1118 585
R9015 gnd.n6516 gnd.n5121 585
R9016 gnd.n6516 gnd.n6515 585
R9017 gnd.n6406 gnd.n5122 585
R9018 gnd.n5131 gnd.n5122 585
R9019 gnd.n6407 gnd.n5144 585
R9020 gnd.n5144 gnd.n5130 585
R9021 gnd.n6409 gnd.n6408 585
R9022 gnd.n6410 gnd.n6409 585
R9023 gnd.n5145 gnd.n5143 585
R9024 gnd.n5152 gnd.n5143 585
R9025 gnd.n6399 gnd.n6398 585
R9026 gnd.n6398 gnd.n6397 585
R9027 gnd.n5148 gnd.n5147 585
R9028 gnd.n6122 gnd.n5148 585
R9029 gnd.n6108 gnd.n5171 585
R9030 gnd.n5171 gnd.n5161 585
R9031 gnd.n6110 gnd.n6109 585
R9032 gnd.n6111 gnd.n6110 585
R9033 gnd.n5172 gnd.n5170 585
R9034 gnd.n5170 gnd.n5168 585
R9035 gnd.n6103 gnd.n6102 585
R9036 gnd.n6102 gnd.n6101 585
R9037 gnd.n5175 gnd.n5174 585
R9038 gnd.n5185 gnd.n5175 585
R9039 gnd.n6062 gnd.n5198 585
R9040 gnd.n5198 gnd.n5184 585
R9041 gnd.n6064 gnd.n6063 585
R9042 gnd.n6065 gnd.n6064 585
R9043 gnd.n5199 gnd.n5197 585
R9044 gnd.n5205 gnd.n5197 585
R9045 gnd.n6057 gnd.n6056 585
R9046 gnd.n6056 gnd.n6055 585
R9047 gnd.n5202 gnd.n5201 585
R9048 gnd.n6036 gnd.n5202 585
R9049 gnd.n6018 gnd.n5224 585
R9050 gnd.n5224 gnd.n5214 585
R9051 gnd.n6020 gnd.n6019 585
R9052 gnd.n6021 gnd.n6020 585
R9053 gnd.n5225 gnd.n5223 585
R9054 gnd.n5232 gnd.n5223 585
R9055 gnd.n6013 gnd.n6012 585
R9056 gnd.n6012 gnd.n6011 585
R9057 gnd.n5228 gnd.n5227 585
R9058 gnd.n5991 gnd.n5228 585
R9059 gnd.n5977 gnd.n5254 585
R9060 gnd.n5254 gnd.n5243 585
R9061 gnd.n5979 gnd.n5978 585
R9062 gnd.n5980 gnd.n5979 585
R9063 gnd.n5255 gnd.n5253 585
R9064 gnd.n5253 gnd.n5250 585
R9065 gnd.n5972 gnd.n5971 585
R9066 gnd.n5971 gnd.n5970 585
R9067 gnd.n5258 gnd.n5257 585
R9068 gnd.n5348 gnd.n5258 585
R9069 gnd.n5935 gnd.n5361 585
R9070 gnd.n5361 gnd.n5347 585
R9071 gnd.n5937 gnd.n5936 585
R9072 gnd.n5938 gnd.n5937 585
R9073 gnd.n5362 gnd.n5360 585
R9074 gnd.n5369 gnd.n5360 585
R9075 gnd.n5930 gnd.n5929 585
R9076 gnd.n5929 gnd.n5928 585
R9077 gnd.n5365 gnd.n5364 585
R9078 gnd.n5909 gnd.n5365 585
R9079 gnd.n5895 gnd.n5388 585
R9080 gnd.n5388 gnd.n5378 585
R9081 gnd.n5897 gnd.n5896 585
R9082 gnd.n5898 gnd.n5897 585
R9083 gnd.n5389 gnd.n5387 585
R9084 gnd.n5886 gnd.n5387 585
R9085 gnd.n5890 gnd.n5889 585
R9086 gnd.n5889 gnd.n5888 585
R9087 gnd.n5392 gnd.n5391 585
R9088 gnd.n5852 gnd.n5392 585
R9089 gnd.n5836 gnd.n5835 585
R9090 gnd.n5835 gnd.n5402 585
R9091 gnd.n5837 gnd.n5421 585
R9092 gnd.n5421 gnd.n5401 585
R9093 gnd.n5839 gnd.n5838 585
R9094 gnd.n5840 gnd.n5839 585
R9095 gnd.n5422 gnd.n5420 585
R9096 gnd.n5420 gnd.n5417 585
R9097 gnd.n5829 gnd.n5828 585
R9098 gnd.n5828 gnd.n5827 585
R9099 gnd.n5425 gnd.n5424 585
R9100 gnd.n5434 gnd.n5425 585
R9101 gnd.n5800 gnd.n5447 585
R9102 gnd.n5447 gnd.n5433 585
R9103 gnd.n5802 gnd.n5801 585
R9104 gnd.n5803 gnd.n5802 585
R9105 gnd.n5448 gnd.n5446 585
R9106 gnd.n5455 gnd.n5446 585
R9107 gnd.n5795 gnd.n5794 585
R9108 gnd.n5794 gnd.n5793 585
R9109 gnd.n5451 gnd.n5450 585
R9110 gnd.n5774 gnd.n5451 585
R9111 gnd.n5770 gnd.n5769 585
R9112 gnd.n5771 gnd.n5770 585
R9113 gnd.n5469 gnd.n5468 585
R9114 gnd.n5476 gnd.n5468 585
R9115 gnd.n5765 gnd.n5764 585
R9116 gnd.n5764 gnd.n5763 585
R9117 gnd.n5472 gnd.n5471 585
R9118 gnd.n5753 gnd.n5472 585
R9119 gnd.n5740 gnd.n5739 585
R9120 gnd.n5738 gnd.n5691 585
R9121 gnd.n5737 gnd.n5690 585
R9122 gnd.n5742 gnd.n5690 585
R9123 gnd.n5736 gnd.n5735 585
R9124 gnd.n5734 gnd.n5733 585
R9125 gnd.n5732 gnd.n5731 585
R9126 gnd.n5730 gnd.n5729 585
R9127 gnd.n5728 gnd.n5727 585
R9128 gnd.n5726 gnd.n5725 585
R9129 gnd.n5724 gnd.n5723 585
R9130 gnd.n5722 gnd.n5721 585
R9131 gnd.n5720 gnd.n5719 585
R9132 gnd.n5718 gnd.n5717 585
R9133 gnd.n5716 gnd.n5715 585
R9134 gnd.n5714 gnd.n5713 585
R9135 gnd.n5712 gnd.n5711 585
R9136 gnd.n5707 gnd.n5483 585
R9137 gnd.n6568 gnd.n6567 585
R9138 gnd.n6561 gnd.n1131 585
R9139 gnd.n6563 gnd.n6562 585
R9140 gnd.n1134 gnd.n1133 585
R9141 gnd.n6533 gnd.n6532 585
R9142 gnd.n6535 gnd.n6534 585
R9143 gnd.n6537 gnd.n6536 585
R9144 gnd.n6539 gnd.n6538 585
R9145 gnd.n6541 gnd.n6540 585
R9146 gnd.n6543 gnd.n6542 585
R9147 gnd.n6545 gnd.n6544 585
R9148 gnd.n6547 gnd.n6546 585
R9149 gnd.n6549 gnd.n6548 585
R9150 gnd.n6552 gnd.n6551 585
R9151 gnd.n6550 gnd.n6522 585
R9152 gnd.n6556 gnd.n5119 585
R9153 gnd.n6558 gnd.n6557 585
R9154 gnd.n6559 gnd.n6558 585
R9155 gnd.n6570 gnd.n6569 585
R9156 gnd.n6569 gnd.n1120 585
R9157 gnd.n1127 gnd.n1126 585
R9158 gnd.n1127 gnd.n1118 585
R9159 gnd.n6415 gnd.n5124 585
R9160 gnd.n6515 gnd.n5124 585
R9161 gnd.n6414 gnd.n6413 585
R9162 gnd.n6413 gnd.n5131 585
R9163 gnd.n6412 gnd.n5138 585
R9164 gnd.n6412 gnd.n5130 585
R9165 gnd.n6411 gnd.n5140 585
R9166 gnd.n6411 gnd.n6410 585
R9167 gnd.n6131 gnd.n5139 585
R9168 gnd.n5152 gnd.n5139 585
R9169 gnd.n6130 gnd.n5150 585
R9170 gnd.n6397 gnd.n5150 585
R9171 gnd.n6121 gnd.n5157 585
R9172 gnd.n6122 gnd.n6121 585
R9173 gnd.n6120 gnd.n6119 585
R9174 gnd.n6120 gnd.n5161 585
R9175 gnd.n6118 gnd.n5163 585
R9176 gnd.n6111 gnd.n5163 585
R9177 gnd.n5177 gnd.n5164 585
R9178 gnd.n5177 gnd.n5168 585
R9179 gnd.n6070 gnd.n5178 585
R9180 gnd.n6101 gnd.n5178 585
R9181 gnd.n6069 gnd.n6068 585
R9182 gnd.n6068 gnd.n5185 585
R9183 gnd.n6067 gnd.n5192 585
R9184 gnd.n6067 gnd.n5184 585
R9185 gnd.n6066 gnd.n5194 585
R9186 gnd.n6066 gnd.n6065 585
R9187 gnd.n6045 gnd.n5193 585
R9188 gnd.n5205 gnd.n5193 585
R9189 gnd.n6044 gnd.n5203 585
R9190 gnd.n6055 gnd.n5203 585
R9191 gnd.n5216 gnd.n5210 585
R9192 gnd.n6036 gnd.n5216 585
R9193 gnd.n6003 gnd.n6002 585
R9194 gnd.n6002 gnd.n5214 585
R9195 gnd.n6004 gnd.n5222 585
R9196 gnd.n6021 gnd.n5222 585
R9197 gnd.n6001 gnd.n6000 585
R9198 gnd.n6000 gnd.n5232 585
R9199 gnd.n5999 gnd.n5230 585
R9200 gnd.n6011 gnd.n5230 585
R9201 gnd.n5990 gnd.n5239 585
R9202 gnd.n5991 gnd.n5990 585
R9203 gnd.n5989 gnd.n5988 585
R9204 gnd.n5989 gnd.n5243 585
R9205 gnd.n5987 gnd.n5245 585
R9206 gnd.n5980 gnd.n5245 585
R9207 gnd.n5260 gnd.n5246 585
R9208 gnd.n5260 gnd.n5250 585
R9209 gnd.n5943 gnd.n5261 585
R9210 gnd.n5970 gnd.n5261 585
R9211 gnd.n5942 gnd.n5941 585
R9212 gnd.n5941 gnd.n5348 585
R9213 gnd.n5940 gnd.n5355 585
R9214 gnd.n5940 gnd.n5347 585
R9215 gnd.n5939 gnd.n5357 585
R9216 gnd.n5939 gnd.n5938 585
R9217 gnd.n5918 gnd.n5356 585
R9218 gnd.n5369 gnd.n5356 585
R9219 gnd.n5917 gnd.n5367 585
R9220 gnd.n5928 gnd.n5367 585
R9221 gnd.n5908 gnd.n5374 585
R9222 gnd.n5909 gnd.n5908 585
R9223 gnd.n5907 gnd.n5906 585
R9224 gnd.n5907 gnd.n5378 585
R9225 gnd.n5905 gnd.n5380 585
R9226 gnd.n5898 gnd.n5380 585
R9227 gnd.n5885 gnd.n5381 585
R9228 gnd.n5886 gnd.n5885 585
R9229 gnd.n5855 gnd.n5394 585
R9230 gnd.n5888 gnd.n5394 585
R9231 gnd.n5854 gnd.n5853 585
R9232 gnd.n5853 gnd.n5852 585
R9233 gnd.n5850 gnd.n5411 585
R9234 gnd.n5850 gnd.n5402 585
R9235 gnd.n5849 gnd.n5848 585
R9236 gnd.n5849 gnd.n5401 585
R9237 gnd.n5413 gnd.n5412 585
R9238 gnd.n5840 gnd.n5412 585
R9239 gnd.n5809 gnd.n5808 585
R9240 gnd.n5808 gnd.n5417 585
R9241 gnd.n5810 gnd.n5427 585
R9242 gnd.n5827 gnd.n5427 585
R9243 gnd.n5807 gnd.n5806 585
R9244 gnd.n5806 gnd.n5434 585
R9245 gnd.n5805 gnd.n5441 585
R9246 gnd.n5805 gnd.n5433 585
R9247 gnd.n5804 gnd.n5443 585
R9248 gnd.n5804 gnd.n5803 585
R9249 gnd.n5783 gnd.n5442 585
R9250 gnd.n5455 gnd.n5442 585
R9251 gnd.n5782 gnd.n5453 585
R9252 gnd.n5793 gnd.n5453 585
R9253 gnd.n5773 gnd.n5460 585
R9254 gnd.n5774 gnd.n5773 585
R9255 gnd.n5772 gnd.n5466 585
R9256 gnd.n5772 gnd.n5771 585
R9257 gnd.n5757 gnd.n5465 585
R9258 gnd.n5476 gnd.n5465 585
R9259 gnd.n5756 gnd.n5474 585
R9260 gnd.n5763 gnd.n5474 585
R9261 gnd.n5755 gnd.n5754 585
R9262 gnd.n5754 gnd.n5753 585
R9263 gnd.n4154 gnd.n2140 585
R9264 gnd.n2140 gnd.n2126 585
R9265 gnd.n4156 gnd.n4155 585
R9266 gnd.n4157 gnd.n4156 585
R9267 gnd.n2141 gnd.n2139 585
R9268 gnd.n2139 gnd.n2134 585
R9269 gnd.n4025 gnd.n4024 585
R9270 gnd.n4026 gnd.n4025 585
R9271 gnd.n4023 gnd.n2213 585
R9272 gnd.n3944 gnd.n2213 585
R9273 gnd.n4022 gnd.n4021 585
R9274 gnd.n4021 gnd.n4020 585
R9275 gnd.n2215 gnd.n2214 585
R9276 gnd.n3997 gnd.n2215 585
R9277 gnd.n4009 gnd.n4008 585
R9278 gnd.n4010 gnd.n4009 585
R9279 gnd.n4007 gnd.n2228 585
R9280 gnd.n2228 gnd.n2223 585
R9281 gnd.n4006 gnd.n4005 585
R9282 gnd.n4005 gnd.n4004 585
R9283 gnd.n2230 gnd.n2229 585
R9284 gnd.n2236 gnd.n2230 585
R9285 gnd.n3990 gnd.n3989 585
R9286 gnd.n3991 gnd.n3990 585
R9287 gnd.n3988 gnd.n2238 585
R9288 gnd.n2244 gnd.n2238 585
R9289 gnd.n3987 gnd.n3986 585
R9290 gnd.n3986 gnd.n3985 585
R9291 gnd.n2240 gnd.n2239 585
R9292 gnd.n3858 gnd.n2240 585
R9293 gnd.n3972 gnd.n3971 585
R9294 gnd.n3973 gnd.n3972 585
R9295 gnd.n3970 gnd.n2255 585
R9296 gnd.n2255 gnd.n2252 585
R9297 gnd.n3969 gnd.n3968 585
R9298 gnd.n3968 gnd.n3967 585
R9299 gnd.n2257 gnd.n2256 585
R9300 gnd.n3855 gnd.n2257 585
R9301 gnd.n3915 gnd.n3914 585
R9302 gnd.n3915 gnd.n2266 585
R9303 gnd.n3917 gnd.n3916 585
R9304 gnd.n3916 gnd.n2265 585
R9305 gnd.n3918 gnd.n2278 585
R9306 gnd.n3869 gnd.n2278 585
R9307 gnd.n3920 gnd.n3919 585
R9308 gnd.n3921 gnd.n3920 585
R9309 gnd.n3913 gnd.n2277 585
R9310 gnd.n2277 gnd.n2273 585
R9311 gnd.n3912 gnd.n3911 585
R9312 gnd.n3911 gnd.n3910 585
R9313 gnd.n2280 gnd.n2279 585
R9314 gnd.n2281 gnd.n2280 585
R9315 gnd.n3881 gnd.n2303 585
R9316 gnd.n3881 gnd.n3880 585
R9317 gnd.n3883 gnd.n3882 585
R9318 gnd.n3882 gnd.n2289 585
R9319 gnd.n3884 gnd.n2301 585
R9320 gnd.n3848 gnd.n2301 585
R9321 gnd.n3886 gnd.n3885 585
R9322 gnd.n3887 gnd.n3886 585
R9323 gnd.n2302 gnd.n2300 585
R9324 gnd.n2300 gnd.n2296 585
R9325 gnd.n3842 gnd.n3841 585
R9326 gnd.n3843 gnd.n3842 585
R9327 gnd.n3840 gnd.n2309 585
R9328 gnd.n2315 gnd.n2309 585
R9329 gnd.n3839 gnd.n3838 585
R9330 gnd.n3838 gnd.n3837 585
R9331 gnd.n2311 gnd.n2310 585
R9332 gnd.n2312 gnd.n2311 585
R9333 gnd.n3825 gnd.n3824 585
R9334 gnd.n3826 gnd.n3825 585
R9335 gnd.n3823 gnd.n2325 585
R9336 gnd.n2325 gnd.n2321 585
R9337 gnd.n3822 gnd.n3821 585
R9338 gnd.n3821 gnd.n3820 585
R9339 gnd.n2327 gnd.n2326 585
R9340 gnd.n2334 gnd.n2327 585
R9341 gnd.n3807 gnd.n3806 585
R9342 gnd.n3808 gnd.n3807 585
R9343 gnd.n3805 gnd.n2336 585
R9344 gnd.n2336 gnd.n2333 585
R9345 gnd.n3804 gnd.n3803 585
R9346 gnd.n3803 gnd.n3802 585
R9347 gnd.n2338 gnd.n2337 585
R9348 gnd.n2350 gnd.n2338 585
R9349 gnd.n3789 gnd.n3788 585
R9350 gnd.n3790 gnd.n3789 585
R9351 gnd.n3787 gnd.n2351 585
R9352 gnd.n2351 gnd.n2347 585
R9353 gnd.n3786 gnd.n3785 585
R9354 gnd.n3785 gnd.n3784 585
R9355 gnd.n2353 gnd.n2352 585
R9356 gnd.n2354 gnd.n2353 585
R9357 gnd.n3732 gnd.n3731 585
R9358 gnd.n3732 gnd.n2363 585
R9359 gnd.n3734 gnd.n3733 585
R9360 gnd.n3733 gnd.n2362 585
R9361 gnd.n3735 gnd.n2377 585
R9362 gnd.n2377 gnd.n2375 585
R9363 gnd.n3737 gnd.n3736 585
R9364 gnd.n3738 gnd.n3737 585
R9365 gnd.n3730 gnd.n2376 585
R9366 gnd.n3725 gnd.n2376 585
R9367 gnd.n3729 gnd.n3728 585
R9368 gnd.n3728 gnd.n3727 585
R9369 gnd.n2379 gnd.n2378 585
R9370 gnd.n2380 gnd.n2379 585
R9371 gnd.n3701 gnd.n3700 585
R9372 gnd.n3702 gnd.n3701 585
R9373 gnd.n3699 gnd.n2386 585
R9374 gnd.n3695 gnd.n2386 585
R9375 gnd.n3698 gnd.n3697 585
R9376 gnd.n3697 gnd.n3696 585
R9377 gnd.n2388 gnd.n2387 585
R9378 gnd.n2394 gnd.n2388 585
R9379 gnd.n3687 gnd.n3686 585
R9380 gnd.n3688 gnd.n3687 585
R9381 gnd.n3685 gnd.n2396 585
R9382 gnd.n2396 gnd.n2393 585
R9383 gnd.n3684 gnd.n3683 585
R9384 gnd.n3683 gnd.n3682 585
R9385 gnd.n2398 gnd.n2397 585
R9386 gnd.n3630 gnd.n2398 585
R9387 gnd.n2434 gnd.n2433 585
R9388 gnd.n2434 gnd.n2422 585
R9389 gnd.n3638 gnd.n3637 585
R9390 gnd.n3637 gnd.n3636 585
R9391 gnd.n3639 gnd.n2431 585
R9392 gnd.n2436 gnd.n2431 585
R9393 gnd.n3641 gnd.n3640 585
R9394 gnd.n3642 gnd.n3641 585
R9395 gnd.n2432 gnd.n2430 585
R9396 gnd.n3624 gnd.n2430 585
R9397 gnd.n2464 gnd.n2463 585
R9398 gnd.n2463 gnd.n2441 585
R9399 gnd.n3596 gnd.n2465 585
R9400 gnd.n3596 gnd.n3595 585
R9401 gnd.n3597 gnd.n2462 585
R9402 gnd.n3597 gnd.n2449 585
R9403 gnd.n3599 gnd.n3598 585
R9404 gnd.n3598 gnd.n2448 585
R9405 gnd.n3600 gnd.n2460 585
R9406 gnd.n3588 gnd.n2460 585
R9407 gnd.n3602 gnd.n3601 585
R9408 gnd.n3603 gnd.n3602 585
R9409 gnd.n2461 gnd.n2459 585
R9410 gnd.n2459 gnd.n2456 585
R9411 gnd.n3579 gnd.n3578 585
R9412 gnd.n3580 gnd.n3579 585
R9413 gnd.n3577 gnd.n2471 585
R9414 gnd.n2478 gnd.n2471 585
R9415 gnd.n3576 gnd.n3575 585
R9416 gnd.n3575 gnd.n3574 585
R9417 gnd.n2473 gnd.n2472 585
R9418 gnd.n3497 gnd.n2473 585
R9419 gnd.n3563 gnd.n3562 585
R9420 gnd.n3564 gnd.n3563 585
R9421 gnd.n3561 gnd.n2487 585
R9422 gnd.n2487 gnd.n2484 585
R9423 gnd.n3560 gnd.n3559 585
R9424 gnd.n3559 gnd.n3558 585
R9425 gnd.n2489 gnd.n2488 585
R9426 gnd.n3493 gnd.n2489 585
R9427 gnd.n3521 gnd.n3520 585
R9428 gnd.n3521 gnd.n2498 585
R9429 gnd.n3523 gnd.n3522 585
R9430 gnd.n3522 gnd.n2497 585
R9431 gnd.n3524 gnd.n2511 585
R9432 gnd.n3509 gnd.n2511 585
R9433 gnd.n3526 gnd.n3525 585
R9434 gnd.n3527 gnd.n3526 585
R9435 gnd.n3519 gnd.n2510 585
R9436 gnd.n2510 gnd.n2507 585
R9437 gnd.n3518 gnd.n3517 585
R9438 gnd.n3517 gnd.n3516 585
R9439 gnd.n2513 gnd.n2512 585
R9440 gnd.n2519 gnd.n2513 585
R9441 gnd.n3486 gnd.n3485 585
R9442 gnd.n3487 gnd.n3486 585
R9443 gnd.n3484 gnd.n2521 585
R9444 gnd.n2521 gnd.n1698 585
R9445 gnd.n3483 gnd.n3482 585
R9446 gnd.n3482 gnd.n3481 585
R9447 gnd.n2523 gnd.n2522 585
R9448 gnd.n3405 gnd.n2523 585
R9449 gnd.n1683 gnd.n1682 585
R9450 gnd.n1687 gnd.n1683 585
R9451 gnd.n4688 gnd.n4687 585
R9452 gnd.n4687 gnd.n4686 585
R9453 gnd.n4689 gnd.n1661 585
R9454 gnd.n3472 gnd.n1661 585
R9455 gnd.n4754 gnd.n4753 585
R9456 gnd.n4752 gnd.n1660 585
R9457 gnd.n4751 gnd.n1659 585
R9458 gnd.n4756 gnd.n1659 585
R9459 gnd.n4750 gnd.n4749 585
R9460 gnd.n4748 gnd.n4747 585
R9461 gnd.n4746 gnd.n4745 585
R9462 gnd.n4744 gnd.n4743 585
R9463 gnd.n4742 gnd.n4741 585
R9464 gnd.n4740 gnd.n4739 585
R9465 gnd.n4738 gnd.n4737 585
R9466 gnd.n4736 gnd.n4735 585
R9467 gnd.n4734 gnd.n4733 585
R9468 gnd.n4732 gnd.n4731 585
R9469 gnd.n4730 gnd.n4729 585
R9470 gnd.n4728 gnd.n4727 585
R9471 gnd.n4726 gnd.n4725 585
R9472 gnd.n4724 gnd.n4723 585
R9473 gnd.n4722 gnd.n4721 585
R9474 gnd.n4720 gnd.n4719 585
R9475 gnd.n4718 gnd.n4717 585
R9476 gnd.n4716 gnd.n4715 585
R9477 gnd.n4714 gnd.n4713 585
R9478 gnd.n4712 gnd.n4711 585
R9479 gnd.n4710 gnd.n4709 585
R9480 gnd.n4708 gnd.n4707 585
R9481 gnd.n4706 gnd.n4705 585
R9482 gnd.n4704 gnd.n4703 585
R9483 gnd.n4702 gnd.n4701 585
R9484 gnd.n4700 gnd.n4699 585
R9485 gnd.n4698 gnd.n4697 585
R9486 gnd.n4696 gnd.n4695 585
R9487 gnd.n4694 gnd.n1623 585
R9488 gnd.n4759 gnd.n4758 585
R9489 gnd.n1625 gnd.n1622 585
R9490 gnd.n3410 gnd.n3409 585
R9491 gnd.n3412 gnd.n3411 585
R9492 gnd.n3415 gnd.n3414 585
R9493 gnd.n3417 gnd.n3416 585
R9494 gnd.n3419 gnd.n3418 585
R9495 gnd.n3421 gnd.n3420 585
R9496 gnd.n3423 gnd.n3422 585
R9497 gnd.n3425 gnd.n3424 585
R9498 gnd.n3427 gnd.n3426 585
R9499 gnd.n3429 gnd.n3428 585
R9500 gnd.n3431 gnd.n3430 585
R9501 gnd.n3433 gnd.n3432 585
R9502 gnd.n3435 gnd.n3434 585
R9503 gnd.n3437 gnd.n3436 585
R9504 gnd.n3439 gnd.n3438 585
R9505 gnd.n3441 gnd.n3440 585
R9506 gnd.n3443 gnd.n3442 585
R9507 gnd.n3445 gnd.n3444 585
R9508 gnd.n3447 gnd.n3446 585
R9509 gnd.n3449 gnd.n3448 585
R9510 gnd.n3451 gnd.n3450 585
R9511 gnd.n3453 gnd.n3452 585
R9512 gnd.n3455 gnd.n3454 585
R9513 gnd.n3457 gnd.n3456 585
R9514 gnd.n3459 gnd.n3458 585
R9515 gnd.n3461 gnd.n3460 585
R9516 gnd.n3463 gnd.n3462 585
R9517 gnd.n3465 gnd.n3464 585
R9518 gnd.n3467 gnd.n3466 585
R9519 gnd.n3469 gnd.n3468 585
R9520 gnd.n3471 gnd.n3470 585
R9521 gnd.n4035 gnd.n4034 585
R9522 gnd.n4036 gnd.n2210 585
R9523 gnd.n4038 gnd.n4037 585
R9524 gnd.n4040 gnd.n2208 585
R9525 gnd.n4042 gnd.n4041 585
R9526 gnd.n4043 gnd.n2207 585
R9527 gnd.n4045 gnd.n4044 585
R9528 gnd.n4047 gnd.n2205 585
R9529 gnd.n4049 gnd.n4048 585
R9530 gnd.n4050 gnd.n2204 585
R9531 gnd.n4052 gnd.n4051 585
R9532 gnd.n4054 gnd.n2202 585
R9533 gnd.n4056 gnd.n4055 585
R9534 gnd.n4057 gnd.n2201 585
R9535 gnd.n4059 gnd.n4058 585
R9536 gnd.n4061 gnd.n2199 585
R9537 gnd.n4063 gnd.n4062 585
R9538 gnd.n4064 gnd.n2198 585
R9539 gnd.n4066 gnd.n4065 585
R9540 gnd.n4068 gnd.n2196 585
R9541 gnd.n4070 gnd.n4069 585
R9542 gnd.n4071 gnd.n2195 585
R9543 gnd.n4073 gnd.n4072 585
R9544 gnd.n4075 gnd.n2193 585
R9545 gnd.n4077 gnd.n4076 585
R9546 gnd.n4078 gnd.n2192 585
R9547 gnd.n4080 gnd.n4079 585
R9548 gnd.n4082 gnd.n2190 585
R9549 gnd.n4084 gnd.n4083 585
R9550 gnd.n4086 gnd.n2187 585
R9551 gnd.n4088 gnd.n4087 585
R9552 gnd.n4090 gnd.n2186 585
R9553 gnd.n4091 gnd.n2128 585
R9554 gnd.n4094 gnd.n1935 585
R9555 gnd.n4096 gnd.n4095 585
R9556 gnd.n4098 gnd.n2184 585
R9557 gnd.n4100 gnd.n4099 585
R9558 gnd.n4102 gnd.n2181 585
R9559 gnd.n4104 gnd.n4103 585
R9560 gnd.n4106 gnd.n2179 585
R9561 gnd.n4108 gnd.n4107 585
R9562 gnd.n4109 gnd.n2178 585
R9563 gnd.n4111 gnd.n4110 585
R9564 gnd.n4113 gnd.n2176 585
R9565 gnd.n4115 gnd.n4114 585
R9566 gnd.n4116 gnd.n2175 585
R9567 gnd.n4118 gnd.n4117 585
R9568 gnd.n4120 gnd.n2173 585
R9569 gnd.n4122 gnd.n4121 585
R9570 gnd.n4123 gnd.n2172 585
R9571 gnd.n4125 gnd.n4124 585
R9572 gnd.n4127 gnd.n2170 585
R9573 gnd.n4129 gnd.n4128 585
R9574 gnd.n4130 gnd.n2169 585
R9575 gnd.n4132 gnd.n4131 585
R9576 gnd.n4134 gnd.n2167 585
R9577 gnd.n4136 gnd.n4135 585
R9578 gnd.n4137 gnd.n2166 585
R9579 gnd.n4139 gnd.n4138 585
R9580 gnd.n4141 gnd.n2164 585
R9581 gnd.n4143 gnd.n4142 585
R9582 gnd.n4144 gnd.n2163 585
R9583 gnd.n4146 gnd.n4145 585
R9584 gnd.n4148 gnd.n2162 585
R9585 gnd.n4149 gnd.n2161 585
R9586 gnd.n4152 gnd.n4151 585
R9587 gnd.n4033 gnd.n4031 585
R9588 gnd.n4033 gnd.n2126 585
R9589 gnd.n4030 gnd.n2136 585
R9590 gnd.n4157 gnd.n2136 585
R9591 gnd.n4029 gnd.n4028 585
R9592 gnd.n4028 gnd.n2134 585
R9593 gnd.n4027 gnd.n2211 585
R9594 gnd.n4027 gnd.n4026 585
R9595 gnd.n3995 gnd.n2212 585
R9596 gnd.n3944 gnd.n2212 585
R9597 gnd.n3996 gnd.n2216 585
R9598 gnd.n4020 gnd.n2216 585
R9599 gnd.n3999 gnd.n3998 585
R9600 gnd.n3998 gnd.n3997 585
R9601 gnd.n4000 gnd.n2225 585
R9602 gnd.n4010 gnd.n2225 585
R9603 gnd.n4001 gnd.n2233 585
R9604 gnd.n2233 gnd.n2223 585
R9605 gnd.n4003 gnd.n4002 585
R9606 gnd.n4004 gnd.n4003 585
R9607 gnd.n3994 gnd.n2232 585
R9608 gnd.n2236 gnd.n2232 585
R9609 gnd.n3993 gnd.n3992 585
R9610 gnd.n3992 gnd.n3991 585
R9611 gnd.n2235 gnd.n2234 585
R9612 gnd.n2244 gnd.n2235 585
R9613 gnd.n3857 gnd.n2242 585
R9614 gnd.n3985 gnd.n2242 585
R9615 gnd.n3860 gnd.n3859 585
R9616 gnd.n3859 gnd.n3858 585
R9617 gnd.n3861 gnd.n2254 585
R9618 gnd.n3973 gnd.n2254 585
R9619 gnd.n3863 gnd.n3862 585
R9620 gnd.n3862 gnd.n2252 585
R9621 gnd.n3864 gnd.n2258 585
R9622 gnd.n3967 gnd.n2258 585
R9623 gnd.n3865 gnd.n3856 585
R9624 gnd.n3856 gnd.n3855 585
R9625 gnd.n3867 gnd.n3866 585
R9626 gnd.n3867 gnd.n2266 585
R9627 gnd.n3868 gnd.n3852 585
R9628 gnd.n3868 gnd.n2265 585
R9629 gnd.n3871 gnd.n3870 585
R9630 gnd.n3870 gnd.n3869 585
R9631 gnd.n3872 gnd.n2275 585
R9632 gnd.n3921 gnd.n2275 585
R9633 gnd.n3874 gnd.n3873 585
R9634 gnd.n3873 gnd.n2273 585
R9635 gnd.n3875 gnd.n2282 585
R9636 gnd.n3910 gnd.n2282 585
R9637 gnd.n3876 gnd.n2305 585
R9638 gnd.n2305 gnd.n2281 585
R9639 gnd.n3878 gnd.n3877 585
R9640 gnd.n3880 gnd.n3878 585
R9641 gnd.n3851 gnd.n2304 585
R9642 gnd.n2304 gnd.n2289 585
R9643 gnd.n3850 gnd.n3849 585
R9644 gnd.n3849 gnd.n3848 585
R9645 gnd.n3847 gnd.n2298 585
R9646 gnd.n3887 gnd.n2298 585
R9647 gnd.n3846 gnd.n3845 585
R9648 gnd.n3845 gnd.n2296 585
R9649 gnd.n3844 gnd.n2306 585
R9650 gnd.n3844 gnd.n3843 585
R9651 gnd.n3812 gnd.n2307 585
R9652 gnd.n2315 gnd.n2307 585
R9653 gnd.n3813 gnd.n2313 585
R9654 gnd.n3837 gnd.n2313 585
R9655 gnd.n3815 gnd.n3814 585
R9656 gnd.n3814 gnd.n2312 585
R9657 gnd.n3816 gnd.n2323 585
R9658 gnd.n3826 gnd.n2323 585
R9659 gnd.n3817 gnd.n2330 585
R9660 gnd.n2330 gnd.n2321 585
R9661 gnd.n3819 gnd.n3818 585
R9662 gnd.n3820 gnd.n3819 585
R9663 gnd.n3811 gnd.n2329 585
R9664 gnd.n2334 gnd.n2329 585
R9665 gnd.n3810 gnd.n3809 585
R9666 gnd.n3809 gnd.n3808 585
R9667 gnd.n2332 gnd.n2331 585
R9668 gnd.n2333 gnd.n2332 585
R9669 gnd.n3709 gnd.n2339 585
R9670 gnd.n3802 gnd.n2339 585
R9671 gnd.n3711 gnd.n3710 585
R9672 gnd.n3710 gnd.n2350 585
R9673 gnd.n3712 gnd.n2349 585
R9674 gnd.n3790 gnd.n2349 585
R9675 gnd.n3714 gnd.n3713 585
R9676 gnd.n3713 gnd.n2347 585
R9677 gnd.n3715 gnd.n2355 585
R9678 gnd.n3784 gnd.n2355 585
R9679 gnd.n3716 gnd.n3708 585
R9680 gnd.n3708 gnd.n2354 585
R9681 gnd.n3718 gnd.n3717 585
R9682 gnd.n3718 gnd.n2363 585
R9683 gnd.n3719 gnd.n3707 585
R9684 gnd.n3719 gnd.n2362 585
R9685 gnd.n3721 gnd.n3720 585
R9686 gnd.n3720 gnd.n2375 585
R9687 gnd.n3722 gnd.n2373 585
R9688 gnd.n3738 gnd.n2373 585
R9689 gnd.n3724 gnd.n3723 585
R9690 gnd.n3725 gnd.n3724 585
R9691 gnd.n3706 gnd.n2381 585
R9692 gnd.n3727 gnd.n2381 585
R9693 gnd.n3705 gnd.n3704 585
R9694 gnd.n3704 gnd.n2380 585
R9695 gnd.n3703 gnd.n2383 585
R9696 gnd.n3703 gnd.n3702 585
R9697 gnd.n3692 gnd.n2384 585
R9698 gnd.n3695 gnd.n2384 585
R9699 gnd.n3694 gnd.n3693 585
R9700 gnd.n3696 gnd.n3694 585
R9701 gnd.n3691 gnd.n2390 585
R9702 gnd.n2394 gnd.n2390 585
R9703 gnd.n3690 gnd.n3689 585
R9704 gnd.n3689 gnd.n3688 585
R9705 gnd.n2392 gnd.n2391 585
R9706 gnd.n2393 gnd.n2392 585
R9707 gnd.n3629 gnd.n2400 585
R9708 gnd.n3682 gnd.n2400 585
R9709 gnd.n3632 gnd.n3631 585
R9710 gnd.n3631 gnd.n3630 585
R9711 gnd.n3633 gnd.n2438 585
R9712 gnd.n2438 gnd.n2422 585
R9713 gnd.n3635 gnd.n3634 585
R9714 gnd.n3636 gnd.n3635 585
R9715 gnd.n3628 gnd.n2437 585
R9716 gnd.n2437 gnd.n2436 585
R9717 gnd.n3627 gnd.n2429 585
R9718 gnd.n3642 gnd.n2429 585
R9719 gnd.n3626 gnd.n3625 585
R9720 gnd.n3625 gnd.n3624 585
R9721 gnd.n2440 gnd.n2439 585
R9722 gnd.n2441 gnd.n2440 585
R9723 gnd.n3594 gnd.n3593 585
R9724 gnd.n3595 gnd.n3594 585
R9725 gnd.n3592 gnd.n2467 585
R9726 gnd.n2467 gnd.n2449 585
R9727 gnd.n3591 gnd.n3590 585
R9728 gnd.n3590 gnd.n2448 585
R9729 gnd.n3589 gnd.n3585 585
R9730 gnd.n3589 gnd.n3588 585
R9731 gnd.n3584 gnd.n2458 585
R9732 gnd.n3603 gnd.n2458 585
R9733 gnd.n3583 gnd.n3582 585
R9734 gnd.n3582 gnd.n2456 585
R9735 gnd.n3581 gnd.n2468 585
R9736 gnd.n3581 gnd.n3580 585
R9737 gnd.n3495 gnd.n2469 585
R9738 gnd.n2478 gnd.n2469 585
R9739 gnd.n3496 gnd.n2476 585
R9740 gnd.n3574 gnd.n2476 585
R9741 gnd.n3499 gnd.n3498 585
R9742 gnd.n3498 gnd.n3497 585
R9743 gnd.n3500 gnd.n2486 585
R9744 gnd.n3564 gnd.n2486 585
R9745 gnd.n3502 gnd.n3501 585
R9746 gnd.n3501 gnd.n2484 585
R9747 gnd.n3503 gnd.n2490 585
R9748 gnd.n3558 gnd.n2490 585
R9749 gnd.n3504 gnd.n3494 585
R9750 gnd.n3494 gnd.n3493 585
R9751 gnd.n3506 gnd.n3505 585
R9752 gnd.n3506 gnd.n2498 585
R9753 gnd.n3507 gnd.n3491 585
R9754 gnd.n3507 gnd.n2497 585
R9755 gnd.n3511 gnd.n3510 585
R9756 gnd.n3510 gnd.n3509 585
R9757 gnd.n3512 gnd.n2509 585
R9758 gnd.n3527 gnd.n2509 585
R9759 gnd.n3513 gnd.n2516 585
R9760 gnd.n2516 gnd.n2507 585
R9761 gnd.n3515 gnd.n3514 585
R9762 gnd.n3516 gnd.n3515 585
R9763 gnd.n3490 gnd.n2515 585
R9764 gnd.n2519 gnd.n2515 585
R9765 gnd.n3489 gnd.n3488 585
R9766 gnd.n3488 gnd.n3487 585
R9767 gnd.n2518 gnd.n2517 585
R9768 gnd.n2518 gnd.n1698 585
R9769 gnd.n3480 gnd.n3479 585
R9770 gnd.n3481 gnd.n3480 585
R9771 gnd.n3478 gnd.n3406 585
R9772 gnd.n3406 gnd.n3405 585
R9773 gnd.n3477 gnd.n3476 585
R9774 gnd.n3476 gnd.n1687 585
R9775 gnd.n3475 gnd.n1685 585
R9776 gnd.n4686 gnd.n1685 585
R9777 gnd.n3474 gnd.n3473 585
R9778 gnd.n3473 gnd.n3472 585
R9779 gnd.n4815 gnd.n1546 585
R9780 gnd.n3318 gnd.n1546 585
R9781 gnd.n4817 gnd.n4816 585
R9782 gnd.n4818 gnd.n4817 585
R9783 gnd.n1531 gnd.n1530 585
R9784 gnd.n3278 gnd.n1531 585
R9785 gnd.n4826 gnd.n4825 585
R9786 gnd.n4825 gnd.n4824 585
R9787 gnd.n4827 gnd.n1525 585
R9788 gnd.n3026 gnd.n1525 585
R9789 gnd.n4829 gnd.n4828 585
R9790 gnd.n4830 gnd.n4829 585
R9791 gnd.n1511 gnd.n1510 585
R9792 gnd.n3291 gnd.n1511 585
R9793 gnd.n4838 gnd.n4837 585
R9794 gnd.n4837 gnd.n4836 585
R9795 gnd.n4839 gnd.n1505 585
R9796 gnd.n3019 gnd.n1505 585
R9797 gnd.n4841 gnd.n4840 585
R9798 gnd.n4842 gnd.n4841 585
R9799 gnd.n1491 gnd.n1490 585
R9800 gnd.n3011 gnd.n1491 585
R9801 gnd.n4850 gnd.n4849 585
R9802 gnd.n4849 gnd.n4848 585
R9803 gnd.n4851 gnd.n1485 585
R9804 gnd.n2973 gnd.n1485 585
R9805 gnd.n4853 gnd.n4852 585
R9806 gnd.n4854 gnd.n4853 585
R9807 gnd.n1471 gnd.n1470 585
R9808 gnd.n2964 gnd.n1471 585
R9809 gnd.n4862 gnd.n4861 585
R9810 gnd.n4861 gnd.n4860 585
R9811 gnd.n4863 gnd.n1465 585
R9812 gnd.n2959 gnd.n1465 585
R9813 gnd.n4865 gnd.n4864 585
R9814 gnd.n4866 gnd.n4865 585
R9815 gnd.n1451 gnd.n1450 585
R9816 gnd.n2987 gnd.n1451 585
R9817 gnd.n4874 gnd.n4873 585
R9818 gnd.n4873 gnd.n4872 585
R9819 gnd.n4875 gnd.n1445 585
R9820 gnd.n2952 gnd.n1445 585
R9821 gnd.n4877 gnd.n4876 585
R9822 gnd.n4878 gnd.n4877 585
R9823 gnd.n1431 gnd.n1430 585
R9824 gnd.n2944 gnd.n1431 585
R9825 gnd.n4886 gnd.n4885 585
R9826 gnd.n4885 gnd.n4884 585
R9827 gnd.n4887 gnd.n1426 585
R9828 gnd.n2938 gnd.n1426 585
R9829 gnd.n4889 gnd.n4888 585
R9830 gnd.n4890 gnd.n4889 585
R9831 gnd.n1410 gnd.n1408 585
R9832 gnd.n2930 gnd.n1410 585
R9833 gnd.n4898 gnd.n4897 585
R9834 gnd.n4897 gnd.n4896 585
R9835 gnd.n1409 gnd.n1407 585
R9836 gnd.n2899 gnd.n1409 585
R9837 gnd.n2888 gnd.n2887 585
R9838 gnd.n2887 gnd.n2641 585
R9839 gnd.n2890 gnd.n2889 585
R9840 gnd.n2891 gnd.n2890 585
R9841 gnd.n2886 gnd.n2653 585
R9842 gnd.n2886 gnd.n2885 585
R9843 gnd.n2652 gnd.n2651 585
R9844 gnd.n2869 gnd.n2651 585
R9845 gnd.n2725 gnd.n2724 585
R9846 gnd.n2726 gnd.n2725 585
R9847 gnd.n1401 gnd.n1399 585
R9848 gnd.n1399 gnd.n1398 585
R9849 gnd.n4902 gnd.n4901 585
R9850 gnd.n4903 gnd.n4902 585
R9851 gnd.n1400 gnd.n1385 585
R9852 gnd.n1389 gnd.n1385 585
R9853 gnd.n4911 gnd.n4910 585
R9854 gnd.n4910 gnd.n4909 585
R9855 gnd.n4912 gnd.n1380 585
R9856 gnd.n1386 gnd.n1380 585
R9857 gnd.n4914 gnd.n4913 585
R9858 gnd.n4915 gnd.n4914 585
R9859 gnd.n1368 gnd.n1367 585
R9860 gnd.n1371 gnd.n1368 585
R9861 gnd.n4923 gnd.n4922 585
R9862 gnd.n4922 gnd.n4921 585
R9863 gnd.n4924 gnd.n1362 585
R9864 gnd.n1362 gnd.n1361 585
R9865 gnd.n4926 gnd.n4925 585
R9866 gnd.n4927 gnd.n4926 585
R9867 gnd.n1348 gnd.n1347 585
R9868 gnd.n1352 gnd.n1348 585
R9869 gnd.n4935 gnd.n4934 585
R9870 gnd.n4934 gnd.n4933 585
R9871 gnd.n4936 gnd.n1342 585
R9872 gnd.n1349 gnd.n1342 585
R9873 gnd.n4938 gnd.n4937 585
R9874 gnd.n4939 gnd.n4938 585
R9875 gnd.n1330 gnd.n1329 585
R9876 gnd.n1333 gnd.n1330 585
R9877 gnd.n4947 gnd.n4946 585
R9878 gnd.n4946 gnd.n4945 585
R9879 gnd.n4948 gnd.n1324 585
R9880 gnd.n1324 gnd.n1323 585
R9881 gnd.n4950 gnd.n4949 585
R9882 gnd.n4951 gnd.n4950 585
R9883 gnd.n1310 gnd.n1309 585
R9884 gnd.n1314 gnd.n1310 585
R9885 gnd.n4959 gnd.n4958 585
R9886 gnd.n4958 gnd.n4957 585
R9887 gnd.n4960 gnd.n1304 585
R9888 gnd.n1311 gnd.n1304 585
R9889 gnd.n4962 gnd.n4961 585
R9890 gnd.n4963 gnd.n4962 585
R9891 gnd.n1292 gnd.n1291 585
R9892 gnd.n1295 gnd.n1292 585
R9893 gnd.n4971 gnd.n4970 585
R9894 gnd.n4970 gnd.n4969 585
R9895 gnd.n4972 gnd.n1286 585
R9896 gnd.n1286 gnd.n1285 585
R9897 gnd.n4974 gnd.n4973 585
R9898 gnd.n4975 gnd.n4974 585
R9899 gnd.n1269 gnd.n1268 585
R9900 gnd.n1273 gnd.n1269 585
R9901 gnd.n4983 gnd.n4982 585
R9902 gnd.n4982 gnd.n4981 585
R9903 gnd.n4984 gnd.n1262 585
R9904 gnd.n1270 gnd.n1262 585
R9905 gnd.n4986 gnd.n4985 585
R9906 gnd.n4987 gnd.n4986 585
R9907 gnd.n1263 gnd.n1189 585
R9908 gnd.n1189 gnd.n1186 585
R9909 gnd.n5109 gnd.n5108 585
R9910 gnd.n5107 gnd.n1188 585
R9911 gnd.n5106 gnd.n1187 585
R9912 gnd.n5111 gnd.n1187 585
R9913 gnd.n5105 gnd.n5104 585
R9914 gnd.n5103 gnd.n5102 585
R9915 gnd.n5101 gnd.n5100 585
R9916 gnd.n5099 gnd.n5098 585
R9917 gnd.n5097 gnd.n5096 585
R9918 gnd.n5095 gnd.n5094 585
R9919 gnd.n5093 gnd.n5092 585
R9920 gnd.n5091 gnd.n5090 585
R9921 gnd.n5089 gnd.n5088 585
R9922 gnd.n5087 gnd.n5086 585
R9923 gnd.n5085 gnd.n5084 585
R9924 gnd.n5083 gnd.n5082 585
R9925 gnd.n5081 gnd.n5080 585
R9926 gnd.n5079 gnd.n5078 585
R9927 gnd.n5077 gnd.n5076 585
R9928 gnd.n5074 gnd.n5073 585
R9929 gnd.n5072 gnd.n5071 585
R9930 gnd.n5070 gnd.n5069 585
R9931 gnd.n5068 gnd.n5067 585
R9932 gnd.n5066 gnd.n5065 585
R9933 gnd.n5064 gnd.n5063 585
R9934 gnd.n5062 gnd.n5061 585
R9935 gnd.n5060 gnd.n5059 585
R9936 gnd.n5058 gnd.n5057 585
R9937 gnd.n5056 gnd.n5055 585
R9938 gnd.n5054 gnd.n5053 585
R9939 gnd.n5052 gnd.n5051 585
R9940 gnd.n5050 gnd.n5049 585
R9941 gnd.n5048 gnd.n5047 585
R9942 gnd.n5046 gnd.n5045 585
R9943 gnd.n5044 gnd.n5043 585
R9944 gnd.n5042 gnd.n5041 585
R9945 gnd.n5040 gnd.n5039 585
R9946 gnd.n5038 gnd.n5037 585
R9947 gnd.n5036 gnd.n5035 585
R9948 gnd.n5034 gnd.n5033 585
R9949 gnd.n5032 gnd.n5031 585
R9950 gnd.n5030 gnd.n5029 585
R9951 gnd.n5028 gnd.n5027 585
R9952 gnd.n5026 gnd.n5025 585
R9953 gnd.n5024 gnd.n5023 585
R9954 gnd.n5022 gnd.n5021 585
R9955 gnd.n5020 gnd.n5019 585
R9956 gnd.n5018 gnd.n5017 585
R9957 gnd.n5016 gnd.n5015 585
R9958 gnd.n5014 gnd.n5013 585
R9959 gnd.n5012 gnd.n5011 585
R9960 gnd.n5010 gnd.n5009 585
R9961 gnd.n5008 gnd.n5007 585
R9962 gnd.n5006 gnd.n5005 585
R9963 gnd.n5004 gnd.n5003 585
R9964 gnd.n5002 gnd.n5001 585
R9965 gnd.n5000 gnd.n4999 585
R9966 gnd.n4998 gnd.n4997 585
R9967 gnd.n4996 gnd.n4995 585
R9968 gnd.n1258 gnd.n1251 585
R9969 gnd.n3270 gnd.n3269 585
R9970 gnd.n3268 gnd.n3179 585
R9971 gnd.n3267 gnd.n3266 585
R9972 gnd.n3260 gnd.n3180 585
R9973 gnd.n3262 gnd.n3261 585
R9974 gnd.n3259 gnd.n3258 585
R9975 gnd.n3257 gnd.n3256 585
R9976 gnd.n3250 gnd.n3182 585
R9977 gnd.n3252 gnd.n3251 585
R9978 gnd.n3249 gnd.n3248 585
R9979 gnd.n3247 gnd.n3246 585
R9980 gnd.n3240 gnd.n3184 585
R9981 gnd.n3242 gnd.n3241 585
R9982 gnd.n3239 gnd.n3238 585
R9983 gnd.n3237 gnd.n3236 585
R9984 gnd.n3230 gnd.n3186 585
R9985 gnd.n3232 gnd.n3231 585
R9986 gnd.n3229 gnd.n3228 585
R9987 gnd.n3227 gnd.n3226 585
R9988 gnd.n3220 gnd.n3188 585
R9989 gnd.n3222 gnd.n3221 585
R9990 gnd.n3219 gnd.n3192 585
R9991 gnd.n3218 gnd.n3217 585
R9992 gnd.n3211 gnd.n3193 585
R9993 gnd.n3213 gnd.n3212 585
R9994 gnd.n3210 gnd.n3209 585
R9995 gnd.n3208 gnd.n3207 585
R9996 gnd.n3201 gnd.n3195 585
R9997 gnd.n3203 gnd.n3202 585
R9998 gnd.n3200 gnd.n3199 585
R9999 gnd.n3198 gnd.n1619 585
R10000 gnd.n4762 gnd.n4761 585
R10001 gnd.n4764 gnd.n4763 585
R10002 gnd.n4766 gnd.n4765 585
R10003 gnd.n4768 gnd.n4767 585
R10004 gnd.n4770 gnd.n4769 585
R10005 gnd.n4772 gnd.n4771 585
R10006 gnd.n4774 gnd.n4773 585
R10007 gnd.n4776 gnd.n4775 585
R10008 gnd.n4779 gnd.n4778 585
R10009 gnd.n4781 gnd.n4780 585
R10010 gnd.n4783 gnd.n4782 585
R10011 gnd.n4785 gnd.n4784 585
R10012 gnd.n4787 gnd.n4786 585
R10013 gnd.n4789 gnd.n4788 585
R10014 gnd.n4791 gnd.n4790 585
R10015 gnd.n4793 gnd.n4792 585
R10016 gnd.n4795 gnd.n4794 585
R10017 gnd.n4797 gnd.n4796 585
R10018 gnd.n4799 gnd.n4798 585
R10019 gnd.n4801 gnd.n4800 585
R10020 gnd.n4803 gnd.n4802 585
R10021 gnd.n4805 gnd.n4804 585
R10022 gnd.n4806 gnd.n1592 585
R10023 gnd.n4808 gnd.n4807 585
R10024 gnd.n1551 gnd.n1550 585
R10025 gnd.n4812 gnd.n4811 585
R10026 gnd.n4811 gnd.n4810 585
R10027 gnd.n3274 gnd.n2581 585
R10028 gnd.n3318 gnd.n2581 585
R10029 gnd.n3275 gnd.n1543 585
R10030 gnd.n4818 gnd.n1543 585
R10031 gnd.n3277 gnd.n3276 585
R10032 gnd.n3278 gnd.n3277 585
R10033 gnd.n3029 gnd.n1533 585
R10034 gnd.n4824 gnd.n1533 585
R10035 gnd.n3028 gnd.n3027 585
R10036 gnd.n3027 gnd.n3026 585
R10037 gnd.n3024 gnd.n1522 585
R10038 gnd.n4830 gnd.n1522 585
R10039 gnd.n3023 gnd.n2592 585
R10040 gnd.n3291 gnd.n2592 585
R10041 gnd.n3022 gnd.n1513 585
R10042 gnd.n4836 gnd.n1513 585
R10043 gnd.n3021 gnd.n3020 585
R10044 gnd.n3020 gnd.n3019 585
R10045 gnd.n2598 gnd.n1502 585
R10046 gnd.n4842 gnd.n1502 585
R10047 gnd.n2969 gnd.n2603 585
R10048 gnd.n3011 gnd.n2603 585
R10049 gnd.n2970 gnd.n1493 585
R10050 gnd.n4848 gnd.n1493 585
R10051 gnd.n2972 gnd.n2971 585
R10052 gnd.n2973 gnd.n2972 585
R10053 gnd.n2967 gnd.n1482 585
R10054 gnd.n4854 gnd.n1482 585
R10055 gnd.n2966 gnd.n2965 585
R10056 gnd.n2965 gnd.n2964 585
R10057 gnd.n2962 gnd.n1473 585
R10058 gnd.n4860 gnd.n1473 585
R10059 gnd.n2961 gnd.n2960 585
R10060 gnd.n2960 gnd.n2959 585
R10061 gnd.n2957 gnd.n1462 585
R10062 gnd.n4866 gnd.n1462 585
R10063 gnd.n2956 gnd.n2615 585
R10064 gnd.n2987 gnd.n2615 585
R10065 gnd.n2955 gnd.n1453 585
R10066 gnd.n4872 gnd.n1453 585
R10067 gnd.n2954 gnd.n2953 585
R10068 gnd.n2953 gnd.n2952 585
R10069 gnd.n2623 gnd.n1442 585
R10070 gnd.n4878 gnd.n1442 585
R10071 gnd.n2943 gnd.n2942 585
R10072 gnd.n2944 gnd.n2943 585
R10073 gnd.n2941 gnd.n1433 585
R10074 gnd.n4884 gnd.n1433 585
R10075 gnd.n2940 gnd.n2939 585
R10076 gnd.n2939 gnd.n2938 585
R10077 gnd.n2629 gnd.n1423 585
R10078 gnd.n4890 gnd.n1423 585
R10079 gnd.n2874 gnd.n2634 585
R10080 gnd.n2930 gnd.n2634 585
R10081 gnd.n2875 gnd.n1412 585
R10082 gnd.n4896 gnd.n1412 585
R10083 gnd.n2876 gnd.n2642 585
R10084 gnd.n2899 gnd.n2642 585
R10085 gnd.n2878 gnd.n2877 585
R10086 gnd.n2877 gnd.n2641 585
R10087 gnd.n2873 gnd.n2648 585
R10088 gnd.n2891 gnd.n2648 585
R10089 gnd.n2872 gnd.n2661 585
R10090 gnd.n2885 gnd.n2661 585
R10091 gnd.n2871 gnd.n2870 585
R10092 gnd.n2870 gnd.n2869 585
R10093 gnd.n2669 gnd.n2667 585
R10094 gnd.n2726 gnd.n2669 585
R10095 gnd.n2719 gnd.n2718 585
R10096 gnd.n2718 gnd.n1398 585
R10097 gnd.n2717 gnd.n1396 585
R10098 gnd.n4903 gnd.n1396 585
R10099 gnd.n2716 gnd.n2715 585
R10100 gnd.n2715 gnd.n1389 585
R10101 gnd.n2714 gnd.n1387 585
R10102 gnd.n4909 gnd.n1387 585
R10103 gnd.n2713 gnd.n2712 585
R10104 gnd.n2712 gnd.n1386 585
R10105 gnd.n2710 gnd.n1378 585
R10106 gnd.n4915 gnd.n1378 585
R10107 gnd.n2709 gnd.n2708 585
R10108 gnd.n2708 gnd.n1371 585
R10109 gnd.n2707 gnd.n1369 585
R10110 gnd.n4921 gnd.n1369 585
R10111 gnd.n2706 gnd.n2705 585
R10112 gnd.n2705 gnd.n1361 585
R10113 gnd.n2703 gnd.n1359 585
R10114 gnd.n4927 gnd.n1359 585
R10115 gnd.n2702 gnd.n2701 585
R10116 gnd.n2701 gnd.n1352 585
R10117 gnd.n2700 gnd.n1350 585
R10118 gnd.n4933 gnd.n1350 585
R10119 gnd.n2699 gnd.n2698 585
R10120 gnd.n2698 gnd.n1349 585
R10121 gnd.n2696 gnd.n1340 585
R10122 gnd.n4939 gnd.n1340 585
R10123 gnd.n2695 gnd.n2694 585
R10124 gnd.n2694 gnd.n1333 585
R10125 gnd.n2693 gnd.n1331 585
R10126 gnd.n4945 gnd.n1331 585
R10127 gnd.n2692 gnd.n2691 585
R10128 gnd.n2691 gnd.n1323 585
R10129 gnd.n2689 gnd.n1321 585
R10130 gnd.n4951 gnd.n1321 585
R10131 gnd.n2688 gnd.n2687 585
R10132 gnd.n2687 gnd.n1314 585
R10133 gnd.n2686 gnd.n1312 585
R10134 gnd.n4957 gnd.n1312 585
R10135 gnd.n2685 gnd.n2684 585
R10136 gnd.n2684 gnd.n1311 585
R10137 gnd.n2682 gnd.n1302 585
R10138 gnd.n4963 gnd.n1302 585
R10139 gnd.n2681 gnd.n2680 585
R10140 gnd.n2680 gnd.n1295 585
R10141 gnd.n2679 gnd.n1293 585
R10142 gnd.n4969 gnd.n1293 585
R10143 gnd.n2678 gnd.n2677 585
R10144 gnd.n2677 gnd.n1285 585
R10145 gnd.n2675 gnd.n1283 585
R10146 gnd.n4975 gnd.n1283 585
R10147 gnd.n2674 gnd.n2673 585
R10148 gnd.n2673 gnd.n1273 585
R10149 gnd.n2672 gnd.n1271 585
R10150 gnd.n4981 gnd.n1271 585
R10151 gnd.n2671 gnd.n1259 585
R10152 gnd.n1270 gnd.n1259 585
R10153 gnd.n4988 gnd.n1257 585
R10154 gnd.n4988 gnd.n4987 585
R10155 gnd.n4990 gnd.n4989 585
R10156 gnd.n4989 gnd.n1186 585
R10157 gnd.n7668 gnd.n245 585
R10158 gnd.n245 gnd.n244 585
R10159 gnd.n7670 gnd.n7669 585
R10160 gnd.n7671 gnd.n7670 585
R10161 gnd.n232 gnd.n231 585
R10162 gnd.n235 gnd.n232 585
R10163 gnd.n7679 gnd.n7678 585
R10164 gnd.n7678 gnd.n7677 585
R10165 gnd.n7680 gnd.n226 585
R10166 gnd.n226 gnd.n225 585
R10167 gnd.n7682 gnd.n7681 585
R10168 gnd.n7683 gnd.n7682 585
R10169 gnd.n213 gnd.n212 585
R10170 gnd.n222 gnd.n213 585
R10171 gnd.n7691 gnd.n7690 585
R10172 gnd.n7690 gnd.n7689 585
R10173 gnd.n7692 gnd.n207 585
R10174 gnd.n207 gnd.n206 585
R10175 gnd.n7694 gnd.n7693 585
R10176 gnd.n7695 gnd.n7694 585
R10177 gnd.n193 gnd.n192 585
R10178 gnd.n197 gnd.n193 585
R10179 gnd.n7703 gnd.n7702 585
R10180 gnd.n7702 gnd.n7701 585
R10181 gnd.n7704 gnd.n187 585
R10182 gnd.n194 gnd.n187 585
R10183 gnd.n7706 gnd.n7705 585
R10184 gnd.n7707 gnd.n7706 585
R10185 gnd.n175 gnd.n174 585
R10186 gnd.n184 gnd.n175 585
R10187 gnd.n7715 gnd.n7714 585
R10188 gnd.n7714 gnd.n7713 585
R10189 gnd.n7716 gnd.n169 585
R10190 gnd.n169 gnd.n168 585
R10191 gnd.n7718 gnd.n7717 585
R10192 gnd.n7719 gnd.n7718 585
R10193 gnd.n155 gnd.n154 585
R10194 gnd.n159 gnd.n155 585
R10195 gnd.n7727 gnd.n7726 585
R10196 gnd.n7726 gnd.n7725 585
R10197 gnd.n7728 gnd.n149 585
R10198 gnd.n156 gnd.n149 585
R10199 gnd.n7730 gnd.n7729 585
R10200 gnd.n7731 gnd.n7730 585
R10201 gnd.n137 gnd.n136 585
R10202 gnd.n146 gnd.n137 585
R10203 gnd.n7739 gnd.n7738 585
R10204 gnd.n7738 gnd.n7737 585
R10205 gnd.n7740 gnd.n132 585
R10206 gnd.n132 gnd.n131 585
R10207 gnd.n7742 gnd.n7741 585
R10208 gnd.n7743 gnd.n7742 585
R10209 gnd.n116 gnd.n114 585
R10210 gnd.n120 gnd.n116 585
R10211 gnd.n7751 gnd.n7750 585
R10212 gnd.n7750 gnd.n7749 585
R10213 gnd.n115 gnd.n107 585
R10214 gnd.n117 gnd.n115 585
R10215 gnd.n7754 gnd.n105 585
R10216 gnd.n105 gnd.n102 585
R10217 gnd.n7756 gnd.n7755 585
R10218 gnd.n7757 gnd.n7756 585
R10219 gnd.n7467 gnd.n104 585
R10220 gnd.n7482 gnd.n104 585
R10221 gnd.n7469 gnd.n7468 585
R10222 gnd.n7469 gnd.n485 585
R10223 gnd.n7472 gnd.n7471 585
R10224 gnd.n7473 gnd.n7472 585
R10225 gnd.n7470 gnd.n7466 585
R10226 gnd.n7466 gnd.n7465 585
R10227 gnd.n7454 gnd.n495 585
R10228 gnd.n7446 gnd.n495 585
R10229 gnd.n7456 gnd.n7455 585
R10230 gnd.n7457 gnd.n7456 585
R10231 gnd.n7453 gnd.n508 585
R10232 gnd.n7453 gnd.n7452 585
R10233 gnd.n7426 gnd.n507 585
R10234 gnd.n7438 gnd.n507 585
R10235 gnd.n7427 gnd.n531 585
R10236 gnd.n7412 gnd.n531 585
R10237 gnd.n7429 gnd.n7428 585
R10238 gnd.n7430 gnd.n7429 585
R10239 gnd.n532 gnd.n530 585
R10240 gnd.n7406 gnd.n530 585
R10241 gnd.n7421 gnd.n7420 585
R10242 gnd.n7420 gnd.n7419 585
R10243 gnd.n535 gnd.n534 585
R10244 gnd.n7402 gnd.n535 585
R10245 gnd.n7390 gnd.n560 585
R10246 gnd.n7376 gnd.n560 585
R10247 gnd.n7392 gnd.n7391 585
R10248 gnd.n7393 gnd.n7392 585
R10249 gnd.n561 gnd.n559 585
R10250 gnd.n7370 gnd.n559 585
R10251 gnd.n7385 gnd.n7384 585
R10252 gnd.n7384 gnd.n7383 585
R10253 gnd.n564 gnd.n563 585
R10254 gnd.n2055 gnd.n564 585
R10255 gnd.n4333 gnd.n4329 585
R10256 gnd.n4329 gnd.n4328 585
R10257 gnd.n4335 gnd.n4334 585
R10258 gnd.n4336 gnd.n4335 585
R10259 gnd.n2039 gnd.n2038 585
R10260 gnd.n4316 gnd.n2039 585
R10261 gnd.n4344 gnd.n4343 585
R10262 gnd.n4343 gnd.n4342 585
R10263 gnd.n4345 gnd.n2033 585
R10264 gnd.n4300 gnd.n2033 585
R10265 gnd.n4347 gnd.n4346 585
R10266 gnd.n4348 gnd.n4347 585
R10267 gnd.n2018 gnd.n2017 585
R10268 gnd.n4285 gnd.n2018 585
R10269 gnd.n4356 gnd.n4355 585
R10270 gnd.n4355 gnd.n4354 585
R10271 gnd.n4357 gnd.n2012 585
R10272 gnd.n4277 gnd.n2012 585
R10273 gnd.n4359 gnd.n4358 585
R10274 gnd.n4360 gnd.n4359 585
R10275 gnd.n1994 gnd.n1993 585
R10276 gnd.n4270 gnd.n1994 585
R10277 gnd.n4368 gnd.n4367 585
R10278 gnd.n4367 gnd.n4366 585
R10279 gnd.n4369 gnd.n1985 585
R10280 gnd.n4262 gnd.n1985 585
R10281 gnd.n4371 gnd.n4370 585
R10282 gnd.n4372 gnd.n4371 585
R10283 gnd.n1986 gnd.n1984 585
R10284 gnd.n4238 gnd.n1984 585
R10285 gnd.n1987 gnd.n1906 585
R10286 gnd.n4380 gnd.n1906 585
R10287 gnd.n4499 gnd.n4498 585
R10288 gnd.n4497 gnd.n1905 585
R10289 gnd.n4496 gnd.n1904 585
R10290 gnd.n4501 gnd.n1904 585
R10291 gnd.n4495 gnd.n4494 585
R10292 gnd.n4493 gnd.n4492 585
R10293 gnd.n4491 gnd.n4490 585
R10294 gnd.n4489 gnd.n4488 585
R10295 gnd.n4487 gnd.n4486 585
R10296 gnd.n4485 gnd.n4484 585
R10297 gnd.n4483 gnd.n4482 585
R10298 gnd.n4481 gnd.n4480 585
R10299 gnd.n4479 gnd.n4478 585
R10300 gnd.n4477 gnd.n4476 585
R10301 gnd.n4475 gnd.n4474 585
R10302 gnd.n4473 gnd.n4472 585
R10303 gnd.n4471 gnd.n4470 585
R10304 gnd.n4469 gnd.n4468 585
R10305 gnd.n4467 gnd.n4466 585
R10306 gnd.n4464 gnd.n4463 585
R10307 gnd.n4462 gnd.n4461 585
R10308 gnd.n4460 gnd.n4459 585
R10309 gnd.n4458 gnd.n4457 585
R10310 gnd.n4456 gnd.n4455 585
R10311 gnd.n4454 gnd.n4453 585
R10312 gnd.n4452 gnd.n4451 585
R10313 gnd.n4450 gnd.n4449 585
R10314 gnd.n4447 gnd.n4446 585
R10315 gnd.n4445 gnd.n4444 585
R10316 gnd.n4443 gnd.n4442 585
R10317 gnd.n4441 gnd.n4440 585
R10318 gnd.n4439 gnd.n4438 585
R10319 gnd.n4437 gnd.n4436 585
R10320 gnd.n4435 gnd.n4434 585
R10321 gnd.n4433 gnd.n4432 585
R10322 gnd.n4431 gnd.n4430 585
R10323 gnd.n4429 gnd.n4428 585
R10324 gnd.n4427 gnd.n4426 585
R10325 gnd.n4425 gnd.n4424 585
R10326 gnd.n4423 gnd.n4422 585
R10327 gnd.n4421 gnd.n4420 585
R10328 gnd.n4419 gnd.n4418 585
R10329 gnd.n4417 gnd.n4416 585
R10330 gnd.n4415 gnd.n4414 585
R10331 gnd.n4413 gnd.n4412 585
R10332 gnd.n4411 gnd.n4410 585
R10333 gnd.n4409 gnd.n4408 585
R10334 gnd.n4407 gnd.n4406 585
R10335 gnd.n4405 gnd.n4404 585
R10336 gnd.n4403 gnd.n4402 585
R10337 gnd.n4401 gnd.n4400 585
R10338 gnd.n4399 gnd.n4398 585
R10339 gnd.n4397 gnd.n4396 585
R10340 gnd.n4395 gnd.n4394 585
R10341 gnd.n4393 gnd.n4392 585
R10342 gnd.n4391 gnd.n4390 585
R10343 gnd.n4389 gnd.n4388 585
R10344 gnd.n4383 gnd.n4382 585
R10345 gnd.n7539 gnd.n345 585
R10346 gnd.n7547 gnd.n7546 585
R10347 gnd.n7549 gnd.n7548 585
R10348 gnd.n7551 gnd.n7550 585
R10349 gnd.n7553 gnd.n7552 585
R10350 gnd.n7555 gnd.n7554 585
R10351 gnd.n7557 gnd.n7556 585
R10352 gnd.n7559 gnd.n7558 585
R10353 gnd.n7561 gnd.n7560 585
R10354 gnd.n7563 gnd.n7562 585
R10355 gnd.n7565 gnd.n7564 585
R10356 gnd.n7567 gnd.n7566 585
R10357 gnd.n7569 gnd.n7568 585
R10358 gnd.n7571 gnd.n7570 585
R10359 gnd.n7573 gnd.n7572 585
R10360 gnd.n7575 gnd.n7574 585
R10361 gnd.n7577 gnd.n7576 585
R10362 gnd.n7579 gnd.n7578 585
R10363 gnd.n7581 gnd.n7580 585
R10364 gnd.n7584 gnd.n7583 585
R10365 gnd.n7582 gnd.n325 585
R10366 gnd.n7589 gnd.n7588 585
R10367 gnd.n7591 gnd.n7590 585
R10368 gnd.n7593 gnd.n7592 585
R10369 gnd.n7595 gnd.n7594 585
R10370 gnd.n7597 gnd.n7596 585
R10371 gnd.n7599 gnd.n7598 585
R10372 gnd.n7601 gnd.n7600 585
R10373 gnd.n7603 gnd.n7602 585
R10374 gnd.n7605 gnd.n7604 585
R10375 gnd.n7607 gnd.n7606 585
R10376 gnd.n7609 gnd.n7608 585
R10377 gnd.n7611 gnd.n7610 585
R10378 gnd.n7613 gnd.n7612 585
R10379 gnd.n7615 gnd.n7614 585
R10380 gnd.n7617 gnd.n7616 585
R10381 gnd.n7619 gnd.n7618 585
R10382 gnd.n7621 gnd.n7620 585
R10383 gnd.n7623 gnd.n7622 585
R10384 gnd.n7625 gnd.n7624 585
R10385 gnd.n7627 gnd.n7626 585
R10386 gnd.n7632 gnd.n7631 585
R10387 gnd.n7634 gnd.n7633 585
R10388 gnd.n7636 gnd.n7635 585
R10389 gnd.n7638 gnd.n7637 585
R10390 gnd.n7640 gnd.n7639 585
R10391 gnd.n7642 gnd.n7641 585
R10392 gnd.n7644 gnd.n7643 585
R10393 gnd.n7646 gnd.n7645 585
R10394 gnd.n7648 gnd.n7647 585
R10395 gnd.n7650 gnd.n7649 585
R10396 gnd.n7652 gnd.n7651 585
R10397 gnd.n7654 gnd.n7653 585
R10398 gnd.n7656 gnd.n7655 585
R10399 gnd.n7658 gnd.n7657 585
R10400 gnd.n7659 gnd.n289 585
R10401 gnd.n7661 gnd.n7660 585
R10402 gnd.n250 gnd.n249 585
R10403 gnd.n7665 gnd.n7664 585
R10404 gnd.n7664 gnd.n7663 585
R10405 gnd.n7541 gnd.n7540 585
R10406 gnd.n7540 gnd.n244 585
R10407 gnd.n7538 gnd.n242 585
R10408 gnd.n7671 gnd.n242 585
R10409 gnd.n7537 gnd.n7536 585
R10410 gnd.n7536 gnd.n235 585
R10411 gnd.n7535 gnd.n233 585
R10412 gnd.n7677 gnd.n233 585
R10413 gnd.n7534 gnd.n7533 585
R10414 gnd.n7533 gnd.n225 585
R10415 gnd.n7531 gnd.n223 585
R10416 gnd.n7683 gnd.n223 585
R10417 gnd.n7530 gnd.n7529 585
R10418 gnd.n7529 gnd.n222 585
R10419 gnd.n7528 gnd.n214 585
R10420 gnd.n7689 gnd.n214 585
R10421 gnd.n7527 gnd.n7526 585
R10422 gnd.n7526 gnd.n206 585
R10423 gnd.n7524 gnd.n204 585
R10424 gnd.n7695 gnd.n204 585
R10425 gnd.n7523 gnd.n7522 585
R10426 gnd.n7522 gnd.n197 585
R10427 gnd.n7521 gnd.n195 585
R10428 gnd.n7701 gnd.n195 585
R10429 gnd.n7520 gnd.n7519 585
R10430 gnd.n7519 gnd.n194 585
R10431 gnd.n7517 gnd.n185 585
R10432 gnd.n7707 gnd.n185 585
R10433 gnd.n7516 gnd.n7515 585
R10434 gnd.n7515 gnd.n184 585
R10435 gnd.n7514 gnd.n176 585
R10436 gnd.n7713 gnd.n176 585
R10437 gnd.n7513 gnd.n7512 585
R10438 gnd.n7512 gnd.n168 585
R10439 gnd.n7510 gnd.n166 585
R10440 gnd.n7719 gnd.n166 585
R10441 gnd.n7509 gnd.n7508 585
R10442 gnd.n7508 gnd.n159 585
R10443 gnd.n7507 gnd.n157 585
R10444 gnd.n7725 gnd.n157 585
R10445 gnd.n7506 gnd.n7505 585
R10446 gnd.n7505 gnd.n156 585
R10447 gnd.n7503 gnd.n147 585
R10448 gnd.n7731 gnd.n147 585
R10449 gnd.n7502 gnd.n7501 585
R10450 gnd.n7501 gnd.n146 585
R10451 gnd.n7500 gnd.n138 585
R10452 gnd.n7737 gnd.n138 585
R10453 gnd.n7499 gnd.n7498 585
R10454 gnd.n7498 gnd.n131 585
R10455 gnd.n7496 gnd.n129 585
R10456 gnd.n7743 gnd.n129 585
R10457 gnd.n7495 gnd.n7494 585
R10458 gnd.n7494 gnd.n120 585
R10459 gnd.n7493 gnd.n118 585
R10460 gnd.n7749 gnd.n118 585
R10461 gnd.n7492 gnd.n7491 585
R10462 gnd.n7491 gnd.n117 585
R10463 gnd.n7490 gnd.n480 585
R10464 gnd.n7490 gnd.n102 585
R10465 gnd.n7479 gnd.n101 585
R10466 gnd.n7757 gnd.n101 585
R10467 gnd.n7481 gnd.n7480 585
R10468 gnd.n7482 gnd.n7481 585
R10469 gnd.n7478 gnd.n486 585
R10470 gnd.n486 gnd.n485 585
R10471 gnd.n491 gnd.n487 585
R10472 gnd.n7473 gnd.n491 585
R10473 gnd.n7443 gnd.n497 585
R10474 gnd.n7465 gnd.n497 585
R10475 gnd.n7445 gnd.n7444 585
R10476 gnd.n7446 gnd.n7445 585
R10477 gnd.n7442 gnd.n505 585
R10478 gnd.n7457 gnd.n505 585
R10479 gnd.n7441 gnd.n510 585
R10480 gnd.n7452 gnd.n510 585
R10481 gnd.n7440 gnd.n7439 585
R10482 gnd.n7439 gnd.n7438 585
R10483 gnd.n519 gnd.n517 585
R10484 gnd.n7412 gnd.n519 585
R10485 gnd.n7409 gnd.n527 585
R10486 gnd.n7430 gnd.n527 585
R10487 gnd.n7408 gnd.n7407 585
R10488 gnd.n7407 gnd.n7406 585
R10489 gnd.n7405 gnd.n537 585
R10490 gnd.n7419 gnd.n537 585
R10491 gnd.n7404 gnd.n7403 585
R10492 gnd.n7403 gnd.n7402 585
R10493 gnd.n547 gnd.n545 585
R10494 gnd.n7376 gnd.n547 585
R10495 gnd.n7373 gnd.n556 585
R10496 gnd.n7393 gnd.n556 585
R10497 gnd.n7372 gnd.n7371 585
R10498 gnd.n7371 gnd.n7370 585
R10499 gnd.n573 gnd.n566 585
R10500 gnd.n7383 gnd.n566 585
R10501 gnd.n4293 gnd.n4292 585
R10502 gnd.n4292 gnd.n2055 585
R10503 gnd.n4294 gnd.n2053 585
R10504 gnd.n4328 gnd.n2053 585
R10505 gnd.n4295 gnd.n2050 585
R10506 gnd.n4336 gnd.n2050 585
R10507 gnd.n4296 gnd.n2061 585
R10508 gnd.n4316 gnd.n2061 585
R10509 gnd.n4297 gnd.n2041 585
R10510 gnd.n4342 gnd.n2041 585
R10511 gnd.n4299 gnd.n4298 585
R10512 gnd.n4300 gnd.n4299 585
R10513 gnd.n4288 gnd.n2030 585
R10514 gnd.n4348 gnd.n2030 585
R10515 gnd.n4287 gnd.n4286 585
R10516 gnd.n4286 gnd.n4285 585
R10517 gnd.n2066 gnd.n2020 585
R10518 gnd.n4354 gnd.n2020 585
R10519 gnd.n4276 gnd.n4275 585
R10520 gnd.n4277 gnd.n4276 585
R10521 gnd.n4273 gnd.n2009 585
R10522 gnd.n4360 gnd.n2009 585
R10523 gnd.n4272 gnd.n4271 585
R10524 gnd.n4271 gnd.n4270 585
R10525 gnd.n2070 gnd.n1996 585
R10526 gnd.n4366 gnd.n1996 585
R10527 gnd.n1980 gnd.n1979 585
R10528 gnd.n4262 gnd.n1980 585
R10529 gnd.n4374 gnd.n4373 585
R10530 gnd.n4373 gnd.n4372 585
R10531 gnd.n4375 gnd.n1969 585
R10532 gnd.n4238 gnd.n1969 585
R10533 gnd.n4381 gnd.n1970 585
R10534 gnd.n4381 gnd.n4380 585
R10535 gnd.n2659 gnd.n2658 585
R10536 gnd.n2660 gnd.n2659 585
R10537 gnd.n7347 gnd.n7346 585
R10538 gnd.n7347 gnd.n494 585
R10539 gnd.n7348 gnd.n592 585
R10540 gnd.n7348 gnd.n496 585
R10541 gnd.n7350 gnd.n7349 585
R10542 gnd.n7349 gnd.n516 585
R10543 gnd.n7353 gnd.n591 585
R10544 gnd.n591 gnd.n504 585
R10545 gnd.n7354 gnd.n587 585
R10546 gnd.n587 gnd.n509 585
R10547 gnd.n7356 gnd.n7355 585
R10548 gnd.n7356 gnd.n520 585
R10549 gnd.n7357 gnd.n586 585
R10550 gnd.n7357 gnd.n528 585
R10551 gnd.n7359 gnd.n7358 585
R10552 gnd.n7358 gnd.n526 585
R10553 gnd.n7360 gnd.n581 585
R10554 gnd.n581 gnd.n539 585
R10555 gnd.n7362 gnd.n7361 585
R10556 gnd.n7362 gnd.n536 585
R10557 gnd.n7363 gnd.n580 585
R10558 gnd.n7363 gnd.n548 585
R10559 gnd.n7365 gnd.n7364 585
R10560 gnd.n7364 gnd.n557 585
R10561 gnd.n7366 gnd.n575 585
R10562 gnd.n575 gnd.n555 585
R10563 gnd.n7368 gnd.n7367 585
R10564 gnd.n7369 gnd.n7368 585
R10565 gnd.n576 gnd.n574 585
R10566 gnd.n574 gnd.n565 585
R10567 gnd.n4326 gnd.n4325 585
R10568 gnd.n4327 gnd.n4326 585
R10569 gnd.n2057 gnd.n2056 585
R10570 gnd.n2056 gnd.n2052 585
R10571 gnd.n4320 gnd.n4319 585
R10572 gnd.n4319 gnd.n2049 585
R10573 gnd.n4318 gnd.n2059 585
R10574 gnd.n4318 gnd.n4317 585
R10575 gnd.n4223 gnd.n2060 585
R10576 gnd.n2060 gnd.n2040 585
R10577 gnd.n4225 gnd.n4224 585
R10578 gnd.n4225 gnd.n2032 585
R10579 gnd.n4227 gnd.n4226 585
R10580 gnd.n4226 gnd.n2029 585
R10581 gnd.n4228 gnd.n4216 585
R10582 gnd.n4216 gnd.n2022 585
R10583 gnd.n4230 gnd.n4229 585
R10584 gnd.n4230 gnd.n2019 585
R10585 gnd.n4231 gnd.n4215 585
R10586 gnd.n4231 gnd.n2011 585
R10587 gnd.n4233 gnd.n4232 585
R10588 gnd.n4232 gnd.n2008 585
R10589 gnd.n4234 gnd.n4210 585
R10590 gnd.n4210 gnd.n1998 585
R10591 gnd.n4236 gnd.n4235 585
R10592 gnd.n4236 gnd.n1995 585
R10593 gnd.n4237 gnd.n4209 585
R10594 gnd.n4237 gnd.n1982 585
R10595 gnd.n4241 gnd.n4240 585
R10596 gnd.n4240 gnd.n4239 585
R10597 gnd.n4242 gnd.n4204 585
R10598 gnd.n4204 gnd.n1973 585
R10599 gnd.n4244 gnd.n4243 585
R10600 gnd.n4244 gnd.n1971 585
R10601 gnd.n4245 gnd.n4203 585
R10602 gnd.n4245 gnd.n1903 585
R10603 gnd.n4247 gnd.n4246 585
R10604 gnd.n4246 gnd.n1861 585
R10605 gnd.n4248 gnd.n2103 585
R10606 gnd.n2103 gnd.n2101 585
R10607 gnd.n4250 gnd.n4249 585
R10608 gnd.n4251 gnd.n4250 585
R10609 gnd.n2104 gnd.n2102 585
R10610 gnd.n2102 gnd.n1794 585
R10611 gnd.n4197 gnd.n1793 585
R10612 gnd.n4569 gnd.n1793 585
R10613 gnd.n4196 gnd.n4195 585
R10614 gnd.n4195 gnd.n1792 585
R10615 gnd.n4194 gnd.n2106 585
R10616 gnd.n4194 gnd.n4193 585
R10617 gnd.n4182 gnd.n2107 585
R10618 gnd.n2108 gnd.n2107 585
R10619 gnd.n4184 gnd.n4183 585
R10620 gnd.n4185 gnd.n4184 585
R10621 gnd.n2117 gnd.n2116 585
R10622 gnd.n2116 gnd.n2115 585
R10623 gnd.n4176 gnd.n4175 585
R10624 gnd.n4175 gnd.n4174 585
R10625 gnd.n2120 gnd.n2119 585
R10626 gnd.n2127 gnd.n2120 585
R10627 gnd.n4165 gnd.n4164 585
R10628 gnd.n4166 gnd.n4165 585
R10629 gnd.n2130 gnd.n2129 585
R10630 gnd.n2138 gnd.n2129 585
R10631 gnd.n4160 gnd.n4159 585
R10632 gnd.n4159 gnd.n4158 585
R10633 gnd.n2133 gnd.n2132 585
R10634 gnd.n3945 gnd.n2133 585
R10635 gnd.n4018 gnd.n4017 585
R10636 gnd.n4019 gnd.n4018 585
R10637 gnd.n2219 gnd.n2218 585
R10638 gnd.n2227 gnd.n2218 585
R10639 gnd.n4013 gnd.n4012 585
R10640 gnd.n4012 gnd.n4011 585
R10641 gnd.n2222 gnd.n2221 585
R10642 gnd.n2231 gnd.n2222 585
R10643 gnd.n3981 gnd.n2247 585
R10644 gnd.n2247 gnd.n2237 585
R10645 gnd.n3983 gnd.n3982 585
R10646 gnd.n3984 gnd.n3983 585
R10647 gnd.n2248 gnd.n2246 585
R10648 gnd.n2246 gnd.n2241 585
R10649 gnd.n3976 gnd.n3975 585
R10650 gnd.n3975 gnd.n3974 585
R10651 gnd.n2251 gnd.n2250 585
R10652 gnd.n3966 gnd.n2251 585
R10653 gnd.n3929 gnd.n2268 585
R10654 gnd.n3854 gnd.n2268 585
R10655 gnd.n3931 gnd.n3930 585
R10656 gnd.n3932 gnd.n3931 585
R10657 gnd.n2269 gnd.n2267 585
R10658 gnd.n2276 gnd.n2267 585
R10659 gnd.n3924 gnd.n3923 585
R10660 gnd.n3923 gnd.n3922 585
R10661 gnd.n2272 gnd.n2271 585
R10662 gnd.n3909 gnd.n2272 585
R10663 gnd.n3896 gnd.n2291 585
R10664 gnd.n3879 gnd.n2291 585
R10665 gnd.n3898 gnd.n3897 585
R10666 gnd.n3899 gnd.n3898 585
R10667 gnd.n2292 gnd.n2290 585
R10668 gnd.n2299 gnd.n2290 585
R10669 gnd.n3891 gnd.n3890 585
R10670 gnd.n3890 gnd.n3889 585
R10671 gnd.n2295 gnd.n2294 585
R10672 gnd.n2308 gnd.n2295 585
R10673 gnd.n3835 gnd.n3834 585
R10674 gnd.n3836 gnd.n3835 585
R10675 gnd.n2317 gnd.n2316 585
R10676 gnd.n2324 gnd.n2316 585
R10677 gnd.n3830 gnd.n3829 585
R10678 gnd.n3829 gnd.n3828 585
R10679 gnd.n2320 gnd.n2319 585
R10680 gnd.n2328 gnd.n2320 585
R10681 gnd.n3798 gnd.n2342 585
R10682 gnd.n2342 gnd.n2335 585
R10683 gnd.n3800 gnd.n3799 585
R10684 gnd.n3801 gnd.n3800 585
R10685 gnd.n2343 gnd.n2341 585
R10686 gnd.n3756 gnd.n2341 585
R10687 gnd.n3793 gnd.n3792 585
R10688 gnd.n3792 gnd.n3791 585
R10689 gnd.n2346 gnd.n2345 585
R10690 gnd.n3783 gnd.n2346 585
R10691 gnd.n3746 gnd.n2367 585
R10692 gnd.n2367 gnd.n2366 585
R10693 gnd.n3748 gnd.n3747 585
R10694 gnd.n3749 gnd.n3748 585
R10695 gnd.n2368 gnd.n2365 585
R10696 gnd.n2374 gnd.n2365 585
R10697 gnd.n3741 gnd.n3740 585
R10698 gnd.n3740 gnd.n3739 585
R10699 gnd.n2371 gnd.n2370 585
R10700 gnd.n3726 gnd.n2371 585
R10701 gnd.n3674 gnd.n2412 585
R10702 gnd.n3674 gnd.n3673 585
R10703 gnd.n3675 gnd.n2409 585
R10704 gnd.n3675 gnd.n2385 585
R10705 gnd.n3677 gnd.n3676 585
R10706 gnd.n3676 gnd.n2389 585
R10707 gnd.n3678 gnd.n2404 585
R10708 gnd.n2404 gnd.n2395 585
R10709 gnd.n3680 gnd.n3679 585
R10710 gnd.n3681 gnd.n3680 585
R10711 gnd.n2405 gnd.n2403 585
R10712 gnd.n2403 gnd.n2399 585
R10713 gnd.n3652 gnd.n3651 585
R10714 gnd.n3653 gnd.n3652 585
R10715 gnd.n2424 gnd.n2423 585
R10716 gnd.n2435 gnd.n2423 585
R10717 gnd.n3646 gnd.n3645 585
R10718 gnd.n3645 gnd.n3644 585
R10719 gnd.n2427 gnd.n2426 585
R10720 gnd.n3623 gnd.n2427 585
R10721 gnd.n3611 gnd.n2451 585
R10722 gnd.n2466 gnd.n2451 585
R10723 gnd.n3613 gnd.n3612 585
R10724 gnd.n3614 gnd.n3613 585
R10725 gnd.n2452 gnd.n2450 585
R10726 gnd.n3587 gnd.n2450 585
R10727 gnd.n3606 gnd.n3605 585
R10728 gnd.n3605 gnd.n3604 585
R10729 gnd.n2455 gnd.n2454 585
R10730 gnd.n2470 gnd.n2455 585
R10731 gnd.n3572 gnd.n3571 585
R10732 gnd.n3573 gnd.n3572 585
R10733 gnd.n2480 gnd.n2479 585
R10734 gnd.n2479 gnd.n2475 585
R10735 gnd.n3567 gnd.n3566 585
R10736 gnd.n3566 gnd.n3565 585
R10737 gnd.n2483 gnd.n2482 585
R10738 gnd.n3557 gnd.n2483 585
R10739 gnd.n3535 gnd.n2501 585
R10740 gnd.n3492 gnd.n2501 585
R10741 gnd.n3537 gnd.n3536 585
R10742 gnd.n3538 gnd.n3537 585
R10743 gnd.n2502 gnd.n2500 585
R10744 gnd.n3508 gnd.n2500 585
R10745 gnd.n3530 gnd.n3529 585
R10746 gnd.n3529 gnd.n3528 585
R10747 gnd.n2506 gnd.n2505 585
R10748 gnd.n2514 gnd.n2506 585
R10749 gnd.n1696 gnd.n1695 585
R10750 gnd.n2520 gnd.n1696 585
R10751 gnd.n4681 gnd.n4680 585
R10752 gnd.n4680 gnd.n4679 585
R10753 gnd.n4682 gnd.n1690 585
R10754 gnd.n3404 gnd.n1690 585
R10755 gnd.n4684 gnd.n4683 585
R10756 gnd.n4685 gnd.n4684 585
R10757 gnd.n1691 gnd.n1689 585
R10758 gnd.n1689 gnd.n1684 585
R10759 gnd.n3373 gnd.n3372 585
R10760 gnd.n3373 gnd.n1658 585
R10761 gnd.n3375 gnd.n3374 585
R10762 gnd.n3374 gnd.n1626 585
R10763 gnd.n3376 gnd.n2537 585
R10764 gnd.n2537 gnd.n2534 585
R10765 gnd.n3378 gnd.n3377 585
R10766 gnd.n3379 gnd.n3378 585
R10767 gnd.n2538 gnd.n2536 585
R10768 gnd.n2536 gnd.n2533 585
R10769 gnd.n3364 gnd.n3363 585
R10770 gnd.n3363 gnd.n3362 585
R10771 gnd.n2541 gnd.n2540 585
R10772 gnd.n2542 gnd.n2541 585
R10773 gnd.n3336 gnd.n3335 585
R10774 gnd.n3337 gnd.n3336 585
R10775 gnd.n2554 gnd.n2553 585
R10776 gnd.n2553 gnd.n2551 585
R10777 gnd.n3331 gnd.n3330 585
R10778 gnd.n3330 gnd.n3329 585
R10779 gnd.n2557 gnd.n2556 585
R10780 gnd.n3328 gnd.n2557 585
R10781 gnd.n3311 gnd.n3310 585
R10782 gnd.n3311 gnd.n2558 585
R10783 gnd.n3313 gnd.n3312 585
R10784 gnd.n3312 gnd.n1563 585
R10785 gnd.n3314 gnd.n2583 585
R10786 gnd.n2583 gnd.n1552 585
R10787 gnd.n3316 gnd.n3315 585
R10788 gnd.n3317 gnd.n3316 585
R10789 gnd.n2584 gnd.n2582 585
R10790 gnd.n2582 gnd.n1545 585
R10791 gnd.n3303 gnd.n3302 585
R10792 gnd.n3302 gnd.n1542 585
R10793 gnd.n3301 gnd.n2586 585
R10794 gnd.n3301 gnd.n1535 585
R10795 gnd.n3300 gnd.n3299 585
R10796 gnd.n3300 gnd.n1532 585
R10797 gnd.n2588 gnd.n2587 585
R10798 gnd.n2587 gnd.n1524 585
R10799 gnd.n3295 gnd.n3294 585
R10800 gnd.n3294 gnd.n1521 585
R10801 gnd.n3293 gnd.n2590 585
R10802 gnd.n3293 gnd.n3292 585
R10803 gnd.n3006 gnd.n2591 585
R10804 gnd.n2591 gnd.n1512 585
R10805 gnd.n3007 gnd.n2605 585
R10806 gnd.n2605 gnd.n1504 585
R10807 gnd.n3009 gnd.n3008 585
R10808 gnd.n3010 gnd.n3009 585
R10809 gnd.n2606 gnd.n2604 585
R10810 gnd.n2604 gnd.n1495 585
R10811 gnd.n3000 gnd.n2999 585
R10812 gnd.n2999 gnd.n1492 585
R10813 gnd.n2998 gnd.n2608 585
R10814 gnd.n2998 gnd.n1484 585
R10815 gnd.n2997 gnd.n2996 585
R10816 gnd.n2997 gnd.n1481 585
R10817 gnd.n2610 gnd.n2609 585
R10818 gnd.n2963 gnd.n2609 585
R10819 gnd.n2992 gnd.n2991 585
R10820 gnd.n2991 gnd.n1472 585
R10821 gnd.n2990 gnd.n2612 585
R10822 gnd.n2990 gnd.n1464 585
R10823 gnd.n2989 gnd.n2614 585
R10824 gnd.n2989 gnd.n2988 585
R10825 gnd.n2917 gnd.n2613 585
R10826 gnd.n2613 gnd.n1455 585
R10827 gnd.n2919 gnd.n2918 585
R10828 gnd.n2918 gnd.n1452 585
R10829 gnd.n2920 gnd.n2910 585
R10830 gnd.n2910 gnd.n1444 585
R10831 gnd.n2922 gnd.n2921 585
R10832 gnd.n2922 gnd.n1441 585
R10833 gnd.n2923 gnd.n2909 585
R10834 gnd.n2923 gnd.n2628 585
R10835 gnd.n2925 gnd.n2924 585
R10836 gnd.n2924 gnd.n1432 585
R10837 gnd.n2926 gnd.n2636 585
R10838 gnd.n2636 gnd.n1425 585
R10839 gnd.n2928 gnd.n2927 585
R10840 gnd.n2929 gnd.n2928 585
R10841 gnd.n2637 gnd.n2635 585
R10842 gnd.n2635 gnd.n1414 585
R10843 gnd.n2903 gnd.n2902 585
R10844 gnd.n2902 gnd.n1411 585
R10845 gnd.n2901 gnd.n2639 585
R10846 gnd.n2901 gnd.n2900 585
R10847 gnd.n2655 gnd.n2640 585
R10848 gnd.n2649 gnd.n2640 585
R10849 gnd.n4568 gnd.n4567 585
R10850 gnd.n4569 gnd.n4568 585
R10851 gnd.n1797 gnd.n1795 585
R10852 gnd.n1795 gnd.n1792 585
R10853 gnd.n4192 gnd.n4191 585
R10854 gnd.n4193 gnd.n4192 585
R10855 gnd.n2110 gnd.n2109 585
R10856 gnd.n2109 gnd.n2108 585
R10857 gnd.n4187 gnd.n4186 585
R10858 gnd.n4186 gnd.n4185 585
R10859 gnd.n2113 gnd.n2112 585
R10860 gnd.n2115 gnd.n2113 585
R10861 gnd.n4173 gnd.n4172 585
R10862 gnd.n4174 gnd.n4173 585
R10863 gnd.n2122 gnd.n2121 585
R10864 gnd.n2127 gnd.n2121 585
R10865 gnd.n4168 gnd.n4167 585
R10866 gnd.n4167 gnd.n4166 585
R10867 gnd.n2125 gnd.n2124 585
R10868 gnd.n2138 gnd.n2125 585
R10869 gnd.n3948 gnd.n2135 585
R10870 gnd.n4158 gnd.n2135 585
R10871 gnd.n3947 gnd.n3946 585
R10872 gnd.n3946 gnd.n3945 585
R10873 gnd.n3952 gnd.n2217 585
R10874 gnd.n4019 gnd.n2217 585
R10875 gnd.n3953 gnd.n3943 585
R10876 gnd.n3943 gnd.n2227 585
R10877 gnd.n3954 gnd.n2224 585
R10878 gnd.n4011 gnd.n2224 585
R10879 gnd.n3941 gnd.n3940 585
R10880 gnd.n3940 gnd.n2231 585
R10881 gnd.n3958 gnd.n3939 585
R10882 gnd.n3939 gnd.n2237 585
R10883 gnd.n3959 gnd.n2243 585
R10884 gnd.n3984 gnd.n2243 585
R10885 gnd.n3960 gnd.n3938 585
R10886 gnd.n3938 gnd.n2241 585
R10887 gnd.n2261 gnd.n2253 585
R10888 gnd.n3974 gnd.n2253 585
R10889 gnd.n3965 gnd.n3964 585
R10890 gnd.n3966 gnd.n3965 585
R10891 gnd.n2260 gnd.n2259 585
R10892 gnd.n3854 gnd.n2259 585
R10893 gnd.n3934 gnd.n3933 585
R10894 gnd.n3933 gnd.n3932 585
R10895 gnd.n2264 gnd.n2263 585
R10896 gnd.n2276 gnd.n2264 585
R10897 gnd.n2285 gnd.n2274 585
R10898 gnd.n3922 gnd.n2274 585
R10899 gnd.n3907 gnd.n3906 585
R10900 gnd.n3909 gnd.n3907 585
R10901 gnd.n2284 gnd.n2283 585
R10902 gnd.n3879 gnd.n2283 585
R10903 gnd.n3901 gnd.n3900 585
R10904 gnd.n3900 gnd.n3899 585
R10905 gnd.n2288 gnd.n2287 585
R10906 gnd.n2299 gnd.n2288 585
R10907 gnd.n3765 gnd.n2297 585
R10908 gnd.n3889 gnd.n2297 585
R10909 gnd.n3764 gnd.n3763 585
R10910 gnd.n3763 gnd.n2308 585
R10911 gnd.n3769 gnd.n2314 585
R10912 gnd.n3836 gnd.n2314 585
R10913 gnd.n3770 gnd.n3762 585
R10914 gnd.n3762 gnd.n2324 585
R10915 gnd.n3771 gnd.n2322 585
R10916 gnd.n3828 gnd.n2322 585
R10917 gnd.n3760 gnd.n3759 585
R10918 gnd.n3759 gnd.n2328 585
R10919 gnd.n3775 gnd.n3758 585
R10920 gnd.n3758 gnd.n2335 585
R10921 gnd.n3776 gnd.n2340 585
R10922 gnd.n3801 gnd.n2340 585
R10923 gnd.n3777 gnd.n3757 585
R10924 gnd.n3757 gnd.n3756 585
R10925 gnd.n2358 gnd.n2348 585
R10926 gnd.n3791 gnd.n2348 585
R10927 gnd.n3782 gnd.n3781 585
R10928 gnd.n3783 gnd.n3782 585
R10929 gnd.n2357 gnd.n2356 585
R10930 gnd.n2366 gnd.n2356 585
R10931 gnd.n3751 gnd.n3750 585
R10932 gnd.n3750 gnd.n3749 585
R10933 gnd.n2361 gnd.n2360 585
R10934 gnd.n2374 gnd.n2361 585
R10935 gnd.n3666 gnd.n2372 585
R10936 gnd.n3739 gnd.n2372 585
R10937 gnd.n2415 gnd.n2382 585
R10938 gnd.n3726 gnd.n2382 585
R10939 gnd.n3671 gnd.n3670 585
R10940 gnd.n3673 gnd.n3671 585
R10941 gnd.n2414 gnd.n2413 585
R10942 gnd.n2413 gnd.n2385 585
R10943 gnd.n3663 gnd.n3662 585
R10944 gnd.n3662 gnd.n2389 585
R10945 gnd.n3661 gnd.n3660 585
R10946 gnd.n3661 gnd.n2395 585
R10947 gnd.n3659 gnd.n2401 585
R10948 gnd.n3681 gnd.n2401 585
R10949 gnd.n2421 gnd.n2417 585
R10950 gnd.n2421 gnd.n2399 585
R10951 gnd.n3655 gnd.n3654 585
R10952 gnd.n3654 gnd.n3653 585
R10953 gnd.n2420 gnd.n2419 585
R10954 gnd.n2435 gnd.n2420 585
R10955 gnd.n2444 gnd.n2428 585
R10956 gnd.n3644 gnd.n2428 585
R10957 gnd.n3622 gnd.n3621 585
R10958 gnd.n3623 gnd.n3622 585
R10959 gnd.n2443 gnd.n2442 585
R10960 gnd.n2466 gnd.n2442 585
R10961 gnd.n3616 gnd.n3615 585
R10962 gnd.n3615 gnd.n3614 585
R10963 gnd.n2447 gnd.n2446 585
R10964 gnd.n3587 gnd.n2447 585
R10965 gnd.n3546 gnd.n2457 585
R10966 gnd.n3604 gnd.n2457 585
R10967 gnd.n3549 gnd.n3545 585
R10968 gnd.n3545 gnd.n2470 585
R10969 gnd.n3550 gnd.n2477 585
R10970 gnd.n3573 gnd.n2477 585
R10971 gnd.n3551 gnd.n3544 585
R10972 gnd.n3544 gnd.n2475 585
R10973 gnd.n2493 gnd.n2485 585
R10974 gnd.n3565 gnd.n2485 585
R10975 gnd.n3556 gnd.n3555 585
R10976 gnd.n3557 gnd.n3556 585
R10977 gnd.n2492 gnd.n2491 585
R10978 gnd.n3492 gnd.n2491 585
R10979 gnd.n3540 gnd.n3539 585
R10980 gnd.n3539 gnd.n3538 585
R10981 gnd.n2496 gnd.n2495 585
R10982 gnd.n3508 gnd.n2496 585
R10983 gnd.n3396 gnd.n2508 585
R10984 gnd.n3528 gnd.n2508 585
R10985 gnd.n3397 gnd.n3394 585
R10986 gnd.n3394 gnd.n2514 585
R10987 gnd.n3398 gnd.n3393 585
R10988 gnd.n3393 gnd.n2520 585
R10989 gnd.n2525 gnd.n1697 585
R10990 gnd.n4679 gnd.n1697 585
R10991 gnd.n3403 gnd.n3402 585
R10992 gnd.n3404 gnd.n3403 585
R10993 gnd.n2524 gnd.n1686 585
R10994 gnd.n4685 gnd.n1686 585
R10995 gnd.n3389 gnd.n3388 585
R10996 gnd.n3388 gnd.n1684 585
R10997 gnd.n3387 gnd.n2527 585
R10998 gnd.n3387 gnd.n1658 585
R10999 gnd.n3386 gnd.n3385 585
R11000 gnd.n3386 gnd.n1626 585
R11001 gnd.n2529 gnd.n2528 585
R11002 gnd.n2534 gnd.n2528 585
R11003 gnd.n3381 gnd.n3380 585
R11004 gnd.n3380 gnd.n3379 585
R11005 gnd.n2532 gnd.n2531 585
R11006 gnd.n2533 gnd.n2532 585
R11007 gnd.n3040 gnd.n2543 585
R11008 gnd.n3362 gnd.n2543 585
R11009 gnd.n3041 gnd.n3039 585
R11010 gnd.n3039 gnd.n2542 585
R11011 gnd.n3037 gnd.n2552 585
R11012 gnd.n3337 gnd.n2552 585
R11013 gnd.n3046 gnd.n3045 585
R11014 gnd.n3046 gnd.n2551 585
R11015 gnd.n3048 gnd.n3047 585
R11016 gnd.n3050 gnd.n3049 585
R11017 gnd.n3052 gnd.n3051 585
R11018 gnd.n3033 gnd.n3032 585
R11019 gnd.n3056 gnd.n3034 585
R11020 gnd.n3058 gnd.n3057 585
R11021 gnd.n3173 gnd.n3059 585
R11022 gnd.n3172 gnd.n3060 585
R11023 gnd.n3171 gnd.n3061 585
R11024 gnd.n3067 gnd.n3062 585
R11025 gnd.n3164 gnd.n3068 585
R11026 gnd.n3163 gnd.n3069 585
R11027 gnd.n3071 gnd.n3070 585
R11028 gnd.n3156 gnd.n3079 585
R11029 gnd.n3155 gnd.n3080 585
R11030 gnd.n3087 gnd.n3081 585
R11031 gnd.n3148 gnd.n3088 585
R11032 gnd.n3147 gnd.n3089 585
R11033 gnd.n3091 gnd.n3090 585
R11034 gnd.n3140 gnd.n3099 585
R11035 gnd.n3139 gnd.n3100 585
R11036 gnd.n3107 gnd.n3101 585
R11037 gnd.n3132 gnd.n3108 585
R11038 gnd.n3131 gnd.n3109 585
R11039 gnd.n3111 gnd.n3110 585
R11040 gnd.n3124 gnd.n3121 585
R11041 gnd.n3123 gnd.n3122 585
R11042 gnd.n2574 gnd.n2573 585
R11043 gnd.n3327 gnd.n3326 585
R11044 gnd.n3328 gnd.n3327 585
R11045 gnd.n4571 gnd.n4570 585
R11046 gnd.n4570 gnd.n4569 585
R11047 gnd.n1790 gnd.n1788 585
R11048 gnd.n1792 gnd.n1790 585
R11049 gnd.n4575 gnd.n1787 585
R11050 gnd.n4193 gnd.n1787 585
R11051 gnd.n4576 gnd.n1786 585
R11052 gnd.n2108 gnd.n1786 585
R11053 gnd.n4577 gnd.n1785 585
R11054 gnd.n4185 gnd.n1785 585
R11055 gnd.n2114 gnd.n1783 585
R11056 gnd.n2115 gnd.n2114 585
R11057 gnd.n4581 gnd.n1782 585
R11058 gnd.n4174 gnd.n1782 585
R11059 gnd.n4582 gnd.n1781 585
R11060 gnd.n2127 gnd.n1781 585
R11061 gnd.n4583 gnd.n1780 585
R11062 gnd.n4166 gnd.n1780 585
R11063 gnd.n2137 gnd.n1778 585
R11064 gnd.n2138 gnd.n2137 585
R11065 gnd.n4587 gnd.n1777 585
R11066 gnd.n4158 gnd.n1777 585
R11067 gnd.n4588 gnd.n1776 585
R11068 gnd.n3945 gnd.n1776 585
R11069 gnd.n4589 gnd.n1775 585
R11070 gnd.n4019 gnd.n1775 585
R11071 gnd.n2226 gnd.n1773 585
R11072 gnd.n2227 gnd.n2226 585
R11073 gnd.n4593 gnd.n1772 585
R11074 gnd.n4011 gnd.n1772 585
R11075 gnd.n4594 gnd.n1771 585
R11076 gnd.n2231 gnd.n1771 585
R11077 gnd.n4595 gnd.n1770 585
R11078 gnd.n2237 gnd.n1770 585
R11079 gnd.n2245 gnd.n1768 585
R11080 gnd.n3984 gnd.n2245 585
R11081 gnd.n4599 gnd.n1767 585
R11082 gnd.n2241 gnd.n1767 585
R11083 gnd.n4600 gnd.n1766 585
R11084 gnd.n3974 gnd.n1766 585
R11085 gnd.n4601 gnd.n1765 585
R11086 gnd.n3966 gnd.n1765 585
R11087 gnd.n3853 gnd.n1763 585
R11088 gnd.n3854 gnd.n3853 585
R11089 gnd.n4605 gnd.n1762 585
R11090 gnd.n3932 gnd.n1762 585
R11091 gnd.n4606 gnd.n1761 585
R11092 gnd.n2276 gnd.n1761 585
R11093 gnd.n4607 gnd.n1760 585
R11094 gnd.n3922 gnd.n1760 585
R11095 gnd.n3908 gnd.n1758 585
R11096 gnd.n3909 gnd.n3908 585
R11097 gnd.n4611 gnd.n1757 585
R11098 gnd.n3879 gnd.n1757 585
R11099 gnd.n4612 gnd.n1756 585
R11100 gnd.n3899 gnd.n1756 585
R11101 gnd.n4613 gnd.n1755 585
R11102 gnd.n2299 gnd.n1755 585
R11103 gnd.n3888 gnd.n1753 585
R11104 gnd.n3889 gnd.n3888 585
R11105 gnd.n4617 gnd.n1752 585
R11106 gnd.n2308 gnd.n1752 585
R11107 gnd.n4618 gnd.n1751 585
R11108 gnd.n3836 gnd.n1751 585
R11109 gnd.n4619 gnd.n1750 585
R11110 gnd.n2324 gnd.n1750 585
R11111 gnd.n3827 gnd.n1748 585
R11112 gnd.n3828 gnd.n3827 585
R11113 gnd.n4623 gnd.n1747 585
R11114 gnd.n2328 gnd.n1747 585
R11115 gnd.n4624 gnd.n1746 585
R11116 gnd.n2335 gnd.n1746 585
R11117 gnd.n4625 gnd.n1745 585
R11118 gnd.n3801 gnd.n1745 585
R11119 gnd.n3755 gnd.n1743 585
R11120 gnd.n3756 gnd.n3755 585
R11121 gnd.n4629 gnd.n1742 585
R11122 gnd.n3791 gnd.n1742 585
R11123 gnd.n4630 gnd.n1741 585
R11124 gnd.n3783 gnd.n1741 585
R11125 gnd.n4631 gnd.n1740 585
R11126 gnd.n2366 gnd.n1740 585
R11127 gnd.n2364 gnd.n1738 585
R11128 gnd.n3749 gnd.n2364 585
R11129 gnd.n4635 gnd.n1737 585
R11130 gnd.n2374 gnd.n1737 585
R11131 gnd.n4636 gnd.n1736 585
R11132 gnd.n3739 gnd.n1736 585
R11133 gnd.n4637 gnd.n1735 585
R11134 gnd.n3726 gnd.n1735 585
R11135 gnd.n3672 gnd.n1733 585
R11136 gnd.n3673 gnd.n3672 585
R11137 gnd.n4641 gnd.n1732 585
R11138 gnd.n2385 gnd.n1732 585
R11139 gnd.n4642 gnd.n1731 585
R11140 gnd.n2389 gnd.n1731 585
R11141 gnd.n4643 gnd.n1730 585
R11142 gnd.n2395 gnd.n1730 585
R11143 gnd.n2402 gnd.n1728 585
R11144 gnd.n3681 gnd.n2402 585
R11145 gnd.n4647 gnd.n1727 585
R11146 gnd.n2399 gnd.n1727 585
R11147 gnd.n4648 gnd.n1726 585
R11148 gnd.n3653 gnd.n1726 585
R11149 gnd.n4649 gnd.n1725 585
R11150 gnd.n2435 gnd.n1725 585
R11151 gnd.n3643 gnd.n1723 585
R11152 gnd.n3644 gnd.n3643 585
R11153 gnd.n4653 gnd.n1722 585
R11154 gnd.n3623 gnd.n1722 585
R11155 gnd.n4654 gnd.n1721 585
R11156 gnd.n2466 gnd.n1721 585
R11157 gnd.n4655 gnd.n1720 585
R11158 gnd.n3614 gnd.n1720 585
R11159 gnd.n3586 gnd.n1718 585
R11160 gnd.n3587 gnd.n3586 585
R11161 gnd.n4659 gnd.n1717 585
R11162 gnd.n3604 gnd.n1717 585
R11163 gnd.n4660 gnd.n1716 585
R11164 gnd.n2470 gnd.n1716 585
R11165 gnd.n4661 gnd.n1715 585
R11166 gnd.n3573 gnd.n1715 585
R11167 gnd.n2474 gnd.n1713 585
R11168 gnd.n2475 gnd.n2474 585
R11169 gnd.n4665 gnd.n1712 585
R11170 gnd.n3565 gnd.n1712 585
R11171 gnd.n4666 gnd.n1711 585
R11172 gnd.n3557 gnd.n1711 585
R11173 gnd.n4667 gnd.n1710 585
R11174 gnd.n3492 gnd.n1710 585
R11175 gnd.n2499 gnd.n1708 585
R11176 gnd.n3538 gnd.n2499 585
R11177 gnd.n4671 gnd.n1707 585
R11178 gnd.n3508 gnd.n1707 585
R11179 gnd.n4672 gnd.n1706 585
R11180 gnd.n3528 gnd.n1706 585
R11181 gnd.n4673 gnd.n1705 585
R11182 gnd.n2514 gnd.n1705 585
R11183 gnd.n1702 gnd.n1700 585
R11184 gnd.n2520 gnd.n1700 585
R11185 gnd.n4678 gnd.n4677 585
R11186 gnd.n4679 gnd.n4678 585
R11187 gnd.n1701 gnd.n1699 585
R11188 gnd.n3404 gnd.n1699 585
R11189 gnd.n3349 gnd.n1688 585
R11190 gnd.n4685 gnd.n1688 585
R11191 gnd.n3350 gnd.n3348 585
R11192 gnd.n3348 gnd.n1684 585
R11193 gnd.n3347 gnd.n3345 585
R11194 gnd.n3347 gnd.n1658 585
R11195 gnd.n3354 gnd.n3344 585
R11196 gnd.n3344 gnd.n1626 585
R11197 gnd.n3355 gnd.n3343 585
R11198 gnd.n3343 gnd.n2534 585
R11199 gnd.n3356 gnd.n2535 585
R11200 gnd.n3379 gnd.n2535 585
R11201 gnd.n2547 gnd.n2545 585
R11202 gnd.n2545 gnd.n2533 585
R11203 gnd.n3361 gnd.n3360 585
R11204 gnd.n3362 gnd.n3361 585
R11205 gnd.n2546 gnd.n2544 585
R11206 gnd.n2544 gnd.n2542 585
R11207 gnd.n3339 gnd.n3338 585
R11208 gnd.n3338 gnd.n3337 585
R11209 gnd.n2550 gnd.n2549 585
R11210 gnd.n2551 gnd.n2550 585
R11211 gnd.n4510 gnd.n1852 585
R11212 gnd.n4511 gnd.n1851 585
R11213 gnd.n2096 gnd.n1845 585
R11214 gnd.n4518 gnd.n1844 585
R11215 gnd.n4519 gnd.n1843 585
R11216 gnd.n2093 gnd.n1837 585
R11217 gnd.n4526 gnd.n1836 585
R11218 gnd.n4527 gnd.n1835 585
R11219 gnd.n2091 gnd.n1829 585
R11220 gnd.n4534 gnd.n1828 585
R11221 gnd.n4535 gnd.n1827 585
R11222 gnd.n2088 gnd.n1821 585
R11223 gnd.n4542 gnd.n1820 585
R11224 gnd.n4543 gnd.n1819 585
R11225 gnd.n2086 gnd.n1812 585
R11226 gnd.n4550 gnd.n1811 585
R11227 gnd.n4551 gnd.n1810 585
R11228 gnd.n2083 gnd.n1807 585
R11229 gnd.n4556 gnd.n1806 585
R11230 gnd.n4557 gnd.n1805 585
R11231 gnd.n4558 gnd.n1804 585
R11232 gnd.n2080 gnd.n1802 585
R11233 gnd.n4562 gnd.n1801 585
R11234 gnd.n4563 gnd.n1800 585
R11235 gnd.n4564 gnd.n1796 585
R11236 gnd.n4254 gnd.n1791 585
R11237 gnd.n4251 gnd.n1791 585
R11238 gnd.n4255 gnd.n4253 585
R11239 gnd.n2078 gnd.n2077 585
R11240 gnd.n2099 gnd.n2098 585
R11241 gnd.n4151 gnd.n2140 482.89
R11242 gnd.n4034 gnd.n4033 482.89
R11243 gnd.n3473 gnd.n3471 482.89
R11244 gnd.n4754 gnd.n1661 482.89
R11245 gnd.n3407 gnd.t348 443.966
R11246 gnd.n2188 gnd.t374 443.966
R11247 gnd.n4691 gnd.t399 443.966
R11248 gnd.n2182 gnd.t303 443.966
R11249 gnd.n6745 gnd.n6744 414.56
R11250 gnd.n3118 gnd.t338 371.625
R11251 gnd.n4504 gnd.t371 371.625
R11252 gnd.n2577 gnd.t383 371.625
R11253 gnd.n1925 gnd.t364 371.625
R11254 gnd.n1948 gnd.t355 371.625
R11255 gnd.n4384 gnd.t292 371.625
R11256 gnd.n346 gnd.t389 371.625
R11257 gnd.n326 gnd.t307 371.625
R11258 gnd.n7628 gnd.t325 371.625
R11259 gnd.n366 gnd.t345 371.625
R11260 gnd.n1208 gnd.t358 371.625
R11261 gnd.n1230 gnd.t296 371.625
R11262 gnd.n1252 gnd.t315 371.625
R11263 gnd.n2746 gnd.t386 371.625
R11264 gnd.n1609 gnd.t380 371.625
R11265 gnd.n3177 gnd.t311 371.625
R11266 gnd.n3190 gnd.t335 371.625
R11267 gnd.n1853 gnd.t318 371.625
R11268 gnd.n5708 gnd.t331 323.425
R11269 gnd.n1129 gnd.t367 323.425
R11270 gnd.n6383 gnd.n6357 289.615
R11271 gnd.n6351 gnd.n6325 289.615
R11272 gnd.n6319 gnd.n6293 289.615
R11273 gnd.n6288 gnd.n6262 289.615
R11274 gnd.n6256 gnd.n6230 289.615
R11275 gnd.n6224 gnd.n6198 289.615
R11276 gnd.n6192 gnd.n6166 289.615
R11277 gnd.n6161 gnd.n6135 289.615
R11278 gnd.n5558 gnd.t285 279.217
R11279 gnd.n6494 gnd.t392 279.217
R11280 gnd.n1668 gnd.t379 260.649
R11281 gnd.n2153 gnd.t302 260.649
R11282 gnd.n4756 gnd.n4755 256.663
R11283 gnd.n4756 gnd.n1627 256.663
R11284 gnd.n4756 gnd.n1628 256.663
R11285 gnd.n4756 gnd.n1629 256.663
R11286 gnd.n4756 gnd.n1630 256.663
R11287 gnd.n4756 gnd.n1631 256.663
R11288 gnd.n4756 gnd.n1632 256.663
R11289 gnd.n4756 gnd.n1633 256.663
R11290 gnd.n4756 gnd.n1634 256.663
R11291 gnd.n4756 gnd.n1635 256.663
R11292 gnd.n4756 gnd.n1636 256.663
R11293 gnd.n4756 gnd.n1637 256.663
R11294 gnd.n4756 gnd.n1638 256.663
R11295 gnd.n4756 gnd.n1639 256.663
R11296 gnd.n4756 gnd.n1640 256.663
R11297 gnd.n4756 gnd.n1641 256.663
R11298 gnd.n4759 gnd.n1624 256.663
R11299 gnd.n4757 gnd.n4756 256.663
R11300 gnd.n4756 gnd.n1642 256.663
R11301 gnd.n4756 gnd.n1643 256.663
R11302 gnd.n4756 gnd.n1644 256.663
R11303 gnd.n4756 gnd.n1645 256.663
R11304 gnd.n4756 gnd.n1646 256.663
R11305 gnd.n4756 gnd.n1647 256.663
R11306 gnd.n4756 gnd.n1648 256.663
R11307 gnd.n4756 gnd.n1649 256.663
R11308 gnd.n4756 gnd.n1650 256.663
R11309 gnd.n4756 gnd.n1651 256.663
R11310 gnd.n4756 gnd.n1652 256.663
R11311 gnd.n4756 gnd.n1653 256.663
R11312 gnd.n4756 gnd.n1654 256.663
R11313 gnd.n4756 gnd.n1655 256.663
R11314 gnd.n4756 gnd.n1656 256.663
R11315 gnd.n4756 gnd.n1657 256.663
R11316 gnd.n4032 gnd.n2128 256.663
R11317 gnd.n4039 gnd.n2128 256.663
R11318 gnd.n2209 gnd.n2128 256.663
R11319 gnd.n4046 gnd.n2128 256.663
R11320 gnd.n2206 gnd.n2128 256.663
R11321 gnd.n4053 gnd.n2128 256.663
R11322 gnd.n2203 gnd.n2128 256.663
R11323 gnd.n4060 gnd.n2128 256.663
R11324 gnd.n2200 gnd.n2128 256.663
R11325 gnd.n4067 gnd.n2128 256.663
R11326 gnd.n2197 gnd.n2128 256.663
R11327 gnd.n4074 gnd.n2128 256.663
R11328 gnd.n2194 gnd.n2128 256.663
R11329 gnd.n4081 gnd.n2128 256.663
R11330 gnd.n2191 gnd.n2128 256.663
R11331 gnd.n4089 gnd.n2128 256.663
R11332 gnd.n4092 gnd.n1935 256.663
R11333 gnd.n4093 gnd.n2128 256.663
R11334 gnd.n4097 gnd.n2128 256.663
R11335 gnd.n2185 gnd.n2128 256.663
R11336 gnd.n4105 gnd.n2128 256.663
R11337 gnd.n2180 gnd.n2128 256.663
R11338 gnd.n4112 gnd.n2128 256.663
R11339 gnd.n2177 gnd.n2128 256.663
R11340 gnd.n4119 gnd.n2128 256.663
R11341 gnd.n2174 gnd.n2128 256.663
R11342 gnd.n4126 gnd.n2128 256.663
R11343 gnd.n2171 gnd.n2128 256.663
R11344 gnd.n4133 gnd.n2128 256.663
R11345 gnd.n2168 gnd.n2128 256.663
R11346 gnd.n4140 gnd.n2128 256.663
R11347 gnd.n2165 gnd.n2128 256.663
R11348 gnd.n4147 gnd.n2128 256.663
R11349 gnd.n4150 gnd.n2128 256.663
R11350 gnd.n5111 gnd.n1176 242.672
R11351 gnd.n5111 gnd.n1177 242.672
R11352 gnd.n5111 gnd.n1178 242.672
R11353 gnd.n5111 gnd.n1179 242.672
R11354 gnd.n5111 gnd.n1180 242.672
R11355 gnd.n5111 gnd.n1181 242.672
R11356 gnd.n5111 gnd.n1182 242.672
R11357 gnd.n5111 gnd.n1183 242.672
R11358 gnd.n5111 gnd.n1184 242.672
R11359 gnd.n4810 gnd.n1562 242.672
R11360 gnd.n4810 gnd.n1561 242.672
R11361 gnd.n4810 gnd.n1560 242.672
R11362 gnd.n4810 gnd.n1559 242.672
R11363 gnd.n4810 gnd.n1558 242.672
R11364 gnd.n4810 gnd.n1557 242.672
R11365 gnd.n4810 gnd.n1556 242.672
R11366 gnd.n4810 gnd.n1555 242.672
R11367 gnd.n4810 gnd.n1554 242.672
R11368 gnd.n5613 gnd.n5522 242.672
R11369 gnd.n5526 gnd.n5522 242.672
R11370 gnd.n5606 gnd.n5522 242.672
R11371 gnd.n5600 gnd.n5522 242.672
R11372 gnd.n5598 gnd.n5522 242.672
R11373 gnd.n5592 gnd.n5522 242.672
R11374 gnd.n5590 gnd.n5522 242.672
R11375 gnd.n5584 gnd.n5522 242.672
R11376 gnd.n5582 gnd.n5522 242.672
R11377 gnd.n5576 gnd.n5522 242.672
R11378 gnd.n5574 gnd.n5522 242.672
R11379 gnd.n5567 gnd.n5522 242.672
R11380 gnd.n5565 gnd.n5522 242.672
R11381 gnd.n6559 gnd.n1147 242.672
R11382 gnd.n6559 gnd.n1146 242.672
R11383 gnd.n6559 gnd.n1145 242.672
R11384 gnd.n6559 gnd.n1144 242.672
R11385 gnd.n6559 gnd.n1143 242.672
R11386 gnd.n6559 gnd.n1142 242.672
R11387 gnd.n6559 gnd.n1141 242.672
R11388 gnd.n6559 gnd.n1140 242.672
R11389 gnd.n6559 gnd.n1139 242.672
R11390 gnd.n6559 gnd.n1138 242.672
R11391 gnd.n6559 gnd.n1137 242.672
R11392 gnd.n6559 gnd.n1136 242.672
R11393 gnd.n6559 gnd.n1135 242.672
R11394 gnd.n4501 gnd.n1890 242.672
R11395 gnd.n4501 gnd.n1892 242.672
R11396 gnd.n4501 gnd.n1893 242.672
R11397 gnd.n4501 gnd.n1895 242.672
R11398 gnd.n4501 gnd.n1897 242.672
R11399 gnd.n4501 gnd.n1898 242.672
R11400 gnd.n4501 gnd.n1900 242.672
R11401 gnd.n4501 gnd.n1902 242.672
R11402 gnd.n4502 gnd.n4501 242.672
R11403 gnd.n7663 gnd.n260 242.672
R11404 gnd.n7663 gnd.n259 242.672
R11405 gnd.n7663 gnd.n258 242.672
R11406 gnd.n7663 gnd.n257 242.672
R11407 gnd.n7663 gnd.n256 242.672
R11408 gnd.n7663 gnd.n255 242.672
R11409 gnd.n7663 gnd.n254 242.672
R11410 gnd.n7663 gnd.n253 242.672
R11411 gnd.n7663 gnd.n252 242.672
R11412 gnd.n5742 gnd.n5741 242.672
R11413 gnd.n5742 gnd.n5683 242.672
R11414 gnd.n5742 gnd.n5684 242.672
R11415 gnd.n5742 gnd.n5685 242.672
R11416 gnd.n5742 gnd.n5686 242.672
R11417 gnd.n5742 gnd.n5687 242.672
R11418 gnd.n5742 gnd.n5688 242.672
R11419 gnd.n5742 gnd.n5689 242.672
R11420 gnd.n6559 gnd.n1128 242.672
R11421 gnd.n6560 gnd.n6559 242.672
R11422 gnd.n6559 gnd.n5112 242.672
R11423 gnd.n6559 gnd.n5113 242.672
R11424 gnd.n6559 gnd.n5114 242.672
R11425 gnd.n6559 gnd.n5115 242.672
R11426 gnd.n6559 gnd.n5116 242.672
R11427 gnd.n6559 gnd.n5117 242.672
R11428 gnd.n5111 gnd.n5110 242.672
R11429 gnd.n5111 gnd.n1148 242.672
R11430 gnd.n5111 gnd.n1149 242.672
R11431 gnd.n5111 gnd.n1150 242.672
R11432 gnd.n5111 gnd.n1151 242.672
R11433 gnd.n5111 gnd.n1152 242.672
R11434 gnd.n5111 gnd.n1153 242.672
R11435 gnd.n5111 gnd.n1154 242.672
R11436 gnd.n5111 gnd.n1155 242.672
R11437 gnd.n5111 gnd.n1156 242.672
R11438 gnd.n5111 gnd.n1157 242.672
R11439 gnd.n5111 gnd.n1158 242.672
R11440 gnd.n5111 gnd.n1159 242.672
R11441 gnd.n5111 gnd.n1160 242.672
R11442 gnd.n5111 gnd.n1161 242.672
R11443 gnd.n5111 gnd.n1162 242.672
R11444 gnd.n5111 gnd.n1163 242.672
R11445 gnd.n5111 gnd.n1164 242.672
R11446 gnd.n5111 gnd.n1165 242.672
R11447 gnd.n5111 gnd.n1166 242.672
R11448 gnd.n5111 gnd.n1167 242.672
R11449 gnd.n5111 gnd.n1168 242.672
R11450 gnd.n5111 gnd.n1169 242.672
R11451 gnd.n5111 gnd.n1170 242.672
R11452 gnd.n5111 gnd.n1171 242.672
R11453 gnd.n5111 gnd.n1172 242.672
R11454 gnd.n5111 gnd.n1173 242.672
R11455 gnd.n5111 gnd.n1174 242.672
R11456 gnd.n5111 gnd.n1175 242.672
R11457 gnd.n4810 gnd.n1564 242.672
R11458 gnd.n4810 gnd.n1565 242.672
R11459 gnd.n4810 gnd.n1566 242.672
R11460 gnd.n4810 gnd.n1567 242.672
R11461 gnd.n4810 gnd.n1568 242.672
R11462 gnd.n4810 gnd.n1569 242.672
R11463 gnd.n4810 gnd.n1570 242.672
R11464 gnd.n4810 gnd.n1571 242.672
R11465 gnd.n4810 gnd.n1572 242.672
R11466 gnd.n4810 gnd.n1573 242.672
R11467 gnd.n4810 gnd.n1574 242.672
R11468 gnd.n4810 gnd.n1575 242.672
R11469 gnd.n4810 gnd.n1576 242.672
R11470 gnd.n4810 gnd.n1577 242.672
R11471 gnd.n4810 gnd.n1578 242.672
R11472 gnd.n4810 gnd.n1579 242.672
R11473 gnd.n4760 gnd.n1620 242.672
R11474 gnd.n4810 gnd.n1580 242.672
R11475 gnd.n4810 gnd.n1581 242.672
R11476 gnd.n4810 gnd.n1582 242.672
R11477 gnd.n4810 gnd.n1583 242.672
R11478 gnd.n4810 gnd.n1584 242.672
R11479 gnd.n4810 gnd.n1585 242.672
R11480 gnd.n4810 gnd.n1586 242.672
R11481 gnd.n4810 gnd.n1587 242.672
R11482 gnd.n4810 gnd.n1588 242.672
R11483 gnd.n4810 gnd.n1589 242.672
R11484 gnd.n4810 gnd.n1590 242.672
R11485 gnd.n4810 gnd.n1591 242.672
R11486 gnd.n4810 gnd.n4809 242.672
R11487 gnd.n4501 gnd.n4500 242.672
R11488 gnd.n4501 gnd.n1862 242.672
R11489 gnd.n4501 gnd.n1863 242.672
R11490 gnd.n4501 gnd.n1864 242.672
R11491 gnd.n4501 gnd.n1865 242.672
R11492 gnd.n4501 gnd.n1866 242.672
R11493 gnd.n4501 gnd.n1867 242.672
R11494 gnd.n4501 gnd.n1868 242.672
R11495 gnd.n4501 gnd.n1869 242.672
R11496 gnd.n4501 gnd.n1870 242.672
R11497 gnd.n4501 gnd.n1871 242.672
R11498 gnd.n4501 gnd.n1872 242.672
R11499 gnd.n4501 gnd.n1873 242.672
R11500 gnd.n4448 gnd.n1936 242.672
R11501 gnd.n4501 gnd.n1874 242.672
R11502 gnd.n4501 gnd.n1875 242.672
R11503 gnd.n4501 gnd.n1876 242.672
R11504 gnd.n4501 gnd.n1877 242.672
R11505 gnd.n4501 gnd.n1878 242.672
R11506 gnd.n4501 gnd.n1879 242.672
R11507 gnd.n4501 gnd.n1880 242.672
R11508 gnd.n4501 gnd.n1881 242.672
R11509 gnd.n4501 gnd.n1882 242.672
R11510 gnd.n4501 gnd.n1883 242.672
R11511 gnd.n4501 gnd.n1884 242.672
R11512 gnd.n4501 gnd.n1885 242.672
R11513 gnd.n4501 gnd.n1886 242.672
R11514 gnd.n4501 gnd.n1887 242.672
R11515 gnd.n4501 gnd.n1888 242.672
R11516 gnd.n4501 gnd.n1889 242.672
R11517 gnd.n7663 gnd.n261 242.672
R11518 gnd.n7663 gnd.n262 242.672
R11519 gnd.n7663 gnd.n263 242.672
R11520 gnd.n7663 gnd.n264 242.672
R11521 gnd.n7663 gnd.n265 242.672
R11522 gnd.n7663 gnd.n266 242.672
R11523 gnd.n7663 gnd.n267 242.672
R11524 gnd.n7663 gnd.n268 242.672
R11525 gnd.n7663 gnd.n269 242.672
R11526 gnd.n7663 gnd.n270 242.672
R11527 gnd.n7663 gnd.n271 242.672
R11528 gnd.n7663 gnd.n272 242.672
R11529 gnd.n7663 gnd.n273 242.672
R11530 gnd.n7663 gnd.n274 242.672
R11531 gnd.n7663 gnd.n275 242.672
R11532 gnd.n7663 gnd.n276 242.672
R11533 gnd.n7663 gnd.n277 242.672
R11534 gnd.n7663 gnd.n278 242.672
R11535 gnd.n7663 gnd.n279 242.672
R11536 gnd.n7663 gnd.n280 242.672
R11537 gnd.n7663 gnd.n281 242.672
R11538 gnd.n7663 gnd.n282 242.672
R11539 gnd.n7663 gnd.n283 242.672
R11540 gnd.n7663 gnd.n284 242.672
R11541 gnd.n7663 gnd.n285 242.672
R11542 gnd.n7663 gnd.n286 242.672
R11543 gnd.n7663 gnd.n287 242.672
R11544 gnd.n7663 gnd.n288 242.672
R11545 gnd.n7663 gnd.n7662 242.672
R11546 gnd.n3328 gnd.n2559 242.672
R11547 gnd.n3328 gnd.n2560 242.672
R11548 gnd.n3328 gnd.n2561 242.672
R11549 gnd.n3328 gnd.n2562 242.672
R11550 gnd.n3328 gnd.n2563 242.672
R11551 gnd.n3328 gnd.n2564 242.672
R11552 gnd.n3328 gnd.n2565 242.672
R11553 gnd.n3328 gnd.n2566 242.672
R11554 gnd.n3328 gnd.n2567 242.672
R11555 gnd.n3328 gnd.n2568 242.672
R11556 gnd.n3328 gnd.n2569 242.672
R11557 gnd.n3328 gnd.n2570 242.672
R11558 gnd.n3328 gnd.n2571 242.672
R11559 gnd.n3328 gnd.n2572 242.672
R11560 gnd.n4251 gnd.n2100 242.672
R11561 gnd.n4251 gnd.n2097 242.672
R11562 gnd.n4251 gnd.n2095 242.672
R11563 gnd.n4251 gnd.n2094 242.672
R11564 gnd.n4251 gnd.n2092 242.672
R11565 gnd.n4251 gnd.n2090 242.672
R11566 gnd.n4251 gnd.n2089 242.672
R11567 gnd.n4251 gnd.n2087 242.672
R11568 gnd.n4251 gnd.n2085 242.672
R11569 gnd.n4251 gnd.n2084 242.672
R11570 gnd.n4251 gnd.n2082 242.672
R11571 gnd.n4251 gnd.n2081 242.672
R11572 gnd.n4251 gnd.n2079 242.672
R11573 gnd.n4252 gnd.n4251 242.672
R11574 gnd.n7664 gnd.n250 240.244
R11575 gnd.n7661 gnd.n289 240.244
R11576 gnd.n7657 gnd.n7656 240.244
R11577 gnd.n7653 gnd.n7652 240.244
R11578 gnd.n7649 gnd.n7648 240.244
R11579 gnd.n7645 gnd.n7644 240.244
R11580 gnd.n7641 gnd.n7640 240.244
R11581 gnd.n7637 gnd.n7636 240.244
R11582 gnd.n7633 gnd.n7632 240.244
R11583 gnd.n7626 gnd.n7625 240.244
R11584 gnd.n7622 gnd.n7621 240.244
R11585 gnd.n7618 gnd.n7617 240.244
R11586 gnd.n7614 gnd.n7613 240.244
R11587 gnd.n7610 gnd.n7609 240.244
R11588 gnd.n7606 gnd.n7605 240.244
R11589 gnd.n7602 gnd.n7601 240.244
R11590 gnd.n7598 gnd.n7597 240.244
R11591 gnd.n7594 gnd.n7593 240.244
R11592 gnd.n7590 gnd.n7589 240.244
R11593 gnd.n7583 gnd.n7582 240.244
R11594 gnd.n7580 gnd.n7579 240.244
R11595 gnd.n7576 gnd.n7575 240.244
R11596 gnd.n7572 gnd.n7571 240.244
R11597 gnd.n7568 gnd.n7567 240.244
R11598 gnd.n7564 gnd.n7563 240.244
R11599 gnd.n7560 gnd.n7559 240.244
R11600 gnd.n7556 gnd.n7555 240.244
R11601 gnd.n7552 gnd.n7551 240.244
R11602 gnd.n7548 gnd.n7547 240.244
R11603 gnd.n4381 gnd.n1969 240.244
R11604 gnd.n4373 gnd.n1969 240.244
R11605 gnd.n4373 gnd.n1980 240.244
R11606 gnd.n1996 gnd.n1980 240.244
R11607 gnd.n4271 gnd.n1996 240.244
R11608 gnd.n4271 gnd.n2009 240.244
R11609 gnd.n4276 gnd.n2009 240.244
R11610 gnd.n4276 gnd.n2020 240.244
R11611 gnd.n4286 gnd.n2020 240.244
R11612 gnd.n4286 gnd.n2030 240.244
R11613 gnd.n4299 gnd.n2030 240.244
R11614 gnd.n4299 gnd.n2041 240.244
R11615 gnd.n2061 gnd.n2041 240.244
R11616 gnd.n2061 gnd.n2050 240.244
R11617 gnd.n2053 gnd.n2050 240.244
R11618 gnd.n4292 gnd.n2053 240.244
R11619 gnd.n4292 gnd.n566 240.244
R11620 gnd.n7371 gnd.n566 240.244
R11621 gnd.n7371 gnd.n556 240.244
R11622 gnd.n556 gnd.n547 240.244
R11623 gnd.n7403 gnd.n547 240.244
R11624 gnd.n7403 gnd.n537 240.244
R11625 gnd.n7407 gnd.n537 240.244
R11626 gnd.n7407 gnd.n527 240.244
R11627 gnd.n527 gnd.n519 240.244
R11628 gnd.n7439 gnd.n519 240.244
R11629 gnd.n7439 gnd.n510 240.244
R11630 gnd.n510 gnd.n505 240.244
R11631 gnd.n7445 gnd.n505 240.244
R11632 gnd.n7445 gnd.n497 240.244
R11633 gnd.n497 gnd.n491 240.244
R11634 gnd.n491 gnd.n486 240.244
R11635 gnd.n7481 gnd.n486 240.244
R11636 gnd.n7481 gnd.n101 240.244
R11637 gnd.n7490 gnd.n101 240.244
R11638 gnd.n7491 gnd.n7490 240.244
R11639 gnd.n7491 gnd.n118 240.244
R11640 gnd.n7494 gnd.n118 240.244
R11641 gnd.n7494 gnd.n129 240.244
R11642 gnd.n7498 gnd.n129 240.244
R11643 gnd.n7498 gnd.n138 240.244
R11644 gnd.n7501 gnd.n138 240.244
R11645 gnd.n7501 gnd.n147 240.244
R11646 gnd.n7505 gnd.n147 240.244
R11647 gnd.n7505 gnd.n157 240.244
R11648 gnd.n7508 gnd.n157 240.244
R11649 gnd.n7508 gnd.n166 240.244
R11650 gnd.n7512 gnd.n166 240.244
R11651 gnd.n7512 gnd.n176 240.244
R11652 gnd.n7515 gnd.n176 240.244
R11653 gnd.n7515 gnd.n185 240.244
R11654 gnd.n7519 gnd.n185 240.244
R11655 gnd.n7519 gnd.n195 240.244
R11656 gnd.n7522 gnd.n195 240.244
R11657 gnd.n7522 gnd.n204 240.244
R11658 gnd.n7526 gnd.n204 240.244
R11659 gnd.n7526 gnd.n214 240.244
R11660 gnd.n7529 gnd.n214 240.244
R11661 gnd.n7529 gnd.n223 240.244
R11662 gnd.n7533 gnd.n223 240.244
R11663 gnd.n7533 gnd.n233 240.244
R11664 gnd.n7536 gnd.n233 240.244
R11665 gnd.n7536 gnd.n242 240.244
R11666 gnd.n7540 gnd.n242 240.244
R11667 gnd.n1905 gnd.n1904 240.244
R11668 gnd.n4494 gnd.n1904 240.244
R11669 gnd.n4492 gnd.n4491 240.244
R11670 gnd.n4488 gnd.n4487 240.244
R11671 gnd.n4484 gnd.n4483 240.244
R11672 gnd.n4480 gnd.n4479 240.244
R11673 gnd.n4476 gnd.n4475 240.244
R11674 gnd.n4472 gnd.n4471 240.244
R11675 gnd.n4468 gnd.n4467 240.244
R11676 gnd.n4463 gnd.n4462 240.244
R11677 gnd.n4459 gnd.n4458 240.244
R11678 gnd.n4455 gnd.n4454 240.244
R11679 gnd.n4451 gnd.n4450 240.244
R11680 gnd.n4446 gnd.n4445 240.244
R11681 gnd.n4442 gnd.n4441 240.244
R11682 gnd.n4438 gnd.n4437 240.244
R11683 gnd.n4434 gnd.n4433 240.244
R11684 gnd.n4430 gnd.n4429 240.244
R11685 gnd.n4426 gnd.n4425 240.244
R11686 gnd.n4422 gnd.n4421 240.244
R11687 gnd.n4418 gnd.n4417 240.244
R11688 gnd.n4414 gnd.n4413 240.244
R11689 gnd.n4410 gnd.n4409 240.244
R11690 gnd.n4406 gnd.n4405 240.244
R11691 gnd.n4402 gnd.n4401 240.244
R11692 gnd.n4398 gnd.n4397 240.244
R11693 gnd.n4394 gnd.n4393 240.244
R11694 gnd.n4390 gnd.n4389 240.244
R11695 gnd.n1984 gnd.n1906 240.244
R11696 gnd.n4371 gnd.n1984 240.244
R11697 gnd.n4371 gnd.n1985 240.244
R11698 gnd.n4367 gnd.n1985 240.244
R11699 gnd.n4367 gnd.n1994 240.244
R11700 gnd.n4359 gnd.n1994 240.244
R11701 gnd.n4359 gnd.n2012 240.244
R11702 gnd.n4355 gnd.n2012 240.244
R11703 gnd.n4355 gnd.n2018 240.244
R11704 gnd.n4347 gnd.n2018 240.244
R11705 gnd.n4347 gnd.n2033 240.244
R11706 gnd.n4343 gnd.n2033 240.244
R11707 gnd.n4343 gnd.n2039 240.244
R11708 gnd.n4335 gnd.n2039 240.244
R11709 gnd.n4335 gnd.n4329 240.244
R11710 gnd.n4329 gnd.n564 240.244
R11711 gnd.n7384 gnd.n564 240.244
R11712 gnd.n7384 gnd.n559 240.244
R11713 gnd.n7392 gnd.n559 240.244
R11714 gnd.n7392 gnd.n560 240.244
R11715 gnd.n560 gnd.n535 240.244
R11716 gnd.n7420 gnd.n535 240.244
R11717 gnd.n7420 gnd.n530 240.244
R11718 gnd.n7429 gnd.n530 240.244
R11719 gnd.n7429 gnd.n531 240.244
R11720 gnd.n531 gnd.n507 240.244
R11721 gnd.n7453 gnd.n507 240.244
R11722 gnd.n7456 gnd.n7453 240.244
R11723 gnd.n7456 gnd.n495 240.244
R11724 gnd.n7466 gnd.n495 240.244
R11725 gnd.n7472 gnd.n7466 240.244
R11726 gnd.n7472 gnd.n7469 240.244
R11727 gnd.n7469 gnd.n104 240.244
R11728 gnd.n7756 gnd.n104 240.244
R11729 gnd.n7756 gnd.n105 240.244
R11730 gnd.n115 gnd.n105 240.244
R11731 gnd.n7750 gnd.n115 240.244
R11732 gnd.n7750 gnd.n116 240.244
R11733 gnd.n7742 gnd.n116 240.244
R11734 gnd.n7742 gnd.n132 240.244
R11735 gnd.n7738 gnd.n132 240.244
R11736 gnd.n7738 gnd.n137 240.244
R11737 gnd.n7730 gnd.n137 240.244
R11738 gnd.n7730 gnd.n149 240.244
R11739 gnd.n7726 gnd.n149 240.244
R11740 gnd.n7726 gnd.n155 240.244
R11741 gnd.n7718 gnd.n155 240.244
R11742 gnd.n7718 gnd.n169 240.244
R11743 gnd.n7714 gnd.n169 240.244
R11744 gnd.n7714 gnd.n175 240.244
R11745 gnd.n7706 gnd.n175 240.244
R11746 gnd.n7706 gnd.n187 240.244
R11747 gnd.n7702 gnd.n187 240.244
R11748 gnd.n7702 gnd.n193 240.244
R11749 gnd.n7694 gnd.n193 240.244
R11750 gnd.n7694 gnd.n207 240.244
R11751 gnd.n7690 gnd.n207 240.244
R11752 gnd.n7690 gnd.n213 240.244
R11753 gnd.n7682 gnd.n213 240.244
R11754 gnd.n7682 gnd.n226 240.244
R11755 gnd.n7678 gnd.n226 240.244
R11756 gnd.n7678 gnd.n232 240.244
R11757 gnd.n7670 gnd.n232 240.244
R11758 gnd.n7670 gnd.n245 240.244
R11759 gnd.n4811 gnd.n1551 240.244
R11760 gnd.n4808 gnd.n1592 240.244
R11761 gnd.n4804 gnd.n4803 240.244
R11762 gnd.n4800 gnd.n4799 240.244
R11763 gnd.n4796 gnd.n4795 240.244
R11764 gnd.n4792 gnd.n4791 240.244
R11765 gnd.n4788 gnd.n4787 240.244
R11766 gnd.n4784 gnd.n4783 240.244
R11767 gnd.n4780 gnd.n4779 240.244
R11768 gnd.n4775 gnd.n4774 240.244
R11769 gnd.n4771 gnd.n4770 240.244
R11770 gnd.n4767 gnd.n4766 240.244
R11771 gnd.n4763 gnd.n4762 240.244
R11772 gnd.n3199 gnd.n3198 240.244
R11773 gnd.n3202 gnd.n3201 240.244
R11774 gnd.n3209 gnd.n3208 240.244
R11775 gnd.n3212 gnd.n3211 240.244
R11776 gnd.n3217 gnd.n3192 240.244
R11777 gnd.n3221 gnd.n3220 240.244
R11778 gnd.n3228 gnd.n3227 240.244
R11779 gnd.n3231 gnd.n3230 240.244
R11780 gnd.n3238 gnd.n3237 240.244
R11781 gnd.n3241 gnd.n3240 240.244
R11782 gnd.n3248 gnd.n3247 240.244
R11783 gnd.n3251 gnd.n3250 240.244
R11784 gnd.n3258 gnd.n3257 240.244
R11785 gnd.n3261 gnd.n3260 240.244
R11786 gnd.n3266 gnd.n3179 240.244
R11787 gnd.n4989 gnd.n4988 240.244
R11788 gnd.n4988 gnd.n1259 240.244
R11789 gnd.n1271 gnd.n1259 240.244
R11790 gnd.n2673 gnd.n1271 240.244
R11791 gnd.n2673 gnd.n1283 240.244
R11792 gnd.n2677 gnd.n1283 240.244
R11793 gnd.n2677 gnd.n1293 240.244
R11794 gnd.n2680 gnd.n1293 240.244
R11795 gnd.n2680 gnd.n1302 240.244
R11796 gnd.n2684 gnd.n1302 240.244
R11797 gnd.n2684 gnd.n1312 240.244
R11798 gnd.n2687 gnd.n1312 240.244
R11799 gnd.n2687 gnd.n1321 240.244
R11800 gnd.n2691 gnd.n1321 240.244
R11801 gnd.n2691 gnd.n1331 240.244
R11802 gnd.n2694 gnd.n1331 240.244
R11803 gnd.n2694 gnd.n1340 240.244
R11804 gnd.n2698 gnd.n1340 240.244
R11805 gnd.n2698 gnd.n1350 240.244
R11806 gnd.n2701 gnd.n1350 240.244
R11807 gnd.n2701 gnd.n1359 240.244
R11808 gnd.n2705 gnd.n1359 240.244
R11809 gnd.n2705 gnd.n1369 240.244
R11810 gnd.n2708 gnd.n1369 240.244
R11811 gnd.n2708 gnd.n1378 240.244
R11812 gnd.n2712 gnd.n1378 240.244
R11813 gnd.n2712 gnd.n1387 240.244
R11814 gnd.n2715 gnd.n1387 240.244
R11815 gnd.n2715 gnd.n1396 240.244
R11816 gnd.n2718 gnd.n1396 240.244
R11817 gnd.n2718 gnd.n2669 240.244
R11818 gnd.n2870 gnd.n2669 240.244
R11819 gnd.n2870 gnd.n2661 240.244
R11820 gnd.n2661 gnd.n2648 240.244
R11821 gnd.n2877 gnd.n2648 240.244
R11822 gnd.n2877 gnd.n2642 240.244
R11823 gnd.n2642 gnd.n1412 240.244
R11824 gnd.n2634 gnd.n1412 240.244
R11825 gnd.n2634 gnd.n1423 240.244
R11826 gnd.n2939 gnd.n1423 240.244
R11827 gnd.n2939 gnd.n1433 240.244
R11828 gnd.n2943 gnd.n1433 240.244
R11829 gnd.n2943 gnd.n1442 240.244
R11830 gnd.n2953 gnd.n1442 240.244
R11831 gnd.n2953 gnd.n1453 240.244
R11832 gnd.n2615 gnd.n1453 240.244
R11833 gnd.n2615 gnd.n1462 240.244
R11834 gnd.n2960 gnd.n1462 240.244
R11835 gnd.n2960 gnd.n1473 240.244
R11836 gnd.n2965 gnd.n1473 240.244
R11837 gnd.n2965 gnd.n1482 240.244
R11838 gnd.n2972 gnd.n1482 240.244
R11839 gnd.n2972 gnd.n1493 240.244
R11840 gnd.n2603 gnd.n1493 240.244
R11841 gnd.n2603 gnd.n1502 240.244
R11842 gnd.n3020 gnd.n1502 240.244
R11843 gnd.n3020 gnd.n1513 240.244
R11844 gnd.n2592 gnd.n1513 240.244
R11845 gnd.n2592 gnd.n1522 240.244
R11846 gnd.n3027 gnd.n1522 240.244
R11847 gnd.n3027 gnd.n1533 240.244
R11848 gnd.n3277 gnd.n1533 240.244
R11849 gnd.n3277 gnd.n1543 240.244
R11850 gnd.n2581 gnd.n1543 240.244
R11851 gnd.n1188 gnd.n1187 240.244
R11852 gnd.n5104 gnd.n1187 240.244
R11853 gnd.n5102 gnd.n5101 240.244
R11854 gnd.n5098 gnd.n5097 240.244
R11855 gnd.n5094 gnd.n5093 240.244
R11856 gnd.n5090 gnd.n5089 240.244
R11857 gnd.n5086 gnd.n5085 240.244
R11858 gnd.n5082 gnd.n5081 240.244
R11859 gnd.n5078 gnd.n5077 240.244
R11860 gnd.n5073 gnd.n5072 240.244
R11861 gnd.n5069 gnd.n5068 240.244
R11862 gnd.n5065 gnd.n5064 240.244
R11863 gnd.n5061 gnd.n5060 240.244
R11864 gnd.n5057 gnd.n5056 240.244
R11865 gnd.n5053 gnd.n5052 240.244
R11866 gnd.n5049 gnd.n5048 240.244
R11867 gnd.n5045 gnd.n5044 240.244
R11868 gnd.n5041 gnd.n5040 240.244
R11869 gnd.n5037 gnd.n5036 240.244
R11870 gnd.n5033 gnd.n5032 240.244
R11871 gnd.n5029 gnd.n5028 240.244
R11872 gnd.n5025 gnd.n5024 240.244
R11873 gnd.n5021 gnd.n5020 240.244
R11874 gnd.n5017 gnd.n5016 240.244
R11875 gnd.n5013 gnd.n5012 240.244
R11876 gnd.n5009 gnd.n5008 240.244
R11877 gnd.n5005 gnd.n5004 240.244
R11878 gnd.n5001 gnd.n5000 240.244
R11879 gnd.n4997 gnd.n4996 240.244
R11880 gnd.n4986 gnd.n1189 240.244
R11881 gnd.n4986 gnd.n1262 240.244
R11882 gnd.n4982 gnd.n1262 240.244
R11883 gnd.n4982 gnd.n1269 240.244
R11884 gnd.n4974 gnd.n1269 240.244
R11885 gnd.n4974 gnd.n1286 240.244
R11886 gnd.n4970 gnd.n1286 240.244
R11887 gnd.n4970 gnd.n1292 240.244
R11888 gnd.n4962 gnd.n1292 240.244
R11889 gnd.n4962 gnd.n1304 240.244
R11890 gnd.n4958 gnd.n1304 240.244
R11891 gnd.n4958 gnd.n1310 240.244
R11892 gnd.n4950 gnd.n1310 240.244
R11893 gnd.n4950 gnd.n1324 240.244
R11894 gnd.n4946 gnd.n1324 240.244
R11895 gnd.n4946 gnd.n1330 240.244
R11896 gnd.n4938 gnd.n1330 240.244
R11897 gnd.n4938 gnd.n1342 240.244
R11898 gnd.n4934 gnd.n1342 240.244
R11899 gnd.n4934 gnd.n1348 240.244
R11900 gnd.n4926 gnd.n1348 240.244
R11901 gnd.n4926 gnd.n1362 240.244
R11902 gnd.n4922 gnd.n1362 240.244
R11903 gnd.n4922 gnd.n1368 240.244
R11904 gnd.n4914 gnd.n1368 240.244
R11905 gnd.n4914 gnd.n1380 240.244
R11906 gnd.n4910 gnd.n1380 240.244
R11907 gnd.n4910 gnd.n1385 240.244
R11908 gnd.n4902 gnd.n1385 240.244
R11909 gnd.n4902 gnd.n1399 240.244
R11910 gnd.n2725 gnd.n1399 240.244
R11911 gnd.n2725 gnd.n2651 240.244
R11912 gnd.n2886 gnd.n2651 240.244
R11913 gnd.n2890 gnd.n2886 240.244
R11914 gnd.n2890 gnd.n2887 240.244
R11915 gnd.n2887 gnd.n1409 240.244
R11916 gnd.n4897 gnd.n1409 240.244
R11917 gnd.n4897 gnd.n1410 240.244
R11918 gnd.n4889 gnd.n1410 240.244
R11919 gnd.n4889 gnd.n1426 240.244
R11920 gnd.n4885 gnd.n1426 240.244
R11921 gnd.n4885 gnd.n1431 240.244
R11922 gnd.n4877 gnd.n1431 240.244
R11923 gnd.n4877 gnd.n1445 240.244
R11924 gnd.n4873 gnd.n1445 240.244
R11925 gnd.n4873 gnd.n1451 240.244
R11926 gnd.n4865 gnd.n1451 240.244
R11927 gnd.n4865 gnd.n1465 240.244
R11928 gnd.n4861 gnd.n1465 240.244
R11929 gnd.n4861 gnd.n1471 240.244
R11930 gnd.n4853 gnd.n1471 240.244
R11931 gnd.n4853 gnd.n1485 240.244
R11932 gnd.n4849 gnd.n1485 240.244
R11933 gnd.n4849 gnd.n1491 240.244
R11934 gnd.n4841 gnd.n1491 240.244
R11935 gnd.n4841 gnd.n1505 240.244
R11936 gnd.n4837 gnd.n1505 240.244
R11937 gnd.n4837 gnd.n1511 240.244
R11938 gnd.n4829 gnd.n1511 240.244
R11939 gnd.n4829 gnd.n1525 240.244
R11940 gnd.n4825 gnd.n1525 240.244
R11941 gnd.n4825 gnd.n1531 240.244
R11942 gnd.n4817 gnd.n1531 240.244
R11943 gnd.n4817 gnd.n1546 240.244
R11944 gnd.n6558 gnd.n5119 240.244
R11945 gnd.n6551 gnd.n6550 240.244
R11946 gnd.n6548 gnd.n6547 240.244
R11947 gnd.n6544 gnd.n6543 240.244
R11948 gnd.n6540 gnd.n6539 240.244
R11949 gnd.n6536 gnd.n6535 240.244
R11950 gnd.n6532 gnd.n1134 240.244
R11951 gnd.n6562 gnd.n6561 240.244
R11952 gnd.n5754 gnd.n5474 240.244
R11953 gnd.n5474 gnd.n5465 240.244
R11954 gnd.n5772 gnd.n5465 240.244
R11955 gnd.n5773 gnd.n5772 240.244
R11956 gnd.n5773 gnd.n5453 240.244
R11957 gnd.n5453 gnd.n5442 240.244
R11958 gnd.n5804 gnd.n5442 240.244
R11959 gnd.n5805 gnd.n5804 240.244
R11960 gnd.n5806 gnd.n5805 240.244
R11961 gnd.n5806 gnd.n5427 240.244
R11962 gnd.n5808 gnd.n5427 240.244
R11963 gnd.n5808 gnd.n5412 240.244
R11964 gnd.n5849 gnd.n5412 240.244
R11965 gnd.n5850 gnd.n5849 240.244
R11966 gnd.n5853 gnd.n5850 240.244
R11967 gnd.n5853 gnd.n5394 240.244
R11968 gnd.n5885 gnd.n5394 240.244
R11969 gnd.n5885 gnd.n5380 240.244
R11970 gnd.n5907 gnd.n5380 240.244
R11971 gnd.n5908 gnd.n5907 240.244
R11972 gnd.n5908 gnd.n5367 240.244
R11973 gnd.n5367 gnd.n5356 240.244
R11974 gnd.n5939 gnd.n5356 240.244
R11975 gnd.n5940 gnd.n5939 240.244
R11976 gnd.n5941 gnd.n5940 240.244
R11977 gnd.n5941 gnd.n5261 240.244
R11978 gnd.n5261 gnd.n5260 240.244
R11979 gnd.n5260 gnd.n5245 240.244
R11980 gnd.n5989 gnd.n5245 240.244
R11981 gnd.n5990 gnd.n5989 240.244
R11982 gnd.n5990 gnd.n5230 240.244
R11983 gnd.n6000 gnd.n5230 240.244
R11984 gnd.n6000 gnd.n5222 240.244
R11985 gnd.n6002 gnd.n5222 240.244
R11986 gnd.n6002 gnd.n5216 240.244
R11987 gnd.n5216 gnd.n5203 240.244
R11988 gnd.n5203 gnd.n5193 240.244
R11989 gnd.n6066 gnd.n5193 240.244
R11990 gnd.n6067 gnd.n6066 240.244
R11991 gnd.n6068 gnd.n6067 240.244
R11992 gnd.n6068 gnd.n5178 240.244
R11993 gnd.n5178 gnd.n5177 240.244
R11994 gnd.n5177 gnd.n5163 240.244
R11995 gnd.n6120 gnd.n5163 240.244
R11996 gnd.n6121 gnd.n6120 240.244
R11997 gnd.n6121 gnd.n5150 240.244
R11998 gnd.n5150 gnd.n5139 240.244
R11999 gnd.n6411 gnd.n5139 240.244
R12000 gnd.n6412 gnd.n6411 240.244
R12001 gnd.n6413 gnd.n6412 240.244
R12002 gnd.n6413 gnd.n5124 240.244
R12003 gnd.n5124 gnd.n1127 240.244
R12004 gnd.n6569 gnd.n1127 240.244
R12005 gnd.n5691 gnd.n5690 240.244
R12006 gnd.n5735 gnd.n5690 240.244
R12007 gnd.n5733 gnd.n5732 240.244
R12008 gnd.n5729 gnd.n5728 240.244
R12009 gnd.n5725 gnd.n5724 240.244
R12010 gnd.n5721 gnd.n5720 240.244
R12011 gnd.n5717 gnd.n5716 240.244
R12012 gnd.n5713 gnd.n5712 240.244
R12013 gnd.n5764 gnd.n5472 240.244
R12014 gnd.n5764 gnd.n5468 240.244
R12015 gnd.n5770 gnd.n5468 240.244
R12016 gnd.n5770 gnd.n5451 240.244
R12017 gnd.n5794 gnd.n5451 240.244
R12018 gnd.n5794 gnd.n5446 240.244
R12019 gnd.n5802 gnd.n5446 240.244
R12020 gnd.n5802 gnd.n5447 240.244
R12021 gnd.n5447 gnd.n5425 240.244
R12022 gnd.n5828 gnd.n5425 240.244
R12023 gnd.n5828 gnd.n5420 240.244
R12024 gnd.n5839 gnd.n5420 240.244
R12025 gnd.n5839 gnd.n5421 240.244
R12026 gnd.n5835 gnd.n5421 240.244
R12027 gnd.n5835 gnd.n5392 240.244
R12028 gnd.n5889 gnd.n5392 240.244
R12029 gnd.n5889 gnd.n5387 240.244
R12030 gnd.n5897 gnd.n5387 240.244
R12031 gnd.n5897 gnd.n5388 240.244
R12032 gnd.n5388 gnd.n5365 240.244
R12033 gnd.n5929 gnd.n5365 240.244
R12034 gnd.n5929 gnd.n5360 240.244
R12035 gnd.n5937 gnd.n5360 240.244
R12036 gnd.n5937 gnd.n5361 240.244
R12037 gnd.n5361 gnd.n5258 240.244
R12038 gnd.n5971 gnd.n5258 240.244
R12039 gnd.n5971 gnd.n5253 240.244
R12040 gnd.n5979 gnd.n5253 240.244
R12041 gnd.n5979 gnd.n5254 240.244
R12042 gnd.n5254 gnd.n5228 240.244
R12043 gnd.n6012 gnd.n5228 240.244
R12044 gnd.n6012 gnd.n5223 240.244
R12045 gnd.n6020 gnd.n5223 240.244
R12046 gnd.n6020 gnd.n5224 240.244
R12047 gnd.n5224 gnd.n5202 240.244
R12048 gnd.n6056 gnd.n5202 240.244
R12049 gnd.n6056 gnd.n5197 240.244
R12050 gnd.n6064 gnd.n5197 240.244
R12051 gnd.n6064 gnd.n5198 240.244
R12052 gnd.n5198 gnd.n5175 240.244
R12053 gnd.n6102 gnd.n5175 240.244
R12054 gnd.n6102 gnd.n5170 240.244
R12055 gnd.n6110 gnd.n5170 240.244
R12056 gnd.n6110 gnd.n5171 240.244
R12057 gnd.n5171 gnd.n5148 240.244
R12058 gnd.n6398 gnd.n5148 240.244
R12059 gnd.n6398 gnd.n5143 240.244
R12060 gnd.n6409 gnd.n5143 240.244
R12061 gnd.n6409 gnd.n5144 240.244
R12062 gnd.n5144 gnd.n5122 240.244
R12063 gnd.n6516 gnd.n5122 240.244
R12064 gnd.n6517 gnd.n6516 240.244
R12065 gnd.n6517 gnd.n5118 240.244
R12066 gnd.n349 gnd.n251 240.244
R12067 gnd.n475 gnd.n474 240.244
R12068 gnd.n471 gnd.n470 240.244
R12069 gnd.n467 gnd.n466 240.244
R12070 gnd.n463 gnd.n462 240.244
R12071 gnd.n459 gnd.n458 240.244
R12072 gnd.n455 gnd.n454 240.244
R12073 gnd.n451 gnd.n450 240.244
R12074 gnd.n447 gnd.n446 240.244
R12075 gnd.n2074 gnd.n1972 240.244
R12076 gnd.n2074 gnd.n1981 240.244
R12077 gnd.n4263 gnd.n1981 240.244
R12078 gnd.n4263 gnd.n1997 240.244
R12079 gnd.n4269 gnd.n1997 240.244
R12080 gnd.n4269 gnd.n2010 240.244
R12081 gnd.n4278 gnd.n2010 240.244
R12082 gnd.n4278 gnd.n2021 240.244
R12083 gnd.n4284 gnd.n2021 240.244
R12084 gnd.n4284 gnd.n2031 240.244
R12085 gnd.n4301 gnd.n2031 240.244
R12086 gnd.n4301 gnd.n2042 240.244
R12087 gnd.n4315 gnd.n2042 240.244
R12088 gnd.n4315 gnd.n2051 240.244
R12089 gnd.n2054 gnd.n2051 240.244
R12090 gnd.n4306 gnd.n2054 240.244
R12091 gnd.n4306 gnd.n567 240.244
R12092 gnd.n567 gnd.n554 240.244
R12093 gnd.n7394 gnd.n554 240.244
R12094 gnd.n7394 gnd.n549 240.244
R12095 gnd.n7401 gnd.n549 240.244
R12096 gnd.n7401 gnd.n538 240.244
R12097 gnd.n538 gnd.n525 240.244
R12098 gnd.n7431 gnd.n525 240.244
R12099 gnd.n7431 gnd.n521 240.244
R12100 gnd.n7437 gnd.n521 240.244
R12101 gnd.n7437 gnd.n503 240.244
R12102 gnd.n7458 gnd.n503 240.244
R12103 gnd.n7458 gnd.n498 240.244
R12104 gnd.n7464 gnd.n498 240.244
R12105 gnd.n7464 gnd.n493 240.244
R12106 gnd.n493 gnd.n492 240.244
R12107 gnd.n492 gnd.n98 240.244
R12108 gnd.n7758 gnd.n98 240.244
R12109 gnd.n7758 gnd.n100 240.244
R12110 gnd.n383 gnd.n100 240.244
R12111 gnd.n383 gnd.n119 240.244
R12112 gnd.n388 gnd.n119 240.244
R12113 gnd.n388 gnd.n130 240.244
R12114 gnd.n391 gnd.n130 240.244
R12115 gnd.n391 gnd.n139 240.244
R12116 gnd.n396 gnd.n139 240.244
R12117 gnd.n396 gnd.n148 240.244
R12118 gnd.n399 gnd.n148 240.244
R12119 gnd.n399 gnd.n158 240.244
R12120 gnd.n404 gnd.n158 240.244
R12121 gnd.n404 gnd.n167 240.244
R12122 gnd.n407 gnd.n167 240.244
R12123 gnd.n407 gnd.n177 240.244
R12124 gnd.n412 gnd.n177 240.244
R12125 gnd.n412 gnd.n186 240.244
R12126 gnd.n415 gnd.n186 240.244
R12127 gnd.n415 gnd.n196 240.244
R12128 gnd.n420 gnd.n196 240.244
R12129 gnd.n420 gnd.n205 240.244
R12130 gnd.n423 gnd.n205 240.244
R12131 gnd.n423 gnd.n215 240.244
R12132 gnd.n428 gnd.n215 240.244
R12133 gnd.n428 gnd.n224 240.244
R12134 gnd.n431 gnd.n224 240.244
R12135 gnd.n431 gnd.n234 240.244
R12136 gnd.n436 gnd.n234 240.244
R12137 gnd.n436 gnd.n243 240.244
R12138 gnd.n440 gnd.n243 240.244
R12139 gnd.n1816 gnd.n1815 240.244
R12140 gnd.n1891 gnd.n1823 240.244
R12141 gnd.n1894 gnd.n1824 240.244
R12142 gnd.n1832 gnd.n1831 240.244
R12143 gnd.n1896 gnd.n1839 240.244
R12144 gnd.n1899 gnd.n1840 240.244
R12145 gnd.n1848 gnd.n1847 240.244
R12146 gnd.n1901 gnd.n1857 240.244
R12147 gnd.n4503 gnd.n1860 240.244
R12148 gnd.n4379 gnd.n1975 240.244
R12149 gnd.n1983 gnd.n1975 240.244
R12150 gnd.n1999 gnd.n1983 240.244
R12151 gnd.n4365 gnd.n1999 240.244
R12152 gnd.n4365 gnd.n2000 240.244
R12153 gnd.n4361 gnd.n2000 240.244
R12154 gnd.n4361 gnd.n2007 240.244
R12155 gnd.n4353 gnd.n2007 240.244
R12156 gnd.n4353 gnd.n2023 240.244
R12157 gnd.n4349 gnd.n2023 240.244
R12158 gnd.n4349 gnd.n2028 240.244
R12159 gnd.n4341 gnd.n2028 240.244
R12160 gnd.n4341 gnd.n2043 240.244
R12161 gnd.n4337 gnd.n2043 240.244
R12162 gnd.n4337 gnd.n2048 240.244
R12163 gnd.n2048 gnd.n568 240.244
R12164 gnd.n7382 gnd.n568 240.244
R12165 gnd.n7382 gnd.n569 240.244
R12166 gnd.n569 gnd.n558 240.244
R12167 gnd.n7377 gnd.n558 240.244
R12168 gnd.n7377 gnd.n540 240.244
R12169 gnd.n7418 gnd.n540 240.244
R12170 gnd.n7418 gnd.n541 240.244
R12171 gnd.n541 gnd.n529 240.244
R12172 gnd.n7413 gnd.n529 240.244
R12173 gnd.n7413 gnd.n511 240.244
R12174 gnd.n7451 gnd.n511 240.244
R12175 gnd.n7451 gnd.n506 240.244
R12176 gnd.n7447 gnd.n506 240.244
R12177 gnd.n7447 gnd.n490 240.244
R12178 gnd.n7474 gnd.n490 240.244
R12179 gnd.n7474 gnd.n484 240.244
R12180 gnd.n7483 gnd.n484 240.244
R12181 gnd.n7483 gnd.n103 240.244
R12182 gnd.n7486 gnd.n103 240.244
R12183 gnd.n7486 gnd.n121 240.244
R12184 gnd.n7748 gnd.n121 240.244
R12185 gnd.n7748 gnd.n122 240.244
R12186 gnd.n7744 gnd.n122 240.244
R12187 gnd.n7744 gnd.n128 240.244
R12188 gnd.n7736 gnd.n128 240.244
R12189 gnd.n7736 gnd.n140 240.244
R12190 gnd.n7732 gnd.n140 240.244
R12191 gnd.n7732 gnd.n145 240.244
R12192 gnd.n7724 gnd.n145 240.244
R12193 gnd.n7724 gnd.n160 240.244
R12194 gnd.n7720 gnd.n160 240.244
R12195 gnd.n7720 gnd.n165 240.244
R12196 gnd.n7712 gnd.n165 240.244
R12197 gnd.n7712 gnd.n178 240.244
R12198 gnd.n7708 gnd.n178 240.244
R12199 gnd.n7708 gnd.n183 240.244
R12200 gnd.n7700 gnd.n183 240.244
R12201 gnd.n7700 gnd.n198 240.244
R12202 gnd.n7696 gnd.n198 240.244
R12203 gnd.n7696 gnd.n203 240.244
R12204 gnd.n7688 gnd.n203 240.244
R12205 gnd.n7688 gnd.n216 240.244
R12206 gnd.n7684 gnd.n216 240.244
R12207 gnd.n7684 gnd.n221 240.244
R12208 gnd.n7676 gnd.n221 240.244
R12209 gnd.n7676 gnd.n236 240.244
R12210 gnd.n7672 gnd.n236 240.244
R12211 gnd.n7672 gnd.n241 240.244
R12212 gnd.n6442 gnd.n1122 240.244
R12213 gnd.n6445 gnd.n6444 240.244
R12214 gnd.n6452 gnd.n6451 240.244
R12215 gnd.n6455 gnd.n6454 240.244
R12216 gnd.n6462 gnd.n6461 240.244
R12217 gnd.n6465 gnd.n6464 240.244
R12218 gnd.n6472 gnd.n6471 240.244
R12219 gnd.n6475 gnd.n6474 240.244
R12220 gnd.n6482 gnd.n6481 240.244
R12221 gnd.n6485 gnd.n6484 240.244
R12222 gnd.n6492 gnd.n6491 240.244
R12223 gnd.n6498 gnd.n6497 240.244
R12224 gnd.n6505 gnd.n6504 240.244
R12225 gnd.n5622 gnd.n5518 240.244
R12226 gnd.n5628 gnd.n5518 240.244
R12227 gnd.n5628 gnd.n5510 240.244
R12228 gnd.n5638 gnd.n5510 240.244
R12229 gnd.n5638 gnd.n5506 240.244
R12230 gnd.n5644 gnd.n5506 240.244
R12231 gnd.n5644 gnd.n5497 240.244
R12232 gnd.n5654 gnd.n5497 240.244
R12233 gnd.n5654 gnd.n5492 240.244
R12234 gnd.n5682 gnd.n5492 240.244
R12235 gnd.n5682 gnd.n5493 240.244
R12236 gnd.n5493 gnd.n5485 240.244
R12237 gnd.n5677 gnd.n5485 240.244
R12238 gnd.n5677 gnd.n5475 240.244
R12239 gnd.n5674 gnd.n5475 240.244
R12240 gnd.n5674 gnd.n5464 240.244
R12241 gnd.n5671 gnd.n5464 240.244
R12242 gnd.n5671 gnd.n5454 240.244
R12243 gnd.n5668 gnd.n5454 240.244
R12244 gnd.n5668 gnd.n5432 240.244
R12245 gnd.n5817 gnd.n5432 240.244
R12246 gnd.n5817 gnd.n5428 240.244
R12247 gnd.n5825 gnd.n5428 240.244
R12248 gnd.n5825 gnd.n5418 240.244
R12249 gnd.n5418 gnd.n5399 240.244
R12250 gnd.n5864 gnd.n5399 240.244
R12251 gnd.n5864 gnd.n5400 240.244
R12252 gnd.n5400 gnd.n5395 240.244
R12253 gnd.n5884 gnd.n5395 240.244
R12254 gnd.n5884 gnd.n5385 240.244
R12255 gnd.n5879 gnd.n5385 240.244
R12256 gnd.n5879 gnd.n5379 240.244
R12257 gnd.n5875 gnd.n5379 240.244
R12258 gnd.n5875 gnd.n5368 240.244
R12259 gnd.n5871 gnd.n5368 240.244
R12260 gnd.n5871 gnd.n5346 240.244
R12261 gnd.n5950 gnd.n5346 240.244
R12262 gnd.n5950 gnd.n5262 240.244
R12263 gnd.n5968 gnd.n5262 240.244
R12264 gnd.n5968 gnd.n5251 240.244
R12265 gnd.n5964 gnd.n5251 240.244
R12266 gnd.n5964 gnd.n5244 240.244
R12267 gnd.n5961 gnd.n5244 240.244
R12268 gnd.n5961 gnd.n5231 240.244
R12269 gnd.n5231 gnd.n5220 240.244
R12270 gnd.n6023 gnd.n5220 240.244
R12271 gnd.n6023 gnd.n5215 240.244
R12272 gnd.n6034 gnd.n5215 240.244
R12273 gnd.n6034 gnd.n5204 240.244
R12274 gnd.n6030 gnd.n5204 240.244
R12275 gnd.n6030 gnd.n5183 240.244
R12276 gnd.n6077 gnd.n5183 240.244
R12277 gnd.n6077 gnd.n5179 240.244
R12278 gnd.n6099 gnd.n5179 240.244
R12279 gnd.n6099 gnd.n5169 240.244
R12280 gnd.n6095 gnd.n5169 240.244
R12281 gnd.n6095 gnd.n5162 240.244
R12282 gnd.n6091 gnd.n5162 240.244
R12283 gnd.n6091 gnd.n5151 240.244
R12284 gnd.n6088 gnd.n5151 240.244
R12285 gnd.n6088 gnd.n5129 240.244
R12286 gnd.n6422 gnd.n5129 240.244
R12287 gnd.n6422 gnd.n5125 240.244
R12288 gnd.n6513 gnd.n5125 240.244
R12289 gnd.n6513 gnd.n1119 240.244
R12290 gnd.n5614 gnd.n5612 240.244
R12291 gnd.n5612 gnd.n5611 240.244
R12292 gnd.n5608 gnd.n5607 240.244
R12293 gnd.n5605 gnd.n5531 240.244
R12294 gnd.n5601 gnd.n5599 240.244
R12295 gnd.n5597 gnd.n5537 240.244
R12296 gnd.n5593 gnd.n5591 240.244
R12297 gnd.n5589 gnd.n5543 240.244
R12298 gnd.n5585 gnd.n5583 240.244
R12299 gnd.n5581 gnd.n5549 240.244
R12300 gnd.n5577 gnd.n5575 240.244
R12301 gnd.n5573 gnd.n5555 240.244
R12302 gnd.n5568 gnd.n5566 240.244
R12303 gnd.n5620 gnd.n5516 240.244
R12304 gnd.n5630 gnd.n5516 240.244
R12305 gnd.n5630 gnd.n5512 240.244
R12306 gnd.n5636 gnd.n5512 240.244
R12307 gnd.n5636 gnd.n5504 240.244
R12308 gnd.n5646 gnd.n5504 240.244
R12309 gnd.n5646 gnd.n5500 240.244
R12310 gnd.n5652 gnd.n5500 240.244
R12311 gnd.n5652 gnd.n5491 240.244
R12312 gnd.n5744 gnd.n5491 240.244
R12313 gnd.n5744 gnd.n5486 240.244
R12314 gnd.n5751 gnd.n5486 240.244
R12315 gnd.n5751 gnd.n5477 240.244
R12316 gnd.n5761 gnd.n5477 240.244
R12317 gnd.n5761 gnd.n5463 240.244
R12318 gnd.n5776 gnd.n5463 240.244
R12319 gnd.n5776 gnd.n5456 240.244
R12320 gnd.n5791 gnd.n5456 240.244
R12321 gnd.n5791 gnd.n5457 240.244
R12322 gnd.n5457 gnd.n5435 240.244
R12323 gnd.n5815 gnd.n5435 240.244
R12324 gnd.n5815 gnd.n5436 240.244
R12325 gnd.n5436 gnd.n5416 240.244
R12326 gnd.n5842 gnd.n5416 240.244
R12327 gnd.n5842 gnd.n5403 240.244
R12328 gnd.n5862 gnd.n5403 240.244
R12329 gnd.n5862 gnd.n5404 240.244
R12330 gnd.n5858 gnd.n5404 240.244
R12331 gnd.n5858 gnd.n5384 240.244
R12332 gnd.n5900 gnd.n5384 240.244
R12333 gnd.n5900 gnd.n5377 240.244
R12334 gnd.n5911 gnd.n5377 240.244
R12335 gnd.n5911 gnd.n5370 240.244
R12336 gnd.n5926 gnd.n5370 240.244
R12337 gnd.n5926 gnd.n5371 240.244
R12338 gnd.n5371 gnd.n5349 240.244
R12339 gnd.n5948 gnd.n5349 240.244
R12340 gnd.n5948 gnd.n5350 240.244
R12341 gnd.n5350 gnd.n5249 240.244
R12342 gnd.n5982 gnd.n5249 240.244
R12343 gnd.n5982 gnd.n5242 240.244
R12344 gnd.n5993 gnd.n5242 240.244
R12345 gnd.n5993 gnd.n5233 240.244
R12346 gnd.n6009 gnd.n5233 240.244
R12347 gnd.n6009 gnd.n5234 240.244
R12348 gnd.n5234 gnd.n5213 240.244
R12349 gnd.n6038 gnd.n5213 240.244
R12350 gnd.n6038 gnd.n5206 240.244
R12351 gnd.n6053 gnd.n5206 240.244
R12352 gnd.n6053 gnd.n5207 240.244
R12353 gnd.n5207 gnd.n5186 240.244
R12354 gnd.n6075 gnd.n5186 240.244
R12355 gnd.n6075 gnd.n5187 240.244
R12356 gnd.n5187 gnd.n5167 240.244
R12357 gnd.n6113 gnd.n5167 240.244
R12358 gnd.n6113 gnd.n5160 240.244
R12359 gnd.n6124 gnd.n5160 240.244
R12360 gnd.n6124 gnd.n5153 240.244
R12361 gnd.n6395 gnd.n5153 240.244
R12362 gnd.n6395 gnd.n5154 240.244
R12363 gnd.n5154 gnd.n5132 240.244
R12364 gnd.n6420 gnd.n5132 240.244
R12365 gnd.n6420 gnd.n5133 240.244
R12366 gnd.n5133 gnd.n1121 240.244
R12367 gnd.n6574 gnd.n1121 240.244
R12368 gnd.n3064 gnd.n1553 240.244
R12369 gnd.n3074 gnd.n3073 240.244
R12370 gnd.n3076 gnd.n3075 240.244
R12371 gnd.n3084 gnd.n3083 240.244
R12372 gnd.n3094 gnd.n3093 240.244
R12373 gnd.n3096 gnd.n3095 240.244
R12374 gnd.n3104 gnd.n3103 240.244
R12375 gnd.n3114 gnd.n3113 240.244
R12376 gnd.n3116 gnd.n3115 240.244
R12377 gnd.n2803 gnd.n1260 240.244
R12378 gnd.n2806 gnd.n1260 240.244
R12379 gnd.n2806 gnd.n1272 240.244
R12380 gnd.n2811 gnd.n1272 240.244
R12381 gnd.n2811 gnd.n1284 240.244
R12382 gnd.n2814 gnd.n1284 240.244
R12383 gnd.n2814 gnd.n1294 240.244
R12384 gnd.n2819 gnd.n1294 240.244
R12385 gnd.n2819 gnd.n1303 240.244
R12386 gnd.n2822 gnd.n1303 240.244
R12387 gnd.n2822 gnd.n1313 240.244
R12388 gnd.n2827 gnd.n1313 240.244
R12389 gnd.n2827 gnd.n1322 240.244
R12390 gnd.n2830 gnd.n1322 240.244
R12391 gnd.n2830 gnd.n1332 240.244
R12392 gnd.n2835 gnd.n1332 240.244
R12393 gnd.n2835 gnd.n1341 240.244
R12394 gnd.n2838 gnd.n1341 240.244
R12395 gnd.n2838 gnd.n1351 240.244
R12396 gnd.n2843 gnd.n1351 240.244
R12397 gnd.n2843 gnd.n1360 240.244
R12398 gnd.n2846 gnd.n1360 240.244
R12399 gnd.n2846 gnd.n1370 240.244
R12400 gnd.n2851 gnd.n1370 240.244
R12401 gnd.n2851 gnd.n1379 240.244
R12402 gnd.n2854 gnd.n1379 240.244
R12403 gnd.n2854 gnd.n1388 240.244
R12404 gnd.n2859 gnd.n1388 240.244
R12405 gnd.n2859 gnd.n1397 240.244
R12406 gnd.n2862 gnd.n1397 240.244
R12407 gnd.n2862 gnd.n2727 240.244
R12408 gnd.n2868 gnd.n2727 240.244
R12409 gnd.n2868 gnd.n2647 240.244
R12410 gnd.n2892 gnd.n2647 240.244
R12411 gnd.n2892 gnd.n2643 240.244
R12412 gnd.n2898 gnd.n2643 240.244
R12413 gnd.n2898 gnd.n1413 240.244
R12414 gnd.n2931 gnd.n1413 240.244
R12415 gnd.n2931 gnd.n1424 240.244
R12416 gnd.n2937 gnd.n1424 240.244
R12417 gnd.n2937 gnd.n1434 240.244
R12418 gnd.n2945 gnd.n1434 240.244
R12419 gnd.n2945 gnd.n1443 240.244
R12420 gnd.n2951 gnd.n1443 240.244
R12421 gnd.n2951 gnd.n1454 240.244
R12422 gnd.n2986 gnd.n1454 240.244
R12423 gnd.n2986 gnd.n1463 240.244
R12424 gnd.n2620 gnd.n1463 240.244
R12425 gnd.n2620 gnd.n1474 240.244
R12426 gnd.n2621 gnd.n1474 240.244
R12427 gnd.n2621 gnd.n1483 240.244
R12428 gnd.n2974 gnd.n1483 240.244
R12429 gnd.n2974 gnd.n1494 240.244
R12430 gnd.n3012 gnd.n1494 240.244
R12431 gnd.n3012 gnd.n1503 240.244
R12432 gnd.n3018 gnd.n1503 240.244
R12433 gnd.n3018 gnd.n1514 240.244
R12434 gnd.n3290 gnd.n1514 240.244
R12435 gnd.n3290 gnd.n1523 240.244
R12436 gnd.n2597 gnd.n1523 240.244
R12437 gnd.n2597 gnd.n1534 240.244
R12438 gnd.n3279 gnd.n1534 240.244
R12439 gnd.n3279 gnd.n1544 240.244
R12440 gnd.n3319 gnd.n1544 240.244
R12441 gnd.n2763 gnd.n2762 240.244
R12442 gnd.n2769 gnd.n2768 240.244
R12443 gnd.n2773 gnd.n2772 240.244
R12444 gnd.n2779 gnd.n2778 240.244
R12445 gnd.n2783 gnd.n2782 240.244
R12446 gnd.n2789 gnd.n2788 240.244
R12447 gnd.n2793 gnd.n2792 240.244
R12448 gnd.n2750 gnd.n2749 240.244
R12449 gnd.n2745 gnd.n1185 240.244
R12450 gnd.n2758 gnd.n1261 240.244
R12451 gnd.n1274 gnd.n1261 240.244
R12452 gnd.n4980 gnd.n1274 240.244
R12453 gnd.n4980 gnd.n1275 240.244
R12454 gnd.n4976 gnd.n1275 240.244
R12455 gnd.n4976 gnd.n1282 240.244
R12456 gnd.n4968 gnd.n1282 240.244
R12457 gnd.n4968 gnd.n1296 240.244
R12458 gnd.n4964 gnd.n1296 240.244
R12459 gnd.n4964 gnd.n1301 240.244
R12460 gnd.n4956 gnd.n1301 240.244
R12461 gnd.n4956 gnd.n1315 240.244
R12462 gnd.n4952 gnd.n1315 240.244
R12463 gnd.n4952 gnd.n1320 240.244
R12464 gnd.n4944 gnd.n1320 240.244
R12465 gnd.n4944 gnd.n1334 240.244
R12466 gnd.n4940 gnd.n1334 240.244
R12467 gnd.n4940 gnd.n1339 240.244
R12468 gnd.n4932 gnd.n1339 240.244
R12469 gnd.n4932 gnd.n1353 240.244
R12470 gnd.n4928 gnd.n1353 240.244
R12471 gnd.n4928 gnd.n1358 240.244
R12472 gnd.n4920 gnd.n1358 240.244
R12473 gnd.n4920 gnd.n1372 240.244
R12474 gnd.n4916 gnd.n1372 240.244
R12475 gnd.n4916 gnd.n1377 240.244
R12476 gnd.n4908 gnd.n1377 240.244
R12477 gnd.n4908 gnd.n1390 240.244
R12478 gnd.n4904 gnd.n1390 240.244
R12479 gnd.n4904 gnd.n1395 240.244
R12480 gnd.n2723 gnd.n1395 240.244
R12481 gnd.n2723 gnd.n2662 240.244
R12482 gnd.n2884 gnd.n2662 240.244
R12483 gnd.n2884 gnd.n2650 240.244
R12484 gnd.n2880 gnd.n2650 240.244
R12485 gnd.n2880 gnd.n1415 240.244
R12486 gnd.n4895 gnd.n1415 240.244
R12487 gnd.n4895 gnd.n1416 240.244
R12488 gnd.n4891 gnd.n1416 240.244
R12489 gnd.n4891 gnd.n1422 240.244
R12490 gnd.n4883 gnd.n1422 240.244
R12491 gnd.n4883 gnd.n1435 240.244
R12492 gnd.n4879 gnd.n1435 240.244
R12493 gnd.n4879 gnd.n1440 240.244
R12494 gnd.n4871 gnd.n1440 240.244
R12495 gnd.n4871 gnd.n1456 240.244
R12496 gnd.n4867 gnd.n1456 240.244
R12497 gnd.n4867 gnd.n1461 240.244
R12498 gnd.n4859 gnd.n1461 240.244
R12499 gnd.n4859 gnd.n1475 240.244
R12500 gnd.n4855 gnd.n1475 240.244
R12501 gnd.n4855 gnd.n1480 240.244
R12502 gnd.n4847 gnd.n1480 240.244
R12503 gnd.n4847 gnd.n1496 240.244
R12504 gnd.n4843 gnd.n1496 240.244
R12505 gnd.n4843 gnd.n1501 240.244
R12506 gnd.n4835 gnd.n1501 240.244
R12507 gnd.n4835 gnd.n1515 240.244
R12508 gnd.n4831 gnd.n1515 240.244
R12509 gnd.n4831 gnd.n1520 240.244
R12510 gnd.n4823 gnd.n1520 240.244
R12511 gnd.n4823 gnd.n1536 240.244
R12512 gnd.n4819 gnd.n1536 240.244
R12513 gnd.n4819 gnd.n1541 240.244
R12514 gnd.n6747 gnd.n950 240.244
R12515 gnd.n6747 gnd.n946 240.244
R12516 gnd.n6753 gnd.n946 240.244
R12517 gnd.n6753 gnd.n944 240.244
R12518 gnd.n6757 gnd.n944 240.244
R12519 gnd.n6757 gnd.n940 240.244
R12520 gnd.n6763 gnd.n940 240.244
R12521 gnd.n6763 gnd.n938 240.244
R12522 gnd.n6767 gnd.n938 240.244
R12523 gnd.n6767 gnd.n934 240.244
R12524 gnd.n6773 gnd.n934 240.244
R12525 gnd.n6773 gnd.n932 240.244
R12526 gnd.n6777 gnd.n932 240.244
R12527 gnd.n6777 gnd.n928 240.244
R12528 gnd.n6783 gnd.n928 240.244
R12529 gnd.n6783 gnd.n926 240.244
R12530 gnd.n6787 gnd.n926 240.244
R12531 gnd.n6787 gnd.n922 240.244
R12532 gnd.n6793 gnd.n922 240.244
R12533 gnd.n6793 gnd.n920 240.244
R12534 gnd.n6797 gnd.n920 240.244
R12535 gnd.n6797 gnd.n916 240.244
R12536 gnd.n6803 gnd.n916 240.244
R12537 gnd.n6803 gnd.n914 240.244
R12538 gnd.n6807 gnd.n914 240.244
R12539 gnd.n6807 gnd.n910 240.244
R12540 gnd.n6813 gnd.n910 240.244
R12541 gnd.n6813 gnd.n908 240.244
R12542 gnd.n6817 gnd.n908 240.244
R12543 gnd.n6817 gnd.n904 240.244
R12544 gnd.n6823 gnd.n904 240.244
R12545 gnd.n6823 gnd.n902 240.244
R12546 gnd.n6827 gnd.n902 240.244
R12547 gnd.n6827 gnd.n898 240.244
R12548 gnd.n6833 gnd.n898 240.244
R12549 gnd.n6833 gnd.n896 240.244
R12550 gnd.n6837 gnd.n896 240.244
R12551 gnd.n6837 gnd.n892 240.244
R12552 gnd.n6843 gnd.n892 240.244
R12553 gnd.n6843 gnd.n890 240.244
R12554 gnd.n6847 gnd.n890 240.244
R12555 gnd.n6847 gnd.n886 240.244
R12556 gnd.n6853 gnd.n886 240.244
R12557 gnd.n6853 gnd.n884 240.244
R12558 gnd.n6857 gnd.n884 240.244
R12559 gnd.n6857 gnd.n880 240.244
R12560 gnd.n6863 gnd.n880 240.244
R12561 gnd.n6863 gnd.n878 240.244
R12562 gnd.n6867 gnd.n878 240.244
R12563 gnd.n6867 gnd.n874 240.244
R12564 gnd.n6873 gnd.n874 240.244
R12565 gnd.n6873 gnd.n872 240.244
R12566 gnd.n6877 gnd.n872 240.244
R12567 gnd.n6877 gnd.n868 240.244
R12568 gnd.n6883 gnd.n868 240.244
R12569 gnd.n6883 gnd.n866 240.244
R12570 gnd.n6887 gnd.n866 240.244
R12571 gnd.n6887 gnd.n862 240.244
R12572 gnd.n6893 gnd.n862 240.244
R12573 gnd.n6893 gnd.n860 240.244
R12574 gnd.n6897 gnd.n860 240.244
R12575 gnd.n6897 gnd.n856 240.244
R12576 gnd.n6903 gnd.n856 240.244
R12577 gnd.n6903 gnd.n854 240.244
R12578 gnd.n6907 gnd.n854 240.244
R12579 gnd.n6907 gnd.n850 240.244
R12580 gnd.n6913 gnd.n850 240.244
R12581 gnd.n6913 gnd.n848 240.244
R12582 gnd.n6917 gnd.n848 240.244
R12583 gnd.n6917 gnd.n844 240.244
R12584 gnd.n6923 gnd.n844 240.244
R12585 gnd.n6923 gnd.n842 240.244
R12586 gnd.n6927 gnd.n842 240.244
R12587 gnd.n6927 gnd.n838 240.244
R12588 gnd.n6933 gnd.n838 240.244
R12589 gnd.n6933 gnd.n836 240.244
R12590 gnd.n6937 gnd.n836 240.244
R12591 gnd.n6937 gnd.n832 240.244
R12592 gnd.n6943 gnd.n832 240.244
R12593 gnd.n6943 gnd.n830 240.244
R12594 gnd.n6947 gnd.n830 240.244
R12595 gnd.n6947 gnd.n826 240.244
R12596 gnd.n6953 gnd.n826 240.244
R12597 gnd.n6953 gnd.n824 240.244
R12598 gnd.n6957 gnd.n824 240.244
R12599 gnd.n6957 gnd.n820 240.244
R12600 gnd.n6963 gnd.n820 240.244
R12601 gnd.n6963 gnd.n818 240.244
R12602 gnd.n6967 gnd.n818 240.244
R12603 gnd.n6967 gnd.n814 240.244
R12604 gnd.n6973 gnd.n814 240.244
R12605 gnd.n6973 gnd.n812 240.244
R12606 gnd.n6977 gnd.n812 240.244
R12607 gnd.n6977 gnd.n808 240.244
R12608 gnd.n6983 gnd.n808 240.244
R12609 gnd.n6983 gnd.n806 240.244
R12610 gnd.n6987 gnd.n806 240.244
R12611 gnd.n6987 gnd.n802 240.244
R12612 gnd.n6993 gnd.n802 240.244
R12613 gnd.n6993 gnd.n800 240.244
R12614 gnd.n6997 gnd.n800 240.244
R12615 gnd.n6997 gnd.n796 240.244
R12616 gnd.n7003 gnd.n796 240.244
R12617 gnd.n7003 gnd.n794 240.244
R12618 gnd.n7007 gnd.n794 240.244
R12619 gnd.n7007 gnd.n790 240.244
R12620 gnd.n7013 gnd.n790 240.244
R12621 gnd.n7013 gnd.n788 240.244
R12622 gnd.n7017 gnd.n788 240.244
R12623 gnd.n7017 gnd.n784 240.244
R12624 gnd.n7023 gnd.n784 240.244
R12625 gnd.n7023 gnd.n782 240.244
R12626 gnd.n7027 gnd.n782 240.244
R12627 gnd.n7027 gnd.n778 240.244
R12628 gnd.n7033 gnd.n778 240.244
R12629 gnd.n7033 gnd.n776 240.244
R12630 gnd.n7037 gnd.n776 240.244
R12631 gnd.n7037 gnd.n772 240.244
R12632 gnd.n7043 gnd.n772 240.244
R12633 gnd.n7043 gnd.n770 240.244
R12634 gnd.n7047 gnd.n770 240.244
R12635 gnd.n7047 gnd.n766 240.244
R12636 gnd.n7053 gnd.n766 240.244
R12637 gnd.n7053 gnd.n764 240.244
R12638 gnd.n7057 gnd.n764 240.244
R12639 gnd.n7057 gnd.n760 240.244
R12640 gnd.n7063 gnd.n760 240.244
R12641 gnd.n7063 gnd.n758 240.244
R12642 gnd.n7067 gnd.n758 240.244
R12643 gnd.n7067 gnd.n754 240.244
R12644 gnd.n7073 gnd.n754 240.244
R12645 gnd.n7073 gnd.n752 240.244
R12646 gnd.n7077 gnd.n752 240.244
R12647 gnd.n7077 gnd.n748 240.244
R12648 gnd.n7083 gnd.n748 240.244
R12649 gnd.n7083 gnd.n746 240.244
R12650 gnd.n7087 gnd.n746 240.244
R12651 gnd.n7087 gnd.n742 240.244
R12652 gnd.n7093 gnd.n742 240.244
R12653 gnd.n7093 gnd.n740 240.244
R12654 gnd.n7097 gnd.n740 240.244
R12655 gnd.n7097 gnd.n736 240.244
R12656 gnd.n7103 gnd.n736 240.244
R12657 gnd.n7103 gnd.n734 240.244
R12658 gnd.n7107 gnd.n734 240.244
R12659 gnd.n7107 gnd.n730 240.244
R12660 gnd.n7113 gnd.n730 240.244
R12661 gnd.n7113 gnd.n728 240.244
R12662 gnd.n7117 gnd.n728 240.244
R12663 gnd.n7117 gnd.n724 240.244
R12664 gnd.n7124 gnd.n724 240.244
R12665 gnd.n7124 gnd.n722 240.244
R12666 gnd.n7128 gnd.n722 240.244
R12667 gnd.n7128 gnd.n719 240.244
R12668 gnd.n7134 gnd.n717 240.244
R12669 gnd.n7138 gnd.n717 240.244
R12670 gnd.n7138 gnd.n713 240.244
R12671 gnd.n7144 gnd.n713 240.244
R12672 gnd.n7144 gnd.n711 240.244
R12673 gnd.n7148 gnd.n711 240.244
R12674 gnd.n7148 gnd.n707 240.244
R12675 gnd.n7154 gnd.n707 240.244
R12676 gnd.n7154 gnd.n705 240.244
R12677 gnd.n7158 gnd.n705 240.244
R12678 gnd.n7158 gnd.n701 240.244
R12679 gnd.n7164 gnd.n701 240.244
R12680 gnd.n7164 gnd.n699 240.244
R12681 gnd.n7168 gnd.n699 240.244
R12682 gnd.n7168 gnd.n695 240.244
R12683 gnd.n7174 gnd.n695 240.244
R12684 gnd.n7174 gnd.n693 240.244
R12685 gnd.n7178 gnd.n693 240.244
R12686 gnd.n7178 gnd.n689 240.244
R12687 gnd.n7184 gnd.n689 240.244
R12688 gnd.n7184 gnd.n687 240.244
R12689 gnd.n7188 gnd.n687 240.244
R12690 gnd.n7188 gnd.n683 240.244
R12691 gnd.n7194 gnd.n683 240.244
R12692 gnd.n7194 gnd.n681 240.244
R12693 gnd.n7198 gnd.n681 240.244
R12694 gnd.n7198 gnd.n677 240.244
R12695 gnd.n7204 gnd.n677 240.244
R12696 gnd.n7204 gnd.n675 240.244
R12697 gnd.n7208 gnd.n675 240.244
R12698 gnd.n7208 gnd.n671 240.244
R12699 gnd.n7214 gnd.n671 240.244
R12700 gnd.n7214 gnd.n669 240.244
R12701 gnd.n7218 gnd.n669 240.244
R12702 gnd.n7218 gnd.n665 240.244
R12703 gnd.n7224 gnd.n665 240.244
R12704 gnd.n7224 gnd.n663 240.244
R12705 gnd.n7228 gnd.n663 240.244
R12706 gnd.n7228 gnd.n659 240.244
R12707 gnd.n7234 gnd.n659 240.244
R12708 gnd.n7234 gnd.n657 240.244
R12709 gnd.n7238 gnd.n657 240.244
R12710 gnd.n7238 gnd.n653 240.244
R12711 gnd.n7244 gnd.n653 240.244
R12712 gnd.n7244 gnd.n651 240.244
R12713 gnd.n7248 gnd.n651 240.244
R12714 gnd.n7248 gnd.n647 240.244
R12715 gnd.n7254 gnd.n647 240.244
R12716 gnd.n7254 gnd.n645 240.244
R12717 gnd.n7258 gnd.n645 240.244
R12718 gnd.n7258 gnd.n641 240.244
R12719 gnd.n7264 gnd.n641 240.244
R12720 gnd.n7264 gnd.n639 240.244
R12721 gnd.n7268 gnd.n639 240.244
R12722 gnd.n7268 gnd.n635 240.244
R12723 gnd.n7274 gnd.n635 240.244
R12724 gnd.n7274 gnd.n633 240.244
R12725 gnd.n7278 gnd.n633 240.244
R12726 gnd.n7278 gnd.n629 240.244
R12727 gnd.n7284 gnd.n629 240.244
R12728 gnd.n7284 gnd.n627 240.244
R12729 gnd.n7288 gnd.n627 240.244
R12730 gnd.n7288 gnd.n623 240.244
R12731 gnd.n7294 gnd.n623 240.244
R12732 gnd.n7294 gnd.n621 240.244
R12733 gnd.n7298 gnd.n621 240.244
R12734 gnd.n7298 gnd.n617 240.244
R12735 gnd.n7304 gnd.n617 240.244
R12736 gnd.n7304 gnd.n615 240.244
R12737 gnd.n7308 gnd.n615 240.244
R12738 gnd.n7308 gnd.n611 240.244
R12739 gnd.n7314 gnd.n611 240.244
R12740 gnd.n7314 gnd.n609 240.244
R12741 gnd.n7318 gnd.n609 240.244
R12742 gnd.n7318 gnd.n605 240.244
R12743 gnd.n7324 gnd.n605 240.244
R12744 gnd.n7324 gnd.n603 240.244
R12745 gnd.n7328 gnd.n603 240.244
R12746 gnd.n7328 gnd.n599 240.244
R12747 gnd.n7334 gnd.n599 240.244
R12748 gnd.n7334 gnd.n597 240.244
R12749 gnd.n7340 gnd.n597 240.244
R12750 gnd.n7340 gnd.n593 240.244
R12751 gnd.n7347 gnd.n593 240.244
R12752 gnd.n2901 gnd.n2640 240.244
R12753 gnd.n2902 gnd.n2901 240.244
R12754 gnd.n2902 gnd.n2635 240.244
R12755 gnd.n2928 gnd.n2635 240.244
R12756 gnd.n2928 gnd.n2636 240.244
R12757 gnd.n2924 gnd.n2636 240.244
R12758 gnd.n2924 gnd.n2923 240.244
R12759 gnd.n2923 gnd.n2922 240.244
R12760 gnd.n2922 gnd.n2910 240.244
R12761 gnd.n2918 gnd.n2910 240.244
R12762 gnd.n2918 gnd.n2613 240.244
R12763 gnd.n2989 gnd.n2613 240.244
R12764 gnd.n2990 gnd.n2989 240.244
R12765 gnd.n2991 gnd.n2990 240.244
R12766 gnd.n2991 gnd.n2609 240.244
R12767 gnd.n2997 gnd.n2609 240.244
R12768 gnd.n2998 gnd.n2997 240.244
R12769 gnd.n2999 gnd.n2998 240.244
R12770 gnd.n2999 gnd.n2604 240.244
R12771 gnd.n3009 gnd.n2604 240.244
R12772 gnd.n3009 gnd.n2605 240.244
R12773 gnd.n2605 gnd.n2591 240.244
R12774 gnd.n3293 gnd.n2591 240.244
R12775 gnd.n3294 gnd.n3293 240.244
R12776 gnd.n3294 gnd.n2587 240.244
R12777 gnd.n3300 gnd.n2587 240.244
R12778 gnd.n3301 gnd.n3300 240.244
R12779 gnd.n3302 gnd.n3301 240.244
R12780 gnd.n3302 gnd.n2582 240.244
R12781 gnd.n3316 gnd.n2582 240.244
R12782 gnd.n3316 gnd.n2583 240.244
R12783 gnd.n3312 gnd.n2583 240.244
R12784 gnd.n3312 gnd.n3311 240.244
R12785 gnd.n3311 gnd.n2557 240.244
R12786 gnd.n3330 gnd.n2557 240.244
R12787 gnd.n3330 gnd.n2553 240.244
R12788 gnd.n3336 gnd.n2553 240.244
R12789 gnd.n3336 gnd.n2541 240.244
R12790 gnd.n3363 gnd.n2541 240.244
R12791 gnd.n3363 gnd.n2536 240.244
R12792 gnd.n3378 gnd.n2536 240.244
R12793 gnd.n3378 gnd.n2537 240.244
R12794 gnd.n3374 gnd.n2537 240.244
R12795 gnd.n3374 gnd.n3373 240.244
R12796 gnd.n3373 gnd.n1689 240.244
R12797 gnd.n4684 gnd.n1689 240.244
R12798 gnd.n4684 gnd.n1690 240.244
R12799 gnd.n4680 gnd.n1690 240.244
R12800 gnd.n4680 gnd.n1696 240.244
R12801 gnd.n2506 gnd.n1696 240.244
R12802 gnd.n3529 gnd.n2506 240.244
R12803 gnd.n3529 gnd.n2500 240.244
R12804 gnd.n3537 gnd.n2500 240.244
R12805 gnd.n3537 gnd.n2501 240.244
R12806 gnd.n2501 gnd.n2483 240.244
R12807 gnd.n3566 gnd.n2483 240.244
R12808 gnd.n3566 gnd.n2479 240.244
R12809 gnd.n3572 gnd.n2479 240.244
R12810 gnd.n3572 gnd.n2455 240.244
R12811 gnd.n3605 gnd.n2455 240.244
R12812 gnd.n3605 gnd.n2450 240.244
R12813 gnd.n3613 gnd.n2450 240.244
R12814 gnd.n3613 gnd.n2451 240.244
R12815 gnd.n2451 gnd.n2427 240.244
R12816 gnd.n3645 gnd.n2427 240.244
R12817 gnd.n3645 gnd.n2423 240.244
R12818 gnd.n3652 gnd.n2423 240.244
R12819 gnd.n3652 gnd.n2403 240.244
R12820 gnd.n3680 gnd.n2403 240.244
R12821 gnd.n3680 gnd.n2404 240.244
R12822 gnd.n3676 gnd.n2404 240.244
R12823 gnd.n3676 gnd.n3675 240.244
R12824 gnd.n3675 gnd.n3674 240.244
R12825 gnd.n3674 gnd.n2371 240.244
R12826 gnd.n3740 gnd.n2371 240.244
R12827 gnd.n3740 gnd.n2365 240.244
R12828 gnd.n3748 gnd.n2365 240.244
R12829 gnd.n3748 gnd.n2367 240.244
R12830 gnd.n2367 gnd.n2346 240.244
R12831 gnd.n3792 gnd.n2346 240.244
R12832 gnd.n3792 gnd.n2341 240.244
R12833 gnd.n3800 gnd.n2341 240.244
R12834 gnd.n3800 gnd.n2342 240.244
R12835 gnd.n2342 gnd.n2320 240.244
R12836 gnd.n3829 gnd.n2320 240.244
R12837 gnd.n3829 gnd.n2316 240.244
R12838 gnd.n3835 gnd.n2316 240.244
R12839 gnd.n3835 gnd.n2295 240.244
R12840 gnd.n3890 gnd.n2295 240.244
R12841 gnd.n3890 gnd.n2290 240.244
R12842 gnd.n3898 gnd.n2290 240.244
R12843 gnd.n3898 gnd.n2291 240.244
R12844 gnd.n2291 gnd.n2272 240.244
R12845 gnd.n3923 gnd.n2272 240.244
R12846 gnd.n3923 gnd.n2267 240.244
R12847 gnd.n3931 gnd.n2267 240.244
R12848 gnd.n3931 gnd.n2268 240.244
R12849 gnd.n2268 gnd.n2251 240.244
R12850 gnd.n3975 gnd.n2251 240.244
R12851 gnd.n3975 gnd.n2246 240.244
R12852 gnd.n3983 gnd.n2246 240.244
R12853 gnd.n3983 gnd.n2247 240.244
R12854 gnd.n2247 gnd.n2222 240.244
R12855 gnd.n4012 gnd.n2222 240.244
R12856 gnd.n4012 gnd.n2218 240.244
R12857 gnd.n4018 gnd.n2218 240.244
R12858 gnd.n4018 gnd.n2133 240.244
R12859 gnd.n4159 gnd.n2133 240.244
R12860 gnd.n4159 gnd.n2129 240.244
R12861 gnd.n4165 gnd.n2129 240.244
R12862 gnd.n4165 gnd.n2120 240.244
R12863 gnd.n4175 gnd.n2120 240.244
R12864 gnd.n4175 gnd.n2116 240.244
R12865 gnd.n4184 gnd.n2116 240.244
R12866 gnd.n4184 gnd.n2107 240.244
R12867 gnd.n4194 gnd.n2107 240.244
R12868 gnd.n4195 gnd.n4194 240.244
R12869 gnd.n4195 gnd.n1793 240.244
R12870 gnd.n2102 gnd.n1793 240.244
R12871 gnd.n4250 gnd.n2102 240.244
R12872 gnd.n4250 gnd.n2103 240.244
R12873 gnd.n4246 gnd.n2103 240.244
R12874 gnd.n4246 gnd.n4245 240.244
R12875 gnd.n4245 gnd.n4244 240.244
R12876 gnd.n4244 gnd.n4204 240.244
R12877 gnd.n4240 gnd.n4204 240.244
R12878 gnd.n4240 gnd.n4237 240.244
R12879 gnd.n4237 gnd.n4236 240.244
R12880 gnd.n4236 gnd.n4210 240.244
R12881 gnd.n4232 gnd.n4210 240.244
R12882 gnd.n4232 gnd.n4231 240.244
R12883 gnd.n4231 gnd.n4230 240.244
R12884 gnd.n4230 gnd.n4216 240.244
R12885 gnd.n4226 gnd.n4216 240.244
R12886 gnd.n4226 gnd.n4225 240.244
R12887 gnd.n4225 gnd.n2060 240.244
R12888 gnd.n4318 gnd.n2060 240.244
R12889 gnd.n4319 gnd.n4318 240.244
R12890 gnd.n4319 gnd.n2056 240.244
R12891 gnd.n4326 gnd.n2056 240.244
R12892 gnd.n4326 gnd.n574 240.244
R12893 gnd.n7368 gnd.n574 240.244
R12894 gnd.n7368 gnd.n575 240.244
R12895 gnd.n7364 gnd.n575 240.244
R12896 gnd.n7364 gnd.n7363 240.244
R12897 gnd.n7363 gnd.n7362 240.244
R12898 gnd.n7362 gnd.n581 240.244
R12899 gnd.n7358 gnd.n581 240.244
R12900 gnd.n7358 gnd.n7357 240.244
R12901 gnd.n7357 gnd.n7356 240.244
R12902 gnd.n7356 gnd.n587 240.244
R12903 gnd.n591 gnd.n587 240.244
R12904 gnd.n7349 gnd.n591 240.244
R12905 gnd.n7349 gnd.n7348 240.244
R12906 gnd.n6743 gnd.n952 240.244
R12907 gnd.n6739 gnd.n952 240.244
R12908 gnd.n6739 gnd.n957 240.244
R12909 gnd.n6735 gnd.n957 240.244
R12910 gnd.n6735 gnd.n959 240.244
R12911 gnd.n6731 gnd.n959 240.244
R12912 gnd.n6731 gnd.n965 240.244
R12913 gnd.n6727 gnd.n965 240.244
R12914 gnd.n6727 gnd.n967 240.244
R12915 gnd.n6723 gnd.n967 240.244
R12916 gnd.n6723 gnd.n973 240.244
R12917 gnd.n6719 gnd.n973 240.244
R12918 gnd.n6719 gnd.n975 240.244
R12919 gnd.n6715 gnd.n975 240.244
R12920 gnd.n6715 gnd.n981 240.244
R12921 gnd.n6711 gnd.n981 240.244
R12922 gnd.n6711 gnd.n983 240.244
R12923 gnd.n6707 gnd.n983 240.244
R12924 gnd.n6707 gnd.n989 240.244
R12925 gnd.n6703 gnd.n989 240.244
R12926 gnd.n6703 gnd.n991 240.244
R12927 gnd.n6699 gnd.n991 240.244
R12928 gnd.n6699 gnd.n997 240.244
R12929 gnd.n6695 gnd.n997 240.244
R12930 gnd.n6695 gnd.n999 240.244
R12931 gnd.n6691 gnd.n999 240.244
R12932 gnd.n6691 gnd.n1005 240.244
R12933 gnd.n6687 gnd.n1005 240.244
R12934 gnd.n6687 gnd.n1007 240.244
R12935 gnd.n6683 gnd.n1007 240.244
R12936 gnd.n6683 gnd.n1013 240.244
R12937 gnd.n6679 gnd.n1013 240.244
R12938 gnd.n6679 gnd.n1015 240.244
R12939 gnd.n6675 gnd.n1015 240.244
R12940 gnd.n6675 gnd.n1021 240.244
R12941 gnd.n6671 gnd.n1021 240.244
R12942 gnd.n6671 gnd.n1023 240.244
R12943 gnd.n6667 gnd.n1023 240.244
R12944 gnd.n6667 gnd.n1029 240.244
R12945 gnd.n6663 gnd.n1029 240.244
R12946 gnd.n6663 gnd.n1031 240.244
R12947 gnd.n6659 gnd.n1031 240.244
R12948 gnd.n6659 gnd.n1037 240.244
R12949 gnd.n6655 gnd.n1037 240.244
R12950 gnd.n6655 gnd.n1039 240.244
R12951 gnd.n6651 gnd.n1039 240.244
R12952 gnd.n6651 gnd.n1045 240.244
R12953 gnd.n6647 gnd.n1045 240.244
R12954 gnd.n6647 gnd.n1047 240.244
R12955 gnd.n6643 gnd.n1047 240.244
R12956 gnd.n6643 gnd.n1053 240.244
R12957 gnd.n6639 gnd.n1053 240.244
R12958 gnd.n6639 gnd.n1055 240.244
R12959 gnd.n6635 gnd.n1055 240.244
R12960 gnd.n6635 gnd.n1061 240.244
R12961 gnd.n6631 gnd.n1061 240.244
R12962 gnd.n6631 gnd.n1063 240.244
R12963 gnd.n6627 gnd.n1063 240.244
R12964 gnd.n6627 gnd.n1069 240.244
R12965 gnd.n6623 gnd.n1069 240.244
R12966 gnd.n6623 gnd.n1071 240.244
R12967 gnd.n6619 gnd.n1071 240.244
R12968 gnd.n6619 gnd.n1077 240.244
R12969 gnd.n6615 gnd.n1077 240.244
R12970 gnd.n6615 gnd.n1079 240.244
R12971 gnd.n6611 gnd.n1079 240.244
R12972 gnd.n6611 gnd.n1085 240.244
R12973 gnd.n6607 gnd.n1085 240.244
R12974 gnd.n6607 gnd.n1087 240.244
R12975 gnd.n6603 gnd.n1087 240.244
R12976 gnd.n6603 gnd.n1093 240.244
R12977 gnd.n6599 gnd.n1093 240.244
R12978 gnd.n6599 gnd.n1095 240.244
R12979 gnd.n6595 gnd.n1095 240.244
R12980 gnd.n6595 gnd.n1101 240.244
R12981 gnd.n6591 gnd.n1101 240.244
R12982 gnd.n6591 gnd.n1103 240.244
R12983 gnd.n6587 gnd.n1103 240.244
R12984 gnd.n6587 gnd.n1109 240.244
R12985 gnd.n6583 gnd.n1109 240.244
R12986 gnd.n6583 gnd.n1111 240.244
R12987 gnd.n6579 gnd.n1111 240.244
R12988 gnd.n6579 gnd.n1117 240.244
R12989 gnd.n2659 gnd.n1117 240.244
R12990 gnd.n3046 gnd.n2552 240.244
R12991 gnd.n3039 gnd.n2552 240.244
R12992 gnd.n3039 gnd.n2543 240.244
R12993 gnd.n2543 gnd.n2532 240.244
R12994 gnd.n3380 gnd.n2532 240.244
R12995 gnd.n3380 gnd.n2528 240.244
R12996 gnd.n3386 gnd.n2528 240.244
R12997 gnd.n3387 gnd.n3386 240.244
R12998 gnd.n3388 gnd.n3387 240.244
R12999 gnd.n3388 gnd.n1686 240.244
R13000 gnd.n3403 gnd.n1686 240.244
R13001 gnd.n3403 gnd.n1697 240.244
R13002 gnd.n3393 gnd.n1697 240.244
R13003 gnd.n3394 gnd.n3393 240.244
R13004 gnd.n3394 gnd.n2508 240.244
R13005 gnd.n2508 gnd.n2496 240.244
R13006 gnd.n3539 gnd.n2496 240.244
R13007 gnd.n3539 gnd.n2491 240.244
R13008 gnd.n3556 gnd.n2491 240.244
R13009 gnd.n3556 gnd.n2485 240.244
R13010 gnd.n3544 gnd.n2485 240.244
R13011 gnd.n3544 gnd.n2477 240.244
R13012 gnd.n3545 gnd.n2477 240.244
R13013 gnd.n3545 gnd.n2457 240.244
R13014 gnd.n2457 gnd.n2447 240.244
R13015 gnd.n3615 gnd.n2447 240.244
R13016 gnd.n3615 gnd.n2442 240.244
R13017 gnd.n3622 gnd.n2442 240.244
R13018 gnd.n3622 gnd.n2428 240.244
R13019 gnd.n2428 gnd.n2420 240.244
R13020 gnd.n3654 gnd.n2420 240.244
R13021 gnd.n3654 gnd.n2421 240.244
R13022 gnd.n2421 gnd.n2401 240.244
R13023 gnd.n3661 gnd.n2401 240.244
R13024 gnd.n3662 gnd.n3661 240.244
R13025 gnd.n3662 gnd.n2413 240.244
R13026 gnd.n3671 gnd.n2413 240.244
R13027 gnd.n3671 gnd.n2382 240.244
R13028 gnd.n2382 gnd.n2372 240.244
R13029 gnd.n2372 gnd.n2361 240.244
R13030 gnd.n3750 gnd.n2361 240.244
R13031 gnd.n3750 gnd.n2356 240.244
R13032 gnd.n3782 gnd.n2356 240.244
R13033 gnd.n3782 gnd.n2348 240.244
R13034 gnd.n3757 gnd.n2348 240.244
R13035 gnd.n3757 gnd.n2340 240.244
R13036 gnd.n3758 gnd.n2340 240.244
R13037 gnd.n3759 gnd.n3758 240.244
R13038 gnd.n3759 gnd.n2322 240.244
R13039 gnd.n3762 gnd.n2322 240.244
R13040 gnd.n3762 gnd.n2314 240.244
R13041 gnd.n3763 gnd.n2314 240.244
R13042 gnd.n3763 gnd.n2297 240.244
R13043 gnd.n2297 gnd.n2288 240.244
R13044 gnd.n3900 gnd.n2288 240.244
R13045 gnd.n3900 gnd.n2283 240.244
R13046 gnd.n3907 gnd.n2283 240.244
R13047 gnd.n3907 gnd.n2274 240.244
R13048 gnd.n2274 gnd.n2264 240.244
R13049 gnd.n3933 gnd.n2264 240.244
R13050 gnd.n3933 gnd.n2259 240.244
R13051 gnd.n3965 gnd.n2259 240.244
R13052 gnd.n3965 gnd.n2253 240.244
R13053 gnd.n3938 gnd.n2253 240.244
R13054 gnd.n3938 gnd.n2243 240.244
R13055 gnd.n3939 gnd.n2243 240.244
R13056 gnd.n3940 gnd.n3939 240.244
R13057 gnd.n3940 gnd.n2224 240.244
R13058 gnd.n3943 gnd.n2224 240.244
R13059 gnd.n3943 gnd.n2217 240.244
R13060 gnd.n3946 gnd.n2217 240.244
R13061 gnd.n3946 gnd.n2135 240.244
R13062 gnd.n2135 gnd.n2125 240.244
R13063 gnd.n4167 gnd.n2125 240.244
R13064 gnd.n4167 gnd.n2121 240.244
R13065 gnd.n4173 gnd.n2121 240.244
R13066 gnd.n4173 gnd.n2113 240.244
R13067 gnd.n4186 gnd.n2113 240.244
R13068 gnd.n4186 gnd.n2109 240.244
R13069 gnd.n4192 gnd.n2109 240.244
R13070 gnd.n4192 gnd.n1795 240.244
R13071 gnd.n4568 gnd.n1795 240.244
R13072 gnd.n3051 gnd.n3050 240.244
R13073 gnd.n3034 gnd.n3033 240.244
R13074 gnd.n3059 gnd.n3058 240.244
R13075 gnd.n3061 gnd.n3060 240.244
R13076 gnd.n3068 gnd.n3067 240.244
R13077 gnd.n3070 gnd.n3069 240.244
R13078 gnd.n3080 gnd.n3079 240.244
R13079 gnd.n3088 gnd.n3087 240.244
R13080 gnd.n3090 gnd.n3089 240.244
R13081 gnd.n3100 gnd.n3099 240.244
R13082 gnd.n3108 gnd.n3107 240.244
R13083 gnd.n3110 gnd.n3109 240.244
R13084 gnd.n3122 gnd.n3121 240.244
R13085 gnd.n3327 gnd.n2573 240.244
R13086 gnd.n3338 gnd.n2550 240.244
R13087 gnd.n3338 gnd.n2544 240.244
R13088 gnd.n3361 gnd.n2544 240.244
R13089 gnd.n3361 gnd.n2545 240.244
R13090 gnd.n2545 gnd.n2535 240.244
R13091 gnd.n3343 gnd.n2535 240.244
R13092 gnd.n3344 gnd.n3343 240.244
R13093 gnd.n3347 gnd.n3344 240.244
R13094 gnd.n3348 gnd.n3347 240.244
R13095 gnd.n3348 gnd.n1688 240.244
R13096 gnd.n1699 gnd.n1688 240.244
R13097 gnd.n4678 gnd.n1699 240.244
R13098 gnd.n4678 gnd.n1700 240.244
R13099 gnd.n1705 gnd.n1700 240.244
R13100 gnd.n1706 gnd.n1705 240.244
R13101 gnd.n1707 gnd.n1706 240.244
R13102 gnd.n2499 gnd.n1707 240.244
R13103 gnd.n2499 gnd.n1710 240.244
R13104 gnd.n1711 gnd.n1710 240.244
R13105 gnd.n1712 gnd.n1711 240.244
R13106 gnd.n2474 gnd.n1712 240.244
R13107 gnd.n2474 gnd.n1715 240.244
R13108 gnd.n1716 gnd.n1715 240.244
R13109 gnd.n1717 gnd.n1716 240.244
R13110 gnd.n3586 gnd.n1717 240.244
R13111 gnd.n3586 gnd.n1720 240.244
R13112 gnd.n1721 gnd.n1720 240.244
R13113 gnd.n1722 gnd.n1721 240.244
R13114 gnd.n3643 gnd.n1722 240.244
R13115 gnd.n3643 gnd.n1725 240.244
R13116 gnd.n1726 gnd.n1725 240.244
R13117 gnd.n1727 gnd.n1726 240.244
R13118 gnd.n2402 gnd.n1727 240.244
R13119 gnd.n2402 gnd.n1730 240.244
R13120 gnd.n1731 gnd.n1730 240.244
R13121 gnd.n1732 gnd.n1731 240.244
R13122 gnd.n3672 gnd.n1732 240.244
R13123 gnd.n3672 gnd.n1735 240.244
R13124 gnd.n1736 gnd.n1735 240.244
R13125 gnd.n1737 gnd.n1736 240.244
R13126 gnd.n2364 gnd.n1737 240.244
R13127 gnd.n2364 gnd.n1740 240.244
R13128 gnd.n1741 gnd.n1740 240.244
R13129 gnd.n1742 gnd.n1741 240.244
R13130 gnd.n3755 gnd.n1742 240.244
R13131 gnd.n3755 gnd.n1745 240.244
R13132 gnd.n1746 gnd.n1745 240.244
R13133 gnd.n1747 gnd.n1746 240.244
R13134 gnd.n3827 gnd.n1747 240.244
R13135 gnd.n3827 gnd.n1750 240.244
R13136 gnd.n1751 gnd.n1750 240.244
R13137 gnd.n1752 gnd.n1751 240.244
R13138 gnd.n3888 gnd.n1752 240.244
R13139 gnd.n3888 gnd.n1755 240.244
R13140 gnd.n1756 gnd.n1755 240.244
R13141 gnd.n1757 gnd.n1756 240.244
R13142 gnd.n3908 gnd.n1757 240.244
R13143 gnd.n3908 gnd.n1760 240.244
R13144 gnd.n1761 gnd.n1760 240.244
R13145 gnd.n1762 gnd.n1761 240.244
R13146 gnd.n3853 gnd.n1762 240.244
R13147 gnd.n3853 gnd.n1765 240.244
R13148 gnd.n1766 gnd.n1765 240.244
R13149 gnd.n1767 gnd.n1766 240.244
R13150 gnd.n2245 gnd.n1767 240.244
R13151 gnd.n2245 gnd.n1770 240.244
R13152 gnd.n1771 gnd.n1770 240.244
R13153 gnd.n1772 gnd.n1771 240.244
R13154 gnd.n2226 gnd.n1772 240.244
R13155 gnd.n2226 gnd.n1775 240.244
R13156 gnd.n1776 gnd.n1775 240.244
R13157 gnd.n1777 gnd.n1776 240.244
R13158 gnd.n2137 gnd.n1777 240.244
R13159 gnd.n2137 gnd.n1780 240.244
R13160 gnd.n1781 gnd.n1780 240.244
R13161 gnd.n1782 gnd.n1781 240.244
R13162 gnd.n2114 gnd.n1782 240.244
R13163 gnd.n2114 gnd.n1785 240.244
R13164 gnd.n1786 gnd.n1785 240.244
R13165 gnd.n1787 gnd.n1786 240.244
R13166 gnd.n1790 gnd.n1787 240.244
R13167 gnd.n4570 gnd.n1790 240.244
R13168 gnd.n1801 gnd.n1800 240.244
R13169 gnd.n2080 gnd.n1804 240.244
R13170 gnd.n1806 gnd.n1805 240.244
R13171 gnd.n2083 gnd.n1810 240.244
R13172 gnd.n2086 gnd.n1811 240.244
R13173 gnd.n1820 gnd.n1819 240.244
R13174 gnd.n2088 gnd.n1827 240.244
R13175 gnd.n2091 gnd.n1828 240.244
R13176 gnd.n1836 gnd.n1835 240.244
R13177 gnd.n2093 gnd.n1843 240.244
R13178 gnd.n2096 gnd.n1844 240.244
R13179 gnd.n1852 gnd.n1851 240.244
R13180 gnd.n2099 gnd.n2078 240.244
R13181 gnd.n4253 gnd.n1791 240.244
R13182 gnd.n1668 gnd.n1667 240.132
R13183 gnd.n2153 gnd.n2152 240.132
R13184 gnd.n6746 gnd.n6745 225.874
R13185 gnd.n6746 gnd.n945 225.874
R13186 gnd.n6754 gnd.n945 225.874
R13187 gnd.n6755 gnd.n6754 225.874
R13188 gnd.n6756 gnd.n6755 225.874
R13189 gnd.n6756 gnd.n939 225.874
R13190 gnd.n6764 gnd.n939 225.874
R13191 gnd.n6765 gnd.n6764 225.874
R13192 gnd.n6766 gnd.n6765 225.874
R13193 gnd.n6766 gnd.n933 225.874
R13194 gnd.n6774 gnd.n933 225.874
R13195 gnd.n6775 gnd.n6774 225.874
R13196 gnd.n6776 gnd.n6775 225.874
R13197 gnd.n6776 gnd.n927 225.874
R13198 gnd.n6784 gnd.n927 225.874
R13199 gnd.n6785 gnd.n6784 225.874
R13200 gnd.n6786 gnd.n6785 225.874
R13201 gnd.n6786 gnd.n921 225.874
R13202 gnd.n6794 gnd.n921 225.874
R13203 gnd.n6795 gnd.n6794 225.874
R13204 gnd.n6796 gnd.n6795 225.874
R13205 gnd.n6796 gnd.n915 225.874
R13206 gnd.n6804 gnd.n915 225.874
R13207 gnd.n6805 gnd.n6804 225.874
R13208 gnd.n6806 gnd.n6805 225.874
R13209 gnd.n6806 gnd.n909 225.874
R13210 gnd.n6814 gnd.n909 225.874
R13211 gnd.n6815 gnd.n6814 225.874
R13212 gnd.n6816 gnd.n6815 225.874
R13213 gnd.n6816 gnd.n903 225.874
R13214 gnd.n6824 gnd.n903 225.874
R13215 gnd.n6825 gnd.n6824 225.874
R13216 gnd.n6826 gnd.n6825 225.874
R13217 gnd.n6826 gnd.n897 225.874
R13218 gnd.n6834 gnd.n897 225.874
R13219 gnd.n6835 gnd.n6834 225.874
R13220 gnd.n6836 gnd.n6835 225.874
R13221 gnd.n6836 gnd.n891 225.874
R13222 gnd.n6844 gnd.n891 225.874
R13223 gnd.n6845 gnd.n6844 225.874
R13224 gnd.n6846 gnd.n6845 225.874
R13225 gnd.n6846 gnd.n885 225.874
R13226 gnd.n6854 gnd.n885 225.874
R13227 gnd.n6855 gnd.n6854 225.874
R13228 gnd.n6856 gnd.n6855 225.874
R13229 gnd.n6856 gnd.n879 225.874
R13230 gnd.n6864 gnd.n879 225.874
R13231 gnd.n6865 gnd.n6864 225.874
R13232 gnd.n6866 gnd.n6865 225.874
R13233 gnd.n6866 gnd.n873 225.874
R13234 gnd.n6874 gnd.n873 225.874
R13235 gnd.n6875 gnd.n6874 225.874
R13236 gnd.n6876 gnd.n6875 225.874
R13237 gnd.n6876 gnd.n867 225.874
R13238 gnd.n6884 gnd.n867 225.874
R13239 gnd.n6885 gnd.n6884 225.874
R13240 gnd.n6886 gnd.n6885 225.874
R13241 gnd.n6886 gnd.n861 225.874
R13242 gnd.n6894 gnd.n861 225.874
R13243 gnd.n6895 gnd.n6894 225.874
R13244 gnd.n6896 gnd.n6895 225.874
R13245 gnd.n6896 gnd.n855 225.874
R13246 gnd.n6904 gnd.n855 225.874
R13247 gnd.n6905 gnd.n6904 225.874
R13248 gnd.n6906 gnd.n6905 225.874
R13249 gnd.n6906 gnd.n849 225.874
R13250 gnd.n6914 gnd.n849 225.874
R13251 gnd.n6915 gnd.n6914 225.874
R13252 gnd.n6916 gnd.n6915 225.874
R13253 gnd.n6916 gnd.n843 225.874
R13254 gnd.n6924 gnd.n843 225.874
R13255 gnd.n6925 gnd.n6924 225.874
R13256 gnd.n6926 gnd.n6925 225.874
R13257 gnd.n6926 gnd.n837 225.874
R13258 gnd.n6934 gnd.n837 225.874
R13259 gnd.n6935 gnd.n6934 225.874
R13260 gnd.n6936 gnd.n6935 225.874
R13261 gnd.n6936 gnd.n831 225.874
R13262 gnd.n6944 gnd.n831 225.874
R13263 gnd.n6945 gnd.n6944 225.874
R13264 gnd.n6946 gnd.n6945 225.874
R13265 gnd.n6946 gnd.n825 225.874
R13266 gnd.n6954 gnd.n825 225.874
R13267 gnd.n6955 gnd.n6954 225.874
R13268 gnd.n6956 gnd.n6955 225.874
R13269 gnd.n6956 gnd.n819 225.874
R13270 gnd.n6964 gnd.n819 225.874
R13271 gnd.n6965 gnd.n6964 225.874
R13272 gnd.n6966 gnd.n6965 225.874
R13273 gnd.n6966 gnd.n813 225.874
R13274 gnd.n6974 gnd.n813 225.874
R13275 gnd.n6975 gnd.n6974 225.874
R13276 gnd.n6976 gnd.n6975 225.874
R13277 gnd.n6976 gnd.n807 225.874
R13278 gnd.n6984 gnd.n807 225.874
R13279 gnd.n6985 gnd.n6984 225.874
R13280 gnd.n6986 gnd.n6985 225.874
R13281 gnd.n6986 gnd.n801 225.874
R13282 gnd.n6994 gnd.n801 225.874
R13283 gnd.n6995 gnd.n6994 225.874
R13284 gnd.n6996 gnd.n6995 225.874
R13285 gnd.n6996 gnd.n795 225.874
R13286 gnd.n7004 gnd.n795 225.874
R13287 gnd.n7005 gnd.n7004 225.874
R13288 gnd.n7006 gnd.n7005 225.874
R13289 gnd.n7006 gnd.n789 225.874
R13290 gnd.n7014 gnd.n789 225.874
R13291 gnd.n7015 gnd.n7014 225.874
R13292 gnd.n7016 gnd.n7015 225.874
R13293 gnd.n7016 gnd.n783 225.874
R13294 gnd.n7024 gnd.n783 225.874
R13295 gnd.n7025 gnd.n7024 225.874
R13296 gnd.n7026 gnd.n7025 225.874
R13297 gnd.n7026 gnd.n777 225.874
R13298 gnd.n7034 gnd.n777 225.874
R13299 gnd.n7035 gnd.n7034 225.874
R13300 gnd.n7036 gnd.n7035 225.874
R13301 gnd.n7036 gnd.n771 225.874
R13302 gnd.n7044 gnd.n771 225.874
R13303 gnd.n7045 gnd.n7044 225.874
R13304 gnd.n7046 gnd.n7045 225.874
R13305 gnd.n7046 gnd.n765 225.874
R13306 gnd.n7054 gnd.n765 225.874
R13307 gnd.n7055 gnd.n7054 225.874
R13308 gnd.n7056 gnd.n7055 225.874
R13309 gnd.n7056 gnd.n759 225.874
R13310 gnd.n7064 gnd.n759 225.874
R13311 gnd.n7065 gnd.n7064 225.874
R13312 gnd.n7066 gnd.n7065 225.874
R13313 gnd.n7066 gnd.n753 225.874
R13314 gnd.n7074 gnd.n753 225.874
R13315 gnd.n7075 gnd.n7074 225.874
R13316 gnd.n7076 gnd.n7075 225.874
R13317 gnd.n7076 gnd.n747 225.874
R13318 gnd.n7084 gnd.n747 225.874
R13319 gnd.n7085 gnd.n7084 225.874
R13320 gnd.n7086 gnd.n7085 225.874
R13321 gnd.n7086 gnd.n741 225.874
R13322 gnd.n7094 gnd.n741 225.874
R13323 gnd.n7095 gnd.n7094 225.874
R13324 gnd.n7096 gnd.n7095 225.874
R13325 gnd.n7096 gnd.n735 225.874
R13326 gnd.n7104 gnd.n735 225.874
R13327 gnd.n7105 gnd.n7104 225.874
R13328 gnd.n7106 gnd.n7105 225.874
R13329 gnd.n7106 gnd.n729 225.874
R13330 gnd.n7114 gnd.n729 225.874
R13331 gnd.n7115 gnd.n7114 225.874
R13332 gnd.n7116 gnd.n7115 225.874
R13333 gnd.n7116 gnd.n723 225.874
R13334 gnd.n7125 gnd.n723 225.874
R13335 gnd.n7126 gnd.n7125 225.874
R13336 gnd.n7127 gnd.n7126 225.874
R13337 gnd.n7127 gnd.n718 225.874
R13338 gnd.n5558 gnd.t288 224.174
R13339 gnd.n6494 gnd.t394 224.174
R13340 gnd.n1936 gnd.n1873 199.319
R13341 gnd.n1936 gnd.n1874 199.319
R13342 gnd.n1620 gnd.n1580 199.319
R13343 gnd.n1620 gnd.n1579 199.319
R13344 gnd.n1669 gnd.n1666 186.49
R13345 gnd.n2154 gnd.n2151 186.49
R13346 gnd.n6384 gnd.n6383 185
R13347 gnd.n6382 gnd.n6381 185
R13348 gnd.n6361 gnd.n6360 185
R13349 gnd.n6376 gnd.n6375 185
R13350 gnd.n6374 gnd.n6373 185
R13351 gnd.n6365 gnd.n6364 185
R13352 gnd.n6368 gnd.n6367 185
R13353 gnd.n6352 gnd.n6351 185
R13354 gnd.n6350 gnd.n6349 185
R13355 gnd.n6329 gnd.n6328 185
R13356 gnd.n6344 gnd.n6343 185
R13357 gnd.n6342 gnd.n6341 185
R13358 gnd.n6333 gnd.n6332 185
R13359 gnd.n6336 gnd.n6335 185
R13360 gnd.n6320 gnd.n6319 185
R13361 gnd.n6318 gnd.n6317 185
R13362 gnd.n6297 gnd.n6296 185
R13363 gnd.n6312 gnd.n6311 185
R13364 gnd.n6310 gnd.n6309 185
R13365 gnd.n6301 gnd.n6300 185
R13366 gnd.n6304 gnd.n6303 185
R13367 gnd.n6289 gnd.n6288 185
R13368 gnd.n6287 gnd.n6286 185
R13369 gnd.n6266 gnd.n6265 185
R13370 gnd.n6281 gnd.n6280 185
R13371 gnd.n6279 gnd.n6278 185
R13372 gnd.n6270 gnd.n6269 185
R13373 gnd.n6273 gnd.n6272 185
R13374 gnd.n6257 gnd.n6256 185
R13375 gnd.n6255 gnd.n6254 185
R13376 gnd.n6234 gnd.n6233 185
R13377 gnd.n6249 gnd.n6248 185
R13378 gnd.n6247 gnd.n6246 185
R13379 gnd.n6238 gnd.n6237 185
R13380 gnd.n6241 gnd.n6240 185
R13381 gnd.n6225 gnd.n6224 185
R13382 gnd.n6223 gnd.n6222 185
R13383 gnd.n6202 gnd.n6201 185
R13384 gnd.n6217 gnd.n6216 185
R13385 gnd.n6215 gnd.n6214 185
R13386 gnd.n6206 gnd.n6205 185
R13387 gnd.n6209 gnd.n6208 185
R13388 gnd.n6193 gnd.n6192 185
R13389 gnd.n6191 gnd.n6190 185
R13390 gnd.n6170 gnd.n6169 185
R13391 gnd.n6185 gnd.n6184 185
R13392 gnd.n6183 gnd.n6182 185
R13393 gnd.n6174 gnd.n6173 185
R13394 gnd.n6177 gnd.n6176 185
R13395 gnd.n6162 gnd.n6161 185
R13396 gnd.n6160 gnd.n6159 185
R13397 gnd.n6139 gnd.n6138 185
R13398 gnd.n6154 gnd.n6153 185
R13399 gnd.n6152 gnd.n6151 185
R13400 gnd.n6143 gnd.n6142 185
R13401 gnd.n6146 gnd.n6145 185
R13402 gnd.n5559 gnd.t287 178.987
R13403 gnd.n6495 gnd.t395 178.987
R13404 gnd.n1 gnd.t50 170.774
R13405 gnd.n7 gnd.t262 170.103
R13406 gnd.n6 gnd.t56 170.103
R13407 gnd.n5 gnd.t149 170.103
R13408 gnd.n4 gnd.t81 170.103
R13409 gnd.n3 gnd.t94 170.103
R13410 gnd.n2 gnd.t169 170.103
R13411 gnd.n1 gnd.t88 170.103
R13412 gnd.n4149 gnd.n4148 163.367
R13413 gnd.n4146 gnd.n2163 163.367
R13414 gnd.n4142 gnd.n4141 163.367
R13415 gnd.n4139 gnd.n2166 163.367
R13416 gnd.n4135 gnd.n4134 163.367
R13417 gnd.n4132 gnd.n2169 163.367
R13418 gnd.n4128 gnd.n4127 163.367
R13419 gnd.n4125 gnd.n2172 163.367
R13420 gnd.n4121 gnd.n4120 163.367
R13421 gnd.n4118 gnd.n2175 163.367
R13422 gnd.n4114 gnd.n4113 163.367
R13423 gnd.n4111 gnd.n2178 163.367
R13424 gnd.n4107 gnd.n4106 163.367
R13425 gnd.n4104 gnd.n2181 163.367
R13426 gnd.n4099 gnd.n4098 163.367
R13427 gnd.n4096 gnd.n4094 163.367
R13428 gnd.n4091 gnd.n4090 163.367
R13429 gnd.n4088 gnd.n2187 163.367
R13430 gnd.n4083 gnd.n4082 163.367
R13431 gnd.n4080 gnd.n2192 163.367
R13432 gnd.n4076 gnd.n4075 163.367
R13433 gnd.n4073 gnd.n2195 163.367
R13434 gnd.n4069 gnd.n4068 163.367
R13435 gnd.n4066 gnd.n2198 163.367
R13436 gnd.n4062 gnd.n4061 163.367
R13437 gnd.n4059 gnd.n2201 163.367
R13438 gnd.n4055 gnd.n4054 163.367
R13439 gnd.n4052 gnd.n2204 163.367
R13440 gnd.n4048 gnd.n4047 163.367
R13441 gnd.n4045 gnd.n2207 163.367
R13442 gnd.n4041 gnd.n4040 163.367
R13443 gnd.n4038 gnd.n2210 163.367
R13444 gnd.n3473 gnd.n1685 163.367
R13445 gnd.n3476 gnd.n1685 163.367
R13446 gnd.n3476 gnd.n3406 163.367
R13447 gnd.n3480 gnd.n3406 163.367
R13448 gnd.n3480 gnd.n2518 163.367
R13449 gnd.n3488 gnd.n2518 163.367
R13450 gnd.n3488 gnd.n2515 163.367
R13451 gnd.n3515 gnd.n2515 163.367
R13452 gnd.n3515 gnd.n2516 163.367
R13453 gnd.n2516 gnd.n2509 163.367
R13454 gnd.n3510 gnd.n2509 163.367
R13455 gnd.n3510 gnd.n3507 163.367
R13456 gnd.n3507 gnd.n3506 163.367
R13457 gnd.n3506 gnd.n3494 163.367
R13458 gnd.n3494 gnd.n2490 163.367
R13459 gnd.n3501 gnd.n2490 163.367
R13460 gnd.n3501 gnd.n2486 163.367
R13461 gnd.n3498 gnd.n2486 163.367
R13462 gnd.n3498 gnd.n2476 163.367
R13463 gnd.n2476 gnd.n2469 163.367
R13464 gnd.n3581 gnd.n2469 163.367
R13465 gnd.n3582 gnd.n3581 163.367
R13466 gnd.n3582 gnd.n2458 163.367
R13467 gnd.n3589 gnd.n2458 163.367
R13468 gnd.n3590 gnd.n3589 163.367
R13469 gnd.n3590 gnd.n2467 163.367
R13470 gnd.n3594 gnd.n2467 163.367
R13471 gnd.n3594 gnd.n2440 163.367
R13472 gnd.n3625 gnd.n2440 163.367
R13473 gnd.n3625 gnd.n2429 163.367
R13474 gnd.n2437 gnd.n2429 163.367
R13475 gnd.n3635 gnd.n2437 163.367
R13476 gnd.n3635 gnd.n2438 163.367
R13477 gnd.n3631 gnd.n2438 163.367
R13478 gnd.n3631 gnd.n2400 163.367
R13479 gnd.n2400 gnd.n2392 163.367
R13480 gnd.n3689 gnd.n2392 163.367
R13481 gnd.n3689 gnd.n2390 163.367
R13482 gnd.n3694 gnd.n2390 163.367
R13483 gnd.n3694 gnd.n2384 163.367
R13484 gnd.n3703 gnd.n2384 163.367
R13485 gnd.n3704 gnd.n3703 163.367
R13486 gnd.n3704 gnd.n2381 163.367
R13487 gnd.n3724 gnd.n2381 163.367
R13488 gnd.n3724 gnd.n2373 163.367
R13489 gnd.n3720 gnd.n2373 163.367
R13490 gnd.n3720 gnd.n3719 163.367
R13491 gnd.n3719 gnd.n3718 163.367
R13492 gnd.n3718 gnd.n3708 163.367
R13493 gnd.n3708 gnd.n2355 163.367
R13494 gnd.n3713 gnd.n2355 163.367
R13495 gnd.n3713 gnd.n2349 163.367
R13496 gnd.n3710 gnd.n2349 163.367
R13497 gnd.n3710 gnd.n2339 163.367
R13498 gnd.n2339 gnd.n2332 163.367
R13499 gnd.n3809 gnd.n2332 163.367
R13500 gnd.n3809 gnd.n2329 163.367
R13501 gnd.n3819 gnd.n2329 163.367
R13502 gnd.n3819 gnd.n2330 163.367
R13503 gnd.n2330 gnd.n2323 163.367
R13504 gnd.n3814 gnd.n2323 163.367
R13505 gnd.n3814 gnd.n2313 163.367
R13506 gnd.n2313 gnd.n2307 163.367
R13507 gnd.n3844 gnd.n2307 163.367
R13508 gnd.n3845 gnd.n3844 163.367
R13509 gnd.n3845 gnd.n2298 163.367
R13510 gnd.n3849 gnd.n2298 163.367
R13511 gnd.n3849 gnd.n2304 163.367
R13512 gnd.n3878 gnd.n2304 163.367
R13513 gnd.n3878 gnd.n2305 163.367
R13514 gnd.n2305 gnd.n2282 163.367
R13515 gnd.n3873 gnd.n2282 163.367
R13516 gnd.n3873 gnd.n2275 163.367
R13517 gnd.n3870 gnd.n2275 163.367
R13518 gnd.n3870 gnd.n3868 163.367
R13519 gnd.n3868 gnd.n3867 163.367
R13520 gnd.n3867 gnd.n3856 163.367
R13521 gnd.n3856 gnd.n2258 163.367
R13522 gnd.n3862 gnd.n2258 163.367
R13523 gnd.n3862 gnd.n2254 163.367
R13524 gnd.n3859 gnd.n2254 163.367
R13525 gnd.n3859 gnd.n2242 163.367
R13526 gnd.n2242 gnd.n2235 163.367
R13527 gnd.n3992 gnd.n2235 163.367
R13528 gnd.n3992 gnd.n2232 163.367
R13529 gnd.n4003 gnd.n2232 163.367
R13530 gnd.n4003 gnd.n2233 163.367
R13531 gnd.n2233 gnd.n2225 163.367
R13532 gnd.n3998 gnd.n2225 163.367
R13533 gnd.n3998 gnd.n2216 163.367
R13534 gnd.n2216 gnd.n2212 163.367
R13535 gnd.n4027 gnd.n2212 163.367
R13536 gnd.n4028 gnd.n4027 163.367
R13537 gnd.n4028 gnd.n2136 163.367
R13538 gnd.n4033 gnd.n2136 163.367
R13539 gnd.n1660 gnd.n1659 163.367
R13540 gnd.n4749 gnd.n1659 163.367
R13541 gnd.n4747 gnd.n4746 163.367
R13542 gnd.n4743 gnd.n4742 163.367
R13543 gnd.n4739 gnd.n4738 163.367
R13544 gnd.n4735 gnd.n4734 163.367
R13545 gnd.n4731 gnd.n4730 163.367
R13546 gnd.n4727 gnd.n4726 163.367
R13547 gnd.n4723 gnd.n4722 163.367
R13548 gnd.n4719 gnd.n4718 163.367
R13549 gnd.n4715 gnd.n4714 163.367
R13550 gnd.n4711 gnd.n4710 163.367
R13551 gnd.n4707 gnd.n4706 163.367
R13552 gnd.n4703 gnd.n4702 163.367
R13553 gnd.n4699 gnd.n4698 163.367
R13554 gnd.n4695 gnd.n4694 163.367
R13555 gnd.n4758 gnd.n1625 163.367
R13556 gnd.n3411 gnd.n3410 163.367
R13557 gnd.n3416 gnd.n3415 163.367
R13558 gnd.n3420 gnd.n3419 163.367
R13559 gnd.n3424 gnd.n3423 163.367
R13560 gnd.n3428 gnd.n3427 163.367
R13561 gnd.n3432 gnd.n3431 163.367
R13562 gnd.n3436 gnd.n3435 163.367
R13563 gnd.n3440 gnd.n3439 163.367
R13564 gnd.n3444 gnd.n3443 163.367
R13565 gnd.n3448 gnd.n3447 163.367
R13566 gnd.n3452 gnd.n3451 163.367
R13567 gnd.n3456 gnd.n3455 163.367
R13568 gnd.n3460 gnd.n3459 163.367
R13569 gnd.n3464 gnd.n3463 163.367
R13570 gnd.n3468 gnd.n3467 163.367
R13571 gnd.n4687 gnd.n1661 163.367
R13572 gnd.n4687 gnd.n1683 163.367
R13573 gnd.n2523 gnd.n1683 163.367
R13574 gnd.n3482 gnd.n2523 163.367
R13575 gnd.n3482 gnd.n2521 163.367
R13576 gnd.n3486 gnd.n2521 163.367
R13577 gnd.n3486 gnd.n2513 163.367
R13578 gnd.n3517 gnd.n2513 163.367
R13579 gnd.n3517 gnd.n2510 163.367
R13580 gnd.n3526 gnd.n2510 163.367
R13581 gnd.n3526 gnd.n2511 163.367
R13582 gnd.n3522 gnd.n2511 163.367
R13583 gnd.n3522 gnd.n3521 163.367
R13584 gnd.n3521 gnd.n2489 163.367
R13585 gnd.n3559 gnd.n2489 163.367
R13586 gnd.n3559 gnd.n2487 163.367
R13587 gnd.n3563 gnd.n2487 163.367
R13588 gnd.n3563 gnd.n2473 163.367
R13589 gnd.n3575 gnd.n2473 163.367
R13590 gnd.n3575 gnd.n2471 163.367
R13591 gnd.n3579 gnd.n2471 163.367
R13592 gnd.n3579 gnd.n2459 163.367
R13593 gnd.n3602 gnd.n2459 163.367
R13594 gnd.n3602 gnd.n2460 163.367
R13595 gnd.n3598 gnd.n2460 163.367
R13596 gnd.n3598 gnd.n3597 163.367
R13597 gnd.n3597 gnd.n3596 163.367
R13598 gnd.n3596 gnd.n2463 163.367
R13599 gnd.n2463 gnd.n2430 163.367
R13600 gnd.n3641 gnd.n2430 163.367
R13601 gnd.n3641 gnd.n2431 163.367
R13602 gnd.n3637 gnd.n2431 163.367
R13603 gnd.n3637 gnd.n2434 163.367
R13604 gnd.n2434 gnd.n2398 163.367
R13605 gnd.n3683 gnd.n2398 163.367
R13606 gnd.n3683 gnd.n2396 163.367
R13607 gnd.n3687 gnd.n2396 163.367
R13608 gnd.n3687 gnd.n2388 163.367
R13609 gnd.n3697 gnd.n2388 163.367
R13610 gnd.n3697 gnd.n2386 163.367
R13611 gnd.n3701 gnd.n2386 163.367
R13612 gnd.n3701 gnd.n2379 163.367
R13613 gnd.n3728 gnd.n2379 163.367
R13614 gnd.n3728 gnd.n2376 163.367
R13615 gnd.n3737 gnd.n2376 163.367
R13616 gnd.n3737 gnd.n2377 163.367
R13617 gnd.n3733 gnd.n2377 163.367
R13618 gnd.n3733 gnd.n3732 163.367
R13619 gnd.n3732 gnd.n2353 163.367
R13620 gnd.n3785 gnd.n2353 163.367
R13621 gnd.n3785 gnd.n2351 163.367
R13622 gnd.n3789 gnd.n2351 163.367
R13623 gnd.n3789 gnd.n2338 163.367
R13624 gnd.n3803 gnd.n2338 163.367
R13625 gnd.n3803 gnd.n2336 163.367
R13626 gnd.n3807 gnd.n2336 163.367
R13627 gnd.n3807 gnd.n2327 163.367
R13628 gnd.n3821 gnd.n2327 163.367
R13629 gnd.n3821 gnd.n2325 163.367
R13630 gnd.n3825 gnd.n2325 163.367
R13631 gnd.n3825 gnd.n2311 163.367
R13632 gnd.n3838 gnd.n2311 163.367
R13633 gnd.n3838 gnd.n2309 163.367
R13634 gnd.n3842 gnd.n2309 163.367
R13635 gnd.n3842 gnd.n2300 163.367
R13636 gnd.n3886 gnd.n2300 163.367
R13637 gnd.n3886 gnd.n2301 163.367
R13638 gnd.n3882 gnd.n2301 163.367
R13639 gnd.n3882 gnd.n3881 163.367
R13640 gnd.n3881 gnd.n2280 163.367
R13641 gnd.n3911 gnd.n2280 163.367
R13642 gnd.n3911 gnd.n2277 163.367
R13643 gnd.n3920 gnd.n2277 163.367
R13644 gnd.n3920 gnd.n2278 163.367
R13645 gnd.n3916 gnd.n2278 163.367
R13646 gnd.n3916 gnd.n3915 163.367
R13647 gnd.n3915 gnd.n2257 163.367
R13648 gnd.n3968 gnd.n2257 163.367
R13649 gnd.n3968 gnd.n2255 163.367
R13650 gnd.n3972 gnd.n2255 163.367
R13651 gnd.n3972 gnd.n2240 163.367
R13652 gnd.n3986 gnd.n2240 163.367
R13653 gnd.n3986 gnd.n2238 163.367
R13654 gnd.n3990 gnd.n2238 163.367
R13655 gnd.n3990 gnd.n2230 163.367
R13656 gnd.n4005 gnd.n2230 163.367
R13657 gnd.n4005 gnd.n2228 163.367
R13658 gnd.n4009 gnd.n2228 163.367
R13659 gnd.n4009 gnd.n2215 163.367
R13660 gnd.n4021 gnd.n2215 163.367
R13661 gnd.n4021 gnd.n2213 163.367
R13662 gnd.n4025 gnd.n2213 163.367
R13663 gnd.n4025 gnd.n2139 163.367
R13664 gnd.n4156 gnd.n2139 163.367
R13665 gnd.n4156 gnd.n2140 163.367
R13666 gnd.n2160 gnd.n2159 156.462
R13667 gnd.n6324 gnd.n6292 153.042
R13668 gnd.n6388 gnd.n6387 152.079
R13669 gnd.n6356 gnd.n6355 152.079
R13670 gnd.n6324 gnd.n6323 152.079
R13671 gnd.n1674 gnd.n1673 152
R13672 gnd.n1675 gnd.n1664 152
R13673 gnd.n1677 gnd.n1676 152
R13674 gnd.n1679 gnd.n1662 152
R13675 gnd.n1681 gnd.n1680 152
R13676 gnd.n2158 gnd.n2142 152
R13677 gnd.n2150 gnd.n2143 152
R13678 gnd.n2149 gnd.n2148 152
R13679 gnd.n2147 gnd.n2144 152
R13680 gnd.n2145 gnd.t300 150.546
R13681 gnd.t219 gnd.n6366 147.661
R13682 gnd.t280 gnd.n6334 147.661
R13683 gnd.t164 gnd.n6302 147.661
R13684 gnd.t208 gnd.n6271 147.661
R13685 gnd.t243 gnd.n6239 147.661
R13686 gnd.t187 gnd.n6207 147.661
R13687 gnd.t90 gnd.n6175 147.661
R13688 gnd.t271 gnd.n6144 147.661
R13689 gnd.n4093 gnd.n4092 143.351
R13690 gnd.n1641 gnd.n1624 143.351
R13691 gnd.n4757 gnd.n1624 143.351
R13692 gnd.n1671 gnd.t352 130.484
R13693 gnd.n1680 gnd.t377 126.766
R13694 gnd.n1678 gnd.t289 126.766
R13695 gnd.n1664 gnd.t361 126.766
R13696 gnd.n1672 gnd.t328 126.766
R13697 gnd.n2146 gnd.t282 126.766
R13698 gnd.n2148 gnd.t396 126.766
R13699 gnd.n2157 gnd.t342 126.766
R13700 gnd.n2159 gnd.t322 126.766
R13701 gnd.n6383 gnd.n6382 104.615
R13702 gnd.n6382 gnd.n6360 104.615
R13703 gnd.n6375 gnd.n6360 104.615
R13704 gnd.n6375 gnd.n6374 104.615
R13705 gnd.n6374 gnd.n6364 104.615
R13706 gnd.n6367 gnd.n6364 104.615
R13707 gnd.n6351 gnd.n6350 104.615
R13708 gnd.n6350 gnd.n6328 104.615
R13709 gnd.n6343 gnd.n6328 104.615
R13710 gnd.n6343 gnd.n6342 104.615
R13711 gnd.n6342 gnd.n6332 104.615
R13712 gnd.n6335 gnd.n6332 104.615
R13713 gnd.n6319 gnd.n6318 104.615
R13714 gnd.n6318 gnd.n6296 104.615
R13715 gnd.n6311 gnd.n6296 104.615
R13716 gnd.n6311 gnd.n6310 104.615
R13717 gnd.n6310 gnd.n6300 104.615
R13718 gnd.n6303 gnd.n6300 104.615
R13719 gnd.n6288 gnd.n6287 104.615
R13720 gnd.n6287 gnd.n6265 104.615
R13721 gnd.n6280 gnd.n6265 104.615
R13722 gnd.n6280 gnd.n6279 104.615
R13723 gnd.n6279 gnd.n6269 104.615
R13724 gnd.n6272 gnd.n6269 104.615
R13725 gnd.n6256 gnd.n6255 104.615
R13726 gnd.n6255 gnd.n6233 104.615
R13727 gnd.n6248 gnd.n6233 104.615
R13728 gnd.n6248 gnd.n6247 104.615
R13729 gnd.n6247 gnd.n6237 104.615
R13730 gnd.n6240 gnd.n6237 104.615
R13731 gnd.n6224 gnd.n6223 104.615
R13732 gnd.n6223 gnd.n6201 104.615
R13733 gnd.n6216 gnd.n6201 104.615
R13734 gnd.n6216 gnd.n6215 104.615
R13735 gnd.n6215 gnd.n6205 104.615
R13736 gnd.n6208 gnd.n6205 104.615
R13737 gnd.n6192 gnd.n6191 104.615
R13738 gnd.n6191 gnd.n6169 104.615
R13739 gnd.n6184 gnd.n6169 104.615
R13740 gnd.n6184 gnd.n6183 104.615
R13741 gnd.n6183 gnd.n6173 104.615
R13742 gnd.n6176 gnd.n6173 104.615
R13743 gnd.n6161 gnd.n6160 104.615
R13744 gnd.n6160 gnd.n6138 104.615
R13745 gnd.n6153 gnd.n6138 104.615
R13746 gnd.n6153 gnd.n6152 104.615
R13747 gnd.n6152 gnd.n6142 104.615
R13748 gnd.n6145 gnd.n6142 104.615
R13749 gnd.n5708 gnd.t334 100.632
R13750 gnd.n1129 gnd.t369 100.632
R13751 gnd.n7662 gnd.n7661 99.6594
R13752 gnd.n7657 gnd.n288 99.6594
R13753 gnd.n7653 gnd.n287 99.6594
R13754 gnd.n7649 gnd.n286 99.6594
R13755 gnd.n7645 gnd.n285 99.6594
R13756 gnd.n7641 gnd.n284 99.6594
R13757 gnd.n7637 gnd.n283 99.6594
R13758 gnd.n7633 gnd.n282 99.6594
R13759 gnd.n7626 gnd.n281 99.6594
R13760 gnd.n7622 gnd.n280 99.6594
R13761 gnd.n7618 gnd.n279 99.6594
R13762 gnd.n7614 gnd.n278 99.6594
R13763 gnd.n7610 gnd.n277 99.6594
R13764 gnd.n7606 gnd.n276 99.6594
R13765 gnd.n7602 gnd.n275 99.6594
R13766 gnd.n7598 gnd.n274 99.6594
R13767 gnd.n7594 gnd.n273 99.6594
R13768 gnd.n7590 gnd.n272 99.6594
R13769 gnd.n7582 gnd.n271 99.6594
R13770 gnd.n7580 gnd.n270 99.6594
R13771 gnd.n7576 gnd.n269 99.6594
R13772 gnd.n7572 gnd.n268 99.6594
R13773 gnd.n7568 gnd.n267 99.6594
R13774 gnd.n7564 gnd.n266 99.6594
R13775 gnd.n7560 gnd.n265 99.6594
R13776 gnd.n7556 gnd.n264 99.6594
R13777 gnd.n7552 gnd.n263 99.6594
R13778 gnd.n7548 gnd.n262 99.6594
R13779 gnd.n7539 gnd.n261 99.6594
R13780 gnd.n4500 gnd.n4499 99.6594
R13781 gnd.n4494 gnd.n1862 99.6594
R13782 gnd.n4491 gnd.n1863 99.6594
R13783 gnd.n4487 gnd.n1864 99.6594
R13784 gnd.n4483 gnd.n1865 99.6594
R13785 gnd.n4479 gnd.n1866 99.6594
R13786 gnd.n4475 gnd.n1867 99.6594
R13787 gnd.n4471 gnd.n1868 99.6594
R13788 gnd.n4467 gnd.n1869 99.6594
R13789 gnd.n4462 gnd.n1870 99.6594
R13790 gnd.n4458 gnd.n1871 99.6594
R13791 gnd.n4454 gnd.n1872 99.6594
R13792 gnd.n4450 gnd.n1873 99.6594
R13793 gnd.n4445 gnd.n1875 99.6594
R13794 gnd.n4441 gnd.n1876 99.6594
R13795 gnd.n4437 gnd.n1877 99.6594
R13796 gnd.n4433 gnd.n1878 99.6594
R13797 gnd.n4429 gnd.n1879 99.6594
R13798 gnd.n4425 gnd.n1880 99.6594
R13799 gnd.n4421 gnd.n1881 99.6594
R13800 gnd.n4417 gnd.n1882 99.6594
R13801 gnd.n4413 gnd.n1883 99.6594
R13802 gnd.n4409 gnd.n1884 99.6594
R13803 gnd.n4405 gnd.n1885 99.6594
R13804 gnd.n4401 gnd.n1886 99.6594
R13805 gnd.n4397 gnd.n1887 99.6594
R13806 gnd.n4393 gnd.n1888 99.6594
R13807 gnd.n4389 gnd.n1889 99.6594
R13808 gnd.n4809 gnd.n4808 99.6594
R13809 gnd.n4804 gnd.n1591 99.6594
R13810 gnd.n4800 gnd.n1590 99.6594
R13811 gnd.n4796 gnd.n1589 99.6594
R13812 gnd.n4792 gnd.n1588 99.6594
R13813 gnd.n4788 gnd.n1587 99.6594
R13814 gnd.n4784 gnd.n1586 99.6594
R13815 gnd.n4780 gnd.n1585 99.6594
R13816 gnd.n4775 gnd.n1584 99.6594
R13817 gnd.n4771 gnd.n1583 99.6594
R13818 gnd.n4767 gnd.n1582 99.6594
R13819 gnd.n4763 gnd.n1581 99.6594
R13820 gnd.n3198 gnd.n1579 99.6594
R13821 gnd.n3202 gnd.n1578 99.6594
R13822 gnd.n3208 gnd.n1577 99.6594
R13823 gnd.n3212 gnd.n1576 99.6594
R13824 gnd.n3217 gnd.n1575 99.6594
R13825 gnd.n3221 gnd.n1574 99.6594
R13826 gnd.n3227 gnd.n1573 99.6594
R13827 gnd.n3231 gnd.n1572 99.6594
R13828 gnd.n3237 gnd.n1571 99.6594
R13829 gnd.n3241 gnd.n1570 99.6594
R13830 gnd.n3247 gnd.n1569 99.6594
R13831 gnd.n3251 gnd.n1568 99.6594
R13832 gnd.n3257 gnd.n1567 99.6594
R13833 gnd.n3261 gnd.n1566 99.6594
R13834 gnd.n3266 gnd.n1565 99.6594
R13835 gnd.n3269 gnd.n1564 99.6594
R13836 gnd.n5110 gnd.n5109 99.6594
R13837 gnd.n5104 gnd.n1148 99.6594
R13838 gnd.n5101 gnd.n1149 99.6594
R13839 gnd.n5097 gnd.n1150 99.6594
R13840 gnd.n5093 gnd.n1151 99.6594
R13841 gnd.n5089 gnd.n1152 99.6594
R13842 gnd.n5085 gnd.n1153 99.6594
R13843 gnd.n5081 gnd.n1154 99.6594
R13844 gnd.n5077 gnd.n1155 99.6594
R13845 gnd.n5072 gnd.n1156 99.6594
R13846 gnd.n5068 gnd.n1157 99.6594
R13847 gnd.n5064 gnd.n1158 99.6594
R13848 gnd.n5060 gnd.n1159 99.6594
R13849 gnd.n5056 gnd.n1160 99.6594
R13850 gnd.n5052 gnd.n1161 99.6594
R13851 gnd.n5048 gnd.n1162 99.6594
R13852 gnd.n5044 gnd.n1163 99.6594
R13853 gnd.n5040 gnd.n1164 99.6594
R13854 gnd.n5036 gnd.n1165 99.6594
R13855 gnd.n5032 gnd.n1166 99.6594
R13856 gnd.n5028 gnd.n1167 99.6594
R13857 gnd.n5024 gnd.n1168 99.6594
R13858 gnd.n5020 gnd.n1169 99.6594
R13859 gnd.n5016 gnd.n1170 99.6594
R13860 gnd.n5012 gnd.n1171 99.6594
R13861 gnd.n5008 gnd.n1172 99.6594
R13862 gnd.n5004 gnd.n1173 99.6594
R13863 gnd.n5000 gnd.n1174 99.6594
R13864 gnd.n4996 gnd.n1175 99.6594
R13865 gnd.n6550 gnd.n5117 99.6594
R13866 gnd.n6548 gnd.n5116 99.6594
R13867 gnd.n6544 gnd.n5115 99.6594
R13868 gnd.n6540 gnd.n5114 99.6594
R13869 gnd.n6536 gnd.n5113 99.6594
R13870 gnd.n6532 gnd.n5112 99.6594
R13871 gnd.n6562 gnd.n6560 99.6594
R13872 gnd.n6568 gnd.n1128 99.6594
R13873 gnd.n5741 gnd.n5740 99.6594
R13874 gnd.n5735 gnd.n5683 99.6594
R13875 gnd.n5732 gnd.n5684 99.6594
R13876 gnd.n5728 gnd.n5685 99.6594
R13877 gnd.n5724 gnd.n5686 99.6594
R13878 gnd.n5720 gnd.n5687 99.6594
R13879 gnd.n5716 gnd.n5688 99.6594
R13880 gnd.n5712 gnd.n5689 99.6594
R13881 gnd.n475 gnd.n252 99.6594
R13882 gnd.n471 gnd.n253 99.6594
R13883 gnd.n467 gnd.n254 99.6594
R13884 gnd.n463 gnd.n255 99.6594
R13885 gnd.n459 gnd.n256 99.6594
R13886 gnd.n455 gnd.n257 99.6594
R13887 gnd.n451 gnd.n258 99.6594
R13888 gnd.n447 gnd.n259 99.6594
R13889 gnd.n439 gnd.n260 99.6594
R13890 gnd.n1974 gnd.n1890 99.6594
R13891 gnd.n1892 gnd.n1816 99.6594
R13892 gnd.n1893 gnd.n1823 99.6594
R13893 gnd.n1895 gnd.n1894 99.6594
R13894 gnd.n1897 gnd.n1832 99.6594
R13895 gnd.n1898 gnd.n1839 99.6594
R13896 gnd.n1900 gnd.n1899 99.6594
R13897 gnd.n1902 gnd.n1848 99.6594
R13898 gnd.n4502 gnd.n1857 99.6594
R13899 gnd.n6445 gnd.n1135 99.6594
R13900 gnd.n6451 gnd.n1136 99.6594
R13901 gnd.n6455 gnd.n1137 99.6594
R13902 gnd.n6461 gnd.n1138 99.6594
R13903 gnd.n6465 gnd.n1139 99.6594
R13904 gnd.n6471 gnd.n1140 99.6594
R13905 gnd.n6475 gnd.n1141 99.6594
R13906 gnd.n6481 gnd.n1142 99.6594
R13907 gnd.n6485 gnd.n1143 99.6594
R13908 gnd.n6491 gnd.n1144 99.6594
R13909 gnd.n6498 gnd.n1145 99.6594
R13910 gnd.n6504 gnd.n1146 99.6594
R13911 gnd.n6507 gnd.n1147 99.6594
R13912 gnd.n5613 gnd.n5523 99.6594
R13913 gnd.n5611 gnd.n5526 99.6594
R13914 gnd.n5607 gnd.n5606 99.6594
R13915 gnd.n5600 gnd.n5531 99.6594
R13916 gnd.n5599 gnd.n5598 99.6594
R13917 gnd.n5592 gnd.n5537 99.6594
R13918 gnd.n5591 gnd.n5590 99.6594
R13919 gnd.n5584 gnd.n5543 99.6594
R13920 gnd.n5583 gnd.n5582 99.6594
R13921 gnd.n5576 gnd.n5549 99.6594
R13922 gnd.n5575 gnd.n5574 99.6594
R13923 gnd.n5567 gnd.n5555 99.6594
R13924 gnd.n5566 gnd.n5565 99.6594
R13925 gnd.n3073 gnd.n1554 99.6594
R13926 gnd.n3075 gnd.n1555 99.6594
R13927 gnd.n3083 gnd.n1556 99.6594
R13928 gnd.n3093 gnd.n1557 99.6594
R13929 gnd.n3095 gnd.n1558 99.6594
R13930 gnd.n3103 gnd.n1559 99.6594
R13931 gnd.n3113 gnd.n1560 99.6594
R13932 gnd.n3116 gnd.n1561 99.6594
R13933 gnd.n3320 gnd.n1562 99.6594
R13934 gnd.n2759 gnd.n1176 99.6594
R13935 gnd.n2763 gnd.n1177 99.6594
R13936 gnd.n2769 gnd.n1178 99.6594
R13937 gnd.n2773 gnd.n1179 99.6594
R13938 gnd.n2779 gnd.n1180 99.6594
R13939 gnd.n2783 gnd.n1181 99.6594
R13940 gnd.n2789 gnd.n1182 99.6594
R13941 gnd.n2793 gnd.n1183 99.6594
R13942 gnd.n2750 gnd.n1184 99.6594
R13943 gnd.n2762 gnd.n1176 99.6594
R13944 gnd.n2768 gnd.n1177 99.6594
R13945 gnd.n2772 gnd.n1178 99.6594
R13946 gnd.n2778 gnd.n1179 99.6594
R13947 gnd.n2782 gnd.n1180 99.6594
R13948 gnd.n2788 gnd.n1181 99.6594
R13949 gnd.n2792 gnd.n1182 99.6594
R13950 gnd.n2749 gnd.n1183 99.6594
R13951 gnd.n2745 gnd.n1184 99.6594
R13952 gnd.n3115 gnd.n1562 99.6594
R13953 gnd.n3114 gnd.n1561 99.6594
R13954 gnd.n3104 gnd.n1560 99.6594
R13955 gnd.n3096 gnd.n1559 99.6594
R13956 gnd.n3094 gnd.n1558 99.6594
R13957 gnd.n3084 gnd.n1557 99.6594
R13958 gnd.n3076 gnd.n1556 99.6594
R13959 gnd.n3074 gnd.n1555 99.6594
R13960 gnd.n3064 gnd.n1554 99.6594
R13961 gnd.n5614 gnd.n5613 99.6594
R13962 gnd.n5608 gnd.n5526 99.6594
R13963 gnd.n5606 gnd.n5605 99.6594
R13964 gnd.n5601 gnd.n5600 99.6594
R13965 gnd.n5598 gnd.n5597 99.6594
R13966 gnd.n5593 gnd.n5592 99.6594
R13967 gnd.n5590 gnd.n5589 99.6594
R13968 gnd.n5585 gnd.n5584 99.6594
R13969 gnd.n5582 gnd.n5581 99.6594
R13970 gnd.n5577 gnd.n5576 99.6594
R13971 gnd.n5574 gnd.n5573 99.6594
R13972 gnd.n5568 gnd.n5567 99.6594
R13973 gnd.n5565 gnd.n5521 99.6594
R13974 gnd.n6505 gnd.n1147 99.6594
R13975 gnd.n6497 gnd.n1146 99.6594
R13976 gnd.n6492 gnd.n1145 99.6594
R13977 gnd.n6484 gnd.n1144 99.6594
R13978 gnd.n6482 gnd.n1143 99.6594
R13979 gnd.n6474 gnd.n1142 99.6594
R13980 gnd.n6472 gnd.n1141 99.6594
R13981 gnd.n6464 gnd.n1140 99.6594
R13982 gnd.n6462 gnd.n1139 99.6594
R13983 gnd.n6454 gnd.n1138 99.6594
R13984 gnd.n6452 gnd.n1137 99.6594
R13985 gnd.n6444 gnd.n1136 99.6594
R13986 gnd.n6442 gnd.n1135 99.6594
R13987 gnd.n1890 gnd.n1815 99.6594
R13988 gnd.n1892 gnd.n1891 99.6594
R13989 gnd.n1893 gnd.n1824 99.6594
R13990 gnd.n1895 gnd.n1831 99.6594
R13991 gnd.n1897 gnd.n1896 99.6594
R13992 gnd.n1898 gnd.n1840 99.6594
R13993 gnd.n1900 gnd.n1847 99.6594
R13994 gnd.n1902 gnd.n1901 99.6594
R13995 gnd.n4503 gnd.n4502 99.6594
R13996 gnd.n446 gnd.n260 99.6594
R13997 gnd.n450 gnd.n259 99.6594
R13998 gnd.n454 gnd.n258 99.6594
R13999 gnd.n458 gnd.n257 99.6594
R14000 gnd.n462 gnd.n256 99.6594
R14001 gnd.n466 gnd.n255 99.6594
R14002 gnd.n470 gnd.n254 99.6594
R14003 gnd.n474 gnd.n253 99.6594
R14004 gnd.n349 gnd.n252 99.6594
R14005 gnd.n5741 gnd.n5691 99.6594
R14006 gnd.n5733 gnd.n5683 99.6594
R14007 gnd.n5729 gnd.n5684 99.6594
R14008 gnd.n5725 gnd.n5685 99.6594
R14009 gnd.n5721 gnd.n5686 99.6594
R14010 gnd.n5717 gnd.n5687 99.6594
R14011 gnd.n5713 gnd.n5688 99.6594
R14012 gnd.n5689 gnd.n5483 99.6594
R14013 gnd.n6561 gnd.n1128 99.6594
R14014 gnd.n6560 gnd.n1134 99.6594
R14015 gnd.n6535 gnd.n5112 99.6594
R14016 gnd.n6539 gnd.n5113 99.6594
R14017 gnd.n6543 gnd.n5114 99.6594
R14018 gnd.n6547 gnd.n5115 99.6594
R14019 gnd.n6551 gnd.n5116 99.6594
R14020 gnd.n5119 gnd.n5117 99.6594
R14021 gnd.n5110 gnd.n1188 99.6594
R14022 gnd.n5102 gnd.n1148 99.6594
R14023 gnd.n5098 gnd.n1149 99.6594
R14024 gnd.n5094 gnd.n1150 99.6594
R14025 gnd.n5090 gnd.n1151 99.6594
R14026 gnd.n5086 gnd.n1152 99.6594
R14027 gnd.n5082 gnd.n1153 99.6594
R14028 gnd.n5078 gnd.n1154 99.6594
R14029 gnd.n5073 gnd.n1155 99.6594
R14030 gnd.n5069 gnd.n1156 99.6594
R14031 gnd.n5065 gnd.n1157 99.6594
R14032 gnd.n5061 gnd.n1158 99.6594
R14033 gnd.n5057 gnd.n1159 99.6594
R14034 gnd.n5053 gnd.n1160 99.6594
R14035 gnd.n5049 gnd.n1161 99.6594
R14036 gnd.n5045 gnd.n1162 99.6594
R14037 gnd.n5041 gnd.n1163 99.6594
R14038 gnd.n5037 gnd.n1164 99.6594
R14039 gnd.n5033 gnd.n1165 99.6594
R14040 gnd.n5029 gnd.n1166 99.6594
R14041 gnd.n5025 gnd.n1167 99.6594
R14042 gnd.n5021 gnd.n1168 99.6594
R14043 gnd.n5017 gnd.n1169 99.6594
R14044 gnd.n5013 gnd.n1170 99.6594
R14045 gnd.n5009 gnd.n1171 99.6594
R14046 gnd.n5005 gnd.n1172 99.6594
R14047 gnd.n5001 gnd.n1173 99.6594
R14048 gnd.n4997 gnd.n1174 99.6594
R14049 gnd.n1258 gnd.n1175 99.6594
R14050 gnd.n3179 gnd.n1564 99.6594
R14051 gnd.n3260 gnd.n1565 99.6594
R14052 gnd.n3258 gnd.n1566 99.6594
R14053 gnd.n3250 gnd.n1567 99.6594
R14054 gnd.n3248 gnd.n1568 99.6594
R14055 gnd.n3240 gnd.n1569 99.6594
R14056 gnd.n3238 gnd.n1570 99.6594
R14057 gnd.n3230 gnd.n1571 99.6594
R14058 gnd.n3228 gnd.n1572 99.6594
R14059 gnd.n3220 gnd.n1573 99.6594
R14060 gnd.n3192 gnd.n1574 99.6594
R14061 gnd.n3211 gnd.n1575 99.6594
R14062 gnd.n3209 gnd.n1576 99.6594
R14063 gnd.n3201 gnd.n1577 99.6594
R14064 gnd.n3199 gnd.n1578 99.6594
R14065 gnd.n4762 gnd.n1580 99.6594
R14066 gnd.n4766 gnd.n1581 99.6594
R14067 gnd.n4770 gnd.n1582 99.6594
R14068 gnd.n4774 gnd.n1583 99.6594
R14069 gnd.n4779 gnd.n1584 99.6594
R14070 gnd.n4783 gnd.n1585 99.6594
R14071 gnd.n4787 gnd.n1586 99.6594
R14072 gnd.n4791 gnd.n1587 99.6594
R14073 gnd.n4795 gnd.n1588 99.6594
R14074 gnd.n4799 gnd.n1589 99.6594
R14075 gnd.n4803 gnd.n1590 99.6594
R14076 gnd.n1592 gnd.n1591 99.6594
R14077 gnd.n4809 gnd.n1551 99.6594
R14078 gnd.n4500 gnd.n1905 99.6594
R14079 gnd.n4492 gnd.n1862 99.6594
R14080 gnd.n4488 gnd.n1863 99.6594
R14081 gnd.n4484 gnd.n1864 99.6594
R14082 gnd.n4480 gnd.n1865 99.6594
R14083 gnd.n4476 gnd.n1866 99.6594
R14084 gnd.n4472 gnd.n1867 99.6594
R14085 gnd.n4468 gnd.n1868 99.6594
R14086 gnd.n4463 gnd.n1869 99.6594
R14087 gnd.n4459 gnd.n1870 99.6594
R14088 gnd.n4455 gnd.n1871 99.6594
R14089 gnd.n4451 gnd.n1872 99.6594
R14090 gnd.n4446 gnd.n1874 99.6594
R14091 gnd.n4442 gnd.n1875 99.6594
R14092 gnd.n4438 gnd.n1876 99.6594
R14093 gnd.n4434 gnd.n1877 99.6594
R14094 gnd.n4430 gnd.n1878 99.6594
R14095 gnd.n4426 gnd.n1879 99.6594
R14096 gnd.n4422 gnd.n1880 99.6594
R14097 gnd.n4418 gnd.n1881 99.6594
R14098 gnd.n4414 gnd.n1882 99.6594
R14099 gnd.n4410 gnd.n1883 99.6594
R14100 gnd.n4406 gnd.n1884 99.6594
R14101 gnd.n4402 gnd.n1885 99.6594
R14102 gnd.n4398 gnd.n1886 99.6594
R14103 gnd.n4394 gnd.n1887 99.6594
R14104 gnd.n4390 gnd.n1888 99.6594
R14105 gnd.n4382 gnd.n1889 99.6594
R14106 gnd.n7547 gnd.n261 99.6594
R14107 gnd.n7551 gnd.n262 99.6594
R14108 gnd.n7555 gnd.n263 99.6594
R14109 gnd.n7559 gnd.n264 99.6594
R14110 gnd.n7563 gnd.n265 99.6594
R14111 gnd.n7567 gnd.n266 99.6594
R14112 gnd.n7571 gnd.n267 99.6594
R14113 gnd.n7575 gnd.n268 99.6594
R14114 gnd.n7579 gnd.n269 99.6594
R14115 gnd.n7583 gnd.n270 99.6594
R14116 gnd.n7589 gnd.n271 99.6594
R14117 gnd.n7593 gnd.n272 99.6594
R14118 gnd.n7597 gnd.n273 99.6594
R14119 gnd.n7601 gnd.n274 99.6594
R14120 gnd.n7605 gnd.n275 99.6594
R14121 gnd.n7609 gnd.n276 99.6594
R14122 gnd.n7613 gnd.n277 99.6594
R14123 gnd.n7617 gnd.n278 99.6594
R14124 gnd.n7621 gnd.n279 99.6594
R14125 gnd.n7625 gnd.n280 99.6594
R14126 gnd.n7632 gnd.n281 99.6594
R14127 gnd.n7636 gnd.n282 99.6594
R14128 gnd.n7640 gnd.n283 99.6594
R14129 gnd.n7644 gnd.n284 99.6594
R14130 gnd.n7648 gnd.n285 99.6594
R14131 gnd.n7652 gnd.n286 99.6594
R14132 gnd.n7656 gnd.n287 99.6594
R14133 gnd.n289 gnd.n288 99.6594
R14134 gnd.n7662 gnd.n250 99.6594
R14135 gnd.n3047 gnd.n2559 99.6594
R14136 gnd.n3051 gnd.n2560 99.6594
R14137 gnd.n3034 gnd.n2561 99.6594
R14138 gnd.n3059 gnd.n2562 99.6594
R14139 gnd.n3061 gnd.n2563 99.6594
R14140 gnd.n3068 gnd.n2564 99.6594
R14141 gnd.n3070 gnd.n2565 99.6594
R14142 gnd.n3080 gnd.n2566 99.6594
R14143 gnd.n3088 gnd.n2567 99.6594
R14144 gnd.n3090 gnd.n2568 99.6594
R14145 gnd.n3100 gnd.n2569 99.6594
R14146 gnd.n3108 gnd.n2570 99.6594
R14147 gnd.n3110 gnd.n2571 99.6594
R14148 gnd.n3122 gnd.n2572 99.6594
R14149 gnd.n3050 gnd.n2559 99.6594
R14150 gnd.n3033 gnd.n2560 99.6594
R14151 gnd.n3058 gnd.n2561 99.6594
R14152 gnd.n3060 gnd.n2562 99.6594
R14153 gnd.n3067 gnd.n2563 99.6594
R14154 gnd.n3069 gnd.n2564 99.6594
R14155 gnd.n3079 gnd.n2565 99.6594
R14156 gnd.n3087 gnd.n2566 99.6594
R14157 gnd.n3089 gnd.n2567 99.6594
R14158 gnd.n3099 gnd.n2568 99.6594
R14159 gnd.n3107 gnd.n2569 99.6594
R14160 gnd.n3109 gnd.n2570 99.6594
R14161 gnd.n3121 gnd.n2571 99.6594
R14162 gnd.n2573 gnd.n2572 99.6594
R14163 gnd.n2079 gnd.n1796 99.6594
R14164 gnd.n2081 gnd.n1801 99.6594
R14165 gnd.n2082 gnd.n1804 99.6594
R14166 gnd.n2084 gnd.n1806 99.6594
R14167 gnd.n2085 gnd.n1810 99.6594
R14168 gnd.n2087 gnd.n2086 99.6594
R14169 gnd.n2089 gnd.n1820 99.6594
R14170 gnd.n2090 gnd.n1827 99.6594
R14171 gnd.n2092 gnd.n2091 99.6594
R14172 gnd.n2094 gnd.n1836 99.6594
R14173 gnd.n2095 gnd.n1843 99.6594
R14174 gnd.n2097 gnd.n2096 99.6594
R14175 gnd.n2100 gnd.n1852 99.6594
R14176 gnd.n4252 gnd.n2078 99.6594
R14177 gnd.n2097 gnd.n1851 99.6594
R14178 gnd.n2095 gnd.n1844 99.6594
R14179 gnd.n2094 gnd.n2093 99.6594
R14180 gnd.n2092 gnd.n1835 99.6594
R14181 gnd.n2090 gnd.n1828 99.6594
R14182 gnd.n2089 gnd.n2088 99.6594
R14183 gnd.n2087 gnd.n1819 99.6594
R14184 gnd.n2085 gnd.n1811 99.6594
R14185 gnd.n2084 gnd.n2083 99.6594
R14186 gnd.n2082 gnd.n1805 99.6594
R14187 gnd.n2081 gnd.n2080 99.6594
R14188 gnd.n2079 gnd.n1800 99.6594
R14189 gnd.n4253 gnd.n4252 99.6594
R14190 gnd.n2100 gnd.n2099 99.6594
R14191 gnd.n3118 gnd.t341 98.63
R14192 gnd.n4504 gnd.t373 98.63
R14193 gnd.n2577 gnd.t384 98.63
R14194 gnd.n1925 gnd.t366 98.63
R14195 gnd.n1948 gnd.t357 98.63
R14196 gnd.n4384 gnd.t295 98.63
R14197 gnd.n346 gnd.t390 98.63
R14198 gnd.n326 gnd.t309 98.63
R14199 gnd.n7628 gnd.t326 98.63
R14200 gnd.n366 gnd.t346 98.63
R14201 gnd.n1208 gnd.t360 98.63
R14202 gnd.n1230 gnd.t299 98.63
R14203 gnd.n1252 gnd.t317 98.63
R14204 gnd.n2746 gnd.t388 98.63
R14205 gnd.n1609 gnd.t381 98.63
R14206 gnd.n3177 gnd.t313 98.63
R14207 gnd.n3190 gnd.t336 98.63
R14208 gnd.n1853 gnd.t320 98.63
R14209 gnd.n3407 gnd.t351 92.8196
R14210 gnd.n2188 gnd.t375 92.8196
R14211 gnd.n4691 gnd.t401 92.8118
R14212 gnd.n2182 gnd.t305 92.8118
R14213 gnd.n7136 gnd.n7135 89.3769
R14214 gnd.n7137 gnd.n7136 89.3769
R14215 gnd.n7137 gnd.n712 89.3769
R14216 gnd.n7145 gnd.n712 89.3769
R14217 gnd.n7146 gnd.n7145 89.3769
R14218 gnd.n7147 gnd.n7146 89.3769
R14219 gnd.n7147 gnd.n706 89.3769
R14220 gnd.n7155 gnd.n706 89.3769
R14221 gnd.n7156 gnd.n7155 89.3769
R14222 gnd.n7157 gnd.n7156 89.3769
R14223 gnd.n7157 gnd.n700 89.3769
R14224 gnd.n7165 gnd.n700 89.3769
R14225 gnd.n7166 gnd.n7165 89.3769
R14226 gnd.n7167 gnd.n7166 89.3769
R14227 gnd.n7167 gnd.n694 89.3769
R14228 gnd.n7175 gnd.n694 89.3769
R14229 gnd.n7176 gnd.n7175 89.3769
R14230 gnd.n7177 gnd.n7176 89.3769
R14231 gnd.n7177 gnd.n688 89.3769
R14232 gnd.n7185 gnd.n688 89.3769
R14233 gnd.n7186 gnd.n7185 89.3769
R14234 gnd.n7187 gnd.n7186 89.3769
R14235 gnd.n7187 gnd.n682 89.3769
R14236 gnd.n7195 gnd.n682 89.3769
R14237 gnd.n7196 gnd.n7195 89.3769
R14238 gnd.n7197 gnd.n7196 89.3769
R14239 gnd.n7197 gnd.n676 89.3769
R14240 gnd.n7205 gnd.n676 89.3769
R14241 gnd.n7206 gnd.n7205 89.3769
R14242 gnd.n7207 gnd.n7206 89.3769
R14243 gnd.n7207 gnd.n670 89.3769
R14244 gnd.n7215 gnd.n670 89.3769
R14245 gnd.n7216 gnd.n7215 89.3769
R14246 gnd.n7217 gnd.n7216 89.3769
R14247 gnd.n7217 gnd.n664 89.3769
R14248 gnd.n7225 gnd.n664 89.3769
R14249 gnd.n7226 gnd.n7225 89.3769
R14250 gnd.n7227 gnd.n7226 89.3769
R14251 gnd.n7227 gnd.n658 89.3769
R14252 gnd.n7235 gnd.n658 89.3769
R14253 gnd.n7236 gnd.n7235 89.3769
R14254 gnd.n7237 gnd.n7236 89.3769
R14255 gnd.n7237 gnd.n652 89.3769
R14256 gnd.n7245 gnd.n652 89.3769
R14257 gnd.n7246 gnd.n7245 89.3769
R14258 gnd.n7247 gnd.n7246 89.3769
R14259 gnd.n7247 gnd.n646 89.3769
R14260 gnd.n7255 gnd.n646 89.3769
R14261 gnd.n7256 gnd.n7255 89.3769
R14262 gnd.n7257 gnd.n7256 89.3769
R14263 gnd.n7257 gnd.n640 89.3769
R14264 gnd.n7265 gnd.n640 89.3769
R14265 gnd.n7266 gnd.n7265 89.3769
R14266 gnd.n7267 gnd.n7266 89.3769
R14267 gnd.n7267 gnd.n634 89.3769
R14268 gnd.n7275 gnd.n634 89.3769
R14269 gnd.n7276 gnd.n7275 89.3769
R14270 gnd.n7277 gnd.n7276 89.3769
R14271 gnd.n7277 gnd.n628 89.3769
R14272 gnd.n7285 gnd.n628 89.3769
R14273 gnd.n7286 gnd.n7285 89.3769
R14274 gnd.n7287 gnd.n7286 89.3769
R14275 gnd.n7287 gnd.n622 89.3769
R14276 gnd.n7295 gnd.n622 89.3769
R14277 gnd.n7296 gnd.n7295 89.3769
R14278 gnd.n7297 gnd.n7296 89.3769
R14279 gnd.n7297 gnd.n616 89.3769
R14280 gnd.n7305 gnd.n616 89.3769
R14281 gnd.n7306 gnd.n7305 89.3769
R14282 gnd.n7307 gnd.n7306 89.3769
R14283 gnd.n7307 gnd.n610 89.3769
R14284 gnd.n7315 gnd.n610 89.3769
R14285 gnd.n7316 gnd.n7315 89.3769
R14286 gnd.n7317 gnd.n7316 89.3769
R14287 gnd.n7317 gnd.n604 89.3769
R14288 gnd.n7325 gnd.n604 89.3769
R14289 gnd.n7326 gnd.n7325 89.3769
R14290 gnd.n7327 gnd.n7326 89.3769
R14291 gnd.n7327 gnd.n598 89.3769
R14292 gnd.n7335 gnd.n598 89.3769
R14293 gnd.n7336 gnd.n7335 89.3769
R14294 gnd.n7339 gnd.n7336 89.3769
R14295 gnd.n7339 gnd.n7338 89.3769
R14296 gnd.n1671 gnd.n1670 81.8399
R14297 gnd.n4448 gnd.n1935 78.9125
R14298 gnd.n4760 gnd.n4759 78.9125
R14299 gnd.n5709 gnd.t333 74.8376
R14300 gnd.n1130 gnd.t370 74.8376
R14301 gnd.n3408 gnd.t350 72.8438
R14302 gnd.n2189 gnd.t376 72.8438
R14303 gnd.n1672 gnd.n1665 72.8411
R14304 gnd.n1678 gnd.n1663 72.8411
R14305 gnd.n2157 gnd.n2156 72.8411
R14306 gnd.n3119 gnd.t340 72.836
R14307 gnd.n4692 gnd.t400 72.836
R14308 gnd.n2183 gnd.t306 72.836
R14309 gnd.n4505 gnd.t372 72.836
R14310 gnd.n2578 gnd.t385 72.836
R14311 gnd.n1926 gnd.t365 72.836
R14312 gnd.n1949 gnd.t356 72.836
R14313 gnd.n4385 gnd.t294 72.836
R14314 gnd.n347 gnd.t391 72.836
R14315 gnd.n327 gnd.t310 72.836
R14316 gnd.n7629 gnd.t327 72.836
R14317 gnd.n367 gnd.t347 72.836
R14318 gnd.n1209 gnd.t359 72.836
R14319 gnd.n1231 gnd.t298 72.836
R14320 gnd.n1253 gnd.t316 72.836
R14321 gnd.n2747 gnd.t387 72.836
R14322 gnd.n1610 gnd.t382 72.836
R14323 gnd.n3178 gnd.t314 72.836
R14324 gnd.n3191 gnd.t337 72.836
R14325 gnd.n1854 gnd.t321 72.836
R14326 gnd.n4150 gnd.n4149 71.676
R14327 gnd.n4147 gnd.n4146 71.676
R14328 gnd.n4142 gnd.n2165 71.676
R14329 gnd.n4140 gnd.n4139 71.676
R14330 gnd.n4135 gnd.n2168 71.676
R14331 gnd.n4133 gnd.n4132 71.676
R14332 gnd.n4128 gnd.n2171 71.676
R14333 gnd.n4126 gnd.n4125 71.676
R14334 gnd.n4121 gnd.n2174 71.676
R14335 gnd.n4119 gnd.n4118 71.676
R14336 gnd.n4114 gnd.n2177 71.676
R14337 gnd.n4112 gnd.n4111 71.676
R14338 gnd.n4107 gnd.n2180 71.676
R14339 gnd.n4105 gnd.n4104 71.676
R14340 gnd.n4099 gnd.n2185 71.676
R14341 gnd.n4097 gnd.n4096 71.676
R14342 gnd.n4092 gnd.n4091 71.676
R14343 gnd.n4089 gnd.n4088 71.676
R14344 gnd.n4083 gnd.n2191 71.676
R14345 gnd.n4081 gnd.n4080 71.676
R14346 gnd.n4076 gnd.n2194 71.676
R14347 gnd.n4074 gnd.n4073 71.676
R14348 gnd.n4069 gnd.n2197 71.676
R14349 gnd.n4067 gnd.n4066 71.676
R14350 gnd.n4062 gnd.n2200 71.676
R14351 gnd.n4060 gnd.n4059 71.676
R14352 gnd.n4055 gnd.n2203 71.676
R14353 gnd.n4053 gnd.n4052 71.676
R14354 gnd.n4048 gnd.n2206 71.676
R14355 gnd.n4046 gnd.n4045 71.676
R14356 gnd.n4041 gnd.n2209 71.676
R14357 gnd.n4039 gnd.n4038 71.676
R14358 gnd.n4034 gnd.n4032 71.676
R14359 gnd.n4755 gnd.n4754 71.676
R14360 gnd.n4749 gnd.n1627 71.676
R14361 gnd.n4746 gnd.n1628 71.676
R14362 gnd.n4742 gnd.n1629 71.676
R14363 gnd.n4738 gnd.n1630 71.676
R14364 gnd.n4734 gnd.n1631 71.676
R14365 gnd.n4730 gnd.n1632 71.676
R14366 gnd.n4726 gnd.n1633 71.676
R14367 gnd.n4722 gnd.n1634 71.676
R14368 gnd.n4718 gnd.n1635 71.676
R14369 gnd.n4714 gnd.n1636 71.676
R14370 gnd.n4710 gnd.n1637 71.676
R14371 gnd.n4706 gnd.n1638 71.676
R14372 gnd.n4702 gnd.n1639 71.676
R14373 gnd.n4698 gnd.n1640 71.676
R14374 gnd.n4694 gnd.n1641 71.676
R14375 gnd.n1642 gnd.n1625 71.676
R14376 gnd.n3411 gnd.n1643 71.676
R14377 gnd.n3416 gnd.n1644 71.676
R14378 gnd.n3420 gnd.n1645 71.676
R14379 gnd.n3424 gnd.n1646 71.676
R14380 gnd.n3428 gnd.n1647 71.676
R14381 gnd.n3432 gnd.n1648 71.676
R14382 gnd.n3436 gnd.n1649 71.676
R14383 gnd.n3440 gnd.n1650 71.676
R14384 gnd.n3444 gnd.n1651 71.676
R14385 gnd.n3448 gnd.n1652 71.676
R14386 gnd.n3452 gnd.n1653 71.676
R14387 gnd.n3456 gnd.n1654 71.676
R14388 gnd.n3460 gnd.n1655 71.676
R14389 gnd.n3464 gnd.n1656 71.676
R14390 gnd.n3468 gnd.n1657 71.676
R14391 gnd.n4755 gnd.n1660 71.676
R14392 gnd.n4747 gnd.n1627 71.676
R14393 gnd.n4743 gnd.n1628 71.676
R14394 gnd.n4739 gnd.n1629 71.676
R14395 gnd.n4735 gnd.n1630 71.676
R14396 gnd.n4731 gnd.n1631 71.676
R14397 gnd.n4727 gnd.n1632 71.676
R14398 gnd.n4723 gnd.n1633 71.676
R14399 gnd.n4719 gnd.n1634 71.676
R14400 gnd.n4715 gnd.n1635 71.676
R14401 gnd.n4711 gnd.n1636 71.676
R14402 gnd.n4707 gnd.n1637 71.676
R14403 gnd.n4703 gnd.n1638 71.676
R14404 gnd.n4699 gnd.n1639 71.676
R14405 gnd.n4695 gnd.n1640 71.676
R14406 gnd.n4758 gnd.n4757 71.676
R14407 gnd.n3410 gnd.n1642 71.676
R14408 gnd.n3415 gnd.n1643 71.676
R14409 gnd.n3419 gnd.n1644 71.676
R14410 gnd.n3423 gnd.n1645 71.676
R14411 gnd.n3427 gnd.n1646 71.676
R14412 gnd.n3431 gnd.n1647 71.676
R14413 gnd.n3435 gnd.n1648 71.676
R14414 gnd.n3439 gnd.n1649 71.676
R14415 gnd.n3443 gnd.n1650 71.676
R14416 gnd.n3447 gnd.n1651 71.676
R14417 gnd.n3451 gnd.n1652 71.676
R14418 gnd.n3455 gnd.n1653 71.676
R14419 gnd.n3459 gnd.n1654 71.676
R14420 gnd.n3463 gnd.n1655 71.676
R14421 gnd.n3467 gnd.n1656 71.676
R14422 gnd.n3471 gnd.n1657 71.676
R14423 gnd.n4032 gnd.n2210 71.676
R14424 gnd.n4040 gnd.n4039 71.676
R14425 gnd.n2209 gnd.n2207 71.676
R14426 gnd.n4047 gnd.n4046 71.676
R14427 gnd.n2206 gnd.n2204 71.676
R14428 gnd.n4054 gnd.n4053 71.676
R14429 gnd.n2203 gnd.n2201 71.676
R14430 gnd.n4061 gnd.n4060 71.676
R14431 gnd.n2200 gnd.n2198 71.676
R14432 gnd.n4068 gnd.n4067 71.676
R14433 gnd.n2197 gnd.n2195 71.676
R14434 gnd.n4075 gnd.n4074 71.676
R14435 gnd.n2194 gnd.n2192 71.676
R14436 gnd.n4082 gnd.n4081 71.676
R14437 gnd.n2191 gnd.n2187 71.676
R14438 gnd.n4090 gnd.n4089 71.676
R14439 gnd.n4094 gnd.n4093 71.676
R14440 gnd.n4098 gnd.n4097 71.676
R14441 gnd.n2185 gnd.n2181 71.676
R14442 gnd.n4106 gnd.n4105 71.676
R14443 gnd.n2180 gnd.n2178 71.676
R14444 gnd.n4113 gnd.n4112 71.676
R14445 gnd.n2177 gnd.n2175 71.676
R14446 gnd.n4120 gnd.n4119 71.676
R14447 gnd.n2174 gnd.n2172 71.676
R14448 gnd.n4127 gnd.n4126 71.676
R14449 gnd.n2171 gnd.n2169 71.676
R14450 gnd.n4134 gnd.n4133 71.676
R14451 gnd.n2168 gnd.n2166 71.676
R14452 gnd.n4141 gnd.n4140 71.676
R14453 gnd.n2165 gnd.n2163 71.676
R14454 gnd.n4148 gnd.n4147 71.676
R14455 gnd.n4151 gnd.n4150 71.676
R14456 gnd.n8 gnd.t151 69.1507
R14457 gnd.n14 gnd.t231 68.4792
R14458 gnd.n13 gnd.t72 68.4792
R14459 gnd.n12 gnd.t403 68.4792
R14460 gnd.n11 gnd.t153 68.4792
R14461 gnd.n10 gnd.t9 68.4792
R14462 gnd.n9 gnd.t229 68.4792
R14463 gnd.n8 gnd.t264 68.4792
R14464 gnd.n5621 gnd.n5522 64.369
R14465 gnd.n3413 gnd.n3408 59.5399
R14466 gnd.n4085 gnd.n2189 59.5399
R14467 gnd.n4693 gnd.n4692 59.5399
R14468 gnd.n4101 gnd.n2183 59.5399
R14469 gnd.n4690 gnd.n1681 59.1804
R14470 gnd.n6559 gnd.n1120 57.3586
R14471 gnd.n5324 gnd.t84 56.407
R14472 gnd.n5265 gnd.t268 56.407
R14473 gnd.n5284 gnd.t95 56.407
R14474 gnd.n5304 gnd.t3 56.407
R14475 gnd.n76 gnd.t244 56.407
R14476 gnd.n17 gnd.t61 56.407
R14477 gnd.n36 gnd.t227 56.407
R14478 gnd.n56 gnd.t405 56.407
R14479 gnd.n5341 gnd.t205 55.8337
R14480 gnd.n5282 gnd.t52 55.8337
R14481 gnd.n5301 gnd.t277 55.8337
R14482 gnd.n5321 gnd.t96 55.8337
R14483 gnd.n93 gnd.t260 55.8337
R14484 gnd.n34 gnd.t190 55.8337
R14485 gnd.n53 gnd.t224 55.8337
R14486 gnd.n73 gnd.t235 55.8337
R14487 gnd.n1669 gnd.n1668 54.358
R14488 gnd.n2154 gnd.n2153 54.358
R14489 gnd.n7338 gnd.n7337 53.6263
R14490 gnd.n5324 gnd.n5323 53.0052
R14491 gnd.n5326 gnd.n5325 53.0052
R14492 gnd.n5328 gnd.n5327 53.0052
R14493 gnd.n5330 gnd.n5329 53.0052
R14494 gnd.n5332 gnd.n5331 53.0052
R14495 gnd.n5334 gnd.n5333 53.0052
R14496 gnd.n5336 gnd.n5335 53.0052
R14497 gnd.n5338 gnd.n5337 53.0052
R14498 gnd.n5340 gnd.n5339 53.0052
R14499 gnd.n5265 gnd.n5264 53.0052
R14500 gnd.n5267 gnd.n5266 53.0052
R14501 gnd.n5269 gnd.n5268 53.0052
R14502 gnd.n5271 gnd.n5270 53.0052
R14503 gnd.n5273 gnd.n5272 53.0052
R14504 gnd.n5275 gnd.n5274 53.0052
R14505 gnd.n5277 gnd.n5276 53.0052
R14506 gnd.n5279 gnd.n5278 53.0052
R14507 gnd.n5281 gnd.n5280 53.0052
R14508 gnd.n5284 gnd.n5283 53.0052
R14509 gnd.n5286 gnd.n5285 53.0052
R14510 gnd.n5288 gnd.n5287 53.0052
R14511 gnd.n5290 gnd.n5289 53.0052
R14512 gnd.n5292 gnd.n5291 53.0052
R14513 gnd.n5294 gnd.n5293 53.0052
R14514 gnd.n5296 gnd.n5295 53.0052
R14515 gnd.n5298 gnd.n5297 53.0052
R14516 gnd.n5300 gnd.n5299 53.0052
R14517 gnd.n5304 gnd.n5303 53.0052
R14518 gnd.n5306 gnd.n5305 53.0052
R14519 gnd.n5308 gnd.n5307 53.0052
R14520 gnd.n5310 gnd.n5309 53.0052
R14521 gnd.n5312 gnd.n5311 53.0052
R14522 gnd.n5314 gnd.n5313 53.0052
R14523 gnd.n5316 gnd.n5315 53.0052
R14524 gnd.n5318 gnd.n5317 53.0052
R14525 gnd.n5320 gnd.n5319 53.0052
R14526 gnd.n92 gnd.n91 53.0052
R14527 gnd.n90 gnd.n89 53.0052
R14528 gnd.n88 gnd.n87 53.0052
R14529 gnd.n86 gnd.n85 53.0052
R14530 gnd.n84 gnd.n83 53.0052
R14531 gnd.n82 gnd.n81 53.0052
R14532 gnd.n80 gnd.n79 53.0052
R14533 gnd.n78 gnd.n77 53.0052
R14534 gnd.n76 gnd.n75 53.0052
R14535 gnd.n33 gnd.n32 53.0052
R14536 gnd.n31 gnd.n30 53.0052
R14537 gnd.n29 gnd.n28 53.0052
R14538 gnd.n27 gnd.n26 53.0052
R14539 gnd.n25 gnd.n24 53.0052
R14540 gnd.n23 gnd.n22 53.0052
R14541 gnd.n21 gnd.n20 53.0052
R14542 gnd.n19 gnd.n18 53.0052
R14543 gnd.n17 gnd.n16 53.0052
R14544 gnd.n52 gnd.n51 53.0052
R14545 gnd.n50 gnd.n49 53.0052
R14546 gnd.n48 gnd.n47 53.0052
R14547 gnd.n46 gnd.n45 53.0052
R14548 gnd.n44 gnd.n43 53.0052
R14549 gnd.n42 gnd.n41 53.0052
R14550 gnd.n40 gnd.n39 53.0052
R14551 gnd.n38 gnd.n37 53.0052
R14552 gnd.n36 gnd.n35 53.0052
R14553 gnd.n72 gnd.n71 53.0052
R14554 gnd.n70 gnd.n69 53.0052
R14555 gnd.n68 gnd.n67 53.0052
R14556 gnd.n66 gnd.n65 53.0052
R14557 gnd.n64 gnd.n63 53.0052
R14558 gnd.n62 gnd.n61 53.0052
R14559 gnd.n60 gnd.n59 53.0052
R14560 gnd.n58 gnd.n57 53.0052
R14561 gnd.n56 gnd.n55 53.0052
R14562 gnd.n2145 gnd.n2144 52.4801
R14563 gnd.n6367 gnd.t219 52.3082
R14564 gnd.n6335 gnd.t280 52.3082
R14565 gnd.n6303 gnd.t164 52.3082
R14566 gnd.n6272 gnd.t208 52.3082
R14567 gnd.n6240 gnd.t243 52.3082
R14568 gnd.n6208 gnd.t187 52.3082
R14569 gnd.n6176 gnd.t90 52.3082
R14570 gnd.n6145 gnd.t271 52.3082
R14571 gnd.n5111 gnd.n1186 51.6227
R14572 gnd.n7663 gnd.n244 51.6227
R14573 gnd.n6197 gnd.n6165 51.4173
R14574 gnd.n6261 gnd.n6260 50.455
R14575 gnd.n6229 gnd.n6228 50.455
R14576 gnd.n6197 gnd.n6196 50.455
R14577 gnd.n5559 gnd.n5558 45.1884
R14578 gnd.n6495 gnd.n6494 45.1884
R14579 gnd.n4153 gnd.n2160 44.3322
R14580 gnd.n1672 gnd.n1671 44.3189
R14581 gnd.n3120 gnd.n3119 42.2793
R14582 gnd.n4506 gnd.n4505 42.2793
R14583 gnd.n5571 gnd.n5559 42.2793
R14584 gnd.n6496 gnd.n6495 42.2793
R14585 gnd.n5711 gnd.n5709 42.2793
R14586 gnd.n1131 gnd.n1130 42.2793
R14587 gnd.n2579 gnd.n2578 42.2793
R14588 gnd.n4465 gnd.n1926 42.2793
R14589 gnd.n4428 gnd.n1949 42.2793
R14590 gnd.n4388 gnd.n4385 42.2793
R14591 gnd.n7546 gnd.n347 42.2793
R14592 gnd.n7588 gnd.n327 42.2793
R14593 gnd.n7630 gnd.n7629 42.2793
R14594 gnd.n445 gnd.n367 42.2793
R14595 gnd.n5075 gnd.n1209 42.2793
R14596 gnd.n5035 gnd.n1231 42.2793
R14597 gnd.n4995 gnd.n1253 42.2793
R14598 gnd.n2799 gnd.n2747 42.2793
R14599 gnd.n4777 gnd.n1610 42.2793
R14600 gnd.n3268 gnd.n3178 42.2793
R14601 gnd.n3219 gnd.n3191 42.2793
R14602 gnd.n1855 gnd.n1854 42.2793
R14603 gnd.n1670 gnd.n1669 41.6274
R14604 gnd.n2155 gnd.n2154 41.6274
R14605 gnd.n1679 gnd.n1678 40.8975
R14606 gnd.n2158 gnd.n2157 40.8975
R14607 gnd.n1678 gnd.n1677 35.055
R14608 gnd.n1673 gnd.n1672 35.055
R14609 gnd.n2147 gnd.n2146 35.055
R14610 gnd.n2157 gnd.n2143 35.055
R14611 gnd.n6744 gnd.n951 32.6173
R14612 gnd.n6738 gnd.n951 32.6173
R14613 gnd.n6738 gnd.n6737 32.6173
R14614 gnd.n6737 gnd.n6736 32.6173
R14615 gnd.n6736 gnd.n958 32.6173
R14616 gnd.n6730 gnd.n958 32.6173
R14617 gnd.n6730 gnd.n6729 32.6173
R14618 gnd.n6729 gnd.n6728 32.6173
R14619 gnd.n6728 gnd.n966 32.6173
R14620 gnd.n6722 gnd.n966 32.6173
R14621 gnd.n6722 gnd.n6721 32.6173
R14622 gnd.n6721 gnd.n6720 32.6173
R14623 gnd.n6720 gnd.n974 32.6173
R14624 gnd.n6714 gnd.n974 32.6173
R14625 gnd.n6714 gnd.n6713 32.6173
R14626 gnd.n6713 gnd.n6712 32.6173
R14627 gnd.n6712 gnd.n982 32.6173
R14628 gnd.n6706 gnd.n982 32.6173
R14629 gnd.n6706 gnd.n6705 32.6173
R14630 gnd.n6705 gnd.n6704 32.6173
R14631 gnd.n6704 gnd.n990 32.6173
R14632 gnd.n6698 gnd.n990 32.6173
R14633 gnd.n6698 gnd.n6697 32.6173
R14634 gnd.n6697 gnd.n6696 32.6173
R14635 gnd.n6696 gnd.n998 32.6173
R14636 gnd.n6690 gnd.n998 32.6173
R14637 gnd.n6690 gnd.n6689 32.6173
R14638 gnd.n6689 gnd.n6688 32.6173
R14639 gnd.n6688 gnd.n1006 32.6173
R14640 gnd.n6682 gnd.n1006 32.6173
R14641 gnd.n6682 gnd.n6681 32.6173
R14642 gnd.n6681 gnd.n6680 32.6173
R14643 gnd.n6680 gnd.n1014 32.6173
R14644 gnd.n6674 gnd.n1014 32.6173
R14645 gnd.n6674 gnd.n6673 32.6173
R14646 gnd.n6673 gnd.n6672 32.6173
R14647 gnd.n6672 gnd.n1022 32.6173
R14648 gnd.n6666 gnd.n1022 32.6173
R14649 gnd.n6666 gnd.n6665 32.6173
R14650 gnd.n6665 gnd.n6664 32.6173
R14651 gnd.n6664 gnd.n1030 32.6173
R14652 gnd.n6658 gnd.n1030 32.6173
R14653 gnd.n6658 gnd.n6657 32.6173
R14654 gnd.n6657 gnd.n6656 32.6173
R14655 gnd.n6656 gnd.n1038 32.6173
R14656 gnd.n6650 gnd.n1038 32.6173
R14657 gnd.n6650 gnd.n6649 32.6173
R14658 gnd.n6649 gnd.n6648 32.6173
R14659 gnd.n6648 gnd.n1046 32.6173
R14660 gnd.n6642 gnd.n1046 32.6173
R14661 gnd.n6642 gnd.n6641 32.6173
R14662 gnd.n6641 gnd.n6640 32.6173
R14663 gnd.n6640 gnd.n1054 32.6173
R14664 gnd.n6634 gnd.n1054 32.6173
R14665 gnd.n6634 gnd.n6633 32.6173
R14666 gnd.n6633 gnd.n6632 32.6173
R14667 gnd.n6632 gnd.n1062 32.6173
R14668 gnd.n6626 gnd.n1062 32.6173
R14669 gnd.n6626 gnd.n6625 32.6173
R14670 gnd.n6625 gnd.n6624 32.6173
R14671 gnd.n6624 gnd.n1070 32.6173
R14672 gnd.n6618 gnd.n1070 32.6173
R14673 gnd.n6618 gnd.n6617 32.6173
R14674 gnd.n6617 gnd.n6616 32.6173
R14675 gnd.n6616 gnd.n1078 32.6173
R14676 gnd.n6610 gnd.n1078 32.6173
R14677 gnd.n6610 gnd.n6609 32.6173
R14678 gnd.n6609 gnd.n6608 32.6173
R14679 gnd.n6608 gnd.n1086 32.6173
R14680 gnd.n6602 gnd.n1086 32.6173
R14681 gnd.n6602 gnd.n6601 32.6173
R14682 gnd.n6601 gnd.n6600 32.6173
R14683 gnd.n6600 gnd.n1094 32.6173
R14684 gnd.n6594 gnd.n1094 32.6173
R14685 gnd.n6594 gnd.n6593 32.6173
R14686 gnd.n6593 gnd.n6592 32.6173
R14687 gnd.n6592 gnd.n1102 32.6173
R14688 gnd.n6586 gnd.n1102 32.6173
R14689 gnd.n6586 gnd.n6585 32.6173
R14690 gnd.n6585 gnd.n6584 32.6173
R14691 gnd.n6584 gnd.n1110 32.6173
R14692 gnd.n6578 gnd.n1110 32.6173
R14693 gnd.n6578 gnd.n6577 32.6173
R14694 gnd.n5621 gnd.n5517 31.8661
R14695 gnd.n5629 gnd.n5517 31.8661
R14696 gnd.n5637 gnd.n5511 31.8661
R14697 gnd.n5637 gnd.n5505 31.8661
R14698 gnd.n5645 gnd.n5505 31.8661
R14699 gnd.n5645 gnd.n5498 31.8661
R14700 gnd.n5653 gnd.n5498 31.8661
R14701 gnd.n5653 gnd.n5499 31.8661
R14702 gnd.n5752 gnd.n5484 31.8661
R14703 gnd.n4987 gnd.n1186 31.8661
R14704 gnd.n4981 gnd.n1270 31.8661
R14705 gnd.n4981 gnd.n1273 31.8661
R14706 gnd.n4975 gnd.n1273 31.8661
R14707 gnd.n4975 gnd.n1285 31.8661
R14708 gnd.n4969 gnd.n1295 31.8661
R14709 gnd.n4963 gnd.n1295 31.8661
R14710 gnd.n4957 gnd.n1311 31.8661
R14711 gnd.n4957 gnd.n1314 31.8661
R14712 gnd.n4951 gnd.n1323 31.8661
R14713 gnd.n4945 gnd.n1333 31.8661
R14714 gnd.n4939 gnd.n1333 31.8661
R14715 gnd.n4933 gnd.n1349 31.8661
R14716 gnd.n4933 gnd.n1352 31.8661
R14717 gnd.n4927 gnd.n1361 31.8661
R14718 gnd.n4921 gnd.n1371 31.8661
R14719 gnd.n4915 gnd.n1371 31.8661
R14720 gnd.n4909 gnd.n1386 31.8661
R14721 gnd.n4909 gnd.n1389 31.8661
R14722 gnd.n4903 gnd.n1398 31.8661
R14723 gnd.n2869 gnd.n2726 31.8661
R14724 gnd.n3317 gnd.n1552 31.8661
R14725 gnd.n2558 gnd.n1563 31.8661
R14726 gnd.n3328 gnd.n2558 31.8661
R14727 gnd.n3329 gnd.n3328 31.8661
R14728 gnd.n3329 gnd.n2551 31.8661
R14729 gnd.n3337 gnd.n2551 31.8661
R14730 gnd.n3362 gnd.n2542 31.8661
R14731 gnd.n3362 gnd.n2533 31.8661
R14732 gnd.n3379 gnd.n2533 31.8661
R14733 gnd.n3379 gnd.n2534 31.8661
R14734 gnd.n4174 gnd.n2115 31.8661
R14735 gnd.n4185 gnd.n2115 31.8661
R14736 gnd.n4185 gnd.n2108 31.8661
R14737 gnd.n4193 gnd.n2108 31.8661
R14738 gnd.n4569 gnd.n1792 31.8661
R14739 gnd.n4569 gnd.n1794 31.8661
R14740 gnd.n4251 gnd.n1794 31.8661
R14741 gnd.n4251 gnd.n2101 31.8661
R14742 gnd.n2101 gnd.n1861 31.8661
R14743 gnd.n1971 gnd.n1903 31.8661
R14744 gnd.n7482 gnd.n485 31.8661
R14745 gnd.n7757 gnd.n102 31.8661
R14746 gnd.n7749 gnd.n117 31.8661
R14747 gnd.n7749 gnd.n120 31.8661
R14748 gnd.n7743 gnd.n131 31.8661
R14749 gnd.n7737 gnd.n131 31.8661
R14750 gnd.n7731 gnd.n146 31.8661
R14751 gnd.n7725 gnd.n156 31.8661
R14752 gnd.n7725 gnd.n159 31.8661
R14753 gnd.n7719 gnd.n168 31.8661
R14754 gnd.n7713 gnd.n168 31.8661
R14755 gnd.n7707 gnd.n184 31.8661
R14756 gnd.n7701 gnd.n194 31.8661
R14757 gnd.n7701 gnd.n197 31.8661
R14758 gnd.n7695 gnd.n206 31.8661
R14759 gnd.n7689 gnd.n206 31.8661
R14760 gnd.n7683 gnd.n222 31.8661
R14761 gnd.n7683 gnd.n225 31.8661
R14762 gnd.n7677 gnd.n225 31.8661
R14763 gnd.n7677 gnd.n235 31.8661
R14764 gnd.n7671 gnd.n244 31.8661
R14765 gnd.n4903 gnd.t172 31.5474
R14766 gnd.t45 gnd.n102 31.5474
R14767 gnd.n4035 gnd.n4031 31.3761
R14768 gnd.n3474 gnd.n3470 31.3761
R14769 gnd.n4927 gnd.t67 30.9101
R14770 gnd.n7731 gnd.t101 30.9101
R14771 gnd.n4951 gnd.t47 30.2728
R14772 gnd.n7707 gnd.t43 30.2728
R14773 gnd.n4987 gnd.t297 28.3609
R14774 gnd.n7671 gnd.t308 28.3609
R14775 gnd.n4810 gnd.n1563 27.4049
R14776 gnd.n4501 gnd.n1861 27.4049
R14777 gnd.n3119 gnd.n3118 25.7944
R14778 gnd.n4505 gnd.n4504 25.7944
R14779 gnd.n5709 gnd.n5708 25.7944
R14780 gnd.n1130 gnd.n1129 25.7944
R14781 gnd.n2578 gnd.n2577 25.7944
R14782 gnd.n1926 gnd.n1925 25.7944
R14783 gnd.n1949 gnd.n1948 25.7944
R14784 gnd.n4385 gnd.n4384 25.7944
R14785 gnd.n347 gnd.n346 25.7944
R14786 gnd.n327 gnd.n326 25.7944
R14787 gnd.n7629 gnd.n7628 25.7944
R14788 gnd.n367 gnd.n366 25.7944
R14789 gnd.n1209 gnd.n1208 25.7944
R14790 gnd.n1231 gnd.n1230 25.7944
R14791 gnd.n1253 gnd.n1252 25.7944
R14792 gnd.n2747 gnd.n2746 25.7944
R14793 gnd.n1610 gnd.n1609 25.7944
R14794 gnd.n3178 gnd.n3177 25.7944
R14795 gnd.n3191 gnd.n3190 25.7944
R14796 gnd.n1854 gnd.n1853 25.7944
R14797 gnd.n5753 gnd.n5473 24.8557
R14798 gnd.n5476 gnd.n5467 24.8557
R14799 gnd.n5774 gnd.n5452 24.8557
R14800 gnd.n5793 gnd.n5792 24.8557
R14801 gnd.n5803 gnd.n5445 24.8557
R14802 gnd.n5816 gnd.n5433 24.8557
R14803 gnd.n5841 gnd.n5417 24.8557
R14804 gnd.n5840 gnd.n5419 24.8557
R14805 gnd.n5863 gnd.n5401 24.8557
R14806 gnd.n5852 gnd.n5393 24.8557
R14807 gnd.n5888 gnd.n5887 24.8557
R14808 gnd.n5898 gnd.n5386 24.8557
R14809 gnd.n5910 gnd.n5378 24.8557
R14810 gnd.n5909 gnd.n5366 24.8557
R14811 gnd.n5928 gnd.n5927 24.8557
R14812 gnd.n5949 gnd.n5347 24.8557
R14813 gnd.n5970 gnd.n5969 24.8557
R14814 gnd.n5981 gnd.n5250 24.8557
R14815 gnd.n5980 gnd.n5252 24.8557
R14816 gnd.n5992 gnd.n5243 24.8557
R14817 gnd.n6011 gnd.n6010 24.8557
R14818 gnd.n5232 gnd.n5221 24.8557
R14819 gnd.n6037 gnd.n5214 24.8557
R14820 gnd.n6036 gnd.n6035 24.8557
R14821 gnd.n6055 gnd.n6054 24.8557
R14822 gnd.n5205 gnd.n5195 24.8557
R14823 gnd.n6076 gnd.n5184 24.8557
R14824 gnd.n5185 gnd.n5176 24.8557
R14825 gnd.n6112 gnd.n5168 24.8557
R14826 gnd.n6123 gnd.n5161 24.8557
R14827 gnd.n6122 gnd.n5149 24.8557
R14828 gnd.n5152 gnd.n5141 24.8557
R14829 gnd.n6410 gnd.n5142 24.8557
R14830 gnd.n6421 gnd.n5130 24.8557
R14831 gnd.n5771 gnd.t270 23.2624
R14832 gnd.t51 gnd.n1285 23.2624
R14833 gnd.n222 gnd.t189 23.2624
R14834 gnd.n5763 gnd.t332 22.6251
R14835 gnd.t137 gnd.n1323 22.6251
R14836 gnd.n184 gnd.t27 22.6251
R14837 gnd.n4166 gnd.n2126 22.3064
R14838 gnd.t22 gnd.n1361 21.9878
R14839 gnd.n146 gnd.t24 21.9878
R14840 gnd.n3487 gnd.n1698 21.6691
R14841 gnd.n3516 gnd.n2507 21.6691
R14842 gnd.n3588 gnd.n2448 21.6691
R14843 gnd.n3595 gnd.n2441 21.6691
R14844 gnd.n3630 gnd.n2422 21.6691
R14845 gnd.n3688 gnd.n2393 21.6691
R14846 gnd.n3696 gnd.n3695 21.6691
R14847 gnd.n3727 gnd.n2380 21.6691
R14848 gnd.n3738 gnd.n2375 21.6691
R14849 gnd.n3784 gnd.n2354 21.6691
R14850 gnd.n3790 gnd.n2350 21.6691
R14851 gnd.n3808 gnd.n2333 21.6691
R14852 gnd.n3820 gnd.n2321 21.6691
R14853 gnd.n3837 gnd.n2312 21.6691
R14854 gnd.n3848 gnd.n2289 21.6691
R14855 gnd.n3910 gnd.n2281 21.6691
R14856 gnd.n4004 gnd.n2223 21.6691
R14857 gnd.n5743 gnd.t207 21.3504
R14858 gnd.t139 gnd.n1398 21.3504
R14859 gnd.n2869 gnd.n2660 21.3504
R14860 gnd.n2891 gnd.t12 21.3504
R14861 gnd.n7465 gnd.t141 21.3504
R14862 gnd.n494 gnd.n485 21.3504
R14863 gnd.n7757 gnd.t63 21.3504
R14864 gnd.n2470 gnd.n2456 21.0318
R14865 gnd.n2374 gnd.n2362 21.0318
R14866 gnd.n2366 gnd.n2363 21.0318
R14867 gnd.n3921 gnd.n2276 21.0318
R14868 gnd.t128 gnd.n6100 20.7131
R14869 gnd.n1386 gnd.t39 20.7131
R14870 gnd.t49 gnd.n1626 20.7131
R14871 gnd.n2127 gnd.t230 20.7131
R14872 gnd.t196 gnd.n120 20.7131
R14873 gnd.t108 gnd.n2497 20.3945
R14874 gnd.n2244 gnd.t116 20.3945
R14875 gnd.n6022 gnd.t130 20.0758
R14876 gnd.n1349 gnd.t4 20.0758
R14877 gnd.t135 gnd.n159 20.0758
R14878 gnd.n3408 gnd.n3407 19.9763
R14879 gnd.n2189 gnd.n2188 19.9763
R14880 gnd.n4692 gnd.n4691 19.9763
R14881 gnd.n2183 gnd.n2182 19.9763
R14882 gnd.n1667 gnd.t291 19.8005
R14883 gnd.n1667 gnd.t363 19.8005
R14884 gnd.n1666 gnd.t330 19.8005
R14885 gnd.n1666 gnd.t354 19.8005
R14886 gnd.n2152 gnd.t284 19.8005
R14887 gnd.n2152 gnd.t398 19.8005
R14888 gnd.n2151 gnd.t344 19.8005
R14889 gnd.n2151 gnd.t324 19.8005
R14890 gnd.n4686 gnd.n4685 19.7572
R14891 gnd.n3405 gnd.t290 19.7572
R14892 gnd.n3558 gnd.t85 19.7572
R14893 gnd.n3574 gnd.n2475 19.7572
R14894 gnd.n3726 gnd.n3725 19.7572
R14895 gnd.n3791 gnd.n2347 19.7572
R14896 gnd.n3854 gnd.n2266 19.7572
R14897 gnd.n3973 gnd.t91 19.7572
R14898 gnd.n4158 gnd.n4157 19.7572
R14899 gnd.n6577 gnd.n6576 19.5706
R14900 gnd.n1663 gnd.n1662 19.5087
R14901 gnd.n1676 gnd.n1663 19.5087
R14902 gnd.n1674 gnd.n1665 19.5087
R14903 gnd.n2156 gnd.n2150 19.5087
R14904 gnd.t132 gnd.n5259 19.4385
R14905 gnd.n1311 gnd.t16 19.4385
R14906 gnd.n3339 gnd.n2549 19.3944
R14907 gnd.n3339 gnd.n2546 19.3944
R14908 gnd.n3360 gnd.n2546 19.3944
R14909 gnd.n3360 gnd.n2547 19.3944
R14910 gnd.n3356 gnd.n2547 19.3944
R14911 gnd.n3356 gnd.n3355 19.3944
R14912 gnd.n3355 gnd.n3354 19.3944
R14913 gnd.n3354 gnd.n3345 19.3944
R14914 gnd.n3350 gnd.n3345 19.3944
R14915 gnd.n3350 gnd.n3349 19.3944
R14916 gnd.n3349 gnd.n1701 19.3944
R14917 gnd.n4677 gnd.n1701 19.3944
R14918 gnd.n4677 gnd.n1702 19.3944
R14919 gnd.n4673 gnd.n1702 19.3944
R14920 gnd.n4673 gnd.n4672 19.3944
R14921 gnd.n4672 gnd.n4671 19.3944
R14922 gnd.n4671 gnd.n1708 19.3944
R14923 gnd.n4667 gnd.n1708 19.3944
R14924 gnd.n4667 gnd.n4666 19.3944
R14925 gnd.n4666 gnd.n4665 19.3944
R14926 gnd.n4665 gnd.n1713 19.3944
R14927 gnd.n4661 gnd.n1713 19.3944
R14928 gnd.n4661 gnd.n4660 19.3944
R14929 gnd.n4660 gnd.n4659 19.3944
R14930 gnd.n4659 gnd.n1718 19.3944
R14931 gnd.n4655 gnd.n1718 19.3944
R14932 gnd.n4655 gnd.n4654 19.3944
R14933 gnd.n4654 gnd.n4653 19.3944
R14934 gnd.n4653 gnd.n1723 19.3944
R14935 gnd.n4649 gnd.n1723 19.3944
R14936 gnd.n4649 gnd.n4648 19.3944
R14937 gnd.n4648 gnd.n4647 19.3944
R14938 gnd.n4647 gnd.n1728 19.3944
R14939 gnd.n4643 gnd.n1728 19.3944
R14940 gnd.n4643 gnd.n4642 19.3944
R14941 gnd.n4642 gnd.n4641 19.3944
R14942 gnd.n4641 gnd.n1733 19.3944
R14943 gnd.n4637 gnd.n1733 19.3944
R14944 gnd.n4637 gnd.n4636 19.3944
R14945 gnd.n4636 gnd.n4635 19.3944
R14946 gnd.n4635 gnd.n1738 19.3944
R14947 gnd.n4631 gnd.n1738 19.3944
R14948 gnd.n4631 gnd.n4630 19.3944
R14949 gnd.n4630 gnd.n4629 19.3944
R14950 gnd.n4629 gnd.n1743 19.3944
R14951 gnd.n4625 gnd.n1743 19.3944
R14952 gnd.n4625 gnd.n4624 19.3944
R14953 gnd.n4624 gnd.n4623 19.3944
R14954 gnd.n4623 gnd.n1748 19.3944
R14955 gnd.n4619 gnd.n1748 19.3944
R14956 gnd.n4619 gnd.n4618 19.3944
R14957 gnd.n4618 gnd.n4617 19.3944
R14958 gnd.n4617 gnd.n1753 19.3944
R14959 gnd.n4613 gnd.n1753 19.3944
R14960 gnd.n4613 gnd.n4612 19.3944
R14961 gnd.n4612 gnd.n4611 19.3944
R14962 gnd.n4611 gnd.n1758 19.3944
R14963 gnd.n4607 gnd.n1758 19.3944
R14964 gnd.n4607 gnd.n4606 19.3944
R14965 gnd.n4606 gnd.n4605 19.3944
R14966 gnd.n4605 gnd.n1763 19.3944
R14967 gnd.n4601 gnd.n1763 19.3944
R14968 gnd.n4601 gnd.n4600 19.3944
R14969 gnd.n4600 gnd.n4599 19.3944
R14970 gnd.n4599 gnd.n1768 19.3944
R14971 gnd.n4595 gnd.n1768 19.3944
R14972 gnd.n4595 gnd.n4594 19.3944
R14973 gnd.n4594 gnd.n4593 19.3944
R14974 gnd.n4593 gnd.n1773 19.3944
R14975 gnd.n4589 gnd.n1773 19.3944
R14976 gnd.n4589 gnd.n4588 19.3944
R14977 gnd.n4588 gnd.n4587 19.3944
R14978 gnd.n4587 gnd.n1778 19.3944
R14979 gnd.n4583 gnd.n1778 19.3944
R14980 gnd.n4583 gnd.n4582 19.3944
R14981 gnd.n4582 gnd.n4581 19.3944
R14982 gnd.n4581 gnd.n1783 19.3944
R14983 gnd.n4577 gnd.n1783 19.3944
R14984 gnd.n4577 gnd.n4576 19.3944
R14985 gnd.n4576 gnd.n4575 19.3944
R14986 gnd.n4575 gnd.n1788 19.3944
R14987 gnd.n4571 gnd.n1788 19.3944
R14988 gnd.n3124 gnd.n3123 19.3944
R14989 gnd.n3123 gnd.n2574 19.3944
R14990 gnd.n3326 gnd.n2574 19.3944
R14991 gnd.n3049 gnd.n3048 19.3944
R14992 gnd.n3052 gnd.n3049 19.3944
R14993 gnd.n3052 gnd.n3032 19.3944
R14994 gnd.n3056 gnd.n3032 19.3944
R14995 gnd.n3057 gnd.n3056 19.3944
R14996 gnd.n3173 gnd.n3057 19.3944
R14997 gnd.n3173 gnd.n3172 19.3944
R14998 gnd.n3172 gnd.n3171 19.3944
R14999 gnd.n3171 gnd.n3062 19.3944
R15000 gnd.n3164 gnd.n3062 19.3944
R15001 gnd.n3164 gnd.n3163 19.3944
R15002 gnd.n3163 gnd.n3071 19.3944
R15003 gnd.n3156 gnd.n3071 19.3944
R15004 gnd.n3156 gnd.n3155 19.3944
R15005 gnd.n3155 gnd.n3081 19.3944
R15006 gnd.n3148 gnd.n3081 19.3944
R15007 gnd.n3148 gnd.n3147 19.3944
R15008 gnd.n3147 gnd.n3091 19.3944
R15009 gnd.n3140 gnd.n3091 19.3944
R15010 gnd.n3140 gnd.n3139 19.3944
R15011 gnd.n3139 gnd.n3101 19.3944
R15012 gnd.n3132 gnd.n3101 19.3944
R15013 gnd.n3132 gnd.n3131 19.3944
R15014 gnd.n3131 gnd.n3111 19.3944
R15015 gnd.n4547 gnd.n1814 19.3944
R15016 gnd.n4547 gnd.n4546 19.3944
R15017 gnd.n4546 gnd.n1817 19.3944
R15018 gnd.n4539 gnd.n1817 19.3944
R15019 gnd.n4539 gnd.n4538 19.3944
R15020 gnd.n4538 gnd.n1825 19.3944
R15021 gnd.n4531 gnd.n1825 19.3944
R15022 gnd.n4531 gnd.n4530 19.3944
R15023 gnd.n4530 gnd.n1833 19.3944
R15024 gnd.n4523 gnd.n1833 19.3944
R15025 gnd.n4523 gnd.n4522 19.3944
R15026 gnd.n4522 gnd.n1841 19.3944
R15027 gnd.n4515 gnd.n1841 19.3944
R15028 gnd.n4515 gnd.n4514 19.3944
R15029 gnd.n4514 gnd.n1849 19.3944
R15030 gnd.n4507 gnd.n1849 19.3944
R15031 gnd.n5616 gnd.n5615 19.3944
R15032 gnd.n5615 gnd.n5525 19.3944
R15033 gnd.n5610 gnd.n5525 19.3944
R15034 gnd.n5610 gnd.n5609 19.3944
R15035 gnd.n5609 gnd.n5530 19.3944
R15036 gnd.n5604 gnd.n5530 19.3944
R15037 gnd.n5604 gnd.n5603 19.3944
R15038 gnd.n5603 gnd.n5602 19.3944
R15039 gnd.n5602 gnd.n5536 19.3944
R15040 gnd.n5596 gnd.n5536 19.3944
R15041 gnd.n5596 gnd.n5595 19.3944
R15042 gnd.n5595 gnd.n5594 19.3944
R15043 gnd.n5594 gnd.n5542 19.3944
R15044 gnd.n5588 gnd.n5542 19.3944
R15045 gnd.n5588 gnd.n5587 19.3944
R15046 gnd.n5587 gnd.n5586 19.3944
R15047 gnd.n5586 gnd.n5548 19.3944
R15048 gnd.n5580 gnd.n5548 19.3944
R15049 gnd.n5580 gnd.n5579 19.3944
R15050 gnd.n5579 gnd.n5578 19.3944
R15051 gnd.n5578 gnd.n5554 19.3944
R15052 gnd.n5572 gnd.n5554 19.3944
R15053 gnd.n5570 gnd.n5569 19.3944
R15054 gnd.n5569 gnd.n5564 19.3944
R15055 gnd.n5564 gnd.n5562 19.3944
R15056 gnd.n6503 gnd.n6428 19.3944
R15057 gnd.n6506 gnd.n6503 19.3944
R15058 gnd.n6508 gnd.n6506 19.3944
R15059 gnd.n6443 gnd.n6441 19.3944
R15060 gnd.n6446 gnd.n6443 19.3944
R15061 gnd.n6446 gnd.n6438 19.3944
R15062 gnd.n6450 gnd.n6438 19.3944
R15063 gnd.n6453 gnd.n6450 19.3944
R15064 gnd.n6456 gnd.n6453 19.3944
R15065 gnd.n6456 gnd.n6436 19.3944
R15066 gnd.n6460 gnd.n6436 19.3944
R15067 gnd.n6463 gnd.n6460 19.3944
R15068 gnd.n6466 gnd.n6463 19.3944
R15069 gnd.n6466 gnd.n6434 19.3944
R15070 gnd.n6470 gnd.n6434 19.3944
R15071 gnd.n6473 gnd.n6470 19.3944
R15072 gnd.n6476 gnd.n6473 19.3944
R15073 gnd.n6476 gnd.n6432 19.3944
R15074 gnd.n6480 gnd.n6432 19.3944
R15075 gnd.n6483 gnd.n6480 19.3944
R15076 gnd.n6486 gnd.n6483 19.3944
R15077 gnd.n6486 gnd.n6430 19.3944
R15078 gnd.n6490 gnd.n6430 19.3944
R15079 gnd.n6493 gnd.n6490 19.3944
R15080 gnd.n6499 gnd.n6493 19.3944
R15081 gnd.n5756 gnd.n5755 19.3944
R15082 gnd.n5757 gnd.n5756 19.3944
R15083 gnd.n5757 gnd.n5466 19.3944
R15084 gnd.n5466 gnd.n5460 19.3944
R15085 gnd.n5782 gnd.n5460 19.3944
R15086 gnd.n5783 gnd.n5782 19.3944
R15087 gnd.n5783 gnd.n5443 19.3944
R15088 gnd.n5443 gnd.n5441 19.3944
R15089 gnd.n5807 gnd.n5441 19.3944
R15090 gnd.n5810 gnd.n5807 19.3944
R15091 gnd.n5810 gnd.n5809 19.3944
R15092 gnd.n5809 gnd.n5413 19.3944
R15093 gnd.n5848 gnd.n5413 19.3944
R15094 gnd.n5848 gnd.n5411 19.3944
R15095 gnd.n5854 gnd.n5411 19.3944
R15096 gnd.n5855 gnd.n5854 19.3944
R15097 gnd.n5855 gnd.n5381 19.3944
R15098 gnd.n5905 gnd.n5381 19.3944
R15099 gnd.n5906 gnd.n5905 19.3944
R15100 gnd.n5906 gnd.n5374 19.3944
R15101 gnd.n5917 gnd.n5374 19.3944
R15102 gnd.n5918 gnd.n5917 19.3944
R15103 gnd.n5918 gnd.n5357 19.3944
R15104 gnd.n5357 gnd.n5355 19.3944
R15105 gnd.n5942 gnd.n5355 19.3944
R15106 gnd.n5943 gnd.n5942 19.3944
R15107 gnd.n5943 gnd.n5246 19.3944
R15108 gnd.n5987 gnd.n5246 19.3944
R15109 gnd.n5988 gnd.n5987 19.3944
R15110 gnd.n5988 gnd.n5239 19.3944
R15111 gnd.n5999 gnd.n5239 19.3944
R15112 gnd.n6001 gnd.n5999 19.3944
R15113 gnd.n6004 gnd.n6001 19.3944
R15114 gnd.n6004 gnd.n6003 19.3944
R15115 gnd.n6003 gnd.n5210 19.3944
R15116 gnd.n6044 gnd.n5210 19.3944
R15117 gnd.n6045 gnd.n6044 19.3944
R15118 gnd.n6045 gnd.n5194 19.3944
R15119 gnd.n5194 gnd.n5192 19.3944
R15120 gnd.n6069 gnd.n5192 19.3944
R15121 gnd.n6070 gnd.n6069 19.3944
R15122 gnd.n6070 gnd.n5164 19.3944
R15123 gnd.n6118 gnd.n5164 19.3944
R15124 gnd.n6119 gnd.n6118 19.3944
R15125 gnd.n6119 gnd.n5157 19.3944
R15126 gnd.n6130 gnd.n5157 19.3944
R15127 gnd.n6131 gnd.n6130 19.3944
R15128 gnd.n6131 gnd.n5140 19.3944
R15129 gnd.n5140 gnd.n5138 19.3944
R15130 gnd.n6414 gnd.n5138 19.3944
R15131 gnd.n6415 gnd.n6414 19.3944
R15132 gnd.n6415 gnd.n1126 19.3944
R15133 gnd.n6570 gnd.n1126 19.3944
R15134 gnd.n5739 gnd.n5738 19.3944
R15135 gnd.n5738 gnd.n5737 19.3944
R15136 gnd.n5737 gnd.n5736 19.3944
R15137 gnd.n5736 gnd.n5734 19.3944
R15138 gnd.n5734 gnd.n5731 19.3944
R15139 gnd.n5731 gnd.n5730 19.3944
R15140 gnd.n5730 gnd.n5727 19.3944
R15141 gnd.n5727 gnd.n5726 19.3944
R15142 gnd.n5726 gnd.n5723 19.3944
R15143 gnd.n5723 gnd.n5722 19.3944
R15144 gnd.n5722 gnd.n5719 19.3944
R15145 gnd.n5719 gnd.n5718 19.3944
R15146 gnd.n5718 gnd.n5715 19.3944
R15147 gnd.n5715 gnd.n5714 19.3944
R15148 gnd.n5765 gnd.n5471 19.3944
R15149 gnd.n5765 gnd.n5469 19.3944
R15150 gnd.n5769 gnd.n5469 19.3944
R15151 gnd.n5769 gnd.n5450 19.3944
R15152 gnd.n5795 gnd.n5450 19.3944
R15153 gnd.n5795 gnd.n5448 19.3944
R15154 gnd.n5801 gnd.n5448 19.3944
R15155 gnd.n5801 gnd.n5800 19.3944
R15156 gnd.n5800 gnd.n5424 19.3944
R15157 gnd.n5829 gnd.n5424 19.3944
R15158 gnd.n5829 gnd.n5422 19.3944
R15159 gnd.n5838 gnd.n5422 19.3944
R15160 gnd.n5838 gnd.n5837 19.3944
R15161 gnd.n5837 gnd.n5836 19.3944
R15162 gnd.n5836 gnd.n5391 19.3944
R15163 gnd.n5890 gnd.n5391 19.3944
R15164 gnd.n5890 gnd.n5389 19.3944
R15165 gnd.n5896 gnd.n5389 19.3944
R15166 gnd.n5896 gnd.n5895 19.3944
R15167 gnd.n5895 gnd.n5364 19.3944
R15168 gnd.n5930 gnd.n5364 19.3944
R15169 gnd.n5930 gnd.n5362 19.3944
R15170 gnd.n5936 gnd.n5362 19.3944
R15171 gnd.n5936 gnd.n5935 19.3944
R15172 gnd.n5935 gnd.n5257 19.3944
R15173 gnd.n5972 gnd.n5257 19.3944
R15174 gnd.n5972 gnd.n5255 19.3944
R15175 gnd.n5978 gnd.n5255 19.3944
R15176 gnd.n5978 gnd.n5977 19.3944
R15177 gnd.n5977 gnd.n5227 19.3944
R15178 gnd.n6013 gnd.n5227 19.3944
R15179 gnd.n6013 gnd.n5225 19.3944
R15180 gnd.n6019 gnd.n5225 19.3944
R15181 gnd.n6019 gnd.n6018 19.3944
R15182 gnd.n6018 gnd.n5201 19.3944
R15183 gnd.n6057 gnd.n5201 19.3944
R15184 gnd.n6057 gnd.n5199 19.3944
R15185 gnd.n6063 gnd.n5199 19.3944
R15186 gnd.n6063 gnd.n6062 19.3944
R15187 gnd.n6062 gnd.n5174 19.3944
R15188 gnd.n6103 gnd.n5174 19.3944
R15189 gnd.n6103 gnd.n5172 19.3944
R15190 gnd.n6109 gnd.n5172 19.3944
R15191 gnd.n6109 gnd.n6108 19.3944
R15192 gnd.n6108 gnd.n5147 19.3944
R15193 gnd.n6399 gnd.n5147 19.3944
R15194 gnd.n6399 gnd.n5145 19.3944
R15195 gnd.n6408 gnd.n5145 19.3944
R15196 gnd.n6408 gnd.n6407 19.3944
R15197 gnd.n6407 gnd.n6406 19.3944
R15198 gnd.n6406 gnd.n5121 19.3944
R15199 gnd.n6518 gnd.n5121 19.3944
R15200 gnd.n6519 gnd.n6518 19.3944
R15201 gnd.n6557 gnd.n6556 19.3944
R15202 gnd.n6556 gnd.n6522 19.3944
R15203 gnd.n6552 gnd.n6522 19.3944
R15204 gnd.n6552 gnd.n6549 19.3944
R15205 gnd.n6549 gnd.n6546 19.3944
R15206 gnd.n6546 gnd.n6545 19.3944
R15207 gnd.n6545 gnd.n6542 19.3944
R15208 gnd.n6542 gnd.n6541 19.3944
R15209 gnd.n6541 gnd.n6538 19.3944
R15210 gnd.n6538 gnd.n6537 19.3944
R15211 gnd.n6537 gnd.n6534 19.3944
R15212 gnd.n6534 gnd.n6533 19.3944
R15213 gnd.n6533 gnd.n1133 19.3944
R15214 gnd.n6563 gnd.n1133 19.3944
R15215 gnd.n5623 gnd.n5519 19.3944
R15216 gnd.n5627 gnd.n5519 19.3944
R15217 gnd.n5627 gnd.n5509 19.3944
R15218 gnd.n5639 gnd.n5509 19.3944
R15219 gnd.n5639 gnd.n5507 19.3944
R15220 gnd.n5643 gnd.n5507 19.3944
R15221 gnd.n5643 gnd.n5496 19.3944
R15222 gnd.n5655 gnd.n5496 19.3944
R15223 gnd.n5655 gnd.n5494 19.3944
R15224 gnd.n5681 gnd.n5494 19.3944
R15225 gnd.n5681 gnd.n5680 19.3944
R15226 gnd.n5680 gnd.n5679 19.3944
R15227 gnd.n5679 gnd.n5678 19.3944
R15228 gnd.n5678 gnd.n5676 19.3944
R15229 gnd.n5676 gnd.n5675 19.3944
R15230 gnd.n5675 gnd.n5673 19.3944
R15231 gnd.n5673 gnd.n5672 19.3944
R15232 gnd.n5672 gnd.n5670 19.3944
R15233 gnd.n5670 gnd.n5669 19.3944
R15234 gnd.n5669 gnd.n5431 19.3944
R15235 gnd.n5818 gnd.n5431 19.3944
R15236 gnd.n5818 gnd.n5429 19.3944
R15237 gnd.n5824 gnd.n5429 19.3944
R15238 gnd.n5824 gnd.n5823 19.3944
R15239 gnd.n5823 gnd.n5398 19.3944
R15240 gnd.n5865 gnd.n5398 19.3944
R15241 gnd.n5865 gnd.n5396 19.3944
R15242 gnd.n5869 gnd.n5396 19.3944
R15243 gnd.n5883 gnd.n5869 19.3944
R15244 gnd.n5881 gnd.n5880 19.3944
R15245 gnd.n5877 gnd.n5876 19.3944
R15246 gnd.n5873 gnd.n5872 19.3944
R15247 gnd.n5951 gnd.n5345 19.3944
R15248 gnd.n5951 gnd.n5263 19.3944
R15249 gnd.n5967 gnd.n5263 19.3944
R15250 gnd.n5967 gnd.n5966 19.3944
R15251 gnd.n5966 gnd.n5965 19.3944
R15252 gnd.n5965 gnd.n5963 19.3944
R15253 gnd.n5963 gnd.n5962 19.3944
R15254 gnd.n5962 gnd.n5960 19.3944
R15255 gnd.n5960 gnd.n5219 19.3944
R15256 gnd.n6024 gnd.n5219 19.3944
R15257 gnd.n6024 gnd.n5217 19.3944
R15258 gnd.n6033 gnd.n5217 19.3944
R15259 gnd.n6033 gnd.n6032 19.3944
R15260 gnd.n6032 gnd.n6031 19.3944
R15261 gnd.n6031 gnd.n5182 19.3944
R15262 gnd.n6078 gnd.n5182 19.3944
R15263 gnd.n6078 gnd.n5180 19.3944
R15264 gnd.n6098 gnd.n5180 19.3944
R15265 gnd.n6098 gnd.n6097 19.3944
R15266 gnd.n6097 gnd.n6096 19.3944
R15267 gnd.n6096 gnd.n6093 19.3944
R15268 gnd.n6093 gnd.n6092 19.3944
R15269 gnd.n6092 gnd.n6090 19.3944
R15270 gnd.n6090 gnd.n6089 19.3944
R15271 gnd.n6089 gnd.n5128 19.3944
R15272 gnd.n6423 gnd.n5128 19.3944
R15273 gnd.n6423 gnd.n5126 19.3944
R15274 gnd.n6512 gnd.n5126 19.3944
R15275 gnd.n6512 gnd.n6511 19.3944
R15276 gnd.n5619 gnd.n5515 19.3944
R15277 gnd.n5631 gnd.n5515 19.3944
R15278 gnd.n5631 gnd.n5513 19.3944
R15279 gnd.n5635 gnd.n5513 19.3944
R15280 gnd.n5635 gnd.n5503 19.3944
R15281 gnd.n5647 gnd.n5503 19.3944
R15282 gnd.n5647 gnd.n5501 19.3944
R15283 gnd.n5651 gnd.n5501 19.3944
R15284 gnd.n5651 gnd.n5490 19.3944
R15285 gnd.n5745 gnd.n5490 19.3944
R15286 gnd.n5745 gnd.n5487 19.3944
R15287 gnd.n5750 gnd.n5487 19.3944
R15288 gnd.n5750 gnd.n5478 19.3944
R15289 gnd.n5760 gnd.n5478 19.3944
R15290 gnd.n5760 gnd.n5462 19.3944
R15291 gnd.n5777 gnd.n5462 19.3944
R15292 gnd.n5777 gnd.n5458 19.3944
R15293 gnd.n5790 gnd.n5458 19.3944
R15294 gnd.n5790 gnd.n5789 19.3944
R15295 gnd.n5789 gnd.n5437 19.3944
R15296 gnd.n5814 gnd.n5437 19.3944
R15297 gnd.n5814 gnd.n5813 19.3944
R15298 gnd.n5813 gnd.n5415 19.3944
R15299 gnd.n5843 gnd.n5415 19.3944
R15300 gnd.n5843 gnd.n5405 19.3944
R15301 gnd.n5861 gnd.n5405 19.3944
R15302 gnd.n5861 gnd.n5860 19.3944
R15303 gnd.n5860 gnd.n5859 19.3944
R15304 gnd.n5859 gnd.n5383 19.3944
R15305 gnd.n5901 gnd.n5383 19.3944
R15306 gnd.n5901 gnd.n5376 19.3944
R15307 gnd.n5912 gnd.n5376 19.3944
R15308 gnd.n5912 gnd.n5372 19.3944
R15309 gnd.n5925 gnd.n5372 19.3944
R15310 gnd.n5925 gnd.n5924 19.3944
R15311 gnd.n5924 gnd.n5351 19.3944
R15312 gnd.n5947 gnd.n5351 19.3944
R15313 gnd.n5947 gnd.n5946 19.3944
R15314 gnd.n5946 gnd.n5248 19.3944
R15315 gnd.n5983 gnd.n5248 19.3944
R15316 gnd.n5983 gnd.n5241 19.3944
R15317 gnd.n5994 gnd.n5241 19.3944
R15318 gnd.n5994 gnd.n5235 19.3944
R15319 gnd.n6008 gnd.n5235 19.3944
R15320 gnd.n6008 gnd.n6007 19.3944
R15321 gnd.n6007 gnd.n5212 19.3944
R15322 gnd.n6039 gnd.n5212 19.3944
R15323 gnd.n6039 gnd.n5208 19.3944
R15324 gnd.n6052 gnd.n5208 19.3944
R15325 gnd.n6052 gnd.n6051 19.3944
R15326 gnd.n6051 gnd.n5188 19.3944
R15327 gnd.n6074 gnd.n5188 19.3944
R15328 gnd.n6074 gnd.n6073 19.3944
R15329 gnd.n6073 gnd.n5166 19.3944
R15330 gnd.n6114 gnd.n5166 19.3944
R15331 gnd.n6114 gnd.n5159 19.3944
R15332 gnd.n6125 gnd.n5159 19.3944
R15333 gnd.n6125 gnd.n5155 19.3944
R15334 gnd.n6394 gnd.n5155 19.3944
R15335 gnd.n6394 gnd.n6393 19.3944
R15336 gnd.n6393 gnd.n5134 19.3944
R15337 gnd.n6419 gnd.n5134 19.3944
R15338 gnd.n6419 gnd.n6418 19.3944
R15339 gnd.n6418 gnd.n1123 19.3944
R15340 gnd.n6573 gnd.n1123 19.3944
R15341 gnd.n3168 gnd.n3167 19.3944
R15342 gnd.n3167 gnd.n3065 19.3944
R15343 gnd.n3160 gnd.n3065 19.3944
R15344 gnd.n3160 gnd.n3159 19.3944
R15345 gnd.n3159 gnd.n3077 19.3944
R15346 gnd.n3152 gnd.n3077 19.3944
R15347 gnd.n3152 gnd.n3151 19.3944
R15348 gnd.n3151 gnd.n3085 19.3944
R15349 gnd.n3144 gnd.n3085 19.3944
R15350 gnd.n3144 gnd.n3143 19.3944
R15351 gnd.n3143 gnd.n3097 19.3944
R15352 gnd.n3136 gnd.n3097 19.3944
R15353 gnd.n3136 gnd.n3135 19.3944
R15354 gnd.n3135 gnd.n3105 19.3944
R15355 gnd.n3128 gnd.n3105 19.3944
R15356 gnd.n3128 gnd.n3127 19.3944
R15357 gnd.n2655 gnd.n2639 19.3944
R15358 gnd.n2903 gnd.n2639 19.3944
R15359 gnd.n2903 gnd.n2637 19.3944
R15360 gnd.n2927 gnd.n2637 19.3944
R15361 gnd.n2927 gnd.n2926 19.3944
R15362 gnd.n2926 gnd.n2925 19.3944
R15363 gnd.n2925 gnd.n2909 19.3944
R15364 gnd.n2921 gnd.n2909 19.3944
R15365 gnd.n2921 gnd.n2920 19.3944
R15366 gnd.n2920 gnd.n2919 19.3944
R15367 gnd.n2919 gnd.n2917 19.3944
R15368 gnd.n2917 gnd.n2614 19.3944
R15369 gnd.n2614 gnd.n2612 19.3944
R15370 gnd.n2992 gnd.n2612 19.3944
R15371 gnd.n2992 gnd.n2610 19.3944
R15372 gnd.n2996 gnd.n2610 19.3944
R15373 gnd.n2996 gnd.n2608 19.3944
R15374 gnd.n3000 gnd.n2608 19.3944
R15375 gnd.n3000 gnd.n2606 19.3944
R15376 gnd.n3008 gnd.n2606 19.3944
R15377 gnd.n3008 gnd.n3007 19.3944
R15378 gnd.n3007 gnd.n3006 19.3944
R15379 gnd.n3006 gnd.n2590 19.3944
R15380 gnd.n3295 gnd.n2590 19.3944
R15381 gnd.n3295 gnd.n2588 19.3944
R15382 gnd.n3299 gnd.n2588 19.3944
R15383 gnd.n3299 gnd.n2586 19.3944
R15384 gnd.n3303 gnd.n2586 19.3944
R15385 gnd.n3303 gnd.n2584 19.3944
R15386 gnd.n3315 gnd.n2584 19.3944
R15387 gnd.n3315 gnd.n3314 19.3944
R15388 gnd.n3314 gnd.n3313 19.3944
R15389 gnd.n3313 gnd.n3310 19.3944
R15390 gnd.n3310 gnd.n2556 19.3944
R15391 gnd.n3331 gnd.n2556 19.3944
R15392 gnd.n3331 gnd.n2554 19.3944
R15393 gnd.n3335 gnd.n2554 19.3944
R15394 gnd.n3335 gnd.n2540 19.3944
R15395 gnd.n3364 gnd.n2540 19.3944
R15396 gnd.n3364 gnd.n2538 19.3944
R15397 gnd.n3377 gnd.n2538 19.3944
R15398 gnd.n3377 gnd.n3376 19.3944
R15399 gnd.n3376 gnd.n3375 19.3944
R15400 gnd.n3375 gnd.n3372 19.3944
R15401 gnd.n3372 gnd.n1691 19.3944
R15402 gnd.n4683 gnd.n1691 19.3944
R15403 gnd.n4683 gnd.n4682 19.3944
R15404 gnd.n4682 gnd.n4681 19.3944
R15405 gnd.n4681 gnd.n1695 19.3944
R15406 gnd.n2505 gnd.n1695 19.3944
R15407 gnd.n3530 gnd.n2505 19.3944
R15408 gnd.n3530 gnd.n2502 19.3944
R15409 gnd.n3536 gnd.n2502 19.3944
R15410 gnd.n3536 gnd.n3535 19.3944
R15411 gnd.n3535 gnd.n2482 19.3944
R15412 gnd.n3567 gnd.n2482 19.3944
R15413 gnd.n3567 gnd.n2480 19.3944
R15414 gnd.n3571 gnd.n2480 19.3944
R15415 gnd.n3571 gnd.n2454 19.3944
R15416 gnd.n3606 gnd.n2454 19.3944
R15417 gnd.n3606 gnd.n2452 19.3944
R15418 gnd.n3612 gnd.n2452 19.3944
R15419 gnd.n3612 gnd.n3611 19.3944
R15420 gnd.n3611 gnd.n2426 19.3944
R15421 gnd.n3646 gnd.n2426 19.3944
R15422 gnd.n3646 gnd.n2424 19.3944
R15423 gnd.n3651 gnd.n2424 19.3944
R15424 gnd.n3651 gnd.n2405 19.3944
R15425 gnd.n3679 gnd.n2405 19.3944
R15426 gnd.n3679 gnd.n3678 19.3944
R15427 gnd.n3678 gnd.n3677 19.3944
R15428 gnd.n3677 gnd.n2409 19.3944
R15429 gnd.n2412 gnd.n2409 19.3944
R15430 gnd.n2412 gnd.n2370 19.3944
R15431 gnd.n3741 gnd.n2370 19.3944
R15432 gnd.n3741 gnd.n2368 19.3944
R15433 gnd.n3747 gnd.n2368 19.3944
R15434 gnd.n3747 gnd.n3746 19.3944
R15435 gnd.n3746 gnd.n2345 19.3944
R15436 gnd.n3793 gnd.n2345 19.3944
R15437 gnd.n3793 gnd.n2343 19.3944
R15438 gnd.n3799 gnd.n2343 19.3944
R15439 gnd.n3799 gnd.n3798 19.3944
R15440 gnd.n3798 gnd.n2319 19.3944
R15441 gnd.n3830 gnd.n2319 19.3944
R15442 gnd.n3830 gnd.n2317 19.3944
R15443 gnd.n3834 gnd.n2317 19.3944
R15444 gnd.n3834 gnd.n2294 19.3944
R15445 gnd.n3891 gnd.n2294 19.3944
R15446 gnd.n3891 gnd.n2292 19.3944
R15447 gnd.n3897 gnd.n2292 19.3944
R15448 gnd.n3897 gnd.n3896 19.3944
R15449 gnd.n3896 gnd.n2271 19.3944
R15450 gnd.n3924 gnd.n2271 19.3944
R15451 gnd.n3924 gnd.n2269 19.3944
R15452 gnd.n3930 gnd.n2269 19.3944
R15453 gnd.n3930 gnd.n3929 19.3944
R15454 gnd.n3929 gnd.n2250 19.3944
R15455 gnd.n3976 gnd.n2250 19.3944
R15456 gnd.n3976 gnd.n2248 19.3944
R15457 gnd.n3982 gnd.n2248 19.3944
R15458 gnd.n3982 gnd.n3981 19.3944
R15459 gnd.n3981 gnd.n2221 19.3944
R15460 gnd.n4013 gnd.n2221 19.3944
R15461 gnd.n4013 gnd.n2219 19.3944
R15462 gnd.n4017 gnd.n2219 19.3944
R15463 gnd.n4017 gnd.n2132 19.3944
R15464 gnd.n4160 gnd.n2132 19.3944
R15465 gnd.n4160 gnd.n2130 19.3944
R15466 gnd.n4164 gnd.n2130 19.3944
R15467 gnd.n4164 gnd.n2119 19.3944
R15468 gnd.n4176 gnd.n2119 19.3944
R15469 gnd.n4176 gnd.n2117 19.3944
R15470 gnd.n4183 gnd.n2117 19.3944
R15471 gnd.n4183 gnd.n4182 19.3944
R15472 gnd.n4182 gnd.n2106 19.3944
R15473 gnd.n4196 gnd.n2106 19.3944
R15474 gnd.n4197 gnd.n4196 19.3944
R15475 gnd.n4197 gnd.n2104 19.3944
R15476 gnd.n4249 gnd.n2104 19.3944
R15477 gnd.n4249 gnd.n4248 19.3944
R15478 gnd.n4248 gnd.n4247 19.3944
R15479 gnd.n4247 gnd.n4203 19.3944
R15480 gnd.n4243 gnd.n4203 19.3944
R15481 gnd.n4243 gnd.n4242 19.3944
R15482 gnd.n4242 gnd.n4241 19.3944
R15483 gnd.n4241 gnd.n4209 19.3944
R15484 gnd.n4235 gnd.n4209 19.3944
R15485 gnd.n4235 gnd.n4234 19.3944
R15486 gnd.n4234 gnd.n4233 19.3944
R15487 gnd.n4233 gnd.n4215 19.3944
R15488 gnd.n4229 gnd.n4215 19.3944
R15489 gnd.n4229 gnd.n4228 19.3944
R15490 gnd.n4228 gnd.n4227 19.3944
R15491 gnd.n4227 gnd.n4224 19.3944
R15492 gnd.n4224 gnd.n4223 19.3944
R15493 gnd.n4223 gnd.n2059 19.3944
R15494 gnd.n4320 gnd.n2059 19.3944
R15495 gnd.n4320 gnd.n2057 19.3944
R15496 gnd.n4325 gnd.n2057 19.3944
R15497 gnd.n4325 gnd.n576 19.3944
R15498 gnd.n7367 gnd.n576 19.3944
R15499 gnd.n7367 gnd.n7366 19.3944
R15500 gnd.n7366 gnd.n7365 19.3944
R15501 gnd.n7365 gnd.n580 19.3944
R15502 gnd.n7361 gnd.n580 19.3944
R15503 gnd.n7361 gnd.n7360 19.3944
R15504 gnd.n7360 gnd.n7359 19.3944
R15505 gnd.n7359 gnd.n586 19.3944
R15506 gnd.n7355 gnd.n586 19.3944
R15507 gnd.n7355 gnd.n7354 19.3944
R15508 gnd.n7354 gnd.n7353 19.3944
R15509 gnd.n7353 gnd.n7350 19.3944
R15510 gnd.n7350 gnd.n592 19.3944
R15511 gnd.n7133 gnd.n716 19.3944
R15512 gnd.n7139 gnd.n716 19.3944
R15513 gnd.n7139 gnd.n714 19.3944
R15514 gnd.n7143 gnd.n714 19.3944
R15515 gnd.n7143 gnd.n710 19.3944
R15516 gnd.n7149 gnd.n710 19.3944
R15517 gnd.n7149 gnd.n708 19.3944
R15518 gnd.n7153 gnd.n708 19.3944
R15519 gnd.n7153 gnd.n704 19.3944
R15520 gnd.n7159 gnd.n704 19.3944
R15521 gnd.n7159 gnd.n702 19.3944
R15522 gnd.n7163 gnd.n702 19.3944
R15523 gnd.n7163 gnd.n698 19.3944
R15524 gnd.n7169 gnd.n698 19.3944
R15525 gnd.n7169 gnd.n696 19.3944
R15526 gnd.n7173 gnd.n696 19.3944
R15527 gnd.n7173 gnd.n692 19.3944
R15528 gnd.n7179 gnd.n692 19.3944
R15529 gnd.n7179 gnd.n690 19.3944
R15530 gnd.n7183 gnd.n690 19.3944
R15531 gnd.n7183 gnd.n686 19.3944
R15532 gnd.n7189 gnd.n686 19.3944
R15533 gnd.n7189 gnd.n684 19.3944
R15534 gnd.n7193 gnd.n684 19.3944
R15535 gnd.n7193 gnd.n680 19.3944
R15536 gnd.n7199 gnd.n680 19.3944
R15537 gnd.n7199 gnd.n678 19.3944
R15538 gnd.n7203 gnd.n678 19.3944
R15539 gnd.n7203 gnd.n674 19.3944
R15540 gnd.n7209 gnd.n674 19.3944
R15541 gnd.n7209 gnd.n672 19.3944
R15542 gnd.n7213 gnd.n672 19.3944
R15543 gnd.n7213 gnd.n668 19.3944
R15544 gnd.n7219 gnd.n668 19.3944
R15545 gnd.n7219 gnd.n666 19.3944
R15546 gnd.n7223 gnd.n666 19.3944
R15547 gnd.n7223 gnd.n662 19.3944
R15548 gnd.n7229 gnd.n662 19.3944
R15549 gnd.n7229 gnd.n660 19.3944
R15550 gnd.n7233 gnd.n660 19.3944
R15551 gnd.n7233 gnd.n656 19.3944
R15552 gnd.n7239 gnd.n656 19.3944
R15553 gnd.n7239 gnd.n654 19.3944
R15554 gnd.n7243 gnd.n654 19.3944
R15555 gnd.n7243 gnd.n650 19.3944
R15556 gnd.n7249 gnd.n650 19.3944
R15557 gnd.n7249 gnd.n648 19.3944
R15558 gnd.n7253 gnd.n648 19.3944
R15559 gnd.n7253 gnd.n644 19.3944
R15560 gnd.n7259 gnd.n644 19.3944
R15561 gnd.n7259 gnd.n642 19.3944
R15562 gnd.n7263 gnd.n642 19.3944
R15563 gnd.n7263 gnd.n638 19.3944
R15564 gnd.n7269 gnd.n638 19.3944
R15565 gnd.n7269 gnd.n636 19.3944
R15566 gnd.n7273 gnd.n636 19.3944
R15567 gnd.n7273 gnd.n632 19.3944
R15568 gnd.n7279 gnd.n632 19.3944
R15569 gnd.n7279 gnd.n630 19.3944
R15570 gnd.n7283 gnd.n630 19.3944
R15571 gnd.n7283 gnd.n626 19.3944
R15572 gnd.n7289 gnd.n626 19.3944
R15573 gnd.n7289 gnd.n624 19.3944
R15574 gnd.n7293 gnd.n624 19.3944
R15575 gnd.n7293 gnd.n620 19.3944
R15576 gnd.n7299 gnd.n620 19.3944
R15577 gnd.n7299 gnd.n618 19.3944
R15578 gnd.n7303 gnd.n618 19.3944
R15579 gnd.n7303 gnd.n614 19.3944
R15580 gnd.n7309 gnd.n614 19.3944
R15581 gnd.n7309 gnd.n612 19.3944
R15582 gnd.n7313 gnd.n612 19.3944
R15583 gnd.n7313 gnd.n608 19.3944
R15584 gnd.n7319 gnd.n608 19.3944
R15585 gnd.n7319 gnd.n606 19.3944
R15586 gnd.n7323 gnd.n606 19.3944
R15587 gnd.n7323 gnd.n602 19.3944
R15588 gnd.n7329 gnd.n602 19.3944
R15589 gnd.n7329 gnd.n600 19.3944
R15590 gnd.n7333 gnd.n600 19.3944
R15591 gnd.n7333 gnd.n596 19.3944
R15592 gnd.n7341 gnd.n596 19.3944
R15593 gnd.n7341 gnd.n594 19.3944
R15594 gnd.n7346 gnd.n594 19.3944
R15595 gnd.n6748 gnd.n949 19.3944
R15596 gnd.n6748 gnd.n947 19.3944
R15597 gnd.n6752 gnd.n947 19.3944
R15598 gnd.n6752 gnd.n943 19.3944
R15599 gnd.n6758 gnd.n943 19.3944
R15600 gnd.n6758 gnd.n941 19.3944
R15601 gnd.n6762 gnd.n941 19.3944
R15602 gnd.n6762 gnd.n937 19.3944
R15603 gnd.n6768 gnd.n937 19.3944
R15604 gnd.n6768 gnd.n935 19.3944
R15605 gnd.n6772 gnd.n935 19.3944
R15606 gnd.n6772 gnd.n931 19.3944
R15607 gnd.n6778 gnd.n931 19.3944
R15608 gnd.n6778 gnd.n929 19.3944
R15609 gnd.n6782 gnd.n929 19.3944
R15610 gnd.n6782 gnd.n925 19.3944
R15611 gnd.n6788 gnd.n925 19.3944
R15612 gnd.n6788 gnd.n923 19.3944
R15613 gnd.n6792 gnd.n923 19.3944
R15614 gnd.n6792 gnd.n919 19.3944
R15615 gnd.n6798 gnd.n919 19.3944
R15616 gnd.n6798 gnd.n917 19.3944
R15617 gnd.n6802 gnd.n917 19.3944
R15618 gnd.n6802 gnd.n913 19.3944
R15619 gnd.n6808 gnd.n913 19.3944
R15620 gnd.n6808 gnd.n911 19.3944
R15621 gnd.n6812 gnd.n911 19.3944
R15622 gnd.n6812 gnd.n907 19.3944
R15623 gnd.n6818 gnd.n907 19.3944
R15624 gnd.n6818 gnd.n905 19.3944
R15625 gnd.n6822 gnd.n905 19.3944
R15626 gnd.n6822 gnd.n901 19.3944
R15627 gnd.n6828 gnd.n901 19.3944
R15628 gnd.n6828 gnd.n899 19.3944
R15629 gnd.n6832 gnd.n899 19.3944
R15630 gnd.n6832 gnd.n895 19.3944
R15631 gnd.n6838 gnd.n895 19.3944
R15632 gnd.n6838 gnd.n893 19.3944
R15633 gnd.n6842 gnd.n893 19.3944
R15634 gnd.n6842 gnd.n889 19.3944
R15635 gnd.n6848 gnd.n889 19.3944
R15636 gnd.n6848 gnd.n887 19.3944
R15637 gnd.n6852 gnd.n887 19.3944
R15638 gnd.n6852 gnd.n883 19.3944
R15639 gnd.n6858 gnd.n883 19.3944
R15640 gnd.n6858 gnd.n881 19.3944
R15641 gnd.n6862 gnd.n881 19.3944
R15642 gnd.n6862 gnd.n877 19.3944
R15643 gnd.n6868 gnd.n877 19.3944
R15644 gnd.n6868 gnd.n875 19.3944
R15645 gnd.n6872 gnd.n875 19.3944
R15646 gnd.n6872 gnd.n871 19.3944
R15647 gnd.n6878 gnd.n871 19.3944
R15648 gnd.n6878 gnd.n869 19.3944
R15649 gnd.n6882 gnd.n869 19.3944
R15650 gnd.n6882 gnd.n865 19.3944
R15651 gnd.n6888 gnd.n865 19.3944
R15652 gnd.n6888 gnd.n863 19.3944
R15653 gnd.n6892 gnd.n863 19.3944
R15654 gnd.n6892 gnd.n859 19.3944
R15655 gnd.n6898 gnd.n859 19.3944
R15656 gnd.n6898 gnd.n857 19.3944
R15657 gnd.n6902 gnd.n857 19.3944
R15658 gnd.n6902 gnd.n853 19.3944
R15659 gnd.n6908 gnd.n853 19.3944
R15660 gnd.n6908 gnd.n851 19.3944
R15661 gnd.n6912 gnd.n851 19.3944
R15662 gnd.n6912 gnd.n847 19.3944
R15663 gnd.n6918 gnd.n847 19.3944
R15664 gnd.n6918 gnd.n845 19.3944
R15665 gnd.n6922 gnd.n845 19.3944
R15666 gnd.n6922 gnd.n841 19.3944
R15667 gnd.n6928 gnd.n841 19.3944
R15668 gnd.n6928 gnd.n839 19.3944
R15669 gnd.n6932 gnd.n839 19.3944
R15670 gnd.n6932 gnd.n835 19.3944
R15671 gnd.n6938 gnd.n835 19.3944
R15672 gnd.n6938 gnd.n833 19.3944
R15673 gnd.n6942 gnd.n833 19.3944
R15674 gnd.n6942 gnd.n829 19.3944
R15675 gnd.n6948 gnd.n829 19.3944
R15676 gnd.n6948 gnd.n827 19.3944
R15677 gnd.n6952 gnd.n827 19.3944
R15678 gnd.n6952 gnd.n823 19.3944
R15679 gnd.n6958 gnd.n823 19.3944
R15680 gnd.n6958 gnd.n821 19.3944
R15681 gnd.n6962 gnd.n821 19.3944
R15682 gnd.n6962 gnd.n817 19.3944
R15683 gnd.n6968 gnd.n817 19.3944
R15684 gnd.n6968 gnd.n815 19.3944
R15685 gnd.n6972 gnd.n815 19.3944
R15686 gnd.n6972 gnd.n811 19.3944
R15687 gnd.n6978 gnd.n811 19.3944
R15688 gnd.n6978 gnd.n809 19.3944
R15689 gnd.n6982 gnd.n809 19.3944
R15690 gnd.n6982 gnd.n805 19.3944
R15691 gnd.n6988 gnd.n805 19.3944
R15692 gnd.n6988 gnd.n803 19.3944
R15693 gnd.n6992 gnd.n803 19.3944
R15694 gnd.n6992 gnd.n799 19.3944
R15695 gnd.n6998 gnd.n799 19.3944
R15696 gnd.n6998 gnd.n797 19.3944
R15697 gnd.n7002 gnd.n797 19.3944
R15698 gnd.n7002 gnd.n793 19.3944
R15699 gnd.n7008 gnd.n793 19.3944
R15700 gnd.n7008 gnd.n791 19.3944
R15701 gnd.n7012 gnd.n791 19.3944
R15702 gnd.n7012 gnd.n787 19.3944
R15703 gnd.n7018 gnd.n787 19.3944
R15704 gnd.n7018 gnd.n785 19.3944
R15705 gnd.n7022 gnd.n785 19.3944
R15706 gnd.n7022 gnd.n781 19.3944
R15707 gnd.n7028 gnd.n781 19.3944
R15708 gnd.n7028 gnd.n779 19.3944
R15709 gnd.n7032 gnd.n779 19.3944
R15710 gnd.n7032 gnd.n775 19.3944
R15711 gnd.n7038 gnd.n775 19.3944
R15712 gnd.n7038 gnd.n773 19.3944
R15713 gnd.n7042 gnd.n773 19.3944
R15714 gnd.n7042 gnd.n769 19.3944
R15715 gnd.n7048 gnd.n769 19.3944
R15716 gnd.n7048 gnd.n767 19.3944
R15717 gnd.n7052 gnd.n767 19.3944
R15718 gnd.n7052 gnd.n763 19.3944
R15719 gnd.n7058 gnd.n763 19.3944
R15720 gnd.n7058 gnd.n761 19.3944
R15721 gnd.n7062 gnd.n761 19.3944
R15722 gnd.n7062 gnd.n757 19.3944
R15723 gnd.n7068 gnd.n757 19.3944
R15724 gnd.n7068 gnd.n755 19.3944
R15725 gnd.n7072 gnd.n755 19.3944
R15726 gnd.n7072 gnd.n751 19.3944
R15727 gnd.n7078 gnd.n751 19.3944
R15728 gnd.n7078 gnd.n749 19.3944
R15729 gnd.n7082 gnd.n749 19.3944
R15730 gnd.n7082 gnd.n745 19.3944
R15731 gnd.n7088 gnd.n745 19.3944
R15732 gnd.n7088 gnd.n743 19.3944
R15733 gnd.n7092 gnd.n743 19.3944
R15734 gnd.n7092 gnd.n739 19.3944
R15735 gnd.n7098 gnd.n739 19.3944
R15736 gnd.n7098 gnd.n737 19.3944
R15737 gnd.n7102 gnd.n737 19.3944
R15738 gnd.n7102 gnd.n733 19.3944
R15739 gnd.n7108 gnd.n733 19.3944
R15740 gnd.n7108 gnd.n731 19.3944
R15741 gnd.n7112 gnd.n731 19.3944
R15742 gnd.n7112 gnd.n727 19.3944
R15743 gnd.n7118 gnd.n727 19.3944
R15744 gnd.n7118 gnd.n725 19.3944
R15745 gnd.n7123 gnd.n725 19.3944
R15746 gnd.n7123 gnd.n721 19.3944
R15747 gnd.n7129 gnd.n721 19.3944
R15748 gnd.n7130 gnd.n7129 19.3944
R15749 gnd.n4498 gnd.n4497 19.3944
R15750 gnd.n4497 gnd.n4496 19.3944
R15751 gnd.n4496 gnd.n4495 19.3944
R15752 gnd.n4495 gnd.n4493 19.3944
R15753 gnd.n4493 gnd.n4490 19.3944
R15754 gnd.n4490 gnd.n4489 19.3944
R15755 gnd.n4489 gnd.n4486 19.3944
R15756 gnd.n4486 gnd.n4485 19.3944
R15757 gnd.n4485 gnd.n4482 19.3944
R15758 gnd.n4482 gnd.n4481 19.3944
R15759 gnd.n4481 gnd.n4478 19.3944
R15760 gnd.n4478 gnd.n4477 19.3944
R15761 gnd.n4477 gnd.n4474 19.3944
R15762 gnd.n4474 gnd.n4473 19.3944
R15763 gnd.n4473 gnd.n4470 19.3944
R15764 gnd.n4470 gnd.n4469 19.3944
R15765 gnd.n4469 gnd.n4466 19.3944
R15766 gnd.n4464 gnd.n4461 19.3944
R15767 gnd.n4461 gnd.n4460 19.3944
R15768 gnd.n4460 gnd.n4457 19.3944
R15769 gnd.n4457 gnd.n4456 19.3944
R15770 gnd.n4456 gnd.n4453 19.3944
R15771 gnd.n4453 gnd.n4452 19.3944
R15772 gnd.n4452 gnd.n4449 19.3944
R15773 gnd.n4447 gnd.n4444 19.3944
R15774 gnd.n4444 gnd.n4443 19.3944
R15775 gnd.n4443 gnd.n4440 19.3944
R15776 gnd.n4440 gnd.n4439 19.3944
R15777 gnd.n4439 gnd.n4436 19.3944
R15778 gnd.n4436 gnd.n4435 19.3944
R15779 gnd.n4435 gnd.n4432 19.3944
R15780 gnd.n4432 gnd.n4431 19.3944
R15781 gnd.n4427 gnd.n4424 19.3944
R15782 gnd.n4424 gnd.n4423 19.3944
R15783 gnd.n4423 gnd.n4420 19.3944
R15784 gnd.n4420 gnd.n4419 19.3944
R15785 gnd.n4419 gnd.n4416 19.3944
R15786 gnd.n4416 gnd.n4415 19.3944
R15787 gnd.n4415 gnd.n4412 19.3944
R15788 gnd.n4412 gnd.n4411 19.3944
R15789 gnd.n4411 gnd.n4408 19.3944
R15790 gnd.n4408 gnd.n4407 19.3944
R15791 gnd.n4407 gnd.n4404 19.3944
R15792 gnd.n4404 gnd.n4403 19.3944
R15793 gnd.n4403 gnd.n4400 19.3944
R15794 gnd.n4400 gnd.n4399 19.3944
R15795 gnd.n4399 gnd.n4396 19.3944
R15796 gnd.n4396 gnd.n4395 19.3944
R15797 gnd.n4395 gnd.n4392 19.3944
R15798 gnd.n4392 gnd.n4391 19.3944
R15799 gnd.n4375 gnd.n1970 19.3944
R15800 gnd.n4375 gnd.n4374 19.3944
R15801 gnd.n4374 gnd.n1979 19.3944
R15802 gnd.n2070 gnd.n1979 19.3944
R15803 gnd.n4272 gnd.n2070 19.3944
R15804 gnd.n4273 gnd.n4272 19.3944
R15805 gnd.n4275 gnd.n4273 19.3944
R15806 gnd.n4275 gnd.n2066 19.3944
R15807 gnd.n4287 gnd.n2066 19.3944
R15808 gnd.n4288 gnd.n4287 19.3944
R15809 gnd.n4298 gnd.n4288 19.3944
R15810 gnd.n4298 gnd.n4297 19.3944
R15811 gnd.n4297 gnd.n4296 19.3944
R15812 gnd.n4296 gnd.n4295 19.3944
R15813 gnd.n4295 gnd.n4294 19.3944
R15814 gnd.n4294 gnd.n4293 19.3944
R15815 gnd.n4293 gnd.n573 19.3944
R15816 gnd.n7372 gnd.n573 19.3944
R15817 gnd.n7373 gnd.n7372 19.3944
R15818 gnd.n7373 gnd.n545 19.3944
R15819 gnd.n7404 gnd.n545 19.3944
R15820 gnd.n7405 gnd.n7404 19.3944
R15821 gnd.n7408 gnd.n7405 19.3944
R15822 gnd.n7409 gnd.n7408 19.3944
R15823 gnd.n7409 gnd.n517 19.3944
R15824 gnd.n7440 gnd.n517 19.3944
R15825 gnd.n7441 gnd.n7440 19.3944
R15826 gnd.n7442 gnd.n7441 19.3944
R15827 gnd.n7444 gnd.n7442 19.3944
R15828 gnd.n7444 gnd.n7443 19.3944
R15829 gnd.n7443 gnd.n487 19.3944
R15830 gnd.n7478 gnd.n487 19.3944
R15831 gnd.n7480 gnd.n7478 19.3944
R15832 gnd.n7480 gnd.n7479 19.3944
R15833 gnd.n7479 gnd.n480 19.3944
R15834 gnd.n7492 gnd.n480 19.3944
R15835 gnd.n7493 gnd.n7492 19.3944
R15836 gnd.n7495 gnd.n7493 19.3944
R15837 gnd.n7496 gnd.n7495 19.3944
R15838 gnd.n7499 gnd.n7496 19.3944
R15839 gnd.n7500 gnd.n7499 19.3944
R15840 gnd.n7502 gnd.n7500 19.3944
R15841 gnd.n7503 gnd.n7502 19.3944
R15842 gnd.n7506 gnd.n7503 19.3944
R15843 gnd.n7507 gnd.n7506 19.3944
R15844 gnd.n7509 gnd.n7507 19.3944
R15845 gnd.n7510 gnd.n7509 19.3944
R15846 gnd.n7513 gnd.n7510 19.3944
R15847 gnd.n7514 gnd.n7513 19.3944
R15848 gnd.n7516 gnd.n7514 19.3944
R15849 gnd.n7517 gnd.n7516 19.3944
R15850 gnd.n7520 gnd.n7517 19.3944
R15851 gnd.n7521 gnd.n7520 19.3944
R15852 gnd.n7523 gnd.n7521 19.3944
R15853 gnd.n7524 gnd.n7523 19.3944
R15854 gnd.n7527 gnd.n7524 19.3944
R15855 gnd.n7528 gnd.n7527 19.3944
R15856 gnd.n7530 gnd.n7528 19.3944
R15857 gnd.n7531 gnd.n7530 19.3944
R15858 gnd.n7534 gnd.n7531 19.3944
R15859 gnd.n7535 gnd.n7534 19.3944
R15860 gnd.n7537 gnd.n7535 19.3944
R15861 gnd.n7538 gnd.n7537 19.3944
R15862 gnd.n7541 gnd.n7538 19.3944
R15863 gnd.n4378 gnd.n4377 19.3944
R15864 gnd.n4377 gnd.n1977 19.3944
R15865 gnd.n2001 gnd.n1977 19.3944
R15866 gnd.n4364 gnd.n2001 19.3944
R15867 gnd.n4364 gnd.n4363 19.3944
R15868 gnd.n4363 gnd.n4362 19.3944
R15869 gnd.n4362 gnd.n2006 19.3944
R15870 gnd.n4352 gnd.n2006 19.3944
R15871 gnd.n4352 gnd.n4351 19.3944
R15872 gnd.n4351 gnd.n4350 19.3944
R15873 gnd.n4350 gnd.n2027 19.3944
R15874 gnd.n4340 gnd.n2027 19.3944
R15875 gnd.n4340 gnd.n4339 19.3944
R15876 gnd.n4339 gnd.n4338 19.3944
R15877 gnd.n4338 gnd.n2047 19.3944
R15878 gnd.n2047 gnd.n570 19.3944
R15879 gnd.n7381 gnd.n570 19.3944
R15880 gnd.n7381 gnd.n7380 19.3944
R15881 gnd.n7380 gnd.n7379 19.3944
R15882 gnd.n7379 gnd.n7378 19.3944
R15883 gnd.n7378 gnd.n542 19.3944
R15884 gnd.n7417 gnd.n542 19.3944
R15885 gnd.n7417 gnd.n7416 19.3944
R15886 gnd.n7416 gnd.n7415 19.3944
R15887 gnd.n7415 gnd.n7414 19.3944
R15888 gnd.n7414 gnd.n512 19.3944
R15889 gnd.n7450 gnd.n512 19.3944
R15890 gnd.n7450 gnd.n7449 19.3944
R15891 gnd.n7449 gnd.n7448 19.3944
R15892 gnd.n7448 gnd.n489 19.3944
R15893 gnd.n7475 gnd.n489 19.3944
R15894 gnd.n7475 gnd.n482 19.3944
R15895 gnd.n7484 gnd.n482 19.3944
R15896 gnd.n7485 gnd.n7484 19.3944
R15897 gnd.n7487 gnd.n7485 19.3944
R15898 gnd.n7487 gnd.n123 19.3944
R15899 gnd.n7747 gnd.n123 19.3944
R15900 gnd.n7747 gnd.n7746 19.3944
R15901 gnd.n7746 gnd.n7745 19.3944
R15902 gnd.n7745 gnd.n127 19.3944
R15903 gnd.n7735 gnd.n127 19.3944
R15904 gnd.n7735 gnd.n7734 19.3944
R15905 gnd.n7734 gnd.n7733 19.3944
R15906 gnd.n7733 gnd.n144 19.3944
R15907 gnd.n7723 gnd.n144 19.3944
R15908 gnd.n7723 gnd.n7722 19.3944
R15909 gnd.n7722 gnd.n7721 19.3944
R15910 gnd.n7721 gnd.n164 19.3944
R15911 gnd.n7711 gnd.n164 19.3944
R15912 gnd.n7711 gnd.n7710 19.3944
R15913 gnd.n7710 gnd.n7709 19.3944
R15914 gnd.n7709 gnd.n182 19.3944
R15915 gnd.n7699 gnd.n182 19.3944
R15916 gnd.n7699 gnd.n7698 19.3944
R15917 gnd.n7698 gnd.n7697 19.3944
R15918 gnd.n7697 gnd.n202 19.3944
R15919 gnd.n7687 gnd.n202 19.3944
R15920 gnd.n7687 gnd.n7686 19.3944
R15921 gnd.n7686 gnd.n7685 19.3944
R15922 gnd.n7685 gnd.n220 19.3944
R15923 gnd.n7675 gnd.n220 19.3944
R15924 gnd.n7675 gnd.n7674 19.3944
R15925 gnd.n7674 gnd.n7673 19.3944
R15926 gnd.n7673 gnd.n240 19.3944
R15927 gnd.n7584 gnd.n325 19.3944
R15928 gnd.n7584 gnd.n7581 19.3944
R15929 gnd.n7581 gnd.n7578 19.3944
R15930 gnd.n7578 gnd.n7577 19.3944
R15931 gnd.n7577 gnd.n7574 19.3944
R15932 gnd.n7574 gnd.n7573 19.3944
R15933 gnd.n7573 gnd.n7570 19.3944
R15934 gnd.n7570 gnd.n7569 19.3944
R15935 gnd.n7569 gnd.n7566 19.3944
R15936 gnd.n7566 gnd.n7565 19.3944
R15937 gnd.n7565 gnd.n7562 19.3944
R15938 gnd.n7562 gnd.n7561 19.3944
R15939 gnd.n7561 gnd.n7558 19.3944
R15940 gnd.n7558 gnd.n7557 19.3944
R15941 gnd.n7557 gnd.n7554 19.3944
R15942 gnd.n7554 gnd.n7553 19.3944
R15943 gnd.n7553 gnd.n7550 19.3944
R15944 gnd.n7550 gnd.n7549 19.3944
R15945 gnd.n7627 gnd.n7624 19.3944
R15946 gnd.n7624 gnd.n7623 19.3944
R15947 gnd.n7623 gnd.n7620 19.3944
R15948 gnd.n7620 gnd.n7619 19.3944
R15949 gnd.n7619 gnd.n7616 19.3944
R15950 gnd.n7616 gnd.n7615 19.3944
R15951 gnd.n7615 gnd.n7612 19.3944
R15952 gnd.n7612 gnd.n7611 19.3944
R15953 gnd.n7611 gnd.n7608 19.3944
R15954 gnd.n7608 gnd.n7607 19.3944
R15955 gnd.n7607 gnd.n7604 19.3944
R15956 gnd.n7604 gnd.n7603 19.3944
R15957 gnd.n7603 gnd.n7600 19.3944
R15958 gnd.n7600 gnd.n7599 19.3944
R15959 gnd.n7599 gnd.n7596 19.3944
R15960 gnd.n7596 gnd.n7595 19.3944
R15961 gnd.n7595 gnd.n7592 19.3944
R15962 gnd.n7592 gnd.n7591 19.3944
R15963 gnd.n7665 gnd.n249 19.3944
R15964 gnd.n7660 gnd.n249 19.3944
R15965 gnd.n7660 gnd.n7659 19.3944
R15966 gnd.n7659 gnd.n7658 19.3944
R15967 gnd.n7658 gnd.n7655 19.3944
R15968 gnd.n7655 gnd.n7654 19.3944
R15969 gnd.n7654 gnd.n7651 19.3944
R15970 gnd.n7651 gnd.n7650 19.3944
R15971 gnd.n7650 gnd.n7647 19.3944
R15972 gnd.n7647 gnd.n7646 19.3944
R15973 gnd.n7646 gnd.n7643 19.3944
R15974 gnd.n7643 gnd.n7642 19.3944
R15975 gnd.n7642 gnd.n7639 19.3944
R15976 gnd.n7639 gnd.n7638 19.3944
R15977 gnd.n7638 gnd.n7635 19.3944
R15978 gnd.n7635 gnd.n7634 19.3944
R15979 gnd.n7634 gnd.n7631 19.3944
R15980 gnd.n478 gnd.n477 19.3944
R15981 gnd.n477 gnd.n476 19.3944
R15982 gnd.n476 gnd.n473 19.3944
R15983 gnd.n473 gnd.n472 19.3944
R15984 gnd.n472 gnd.n469 19.3944
R15985 gnd.n469 gnd.n468 19.3944
R15986 gnd.n468 gnd.n465 19.3944
R15987 gnd.n465 gnd.n464 19.3944
R15988 gnd.n464 gnd.n461 19.3944
R15989 gnd.n461 gnd.n460 19.3944
R15990 gnd.n460 gnd.n457 19.3944
R15991 gnd.n457 gnd.n456 19.3944
R15992 gnd.n456 gnd.n453 19.3944
R15993 gnd.n453 gnd.n452 19.3944
R15994 gnd.n452 gnd.n449 19.3944
R15995 gnd.n449 gnd.n448 19.3944
R15996 gnd.n4260 gnd.n2073 19.3944
R15997 gnd.n4261 gnd.n4260 19.3944
R15998 gnd.n4264 gnd.n4261 19.3944
R15999 gnd.n4264 gnd.n2071 19.3944
R16000 gnd.n4268 gnd.n2071 19.3944
R16001 gnd.n4268 gnd.n2069 19.3944
R16002 gnd.n4279 gnd.n2069 19.3944
R16003 gnd.n4279 gnd.n2067 19.3944
R16004 gnd.n4283 gnd.n2067 19.3944
R16005 gnd.n4283 gnd.n2065 19.3944
R16006 gnd.n4302 gnd.n2065 19.3944
R16007 gnd.n4302 gnd.n2062 19.3944
R16008 gnd.n4314 gnd.n2062 19.3944
R16009 gnd.n4314 gnd.n2063 19.3944
R16010 gnd.n4310 gnd.n2063 19.3944
R16011 gnd.n4310 gnd.n4309 19.3944
R16012 gnd.n4309 gnd.n4308 19.3944
R16013 gnd.n4308 gnd.n553 19.3944
R16014 gnd.n7395 gnd.n553 19.3944
R16015 gnd.n7395 gnd.n550 19.3944
R16016 gnd.n7400 gnd.n550 19.3944
R16017 gnd.n7400 gnd.n551 19.3944
R16018 gnd.n551 gnd.n524 19.3944
R16019 gnd.n7432 gnd.n524 19.3944
R16020 gnd.n7432 gnd.n522 19.3944
R16021 gnd.n7436 gnd.n522 19.3944
R16022 gnd.n7436 gnd.n502 19.3944
R16023 gnd.n7459 gnd.n502 19.3944
R16024 gnd.n7459 gnd.n499 19.3944
R16025 gnd.n7463 gnd.n499 19.3944
R16026 gnd.n7463 gnd.n500 19.3944
R16027 gnd.n500 gnd.n96 19.3944
R16028 gnd.n7760 gnd.n96 19.3944
R16029 gnd.n7760 gnd.n7759 19.3944
R16030 gnd.n7759 gnd.n99 19.3944
R16031 gnd.n384 gnd.n99 19.3944
R16032 gnd.n384 gnd.n381 19.3944
R16033 gnd.n389 gnd.n381 19.3944
R16034 gnd.n390 gnd.n389 19.3944
R16035 gnd.n392 gnd.n390 19.3944
R16036 gnd.n392 gnd.n379 19.3944
R16037 gnd.n397 gnd.n379 19.3944
R16038 gnd.n398 gnd.n397 19.3944
R16039 gnd.n400 gnd.n398 19.3944
R16040 gnd.n400 gnd.n377 19.3944
R16041 gnd.n405 gnd.n377 19.3944
R16042 gnd.n406 gnd.n405 19.3944
R16043 gnd.n408 gnd.n406 19.3944
R16044 gnd.n408 gnd.n375 19.3944
R16045 gnd.n413 gnd.n375 19.3944
R16046 gnd.n414 gnd.n413 19.3944
R16047 gnd.n416 gnd.n414 19.3944
R16048 gnd.n416 gnd.n373 19.3944
R16049 gnd.n421 gnd.n373 19.3944
R16050 gnd.n422 gnd.n421 19.3944
R16051 gnd.n424 gnd.n422 19.3944
R16052 gnd.n424 gnd.n371 19.3944
R16053 gnd.n429 gnd.n371 19.3944
R16054 gnd.n430 gnd.n429 19.3944
R16055 gnd.n432 gnd.n430 19.3944
R16056 gnd.n432 gnd.n369 19.3944
R16057 gnd.n437 gnd.n369 19.3944
R16058 gnd.n438 gnd.n437 19.3944
R16059 gnd.n441 gnd.n438 19.3944
R16060 gnd.n1987 gnd.n1986 19.3944
R16061 gnd.n4370 gnd.n1986 19.3944
R16062 gnd.n4370 gnd.n4369 19.3944
R16063 gnd.n4369 gnd.n4368 19.3944
R16064 gnd.n4368 gnd.n1993 19.3944
R16065 gnd.n4358 gnd.n1993 19.3944
R16066 gnd.n4358 gnd.n4357 19.3944
R16067 gnd.n4357 gnd.n4356 19.3944
R16068 gnd.n4356 gnd.n2017 19.3944
R16069 gnd.n4346 gnd.n2017 19.3944
R16070 gnd.n4346 gnd.n4345 19.3944
R16071 gnd.n4345 gnd.n4344 19.3944
R16072 gnd.n4344 gnd.n2038 19.3944
R16073 gnd.n4334 gnd.n2038 19.3944
R16074 gnd.n4334 gnd.n4333 19.3944
R16075 gnd.n4333 gnd.n563 19.3944
R16076 gnd.n7385 gnd.n563 19.3944
R16077 gnd.n7385 gnd.n561 19.3944
R16078 gnd.n7391 gnd.n561 19.3944
R16079 gnd.n7391 gnd.n7390 19.3944
R16080 gnd.n7390 gnd.n534 19.3944
R16081 gnd.n7421 gnd.n534 19.3944
R16082 gnd.n7421 gnd.n532 19.3944
R16083 gnd.n7428 gnd.n532 19.3944
R16084 gnd.n7428 gnd.n7427 19.3944
R16085 gnd.n7427 gnd.n7426 19.3944
R16086 gnd.n7426 gnd.n508 19.3944
R16087 gnd.n7455 gnd.n7454 19.3944
R16088 gnd.n7471 gnd.n7470 19.3944
R16089 gnd.n7468 gnd.n7467 19.3944
R16090 gnd.n7755 gnd.n7754 19.3944
R16091 gnd.n7751 gnd.n107 19.3944
R16092 gnd.n7751 gnd.n114 19.3944
R16093 gnd.n7741 gnd.n114 19.3944
R16094 gnd.n7741 gnd.n7740 19.3944
R16095 gnd.n7740 gnd.n7739 19.3944
R16096 gnd.n7739 gnd.n136 19.3944
R16097 gnd.n7729 gnd.n136 19.3944
R16098 gnd.n7729 gnd.n7728 19.3944
R16099 gnd.n7728 gnd.n7727 19.3944
R16100 gnd.n7727 gnd.n154 19.3944
R16101 gnd.n7717 gnd.n154 19.3944
R16102 gnd.n7717 gnd.n7716 19.3944
R16103 gnd.n7716 gnd.n7715 19.3944
R16104 gnd.n7715 gnd.n174 19.3944
R16105 gnd.n7705 gnd.n174 19.3944
R16106 gnd.n7705 gnd.n7704 19.3944
R16107 gnd.n7704 gnd.n7703 19.3944
R16108 gnd.n7703 gnd.n192 19.3944
R16109 gnd.n7693 gnd.n192 19.3944
R16110 gnd.n7693 gnd.n7692 19.3944
R16111 gnd.n7692 gnd.n7691 19.3944
R16112 gnd.n7691 gnd.n212 19.3944
R16113 gnd.n7681 gnd.n212 19.3944
R16114 gnd.n7681 gnd.n7680 19.3944
R16115 gnd.n7680 gnd.n7679 19.3944
R16116 gnd.n7679 gnd.n231 19.3944
R16117 gnd.n7669 gnd.n231 19.3944
R16118 gnd.n7669 gnd.n7668 19.3944
R16119 gnd.n5108 gnd.n5107 19.3944
R16120 gnd.n5107 gnd.n5106 19.3944
R16121 gnd.n5106 gnd.n5105 19.3944
R16122 gnd.n5105 gnd.n5103 19.3944
R16123 gnd.n5103 gnd.n5100 19.3944
R16124 gnd.n5100 gnd.n5099 19.3944
R16125 gnd.n5099 gnd.n5096 19.3944
R16126 gnd.n5096 gnd.n5095 19.3944
R16127 gnd.n5095 gnd.n5092 19.3944
R16128 gnd.n5092 gnd.n5091 19.3944
R16129 gnd.n5091 gnd.n5088 19.3944
R16130 gnd.n5088 gnd.n5087 19.3944
R16131 gnd.n5087 gnd.n5084 19.3944
R16132 gnd.n5084 gnd.n5083 19.3944
R16133 gnd.n5083 gnd.n5080 19.3944
R16134 gnd.n5080 gnd.n5079 19.3944
R16135 gnd.n5079 gnd.n5076 19.3944
R16136 gnd.n5074 gnd.n5071 19.3944
R16137 gnd.n5071 gnd.n5070 19.3944
R16138 gnd.n5070 gnd.n5067 19.3944
R16139 gnd.n5067 gnd.n5066 19.3944
R16140 gnd.n5066 gnd.n5063 19.3944
R16141 gnd.n5063 gnd.n5062 19.3944
R16142 gnd.n5062 gnd.n5059 19.3944
R16143 gnd.n5059 gnd.n5058 19.3944
R16144 gnd.n5058 gnd.n5055 19.3944
R16145 gnd.n5055 gnd.n5054 19.3944
R16146 gnd.n5054 gnd.n5051 19.3944
R16147 gnd.n5051 gnd.n5050 19.3944
R16148 gnd.n5050 gnd.n5047 19.3944
R16149 gnd.n5047 gnd.n5046 19.3944
R16150 gnd.n5046 gnd.n5043 19.3944
R16151 gnd.n5043 gnd.n5042 19.3944
R16152 gnd.n5042 gnd.n5039 19.3944
R16153 gnd.n5039 gnd.n5038 19.3944
R16154 gnd.n5034 gnd.n5031 19.3944
R16155 gnd.n5031 gnd.n5030 19.3944
R16156 gnd.n5030 gnd.n5027 19.3944
R16157 gnd.n5027 gnd.n5026 19.3944
R16158 gnd.n5026 gnd.n5023 19.3944
R16159 gnd.n5023 gnd.n5022 19.3944
R16160 gnd.n5022 gnd.n5019 19.3944
R16161 gnd.n5019 gnd.n5018 19.3944
R16162 gnd.n5018 gnd.n5015 19.3944
R16163 gnd.n5015 gnd.n5014 19.3944
R16164 gnd.n5014 gnd.n5011 19.3944
R16165 gnd.n5011 gnd.n5010 19.3944
R16166 gnd.n5010 gnd.n5007 19.3944
R16167 gnd.n5007 gnd.n5006 19.3944
R16168 gnd.n5006 gnd.n5003 19.3944
R16169 gnd.n5003 gnd.n5002 19.3944
R16170 gnd.n5002 gnd.n4999 19.3944
R16171 gnd.n4999 gnd.n4998 19.3944
R16172 gnd.n2761 gnd.n2760 19.3944
R16173 gnd.n2764 gnd.n2761 19.3944
R16174 gnd.n2764 gnd.n2756 19.3944
R16175 gnd.n2770 gnd.n2756 19.3944
R16176 gnd.n2771 gnd.n2770 19.3944
R16177 gnd.n2774 gnd.n2771 19.3944
R16178 gnd.n2774 gnd.n2754 19.3944
R16179 gnd.n2780 gnd.n2754 19.3944
R16180 gnd.n2781 gnd.n2780 19.3944
R16181 gnd.n2784 gnd.n2781 19.3944
R16182 gnd.n2784 gnd.n2752 19.3944
R16183 gnd.n2790 gnd.n2752 19.3944
R16184 gnd.n2791 gnd.n2790 19.3944
R16185 gnd.n2794 gnd.n2791 19.3944
R16186 gnd.n2794 gnd.n2748 19.3944
R16187 gnd.n2798 gnd.n2748 19.3944
R16188 gnd.n2805 gnd.n2804 19.3944
R16189 gnd.n2807 gnd.n2805 19.3944
R16190 gnd.n2807 gnd.n2742 19.3944
R16191 gnd.n2812 gnd.n2742 19.3944
R16192 gnd.n2813 gnd.n2812 19.3944
R16193 gnd.n2815 gnd.n2813 19.3944
R16194 gnd.n2815 gnd.n2740 19.3944
R16195 gnd.n2820 gnd.n2740 19.3944
R16196 gnd.n2821 gnd.n2820 19.3944
R16197 gnd.n2823 gnd.n2821 19.3944
R16198 gnd.n2823 gnd.n2738 19.3944
R16199 gnd.n2828 gnd.n2738 19.3944
R16200 gnd.n2829 gnd.n2828 19.3944
R16201 gnd.n2831 gnd.n2829 19.3944
R16202 gnd.n2831 gnd.n2736 19.3944
R16203 gnd.n2836 gnd.n2736 19.3944
R16204 gnd.n2837 gnd.n2836 19.3944
R16205 gnd.n2839 gnd.n2837 19.3944
R16206 gnd.n2839 gnd.n2734 19.3944
R16207 gnd.n2844 gnd.n2734 19.3944
R16208 gnd.n2845 gnd.n2844 19.3944
R16209 gnd.n2847 gnd.n2845 19.3944
R16210 gnd.n2847 gnd.n2732 19.3944
R16211 gnd.n2852 gnd.n2732 19.3944
R16212 gnd.n2853 gnd.n2852 19.3944
R16213 gnd.n2855 gnd.n2853 19.3944
R16214 gnd.n2855 gnd.n2730 19.3944
R16215 gnd.n2860 gnd.n2730 19.3944
R16216 gnd.n2861 gnd.n2860 19.3944
R16217 gnd.n2863 gnd.n2861 19.3944
R16218 gnd.n2863 gnd.n2728 19.3944
R16219 gnd.n2867 gnd.n2728 19.3944
R16220 gnd.n2867 gnd.n2646 19.3944
R16221 gnd.n2893 gnd.n2646 19.3944
R16222 gnd.n2893 gnd.n2644 19.3944
R16223 gnd.n2897 gnd.n2644 19.3944
R16224 gnd.n2897 gnd.n2633 19.3944
R16225 gnd.n2932 gnd.n2633 19.3944
R16226 gnd.n2932 gnd.n2631 19.3944
R16227 gnd.n2936 gnd.n2631 19.3944
R16228 gnd.n2936 gnd.n2627 19.3944
R16229 gnd.n2946 gnd.n2627 19.3944
R16230 gnd.n2946 gnd.n2625 19.3944
R16231 gnd.n2950 gnd.n2625 19.3944
R16232 gnd.n2950 gnd.n2616 19.3944
R16233 gnd.n2985 gnd.n2616 19.3944
R16234 gnd.n2985 gnd.n2617 19.3944
R16235 gnd.n2981 gnd.n2617 19.3944
R16236 gnd.n2981 gnd.n2980 19.3944
R16237 gnd.n2980 gnd.n2979 19.3944
R16238 gnd.n2979 gnd.n2622 19.3944
R16239 gnd.n2975 gnd.n2622 19.3944
R16240 gnd.n2975 gnd.n2602 19.3944
R16241 gnd.n3013 gnd.n2602 19.3944
R16242 gnd.n3013 gnd.n2600 19.3944
R16243 gnd.n3017 gnd.n2600 19.3944
R16244 gnd.n3017 gnd.n2593 19.3944
R16245 gnd.n3289 gnd.n2593 19.3944
R16246 gnd.n3289 gnd.n2594 19.3944
R16247 gnd.n3285 gnd.n2594 19.3944
R16248 gnd.n3285 gnd.n3284 19.3944
R16249 gnd.n3284 gnd.n3283 19.3944
R16250 gnd.n3283 gnd.n3280 19.3944
R16251 gnd.n3280 gnd.n2580 19.3944
R16252 gnd.n4990 gnd.n1257 19.3944
R16253 gnd.n2671 gnd.n1257 19.3944
R16254 gnd.n2672 gnd.n2671 19.3944
R16255 gnd.n2674 gnd.n2672 19.3944
R16256 gnd.n2675 gnd.n2674 19.3944
R16257 gnd.n2678 gnd.n2675 19.3944
R16258 gnd.n2679 gnd.n2678 19.3944
R16259 gnd.n2681 gnd.n2679 19.3944
R16260 gnd.n2682 gnd.n2681 19.3944
R16261 gnd.n2685 gnd.n2682 19.3944
R16262 gnd.n2686 gnd.n2685 19.3944
R16263 gnd.n2688 gnd.n2686 19.3944
R16264 gnd.n2689 gnd.n2688 19.3944
R16265 gnd.n2692 gnd.n2689 19.3944
R16266 gnd.n2693 gnd.n2692 19.3944
R16267 gnd.n2695 gnd.n2693 19.3944
R16268 gnd.n2696 gnd.n2695 19.3944
R16269 gnd.n2699 gnd.n2696 19.3944
R16270 gnd.n2700 gnd.n2699 19.3944
R16271 gnd.n2702 gnd.n2700 19.3944
R16272 gnd.n2703 gnd.n2702 19.3944
R16273 gnd.n2706 gnd.n2703 19.3944
R16274 gnd.n2707 gnd.n2706 19.3944
R16275 gnd.n2709 gnd.n2707 19.3944
R16276 gnd.n2710 gnd.n2709 19.3944
R16277 gnd.n2713 gnd.n2710 19.3944
R16278 gnd.n2714 gnd.n2713 19.3944
R16279 gnd.n2716 gnd.n2714 19.3944
R16280 gnd.n2717 gnd.n2716 19.3944
R16281 gnd.n2719 gnd.n2717 19.3944
R16282 gnd.n2719 gnd.n2667 19.3944
R16283 gnd.n2871 gnd.n2667 19.3944
R16284 gnd.n2872 gnd.n2871 19.3944
R16285 gnd.n2873 gnd.n2872 19.3944
R16286 gnd.n2878 gnd.n2873 19.3944
R16287 gnd.n2878 gnd.n2876 19.3944
R16288 gnd.n2876 gnd.n2875 19.3944
R16289 gnd.n2875 gnd.n2874 19.3944
R16290 gnd.n2874 gnd.n2629 19.3944
R16291 gnd.n2940 gnd.n2629 19.3944
R16292 gnd.n2941 gnd.n2940 19.3944
R16293 gnd.n2942 gnd.n2941 19.3944
R16294 gnd.n2942 gnd.n2623 19.3944
R16295 gnd.n2954 gnd.n2623 19.3944
R16296 gnd.n2955 gnd.n2954 19.3944
R16297 gnd.n2956 gnd.n2955 19.3944
R16298 gnd.n2957 gnd.n2956 19.3944
R16299 gnd.n2961 gnd.n2957 19.3944
R16300 gnd.n2962 gnd.n2961 19.3944
R16301 gnd.n2966 gnd.n2962 19.3944
R16302 gnd.n2967 gnd.n2966 19.3944
R16303 gnd.n2971 gnd.n2967 19.3944
R16304 gnd.n2971 gnd.n2970 19.3944
R16305 gnd.n2970 gnd.n2969 19.3944
R16306 gnd.n2969 gnd.n2598 19.3944
R16307 gnd.n3021 gnd.n2598 19.3944
R16308 gnd.n3022 gnd.n3021 19.3944
R16309 gnd.n3023 gnd.n3022 19.3944
R16310 gnd.n3024 gnd.n3023 19.3944
R16311 gnd.n3028 gnd.n3024 19.3944
R16312 gnd.n3029 gnd.n3028 19.3944
R16313 gnd.n3276 gnd.n3029 19.3944
R16314 gnd.n3276 gnd.n3275 19.3944
R16315 gnd.n3275 gnd.n3274 19.3944
R16316 gnd.n1276 gnd.n1255 19.3944
R16317 gnd.n1277 gnd.n1276 19.3944
R16318 gnd.n4979 gnd.n1277 19.3944
R16319 gnd.n4979 gnd.n4978 19.3944
R16320 gnd.n4978 gnd.n4977 19.3944
R16321 gnd.n4977 gnd.n1281 19.3944
R16322 gnd.n4967 gnd.n1281 19.3944
R16323 gnd.n4967 gnd.n4966 19.3944
R16324 gnd.n4966 gnd.n4965 19.3944
R16325 gnd.n4965 gnd.n1300 19.3944
R16326 gnd.n4955 gnd.n1300 19.3944
R16327 gnd.n4955 gnd.n4954 19.3944
R16328 gnd.n4954 gnd.n4953 19.3944
R16329 gnd.n4953 gnd.n1319 19.3944
R16330 gnd.n4943 gnd.n1319 19.3944
R16331 gnd.n4943 gnd.n4942 19.3944
R16332 gnd.n4942 gnd.n4941 19.3944
R16333 gnd.n4941 gnd.n1338 19.3944
R16334 gnd.n4931 gnd.n1338 19.3944
R16335 gnd.n4931 gnd.n4930 19.3944
R16336 gnd.n4930 gnd.n4929 19.3944
R16337 gnd.n4929 gnd.n1357 19.3944
R16338 gnd.n4919 gnd.n1357 19.3944
R16339 gnd.n4919 gnd.n4918 19.3944
R16340 gnd.n4918 gnd.n4917 19.3944
R16341 gnd.n4917 gnd.n1376 19.3944
R16342 gnd.n4907 gnd.n1376 19.3944
R16343 gnd.n4907 gnd.n4906 19.3944
R16344 gnd.n4906 gnd.n4905 19.3944
R16345 gnd.n4905 gnd.n1394 19.3944
R16346 gnd.n2722 gnd.n1394 19.3944
R16347 gnd.n2722 gnd.n2663 19.3944
R16348 gnd.n2883 gnd.n2663 19.3944
R16349 gnd.n2883 gnd.n2882 19.3944
R16350 gnd.n2882 gnd.n2881 19.3944
R16351 gnd.n2881 gnd.n1417 19.3944
R16352 gnd.n4894 gnd.n1417 19.3944
R16353 gnd.n4894 gnd.n4893 19.3944
R16354 gnd.n4893 gnd.n4892 19.3944
R16355 gnd.n4892 gnd.n1421 19.3944
R16356 gnd.n4882 gnd.n1421 19.3944
R16357 gnd.n4882 gnd.n4881 19.3944
R16358 gnd.n4881 gnd.n4880 19.3944
R16359 gnd.n4880 gnd.n1439 19.3944
R16360 gnd.n4870 gnd.n1439 19.3944
R16361 gnd.n4870 gnd.n4869 19.3944
R16362 gnd.n4869 gnd.n4868 19.3944
R16363 gnd.n4868 gnd.n1460 19.3944
R16364 gnd.n4858 gnd.n1460 19.3944
R16365 gnd.n4858 gnd.n4857 19.3944
R16366 gnd.n4857 gnd.n4856 19.3944
R16367 gnd.n4856 gnd.n1479 19.3944
R16368 gnd.n4846 gnd.n1479 19.3944
R16369 gnd.n4846 gnd.n4845 19.3944
R16370 gnd.n4845 gnd.n4844 19.3944
R16371 gnd.n4844 gnd.n1500 19.3944
R16372 gnd.n4834 gnd.n1500 19.3944
R16373 gnd.n4834 gnd.n4833 19.3944
R16374 gnd.n4833 gnd.n4832 19.3944
R16375 gnd.n4832 gnd.n1519 19.3944
R16376 gnd.n4822 gnd.n1519 19.3944
R16377 gnd.n4822 gnd.n4821 19.3944
R16378 gnd.n4821 gnd.n4820 19.3944
R16379 gnd.n4820 gnd.n1540 19.3944
R16380 gnd.n4812 gnd.n1550 19.3944
R16381 gnd.n4807 gnd.n1550 19.3944
R16382 gnd.n4807 gnd.n4806 19.3944
R16383 gnd.n4806 gnd.n4805 19.3944
R16384 gnd.n4805 gnd.n4802 19.3944
R16385 gnd.n4802 gnd.n4801 19.3944
R16386 gnd.n4801 gnd.n4798 19.3944
R16387 gnd.n4798 gnd.n4797 19.3944
R16388 gnd.n4797 gnd.n4794 19.3944
R16389 gnd.n4794 gnd.n4793 19.3944
R16390 gnd.n4793 gnd.n4790 19.3944
R16391 gnd.n4790 gnd.n4789 19.3944
R16392 gnd.n4789 gnd.n4786 19.3944
R16393 gnd.n4786 gnd.n4785 19.3944
R16394 gnd.n4785 gnd.n4782 19.3944
R16395 gnd.n4782 gnd.n4781 19.3944
R16396 gnd.n4781 gnd.n4778 19.3944
R16397 gnd.n3222 gnd.n3188 19.3944
R16398 gnd.n3226 gnd.n3188 19.3944
R16399 gnd.n3229 gnd.n3226 19.3944
R16400 gnd.n3232 gnd.n3229 19.3944
R16401 gnd.n3232 gnd.n3186 19.3944
R16402 gnd.n3236 gnd.n3186 19.3944
R16403 gnd.n3239 gnd.n3236 19.3944
R16404 gnd.n3242 gnd.n3239 19.3944
R16405 gnd.n3242 gnd.n3184 19.3944
R16406 gnd.n3246 gnd.n3184 19.3944
R16407 gnd.n3249 gnd.n3246 19.3944
R16408 gnd.n3252 gnd.n3249 19.3944
R16409 gnd.n3252 gnd.n3182 19.3944
R16410 gnd.n3256 gnd.n3182 19.3944
R16411 gnd.n3259 gnd.n3256 19.3944
R16412 gnd.n3262 gnd.n3259 19.3944
R16413 gnd.n3262 gnd.n3180 19.3944
R16414 gnd.n3267 gnd.n3180 19.3944
R16415 gnd.n3200 gnd.n1619 19.3944
R16416 gnd.n3203 gnd.n3200 19.3944
R16417 gnd.n3203 gnd.n3195 19.3944
R16418 gnd.n3207 gnd.n3195 19.3944
R16419 gnd.n3210 gnd.n3207 19.3944
R16420 gnd.n3213 gnd.n3210 19.3944
R16421 gnd.n3213 gnd.n3193 19.3944
R16422 gnd.n3218 gnd.n3193 19.3944
R16423 gnd.n4776 gnd.n4773 19.3944
R16424 gnd.n4773 gnd.n4772 19.3944
R16425 gnd.n4772 gnd.n4769 19.3944
R16426 gnd.n4769 gnd.n4768 19.3944
R16427 gnd.n4768 gnd.n4765 19.3944
R16428 gnd.n4765 gnd.n4764 19.3944
R16429 gnd.n4764 gnd.n4761 19.3944
R16430 gnd.n4985 gnd.n1263 19.3944
R16431 gnd.n4985 gnd.n4984 19.3944
R16432 gnd.n4984 gnd.n4983 19.3944
R16433 gnd.n4983 gnd.n1268 19.3944
R16434 gnd.n4973 gnd.n1268 19.3944
R16435 gnd.n4973 gnd.n4972 19.3944
R16436 gnd.n4972 gnd.n4971 19.3944
R16437 gnd.n4971 gnd.n1291 19.3944
R16438 gnd.n4961 gnd.n1291 19.3944
R16439 gnd.n4961 gnd.n4960 19.3944
R16440 gnd.n4960 gnd.n4959 19.3944
R16441 gnd.n4959 gnd.n1309 19.3944
R16442 gnd.n4949 gnd.n1309 19.3944
R16443 gnd.n4949 gnd.n4948 19.3944
R16444 gnd.n4948 gnd.n4947 19.3944
R16445 gnd.n4947 gnd.n1329 19.3944
R16446 gnd.n4937 gnd.n1329 19.3944
R16447 gnd.n4937 gnd.n4936 19.3944
R16448 gnd.n4936 gnd.n4935 19.3944
R16449 gnd.n4935 gnd.n1347 19.3944
R16450 gnd.n4925 gnd.n1347 19.3944
R16451 gnd.n4925 gnd.n4924 19.3944
R16452 gnd.n4924 gnd.n4923 19.3944
R16453 gnd.n4923 gnd.n1367 19.3944
R16454 gnd.n4913 gnd.n1367 19.3944
R16455 gnd.n4913 gnd.n4912 19.3944
R16456 gnd.n4912 gnd.n4911 19.3944
R16457 gnd.n4901 gnd.n1400 19.3944
R16458 gnd.n2724 gnd.n1401 19.3944
R16459 gnd.n2653 gnd.n2652 19.3944
R16460 gnd.n2889 gnd.n2888 19.3944
R16461 gnd.n4898 gnd.n1407 19.3944
R16462 gnd.n4898 gnd.n1408 19.3944
R16463 gnd.n4888 gnd.n1408 19.3944
R16464 gnd.n4888 gnd.n4887 19.3944
R16465 gnd.n4887 gnd.n4886 19.3944
R16466 gnd.n4886 gnd.n1430 19.3944
R16467 gnd.n4876 gnd.n1430 19.3944
R16468 gnd.n4876 gnd.n4875 19.3944
R16469 gnd.n4875 gnd.n4874 19.3944
R16470 gnd.n4874 gnd.n1450 19.3944
R16471 gnd.n4864 gnd.n1450 19.3944
R16472 gnd.n4864 gnd.n4863 19.3944
R16473 gnd.n4863 gnd.n4862 19.3944
R16474 gnd.n4862 gnd.n1470 19.3944
R16475 gnd.n4852 gnd.n1470 19.3944
R16476 gnd.n4852 gnd.n4851 19.3944
R16477 gnd.n4851 gnd.n4850 19.3944
R16478 gnd.n4850 gnd.n1490 19.3944
R16479 gnd.n4840 gnd.n1490 19.3944
R16480 gnd.n4840 gnd.n4839 19.3944
R16481 gnd.n4839 gnd.n4838 19.3944
R16482 gnd.n4838 gnd.n1510 19.3944
R16483 gnd.n4828 gnd.n1510 19.3944
R16484 gnd.n4828 gnd.n4827 19.3944
R16485 gnd.n4827 gnd.n4826 19.3944
R16486 gnd.n4826 gnd.n1530 19.3944
R16487 gnd.n4816 gnd.n1530 19.3944
R16488 gnd.n4816 gnd.n4815 19.3944
R16489 gnd.n6742 gnd.n6741 19.3944
R16490 gnd.n6741 gnd.n6740 19.3944
R16491 gnd.n6740 gnd.n956 19.3944
R16492 gnd.n6734 gnd.n956 19.3944
R16493 gnd.n6734 gnd.n6733 19.3944
R16494 gnd.n6733 gnd.n6732 19.3944
R16495 gnd.n6732 gnd.n964 19.3944
R16496 gnd.n6726 gnd.n964 19.3944
R16497 gnd.n6726 gnd.n6725 19.3944
R16498 gnd.n6725 gnd.n6724 19.3944
R16499 gnd.n6724 gnd.n972 19.3944
R16500 gnd.n6718 gnd.n972 19.3944
R16501 gnd.n6718 gnd.n6717 19.3944
R16502 gnd.n6717 gnd.n6716 19.3944
R16503 gnd.n6716 gnd.n980 19.3944
R16504 gnd.n6710 gnd.n980 19.3944
R16505 gnd.n6710 gnd.n6709 19.3944
R16506 gnd.n6709 gnd.n6708 19.3944
R16507 gnd.n6708 gnd.n988 19.3944
R16508 gnd.n6702 gnd.n988 19.3944
R16509 gnd.n6702 gnd.n6701 19.3944
R16510 gnd.n6701 gnd.n6700 19.3944
R16511 gnd.n6700 gnd.n996 19.3944
R16512 gnd.n6694 gnd.n996 19.3944
R16513 gnd.n6694 gnd.n6693 19.3944
R16514 gnd.n6693 gnd.n6692 19.3944
R16515 gnd.n6692 gnd.n1004 19.3944
R16516 gnd.n6686 gnd.n1004 19.3944
R16517 gnd.n6686 gnd.n6685 19.3944
R16518 gnd.n6685 gnd.n6684 19.3944
R16519 gnd.n6684 gnd.n1012 19.3944
R16520 gnd.n6678 gnd.n1012 19.3944
R16521 gnd.n6678 gnd.n6677 19.3944
R16522 gnd.n6677 gnd.n6676 19.3944
R16523 gnd.n6676 gnd.n1020 19.3944
R16524 gnd.n6670 gnd.n1020 19.3944
R16525 gnd.n6670 gnd.n6669 19.3944
R16526 gnd.n6669 gnd.n6668 19.3944
R16527 gnd.n6668 gnd.n1028 19.3944
R16528 gnd.n6662 gnd.n1028 19.3944
R16529 gnd.n6662 gnd.n6661 19.3944
R16530 gnd.n6661 gnd.n6660 19.3944
R16531 gnd.n6660 gnd.n1036 19.3944
R16532 gnd.n6654 gnd.n1036 19.3944
R16533 gnd.n6654 gnd.n6653 19.3944
R16534 gnd.n6653 gnd.n6652 19.3944
R16535 gnd.n6652 gnd.n1044 19.3944
R16536 gnd.n6646 gnd.n1044 19.3944
R16537 gnd.n6646 gnd.n6645 19.3944
R16538 gnd.n6645 gnd.n6644 19.3944
R16539 gnd.n6644 gnd.n1052 19.3944
R16540 gnd.n6638 gnd.n1052 19.3944
R16541 gnd.n6638 gnd.n6637 19.3944
R16542 gnd.n6637 gnd.n6636 19.3944
R16543 gnd.n6636 gnd.n1060 19.3944
R16544 gnd.n6630 gnd.n1060 19.3944
R16545 gnd.n6630 gnd.n6629 19.3944
R16546 gnd.n6629 gnd.n6628 19.3944
R16547 gnd.n6628 gnd.n1068 19.3944
R16548 gnd.n6622 gnd.n1068 19.3944
R16549 gnd.n6622 gnd.n6621 19.3944
R16550 gnd.n6621 gnd.n6620 19.3944
R16551 gnd.n6620 gnd.n1076 19.3944
R16552 gnd.n6614 gnd.n1076 19.3944
R16553 gnd.n6614 gnd.n6613 19.3944
R16554 gnd.n6613 gnd.n6612 19.3944
R16555 gnd.n6612 gnd.n1084 19.3944
R16556 gnd.n6606 gnd.n1084 19.3944
R16557 gnd.n6606 gnd.n6605 19.3944
R16558 gnd.n6605 gnd.n6604 19.3944
R16559 gnd.n6604 gnd.n1092 19.3944
R16560 gnd.n6598 gnd.n1092 19.3944
R16561 gnd.n6598 gnd.n6597 19.3944
R16562 gnd.n6597 gnd.n6596 19.3944
R16563 gnd.n6596 gnd.n1100 19.3944
R16564 gnd.n6590 gnd.n1100 19.3944
R16565 gnd.n6590 gnd.n6589 19.3944
R16566 gnd.n6589 gnd.n6588 19.3944
R16567 gnd.n6588 gnd.n1108 19.3944
R16568 gnd.n6582 gnd.n1108 19.3944
R16569 gnd.n6582 gnd.n6581 19.3944
R16570 gnd.n6581 gnd.n6580 19.3944
R16571 gnd.n6580 gnd.n1116 19.3944
R16572 gnd.n2658 gnd.n1116 19.3944
R16573 gnd.n3045 gnd.n3037 19.3944
R16574 gnd.n3041 gnd.n3037 19.3944
R16575 gnd.n3041 gnd.n3040 19.3944
R16576 gnd.n3040 gnd.n2531 19.3944
R16577 gnd.n3381 gnd.n2531 19.3944
R16578 gnd.n3381 gnd.n2529 19.3944
R16579 gnd.n3385 gnd.n2529 19.3944
R16580 gnd.n3385 gnd.n2527 19.3944
R16581 gnd.n3389 gnd.n2527 19.3944
R16582 gnd.n3389 gnd.n2524 19.3944
R16583 gnd.n3402 gnd.n2524 19.3944
R16584 gnd.n3402 gnd.n2525 19.3944
R16585 gnd.n3398 gnd.n2525 19.3944
R16586 gnd.n3398 gnd.n3397 19.3944
R16587 gnd.n3397 gnd.n3396 19.3944
R16588 gnd.n3396 gnd.n2495 19.3944
R16589 gnd.n3540 gnd.n2495 19.3944
R16590 gnd.n3540 gnd.n2492 19.3944
R16591 gnd.n3555 gnd.n2492 19.3944
R16592 gnd.n3555 gnd.n2493 19.3944
R16593 gnd.n3551 gnd.n2493 19.3944
R16594 gnd.n3551 gnd.n3550 19.3944
R16595 gnd.n3550 gnd.n3549 19.3944
R16596 gnd.n3549 gnd.n3546 19.3944
R16597 gnd.n3546 gnd.n2446 19.3944
R16598 gnd.n3616 gnd.n2446 19.3944
R16599 gnd.n3616 gnd.n2443 19.3944
R16600 gnd.n3621 gnd.n2443 19.3944
R16601 gnd.n3621 gnd.n2444 19.3944
R16602 gnd.n2444 gnd.n2419 19.3944
R16603 gnd.n3655 gnd.n2419 19.3944
R16604 gnd.n3655 gnd.n2417 19.3944
R16605 gnd.n3659 gnd.n2417 19.3944
R16606 gnd.n3660 gnd.n3659 19.3944
R16607 gnd.n3663 gnd.n3660 19.3944
R16608 gnd.n3663 gnd.n2414 19.3944
R16609 gnd.n3670 gnd.n2414 19.3944
R16610 gnd.n3670 gnd.n2415 19.3944
R16611 gnd.n3666 gnd.n2415 19.3944
R16612 gnd.n3666 gnd.n2360 19.3944
R16613 gnd.n3751 gnd.n2360 19.3944
R16614 gnd.n3751 gnd.n2357 19.3944
R16615 gnd.n3781 gnd.n2357 19.3944
R16616 gnd.n3781 gnd.n2358 19.3944
R16617 gnd.n3777 gnd.n2358 19.3944
R16618 gnd.n3777 gnd.n3776 19.3944
R16619 gnd.n3776 gnd.n3775 19.3944
R16620 gnd.n3775 gnd.n3760 19.3944
R16621 gnd.n3771 gnd.n3760 19.3944
R16622 gnd.n3771 gnd.n3770 19.3944
R16623 gnd.n3770 gnd.n3769 19.3944
R16624 gnd.n3769 gnd.n3764 19.3944
R16625 gnd.n3765 gnd.n3764 19.3944
R16626 gnd.n3765 gnd.n2287 19.3944
R16627 gnd.n3901 gnd.n2287 19.3944
R16628 gnd.n3901 gnd.n2284 19.3944
R16629 gnd.n3906 gnd.n2284 19.3944
R16630 gnd.n3906 gnd.n2285 19.3944
R16631 gnd.n2285 gnd.n2263 19.3944
R16632 gnd.n3934 gnd.n2263 19.3944
R16633 gnd.n3934 gnd.n2260 19.3944
R16634 gnd.n3964 gnd.n2260 19.3944
R16635 gnd.n3964 gnd.n2261 19.3944
R16636 gnd.n3960 gnd.n2261 19.3944
R16637 gnd.n3960 gnd.n3959 19.3944
R16638 gnd.n3959 gnd.n3958 19.3944
R16639 gnd.n3958 gnd.n3941 19.3944
R16640 gnd.n3954 gnd.n3941 19.3944
R16641 gnd.n3954 gnd.n3953 19.3944
R16642 gnd.n3953 gnd.n3952 19.3944
R16643 gnd.n3952 gnd.n3947 19.3944
R16644 gnd.n3948 gnd.n3947 19.3944
R16645 gnd.n3948 gnd.n2124 19.3944
R16646 gnd.n4168 gnd.n2124 19.3944
R16647 gnd.n4168 gnd.n2122 19.3944
R16648 gnd.n4172 gnd.n2122 19.3944
R16649 gnd.n4172 gnd.n2112 19.3944
R16650 gnd.n4187 gnd.n2112 19.3944
R16651 gnd.n4187 gnd.n2110 19.3944
R16652 gnd.n4191 gnd.n2110 19.3944
R16653 gnd.n4191 gnd.n1797 19.3944
R16654 gnd.n4567 gnd.n1797 19.3944
R16655 gnd.n4564 gnd.n4563 19.3944
R16656 gnd.n4563 gnd.n4562 19.3944
R16657 gnd.n4562 gnd.n1802 19.3944
R16658 gnd.n4558 gnd.n1802 19.3944
R16659 gnd.n4558 gnd.n4557 19.3944
R16660 gnd.n4557 gnd.n4556 19.3944
R16661 gnd.n4556 gnd.n1807 19.3944
R16662 gnd.n4551 gnd.n1807 19.3944
R16663 gnd.n4551 gnd.n4550 19.3944
R16664 gnd.n4550 gnd.n1812 19.3944
R16665 gnd.n4543 gnd.n1812 19.3944
R16666 gnd.n4543 gnd.n4542 19.3944
R16667 gnd.n4542 gnd.n1821 19.3944
R16668 gnd.n4535 gnd.n1821 19.3944
R16669 gnd.n4535 gnd.n4534 19.3944
R16670 gnd.n4534 gnd.n1829 19.3944
R16671 gnd.n4527 gnd.n1829 19.3944
R16672 gnd.n4527 gnd.n4526 19.3944
R16673 gnd.n4526 gnd.n1837 19.3944
R16674 gnd.n4519 gnd.n1837 19.3944
R16675 gnd.n4519 gnd.n4518 19.3944
R16676 gnd.n4518 gnd.n1845 19.3944
R16677 gnd.n4511 gnd.n1845 19.3944
R16678 gnd.n4511 gnd.n4510 19.3944
R16679 gnd.n2098 gnd.n2077 19.3944
R16680 gnd.n4255 gnd.n2077 19.3944
R16681 gnd.n4255 gnd.n4254 19.3944
R16682 gnd.n4690 gnd.n4689 19.2005
R16683 gnd.n4154 gnd.n4153 19.2005
R16684 gnd.n3497 gnd.t100 19.1199
R16685 gnd.n3855 gnd.t99 19.1199
R16686 gnd.n5899 gnd.t121 18.8012
R16687 gnd.n5938 gnd.t279 18.8012
R16688 gnd.n5742 gnd.n5484 18.4825
R16689 gnd.n3557 gnd.n2484 18.4825
R16690 gnd.n3580 gnd.t111 18.4825
R16691 gnd.n3702 gnd.n2385 18.4825
R16692 gnd.n3802 gnd.n3801 18.4825
R16693 gnd.n3869 gnd.t78 18.4825
R16694 gnd.n3974 gnd.n2252 18.4825
R16695 gnd.t397 gnd.n2134 18.4825
R16696 gnd.n4449 gnd.n4448 18.4247
R16697 gnd.n4761 gnd.n4760 18.4247
R16698 gnd.n4507 gnd.n4506 18.2308
R16699 gnd.n3127 gnd.n2579 18.2308
R16700 gnd.n448 gnd.n445 18.2308
R16701 gnd.n2799 gnd.n2798 18.2308
R16702 gnd.t127 gnd.n5426 18.1639
R16703 gnd.n3944 gnd.t304 17.8452
R16704 gnd.n5455 gnd.t119 17.5266
R16705 gnd.n6576 gnd.n1118 17.2079
R16706 gnd.n2519 gnd.n2514 17.2079
R16707 gnd.n3538 gnd.n2498 17.2079
R16708 gnd.n3985 gnd.n3984 17.2079
R16709 gnd.n7337 gnd.n197 17.2079
R16710 gnd.t131 gnd.n5402 16.8893
R16711 gnd.n4756 gnd.n1658 16.8893
R16712 gnd.n4166 gnd.n2128 16.8893
R16713 gnd.n4431 gnd.n4428 16.6793
R16714 gnd.n7591 gnd.n7588 16.6793
R16715 gnd.n5038 gnd.n5035 16.6793
R16716 gnd.n3219 gnd.n3218 16.6793
R16717 gnd.n2649 gnd.n2641 16.5706
R16718 gnd.n4896 gnd.n1411 16.5706
R16719 gnd.n2930 gnd.n1414 16.5706
R16720 gnd.n2938 gnd.n1425 16.5706
R16721 gnd.n4884 gnd.n1432 16.5706
R16722 gnd.n2944 gnd.n2628 16.5706
R16723 gnd.n4878 gnd.n1441 16.5706
R16724 gnd.n4872 gnd.n1452 16.5706
R16725 gnd.n2987 gnd.n1455 16.5706
R16726 gnd.n2959 gnd.n1464 16.5706
R16727 gnd.n4860 gnd.n1472 16.5706
R16728 gnd.n2964 gnd.n2963 16.5706
R16729 gnd.n4854 gnd.n1481 16.5706
R16730 gnd.n4848 gnd.n1492 16.5706
R16731 gnd.n3011 gnd.n1495 16.5706
R16732 gnd.n3019 gnd.n1504 16.5706
R16733 gnd.n4836 gnd.n1512 16.5706
R16734 gnd.n3292 gnd.n3291 16.5706
R16735 gnd.n4830 gnd.n1521 16.5706
R16736 gnd.n3026 gnd.n1524 16.5706
R16737 gnd.n4824 gnd.n1532 16.5706
R16738 gnd.n3278 gnd.n1535 16.5706
R16739 gnd.n4818 gnd.n1542 16.5706
R16740 gnd.n3318 gnd.n1545 16.5706
R16741 gnd.n4380 gnd.n1973 16.5706
R16742 gnd.n4239 gnd.n4238 16.5706
R16743 gnd.n4372 gnd.n1982 16.5706
R16744 gnd.n4262 gnd.n1995 16.5706
R16745 gnd.n4366 gnd.n1998 16.5706
R16746 gnd.n4270 gnd.n2008 16.5706
R16747 gnd.n4360 gnd.n2011 16.5706
R16748 gnd.n4277 gnd.n2019 16.5706
R16749 gnd.n4354 gnd.n2022 16.5706
R16750 gnd.n4348 gnd.n2032 16.5706
R16751 gnd.n4300 gnd.n2040 16.5706
R16752 gnd.n4316 gnd.n2049 16.5706
R16753 gnd.n4336 gnd.n2052 16.5706
R16754 gnd.n4328 gnd.n4327 16.5706
R16755 gnd.n2055 gnd.n565 16.5706
R16756 gnd.n7370 gnd.n555 16.5706
R16757 gnd.n7393 gnd.n557 16.5706
R16758 gnd.n7402 gnd.n536 16.5706
R16759 gnd.n7419 gnd.n539 16.5706
R16760 gnd.n7406 gnd.n526 16.5706
R16761 gnd.n7430 gnd.n528 16.5706
R16762 gnd.n7438 gnd.n509 16.5706
R16763 gnd.n7452 gnd.n504 16.5706
R16764 gnd.n7446 gnd.n496 16.5706
R16765 gnd.t286 gnd.n5511 16.2519
R16766 gnd.n5369 gnd.t129 16.2519
R16767 gnd.n2900 gnd.t165 16.2519
R16768 gnd.n3337 gnd.t339 16.2519
R16769 gnd.t319 gnd.n1792 16.2519
R16770 gnd.n516 gnd.t35 16.2519
R16771 gnd.n3682 gnd.n2399 15.9333
R16772 gnd.n3826 gnd.n2324 15.9333
R16773 gnd.n2236 gnd.n2231 15.9333
R16774 gnd.t301 gnd.n4010 15.9333
R16775 gnd.n6368 gnd.n6366 15.6674
R16776 gnd.n6336 gnd.n6334 15.6674
R16777 gnd.n6304 gnd.n6302 15.6674
R16778 gnd.n6273 gnd.n6271 15.6674
R16779 gnd.n6241 gnd.n6239 15.6674
R16780 gnd.n6209 gnd.n6207 15.6674
R16781 gnd.n6177 gnd.n6175 15.6674
R16782 gnd.n6146 gnd.n6144 15.6674
R16783 gnd.n5629 gnd.t286 15.6146
R16784 gnd.t393 gnd.n5123 15.6146
R16785 gnd.t368 gnd.n6514 15.6146
R16786 gnd.t103 gnd.n1444 15.6146
R16787 gnd.t339 gnd.n2542 15.6146
R16788 gnd.n4193 gnd.t319 15.6146
R16789 gnd.t29 gnd.n548 15.6146
R16790 gnd.n4388 gnd.n4383 15.3217
R16791 gnd.n7546 gnd.n345 15.3217
R16792 gnd.n4995 gnd.n1251 15.3217
R16793 gnd.n3270 gnd.n3268 15.3217
R16794 gnd.n2891 gnd.n2649 15.296
R16795 gnd.n2900 gnd.n2641 15.296
R16796 gnd.n2899 gnd.n1411 15.296
R16797 gnd.n4896 gnd.n1414 15.296
R16798 gnd.n2930 gnd.n2929 15.296
R16799 gnd.n4890 gnd.n1425 15.296
R16800 gnd.n2938 gnd.n1432 15.296
R16801 gnd.n2944 gnd.n1441 15.296
R16802 gnd.n4878 gnd.n1444 15.296
R16803 gnd.n2952 gnd.n1452 15.296
R16804 gnd.n4872 gnd.n1455 15.296
R16805 gnd.n2988 gnd.n2987 15.296
R16806 gnd.n4866 gnd.n1464 15.296
R16807 gnd.n2959 gnd.n1472 15.296
R16808 gnd.n2964 gnd.n1481 15.296
R16809 gnd.n4854 gnd.n1484 15.296
R16810 gnd.n2973 gnd.n1492 15.296
R16811 gnd.n4848 gnd.n1495 15.296
R16812 gnd.n3011 gnd.n3010 15.296
R16813 gnd.n4842 gnd.n1504 15.296
R16814 gnd.n3019 gnd.n1512 15.296
R16815 gnd.n3291 gnd.n1521 15.296
R16816 gnd.n4830 gnd.n1524 15.296
R16817 gnd.n3026 gnd.n1532 15.296
R16818 gnd.n4824 gnd.n1535 15.296
R16819 gnd.n4818 gnd.n1545 15.296
R16820 gnd.n3318 gnd.n3317 15.296
R16821 gnd.n2466 gnd.t53 15.296
R16822 gnd.n3899 gnd.t117 15.296
R16823 gnd.n3997 gnd.t283 15.296
R16824 gnd.n4380 gnd.n1971 15.296
R16825 gnd.n4238 gnd.n1973 15.296
R16826 gnd.n4262 gnd.n1982 15.296
R16827 gnd.n4366 gnd.n1995 15.296
R16828 gnd.n4270 gnd.n1998 15.296
R16829 gnd.n4360 gnd.n2008 15.296
R16830 gnd.n4354 gnd.n2019 15.296
R16831 gnd.n4285 gnd.n2022 15.296
R16832 gnd.n4348 gnd.n2029 15.296
R16833 gnd.n4300 gnd.n2032 15.296
R16834 gnd.n4342 gnd.n2040 15.296
R16835 gnd.n4317 gnd.n4316 15.296
R16836 gnd.n4336 gnd.n2049 15.296
R16837 gnd.n4327 gnd.n2055 15.296
R16838 gnd.n7383 gnd.n565 15.296
R16839 gnd.n7370 gnd.n7369 15.296
R16840 gnd.n7393 gnd.n555 15.296
R16841 gnd.n7376 gnd.n557 15.296
R16842 gnd.n7402 gnd.n548 15.296
R16843 gnd.n7419 gnd.n536 15.296
R16844 gnd.n7430 gnd.n526 15.296
R16845 gnd.n7412 gnd.n528 15.296
R16846 gnd.n7438 gnd.n520 15.296
R16847 gnd.n7452 gnd.n509 15.296
R16848 gnd.n7457 gnd.n504 15.296
R16849 gnd.n7446 gnd.n516 15.296
R16850 gnd.n7465 gnd.n496 15.296
R16851 gnd.n2146 gnd.n2145 15.0827
R16852 gnd.n1670 gnd.n1665 15.0481
R16853 gnd.n2156 gnd.n2155 15.0481
R16854 gnd.n6065 gnd.t120 14.9773
R16855 gnd.t20 gnd.n1484 14.9773
R16856 gnd.n4756 gnd.n1626 14.9773
R16857 gnd.t93 gnd.n2394 14.9773
R16858 gnd.n2334 gnd.t152 14.9773
R16859 gnd.n4317 gnd.t37 14.9773
R16860 gnd.t378 gnd.n1658 14.6587
R16861 gnd.n3492 gnd.n2498 14.6587
R16862 gnd.n3636 gnd.n2435 14.6587
R16863 gnd.n2315 gnd.n2308 14.6587
R16864 gnd.n3985 gnd.n2241 14.6587
R16865 gnd.n4010 gnd.n2227 14.6587
R16866 gnd.n6111 gnd.t242 14.34
R16867 gnd.n6397 gnd.t118 14.34
R16868 gnd.n2520 gnd.t329 14.0214
R16869 gnd.t163 gnd.n5826 13.7027
R16870 gnd.n5711 gnd.n5707 13.5763
R16871 gnd.n6567 gnd.n1131 13.5763
R16872 gnd.n5743 gnd.n5742 13.384
R16873 gnd.n3481 gnd.n3404 13.384
R16874 gnd.n3565 gnd.n2484 13.384
R16875 gnd.n3624 gnd.n3623 13.384
R16876 gnd.n3644 gnd.t54 13.384
R16877 gnd.n3889 gnd.t115 13.384
R16878 gnd.n3887 gnd.n2299 13.384
R16879 gnd.n3966 gnd.n2252 13.384
R16880 gnd.n3945 gnd.n3944 13.384
R16881 gnd.n1681 gnd.n1662 13.1884
R16882 gnd.n1676 gnd.n1675 13.1884
R16883 gnd.n1675 gnd.n1674 13.1884
R16884 gnd.n2149 gnd.n2144 13.1884
R16885 gnd.n2150 gnd.n2149 13.1884
R16886 gnd.n1677 gnd.n1664 13.146
R16887 gnd.n1673 gnd.n1664 13.146
R16888 gnd.n2148 gnd.n2147 13.146
R16889 gnd.n2148 gnd.n2143 13.146
R16890 gnd.n3508 gnd.t87 13.0654
R16891 gnd.n2237 gnd.t71 13.0654
R16892 gnd.n6369 gnd.n6365 12.8005
R16893 gnd.n6337 gnd.n6333 12.8005
R16894 gnd.n6305 gnd.n6301 12.8005
R16895 gnd.n6274 gnd.n6270 12.8005
R16896 gnd.n6242 gnd.n6238 12.8005
R16897 gnd.n6210 gnd.n6206 12.8005
R16898 gnd.n6178 gnd.n6174 12.8005
R16899 gnd.n6147 gnd.n6143 12.8005
R16900 gnd.t353 gnd.n3527 12.7467
R16901 gnd.n4963 gnd.t16 12.4281
R16902 gnd.n4842 gnd.t69 12.4281
R16903 gnd.n4285 gnd.t184 12.4281
R16904 gnd.n7695 gnd.t32 12.4281
R16905 gnd.n5714 gnd.n5711 12.4126
R16906 gnd.n6563 gnd.n1131 12.4126
R16907 gnd.n4753 gnd.n4690 12.1761
R16908 gnd.n4153 gnd.n4152 12.1761
R16909 gnd.n4686 gnd.n1684 12.1094
R16910 gnd.n3574 gnd.n3573 12.1094
R16911 gnd.n3614 gnd.n2449 12.1094
R16912 gnd.n3880 gnd.n3879 12.1094
R16913 gnd.n3932 gnd.n2266 12.1094
R16914 gnd.n4157 gnd.n2138 12.1094
R16915 gnd.n6373 gnd.n6372 12.0247
R16916 gnd.n6341 gnd.n6340 12.0247
R16917 gnd.n6309 gnd.n6308 12.0247
R16918 gnd.n6278 gnd.n6277 12.0247
R16919 gnd.n6246 gnd.n6245 12.0247
R16920 gnd.n6214 gnd.n6213 12.0247
R16921 gnd.n6182 gnd.n6181 12.0247
R16922 gnd.n6151 gnd.n6150 12.0247
R16923 gnd.n4939 gnd.t4 11.7908
R16924 gnd.n4866 gnd.t18 11.7908
R16925 gnd.t312 gnd.n1542 11.7908
R16926 gnd.t168 gnd.t114 11.7908
R16927 gnd.t402 gnd.t113 11.7908
R16928 gnd.n4239 gnd.t293 11.7908
R16929 gnd.n7383 gnd.t14 11.7908
R16930 gnd.n7719 gnd.t135 11.7908
R16931 gnd.n3481 gnd.t362 11.4721
R16932 gnd.n3653 gnd.t107 11.4721
R16933 gnd.n3836 gnd.t7 11.4721
R16934 gnd.n6376 gnd.n6363 11.249
R16935 gnd.n6344 gnd.n6331 11.249
R16936 gnd.n6312 gnd.n6299 11.249
R16937 gnd.n6281 gnd.n6268 11.249
R16938 gnd.n6249 gnd.n6236 11.249
R16939 gnd.n6217 gnd.n6204 11.249
R16940 gnd.n6185 gnd.n6172 11.249
R16941 gnd.n6154 gnd.n6141 11.249
R16942 gnd.n5827 gnd.t163 11.1535
R16943 gnd.n4915 gnd.t39 11.1535
R16944 gnd.n4890 gnd.t105 11.1535
R16945 gnd.n2534 gnd.t49 11.1535
R16946 gnd.n3642 gnd.t228 11.1535
R16947 gnd.t148 gnd.n2296 11.1535
R16948 gnd.n4174 gnd.t230 11.1535
R16949 gnd.n7412 gnd.t143 11.1535
R16950 gnd.n7743 gnd.t196 11.1535
R16951 gnd.n3604 gnd.n2456 10.8348
R16952 gnd.n3604 gnd.n3603 10.8348
R16953 gnd.n3749 gnd.n2362 10.8348
R16954 gnd.n3749 gnd.n2363 10.8348
R16955 gnd.n3922 gnd.n2273 10.8348
R16956 gnd.n3922 gnd.n3921 10.8348
R16957 gnd.n4391 gnd.n4388 10.6672
R16958 gnd.n7549 gnd.n7546 10.6672
R16959 gnd.n4998 gnd.n4995 10.6672
R16960 gnd.n3268 gnd.n3267 10.6672
R16961 gnd.n4087 gnd.n2186 10.6151
R16962 gnd.n4087 gnd.n4086 10.6151
R16963 gnd.n4084 gnd.n2190 10.6151
R16964 gnd.n4079 gnd.n2190 10.6151
R16965 gnd.n4079 gnd.n4078 10.6151
R16966 gnd.n4078 gnd.n4077 10.6151
R16967 gnd.n4077 gnd.n2193 10.6151
R16968 gnd.n4072 gnd.n2193 10.6151
R16969 gnd.n4072 gnd.n4071 10.6151
R16970 gnd.n4071 gnd.n4070 10.6151
R16971 gnd.n4070 gnd.n2196 10.6151
R16972 gnd.n4065 gnd.n2196 10.6151
R16973 gnd.n4065 gnd.n4064 10.6151
R16974 gnd.n4064 gnd.n4063 10.6151
R16975 gnd.n4063 gnd.n2199 10.6151
R16976 gnd.n4058 gnd.n2199 10.6151
R16977 gnd.n4058 gnd.n4057 10.6151
R16978 gnd.n4057 gnd.n4056 10.6151
R16979 gnd.n4056 gnd.n2202 10.6151
R16980 gnd.n4051 gnd.n2202 10.6151
R16981 gnd.n4051 gnd.n4050 10.6151
R16982 gnd.n4050 gnd.n4049 10.6151
R16983 gnd.n4049 gnd.n2205 10.6151
R16984 gnd.n4044 gnd.n2205 10.6151
R16985 gnd.n4044 gnd.n4043 10.6151
R16986 gnd.n4043 gnd.n4042 10.6151
R16987 gnd.n4042 gnd.n2208 10.6151
R16988 gnd.n4037 gnd.n2208 10.6151
R16989 gnd.n4037 gnd.n4036 10.6151
R16990 gnd.n4036 gnd.n4035 10.6151
R16991 gnd.n3475 gnd.n3474 10.6151
R16992 gnd.n3477 gnd.n3475 10.6151
R16993 gnd.n3478 gnd.n3477 10.6151
R16994 gnd.n3479 gnd.n3478 10.6151
R16995 gnd.n3479 gnd.n2517 10.6151
R16996 gnd.n3489 gnd.n2517 10.6151
R16997 gnd.n3490 gnd.n3489 10.6151
R16998 gnd.n3514 gnd.n3490 10.6151
R16999 gnd.n3514 gnd.n3513 10.6151
R17000 gnd.n3513 gnd.n3512 10.6151
R17001 gnd.n3512 gnd.n3511 10.6151
R17002 gnd.n3511 gnd.n3491 10.6151
R17003 gnd.n3505 gnd.n3491 10.6151
R17004 gnd.n3505 gnd.n3504 10.6151
R17005 gnd.n3504 gnd.n3503 10.6151
R17006 gnd.n3503 gnd.n3502 10.6151
R17007 gnd.n3502 gnd.n3500 10.6151
R17008 gnd.n3500 gnd.n3499 10.6151
R17009 gnd.n3499 gnd.n3496 10.6151
R17010 gnd.n3496 gnd.n3495 10.6151
R17011 gnd.n3495 gnd.n2468 10.6151
R17012 gnd.n3583 gnd.n2468 10.6151
R17013 gnd.n3584 gnd.n3583 10.6151
R17014 gnd.n3585 gnd.n3584 10.6151
R17015 gnd.n3591 gnd.n3585 10.6151
R17016 gnd.n3592 gnd.n3591 10.6151
R17017 gnd.n3593 gnd.n3592 10.6151
R17018 gnd.n3593 gnd.n2439 10.6151
R17019 gnd.n3626 gnd.n2439 10.6151
R17020 gnd.n3627 gnd.n3626 10.6151
R17021 gnd.n3628 gnd.n3627 10.6151
R17022 gnd.n3634 gnd.n3628 10.6151
R17023 gnd.n3634 gnd.n3633 10.6151
R17024 gnd.n3633 gnd.n3632 10.6151
R17025 gnd.n3632 gnd.n3629 10.6151
R17026 gnd.n3629 gnd.n2391 10.6151
R17027 gnd.n3690 gnd.n2391 10.6151
R17028 gnd.n3691 gnd.n3690 10.6151
R17029 gnd.n3693 gnd.n3691 10.6151
R17030 gnd.n3693 gnd.n3692 10.6151
R17031 gnd.n3692 gnd.n2383 10.6151
R17032 gnd.n3705 gnd.n2383 10.6151
R17033 gnd.n3706 gnd.n3705 10.6151
R17034 gnd.n3723 gnd.n3706 10.6151
R17035 gnd.n3723 gnd.n3722 10.6151
R17036 gnd.n3722 gnd.n3721 10.6151
R17037 gnd.n3721 gnd.n3707 10.6151
R17038 gnd.n3717 gnd.n3707 10.6151
R17039 gnd.n3717 gnd.n3716 10.6151
R17040 gnd.n3716 gnd.n3715 10.6151
R17041 gnd.n3715 gnd.n3714 10.6151
R17042 gnd.n3714 gnd.n3712 10.6151
R17043 gnd.n3712 gnd.n3711 10.6151
R17044 gnd.n3711 gnd.n3709 10.6151
R17045 gnd.n3709 gnd.n2331 10.6151
R17046 gnd.n3810 gnd.n2331 10.6151
R17047 gnd.n3811 gnd.n3810 10.6151
R17048 gnd.n3818 gnd.n3811 10.6151
R17049 gnd.n3818 gnd.n3817 10.6151
R17050 gnd.n3817 gnd.n3816 10.6151
R17051 gnd.n3816 gnd.n3815 10.6151
R17052 gnd.n3815 gnd.n3813 10.6151
R17053 gnd.n3813 gnd.n3812 10.6151
R17054 gnd.n3812 gnd.n2306 10.6151
R17055 gnd.n3846 gnd.n2306 10.6151
R17056 gnd.n3847 gnd.n3846 10.6151
R17057 gnd.n3850 gnd.n3847 10.6151
R17058 gnd.n3851 gnd.n3850 10.6151
R17059 gnd.n3877 gnd.n3851 10.6151
R17060 gnd.n3877 gnd.n3876 10.6151
R17061 gnd.n3876 gnd.n3875 10.6151
R17062 gnd.n3875 gnd.n3874 10.6151
R17063 gnd.n3874 gnd.n3872 10.6151
R17064 gnd.n3872 gnd.n3871 10.6151
R17065 gnd.n3871 gnd.n3852 10.6151
R17066 gnd.n3866 gnd.n3852 10.6151
R17067 gnd.n3866 gnd.n3865 10.6151
R17068 gnd.n3865 gnd.n3864 10.6151
R17069 gnd.n3864 gnd.n3863 10.6151
R17070 gnd.n3863 gnd.n3861 10.6151
R17071 gnd.n3861 gnd.n3860 10.6151
R17072 gnd.n3860 gnd.n3857 10.6151
R17073 gnd.n3857 gnd.n2234 10.6151
R17074 gnd.n3993 gnd.n2234 10.6151
R17075 gnd.n3994 gnd.n3993 10.6151
R17076 gnd.n4002 gnd.n3994 10.6151
R17077 gnd.n4002 gnd.n4001 10.6151
R17078 gnd.n4001 gnd.n4000 10.6151
R17079 gnd.n4000 gnd.n3999 10.6151
R17080 gnd.n3999 gnd.n3996 10.6151
R17081 gnd.n3996 gnd.n3995 10.6151
R17082 gnd.n3995 gnd.n2211 10.6151
R17083 gnd.n4029 gnd.n2211 10.6151
R17084 gnd.n4030 gnd.n4029 10.6151
R17085 gnd.n4031 gnd.n4030 10.6151
R17086 gnd.n3409 gnd.n1622 10.6151
R17087 gnd.n3412 gnd.n3409 10.6151
R17088 gnd.n3417 gnd.n3414 10.6151
R17089 gnd.n3418 gnd.n3417 10.6151
R17090 gnd.n3421 gnd.n3418 10.6151
R17091 gnd.n3422 gnd.n3421 10.6151
R17092 gnd.n3425 gnd.n3422 10.6151
R17093 gnd.n3426 gnd.n3425 10.6151
R17094 gnd.n3429 gnd.n3426 10.6151
R17095 gnd.n3430 gnd.n3429 10.6151
R17096 gnd.n3433 gnd.n3430 10.6151
R17097 gnd.n3434 gnd.n3433 10.6151
R17098 gnd.n3437 gnd.n3434 10.6151
R17099 gnd.n3438 gnd.n3437 10.6151
R17100 gnd.n3441 gnd.n3438 10.6151
R17101 gnd.n3442 gnd.n3441 10.6151
R17102 gnd.n3445 gnd.n3442 10.6151
R17103 gnd.n3446 gnd.n3445 10.6151
R17104 gnd.n3449 gnd.n3446 10.6151
R17105 gnd.n3450 gnd.n3449 10.6151
R17106 gnd.n3453 gnd.n3450 10.6151
R17107 gnd.n3454 gnd.n3453 10.6151
R17108 gnd.n3457 gnd.n3454 10.6151
R17109 gnd.n3458 gnd.n3457 10.6151
R17110 gnd.n3461 gnd.n3458 10.6151
R17111 gnd.n3462 gnd.n3461 10.6151
R17112 gnd.n3465 gnd.n3462 10.6151
R17113 gnd.n3466 gnd.n3465 10.6151
R17114 gnd.n3469 gnd.n3466 10.6151
R17115 gnd.n3470 gnd.n3469 10.6151
R17116 gnd.n4753 gnd.n4752 10.6151
R17117 gnd.n4752 gnd.n4751 10.6151
R17118 gnd.n4751 gnd.n4750 10.6151
R17119 gnd.n4750 gnd.n4748 10.6151
R17120 gnd.n4748 gnd.n4745 10.6151
R17121 gnd.n4745 gnd.n4744 10.6151
R17122 gnd.n4744 gnd.n4741 10.6151
R17123 gnd.n4741 gnd.n4740 10.6151
R17124 gnd.n4740 gnd.n4737 10.6151
R17125 gnd.n4737 gnd.n4736 10.6151
R17126 gnd.n4736 gnd.n4733 10.6151
R17127 gnd.n4733 gnd.n4732 10.6151
R17128 gnd.n4732 gnd.n4729 10.6151
R17129 gnd.n4729 gnd.n4728 10.6151
R17130 gnd.n4728 gnd.n4725 10.6151
R17131 gnd.n4725 gnd.n4724 10.6151
R17132 gnd.n4724 gnd.n4721 10.6151
R17133 gnd.n4721 gnd.n4720 10.6151
R17134 gnd.n4720 gnd.n4717 10.6151
R17135 gnd.n4717 gnd.n4716 10.6151
R17136 gnd.n4716 gnd.n4713 10.6151
R17137 gnd.n4713 gnd.n4712 10.6151
R17138 gnd.n4712 gnd.n4709 10.6151
R17139 gnd.n4709 gnd.n4708 10.6151
R17140 gnd.n4708 gnd.n4705 10.6151
R17141 gnd.n4705 gnd.n4704 10.6151
R17142 gnd.n4704 gnd.n4701 10.6151
R17143 gnd.n4701 gnd.n4700 10.6151
R17144 gnd.n4697 gnd.n4696 10.6151
R17145 gnd.n4696 gnd.n1623 10.6151
R17146 gnd.n4152 gnd.n2161 10.6151
R17147 gnd.n2162 gnd.n2161 10.6151
R17148 gnd.n4145 gnd.n2162 10.6151
R17149 gnd.n4145 gnd.n4144 10.6151
R17150 gnd.n4144 gnd.n4143 10.6151
R17151 gnd.n4143 gnd.n2164 10.6151
R17152 gnd.n4138 gnd.n2164 10.6151
R17153 gnd.n4138 gnd.n4137 10.6151
R17154 gnd.n4137 gnd.n4136 10.6151
R17155 gnd.n4136 gnd.n2167 10.6151
R17156 gnd.n4131 gnd.n2167 10.6151
R17157 gnd.n4131 gnd.n4130 10.6151
R17158 gnd.n4130 gnd.n4129 10.6151
R17159 gnd.n4129 gnd.n2170 10.6151
R17160 gnd.n4124 gnd.n2170 10.6151
R17161 gnd.n4124 gnd.n4123 10.6151
R17162 gnd.n4123 gnd.n4122 10.6151
R17163 gnd.n4122 gnd.n2173 10.6151
R17164 gnd.n4117 gnd.n2173 10.6151
R17165 gnd.n4117 gnd.n4116 10.6151
R17166 gnd.n4116 gnd.n4115 10.6151
R17167 gnd.n4115 gnd.n2176 10.6151
R17168 gnd.n4110 gnd.n2176 10.6151
R17169 gnd.n4110 gnd.n4109 10.6151
R17170 gnd.n4109 gnd.n4108 10.6151
R17171 gnd.n4108 gnd.n2179 10.6151
R17172 gnd.n4103 gnd.n2179 10.6151
R17173 gnd.n4103 gnd.n4102 10.6151
R17174 gnd.n4100 gnd.n2184 10.6151
R17175 gnd.n4095 gnd.n2184 10.6151
R17176 gnd.n4689 gnd.n4688 10.6151
R17177 gnd.n4688 gnd.n1682 10.6151
R17178 gnd.n2522 gnd.n1682 10.6151
R17179 gnd.n3483 gnd.n2522 10.6151
R17180 gnd.n3484 gnd.n3483 10.6151
R17181 gnd.n3485 gnd.n3484 10.6151
R17182 gnd.n3485 gnd.n2512 10.6151
R17183 gnd.n3518 gnd.n2512 10.6151
R17184 gnd.n3519 gnd.n3518 10.6151
R17185 gnd.n3525 gnd.n3519 10.6151
R17186 gnd.n3525 gnd.n3524 10.6151
R17187 gnd.n3524 gnd.n3523 10.6151
R17188 gnd.n3523 gnd.n3520 10.6151
R17189 gnd.n3520 gnd.n2488 10.6151
R17190 gnd.n3560 gnd.n2488 10.6151
R17191 gnd.n3561 gnd.n3560 10.6151
R17192 gnd.n3562 gnd.n3561 10.6151
R17193 gnd.n3562 gnd.n2472 10.6151
R17194 gnd.n3576 gnd.n2472 10.6151
R17195 gnd.n3577 gnd.n3576 10.6151
R17196 gnd.n3578 gnd.n3577 10.6151
R17197 gnd.n3578 gnd.n2461 10.6151
R17198 gnd.n3601 gnd.n2461 10.6151
R17199 gnd.n3601 gnd.n3600 10.6151
R17200 gnd.n3600 gnd.n3599 10.6151
R17201 gnd.n3599 gnd.n2462 10.6151
R17202 gnd.n2465 gnd.n2462 10.6151
R17203 gnd.n2465 gnd.n2464 10.6151
R17204 gnd.n2464 gnd.n2432 10.6151
R17205 gnd.n3640 gnd.n2432 10.6151
R17206 gnd.n3640 gnd.n3639 10.6151
R17207 gnd.n3639 gnd.n3638 10.6151
R17208 gnd.n3638 gnd.n2433 10.6151
R17209 gnd.n2433 gnd.n2397 10.6151
R17210 gnd.n3684 gnd.n2397 10.6151
R17211 gnd.n3685 gnd.n3684 10.6151
R17212 gnd.n3686 gnd.n3685 10.6151
R17213 gnd.n3686 gnd.n2387 10.6151
R17214 gnd.n3698 gnd.n2387 10.6151
R17215 gnd.n3699 gnd.n3698 10.6151
R17216 gnd.n3700 gnd.n3699 10.6151
R17217 gnd.n3700 gnd.n2378 10.6151
R17218 gnd.n3729 gnd.n2378 10.6151
R17219 gnd.n3730 gnd.n3729 10.6151
R17220 gnd.n3736 gnd.n3730 10.6151
R17221 gnd.n3736 gnd.n3735 10.6151
R17222 gnd.n3735 gnd.n3734 10.6151
R17223 gnd.n3734 gnd.n3731 10.6151
R17224 gnd.n3731 gnd.n2352 10.6151
R17225 gnd.n3786 gnd.n2352 10.6151
R17226 gnd.n3787 gnd.n3786 10.6151
R17227 gnd.n3788 gnd.n3787 10.6151
R17228 gnd.n3788 gnd.n2337 10.6151
R17229 gnd.n3804 gnd.n2337 10.6151
R17230 gnd.n3805 gnd.n3804 10.6151
R17231 gnd.n3806 gnd.n3805 10.6151
R17232 gnd.n3806 gnd.n2326 10.6151
R17233 gnd.n3822 gnd.n2326 10.6151
R17234 gnd.n3823 gnd.n3822 10.6151
R17235 gnd.n3824 gnd.n3823 10.6151
R17236 gnd.n3824 gnd.n2310 10.6151
R17237 gnd.n3839 gnd.n2310 10.6151
R17238 gnd.n3840 gnd.n3839 10.6151
R17239 gnd.n3841 gnd.n3840 10.6151
R17240 gnd.n3841 gnd.n2302 10.6151
R17241 gnd.n3885 gnd.n2302 10.6151
R17242 gnd.n3885 gnd.n3884 10.6151
R17243 gnd.n3884 gnd.n3883 10.6151
R17244 gnd.n3883 gnd.n2303 10.6151
R17245 gnd.n2303 gnd.n2279 10.6151
R17246 gnd.n3912 gnd.n2279 10.6151
R17247 gnd.n3913 gnd.n3912 10.6151
R17248 gnd.n3919 gnd.n3913 10.6151
R17249 gnd.n3919 gnd.n3918 10.6151
R17250 gnd.n3918 gnd.n3917 10.6151
R17251 gnd.n3917 gnd.n3914 10.6151
R17252 gnd.n3914 gnd.n2256 10.6151
R17253 gnd.n3969 gnd.n2256 10.6151
R17254 gnd.n3970 gnd.n3969 10.6151
R17255 gnd.n3971 gnd.n3970 10.6151
R17256 gnd.n3971 gnd.n2239 10.6151
R17257 gnd.n3987 gnd.n2239 10.6151
R17258 gnd.n3988 gnd.n3987 10.6151
R17259 gnd.n3989 gnd.n3988 10.6151
R17260 gnd.n3989 gnd.n2229 10.6151
R17261 gnd.n4006 gnd.n2229 10.6151
R17262 gnd.n4007 gnd.n4006 10.6151
R17263 gnd.n4008 gnd.n4007 10.6151
R17264 gnd.n4008 gnd.n2214 10.6151
R17265 gnd.n4022 gnd.n2214 10.6151
R17266 gnd.n4023 gnd.n4022 10.6151
R17267 gnd.n4024 gnd.n4023 10.6151
R17268 gnd.n4024 gnd.n2141 10.6151
R17269 gnd.n4155 gnd.n2141 10.6151
R17270 gnd.n4155 gnd.n4154 10.6151
R17271 gnd.n5499 gnd.t207 10.5161
R17272 gnd.n6094 gnd.t242 10.5161
R17273 gnd.t118 gnd.n6396 10.5161
R17274 gnd.n2726 gnd.t139 10.5161
R17275 gnd.n2885 gnd.n2660 10.5161
R17276 gnd.n2885 gnd.t12 10.5161
R17277 gnd.n2436 gnd.t228 10.5161
R17278 gnd.n3843 gnd.t148 10.5161
R17279 gnd.n7473 gnd.t141 10.5161
R17280 gnd.n7473 gnd.n494 10.5161
R17281 gnd.n7482 gnd.t63 10.5161
R17282 gnd.n6377 gnd.n6361 10.4732
R17283 gnd.n6345 gnd.n6329 10.4732
R17284 gnd.n6313 gnd.n6297 10.4732
R17285 gnd.n6282 gnd.n6266 10.4732
R17286 gnd.n6250 gnd.n6234 10.4732
R17287 gnd.n6218 gnd.n6202 10.4732
R17288 gnd.n6186 gnd.n6170 10.4732
R17289 gnd.n6155 gnd.n6139 10.4732
R17290 gnd.t323 gnd.n2127 10.1975
R17291 gnd.t120 gnd.n5196 9.87883
R17292 gnd.n4921 gnd.t22 9.87883
R17293 gnd.n4884 gnd.t0 9.87883
R17294 gnd.n7406 gnd.t58 9.87883
R17295 gnd.n7737 gnd.t24 9.87883
R17296 gnd.n6381 gnd.n6380 9.69747
R17297 gnd.n6349 gnd.n6348 9.69747
R17298 gnd.n6317 gnd.n6316 9.69747
R17299 gnd.n6286 gnd.n6285 9.69747
R17300 gnd.n6254 gnd.n6253 9.69747
R17301 gnd.n6222 gnd.n6221 9.69747
R17302 gnd.n6190 gnd.n6189 9.69747
R17303 gnd.n6159 gnd.n6158 9.69747
R17304 gnd.n3472 gnd.n1684 9.56018
R17305 gnd.n3573 gnd.n2478 9.56018
R17306 gnd.n3614 gnd.n2448 9.56018
R17307 gnd.t92 gnd.n3681 9.56018
R17308 gnd.n3739 gnd.n3738 9.56018
R17309 gnd.n3784 gnd.n3783 9.56018
R17310 gnd.n3828 gnd.t79 9.56018
R17311 gnd.n3879 gnd.n2281 9.56018
R17312 gnd.n3932 gnd.n2265 9.56018
R17313 gnd.n6387 gnd.n6386 9.45567
R17314 gnd.n6355 gnd.n6354 9.45567
R17315 gnd.n6323 gnd.n6322 9.45567
R17316 gnd.n6292 gnd.n6291 9.45567
R17317 gnd.n6260 gnd.n6259 9.45567
R17318 gnd.n6228 gnd.n6227 9.45567
R17319 gnd.n6196 gnd.n6195 9.45567
R17320 gnd.n6165 gnd.n6164 9.45567
R17321 gnd.n4428 gnd.n4427 9.30959
R17322 gnd.n7588 gnd.n325 9.30959
R17323 gnd.n5035 gnd.n5034 9.30959
R17324 gnd.n3222 gnd.n3219 9.30959
R17325 gnd.n6386 gnd.n6385 9.3005
R17326 gnd.n6359 gnd.n6358 9.3005
R17327 gnd.n6380 gnd.n6379 9.3005
R17328 gnd.n6378 gnd.n6377 9.3005
R17329 gnd.n6363 gnd.n6362 9.3005
R17330 gnd.n6372 gnd.n6371 9.3005
R17331 gnd.n6370 gnd.n6369 9.3005
R17332 gnd.n6354 gnd.n6353 9.3005
R17333 gnd.n6327 gnd.n6326 9.3005
R17334 gnd.n6348 gnd.n6347 9.3005
R17335 gnd.n6346 gnd.n6345 9.3005
R17336 gnd.n6331 gnd.n6330 9.3005
R17337 gnd.n6340 gnd.n6339 9.3005
R17338 gnd.n6338 gnd.n6337 9.3005
R17339 gnd.n6322 gnd.n6321 9.3005
R17340 gnd.n6295 gnd.n6294 9.3005
R17341 gnd.n6316 gnd.n6315 9.3005
R17342 gnd.n6314 gnd.n6313 9.3005
R17343 gnd.n6299 gnd.n6298 9.3005
R17344 gnd.n6308 gnd.n6307 9.3005
R17345 gnd.n6306 gnd.n6305 9.3005
R17346 gnd.n6291 gnd.n6290 9.3005
R17347 gnd.n6264 gnd.n6263 9.3005
R17348 gnd.n6285 gnd.n6284 9.3005
R17349 gnd.n6283 gnd.n6282 9.3005
R17350 gnd.n6268 gnd.n6267 9.3005
R17351 gnd.n6277 gnd.n6276 9.3005
R17352 gnd.n6275 gnd.n6274 9.3005
R17353 gnd.n6259 gnd.n6258 9.3005
R17354 gnd.n6232 gnd.n6231 9.3005
R17355 gnd.n6253 gnd.n6252 9.3005
R17356 gnd.n6251 gnd.n6250 9.3005
R17357 gnd.n6236 gnd.n6235 9.3005
R17358 gnd.n6245 gnd.n6244 9.3005
R17359 gnd.n6243 gnd.n6242 9.3005
R17360 gnd.n6227 gnd.n6226 9.3005
R17361 gnd.n6200 gnd.n6199 9.3005
R17362 gnd.n6221 gnd.n6220 9.3005
R17363 gnd.n6219 gnd.n6218 9.3005
R17364 gnd.n6204 gnd.n6203 9.3005
R17365 gnd.n6213 gnd.n6212 9.3005
R17366 gnd.n6211 gnd.n6210 9.3005
R17367 gnd.n6195 gnd.n6194 9.3005
R17368 gnd.n6168 gnd.n6167 9.3005
R17369 gnd.n6189 gnd.n6188 9.3005
R17370 gnd.n6187 gnd.n6186 9.3005
R17371 gnd.n6172 gnd.n6171 9.3005
R17372 gnd.n6181 gnd.n6180 9.3005
R17373 gnd.n6179 gnd.n6178 9.3005
R17374 gnd.n6164 gnd.n6163 9.3005
R17375 gnd.n6137 gnd.n6136 9.3005
R17376 gnd.n6158 gnd.n6157 9.3005
R17377 gnd.n6156 gnd.n6155 9.3005
R17378 gnd.n6141 gnd.n6140 9.3005
R17379 gnd.n6150 gnd.n6149 9.3005
R17380 gnd.n6148 gnd.n6147 9.3005
R17381 gnd.n6556 gnd.n6555 9.3005
R17382 gnd.n6554 gnd.n6522 9.3005
R17383 gnd.n6553 gnd.n6552 9.3005
R17384 gnd.n6549 gnd.n6523 9.3005
R17385 gnd.n6546 gnd.n6524 9.3005
R17386 gnd.n6545 gnd.n6525 9.3005
R17387 gnd.n6542 gnd.n6526 9.3005
R17388 gnd.n6541 gnd.n6527 9.3005
R17389 gnd.n6538 gnd.n6528 9.3005
R17390 gnd.n6537 gnd.n6529 9.3005
R17391 gnd.n6534 gnd.n6530 9.3005
R17392 gnd.n6533 gnd.n6531 9.3005
R17393 gnd.n1133 gnd.n1132 9.3005
R17394 gnd.n6564 gnd.n6563 9.3005
R17395 gnd.n6565 gnd.n1131 9.3005
R17396 gnd.n6567 gnd.n6566 9.3005
R17397 gnd.n6557 gnd.n6521 9.3005
R17398 gnd.n5766 gnd.n5765 9.3005
R17399 gnd.n5767 gnd.n5469 9.3005
R17400 gnd.n5769 gnd.n5768 9.3005
R17401 gnd.n5450 gnd.n5449 9.3005
R17402 gnd.n5796 gnd.n5795 9.3005
R17403 gnd.n5797 gnd.n5448 9.3005
R17404 gnd.n5801 gnd.n5798 9.3005
R17405 gnd.n5800 gnd.n5799 9.3005
R17406 gnd.n5424 gnd.n5423 9.3005
R17407 gnd.n5830 gnd.n5829 9.3005
R17408 gnd.n5831 gnd.n5422 9.3005
R17409 gnd.n5838 gnd.n5832 9.3005
R17410 gnd.n5837 gnd.n5833 9.3005
R17411 gnd.n5836 gnd.n5834 9.3005
R17412 gnd.n5391 gnd.n5390 9.3005
R17413 gnd.n5891 gnd.n5890 9.3005
R17414 gnd.n5892 gnd.n5389 9.3005
R17415 gnd.n5896 gnd.n5893 9.3005
R17416 gnd.n5895 gnd.n5894 9.3005
R17417 gnd.n5364 gnd.n5363 9.3005
R17418 gnd.n5931 gnd.n5930 9.3005
R17419 gnd.n5932 gnd.n5362 9.3005
R17420 gnd.n5936 gnd.n5933 9.3005
R17421 gnd.n5935 gnd.n5934 9.3005
R17422 gnd.n5257 gnd.n5256 9.3005
R17423 gnd.n5973 gnd.n5972 9.3005
R17424 gnd.n5974 gnd.n5255 9.3005
R17425 gnd.n5978 gnd.n5975 9.3005
R17426 gnd.n5977 gnd.n5976 9.3005
R17427 gnd.n5227 gnd.n5226 9.3005
R17428 gnd.n6014 gnd.n6013 9.3005
R17429 gnd.n6015 gnd.n5225 9.3005
R17430 gnd.n6019 gnd.n6016 9.3005
R17431 gnd.n6018 gnd.n6017 9.3005
R17432 gnd.n5201 gnd.n5200 9.3005
R17433 gnd.n6058 gnd.n6057 9.3005
R17434 gnd.n6059 gnd.n5199 9.3005
R17435 gnd.n6063 gnd.n6060 9.3005
R17436 gnd.n6062 gnd.n6061 9.3005
R17437 gnd.n5174 gnd.n5173 9.3005
R17438 gnd.n6104 gnd.n6103 9.3005
R17439 gnd.n6105 gnd.n5172 9.3005
R17440 gnd.n6109 gnd.n6106 9.3005
R17441 gnd.n6108 gnd.n6107 9.3005
R17442 gnd.n5147 gnd.n5146 9.3005
R17443 gnd.n6400 gnd.n6399 9.3005
R17444 gnd.n6401 gnd.n5145 9.3005
R17445 gnd.n6408 gnd.n6402 9.3005
R17446 gnd.n6407 gnd.n6403 9.3005
R17447 gnd.n6406 gnd.n6405 9.3005
R17448 gnd.n6404 gnd.n5121 9.3005
R17449 gnd.n6518 gnd.n5120 9.3005
R17450 gnd.n6520 gnd.n6519 9.3005
R17451 gnd.n5471 gnd.n5470 9.3005
R17452 gnd.n5711 gnd.n5710 9.3005
R17453 gnd.n5714 gnd.n5706 9.3005
R17454 gnd.n5715 gnd.n5705 9.3005
R17455 gnd.n5718 gnd.n5704 9.3005
R17456 gnd.n5719 gnd.n5703 9.3005
R17457 gnd.n5722 gnd.n5702 9.3005
R17458 gnd.n5723 gnd.n5701 9.3005
R17459 gnd.n5726 gnd.n5700 9.3005
R17460 gnd.n5727 gnd.n5699 9.3005
R17461 gnd.n5730 gnd.n5698 9.3005
R17462 gnd.n5731 gnd.n5697 9.3005
R17463 gnd.n5734 gnd.n5696 9.3005
R17464 gnd.n5736 gnd.n5695 9.3005
R17465 gnd.n5737 gnd.n5694 9.3005
R17466 gnd.n5738 gnd.n5693 9.3005
R17467 gnd.n5739 gnd.n5692 9.3005
R17468 gnd.n5707 gnd.n5488 9.3005
R17469 gnd.n5756 gnd.n5479 9.3005
R17470 gnd.n5758 gnd.n5757 9.3005
R17471 gnd.n5466 gnd.n5461 9.3005
R17472 gnd.n5779 gnd.n5460 9.3005
R17473 gnd.n5782 gnd.n5781 9.3005
R17474 gnd.n5784 gnd.n5783 9.3005
R17475 gnd.n5787 gnd.n5443 9.3005
R17476 gnd.n5785 gnd.n5441 9.3005
R17477 gnd.n5807 gnd.n5439 9.3005
R17478 gnd.n5811 gnd.n5810 9.3005
R17479 gnd.n5809 gnd.n5414 9.3005
R17480 gnd.n5845 gnd.n5413 9.3005
R17481 gnd.n5848 gnd.n5847 9.3005
R17482 gnd.n5411 gnd.n5410 9.3005
R17483 gnd.n5854 gnd.n5408 9.3005
R17484 gnd.n5856 gnd.n5855 9.3005
R17485 gnd.n5382 gnd.n5381 9.3005
R17486 gnd.n5905 gnd.n5904 9.3005
R17487 gnd.n5906 gnd.n5375 9.3005
R17488 gnd.n5914 gnd.n5374 9.3005
R17489 gnd.n5917 gnd.n5916 9.3005
R17490 gnd.n5919 gnd.n5918 9.3005
R17491 gnd.n5922 gnd.n5357 9.3005
R17492 gnd.n5920 gnd.n5355 9.3005
R17493 gnd.n5942 gnd.n5353 9.3005
R17494 gnd.n5944 gnd.n5943 9.3005
R17495 gnd.n5247 gnd.n5246 9.3005
R17496 gnd.n5987 gnd.n5986 9.3005
R17497 gnd.n5988 gnd.n5240 9.3005
R17498 gnd.n5996 gnd.n5239 9.3005
R17499 gnd.n5999 gnd.n5998 9.3005
R17500 gnd.n6001 gnd.n5237 9.3005
R17501 gnd.n6005 gnd.n6004 9.3005
R17502 gnd.n6003 gnd.n5211 9.3005
R17503 gnd.n6041 gnd.n5210 9.3005
R17504 gnd.n6044 gnd.n6043 9.3005
R17505 gnd.n6046 gnd.n6045 9.3005
R17506 gnd.n6049 gnd.n5194 9.3005
R17507 gnd.n6047 gnd.n5192 9.3005
R17508 gnd.n6069 gnd.n5190 9.3005
R17509 gnd.n6071 gnd.n6070 9.3005
R17510 gnd.n5165 gnd.n5164 9.3005
R17511 gnd.n6118 gnd.n6117 9.3005
R17512 gnd.n6119 gnd.n5158 9.3005
R17513 gnd.n6127 gnd.n5157 9.3005
R17514 gnd.n6130 gnd.n6129 9.3005
R17515 gnd.n6132 gnd.n6131 9.3005
R17516 gnd.n6391 gnd.n5140 9.3005
R17517 gnd.n6133 gnd.n5138 9.3005
R17518 gnd.n6414 gnd.n5136 9.3005
R17519 gnd.n6416 gnd.n6415 9.3005
R17520 gnd.n1126 gnd.n1124 9.3005
R17521 gnd.n6571 gnd.n6570 9.3005
R17522 gnd.n5755 gnd.n5482 9.3005
R17523 gnd.n6443 gnd.n6439 9.3005
R17524 gnd.n6447 gnd.n6446 9.3005
R17525 gnd.n6448 gnd.n6438 9.3005
R17526 gnd.n6450 gnd.n6449 9.3005
R17527 gnd.n6453 gnd.n6437 9.3005
R17528 gnd.n6457 gnd.n6456 9.3005
R17529 gnd.n6458 gnd.n6436 9.3005
R17530 gnd.n6460 gnd.n6459 9.3005
R17531 gnd.n6463 gnd.n6435 9.3005
R17532 gnd.n6467 gnd.n6466 9.3005
R17533 gnd.n6468 gnd.n6434 9.3005
R17534 gnd.n6470 gnd.n6469 9.3005
R17535 gnd.n6473 gnd.n6433 9.3005
R17536 gnd.n6477 gnd.n6476 9.3005
R17537 gnd.n6478 gnd.n6432 9.3005
R17538 gnd.n6480 gnd.n6479 9.3005
R17539 gnd.n6483 gnd.n6431 9.3005
R17540 gnd.n6487 gnd.n6486 9.3005
R17541 gnd.n6488 gnd.n6430 9.3005
R17542 gnd.n6490 gnd.n6489 9.3005
R17543 gnd.n6493 gnd.n6429 9.3005
R17544 gnd.n6500 gnd.n6499 9.3005
R17545 gnd.n6501 gnd.n6428 9.3005
R17546 gnd.n6503 gnd.n6502 9.3005
R17547 gnd.n6506 gnd.n6427 9.3005
R17548 gnd.n6509 gnd.n6508 9.3005
R17549 gnd.n6441 gnd.n6440 9.3005
R17550 gnd.n5952 gnd.n5951 9.3005
R17551 gnd.n5953 gnd.n5263 9.3005
R17552 gnd.n5967 gnd.n5954 9.3005
R17553 gnd.n5966 gnd.n5955 9.3005
R17554 gnd.n5965 gnd.n5956 9.3005
R17555 gnd.n5963 gnd.n5957 9.3005
R17556 gnd.n5962 gnd.n5958 9.3005
R17557 gnd.n5960 gnd.n5959 9.3005
R17558 gnd.n5219 gnd.n5218 9.3005
R17559 gnd.n6025 gnd.n6024 9.3005
R17560 gnd.n6026 gnd.n5217 9.3005
R17561 gnd.n6033 gnd.n6027 9.3005
R17562 gnd.n6032 gnd.n6028 9.3005
R17563 gnd.n6031 gnd.n6029 9.3005
R17564 gnd.n5182 gnd.n5181 9.3005
R17565 gnd.n6079 gnd.n6078 9.3005
R17566 gnd.n6080 gnd.n5180 9.3005
R17567 gnd.n6098 gnd.n6081 9.3005
R17568 gnd.n6097 gnd.n6082 9.3005
R17569 gnd.n6096 gnd.n6083 9.3005
R17570 gnd.n6093 gnd.n6084 9.3005
R17571 gnd.n6092 gnd.n6085 9.3005
R17572 gnd.n6090 gnd.n6086 9.3005
R17573 gnd.n6089 gnd.n6087 9.3005
R17574 gnd.n5128 gnd.n5127 9.3005
R17575 gnd.n6424 gnd.n6423 9.3005
R17576 gnd.n6425 gnd.n5126 9.3005
R17577 gnd.n6512 gnd.n6426 9.3005
R17578 gnd.n6511 gnd.n6510 9.3005
R17579 gnd.n5625 gnd.n5519 9.3005
R17580 gnd.n5627 gnd.n5626 9.3005
R17581 gnd.n5509 gnd.n5508 9.3005
R17582 gnd.n5640 gnd.n5639 9.3005
R17583 gnd.n5641 gnd.n5507 9.3005
R17584 gnd.n5643 gnd.n5642 9.3005
R17585 gnd.n5496 gnd.n5495 9.3005
R17586 gnd.n5656 gnd.n5655 9.3005
R17587 gnd.n5657 gnd.n5494 9.3005
R17588 gnd.n5681 gnd.n5658 9.3005
R17589 gnd.n5680 gnd.n5659 9.3005
R17590 gnd.n5679 gnd.n5660 9.3005
R17591 gnd.n5678 gnd.n5661 9.3005
R17592 gnd.n5676 gnd.n5662 9.3005
R17593 gnd.n5675 gnd.n5663 9.3005
R17594 gnd.n5673 gnd.n5664 9.3005
R17595 gnd.n5672 gnd.n5665 9.3005
R17596 gnd.n5670 gnd.n5666 9.3005
R17597 gnd.n5669 gnd.n5667 9.3005
R17598 gnd.n5431 gnd.n5430 9.3005
R17599 gnd.n5819 gnd.n5818 9.3005
R17600 gnd.n5820 gnd.n5429 9.3005
R17601 gnd.n5824 gnd.n5821 9.3005
R17602 gnd.n5823 gnd.n5822 9.3005
R17603 gnd.n5398 gnd.n5397 9.3005
R17604 gnd.n5866 gnd.n5865 9.3005
R17605 gnd.n5867 gnd.n5396 9.3005
R17606 gnd.n5869 gnd.n5868 9.3005
R17607 gnd.n5624 gnd.n5623 9.3005
R17608 gnd.n5564 gnd.n5563 9.3005
R17609 gnd.n5569 gnd.n5561 9.3005
R17610 gnd.n5570 gnd.n5560 9.3005
R17611 gnd.n5572 gnd.n5557 9.3005
R17612 gnd.n5556 gnd.n5554 9.3005
R17613 gnd.n5578 gnd.n5553 9.3005
R17614 gnd.n5579 gnd.n5552 9.3005
R17615 gnd.n5580 gnd.n5551 9.3005
R17616 gnd.n5550 gnd.n5548 9.3005
R17617 gnd.n5586 gnd.n5547 9.3005
R17618 gnd.n5587 gnd.n5546 9.3005
R17619 gnd.n5588 gnd.n5545 9.3005
R17620 gnd.n5544 gnd.n5542 9.3005
R17621 gnd.n5594 gnd.n5541 9.3005
R17622 gnd.n5595 gnd.n5540 9.3005
R17623 gnd.n5596 gnd.n5539 9.3005
R17624 gnd.n5538 gnd.n5536 9.3005
R17625 gnd.n5602 gnd.n5535 9.3005
R17626 gnd.n5603 gnd.n5534 9.3005
R17627 gnd.n5604 gnd.n5533 9.3005
R17628 gnd.n5532 gnd.n5530 9.3005
R17629 gnd.n5609 gnd.n5529 9.3005
R17630 gnd.n5610 gnd.n5528 9.3005
R17631 gnd.n5527 gnd.n5525 9.3005
R17632 gnd.n5615 gnd.n5524 9.3005
R17633 gnd.n5617 gnd.n5616 9.3005
R17634 gnd.n5562 gnd.n5520 9.3005
R17635 gnd.n5515 gnd.n5514 9.3005
R17636 gnd.n5632 gnd.n5631 9.3005
R17637 gnd.n5633 gnd.n5513 9.3005
R17638 gnd.n5635 gnd.n5634 9.3005
R17639 gnd.n5503 gnd.n5502 9.3005
R17640 gnd.n5648 gnd.n5647 9.3005
R17641 gnd.n5649 gnd.n5501 9.3005
R17642 gnd.n5651 gnd.n5650 9.3005
R17643 gnd.n5490 gnd.n5489 9.3005
R17644 gnd.n5746 gnd.n5745 9.3005
R17645 gnd.n5748 gnd.n5487 9.3005
R17646 gnd.n5750 gnd.n5749 9.3005
R17647 gnd.n5481 gnd.n5478 9.3005
R17648 gnd.n5760 gnd.n5759 9.3005
R17649 gnd.n5480 gnd.n5462 9.3005
R17650 gnd.n5778 gnd.n5777 9.3005
R17651 gnd.n5780 gnd.n5458 9.3005
R17652 gnd.n5790 gnd.n5459 9.3005
R17653 gnd.n5789 gnd.n5788 9.3005
R17654 gnd.n5786 gnd.n5437 9.3005
R17655 gnd.n5814 gnd.n5438 9.3005
R17656 gnd.n5813 gnd.n5812 9.3005
R17657 gnd.n5440 gnd.n5415 9.3005
R17658 gnd.n5844 gnd.n5843 9.3005
R17659 gnd.n5846 gnd.n5405 9.3005
R17660 gnd.n5861 gnd.n5406 9.3005
R17661 gnd.n5860 gnd.n5407 9.3005
R17662 gnd.n5859 gnd.n5857 9.3005
R17663 gnd.n5409 gnd.n5383 9.3005
R17664 gnd.n5902 gnd.n5901 9.3005
R17665 gnd.n5903 gnd.n5376 9.3005
R17666 gnd.n5913 gnd.n5912 9.3005
R17667 gnd.n5915 gnd.n5372 9.3005
R17668 gnd.n5925 gnd.n5373 9.3005
R17669 gnd.n5924 gnd.n5923 9.3005
R17670 gnd.n5921 gnd.n5351 9.3005
R17671 gnd.n5947 gnd.n5352 9.3005
R17672 gnd.n5946 gnd.n5945 9.3005
R17673 gnd.n5354 gnd.n5248 9.3005
R17674 gnd.n5984 gnd.n5983 9.3005
R17675 gnd.n5985 gnd.n5241 9.3005
R17676 gnd.n5995 gnd.n5994 9.3005
R17677 gnd.n5997 gnd.n5235 9.3005
R17678 gnd.n6008 gnd.n5236 9.3005
R17679 gnd.n6007 gnd.n6006 9.3005
R17680 gnd.n5238 gnd.n5212 9.3005
R17681 gnd.n6040 gnd.n6039 9.3005
R17682 gnd.n6042 gnd.n5208 9.3005
R17683 gnd.n6052 gnd.n5209 9.3005
R17684 gnd.n6051 gnd.n6050 9.3005
R17685 gnd.n6048 gnd.n5188 9.3005
R17686 gnd.n6074 gnd.n5189 9.3005
R17687 gnd.n6073 gnd.n6072 9.3005
R17688 gnd.n5191 gnd.n5166 9.3005
R17689 gnd.n6115 gnd.n6114 9.3005
R17690 gnd.n6116 gnd.n5159 9.3005
R17691 gnd.n6126 gnd.n6125 9.3005
R17692 gnd.n6128 gnd.n5155 9.3005
R17693 gnd.n6394 gnd.n5156 9.3005
R17694 gnd.n6393 gnd.n6392 9.3005
R17695 gnd.n6134 gnd.n5134 9.3005
R17696 gnd.n6419 gnd.n5135 9.3005
R17697 gnd.n6418 gnd.n6417 9.3005
R17698 gnd.n5137 gnd.n1123 9.3005
R17699 gnd.n6573 gnd.n6572 9.3005
R17700 gnd.n5619 gnd.n5618 9.3005
R17701 gnd.n949 gnd.n948 9.3005
R17702 gnd.n6749 gnd.n6748 9.3005
R17703 gnd.n6750 gnd.n947 9.3005
R17704 gnd.n6752 gnd.n6751 9.3005
R17705 gnd.n943 gnd.n942 9.3005
R17706 gnd.n6759 gnd.n6758 9.3005
R17707 gnd.n6760 gnd.n941 9.3005
R17708 gnd.n6762 gnd.n6761 9.3005
R17709 gnd.n937 gnd.n936 9.3005
R17710 gnd.n6769 gnd.n6768 9.3005
R17711 gnd.n6770 gnd.n935 9.3005
R17712 gnd.n6772 gnd.n6771 9.3005
R17713 gnd.n931 gnd.n930 9.3005
R17714 gnd.n6779 gnd.n6778 9.3005
R17715 gnd.n6780 gnd.n929 9.3005
R17716 gnd.n6782 gnd.n6781 9.3005
R17717 gnd.n925 gnd.n924 9.3005
R17718 gnd.n6789 gnd.n6788 9.3005
R17719 gnd.n6790 gnd.n923 9.3005
R17720 gnd.n6792 gnd.n6791 9.3005
R17721 gnd.n919 gnd.n918 9.3005
R17722 gnd.n6799 gnd.n6798 9.3005
R17723 gnd.n6800 gnd.n917 9.3005
R17724 gnd.n6802 gnd.n6801 9.3005
R17725 gnd.n913 gnd.n912 9.3005
R17726 gnd.n6809 gnd.n6808 9.3005
R17727 gnd.n6810 gnd.n911 9.3005
R17728 gnd.n6812 gnd.n6811 9.3005
R17729 gnd.n907 gnd.n906 9.3005
R17730 gnd.n6819 gnd.n6818 9.3005
R17731 gnd.n6820 gnd.n905 9.3005
R17732 gnd.n6822 gnd.n6821 9.3005
R17733 gnd.n901 gnd.n900 9.3005
R17734 gnd.n6829 gnd.n6828 9.3005
R17735 gnd.n6830 gnd.n899 9.3005
R17736 gnd.n6832 gnd.n6831 9.3005
R17737 gnd.n895 gnd.n894 9.3005
R17738 gnd.n6839 gnd.n6838 9.3005
R17739 gnd.n6840 gnd.n893 9.3005
R17740 gnd.n6842 gnd.n6841 9.3005
R17741 gnd.n889 gnd.n888 9.3005
R17742 gnd.n6849 gnd.n6848 9.3005
R17743 gnd.n6850 gnd.n887 9.3005
R17744 gnd.n6852 gnd.n6851 9.3005
R17745 gnd.n883 gnd.n882 9.3005
R17746 gnd.n6859 gnd.n6858 9.3005
R17747 gnd.n6860 gnd.n881 9.3005
R17748 gnd.n6862 gnd.n6861 9.3005
R17749 gnd.n877 gnd.n876 9.3005
R17750 gnd.n6869 gnd.n6868 9.3005
R17751 gnd.n6870 gnd.n875 9.3005
R17752 gnd.n6872 gnd.n6871 9.3005
R17753 gnd.n871 gnd.n870 9.3005
R17754 gnd.n6879 gnd.n6878 9.3005
R17755 gnd.n6880 gnd.n869 9.3005
R17756 gnd.n6882 gnd.n6881 9.3005
R17757 gnd.n865 gnd.n864 9.3005
R17758 gnd.n6889 gnd.n6888 9.3005
R17759 gnd.n6890 gnd.n863 9.3005
R17760 gnd.n6892 gnd.n6891 9.3005
R17761 gnd.n859 gnd.n858 9.3005
R17762 gnd.n6899 gnd.n6898 9.3005
R17763 gnd.n6900 gnd.n857 9.3005
R17764 gnd.n6902 gnd.n6901 9.3005
R17765 gnd.n853 gnd.n852 9.3005
R17766 gnd.n6909 gnd.n6908 9.3005
R17767 gnd.n6910 gnd.n851 9.3005
R17768 gnd.n6912 gnd.n6911 9.3005
R17769 gnd.n847 gnd.n846 9.3005
R17770 gnd.n6919 gnd.n6918 9.3005
R17771 gnd.n6920 gnd.n845 9.3005
R17772 gnd.n6922 gnd.n6921 9.3005
R17773 gnd.n841 gnd.n840 9.3005
R17774 gnd.n6929 gnd.n6928 9.3005
R17775 gnd.n6930 gnd.n839 9.3005
R17776 gnd.n6932 gnd.n6931 9.3005
R17777 gnd.n835 gnd.n834 9.3005
R17778 gnd.n6939 gnd.n6938 9.3005
R17779 gnd.n6940 gnd.n833 9.3005
R17780 gnd.n6942 gnd.n6941 9.3005
R17781 gnd.n829 gnd.n828 9.3005
R17782 gnd.n6949 gnd.n6948 9.3005
R17783 gnd.n6950 gnd.n827 9.3005
R17784 gnd.n6952 gnd.n6951 9.3005
R17785 gnd.n823 gnd.n822 9.3005
R17786 gnd.n6959 gnd.n6958 9.3005
R17787 gnd.n6960 gnd.n821 9.3005
R17788 gnd.n6962 gnd.n6961 9.3005
R17789 gnd.n817 gnd.n816 9.3005
R17790 gnd.n6969 gnd.n6968 9.3005
R17791 gnd.n6970 gnd.n815 9.3005
R17792 gnd.n6972 gnd.n6971 9.3005
R17793 gnd.n811 gnd.n810 9.3005
R17794 gnd.n6979 gnd.n6978 9.3005
R17795 gnd.n6980 gnd.n809 9.3005
R17796 gnd.n6982 gnd.n6981 9.3005
R17797 gnd.n805 gnd.n804 9.3005
R17798 gnd.n6989 gnd.n6988 9.3005
R17799 gnd.n6990 gnd.n803 9.3005
R17800 gnd.n6992 gnd.n6991 9.3005
R17801 gnd.n799 gnd.n798 9.3005
R17802 gnd.n6999 gnd.n6998 9.3005
R17803 gnd.n7000 gnd.n797 9.3005
R17804 gnd.n7002 gnd.n7001 9.3005
R17805 gnd.n793 gnd.n792 9.3005
R17806 gnd.n7009 gnd.n7008 9.3005
R17807 gnd.n7010 gnd.n791 9.3005
R17808 gnd.n7012 gnd.n7011 9.3005
R17809 gnd.n787 gnd.n786 9.3005
R17810 gnd.n7019 gnd.n7018 9.3005
R17811 gnd.n7020 gnd.n785 9.3005
R17812 gnd.n7022 gnd.n7021 9.3005
R17813 gnd.n781 gnd.n780 9.3005
R17814 gnd.n7029 gnd.n7028 9.3005
R17815 gnd.n7030 gnd.n779 9.3005
R17816 gnd.n7032 gnd.n7031 9.3005
R17817 gnd.n775 gnd.n774 9.3005
R17818 gnd.n7039 gnd.n7038 9.3005
R17819 gnd.n7040 gnd.n773 9.3005
R17820 gnd.n7042 gnd.n7041 9.3005
R17821 gnd.n769 gnd.n768 9.3005
R17822 gnd.n7049 gnd.n7048 9.3005
R17823 gnd.n7050 gnd.n767 9.3005
R17824 gnd.n7052 gnd.n7051 9.3005
R17825 gnd.n763 gnd.n762 9.3005
R17826 gnd.n7059 gnd.n7058 9.3005
R17827 gnd.n7060 gnd.n761 9.3005
R17828 gnd.n7062 gnd.n7061 9.3005
R17829 gnd.n757 gnd.n756 9.3005
R17830 gnd.n7069 gnd.n7068 9.3005
R17831 gnd.n7070 gnd.n755 9.3005
R17832 gnd.n7072 gnd.n7071 9.3005
R17833 gnd.n751 gnd.n750 9.3005
R17834 gnd.n7079 gnd.n7078 9.3005
R17835 gnd.n7080 gnd.n749 9.3005
R17836 gnd.n7082 gnd.n7081 9.3005
R17837 gnd.n745 gnd.n744 9.3005
R17838 gnd.n7089 gnd.n7088 9.3005
R17839 gnd.n7090 gnd.n743 9.3005
R17840 gnd.n7092 gnd.n7091 9.3005
R17841 gnd.n739 gnd.n738 9.3005
R17842 gnd.n7099 gnd.n7098 9.3005
R17843 gnd.n7100 gnd.n737 9.3005
R17844 gnd.n7102 gnd.n7101 9.3005
R17845 gnd.n733 gnd.n732 9.3005
R17846 gnd.n7109 gnd.n7108 9.3005
R17847 gnd.n7110 gnd.n731 9.3005
R17848 gnd.n7112 gnd.n7111 9.3005
R17849 gnd.n727 gnd.n726 9.3005
R17850 gnd.n7119 gnd.n7118 9.3005
R17851 gnd.n7120 gnd.n725 9.3005
R17852 gnd.n7123 gnd.n7122 9.3005
R17853 gnd.n7121 gnd.n721 9.3005
R17854 gnd.n7129 gnd.n720 9.3005
R17855 gnd.n7131 gnd.n7130 9.3005
R17856 gnd.n716 gnd.n715 9.3005
R17857 gnd.n7140 gnd.n7139 9.3005
R17858 gnd.n7141 gnd.n714 9.3005
R17859 gnd.n7143 gnd.n7142 9.3005
R17860 gnd.n710 gnd.n709 9.3005
R17861 gnd.n7150 gnd.n7149 9.3005
R17862 gnd.n7151 gnd.n708 9.3005
R17863 gnd.n7153 gnd.n7152 9.3005
R17864 gnd.n704 gnd.n703 9.3005
R17865 gnd.n7160 gnd.n7159 9.3005
R17866 gnd.n7161 gnd.n702 9.3005
R17867 gnd.n7163 gnd.n7162 9.3005
R17868 gnd.n698 gnd.n697 9.3005
R17869 gnd.n7170 gnd.n7169 9.3005
R17870 gnd.n7171 gnd.n696 9.3005
R17871 gnd.n7173 gnd.n7172 9.3005
R17872 gnd.n692 gnd.n691 9.3005
R17873 gnd.n7180 gnd.n7179 9.3005
R17874 gnd.n7181 gnd.n690 9.3005
R17875 gnd.n7183 gnd.n7182 9.3005
R17876 gnd.n686 gnd.n685 9.3005
R17877 gnd.n7190 gnd.n7189 9.3005
R17878 gnd.n7191 gnd.n684 9.3005
R17879 gnd.n7193 gnd.n7192 9.3005
R17880 gnd.n680 gnd.n679 9.3005
R17881 gnd.n7200 gnd.n7199 9.3005
R17882 gnd.n7201 gnd.n678 9.3005
R17883 gnd.n7203 gnd.n7202 9.3005
R17884 gnd.n674 gnd.n673 9.3005
R17885 gnd.n7210 gnd.n7209 9.3005
R17886 gnd.n7211 gnd.n672 9.3005
R17887 gnd.n7213 gnd.n7212 9.3005
R17888 gnd.n668 gnd.n667 9.3005
R17889 gnd.n7220 gnd.n7219 9.3005
R17890 gnd.n7221 gnd.n666 9.3005
R17891 gnd.n7223 gnd.n7222 9.3005
R17892 gnd.n662 gnd.n661 9.3005
R17893 gnd.n7230 gnd.n7229 9.3005
R17894 gnd.n7231 gnd.n660 9.3005
R17895 gnd.n7233 gnd.n7232 9.3005
R17896 gnd.n656 gnd.n655 9.3005
R17897 gnd.n7240 gnd.n7239 9.3005
R17898 gnd.n7241 gnd.n654 9.3005
R17899 gnd.n7243 gnd.n7242 9.3005
R17900 gnd.n650 gnd.n649 9.3005
R17901 gnd.n7250 gnd.n7249 9.3005
R17902 gnd.n7251 gnd.n648 9.3005
R17903 gnd.n7253 gnd.n7252 9.3005
R17904 gnd.n644 gnd.n643 9.3005
R17905 gnd.n7260 gnd.n7259 9.3005
R17906 gnd.n7261 gnd.n642 9.3005
R17907 gnd.n7263 gnd.n7262 9.3005
R17908 gnd.n638 gnd.n637 9.3005
R17909 gnd.n7270 gnd.n7269 9.3005
R17910 gnd.n7271 gnd.n636 9.3005
R17911 gnd.n7273 gnd.n7272 9.3005
R17912 gnd.n632 gnd.n631 9.3005
R17913 gnd.n7280 gnd.n7279 9.3005
R17914 gnd.n7281 gnd.n630 9.3005
R17915 gnd.n7283 gnd.n7282 9.3005
R17916 gnd.n626 gnd.n625 9.3005
R17917 gnd.n7290 gnd.n7289 9.3005
R17918 gnd.n7291 gnd.n624 9.3005
R17919 gnd.n7293 gnd.n7292 9.3005
R17920 gnd.n620 gnd.n619 9.3005
R17921 gnd.n7300 gnd.n7299 9.3005
R17922 gnd.n7301 gnd.n618 9.3005
R17923 gnd.n7303 gnd.n7302 9.3005
R17924 gnd.n614 gnd.n613 9.3005
R17925 gnd.n7310 gnd.n7309 9.3005
R17926 gnd.n7311 gnd.n612 9.3005
R17927 gnd.n7313 gnd.n7312 9.3005
R17928 gnd.n608 gnd.n607 9.3005
R17929 gnd.n7320 gnd.n7319 9.3005
R17930 gnd.n7321 gnd.n606 9.3005
R17931 gnd.n7323 gnd.n7322 9.3005
R17932 gnd.n602 gnd.n601 9.3005
R17933 gnd.n7330 gnd.n7329 9.3005
R17934 gnd.n7331 gnd.n600 9.3005
R17935 gnd.n7333 gnd.n7332 9.3005
R17936 gnd.n596 gnd.n595 9.3005
R17937 gnd.n7342 gnd.n7341 9.3005
R17938 gnd.n7343 gnd.n594 9.3005
R17939 gnd.n7346 gnd.n7345 9.3005
R17940 gnd.n7133 gnd.n7132 9.3005
R17941 gnd.n7761 gnd.n7760 9.3005
R17942 gnd.n7759 gnd.n97 9.3005
R17943 gnd.n382 gnd.n99 9.3005
R17944 gnd.n385 gnd.n384 9.3005
R17945 gnd.n386 gnd.n381 9.3005
R17946 gnd.n389 gnd.n387 9.3005
R17947 gnd.n390 gnd.n380 9.3005
R17948 gnd.n393 gnd.n392 9.3005
R17949 gnd.n394 gnd.n379 9.3005
R17950 gnd.n397 gnd.n395 9.3005
R17951 gnd.n398 gnd.n378 9.3005
R17952 gnd.n401 gnd.n400 9.3005
R17953 gnd.n402 gnd.n377 9.3005
R17954 gnd.n405 gnd.n403 9.3005
R17955 gnd.n406 gnd.n376 9.3005
R17956 gnd.n409 gnd.n408 9.3005
R17957 gnd.n410 gnd.n375 9.3005
R17958 gnd.n413 gnd.n411 9.3005
R17959 gnd.n414 gnd.n374 9.3005
R17960 gnd.n417 gnd.n416 9.3005
R17961 gnd.n418 gnd.n373 9.3005
R17962 gnd.n421 gnd.n419 9.3005
R17963 gnd.n422 gnd.n372 9.3005
R17964 gnd.n425 gnd.n424 9.3005
R17965 gnd.n426 gnd.n371 9.3005
R17966 gnd.n429 gnd.n427 9.3005
R17967 gnd.n430 gnd.n370 9.3005
R17968 gnd.n433 gnd.n432 9.3005
R17969 gnd.n434 gnd.n369 9.3005
R17970 gnd.n437 gnd.n435 9.3005
R17971 gnd.n438 gnd.n368 9.3005
R17972 gnd.n442 gnd.n441 9.3005
R17973 gnd.n477 gnd.n348 9.3005
R17974 gnd.n476 gnd.n350 9.3005
R17975 gnd.n473 gnd.n351 9.3005
R17976 gnd.n472 gnd.n352 9.3005
R17977 gnd.n469 gnd.n353 9.3005
R17978 gnd.n468 gnd.n354 9.3005
R17979 gnd.n465 gnd.n355 9.3005
R17980 gnd.n464 gnd.n356 9.3005
R17981 gnd.n461 gnd.n357 9.3005
R17982 gnd.n460 gnd.n358 9.3005
R17983 gnd.n457 gnd.n359 9.3005
R17984 gnd.n456 gnd.n360 9.3005
R17985 gnd.n453 gnd.n361 9.3005
R17986 gnd.n452 gnd.n362 9.3005
R17987 gnd.n449 gnd.n363 9.3005
R17988 gnd.n448 gnd.n364 9.3005
R17989 gnd.n445 gnd.n444 9.3005
R17990 gnd.n443 gnd.n365 9.3005
R17991 gnd.n479 gnd.n478 9.3005
R17992 gnd.n249 gnd.n248 9.3005
R17993 gnd.n7660 gnd.n290 9.3005
R17994 gnd.n7659 gnd.n291 9.3005
R17995 gnd.n7658 gnd.n292 9.3005
R17996 gnd.n7655 gnd.n293 9.3005
R17997 gnd.n7654 gnd.n294 9.3005
R17998 gnd.n7651 gnd.n295 9.3005
R17999 gnd.n7650 gnd.n296 9.3005
R18000 gnd.n7647 gnd.n297 9.3005
R18001 gnd.n7646 gnd.n298 9.3005
R18002 gnd.n7643 gnd.n299 9.3005
R18003 gnd.n7642 gnd.n300 9.3005
R18004 gnd.n7639 gnd.n301 9.3005
R18005 gnd.n7638 gnd.n302 9.3005
R18006 gnd.n7635 gnd.n303 9.3005
R18007 gnd.n7634 gnd.n304 9.3005
R18008 gnd.n7631 gnd.n305 9.3005
R18009 gnd.n7627 gnd.n306 9.3005
R18010 gnd.n7624 gnd.n307 9.3005
R18011 gnd.n7623 gnd.n308 9.3005
R18012 gnd.n7620 gnd.n309 9.3005
R18013 gnd.n7619 gnd.n310 9.3005
R18014 gnd.n7616 gnd.n311 9.3005
R18015 gnd.n7615 gnd.n312 9.3005
R18016 gnd.n7612 gnd.n313 9.3005
R18017 gnd.n7611 gnd.n314 9.3005
R18018 gnd.n7608 gnd.n315 9.3005
R18019 gnd.n7607 gnd.n316 9.3005
R18020 gnd.n7604 gnd.n317 9.3005
R18021 gnd.n7603 gnd.n318 9.3005
R18022 gnd.n7600 gnd.n319 9.3005
R18023 gnd.n7599 gnd.n320 9.3005
R18024 gnd.n7596 gnd.n321 9.3005
R18025 gnd.n7595 gnd.n322 9.3005
R18026 gnd.n7592 gnd.n323 9.3005
R18027 gnd.n7591 gnd.n324 9.3005
R18028 gnd.n7588 gnd.n7587 9.3005
R18029 gnd.n7586 gnd.n325 9.3005
R18030 gnd.n7585 gnd.n7584 9.3005
R18031 gnd.n7581 gnd.n328 9.3005
R18032 gnd.n7578 gnd.n329 9.3005
R18033 gnd.n7577 gnd.n330 9.3005
R18034 gnd.n7574 gnd.n331 9.3005
R18035 gnd.n7573 gnd.n332 9.3005
R18036 gnd.n7570 gnd.n333 9.3005
R18037 gnd.n7569 gnd.n334 9.3005
R18038 gnd.n7566 gnd.n335 9.3005
R18039 gnd.n7565 gnd.n336 9.3005
R18040 gnd.n7562 gnd.n337 9.3005
R18041 gnd.n7561 gnd.n338 9.3005
R18042 gnd.n7558 gnd.n339 9.3005
R18043 gnd.n7557 gnd.n340 9.3005
R18044 gnd.n7554 gnd.n341 9.3005
R18045 gnd.n7553 gnd.n342 9.3005
R18046 gnd.n7550 gnd.n343 9.3005
R18047 gnd.n7549 gnd.n344 9.3005
R18048 gnd.n7546 gnd.n7545 9.3005
R18049 gnd.n7544 gnd.n345 9.3005
R18050 gnd.n7666 gnd.n7665 9.3005
R18051 gnd.n4377 gnd.n4376 9.3005
R18052 gnd.n1978 gnd.n1977 9.3005
R18053 gnd.n2002 gnd.n2001 9.3005
R18054 gnd.n4364 gnd.n2003 9.3005
R18055 gnd.n4363 gnd.n2004 9.3005
R18056 gnd.n4362 gnd.n2005 9.3005
R18057 gnd.n4274 gnd.n2006 9.3005
R18058 gnd.n4352 gnd.n2024 9.3005
R18059 gnd.n4351 gnd.n2025 9.3005
R18060 gnd.n4350 gnd.n2026 9.3005
R18061 gnd.n4289 gnd.n2027 9.3005
R18062 gnd.n4340 gnd.n2044 9.3005
R18063 gnd.n4339 gnd.n2045 9.3005
R18064 gnd.n4338 gnd.n2046 9.3005
R18065 gnd.n4290 gnd.n2047 9.3005
R18066 gnd.n4291 gnd.n570 9.3005
R18067 gnd.n7381 gnd.n571 9.3005
R18068 gnd.n7380 gnd.n572 9.3005
R18069 gnd.n7379 gnd.n7374 9.3005
R18070 gnd.n7378 gnd.n7375 9.3005
R18071 gnd.n546 gnd.n542 9.3005
R18072 gnd.n7417 gnd.n543 9.3005
R18073 gnd.n7416 gnd.n544 9.3005
R18074 gnd.n7415 gnd.n7410 9.3005
R18075 gnd.n7414 gnd.n7411 9.3005
R18076 gnd.n518 gnd.n512 9.3005
R18077 gnd.n7450 gnd.n513 9.3005
R18078 gnd.n7449 gnd.n514 9.3005
R18079 gnd.n7448 gnd.n515 9.3005
R18080 gnd.n489 gnd.n488 9.3005
R18081 gnd.n7476 gnd.n7475 9.3005
R18082 gnd.n7477 gnd.n482 9.3005
R18083 gnd.n7484 gnd.n483 9.3005
R18084 gnd.n7485 gnd.n481 9.3005
R18085 gnd.n7488 gnd.n7487 9.3005
R18086 gnd.n7489 gnd.n123 9.3005
R18087 gnd.n7747 gnd.n124 9.3005
R18088 gnd.n7746 gnd.n125 9.3005
R18089 gnd.n7745 gnd.n126 9.3005
R18090 gnd.n7497 gnd.n127 9.3005
R18091 gnd.n7735 gnd.n141 9.3005
R18092 gnd.n7734 gnd.n142 9.3005
R18093 gnd.n7733 gnd.n143 9.3005
R18094 gnd.n7504 gnd.n144 9.3005
R18095 gnd.n7723 gnd.n161 9.3005
R18096 gnd.n7722 gnd.n162 9.3005
R18097 gnd.n7721 gnd.n163 9.3005
R18098 gnd.n7511 gnd.n164 9.3005
R18099 gnd.n7711 gnd.n179 9.3005
R18100 gnd.n7710 gnd.n180 9.3005
R18101 gnd.n7709 gnd.n181 9.3005
R18102 gnd.n7518 gnd.n182 9.3005
R18103 gnd.n7699 gnd.n199 9.3005
R18104 gnd.n7698 gnd.n200 9.3005
R18105 gnd.n7697 gnd.n201 9.3005
R18106 gnd.n7525 gnd.n202 9.3005
R18107 gnd.n7687 gnd.n217 9.3005
R18108 gnd.n7686 gnd.n218 9.3005
R18109 gnd.n7685 gnd.n219 9.3005
R18110 gnd.n7532 gnd.n220 9.3005
R18111 gnd.n7675 gnd.n237 9.3005
R18112 gnd.n7674 gnd.n238 9.3005
R18113 gnd.n7673 gnd.n239 9.3005
R18114 gnd.n7542 gnd.n240 9.3005
R18115 gnd.n4378 gnd.n1976 9.3005
R18116 gnd.n4376 gnd.n4375 9.3005
R18117 gnd.n4374 gnd.n1978 9.3005
R18118 gnd.n2002 gnd.n1979 9.3005
R18119 gnd.n2070 gnd.n2003 9.3005
R18120 gnd.n4272 gnd.n2004 9.3005
R18121 gnd.n4273 gnd.n2005 9.3005
R18122 gnd.n4275 gnd.n4274 9.3005
R18123 gnd.n2066 gnd.n2024 9.3005
R18124 gnd.n4287 gnd.n2025 9.3005
R18125 gnd.n4288 gnd.n2026 9.3005
R18126 gnd.n4298 gnd.n4289 9.3005
R18127 gnd.n4297 gnd.n2044 9.3005
R18128 gnd.n4296 gnd.n2045 9.3005
R18129 gnd.n4295 gnd.n2046 9.3005
R18130 gnd.n4294 gnd.n4290 9.3005
R18131 gnd.n4293 gnd.n4291 9.3005
R18132 gnd.n573 gnd.n571 9.3005
R18133 gnd.n7372 gnd.n572 9.3005
R18134 gnd.n7374 gnd.n7373 9.3005
R18135 gnd.n7375 gnd.n545 9.3005
R18136 gnd.n7404 gnd.n546 9.3005
R18137 gnd.n7405 gnd.n543 9.3005
R18138 gnd.n7408 gnd.n544 9.3005
R18139 gnd.n7410 gnd.n7409 9.3005
R18140 gnd.n7411 gnd.n517 9.3005
R18141 gnd.n7440 gnd.n518 9.3005
R18142 gnd.n7441 gnd.n513 9.3005
R18143 gnd.n7442 gnd.n514 9.3005
R18144 gnd.n7444 gnd.n515 9.3005
R18145 gnd.n7443 gnd.n488 9.3005
R18146 gnd.n7476 gnd.n487 9.3005
R18147 gnd.n7478 gnd.n7477 9.3005
R18148 gnd.n7480 gnd.n483 9.3005
R18149 gnd.n7479 gnd.n481 9.3005
R18150 gnd.n7488 gnd.n480 9.3005
R18151 gnd.n7492 gnd.n7489 9.3005
R18152 gnd.n7493 gnd.n124 9.3005
R18153 gnd.n7495 gnd.n125 9.3005
R18154 gnd.n7496 gnd.n126 9.3005
R18155 gnd.n7499 gnd.n7497 9.3005
R18156 gnd.n7500 gnd.n141 9.3005
R18157 gnd.n7502 gnd.n142 9.3005
R18158 gnd.n7503 gnd.n143 9.3005
R18159 gnd.n7506 gnd.n7504 9.3005
R18160 gnd.n7507 gnd.n161 9.3005
R18161 gnd.n7509 gnd.n162 9.3005
R18162 gnd.n7510 gnd.n163 9.3005
R18163 gnd.n7513 gnd.n7511 9.3005
R18164 gnd.n7514 gnd.n179 9.3005
R18165 gnd.n7516 gnd.n180 9.3005
R18166 gnd.n7517 gnd.n181 9.3005
R18167 gnd.n7520 gnd.n7518 9.3005
R18168 gnd.n7521 gnd.n199 9.3005
R18169 gnd.n7523 gnd.n200 9.3005
R18170 gnd.n7524 gnd.n201 9.3005
R18171 gnd.n7527 gnd.n7525 9.3005
R18172 gnd.n7528 gnd.n217 9.3005
R18173 gnd.n7530 gnd.n218 9.3005
R18174 gnd.n7531 gnd.n219 9.3005
R18175 gnd.n7534 gnd.n7532 9.3005
R18176 gnd.n7535 gnd.n237 9.3005
R18177 gnd.n7537 gnd.n238 9.3005
R18178 gnd.n7538 gnd.n239 9.3005
R18179 gnd.n7542 gnd.n7541 9.3005
R18180 gnd.n1976 gnd.n1970 9.3005
R18181 gnd.n4388 gnd.n4387 9.3005
R18182 gnd.n4391 gnd.n1968 9.3005
R18183 gnd.n4392 gnd.n1967 9.3005
R18184 gnd.n4395 gnd.n1966 9.3005
R18185 gnd.n4396 gnd.n1965 9.3005
R18186 gnd.n4399 gnd.n1964 9.3005
R18187 gnd.n4400 gnd.n1963 9.3005
R18188 gnd.n4403 gnd.n1962 9.3005
R18189 gnd.n4404 gnd.n1961 9.3005
R18190 gnd.n4407 gnd.n1960 9.3005
R18191 gnd.n4408 gnd.n1959 9.3005
R18192 gnd.n4411 gnd.n1958 9.3005
R18193 gnd.n4412 gnd.n1957 9.3005
R18194 gnd.n4415 gnd.n1956 9.3005
R18195 gnd.n4416 gnd.n1955 9.3005
R18196 gnd.n4419 gnd.n1954 9.3005
R18197 gnd.n4420 gnd.n1953 9.3005
R18198 gnd.n4423 gnd.n1952 9.3005
R18199 gnd.n4424 gnd.n1951 9.3005
R18200 gnd.n4427 gnd.n1950 9.3005
R18201 gnd.n4431 gnd.n1946 9.3005
R18202 gnd.n4432 gnd.n1945 9.3005
R18203 gnd.n4435 gnd.n1944 9.3005
R18204 gnd.n4436 gnd.n1943 9.3005
R18205 gnd.n4439 gnd.n1942 9.3005
R18206 gnd.n4440 gnd.n1941 9.3005
R18207 gnd.n4443 gnd.n1940 9.3005
R18208 gnd.n4444 gnd.n1939 9.3005
R18209 gnd.n4447 gnd.n1938 9.3005
R18210 gnd.n4449 gnd.n1934 9.3005
R18211 gnd.n4452 gnd.n1933 9.3005
R18212 gnd.n4453 gnd.n1932 9.3005
R18213 gnd.n4456 gnd.n1931 9.3005
R18214 gnd.n4457 gnd.n1930 9.3005
R18215 gnd.n4460 gnd.n1929 9.3005
R18216 gnd.n4461 gnd.n1928 9.3005
R18217 gnd.n4464 gnd.n1927 9.3005
R18218 gnd.n4466 gnd.n1924 9.3005
R18219 gnd.n4469 gnd.n1923 9.3005
R18220 gnd.n4470 gnd.n1922 9.3005
R18221 gnd.n4473 gnd.n1921 9.3005
R18222 gnd.n4474 gnd.n1920 9.3005
R18223 gnd.n4477 gnd.n1919 9.3005
R18224 gnd.n4478 gnd.n1918 9.3005
R18225 gnd.n4481 gnd.n1917 9.3005
R18226 gnd.n4482 gnd.n1916 9.3005
R18227 gnd.n4485 gnd.n1915 9.3005
R18228 gnd.n4486 gnd.n1914 9.3005
R18229 gnd.n4489 gnd.n1913 9.3005
R18230 gnd.n4490 gnd.n1912 9.3005
R18231 gnd.n4493 gnd.n1911 9.3005
R18232 gnd.n4495 gnd.n1910 9.3005
R18233 gnd.n4496 gnd.n1909 9.3005
R18234 gnd.n4497 gnd.n1908 9.3005
R18235 gnd.n4498 gnd.n1907 9.3005
R18236 gnd.n4428 gnd.n1947 9.3005
R18237 gnd.n4386 gnd.n4383 9.3005
R18238 gnd.n1989 gnd.n1986 9.3005
R18239 gnd.n4370 gnd.n1990 9.3005
R18240 gnd.n4369 gnd.n1991 9.3005
R18241 gnd.n4368 gnd.n1992 9.3005
R18242 gnd.n2013 gnd.n1993 9.3005
R18243 gnd.n4358 gnd.n2014 9.3005
R18244 gnd.n4357 gnd.n2015 9.3005
R18245 gnd.n4356 gnd.n2016 9.3005
R18246 gnd.n2034 gnd.n2017 9.3005
R18247 gnd.n4346 gnd.n2035 9.3005
R18248 gnd.n4345 gnd.n2036 9.3005
R18249 gnd.n4344 gnd.n2037 9.3005
R18250 gnd.n4330 gnd.n2038 9.3005
R18251 gnd.n4334 gnd.n4331 9.3005
R18252 gnd.n4333 gnd.n4332 9.3005
R18253 gnd.n563 gnd.n562 9.3005
R18254 gnd.n7386 gnd.n7385 9.3005
R18255 gnd.n7387 gnd.n561 9.3005
R18256 gnd.n7391 gnd.n7388 9.3005
R18257 gnd.n7390 gnd.n7389 9.3005
R18258 gnd.n534 gnd.n533 9.3005
R18259 gnd.n7422 gnd.n7421 9.3005
R18260 gnd.n7423 gnd.n532 9.3005
R18261 gnd.n7428 gnd.n7424 9.3005
R18262 gnd.n7427 gnd.n7425 9.3005
R18263 gnd.n7426 gnd.n109 9.3005
R18264 gnd.n114 gnd.n108 9.3005
R18265 gnd.n7741 gnd.n133 9.3005
R18266 gnd.n7740 gnd.n134 9.3005
R18267 gnd.n7739 gnd.n135 9.3005
R18268 gnd.n150 gnd.n136 9.3005
R18269 gnd.n7729 gnd.n151 9.3005
R18270 gnd.n7728 gnd.n152 9.3005
R18271 gnd.n7727 gnd.n153 9.3005
R18272 gnd.n170 gnd.n154 9.3005
R18273 gnd.n7717 gnd.n171 9.3005
R18274 gnd.n7716 gnd.n172 9.3005
R18275 gnd.n7715 gnd.n173 9.3005
R18276 gnd.n188 gnd.n174 9.3005
R18277 gnd.n7705 gnd.n189 9.3005
R18278 gnd.n7704 gnd.n190 9.3005
R18279 gnd.n7703 gnd.n191 9.3005
R18280 gnd.n208 gnd.n192 9.3005
R18281 gnd.n7693 gnd.n209 9.3005
R18282 gnd.n7692 gnd.n210 9.3005
R18283 gnd.n7691 gnd.n211 9.3005
R18284 gnd.n227 gnd.n212 9.3005
R18285 gnd.n7681 gnd.n228 9.3005
R18286 gnd.n7680 gnd.n229 9.3005
R18287 gnd.n7679 gnd.n230 9.3005
R18288 gnd.n246 gnd.n231 9.3005
R18289 gnd.n7669 gnd.n247 9.3005
R18290 gnd.n7668 gnd.n7667 9.3005
R18291 gnd.n1988 gnd.n1987 9.3005
R18292 gnd.n7752 gnd.n7751 9.3005
R18293 gnd.n7353 gnd.n7352 9.3005
R18294 gnd.n7351 gnd.n7350 9.3005
R18295 gnd.n7344 gnd.n592 9.3005
R18296 gnd.n2905 gnd.n2637 9.3005
R18297 gnd.n2927 gnd.n2906 9.3005
R18298 gnd.n2926 gnd.n2907 9.3005
R18299 gnd.n2925 gnd.n2908 9.3005
R18300 gnd.n2911 gnd.n2909 9.3005
R18301 gnd.n2921 gnd.n2912 9.3005
R18302 gnd.n2920 gnd.n2913 9.3005
R18303 gnd.n2919 gnd.n2914 9.3005
R18304 gnd.n2917 gnd.n2916 9.3005
R18305 gnd.n2915 gnd.n2614 9.3005
R18306 gnd.n2612 gnd.n2611 9.3005
R18307 gnd.n2993 gnd.n2992 9.3005
R18308 gnd.n2994 gnd.n2610 9.3005
R18309 gnd.n2996 gnd.n2995 9.3005
R18310 gnd.n2608 gnd.n2607 9.3005
R18311 gnd.n3001 gnd.n3000 9.3005
R18312 gnd.n3002 gnd.n2606 9.3005
R18313 gnd.n3008 gnd.n3003 9.3005
R18314 gnd.n3007 gnd.n3004 9.3005
R18315 gnd.n3006 gnd.n3005 9.3005
R18316 gnd.n2590 gnd.n2589 9.3005
R18317 gnd.n3296 gnd.n3295 9.3005
R18318 gnd.n3297 gnd.n2588 9.3005
R18319 gnd.n3299 gnd.n3298 9.3005
R18320 gnd.n2586 gnd.n2585 9.3005
R18321 gnd.n3304 gnd.n3303 9.3005
R18322 gnd.n3305 gnd.n2584 9.3005
R18323 gnd.n3315 gnd.n3306 9.3005
R18324 gnd.n3314 gnd.n3307 9.3005
R18325 gnd.n3313 gnd.n3308 9.3005
R18326 gnd.n3310 gnd.n3309 9.3005
R18327 gnd.n2556 gnd.n2555 9.3005
R18328 gnd.n3332 gnd.n3331 9.3005
R18329 gnd.n3333 gnd.n2554 9.3005
R18330 gnd.n3335 gnd.n3334 9.3005
R18331 gnd.n2540 gnd.n2539 9.3005
R18332 gnd.n3365 gnd.n3364 9.3005
R18333 gnd.n3366 gnd.n2538 9.3005
R18334 gnd.n3377 gnd.n3367 9.3005
R18335 gnd.n3376 gnd.n3368 9.3005
R18336 gnd.n3375 gnd.n3369 9.3005
R18337 gnd.n3372 gnd.n3371 9.3005
R18338 gnd.n3370 gnd.n1691 9.3005
R18339 gnd.n4683 gnd.n1692 9.3005
R18340 gnd.n4682 gnd.n1693 9.3005
R18341 gnd.n4681 gnd.n1694 9.3005
R18342 gnd.n2503 gnd.n1695 9.3005
R18343 gnd.n2505 gnd.n2504 9.3005
R18344 gnd.n3531 gnd.n3530 9.3005
R18345 gnd.n3532 gnd.n2502 9.3005
R18346 gnd.n3536 gnd.n3533 9.3005
R18347 gnd.n3535 gnd.n3534 9.3005
R18348 gnd.n2482 gnd.n2481 9.3005
R18349 gnd.n3568 gnd.n3567 9.3005
R18350 gnd.n3569 gnd.n2480 9.3005
R18351 gnd.n3571 gnd.n3570 9.3005
R18352 gnd.n2454 gnd.n2453 9.3005
R18353 gnd.n3607 gnd.n3606 9.3005
R18354 gnd.n3608 gnd.n2452 9.3005
R18355 gnd.n3612 gnd.n3609 9.3005
R18356 gnd.n3611 gnd.n3610 9.3005
R18357 gnd.n2426 gnd.n2425 9.3005
R18358 gnd.n3647 gnd.n3646 9.3005
R18359 gnd.n3648 gnd.n2424 9.3005
R18360 gnd.n3651 gnd.n3650 9.3005
R18361 gnd.n3649 gnd.n2405 9.3005
R18362 gnd.n3679 gnd.n2406 9.3005
R18363 gnd.n3678 gnd.n2407 9.3005
R18364 gnd.n3677 gnd.n2408 9.3005
R18365 gnd.n2410 gnd.n2409 9.3005
R18366 gnd.n2412 gnd.n2411 9.3005
R18367 gnd.n2370 gnd.n2369 9.3005
R18368 gnd.n3742 gnd.n3741 9.3005
R18369 gnd.n3743 gnd.n2368 9.3005
R18370 gnd.n3747 gnd.n3744 9.3005
R18371 gnd.n3746 gnd.n3745 9.3005
R18372 gnd.n2345 gnd.n2344 9.3005
R18373 gnd.n3794 gnd.n3793 9.3005
R18374 gnd.n3795 gnd.n2343 9.3005
R18375 gnd.n3799 gnd.n3796 9.3005
R18376 gnd.n3798 gnd.n3797 9.3005
R18377 gnd.n2319 gnd.n2318 9.3005
R18378 gnd.n3831 gnd.n3830 9.3005
R18379 gnd.n3832 gnd.n2317 9.3005
R18380 gnd.n3834 gnd.n3833 9.3005
R18381 gnd.n2294 gnd.n2293 9.3005
R18382 gnd.n3892 gnd.n3891 9.3005
R18383 gnd.n3893 gnd.n2292 9.3005
R18384 gnd.n3897 gnd.n3894 9.3005
R18385 gnd.n3896 gnd.n3895 9.3005
R18386 gnd.n2271 gnd.n2270 9.3005
R18387 gnd.n3925 gnd.n3924 9.3005
R18388 gnd.n3926 gnd.n2269 9.3005
R18389 gnd.n3930 gnd.n3927 9.3005
R18390 gnd.n3929 gnd.n3928 9.3005
R18391 gnd.n2250 gnd.n2249 9.3005
R18392 gnd.n3977 gnd.n3976 9.3005
R18393 gnd.n3978 gnd.n2248 9.3005
R18394 gnd.n3982 gnd.n3979 9.3005
R18395 gnd.n3981 gnd.n3980 9.3005
R18396 gnd.n2221 gnd.n2220 9.3005
R18397 gnd.n4014 gnd.n4013 9.3005
R18398 gnd.n4015 gnd.n2219 9.3005
R18399 gnd.n4017 gnd.n4016 9.3005
R18400 gnd.n2132 gnd.n2131 9.3005
R18401 gnd.n4161 gnd.n4160 9.3005
R18402 gnd.n4162 gnd.n2130 9.3005
R18403 gnd.n4164 gnd.n4163 9.3005
R18404 gnd.n2119 gnd.n2118 9.3005
R18405 gnd.n4177 gnd.n4176 9.3005
R18406 gnd.n4178 gnd.n2117 9.3005
R18407 gnd.n4183 gnd.n4179 9.3005
R18408 gnd.n4182 gnd.n4181 9.3005
R18409 gnd.n4180 gnd.n2106 9.3005
R18410 gnd.n4196 gnd.n2105 9.3005
R18411 gnd.n4198 gnd.n4197 9.3005
R18412 gnd.n4199 gnd.n2104 9.3005
R18413 gnd.n4249 gnd.n4200 9.3005
R18414 gnd.n4248 gnd.n4201 9.3005
R18415 gnd.n4247 gnd.n4202 9.3005
R18416 gnd.n4205 gnd.n4203 9.3005
R18417 gnd.n4243 gnd.n4206 9.3005
R18418 gnd.n4242 gnd.n4207 9.3005
R18419 gnd.n4241 gnd.n4208 9.3005
R18420 gnd.n4211 gnd.n4209 9.3005
R18421 gnd.n4235 gnd.n4212 9.3005
R18422 gnd.n4234 gnd.n4213 9.3005
R18423 gnd.n4233 gnd.n4214 9.3005
R18424 gnd.n4217 gnd.n4215 9.3005
R18425 gnd.n4229 gnd.n4218 9.3005
R18426 gnd.n4228 gnd.n4219 9.3005
R18427 gnd.n4227 gnd.n4220 9.3005
R18428 gnd.n4224 gnd.n4221 9.3005
R18429 gnd.n4223 gnd.n4222 9.3005
R18430 gnd.n2059 gnd.n2058 9.3005
R18431 gnd.n4321 gnd.n4320 9.3005
R18432 gnd.n4322 gnd.n2057 9.3005
R18433 gnd.n4325 gnd.n4324 9.3005
R18434 gnd.n4323 gnd.n576 9.3005
R18435 gnd.n7367 gnd.n577 9.3005
R18436 gnd.n7366 gnd.n578 9.3005
R18437 gnd.n7365 gnd.n579 9.3005
R18438 gnd.n582 gnd.n580 9.3005
R18439 gnd.n7361 gnd.n583 9.3005
R18440 gnd.n7360 gnd.n584 9.3005
R18441 gnd.n7359 gnd.n585 9.3005
R18442 gnd.n588 gnd.n586 9.3005
R18443 gnd.n7355 gnd.n589 9.3005
R18444 gnd.n7354 gnd.n590 9.3005
R18445 gnd.n2867 gnd.n2866 9.3005
R18446 gnd.n2805 gnd.n2743 9.3005
R18447 gnd.n2808 gnd.n2807 9.3005
R18448 gnd.n2809 gnd.n2742 9.3005
R18449 gnd.n2812 gnd.n2810 9.3005
R18450 gnd.n2813 gnd.n2741 9.3005
R18451 gnd.n2816 gnd.n2815 9.3005
R18452 gnd.n2817 gnd.n2740 9.3005
R18453 gnd.n2820 gnd.n2818 9.3005
R18454 gnd.n2821 gnd.n2739 9.3005
R18455 gnd.n2824 gnd.n2823 9.3005
R18456 gnd.n2825 gnd.n2738 9.3005
R18457 gnd.n2828 gnd.n2826 9.3005
R18458 gnd.n2829 gnd.n2737 9.3005
R18459 gnd.n2832 gnd.n2831 9.3005
R18460 gnd.n2833 gnd.n2736 9.3005
R18461 gnd.n2836 gnd.n2834 9.3005
R18462 gnd.n2837 gnd.n2735 9.3005
R18463 gnd.n2840 gnd.n2839 9.3005
R18464 gnd.n2841 gnd.n2734 9.3005
R18465 gnd.n2844 gnd.n2842 9.3005
R18466 gnd.n2845 gnd.n2733 9.3005
R18467 gnd.n2848 gnd.n2847 9.3005
R18468 gnd.n2849 gnd.n2732 9.3005
R18469 gnd.n2852 gnd.n2850 9.3005
R18470 gnd.n2853 gnd.n2731 9.3005
R18471 gnd.n2856 gnd.n2855 9.3005
R18472 gnd.n2857 gnd.n2730 9.3005
R18473 gnd.n2860 gnd.n2858 9.3005
R18474 gnd.n2861 gnd.n2729 9.3005
R18475 gnd.n2864 gnd.n2863 9.3005
R18476 gnd.n2865 gnd.n2728 9.3005
R18477 gnd.n2804 gnd.n2802 9.3005
R18478 gnd.n2798 gnd.n2797 9.3005
R18479 gnd.n2796 gnd.n2748 9.3005
R18480 gnd.n2795 gnd.n2794 9.3005
R18481 gnd.n2791 gnd.n2751 9.3005
R18482 gnd.n2790 gnd.n2787 9.3005
R18483 gnd.n2786 gnd.n2752 9.3005
R18484 gnd.n2785 gnd.n2784 9.3005
R18485 gnd.n2781 gnd.n2753 9.3005
R18486 gnd.n2780 gnd.n2777 9.3005
R18487 gnd.n2776 gnd.n2754 9.3005
R18488 gnd.n2775 gnd.n2774 9.3005
R18489 gnd.n2771 gnd.n2755 9.3005
R18490 gnd.n2770 gnd.n2767 9.3005
R18491 gnd.n2766 gnd.n2756 9.3005
R18492 gnd.n2765 gnd.n2764 9.3005
R18493 gnd.n2761 gnd.n2757 9.3005
R18494 gnd.n2760 gnd.n1254 9.3005
R18495 gnd.n2799 gnd.n2744 9.3005
R18496 gnd.n2801 gnd.n2800 9.3005
R18497 gnd.n4761 gnd.n1618 9.3005
R18498 gnd.n4764 gnd.n1617 9.3005
R18499 gnd.n4765 gnd.n1616 9.3005
R18500 gnd.n4768 gnd.n1615 9.3005
R18501 gnd.n4769 gnd.n1614 9.3005
R18502 gnd.n4772 gnd.n1613 9.3005
R18503 gnd.n4773 gnd.n1612 9.3005
R18504 gnd.n4776 gnd.n1611 9.3005
R18505 gnd.n4778 gnd.n1608 9.3005
R18506 gnd.n4781 gnd.n1607 9.3005
R18507 gnd.n4782 gnd.n1606 9.3005
R18508 gnd.n4785 gnd.n1605 9.3005
R18509 gnd.n4786 gnd.n1604 9.3005
R18510 gnd.n4789 gnd.n1603 9.3005
R18511 gnd.n4790 gnd.n1602 9.3005
R18512 gnd.n4793 gnd.n1601 9.3005
R18513 gnd.n4794 gnd.n1600 9.3005
R18514 gnd.n4797 gnd.n1599 9.3005
R18515 gnd.n4798 gnd.n1598 9.3005
R18516 gnd.n4801 gnd.n1597 9.3005
R18517 gnd.n4802 gnd.n1596 9.3005
R18518 gnd.n4805 gnd.n1595 9.3005
R18519 gnd.n4806 gnd.n1594 9.3005
R18520 gnd.n4807 gnd.n1593 9.3005
R18521 gnd.n1550 gnd.n1549 9.3005
R18522 gnd.n4813 gnd.n4812 9.3005
R18523 gnd.n3200 gnd.n3197 9.3005
R18524 gnd.n3204 gnd.n3203 9.3005
R18525 gnd.n3205 gnd.n3195 9.3005
R18526 gnd.n3207 gnd.n3206 9.3005
R18527 gnd.n3210 gnd.n3194 9.3005
R18528 gnd.n3214 gnd.n3213 9.3005
R18529 gnd.n3215 gnd.n3193 9.3005
R18530 gnd.n3218 gnd.n3216 9.3005
R18531 gnd.n3219 gnd.n3189 9.3005
R18532 gnd.n3223 gnd.n3222 9.3005
R18533 gnd.n3224 gnd.n3188 9.3005
R18534 gnd.n3226 gnd.n3225 9.3005
R18535 gnd.n3229 gnd.n3187 9.3005
R18536 gnd.n3233 gnd.n3232 9.3005
R18537 gnd.n3234 gnd.n3186 9.3005
R18538 gnd.n3236 gnd.n3235 9.3005
R18539 gnd.n3239 gnd.n3185 9.3005
R18540 gnd.n3243 gnd.n3242 9.3005
R18541 gnd.n3244 gnd.n3184 9.3005
R18542 gnd.n3246 gnd.n3245 9.3005
R18543 gnd.n3249 gnd.n3183 9.3005
R18544 gnd.n3253 gnd.n3252 9.3005
R18545 gnd.n3254 gnd.n3182 9.3005
R18546 gnd.n3256 gnd.n3255 9.3005
R18547 gnd.n3259 gnd.n3181 9.3005
R18548 gnd.n3263 gnd.n3262 9.3005
R18549 gnd.n3264 gnd.n3180 9.3005
R18550 gnd.n3267 gnd.n3265 9.3005
R18551 gnd.n3268 gnd.n3176 9.3005
R18552 gnd.n3271 gnd.n3270 9.3005
R18553 gnd.n3196 gnd.n1619 9.3005
R18554 gnd.n1276 gnd.n1256 9.3005
R18555 gnd.n2670 gnd.n1277 9.3005
R18556 gnd.n4979 gnd.n1278 9.3005
R18557 gnd.n4978 gnd.n1279 9.3005
R18558 gnd.n4977 gnd.n1280 9.3005
R18559 gnd.n2676 gnd.n1281 9.3005
R18560 gnd.n4967 gnd.n1297 9.3005
R18561 gnd.n4966 gnd.n1298 9.3005
R18562 gnd.n4965 gnd.n1299 9.3005
R18563 gnd.n2683 gnd.n1300 9.3005
R18564 gnd.n4955 gnd.n1316 9.3005
R18565 gnd.n4954 gnd.n1317 9.3005
R18566 gnd.n4953 gnd.n1318 9.3005
R18567 gnd.n2690 gnd.n1319 9.3005
R18568 gnd.n4943 gnd.n1335 9.3005
R18569 gnd.n4942 gnd.n1336 9.3005
R18570 gnd.n4941 gnd.n1337 9.3005
R18571 gnd.n2697 gnd.n1338 9.3005
R18572 gnd.n4931 gnd.n1354 9.3005
R18573 gnd.n4930 gnd.n1355 9.3005
R18574 gnd.n4929 gnd.n1356 9.3005
R18575 gnd.n2704 gnd.n1357 9.3005
R18576 gnd.n4919 gnd.n1373 9.3005
R18577 gnd.n4918 gnd.n1374 9.3005
R18578 gnd.n4917 gnd.n1375 9.3005
R18579 gnd.n2711 gnd.n1376 9.3005
R18580 gnd.n4907 gnd.n1391 9.3005
R18581 gnd.n4906 gnd.n1392 9.3005
R18582 gnd.n4905 gnd.n1393 9.3005
R18583 gnd.n2720 gnd.n1394 9.3005
R18584 gnd.n2722 gnd.n2721 9.3005
R18585 gnd.n2668 gnd.n2663 9.3005
R18586 gnd.n2883 gnd.n2664 9.3005
R18587 gnd.n2882 gnd.n2665 9.3005
R18588 gnd.n2881 gnd.n2879 9.3005
R18589 gnd.n2666 gnd.n1417 9.3005
R18590 gnd.n4894 gnd.n1418 9.3005
R18591 gnd.n4893 gnd.n1419 9.3005
R18592 gnd.n4892 gnd.n1420 9.3005
R18593 gnd.n2630 gnd.n1421 9.3005
R18594 gnd.n4882 gnd.n1436 9.3005
R18595 gnd.n4881 gnd.n1437 9.3005
R18596 gnd.n4880 gnd.n1438 9.3005
R18597 gnd.n2624 gnd.n1439 9.3005
R18598 gnd.n4870 gnd.n1457 9.3005
R18599 gnd.n4869 gnd.n1458 9.3005
R18600 gnd.n4868 gnd.n1459 9.3005
R18601 gnd.n2958 gnd.n1460 9.3005
R18602 gnd.n4858 gnd.n1476 9.3005
R18603 gnd.n4857 gnd.n1477 9.3005
R18604 gnd.n4856 gnd.n1478 9.3005
R18605 gnd.n2968 gnd.n1479 9.3005
R18606 gnd.n4846 gnd.n1497 9.3005
R18607 gnd.n4845 gnd.n1498 9.3005
R18608 gnd.n4844 gnd.n1499 9.3005
R18609 gnd.n2599 gnd.n1500 9.3005
R18610 gnd.n4834 gnd.n1516 9.3005
R18611 gnd.n4833 gnd.n1517 9.3005
R18612 gnd.n4832 gnd.n1518 9.3005
R18613 gnd.n3025 gnd.n1519 9.3005
R18614 gnd.n4822 gnd.n1537 9.3005
R18615 gnd.n4821 gnd.n1538 9.3005
R18616 gnd.n4820 gnd.n1539 9.3005
R18617 gnd.n3273 gnd.n1540 9.3005
R18618 gnd.n4991 gnd.n1255 9.3005
R18619 gnd.n1257 gnd.n1256 9.3005
R18620 gnd.n2671 gnd.n2670 9.3005
R18621 gnd.n2672 gnd.n1278 9.3005
R18622 gnd.n2674 gnd.n1279 9.3005
R18623 gnd.n2675 gnd.n1280 9.3005
R18624 gnd.n2678 gnd.n2676 9.3005
R18625 gnd.n2679 gnd.n1297 9.3005
R18626 gnd.n2681 gnd.n1298 9.3005
R18627 gnd.n2682 gnd.n1299 9.3005
R18628 gnd.n2685 gnd.n2683 9.3005
R18629 gnd.n2686 gnd.n1316 9.3005
R18630 gnd.n2688 gnd.n1317 9.3005
R18631 gnd.n2689 gnd.n1318 9.3005
R18632 gnd.n2692 gnd.n2690 9.3005
R18633 gnd.n2693 gnd.n1335 9.3005
R18634 gnd.n2695 gnd.n1336 9.3005
R18635 gnd.n2696 gnd.n1337 9.3005
R18636 gnd.n2699 gnd.n2697 9.3005
R18637 gnd.n2700 gnd.n1354 9.3005
R18638 gnd.n2702 gnd.n1355 9.3005
R18639 gnd.n2703 gnd.n1356 9.3005
R18640 gnd.n2706 gnd.n2704 9.3005
R18641 gnd.n2707 gnd.n1373 9.3005
R18642 gnd.n2709 gnd.n1374 9.3005
R18643 gnd.n2710 gnd.n1375 9.3005
R18644 gnd.n2713 gnd.n2711 9.3005
R18645 gnd.n2714 gnd.n1391 9.3005
R18646 gnd.n2716 gnd.n1392 9.3005
R18647 gnd.n2717 gnd.n1393 9.3005
R18648 gnd.n2720 gnd.n2719 9.3005
R18649 gnd.n2721 gnd.n2667 9.3005
R18650 gnd.n2871 gnd.n2668 9.3005
R18651 gnd.n2872 gnd.n2664 9.3005
R18652 gnd.n2873 gnd.n2665 9.3005
R18653 gnd.n2879 gnd.n2878 9.3005
R18654 gnd.n2876 gnd.n2666 9.3005
R18655 gnd.n2875 gnd.n1418 9.3005
R18656 gnd.n2874 gnd.n1419 9.3005
R18657 gnd.n2629 gnd.n1420 9.3005
R18658 gnd.n2940 gnd.n2630 9.3005
R18659 gnd.n2941 gnd.n1436 9.3005
R18660 gnd.n2942 gnd.n1437 9.3005
R18661 gnd.n2623 gnd.n1438 9.3005
R18662 gnd.n2954 gnd.n2624 9.3005
R18663 gnd.n2955 gnd.n1457 9.3005
R18664 gnd.n2956 gnd.n1458 9.3005
R18665 gnd.n2957 gnd.n1459 9.3005
R18666 gnd.n2961 gnd.n2958 9.3005
R18667 gnd.n2962 gnd.n1476 9.3005
R18668 gnd.n2966 gnd.n1477 9.3005
R18669 gnd.n2967 gnd.n1478 9.3005
R18670 gnd.n2971 gnd.n2968 9.3005
R18671 gnd.n2970 gnd.n1497 9.3005
R18672 gnd.n2969 gnd.n1498 9.3005
R18673 gnd.n2598 gnd.n1499 9.3005
R18674 gnd.n3021 gnd.n2599 9.3005
R18675 gnd.n3022 gnd.n1516 9.3005
R18676 gnd.n3023 gnd.n1517 9.3005
R18677 gnd.n3024 gnd.n1518 9.3005
R18678 gnd.n3028 gnd.n3025 9.3005
R18679 gnd.n3029 gnd.n1537 9.3005
R18680 gnd.n3276 gnd.n1538 9.3005
R18681 gnd.n3275 gnd.n1539 9.3005
R18682 gnd.n3274 gnd.n3273 9.3005
R18683 gnd.n4991 gnd.n4990 9.3005
R18684 gnd.n4995 gnd.n4994 9.3005
R18685 gnd.n4998 gnd.n1250 9.3005
R18686 gnd.n4999 gnd.n1249 9.3005
R18687 gnd.n5002 gnd.n1248 9.3005
R18688 gnd.n5003 gnd.n1247 9.3005
R18689 gnd.n5006 gnd.n1246 9.3005
R18690 gnd.n5007 gnd.n1245 9.3005
R18691 gnd.n5010 gnd.n1244 9.3005
R18692 gnd.n5011 gnd.n1243 9.3005
R18693 gnd.n5014 gnd.n1242 9.3005
R18694 gnd.n5015 gnd.n1241 9.3005
R18695 gnd.n5018 gnd.n1240 9.3005
R18696 gnd.n5019 gnd.n1239 9.3005
R18697 gnd.n5022 gnd.n1238 9.3005
R18698 gnd.n5023 gnd.n1237 9.3005
R18699 gnd.n5026 gnd.n1236 9.3005
R18700 gnd.n5027 gnd.n1235 9.3005
R18701 gnd.n5030 gnd.n1234 9.3005
R18702 gnd.n5031 gnd.n1233 9.3005
R18703 gnd.n5034 gnd.n1232 9.3005
R18704 gnd.n5038 gnd.n1228 9.3005
R18705 gnd.n5039 gnd.n1227 9.3005
R18706 gnd.n5042 gnd.n1226 9.3005
R18707 gnd.n5043 gnd.n1225 9.3005
R18708 gnd.n5046 gnd.n1224 9.3005
R18709 gnd.n5047 gnd.n1223 9.3005
R18710 gnd.n5050 gnd.n1222 9.3005
R18711 gnd.n5051 gnd.n1221 9.3005
R18712 gnd.n5054 gnd.n1220 9.3005
R18713 gnd.n5055 gnd.n1219 9.3005
R18714 gnd.n5058 gnd.n1218 9.3005
R18715 gnd.n5059 gnd.n1217 9.3005
R18716 gnd.n5062 gnd.n1216 9.3005
R18717 gnd.n5063 gnd.n1215 9.3005
R18718 gnd.n5066 gnd.n1214 9.3005
R18719 gnd.n5067 gnd.n1213 9.3005
R18720 gnd.n5070 gnd.n1212 9.3005
R18721 gnd.n5071 gnd.n1211 9.3005
R18722 gnd.n5074 gnd.n1210 9.3005
R18723 gnd.n5076 gnd.n1207 9.3005
R18724 gnd.n5079 gnd.n1206 9.3005
R18725 gnd.n5080 gnd.n1205 9.3005
R18726 gnd.n5083 gnd.n1204 9.3005
R18727 gnd.n5084 gnd.n1203 9.3005
R18728 gnd.n5087 gnd.n1202 9.3005
R18729 gnd.n5088 gnd.n1201 9.3005
R18730 gnd.n5091 gnd.n1200 9.3005
R18731 gnd.n5092 gnd.n1199 9.3005
R18732 gnd.n5095 gnd.n1198 9.3005
R18733 gnd.n5096 gnd.n1197 9.3005
R18734 gnd.n5099 gnd.n1196 9.3005
R18735 gnd.n5100 gnd.n1195 9.3005
R18736 gnd.n5103 gnd.n1194 9.3005
R18737 gnd.n5105 gnd.n1193 9.3005
R18738 gnd.n5106 gnd.n1192 9.3005
R18739 gnd.n5107 gnd.n1191 9.3005
R18740 gnd.n5108 gnd.n1190 9.3005
R18741 gnd.n5035 gnd.n1229 9.3005
R18742 gnd.n4993 gnd.n1251 9.3005
R18743 gnd.n4985 gnd.n1265 9.3005
R18744 gnd.n4984 gnd.n1266 9.3005
R18745 gnd.n4983 gnd.n1267 9.3005
R18746 gnd.n1287 gnd.n1268 9.3005
R18747 gnd.n4973 gnd.n1288 9.3005
R18748 gnd.n4972 gnd.n1289 9.3005
R18749 gnd.n4971 gnd.n1290 9.3005
R18750 gnd.n1305 gnd.n1291 9.3005
R18751 gnd.n4961 gnd.n1306 9.3005
R18752 gnd.n4960 gnd.n1307 9.3005
R18753 gnd.n4959 gnd.n1308 9.3005
R18754 gnd.n1325 gnd.n1309 9.3005
R18755 gnd.n4949 gnd.n1326 9.3005
R18756 gnd.n4948 gnd.n1327 9.3005
R18757 gnd.n4947 gnd.n1328 9.3005
R18758 gnd.n1343 gnd.n1329 9.3005
R18759 gnd.n4937 gnd.n1344 9.3005
R18760 gnd.n4936 gnd.n1345 9.3005
R18761 gnd.n4935 gnd.n1346 9.3005
R18762 gnd.n1363 gnd.n1347 9.3005
R18763 gnd.n4925 gnd.n1364 9.3005
R18764 gnd.n4924 gnd.n1365 9.3005
R18765 gnd.n4923 gnd.n1366 9.3005
R18766 gnd.n1381 gnd.n1367 9.3005
R18767 gnd.n4913 gnd.n1382 9.3005
R18768 gnd.n4912 gnd.n1383 9.3005
R18769 gnd.n1408 gnd.n1402 9.3005
R18770 gnd.n4888 gnd.n1427 9.3005
R18771 gnd.n4887 gnd.n1428 9.3005
R18772 gnd.n4886 gnd.n1429 9.3005
R18773 gnd.n1446 gnd.n1430 9.3005
R18774 gnd.n4876 gnd.n1447 9.3005
R18775 gnd.n4875 gnd.n1448 9.3005
R18776 gnd.n4874 gnd.n1449 9.3005
R18777 gnd.n1466 gnd.n1450 9.3005
R18778 gnd.n4864 gnd.n1467 9.3005
R18779 gnd.n4863 gnd.n1468 9.3005
R18780 gnd.n4862 gnd.n1469 9.3005
R18781 gnd.n1486 gnd.n1470 9.3005
R18782 gnd.n4852 gnd.n1487 9.3005
R18783 gnd.n4851 gnd.n1488 9.3005
R18784 gnd.n4850 gnd.n1489 9.3005
R18785 gnd.n1506 gnd.n1490 9.3005
R18786 gnd.n4840 gnd.n1507 9.3005
R18787 gnd.n4839 gnd.n1508 9.3005
R18788 gnd.n4838 gnd.n1509 9.3005
R18789 gnd.n1526 gnd.n1510 9.3005
R18790 gnd.n4828 gnd.n1527 9.3005
R18791 gnd.n4827 gnd.n1528 9.3005
R18792 gnd.n4826 gnd.n1529 9.3005
R18793 gnd.n1547 gnd.n1530 9.3005
R18794 gnd.n4816 gnd.n1548 9.3005
R18795 gnd.n4815 gnd.n4814 9.3005
R18796 gnd.n1264 gnd.n1263 9.3005
R18797 gnd.n4899 gnd.n4898 9.3005
R18798 gnd.n2639 gnd.n2638 9.3005
R18799 gnd.n2904 gnd.n2903 9.3005
R18800 gnd.n2656 gnd.n2655 9.3005
R18801 gnd.n2654 gnd.n1116 9.3005
R18802 gnd.n6580 gnd.n1115 9.3005
R18803 gnd.n6581 gnd.n1114 9.3005
R18804 gnd.n6582 gnd.n1113 9.3005
R18805 gnd.n1112 gnd.n1108 9.3005
R18806 gnd.n6588 gnd.n1107 9.3005
R18807 gnd.n6589 gnd.n1106 9.3005
R18808 gnd.n6590 gnd.n1105 9.3005
R18809 gnd.n1104 gnd.n1100 9.3005
R18810 gnd.n6596 gnd.n1099 9.3005
R18811 gnd.n6597 gnd.n1098 9.3005
R18812 gnd.n6598 gnd.n1097 9.3005
R18813 gnd.n1096 gnd.n1092 9.3005
R18814 gnd.n6604 gnd.n1091 9.3005
R18815 gnd.n6605 gnd.n1090 9.3005
R18816 gnd.n6606 gnd.n1089 9.3005
R18817 gnd.n1088 gnd.n1084 9.3005
R18818 gnd.n6612 gnd.n1083 9.3005
R18819 gnd.n6613 gnd.n1082 9.3005
R18820 gnd.n6614 gnd.n1081 9.3005
R18821 gnd.n1080 gnd.n1076 9.3005
R18822 gnd.n6620 gnd.n1075 9.3005
R18823 gnd.n6621 gnd.n1074 9.3005
R18824 gnd.n6622 gnd.n1073 9.3005
R18825 gnd.n1072 gnd.n1068 9.3005
R18826 gnd.n6628 gnd.n1067 9.3005
R18827 gnd.n6629 gnd.n1066 9.3005
R18828 gnd.n6630 gnd.n1065 9.3005
R18829 gnd.n1064 gnd.n1060 9.3005
R18830 gnd.n6636 gnd.n1059 9.3005
R18831 gnd.n6637 gnd.n1058 9.3005
R18832 gnd.n6638 gnd.n1057 9.3005
R18833 gnd.n1056 gnd.n1052 9.3005
R18834 gnd.n6644 gnd.n1051 9.3005
R18835 gnd.n6645 gnd.n1050 9.3005
R18836 gnd.n6646 gnd.n1049 9.3005
R18837 gnd.n1048 gnd.n1044 9.3005
R18838 gnd.n6652 gnd.n1043 9.3005
R18839 gnd.n6653 gnd.n1042 9.3005
R18840 gnd.n6654 gnd.n1041 9.3005
R18841 gnd.n1040 gnd.n1036 9.3005
R18842 gnd.n6660 gnd.n1035 9.3005
R18843 gnd.n6661 gnd.n1034 9.3005
R18844 gnd.n6662 gnd.n1033 9.3005
R18845 gnd.n1032 gnd.n1028 9.3005
R18846 gnd.n6668 gnd.n1027 9.3005
R18847 gnd.n6669 gnd.n1026 9.3005
R18848 gnd.n6670 gnd.n1025 9.3005
R18849 gnd.n1024 gnd.n1020 9.3005
R18850 gnd.n6676 gnd.n1019 9.3005
R18851 gnd.n6677 gnd.n1018 9.3005
R18852 gnd.n6678 gnd.n1017 9.3005
R18853 gnd.n1016 gnd.n1012 9.3005
R18854 gnd.n6684 gnd.n1011 9.3005
R18855 gnd.n6685 gnd.n1010 9.3005
R18856 gnd.n6686 gnd.n1009 9.3005
R18857 gnd.n1008 gnd.n1004 9.3005
R18858 gnd.n6692 gnd.n1003 9.3005
R18859 gnd.n6693 gnd.n1002 9.3005
R18860 gnd.n6694 gnd.n1001 9.3005
R18861 gnd.n1000 gnd.n996 9.3005
R18862 gnd.n6700 gnd.n995 9.3005
R18863 gnd.n6701 gnd.n994 9.3005
R18864 gnd.n6702 gnd.n993 9.3005
R18865 gnd.n992 gnd.n988 9.3005
R18866 gnd.n6708 gnd.n987 9.3005
R18867 gnd.n6709 gnd.n986 9.3005
R18868 gnd.n6710 gnd.n985 9.3005
R18869 gnd.n984 gnd.n980 9.3005
R18870 gnd.n6716 gnd.n979 9.3005
R18871 gnd.n6717 gnd.n978 9.3005
R18872 gnd.n6718 gnd.n977 9.3005
R18873 gnd.n976 gnd.n972 9.3005
R18874 gnd.n6724 gnd.n971 9.3005
R18875 gnd.n6725 gnd.n970 9.3005
R18876 gnd.n6726 gnd.n969 9.3005
R18877 gnd.n968 gnd.n964 9.3005
R18878 gnd.n6732 gnd.n963 9.3005
R18879 gnd.n6733 gnd.n962 9.3005
R18880 gnd.n6734 gnd.n961 9.3005
R18881 gnd.n960 gnd.n956 9.3005
R18882 gnd.n6740 gnd.n955 9.3005
R18883 gnd.n6741 gnd.n954 9.3005
R18884 gnd.n6742 gnd.n953 9.3005
R18885 gnd.n2658 gnd.n2657 9.3005
R18886 gnd.n4254 gnd.n1789 9.3005
R18887 gnd.n3340 gnd.n3339 9.3005
R18888 gnd.n3341 gnd.n2546 9.3005
R18889 gnd.n3360 gnd.n3359 9.3005
R18890 gnd.n3358 gnd.n2547 9.3005
R18891 gnd.n3357 gnd.n3356 9.3005
R18892 gnd.n3355 gnd.n3342 9.3005
R18893 gnd.n3354 gnd.n3353 9.3005
R18894 gnd.n3352 gnd.n3345 9.3005
R18895 gnd.n3351 gnd.n3350 9.3005
R18896 gnd.n3349 gnd.n3346 9.3005
R18897 gnd.n1703 gnd.n1701 9.3005
R18898 gnd.n4677 gnd.n4676 9.3005
R18899 gnd.n4675 gnd.n1702 9.3005
R18900 gnd.n4674 gnd.n4673 9.3005
R18901 gnd.n4672 gnd.n1704 9.3005
R18902 gnd.n4671 gnd.n4670 9.3005
R18903 gnd.n4669 gnd.n1708 9.3005
R18904 gnd.n4668 gnd.n4667 9.3005
R18905 gnd.n4666 gnd.n1709 9.3005
R18906 gnd.n4665 gnd.n4664 9.3005
R18907 gnd.n4663 gnd.n1713 9.3005
R18908 gnd.n4662 gnd.n4661 9.3005
R18909 gnd.n4660 gnd.n1714 9.3005
R18910 gnd.n4659 gnd.n4658 9.3005
R18911 gnd.n4657 gnd.n1718 9.3005
R18912 gnd.n4656 gnd.n4655 9.3005
R18913 gnd.n4654 gnd.n1719 9.3005
R18914 gnd.n4653 gnd.n4652 9.3005
R18915 gnd.n4651 gnd.n1723 9.3005
R18916 gnd.n4650 gnd.n4649 9.3005
R18917 gnd.n4648 gnd.n1724 9.3005
R18918 gnd.n4647 gnd.n4646 9.3005
R18919 gnd.n4645 gnd.n1728 9.3005
R18920 gnd.n4644 gnd.n4643 9.3005
R18921 gnd.n4642 gnd.n1729 9.3005
R18922 gnd.n4641 gnd.n4640 9.3005
R18923 gnd.n4639 gnd.n1733 9.3005
R18924 gnd.n4638 gnd.n4637 9.3005
R18925 gnd.n4636 gnd.n1734 9.3005
R18926 gnd.n4635 gnd.n4634 9.3005
R18927 gnd.n4633 gnd.n1738 9.3005
R18928 gnd.n4632 gnd.n4631 9.3005
R18929 gnd.n4630 gnd.n1739 9.3005
R18930 gnd.n4629 gnd.n4628 9.3005
R18931 gnd.n4627 gnd.n1743 9.3005
R18932 gnd.n4626 gnd.n4625 9.3005
R18933 gnd.n4624 gnd.n1744 9.3005
R18934 gnd.n4623 gnd.n4622 9.3005
R18935 gnd.n4621 gnd.n1748 9.3005
R18936 gnd.n4620 gnd.n4619 9.3005
R18937 gnd.n4618 gnd.n1749 9.3005
R18938 gnd.n4617 gnd.n4616 9.3005
R18939 gnd.n4615 gnd.n1753 9.3005
R18940 gnd.n4614 gnd.n4613 9.3005
R18941 gnd.n4612 gnd.n1754 9.3005
R18942 gnd.n4611 gnd.n4610 9.3005
R18943 gnd.n4609 gnd.n1758 9.3005
R18944 gnd.n4608 gnd.n4607 9.3005
R18945 gnd.n4606 gnd.n1759 9.3005
R18946 gnd.n4605 gnd.n4604 9.3005
R18947 gnd.n4603 gnd.n1763 9.3005
R18948 gnd.n4602 gnd.n4601 9.3005
R18949 gnd.n4600 gnd.n1764 9.3005
R18950 gnd.n4599 gnd.n4598 9.3005
R18951 gnd.n4597 gnd.n1768 9.3005
R18952 gnd.n4596 gnd.n4595 9.3005
R18953 gnd.n4594 gnd.n1769 9.3005
R18954 gnd.n4593 gnd.n4592 9.3005
R18955 gnd.n4591 gnd.n1773 9.3005
R18956 gnd.n4590 gnd.n4589 9.3005
R18957 gnd.n4588 gnd.n1774 9.3005
R18958 gnd.n4587 gnd.n4586 9.3005
R18959 gnd.n4585 gnd.n1778 9.3005
R18960 gnd.n4584 gnd.n4583 9.3005
R18961 gnd.n4582 gnd.n1779 9.3005
R18962 gnd.n4581 gnd.n4580 9.3005
R18963 gnd.n4579 gnd.n1783 9.3005
R18964 gnd.n4578 gnd.n4577 9.3005
R18965 gnd.n4576 gnd.n1784 9.3005
R18966 gnd.n4575 gnd.n4574 9.3005
R18967 gnd.n4573 gnd.n1788 9.3005
R18968 gnd.n4572 gnd.n4571 9.3005
R18969 gnd.n2549 gnd.n2548 9.3005
R18970 gnd.n3326 gnd.n3325 9.3005
R18971 gnd.n2646 gnd.n2645 9.3005
R18972 gnd.n2894 gnd.n2893 9.3005
R18973 gnd.n2895 gnd.n2644 9.3005
R18974 gnd.n2897 gnd.n2896 9.3005
R18975 gnd.n2633 gnd.n2632 9.3005
R18976 gnd.n2933 gnd.n2932 9.3005
R18977 gnd.n2934 gnd.n2631 9.3005
R18978 gnd.n2936 gnd.n2935 9.3005
R18979 gnd.n2627 gnd.n2626 9.3005
R18980 gnd.n2947 gnd.n2946 9.3005
R18981 gnd.n2948 gnd.n2625 9.3005
R18982 gnd.n2950 gnd.n2949 9.3005
R18983 gnd.n2618 gnd.n2616 9.3005
R18984 gnd.n2985 gnd.n2984 9.3005
R18985 gnd.n2983 gnd.n2617 9.3005
R18986 gnd.n2982 gnd.n2981 9.3005
R18987 gnd.n2980 gnd.n2619 9.3005
R18988 gnd.n2979 gnd.n2978 9.3005
R18989 gnd.n2977 gnd.n2622 9.3005
R18990 gnd.n2976 gnd.n2975 9.3005
R18991 gnd.n2602 gnd.n2601 9.3005
R18992 gnd.n3014 gnd.n3013 9.3005
R18993 gnd.n3015 gnd.n2600 9.3005
R18994 gnd.n3017 gnd.n3016 9.3005
R18995 gnd.n2595 gnd.n2593 9.3005
R18996 gnd.n3289 gnd.n3288 9.3005
R18997 gnd.n3287 gnd.n2594 9.3005
R18998 gnd.n3286 gnd.n3285 9.3005
R18999 gnd.n3284 gnd.n2596 9.3005
R19000 gnd.n3283 gnd.n3282 9.3005
R19001 gnd.n3281 gnd.n3280 9.3005
R19002 gnd.n2580 gnd.n2575 9.3005
R19003 gnd.n3167 gnd.n3166 9.3005
R19004 gnd.n3066 gnd.n3065 9.3005
R19005 gnd.n3161 gnd.n3160 9.3005
R19006 gnd.n3159 gnd.n3158 9.3005
R19007 gnd.n3078 gnd.n3077 9.3005
R19008 gnd.n3153 gnd.n3152 9.3005
R19009 gnd.n3151 gnd.n3150 9.3005
R19010 gnd.n3086 gnd.n3085 9.3005
R19011 gnd.n3145 gnd.n3144 9.3005
R19012 gnd.n3143 gnd.n3142 9.3005
R19013 gnd.n3098 gnd.n3097 9.3005
R19014 gnd.n3137 gnd.n3136 9.3005
R19015 gnd.n3135 gnd.n3134 9.3005
R19016 gnd.n3106 gnd.n3105 9.3005
R19017 gnd.n3129 gnd.n3128 9.3005
R19018 gnd.n3127 gnd.n3126 9.3005
R19019 gnd.n3117 gnd.n2579 9.3005
R19020 gnd.n3322 gnd.n3321 9.3005
R19021 gnd.n3169 gnd.n3168 9.3005
R19022 gnd.n3323 gnd.n2574 9.3005
R19023 gnd.n3123 gnd.n2576 9.3005
R19024 gnd.n3125 gnd.n3124 9.3005
R19025 gnd.n3112 gnd.n3111 9.3005
R19026 gnd.n3131 gnd.n3130 9.3005
R19027 gnd.n3133 gnd.n3132 9.3005
R19028 gnd.n3102 gnd.n3101 9.3005
R19029 gnd.n3139 gnd.n3138 9.3005
R19030 gnd.n3141 gnd.n3140 9.3005
R19031 gnd.n3092 gnd.n3091 9.3005
R19032 gnd.n3147 gnd.n3146 9.3005
R19033 gnd.n3149 gnd.n3148 9.3005
R19034 gnd.n3082 gnd.n3081 9.3005
R19035 gnd.n3155 gnd.n3154 9.3005
R19036 gnd.n3157 gnd.n3156 9.3005
R19037 gnd.n3072 gnd.n3071 9.3005
R19038 gnd.n3163 gnd.n3162 9.3005
R19039 gnd.n3165 gnd.n3164 9.3005
R19040 gnd.n3063 gnd.n3062 9.3005
R19041 gnd.n3171 gnd.n3170 9.3005
R19042 gnd.n3172 gnd.n3030 9.3005
R19043 gnd.n3174 gnd.n3173 9.3005
R19044 gnd.n3057 gnd.n3031 9.3005
R19045 gnd.n3056 gnd.n3055 9.3005
R19046 gnd.n3054 gnd.n3032 9.3005
R19047 gnd.n3053 gnd.n3052 9.3005
R19048 gnd.n3049 gnd.n3035 9.3005
R19049 gnd.n3048 gnd.n3036 9.3005
R19050 gnd.n3043 gnd.n3037 9.3005
R19051 gnd.n3042 gnd.n3041 9.3005
R19052 gnd.n3040 gnd.n3038 9.3005
R19053 gnd.n2531 gnd.n2530 9.3005
R19054 gnd.n3382 gnd.n3381 9.3005
R19055 gnd.n3383 gnd.n2529 9.3005
R19056 gnd.n3385 gnd.n3384 9.3005
R19057 gnd.n2527 gnd.n2526 9.3005
R19058 gnd.n3390 gnd.n3389 9.3005
R19059 gnd.n3391 gnd.n2524 9.3005
R19060 gnd.n3402 gnd.n3401 9.3005
R19061 gnd.n3400 gnd.n2525 9.3005
R19062 gnd.n3399 gnd.n3398 9.3005
R19063 gnd.n3397 gnd.n3392 9.3005
R19064 gnd.n3396 gnd.n3395 9.3005
R19065 gnd.n2495 gnd.n2494 9.3005
R19066 gnd.n3541 gnd.n3540 9.3005
R19067 gnd.n3542 gnd.n2492 9.3005
R19068 gnd.n3555 gnd.n3554 9.3005
R19069 gnd.n3553 gnd.n2493 9.3005
R19070 gnd.n3552 gnd.n3551 9.3005
R19071 gnd.n3550 gnd.n3543 9.3005
R19072 gnd.n3549 gnd.n3548 9.3005
R19073 gnd.n3547 gnd.n3546 9.3005
R19074 gnd.n2446 gnd.n2445 9.3005
R19075 gnd.n3617 gnd.n3616 9.3005
R19076 gnd.n3618 gnd.n2443 9.3005
R19077 gnd.n3621 gnd.n3620 9.3005
R19078 gnd.n3619 gnd.n2444 9.3005
R19079 gnd.n2419 gnd.n2418 9.3005
R19080 gnd.n3656 gnd.n3655 9.3005
R19081 gnd.n3657 gnd.n2417 9.3005
R19082 gnd.n3659 gnd.n3658 9.3005
R19083 gnd.n3660 gnd.n2416 9.3005
R19084 gnd.n3664 gnd.n3663 9.3005
R19085 gnd.n3665 gnd.n2414 9.3005
R19086 gnd.n3670 gnd.n3669 9.3005
R19087 gnd.n3668 gnd.n2415 9.3005
R19088 gnd.n3667 gnd.n3666 9.3005
R19089 gnd.n2360 gnd.n2359 9.3005
R19090 gnd.n3752 gnd.n3751 9.3005
R19091 gnd.n3753 gnd.n2357 9.3005
R19092 gnd.n3781 gnd.n3780 9.3005
R19093 gnd.n3779 gnd.n2358 9.3005
R19094 gnd.n3778 gnd.n3777 9.3005
R19095 gnd.n3776 gnd.n3754 9.3005
R19096 gnd.n3775 gnd.n3774 9.3005
R19097 gnd.n3773 gnd.n3760 9.3005
R19098 gnd.n3772 gnd.n3771 9.3005
R19099 gnd.n3770 gnd.n3761 9.3005
R19100 gnd.n3769 gnd.n3768 9.3005
R19101 gnd.n3767 gnd.n3764 9.3005
R19102 gnd.n3766 gnd.n3765 9.3005
R19103 gnd.n2287 gnd.n2286 9.3005
R19104 gnd.n3902 gnd.n3901 9.3005
R19105 gnd.n3903 gnd.n2284 9.3005
R19106 gnd.n3906 gnd.n3905 9.3005
R19107 gnd.n3904 gnd.n2285 9.3005
R19108 gnd.n2263 gnd.n2262 9.3005
R19109 gnd.n3935 gnd.n3934 9.3005
R19110 gnd.n3936 gnd.n2260 9.3005
R19111 gnd.n3964 gnd.n3963 9.3005
R19112 gnd.n3962 gnd.n2261 9.3005
R19113 gnd.n3961 gnd.n3960 9.3005
R19114 gnd.n3959 gnd.n3937 9.3005
R19115 gnd.n3958 gnd.n3957 9.3005
R19116 gnd.n3956 gnd.n3941 9.3005
R19117 gnd.n3955 gnd.n3954 9.3005
R19118 gnd.n3953 gnd.n3942 9.3005
R19119 gnd.n3952 gnd.n3951 9.3005
R19120 gnd.n3950 gnd.n3947 9.3005
R19121 gnd.n3949 gnd.n3948 9.3005
R19122 gnd.n2124 gnd.n2123 9.3005
R19123 gnd.n4169 gnd.n4168 9.3005
R19124 gnd.n4170 gnd.n2122 9.3005
R19125 gnd.n4172 gnd.n4171 9.3005
R19126 gnd.n2112 gnd.n2111 9.3005
R19127 gnd.n4188 gnd.n4187 9.3005
R19128 gnd.n4189 gnd.n2110 9.3005
R19129 gnd.n4191 gnd.n4190 9.3005
R19130 gnd.n1798 gnd.n1797 9.3005
R19131 gnd.n4567 gnd.n4566 9.3005
R19132 gnd.n3045 gnd.n3044 9.3005
R19133 gnd.n4563 gnd.n1799 9.3005
R19134 gnd.n4562 gnd.n4561 9.3005
R19135 gnd.n4560 gnd.n1802 9.3005
R19136 gnd.n4559 gnd.n4558 9.3005
R19137 gnd.n4557 gnd.n1803 9.3005
R19138 gnd.n4556 gnd.n4555 9.3005
R19139 gnd.n4565 gnd.n4564 9.3005
R19140 gnd.n4508 gnd.n4507 9.3005
R19141 gnd.n1850 gnd.n1849 9.3005
R19142 gnd.n4514 gnd.n4513 9.3005
R19143 gnd.n4516 gnd.n4515 9.3005
R19144 gnd.n1842 gnd.n1841 9.3005
R19145 gnd.n4522 gnd.n4521 9.3005
R19146 gnd.n4524 gnd.n4523 9.3005
R19147 gnd.n1834 gnd.n1833 9.3005
R19148 gnd.n4530 gnd.n4529 9.3005
R19149 gnd.n4532 gnd.n4531 9.3005
R19150 gnd.n1826 gnd.n1825 9.3005
R19151 gnd.n4538 gnd.n4537 9.3005
R19152 gnd.n4540 gnd.n4539 9.3005
R19153 gnd.n1818 gnd.n1817 9.3005
R19154 gnd.n4546 gnd.n4545 9.3005
R19155 gnd.n4548 gnd.n4547 9.3005
R19156 gnd.n1814 gnd.n1809 9.3005
R19157 gnd.n4506 gnd.n1859 9.3005
R19158 gnd.n2075 gnd.n1858 9.3005
R19159 gnd.n4553 gnd.n1807 9.3005
R19160 gnd.n4552 gnd.n4551 9.3005
R19161 gnd.n4550 gnd.n4549 9.3005
R19162 gnd.n1813 gnd.n1812 9.3005
R19163 gnd.n4544 gnd.n4543 9.3005
R19164 gnd.n4542 gnd.n4541 9.3005
R19165 gnd.n1822 gnd.n1821 9.3005
R19166 gnd.n4536 gnd.n4535 9.3005
R19167 gnd.n4534 gnd.n4533 9.3005
R19168 gnd.n1830 gnd.n1829 9.3005
R19169 gnd.n4528 gnd.n4527 9.3005
R19170 gnd.n4526 gnd.n4525 9.3005
R19171 gnd.n1838 gnd.n1837 9.3005
R19172 gnd.n4520 gnd.n4519 9.3005
R19173 gnd.n4518 gnd.n4517 9.3005
R19174 gnd.n1846 gnd.n1845 9.3005
R19175 gnd.n4512 gnd.n4511 9.3005
R19176 gnd.n4510 gnd.n4509 9.3005
R19177 gnd.n2098 gnd.n1856 9.3005
R19178 gnd.n2077 gnd.n2076 9.3005
R19179 gnd.n4256 gnd.n4255 9.3005
R19180 gnd.n4260 gnd.n4259 9.3005
R19181 gnd.n4261 gnd.n2072 9.3005
R19182 gnd.n4265 gnd.n4264 9.3005
R19183 gnd.n4266 gnd.n2071 9.3005
R19184 gnd.n4268 gnd.n4267 9.3005
R19185 gnd.n2069 gnd.n2068 9.3005
R19186 gnd.n4280 gnd.n4279 9.3005
R19187 gnd.n4281 gnd.n2067 9.3005
R19188 gnd.n4283 gnd.n4282 9.3005
R19189 gnd.n2065 gnd.n2064 9.3005
R19190 gnd.n4303 gnd.n4302 9.3005
R19191 gnd.n4304 gnd.n2062 9.3005
R19192 gnd.n4314 gnd.n4313 9.3005
R19193 gnd.n4312 gnd.n2063 9.3005
R19194 gnd.n4311 gnd.n4310 9.3005
R19195 gnd.n4309 gnd.n4305 9.3005
R19196 gnd.n4308 gnd.n4307 9.3005
R19197 gnd.n553 gnd.n552 9.3005
R19198 gnd.n7396 gnd.n7395 9.3005
R19199 gnd.n7397 gnd.n550 9.3005
R19200 gnd.n7400 gnd.n7399 9.3005
R19201 gnd.n7398 gnd.n551 9.3005
R19202 gnd.n524 gnd.n523 9.3005
R19203 gnd.n7433 gnd.n7432 9.3005
R19204 gnd.n7434 gnd.n522 9.3005
R19205 gnd.n7436 gnd.n7435 9.3005
R19206 gnd.n502 gnd.n501 9.3005
R19207 gnd.n7460 gnd.n7459 9.3005
R19208 gnd.n7461 gnd.n499 9.3005
R19209 gnd.n7463 gnd.n7462 9.3005
R19210 gnd.n500 gnd.n95 9.3005
R19211 gnd.n4258 gnd.n2073 9.3005
R19212 gnd.n7762 gnd.n96 9.3005
R19213 gnd.t122 gnd.n5229 9.24152
R19214 gnd.n5131 gnd.t393 9.24152
R19215 gnd.n6515 gnd.t368 9.24152
R19216 gnd.n4945 gnd.t137 9.24152
R19217 gnd.n4860 gnd.t10 9.24152
R19218 gnd.n4328 gnd.t74 9.24152
R19219 gnd.n7713 gnd.t27 9.24152
R19220 gnd.t186 gnd.t122 8.92286
R19221 gnd.t343 gnd.n2126 8.92286
R19222 gnd.n6384 gnd.n6359 8.92171
R19223 gnd.n6352 gnd.n6327 8.92171
R19224 gnd.n6320 gnd.n6295 8.92171
R19225 gnd.n6289 gnd.n6264 8.92171
R19226 gnd.n6257 gnd.n6232 8.92171
R19227 gnd.n6225 gnd.n6200 8.92171
R19228 gnd.n6193 gnd.n6168 8.92171
R19229 gnd.n6162 gnd.n6137 8.92171
R19230 gnd.n2160 gnd.n2142 8.72777
R19231 gnd.t129 gnd.n5358 8.60421
R19232 gnd.n4969 gnd.t51 8.60421
R19233 gnd.n4836 gnd.t2 8.60421
R19234 gnd.n4277 gnd.t60 8.60421
R19235 gnd.n7689 gnd.t189 8.60421
R19236 gnd.n5302 gnd.n5282 8.43656
R19237 gnd.n54 gnd.n34 8.43656
R19238 gnd.n3623 gnd.n2441 8.28555
R19239 gnd.n3673 gnd.n2380 8.28555
R19240 gnd.n3756 gnd.n2350 8.28555
R19241 gnd.n3848 gnd.n2299 8.28555
R19242 gnd.n6385 gnd.n6357 8.14595
R19243 gnd.n6353 gnd.n6325 8.14595
R19244 gnd.n6321 gnd.n6293 8.14595
R19245 gnd.n6290 gnd.n6262 8.14595
R19246 gnd.n6258 gnd.n6230 8.14595
R19247 gnd.n6226 gnd.n6198 8.14595
R19248 gnd.n6194 gnd.n6166 8.14595
R19249 gnd.n6163 gnd.n6135 8.14595
R19250 gnd.n2866 gnd.n0 8.10675
R19251 gnd.n7763 gnd.n7762 8.10675
R19252 gnd.n6390 gnd.n6389 7.97301
R19253 gnd.n5851 gnd.t131 7.9669
R19254 gnd.n7763 gnd.n94 7.95236
R19255 gnd.n4506 gnd.n1858 7.75808
R19256 gnd.n3321 gnd.n2579 7.75808
R19257 gnd.n445 gnd.n365 7.75808
R19258 gnd.n2800 gnd.n2799 7.75808
R19259 gnd.n6576 gnd.n6575 7.64824
R19260 gnd.n3472 gnd.t378 7.64824
R19261 gnd.t86 gnd.n2389 7.64824
R19262 gnd.n3702 gnd.t77 7.64824
R19263 gnd.n3802 gnd.t110 7.64824
R19264 gnd.n2335 gnd.t6 7.64824
R19265 gnd.n5343 gnd.n5342 7.53171
R19266 gnd.t119 gnd.n5444 7.32958
R19267 gnd.n3405 gnd.t150 7.32958
R19268 gnd.n4026 gnd.t261 7.32958
R19269 gnd.n1680 gnd.n1679 7.30353
R19270 gnd.n2159 gnd.n2158 7.30353
R19271 gnd.n5753 gnd.n5752 7.01093
R19272 gnd.n5763 gnd.n5473 7.01093
R19273 gnd.n5762 gnd.n5476 7.01093
R19274 gnd.n5771 gnd.n5467 7.01093
R19275 gnd.n5775 gnd.n5774 7.01093
R19276 gnd.n5793 gnd.n5452 7.01093
R19277 gnd.n5792 gnd.n5455 7.01093
R19278 gnd.n5803 gnd.n5444 7.01093
R19279 gnd.n5445 gnd.n5433 7.01093
R19280 gnd.n5816 gnd.n5434 7.01093
R19281 gnd.n5827 gnd.n5426 7.01093
R19282 gnd.n5826 gnd.n5417 7.01093
R19283 gnd.n5419 gnd.n5401 7.01093
R19284 gnd.n5863 gnd.n5402 7.01093
R19285 gnd.n5852 gnd.n5851 7.01093
R19286 gnd.n5888 gnd.n5393 7.01093
R19287 gnd.n5899 gnd.n5898 7.01093
R19288 gnd.n5386 gnd.n5378 7.01093
R19289 gnd.n5928 gnd.n5366 7.01093
R19290 gnd.n5927 gnd.n5369 7.01093
R19291 gnd.n5938 gnd.n5358 7.01093
R19292 gnd.n5359 gnd.n5347 7.01093
R19293 gnd.n5949 gnd.n5348 7.01093
R19294 gnd.n5970 gnd.n5259 7.01093
R19295 gnd.n5969 gnd.n5250 7.01093
R19296 gnd.n5252 gnd.n5243 7.01093
R19297 gnd.n5992 gnd.n5991 7.01093
R19298 gnd.n6011 gnd.n5229 7.01093
R19299 gnd.n6010 gnd.n5232 7.01093
R19300 gnd.n6021 gnd.n5221 7.01093
R19301 gnd.n6022 gnd.n5214 7.01093
R19302 gnd.n6037 gnd.n6036 7.01093
R19303 gnd.n6065 gnd.n5195 7.01093
R19304 gnd.n5196 gnd.n5184 7.01093
R19305 gnd.n6076 gnd.n5185 7.01093
R19306 gnd.n6101 gnd.n5176 7.01093
R19307 gnd.n6100 gnd.n5168 7.01093
R19308 gnd.n6112 gnd.n6111 7.01093
R19309 gnd.n6123 gnd.n6122 7.01093
R19310 gnd.n6397 gnd.n5149 7.01093
R19311 gnd.n6396 gnd.n5152 7.01093
R19312 gnd.n6410 gnd.n5141 7.01093
R19313 gnd.n5142 gnd.n5130 7.01093
R19314 gnd.n6421 gnd.n5131 7.01093
R19315 gnd.n6515 gnd.n5123 7.01093
R19316 gnd.n6514 gnd.n1118 7.01093
R19317 gnd.n6575 gnd.n1120 7.01093
R19318 gnd.n3487 gnd.n2520 7.01093
R19319 gnd.n3493 gnd.n3492 7.01093
R19320 gnd.n2436 gnd.n2435 7.01093
R19321 gnd.n2394 gnd.t86 7.01093
R19322 gnd.n3696 gnd.n2389 7.01093
R19323 gnd.n3808 gnd.n2335 7.01093
R19324 gnd.t6 gnd.n2334 7.01093
R19325 gnd.n3843 gnd.n2308 7.01093
R19326 gnd.n3858 gnd.n2241 7.01093
R19327 gnd.n3997 gnd.n2227 7.01093
R19328 gnd.n5434 gnd.t127 6.69227
R19329 gnd.n5991 gnd.t186 6.69227
R19330 gnd.t126 gnd.n5161 6.69227
R19331 gnd.n3292 gnd.t2 6.69227
R19332 gnd.n3565 gnd.t263 6.69227
R19333 gnd.t55 gnd.n3966 6.69227
R19334 gnd.t60 gnd.n2011 6.69227
R19335 gnd.n4086 gnd.n4085 6.5566
R19336 gnd.n3413 gnd.n3412 6.5566
R19337 gnd.n4697 gnd.n4693 6.5566
R19338 gnd.n4101 gnd.n4100 6.5566
R19339 gnd.t362 gnd.t349 6.37362
R19340 gnd.n3682 gnd.t92 6.37362
R19341 gnd.t79 gnd.n3826 6.37362
R19342 gnd.n4020 gnd.t283 6.37362
R19343 gnd.n3124 gnd.n3120 6.20656
R19344 gnd.n2098 gnd.n1855 6.20656
R19345 gnd.n5887 gnd.t89 6.05496
R19346 gnd.n5886 gnd.t121 6.05496
R19347 gnd.t279 gnd.n5359 6.05496
R19348 gnd.n6055 gnd.t133 6.05496
R19349 gnd.n2963 gnd.t10 6.05496
R19350 gnd.t8 gnd.t112 6.05496
R19351 gnd.t109 gnd.t80 6.05496
R19352 gnd.t74 gnd.n2052 6.05496
R19353 gnd.n6387 gnd.n6357 5.81868
R19354 gnd.n6355 gnd.n6325 5.81868
R19355 gnd.n6323 gnd.n6293 5.81868
R19356 gnd.n6292 gnd.n6262 5.81868
R19357 gnd.n6260 gnd.n6230 5.81868
R19358 gnd.n6228 gnd.n6198 5.81868
R19359 gnd.n6196 gnd.n6166 5.81868
R19360 gnd.n6165 gnd.n6135 5.81868
R19361 gnd.n3528 gnd.n2507 5.73631
R19362 gnd.n3509 gnd.n3508 5.73631
R19363 gnd.n3636 gnd.t107 5.73631
R19364 gnd.n3630 gnd.n2399 5.73631
R19365 gnd.n3681 gnd.n2393 5.73631
R19366 gnd.n3673 gnd.t77 5.73631
R19367 gnd.n3756 gnd.t110 5.73631
R19368 gnd.n3828 gnd.n2321 5.73631
R19369 gnd.n2324 gnd.n2312 5.73631
R19370 gnd.t7 gnd.n2315 5.73631
R19371 gnd.n3991 gnd.n2237 5.73631
R19372 gnd.n4004 gnd.n2231 5.73631
R19373 gnd.n2186 gnd.n1935 5.62001
R19374 gnd.n4759 gnd.n1622 5.62001
R19375 gnd.n4759 gnd.n1623 5.62001
R19376 gnd.n4095 gnd.n1935 5.62001
R19377 gnd.n5571 gnd.n5570 5.4308
R19378 gnd.n6496 gnd.n6428 5.4308
R19379 gnd.n5348 gnd.t132 5.41765
R19380 gnd.t123 gnd.n5980 5.41765
R19381 gnd.t218 gnd.n5205 5.41765
R19382 gnd.n2929 gnd.t105 5.41765
R19383 gnd.n2628 gnd.t0 5.41765
R19384 gnd.n3587 gnd.t168 5.41765
R19385 gnd.n3909 gnd.t402 5.41765
R19386 gnd.t58 gnd.n539 5.41765
R19387 gnd.t143 gnd.n520 5.41765
R19388 gnd.n3624 gnd.t54 5.09899
R19389 gnd.t115 gnd.n3887 5.09899
R19390 gnd.n6385 gnd.n6384 5.04292
R19391 gnd.n6353 gnd.n6352 5.04292
R19392 gnd.n6321 gnd.n6320 5.04292
R19393 gnd.n6290 gnd.n6289 5.04292
R19394 gnd.n6258 gnd.n6257 5.04292
R19395 gnd.n6226 gnd.n6225 5.04292
R19396 gnd.n6194 gnd.n6193 5.04292
R19397 gnd.n6163 gnd.n6162 5.04292
R19398 gnd.t124 gnd.n5909 4.78034
R19399 gnd.t130 gnd.n6021 4.78034
R19400 gnd.n2988 gnd.t18 4.78034
R19401 gnd.n2128 gnd.t323 4.78034
R19402 gnd.n7369 gnd.t14 4.78034
R19403 gnd.n5883 gnd.n5882 4.74817
R19404 gnd.n5878 gnd.n5877 4.74817
R19405 gnd.n5874 gnd.n5873 4.74817
R19406 gnd.n5870 gnd.n5345 4.74817
R19407 gnd.n5882 gnd.n5881 4.74817
R19408 gnd.n5880 gnd.n5878 4.74817
R19409 gnd.n5876 gnd.n5874 4.74817
R19410 gnd.n5872 gnd.n5870 4.74817
R19411 gnd.n7455 gnd.n113 4.74817
R19412 gnd.n7470 gnd.n112 4.74817
R19413 gnd.n7468 gnd.n111 4.74817
R19414 gnd.n7755 gnd.n106 4.74817
R19415 gnd.n7753 gnd.n107 4.74817
R19416 gnd.n508 gnd.n113 4.74817
R19417 gnd.n7454 gnd.n112 4.74817
R19418 gnd.n7471 gnd.n111 4.74817
R19419 gnd.n7467 gnd.n106 4.74817
R19420 gnd.n7754 gnd.n7753 4.74817
R19421 gnd.n1400 gnd.n1384 4.74817
R19422 gnd.n4900 gnd.n1401 4.74817
R19423 gnd.n2652 gnd.n1406 4.74817
R19424 gnd.n2889 gnd.n1405 4.74817
R19425 gnd.n1407 gnd.n1404 4.74817
R19426 gnd.n4911 gnd.n1384 4.74817
R19427 gnd.n4901 gnd.n4900 4.74817
R19428 gnd.n2724 gnd.n1406 4.74817
R19429 gnd.n2653 gnd.n1405 4.74817
R19430 gnd.n2888 gnd.n1404 4.74817
R19431 gnd.n5342 gnd.n5341 4.74296
R19432 gnd.n94 gnd.n93 4.74296
R19433 gnd.n5302 gnd.n5301 4.7074
R19434 gnd.n5322 gnd.n5321 4.7074
R19435 gnd.n54 gnd.n53 4.7074
R19436 gnd.n74 gnd.n73 4.7074
R19437 gnd.n5342 gnd.n5322 4.65959
R19438 gnd.n94 gnd.n74 4.65959
R19439 gnd.n4448 gnd.n1937 4.6132
R19440 gnd.n4760 gnd.n1621 4.6132
R19441 gnd.n4810 gnd.n1552 4.46168
R19442 gnd.n3516 gnd.n2514 4.46168
R19443 gnd.n3538 gnd.n2497 4.46168
R19444 gnd.t53 gnd.n2449 4.46168
R19445 gnd.n3653 gnd.n2422 4.46168
R19446 gnd.n3688 gnd.n2395 4.46168
R19447 gnd.n3820 gnd.n2328 4.46168
R19448 gnd.n3837 gnd.n3836 4.46168
R19449 gnd.n3880 gnd.t117 4.46168
R19450 gnd.n3984 gnd.n2244 4.46168
R19451 gnd.n4011 gnd.n2223 4.46168
R19452 gnd.n4501 gnd.n1903 4.46168
R19453 gnd.n2155 gnd.n2142 4.46111
R19454 gnd.n6370 gnd.n6366 4.38594
R19455 gnd.n6338 gnd.n6334 4.38594
R19456 gnd.n6306 gnd.n6302 4.38594
R19457 gnd.n6275 gnd.n6271 4.38594
R19458 gnd.n6243 gnd.n6239 4.38594
R19459 gnd.n6211 gnd.n6207 4.38594
R19460 gnd.n6179 gnd.n6175 4.38594
R19461 gnd.n6148 gnd.n6144 4.38594
R19462 gnd.n6381 gnd.n6359 4.26717
R19463 gnd.n6349 gnd.n6327 4.26717
R19464 gnd.n6317 gnd.n6295 4.26717
R19465 gnd.n6286 gnd.n6264 4.26717
R19466 gnd.n6254 gnd.n6232 4.26717
R19467 gnd.n6222 gnd.n6200 4.26717
R19468 gnd.n6190 gnd.n6168 4.26717
R19469 gnd.n6159 gnd.n6137 4.26717
R19470 gnd.t125 gnd.n5840 4.14303
R19471 gnd.n6101 gnd.t128 4.14303
R19472 gnd.n3010 gnd.t69 4.14303
R19473 gnd.t184 gnd.n2029 4.14303
R19474 gnd.n6389 gnd.n6388 4.08274
R19475 gnd.n4085 gnd.n4084 4.05904
R19476 gnd.n3414 gnd.n3413 4.05904
R19477 gnd.n4700 gnd.n4693 4.05904
R19478 gnd.n4102 gnd.n4101 4.05904
R19479 gnd.n15 gnd.n7 3.99943
R19480 gnd.n3603 gnd.t114 3.82437
R19481 gnd.n3739 gnd.t112 3.82437
R19482 gnd.n3783 gnd.t109 3.82437
R19483 gnd.t113 gnd.n2273 3.82437
R19484 gnd.n5344 gnd.n5343 3.81325
R19485 gnd.n5322 gnd.n5302 3.72967
R19486 gnd.n74 gnd.n54 3.72967
R19487 gnd.n6389 gnd.n6261 3.70378
R19488 gnd.n15 gnd.n14 3.60163
R19489 gnd.n1270 gnd.t297 3.50571
R19490 gnd.n3278 gnd.t312 3.50571
R19491 gnd.n4372 gnd.t293 3.50571
R19492 gnd.t308 gnd.n235 3.50571
R19493 gnd.n6380 gnd.n6361 3.49141
R19494 gnd.n6348 gnd.n6329 3.49141
R19495 gnd.n6316 gnd.n6297 3.49141
R19496 gnd.n6285 gnd.n6266 3.49141
R19497 gnd.n6253 gnd.n6234 3.49141
R19498 gnd.n6221 gnd.n6202 3.49141
R19499 gnd.n6189 gnd.n6170 3.49141
R19500 gnd.n6158 gnd.n6139 3.49141
R19501 gnd.n4466 gnd.n4465 3.29747
R19502 gnd.n4465 gnd.n4464 3.29747
R19503 gnd.n7630 gnd.n7627 3.29747
R19504 gnd.n7631 gnd.n7630 3.29747
R19505 gnd.n5076 gnd.n5075 3.29747
R19506 gnd.n5075 gnd.n5074 3.29747
R19507 gnd.n4778 gnd.n4777 3.29747
R19508 gnd.n4777 gnd.n4776 3.29747
R19509 gnd.n4679 gnd.n1698 3.18706
R19510 gnd.n3528 gnd.t353 3.18706
R19511 gnd.n3558 gnd.n3557 3.18706
R19512 gnd.n2478 gnd.t111 3.18706
R19513 gnd.n3644 gnd.n3642 3.18706
R19514 gnd.n3695 gnd.n2385 3.18706
R19515 gnd.n3801 gnd.n2333 3.18706
R19516 gnd.n3889 gnd.n2296 3.18706
R19517 gnd.t78 gnd.n2265 3.18706
R19518 gnd.n3974 gnd.n3973 3.18706
R19519 gnd.n4020 gnd.n4019 3.18706
R19520 gnd.n4026 gnd.t397 3.18706
R19521 gnd.n5841 gnd.t125 2.8684
R19522 gnd.n3527 gnd.t87 2.8684
R19523 gnd.t71 gnd.n2236 2.8684
R19524 gnd.n5323 gnd.t234 2.82907
R19525 gnd.n5323 gnd.t70 2.82907
R19526 gnd.n5325 gnd.t147 2.82907
R19527 gnd.n5325 gnd.t98 2.82907
R19528 gnd.n5327 gnd.t34 2.82907
R19529 gnd.n5327 gnd.t104 2.82907
R19530 gnd.n5329 gnd.t166 2.82907
R19531 gnd.n5329 gnd.t106 2.82907
R19532 gnd.n5331 gnd.t269 2.82907
R19533 gnd.n5331 gnd.t258 2.82907
R19534 gnd.n5333 gnd.t220 2.82907
R19535 gnd.n5333 gnd.t206 2.82907
R19536 gnd.n5335 gnd.t257 2.82907
R19537 gnd.n5335 gnd.t259 2.82907
R19538 gnd.n5337 gnd.t216 2.82907
R19539 gnd.n5337 gnd.t281 2.82907
R19540 gnd.n5339 gnd.t167 2.82907
R19541 gnd.n5339 gnd.t48 2.82907
R19542 gnd.n5264 gnd.t21 2.82907
R19543 gnd.n5264 gnd.t177 2.82907
R19544 gnd.n5266 gnd.t26 2.82907
R19545 gnd.n5266 gnd.t249 2.82907
R19546 gnd.n5268 gnd.t1 2.82907
R19547 gnd.n5268 gnd.t191 2.82907
R19548 gnd.n5270 gnd.t182 2.82907
R19549 gnd.n5270 gnd.t180 2.82907
R19550 gnd.n5272 gnd.t274 2.82907
R19551 gnd.n5272 gnd.t157 2.82907
R19552 gnd.n5274 gnd.t194 2.82907
R19553 gnd.n5274 gnd.t247 2.82907
R19554 gnd.n5276 gnd.t73 2.82907
R19555 gnd.n5276 gnd.t23 2.82907
R19556 gnd.n5278 gnd.t138 2.82907
R19557 gnd.n5278 gnd.t5 2.82907
R19558 gnd.n5280 gnd.t145 2.82907
R19559 gnd.n5280 gnd.t266 2.82907
R19560 gnd.n5283 gnd.t159 2.82907
R19561 gnd.n5283 gnd.t82 2.82907
R19562 gnd.n5285 gnd.t154 2.82907
R19563 gnd.n5285 gnd.t11 2.82907
R19564 gnd.n5287 gnd.t199 2.82907
R19565 gnd.n5287 gnd.t146 2.82907
R19566 gnd.n5289 gnd.t204 2.82907
R19567 gnd.n5289 gnd.t134 2.82907
R19568 gnd.n5291 gnd.t255 2.82907
R19569 gnd.n5291 gnd.t178 2.82907
R19570 gnd.n5293 gnd.t276 2.82907
R19571 gnd.n5293 gnd.t195 2.82907
R19572 gnd.n5295 gnd.t68 2.82907
R19573 gnd.n5295 gnd.t66 2.82907
R19574 gnd.n5297 gnd.t238 2.82907
R19575 gnd.n5297 gnd.t253 2.82907
R19576 gnd.n5299 gnd.t162 2.82907
R19577 gnd.n5299 gnd.t192 2.82907
R19578 gnd.n5303 gnd.t62 2.82907
R19579 gnd.n5303 gnd.t155 2.82907
R19580 gnd.n5305 gnd.t19 2.82907
R19581 gnd.n5305 gnd.t193 2.82907
R19582 gnd.n5307 gnd.t31 2.82907
R19583 gnd.n5307 gnd.t179 2.82907
R19584 gnd.n5309 gnd.t226 2.82907
R19585 gnd.n5309 gnd.t236 2.82907
R19586 gnd.n5311 gnd.t140 2.82907
R19587 gnd.n5311 gnd.t13 2.82907
R19588 gnd.n5313 gnd.t40 2.82907
R19589 gnd.n5313 gnd.t173 2.82907
R19590 gnd.n5315 gnd.t250 2.82907
R19591 gnd.n5315 gnd.t158 2.82907
R19592 gnd.n5317 gnd.t222 2.82907
R19593 gnd.n5317 gnd.t198 2.82907
R19594 gnd.n5319 gnd.t17 2.82907
R19595 gnd.n5319 gnd.t212 2.82907
R19596 gnd.n91 gnd.t160 2.82907
R19597 gnd.n91 gnd.t57 2.82907
R19598 gnd.n89 gnd.t221 2.82907
R19599 gnd.n89 gnd.t76 2.82907
R19600 gnd.n87 gnd.t407 2.82907
R19601 gnd.n87 gnd.t217 2.82907
R19602 gnd.n85 gnd.t46 2.82907
R19603 gnd.n85 gnd.t406 2.82907
R19604 gnd.n83 gnd.t241 2.82907
R19605 gnd.n83 gnd.t188 2.82907
R19606 gnd.n81 gnd.t144 2.82907
R19607 gnd.n81 gnd.t36 2.82907
R19608 gnd.n79 gnd.t213 2.82907
R19609 gnd.n79 gnd.t59 2.82907
R19610 gnd.n77 gnd.t161 2.82907
R19611 gnd.n77 gnd.t183 2.82907
R19612 gnd.n75 gnd.t185 2.82907
R19613 gnd.n75 gnd.t38 2.82907
R19614 gnd.n32 gnd.t44 2.82907
R19615 gnd.n32 gnd.t83 2.82907
R19616 gnd.n30 gnd.t211 2.82907
R19617 gnd.n30 gnd.t170 2.82907
R19618 gnd.n28 gnd.t202 2.82907
R19619 gnd.n28 gnd.t176 2.82907
R19620 gnd.n26 gnd.t175 2.82907
R19621 gnd.n26 gnd.t273 2.82907
R19622 gnd.n24 gnd.t142 2.82907
R19623 gnd.n24 gnd.t174 2.82907
R19624 gnd.n22 gnd.t210 2.82907
R19625 gnd.n22 gnd.t42 2.82907
R19626 gnd.n20 gnd.t201 2.82907
R19627 gnd.n20 gnd.t214 2.82907
R19628 gnd.n18 gnd.t156 2.82907
R19629 gnd.n18 gnd.t171 2.82907
R19630 gnd.n16 gnd.t203 2.82907
R19631 gnd.n16 gnd.t251 2.82907
R19632 gnd.n51 gnd.t267 2.82907
R19633 gnd.n51 gnd.t97 2.82907
R19634 gnd.n49 gnd.t136 2.82907
R19635 gnd.n49 gnd.t233 2.82907
R19636 gnd.n47 gnd.t25 2.82907
R19637 gnd.n47 gnd.t237 2.82907
R19638 gnd.n45 gnd.t200 2.82907
R19639 gnd.n45 gnd.t197 2.82907
R19640 gnd.n43 gnd.t232 2.82907
R19641 gnd.n43 gnd.t215 2.82907
R19642 gnd.n41 gnd.t246 2.82907
R19643 gnd.n41 gnd.t65 2.82907
R19644 gnd.n39 gnd.t30 2.82907
R19645 gnd.n39 gnd.t278 2.82907
R19646 gnd.n37 gnd.t181 2.82907
R19647 gnd.n37 gnd.t209 2.82907
R19648 gnd.n35 gnd.t272 2.82907
R19649 gnd.n35 gnd.t248 2.82907
R19650 gnd.n71 gnd.t254 2.82907
R19651 gnd.n71 gnd.t33 2.82907
R19652 gnd.n69 gnd.t275 2.82907
R19653 gnd.n69 gnd.t28 2.82907
R19654 gnd.n67 gnd.t223 2.82907
R19655 gnd.n67 gnd.t102 2.82907
R19656 gnd.n65 gnd.t225 2.82907
R19657 gnd.n65 gnd.t265 2.82907
R19658 gnd.n63 gnd.t256 2.82907
R19659 gnd.n63 gnd.t64 2.82907
R19660 gnd.n61 gnd.t240 2.82907
R19661 gnd.n61 gnd.t245 2.82907
R19662 gnd.n59 gnd.t41 2.82907
R19663 gnd.n59 gnd.t252 2.82907
R19664 gnd.n57 gnd.t75 2.82907
R19665 gnd.n57 gnd.t15 2.82907
R19666 gnd.n55 gnd.t239 2.82907
R19667 gnd.n55 gnd.t404 2.82907
R19668 gnd.n6377 gnd.n6376 2.71565
R19669 gnd.n6345 gnd.n6344 2.71565
R19670 gnd.n6313 gnd.n6312 2.71565
R19671 gnd.n6282 gnd.n6281 2.71565
R19672 gnd.n6250 gnd.n6249 2.71565
R19673 gnd.n6218 gnd.n6217 2.71565
R19674 gnd.n6186 gnd.n6185 2.71565
R19675 gnd.n6155 gnd.n6154 2.71565
R19676 gnd.n3564 gnd.t100 2.54975
R19677 gnd.n3967 gnd.t99 2.54975
R19678 gnd.n5882 gnd.n5344 2.27742
R19679 gnd.n5878 gnd.n5344 2.27742
R19680 gnd.n5874 gnd.n5344 2.27742
R19681 gnd.n5870 gnd.n5344 2.27742
R19682 gnd.n7752 gnd.n113 2.27742
R19683 gnd.n7752 gnd.n112 2.27742
R19684 gnd.n7752 gnd.n111 2.27742
R19685 gnd.n7752 gnd.n106 2.27742
R19686 gnd.n7753 gnd.n7752 2.27742
R19687 gnd.n4899 gnd.n1384 2.27742
R19688 gnd.n4900 gnd.n4899 2.27742
R19689 gnd.n4899 gnd.n1406 2.27742
R19690 gnd.n4899 gnd.n1405 2.27742
R19691 gnd.n4899 gnd.n1404 2.27742
R19692 gnd.t332 gnd.n5762 2.23109
R19693 gnd.n5910 gnd.t124 2.23109
R19694 gnd.n2395 gnd.t93 2.23109
R19695 gnd.n3725 gnd.t8 2.23109
R19696 gnd.t80 gnd.n2347 2.23109
R19697 gnd.t152 gnd.n2328 2.23109
R19698 gnd.n7337 gnd.t32 2.23109
R19699 gnd.n6373 gnd.n6363 1.93989
R19700 gnd.n6341 gnd.n6331 1.93989
R19701 gnd.n6309 gnd.n6299 1.93989
R19702 gnd.n6278 gnd.n6268 1.93989
R19703 gnd.n6246 gnd.n6236 1.93989
R19704 gnd.n6214 gnd.n6204 1.93989
R19705 gnd.n6182 gnd.n6172 1.93989
R19706 gnd.n6151 gnd.n6141 1.93989
R19707 gnd.n4685 gnd.n1687 1.91244
R19708 gnd.t290 gnd.n1687 1.91244
R19709 gnd.n3493 gnd.t85 1.91244
R19710 gnd.n3497 gnd.n2475 1.91244
R19711 gnd.n3595 gnd.n2466 1.91244
R19712 gnd.n3727 gnd.n3726 1.91244
R19713 gnd.n3791 gnd.n3790 1.91244
R19714 gnd.n3899 gnd.n2289 1.91244
R19715 gnd.n3855 gnd.n3854 1.91244
R19716 gnd.n3858 gnd.t91 1.91244
R19717 gnd.n4158 gnd.n2134 1.91244
R19718 gnd.n5775 gnd.t270 1.59378
R19719 gnd.n5981 gnd.t123 1.59378
R19720 gnd.n6054 gnd.t218 1.59378
R19721 gnd.t47 gnd.n1314 1.59378
R19722 gnd.n2973 gnd.t20 1.59378
R19723 gnd.t263 gnd.n3564 1.59378
R19724 gnd.n3967 gnd.t55 1.59378
R19725 gnd.n4342 gnd.t37 1.59378
R19726 gnd.n194 gnd.t43 1.59378
R19727 gnd.n3509 gnd.t108 1.27512
R19728 gnd.n3991 gnd.t116 1.27512
R19729 gnd.n4011 gnd.t301 1.27512
R19730 gnd.n5572 gnd.n5571 1.16414
R19731 gnd.n6499 gnd.n6496 1.16414
R19732 gnd.n6372 gnd.n6365 1.16414
R19733 gnd.n6340 gnd.n6333 1.16414
R19734 gnd.n6308 gnd.n6301 1.16414
R19735 gnd.n6277 gnd.n6270 1.16414
R19736 gnd.n6245 gnd.n6238 1.16414
R19737 gnd.n6213 gnd.n6206 1.16414
R19738 gnd.n6181 gnd.n6174 1.16414
R19739 gnd.n6150 gnd.n6143 1.16414
R19740 gnd.n4448 gnd.n4447 0.970197
R19741 gnd.n4760 gnd.n1619 0.970197
R19742 gnd.n6356 gnd.n6324 0.962709
R19743 gnd.n6388 gnd.n6356 0.962709
R19744 gnd.n6229 gnd.n6197 0.962709
R19745 gnd.n6261 gnd.n6229 0.962709
R19746 gnd.t89 gnd.n5886 0.956468
R19747 gnd.n6035 gnd.t133 0.956468
R19748 gnd.t67 gnd.n1352 0.956468
R19749 gnd.n2952 gnd.t103 0.956468
R19750 gnd.t150 gnd.n3404 0.956468
R19751 gnd.n3945 gnd.t261 0.956468
R19752 gnd.n7376 gnd.t29 0.956468
R19753 gnd.n156 gnd.t101 0.956468
R19754 gnd.n2 gnd.n1 0.672012
R19755 gnd.n3 gnd.n2 0.672012
R19756 gnd.n4 gnd.n3 0.672012
R19757 gnd.n5 gnd.n4 0.672012
R19758 gnd.n6 gnd.n5 0.672012
R19759 gnd.n7 gnd.n6 0.672012
R19760 gnd.n9 gnd.n8 0.672012
R19761 gnd.n10 gnd.n9 0.672012
R19762 gnd.n11 gnd.n10 0.672012
R19763 gnd.n12 gnd.n11 0.672012
R19764 gnd.n13 gnd.n12 0.672012
R19765 gnd.n14 gnd.n13 0.672012
R19766 gnd.n4679 gnd.t349 0.637812
R19767 gnd.t329 gnd.n2519 0.637812
R19768 gnd.n3580 gnd.n2470 0.637812
R19769 gnd.n3588 gnd.n3587 0.637812
R19770 gnd.n2375 gnd.n2374 0.637812
R19771 gnd.n2366 gnd.n2354 0.637812
R19772 gnd.n3910 gnd.n3909 0.637812
R19773 gnd.n3869 gnd.n2276 0.637812
R19774 gnd.n4019 gnd.t304 0.637812
R19775 gnd.n2138 gnd.t343 0.637812
R19776 gnd.n7764 gnd.n7763 0.63688
R19777 gnd gnd.n0 0.634843
R19778 gnd.n5341 gnd.n5340 0.573776
R19779 gnd.n5340 gnd.n5338 0.573776
R19780 gnd.n5338 gnd.n5336 0.573776
R19781 gnd.n5336 gnd.n5334 0.573776
R19782 gnd.n5334 gnd.n5332 0.573776
R19783 gnd.n5332 gnd.n5330 0.573776
R19784 gnd.n5330 gnd.n5328 0.573776
R19785 gnd.n5328 gnd.n5326 0.573776
R19786 gnd.n5326 gnd.n5324 0.573776
R19787 gnd.n5282 gnd.n5281 0.573776
R19788 gnd.n5281 gnd.n5279 0.573776
R19789 gnd.n5279 gnd.n5277 0.573776
R19790 gnd.n5277 gnd.n5275 0.573776
R19791 gnd.n5275 gnd.n5273 0.573776
R19792 gnd.n5273 gnd.n5271 0.573776
R19793 gnd.n5271 gnd.n5269 0.573776
R19794 gnd.n5269 gnd.n5267 0.573776
R19795 gnd.n5267 gnd.n5265 0.573776
R19796 gnd.n5301 gnd.n5300 0.573776
R19797 gnd.n5300 gnd.n5298 0.573776
R19798 gnd.n5298 gnd.n5296 0.573776
R19799 gnd.n5296 gnd.n5294 0.573776
R19800 gnd.n5294 gnd.n5292 0.573776
R19801 gnd.n5292 gnd.n5290 0.573776
R19802 gnd.n5290 gnd.n5288 0.573776
R19803 gnd.n5288 gnd.n5286 0.573776
R19804 gnd.n5286 gnd.n5284 0.573776
R19805 gnd.n5321 gnd.n5320 0.573776
R19806 gnd.n5320 gnd.n5318 0.573776
R19807 gnd.n5318 gnd.n5316 0.573776
R19808 gnd.n5316 gnd.n5314 0.573776
R19809 gnd.n5314 gnd.n5312 0.573776
R19810 gnd.n5312 gnd.n5310 0.573776
R19811 gnd.n5310 gnd.n5308 0.573776
R19812 gnd.n5308 gnd.n5306 0.573776
R19813 gnd.n5306 gnd.n5304 0.573776
R19814 gnd.n78 gnd.n76 0.573776
R19815 gnd.n80 gnd.n78 0.573776
R19816 gnd.n82 gnd.n80 0.573776
R19817 gnd.n84 gnd.n82 0.573776
R19818 gnd.n86 gnd.n84 0.573776
R19819 gnd.n88 gnd.n86 0.573776
R19820 gnd.n90 gnd.n88 0.573776
R19821 gnd.n92 gnd.n90 0.573776
R19822 gnd.n93 gnd.n92 0.573776
R19823 gnd.n19 gnd.n17 0.573776
R19824 gnd.n21 gnd.n19 0.573776
R19825 gnd.n23 gnd.n21 0.573776
R19826 gnd.n25 gnd.n23 0.573776
R19827 gnd.n27 gnd.n25 0.573776
R19828 gnd.n29 gnd.n27 0.573776
R19829 gnd.n31 gnd.n29 0.573776
R19830 gnd.n33 gnd.n31 0.573776
R19831 gnd.n34 gnd.n33 0.573776
R19832 gnd.n38 gnd.n36 0.573776
R19833 gnd.n40 gnd.n38 0.573776
R19834 gnd.n42 gnd.n40 0.573776
R19835 gnd.n44 gnd.n42 0.573776
R19836 gnd.n46 gnd.n44 0.573776
R19837 gnd.n48 gnd.n46 0.573776
R19838 gnd.n50 gnd.n48 0.573776
R19839 gnd.n52 gnd.n50 0.573776
R19840 gnd.n53 gnd.n52 0.573776
R19841 gnd.n58 gnd.n56 0.573776
R19842 gnd.n60 gnd.n58 0.573776
R19843 gnd.n62 gnd.n60 0.573776
R19844 gnd.n64 gnd.n62 0.573776
R19845 gnd.n66 gnd.n64 0.573776
R19846 gnd.n68 gnd.n66 0.573776
R19847 gnd.n70 gnd.n68 0.573776
R19848 gnd.n72 gnd.n70 0.573776
R19849 gnd.n73 gnd.n72 0.573776
R19850 gnd.n4572 gnd.n1789 0.489829
R19851 gnd.n3325 gnd.n2548 0.489829
R19852 gnd.n3044 gnd.n3036 0.489829
R19853 gnd.n4566 gnd.n4565 0.489829
R19854 gnd.n6510 gnd.n6509 0.486781
R19855 gnd.n5624 gnd.n5520 0.48678
R19856 gnd.n6521 gnd.n6520 0.480683
R19857 gnd.n5692 gnd.n5470 0.480683
R19858 gnd.n443 gnd.n442 0.477634
R19859 gnd.n2802 gnd.n2801 0.477634
R19860 gnd.n953 gnd.n948 0.459342
R19861 gnd.n7132 gnd.n7131 0.459342
R19862 gnd.n7345 gnd.n7344 0.459342
R19863 gnd.n2657 gnd.n2656 0.459342
R19864 gnd.n7667 gnd.n7666 0.442573
R19865 gnd.n1988 gnd.n1907 0.442573
R19866 gnd.n4814 gnd.n4813 0.442573
R19867 gnd.n1264 gnd.n1190 0.442573
R19868 gnd.n7752 gnd.n110 0.420375
R19869 gnd.n4899 gnd.n1403 0.420375
R19870 gnd.n3120 gnd.n3111 0.388379
R19871 gnd.n6369 gnd.n6368 0.388379
R19872 gnd.n6337 gnd.n6336 0.388379
R19873 gnd.n6305 gnd.n6304 0.388379
R19874 gnd.n6274 gnd.n6273 0.388379
R19875 gnd.n6242 gnd.n6241 0.388379
R19876 gnd.n6210 gnd.n6209 0.388379
R19877 gnd.n6178 gnd.n6177 0.388379
R19878 gnd.n6147 gnd.n6146 0.388379
R19879 gnd.n4510 gnd.n1855 0.388379
R19880 gnd.n7764 gnd.n15 0.374463
R19881 gnd.n6094 gnd.t126 0.319156
R19882 gnd.t172 gnd.n1389 0.319156
R19883 gnd.t165 gnd.n2899 0.319156
R19884 gnd.n7457 gnd.t35 0.319156
R19885 gnd.n117 gnd.t45 0.319156
R19886 gnd.n5618 gnd.n5617 0.311721
R19887 gnd gnd.n7764 0.295112
R19888 gnd.n7543 gnd.n479 0.293183
R19889 gnd.n4992 gnd.n1254 0.293183
R19890 gnd.n6566 gnd.n1125 0.268793
R19891 gnd.n7544 gnd.n7543 0.258122
R19892 gnd.n4386 gnd.n1808 0.258122
R19893 gnd.n3272 gnd.n3271 0.258122
R19894 gnd.n4993 gnd.n4992 0.258122
R19895 gnd.n3324 gnd.n2575 0.247451
R19896 gnd.n4258 gnd.n4257 0.247451
R19897 gnd.n6440 gnd.n1125 0.241354
R19898 gnd.n1937 gnd.n1934 0.229039
R19899 gnd.n1938 gnd.n1937 0.229039
R19900 gnd.n1621 gnd.n1618 0.229039
R19901 gnd.n3196 gnd.n1621 0.229039
R19902 gnd.n5343 gnd.n0 0.210825
R19903 gnd.n5747 gnd.n5488 0.206293
R19904 gnd.n6386 gnd.n6358 0.155672
R19905 gnd.n6379 gnd.n6358 0.155672
R19906 gnd.n6379 gnd.n6378 0.155672
R19907 gnd.n6378 gnd.n6362 0.155672
R19908 gnd.n6371 gnd.n6362 0.155672
R19909 gnd.n6371 gnd.n6370 0.155672
R19910 gnd.n6354 gnd.n6326 0.155672
R19911 gnd.n6347 gnd.n6326 0.155672
R19912 gnd.n6347 gnd.n6346 0.155672
R19913 gnd.n6346 gnd.n6330 0.155672
R19914 gnd.n6339 gnd.n6330 0.155672
R19915 gnd.n6339 gnd.n6338 0.155672
R19916 gnd.n6322 gnd.n6294 0.155672
R19917 gnd.n6315 gnd.n6294 0.155672
R19918 gnd.n6315 gnd.n6314 0.155672
R19919 gnd.n6314 gnd.n6298 0.155672
R19920 gnd.n6307 gnd.n6298 0.155672
R19921 gnd.n6307 gnd.n6306 0.155672
R19922 gnd.n6291 gnd.n6263 0.155672
R19923 gnd.n6284 gnd.n6263 0.155672
R19924 gnd.n6284 gnd.n6283 0.155672
R19925 gnd.n6283 gnd.n6267 0.155672
R19926 gnd.n6276 gnd.n6267 0.155672
R19927 gnd.n6276 gnd.n6275 0.155672
R19928 gnd.n6259 gnd.n6231 0.155672
R19929 gnd.n6252 gnd.n6231 0.155672
R19930 gnd.n6252 gnd.n6251 0.155672
R19931 gnd.n6251 gnd.n6235 0.155672
R19932 gnd.n6244 gnd.n6235 0.155672
R19933 gnd.n6244 gnd.n6243 0.155672
R19934 gnd.n6227 gnd.n6199 0.155672
R19935 gnd.n6220 gnd.n6199 0.155672
R19936 gnd.n6220 gnd.n6219 0.155672
R19937 gnd.n6219 gnd.n6203 0.155672
R19938 gnd.n6212 gnd.n6203 0.155672
R19939 gnd.n6212 gnd.n6211 0.155672
R19940 gnd.n6195 gnd.n6167 0.155672
R19941 gnd.n6188 gnd.n6167 0.155672
R19942 gnd.n6188 gnd.n6187 0.155672
R19943 gnd.n6187 gnd.n6171 0.155672
R19944 gnd.n6180 gnd.n6171 0.155672
R19945 gnd.n6180 gnd.n6179 0.155672
R19946 gnd.n6164 gnd.n6136 0.155672
R19947 gnd.n6157 gnd.n6136 0.155672
R19948 gnd.n6157 gnd.n6156 0.155672
R19949 gnd.n6156 gnd.n6140 0.155672
R19950 gnd.n6149 gnd.n6140 0.155672
R19951 gnd.n6149 gnd.n6148 0.155672
R19952 gnd.n6555 gnd.n6521 0.152939
R19953 gnd.n6555 gnd.n6554 0.152939
R19954 gnd.n6554 gnd.n6553 0.152939
R19955 gnd.n6553 gnd.n6523 0.152939
R19956 gnd.n6524 gnd.n6523 0.152939
R19957 gnd.n6525 gnd.n6524 0.152939
R19958 gnd.n6526 gnd.n6525 0.152939
R19959 gnd.n6527 gnd.n6526 0.152939
R19960 gnd.n6528 gnd.n6527 0.152939
R19961 gnd.n6529 gnd.n6528 0.152939
R19962 gnd.n6530 gnd.n6529 0.152939
R19963 gnd.n6531 gnd.n6530 0.152939
R19964 gnd.n6531 gnd.n1132 0.152939
R19965 gnd.n6564 gnd.n1132 0.152939
R19966 gnd.n6565 gnd.n6564 0.152939
R19967 gnd.n6566 gnd.n6565 0.152939
R19968 gnd.n5766 gnd.n5470 0.152939
R19969 gnd.n5767 gnd.n5766 0.152939
R19970 gnd.n5768 gnd.n5767 0.152939
R19971 gnd.n5768 gnd.n5449 0.152939
R19972 gnd.n5796 gnd.n5449 0.152939
R19973 gnd.n5797 gnd.n5796 0.152939
R19974 gnd.n5798 gnd.n5797 0.152939
R19975 gnd.n5799 gnd.n5798 0.152939
R19976 gnd.n5799 gnd.n5423 0.152939
R19977 gnd.n5830 gnd.n5423 0.152939
R19978 gnd.n5831 gnd.n5830 0.152939
R19979 gnd.n5832 gnd.n5831 0.152939
R19980 gnd.n5833 gnd.n5832 0.152939
R19981 gnd.n5834 gnd.n5833 0.152939
R19982 gnd.n5834 gnd.n5390 0.152939
R19983 gnd.n5891 gnd.n5390 0.152939
R19984 gnd.n5892 gnd.n5891 0.152939
R19985 gnd.n5893 gnd.n5892 0.152939
R19986 gnd.n5894 gnd.n5893 0.152939
R19987 gnd.n5894 gnd.n5363 0.152939
R19988 gnd.n5931 gnd.n5363 0.152939
R19989 gnd.n5932 gnd.n5931 0.152939
R19990 gnd.n5933 gnd.n5932 0.152939
R19991 gnd.n5934 gnd.n5933 0.152939
R19992 gnd.n5934 gnd.n5256 0.152939
R19993 gnd.n5973 gnd.n5256 0.152939
R19994 gnd.n5974 gnd.n5973 0.152939
R19995 gnd.n5975 gnd.n5974 0.152939
R19996 gnd.n5976 gnd.n5975 0.152939
R19997 gnd.n5976 gnd.n5226 0.152939
R19998 gnd.n6014 gnd.n5226 0.152939
R19999 gnd.n6015 gnd.n6014 0.152939
R20000 gnd.n6016 gnd.n6015 0.152939
R20001 gnd.n6017 gnd.n6016 0.152939
R20002 gnd.n6017 gnd.n5200 0.152939
R20003 gnd.n6058 gnd.n5200 0.152939
R20004 gnd.n6059 gnd.n6058 0.152939
R20005 gnd.n6060 gnd.n6059 0.152939
R20006 gnd.n6061 gnd.n6060 0.152939
R20007 gnd.n6061 gnd.n5173 0.152939
R20008 gnd.n6104 gnd.n5173 0.152939
R20009 gnd.n6105 gnd.n6104 0.152939
R20010 gnd.n6106 gnd.n6105 0.152939
R20011 gnd.n6107 gnd.n6106 0.152939
R20012 gnd.n6107 gnd.n5146 0.152939
R20013 gnd.n6400 gnd.n5146 0.152939
R20014 gnd.n6401 gnd.n6400 0.152939
R20015 gnd.n6402 gnd.n6401 0.152939
R20016 gnd.n6403 gnd.n6402 0.152939
R20017 gnd.n6405 gnd.n6403 0.152939
R20018 gnd.n6405 gnd.n6404 0.152939
R20019 gnd.n6404 gnd.n5120 0.152939
R20020 gnd.n6520 gnd.n5120 0.152939
R20021 gnd.n5693 gnd.n5692 0.152939
R20022 gnd.n5694 gnd.n5693 0.152939
R20023 gnd.n5695 gnd.n5694 0.152939
R20024 gnd.n5696 gnd.n5695 0.152939
R20025 gnd.n5697 gnd.n5696 0.152939
R20026 gnd.n5698 gnd.n5697 0.152939
R20027 gnd.n5699 gnd.n5698 0.152939
R20028 gnd.n5700 gnd.n5699 0.152939
R20029 gnd.n5701 gnd.n5700 0.152939
R20030 gnd.n5702 gnd.n5701 0.152939
R20031 gnd.n5703 gnd.n5702 0.152939
R20032 gnd.n5704 gnd.n5703 0.152939
R20033 gnd.n5705 gnd.n5704 0.152939
R20034 gnd.n5706 gnd.n5705 0.152939
R20035 gnd.n5710 gnd.n5706 0.152939
R20036 gnd.n5710 gnd.n5488 0.152939
R20037 gnd.n6440 gnd.n6439 0.152939
R20038 gnd.n6447 gnd.n6439 0.152939
R20039 gnd.n6448 gnd.n6447 0.152939
R20040 gnd.n6449 gnd.n6448 0.152939
R20041 gnd.n6449 gnd.n6437 0.152939
R20042 gnd.n6457 gnd.n6437 0.152939
R20043 gnd.n6458 gnd.n6457 0.152939
R20044 gnd.n6459 gnd.n6458 0.152939
R20045 gnd.n6459 gnd.n6435 0.152939
R20046 gnd.n6467 gnd.n6435 0.152939
R20047 gnd.n6468 gnd.n6467 0.152939
R20048 gnd.n6469 gnd.n6468 0.152939
R20049 gnd.n6469 gnd.n6433 0.152939
R20050 gnd.n6477 gnd.n6433 0.152939
R20051 gnd.n6478 gnd.n6477 0.152939
R20052 gnd.n6479 gnd.n6478 0.152939
R20053 gnd.n6479 gnd.n6431 0.152939
R20054 gnd.n6487 gnd.n6431 0.152939
R20055 gnd.n6488 gnd.n6487 0.152939
R20056 gnd.n6489 gnd.n6488 0.152939
R20057 gnd.n6489 gnd.n6429 0.152939
R20058 gnd.n6500 gnd.n6429 0.152939
R20059 gnd.n6501 gnd.n6500 0.152939
R20060 gnd.n6502 gnd.n6501 0.152939
R20061 gnd.n6502 gnd.n6427 0.152939
R20062 gnd.n6509 gnd.n6427 0.152939
R20063 gnd.n5953 gnd.n5952 0.152939
R20064 gnd.n5954 gnd.n5953 0.152939
R20065 gnd.n5955 gnd.n5954 0.152939
R20066 gnd.n5956 gnd.n5955 0.152939
R20067 gnd.n5957 gnd.n5956 0.152939
R20068 gnd.n5958 gnd.n5957 0.152939
R20069 gnd.n5959 gnd.n5958 0.152939
R20070 gnd.n5959 gnd.n5218 0.152939
R20071 gnd.n6025 gnd.n5218 0.152939
R20072 gnd.n6026 gnd.n6025 0.152939
R20073 gnd.n6027 gnd.n6026 0.152939
R20074 gnd.n6028 gnd.n6027 0.152939
R20075 gnd.n6029 gnd.n6028 0.152939
R20076 gnd.n6029 gnd.n5181 0.152939
R20077 gnd.n6079 gnd.n5181 0.152939
R20078 gnd.n6080 gnd.n6079 0.152939
R20079 gnd.n6081 gnd.n6080 0.152939
R20080 gnd.n6082 gnd.n6081 0.152939
R20081 gnd.n6083 gnd.n6082 0.152939
R20082 gnd.n6084 gnd.n6083 0.152939
R20083 gnd.n6085 gnd.n6084 0.152939
R20084 gnd.n6086 gnd.n6085 0.152939
R20085 gnd.n6087 gnd.n6086 0.152939
R20086 gnd.n6087 gnd.n5127 0.152939
R20087 gnd.n6424 gnd.n5127 0.152939
R20088 gnd.n6425 gnd.n6424 0.152939
R20089 gnd.n6426 gnd.n6425 0.152939
R20090 gnd.n6510 gnd.n6426 0.152939
R20091 gnd.n5625 gnd.n5624 0.152939
R20092 gnd.n5626 gnd.n5625 0.152939
R20093 gnd.n5626 gnd.n5508 0.152939
R20094 gnd.n5640 gnd.n5508 0.152939
R20095 gnd.n5641 gnd.n5640 0.152939
R20096 gnd.n5642 gnd.n5641 0.152939
R20097 gnd.n5642 gnd.n5495 0.152939
R20098 gnd.n5656 gnd.n5495 0.152939
R20099 gnd.n5657 gnd.n5656 0.152939
R20100 gnd.n5658 gnd.n5657 0.152939
R20101 gnd.n5659 gnd.n5658 0.152939
R20102 gnd.n5660 gnd.n5659 0.152939
R20103 gnd.n5661 gnd.n5660 0.152939
R20104 gnd.n5662 gnd.n5661 0.152939
R20105 gnd.n5663 gnd.n5662 0.152939
R20106 gnd.n5664 gnd.n5663 0.152939
R20107 gnd.n5665 gnd.n5664 0.152939
R20108 gnd.n5666 gnd.n5665 0.152939
R20109 gnd.n5667 gnd.n5666 0.152939
R20110 gnd.n5667 gnd.n5430 0.152939
R20111 gnd.n5819 gnd.n5430 0.152939
R20112 gnd.n5820 gnd.n5819 0.152939
R20113 gnd.n5821 gnd.n5820 0.152939
R20114 gnd.n5822 gnd.n5821 0.152939
R20115 gnd.n5822 gnd.n5397 0.152939
R20116 gnd.n5866 gnd.n5397 0.152939
R20117 gnd.n5867 gnd.n5866 0.152939
R20118 gnd.n5868 gnd.n5867 0.152939
R20119 gnd.n5617 gnd.n5524 0.152939
R20120 gnd.n5527 gnd.n5524 0.152939
R20121 gnd.n5528 gnd.n5527 0.152939
R20122 gnd.n5529 gnd.n5528 0.152939
R20123 gnd.n5532 gnd.n5529 0.152939
R20124 gnd.n5533 gnd.n5532 0.152939
R20125 gnd.n5534 gnd.n5533 0.152939
R20126 gnd.n5535 gnd.n5534 0.152939
R20127 gnd.n5538 gnd.n5535 0.152939
R20128 gnd.n5539 gnd.n5538 0.152939
R20129 gnd.n5540 gnd.n5539 0.152939
R20130 gnd.n5541 gnd.n5540 0.152939
R20131 gnd.n5544 gnd.n5541 0.152939
R20132 gnd.n5545 gnd.n5544 0.152939
R20133 gnd.n5546 gnd.n5545 0.152939
R20134 gnd.n5547 gnd.n5546 0.152939
R20135 gnd.n5550 gnd.n5547 0.152939
R20136 gnd.n5551 gnd.n5550 0.152939
R20137 gnd.n5552 gnd.n5551 0.152939
R20138 gnd.n5553 gnd.n5552 0.152939
R20139 gnd.n5556 gnd.n5553 0.152939
R20140 gnd.n5557 gnd.n5556 0.152939
R20141 gnd.n5560 gnd.n5557 0.152939
R20142 gnd.n5561 gnd.n5560 0.152939
R20143 gnd.n5563 gnd.n5561 0.152939
R20144 gnd.n5563 gnd.n5520 0.152939
R20145 gnd.n6749 gnd.n948 0.152939
R20146 gnd.n6750 gnd.n6749 0.152939
R20147 gnd.n6751 gnd.n6750 0.152939
R20148 gnd.n6751 gnd.n942 0.152939
R20149 gnd.n6759 gnd.n942 0.152939
R20150 gnd.n6760 gnd.n6759 0.152939
R20151 gnd.n6761 gnd.n6760 0.152939
R20152 gnd.n6761 gnd.n936 0.152939
R20153 gnd.n6769 gnd.n936 0.152939
R20154 gnd.n6770 gnd.n6769 0.152939
R20155 gnd.n6771 gnd.n6770 0.152939
R20156 gnd.n6771 gnd.n930 0.152939
R20157 gnd.n6779 gnd.n930 0.152939
R20158 gnd.n6780 gnd.n6779 0.152939
R20159 gnd.n6781 gnd.n6780 0.152939
R20160 gnd.n6781 gnd.n924 0.152939
R20161 gnd.n6789 gnd.n924 0.152939
R20162 gnd.n6790 gnd.n6789 0.152939
R20163 gnd.n6791 gnd.n6790 0.152939
R20164 gnd.n6791 gnd.n918 0.152939
R20165 gnd.n6799 gnd.n918 0.152939
R20166 gnd.n6800 gnd.n6799 0.152939
R20167 gnd.n6801 gnd.n6800 0.152939
R20168 gnd.n6801 gnd.n912 0.152939
R20169 gnd.n6809 gnd.n912 0.152939
R20170 gnd.n6810 gnd.n6809 0.152939
R20171 gnd.n6811 gnd.n6810 0.152939
R20172 gnd.n6811 gnd.n906 0.152939
R20173 gnd.n6819 gnd.n906 0.152939
R20174 gnd.n6820 gnd.n6819 0.152939
R20175 gnd.n6821 gnd.n6820 0.152939
R20176 gnd.n6821 gnd.n900 0.152939
R20177 gnd.n6829 gnd.n900 0.152939
R20178 gnd.n6830 gnd.n6829 0.152939
R20179 gnd.n6831 gnd.n6830 0.152939
R20180 gnd.n6831 gnd.n894 0.152939
R20181 gnd.n6839 gnd.n894 0.152939
R20182 gnd.n6840 gnd.n6839 0.152939
R20183 gnd.n6841 gnd.n6840 0.152939
R20184 gnd.n6841 gnd.n888 0.152939
R20185 gnd.n6849 gnd.n888 0.152939
R20186 gnd.n6850 gnd.n6849 0.152939
R20187 gnd.n6851 gnd.n6850 0.152939
R20188 gnd.n6851 gnd.n882 0.152939
R20189 gnd.n6859 gnd.n882 0.152939
R20190 gnd.n6860 gnd.n6859 0.152939
R20191 gnd.n6861 gnd.n6860 0.152939
R20192 gnd.n6861 gnd.n876 0.152939
R20193 gnd.n6869 gnd.n876 0.152939
R20194 gnd.n6870 gnd.n6869 0.152939
R20195 gnd.n6871 gnd.n6870 0.152939
R20196 gnd.n6871 gnd.n870 0.152939
R20197 gnd.n6879 gnd.n870 0.152939
R20198 gnd.n6880 gnd.n6879 0.152939
R20199 gnd.n6881 gnd.n6880 0.152939
R20200 gnd.n6881 gnd.n864 0.152939
R20201 gnd.n6889 gnd.n864 0.152939
R20202 gnd.n6890 gnd.n6889 0.152939
R20203 gnd.n6891 gnd.n6890 0.152939
R20204 gnd.n6891 gnd.n858 0.152939
R20205 gnd.n6899 gnd.n858 0.152939
R20206 gnd.n6900 gnd.n6899 0.152939
R20207 gnd.n6901 gnd.n6900 0.152939
R20208 gnd.n6901 gnd.n852 0.152939
R20209 gnd.n6909 gnd.n852 0.152939
R20210 gnd.n6910 gnd.n6909 0.152939
R20211 gnd.n6911 gnd.n6910 0.152939
R20212 gnd.n6911 gnd.n846 0.152939
R20213 gnd.n6919 gnd.n846 0.152939
R20214 gnd.n6920 gnd.n6919 0.152939
R20215 gnd.n6921 gnd.n6920 0.152939
R20216 gnd.n6921 gnd.n840 0.152939
R20217 gnd.n6929 gnd.n840 0.152939
R20218 gnd.n6930 gnd.n6929 0.152939
R20219 gnd.n6931 gnd.n6930 0.152939
R20220 gnd.n6931 gnd.n834 0.152939
R20221 gnd.n6939 gnd.n834 0.152939
R20222 gnd.n6940 gnd.n6939 0.152939
R20223 gnd.n6941 gnd.n6940 0.152939
R20224 gnd.n6941 gnd.n828 0.152939
R20225 gnd.n6949 gnd.n828 0.152939
R20226 gnd.n6950 gnd.n6949 0.152939
R20227 gnd.n6951 gnd.n6950 0.152939
R20228 gnd.n6951 gnd.n822 0.152939
R20229 gnd.n6959 gnd.n822 0.152939
R20230 gnd.n6960 gnd.n6959 0.152939
R20231 gnd.n6961 gnd.n6960 0.152939
R20232 gnd.n6961 gnd.n816 0.152939
R20233 gnd.n6969 gnd.n816 0.152939
R20234 gnd.n6970 gnd.n6969 0.152939
R20235 gnd.n6971 gnd.n6970 0.152939
R20236 gnd.n6971 gnd.n810 0.152939
R20237 gnd.n6979 gnd.n810 0.152939
R20238 gnd.n6980 gnd.n6979 0.152939
R20239 gnd.n6981 gnd.n6980 0.152939
R20240 gnd.n6981 gnd.n804 0.152939
R20241 gnd.n6989 gnd.n804 0.152939
R20242 gnd.n6990 gnd.n6989 0.152939
R20243 gnd.n6991 gnd.n6990 0.152939
R20244 gnd.n6991 gnd.n798 0.152939
R20245 gnd.n6999 gnd.n798 0.152939
R20246 gnd.n7000 gnd.n6999 0.152939
R20247 gnd.n7001 gnd.n7000 0.152939
R20248 gnd.n7001 gnd.n792 0.152939
R20249 gnd.n7009 gnd.n792 0.152939
R20250 gnd.n7010 gnd.n7009 0.152939
R20251 gnd.n7011 gnd.n7010 0.152939
R20252 gnd.n7011 gnd.n786 0.152939
R20253 gnd.n7019 gnd.n786 0.152939
R20254 gnd.n7020 gnd.n7019 0.152939
R20255 gnd.n7021 gnd.n7020 0.152939
R20256 gnd.n7021 gnd.n780 0.152939
R20257 gnd.n7029 gnd.n780 0.152939
R20258 gnd.n7030 gnd.n7029 0.152939
R20259 gnd.n7031 gnd.n7030 0.152939
R20260 gnd.n7031 gnd.n774 0.152939
R20261 gnd.n7039 gnd.n774 0.152939
R20262 gnd.n7040 gnd.n7039 0.152939
R20263 gnd.n7041 gnd.n7040 0.152939
R20264 gnd.n7041 gnd.n768 0.152939
R20265 gnd.n7049 gnd.n768 0.152939
R20266 gnd.n7050 gnd.n7049 0.152939
R20267 gnd.n7051 gnd.n7050 0.152939
R20268 gnd.n7051 gnd.n762 0.152939
R20269 gnd.n7059 gnd.n762 0.152939
R20270 gnd.n7060 gnd.n7059 0.152939
R20271 gnd.n7061 gnd.n7060 0.152939
R20272 gnd.n7061 gnd.n756 0.152939
R20273 gnd.n7069 gnd.n756 0.152939
R20274 gnd.n7070 gnd.n7069 0.152939
R20275 gnd.n7071 gnd.n7070 0.152939
R20276 gnd.n7071 gnd.n750 0.152939
R20277 gnd.n7079 gnd.n750 0.152939
R20278 gnd.n7080 gnd.n7079 0.152939
R20279 gnd.n7081 gnd.n7080 0.152939
R20280 gnd.n7081 gnd.n744 0.152939
R20281 gnd.n7089 gnd.n744 0.152939
R20282 gnd.n7090 gnd.n7089 0.152939
R20283 gnd.n7091 gnd.n7090 0.152939
R20284 gnd.n7091 gnd.n738 0.152939
R20285 gnd.n7099 gnd.n738 0.152939
R20286 gnd.n7100 gnd.n7099 0.152939
R20287 gnd.n7101 gnd.n7100 0.152939
R20288 gnd.n7101 gnd.n732 0.152939
R20289 gnd.n7109 gnd.n732 0.152939
R20290 gnd.n7110 gnd.n7109 0.152939
R20291 gnd.n7111 gnd.n7110 0.152939
R20292 gnd.n7111 gnd.n726 0.152939
R20293 gnd.n7119 gnd.n726 0.152939
R20294 gnd.n7120 gnd.n7119 0.152939
R20295 gnd.n7122 gnd.n7120 0.152939
R20296 gnd.n7122 gnd.n7121 0.152939
R20297 gnd.n7121 gnd.n720 0.152939
R20298 gnd.n7131 gnd.n720 0.152939
R20299 gnd.n7132 gnd.n715 0.152939
R20300 gnd.n7140 gnd.n715 0.152939
R20301 gnd.n7141 gnd.n7140 0.152939
R20302 gnd.n7142 gnd.n7141 0.152939
R20303 gnd.n7142 gnd.n709 0.152939
R20304 gnd.n7150 gnd.n709 0.152939
R20305 gnd.n7151 gnd.n7150 0.152939
R20306 gnd.n7152 gnd.n7151 0.152939
R20307 gnd.n7152 gnd.n703 0.152939
R20308 gnd.n7160 gnd.n703 0.152939
R20309 gnd.n7161 gnd.n7160 0.152939
R20310 gnd.n7162 gnd.n7161 0.152939
R20311 gnd.n7162 gnd.n697 0.152939
R20312 gnd.n7170 gnd.n697 0.152939
R20313 gnd.n7171 gnd.n7170 0.152939
R20314 gnd.n7172 gnd.n7171 0.152939
R20315 gnd.n7172 gnd.n691 0.152939
R20316 gnd.n7180 gnd.n691 0.152939
R20317 gnd.n7181 gnd.n7180 0.152939
R20318 gnd.n7182 gnd.n7181 0.152939
R20319 gnd.n7182 gnd.n685 0.152939
R20320 gnd.n7190 gnd.n685 0.152939
R20321 gnd.n7191 gnd.n7190 0.152939
R20322 gnd.n7192 gnd.n7191 0.152939
R20323 gnd.n7192 gnd.n679 0.152939
R20324 gnd.n7200 gnd.n679 0.152939
R20325 gnd.n7201 gnd.n7200 0.152939
R20326 gnd.n7202 gnd.n7201 0.152939
R20327 gnd.n7202 gnd.n673 0.152939
R20328 gnd.n7210 gnd.n673 0.152939
R20329 gnd.n7211 gnd.n7210 0.152939
R20330 gnd.n7212 gnd.n7211 0.152939
R20331 gnd.n7212 gnd.n667 0.152939
R20332 gnd.n7220 gnd.n667 0.152939
R20333 gnd.n7221 gnd.n7220 0.152939
R20334 gnd.n7222 gnd.n7221 0.152939
R20335 gnd.n7222 gnd.n661 0.152939
R20336 gnd.n7230 gnd.n661 0.152939
R20337 gnd.n7231 gnd.n7230 0.152939
R20338 gnd.n7232 gnd.n7231 0.152939
R20339 gnd.n7232 gnd.n655 0.152939
R20340 gnd.n7240 gnd.n655 0.152939
R20341 gnd.n7241 gnd.n7240 0.152939
R20342 gnd.n7242 gnd.n7241 0.152939
R20343 gnd.n7242 gnd.n649 0.152939
R20344 gnd.n7250 gnd.n649 0.152939
R20345 gnd.n7251 gnd.n7250 0.152939
R20346 gnd.n7252 gnd.n7251 0.152939
R20347 gnd.n7252 gnd.n643 0.152939
R20348 gnd.n7260 gnd.n643 0.152939
R20349 gnd.n7261 gnd.n7260 0.152939
R20350 gnd.n7262 gnd.n7261 0.152939
R20351 gnd.n7262 gnd.n637 0.152939
R20352 gnd.n7270 gnd.n637 0.152939
R20353 gnd.n7271 gnd.n7270 0.152939
R20354 gnd.n7272 gnd.n7271 0.152939
R20355 gnd.n7272 gnd.n631 0.152939
R20356 gnd.n7280 gnd.n631 0.152939
R20357 gnd.n7281 gnd.n7280 0.152939
R20358 gnd.n7282 gnd.n7281 0.152939
R20359 gnd.n7282 gnd.n625 0.152939
R20360 gnd.n7290 gnd.n625 0.152939
R20361 gnd.n7291 gnd.n7290 0.152939
R20362 gnd.n7292 gnd.n7291 0.152939
R20363 gnd.n7292 gnd.n619 0.152939
R20364 gnd.n7300 gnd.n619 0.152939
R20365 gnd.n7301 gnd.n7300 0.152939
R20366 gnd.n7302 gnd.n7301 0.152939
R20367 gnd.n7302 gnd.n613 0.152939
R20368 gnd.n7310 gnd.n613 0.152939
R20369 gnd.n7311 gnd.n7310 0.152939
R20370 gnd.n7312 gnd.n7311 0.152939
R20371 gnd.n7312 gnd.n607 0.152939
R20372 gnd.n7320 gnd.n607 0.152939
R20373 gnd.n7321 gnd.n7320 0.152939
R20374 gnd.n7322 gnd.n7321 0.152939
R20375 gnd.n7322 gnd.n601 0.152939
R20376 gnd.n7330 gnd.n601 0.152939
R20377 gnd.n7331 gnd.n7330 0.152939
R20378 gnd.n7332 gnd.n7331 0.152939
R20379 gnd.n7332 gnd.n595 0.152939
R20380 gnd.n7342 gnd.n595 0.152939
R20381 gnd.n7343 gnd.n7342 0.152939
R20382 gnd.n7345 gnd.n7343 0.152939
R20383 gnd.n7752 gnd.n108 0.152939
R20384 gnd.n133 gnd.n108 0.152939
R20385 gnd.n134 gnd.n133 0.152939
R20386 gnd.n135 gnd.n134 0.152939
R20387 gnd.n150 gnd.n135 0.152939
R20388 gnd.n151 gnd.n150 0.152939
R20389 gnd.n152 gnd.n151 0.152939
R20390 gnd.n153 gnd.n152 0.152939
R20391 gnd.n170 gnd.n153 0.152939
R20392 gnd.n171 gnd.n170 0.152939
R20393 gnd.n172 gnd.n171 0.152939
R20394 gnd.n173 gnd.n172 0.152939
R20395 gnd.n188 gnd.n173 0.152939
R20396 gnd.n189 gnd.n188 0.152939
R20397 gnd.n190 gnd.n189 0.152939
R20398 gnd.n191 gnd.n190 0.152939
R20399 gnd.n208 gnd.n191 0.152939
R20400 gnd.n209 gnd.n208 0.152939
R20401 gnd.n210 gnd.n209 0.152939
R20402 gnd.n211 gnd.n210 0.152939
R20403 gnd.n227 gnd.n211 0.152939
R20404 gnd.n228 gnd.n227 0.152939
R20405 gnd.n229 gnd.n228 0.152939
R20406 gnd.n230 gnd.n229 0.152939
R20407 gnd.n246 gnd.n230 0.152939
R20408 gnd.n247 gnd.n246 0.152939
R20409 gnd.n7667 gnd.n247 0.152939
R20410 gnd.n7761 gnd.n97 0.152939
R20411 gnd.n382 gnd.n97 0.152939
R20412 gnd.n385 gnd.n382 0.152939
R20413 gnd.n386 gnd.n385 0.152939
R20414 gnd.n387 gnd.n386 0.152939
R20415 gnd.n387 gnd.n380 0.152939
R20416 gnd.n393 gnd.n380 0.152939
R20417 gnd.n394 gnd.n393 0.152939
R20418 gnd.n395 gnd.n394 0.152939
R20419 gnd.n395 gnd.n378 0.152939
R20420 gnd.n401 gnd.n378 0.152939
R20421 gnd.n402 gnd.n401 0.152939
R20422 gnd.n403 gnd.n402 0.152939
R20423 gnd.n403 gnd.n376 0.152939
R20424 gnd.n409 gnd.n376 0.152939
R20425 gnd.n410 gnd.n409 0.152939
R20426 gnd.n411 gnd.n410 0.152939
R20427 gnd.n411 gnd.n374 0.152939
R20428 gnd.n417 gnd.n374 0.152939
R20429 gnd.n418 gnd.n417 0.152939
R20430 gnd.n419 gnd.n418 0.152939
R20431 gnd.n419 gnd.n372 0.152939
R20432 gnd.n425 gnd.n372 0.152939
R20433 gnd.n426 gnd.n425 0.152939
R20434 gnd.n427 gnd.n426 0.152939
R20435 gnd.n427 gnd.n370 0.152939
R20436 gnd.n433 gnd.n370 0.152939
R20437 gnd.n434 gnd.n433 0.152939
R20438 gnd.n435 gnd.n434 0.152939
R20439 gnd.n435 gnd.n368 0.152939
R20440 gnd.n442 gnd.n368 0.152939
R20441 gnd.n479 gnd.n348 0.152939
R20442 gnd.n350 gnd.n348 0.152939
R20443 gnd.n351 gnd.n350 0.152939
R20444 gnd.n352 gnd.n351 0.152939
R20445 gnd.n353 gnd.n352 0.152939
R20446 gnd.n354 gnd.n353 0.152939
R20447 gnd.n355 gnd.n354 0.152939
R20448 gnd.n356 gnd.n355 0.152939
R20449 gnd.n357 gnd.n356 0.152939
R20450 gnd.n358 gnd.n357 0.152939
R20451 gnd.n359 gnd.n358 0.152939
R20452 gnd.n360 gnd.n359 0.152939
R20453 gnd.n361 gnd.n360 0.152939
R20454 gnd.n362 gnd.n361 0.152939
R20455 gnd.n363 gnd.n362 0.152939
R20456 gnd.n364 gnd.n363 0.152939
R20457 gnd.n444 gnd.n364 0.152939
R20458 gnd.n444 gnd.n443 0.152939
R20459 gnd.n7666 gnd.n248 0.152939
R20460 gnd.n290 gnd.n248 0.152939
R20461 gnd.n291 gnd.n290 0.152939
R20462 gnd.n292 gnd.n291 0.152939
R20463 gnd.n293 gnd.n292 0.152939
R20464 gnd.n294 gnd.n293 0.152939
R20465 gnd.n295 gnd.n294 0.152939
R20466 gnd.n296 gnd.n295 0.152939
R20467 gnd.n297 gnd.n296 0.152939
R20468 gnd.n298 gnd.n297 0.152939
R20469 gnd.n299 gnd.n298 0.152939
R20470 gnd.n300 gnd.n299 0.152939
R20471 gnd.n301 gnd.n300 0.152939
R20472 gnd.n302 gnd.n301 0.152939
R20473 gnd.n303 gnd.n302 0.152939
R20474 gnd.n304 gnd.n303 0.152939
R20475 gnd.n305 gnd.n304 0.152939
R20476 gnd.n306 gnd.n305 0.152939
R20477 gnd.n307 gnd.n306 0.152939
R20478 gnd.n308 gnd.n307 0.152939
R20479 gnd.n309 gnd.n308 0.152939
R20480 gnd.n310 gnd.n309 0.152939
R20481 gnd.n311 gnd.n310 0.152939
R20482 gnd.n312 gnd.n311 0.152939
R20483 gnd.n313 gnd.n312 0.152939
R20484 gnd.n314 gnd.n313 0.152939
R20485 gnd.n315 gnd.n314 0.152939
R20486 gnd.n316 gnd.n315 0.152939
R20487 gnd.n317 gnd.n316 0.152939
R20488 gnd.n318 gnd.n317 0.152939
R20489 gnd.n319 gnd.n318 0.152939
R20490 gnd.n320 gnd.n319 0.152939
R20491 gnd.n321 gnd.n320 0.152939
R20492 gnd.n322 gnd.n321 0.152939
R20493 gnd.n323 gnd.n322 0.152939
R20494 gnd.n324 gnd.n323 0.152939
R20495 gnd.n7587 gnd.n324 0.152939
R20496 gnd.n7587 gnd.n7586 0.152939
R20497 gnd.n7586 gnd.n7585 0.152939
R20498 gnd.n7585 gnd.n328 0.152939
R20499 gnd.n329 gnd.n328 0.152939
R20500 gnd.n330 gnd.n329 0.152939
R20501 gnd.n331 gnd.n330 0.152939
R20502 gnd.n332 gnd.n331 0.152939
R20503 gnd.n333 gnd.n332 0.152939
R20504 gnd.n334 gnd.n333 0.152939
R20505 gnd.n335 gnd.n334 0.152939
R20506 gnd.n336 gnd.n335 0.152939
R20507 gnd.n337 gnd.n336 0.152939
R20508 gnd.n338 gnd.n337 0.152939
R20509 gnd.n339 gnd.n338 0.152939
R20510 gnd.n340 gnd.n339 0.152939
R20511 gnd.n341 gnd.n340 0.152939
R20512 gnd.n342 gnd.n341 0.152939
R20513 gnd.n343 gnd.n342 0.152939
R20514 gnd.n344 gnd.n343 0.152939
R20515 gnd.n7545 gnd.n344 0.152939
R20516 gnd.n7545 gnd.n7544 0.152939
R20517 gnd.n1908 gnd.n1907 0.152939
R20518 gnd.n1909 gnd.n1908 0.152939
R20519 gnd.n1910 gnd.n1909 0.152939
R20520 gnd.n1911 gnd.n1910 0.152939
R20521 gnd.n1912 gnd.n1911 0.152939
R20522 gnd.n1913 gnd.n1912 0.152939
R20523 gnd.n1914 gnd.n1913 0.152939
R20524 gnd.n1915 gnd.n1914 0.152939
R20525 gnd.n1916 gnd.n1915 0.152939
R20526 gnd.n1917 gnd.n1916 0.152939
R20527 gnd.n1918 gnd.n1917 0.152939
R20528 gnd.n1919 gnd.n1918 0.152939
R20529 gnd.n1920 gnd.n1919 0.152939
R20530 gnd.n1921 gnd.n1920 0.152939
R20531 gnd.n1922 gnd.n1921 0.152939
R20532 gnd.n1923 gnd.n1922 0.152939
R20533 gnd.n1924 gnd.n1923 0.152939
R20534 gnd.n1927 gnd.n1924 0.152939
R20535 gnd.n1928 gnd.n1927 0.152939
R20536 gnd.n1929 gnd.n1928 0.152939
R20537 gnd.n1930 gnd.n1929 0.152939
R20538 gnd.n1931 gnd.n1930 0.152939
R20539 gnd.n1932 gnd.n1931 0.152939
R20540 gnd.n1933 gnd.n1932 0.152939
R20541 gnd.n1934 gnd.n1933 0.152939
R20542 gnd.n1939 gnd.n1938 0.152939
R20543 gnd.n1940 gnd.n1939 0.152939
R20544 gnd.n1941 gnd.n1940 0.152939
R20545 gnd.n1942 gnd.n1941 0.152939
R20546 gnd.n1943 gnd.n1942 0.152939
R20547 gnd.n1944 gnd.n1943 0.152939
R20548 gnd.n1945 gnd.n1944 0.152939
R20549 gnd.n1946 gnd.n1945 0.152939
R20550 gnd.n1947 gnd.n1946 0.152939
R20551 gnd.n1950 gnd.n1947 0.152939
R20552 gnd.n1951 gnd.n1950 0.152939
R20553 gnd.n1952 gnd.n1951 0.152939
R20554 gnd.n1953 gnd.n1952 0.152939
R20555 gnd.n1954 gnd.n1953 0.152939
R20556 gnd.n1955 gnd.n1954 0.152939
R20557 gnd.n1956 gnd.n1955 0.152939
R20558 gnd.n1957 gnd.n1956 0.152939
R20559 gnd.n1958 gnd.n1957 0.152939
R20560 gnd.n1959 gnd.n1958 0.152939
R20561 gnd.n1960 gnd.n1959 0.152939
R20562 gnd.n1961 gnd.n1960 0.152939
R20563 gnd.n1962 gnd.n1961 0.152939
R20564 gnd.n1963 gnd.n1962 0.152939
R20565 gnd.n1964 gnd.n1963 0.152939
R20566 gnd.n1965 gnd.n1964 0.152939
R20567 gnd.n1966 gnd.n1965 0.152939
R20568 gnd.n1967 gnd.n1966 0.152939
R20569 gnd.n1968 gnd.n1967 0.152939
R20570 gnd.n4387 gnd.n1968 0.152939
R20571 gnd.n4387 gnd.n4386 0.152939
R20572 gnd.n1989 gnd.n1988 0.152939
R20573 gnd.n1990 gnd.n1989 0.152939
R20574 gnd.n1991 gnd.n1990 0.152939
R20575 gnd.n1992 gnd.n1991 0.152939
R20576 gnd.n2013 gnd.n1992 0.152939
R20577 gnd.n2014 gnd.n2013 0.152939
R20578 gnd.n2015 gnd.n2014 0.152939
R20579 gnd.n2016 gnd.n2015 0.152939
R20580 gnd.n2034 gnd.n2016 0.152939
R20581 gnd.n2035 gnd.n2034 0.152939
R20582 gnd.n2036 gnd.n2035 0.152939
R20583 gnd.n2037 gnd.n2036 0.152939
R20584 gnd.n4330 gnd.n2037 0.152939
R20585 gnd.n4331 gnd.n4330 0.152939
R20586 gnd.n4332 gnd.n4331 0.152939
R20587 gnd.n4332 gnd.n562 0.152939
R20588 gnd.n7386 gnd.n562 0.152939
R20589 gnd.n7387 gnd.n7386 0.152939
R20590 gnd.n7388 gnd.n7387 0.152939
R20591 gnd.n7389 gnd.n7388 0.152939
R20592 gnd.n7389 gnd.n533 0.152939
R20593 gnd.n7422 gnd.n533 0.152939
R20594 gnd.n7423 gnd.n7422 0.152939
R20595 gnd.n7424 gnd.n7423 0.152939
R20596 gnd.n7425 gnd.n7424 0.152939
R20597 gnd.n7425 gnd.n109 0.152939
R20598 gnd.n7752 gnd.n109 0.152939
R20599 gnd.n7352 gnd.n590 0.152939
R20600 gnd.n7352 gnd.n7351 0.152939
R20601 gnd.n2905 gnd.n2904 0.152939
R20602 gnd.n2906 gnd.n2905 0.152939
R20603 gnd.n2907 gnd.n2906 0.152939
R20604 gnd.n2908 gnd.n2907 0.152939
R20605 gnd.n2911 gnd.n2908 0.152939
R20606 gnd.n2912 gnd.n2911 0.152939
R20607 gnd.n2913 gnd.n2912 0.152939
R20608 gnd.n2914 gnd.n2913 0.152939
R20609 gnd.n2916 gnd.n2914 0.152939
R20610 gnd.n2916 gnd.n2915 0.152939
R20611 gnd.n2915 gnd.n2611 0.152939
R20612 gnd.n2993 gnd.n2611 0.152939
R20613 gnd.n2994 gnd.n2993 0.152939
R20614 gnd.n2995 gnd.n2994 0.152939
R20615 gnd.n2995 gnd.n2607 0.152939
R20616 gnd.n3001 gnd.n2607 0.152939
R20617 gnd.n3002 gnd.n3001 0.152939
R20618 gnd.n3003 gnd.n3002 0.152939
R20619 gnd.n3004 gnd.n3003 0.152939
R20620 gnd.n3005 gnd.n3004 0.152939
R20621 gnd.n3005 gnd.n2589 0.152939
R20622 gnd.n3296 gnd.n2589 0.152939
R20623 gnd.n3297 gnd.n3296 0.152939
R20624 gnd.n3298 gnd.n3297 0.152939
R20625 gnd.n3298 gnd.n2585 0.152939
R20626 gnd.n3304 gnd.n2585 0.152939
R20627 gnd.n3305 gnd.n3304 0.152939
R20628 gnd.n3306 gnd.n3305 0.152939
R20629 gnd.n3307 gnd.n3306 0.152939
R20630 gnd.n3308 gnd.n3307 0.152939
R20631 gnd.n3309 gnd.n3308 0.152939
R20632 gnd.n3309 gnd.n2555 0.152939
R20633 gnd.n3332 gnd.n2555 0.152939
R20634 gnd.n3333 gnd.n3332 0.152939
R20635 gnd.n3334 gnd.n3333 0.152939
R20636 gnd.n3334 gnd.n2539 0.152939
R20637 gnd.n3365 gnd.n2539 0.152939
R20638 gnd.n3366 gnd.n3365 0.152939
R20639 gnd.n3367 gnd.n3366 0.152939
R20640 gnd.n3368 gnd.n3367 0.152939
R20641 gnd.n3369 gnd.n3368 0.152939
R20642 gnd.n3371 gnd.n3369 0.152939
R20643 gnd.n3371 gnd.n3370 0.152939
R20644 gnd.n3370 gnd.n1692 0.152939
R20645 gnd.n1693 gnd.n1692 0.152939
R20646 gnd.n1694 gnd.n1693 0.152939
R20647 gnd.n2503 gnd.n1694 0.152939
R20648 gnd.n2504 gnd.n2503 0.152939
R20649 gnd.n3531 gnd.n2504 0.152939
R20650 gnd.n3532 gnd.n3531 0.152939
R20651 gnd.n3533 gnd.n3532 0.152939
R20652 gnd.n3534 gnd.n3533 0.152939
R20653 gnd.n3534 gnd.n2481 0.152939
R20654 gnd.n3568 gnd.n2481 0.152939
R20655 gnd.n3569 gnd.n3568 0.152939
R20656 gnd.n3570 gnd.n3569 0.152939
R20657 gnd.n3570 gnd.n2453 0.152939
R20658 gnd.n3607 gnd.n2453 0.152939
R20659 gnd.n3608 gnd.n3607 0.152939
R20660 gnd.n3609 gnd.n3608 0.152939
R20661 gnd.n3610 gnd.n3609 0.152939
R20662 gnd.n3610 gnd.n2425 0.152939
R20663 gnd.n3647 gnd.n2425 0.152939
R20664 gnd.n3648 gnd.n3647 0.152939
R20665 gnd.n3650 gnd.n3648 0.152939
R20666 gnd.n3650 gnd.n3649 0.152939
R20667 gnd.n3649 gnd.n2406 0.152939
R20668 gnd.n2407 gnd.n2406 0.152939
R20669 gnd.n2408 gnd.n2407 0.152939
R20670 gnd.n2410 gnd.n2408 0.152939
R20671 gnd.n2411 gnd.n2410 0.152939
R20672 gnd.n2411 gnd.n2369 0.152939
R20673 gnd.n3742 gnd.n2369 0.152939
R20674 gnd.n3743 gnd.n3742 0.152939
R20675 gnd.n3744 gnd.n3743 0.152939
R20676 gnd.n3745 gnd.n3744 0.152939
R20677 gnd.n3745 gnd.n2344 0.152939
R20678 gnd.n3794 gnd.n2344 0.152939
R20679 gnd.n3795 gnd.n3794 0.152939
R20680 gnd.n3796 gnd.n3795 0.152939
R20681 gnd.n3797 gnd.n3796 0.152939
R20682 gnd.n3797 gnd.n2318 0.152939
R20683 gnd.n3831 gnd.n2318 0.152939
R20684 gnd.n3832 gnd.n3831 0.152939
R20685 gnd.n3833 gnd.n3832 0.152939
R20686 gnd.n3833 gnd.n2293 0.152939
R20687 gnd.n3892 gnd.n2293 0.152939
R20688 gnd.n3893 gnd.n3892 0.152939
R20689 gnd.n3894 gnd.n3893 0.152939
R20690 gnd.n3895 gnd.n3894 0.152939
R20691 gnd.n3895 gnd.n2270 0.152939
R20692 gnd.n3925 gnd.n2270 0.152939
R20693 gnd.n3926 gnd.n3925 0.152939
R20694 gnd.n3927 gnd.n3926 0.152939
R20695 gnd.n3928 gnd.n3927 0.152939
R20696 gnd.n3928 gnd.n2249 0.152939
R20697 gnd.n3977 gnd.n2249 0.152939
R20698 gnd.n3978 gnd.n3977 0.152939
R20699 gnd.n3979 gnd.n3978 0.152939
R20700 gnd.n3980 gnd.n3979 0.152939
R20701 gnd.n3980 gnd.n2220 0.152939
R20702 gnd.n4014 gnd.n2220 0.152939
R20703 gnd.n4015 gnd.n4014 0.152939
R20704 gnd.n4016 gnd.n4015 0.152939
R20705 gnd.n4016 gnd.n2131 0.152939
R20706 gnd.n4161 gnd.n2131 0.152939
R20707 gnd.n4162 gnd.n4161 0.152939
R20708 gnd.n4163 gnd.n4162 0.152939
R20709 gnd.n4163 gnd.n2118 0.152939
R20710 gnd.n4177 gnd.n2118 0.152939
R20711 gnd.n4178 gnd.n4177 0.152939
R20712 gnd.n4179 gnd.n4178 0.152939
R20713 gnd.n4181 gnd.n4179 0.152939
R20714 gnd.n4181 gnd.n4180 0.152939
R20715 gnd.n4180 gnd.n2105 0.152939
R20716 gnd.n4198 gnd.n2105 0.152939
R20717 gnd.n4199 gnd.n4198 0.152939
R20718 gnd.n4200 gnd.n4199 0.152939
R20719 gnd.n4201 gnd.n4200 0.152939
R20720 gnd.n4202 gnd.n4201 0.152939
R20721 gnd.n4205 gnd.n4202 0.152939
R20722 gnd.n4206 gnd.n4205 0.152939
R20723 gnd.n4207 gnd.n4206 0.152939
R20724 gnd.n4208 gnd.n4207 0.152939
R20725 gnd.n4211 gnd.n4208 0.152939
R20726 gnd.n4212 gnd.n4211 0.152939
R20727 gnd.n4213 gnd.n4212 0.152939
R20728 gnd.n4214 gnd.n4213 0.152939
R20729 gnd.n4217 gnd.n4214 0.152939
R20730 gnd.n4218 gnd.n4217 0.152939
R20731 gnd.n4219 gnd.n4218 0.152939
R20732 gnd.n4220 gnd.n4219 0.152939
R20733 gnd.n4221 gnd.n4220 0.152939
R20734 gnd.n4222 gnd.n4221 0.152939
R20735 gnd.n4222 gnd.n2058 0.152939
R20736 gnd.n4321 gnd.n2058 0.152939
R20737 gnd.n4322 gnd.n4321 0.152939
R20738 gnd.n4324 gnd.n4322 0.152939
R20739 gnd.n4324 gnd.n4323 0.152939
R20740 gnd.n4323 gnd.n577 0.152939
R20741 gnd.n578 gnd.n577 0.152939
R20742 gnd.n579 gnd.n578 0.152939
R20743 gnd.n582 gnd.n579 0.152939
R20744 gnd.n583 gnd.n582 0.152939
R20745 gnd.n584 gnd.n583 0.152939
R20746 gnd.n585 gnd.n584 0.152939
R20747 gnd.n588 gnd.n585 0.152939
R20748 gnd.n589 gnd.n588 0.152939
R20749 gnd.n590 gnd.n589 0.152939
R20750 gnd.n2802 gnd.n2743 0.152939
R20751 gnd.n2808 gnd.n2743 0.152939
R20752 gnd.n2809 gnd.n2808 0.152939
R20753 gnd.n2810 gnd.n2809 0.152939
R20754 gnd.n2810 gnd.n2741 0.152939
R20755 gnd.n2816 gnd.n2741 0.152939
R20756 gnd.n2817 gnd.n2816 0.152939
R20757 gnd.n2818 gnd.n2817 0.152939
R20758 gnd.n2818 gnd.n2739 0.152939
R20759 gnd.n2824 gnd.n2739 0.152939
R20760 gnd.n2825 gnd.n2824 0.152939
R20761 gnd.n2826 gnd.n2825 0.152939
R20762 gnd.n2826 gnd.n2737 0.152939
R20763 gnd.n2832 gnd.n2737 0.152939
R20764 gnd.n2833 gnd.n2832 0.152939
R20765 gnd.n2834 gnd.n2833 0.152939
R20766 gnd.n2834 gnd.n2735 0.152939
R20767 gnd.n2840 gnd.n2735 0.152939
R20768 gnd.n2841 gnd.n2840 0.152939
R20769 gnd.n2842 gnd.n2841 0.152939
R20770 gnd.n2842 gnd.n2733 0.152939
R20771 gnd.n2848 gnd.n2733 0.152939
R20772 gnd.n2849 gnd.n2848 0.152939
R20773 gnd.n2850 gnd.n2849 0.152939
R20774 gnd.n2850 gnd.n2731 0.152939
R20775 gnd.n2856 gnd.n2731 0.152939
R20776 gnd.n2857 gnd.n2856 0.152939
R20777 gnd.n2858 gnd.n2857 0.152939
R20778 gnd.n2858 gnd.n2729 0.152939
R20779 gnd.n2864 gnd.n2729 0.152939
R20780 gnd.n2865 gnd.n2864 0.152939
R20781 gnd.n2757 gnd.n1254 0.152939
R20782 gnd.n2765 gnd.n2757 0.152939
R20783 gnd.n2766 gnd.n2765 0.152939
R20784 gnd.n2767 gnd.n2766 0.152939
R20785 gnd.n2767 gnd.n2755 0.152939
R20786 gnd.n2775 gnd.n2755 0.152939
R20787 gnd.n2776 gnd.n2775 0.152939
R20788 gnd.n2777 gnd.n2776 0.152939
R20789 gnd.n2777 gnd.n2753 0.152939
R20790 gnd.n2785 gnd.n2753 0.152939
R20791 gnd.n2786 gnd.n2785 0.152939
R20792 gnd.n2787 gnd.n2786 0.152939
R20793 gnd.n2787 gnd.n2751 0.152939
R20794 gnd.n2795 gnd.n2751 0.152939
R20795 gnd.n2796 gnd.n2795 0.152939
R20796 gnd.n2797 gnd.n2796 0.152939
R20797 gnd.n2797 gnd.n2744 0.152939
R20798 gnd.n2801 gnd.n2744 0.152939
R20799 gnd.n4899 gnd.n1402 0.152939
R20800 gnd.n1427 gnd.n1402 0.152939
R20801 gnd.n1428 gnd.n1427 0.152939
R20802 gnd.n1429 gnd.n1428 0.152939
R20803 gnd.n1446 gnd.n1429 0.152939
R20804 gnd.n1447 gnd.n1446 0.152939
R20805 gnd.n1448 gnd.n1447 0.152939
R20806 gnd.n1449 gnd.n1448 0.152939
R20807 gnd.n1466 gnd.n1449 0.152939
R20808 gnd.n1467 gnd.n1466 0.152939
R20809 gnd.n1468 gnd.n1467 0.152939
R20810 gnd.n1469 gnd.n1468 0.152939
R20811 gnd.n1486 gnd.n1469 0.152939
R20812 gnd.n1487 gnd.n1486 0.152939
R20813 gnd.n1488 gnd.n1487 0.152939
R20814 gnd.n1489 gnd.n1488 0.152939
R20815 gnd.n1506 gnd.n1489 0.152939
R20816 gnd.n1507 gnd.n1506 0.152939
R20817 gnd.n1508 gnd.n1507 0.152939
R20818 gnd.n1509 gnd.n1508 0.152939
R20819 gnd.n1526 gnd.n1509 0.152939
R20820 gnd.n1527 gnd.n1526 0.152939
R20821 gnd.n1528 gnd.n1527 0.152939
R20822 gnd.n1529 gnd.n1528 0.152939
R20823 gnd.n1547 gnd.n1529 0.152939
R20824 gnd.n1548 gnd.n1547 0.152939
R20825 gnd.n4814 gnd.n1548 0.152939
R20826 gnd.n4813 gnd.n1549 0.152939
R20827 gnd.n1593 gnd.n1549 0.152939
R20828 gnd.n1594 gnd.n1593 0.152939
R20829 gnd.n1595 gnd.n1594 0.152939
R20830 gnd.n1596 gnd.n1595 0.152939
R20831 gnd.n1597 gnd.n1596 0.152939
R20832 gnd.n1598 gnd.n1597 0.152939
R20833 gnd.n1599 gnd.n1598 0.152939
R20834 gnd.n1600 gnd.n1599 0.152939
R20835 gnd.n1601 gnd.n1600 0.152939
R20836 gnd.n1602 gnd.n1601 0.152939
R20837 gnd.n1603 gnd.n1602 0.152939
R20838 gnd.n1604 gnd.n1603 0.152939
R20839 gnd.n1605 gnd.n1604 0.152939
R20840 gnd.n1606 gnd.n1605 0.152939
R20841 gnd.n1607 gnd.n1606 0.152939
R20842 gnd.n1608 gnd.n1607 0.152939
R20843 gnd.n1611 gnd.n1608 0.152939
R20844 gnd.n1612 gnd.n1611 0.152939
R20845 gnd.n1613 gnd.n1612 0.152939
R20846 gnd.n1614 gnd.n1613 0.152939
R20847 gnd.n1615 gnd.n1614 0.152939
R20848 gnd.n1616 gnd.n1615 0.152939
R20849 gnd.n1617 gnd.n1616 0.152939
R20850 gnd.n1618 gnd.n1617 0.152939
R20851 gnd.n3197 gnd.n3196 0.152939
R20852 gnd.n3204 gnd.n3197 0.152939
R20853 gnd.n3205 gnd.n3204 0.152939
R20854 gnd.n3206 gnd.n3205 0.152939
R20855 gnd.n3206 gnd.n3194 0.152939
R20856 gnd.n3214 gnd.n3194 0.152939
R20857 gnd.n3215 gnd.n3214 0.152939
R20858 gnd.n3216 gnd.n3215 0.152939
R20859 gnd.n3216 gnd.n3189 0.152939
R20860 gnd.n3223 gnd.n3189 0.152939
R20861 gnd.n3224 gnd.n3223 0.152939
R20862 gnd.n3225 gnd.n3224 0.152939
R20863 gnd.n3225 gnd.n3187 0.152939
R20864 gnd.n3233 gnd.n3187 0.152939
R20865 gnd.n3234 gnd.n3233 0.152939
R20866 gnd.n3235 gnd.n3234 0.152939
R20867 gnd.n3235 gnd.n3185 0.152939
R20868 gnd.n3243 gnd.n3185 0.152939
R20869 gnd.n3244 gnd.n3243 0.152939
R20870 gnd.n3245 gnd.n3244 0.152939
R20871 gnd.n3245 gnd.n3183 0.152939
R20872 gnd.n3253 gnd.n3183 0.152939
R20873 gnd.n3254 gnd.n3253 0.152939
R20874 gnd.n3255 gnd.n3254 0.152939
R20875 gnd.n3255 gnd.n3181 0.152939
R20876 gnd.n3263 gnd.n3181 0.152939
R20877 gnd.n3264 gnd.n3263 0.152939
R20878 gnd.n3265 gnd.n3264 0.152939
R20879 gnd.n3265 gnd.n3176 0.152939
R20880 gnd.n3271 gnd.n3176 0.152939
R20881 gnd.n1191 gnd.n1190 0.152939
R20882 gnd.n1192 gnd.n1191 0.152939
R20883 gnd.n1193 gnd.n1192 0.152939
R20884 gnd.n1194 gnd.n1193 0.152939
R20885 gnd.n1195 gnd.n1194 0.152939
R20886 gnd.n1196 gnd.n1195 0.152939
R20887 gnd.n1197 gnd.n1196 0.152939
R20888 gnd.n1198 gnd.n1197 0.152939
R20889 gnd.n1199 gnd.n1198 0.152939
R20890 gnd.n1200 gnd.n1199 0.152939
R20891 gnd.n1201 gnd.n1200 0.152939
R20892 gnd.n1202 gnd.n1201 0.152939
R20893 gnd.n1203 gnd.n1202 0.152939
R20894 gnd.n1204 gnd.n1203 0.152939
R20895 gnd.n1205 gnd.n1204 0.152939
R20896 gnd.n1206 gnd.n1205 0.152939
R20897 gnd.n1207 gnd.n1206 0.152939
R20898 gnd.n1210 gnd.n1207 0.152939
R20899 gnd.n1211 gnd.n1210 0.152939
R20900 gnd.n1212 gnd.n1211 0.152939
R20901 gnd.n1213 gnd.n1212 0.152939
R20902 gnd.n1214 gnd.n1213 0.152939
R20903 gnd.n1215 gnd.n1214 0.152939
R20904 gnd.n1216 gnd.n1215 0.152939
R20905 gnd.n1217 gnd.n1216 0.152939
R20906 gnd.n1218 gnd.n1217 0.152939
R20907 gnd.n1219 gnd.n1218 0.152939
R20908 gnd.n1220 gnd.n1219 0.152939
R20909 gnd.n1221 gnd.n1220 0.152939
R20910 gnd.n1222 gnd.n1221 0.152939
R20911 gnd.n1223 gnd.n1222 0.152939
R20912 gnd.n1224 gnd.n1223 0.152939
R20913 gnd.n1225 gnd.n1224 0.152939
R20914 gnd.n1226 gnd.n1225 0.152939
R20915 gnd.n1227 gnd.n1226 0.152939
R20916 gnd.n1228 gnd.n1227 0.152939
R20917 gnd.n1229 gnd.n1228 0.152939
R20918 gnd.n1232 gnd.n1229 0.152939
R20919 gnd.n1233 gnd.n1232 0.152939
R20920 gnd.n1234 gnd.n1233 0.152939
R20921 gnd.n1235 gnd.n1234 0.152939
R20922 gnd.n1236 gnd.n1235 0.152939
R20923 gnd.n1237 gnd.n1236 0.152939
R20924 gnd.n1238 gnd.n1237 0.152939
R20925 gnd.n1239 gnd.n1238 0.152939
R20926 gnd.n1240 gnd.n1239 0.152939
R20927 gnd.n1241 gnd.n1240 0.152939
R20928 gnd.n1242 gnd.n1241 0.152939
R20929 gnd.n1243 gnd.n1242 0.152939
R20930 gnd.n1244 gnd.n1243 0.152939
R20931 gnd.n1245 gnd.n1244 0.152939
R20932 gnd.n1246 gnd.n1245 0.152939
R20933 gnd.n1247 gnd.n1246 0.152939
R20934 gnd.n1248 gnd.n1247 0.152939
R20935 gnd.n1249 gnd.n1248 0.152939
R20936 gnd.n1250 gnd.n1249 0.152939
R20937 gnd.n4994 gnd.n1250 0.152939
R20938 gnd.n4994 gnd.n4993 0.152939
R20939 gnd.n1265 gnd.n1264 0.152939
R20940 gnd.n1266 gnd.n1265 0.152939
R20941 gnd.n1267 gnd.n1266 0.152939
R20942 gnd.n1287 gnd.n1267 0.152939
R20943 gnd.n1288 gnd.n1287 0.152939
R20944 gnd.n1289 gnd.n1288 0.152939
R20945 gnd.n1290 gnd.n1289 0.152939
R20946 gnd.n1305 gnd.n1290 0.152939
R20947 gnd.n1306 gnd.n1305 0.152939
R20948 gnd.n1307 gnd.n1306 0.152939
R20949 gnd.n1308 gnd.n1307 0.152939
R20950 gnd.n1325 gnd.n1308 0.152939
R20951 gnd.n1326 gnd.n1325 0.152939
R20952 gnd.n1327 gnd.n1326 0.152939
R20953 gnd.n1328 gnd.n1327 0.152939
R20954 gnd.n1343 gnd.n1328 0.152939
R20955 gnd.n1344 gnd.n1343 0.152939
R20956 gnd.n1345 gnd.n1344 0.152939
R20957 gnd.n1346 gnd.n1345 0.152939
R20958 gnd.n1363 gnd.n1346 0.152939
R20959 gnd.n1364 gnd.n1363 0.152939
R20960 gnd.n1365 gnd.n1364 0.152939
R20961 gnd.n1366 gnd.n1365 0.152939
R20962 gnd.n1381 gnd.n1366 0.152939
R20963 gnd.n1382 gnd.n1381 0.152939
R20964 gnd.n1383 gnd.n1382 0.152939
R20965 gnd.n4899 gnd.n1383 0.152939
R20966 gnd.n2904 gnd.n2638 0.152939
R20967 gnd.n954 gnd.n953 0.152939
R20968 gnd.n955 gnd.n954 0.152939
R20969 gnd.n960 gnd.n955 0.152939
R20970 gnd.n961 gnd.n960 0.152939
R20971 gnd.n962 gnd.n961 0.152939
R20972 gnd.n963 gnd.n962 0.152939
R20973 gnd.n968 gnd.n963 0.152939
R20974 gnd.n969 gnd.n968 0.152939
R20975 gnd.n970 gnd.n969 0.152939
R20976 gnd.n971 gnd.n970 0.152939
R20977 gnd.n976 gnd.n971 0.152939
R20978 gnd.n977 gnd.n976 0.152939
R20979 gnd.n978 gnd.n977 0.152939
R20980 gnd.n979 gnd.n978 0.152939
R20981 gnd.n984 gnd.n979 0.152939
R20982 gnd.n985 gnd.n984 0.152939
R20983 gnd.n986 gnd.n985 0.152939
R20984 gnd.n987 gnd.n986 0.152939
R20985 gnd.n992 gnd.n987 0.152939
R20986 gnd.n993 gnd.n992 0.152939
R20987 gnd.n994 gnd.n993 0.152939
R20988 gnd.n995 gnd.n994 0.152939
R20989 gnd.n1000 gnd.n995 0.152939
R20990 gnd.n1001 gnd.n1000 0.152939
R20991 gnd.n1002 gnd.n1001 0.152939
R20992 gnd.n1003 gnd.n1002 0.152939
R20993 gnd.n1008 gnd.n1003 0.152939
R20994 gnd.n1009 gnd.n1008 0.152939
R20995 gnd.n1010 gnd.n1009 0.152939
R20996 gnd.n1011 gnd.n1010 0.152939
R20997 gnd.n1016 gnd.n1011 0.152939
R20998 gnd.n1017 gnd.n1016 0.152939
R20999 gnd.n1018 gnd.n1017 0.152939
R21000 gnd.n1019 gnd.n1018 0.152939
R21001 gnd.n1024 gnd.n1019 0.152939
R21002 gnd.n1025 gnd.n1024 0.152939
R21003 gnd.n1026 gnd.n1025 0.152939
R21004 gnd.n1027 gnd.n1026 0.152939
R21005 gnd.n1032 gnd.n1027 0.152939
R21006 gnd.n1033 gnd.n1032 0.152939
R21007 gnd.n1034 gnd.n1033 0.152939
R21008 gnd.n1035 gnd.n1034 0.152939
R21009 gnd.n1040 gnd.n1035 0.152939
R21010 gnd.n1041 gnd.n1040 0.152939
R21011 gnd.n1042 gnd.n1041 0.152939
R21012 gnd.n1043 gnd.n1042 0.152939
R21013 gnd.n1048 gnd.n1043 0.152939
R21014 gnd.n1049 gnd.n1048 0.152939
R21015 gnd.n1050 gnd.n1049 0.152939
R21016 gnd.n1051 gnd.n1050 0.152939
R21017 gnd.n1056 gnd.n1051 0.152939
R21018 gnd.n1057 gnd.n1056 0.152939
R21019 gnd.n1058 gnd.n1057 0.152939
R21020 gnd.n1059 gnd.n1058 0.152939
R21021 gnd.n1064 gnd.n1059 0.152939
R21022 gnd.n1065 gnd.n1064 0.152939
R21023 gnd.n1066 gnd.n1065 0.152939
R21024 gnd.n1067 gnd.n1066 0.152939
R21025 gnd.n1072 gnd.n1067 0.152939
R21026 gnd.n1073 gnd.n1072 0.152939
R21027 gnd.n1074 gnd.n1073 0.152939
R21028 gnd.n1075 gnd.n1074 0.152939
R21029 gnd.n1080 gnd.n1075 0.152939
R21030 gnd.n1081 gnd.n1080 0.152939
R21031 gnd.n1082 gnd.n1081 0.152939
R21032 gnd.n1083 gnd.n1082 0.152939
R21033 gnd.n1088 gnd.n1083 0.152939
R21034 gnd.n1089 gnd.n1088 0.152939
R21035 gnd.n1090 gnd.n1089 0.152939
R21036 gnd.n1091 gnd.n1090 0.152939
R21037 gnd.n1096 gnd.n1091 0.152939
R21038 gnd.n1097 gnd.n1096 0.152939
R21039 gnd.n1098 gnd.n1097 0.152939
R21040 gnd.n1099 gnd.n1098 0.152939
R21041 gnd.n1104 gnd.n1099 0.152939
R21042 gnd.n1105 gnd.n1104 0.152939
R21043 gnd.n1106 gnd.n1105 0.152939
R21044 gnd.n1107 gnd.n1106 0.152939
R21045 gnd.n1112 gnd.n1107 0.152939
R21046 gnd.n1113 gnd.n1112 0.152939
R21047 gnd.n1114 gnd.n1113 0.152939
R21048 gnd.n1115 gnd.n1114 0.152939
R21049 gnd.n2654 gnd.n1115 0.152939
R21050 gnd.n2657 gnd.n2654 0.152939
R21051 gnd.n3340 gnd.n2548 0.152939
R21052 gnd.n3341 gnd.n3340 0.152939
R21053 gnd.n3359 gnd.n3341 0.152939
R21054 gnd.n3359 gnd.n3358 0.152939
R21055 gnd.n3358 gnd.n3357 0.152939
R21056 gnd.n3357 gnd.n3342 0.152939
R21057 gnd.n3353 gnd.n3342 0.152939
R21058 gnd.n3353 gnd.n3352 0.152939
R21059 gnd.n3352 gnd.n3351 0.152939
R21060 gnd.n3351 gnd.n3346 0.152939
R21061 gnd.n3346 gnd.n1703 0.152939
R21062 gnd.n4676 gnd.n1703 0.152939
R21063 gnd.n4676 gnd.n4675 0.152939
R21064 gnd.n4675 gnd.n4674 0.152939
R21065 gnd.n4674 gnd.n1704 0.152939
R21066 gnd.n4670 gnd.n1704 0.152939
R21067 gnd.n4670 gnd.n4669 0.152939
R21068 gnd.n4669 gnd.n4668 0.152939
R21069 gnd.n4668 gnd.n1709 0.152939
R21070 gnd.n4664 gnd.n1709 0.152939
R21071 gnd.n4664 gnd.n4663 0.152939
R21072 gnd.n4663 gnd.n4662 0.152939
R21073 gnd.n4662 gnd.n1714 0.152939
R21074 gnd.n4658 gnd.n1714 0.152939
R21075 gnd.n4658 gnd.n4657 0.152939
R21076 gnd.n4657 gnd.n4656 0.152939
R21077 gnd.n4656 gnd.n1719 0.152939
R21078 gnd.n4652 gnd.n1719 0.152939
R21079 gnd.n4652 gnd.n4651 0.152939
R21080 gnd.n4651 gnd.n4650 0.152939
R21081 gnd.n4650 gnd.n1724 0.152939
R21082 gnd.n4646 gnd.n1724 0.152939
R21083 gnd.n4646 gnd.n4645 0.152939
R21084 gnd.n4645 gnd.n4644 0.152939
R21085 gnd.n4644 gnd.n1729 0.152939
R21086 gnd.n4640 gnd.n1729 0.152939
R21087 gnd.n4640 gnd.n4639 0.152939
R21088 gnd.n4639 gnd.n4638 0.152939
R21089 gnd.n4638 gnd.n1734 0.152939
R21090 gnd.n4634 gnd.n1734 0.152939
R21091 gnd.n4634 gnd.n4633 0.152939
R21092 gnd.n4633 gnd.n4632 0.152939
R21093 gnd.n4632 gnd.n1739 0.152939
R21094 gnd.n4628 gnd.n1739 0.152939
R21095 gnd.n4628 gnd.n4627 0.152939
R21096 gnd.n4627 gnd.n4626 0.152939
R21097 gnd.n4626 gnd.n1744 0.152939
R21098 gnd.n4622 gnd.n1744 0.152939
R21099 gnd.n4622 gnd.n4621 0.152939
R21100 gnd.n4621 gnd.n4620 0.152939
R21101 gnd.n4620 gnd.n1749 0.152939
R21102 gnd.n4616 gnd.n1749 0.152939
R21103 gnd.n4616 gnd.n4615 0.152939
R21104 gnd.n4615 gnd.n4614 0.152939
R21105 gnd.n4614 gnd.n1754 0.152939
R21106 gnd.n4610 gnd.n1754 0.152939
R21107 gnd.n4610 gnd.n4609 0.152939
R21108 gnd.n4609 gnd.n4608 0.152939
R21109 gnd.n4608 gnd.n1759 0.152939
R21110 gnd.n4604 gnd.n1759 0.152939
R21111 gnd.n4604 gnd.n4603 0.152939
R21112 gnd.n4603 gnd.n4602 0.152939
R21113 gnd.n4602 gnd.n1764 0.152939
R21114 gnd.n4598 gnd.n1764 0.152939
R21115 gnd.n4598 gnd.n4597 0.152939
R21116 gnd.n4597 gnd.n4596 0.152939
R21117 gnd.n4596 gnd.n1769 0.152939
R21118 gnd.n4592 gnd.n1769 0.152939
R21119 gnd.n4592 gnd.n4591 0.152939
R21120 gnd.n4591 gnd.n4590 0.152939
R21121 gnd.n4590 gnd.n1774 0.152939
R21122 gnd.n4586 gnd.n1774 0.152939
R21123 gnd.n4586 gnd.n4585 0.152939
R21124 gnd.n4585 gnd.n4584 0.152939
R21125 gnd.n4584 gnd.n1779 0.152939
R21126 gnd.n4580 gnd.n1779 0.152939
R21127 gnd.n4580 gnd.n4579 0.152939
R21128 gnd.n4579 gnd.n4578 0.152939
R21129 gnd.n4578 gnd.n1784 0.152939
R21130 gnd.n4574 gnd.n1784 0.152939
R21131 gnd.n4574 gnd.n4573 0.152939
R21132 gnd.n4573 gnd.n4572 0.152939
R21133 gnd.n2894 gnd.n2645 0.152939
R21134 gnd.n2895 gnd.n2894 0.152939
R21135 gnd.n2896 gnd.n2895 0.152939
R21136 gnd.n2896 gnd.n2632 0.152939
R21137 gnd.n2933 gnd.n2632 0.152939
R21138 gnd.n2934 gnd.n2933 0.152939
R21139 gnd.n2935 gnd.n2934 0.152939
R21140 gnd.n2935 gnd.n2626 0.152939
R21141 gnd.n2947 gnd.n2626 0.152939
R21142 gnd.n2948 gnd.n2947 0.152939
R21143 gnd.n2949 gnd.n2948 0.152939
R21144 gnd.n2949 gnd.n2618 0.152939
R21145 gnd.n2984 gnd.n2618 0.152939
R21146 gnd.n2984 gnd.n2983 0.152939
R21147 gnd.n2983 gnd.n2982 0.152939
R21148 gnd.n2982 gnd.n2619 0.152939
R21149 gnd.n2978 gnd.n2619 0.152939
R21150 gnd.n2978 gnd.n2977 0.152939
R21151 gnd.n2977 gnd.n2976 0.152939
R21152 gnd.n2976 gnd.n2601 0.152939
R21153 gnd.n3014 gnd.n2601 0.152939
R21154 gnd.n3015 gnd.n3014 0.152939
R21155 gnd.n3016 gnd.n3015 0.152939
R21156 gnd.n3016 gnd.n2595 0.152939
R21157 gnd.n3288 gnd.n2595 0.152939
R21158 gnd.n3288 gnd.n3287 0.152939
R21159 gnd.n3287 gnd.n3286 0.152939
R21160 gnd.n3286 gnd.n2596 0.152939
R21161 gnd.n3282 gnd.n2596 0.152939
R21162 gnd.n3282 gnd.n3281 0.152939
R21163 gnd.n3281 gnd.n2575 0.152939
R21164 gnd.n3036 gnd.n3035 0.152939
R21165 gnd.n3053 gnd.n3035 0.152939
R21166 gnd.n3054 gnd.n3053 0.152939
R21167 gnd.n3055 gnd.n3054 0.152939
R21168 gnd.n3055 gnd.n3031 0.152939
R21169 gnd.n3174 gnd.n3031 0.152939
R21170 gnd.n3044 gnd.n3043 0.152939
R21171 gnd.n3043 gnd.n3042 0.152939
R21172 gnd.n3042 gnd.n3038 0.152939
R21173 gnd.n3038 gnd.n2530 0.152939
R21174 gnd.n3382 gnd.n2530 0.152939
R21175 gnd.n3383 gnd.n3382 0.152939
R21176 gnd.n3384 gnd.n3383 0.152939
R21177 gnd.n3384 gnd.n2526 0.152939
R21178 gnd.n3390 gnd.n2526 0.152939
R21179 gnd.n3391 gnd.n3390 0.152939
R21180 gnd.n3401 gnd.n3391 0.152939
R21181 gnd.n3401 gnd.n3400 0.152939
R21182 gnd.n3400 gnd.n3399 0.152939
R21183 gnd.n3399 gnd.n3392 0.152939
R21184 gnd.n3395 gnd.n3392 0.152939
R21185 gnd.n3395 gnd.n2494 0.152939
R21186 gnd.n3541 gnd.n2494 0.152939
R21187 gnd.n3542 gnd.n3541 0.152939
R21188 gnd.n3554 gnd.n3542 0.152939
R21189 gnd.n3554 gnd.n3553 0.152939
R21190 gnd.n3553 gnd.n3552 0.152939
R21191 gnd.n3552 gnd.n3543 0.152939
R21192 gnd.n3548 gnd.n3543 0.152939
R21193 gnd.n3548 gnd.n3547 0.152939
R21194 gnd.n3547 gnd.n2445 0.152939
R21195 gnd.n3617 gnd.n2445 0.152939
R21196 gnd.n3618 gnd.n3617 0.152939
R21197 gnd.n3620 gnd.n3618 0.152939
R21198 gnd.n3620 gnd.n3619 0.152939
R21199 gnd.n3619 gnd.n2418 0.152939
R21200 gnd.n3656 gnd.n2418 0.152939
R21201 gnd.n3657 gnd.n3656 0.152939
R21202 gnd.n3658 gnd.n3657 0.152939
R21203 gnd.n3658 gnd.n2416 0.152939
R21204 gnd.n3664 gnd.n2416 0.152939
R21205 gnd.n3665 gnd.n3664 0.152939
R21206 gnd.n3669 gnd.n3665 0.152939
R21207 gnd.n3669 gnd.n3668 0.152939
R21208 gnd.n3668 gnd.n3667 0.152939
R21209 gnd.n3667 gnd.n2359 0.152939
R21210 gnd.n3752 gnd.n2359 0.152939
R21211 gnd.n3753 gnd.n3752 0.152939
R21212 gnd.n3780 gnd.n3753 0.152939
R21213 gnd.n3780 gnd.n3779 0.152939
R21214 gnd.n3779 gnd.n3778 0.152939
R21215 gnd.n3778 gnd.n3754 0.152939
R21216 gnd.n3774 gnd.n3754 0.152939
R21217 gnd.n3774 gnd.n3773 0.152939
R21218 gnd.n3773 gnd.n3772 0.152939
R21219 gnd.n3772 gnd.n3761 0.152939
R21220 gnd.n3768 gnd.n3761 0.152939
R21221 gnd.n3768 gnd.n3767 0.152939
R21222 gnd.n3767 gnd.n3766 0.152939
R21223 gnd.n3766 gnd.n2286 0.152939
R21224 gnd.n3902 gnd.n2286 0.152939
R21225 gnd.n3903 gnd.n3902 0.152939
R21226 gnd.n3905 gnd.n3903 0.152939
R21227 gnd.n3905 gnd.n3904 0.152939
R21228 gnd.n3904 gnd.n2262 0.152939
R21229 gnd.n3935 gnd.n2262 0.152939
R21230 gnd.n3936 gnd.n3935 0.152939
R21231 gnd.n3963 gnd.n3936 0.152939
R21232 gnd.n3963 gnd.n3962 0.152939
R21233 gnd.n3962 gnd.n3961 0.152939
R21234 gnd.n3961 gnd.n3937 0.152939
R21235 gnd.n3957 gnd.n3937 0.152939
R21236 gnd.n3957 gnd.n3956 0.152939
R21237 gnd.n3956 gnd.n3955 0.152939
R21238 gnd.n3955 gnd.n3942 0.152939
R21239 gnd.n3951 gnd.n3942 0.152939
R21240 gnd.n3951 gnd.n3950 0.152939
R21241 gnd.n3950 gnd.n3949 0.152939
R21242 gnd.n3949 gnd.n2123 0.152939
R21243 gnd.n4169 gnd.n2123 0.152939
R21244 gnd.n4170 gnd.n4169 0.152939
R21245 gnd.n4171 gnd.n4170 0.152939
R21246 gnd.n4171 gnd.n2111 0.152939
R21247 gnd.n4188 gnd.n2111 0.152939
R21248 gnd.n4189 gnd.n4188 0.152939
R21249 gnd.n4190 gnd.n4189 0.152939
R21250 gnd.n4190 gnd.n1798 0.152939
R21251 gnd.n4566 gnd.n1798 0.152939
R21252 gnd.n4565 gnd.n1799 0.152939
R21253 gnd.n4561 gnd.n1799 0.152939
R21254 gnd.n4561 gnd.n4560 0.152939
R21255 gnd.n4560 gnd.n4559 0.152939
R21256 gnd.n4559 gnd.n1803 0.152939
R21257 gnd.n4555 gnd.n1803 0.152939
R21258 gnd.n4259 gnd.n4258 0.152939
R21259 gnd.n4259 gnd.n2072 0.152939
R21260 gnd.n4265 gnd.n2072 0.152939
R21261 gnd.n4266 gnd.n4265 0.152939
R21262 gnd.n4267 gnd.n4266 0.152939
R21263 gnd.n4267 gnd.n2068 0.152939
R21264 gnd.n4280 gnd.n2068 0.152939
R21265 gnd.n4281 gnd.n4280 0.152939
R21266 gnd.n4282 gnd.n4281 0.152939
R21267 gnd.n4282 gnd.n2064 0.152939
R21268 gnd.n4303 gnd.n2064 0.152939
R21269 gnd.n4304 gnd.n4303 0.152939
R21270 gnd.n4313 gnd.n4304 0.152939
R21271 gnd.n4313 gnd.n4312 0.152939
R21272 gnd.n4312 gnd.n4311 0.152939
R21273 gnd.n4311 gnd.n4305 0.152939
R21274 gnd.n4307 gnd.n4305 0.152939
R21275 gnd.n4307 gnd.n552 0.152939
R21276 gnd.n7396 gnd.n552 0.152939
R21277 gnd.n7397 gnd.n7396 0.152939
R21278 gnd.n7399 gnd.n7397 0.152939
R21279 gnd.n7399 gnd.n7398 0.152939
R21280 gnd.n7398 gnd.n523 0.152939
R21281 gnd.n7433 gnd.n523 0.152939
R21282 gnd.n7434 gnd.n7433 0.152939
R21283 gnd.n7435 gnd.n7434 0.152939
R21284 gnd.n7435 gnd.n501 0.152939
R21285 gnd.n7460 gnd.n501 0.152939
R21286 gnd.n7461 gnd.n7460 0.152939
R21287 gnd.n7462 gnd.n7461 0.152939
R21288 gnd.n7462 gnd.n95 0.152939
R21289 gnd.n7762 gnd.n7761 0.145814
R21290 gnd.n2866 gnd.n2865 0.145814
R21291 gnd.n2866 gnd.n2645 0.145814
R21292 gnd.n7762 gnd.n95 0.145814
R21293 gnd.n7351 gnd.n110 0.130073
R21294 gnd.n2638 gnd.n1403 0.130073
R21295 gnd.n3175 gnd.n3174 0.128549
R21296 gnd.n4555 gnd.n4554 0.128549
R21297 gnd.n5952 gnd.n5344 0.0767195
R21298 gnd.n5868 gnd.n5344 0.0767195
R21299 gnd.n3272 gnd.n3175 0.063
R21300 gnd.n4554 gnd.n1808 0.063
R21301 gnd.n6571 gnd.n1125 0.0477147
R21302 gnd.n5618 gnd.n5514 0.0442063
R21303 gnd.n5632 gnd.n5514 0.0442063
R21304 gnd.n5633 gnd.n5632 0.0442063
R21305 gnd.n5634 gnd.n5633 0.0442063
R21306 gnd.n5634 gnd.n5502 0.0442063
R21307 gnd.n5648 gnd.n5502 0.0442063
R21308 gnd.n5649 gnd.n5648 0.0442063
R21309 gnd.n5650 gnd.n5649 0.0442063
R21310 gnd.n5650 gnd.n5489 0.0442063
R21311 gnd.n5746 gnd.n5489 0.0442063
R21312 gnd.n1976 gnd.n1808 0.0416005
R21313 gnd.n7543 gnd.n7542 0.0416005
R21314 gnd.n4992 gnd.n4991 0.0416005
R21315 gnd.n3273 gnd.n3272 0.0416005
R21316 gnd.n5749 gnd.n5748 0.0344674
R21317 gnd.n4376 gnd.n1976 0.0344674
R21318 gnd.n4376 gnd.n1978 0.0344674
R21319 gnd.n2002 gnd.n1978 0.0344674
R21320 gnd.n2003 gnd.n2002 0.0344674
R21321 gnd.n2004 gnd.n2003 0.0344674
R21322 gnd.n2005 gnd.n2004 0.0344674
R21323 gnd.n4274 gnd.n2005 0.0344674
R21324 gnd.n4274 gnd.n2024 0.0344674
R21325 gnd.n2025 gnd.n2024 0.0344674
R21326 gnd.n2026 gnd.n2025 0.0344674
R21327 gnd.n4289 gnd.n2026 0.0344674
R21328 gnd.n4289 gnd.n2044 0.0344674
R21329 gnd.n2045 gnd.n2044 0.0344674
R21330 gnd.n2046 gnd.n2045 0.0344674
R21331 gnd.n4290 gnd.n2046 0.0344674
R21332 gnd.n4291 gnd.n4290 0.0344674
R21333 gnd.n4291 gnd.n571 0.0344674
R21334 gnd.n572 gnd.n571 0.0344674
R21335 gnd.n7374 gnd.n572 0.0344674
R21336 gnd.n7375 gnd.n7374 0.0344674
R21337 gnd.n7375 gnd.n546 0.0344674
R21338 gnd.n546 gnd.n543 0.0344674
R21339 gnd.n544 gnd.n543 0.0344674
R21340 gnd.n7410 gnd.n544 0.0344674
R21341 gnd.n7411 gnd.n7410 0.0344674
R21342 gnd.n7411 gnd.n518 0.0344674
R21343 gnd.n518 gnd.n513 0.0344674
R21344 gnd.n514 gnd.n513 0.0344674
R21345 gnd.n515 gnd.n514 0.0344674
R21346 gnd.n515 gnd.n488 0.0344674
R21347 gnd.n7476 gnd.n488 0.0344674
R21348 gnd.n7477 gnd.n7476 0.0344674
R21349 gnd.n7477 gnd.n483 0.0344674
R21350 gnd.n483 gnd.n481 0.0344674
R21351 gnd.n7488 gnd.n481 0.0344674
R21352 gnd.n7489 gnd.n7488 0.0344674
R21353 gnd.n7489 gnd.n124 0.0344674
R21354 gnd.n125 gnd.n124 0.0344674
R21355 gnd.n126 gnd.n125 0.0344674
R21356 gnd.n7497 gnd.n126 0.0344674
R21357 gnd.n7497 gnd.n141 0.0344674
R21358 gnd.n142 gnd.n141 0.0344674
R21359 gnd.n143 gnd.n142 0.0344674
R21360 gnd.n7504 gnd.n143 0.0344674
R21361 gnd.n7504 gnd.n161 0.0344674
R21362 gnd.n162 gnd.n161 0.0344674
R21363 gnd.n163 gnd.n162 0.0344674
R21364 gnd.n7511 gnd.n163 0.0344674
R21365 gnd.n7511 gnd.n179 0.0344674
R21366 gnd.n180 gnd.n179 0.0344674
R21367 gnd.n181 gnd.n180 0.0344674
R21368 gnd.n7518 gnd.n181 0.0344674
R21369 gnd.n7518 gnd.n199 0.0344674
R21370 gnd.n200 gnd.n199 0.0344674
R21371 gnd.n201 gnd.n200 0.0344674
R21372 gnd.n7525 gnd.n201 0.0344674
R21373 gnd.n7525 gnd.n217 0.0344674
R21374 gnd.n218 gnd.n217 0.0344674
R21375 gnd.n219 gnd.n218 0.0344674
R21376 gnd.n7532 gnd.n219 0.0344674
R21377 gnd.n7532 gnd.n237 0.0344674
R21378 gnd.n238 gnd.n237 0.0344674
R21379 gnd.n239 gnd.n238 0.0344674
R21380 gnd.n7542 gnd.n239 0.0344674
R21381 gnd.n4991 gnd.n1256 0.0344674
R21382 gnd.n2670 gnd.n1256 0.0344674
R21383 gnd.n2670 gnd.n1278 0.0344674
R21384 gnd.n1279 gnd.n1278 0.0344674
R21385 gnd.n1280 gnd.n1279 0.0344674
R21386 gnd.n2676 gnd.n1280 0.0344674
R21387 gnd.n2676 gnd.n1297 0.0344674
R21388 gnd.n1298 gnd.n1297 0.0344674
R21389 gnd.n1299 gnd.n1298 0.0344674
R21390 gnd.n2683 gnd.n1299 0.0344674
R21391 gnd.n2683 gnd.n1316 0.0344674
R21392 gnd.n1317 gnd.n1316 0.0344674
R21393 gnd.n1318 gnd.n1317 0.0344674
R21394 gnd.n2690 gnd.n1318 0.0344674
R21395 gnd.n2690 gnd.n1335 0.0344674
R21396 gnd.n1336 gnd.n1335 0.0344674
R21397 gnd.n1337 gnd.n1336 0.0344674
R21398 gnd.n2697 gnd.n1337 0.0344674
R21399 gnd.n2697 gnd.n1354 0.0344674
R21400 gnd.n1355 gnd.n1354 0.0344674
R21401 gnd.n1356 gnd.n1355 0.0344674
R21402 gnd.n2704 gnd.n1356 0.0344674
R21403 gnd.n2704 gnd.n1373 0.0344674
R21404 gnd.n1374 gnd.n1373 0.0344674
R21405 gnd.n1375 gnd.n1374 0.0344674
R21406 gnd.n2711 gnd.n1375 0.0344674
R21407 gnd.n2711 gnd.n1391 0.0344674
R21408 gnd.n1392 gnd.n1391 0.0344674
R21409 gnd.n1393 gnd.n1392 0.0344674
R21410 gnd.n2720 gnd.n1393 0.0344674
R21411 gnd.n2721 gnd.n2720 0.0344674
R21412 gnd.n2721 gnd.n2668 0.0344674
R21413 gnd.n2668 gnd.n2664 0.0344674
R21414 gnd.n2665 gnd.n2664 0.0344674
R21415 gnd.n2879 gnd.n2665 0.0344674
R21416 gnd.n2879 gnd.n2666 0.0344674
R21417 gnd.n2666 gnd.n1418 0.0344674
R21418 gnd.n1419 gnd.n1418 0.0344674
R21419 gnd.n1420 gnd.n1419 0.0344674
R21420 gnd.n2630 gnd.n1420 0.0344674
R21421 gnd.n2630 gnd.n1436 0.0344674
R21422 gnd.n1437 gnd.n1436 0.0344674
R21423 gnd.n1438 gnd.n1437 0.0344674
R21424 gnd.n2624 gnd.n1438 0.0344674
R21425 gnd.n2624 gnd.n1457 0.0344674
R21426 gnd.n1458 gnd.n1457 0.0344674
R21427 gnd.n1459 gnd.n1458 0.0344674
R21428 gnd.n2958 gnd.n1459 0.0344674
R21429 gnd.n2958 gnd.n1476 0.0344674
R21430 gnd.n1477 gnd.n1476 0.0344674
R21431 gnd.n1478 gnd.n1477 0.0344674
R21432 gnd.n2968 gnd.n1478 0.0344674
R21433 gnd.n2968 gnd.n1497 0.0344674
R21434 gnd.n1498 gnd.n1497 0.0344674
R21435 gnd.n1499 gnd.n1498 0.0344674
R21436 gnd.n2599 gnd.n1499 0.0344674
R21437 gnd.n2599 gnd.n1516 0.0344674
R21438 gnd.n1517 gnd.n1516 0.0344674
R21439 gnd.n1518 gnd.n1517 0.0344674
R21440 gnd.n3025 gnd.n1518 0.0344674
R21441 gnd.n3025 gnd.n1537 0.0344674
R21442 gnd.n1538 gnd.n1537 0.0344674
R21443 gnd.n1539 gnd.n1538 0.0344674
R21444 gnd.n3273 gnd.n1539 0.0344674
R21445 gnd.n3170 gnd.n3030 0.0344674
R21446 gnd.n4553 gnd.n4552 0.0344674
R21447 gnd.n3324 gnd.n3323 0.029712
R21448 gnd.n4257 gnd.n4256 0.029712
R21449 gnd.n5482 gnd.n5481 0.0269946
R21450 gnd.n5759 gnd.n5479 0.0269946
R21451 gnd.n5758 gnd.n5480 0.0269946
R21452 gnd.n5778 gnd.n5461 0.0269946
R21453 gnd.n5780 gnd.n5779 0.0269946
R21454 gnd.n5781 gnd.n5459 0.0269946
R21455 gnd.n5788 gnd.n5784 0.0269946
R21456 gnd.n5787 gnd.n5786 0.0269946
R21457 gnd.n5785 gnd.n5438 0.0269946
R21458 gnd.n5812 gnd.n5439 0.0269946
R21459 gnd.n5811 gnd.n5440 0.0269946
R21460 gnd.n5844 gnd.n5414 0.0269946
R21461 gnd.n5846 gnd.n5845 0.0269946
R21462 gnd.n5847 gnd.n5406 0.0269946
R21463 gnd.n5410 gnd.n5407 0.0269946
R21464 gnd.n5857 gnd.n5408 0.0269946
R21465 gnd.n5856 gnd.n5409 0.0269946
R21466 gnd.n5902 gnd.n5382 0.0269946
R21467 gnd.n5904 gnd.n5903 0.0269946
R21468 gnd.n5913 gnd.n5375 0.0269946
R21469 gnd.n5915 gnd.n5914 0.0269946
R21470 gnd.n5916 gnd.n5373 0.0269946
R21471 gnd.n5923 gnd.n5919 0.0269946
R21472 gnd.n5922 gnd.n5921 0.0269946
R21473 gnd.n5920 gnd.n5352 0.0269946
R21474 gnd.n5945 gnd.n5353 0.0269946
R21475 gnd.n5944 gnd.n5354 0.0269946
R21476 gnd.n5984 gnd.n5247 0.0269946
R21477 gnd.n5986 gnd.n5985 0.0269946
R21478 gnd.n5995 gnd.n5240 0.0269946
R21479 gnd.n5997 gnd.n5996 0.0269946
R21480 gnd.n5998 gnd.n5236 0.0269946
R21481 gnd.n6006 gnd.n5237 0.0269946
R21482 gnd.n6005 gnd.n5238 0.0269946
R21483 gnd.n6040 gnd.n5211 0.0269946
R21484 gnd.n6042 gnd.n6041 0.0269946
R21485 gnd.n6043 gnd.n5209 0.0269946
R21486 gnd.n6050 gnd.n6046 0.0269946
R21487 gnd.n6049 gnd.n6048 0.0269946
R21488 gnd.n6047 gnd.n5189 0.0269946
R21489 gnd.n6072 gnd.n5190 0.0269946
R21490 gnd.n6071 gnd.n5191 0.0269946
R21491 gnd.n6115 gnd.n5165 0.0269946
R21492 gnd.n6117 gnd.n6116 0.0269946
R21493 gnd.n6126 gnd.n5158 0.0269946
R21494 gnd.n6128 gnd.n6127 0.0269946
R21495 gnd.n6129 gnd.n5156 0.0269946
R21496 gnd.n6392 gnd.n6132 0.0269946
R21497 gnd.n6133 gnd.n5135 0.0269946
R21498 gnd.n6417 gnd.n5136 0.0269946
R21499 gnd.n6416 gnd.n5137 0.0269946
R21500 gnd.n6572 gnd.n1124 0.0269946
R21501 gnd.n7344 gnd.n110 0.0233659
R21502 gnd.n2656 gnd.n1403 0.0233659
R21503 gnd.n3169 gnd.n3063 0.0225788
R21504 gnd.n3166 gnd.n3165 0.0225788
R21505 gnd.n3162 gnd.n3066 0.0225788
R21506 gnd.n3161 gnd.n3072 0.0225788
R21507 gnd.n3158 gnd.n3157 0.0225788
R21508 gnd.n3154 gnd.n3078 0.0225788
R21509 gnd.n3153 gnd.n3082 0.0225788
R21510 gnd.n3150 gnd.n3149 0.0225788
R21511 gnd.n3146 gnd.n3086 0.0225788
R21512 gnd.n3145 gnd.n3092 0.0225788
R21513 gnd.n3142 gnd.n3141 0.0225788
R21514 gnd.n3138 gnd.n3098 0.0225788
R21515 gnd.n3137 gnd.n3102 0.0225788
R21516 gnd.n3134 gnd.n3133 0.0225788
R21517 gnd.n3130 gnd.n3106 0.0225788
R21518 gnd.n3129 gnd.n3112 0.0225788
R21519 gnd.n3126 gnd.n3125 0.0225788
R21520 gnd.n3117 gnd.n2576 0.0225788
R21521 gnd.n3323 gnd.n3322 0.0225788
R21522 gnd.n4549 gnd.n1809 0.0225788
R21523 gnd.n4548 gnd.n1813 0.0225788
R21524 gnd.n4545 gnd.n4544 0.0225788
R21525 gnd.n4541 gnd.n1818 0.0225788
R21526 gnd.n4540 gnd.n1822 0.0225788
R21527 gnd.n4537 gnd.n4536 0.0225788
R21528 gnd.n4533 gnd.n1826 0.0225788
R21529 gnd.n4532 gnd.n1830 0.0225788
R21530 gnd.n4529 gnd.n4528 0.0225788
R21531 gnd.n4525 gnd.n1834 0.0225788
R21532 gnd.n4524 gnd.n1838 0.0225788
R21533 gnd.n4521 gnd.n4520 0.0225788
R21534 gnd.n4517 gnd.n1842 0.0225788
R21535 gnd.n4516 gnd.n1846 0.0225788
R21536 gnd.n4513 gnd.n4512 0.0225788
R21537 gnd.n4509 gnd.n1850 0.0225788
R21538 gnd.n4508 gnd.n1856 0.0225788
R21539 gnd.n2076 gnd.n1859 0.0225788
R21540 gnd.n4256 gnd.n2075 0.0225788
R21541 gnd.n4257 gnd.n1789 0.0218415
R21542 gnd.n3325 gnd.n3324 0.0218415
R21543 gnd.n5748 gnd.n5747 0.0202011
R21544 gnd.n5747 gnd.n5746 0.0148637
R21545 gnd.n6391 gnd.n6390 0.0144266
R21546 gnd.n6390 gnd.n6134 0.0130679
R21547 gnd.n3170 gnd.n3169 0.0123886
R21548 gnd.n3166 gnd.n3063 0.0123886
R21549 gnd.n3165 gnd.n3066 0.0123886
R21550 gnd.n3162 gnd.n3161 0.0123886
R21551 gnd.n3158 gnd.n3072 0.0123886
R21552 gnd.n3157 gnd.n3078 0.0123886
R21553 gnd.n3154 gnd.n3153 0.0123886
R21554 gnd.n3150 gnd.n3082 0.0123886
R21555 gnd.n3149 gnd.n3086 0.0123886
R21556 gnd.n3146 gnd.n3145 0.0123886
R21557 gnd.n3142 gnd.n3092 0.0123886
R21558 gnd.n3141 gnd.n3098 0.0123886
R21559 gnd.n3138 gnd.n3137 0.0123886
R21560 gnd.n3134 gnd.n3102 0.0123886
R21561 gnd.n3133 gnd.n3106 0.0123886
R21562 gnd.n3130 gnd.n3129 0.0123886
R21563 gnd.n3126 gnd.n3112 0.0123886
R21564 gnd.n3125 gnd.n3117 0.0123886
R21565 gnd.n3322 gnd.n2576 0.0123886
R21566 gnd.n4552 gnd.n1809 0.0123886
R21567 gnd.n4549 gnd.n4548 0.0123886
R21568 gnd.n4545 gnd.n1813 0.0123886
R21569 gnd.n4544 gnd.n1818 0.0123886
R21570 gnd.n4541 gnd.n4540 0.0123886
R21571 gnd.n4537 gnd.n1822 0.0123886
R21572 gnd.n4536 gnd.n1826 0.0123886
R21573 gnd.n4533 gnd.n4532 0.0123886
R21574 gnd.n4529 gnd.n1830 0.0123886
R21575 gnd.n4528 gnd.n1834 0.0123886
R21576 gnd.n4525 gnd.n4524 0.0123886
R21577 gnd.n4521 gnd.n1838 0.0123886
R21578 gnd.n4520 gnd.n1842 0.0123886
R21579 gnd.n4517 gnd.n4516 0.0123886
R21580 gnd.n4513 gnd.n1846 0.0123886
R21581 gnd.n4512 gnd.n1850 0.0123886
R21582 gnd.n4509 gnd.n4508 0.0123886
R21583 gnd.n1859 gnd.n1856 0.0123886
R21584 gnd.n2076 gnd.n2075 0.0123886
R21585 gnd.n5749 gnd.n5482 0.00797283
R21586 gnd.n5481 gnd.n5479 0.00797283
R21587 gnd.n5759 gnd.n5758 0.00797283
R21588 gnd.n5480 gnd.n5461 0.00797283
R21589 gnd.n5779 gnd.n5778 0.00797283
R21590 gnd.n5781 gnd.n5780 0.00797283
R21591 gnd.n5784 gnd.n5459 0.00797283
R21592 gnd.n5788 gnd.n5787 0.00797283
R21593 gnd.n5786 gnd.n5785 0.00797283
R21594 gnd.n5439 gnd.n5438 0.00797283
R21595 gnd.n5812 gnd.n5811 0.00797283
R21596 gnd.n5440 gnd.n5414 0.00797283
R21597 gnd.n5845 gnd.n5844 0.00797283
R21598 gnd.n5847 gnd.n5846 0.00797283
R21599 gnd.n5410 gnd.n5406 0.00797283
R21600 gnd.n5408 gnd.n5407 0.00797283
R21601 gnd.n5857 gnd.n5856 0.00797283
R21602 gnd.n5409 gnd.n5382 0.00797283
R21603 gnd.n5904 gnd.n5902 0.00797283
R21604 gnd.n5903 gnd.n5375 0.00797283
R21605 gnd.n5914 gnd.n5913 0.00797283
R21606 gnd.n5916 gnd.n5915 0.00797283
R21607 gnd.n5919 gnd.n5373 0.00797283
R21608 gnd.n5923 gnd.n5922 0.00797283
R21609 gnd.n5921 gnd.n5920 0.00797283
R21610 gnd.n5353 gnd.n5352 0.00797283
R21611 gnd.n5945 gnd.n5944 0.00797283
R21612 gnd.n5354 gnd.n5247 0.00797283
R21613 gnd.n5986 gnd.n5984 0.00797283
R21614 gnd.n5985 gnd.n5240 0.00797283
R21615 gnd.n5996 gnd.n5995 0.00797283
R21616 gnd.n5998 gnd.n5997 0.00797283
R21617 gnd.n5237 gnd.n5236 0.00797283
R21618 gnd.n6006 gnd.n6005 0.00797283
R21619 gnd.n5238 gnd.n5211 0.00797283
R21620 gnd.n6041 gnd.n6040 0.00797283
R21621 gnd.n6043 gnd.n6042 0.00797283
R21622 gnd.n6046 gnd.n5209 0.00797283
R21623 gnd.n6050 gnd.n6049 0.00797283
R21624 gnd.n6048 gnd.n6047 0.00797283
R21625 gnd.n5190 gnd.n5189 0.00797283
R21626 gnd.n6072 gnd.n6071 0.00797283
R21627 gnd.n5191 gnd.n5165 0.00797283
R21628 gnd.n6117 gnd.n6115 0.00797283
R21629 gnd.n6116 gnd.n5158 0.00797283
R21630 gnd.n6127 gnd.n6126 0.00797283
R21631 gnd.n6129 gnd.n6128 0.00797283
R21632 gnd.n6132 gnd.n5156 0.00797283
R21633 gnd.n6392 gnd.n6391 0.00797283
R21634 gnd.n6134 gnd.n6133 0.00797283
R21635 gnd.n5136 gnd.n5135 0.00797283
R21636 gnd.n6417 gnd.n6416 0.00797283
R21637 gnd.n5137 gnd.n1124 0.00797283
R21638 gnd.n6572 gnd.n6571 0.00797283
R21639 gnd.n3175 gnd.n3030 0.00593478
R21640 gnd.n4554 gnd.n4553 0.00593478
R21641 a_n2408_n452.n95 a_n2408_n452.t73 512.366
R21642 a_n2408_n452.n85 a_n2408_n452.t64 512.366
R21643 a_n2408_n452.n96 a_n2408_n452.t56 512.366
R21644 a_n2408_n452.n93 a_n2408_n452.t81 512.366
R21645 a_n2408_n452.n86 a_n2408_n452.t70 512.366
R21646 a_n2408_n452.n94 a_n2408_n452.t69 512.366
R21647 a_n2408_n452.n91 a_n2408_n452.t77 512.366
R21648 a_n2408_n452.n87 a_n2408_n452.t62 512.366
R21649 a_n2408_n452.n92 a_n2408_n452.t63 512.366
R21650 a_n2408_n452.n89 a_n2408_n452.t65 512.366
R21651 a_n2408_n452.n88 a_n2408_n452.t75 512.366
R21652 a_n2408_n452.n90 a_n2408_n452.t87 512.366
R21653 a_n2408_n452.n36 a_n2408_n452.t86 533.335
R21654 a_n2408_n452.n101 a_n2408_n452.t67 512.366
R21655 a_n2408_n452.n67 a_n2408_n452.t71 512.366
R21656 a_n2408_n452.n100 a_n2408_n452.t61 512.366
R21657 a_n2408_n452.n99 a_n2408_n452.t76 512.366
R21658 a_n2408_n452.n68 a_n2408_n452.t83 512.366
R21659 a_n2408_n452.n98 a_n2408_n452.t84 512.366
R21660 a_n2408_n452.n35 a_n2408_n452.t12 533.335
R21661 a_n2408_n452.n102 a_n2408_n452.t4 512.366
R21662 a_n2408_n452.n65 a_n2408_n452.t22 512.366
R21663 a_n2408_n452.n31 a_n2408_n452.t8 533.335
R21664 a_n2408_n452.n117 a_n2408_n452.t16 512.366
R21665 a_n2408_n452.n66 a_n2408_n452.t6 512.366
R21666 a_n2408_n452.n116 a_n2408_n452.t14 512.366
R21667 a_n2408_n452.n115 a_n2408_n452.t2 512.366
R21668 a_n2408_n452.n49 a_n2408_n452.t18 533.335
R21669 a_n2408_n452.n79 a_n2408_n452.t24 512.366
R21670 a_n2408_n452.n80 a_n2408_n452.t30 512.366
R21671 a_n2408_n452.n81 a_n2408_n452.t32 512.366
R21672 a_n2408_n452.n82 a_n2408_n452.t20 512.366
R21673 a_n2408_n452.n72 a_n2408_n452.t10 512.366
R21674 a_n2408_n452.n83 a_n2408_n452.t28 512.366
R21675 a_n2408_n452.n42 a_n2408_n452.t82 533.335
R21676 a_n2408_n452.n74 a_n2408_n452.t60 512.366
R21677 a_n2408_n452.n75 a_n2408_n452.t79 512.366
R21678 a_n2408_n452.n76 a_n2408_n452.t80 512.366
R21679 a_n2408_n452.n77 a_n2408_n452.t57 512.366
R21680 a_n2408_n452.n73 a_n2408_n452.t66 512.366
R21681 a_n2408_n452.n78 a_n2408_n452.t74 512.366
R21682 a_n2408_n452.n5 a_n2408_n452.n63 70.1674
R21683 a_n2408_n452.n7 a_n2408_n452.n61 70.1674
R21684 a_n2408_n452.n9 a_n2408_n452.n59 70.1674
R21685 a_n2408_n452.n12 a_n2408_n452.n57 70.1674
R21686 a_n2408_n452.n41 a_n2408_n452.n21 70.1674
R21687 a_n2408_n452.n34 a_n2408_n452.n24 77.6622
R21688 a_n2408_n452.n115 a_n2408_n452.n34 5.97853
R21689 a_n2408_n452.n33 a_n2408_n452.n26 77.6622
R21690 a_n2408_n452.n26 a_n2408_n452.n32 72.3034
R21691 a_n2408_n452.n117 a_n2408_n452.n31 20.9683
R21692 a_n2408_n452.n25 a_n2408_n452.n31 70.1674
R21693 a_n2408_n452.n64 a_n2408_n452.n65 16.6962
R21694 a_n2408_n452.n35 a_n2408_n452.n24 70.1674
R21695 a_n2408_n452.n102 a_n2408_n452.n35 20.9683
R21696 a_n2408_n452.n24 a_n2408_n452.n64 72.3034
R21697 a_n2408_n452.n98 a_n2408_n452.n41 20.9683
R21698 a_n2408_n452.n22 a_n2408_n452.n40 72.3034
R21699 a_n2408_n452.n40 a_n2408_n452.n68 16.6962
R21700 a_n2408_n452.n39 a_n2408_n452.n22 77.6622
R21701 a_n2408_n452.n99 a_n2408_n452.n39 5.97853
R21702 a_n2408_n452.n38 a_n2408_n452.n20 77.6622
R21703 a_n2408_n452.n20 a_n2408_n452.n37 72.3034
R21704 a_n2408_n452.n101 a_n2408_n452.n36 20.9683
R21705 a_n2408_n452.n23 a_n2408_n452.n36 70.1674
R21706 a_n2408_n452.n14 a_n2408_n452.n55 70.1674
R21707 a_n2408_n452.n17 a_n2408_n452.n48 70.1674
R21708 a_n2408_n452.n78 a_n2408_n452.n48 20.9683
R21709 a_n2408_n452.n47 a_n2408_n452.n18 72.3034
R21710 a_n2408_n452.n47 a_n2408_n452.n73 16.6962
R21711 a_n2408_n452.n18 a_n2408_n452.n46 77.6622
R21712 a_n2408_n452.n77 a_n2408_n452.n46 5.97853
R21713 a_n2408_n452.n45 a_n2408_n452.n19 77.6622
R21714 a_n2408_n452.n19 a_n2408_n452.n44 72.3034
R21715 a_n2408_n452.n74 a_n2408_n452.n42 20.9683
R21716 a_n2408_n452.n43 a_n2408_n452.n42 70.1674
R21717 a_n2408_n452.n83 a_n2408_n452.n55 20.9683
R21718 a_n2408_n452.n54 a_n2408_n452.n15 72.3034
R21719 a_n2408_n452.n54 a_n2408_n452.n72 16.6962
R21720 a_n2408_n452.n15 a_n2408_n452.n53 77.6622
R21721 a_n2408_n452.n82 a_n2408_n452.n53 5.97853
R21722 a_n2408_n452.n52 a_n2408_n452.n16 77.6622
R21723 a_n2408_n452.n16 a_n2408_n452.n51 72.3034
R21724 a_n2408_n452.n79 a_n2408_n452.n49 20.9683
R21725 a_n2408_n452.n50 a_n2408_n452.n49 70.1674
R21726 a_n2408_n452.n90 a_n2408_n452.n57 20.9683
R21727 a_n2408_n452.n56 a_n2408_n452.n13 75.0448
R21728 a_n2408_n452.n56 a_n2408_n452.n88 11.2134
R21729 a_n2408_n452.n13 a_n2408_n452.n89 161.3
R21730 a_n2408_n452.n92 a_n2408_n452.n59 20.9683
R21731 a_n2408_n452.n58 a_n2408_n452.n10 75.0448
R21732 a_n2408_n452.n58 a_n2408_n452.n87 11.2134
R21733 a_n2408_n452.n10 a_n2408_n452.n91 161.3
R21734 a_n2408_n452.n94 a_n2408_n452.n61 20.9683
R21735 a_n2408_n452.n60 a_n2408_n452.n8 75.0448
R21736 a_n2408_n452.n60 a_n2408_n452.n86 11.2134
R21737 a_n2408_n452.n8 a_n2408_n452.n93 161.3
R21738 a_n2408_n452.n96 a_n2408_n452.n63 20.9683
R21739 a_n2408_n452.n62 a_n2408_n452.n6 75.0448
R21740 a_n2408_n452.n62 a_n2408_n452.n85 11.2134
R21741 a_n2408_n452.n6 a_n2408_n452.n95 161.3
R21742 a_n2408_n452.n3 a_n2408_n452.n112 81.3764
R21743 a_n2408_n452.n4 a_n2408_n452.n106 81.3764
R21744 a_n2408_n452.n0 a_n2408_n452.n103 81.3764
R21745 a_n2408_n452.n3 a_n2408_n452.n113 80.9324
R21746 a_n2408_n452.n2 a_n2408_n452.n114 80.9324
R21747 a_n2408_n452.n2 a_n2408_n452.n111 80.9324
R21748 a_n2408_n452.n2 a_n2408_n452.n110 80.9324
R21749 a_n2408_n452.n1 a_n2408_n452.n109 80.9324
R21750 a_n2408_n452.n4 a_n2408_n452.n107 80.9324
R21751 a_n2408_n452.n0 a_n2408_n452.n108 80.9324
R21752 a_n2408_n452.n0 a_n2408_n452.n105 80.9324
R21753 a_n2408_n452.n0 a_n2408_n452.n104 80.9324
R21754 a_n2408_n452.n30 a_n2408_n452.t13 74.6477
R21755 a_n2408_n452.n27 a_n2408_n452.t19 74.6477
R21756 a_n2408_n452.n29 a_n2408_n452.t9 74.2899
R21757 a_n2408_n452.n28 a_n2408_n452.t27 74.2897
R21758 a_n2408_n452.n30 a_n2408_n452.n120 70.6783
R21759 a_n2408_n452.n29 a_n2408_n452.n119 70.6783
R21760 a_n2408_n452.n28 a_n2408_n452.n71 70.6783
R21761 a_n2408_n452.n27 a_n2408_n452.n70 70.6783
R21762 a_n2408_n452.n27 a_n2408_n452.n69 70.6783
R21763 a_n2408_n452.n121 a_n2408_n452.n30 70.6782
R21764 a_n2408_n452.n95 a_n2408_n452.n85 48.2005
R21765 a_n2408_n452.t78 a_n2408_n452.n63 533.335
R21766 a_n2408_n452.n93 a_n2408_n452.n86 48.2005
R21767 a_n2408_n452.t85 a_n2408_n452.n61 533.335
R21768 a_n2408_n452.n91 a_n2408_n452.n87 48.2005
R21769 a_n2408_n452.t72 a_n2408_n452.n59 533.335
R21770 a_n2408_n452.n89 a_n2408_n452.n88 48.2005
R21771 a_n2408_n452.t68 a_n2408_n452.n57 533.335
R21772 a_n2408_n452.n100 a_n2408_n452.n99 48.2005
R21773 a_n2408_n452.n41 a_n2408_n452.t58 533.335
R21774 a_n2408_n452.n116 a_n2408_n452.n115 48.2005
R21775 a_n2408_n452.n82 a_n2408_n452.n81 48.2005
R21776 a_n2408_n452.t26 a_n2408_n452.n55 533.335
R21777 a_n2408_n452.n77 a_n2408_n452.n76 48.2005
R21778 a_n2408_n452.t59 a_n2408_n452.n48 533.335
R21779 a_n2408_n452.n37 a_n2408_n452.n67 16.6962
R21780 a_n2408_n452.n98 a_n2408_n452.n40 27.6507
R21781 a_n2408_n452.n102 a_n2408_n452.n64 27.6507
R21782 a_n2408_n452.n32 a_n2408_n452.n66 16.6962
R21783 a_n2408_n452.n80 a_n2408_n452.n51 16.6962
R21784 a_n2408_n452.n83 a_n2408_n452.n54 27.6507
R21785 a_n2408_n452.n75 a_n2408_n452.n44 16.6962
R21786 a_n2408_n452.n78 a_n2408_n452.n47 27.6507
R21787 a_n2408_n452.n38 a_n2408_n452.n67 41.7634
R21788 a_n2408_n452.n33 a_n2408_n452.n66 41.7634
R21789 a_n2408_n452.n80 a_n2408_n452.n52 41.7634
R21790 a_n2408_n452.n75 a_n2408_n452.n45 41.7634
R21791 a_n2408_n452.n1 a_n2408_n452.n0 32.6799
R21792 a_n2408_n452.n96 a_n2408_n452.n62 35.3134
R21793 a_n2408_n452.n94 a_n2408_n452.n60 35.3134
R21794 a_n2408_n452.n92 a_n2408_n452.n58 35.3134
R21795 a_n2408_n452.n90 a_n2408_n452.n56 35.3134
R21796 a_n2408_n452.n24 a_n2408_n452.n2 23.891
R21797 a_n2408_n452.n43 a_n2408_n452.n11 12.705
R21798 a_n2408_n452.n21 a_n2408_n452.n97 12.5005
R21799 a_n2408_n452.n38 a_n2408_n452.n100 5.97853
R21800 a_n2408_n452.n39 a_n2408_n452.n68 41.7634
R21801 a_n2408_n452.n33 a_n2408_n452.n116 5.97853
R21802 a_n2408_n452.n34 a_n2408_n452.n65 41.7634
R21803 a_n2408_n452.n81 a_n2408_n452.n52 5.97853
R21804 a_n2408_n452.n72 a_n2408_n452.n53 41.7634
R21805 a_n2408_n452.n76 a_n2408_n452.n45 5.97853
R21806 a_n2408_n452.n73 a_n2408_n452.n46 41.7634
R21807 a_n2408_n452.n118 a_n2408_n452.n25 11.1956
R21808 a_n2408_n452.n101 a_n2408_n452.n37 27.6507
R21809 a_n2408_n452.n117 a_n2408_n452.n32 27.6507
R21810 a_n2408_n452.n51 a_n2408_n452.n79 27.6507
R21811 a_n2408_n452.n44 a_n2408_n452.n74 27.6507
R21812 a_n2408_n452.n84 a_n2408_n452.n28 9.85898
R21813 a_n2408_n452.n97 a_n2408_n452.n5 8.73345
R21814 a_n2408_n452.n13 a_n2408_n452.n11 8.73345
R21815 a_n2408_n452.n84 a_n2408_n452.n14 7.36035
R21816 a_n2408_n452.n29 a_n2408_n452.n118 6.01559
R21817 a_n2408_n452.n97 a_n2408_n452.n84 5.3452
R21818 a_n2408_n452.n24 a_n2408_n452.n23 4.01186
R21819 a_n2408_n452.n50 a_n2408_n452.n17 4.01186
R21820 a_n2408_n452.n120 a_n2408_n452.t23 3.61217
R21821 a_n2408_n452.n120 a_n2408_n452.t5 3.61217
R21822 a_n2408_n452.n119 a_n2408_n452.t17 3.61217
R21823 a_n2408_n452.n119 a_n2408_n452.t7 3.61217
R21824 a_n2408_n452.n71 a_n2408_n452.t11 3.61217
R21825 a_n2408_n452.n71 a_n2408_n452.t29 3.61217
R21826 a_n2408_n452.n70 a_n2408_n452.t33 3.61217
R21827 a_n2408_n452.n70 a_n2408_n452.t21 3.61217
R21828 a_n2408_n452.n69 a_n2408_n452.t25 3.61217
R21829 a_n2408_n452.n69 a_n2408_n452.t31 3.61217
R21830 a_n2408_n452.n121 a_n2408_n452.t15 3.61217
R21831 a_n2408_n452.t3 a_n2408_n452.n121 3.61217
R21832 a_n2408_n452.n112 a_n2408_n452.t36 2.82907
R21833 a_n2408_n452.n112 a_n2408_n452.t45 2.82907
R21834 a_n2408_n452.n113 a_n2408_n452.t42 2.82907
R21835 a_n2408_n452.n113 a_n2408_n452.t40 2.82907
R21836 a_n2408_n452.n114 a_n2408_n452.t35 2.82907
R21837 a_n2408_n452.n114 a_n2408_n452.t51 2.82907
R21838 a_n2408_n452.n111 a_n2408_n452.t54 2.82907
R21839 a_n2408_n452.n111 a_n2408_n452.t34 2.82907
R21840 a_n2408_n452.n110 a_n2408_n452.t44 2.82907
R21841 a_n2408_n452.n110 a_n2408_n452.t47 2.82907
R21842 a_n2408_n452.n109 a_n2408_n452.t53 2.82907
R21843 a_n2408_n452.n109 a_n2408_n452.t39 2.82907
R21844 a_n2408_n452.n106 a_n2408_n452.t41 2.82907
R21845 a_n2408_n452.n106 a_n2408_n452.t46 2.82907
R21846 a_n2408_n452.n107 a_n2408_n452.t37 2.82907
R21847 a_n2408_n452.n107 a_n2408_n452.t43 2.82907
R21848 a_n2408_n452.n108 a_n2408_n452.t48 2.82907
R21849 a_n2408_n452.n108 a_n2408_n452.t55 2.82907
R21850 a_n2408_n452.n105 a_n2408_n452.t1 2.82907
R21851 a_n2408_n452.n105 a_n2408_n452.t50 2.82907
R21852 a_n2408_n452.n104 a_n2408_n452.t0 2.82907
R21853 a_n2408_n452.n104 a_n2408_n452.t38 2.82907
R21854 a_n2408_n452.n103 a_n2408_n452.t49 2.82907
R21855 a_n2408_n452.n103 a_n2408_n452.t52 2.82907
R21856 a_n2408_n452.n0 a_n2408_n452.n4 1.3324
R21857 a_n2408_n452.n118 a_n2408_n452.n11 1.30542
R21858 a_n2408_n452.n24 a_n2408_n452.n26 1.09898
R21859 a_n2408_n452.n30 a_n2408_n452.n29 1.07378
R21860 a_n2408_n452.n28 a_n2408_n452.n27 1.07378
R21861 a_n2408_n452.n8 a_n2408_n452.n9 1.04595
R21862 a_n2408_n452.n26 a_n2408_n452.n25 0.94747
R21863 a_n2408_n452.n2 a_n2408_n452.n3 0.888431
R21864 a_n2408_n452.n2 a_n2408_n452.n1 0.888431
R21865 a_n2408_n452.n22 a_n2408_n452.n20 0.758076
R21866 a_n2408_n452.n22 a_n2408_n452.n21 0.758076
R21867 a_n2408_n452.n19 a_n2408_n452.n18 0.758076
R21868 a_n2408_n452.n18 a_n2408_n452.n17 0.758076
R21869 a_n2408_n452.n16 a_n2408_n452.n15 0.758076
R21870 a_n2408_n452.n15 a_n2408_n452.n14 0.758076
R21871 a_n2408_n452.n13 a_n2408_n452.n12 0.758076
R21872 a_n2408_n452.n10 a_n2408_n452.n9 0.758076
R21873 a_n2408_n452.n8 a_n2408_n452.n7 0.758076
R21874 a_n2408_n452.n6 a_n2408_n452.n5 0.758076
R21875 a_n2408_n452.n10 a_n2408_n452.n12 0.67853
R21876 a_n2408_n452.n6 a_n2408_n452.n7 0.67853
R21877 a_n2408_n452.n50 a_n2408_n452.n16 0.568682
R21878 a_n2408_n452.n43 a_n2408_n452.n19 0.568682
R21879 a_n2408_n452.n20 a_n2408_n452.n23 0.568682
R21880 a_n2140_13878.n21 a_n2140_13878.n20 98.9632
R21881 a_n2140_13878.n2 a_n2140_13878.n0 98.7517
R21882 a_n2140_13878.n18 a_n2140_13878.n17 98.6055
R21883 a_n2140_13878.n20 a_n2140_13878.n19 98.6055
R21884 a_n2140_13878.n6 a_n2140_13878.n5 98.6055
R21885 a_n2140_13878.n4 a_n2140_13878.n3 98.6055
R21886 a_n2140_13878.n2 a_n2140_13878.n1 98.6055
R21887 a_n2140_13878.n16 a_n2140_13878.n15 98.6054
R21888 a_n2140_13878.n8 a_n2140_13878.t17 74.6477
R21889 a_n2140_13878.n13 a_n2140_13878.t18 74.2899
R21890 a_n2140_13878.n10 a_n2140_13878.t19 74.2899
R21891 a_n2140_13878.n9 a_n2140_13878.t16 74.2899
R21892 a_n2140_13878.n12 a_n2140_13878.n11 70.6783
R21893 a_n2140_13878.n8 a_n2140_13878.n7 70.6783
R21894 a_n2140_13878.n14 a_n2140_13878.n6 14.2849
R21895 a_n2140_13878.n16 a_n2140_13878.n14 11.9339
R21896 a_n2140_13878.n14 a_n2140_13878.n13 6.95632
R21897 a_n2140_13878.n15 a_n2140_13878.t6 3.61217
R21898 a_n2140_13878.n15 a_n2140_13878.t7 3.61217
R21899 a_n2140_13878.n17 a_n2140_13878.t13 3.61217
R21900 a_n2140_13878.n17 a_n2140_13878.t14 3.61217
R21901 a_n2140_13878.n19 a_n2140_13878.t0 3.61217
R21902 a_n2140_13878.n19 a_n2140_13878.t8 3.61217
R21903 a_n2140_13878.n11 a_n2140_13878.t22 3.61217
R21904 a_n2140_13878.n11 a_n2140_13878.t23 3.61217
R21905 a_n2140_13878.n7 a_n2140_13878.t20 3.61217
R21906 a_n2140_13878.n7 a_n2140_13878.t21 3.61217
R21907 a_n2140_13878.n5 a_n2140_13878.t9 3.61217
R21908 a_n2140_13878.n5 a_n2140_13878.t1 3.61217
R21909 a_n2140_13878.n3 a_n2140_13878.t12 3.61217
R21910 a_n2140_13878.n3 a_n2140_13878.t3 3.61217
R21911 a_n2140_13878.n1 a_n2140_13878.t2 3.61217
R21912 a_n2140_13878.n1 a_n2140_13878.t4 3.61217
R21913 a_n2140_13878.n0 a_n2140_13878.t10 3.61217
R21914 a_n2140_13878.n0 a_n2140_13878.t5 3.61217
R21915 a_n2140_13878.n21 a_n2140_13878.t11 3.61217
R21916 a_n2140_13878.t15 a_n2140_13878.n21 3.61217
R21917 a_n2140_13878.n9 a_n2140_13878.n8 0.358259
R21918 a_n2140_13878.n12 a_n2140_13878.n10 0.358259
R21919 a_n2140_13878.n13 a_n2140_13878.n12 0.358259
R21920 a_n2140_13878.n20 a_n2140_13878.n18 0.358259
R21921 a_n2140_13878.n18 a_n2140_13878.n16 0.358259
R21922 a_n2140_13878.n4 a_n2140_13878.n2 0.146627
R21923 a_n2140_13878.n6 a_n2140_13878.n4 0.146627
R21924 a_n2140_13878.n10 a_n2140_13878.n9 0.101793
R21925 commonsourceibias.n397 commonsourceibias.t184 222.032
R21926 commonsourceibias.n281 commonsourceibias.t134 222.032
R21927 commonsourceibias.n44 commonsourceibias.t26 222.032
R21928 commonsourceibias.n166 commonsourceibias.t140 222.032
R21929 commonsourceibias.n875 commonsourceibias.t191 222.032
R21930 commonsourceibias.n759 commonsourceibias.t98 222.032
R21931 commonsourceibias.n529 commonsourceibias.t68 222.032
R21932 commonsourceibias.n645 commonsourceibias.t177 222.032
R21933 commonsourceibias.n480 commonsourceibias.t183 207.983
R21934 commonsourceibias.n364 commonsourceibias.t88 207.983
R21935 commonsourceibias.n127 commonsourceibias.t16 207.983
R21936 commonsourceibias.n249 commonsourceibias.t151 207.983
R21937 commonsourceibias.n963 commonsourceibias.t101 207.983
R21938 commonsourceibias.n847 commonsourceibias.t189 207.983
R21939 commonsourceibias.n617 commonsourceibias.t40 207.983
R21940 commonsourceibias.n732 commonsourceibias.t112 207.983
R21941 commonsourceibias.n396 commonsourceibias.t150 168.701
R21942 commonsourceibias.n402 commonsourceibias.t155 168.701
R21943 commonsourceibias.n408 commonsourceibias.t199 168.701
R21944 commonsourceibias.n392 commonsourceibias.t175 168.701
R21945 commonsourceibias.n416 commonsourceibias.t165 168.701
R21946 commonsourceibias.n422 commonsourceibias.t96 168.701
R21947 commonsourceibias.n387 commonsourceibias.t187 168.701
R21948 commonsourceibias.n430 commonsourceibias.t168 168.701
R21949 commonsourceibias.n436 commonsourceibias.t172 168.701
R21950 commonsourceibias.n382 commonsourceibias.t80 168.701
R21951 commonsourceibias.n444 commonsourceibias.t173 168.701
R21952 commonsourceibias.n450 commonsourceibias.t182 168.701
R21953 commonsourceibias.n377 commonsourceibias.t149 168.701
R21954 commonsourceibias.n458 commonsourceibias.t110 168.701
R21955 commonsourceibias.n464 commonsourceibias.t194 168.701
R21956 commonsourceibias.n372 commonsourceibias.t157 168.701
R21957 commonsourceibias.n472 commonsourceibias.t163 168.701
R21958 commonsourceibias.n478 commonsourceibias.t92 168.701
R21959 commonsourceibias.n362 commonsourceibias.t198 168.701
R21960 commonsourceibias.n356 commonsourceibias.t186 168.701
R21961 commonsourceibias.n256 commonsourceibias.t95 168.701
R21962 commonsourceibias.n348 commonsourceibias.t196 168.701
R21963 commonsourceibias.n342 commonsourceibias.t105 168.701
R21964 commonsourceibias.n261 commonsourceibias.t94 168.701
R21965 commonsourceibias.n334 commonsourceibias.t197 168.701
R21966 commonsourceibias.n328 commonsourceibias.t115 168.701
R21967 commonsourceibias.n266 commonsourceibias.t141 168.701
R21968 commonsourceibias.n320 commonsourceibias.t195 168.701
R21969 commonsourceibias.n314 commonsourceibias.t113 168.701
R21970 commonsourceibias.n271 commonsourceibias.t138 168.701
R21971 commonsourceibias.n306 commonsourceibias.t130 168.701
R21972 commonsourceibias.n300 commonsourceibias.t114 168.701
R21973 commonsourceibias.n276 commonsourceibias.t139 168.701
R21974 commonsourceibias.n292 commonsourceibias.t129 168.701
R21975 commonsourceibias.n286 commonsourceibias.t125 168.701
R21976 commonsourceibias.n280 commonsourceibias.t147 168.701
R21977 commonsourceibias.n125 commonsourceibias.t60 168.701
R21978 commonsourceibias.n119 commonsourceibias.t4 168.701
R21979 commonsourceibias.n19 commonsourceibias.t14 168.701
R21980 commonsourceibias.n111 commonsourceibias.t74 168.701
R21981 commonsourceibias.n105 commonsourceibias.t20 168.701
R21982 commonsourceibias.n24 commonsourceibias.t34 168.701
R21983 commonsourceibias.n97 commonsourceibias.t10 168.701
R21984 commonsourceibias.n91 commonsourceibias.t18 168.701
R21985 commonsourceibias.n29 commonsourceibias.t54 168.701
R21986 commonsourceibias.n83 commonsourceibias.t30 168.701
R21987 commonsourceibias.n77 commonsourceibias.t36 168.701
R21988 commonsourceibias.n34 commonsourceibias.t70 168.701
R21989 commonsourceibias.n69 commonsourceibias.t22 168.701
R21990 commonsourceibias.n63 commonsourceibias.t62 168.701
R21991 commonsourceibias.n39 commonsourceibias.t0 168.701
R21992 commonsourceibias.n55 commonsourceibias.t42 168.701
R21993 commonsourceibias.n49 commonsourceibias.t52 168.701
R21994 commonsourceibias.n43 commonsourceibias.t58 168.701
R21995 commonsourceibias.n247 commonsourceibias.t83 168.701
R21996 commonsourceibias.n241 commonsourceibias.t161 168.701
R21997 commonsourceibias.n5 commonsourceibias.t152 168.701
R21998 commonsourceibias.n233 commonsourceibias.t171 168.701
R21999 commonsourceibias.n227 commonsourceibias.t145 168.701
R22000 commonsourceibias.n10 commonsourceibias.t124 168.701
R22001 commonsourceibias.n219 commonsourceibias.t158 168.701
R22002 commonsourceibias.n213 commonsourceibias.t148 168.701
R22003 commonsourceibias.n150 commonsourceibias.t93 168.701
R22004 commonsourceibias.n151 commonsourceibias.t131 168.701
R22005 commonsourceibias.n153 commonsourceibias.t117 168.701
R22006 commonsourceibias.n155 commonsourceibias.t176 168.701
R22007 commonsourceibias.n191 commonsourceibias.t144 168.701
R22008 commonsourceibias.n185 commonsourceibias.t190 168.701
R22009 commonsourceibias.n161 commonsourceibias.t164 168.701
R22010 commonsourceibias.n177 commonsourceibias.t111 168.701
R22011 commonsourceibias.n171 commonsourceibias.t100 168.701
R22012 commonsourceibias.n165 commonsourceibias.t84 168.701
R22013 commonsourceibias.n874 commonsourceibias.t156 168.701
R22014 commonsourceibias.n880 commonsourceibias.t146 168.701
R22015 commonsourceibias.n886 commonsourceibias.t126 168.701
R22016 commonsourceibias.n888 commonsourceibias.t91 168.701
R22017 commonsourceibias.n895 commonsourceibias.t181 168.701
R22018 commonsourceibias.n901 commonsourceibias.t136 168.701
R22019 commonsourceibias.n903 commonsourceibias.t107 168.701
R22020 commonsourceibias.n910 commonsourceibias.t192 168.701
R22021 commonsourceibias.n916 commonsourceibias.t167 168.701
R22022 commonsourceibias.n918 commonsourceibias.t127 168.701
R22023 commonsourceibias.n925 commonsourceibias.t87 168.701
R22024 commonsourceibias.n931 commonsourceibias.t99 168.701
R22025 commonsourceibias.n933 commonsourceibias.t137 168.701
R22026 commonsourceibias.n940 commonsourceibias.t143 168.701
R22027 commonsourceibias.n946 commonsourceibias.t122 168.701
R22028 commonsourceibias.n948 commonsourceibias.t170 168.701
R22029 commonsourceibias.n955 commonsourceibias.t153 168.701
R22030 commonsourceibias.n961 commonsourceibias.t133 168.701
R22031 commonsourceibias.n758 commonsourceibias.t123 168.701
R22032 commonsourceibias.n764 commonsourceibias.t132 168.701
R22033 commonsourceibias.n770 commonsourceibias.t104 168.701
R22034 commonsourceibias.n772 commonsourceibias.t118 168.701
R22035 commonsourceibias.n779 commonsourceibias.t85 168.701
R22036 commonsourceibias.n785 commonsourceibias.t106 168.701
R22037 commonsourceibias.n787 commonsourceibias.t119 168.701
R22038 commonsourceibias.n794 commonsourceibias.t86 168.701
R22039 commonsourceibias.n800 commonsourceibias.t97 168.701
R22040 commonsourceibias.n802 commonsourceibias.t120 168.701
R22041 commonsourceibias.n809 commonsourceibias.t89 168.701
R22042 commonsourceibias.n815 commonsourceibias.t178 168.701
R22043 commonsourceibias.n817 commonsourceibias.t121 168.701
R22044 commonsourceibias.n824 commonsourceibias.t81 168.701
R22045 commonsourceibias.n830 commonsourceibias.t179 168.701
R22046 commonsourceibias.n832 commonsourceibias.t193 168.701
R22047 commonsourceibias.n839 commonsourceibias.t82 168.701
R22048 commonsourceibias.n845 commonsourceibias.t180 168.701
R22049 commonsourceibias.n528 commonsourceibias.t8 168.701
R22050 commonsourceibias.n534 commonsourceibias.t6 168.701
R22051 commonsourceibias.n540 commonsourceibias.t66 168.701
R22052 commonsourceibias.n542 commonsourceibias.t28 168.701
R22053 commonsourceibias.n549 commonsourceibias.t78 168.701
R22054 commonsourceibias.n555 commonsourceibias.t48 168.701
R22055 commonsourceibias.n557 commonsourceibias.t2 168.701
R22056 commonsourceibias.n564 commonsourceibias.t64 168.701
R22057 commonsourceibias.n570 commonsourceibias.t50 168.701
R22058 commonsourceibias.n572 commonsourceibias.t72 168.701
R22059 commonsourceibias.n579 commonsourceibias.t44 168.701
R22060 commonsourceibias.n585 commonsourceibias.t32 168.701
R22061 commonsourceibias.n587 commonsourceibias.t56 168.701
R22062 commonsourceibias.n594 commonsourceibias.t46 168.701
R22063 commonsourceibias.n600 commonsourceibias.t12 168.701
R22064 commonsourceibias.n602 commonsourceibias.t38 168.701
R22065 commonsourceibias.n609 commonsourceibias.t24 168.701
R22066 commonsourceibias.n615 commonsourceibias.t76 168.701
R22067 commonsourceibias.n730 commonsourceibias.t169 168.701
R22068 commonsourceibias.n724 commonsourceibias.t142 168.701
R22069 commonsourceibias.n717 commonsourceibias.t116 168.701
R22070 commonsourceibias.n715 commonsourceibias.t154 168.701
R22071 commonsourceibias.n709 commonsourceibias.t108 168.701
R22072 commonsourceibias.n702 commonsourceibias.t90 168.701
R22073 commonsourceibias.n700 commonsourceibias.t128 168.701
R22074 commonsourceibias.n694 commonsourceibias.t109 168.701
R22075 commonsourceibias.n687 commonsourceibias.t174 168.701
R22076 commonsourceibias.n644 commonsourceibias.t159 168.701
R22077 commonsourceibias.n650 commonsourceibias.t160 168.701
R22078 commonsourceibias.n656 commonsourceibias.t185 168.701
R22079 commonsourceibias.n658 commonsourceibias.t135 168.701
R22080 commonsourceibias.n665 commonsourceibias.t166 168.701
R22081 commonsourceibias.n671 commonsourceibias.t103 168.701
R22082 commonsourceibias.n635 commonsourceibias.t162 168.701
R22083 commonsourceibias.n633 commonsourceibias.t188 168.701
R22084 commonsourceibias.n631 commonsourceibias.t102 168.701
R22085 commonsourceibias.n479 commonsourceibias.n367 161.3
R22086 commonsourceibias.n477 commonsourceibias.n476 161.3
R22087 commonsourceibias.n475 commonsourceibias.n368 161.3
R22088 commonsourceibias.n474 commonsourceibias.n473 161.3
R22089 commonsourceibias.n471 commonsourceibias.n369 161.3
R22090 commonsourceibias.n470 commonsourceibias.n469 161.3
R22091 commonsourceibias.n468 commonsourceibias.n370 161.3
R22092 commonsourceibias.n467 commonsourceibias.n466 161.3
R22093 commonsourceibias.n465 commonsourceibias.n371 161.3
R22094 commonsourceibias.n463 commonsourceibias.n462 161.3
R22095 commonsourceibias.n461 commonsourceibias.n373 161.3
R22096 commonsourceibias.n460 commonsourceibias.n459 161.3
R22097 commonsourceibias.n457 commonsourceibias.n374 161.3
R22098 commonsourceibias.n456 commonsourceibias.n455 161.3
R22099 commonsourceibias.n454 commonsourceibias.n375 161.3
R22100 commonsourceibias.n453 commonsourceibias.n452 161.3
R22101 commonsourceibias.n451 commonsourceibias.n376 161.3
R22102 commonsourceibias.n449 commonsourceibias.n448 161.3
R22103 commonsourceibias.n447 commonsourceibias.n378 161.3
R22104 commonsourceibias.n446 commonsourceibias.n445 161.3
R22105 commonsourceibias.n443 commonsourceibias.n379 161.3
R22106 commonsourceibias.n442 commonsourceibias.n441 161.3
R22107 commonsourceibias.n440 commonsourceibias.n380 161.3
R22108 commonsourceibias.n439 commonsourceibias.n438 161.3
R22109 commonsourceibias.n437 commonsourceibias.n381 161.3
R22110 commonsourceibias.n435 commonsourceibias.n434 161.3
R22111 commonsourceibias.n433 commonsourceibias.n383 161.3
R22112 commonsourceibias.n432 commonsourceibias.n431 161.3
R22113 commonsourceibias.n429 commonsourceibias.n384 161.3
R22114 commonsourceibias.n428 commonsourceibias.n427 161.3
R22115 commonsourceibias.n426 commonsourceibias.n385 161.3
R22116 commonsourceibias.n425 commonsourceibias.n424 161.3
R22117 commonsourceibias.n423 commonsourceibias.n386 161.3
R22118 commonsourceibias.n421 commonsourceibias.n420 161.3
R22119 commonsourceibias.n419 commonsourceibias.n388 161.3
R22120 commonsourceibias.n418 commonsourceibias.n417 161.3
R22121 commonsourceibias.n415 commonsourceibias.n389 161.3
R22122 commonsourceibias.n414 commonsourceibias.n413 161.3
R22123 commonsourceibias.n412 commonsourceibias.n390 161.3
R22124 commonsourceibias.n411 commonsourceibias.n410 161.3
R22125 commonsourceibias.n409 commonsourceibias.n391 161.3
R22126 commonsourceibias.n407 commonsourceibias.n406 161.3
R22127 commonsourceibias.n405 commonsourceibias.n393 161.3
R22128 commonsourceibias.n404 commonsourceibias.n403 161.3
R22129 commonsourceibias.n401 commonsourceibias.n394 161.3
R22130 commonsourceibias.n400 commonsourceibias.n399 161.3
R22131 commonsourceibias.n398 commonsourceibias.n395 161.3
R22132 commonsourceibias.n282 commonsourceibias.n279 161.3
R22133 commonsourceibias.n284 commonsourceibias.n283 161.3
R22134 commonsourceibias.n285 commonsourceibias.n278 161.3
R22135 commonsourceibias.n288 commonsourceibias.n287 161.3
R22136 commonsourceibias.n289 commonsourceibias.n277 161.3
R22137 commonsourceibias.n291 commonsourceibias.n290 161.3
R22138 commonsourceibias.n293 commonsourceibias.n275 161.3
R22139 commonsourceibias.n295 commonsourceibias.n294 161.3
R22140 commonsourceibias.n296 commonsourceibias.n274 161.3
R22141 commonsourceibias.n298 commonsourceibias.n297 161.3
R22142 commonsourceibias.n299 commonsourceibias.n273 161.3
R22143 commonsourceibias.n302 commonsourceibias.n301 161.3
R22144 commonsourceibias.n303 commonsourceibias.n272 161.3
R22145 commonsourceibias.n305 commonsourceibias.n304 161.3
R22146 commonsourceibias.n307 commonsourceibias.n270 161.3
R22147 commonsourceibias.n309 commonsourceibias.n308 161.3
R22148 commonsourceibias.n310 commonsourceibias.n269 161.3
R22149 commonsourceibias.n312 commonsourceibias.n311 161.3
R22150 commonsourceibias.n313 commonsourceibias.n268 161.3
R22151 commonsourceibias.n316 commonsourceibias.n315 161.3
R22152 commonsourceibias.n317 commonsourceibias.n267 161.3
R22153 commonsourceibias.n319 commonsourceibias.n318 161.3
R22154 commonsourceibias.n321 commonsourceibias.n265 161.3
R22155 commonsourceibias.n323 commonsourceibias.n322 161.3
R22156 commonsourceibias.n324 commonsourceibias.n264 161.3
R22157 commonsourceibias.n326 commonsourceibias.n325 161.3
R22158 commonsourceibias.n327 commonsourceibias.n263 161.3
R22159 commonsourceibias.n330 commonsourceibias.n329 161.3
R22160 commonsourceibias.n331 commonsourceibias.n262 161.3
R22161 commonsourceibias.n333 commonsourceibias.n332 161.3
R22162 commonsourceibias.n335 commonsourceibias.n260 161.3
R22163 commonsourceibias.n337 commonsourceibias.n336 161.3
R22164 commonsourceibias.n338 commonsourceibias.n259 161.3
R22165 commonsourceibias.n340 commonsourceibias.n339 161.3
R22166 commonsourceibias.n341 commonsourceibias.n258 161.3
R22167 commonsourceibias.n344 commonsourceibias.n343 161.3
R22168 commonsourceibias.n345 commonsourceibias.n257 161.3
R22169 commonsourceibias.n347 commonsourceibias.n346 161.3
R22170 commonsourceibias.n349 commonsourceibias.n255 161.3
R22171 commonsourceibias.n351 commonsourceibias.n350 161.3
R22172 commonsourceibias.n352 commonsourceibias.n254 161.3
R22173 commonsourceibias.n354 commonsourceibias.n353 161.3
R22174 commonsourceibias.n355 commonsourceibias.n253 161.3
R22175 commonsourceibias.n358 commonsourceibias.n357 161.3
R22176 commonsourceibias.n359 commonsourceibias.n252 161.3
R22177 commonsourceibias.n361 commonsourceibias.n360 161.3
R22178 commonsourceibias.n363 commonsourceibias.n251 161.3
R22179 commonsourceibias.n45 commonsourceibias.n42 161.3
R22180 commonsourceibias.n47 commonsourceibias.n46 161.3
R22181 commonsourceibias.n48 commonsourceibias.n41 161.3
R22182 commonsourceibias.n51 commonsourceibias.n50 161.3
R22183 commonsourceibias.n52 commonsourceibias.n40 161.3
R22184 commonsourceibias.n54 commonsourceibias.n53 161.3
R22185 commonsourceibias.n56 commonsourceibias.n38 161.3
R22186 commonsourceibias.n58 commonsourceibias.n57 161.3
R22187 commonsourceibias.n59 commonsourceibias.n37 161.3
R22188 commonsourceibias.n61 commonsourceibias.n60 161.3
R22189 commonsourceibias.n62 commonsourceibias.n36 161.3
R22190 commonsourceibias.n65 commonsourceibias.n64 161.3
R22191 commonsourceibias.n66 commonsourceibias.n35 161.3
R22192 commonsourceibias.n68 commonsourceibias.n67 161.3
R22193 commonsourceibias.n70 commonsourceibias.n33 161.3
R22194 commonsourceibias.n72 commonsourceibias.n71 161.3
R22195 commonsourceibias.n73 commonsourceibias.n32 161.3
R22196 commonsourceibias.n75 commonsourceibias.n74 161.3
R22197 commonsourceibias.n76 commonsourceibias.n31 161.3
R22198 commonsourceibias.n79 commonsourceibias.n78 161.3
R22199 commonsourceibias.n80 commonsourceibias.n30 161.3
R22200 commonsourceibias.n82 commonsourceibias.n81 161.3
R22201 commonsourceibias.n84 commonsourceibias.n28 161.3
R22202 commonsourceibias.n86 commonsourceibias.n85 161.3
R22203 commonsourceibias.n87 commonsourceibias.n27 161.3
R22204 commonsourceibias.n89 commonsourceibias.n88 161.3
R22205 commonsourceibias.n90 commonsourceibias.n26 161.3
R22206 commonsourceibias.n93 commonsourceibias.n92 161.3
R22207 commonsourceibias.n94 commonsourceibias.n25 161.3
R22208 commonsourceibias.n96 commonsourceibias.n95 161.3
R22209 commonsourceibias.n98 commonsourceibias.n23 161.3
R22210 commonsourceibias.n100 commonsourceibias.n99 161.3
R22211 commonsourceibias.n101 commonsourceibias.n22 161.3
R22212 commonsourceibias.n103 commonsourceibias.n102 161.3
R22213 commonsourceibias.n104 commonsourceibias.n21 161.3
R22214 commonsourceibias.n107 commonsourceibias.n106 161.3
R22215 commonsourceibias.n108 commonsourceibias.n20 161.3
R22216 commonsourceibias.n110 commonsourceibias.n109 161.3
R22217 commonsourceibias.n112 commonsourceibias.n18 161.3
R22218 commonsourceibias.n114 commonsourceibias.n113 161.3
R22219 commonsourceibias.n115 commonsourceibias.n17 161.3
R22220 commonsourceibias.n117 commonsourceibias.n116 161.3
R22221 commonsourceibias.n118 commonsourceibias.n16 161.3
R22222 commonsourceibias.n121 commonsourceibias.n120 161.3
R22223 commonsourceibias.n122 commonsourceibias.n15 161.3
R22224 commonsourceibias.n124 commonsourceibias.n123 161.3
R22225 commonsourceibias.n126 commonsourceibias.n14 161.3
R22226 commonsourceibias.n167 commonsourceibias.n164 161.3
R22227 commonsourceibias.n169 commonsourceibias.n168 161.3
R22228 commonsourceibias.n170 commonsourceibias.n163 161.3
R22229 commonsourceibias.n173 commonsourceibias.n172 161.3
R22230 commonsourceibias.n174 commonsourceibias.n162 161.3
R22231 commonsourceibias.n176 commonsourceibias.n175 161.3
R22232 commonsourceibias.n178 commonsourceibias.n160 161.3
R22233 commonsourceibias.n180 commonsourceibias.n179 161.3
R22234 commonsourceibias.n181 commonsourceibias.n159 161.3
R22235 commonsourceibias.n183 commonsourceibias.n182 161.3
R22236 commonsourceibias.n184 commonsourceibias.n158 161.3
R22237 commonsourceibias.n187 commonsourceibias.n186 161.3
R22238 commonsourceibias.n188 commonsourceibias.n157 161.3
R22239 commonsourceibias.n190 commonsourceibias.n189 161.3
R22240 commonsourceibias.n192 commonsourceibias.n156 161.3
R22241 commonsourceibias.n194 commonsourceibias.n193 161.3
R22242 commonsourceibias.n196 commonsourceibias.n195 161.3
R22243 commonsourceibias.n197 commonsourceibias.n154 161.3
R22244 commonsourceibias.n199 commonsourceibias.n198 161.3
R22245 commonsourceibias.n201 commonsourceibias.n200 161.3
R22246 commonsourceibias.n202 commonsourceibias.n152 161.3
R22247 commonsourceibias.n204 commonsourceibias.n203 161.3
R22248 commonsourceibias.n206 commonsourceibias.n205 161.3
R22249 commonsourceibias.n208 commonsourceibias.n207 161.3
R22250 commonsourceibias.n209 commonsourceibias.n13 161.3
R22251 commonsourceibias.n211 commonsourceibias.n210 161.3
R22252 commonsourceibias.n212 commonsourceibias.n12 161.3
R22253 commonsourceibias.n215 commonsourceibias.n214 161.3
R22254 commonsourceibias.n216 commonsourceibias.n11 161.3
R22255 commonsourceibias.n218 commonsourceibias.n217 161.3
R22256 commonsourceibias.n220 commonsourceibias.n9 161.3
R22257 commonsourceibias.n222 commonsourceibias.n221 161.3
R22258 commonsourceibias.n223 commonsourceibias.n8 161.3
R22259 commonsourceibias.n225 commonsourceibias.n224 161.3
R22260 commonsourceibias.n226 commonsourceibias.n7 161.3
R22261 commonsourceibias.n229 commonsourceibias.n228 161.3
R22262 commonsourceibias.n230 commonsourceibias.n6 161.3
R22263 commonsourceibias.n232 commonsourceibias.n231 161.3
R22264 commonsourceibias.n234 commonsourceibias.n4 161.3
R22265 commonsourceibias.n236 commonsourceibias.n235 161.3
R22266 commonsourceibias.n237 commonsourceibias.n3 161.3
R22267 commonsourceibias.n239 commonsourceibias.n238 161.3
R22268 commonsourceibias.n240 commonsourceibias.n2 161.3
R22269 commonsourceibias.n243 commonsourceibias.n242 161.3
R22270 commonsourceibias.n244 commonsourceibias.n1 161.3
R22271 commonsourceibias.n246 commonsourceibias.n245 161.3
R22272 commonsourceibias.n248 commonsourceibias.n0 161.3
R22273 commonsourceibias.n962 commonsourceibias.n850 161.3
R22274 commonsourceibias.n960 commonsourceibias.n959 161.3
R22275 commonsourceibias.n958 commonsourceibias.n851 161.3
R22276 commonsourceibias.n957 commonsourceibias.n956 161.3
R22277 commonsourceibias.n954 commonsourceibias.n852 161.3
R22278 commonsourceibias.n953 commonsourceibias.n952 161.3
R22279 commonsourceibias.n951 commonsourceibias.n853 161.3
R22280 commonsourceibias.n950 commonsourceibias.n949 161.3
R22281 commonsourceibias.n947 commonsourceibias.n854 161.3
R22282 commonsourceibias.n945 commonsourceibias.n944 161.3
R22283 commonsourceibias.n943 commonsourceibias.n855 161.3
R22284 commonsourceibias.n942 commonsourceibias.n941 161.3
R22285 commonsourceibias.n939 commonsourceibias.n856 161.3
R22286 commonsourceibias.n938 commonsourceibias.n937 161.3
R22287 commonsourceibias.n936 commonsourceibias.n857 161.3
R22288 commonsourceibias.n935 commonsourceibias.n934 161.3
R22289 commonsourceibias.n932 commonsourceibias.n858 161.3
R22290 commonsourceibias.n930 commonsourceibias.n929 161.3
R22291 commonsourceibias.n928 commonsourceibias.n859 161.3
R22292 commonsourceibias.n927 commonsourceibias.n926 161.3
R22293 commonsourceibias.n924 commonsourceibias.n860 161.3
R22294 commonsourceibias.n923 commonsourceibias.n922 161.3
R22295 commonsourceibias.n921 commonsourceibias.n861 161.3
R22296 commonsourceibias.n920 commonsourceibias.n919 161.3
R22297 commonsourceibias.n917 commonsourceibias.n862 161.3
R22298 commonsourceibias.n915 commonsourceibias.n914 161.3
R22299 commonsourceibias.n913 commonsourceibias.n863 161.3
R22300 commonsourceibias.n912 commonsourceibias.n911 161.3
R22301 commonsourceibias.n909 commonsourceibias.n864 161.3
R22302 commonsourceibias.n908 commonsourceibias.n907 161.3
R22303 commonsourceibias.n906 commonsourceibias.n865 161.3
R22304 commonsourceibias.n905 commonsourceibias.n904 161.3
R22305 commonsourceibias.n902 commonsourceibias.n866 161.3
R22306 commonsourceibias.n900 commonsourceibias.n899 161.3
R22307 commonsourceibias.n898 commonsourceibias.n867 161.3
R22308 commonsourceibias.n897 commonsourceibias.n896 161.3
R22309 commonsourceibias.n894 commonsourceibias.n868 161.3
R22310 commonsourceibias.n893 commonsourceibias.n892 161.3
R22311 commonsourceibias.n891 commonsourceibias.n869 161.3
R22312 commonsourceibias.n890 commonsourceibias.n889 161.3
R22313 commonsourceibias.n887 commonsourceibias.n870 161.3
R22314 commonsourceibias.n885 commonsourceibias.n884 161.3
R22315 commonsourceibias.n883 commonsourceibias.n871 161.3
R22316 commonsourceibias.n882 commonsourceibias.n881 161.3
R22317 commonsourceibias.n879 commonsourceibias.n872 161.3
R22318 commonsourceibias.n878 commonsourceibias.n877 161.3
R22319 commonsourceibias.n876 commonsourceibias.n873 161.3
R22320 commonsourceibias.n846 commonsourceibias.n734 161.3
R22321 commonsourceibias.n844 commonsourceibias.n843 161.3
R22322 commonsourceibias.n842 commonsourceibias.n735 161.3
R22323 commonsourceibias.n841 commonsourceibias.n840 161.3
R22324 commonsourceibias.n838 commonsourceibias.n736 161.3
R22325 commonsourceibias.n837 commonsourceibias.n836 161.3
R22326 commonsourceibias.n835 commonsourceibias.n737 161.3
R22327 commonsourceibias.n834 commonsourceibias.n833 161.3
R22328 commonsourceibias.n831 commonsourceibias.n738 161.3
R22329 commonsourceibias.n829 commonsourceibias.n828 161.3
R22330 commonsourceibias.n827 commonsourceibias.n739 161.3
R22331 commonsourceibias.n826 commonsourceibias.n825 161.3
R22332 commonsourceibias.n823 commonsourceibias.n740 161.3
R22333 commonsourceibias.n822 commonsourceibias.n821 161.3
R22334 commonsourceibias.n820 commonsourceibias.n741 161.3
R22335 commonsourceibias.n819 commonsourceibias.n818 161.3
R22336 commonsourceibias.n816 commonsourceibias.n742 161.3
R22337 commonsourceibias.n814 commonsourceibias.n813 161.3
R22338 commonsourceibias.n812 commonsourceibias.n743 161.3
R22339 commonsourceibias.n811 commonsourceibias.n810 161.3
R22340 commonsourceibias.n808 commonsourceibias.n744 161.3
R22341 commonsourceibias.n807 commonsourceibias.n806 161.3
R22342 commonsourceibias.n805 commonsourceibias.n745 161.3
R22343 commonsourceibias.n804 commonsourceibias.n803 161.3
R22344 commonsourceibias.n801 commonsourceibias.n746 161.3
R22345 commonsourceibias.n799 commonsourceibias.n798 161.3
R22346 commonsourceibias.n797 commonsourceibias.n747 161.3
R22347 commonsourceibias.n796 commonsourceibias.n795 161.3
R22348 commonsourceibias.n793 commonsourceibias.n748 161.3
R22349 commonsourceibias.n792 commonsourceibias.n791 161.3
R22350 commonsourceibias.n790 commonsourceibias.n749 161.3
R22351 commonsourceibias.n789 commonsourceibias.n788 161.3
R22352 commonsourceibias.n786 commonsourceibias.n750 161.3
R22353 commonsourceibias.n784 commonsourceibias.n783 161.3
R22354 commonsourceibias.n782 commonsourceibias.n751 161.3
R22355 commonsourceibias.n781 commonsourceibias.n780 161.3
R22356 commonsourceibias.n778 commonsourceibias.n752 161.3
R22357 commonsourceibias.n777 commonsourceibias.n776 161.3
R22358 commonsourceibias.n775 commonsourceibias.n753 161.3
R22359 commonsourceibias.n774 commonsourceibias.n773 161.3
R22360 commonsourceibias.n771 commonsourceibias.n754 161.3
R22361 commonsourceibias.n769 commonsourceibias.n768 161.3
R22362 commonsourceibias.n767 commonsourceibias.n755 161.3
R22363 commonsourceibias.n766 commonsourceibias.n765 161.3
R22364 commonsourceibias.n763 commonsourceibias.n756 161.3
R22365 commonsourceibias.n762 commonsourceibias.n761 161.3
R22366 commonsourceibias.n760 commonsourceibias.n757 161.3
R22367 commonsourceibias.n616 commonsourceibias.n504 161.3
R22368 commonsourceibias.n614 commonsourceibias.n613 161.3
R22369 commonsourceibias.n612 commonsourceibias.n505 161.3
R22370 commonsourceibias.n611 commonsourceibias.n610 161.3
R22371 commonsourceibias.n608 commonsourceibias.n506 161.3
R22372 commonsourceibias.n607 commonsourceibias.n606 161.3
R22373 commonsourceibias.n605 commonsourceibias.n507 161.3
R22374 commonsourceibias.n604 commonsourceibias.n603 161.3
R22375 commonsourceibias.n601 commonsourceibias.n508 161.3
R22376 commonsourceibias.n599 commonsourceibias.n598 161.3
R22377 commonsourceibias.n597 commonsourceibias.n509 161.3
R22378 commonsourceibias.n596 commonsourceibias.n595 161.3
R22379 commonsourceibias.n593 commonsourceibias.n510 161.3
R22380 commonsourceibias.n592 commonsourceibias.n591 161.3
R22381 commonsourceibias.n590 commonsourceibias.n511 161.3
R22382 commonsourceibias.n589 commonsourceibias.n588 161.3
R22383 commonsourceibias.n586 commonsourceibias.n512 161.3
R22384 commonsourceibias.n584 commonsourceibias.n583 161.3
R22385 commonsourceibias.n582 commonsourceibias.n513 161.3
R22386 commonsourceibias.n581 commonsourceibias.n580 161.3
R22387 commonsourceibias.n578 commonsourceibias.n514 161.3
R22388 commonsourceibias.n577 commonsourceibias.n576 161.3
R22389 commonsourceibias.n575 commonsourceibias.n515 161.3
R22390 commonsourceibias.n574 commonsourceibias.n573 161.3
R22391 commonsourceibias.n571 commonsourceibias.n516 161.3
R22392 commonsourceibias.n569 commonsourceibias.n568 161.3
R22393 commonsourceibias.n567 commonsourceibias.n517 161.3
R22394 commonsourceibias.n566 commonsourceibias.n565 161.3
R22395 commonsourceibias.n563 commonsourceibias.n518 161.3
R22396 commonsourceibias.n562 commonsourceibias.n561 161.3
R22397 commonsourceibias.n560 commonsourceibias.n519 161.3
R22398 commonsourceibias.n559 commonsourceibias.n558 161.3
R22399 commonsourceibias.n556 commonsourceibias.n520 161.3
R22400 commonsourceibias.n554 commonsourceibias.n553 161.3
R22401 commonsourceibias.n552 commonsourceibias.n521 161.3
R22402 commonsourceibias.n551 commonsourceibias.n550 161.3
R22403 commonsourceibias.n548 commonsourceibias.n522 161.3
R22404 commonsourceibias.n547 commonsourceibias.n546 161.3
R22405 commonsourceibias.n545 commonsourceibias.n523 161.3
R22406 commonsourceibias.n544 commonsourceibias.n543 161.3
R22407 commonsourceibias.n541 commonsourceibias.n524 161.3
R22408 commonsourceibias.n539 commonsourceibias.n538 161.3
R22409 commonsourceibias.n537 commonsourceibias.n525 161.3
R22410 commonsourceibias.n536 commonsourceibias.n535 161.3
R22411 commonsourceibias.n533 commonsourceibias.n526 161.3
R22412 commonsourceibias.n532 commonsourceibias.n531 161.3
R22413 commonsourceibias.n530 commonsourceibias.n527 161.3
R22414 commonsourceibias.n686 commonsourceibias.n685 161.3
R22415 commonsourceibias.n684 commonsourceibias.n683 161.3
R22416 commonsourceibias.n682 commonsourceibias.n632 161.3
R22417 commonsourceibias.n681 commonsourceibias.n680 161.3
R22418 commonsourceibias.n679 commonsourceibias.n678 161.3
R22419 commonsourceibias.n677 commonsourceibias.n634 161.3
R22420 commonsourceibias.n676 commonsourceibias.n675 161.3
R22421 commonsourceibias.n674 commonsourceibias.n673 161.3
R22422 commonsourceibias.n672 commonsourceibias.n636 161.3
R22423 commonsourceibias.n670 commonsourceibias.n669 161.3
R22424 commonsourceibias.n668 commonsourceibias.n637 161.3
R22425 commonsourceibias.n667 commonsourceibias.n666 161.3
R22426 commonsourceibias.n664 commonsourceibias.n638 161.3
R22427 commonsourceibias.n663 commonsourceibias.n662 161.3
R22428 commonsourceibias.n661 commonsourceibias.n639 161.3
R22429 commonsourceibias.n660 commonsourceibias.n659 161.3
R22430 commonsourceibias.n657 commonsourceibias.n640 161.3
R22431 commonsourceibias.n655 commonsourceibias.n654 161.3
R22432 commonsourceibias.n653 commonsourceibias.n641 161.3
R22433 commonsourceibias.n652 commonsourceibias.n651 161.3
R22434 commonsourceibias.n649 commonsourceibias.n642 161.3
R22435 commonsourceibias.n648 commonsourceibias.n647 161.3
R22436 commonsourceibias.n646 commonsourceibias.n643 161.3
R22437 commonsourceibias.n731 commonsourceibias.n483 161.3
R22438 commonsourceibias.n729 commonsourceibias.n728 161.3
R22439 commonsourceibias.n727 commonsourceibias.n484 161.3
R22440 commonsourceibias.n726 commonsourceibias.n725 161.3
R22441 commonsourceibias.n723 commonsourceibias.n485 161.3
R22442 commonsourceibias.n722 commonsourceibias.n721 161.3
R22443 commonsourceibias.n720 commonsourceibias.n486 161.3
R22444 commonsourceibias.n719 commonsourceibias.n718 161.3
R22445 commonsourceibias.n716 commonsourceibias.n487 161.3
R22446 commonsourceibias.n714 commonsourceibias.n713 161.3
R22447 commonsourceibias.n712 commonsourceibias.n488 161.3
R22448 commonsourceibias.n711 commonsourceibias.n710 161.3
R22449 commonsourceibias.n708 commonsourceibias.n489 161.3
R22450 commonsourceibias.n707 commonsourceibias.n706 161.3
R22451 commonsourceibias.n705 commonsourceibias.n490 161.3
R22452 commonsourceibias.n704 commonsourceibias.n703 161.3
R22453 commonsourceibias.n701 commonsourceibias.n491 161.3
R22454 commonsourceibias.n699 commonsourceibias.n698 161.3
R22455 commonsourceibias.n697 commonsourceibias.n492 161.3
R22456 commonsourceibias.n696 commonsourceibias.n695 161.3
R22457 commonsourceibias.n693 commonsourceibias.n493 161.3
R22458 commonsourceibias.n692 commonsourceibias.n691 161.3
R22459 commonsourceibias.n690 commonsourceibias.n494 161.3
R22460 commonsourceibias.n689 commonsourceibias.n688 161.3
R22461 commonsourceibias.n141 commonsourceibias.n139 81.5057
R22462 commonsourceibias.n497 commonsourceibias.n495 81.5057
R22463 commonsourceibias.n141 commonsourceibias.n140 80.9324
R22464 commonsourceibias.n143 commonsourceibias.n142 80.9324
R22465 commonsourceibias.n145 commonsourceibias.n144 80.9324
R22466 commonsourceibias.n147 commonsourceibias.n146 80.9324
R22467 commonsourceibias.n138 commonsourceibias.n137 80.9324
R22468 commonsourceibias.n136 commonsourceibias.n135 80.9324
R22469 commonsourceibias.n134 commonsourceibias.n133 80.9324
R22470 commonsourceibias.n132 commonsourceibias.n131 80.9324
R22471 commonsourceibias.n130 commonsourceibias.n129 80.9324
R22472 commonsourceibias.n620 commonsourceibias.n619 80.9324
R22473 commonsourceibias.n622 commonsourceibias.n621 80.9324
R22474 commonsourceibias.n624 commonsourceibias.n623 80.9324
R22475 commonsourceibias.n626 commonsourceibias.n625 80.9324
R22476 commonsourceibias.n628 commonsourceibias.n627 80.9324
R22477 commonsourceibias.n503 commonsourceibias.n502 80.9324
R22478 commonsourceibias.n501 commonsourceibias.n500 80.9324
R22479 commonsourceibias.n499 commonsourceibias.n498 80.9324
R22480 commonsourceibias.n497 commonsourceibias.n496 80.9324
R22481 commonsourceibias.n481 commonsourceibias.n480 80.6037
R22482 commonsourceibias.n365 commonsourceibias.n364 80.6037
R22483 commonsourceibias.n128 commonsourceibias.n127 80.6037
R22484 commonsourceibias.n250 commonsourceibias.n249 80.6037
R22485 commonsourceibias.n964 commonsourceibias.n963 80.6037
R22486 commonsourceibias.n848 commonsourceibias.n847 80.6037
R22487 commonsourceibias.n618 commonsourceibias.n617 80.6037
R22488 commonsourceibias.n733 commonsourceibias.n732 80.6037
R22489 commonsourceibias.n438 commonsourceibias.n437 56.5617
R22490 commonsourceibias.n452 commonsourceibias.n451 56.5617
R22491 commonsourceibias.n322 commonsourceibias.n321 56.5617
R22492 commonsourceibias.n308 commonsourceibias.n307 56.5617
R22493 commonsourceibias.n85 commonsourceibias.n84 56.5617
R22494 commonsourceibias.n71 commonsourceibias.n70 56.5617
R22495 commonsourceibias.n207 commonsourceibias.n206 56.5617
R22496 commonsourceibias.n193 commonsourceibias.n192 56.5617
R22497 commonsourceibias.n919 commonsourceibias.n917 56.5617
R22498 commonsourceibias.n934 commonsourceibias.n932 56.5617
R22499 commonsourceibias.n803 commonsourceibias.n801 56.5617
R22500 commonsourceibias.n818 commonsourceibias.n816 56.5617
R22501 commonsourceibias.n573 commonsourceibias.n571 56.5617
R22502 commonsourceibias.n588 commonsourceibias.n586 56.5617
R22503 commonsourceibias.n688 commonsourceibias.n686 56.5617
R22504 commonsourceibias.n410 commonsourceibias.n409 56.5617
R22505 commonsourceibias.n424 commonsourceibias.n423 56.5617
R22506 commonsourceibias.n466 commonsourceibias.n465 56.5617
R22507 commonsourceibias.n350 commonsourceibias.n349 56.5617
R22508 commonsourceibias.n336 commonsourceibias.n335 56.5617
R22509 commonsourceibias.n294 commonsourceibias.n293 56.5617
R22510 commonsourceibias.n113 commonsourceibias.n112 56.5617
R22511 commonsourceibias.n99 commonsourceibias.n98 56.5617
R22512 commonsourceibias.n57 commonsourceibias.n56 56.5617
R22513 commonsourceibias.n235 commonsourceibias.n234 56.5617
R22514 commonsourceibias.n221 commonsourceibias.n220 56.5617
R22515 commonsourceibias.n179 commonsourceibias.n178 56.5617
R22516 commonsourceibias.n889 commonsourceibias.n887 56.5617
R22517 commonsourceibias.n904 commonsourceibias.n902 56.5617
R22518 commonsourceibias.n949 commonsourceibias.n947 56.5617
R22519 commonsourceibias.n773 commonsourceibias.n771 56.5617
R22520 commonsourceibias.n788 commonsourceibias.n786 56.5617
R22521 commonsourceibias.n833 commonsourceibias.n831 56.5617
R22522 commonsourceibias.n543 commonsourceibias.n541 56.5617
R22523 commonsourceibias.n558 commonsourceibias.n556 56.5617
R22524 commonsourceibias.n603 commonsourceibias.n601 56.5617
R22525 commonsourceibias.n718 commonsourceibias.n716 56.5617
R22526 commonsourceibias.n703 commonsourceibias.n701 56.5617
R22527 commonsourceibias.n659 commonsourceibias.n657 56.5617
R22528 commonsourceibias.n673 commonsourceibias.n672 56.5617
R22529 commonsourceibias.n401 commonsourceibias.n400 51.2335
R22530 commonsourceibias.n473 commonsourceibias.n368 51.2335
R22531 commonsourceibias.n357 commonsourceibias.n252 51.2335
R22532 commonsourceibias.n285 commonsourceibias.n284 51.2335
R22533 commonsourceibias.n120 commonsourceibias.n15 51.2335
R22534 commonsourceibias.n48 commonsourceibias.n47 51.2335
R22535 commonsourceibias.n242 commonsourceibias.n1 51.2335
R22536 commonsourceibias.n170 commonsourceibias.n169 51.2335
R22537 commonsourceibias.n879 commonsourceibias.n878 51.2335
R22538 commonsourceibias.n956 commonsourceibias.n851 51.2335
R22539 commonsourceibias.n763 commonsourceibias.n762 51.2335
R22540 commonsourceibias.n840 commonsourceibias.n735 51.2335
R22541 commonsourceibias.n533 commonsourceibias.n532 51.2335
R22542 commonsourceibias.n610 commonsourceibias.n505 51.2335
R22543 commonsourceibias.n725 commonsourceibias.n484 51.2335
R22544 commonsourceibias.n649 commonsourceibias.n648 51.2335
R22545 commonsourceibias.n480 commonsourceibias.n479 50.9056
R22546 commonsourceibias.n364 commonsourceibias.n363 50.9056
R22547 commonsourceibias.n127 commonsourceibias.n126 50.9056
R22548 commonsourceibias.n249 commonsourceibias.n248 50.9056
R22549 commonsourceibias.n963 commonsourceibias.n962 50.9056
R22550 commonsourceibias.n847 commonsourceibias.n846 50.9056
R22551 commonsourceibias.n617 commonsourceibias.n616 50.9056
R22552 commonsourceibias.n732 commonsourceibias.n731 50.9056
R22553 commonsourceibias.n415 commonsourceibias.n414 50.2647
R22554 commonsourceibias.n459 commonsourceibias.n373 50.2647
R22555 commonsourceibias.n343 commonsourceibias.n257 50.2647
R22556 commonsourceibias.n299 commonsourceibias.n298 50.2647
R22557 commonsourceibias.n106 commonsourceibias.n20 50.2647
R22558 commonsourceibias.n62 commonsourceibias.n61 50.2647
R22559 commonsourceibias.n228 commonsourceibias.n6 50.2647
R22560 commonsourceibias.n184 commonsourceibias.n183 50.2647
R22561 commonsourceibias.n894 commonsourceibias.n893 50.2647
R22562 commonsourceibias.n941 commonsourceibias.n855 50.2647
R22563 commonsourceibias.n778 commonsourceibias.n777 50.2647
R22564 commonsourceibias.n825 commonsourceibias.n739 50.2647
R22565 commonsourceibias.n548 commonsourceibias.n547 50.2647
R22566 commonsourceibias.n595 commonsourceibias.n509 50.2647
R22567 commonsourceibias.n710 commonsourceibias.n488 50.2647
R22568 commonsourceibias.n664 commonsourceibias.n663 50.2647
R22569 commonsourceibias.n397 commonsourceibias.n396 49.9027
R22570 commonsourceibias.n281 commonsourceibias.n280 49.9027
R22571 commonsourceibias.n44 commonsourceibias.n43 49.9027
R22572 commonsourceibias.n166 commonsourceibias.n165 49.9027
R22573 commonsourceibias.n875 commonsourceibias.n874 49.9027
R22574 commonsourceibias.n759 commonsourceibias.n758 49.9027
R22575 commonsourceibias.n529 commonsourceibias.n528 49.9027
R22576 commonsourceibias.n645 commonsourceibias.n644 49.9027
R22577 commonsourceibias.n429 commonsourceibias.n428 49.296
R22578 commonsourceibias.n445 commonsourceibias.n378 49.296
R22579 commonsourceibias.n329 commonsourceibias.n262 49.296
R22580 commonsourceibias.n313 commonsourceibias.n312 49.296
R22581 commonsourceibias.n92 commonsourceibias.n25 49.296
R22582 commonsourceibias.n76 commonsourceibias.n75 49.296
R22583 commonsourceibias.n214 commonsourceibias.n11 49.296
R22584 commonsourceibias.n198 commonsourceibias.n197 49.296
R22585 commonsourceibias.n909 commonsourceibias.n908 49.296
R22586 commonsourceibias.n926 commonsourceibias.n859 49.296
R22587 commonsourceibias.n793 commonsourceibias.n792 49.296
R22588 commonsourceibias.n810 commonsourceibias.n743 49.296
R22589 commonsourceibias.n563 commonsourceibias.n562 49.296
R22590 commonsourceibias.n580 commonsourceibias.n513 49.296
R22591 commonsourceibias.n695 commonsourceibias.n492 49.296
R22592 commonsourceibias.n678 commonsourceibias.n677 49.296
R22593 commonsourceibias.n431 commonsourceibias.n383 48.3272
R22594 commonsourceibias.n443 commonsourceibias.n442 48.3272
R22595 commonsourceibias.n327 commonsourceibias.n326 48.3272
R22596 commonsourceibias.n315 commonsourceibias.n267 48.3272
R22597 commonsourceibias.n90 commonsourceibias.n89 48.3272
R22598 commonsourceibias.n78 commonsourceibias.n30 48.3272
R22599 commonsourceibias.n212 commonsourceibias.n211 48.3272
R22600 commonsourceibias.n202 commonsourceibias.n201 48.3272
R22601 commonsourceibias.n911 commonsourceibias.n863 48.3272
R22602 commonsourceibias.n924 commonsourceibias.n923 48.3272
R22603 commonsourceibias.n795 commonsourceibias.n747 48.3272
R22604 commonsourceibias.n808 commonsourceibias.n807 48.3272
R22605 commonsourceibias.n565 commonsourceibias.n517 48.3272
R22606 commonsourceibias.n578 commonsourceibias.n577 48.3272
R22607 commonsourceibias.n693 commonsourceibias.n692 48.3272
R22608 commonsourceibias.n682 commonsourceibias.n681 48.3272
R22609 commonsourceibias.n417 commonsourceibias.n388 47.3584
R22610 commonsourceibias.n457 commonsourceibias.n456 47.3584
R22611 commonsourceibias.n341 commonsourceibias.n340 47.3584
R22612 commonsourceibias.n301 commonsourceibias.n272 47.3584
R22613 commonsourceibias.n104 commonsourceibias.n103 47.3584
R22614 commonsourceibias.n64 commonsourceibias.n35 47.3584
R22615 commonsourceibias.n226 commonsourceibias.n225 47.3584
R22616 commonsourceibias.n186 commonsourceibias.n157 47.3584
R22617 commonsourceibias.n896 commonsourceibias.n867 47.3584
R22618 commonsourceibias.n939 commonsourceibias.n938 47.3584
R22619 commonsourceibias.n780 commonsourceibias.n751 47.3584
R22620 commonsourceibias.n823 commonsourceibias.n822 47.3584
R22621 commonsourceibias.n550 commonsourceibias.n521 47.3584
R22622 commonsourceibias.n593 commonsourceibias.n592 47.3584
R22623 commonsourceibias.n708 commonsourceibias.n707 47.3584
R22624 commonsourceibias.n666 commonsourceibias.n637 47.3584
R22625 commonsourceibias.n403 commonsourceibias.n393 46.3896
R22626 commonsourceibias.n471 commonsourceibias.n470 46.3896
R22627 commonsourceibias.n355 commonsourceibias.n354 46.3896
R22628 commonsourceibias.n287 commonsourceibias.n277 46.3896
R22629 commonsourceibias.n118 commonsourceibias.n117 46.3896
R22630 commonsourceibias.n50 commonsourceibias.n40 46.3896
R22631 commonsourceibias.n240 commonsourceibias.n239 46.3896
R22632 commonsourceibias.n172 commonsourceibias.n162 46.3896
R22633 commonsourceibias.n881 commonsourceibias.n871 46.3896
R22634 commonsourceibias.n954 commonsourceibias.n953 46.3896
R22635 commonsourceibias.n765 commonsourceibias.n755 46.3896
R22636 commonsourceibias.n838 commonsourceibias.n837 46.3896
R22637 commonsourceibias.n535 commonsourceibias.n525 46.3896
R22638 commonsourceibias.n608 commonsourceibias.n607 46.3896
R22639 commonsourceibias.n723 commonsourceibias.n722 46.3896
R22640 commonsourceibias.n651 commonsourceibias.n641 46.3896
R22641 commonsourceibias.n398 commonsourceibias.n397 44.7059
R22642 commonsourceibias.n876 commonsourceibias.n875 44.7059
R22643 commonsourceibias.n760 commonsourceibias.n759 44.7059
R22644 commonsourceibias.n530 commonsourceibias.n529 44.7059
R22645 commonsourceibias.n646 commonsourceibias.n645 44.7059
R22646 commonsourceibias.n282 commonsourceibias.n281 44.7059
R22647 commonsourceibias.n45 commonsourceibias.n44 44.7059
R22648 commonsourceibias.n167 commonsourceibias.n166 44.7059
R22649 commonsourceibias.n407 commonsourceibias.n393 34.7644
R22650 commonsourceibias.n470 commonsourceibias.n370 34.7644
R22651 commonsourceibias.n354 commonsourceibias.n254 34.7644
R22652 commonsourceibias.n291 commonsourceibias.n277 34.7644
R22653 commonsourceibias.n117 commonsourceibias.n17 34.7644
R22654 commonsourceibias.n54 commonsourceibias.n40 34.7644
R22655 commonsourceibias.n239 commonsourceibias.n3 34.7644
R22656 commonsourceibias.n176 commonsourceibias.n162 34.7644
R22657 commonsourceibias.n885 commonsourceibias.n871 34.7644
R22658 commonsourceibias.n953 commonsourceibias.n853 34.7644
R22659 commonsourceibias.n769 commonsourceibias.n755 34.7644
R22660 commonsourceibias.n837 commonsourceibias.n737 34.7644
R22661 commonsourceibias.n539 commonsourceibias.n525 34.7644
R22662 commonsourceibias.n607 commonsourceibias.n507 34.7644
R22663 commonsourceibias.n722 commonsourceibias.n486 34.7644
R22664 commonsourceibias.n655 commonsourceibias.n641 34.7644
R22665 commonsourceibias.n421 commonsourceibias.n388 33.7956
R22666 commonsourceibias.n456 commonsourceibias.n375 33.7956
R22667 commonsourceibias.n340 commonsourceibias.n259 33.7956
R22668 commonsourceibias.n305 commonsourceibias.n272 33.7956
R22669 commonsourceibias.n103 commonsourceibias.n22 33.7956
R22670 commonsourceibias.n68 commonsourceibias.n35 33.7956
R22671 commonsourceibias.n225 commonsourceibias.n8 33.7956
R22672 commonsourceibias.n190 commonsourceibias.n157 33.7956
R22673 commonsourceibias.n900 commonsourceibias.n867 33.7956
R22674 commonsourceibias.n938 commonsourceibias.n857 33.7956
R22675 commonsourceibias.n784 commonsourceibias.n751 33.7956
R22676 commonsourceibias.n822 commonsourceibias.n741 33.7956
R22677 commonsourceibias.n554 commonsourceibias.n521 33.7956
R22678 commonsourceibias.n592 commonsourceibias.n511 33.7956
R22679 commonsourceibias.n707 commonsourceibias.n490 33.7956
R22680 commonsourceibias.n670 commonsourceibias.n637 33.7956
R22681 commonsourceibias.n435 commonsourceibias.n383 32.8269
R22682 commonsourceibias.n442 commonsourceibias.n380 32.8269
R22683 commonsourceibias.n326 commonsourceibias.n264 32.8269
R22684 commonsourceibias.n319 commonsourceibias.n267 32.8269
R22685 commonsourceibias.n89 commonsourceibias.n27 32.8269
R22686 commonsourceibias.n82 commonsourceibias.n30 32.8269
R22687 commonsourceibias.n211 commonsourceibias.n13 32.8269
R22688 commonsourceibias.n203 commonsourceibias.n202 32.8269
R22689 commonsourceibias.n915 commonsourceibias.n863 32.8269
R22690 commonsourceibias.n923 commonsourceibias.n861 32.8269
R22691 commonsourceibias.n799 commonsourceibias.n747 32.8269
R22692 commonsourceibias.n807 commonsourceibias.n745 32.8269
R22693 commonsourceibias.n569 commonsourceibias.n517 32.8269
R22694 commonsourceibias.n577 commonsourceibias.n515 32.8269
R22695 commonsourceibias.n692 commonsourceibias.n494 32.8269
R22696 commonsourceibias.n683 commonsourceibias.n682 32.8269
R22697 commonsourceibias.n428 commonsourceibias.n385 31.8581
R22698 commonsourceibias.n449 commonsourceibias.n378 31.8581
R22699 commonsourceibias.n333 commonsourceibias.n262 31.8581
R22700 commonsourceibias.n312 commonsourceibias.n269 31.8581
R22701 commonsourceibias.n96 commonsourceibias.n25 31.8581
R22702 commonsourceibias.n75 commonsourceibias.n32 31.8581
R22703 commonsourceibias.n218 commonsourceibias.n11 31.8581
R22704 commonsourceibias.n197 commonsourceibias.n196 31.8581
R22705 commonsourceibias.n908 commonsourceibias.n865 31.8581
R22706 commonsourceibias.n930 commonsourceibias.n859 31.8581
R22707 commonsourceibias.n792 commonsourceibias.n749 31.8581
R22708 commonsourceibias.n814 commonsourceibias.n743 31.8581
R22709 commonsourceibias.n562 commonsourceibias.n519 31.8581
R22710 commonsourceibias.n584 commonsourceibias.n513 31.8581
R22711 commonsourceibias.n699 commonsourceibias.n492 31.8581
R22712 commonsourceibias.n677 commonsourceibias.n676 31.8581
R22713 commonsourceibias.n414 commonsourceibias.n390 30.8893
R22714 commonsourceibias.n463 commonsourceibias.n373 30.8893
R22715 commonsourceibias.n347 commonsourceibias.n257 30.8893
R22716 commonsourceibias.n298 commonsourceibias.n274 30.8893
R22717 commonsourceibias.n110 commonsourceibias.n20 30.8893
R22718 commonsourceibias.n61 commonsourceibias.n37 30.8893
R22719 commonsourceibias.n232 commonsourceibias.n6 30.8893
R22720 commonsourceibias.n183 commonsourceibias.n159 30.8893
R22721 commonsourceibias.n893 commonsourceibias.n869 30.8893
R22722 commonsourceibias.n945 commonsourceibias.n855 30.8893
R22723 commonsourceibias.n777 commonsourceibias.n753 30.8893
R22724 commonsourceibias.n829 commonsourceibias.n739 30.8893
R22725 commonsourceibias.n547 commonsourceibias.n523 30.8893
R22726 commonsourceibias.n599 commonsourceibias.n509 30.8893
R22727 commonsourceibias.n714 commonsourceibias.n488 30.8893
R22728 commonsourceibias.n663 commonsourceibias.n639 30.8893
R22729 commonsourceibias.n400 commonsourceibias.n395 29.9206
R22730 commonsourceibias.n477 commonsourceibias.n368 29.9206
R22731 commonsourceibias.n361 commonsourceibias.n252 29.9206
R22732 commonsourceibias.n284 commonsourceibias.n279 29.9206
R22733 commonsourceibias.n124 commonsourceibias.n15 29.9206
R22734 commonsourceibias.n47 commonsourceibias.n42 29.9206
R22735 commonsourceibias.n246 commonsourceibias.n1 29.9206
R22736 commonsourceibias.n169 commonsourceibias.n164 29.9206
R22737 commonsourceibias.n878 commonsourceibias.n873 29.9206
R22738 commonsourceibias.n960 commonsourceibias.n851 29.9206
R22739 commonsourceibias.n762 commonsourceibias.n757 29.9206
R22740 commonsourceibias.n844 commonsourceibias.n735 29.9206
R22741 commonsourceibias.n532 commonsourceibias.n527 29.9206
R22742 commonsourceibias.n614 commonsourceibias.n505 29.9206
R22743 commonsourceibias.n729 commonsourceibias.n484 29.9206
R22744 commonsourceibias.n648 commonsourceibias.n643 29.9206
R22745 commonsourceibias.n479 commonsourceibias.n478 21.8872
R22746 commonsourceibias.n363 commonsourceibias.n362 21.8872
R22747 commonsourceibias.n126 commonsourceibias.n125 21.8872
R22748 commonsourceibias.n248 commonsourceibias.n247 21.8872
R22749 commonsourceibias.n962 commonsourceibias.n961 21.8872
R22750 commonsourceibias.n846 commonsourceibias.n845 21.8872
R22751 commonsourceibias.n616 commonsourceibias.n615 21.8872
R22752 commonsourceibias.n731 commonsourceibias.n730 21.8872
R22753 commonsourceibias.n410 commonsourceibias.n392 21.3954
R22754 commonsourceibias.n465 commonsourceibias.n464 21.3954
R22755 commonsourceibias.n349 commonsourceibias.n348 21.3954
R22756 commonsourceibias.n294 commonsourceibias.n276 21.3954
R22757 commonsourceibias.n112 commonsourceibias.n111 21.3954
R22758 commonsourceibias.n57 commonsourceibias.n39 21.3954
R22759 commonsourceibias.n234 commonsourceibias.n233 21.3954
R22760 commonsourceibias.n179 commonsourceibias.n161 21.3954
R22761 commonsourceibias.n889 commonsourceibias.n888 21.3954
R22762 commonsourceibias.n947 commonsourceibias.n946 21.3954
R22763 commonsourceibias.n773 commonsourceibias.n772 21.3954
R22764 commonsourceibias.n831 commonsourceibias.n830 21.3954
R22765 commonsourceibias.n543 commonsourceibias.n542 21.3954
R22766 commonsourceibias.n601 commonsourceibias.n600 21.3954
R22767 commonsourceibias.n716 commonsourceibias.n715 21.3954
R22768 commonsourceibias.n659 commonsourceibias.n658 21.3954
R22769 commonsourceibias.n424 commonsourceibias.n387 20.9036
R22770 commonsourceibias.n451 commonsourceibias.n450 20.9036
R22771 commonsourceibias.n335 commonsourceibias.n334 20.9036
R22772 commonsourceibias.n308 commonsourceibias.n271 20.9036
R22773 commonsourceibias.n98 commonsourceibias.n97 20.9036
R22774 commonsourceibias.n71 commonsourceibias.n34 20.9036
R22775 commonsourceibias.n220 commonsourceibias.n219 20.9036
R22776 commonsourceibias.n193 commonsourceibias.n155 20.9036
R22777 commonsourceibias.n904 commonsourceibias.n903 20.9036
R22778 commonsourceibias.n932 commonsourceibias.n931 20.9036
R22779 commonsourceibias.n788 commonsourceibias.n787 20.9036
R22780 commonsourceibias.n816 commonsourceibias.n815 20.9036
R22781 commonsourceibias.n558 commonsourceibias.n557 20.9036
R22782 commonsourceibias.n586 commonsourceibias.n585 20.9036
R22783 commonsourceibias.n701 commonsourceibias.n700 20.9036
R22784 commonsourceibias.n673 commonsourceibias.n635 20.9036
R22785 commonsourceibias.n437 commonsourceibias.n436 20.4117
R22786 commonsourceibias.n438 commonsourceibias.n382 20.4117
R22787 commonsourceibias.n322 commonsourceibias.n266 20.4117
R22788 commonsourceibias.n321 commonsourceibias.n320 20.4117
R22789 commonsourceibias.n85 commonsourceibias.n29 20.4117
R22790 commonsourceibias.n84 commonsourceibias.n83 20.4117
R22791 commonsourceibias.n207 commonsourceibias.n150 20.4117
R22792 commonsourceibias.n206 commonsourceibias.n151 20.4117
R22793 commonsourceibias.n917 commonsourceibias.n916 20.4117
R22794 commonsourceibias.n919 commonsourceibias.n918 20.4117
R22795 commonsourceibias.n801 commonsourceibias.n800 20.4117
R22796 commonsourceibias.n803 commonsourceibias.n802 20.4117
R22797 commonsourceibias.n571 commonsourceibias.n570 20.4117
R22798 commonsourceibias.n573 commonsourceibias.n572 20.4117
R22799 commonsourceibias.n688 commonsourceibias.n687 20.4117
R22800 commonsourceibias.n686 commonsourceibias.n631 20.4117
R22801 commonsourceibias.n423 commonsourceibias.n422 19.9199
R22802 commonsourceibias.n452 commonsourceibias.n377 19.9199
R22803 commonsourceibias.n336 commonsourceibias.n261 19.9199
R22804 commonsourceibias.n307 commonsourceibias.n306 19.9199
R22805 commonsourceibias.n99 commonsourceibias.n24 19.9199
R22806 commonsourceibias.n70 commonsourceibias.n69 19.9199
R22807 commonsourceibias.n221 commonsourceibias.n10 19.9199
R22808 commonsourceibias.n192 commonsourceibias.n191 19.9199
R22809 commonsourceibias.n902 commonsourceibias.n901 19.9199
R22810 commonsourceibias.n934 commonsourceibias.n933 19.9199
R22811 commonsourceibias.n786 commonsourceibias.n785 19.9199
R22812 commonsourceibias.n818 commonsourceibias.n817 19.9199
R22813 commonsourceibias.n556 commonsourceibias.n555 19.9199
R22814 commonsourceibias.n588 commonsourceibias.n587 19.9199
R22815 commonsourceibias.n703 commonsourceibias.n702 19.9199
R22816 commonsourceibias.n672 commonsourceibias.n671 19.9199
R22817 commonsourceibias.n409 commonsourceibias.n408 19.4281
R22818 commonsourceibias.n466 commonsourceibias.n372 19.4281
R22819 commonsourceibias.n350 commonsourceibias.n256 19.4281
R22820 commonsourceibias.n293 commonsourceibias.n292 19.4281
R22821 commonsourceibias.n113 commonsourceibias.n19 19.4281
R22822 commonsourceibias.n56 commonsourceibias.n55 19.4281
R22823 commonsourceibias.n235 commonsourceibias.n5 19.4281
R22824 commonsourceibias.n178 commonsourceibias.n177 19.4281
R22825 commonsourceibias.n887 commonsourceibias.n886 19.4281
R22826 commonsourceibias.n949 commonsourceibias.n948 19.4281
R22827 commonsourceibias.n771 commonsourceibias.n770 19.4281
R22828 commonsourceibias.n833 commonsourceibias.n832 19.4281
R22829 commonsourceibias.n541 commonsourceibias.n540 19.4281
R22830 commonsourceibias.n603 commonsourceibias.n602 19.4281
R22831 commonsourceibias.n718 commonsourceibias.n717 19.4281
R22832 commonsourceibias.n657 commonsourceibias.n656 19.4281
R22833 commonsourceibias.n402 commonsourceibias.n401 13.526
R22834 commonsourceibias.n473 commonsourceibias.n472 13.526
R22835 commonsourceibias.n357 commonsourceibias.n356 13.526
R22836 commonsourceibias.n286 commonsourceibias.n285 13.526
R22837 commonsourceibias.n120 commonsourceibias.n119 13.526
R22838 commonsourceibias.n49 commonsourceibias.n48 13.526
R22839 commonsourceibias.n242 commonsourceibias.n241 13.526
R22840 commonsourceibias.n171 commonsourceibias.n170 13.526
R22841 commonsourceibias.n880 commonsourceibias.n879 13.526
R22842 commonsourceibias.n956 commonsourceibias.n955 13.526
R22843 commonsourceibias.n764 commonsourceibias.n763 13.526
R22844 commonsourceibias.n840 commonsourceibias.n839 13.526
R22845 commonsourceibias.n534 commonsourceibias.n533 13.526
R22846 commonsourceibias.n610 commonsourceibias.n609 13.526
R22847 commonsourceibias.n725 commonsourceibias.n724 13.526
R22848 commonsourceibias.n650 commonsourceibias.n649 13.526
R22849 commonsourceibias.n130 commonsourceibias.n128 13.2322
R22850 commonsourceibias.n620 commonsourceibias.n618 13.2322
R22851 commonsourceibias.n416 commonsourceibias.n415 13.0342
R22852 commonsourceibias.n459 commonsourceibias.n458 13.0342
R22853 commonsourceibias.n343 commonsourceibias.n342 13.0342
R22854 commonsourceibias.n300 commonsourceibias.n299 13.0342
R22855 commonsourceibias.n106 commonsourceibias.n105 13.0342
R22856 commonsourceibias.n63 commonsourceibias.n62 13.0342
R22857 commonsourceibias.n228 commonsourceibias.n227 13.0342
R22858 commonsourceibias.n185 commonsourceibias.n184 13.0342
R22859 commonsourceibias.n895 commonsourceibias.n894 13.0342
R22860 commonsourceibias.n941 commonsourceibias.n940 13.0342
R22861 commonsourceibias.n779 commonsourceibias.n778 13.0342
R22862 commonsourceibias.n825 commonsourceibias.n824 13.0342
R22863 commonsourceibias.n549 commonsourceibias.n548 13.0342
R22864 commonsourceibias.n595 commonsourceibias.n594 13.0342
R22865 commonsourceibias.n710 commonsourceibias.n709 13.0342
R22866 commonsourceibias.n665 commonsourceibias.n664 13.0342
R22867 commonsourceibias.n430 commonsourceibias.n429 12.5423
R22868 commonsourceibias.n445 commonsourceibias.n444 12.5423
R22869 commonsourceibias.n329 commonsourceibias.n328 12.5423
R22870 commonsourceibias.n314 commonsourceibias.n313 12.5423
R22871 commonsourceibias.n92 commonsourceibias.n91 12.5423
R22872 commonsourceibias.n77 commonsourceibias.n76 12.5423
R22873 commonsourceibias.n214 commonsourceibias.n213 12.5423
R22874 commonsourceibias.n198 commonsourceibias.n153 12.5423
R22875 commonsourceibias.n910 commonsourceibias.n909 12.5423
R22876 commonsourceibias.n926 commonsourceibias.n925 12.5423
R22877 commonsourceibias.n794 commonsourceibias.n793 12.5423
R22878 commonsourceibias.n810 commonsourceibias.n809 12.5423
R22879 commonsourceibias.n564 commonsourceibias.n563 12.5423
R22880 commonsourceibias.n580 commonsourceibias.n579 12.5423
R22881 commonsourceibias.n695 commonsourceibias.n694 12.5423
R22882 commonsourceibias.n678 commonsourceibias.n633 12.5423
R22883 commonsourceibias.n431 commonsourceibias.n430 12.0505
R22884 commonsourceibias.n444 commonsourceibias.n443 12.0505
R22885 commonsourceibias.n328 commonsourceibias.n327 12.0505
R22886 commonsourceibias.n315 commonsourceibias.n314 12.0505
R22887 commonsourceibias.n91 commonsourceibias.n90 12.0505
R22888 commonsourceibias.n78 commonsourceibias.n77 12.0505
R22889 commonsourceibias.n213 commonsourceibias.n212 12.0505
R22890 commonsourceibias.n201 commonsourceibias.n153 12.0505
R22891 commonsourceibias.n911 commonsourceibias.n910 12.0505
R22892 commonsourceibias.n925 commonsourceibias.n924 12.0505
R22893 commonsourceibias.n795 commonsourceibias.n794 12.0505
R22894 commonsourceibias.n809 commonsourceibias.n808 12.0505
R22895 commonsourceibias.n565 commonsourceibias.n564 12.0505
R22896 commonsourceibias.n579 commonsourceibias.n578 12.0505
R22897 commonsourceibias.n694 commonsourceibias.n693 12.0505
R22898 commonsourceibias.n681 commonsourceibias.n633 12.0505
R22899 commonsourceibias.n417 commonsourceibias.n416 11.5587
R22900 commonsourceibias.n458 commonsourceibias.n457 11.5587
R22901 commonsourceibias.n342 commonsourceibias.n341 11.5587
R22902 commonsourceibias.n301 commonsourceibias.n300 11.5587
R22903 commonsourceibias.n105 commonsourceibias.n104 11.5587
R22904 commonsourceibias.n64 commonsourceibias.n63 11.5587
R22905 commonsourceibias.n227 commonsourceibias.n226 11.5587
R22906 commonsourceibias.n186 commonsourceibias.n185 11.5587
R22907 commonsourceibias.n896 commonsourceibias.n895 11.5587
R22908 commonsourceibias.n940 commonsourceibias.n939 11.5587
R22909 commonsourceibias.n780 commonsourceibias.n779 11.5587
R22910 commonsourceibias.n824 commonsourceibias.n823 11.5587
R22911 commonsourceibias.n550 commonsourceibias.n549 11.5587
R22912 commonsourceibias.n594 commonsourceibias.n593 11.5587
R22913 commonsourceibias.n709 commonsourceibias.n708 11.5587
R22914 commonsourceibias.n666 commonsourceibias.n665 11.5587
R22915 commonsourceibias.n403 commonsourceibias.n402 11.0668
R22916 commonsourceibias.n472 commonsourceibias.n471 11.0668
R22917 commonsourceibias.n356 commonsourceibias.n355 11.0668
R22918 commonsourceibias.n287 commonsourceibias.n286 11.0668
R22919 commonsourceibias.n119 commonsourceibias.n118 11.0668
R22920 commonsourceibias.n50 commonsourceibias.n49 11.0668
R22921 commonsourceibias.n241 commonsourceibias.n240 11.0668
R22922 commonsourceibias.n172 commonsourceibias.n171 11.0668
R22923 commonsourceibias.n881 commonsourceibias.n880 11.0668
R22924 commonsourceibias.n955 commonsourceibias.n954 11.0668
R22925 commonsourceibias.n765 commonsourceibias.n764 11.0668
R22926 commonsourceibias.n839 commonsourceibias.n838 11.0668
R22927 commonsourceibias.n535 commonsourceibias.n534 11.0668
R22928 commonsourceibias.n609 commonsourceibias.n608 11.0668
R22929 commonsourceibias.n724 commonsourceibias.n723 11.0668
R22930 commonsourceibias.n651 commonsourceibias.n650 11.0668
R22931 commonsourceibias.n966 commonsourceibias.n482 10.122
R22932 commonsourceibias.n149 commonsourceibias.n148 9.50363
R22933 commonsourceibias.n630 commonsourceibias.n629 9.50363
R22934 commonsourceibias.n366 commonsourceibias.n250 8.76042
R22935 commonsourceibias.n849 commonsourceibias.n733 8.76042
R22936 commonsourceibias.n966 commonsourceibias.n965 8.46921
R22937 commonsourceibias.n408 commonsourceibias.n407 5.16479
R22938 commonsourceibias.n372 commonsourceibias.n370 5.16479
R22939 commonsourceibias.n256 commonsourceibias.n254 5.16479
R22940 commonsourceibias.n292 commonsourceibias.n291 5.16479
R22941 commonsourceibias.n19 commonsourceibias.n17 5.16479
R22942 commonsourceibias.n55 commonsourceibias.n54 5.16479
R22943 commonsourceibias.n5 commonsourceibias.n3 5.16479
R22944 commonsourceibias.n177 commonsourceibias.n176 5.16479
R22945 commonsourceibias.n886 commonsourceibias.n885 5.16479
R22946 commonsourceibias.n948 commonsourceibias.n853 5.16479
R22947 commonsourceibias.n770 commonsourceibias.n769 5.16479
R22948 commonsourceibias.n832 commonsourceibias.n737 5.16479
R22949 commonsourceibias.n540 commonsourceibias.n539 5.16479
R22950 commonsourceibias.n602 commonsourceibias.n507 5.16479
R22951 commonsourceibias.n717 commonsourceibias.n486 5.16479
R22952 commonsourceibias.n656 commonsourceibias.n655 5.16479
R22953 commonsourceibias.n482 commonsourceibias.n481 5.03125
R22954 commonsourceibias.n366 commonsourceibias.n365 5.03125
R22955 commonsourceibias.n965 commonsourceibias.n964 5.03125
R22956 commonsourceibias.n849 commonsourceibias.n848 5.03125
R22957 commonsourceibias.n422 commonsourceibias.n421 4.67295
R22958 commonsourceibias.n377 commonsourceibias.n375 4.67295
R22959 commonsourceibias.n261 commonsourceibias.n259 4.67295
R22960 commonsourceibias.n306 commonsourceibias.n305 4.67295
R22961 commonsourceibias.n24 commonsourceibias.n22 4.67295
R22962 commonsourceibias.n69 commonsourceibias.n68 4.67295
R22963 commonsourceibias.n10 commonsourceibias.n8 4.67295
R22964 commonsourceibias.n191 commonsourceibias.n190 4.67295
R22965 commonsourceibias.n901 commonsourceibias.n900 4.67295
R22966 commonsourceibias.n933 commonsourceibias.n857 4.67295
R22967 commonsourceibias.n785 commonsourceibias.n784 4.67295
R22968 commonsourceibias.n817 commonsourceibias.n741 4.67295
R22969 commonsourceibias.n555 commonsourceibias.n554 4.67295
R22970 commonsourceibias.n587 commonsourceibias.n511 4.67295
R22971 commonsourceibias.n702 commonsourceibias.n490 4.67295
R22972 commonsourceibias.n671 commonsourceibias.n670 4.67295
R22973 commonsourceibias commonsourceibias.n966 4.20978
R22974 commonsourceibias.n436 commonsourceibias.n435 4.18111
R22975 commonsourceibias.n382 commonsourceibias.n380 4.18111
R22976 commonsourceibias.n266 commonsourceibias.n264 4.18111
R22977 commonsourceibias.n320 commonsourceibias.n319 4.18111
R22978 commonsourceibias.n29 commonsourceibias.n27 4.18111
R22979 commonsourceibias.n83 commonsourceibias.n82 4.18111
R22980 commonsourceibias.n150 commonsourceibias.n13 4.18111
R22981 commonsourceibias.n203 commonsourceibias.n151 4.18111
R22982 commonsourceibias.n916 commonsourceibias.n915 4.18111
R22983 commonsourceibias.n918 commonsourceibias.n861 4.18111
R22984 commonsourceibias.n800 commonsourceibias.n799 4.18111
R22985 commonsourceibias.n802 commonsourceibias.n745 4.18111
R22986 commonsourceibias.n570 commonsourceibias.n569 4.18111
R22987 commonsourceibias.n572 commonsourceibias.n515 4.18111
R22988 commonsourceibias.n687 commonsourceibias.n494 4.18111
R22989 commonsourceibias.n683 commonsourceibias.n631 4.18111
R22990 commonsourceibias.n482 commonsourceibias.n366 3.72967
R22991 commonsourceibias.n965 commonsourceibias.n849 3.72967
R22992 commonsourceibias.n387 commonsourceibias.n385 3.68928
R22993 commonsourceibias.n450 commonsourceibias.n449 3.68928
R22994 commonsourceibias.n334 commonsourceibias.n333 3.68928
R22995 commonsourceibias.n271 commonsourceibias.n269 3.68928
R22996 commonsourceibias.n97 commonsourceibias.n96 3.68928
R22997 commonsourceibias.n34 commonsourceibias.n32 3.68928
R22998 commonsourceibias.n219 commonsourceibias.n218 3.68928
R22999 commonsourceibias.n196 commonsourceibias.n155 3.68928
R23000 commonsourceibias.n903 commonsourceibias.n865 3.68928
R23001 commonsourceibias.n931 commonsourceibias.n930 3.68928
R23002 commonsourceibias.n787 commonsourceibias.n749 3.68928
R23003 commonsourceibias.n815 commonsourceibias.n814 3.68928
R23004 commonsourceibias.n557 commonsourceibias.n519 3.68928
R23005 commonsourceibias.n585 commonsourceibias.n584 3.68928
R23006 commonsourceibias.n700 commonsourceibias.n699 3.68928
R23007 commonsourceibias.n676 commonsourceibias.n635 3.68928
R23008 commonsourceibias.n392 commonsourceibias.n390 3.19744
R23009 commonsourceibias.n464 commonsourceibias.n463 3.19744
R23010 commonsourceibias.n348 commonsourceibias.n347 3.19744
R23011 commonsourceibias.n276 commonsourceibias.n274 3.19744
R23012 commonsourceibias.n111 commonsourceibias.n110 3.19744
R23013 commonsourceibias.n39 commonsourceibias.n37 3.19744
R23014 commonsourceibias.n233 commonsourceibias.n232 3.19744
R23015 commonsourceibias.n161 commonsourceibias.n159 3.19744
R23016 commonsourceibias.n888 commonsourceibias.n869 3.19744
R23017 commonsourceibias.n946 commonsourceibias.n945 3.19744
R23018 commonsourceibias.n772 commonsourceibias.n753 3.19744
R23019 commonsourceibias.n830 commonsourceibias.n829 3.19744
R23020 commonsourceibias.n542 commonsourceibias.n523 3.19744
R23021 commonsourceibias.n600 commonsourceibias.n599 3.19744
R23022 commonsourceibias.n715 commonsourceibias.n714 3.19744
R23023 commonsourceibias.n658 commonsourceibias.n639 3.19744
R23024 commonsourceibias.n139 commonsourceibias.t59 2.82907
R23025 commonsourceibias.n139 commonsourceibias.t27 2.82907
R23026 commonsourceibias.n140 commonsourceibias.t43 2.82907
R23027 commonsourceibias.n140 commonsourceibias.t53 2.82907
R23028 commonsourceibias.n142 commonsourceibias.t63 2.82907
R23029 commonsourceibias.n142 commonsourceibias.t1 2.82907
R23030 commonsourceibias.n144 commonsourceibias.t71 2.82907
R23031 commonsourceibias.n144 commonsourceibias.t23 2.82907
R23032 commonsourceibias.n146 commonsourceibias.t31 2.82907
R23033 commonsourceibias.n146 commonsourceibias.t37 2.82907
R23034 commonsourceibias.n137 commonsourceibias.t19 2.82907
R23035 commonsourceibias.n137 commonsourceibias.t55 2.82907
R23036 commonsourceibias.n135 commonsourceibias.t35 2.82907
R23037 commonsourceibias.n135 commonsourceibias.t11 2.82907
R23038 commonsourceibias.n133 commonsourceibias.t75 2.82907
R23039 commonsourceibias.n133 commonsourceibias.t21 2.82907
R23040 commonsourceibias.n131 commonsourceibias.t5 2.82907
R23041 commonsourceibias.n131 commonsourceibias.t15 2.82907
R23042 commonsourceibias.n129 commonsourceibias.t17 2.82907
R23043 commonsourceibias.n129 commonsourceibias.t61 2.82907
R23044 commonsourceibias.n619 commonsourceibias.t77 2.82907
R23045 commonsourceibias.n619 commonsourceibias.t41 2.82907
R23046 commonsourceibias.n621 commonsourceibias.t39 2.82907
R23047 commonsourceibias.n621 commonsourceibias.t25 2.82907
R23048 commonsourceibias.n623 commonsourceibias.t47 2.82907
R23049 commonsourceibias.n623 commonsourceibias.t13 2.82907
R23050 commonsourceibias.n625 commonsourceibias.t33 2.82907
R23051 commonsourceibias.n625 commonsourceibias.t57 2.82907
R23052 commonsourceibias.n627 commonsourceibias.t73 2.82907
R23053 commonsourceibias.n627 commonsourceibias.t45 2.82907
R23054 commonsourceibias.n502 commonsourceibias.t65 2.82907
R23055 commonsourceibias.n502 commonsourceibias.t51 2.82907
R23056 commonsourceibias.n500 commonsourceibias.t49 2.82907
R23057 commonsourceibias.n500 commonsourceibias.t3 2.82907
R23058 commonsourceibias.n498 commonsourceibias.t29 2.82907
R23059 commonsourceibias.n498 commonsourceibias.t79 2.82907
R23060 commonsourceibias.n496 commonsourceibias.t7 2.82907
R23061 commonsourceibias.n496 commonsourceibias.t67 2.82907
R23062 commonsourceibias.n495 commonsourceibias.t69 2.82907
R23063 commonsourceibias.n495 commonsourceibias.t9 2.82907
R23064 commonsourceibias.n396 commonsourceibias.n395 2.7056
R23065 commonsourceibias.n478 commonsourceibias.n477 2.7056
R23066 commonsourceibias.n362 commonsourceibias.n361 2.7056
R23067 commonsourceibias.n280 commonsourceibias.n279 2.7056
R23068 commonsourceibias.n125 commonsourceibias.n124 2.7056
R23069 commonsourceibias.n43 commonsourceibias.n42 2.7056
R23070 commonsourceibias.n247 commonsourceibias.n246 2.7056
R23071 commonsourceibias.n165 commonsourceibias.n164 2.7056
R23072 commonsourceibias.n874 commonsourceibias.n873 2.7056
R23073 commonsourceibias.n961 commonsourceibias.n960 2.7056
R23074 commonsourceibias.n758 commonsourceibias.n757 2.7056
R23075 commonsourceibias.n845 commonsourceibias.n844 2.7056
R23076 commonsourceibias.n528 commonsourceibias.n527 2.7056
R23077 commonsourceibias.n615 commonsourceibias.n614 2.7056
R23078 commonsourceibias.n730 commonsourceibias.n729 2.7056
R23079 commonsourceibias.n644 commonsourceibias.n643 2.7056
R23080 commonsourceibias.n132 commonsourceibias.n130 0.573776
R23081 commonsourceibias.n134 commonsourceibias.n132 0.573776
R23082 commonsourceibias.n136 commonsourceibias.n134 0.573776
R23083 commonsourceibias.n138 commonsourceibias.n136 0.573776
R23084 commonsourceibias.n147 commonsourceibias.n145 0.573776
R23085 commonsourceibias.n145 commonsourceibias.n143 0.573776
R23086 commonsourceibias.n143 commonsourceibias.n141 0.573776
R23087 commonsourceibias.n499 commonsourceibias.n497 0.573776
R23088 commonsourceibias.n501 commonsourceibias.n499 0.573776
R23089 commonsourceibias.n503 commonsourceibias.n501 0.573776
R23090 commonsourceibias.n628 commonsourceibias.n626 0.573776
R23091 commonsourceibias.n626 commonsourceibias.n624 0.573776
R23092 commonsourceibias.n624 commonsourceibias.n622 0.573776
R23093 commonsourceibias.n622 commonsourceibias.n620 0.573776
R23094 commonsourceibias.n148 commonsourceibias.n138 0.287138
R23095 commonsourceibias.n148 commonsourceibias.n147 0.287138
R23096 commonsourceibias.n629 commonsourceibias.n503 0.287138
R23097 commonsourceibias.n629 commonsourceibias.n628 0.287138
R23098 commonsourceibias.n481 commonsourceibias.n367 0.285035
R23099 commonsourceibias.n365 commonsourceibias.n251 0.285035
R23100 commonsourceibias.n128 commonsourceibias.n14 0.285035
R23101 commonsourceibias.n250 commonsourceibias.n0 0.285035
R23102 commonsourceibias.n964 commonsourceibias.n850 0.285035
R23103 commonsourceibias.n848 commonsourceibias.n734 0.285035
R23104 commonsourceibias.n618 commonsourceibias.n504 0.285035
R23105 commonsourceibias.n733 commonsourceibias.n483 0.285035
R23106 commonsourceibias.n476 commonsourceibias.n367 0.189894
R23107 commonsourceibias.n476 commonsourceibias.n475 0.189894
R23108 commonsourceibias.n475 commonsourceibias.n474 0.189894
R23109 commonsourceibias.n474 commonsourceibias.n369 0.189894
R23110 commonsourceibias.n469 commonsourceibias.n369 0.189894
R23111 commonsourceibias.n469 commonsourceibias.n468 0.189894
R23112 commonsourceibias.n468 commonsourceibias.n467 0.189894
R23113 commonsourceibias.n467 commonsourceibias.n371 0.189894
R23114 commonsourceibias.n462 commonsourceibias.n371 0.189894
R23115 commonsourceibias.n462 commonsourceibias.n461 0.189894
R23116 commonsourceibias.n461 commonsourceibias.n460 0.189894
R23117 commonsourceibias.n460 commonsourceibias.n374 0.189894
R23118 commonsourceibias.n455 commonsourceibias.n374 0.189894
R23119 commonsourceibias.n455 commonsourceibias.n454 0.189894
R23120 commonsourceibias.n454 commonsourceibias.n453 0.189894
R23121 commonsourceibias.n453 commonsourceibias.n376 0.189894
R23122 commonsourceibias.n448 commonsourceibias.n376 0.189894
R23123 commonsourceibias.n448 commonsourceibias.n447 0.189894
R23124 commonsourceibias.n447 commonsourceibias.n446 0.189894
R23125 commonsourceibias.n446 commonsourceibias.n379 0.189894
R23126 commonsourceibias.n441 commonsourceibias.n379 0.189894
R23127 commonsourceibias.n441 commonsourceibias.n440 0.189894
R23128 commonsourceibias.n440 commonsourceibias.n439 0.189894
R23129 commonsourceibias.n439 commonsourceibias.n381 0.189894
R23130 commonsourceibias.n434 commonsourceibias.n381 0.189894
R23131 commonsourceibias.n434 commonsourceibias.n433 0.189894
R23132 commonsourceibias.n433 commonsourceibias.n432 0.189894
R23133 commonsourceibias.n432 commonsourceibias.n384 0.189894
R23134 commonsourceibias.n427 commonsourceibias.n384 0.189894
R23135 commonsourceibias.n427 commonsourceibias.n426 0.189894
R23136 commonsourceibias.n426 commonsourceibias.n425 0.189894
R23137 commonsourceibias.n425 commonsourceibias.n386 0.189894
R23138 commonsourceibias.n420 commonsourceibias.n386 0.189894
R23139 commonsourceibias.n420 commonsourceibias.n419 0.189894
R23140 commonsourceibias.n419 commonsourceibias.n418 0.189894
R23141 commonsourceibias.n418 commonsourceibias.n389 0.189894
R23142 commonsourceibias.n413 commonsourceibias.n389 0.189894
R23143 commonsourceibias.n413 commonsourceibias.n412 0.189894
R23144 commonsourceibias.n412 commonsourceibias.n411 0.189894
R23145 commonsourceibias.n411 commonsourceibias.n391 0.189894
R23146 commonsourceibias.n406 commonsourceibias.n391 0.189894
R23147 commonsourceibias.n406 commonsourceibias.n405 0.189894
R23148 commonsourceibias.n405 commonsourceibias.n404 0.189894
R23149 commonsourceibias.n404 commonsourceibias.n394 0.189894
R23150 commonsourceibias.n399 commonsourceibias.n394 0.189894
R23151 commonsourceibias.n399 commonsourceibias.n398 0.189894
R23152 commonsourceibias.n360 commonsourceibias.n251 0.189894
R23153 commonsourceibias.n360 commonsourceibias.n359 0.189894
R23154 commonsourceibias.n359 commonsourceibias.n358 0.189894
R23155 commonsourceibias.n358 commonsourceibias.n253 0.189894
R23156 commonsourceibias.n353 commonsourceibias.n253 0.189894
R23157 commonsourceibias.n353 commonsourceibias.n352 0.189894
R23158 commonsourceibias.n352 commonsourceibias.n351 0.189894
R23159 commonsourceibias.n351 commonsourceibias.n255 0.189894
R23160 commonsourceibias.n346 commonsourceibias.n255 0.189894
R23161 commonsourceibias.n346 commonsourceibias.n345 0.189894
R23162 commonsourceibias.n345 commonsourceibias.n344 0.189894
R23163 commonsourceibias.n344 commonsourceibias.n258 0.189894
R23164 commonsourceibias.n339 commonsourceibias.n258 0.189894
R23165 commonsourceibias.n339 commonsourceibias.n338 0.189894
R23166 commonsourceibias.n338 commonsourceibias.n337 0.189894
R23167 commonsourceibias.n337 commonsourceibias.n260 0.189894
R23168 commonsourceibias.n332 commonsourceibias.n260 0.189894
R23169 commonsourceibias.n332 commonsourceibias.n331 0.189894
R23170 commonsourceibias.n331 commonsourceibias.n330 0.189894
R23171 commonsourceibias.n330 commonsourceibias.n263 0.189894
R23172 commonsourceibias.n325 commonsourceibias.n263 0.189894
R23173 commonsourceibias.n325 commonsourceibias.n324 0.189894
R23174 commonsourceibias.n324 commonsourceibias.n323 0.189894
R23175 commonsourceibias.n323 commonsourceibias.n265 0.189894
R23176 commonsourceibias.n318 commonsourceibias.n265 0.189894
R23177 commonsourceibias.n318 commonsourceibias.n317 0.189894
R23178 commonsourceibias.n317 commonsourceibias.n316 0.189894
R23179 commonsourceibias.n316 commonsourceibias.n268 0.189894
R23180 commonsourceibias.n311 commonsourceibias.n268 0.189894
R23181 commonsourceibias.n311 commonsourceibias.n310 0.189894
R23182 commonsourceibias.n310 commonsourceibias.n309 0.189894
R23183 commonsourceibias.n309 commonsourceibias.n270 0.189894
R23184 commonsourceibias.n304 commonsourceibias.n270 0.189894
R23185 commonsourceibias.n304 commonsourceibias.n303 0.189894
R23186 commonsourceibias.n303 commonsourceibias.n302 0.189894
R23187 commonsourceibias.n302 commonsourceibias.n273 0.189894
R23188 commonsourceibias.n297 commonsourceibias.n273 0.189894
R23189 commonsourceibias.n297 commonsourceibias.n296 0.189894
R23190 commonsourceibias.n296 commonsourceibias.n295 0.189894
R23191 commonsourceibias.n295 commonsourceibias.n275 0.189894
R23192 commonsourceibias.n290 commonsourceibias.n275 0.189894
R23193 commonsourceibias.n290 commonsourceibias.n289 0.189894
R23194 commonsourceibias.n289 commonsourceibias.n288 0.189894
R23195 commonsourceibias.n288 commonsourceibias.n278 0.189894
R23196 commonsourceibias.n283 commonsourceibias.n278 0.189894
R23197 commonsourceibias.n283 commonsourceibias.n282 0.189894
R23198 commonsourceibias.n123 commonsourceibias.n14 0.189894
R23199 commonsourceibias.n123 commonsourceibias.n122 0.189894
R23200 commonsourceibias.n122 commonsourceibias.n121 0.189894
R23201 commonsourceibias.n121 commonsourceibias.n16 0.189894
R23202 commonsourceibias.n116 commonsourceibias.n16 0.189894
R23203 commonsourceibias.n116 commonsourceibias.n115 0.189894
R23204 commonsourceibias.n115 commonsourceibias.n114 0.189894
R23205 commonsourceibias.n114 commonsourceibias.n18 0.189894
R23206 commonsourceibias.n109 commonsourceibias.n18 0.189894
R23207 commonsourceibias.n109 commonsourceibias.n108 0.189894
R23208 commonsourceibias.n108 commonsourceibias.n107 0.189894
R23209 commonsourceibias.n107 commonsourceibias.n21 0.189894
R23210 commonsourceibias.n102 commonsourceibias.n21 0.189894
R23211 commonsourceibias.n102 commonsourceibias.n101 0.189894
R23212 commonsourceibias.n101 commonsourceibias.n100 0.189894
R23213 commonsourceibias.n100 commonsourceibias.n23 0.189894
R23214 commonsourceibias.n95 commonsourceibias.n23 0.189894
R23215 commonsourceibias.n95 commonsourceibias.n94 0.189894
R23216 commonsourceibias.n94 commonsourceibias.n93 0.189894
R23217 commonsourceibias.n93 commonsourceibias.n26 0.189894
R23218 commonsourceibias.n88 commonsourceibias.n26 0.189894
R23219 commonsourceibias.n88 commonsourceibias.n87 0.189894
R23220 commonsourceibias.n87 commonsourceibias.n86 0.189894
R23221 commonsourceibias.n86 commonsourceibias.n28 0.189894
R23222 commonsourceibias.n81 commonsourceibias.n28 0.189894
R23223 commonsourceibias.n81 commonsourceibias.n80 0.189894
R23224 commonsourceibias.n80 commonsourceibias.n79 0.189894
R23225 commonsourceibias.n79 commonsourceibias.n31 0.189894
R23226 commonsourceibias.n74 commonsourceibias.n31 0.189894
R23227 commonsourceibias.n74 commonsourceibias.n73 0.189894
R23228 commonsourceibias.n73 commonsourceibias.n72 0.189894
R23229 commonsourceibias.n72 commonsourceibias.n33 0.189894
R23230 commonsourceibias.n67 commonsourceibias.n33 0.189894
R23231 commonsourceibias.n67 commonsourceibias.n66 0.189894
R23232 commonsourceibias.n66 commonsourceibias.n65 0.189894
R23233 commonsourceibias.n65 commonsourceibias.n36 0.189894
R23234 commonsourceibias.n60 commonsourceibias.n36 0.189894
R23235 commonsourceibias.n60 commonsourceibias.n59 0.189894
R23236 commonsourceibias.n59 commonsourceibias.n58 0.189894
R23237 commonsourceibias.n58 commonsourceibias.n38 0.189894
R23238 commonsourceibias.n53 commonsourceibias.n38 0.189894
R23239 commonsourceibias.n53 commonsourceibias.n52 0.189894
R23240 commonsourceibias.n52 commonsourceibias.n51 0.189894
R23241 commonsourceibias.n51 commonsourceibias.n41 0.189894
R23242 commonsourceibias.n46 commonsourceibias.n41 0.189894
R23243 commonsourceibias.n46 commonsourceibias.n45 0.189894
R23244 commonsourceibias.n205 commonsourceibias.n204 0.189894
R23245 commonsourceibias.n204 commonsourceibias.n152 0.189894
R23246 commonsourceibias.n200 commonsourceibias.n152 0.189894
R23247 commonsourceibias.n200 commonsourceibias.n199 0.189894
R23248 commonsourceibias.n199 commonsourceibias.n154 0.189894
R23249 commonsourceibias.n195 commonsourceibias.n154 0.189894
R23250 commonsourceibias.n195 commonsourceibias.n194 0.189894
R23251 commonsourceibias.n194 commonsourceibias.n156 0.189894
R23252 commonsourceibias.n189 commonsourceibias.n156 0.189894
R23253 commonsourceibias.n189 commonsourceibias.n188 0.189894
R23254 commonsourceibias.n188 commonsourceibias.n187 0.189894
R23255 commonsourceibias.n187 commonsourceibias.n158 0.189894
R23256 commonsourceibias.n182 commonsourceibias.n158 0.189894
R23257 commonsourceibias.n182 commonsourceibias.n181 0.189894
R23258 commonsourceibias.n181 commonsourceibias.n180 0.189894
R23259 commonsourceibias.n180 commonsourceibias.n160 0.189894
R23260 commonsourceibias.n175 commonsourceibias.n160 0.189894
R23261 commonsourceibias.n175 commonsourceibias.n174 0.189894
R23262 commonsourceibias.n174 commonsourceibias.n173 0.189894
R23263 commonsourceibias.n173 commonsourceibias.n163 0.189894
R23264 commonsourceibias.n168 commonsourceibias.n163 0.189894
R23265 commonsourceibias.n168 commonsourceibias.n167 0.189894
R23266 commonsourceibias.n245 commonsourceibias.n0 0.189894
R23267 commonsourceibias.n245 commonsourceibias.n244 0.189894
R23268 commonsourceibias.n244 commonsourceibias.n243 0.189894
R23269 commonsourceibias.n243 commonsourceibias.n2 0.189894
R23270 commonsourceibias.n238 commonsourceibias.n2 0.189894
R23271 commonsourceibias.n238 commonsourceibias.n237 0.189894
R23272 commonsourceibias.n237 commonsourceibias.n236 0.189894
R23273 commonsourceibias.n236 commonsourceibias.n4 0.189894
R23274 commonsourceibias.n231 commonsourceibias.n4 0.189894
R23275 commonsourceibias.n231 commonsourceibias.n230 0.189894
R23276 commonsourceibias.n230 commonsourceibias.n229 0.189894
R23277 commonsourceibias.n229 commonsourceibias.n7 0.189894
R23278 commonsourceibias.n224 commonsourceibias.n7 0.189894
R23279 commonsourceibias.n224 commonsourceibias.n223 0.189894
R23280 commonsourceibias.n223 commonsourceibias.n222 0.189894
R23281 commonsourceibias.n222 commonsourceibias.n9 0.189894
R23282 commonsourceibias.n217 commonsourceibias.n9 0.189894
R23283 commonsourceibias.n217 commonsourceibias.n216 0.189894
R23284 commonsourceibias.n216 commonsourceibias.n215 0.189894
R23285 commonsourceibias.n215 commonsourceibias.n12 0.189894
R23286 commonsourceibias.n210 commonsourceibias.n12 0.189894
R23287 commonsourceibias.n210 commonsourceibias.n209 0.189894
R23288 commonsourceibias.n209 commonsourceibias.n208 0.189894
R23289 commonsourceibias.n877 commonsourceibias.n876 0.189894
R23290 commonsourceibias.n877 commonsourceibias.n872 0.189894
R23291 commonsourceibias.n882 commonsourceibias.n872 0.189894
R23292 commonsourceibias.n883 commonsourceibias.n882 0.189894
R23293 commonsourceibias.n884 commonsourceibias.n883 0.189894
R23294 commonsourceibias.n884 commonsourceibias.n870 0.189894
R23295 commonsourceibias.n890 commonsourceibias.n870 0.189894
R23296 commonsourceibias.n891 commonsourceibias.n890 0.189894
R23297 commonsourceibias.n892 commonsourceibias.n891 0.189894
R23298 commonsourceibias.n892 commonsourceibias.n868 0.189894
R23299 commonsourceibias.n897 commonsourceibias.n868 0.189894
R23300 commonsourceibias.n898 commonsourceibias.n897 0.189894
R23301 commonsourceibias.n899 commonsourceibias.n898 0.189894
R23302 commonsourceibias.n899 commonsourceibias.n866 0.189894
R23303 commonsourceibias.n905 commonsourceibias.n866 0.189894
R23304 commonsourceibias.n906 commonsourceibias.n905 0.189894
R23305 commonsourceibias.n907 commonsourceibias.n906 0.189894
R23306 commonsourceibias.n907 commonsourceibias.n864 0.189894
R23307 commonsourceibias.n912 commonsourceibias.n864 0.189894
R23308 commonsourceibias.n913 commonsourceibias.n912 0.189894
R23309 commonsourceibias.n914 commonsourceibias.n913 0.189894
R23310 commonsourceibias.n914 commonsourceibias.n862 0.189894
R23311 commonsourceibias.n920 commonsourceibias.n862 0.189894
R23312 commonsourceibias.n921 commonsourceibias.n920 0.189894
R23313 commonsourceibias.n922 commonsourceibias.n921 0.189894
R23314 commonsourceibias.n922 commonsourceibias.n860 0.189894
R23315 commonsourceibias.n927 commonsourceibias.n860 0.189894
R23316 commonsourceibias.n928 commonsourceibias.n927 0.189894
R23317 commonsourceibias.n929 commonsourceibias.n928 0.189894
R23318 commonsourceibias.n929 commonsourceibias.n858 0.189894
R23319 commonsourceibias.n935 commonsourceibias.n858 0.189894
R23320 commonsourceibias.n936 commonsourceibias.n935 0.189894
R23321 commonsourceibias.n937 commonsourceibias.n936 0.189894
R23322 commonsourceibias.n937 commonsourceibias.n856 0.189894
R23323 commonsourceibias.n942 commonsourceibias.n856 0.189894
R23324 commonsourceibias.n943 commonsourceibias.n942 0.189894
R23325 commonsourceibias.n944 commonsourceibias.n943 0.189894
R23326 commonsourceibias.n944 commonsourceibias.n854 0.189894
R23327 commonsourceibias.n950 commonsourceibias.n854 0.189894
R23328 commonsourceibias.n951 commonsourceibias.n950 0.189894
R23329 commonsourceibias.n952 commonsourceibias.n951 0.189894
R23330 commonsourceibias.n952 commonsourceibias.n852 0.189894
R23331 commonsourceibias.n957 commonsourceibias.n852 0.189894
R23332 commonsourceibias.n958 commonsourceibias.n957 0.189894
R23333 commonsourceibias.n959 commonsourceibias.n958 0.189894
R23334 commonsourceibias.n959 commonsourceibias.n850 0.189894
R23335 commonsourceibias.n761 commonsourceibias.n760 0.189894
R23336 commonsourceibias.n761 commonsourceibias.n756 0.189894
R23337 commonsourceibias.n766 commonsourceibias.n756 0.189894
R23338 commonsourceibias.n767 commonsourceibias.n766 0.189894
R23339 commonsourceibias.n768 commonsourceibias.n767 0.189894
R23340 commonsourceibias.n768 commonsourceibias.n754 0.189894
R23341 commonsourceibias.n774 commonsourceibias.n754 0.189894
R23342 commonsourceibias.n775 commonsourceibias.n774 0.189894
R23343 commonsourceibias.n776 commonsourceibias.n775 0.189894
R23344 commonsourceibias.n776 commonsourceibias.n752 0.189894
R23345 commonsourceibias.n781 commonsourceibias.n752 0.189894
R23346 commonsourceibias.n782 commonsourceibias.n781 0.189894
R23347 commonsourceibias.n783 commonsourceibias.n782 0.189894
R23348 commonsourceibias.n783 commonsourceibias.n750 0.189894
R23349 commonsourceibias.n789 commonsourceibias.n750 0.189894
R23350 commonsourceibias.n790 commonsourceibias.n789 0.189894
R23351 commonsourceibias.n791 commonsourceibias.n790 0.189894
R23352 commonsourceibias.n791 commonsourceibias.n748 0.189894
R23353 commonsourceibias.n796 commonsourceibias.n748 0.189894
R23354 commonsourceibias.n797 commonsourceibias.n796 0.189894
R23355 commonsourceibias.n798 commonsourceibias.n797 0.189894
R23356 commonsourceibias.n798 commonsourceibias.n746 0.189894
R23357 commonsourceibias.n804 commonsourceibias.n746 0.189894
R23358 commonsourceibias.n805 commonsourceibias.n804 0.189894
R23359 commonsourceibias.n806 commonsourceibias.n805 0.189894
R23360 commonsourceibias.n806 commonsourceibias.n744 0.189894
R23361 commonsourceibias.n811 commonsourceibias.n744 0.189894
R23362 commonsourceibias.n812 commonsourceibias.n811 0.189894
R23363 commonsourceibias.n813 commonsourceibias.n812 0.189894
R23364 commonsourceibias.n813 commonsourceibias.n742 0.189894
R23365 commonsourceibias.n819 commonsourceibias.n742 0.189894
R23366 commonsourceibias.n820 commonsourceibias.n819 0.189894
R23367 commonsourceibias.n821 commonsourceibias.n820 0.189894
R23368 commonsourceibias.n821 commonsourceibias.n740 0.189894
R23369 commonsourceibias.n826 commonsourceibias.n740 0.189894
R23370 commonsourceibias.n827 commonsourceibias.n826 0.189894
R23371 commonsourceibias.n828 commonsourceibias.n827 0.189894
R23372 commonsourceibias.n828 commonsourceibias.n738 0.189894
R23373 commonsourceibias.n834 commonsourceibias.n738 0.189894
R23374 commonsourceibias.n835 commonsourceibias.n834 0.189894
R23375 commonsourceibias.n836 commonsourceibias.n835 0.189894
R23376 commonsourceibias.n836 commonsourceibias.n736 0.189894
R23377 commonsourceibias.n841 commonsourceibias.n736 0.189894
R23378 commonsourceibias.n842 commonsourceibias.n841 0.189894
R23379 commonsourceibias.n843 commonsourceibias.n842 0.189894
R23380 commonsourceibias.n843 commonsourceibias.n734 0.189894
R23381 commonsourceibias.n531 commonsourceibias.n530 0.189894
R23382 commonsourceibias.n531 commonsourceibias.n526 0.189894
R23383 commonsourceibias.n536 commonsourceibias.n526 0.189894
R23384 commonsourceibias.n537 commonsourceibias.n536 0.189894
R23385 commonsourceibias.n538 commonsourceibias.n537 0.189894
R23386 commonsourceibias.n538 commonsourceibias.n524 0.189894
R23387 commonsourceibias.n544 commonsourceibias.n524 0.189894
R23388 commonsourceibias.n545 commonsourceibias.n544 0.189894
R23389 commonsourceibias.n546 commonsourceibias.n545 0.189894
R23390 commonsourceibias.n546 commonsourceibias.n522 0.189894
R23391 commonsourceibias.n551 commonsourceibias.n522 0.189894
R23392 commonsourceibias.n552 commonsourceibias.n551 0.189894
R23393 commonsourceibias.n553 commonsourceibias.n552 0.189894
R23394 commonsourceibias.n553 commonsourceibias.n520 0.189894
R23395 commonsourceibias.n559 commonsourceibias.n520 0.189894
R23396 commonsourceibias.n560 commonsourceibias.n559 0.189894
R23397 commonsourceibias.n561 commonsourceibias.n560 0.189894
R23398 commonsourceibias.n561 commonsourceibias.n518 0.189894
R23399 commonsourceibias.n566 commonsourceibias.n518 0.189894
R23400 commonsourceibias.n567 commonsourceibias.n566 0.189894
R23401 commonsourceibias.n568 commonsourceibias.n567 0.189894
R23402 commonsourceibias.n568 commonsourceibias.n516 0.189894
R23403 commonsourceibias.n574 commonsourceibias.n516 0.189894
R23404 commonsourceibias.n575 commonsourceibias.n574 0.189894
R23405 commonsourceibias.n576 commonsourceibias.n575 0.189894
R23406 commonsourceibias.n576 commonsourceibias.n514 0.189894
R23407 commonsourceibias.n581 commonsourceibias.n514 0.189894
R23408 commonsourceibias.n582 commonsourceibias.n581 0.189894
R23409 commonsourceibias.n583 commonsourceibias.n582 0.189894
R23410 commonsourceibias.n583 commonsourceibias.n512 0.189894
R23411 commonsourceibias.n589 commonsourceibias.n512 0.189894
R23412 commonsourceibias.n590 commonsourceibias.n589 0.189894
R23413 commonsourceibias.n591 commonsourceibias.n590 0.189894
R23414 commonsourceibias.n591 commonsourceibias.n510 0.189894
R23415 commonsourceibias.n596 commonsourceibias.n510 0.189894
R23416 commonsourceibias.n597 commonsourceibias.n596 0.189894
R23417 commonsourceibias.n598 commonsourceibias.n597 0.189894
R23418 commonsourceibias.n598 commonsourceibias.n508 0.189894
R23419 commonsourceibias.n604 commonsourceibias.n508 0.189894
R23420 commonsourceibias.n605 commonsourceibias.n604 0.189894
R23421 commonsourceibias.n606 commonsourceibias.n605 0.189894
R23422 commonsourceibias.n606 commonsourceibias.n506 0.189894
R23423 commonsourceibias.n611 commonsourceibias.n506 0.189894
R23424 commonsourceibias.n612 commonsourceibias.n611 0.189894
R23425 commonsourceibias.n613 commonsourceibias.n612 0.189894
R23426 commonsourceibias.n613 commonsourceibias.n504 0.189894
R23427 commonsourceibias.n647 commonsourceibias.n646 0.189894
R23428 commonsourceibias.n647 commonsourceibias.n642 0.189894
R23429 commonsourceibias.n652 commonsourceibias.n642 0.189894
R23430 commonsourceibias.n653 commonsourceibias.n652 0.189894
R23431 commonsourceibias.n654 commonsourceibias.n653 0.189894
R23432 commonsourceibias.n654 commonsourceibias.n640 0.189894
R23433 commonsourceibias.n660 commonsourceibias.n640 0.189894
R23434 commonsourceibias.n661 commonsourceibias.n660 0.189894
R23435 commonsourceibias.n662 commonsourceibias.n661 0.189894
R23436 commonsourceibias.n662 commonsourceibias.n638 0.189894
R23437 commonsourceibias.n667 commonsourceibias.n638 0.189894
R23438 commonsourceibias.n668 commonsourceibias.n667 0.189894
R23439 commonsourceibias.n669 commonsourceibias.n668 0.189894
R23440 commonsourceibias.n669 commonsourceibias.n636 0.189894
R23441 commonsourceibias.n674 commonsourceibias.n636 0.189894
R23442 commonsourceibias.n675 commonsourceibias.n674 0.189894
R23443 commonsourceibias.n675 commonsourceibias.n634 0.189894
R23444 commonsourceibias.n679 commonsourceibias.n634 0.189894
R23445 commonsourceibias.n680 commonsourceibias.n679 0.189894
R23446 commonsourceibias.n680 commonsourceibias.n632 0.189894
R23447 commonsourceibias.n684 commonsourceibias.n632 0.189894
R23448 commonsourceibias.n685 commonsourceibias.n684 0.189894
R23449 commonsourceibias.n690 commonsourceibias.n689 0.189894
R23450 commonsourceibias.n691 commonsourceibias.n690 0.189894
R23451 commonsourceibias.n691 commonsourceibias.n493 0.189894
R23452 commonsourceibias.n696 commonsourceibias.n493 0.189894
R23453 commonsourceibias.n697 commonsourceibias.n696 0.189894
R23454 commonsourceibias.n698 commonsourceibias.n697 0.189894
R23455 commonsourceibias.n698 commonsourceibias.n491 0.189894
R23456 commonsourceibias.n704 commonsourceibias.n491 0.189894
R23457 commonsourceibias.n705 commonsourceibias.n704 0.189894
R23458 commonsourceibias.n706 commonsourceibias.n705 0.189894
R23459 commonsourceibias.n706 commonsourceibias.n489 0.189894
R23460 commonsourceibias.n711 commonsourceibias.n489 0.189894
R23461 commonsourceibias.n712 commonsourceibias.n711 0.189894
R23462 commonsourceibias.n713 commonsourceibias.n712 0.189894
R23463 commonsourceibias.n713 commonsourceibias.n487 0.189894
R23464 commonsourceibias.n719 commonsourceibias.n487 0.189894
R23465 commonsourceibias.n720 commonsourceibias.n719 0.189894
R23466 commonsourceibias.n721 commonsourceibias.n720 0.189894
R23467 commonsourceibias.n721 commonsourceibias.n485 0.189894
R23468 commonsourceibias.n726 commonsourceibias.n485 0.189894
R23469 commonsourceibias.n727 commonsourceibias.n726 0.189894
R23470 commonsourceibias.n728 commonsourceibias.n727 0.189894
R23471 commonsourceibias.n728 commonsourceibias.n483 0.189894
R23472 commonsourceibias.n205 commonsourceibias.n149 0.0762576
R23473 commonsourceibias.n208 commonsourceibias.n149 0.0762576
R23474 commonsourceibias.n685 commonsourceibias.n630 0.0762576
R23475 commonsourceibias.n689 commonsourceibias.n630 0.0762576
R23476 minus.n53 minus.t28 323.478
R23477 minus.n11 minus.t8 323.478
R23478 minus.n82 minus.t13 297.12
R23479 minus.n80 minus.t15 297.12
R23480 minus.n44 minus.t5 297.12
R23481 minus.n74 minus.t6 297.12
R23482 minus.n46 minus.t26 297.12
R23483 minus.n68 minus.t21 297.12
R23484 minus.n48 minus.t23 297.12
R23485 minus.n62 minus.t16 297.12
R23486 minus.n50 minus.t17 297.12
R23487 minus.n56 minus.t9 297.12
R23488 minus.n52 minus.t27 297.12
R23489 minus.n10 minus.t7 297.12
R23490 minus.n14 minus.t11 297.12
R23491 minus.n16 minus.t10 297.12
R23492 minus.n20 minus.t12 297.12
R23493 minus.n22 minus.t20 297.12
R23494 minus.n26 minus.t18 297.12
R23495 minus.n28 minus.t25 297.12
R23496 minus.n32 minus.t24 297.12
R23497 minus.n34 minus.t14 297.12
R23498 minus.n38 minus.t22 297.12
R23499 minus.n40 minus.t19 297.12
R23500 minus.n88 minus.t2 243.255
R23501 minus.n87 minus.n85 224.169
R23502 minus.n87 minus.n86 223.454
R23503 minus.n55 minus.n54 161.3
R23504 minus.n56 minus.n51 161.3
R23505 minus.n58 minus.n57 161.3
R23506 minus.n59 minus.n50 161.3
R23507 minus.n61 minus.n60 161.3
R23508 minus.n62 minus.n49 161.3
R23509 minus.n64 minus.n63 161.3
R23510 minus.n65 minus.n48 161.3
R23511 minus.n67 minus.n66 161.3
R23512 minus.n68 minus.n47 161.3
R23513 minus.n70 minus.n69 161.3
R23514 minus.n71 minus.n46 161.3
R23515 minus.n73 minus.n72 161.3
R23516 minus.n74 minus.n45 161.3
R23517 minus.n76 minus.n75 161.3
R23518 minus.n77 minus.n44 161.3
R23519 minus.n79 minus.n78 161.3
R23520 minus.n80 minus.n43 161.3
R23521 minus.n81 minus.n42 161.3
R23522 minus.n83 minus.n82 161.3
R23523 minus.n41 minus.n40 161.3
R23524 minus.n39 minus.n0 161.3
R23525 minus.n38 minus.n37 161.3
R23526 minus.n36 minus.n1 161.3
R23527 minus.n35 minus.n34 161.3
R23528 minus.n33 minus.n2 161.3
R23529 minus.n32 minus.n31 161.3
R23530 minus.n30 minus.n3 161.3
R23531 minus.n29 minus.n28 161.3
R23532 minus.n27 minus.n4 161.3
R23533 minus.n26 minus.n25 161.3
R23534 minus.n24 minus.n5 161.3
R23535 minus.n23 minus.n22 161.3
R23536 minus.n21 minus.n6 161.3
R23537 minus.n20 minus.n19 161.3
R23538 minus.n18 minus.n7 161.3
R23539 minus.n17 minus.n16 161.3
R23540 minus.n15 minus.n8 161.3
R23541 minus.n14 minus.n13 161.3
R23542 minus.n12 minus.n9 161.3
R23543 minus.n82 minus.n81 46.0096
R23544 minus.n40 minus.n39 46.0096
R23545 minus.n12 minus.n11 45.0871
R23546 minus.n54 minus.n53 45.0871
R23547 minus.n80 minus.n79 41.6278
R23548 minus.n55 minus.n52 41.6278
R23549 minus.n10 minus.n9 41.6278
R23550 minus.n38 minus.n1 41.6278
R23551 minus.n75 minus.n44 37.246
R23552 minus.n57 minus.n56 37.246
R23553 minus.n15 minus.n14 37.246
R23554 minus.n34 minus.n33 37.246
R23555 minus.n84 minus.n83 33.3925
R23556 minus.n74 minus.n73 32.8641
R23557 minus.n61 minus.n50 32.8641
R23558 minus.n16 minus.n7 32.8641
R23559 minus.n32 minus.n3 32.8641
R23560 minus.n69 minus.n46 28.4823
R23561 minus.n63 minus.n62 28.4823
R23562 minus.n21 minus.n20 28.4823
R23563 minus.n28 minus.n27 28.4823
R23564 minus.n68 minus.n67 24.1005
R23565 minus.n67 minus.n48 24.1005
R23566 minus.n22 minus.n5 24.1005
R23567 minus.n26 minus.n5 24.1005
R23568 minus.n86 minus.t4 19.8005
R23569 minus.n86 minus.t3 19.8005
R23570 minus.n85 minus.t1 19.8005
R23571 minus.n85 minus.t0 19.8005
R23572 minus.n69 minus.n68 19.7187
R23573 minus.n63 minus.n48 19.7187
R23574 minus.n22 minus.n21 19.7187
R23575 minus.n27 minus.n26 19.7187
R23576 minus.n73 minus.n46 15.3369
R23577 minus.n62 minus.n61 15.3369
R23578 minus.n20 minus.n7 15.3369
R23579 minus.n28 minus.n3 15.3369
R23580 minus.n53 minus.n52 14.1472
R23581 minus.n11 minus.n10 14.1472
R23582 minus.n84 minus.n41 12.0933
R23583 minus minus.n89 11.7437
R23584 minus.n75 minus.n74 10.955
R23585 minus.n57 minus.n50 10.955
R23586 minus.n16 minus.n15 10.955
R23587 minus.n33 minus.n32 10.955
R23588 minus.n79 minus.n44 6.57323
R23589 minus.n56 minus.n55 6.57323
R23590 minus.n14 minus.n9 6.57323
R23591 minus.n34 minus.n1 6.57323
R23592 minus.n89 minus.n88 4.80222
R23593 minus.n81 minus.n80 2.19141
R23594 minus.n39 minus.n38 2.19141
R23595 minus.n89 minus.n84 0.972091
R23596 minus.n88 minus.n87 0.716017
R23597 minus.n83 minus.n42 0.189894
R23598 minus.n43 minus.n42 0.189894
R23599 minus.n78 minus.n43 0.189894
R23600 minus.n78 minus.n77 0.189894
R23601 minus.n77 minus.n76 0.189894
R23602 minus.n76 minus.n45 0.189894
R23603 minus.n72 minus.n45 0.189894
R23604 minus.n72 minus.n71 0.189894
R23605 minus.n71 minus.n70 0.189894
R23606 minus.n70 minus.n47 0.189894
R23607 minus.n66 minus.n47 0.189894
R23608 minus.n66 minus.n65 0.189894
R23609 minus.n65 minus.n64 0.189894
R23610 minus.n64 minus.n49 0.189894
R23611 minus.n60 minus.n49 0.189894
R23612 minus.n60 minus.n59 0.189894
R23613 minus.n59 minus.n58 0.189894
R23614 minus.n58 minus.n51 0.189894
R23615 minus.n54 minus.n51 0.189894
R23616 minus.n13 minus.n12 0.189894
R23617 minus.n13 minus.n8 0.189894
R23618 minus.n17 minus.n8 0.189894
R23619 minus.n18 minus.n17 0.189894
R23620 minus.n19 minus.n18 0.189894
R23621 minus.n19 minus.n6 0.189894
R23622 minus.n23 minus.n6 0.189894
R23623 minus.n24 minus.n23 0.189894
R23624 minus.n25 minus.n24 0.189894
R23625 minus.n25 minus.n4 0.189894
R23626 minus.n29 minus.n4 0.189894
R23627 minus.n30 minus.n29 0.189894
R23628 minus.n31 minus.n30 0.189894
R23629 minus.n31 minus.n2 0.189894
R23630 minus.n35 minus.n2 0.189894
R23631 minus.n36 minus.n35 0.189894
R23632 minus.n37 minus.n36 0.189894
R23633 minus.n37 minus.n0 0.189894
R23634 minus.n41 minus.n0 0.189894
R23635 a_n2318_8322.n8 a_n2318_8322.t3 74.6477
R23636 a_n2318_8322.n1 a_n2318_8322.t22 74.6477
R23637 a_n2318_8322.n20 a_n2318_8322.t21 74.6474
R23638 a_n2318_8322.n16 a_n2318_8322.t11 74.2899
R23639 a_n2318_8322.n9 a_n2318_8322.t1 74.2899
R23640 a_n2318_8322.n10 a_n2318_8322.t4 74.2899
R23641 a_n2318_8322.n13 a_n2318_8322.t5 74.2899
R23642 a_n2318_8322.n6 a_n2318_8322.t8 74.2899
R23643 a_n2318_8322.n20 a_n2318_8322.n19 70.6783
R23644 a_n2318_8322.n18 a_n2318_8322.n17 70.6783
R23645 a_n2318_8322.n8 a_n2318_8322.n7 70.6783
R23646 a_n2318_8322.n12 a_n2318_8322.n11 70.6783
R23647 a_n2318_8322.n1 a_n2318_8322.n0 70.6783
R23648 a_n2318_8322.n3 a_n2318_8322.n2 70.6783
R23649 a_n2318_8322.n5 a_n2318_8322.n4 70.6783
R23650 a_n2318_8322.n22 a_n2318_8322.n21 70.6782
R23651 a_n2318_8322.n14 a_n2318_8322.n6 23.4712
R23652 a_n2318_8322.n15 a_n2318_8322.t27 10.0266
R23653 a_n2318_8322.n14 a_n2318_8322.n13 6.95632
R23654 a_n2318_8322.n16 a_n2318_8322.n15 6.19447
R23655 a_n2318_8322.n15 a_n2318_8322.n14 5.3452
R23656 a_n2318_8322.n19 a_n2318_8322.t18 3.61217
R23657 a_n2318_8322.n19 a_n2318_8322.t15 3.61217
R23658 a_n2318_8322.n17 a_n2318_8322.t20 3.61217
R23659 a_n2318_8322.n17 a_n2318_8322.t13 3.61217
R23660 a_n2318_8322.n7 a_n2318_8322.t7 3.61217
R23661 a_n2318_8322.n7 a_n2318_8322.t6 3.61217
R23662 a_n2318_8322.n11 a_n2318_8322.t2 3.61217
R23663 a_n2318_8322.n11 a_n2318_8322.t0 3.61217
R23664 a_n2318_8322.n0 a_n2318_8322.t10 3.61217
R23665 a_n2318_8322.n0 a_n2318_8322.t9 3.61217
R23666 a_n2318_8322.n2 a_n2318_8322.t19 3.61217
R23667 a_n2318_8322.n2 a_n2318_8322.t14 3.61217
R23668 a_n2318_8322.n4 a_n2318_8322.t17 3.61217
R23669 a_n2318_8322.n4 a_n2318_8322.t16 3.61217
R23670 a_n2318_8322.n22 a_n2318_8322.t12 3.61217
R23671 a_n2318_8322.t23 a_n2318_8322.n22 3.61217
R23672 a_n2318_8322.n13 a_n2318_8322.n12 0.358259
R23673 a_n2318_8322.n12 a_n2318_8322.n10 0.358259
R23674 a_n2318_8322.n9 a_n2318_8322.n8 0.358259
R23675 a_n2318_8322.n6 a_n2318_8322.n5 0.358259
R23676 a_n2318_8322.n5 a_n2318_8322.n3 0.358259
R23677 a_n2318_8322.n3 a_n2318_8322.n1 0.358259
R23678 a_n2318_8322.n18 a_n2318_8322.n16 0.358259
R23679 a_n2318_8322.n21 a_n2318_8322.n18 0.358259
R23680 a_n2318_8322.n21 a_n2318_8322.n20 0.358259
R23681 a_n2318_8322.n10 a_n2318_8322.n9 0.101793
R23682 a_n2318_8322.t26 a_n2318_8322.t25 0.0788333
R23683 a_n2318_8322.t24 a_n2318_8322.t26 0.0631667
R23684 a_n2318_8322.t27 a_n2318_8322.t24 0.0471944
R23685 a_n2318_8322.t27 a_n2318_8322.t25 0.0453889
R23686 output.n41 output.n15 289.615
R23687 output.n72 output.n46 289.615
R23688 output.n104 output.n78 289.615
R23689 output.n136 output.n110 289.615
R23690 output.n77 output.n45 197.26
R23691 output.n77 output.n76 196.298
R23692 output.n109 output.n108 196.298
R23693 output.n141 output.n140 196.298
R23694 output.n42 output.n41 185
R23695 output.n40 output.n39 185
R23696 output.n19 output.n18 185
R23697 output.n34 output.n33 185
R23698 output.n32 output.n31 185
R23699 output.n23 output.n22 185
R23700 output.n26 output.n25 185
R23701 output.n73 output.n72 185
R23702 output.n71 output.n70 185
R23703 output.n50 output.n49 185
R23704 output.n65 output.n64 185
R23705 output.n63 output.n62 185
R23706 output.n54 output.n53 185
R23707 output.n57 output.n56 185
R23708 output.n105 output.n104 185
R23709 output.n103 output.n102 185
R23710 output.n82 output.n81 185
R23711 output.n97 output.n96 185
R23712 output.n95 output.n94 185
R23713 output.n86 output.n85 185
R23714 output.n89 output.n88 185
R23715 output.n137 output.n136 185
R23716 output.n135 output.n134 185
R23717 output.n114 output.n113 185
R23718 output.n129 output.n128 185
R23719 output.n127 output.n126 185
R23720 output.n118 output.n117 185
R23721 output.n121 output.n120 185
R23722 output.t18 output.n24 147.661
R23723 output.t19 output.n55 147.661
R23724 output.t16 output.n87 147.661
R23725 output.t17 output.n119 147.661
R23726 output.n41 output.n40 104.615
R23727 output.n40 output.n18 104.615
R23728 output.n33 output.n18 104.615
R23729 output.n33 output.n32 104.615
R23730 output.n32 output.n22 104.615
R23731 output.n25 output.n22 104.615
R23732 output.n72 output.n71 104.615
R23733 output.n71 output.n49 104.615
R23734 output.n64 output.n49 104.615
R23735 output.n64 output.n63 104.615
R23736 output.n63 output.n53 104.615
R23737 output.n56 output.n53 104.615
R23738 output.n104 output.n103 104.615
R23739 output.n103 output.n81 104.615
R23740 output.n96 output.n81 104.615
R23741 output.n96 output.n95 104.615
R23742 output.n95 output.n85 104.615
R23743 output.n88 output.n85 104.615
R23744 output.n136 output.n135 104.615
R23745 output.n135 output.n113 104.615
R23746 output.n128 output.n113 104.615
R23747 output.n128 output.n127 104.615
R23748 output.n127 output.n117 104.615
R23749 output.n120 output.n117 104.615
R23750 output.n1 output.t0 77.056
R23751 output.n14 output.t1 76.6694
R23752 output.n1 output.n0 72.7095
R23753 output.n3 output.n2 72.7095
R23754 output.n5 output.n4 72.7095
R23755 output.n7 output.n6 72.7095
R23756 output.n9 output.n8 72.7095
R23757 output.n11 output.n10 72.7095
R23758 output.n13 output.n12 72.7095
R23759 output.n25 output.t18 52.3082
R23760 output.n56 output.t19 52.3082
R23761 output.n88 output.t16 52.3082
R23762 output.n120 output.t17 52.3082
R23763 output.n26 output.n24 15.6674
R23764 output.n57 output.n55 15.6674
R23765 output.n89 output.n87 15.6674
R23766 output.n121 output.n119 15.6674
R23767 output.n27 output.n23 12.8005
R23768 output.n58 output.n54 12.8005
R23769 output.n90 output.n86 12.8005
R23770 output.n122 output.n118 12.8005
R23771 output.n31 output.n30 12.0247
R23772 output.n62 output.n61 12.0247
R23773 output.n94 output.n93 12.0247
R23774 output.n126 output.n125 12.0247
R23775 output.n34 output.n21 11.249
R23776 output.n65 output.n52 11.249
R23777 output.n97 output.n84 11.249
R23778 output.n129 output.n116 11.249
R23779 output.n35 output.n19 10.4732
R23780 output.n66 output.n50 10.4732
R23781 output.n98 output.n82 10.4732
R23782 output.n130 output.n114 10.4732
R23783 output.n39 output.n38 9.69747
R23784 output.n70 output.n69 9.69747
R23785 output.n102 output.n101 9.69747
R23786 output.n134 output.n133 9.69747
R23787 output.n45 output.n44 9.45567
R23788 output.n76 output.n75 9.45567
R23789 output.n108 output.n107 9.45567
R23790 output.n140 output.n139 9.45567
R23791 output.n44 output.n43 9.3005
R23792 output.n17 output.n16 9.3005
R23793 output.n38 output.n37 9.3005
R23794 output.n36 output.n35 9.3005
R23795 output.n21 output.n20 9.3005
R23796 output.n30 output.n29 9.3005
R23797 output.n28 output.n27 9.3005
R23798 output.n75 output.n74 9.3005
R23799 output.n48 output.n47 9.3005
R23800 output.n69 output.n68 9.3005
R23801 output.n67 output.n66 9.3005
R23802 output.n52 output.n51 9.3005
R23803 output.n61 output.n60 9.3005
R23804 output.n59 output.n58 9.3005
R23805 output.n107 output.n106 9.3005
R23806 output.n80 output.n79 9.3005
R23807 output.n101 output.n100 9.3005
R23808 output.n99 output.n98 9.3005
R23809 output.n84 output.n83 9.3005
R23810 output.n93 output.n92 9.3005
R23811 output.n91 output.n90 9.3005
R23812 output.n139 output.n138 9.3005
R23813 output.n112 output.n111 9.3005
R23814 output.n133 output.n132 9.3005
R23815 output.n131 output.n130 9.3005
R23816 output.n116 output.n115 9.3005
R23817 output.n125 output.n124 9.3005
R23818 output.n123 output.n122 9.3005
R23819 output.n42 output.n17 8.92171
R23820 output.n73 output.n48 8.92171
R23821 output.n105 output.n80 8.92171
R23822 output.n137 output.n112 8.92171
R23823 output output.n141 8.15037
R23824 output.n43 output.n15 8.14595
R23825 output.n74 output.n46 8.14595
R23826 output.n106 output.n78 8.14595
R23827 output.n138 output.n110 8.14595
R23828 output.n45 output.n15 5.81868
R23829 output.n76 output.n46 5.81868
R23830 output.n108 output.n78 5.81868
R23831 output.n140 output.n110 5.81868
R23832 output.n43 output.n42 5.04292
R23833 output.n74 output.n73 5.04292
R23834 output.n106 output.n105 5.04292
R23835 output.n138 output.n137 5.04292
R23836 output.n28 output.n24 4.38594
R23837 output.n59 output.n55 4.38594
R23838 output.n91 output.n87 4.38594
R23839 output.n123 output.n119 4.38594
R23840 output.n39 output.n17 4.26717
R23841 output.n70 output.n48 4.26717
R23842 output.n102 output.n80 4.26717
R23843 output.n134 output.n112 4.26717
R23844 output.n0 output.t10 3.9605
R23845 output.n0 output.t8 3.9605
R23846 output.n2 output.t15 3.9605
R23847 output.n2 output.t2 3.9605
R23848 output.n4 output.t4 3.9605
R23849 output.n4 output.t12 3.9605
R23850 output.n6 output.t14 3.9605
R23851 output.n6 output.t5 3.9605
R23852 output.n8 output.t6 3.9605
R23853 output.n8 output.t11 3.9605
R23854 output.n10 output.t13 3.9605
R23855 output.n10 output.t3 3.9605
R23856 output.n12 output.t9 3.9605
R23857 output.n12 output.t7 3.9605
R23858 output.n38 output.n19 3.49141
R23859 output.n69 output.n50 3.49141
R23860 output.n101 output.n82 3.49141
R23861 output.n133 output.n114 3.49141
R23862 output.n35 output.n34 2.71565
R23863 output.n66 output.n65 2.71565
R23864 output.n98 output.n97 2.71565
R23865 output.n130 output.n129 2.71565
R23866 output.n31 output.n21 1.93989
R23867 output.n62 output.n52 1.93989
R23868 output.n94 output.n84 1.93989
R23869 output.n126 output.n116 1.93989
R23870 output.n30 output.n23 1.16414
R23871 output.n61 output.n54 1.16414
R23872 output.n93 output.n86 1.16414
R23873 output.n125 output.n118 1.16414
R23874 output.n141 output.n109 0.962709
R23875 output.n109 output.n77 0.962709
R23876 output.n27 output.n26 0.388379
R23877 output.n58 output.n57 0.388379
R23878 output.n90 output.n89 0.388379
R23879 output.n122 output.n121 0.388379
R23880 output.n14 output.n13 0.387128
R23881 output.n13 output.n11 0.387128
R23882 output.n11 output.n9 0.387128
R23883 output.n9 output.n7 0.387128
R23884 output.n7 output.n5 0.387128
R23885 output.n5 output.n3 0.387128
R23886 output.n3 output.n1 0.387128
R23887 output.n44 output.n16 0.155672
R23888 output.n37 output.n16 0.155672
R23889 output.n37 output.n36 0.155672
R23890 output.n36 output.n20 0.155672
R23891 output.n29 output.n20 0.155672
R23892 output.n29 output.n28 0.155672
R23893 output.n75 output.n47 0.155672
R23894 output.n68 output.n47 0.155672
R23895 output.n68 output.n67 0.155672
R23896 output.n67 output.n51 0.155672
R23897 output.n60 output.n51 0.155672
R23898 output.n60 output.n59 0.155672
R23899 output.n107 output.n79 0.155672
R23900 output.n100 output.n79 0.155672
R23901 output.n100 output.n99 0.155672
R23902 output.n99 output.n83 0.155672
R23903 output.n92 output.n83 0.155672
R23904 output.n92 output.n91 0.155672
R23905 output.n139 output.n111 0.155672
R23906 output.n132 output.n111 0.155672
R23907 output.n132 output.n131 0.155672
R23908 output.n131 output.n115 0.155672
R23909 output.n124 output.n115 0.155672
R23910 output.n124 output.n123 0.155672
R23911 output output.n14 0.126227
R23912 diffpairibias.n0 diffpairibias.t18 436.822
R23913 diffpairibias.n21 diffpairibias.t19 435.479
R23914 diffpairibias.n20 diffpairibias.t16 435.479
R23915 diffpairibias.n19 diffpairibias.t17 435.479
R23916 diffpairibias.n18 diffpairibias.t21 435.479
R23917 diffpairibias.n0 diffpairibias.t22 435.479
R23918 diffpairibias.n1 diffpairibias.t20 435.479
R23919 diffpairibias.n2 diffpairibias.t23 435.479
R23920 diffpairibias.n10 diffpairibias.t0 377.536
R23921 diffpairibias.n10 diffpairibias.t8 376.193
R23922 diffpairibias.n11 diffpairibias.t10 376.193
R23923 diffpairibias.n12 diffpairibias.t6 376.193
R23924 diffpairibias.n13 diffpairibias.t2 376.193
R23925 diffpairibias.n14 diffpairibias.t12 376.193
R23926 diffpairibias.n15 diffpairibias.t4 376.193
R23927 diffpairibias.n16 diffpairibias.t14 376.193
R23928 diffpairibias.n3 diffpairibias.t1 113.368
R23929 diffpairibias.n3 diffpairibias.t9 112.698
R23930 diffpairibias.n4 diffpairibias.t11 112.698
R23931 diffpairibias.n5 diffpairibias.t7 112.698
R23932 diffpairibias.n6 diffpairibias.t3 112.698
R23933 diffpairibias.n7 diffpairibias.t13 112.698
R23934 diffpairibias.n8 diffpairibias.t5 112.698
R23935 diffpairibias.n9 diffpairibias.t15 112.698
R23936 diffpairibias.n17 diffpairibias.n16 4.77242
R23937 diffpairibias.n17 diffpairibias.n9 4.30807
R23938 diffpairibias.n18 diffpairibias.n17 4.13945
R23939 diffpairibias.n16 diffpairibias.n15 1.34352
R23940 diffpairibias.n15 diffpairibias.n14 1.34352
R23941 diffpairibias.n14 diffpairibias.n13 1.34352
R23942 diffpairibias.n13 diffpairibias.n12 1.34352
R23943 diffpairibias.n12 diffpairibias.n11 1.34352
R23944 diffpairibias.n11 diffpairibias.n10 1.34352
R23945 diffpairibias.n2 diffpairibias.n1 1.34352
R23946 diffpairibias.n1 diffpairibias.n0 1.34352
R23947 diffpairibias.n19 diffpairibias.n18 1.34352
R23948 diffpairibias.n20 diffpairibias.n19 1.34352
R23949 diffpairibias.n21 diffpairibias.n20 1.34352
R23950 diffpairibias.n22 diffpairibias.n21 0.862419
R23951 diffpairibias diffpairibias.n22 0.684875
R23952 diffpairibias.n9 diffpairibias.n8 0.672012
R23953 diffpairibias.n8 diffpairibias.n7 0.672012
R23954 diffpairibias.n7 diffpairibias.n6 0.672012
R23955 diffpairibias.n6 diffpairibias.n5 0.672012
R23956 diffpairibias.n5 diffpairibias.n4 0.672012
R23957 diffpairibias.n4 diffpairibias.n3 0.672012
R23958 diffpairibias.n22 diffpairibias.n2 0.190907
R23959 outputibias.n27 outputibias.n1 289.615
R23960 outputibias.n58 outputibias.n32 289.615
R23961 outputibias.n90 outputibias.n64 289.615
R23962 outputibias.n122 outputibias.n96 289.615
R23963 outputibias.n28 outputibias.n27 185
R23964 outputibias.n26 outputibias.n25 185
R23965 outputibias.n5 outputibias.n4 185
R23966 outputibias.n20 outputibias.n19 185
R23967 outputibias.n18 outputibias.n17 185
R23968 outputibias.n9 outputibias.n8 185
R23969 outputibias.n12 outputibias.n11 185
R23970 outputibias.n59 outputibias.n58 185
R23971 outputibias.n57 outputibias.n56 185
R23972 outputibias.n36 outputibias.n35 185
R23973 outputibias.n51 outputibias.n50 185
R23974 outputibias.n49 outputibias.n48 185
R23975 outputibias.n40 outputibias.n39 185
R23976 outputibias.n43 outputibias.n42 185
R23977 outputibias.n91 outputibias.n90 185
R23978 outputibias.n89 outputibias.n88 185
R23979 outputibias.n68 outputibias.n67 185
R23980 outputibias.n83 outputibias.n82 185
R23981 outputibias.n81 outputibias.n80 185
R23982 outputibias.n72 outputibias.n71 185
R23983 outputibias.n75 outputibias.n74 185
R23984 outputibias.n123 outputibias.n122 185
R23985 outputibias.n121 outputibias.n120 185
R23986 outputibias.n100 outputibias.n99 185
R23987 outputibias.n115 outputibias.n114 185
R23988 outputibias.n113 outputibias.n112 185
R23989 outputibias.n104 outputibias.n103 185
R23990 outputibias.n107 outputibias.n106 185
R23991 outputibias.n0 outputibias.t8 178.945
R23992 outputibias.n133 outputibias.t11 177.018
R23993 outputibias.n132 outputibias.t9 177.018
R23994 outputibias.n0 outputibias.t10 177.018
R23995 outputibias.t7 outputibias.n10 147.661
R23996 outputibias.t1 outputibias.n41 147.661
R23997 outputibias.t3 outputibias.n73 147.661
R23998 outputibias.t5 outputibias.n105 147.661
R23999 outputibias.n128 outputibias.t6 132.363
R24000 outputibias.n128 outputibias.t0 130.436
R24001 outputibias.n129 outputibias.t2 130.436
R24002 outputibias.n130 outputibias.t4 130.436
R24003 outputibias.n27 outputibias.n26 104.615
R24004 outputibias.n26 outputibias.n4 104.615
R24005 outputibias.n19 outputibias.n4 104.615
R24006 outputibias.n19 outputibias.n18 104.615
R24007 outputibias.n18 outputibias.n8 104.615
R24008 outputibias.n11 outputibias.n8 104.615
R24009 outputibias.n58 outputibias.n57 104.615
R24010 outputibias.n57 outputibias.n35 104.615
R24011 outputibias.n50 outputibias.n35 104.615
R24012 outputibias.n50 outputibias.n49 104.615
R24013 outputibias.n49 outputibias.n39 104.615
R24014 outputibias.n42 outputibias.n39 104.615
R24015 outputibias.n90 outputibias.n89 104.615
R24016 outputibias.n89 outputibias.n67 104.615
R24017 outputibias.n82 outputibias.n67 104.615
R24018 outputibias.n82 outputibias.n81 104.615
R24019 outputibias.n81 outputibias.n71 104.615
R24020 outputibias.n74 outputibias.n71 104.615
R24021 outputibias.n122 outputibias.n121 104.615
R24022 outputibias.n121 outputibias.n99 104.615
R24023 outputibias.n114 outputibias.n99 104.615
R24024 outputibias.n114 outputibias.n113 104.615
R24025 outputibias.n113 outputibias.n103 104.615
R24026 outputibias.n106 outputibias.n103 104.615
R24027 outputibias.n63 outputibias.n31 95.6354
R24028 outputibias.n63 outputibias.n62 94.6732
R24029 outputibias.n95 outputibias.n94 94.6732
R24030 outputibias.n127 outputibias.n126 94.6732
R24031 outputibias.n11 outputibias.t7 52.3082
R24032 outputibias.n42 outputibias.t1 52.3082
R24033 outputibias.n74 outputibias.t3 52.3082
R24034 outputibias.n106 outputibias.t5 52.3082
R24035 outputibias.n12 outputibias.n10 15.6674
R24036 outputibias.n43 outputibias.n41 15.6674
R24037 outputibias.n75 outputibias.n73 15.6674
R24038 outputibias.n107 outputibias.n105 15.6674
R24039 outputibias.n13 outputibias.n9 12.8005
R24040 outputibias.n44 outputibias.n40 12.8005
R24041 outputibias.n76 outputibias.n72 12.8005
R24042 outputibias.n108 outputibias.n104 12.8005
R24043 outputibias.n17 outputibias.n16 12.0247
R24044 outputibias.n48 outputibias.n47 12.0247
R24045 outputibias.n80 outputibias.n79 12.0247
R24046 outputibias.n112 outputibias.n111 12.0247
R24047 outputibias.n20 outputibias.n7 11.249
R24048 outputibias.n51 outputibias.n38 11.249
R24049 outputibias.n83 outputibias.n70 11.249
R24050 outputibias.n115 outputibias.n102 11.249
R24051 outputibias.n21 outputibias.n5 10.4732
R24052 outputibias.n52 outputibias.n36 10.4732
R24053 outputibias.n84 outputibias.n68 10.4732
R24054 outputibias.n116 outputibias.n100 10.4732
R24055 outputibias.n25 outputibias.n24 9.69747
R24056 outputibias.n56 outputibias.n55 9.69747
R24057 outputibias.n88 outputibias.n87 9.69747
R24058 outputibias.n120 outputibias.n119 9.69747
R24059 outputibias.n31 outputibias.n30 9.45567
R24060 outputibias.n62 outputibias.n61 9.45567
R24061 outputibias.n94 outputibias.n93 9.45567
R24062 outputibias.n126 outputibias.n125 9.45567
R24063 outputibias.n30 outputibias.n29 9.3005
R24064 outputibias.n3 outputibias.n2 9.3005
R24065 outputibias.n24 outputibias.n23 9.3005
R24066 outputibias.n22 outputibias.n21 9.3005
R24067 outputibias.n7 outputibias.n6 9.3005
R24068 outputibias.n16 outputibias.n15 9.3005
R24069 outputibias.n14 outputibias.n13 9.3005
R24070 outputibias.n61 outputibias.n60 9.3005
R24071 outputibias.n34 outputibias.n33 9.3005
R24072 outputibias.n55 outputibias.n54 9.3005
R24073 outputibias.n53 outputibias.n52 9.3005
R24074 outputibias.n38 outputibias.n37 9.3005
R24075 outputibias.n47 outputibias.n46 9.3005
R24076 outputibias.n45 outputibias.n44 9.3005
R24077 outputibias.n93 outputibias.n92 9.3005
R24078 outputibias.n66 outputibias.n65 9.3005
R24079 outputibias.n87 outputibias.n86 9.3005
R24080 outputibias.n85 outputibias.n84 9.3005
R24081 outputibias.n70 outputibias.n69 9.3005
R24082 outputibias.n79 outputibias.n78 9.3005
R24083 outputibias.n77 outputibias.n76 9.3005
R24084 outputibias.n125 outputibias.n124 9.3005
R24085 outputibias.n98 outputibias.n97 9.3005
R24086 outputibias.n119 outputibias.n118 9.3005
R24087 outputibias.n117 outputibias.n116 9.3005
R24088 outputibias.n102 outputibias.n101 9.3005
R24089 outputibias.n111 outputibias.n110 9.3005
R24090 outputibias.n109 outputibias.n108 9.3005
R24091 outputibias.n28 outputibias.n3 8.92171
R24092 outputibias.n59 outputibias.n34 8.92171
R24093 outputibias.n91 outputibias.n66 8.92171
R24094 outputibias.n123 outputibias.n98 8.92171
R24095 outputibias.n29 outputibias.n1 8.14595
R24096 outputibias.n60 outputibias.n32 8.14595
R24097 outputibias.n92 outputibias.n64 8.14595
R24098 outputibias.n124 outputibias.n96 8.14595
R24099 outputibias.n31 outputibias.n1 5.81868
R24100 outputibias.n62 outputibias.n32 5.81868
R24101 outputibias.n94 outputibias.n64 5.81868
R24102 outputibias.n126 outputibias.n96 5.81868
R24103 outputibias.n131 outputibias.n130 5.20947
R24104 outputibias.n29 outputibias.n28 5.04292
R24105 outputibias.n60 outputibias.n59 5.04292
R24106 outputibias.n92 outputibias.n91 5.04292
R24107 outputibias.n124 outputibias.n123 5.04292
R24108 outputibias.n131 outputibias.n127 4.42209
R24109 outputibias.n14 outputibias.n10 4.38594
R24110 outputibias.n45 outputibias.n41 4.38594
R24111 outputibias.n77 outputibias.n73 4.38594
R24112 outputibias.n109 outputibias.n105 4.38594
R24113 outputibias.n132 outputibias.n131 4.28454
R24114 outputibias.n25 outputibias.n3 4.26717
R24115 outputibias.n56 outputibias.n34 4.26717
R24116 outputibias.n88 outputibias.n66 4.26717
R24117 outputibias.n120 outputibias.n98 4.26717
R24118 outputibias.n24 outputibias.n5 3.49141
R24119 outputibias.n55 outputibias.n36 3.49141
R24120 outputibias.n87 outputibias.n68 3.49141
R24121 outputibias.n119 outputibias.n100 3.49141
R24122 outputibias.n21 outputibias.n20 2.71565
R24123 outputibias.n52 outputibias.n51 2.71565
R24124 outputibias.n84 outputibias.n83 2.71565
R24125 outputibias.n116 outputibias.n115 2.71565
R24126 outputibias.n17 outputibias.n7 1.93989
R24127 outputibias.n48 outputibias.n38 1.93989
R24128 outputibias.n80 outputibias.n70 1.93989
R24129 outputibias.n112 outputibias.n102 1.93989
R24130 outputibias.n130 outputibias.n129 1.9266
R24131 outputibias.n129 outputibias.n128 1.9266
R24132 outputibias.n133 outputibias.n132 1.92658
R24133 outputibias.n134 outputibias.n133 1.29913
R24134 outputibias.n16 outputibias.n9 1.16414
R24135 outputibias.n47 outputibias.n40 1.16414
R24136 outputibias.n79 outputibias.n72 1.16414
R24137 outputibias.n111 outputibias.n104 1.16414
R24138 outputibias.n127 outputibias.n95 0.962709
R24139 outputibias.n95 outputibias.n63 0.962709
R24140 outputibias.n13 outputibias.n12 0.388379
R24141 outputibias.n44 outputibias.n43 0.388379
R24142 outputibias.n76 outputibias.n75 0.388379
R24143 outputibias.n108 outputibias.n107 0.388379
R24144 outputibias.n134 outputibias.n0 0.337251
R24145 outputibias outputibias.n134 0.302375
R24146 outputibias.n30 outputibias.n2 0.155672
R24147 outputibias.n23 outputibias.n2 0.155672
R24148 outputibias.n23 outputibias.n22 0.155672
R24149 outputibias.n22 outputibias.n6 0.155672
R24150 outputibias.n15 outputibias.n6 0.155672
R24151 outputibias.n15 outputibias.n14 0.155672
R24152 outputibias.n61 outputibias.n33 0.155672
R24153 outputibias.n54 outputibias.n33 0.155672
R24154 outputibias.n54 outputibias.n53 0.155672
R24155 outputibias.n53 outputibias.n37 0.155672
R24156 outputibias.n46 outputibias.n37 0.155672
R24157 outputibias.n46 outputibias.n45 0.155672
R24158 outputibias.n93 outputibias.n65 0.155672
R24159 outputibias.n86 outputibias.n65 0.155672
R24160 outputibias.n86 outputibias.n85 0.155672
R24161 outputibias.n85 outputibias.n69 0.155672
R24162 outputibias.n78 outputibias.n69 0.155672
R24163 outputibias.n78 outputibias.n77 0.155672
R24164 outputibias.n125 outputibias.n97 0.155672
R24165 outputibias.n118 outputibias.n97 0.155672
R24166 outputibias.n118 outputibias.n117 0.155672
R24167 outputibias.n117 outputibias.n101 0.155672
R24168 outputibias.n110 outputibias.n101 0.155672
R24169 outputibias.n110 outputibias.n109 0.155672
C0 commonsourceibias output 0.006808f
C1 minus diffpairibias 4.33e-19
C2 CSoutput minus 2.93202f
C3 vdd plus 0.080199f
C4 plus diffpairibias 4.56e-19
C5 commonsourceibias outputibias 0.003832f
C6 vdd commonsourceibias 0.004218f
C7 CSoutput plus 0.894663f
C8 commonsourceibias diffpairibias 0.06482f
C9 CSoutput commonsourceibias 66.33679f
C10 minus plus 9.97292f
C11 minus commonsourceibias 0.460231f
C12 plus commonsourceibias 0.415048f
C13 output outputibias 2.34152f
C14 vdd output 7.23429f
C15 CSoutput output 6.13881f
C16 CSoutput outputibias 0.032386f
C17 vdd CSoutput 92.295f
C18 diffpairibias gnd 48.980137f
C19 outputibias gnd 32.465668f
C20 output gnd 15.47879f
C21 commonsourceibias gnd 0.222236p
C22 plus gnd 36.812397f
C23 minus gnd 30.0463f
C24 CSoutput gnd 0.143669p
C25 vdd gnd 0.411227p
C26 outputibias.t10 gnd 0.11477f
C27 outputibias.t8 gnd 0.115567f
C28 outputibias.n0 gnd 0.130108f
C29 outputibias.n1 gnd 0.001372f
C30 outputibias.n2 gnd 9.76e-19
C31 outputibias.n3 gnd 5.24e-19
C32 outputibias.n4 gnd 0.001239f
C33 outputibias.n5 gnd 5.55e-19
C34 outputibias.n6 gnd 9.76e-19
C35 outputibias.n7 gnd 5.24e-19
C36 outputibias.n8 gnd 0.001239f
C37 outputibias.n9 gnd 5.55e-19
C38 outputibias.n10 gnd 0.004176f
C39 outputibias.t7 gnd 0.00202f
C40 outputibias.n11 gnd 9.3e-19
C41 outputibias.n12 gnd 7.32e-19
C42 outputibias.n13 gnd 5.24e-19
C43 outputibias.n14 gnd 0.02322f
C44 outputibias.n15 gnd 9.76e-19
C45 outputibias.n16 gnd 5.24e-19
C46 outputibias.n17 gnd 5.55e-19
C47 outputibias.n18 gnd 0.001239f
C48 outputibias.n19 gnd 0.001239f
C49 outputibias.n20 gnd 5.55e-19
C50 outputibias.n21 gnd 5.24e-19
C51 outputibias.n22 gnd 9.76e-19
C52 outputibias.n23 gnd 9.76e-19
C53 outputibias.n24 gnd 5.24e-19
C54 outputibias.n25 gnd 5.55e-19
C55 outputibias.n26 gnd 0.001239f
C56 outputibias.n27 gnd 0.002683f
C57 outputibias.n28 gnd 5.55e-19
C58 outputibias.n29 gnd 5.24e-19
C59 outputibias.n30 gnd 0.002256f
C60 outputibias.n31 gnd 0.005781f
C61 outputibias.n32 gnd 0.001372f
C62 outputibias.n33 gnd 9.76e-19
C63 outputibias.n34 gnd 5.24e-19
C64 outputibias.n35 gnd 0.001239f
C65 outputibias.n36 gnd 5.55e-19
C66 outputibias.n37 gnd 9.76e-19
C67 outputibias.n38 gnd 5.24e-19
C68 outputibias.n39 gnd 0.001239f
C69 outputibias.n40 gnd 5.55e-19
C70 outputibias.n41 gnd 0.004176f
C71 outputibias.t1 gnd 0.00202f
C72 outputibias.n42 gnd 9.3e-19
C73 outputibias.n43 gnd 7.32e-19
C74 outputibias.n44 gnd 5.24e-19
C75 outputibias.n45 gnd 0.02322f
C76 outputibias.n46 gnd 9.76e-19
C77 outputibias.n47 gnd 5.24e-19
C78 outputibias.n48 gnd 5.55e-19
C79 outputibias.n49 gnd 0.001239f
C80 outputibias.n50 gnd 0.001239f
C81 outputibias.n51 gnd 5.55e-19
C82 outputibias.n52 gnd 5.24e-19
C83 outputibias.n53 gnd 9.76e-19
C84 outputibias.n54 gnd 9.76e-19
C85 outputibias.n55 gnd 5.24e-19
C86 outputibias.n56 gnd 5.55e-19
C87 outputibias.n57 gnd 0.001239f
C88 outputibias.n58 gnd 0.002683f
C89 outputibias.n59 gnd 5.55e-19
C90 outputibias.n60 gnd 5.24e-19
C91 outputibias.n61 gnd 0.002256f
C92 outputibias.n62 gnd 0.005197f
C93 outputibias.n63 gnd 0.121892f
C94 outputibias.n64 gnd 0.001372f
C95 outputibias.n65 gnd 9.76e-19
C96 outputibias.n66 gnd 5.24e-19
C97 outputibias.n67 gnd 0.001239f
C98 outputibias.n68 gnd 5.55e-19
C99 outputibias.n69 gnd 9.76e-19
C100 outputibias.n70 gnd 5.24e-19
C101 outputibias.n71 gnd 0.001239f
C102 outputibias.n72 gnd 5.55e-19
C103 outputibias.n73 gnd 0.004176f
C104 outputibias.t3 gnd 0.00202f
C105 outputibias.n74 gnd 9.3e-19
C106 outputibias.n75 gnd 7.32e-19
C107 outputibias.n76 gnd 5.24e-19
C108 outputibias.n77 gnd 0.02322f
C109 outputibias.n78 gnd 9.76e-19
C110 outputibias.n79 gnd 5.24e-19
C111 outputibias.n80 gnd 5.55e-19
C112 outputibias.n81 gnd 0.001239f
C113 outputibias.n82 gnd 0.001239f
C114 outputibias.n83 gnd 5.55e-19
C115 outputibias.n84 gnd 5.24e-19
C116 outputibias.n85 gnd 9.76e-19
C117 outputibias.n86 gnd 9.76e-19
C118 outputibias.n87 gnd 5.24e-19
C119 outputibias.n88 gnd 5.55e-19
C120 outputibias.n89 gnd 0.001239f
C121 outputibias.n90 gnd 0.002683f
C122 outputibias.n91 gnd 5.55e-19
C123 outputibias.n92 gnd 5.24e-19
C124 outputibias.n93 gnd 0.002256f
C125 outputibias.n94 gnd 0.005197f
C126 outputibias.n95 gnd 0.064513f
C127 outputibias.n96 gnd 0.001372f
C128 outputibias.n97 gnd 9.76e-19
C129 outputibias.n98 gnd 5.24e-19
C130 outputibias.n99 gnd 0.001239f
C131 outputibias.n100 gnd 5.55e-19
C132 outputibias.n101 gnd 9.76e-19
C133 outputibias.n102 gnd 5.24e-19
C134 outputibias.n103 gnd 0.001239f
C135 outputibias.n104 gnd 5.55e-19
C136 outputibias.n105 gnd 0.004176f
C137 outputibias.t5 gnd 0.00202f
C138 outputibias.n106 gnd 9.3e-19
C139 outputibias.n107 gnd 7.32e-19
C140 outputibias.n108 gnd 5.24e-19
C141 outputibias.n109 gnd 0.02322f
C142 outputibias.n110 gnd 9.76e-19
C143 outputibias.n111 gnd 5.24e-19
C144 outputibias.n112 gnd 5.55e-19
C145 outputibias.n113 gnd 0.001239f
C146 outputibias.n114 gnd 0.001239f
C147 outputibias.n115 gnd 5.55e-19
C148 outputibias.n116 gnd 5.24e-19
C149 outputibias.n117 gnd 9.76e-19
C150 outputibias.n118 gnd 9.76e-19
C151 outputibias.n119 gnd 5.24e-19
C152 outputibias.n120 gnd 5.55e-19
C153 outputibias.n121 gnd 0.001239f
C154 outputibias.n122 gnd 0.002683f
C155 outputibias.n123 gnd 5.55e-19
C156 outputibias.n124 gnd 5.24e-19
C157 outputibias.n125 gnd 0.002256f
C158 outputibias.n126 gnd 0.005197f
C159 outputibias.n127 gnd 0.084814f
C160 outputibias.t4 gnd 0.108319f
C161 outputibias.t2 gnd 0.108319f
C162 outputibias.t0 gnd 0.108319f
C163 outputibias.t6 gnd 0.109238f
C164 outputibias.n128 gnd 0.134674f
C165 outputibias.n129 gnd 0.07244f
C166 outputibias.n130 gnd 0.079818f
C167 outputibias.n131 gnd 0.164901f
C168 outputibias.t9 gnd 0.11477f
C169 outputibias.n132 gnd 0.067481f
C170 outputibias.t11 gnd 0.11477f
C171 outputibias.n133 gnd 0.065115f
C172 outputibias.n134 gnd 0.029159f
C173 diffpairibias.t18 gnd 0.087401f
C174 diffpairibias.t22 gnd 0.087239f
C175 diffpairibias.n0 gnd 0.102784f
C176 diffpairibias.t20 gnd 0.087239f
C177 diffpairibias.n1 gnd 0.050171f
C178 diffpairibias.t23 gnd 0.087239f
C179 diffpairibias.n2 gnd 0.039841f
C180 diffpairibias.t1 gnd 0.083757f
C181 diffpairibias.t9 gnd 0.083392f
C182 diffpairibias.n3 gnd 0.131682f
C183 diffpairibias.t11 gnd 0.083392f
C184 diffpairibias.n4 gnd 0.07027f
C185 diffpairibias.t7 gnd 0.083392f
C186 diffpairibias.n5 gnd 0.07027f
C187 diffpairibias.t3 gnd 0.083392f
C188 diffpairibias.n6 gnd 0.07027f
C189 diffpairibias.t13 gnd 0.083392f
C190 diffpairibias.n7 gnd 0.07027f
C191 diffpairibias.t5 gnd 0.083392f
C192 diffpairibias.n8 gnd 0.07027f
C193 diffpairibias.t15 gnd 0.083392f
C194 diffpairibias.n9 gnd 0.099771f
C195 diffpairibias.t0 gnd 0.08427f
C196 diffpairibias.t8 gnd 0.084123f
C197 diffpairibias.n10 gnd 0.091784f
C198 diffpairibias.t10 gnd 0.084123f
C199 diffpairibias.n11 gnd 0.050681f
C200 diffpairibias.t6 gnd 0.084123f
C201 diffpairibias.n12 gnd 0.050681f
C202 diffpairibias.t2 gnd 0.084123f
C203 diffpairibias.n13 gnd 0.050681f
C204 diffpairibias.t12 gnd 0.084123f
C205 diffpairibias.n14 gnd 0.050681f
C206 diffpairibias.t4 gnd 0.084123f
C207 diffpairibias.n15 gnd 0.050681f
C208 diffpairibias.t14 gnd 0.084123f
C209 diffpairibias.n16 gnd 0.059977f
C210 diffpairibias.n17 gnd 0.226448f
C211 diffpairibias.t21 gnd 0.087239f
C212 diffpairibias.n18 gnd 0.050181f
C213 diffpairibias.t17 gnd 0.087239f
C214 diffpairibias.n19 gnd 0.050171f
C215 diffpairibias.t16 gnd 0.087239f
C216 diffpairibias.n20 gnd 0.050171f
C217 diffpairibias.t19 gnd 0.087239f
C218 diffpairibias.n21 gnd 0.045859f
C219 diffpairibias.n22 gnd 0.046268f
C220 output.t0 gnd 0.464308f
C221 output.t10 gnd 0.044422f
C222 output.t8 gnd 0.044422f
C223 output.n0 gnd 0.364624f
C224 output.n1 gnd 0.614102f
C225 output.t15 gnd 0.044422f
C226 output.t2 gnd 0.044422f
C227 output.n2 gnd 0.364624f
C228 output.n3 gnd 0.350265f
C229 output.t4 gnd 0.044422f
C230 output.t12 gnd 0.044422f
C231 output.n4 gnd 0.364624f
C232 output.n5 gnd 0.350265f
C233 output.t14 gnd 0.044422f
C234 output.t5 gnd 0.044422f
C235 output.n6 gnd 0.364624f
C236 output.n7 gnd 0.350265f
C237 output.t6 gnd 0.044422f
C238 output.t11 gnd 0.044422f
C239 output.n8 gnd 0.364624f
C240 output.n9 gnd 0.350265f
C241 output.t13 gnd 0.044422f
C242 output.t3 gnd 0.044422f
C243 output.n10 gnd 0.364624f
C244 output.n11 gnd 0.350265f
C245 output.t9 gnd 0.044422f
C246 output.t7 gnd 0.044422f
C247 output.n12 gnd 0.364624f
C248 output.n13 gnd 0.350265f
C249 output.t1 gnd 0.462979f
C250 output.n14 gnd 0.28994f
C251 output.n15 gnd 0.015803f
C252 output.n16 gnd 0.011243f
C253 output.n17 gnd 0.006041f
C254 output.n18 gnd 0.01428f
C255 output.n19 gnd 0.006397f
C256 output.n20 gnd 0.011243f
C257 output.n21 gnd 0.006041f
C258 output.n22 gnd 0.01428f
C259 output.n23 gnd 0.006397f
C260 output.n24 gnd 0.048111f
C261 output.t18 gnd 0.023274f
C262 output.n25 gnd 0.01071f
C263 output.n26 gnd 0.008435f
C264 output.n27 gnd 0.006041f
C265 output.n28 gnd 0.267512f
C266 output.n29 gnd 0.011243f
C267 output.n30 gnd 0.006041f
C268 output.n31 gnd 0.006397f
C269 output.n32 gnd 0.01428f
C270 output.n33 gnd 0.01428f
C271 output.n34 gnd 0.006397f
C272 output.n35 gnd 0.006041f
C273 output.n36 gnd 0.011243f
C274 output.n37 gnd 0.011243f
C275 output.n38 gnd 0.006041f
C276 output.n39 gnd 0.006397f
C277 output.n40 gnd 0.01428f
C278 output.n41 gnd 0.030913f
C279 output.n42 gnd 0.006397f
C280 output.n43 gnd 0.006041f
C281 output.n44 gnd 0.025987f
C282 output.n45 gnd 0.097665f
C283 output.n46 gnd 0.015803f
C284 output.n47 gnd 0.011243f
C285 output.n48 gnd 0.006041f
C286 output.n49 gnd 0.01428f
C287 output.n50 gnd 0.006397f
C288 output.n51 gnd 0.011243f
C289 output.n52 gnd 0.006041f
C290 output.n53 gnd 0.01428f
C291 output.n54 gnd 0.006397f
C292 output.n55 gnd 0.048111f
C293 output.t19 gnd 0.023274f
C294 output.n56 gnd 0.01071f
C295 output.n57 gnd 0.008435f
C296 output.n58 gnd 0.006041f
C297 output.n59 gnd 0.267512f
C298 output.n60 gnd 0.011243f
C299 output.n61 gnd 0.006041f
C300 output.n62 gnd 0.006397f
C301 output.n63 gnd 0.01428f
C302 output.n64 gnd 0.01428f
C303 output.n65 gnd 0.006397f
C304 output.n66 gnd 0.006041f
C305 output.n67 gnd 0.011243f
C306 output.n68 gnd 0.011243f
C307 output.n69 gnd 0.006041f
C308 output.n70 gnd 0.006397f
C309 output.n71 gnd 0.01428f
C310 output.n72 gnd 0.030913f
C311 output.n73 gnd 0.006397f
C312 output.n74 gnd 0.006041f
C313 output.n75 gnd 0.025987f
C314 output.n76 gnd 0.09306f
C315 output.n77 gnd 1.65264f
C316 output.n78 gnd 0.015803f
C317 output.n79 gnd 0.011243f
C318 output.n80 gnd 0.006041f
C319 output.n81 gnd 0.01428f
C320 output.n82 gnd 0.006397f
C321 output.n83 gnd 0.011243f
C322 output.n84 gnd 0.006041f
C323 output.n85 gnd 0.01428f
C324 output.n86 gnd 0.006397f
C325 output.n87 gnd 0.048111f
C326 output.t16 gnd 0.023274f
C327 output.n88 gnd 0.01071f
C328 output.n89 gnd 0.008435f
C329 output.n90 gnd 0.006041f
C330 output.n91 gnd 0.267512f
C331 output.n92 gnd 0.011243f
C332 output.n93 gnd 0.006041f
C333 output.n94 gnd 0.006397f
C334 output.n95 gnd 0.01428f
C335 output.n96 gnd 0.01428f
C336 output.n97 gnd 0.006397f
C337 output.n98 gnd 0.006041f
C338 output.n99 gnd 0.011243f
C339 output.n100 gnd 0.011243f
C340 output.n101 gnd 0.006041f
C341 output.n102 gnd 0.006397f
C342 output.n103 gnd 0.01428f
C343 output.n104 gnd 0.030913f
C344 output.n105 gnd 0.006397f
C345 output.n106 gnd 0.006041f
C346 output.n107 gnd 0.025987f
C347 output.n108 gnd 0.09306f
C348 output.n109 gnd 0.713089f
C349 output.n110 gnd 0.015803f
C350 output.n111 gnd 0.011243f
C351 output.n112 gnd 0.006041f
C352 output.n113 gnd 0.01428f
C353 output.n114 gnd 0.006397f
C354 output.n115 gnd 0.011243f
C355 output.n116 gnd 0.006041f
C356 output.n117 gnd 0.01428f
C357 output.n118 gnd 0.006397f
C358 output.n119 gnd 0.048111f
C359 output.t17 gnd 0.023274f
C360 output.n120 gnd 0.01071f
C361 output.n121 gnd 0.008435f
C362 output.n122 gnd 0.006041f
C363 output.n123 gnd 0.267512f
C364 output.n124 gnd 0.011243f
C365 output.n125 gnd 0.006041f
C366 output.n126 gnd 0.006397f
C367 output.n127 gnd 0.01428f
C368 output.n128 gnd 0.01428f
C369 output.n129 gnd 0.006397f
C370 output.n130 gnd 0.006041f
C371 output.n131 gnd 0.011243f
C372 output.n132 gnd 0.011243f
C373 output.n133 gnd 0.006041f
C374 output.n134 gnd 0.006397f
C375 output.n135 gnd 0.01428f
C376 output.n136 gnd 0.030913f
C377 output.n137 gnd 0.006397f
C378 output.n138 gnd 0.006041f
C379 output.n139 gnd 0.025987f
C380 output.n140 gnd 0.09306f
C381 output.n141 gnd 1.67353f
C382 a_n2318_8322.t25 gnd 39.602997f
C383 a_n2318_8322.t27 gnd 29.1868f
C384 a_n2318_8322.t26 gnd 19.7318f
C385 a_n2318_8322.t24 gnd 39.602997f
C386 a_n2318_8322.t12 gnd 0.095784f
C387 a_n2318_8322.t22 gnd 0.896867f
C388 a_n2318_8322.t10 gnd 0.095784f
C389 a_n2318_8322.t9 gnd 0.095784f
C390 a_n2318_8322.n0 gnd 0.674698f
C391 a_n2318_8322.n1 gnd 0.753876f
C392 a_n2318_8322.t19 gnd 0.095784f
C393 a_n2318_8322.t14 gnd 0.095784f
C394 a_n2318_8322.n2 gnd 0.674698f
C395 a_n2318_8322.n3 gnd 0.383035f
C396 a_n2318_8322.t17 gnd 0.095784f
C397 a_n2318_8322.t16 gnd 0.095784f
C398 a_n2318_8322.n4 gnd 0.674698f
C399 a_n2318_8322.n5 gnd 0.383035f
C400 a_n2318_8322.t8 gnd 0.895081f
C401 a_n2318_8322.n6 gnd 1.55131f
C402 a_n2318_8322.t3 gnd 0.896867f
C403 a_n2318_8322.t7 gnd 0.095784f
C404 a_n2318_8322.t6 gnd 0.095784f
C405 a_n2318_8322.n7 gnd 0.674698f
C406 a_n2318_8322.n8 gnd 0.753876f
C407 a_n2318_8322.t1 gnd 0.895081f
C408 a_n2318_8322.n9 gnd 0.379361f
C409 a_n2318_8322.t4 gnd 0.895081f
C410 a_n2318_8322.n10 gnd 0.379361f
C411 a_n2318_8322.t2 gnd 0.095784f
C412 a_n2318_8322.t0 gnd 0.095784f
C413 a_n2318_8322.n11 gnd 0.674698f
C414 a_n2318_8322.n12 gnd 0.383035f
C415 a_n2318_8322.t5 gnd 0.895081f
C416 a_n2318_8322.n13 gnd 1.07426f
C417 a_n2318_8322.n14 gnd 1.82616f
C418 a_n2318_8322.n15 gnd 3.71089f
C419 a_n2318_8322.t11 gnd 0.895081f
C420 a_n2318_8322.n16 gnd 0.881139f
C421 a_n2318_8322.t20 gnd 0.095784f
C422 a_n2318_8322.t13 gnd 0.095784f
C423 a_n2318_8322.n17 gnd 0.674698f
C424 a_n2318_8322.n18 gnd 0.383035f
C425 a_n2318_8322.t21 gnd 0.896865f
C426 a_n2318_8322.t18 gnd 0.095784f
C427 a_n2318_8322.t15 gnd 0.095784f
C428 a_n2318_8322.n19 gnd 0.674698f
C429 a_n2318_8322.n20 gnd 0.753878f
C430 a_n2318_8322.n21 gnd 0.383033f
C431 a_n2318_8322.n22 gnd 0.6747f
C432 a_n2318_8322.t23 gnd 0.095784f
C433 minus.n0 gnd 0.031734f
C434 minus.n1 gnd 0.007201f
C435 minus.n2 gnd 0.031734f
C436 minus.n3 gnd 0.007201f
C437 minus.n4 gnd 0.031734f
C438 minus.n5 gnd 0.007201f
C439 minus.n6 gnd 0.031734f
C440 minus.n7 gnd 0.007201f
C441 minus.n8 gnd 0.031734f
C442 minus.n9 gnd 0.007201f
C443 minus.t8 gnd 0.465132f
C444 minus.t7 gnd 0.44884f
C445 minus.n10 gnd 0.205883f
C446 minus.n11 gnd 0.184786f
C447 minus.n12 gnd 0.136614f
C448 minus.n13 gnd 0.031734f
C449 minus.t11 gnd 0.44884f
C450 minus.n14 gnd 0.199389f
C451 minus.n15 gnd 0.007201f
C452 minus.t10 gnd 0.44884f
C453 minus.n16 gnd 0.199389f
C454 minus.n17 gnd 0.031734f
C455 minus.n18 gnd 0.031734f
C456 minus.n19 gnd 0.031734f
C457 minus.t12 gnd 0.44884f
C458 minus.n20 gnd 0.199389f
C459 minus.n21 gnd 0.007201f
C460 minus.t20 gnd 0.44884f
C461 minus.n22 gnd 0.199389f
C462 minus.n23 gnd 0.031734f
C463 minus.n24 gnd 0.031734f
C464 minus.n25 gnd 0.031734f
C465 minus.t18 gnd 0.44884f
C466 minus.n26 gnd 0.199389f
C467 minus.n27 gnd 0.007201f
C468 minus.t25 gnd 0.44884f
C469 minus.n28 gnd 0.199389f
C470 minus.n29 gnd 0.031734f
C471 minus.n30 gnd 0.031734f
C472 minus.n31 gnd 0.031734f
C473 minus.t24 gnd 0.44884f
C474 minus.n32 gnd 0.199389f
C475 minus.n33 gnd 0.007201f
C476 minus.t14 gnd 0.44884f
C477 minus.n34 gnd 0.199389f
C478 minus.n35 gnd 0.031734f
C479 minus.n36 gnd 0.031734f
C480 minus.n37 gnd 0.031734f
C481 minus.t22 gnd 0.44884f
C482 minus.n38 gnd 0.199389f
C483 minus.n39 gnd 0.007201f
C484 minus.t19 gnd 0.44884f
C485 minus.n40 gnd 0.199682f
C486 minus.n41 gnd 0.367505f
C487 minus.n42 gnd 0.031734f
C488 minus.t13 gnd 0.44884f
C489 minus.t15 gnd 0.44884f
C490 minus.n43 gnd 0.031734f
C491 minus.t5 gnd 0.44884f
C492 minus.n44 gnd 0.199389f
C493 minus.n45 gnd 0.031734f
C494 minus.t6 gnd 0.44884f
C495 minus.t26 gnd 0.44884f
C496 minus.n46 gnd 0.199389f
C497 minus.n47 gnd 0.031734f
C498 minus.t21 gnd 0.44884f
C499 minus.t23 gnd 0.44884f
C500 minus.n48 gnd 0.199389f
C501 minus.n49 gnd 0.031734f
C502 minus.t16 gnd 0.44884f
C503 minus.t17 gnd 0.44884f
C504 minus.n50 gnd 0.199389f
C505 minus.n51 gnd 0.031734f
C506 minus.t9 gnd 0.44884f
C507 minus.t27 gnd 0.44884f
C508 minus.n52 gnd 0.205883f
C509 minus.t28 gnd 0.465132f
C510 minus.n53 gnd 0.184786f
C511 minus.n54 gnd 0.136614f
C512 minus.n55 gnd 0.007201f
C513 minus.n56 gnd 0.199389f
C514 minus.n57 gnd 0.007201f
C515 minus.n58 gnd 0.031734f
C516 minus.n59 gnd 0.031734f
C517 minus.n60 gnd 0.031734f
C518 minus.n61 gnd 0.007201f
C519 minus.n62 gnd 0.199389f
C520 minus.n63 gnd 0.007201f
C521 minus.n64 gnd 0.031734f
C522 minus.n65 gnd 0.031734f
C523 minus.n66 gnd 0.031734f
C524 minus.n67 gnd 0.007201f
C525 minus.n68 gnd 0.199389f
C526 minus.n69 gnd 0.007201f
C527 minus.n70 gnd 0.031734f
C528 minus.n71 gnd 0.031734f
C529 minus.n72 gnd 0.031734f
C530 minus.n73 gnd 0.007201f
C531 minus.n74 gnd 0.199389f
C532 minus.n75 gnd 0.007201f
C533 minus.n76 gnd 0.031734f
C534 minus.n77 gnd 0.031734f
C535 minus.n78 gnd 0.031734f
C536 minus.n79 gnd 0.007201f
C537 minus.n80 gnd 0.199389f
C538 minus.n81 gnd 0.007201f
C539 minus.n82 gnd 0.199682f
C540 minus.n83 gnd 1.0631f
C541 minus.n84 gnd 1.584f
C542 minus.t1 gnd 0.009783f
C543 minus.t0 gnd 0.009783f
C544 minus.n85 gnd 0.032167f
C545 minus.t4 gnd 0.009783f
C546 minus.t3 gnd 0.009783f
C547 minus.n86 gnd 0.031726f
C548 minus.n87 gnd 0.27077f
C549 minus.t2 gnd 0.054448f
C550 minus.n88 gnd 0.147756f
C551 minus.n89 gnd 2.136f
C552 commonsourceibias.n0 gnd 0.012817f
C553 commonsourceibias.t151 gnd 0.194086f
C554 commonsourceibias.t83 gnd 0.17946f
C555 commonsourceibias.n1 gnd 0.009349f
C556 commonsourceibias.n2 gnd 0.009605f
C557 commonsourceibias.t161 gnd 0.17946f
C558 commonsourceibias.n3 gnd 0.012358f
C559 commonsourceibias.n4 gnd 0.009605f
C560 commonsourceibias.t152 gnd 0.17946f
C561 commonsourceibias.n5 gnd 0.071604f
C562 commonsourceibias.t171 gnd 0.17946f
C563 commonsourceibias.n6 gnd 0.009057f
C564 commonsourceibias.n7 gnd 0.009605f
C565 commonsourceibias.t145 gnd 0.17946f
C566 commonsourceibias.n8 gnd 0.012174f
C567 commonsourceibias.n9 gnd 0.009605f
C568 commonsourceibias.t124 gnd 0.17946f
C569 commonsourceibias.n10 gnd 0.071604f
C570 commonsourceibias.t158 gnd 0.17946f
C571 commonsourceibias.n11 gnd 0.008798f
C572 commonsourceibias.n12 gnd 0.009605f
C573 commonsourceibias.t148 gnd 0.17946f
C574 commonsourceibias.n13 gnd 0.01197f
C575 commonsourceibias.n14 gnd 0.012817f
C576 commonsourceibias.t16 gnd 0.194086f
C577 commonsourceibias.t60 gnd 0.17946f
C578 commonsourceibias.n15 gnd 0.009349f
C579 commonsourceibias.n16 gnd 0.009605f
C580 commonsourceibias.t4 gnd 0.17946f
C581 commonsourceibias.n17 gnd 0.012358f
C582 commonsourceibias.n18 gnd 0.009605f
C583 commonsourceibias.t14 gnd 0.17946f
C584 commonsourceibias.n19 gnd 0.071604f
C585 commonsourceibias.t74 gnd 0.17946f
C586 commonsourceibias.n20 gnd 0.009057f
C587 commonsourceibias.n21 gnd 0.009605f
C588 commonsourceibias.t20 gnd 0.17946f
C589 commonsourceibias.n22 gnd 0.012174f
C590 commonsourceibias.n23 gnd 0.009605f
C591 commonsourceibias.t34 gnd 0.17946f
C592 commonsourceibias.n24 gnd 0.071604f
C593 commonsourceibias.t10 gnd 0.17946f
C594 commonsourceibias.n25 gnd 0.008798f
C595 commonsourceibias.n26 gnd 0.009605f
C596 commonsourceibias.t18 gnd 0.17946f
C597 commonsourceibias.n27 gnd 0.01197f
C598 commonsourceibias.n28 gnd 0.009605f
C599 commonsourceibias.t54 gnd 0.17946f
C600 commonsourceibias.n29 gnd 0.071604f
C601 commonsourceibias.t30 gnd 0.17946f
C602 commonsourceibias.n30 gnd 0.008571f
C603 commonsourceibias.n31 gnd 0.009605f
C604 commonsourceibias.t36 gnd 0.17946f
C605 commonsourceibias.n32 gnd 0.011742f
C606 commonsourceibias.n33 gnd 0.009605f
C607 commonsourceibias.t70 gnd 0.17946f
C608 commonsourceibias.n34 gnd 0.071604f
C609 commonsourceibias.t22 gnd 0.17946f
C610 commonsourceibias.n35 gnd 0.008375f
C611 commonsourceibias.n36 gnd 0.009605f
C612 commonsourceibias.t62 gnd 0.17946f
C613 commonsourceibias.n37 gnd 0.011489f
C614 commonsourceibias.n38 gnd 0.009605f
C615 commonsourceibias.t0 gnd 0.17946f
C616 commonsourceibias.n39 gnd 0.071604f
C617 commonsourceibias.t42 gnd 0.17946f
C618 commonsourceibias.n40 gnd 0.008208f
C619 commonsourceibias.n41 gnd 0.009605f
C620 commonsourceibias.t52 gnd 0.17946f
C621 commonsourceibias.n42 gnd 0.011208f
C622 commonsourceibias.t26 gnd 0.199526f
C623 commonsourceibias.t58 gnd 0.17946f
C624 commonsourceibias.n43 gnd 0.078221f
C625 commonsourceibias.n44 gnd 0.085838f
C626 commonsourceibias.n45 gnd 0.03983f
C627 commonsourceibias.n46 gnd 0.009605f
C628 commonsourceibias.n47 gnd 0.009349f
C629 commonsourceibias.n48 gnd 0.013398f
C630 commonsourceibias.n49 gnd 0.071604f
C631 commonsourceibias.n50 gnd 0.013389f
C632 commonsourceibias.n51 gnd 0.009605f
C633 commonsourceibias.n52 gnd 0.009605f
C634 commonsourceibias.n53 gnd 0.009605f
C635 commonsourceibias.n54 gnd 0.012358f
C636 commonsourceibias.n55 gnd 0.071604f
C637 commonsourceibias.n56 gnd 0.012648f
C638 commonsourceibias.n57 gnd 0.012288f
C639 commonsourceibias.n58 gnd 0.009605f
C640 commonsourceibias.n59 gnd 0.009605f
C641 commonsourceibias.n60 gnd 0.009605f
C642 commonsourceibias.n61 gnd 0.009057f
C643 commonsourceibias.n62 gnd 0.01341f
C644 commonsourceibias.n63 gnd 0.071604f
C645 commonsourceibias.n64 gnd 0.013406f
C646 commonsourceibias.n65 gnd 0.009605f
C647 commonsourceibias.n66 gnd 0.009605f
C648 commonsourceibias.n67 gnd 0.009605f
C649 commonsourceibias.n68 gnd 0.012174f
C650 commonsourceibias.n69 gnd 0.071604f
C651 commonsourceibias.n70 gnd 0.012558f
C652 commonsourceibias.n71 gnd 0.012378f
C653 commonsourceibias.n72 gnd 0.009605f
C654 commonsourceibias.n73 gnd 0.009605f
C655 commonsourceibias.n74 gnd 0.009605f
C656 commonsourceibias.n75 gnd 0.008798f
C657 commonsourceibias.n76 gnd 0.013415f
C658 commonsourceibias.n77 gnd 0.071604f
C659 commonsourceibias.n78 gnd 0.013414f
C660 commonsourceibias.n79 gnd 0.009605f
C661 commonsourceibias.n80 gnd 0.009605f
C662 commonsourceibias.n81 gnd 0.009605f
C663 commonsourceibias.n82 gnd 0.01197f
C664 commonsourceibias.n83 gnd 0.071604f
C665 commonsourceibias.n84 gnd 0.012468f
C666 commonsourceibias.n85 gnd 0.012468f
C667 commonsourceibias.n86 gnd 0.009605f
C668 commonsourceibias.n87 gnd 0.009605f
C669 commonsourceibias.n88 gnd 0.009605f
C670 commonsourceibias.n89 gnd 0.008571f
C671 commonsourceibias.n90 gnd 0.013414f
C672 commonsourceibias.n91 gnd 0.071604f
C673 commonsourceibias.n92 gnd 0.013415f
C674 commonsourceibias.n93 gnd 0.009605f
C675 commonsourceibias.n94 gnd 0.009605f
C676 commonsourceibias.n95 gnd 0.009605f
C677 commonsourceibias.n96 gnd 0.011742f
C678 commonsourceibias.n97 gnd 0.071604f
C679 commonsourceibias.n98 gnd 0.012378f
C680 commonsourceibias.n99 gnd 0.012558f
C681 commonsourceibias.n100 gnd 0.009605f
C682 commonsourceibias.n101 gnd 0.009605f
C683 commonsourceibias.n102 gnd 0.009605f
C684 commonsourceibias.n103 gnd 0.008375f
C685 commonsourceibias.n104 gnd 0.013406f
C686 commonsourceibias.n105 gnd 0.071604f
C687 commonsourceibias.n106 gnd 0.01341f
C688 commonsourceibias.n107 gnd 0.009605f
C689 commonsourceibias.n108 gnd 0.009605f
C690 commonsourceibias.n109 gnd 0.009605f
C691 commonsourceibias.n110 gnd 0.011489f
C692 commonsourceibias.n111 gnd 0.071604f
C693 commonsourceibias.n112 gnd 0.012288f
C694 commonsourceibias.n113 gnd 0.012648f
C695 commonsourceibias.n114 gnd 0.009605f
C696 commonsourceibias.n115 gnd 0.009605f
C697 commonsourceibias.n116 gnd 0.009605f
C698 commonsourceibias.n117 gnd 0.008208f
C699 commonsourceibias.n118 gnd 0.013389f
C700 commonsourceibias.n119 gnd 0.071604f
C701 commonsourceibias.n120 gnd 0.013398f
C702 commonsourceibias.n121 gnd 0.009605f
C703 commonsourceibias.n122 gnd 0.009605f
C704 commonsourceibias.n123 gnd 0.009605f
C705 commonsourceibias.n124 gnd 0.011208f
C706 commonsourceibias.n125 gnd 0.071604f
C707 commonsourceibias.n126 gnd 0.011785f
C708 commonsourceibias.n127 gnd 0.085919f
C709 commonsourceibias.n128 gnd 0.095702f
C710 commonsourceibias.t17 gnd 0.020728f
C711 commonsourceibias.t61 gnd 0.020728f
C712 commonsourceibias.n129 gnd 0.183157f
C713 commonsourceibias.n130 gnd 0.158432f
C714 commonsourceibias.t5 gnd 0.020728f
C715 commonsourceibias.t15 gnd 0.020728f
C716 commonsourceibias.n131 gnd 0.183157f
C717 commonsourceibias.n132 gnd 0.084131f
C718 commonsourceibias.t75 gnd 0.020728f
C719 commonsourceibias.t21 gnd 0.020728f
C720 commonsourceibias.n133 gnd 0.183157f
C721 commonsourceibias.n134 gnd 0.084131f
C722 commonsourceibias.t35 gnd 0.020728f
C723 commonsourceibias.t11 gnd 0.020728f
C724 commonsourceibias.n135 gnd 0.183157f
C725 commonsourceibias.n136 gnd 0.084131f
C726 commonsourceibias.t19 gnd 0.020728f
C727 commonsourceibias.t55 gnd 0.020728f
C728 commonsourceibias.n137 gnd 0.183157f
C729 commonsourceibias.n138 gnd 0.070287f
C730 commonsourceibias.t59 gnd 0.020728f
C731 commonsourceibias.t27 gnd 0.020728f
C732 commonsourceibias.n139 gnd 0.18377f
C733 commonsourceibias.t43 gnd 0.020728f
C734 commonsourceibias.t53 gnd 0.020728f
C735 commonsourceibias.n140 gnd 0.183157f
C736 commonsourceibias.n141 gnd 0.170668f
C737 commonsourceibias.t63 gnd 0.020728f
C738 commonsourceibias.t1 gnd 0.020728f
C739 commonsourceibias.n142 gnd 0.183157f
C740 commonsourceibias.n143 gnd 0.084131f
C741 commonsourceibias.t71 gnd 0.020728f
C742 commonsourceibias.t23 gnd 0.020728f
C743 commonsourceibias.n144 gnd 0.183157f
C744 commonsourceibias.n145 gnd 0.084131f
C745 commonsourceibias.t31 gnd 0.020728f
C746 commonsourceibias.t37 gnd 0.020728f
C747 commonsourceibias.n146 gnd 0.183157f
C748 commonsourceibias.n147 gnd 0.070287f
C749 commonsourceibias.n148 gnd 0.085111f
C750 commonsourceibias.n149 gnd 0.062167f
C751 commonsourceibias.t93 gnd 0.17946f
C752 commonsourceibias.n150 gnd 0.071604f
C753 commonsourceibias.t131 gnd 0.17946f
C754 commonsourceibias.n151 gnd 0.071604f
C755 commonsourceibias.n152 gnd 0.009605f
C756 commonsourceibias.t117 gnd 0.17946f
C757 commonsourceibias.n153 gnd 0.071604f
C758 commonsourceibias.n154 gnd 0.009605f
C759 commonsourceibias.t176 gnd 0.17946f
C760 commonsourceibias.n155 gnd 0.071604f
C761 commonsourceibias.n156 gnd 0.009605f
C762 commonsourceibias.t144 gnd 0.17946f
C763 commonsourceibias.n157 gnd 0.008375f
C764 commonsourceibias.n158 gnd 0.009605f
C765 commonsourceibias.t190 gnd 0.17946f
C766 commonsourceibias.n159 gnd 0.011489f
C767 commonsourceibias.n160 gnd 0.009605f
C768 commonsourceibias.t164 gnd 0.17946f
C769 commonsourceibias.n161 gnd 0.071604f
C770 commonsourceibias.t111 gnd 0.17946f
C771 commonsourceibias.n162 gnd 0.008208f
C772 commonsourceibias.n163 gnd 0.009605f
C773 commonsourceibias.t100 gnd 0.17946f
C774 commonsourceibias.n164 gnd 0.011208f
C775 commonsourceibias.t140 gnd 0.199526f
C776 commonsourceibias.t84 gnd 0.17946f
C777 commonsourceibias.n165 gnd 0.078221f
C778 commonsourceibias.n166 gnd 0.085838f
C779 commonsourceibias.n167 gnd 0.03983f
C780 commonsourceibias.n168 gnd 0.009605f
C781 commonsourceibias.n169 gnd 0.009349f
C782 commonsourceibias.n170 gnd 0.013398f
C783 commonsourceibias.n171 gnd 0.071604f
C784 commonsourceibias.n172 gnd 0.013389f
C785 commonsourceibias.n173 gnd 0.009605f
C786 commonsourceibias.n174 gnd 0.009605f
C787 commonsourceibias.n175 gnd 0.009605f
C788 commonsourceibias.n176 gnd 0.012358f
C789 commonsourceibias.n177 gnd 0.071604f
C790 commonsourceibias.n178 gnd 0.012648f
C791 commonsourceibias.n179 gnd 0.012288f
C792 commonsourceibias.n180 gnd 0.009605f
C793 commonsourceibias.n181 gnd 0.009605f
C794 commonsourceibias.n182 gnd 0.009605f
C795 commonsourceibias.n183 gnd 0.009057f
C796 commonsourceibias.n184 gnd 0.01341f
C797 commonsourceibias.n185 gnd 0.071604f
C798 commonsourceibias.n186 gnd 0.013406f
C799 commonsourceibias.n187 gnd 0.009605f
C800 commonsourceibias.n188 gnd 0.009605f
C801 commonsourceibias.n189 gnd 0.009605f
C802 commonsourceibias.n190 gnd 0.012174f
C803 commonsourceibias.n191 gnd 0.071604f
C804 commonsourceibias.n192 gnd 0.012558f
C805 commonsourceibias.n193 gnd 0.012378f
C806 commonsourceibias.n194 gnd 0.009605f
C807 commonsourceibias.n195 gnd 0.009605f
C808 commonsourceibias.n196 gnd 0.011742f
C809 commonsourceibias.n197 gnd 0.008798f
C810 commonsourceibias.n198 gnd 0.013415f
C811 commonsourceibias.n199 gnd 0.009605f
C812 commonsourceibias.n200 gnd 0.009605f
C813 commonsourceibias.n201 gnd 0.013414f
C814 commonsourceibias.n202 gnd 0.008571f
C815 commonsourceibias.n203 gnd 0.01197f
C816 commonsourceibias.n204 gnd 0.009605f
C817 commonsourceibias.n205 gnd 0.008391f
C818 commonsourceibias.n206 gnd 0.012468f
C819 commonsourceibias.n207 gnd 0.012468f
C820 commonsourceibias.n208 gnd 0.008391f
C821 commonsourceibias.n209 gnd 0.009605f
C822 commonsourceibias.n210 gnd 0.009605f
C823 commonsourceibias.n211 gnd 0.008571f
C824 commonsourceibias.n212 gnd 0.013414f
C825 commonsourceibias.n213 gnd 0.071604f
C826 commonsourceibias.n214 gnd 0.013415f
C827 commonsourceibias.n215 gnd 0.009605f
C828 commonsourceibias.n216 gnd 0.009605f
C829 commonsourceibias.n217 gnd 0.009605f
C830 commonsourceibias.n218 gnd 0.011742f
C831 commonsourceibias.n219 gnd 0.071604f
C832 commonsourceibias.n220 gnd 0.012378f
C833 commonsourceibias.n221 gnd 0.012558f
C834 commonsourceibias.n222 gnd 0.009605f
C835 commonsourceibias.n223 gnd 0.009605f
C836 commonsourceibias.n224 gnd 0.009605f
C837 commonsourceibias.n225 gnd 0.008375f
C838 commonsourceibias.n226 gnd 0.013406f
C839 commonsourceibias.n227 gnd 0.071604f
C840 commonsourceibias.n228 gnd 0.01341f
C841 commonsourceibias.n229 gnd 0.009605f
C842 commonsourceibias.n230 gnd 0.009605f
C843 commonsourceibias.n231 gnd 0.009605f
C844 commonsourceibias.n232 gnd 0.011489f
C845 commonsourceibias.n233 gnd 0.071604f
C846 commonsourceibias.n234 gnd 0.012288f
C847 commonsourceibias.n235 gnd 0.012648f
C848 commonsourceibias.n236 gnd 0.009605f
C849 commonsourceibias.n237 gnd 0.009605f
C850 commonsourceibias.n238 gnd 0.009605f
C851 commonsourceibias.n239 gnd 0.008208f
C852 commonsourceibias.n240 gnd 0.013389f
C853 commonsourceibias.n241 gnd 0.071604f
C854 commonsourceibias.n242 gnd 0.013398f
C855 commonsourceibias.n243 gnd 0.009605f
C856 commonsourceibias.n244 gnd 0.009605f
C857 commonsourceibias.n245 gnd 0.009605f
C858 commonsourceibias.n246 gnd 0.011208f
C859 commonsourceibias.n247 gnd 0.071604f
C860 commonsourceibias.n248 gnd 0.011785f
C861 commonsourceibias.n249 gnd 0.085919f
C862 commonsourceibias.n250 gnd 0.056156f
C863 commonsourceibias.n251 gnd 0.012817f
C864 commonsourceibias.t88 gnd 0.194086f
C865 commonsourceibias.t198 gnd 0.17946f
C866 commonsourceibias.n252 gnd 0.009349f
C867 commonsourceibias.n253 gnd 0.009605f
C868 commonsourceibias.t186 gnd 0.17946f
C869 commonsourceibias.n254 gnd 0.012358f
C870 commonsourceibias.n255 gnd 0.009605f
C871 commonsourceibias.t95 gnd 0.17946f
C872 commonsourceibias.n256 gnd 0.071604f
C873 commonsourceibias.t196 gnd 0.17946f
C874 commonsourceibias.n257 gnd 0.009057f
C875 commonsourceibias.n258 gnd 0.009605f
C876 commonsourceibias.t105 gnd 0.17946f
C877 commonsourceibias.n259 gnd 0.012174f
C878 commonsourceibias.n260 gnd 0.009605f
C879 commonsourceibias.t94 gnd 0.17946f
C880 commonsourceibias.n261 gnd 0.071604f
C881 commonsourceibias.t197 gnd 0.17946f
C882 commonsourceibias.n262 gnd 0.008798f
C883 commonsourceibias.n263 gnd 0.009605f
C884 commonsourceibias.t115 gnd 0.17946f
C885 commonsourceibias.n264 gnd 0.01197f
C886 commonsourceibias.n265 gnd 0.009605f
C887 commonsourceibias.t141 gnd 0.17946f
C888 commonsourceibias.n266 gnd 0.071604f
C889 commonsourceibias.t195 gnd 0.17946f
C890 commonsourceibias.n267 gnd 0.008571f
C891 commonsourceibias.n268 gnd 0.009605f
C892 commonsourceibias.t113 gnd 0.17946f
C893 commonsourceibias.n269 gnd 0.011742f
C894 commonsourceibias.n270 gnd 0.009605f
C895 commonsourceibias.t138 gnd 0.17946f
C896 commonsourceibias.n271 gnd 0.071604f
C897 commonsourceibias.t130 gnd 0.17946f
C898 commonsourceibias.n272 gnd 0.008375f
C899 commonsourceibias.n273 gnd 0.009605f
C900 commonsourceibias.t114 gnd 0.17946f
C901 commonsourceibias.n274 gnd 0.011489f
C902 commonsourceibias.n275 gnd 0.009605f
C903 commonsourceibias.t139 gnd 0.17946f
C904 commonsourceibias.n276 gnd 0.071604f
C905 commonsourceibias.t129 gnd 0.17946f
C906 commonsourceibias.n277 gnd 0.008208f
C907 commonsourceibias.n278 gnd 0.009605f
C908 commonsourceibias.t125 gnd 0.17946f
C909 commonsourceibias.n279 gnd 0.011208f
C910 commonsourceibias.t134 gnd 0.199526f
C911 commonsourceibias.t147 gnd 0.17946f
C912 commonsourceibias.n280 gnd 0.078221f
C913 commonsourceibias.n281 gnd 0.085838f
C914 commonsourceibias.n282 gnd 0.03983f
C915 commonsourceibias.n283 gnd 0.009605f
C916 commonsourceibias.n284 gnd 0.009349f
C917 commonsourceibias.n285 gnd 0.013398f
C918 commonsourceibias.n286 gnd 0.071604f
C919 commonsourceibias.n287 gnd 0.013389f
C920 commonsourceibias.n288 gnd 0.009605f
C921 commonsourceibias.n289 gnd 0.009605f
C922 commonsourceibias.n290 gnd 0.009605f
C923 commonsourceibias.n291 gnd 0.012358f
C924 commonsourceibias.n292 gnd 0.071604f
C925 commonsourceibias.n293 gnd 0.012648f
C926 commonsourceibias.n294 gnd 0.012288f
C927 commonsourceibias.n295 gnd 0.009605f
C928 commonsourceibias.n296 gnd 0.009605f
C929 commonsourceibias.n297 gnd 0.009605f
C930 commonsourceibias.n298 gnd 0.009057f
C931 commonsourceibias.n299 gnd 0.01341f
C932 commonsourceibias.n300 gnd 0.071604f
C933 commonsourceibias.n301 gnd 0.013406f
C934 commonsourceibias.n302 gnd 0.009605f
C935 commonsourceibias.n303 gnd 0.009605f
C936 commonsourceibias.n304 gnd 0.009605f
C937 commonsourceibias.n305 gnd 0.012174f
C938 commonsourceibias.n306 gnd 0.071604f
C939 commonsourceibias.n307 gnd 0.012558f
C940 commonsourceibias.n308 gnd 0.012378f
C941 commonsourceibias.n309 gnd 0.009605f
C942 commonsourceibias.n310 gnd 0.009605f
C943 commonsourceibias.n311 gnd 0.009605f
C944 commonsourceibias.n312 gnd 0.008798f
C945 commonsourceibias.n313 gnd 0.013415f
C946 commonsourceibias.n314 gnd 0.071604f
C947 commonsourceibias.n315 gnd 0.013414f
C948 commonsourceibias.n316 gnd 0.009605f
C949 commonsourceibias.n317 gnd 0.009605f
C950 commonsourceibias.n318 gnd 0.009605f
C951 commonsourceibias.n319 gnd 0.01197f
C952 commonsourceibias.n320 gnd 0.071604f
C953 commonsourceibias.n321 gnd 0.012468f
C954 commonsourceibias.n322 gnd 0.012468f
C955 commonsourceibias.n323 gnd 0.009605f
C956 commonsourceibias.n324 gnd 0.009605f
C957 commonsourceibias.n325 gnd 0.009605f
C958 commonsourceibias.n326 gnd 0.008571f
C959 commonsourceibias.n327 gnd 0.013414f
C960 commonsourceibias.n328 gnd 0.071604f
C961 commonsourceibias.n329 gnd 0.013415f
C962 commonsourceibias.n330 gnd 0.009605f
C963 commonsourceibias.n331 gnd 0.009605f
C964 commonsourceibias.n332 gnd 0.009605f
C965 commonsourceibias.n333 gnd 0.011742f
C966 commonsourceibias.n334 gnd 0.071604f
C967 commonsourceibias.n335 gnd 0.012378f
C968 commonsourceibias.n336 gnd 0.012558f
C969 commonsourceibias.n337 gnd 0.009605f
C970 commonsourceibias.n338 gnd 0.009605f
C971 commonsourceibias.n339 gnd 0.009605f
C972 commonsourceibias.n340 gnd 0.008375f
C973 commonsourceibias.n341 gnd 0.013406f
C974 commonsourceibias.n342 gnd 0.071604f
C975 commonsourceibias.n343 gnd 0.01341f
C976 commonsourceibias.n344 gnd 0.009605f
C977 commonsourceibias.n345 gnd 0.009605f
C978 commonsourceibias.n346 gnd 0.009605f
C979 commonsourceibias.n347 gnd 0.011489f
C980 commonsourceibias.n348 gnd 0.071604f
C981 commonsourceibias.n349 gnd 0.012288f
C982 commonsourceibias.n350 gnd 0.012648f
C983 commonsourceibias.n351 gnd 0.009605f
C984 commonsourceibias.n352 gnd 0.009605f
C985 commonsourceibias.n353 gnd 0.009605f
C986 commonsourceibias.n354 gnd 0.008208f
C987 commonsourceibias.n355 gnd 0.013389f
C988 commonsourceibias.n356 gnd 0.071604f
C989 commonsourceibias.n357 gnd 0.013398f
C990 commonsourceibias.n358 gnd 0.009605f
C991 commonsourceibias.n359 gnd 0.009605f
C992 commonsourceibias.n360 gnd 0.009605f
C993 commonsourceibias.n361 gnd 0.011208f
C994 commonsourceibias.n362 gnd 0.071604f
C995 commonsourceibias.n363 gnd 0.011785f
C996 commonsourceibias.n364 gnd 0.085919f
C997 commonsourceibias.n365 gnd 0.029883f
C998 commonsourceibias.n366 gnd 0.153509f
C999 commonsourceibias.n367 gnd 0.012817f
C1000 commonsourceibias.t92 gnd 0.17946f
C1001 commonsourceibias.n368 gnd 0.009349f
C1002 commonsourceibias.n369 gnd 0.009605f
C1003 commonsourceibias.t163 gnd 0.17946f
C1004 commonsourceibias.n370 gnd 0.012358f
C1005 commonsourceibias.n371 gnd 0.009605f
C1006 commonsourceibias.t157 gnd 0.17946f
C1007 commonsourceibias.n372 gnd 0.071604f
C1008 commonsourceibias.t194 gnd 0.17946f
C1009 commonsourceibias.n373 gnd 0.009057f
C1010 commonsourceibias.n374 gnd 0.009605f
C1011 commonsourceibias.t110 gnd 0.17946f
C1012 commonsourceibias.n375 gnd 0.012174f
C1013 commonsourceibias.n376 gnd 0.009605f
C1014 commonsourceibias.t149 gnd 0.17946f
C1015 commonsourceibias.n377 gnd 0.071604f
C1016 commonsourceibias.t182 gnd 0.17946f
C1017 commonsourceibias.n378 gnd 0.008798f
C1018 commonsourceibias.n379 gnd 0.009605f
C1019 commonsourceibias.t173 gnd 0.17946f
C1020 commonsourceibias.n380 gnd 0.01197f
C1021 commonsourceibias.n381 gnd 0.009605f
C1022 commonsourceibias.t80 gnd 0.17946f
C1023 commonsourceibias.n382 gnd 0.071604f
C1024 commonsourceibias.t172 gnd 0.17946f
C1025 commonsourceibias.n383 gnd 0.008571f
C1026 commonsourceibias.n384 gnd 0.009605f
C1027 commonsourceibias.t168 gnd 0.17946f
C1028 commonsourceibias.n385 gnd 0.011742f
C1029 commonsourceibias.n386 gnd 0.009605f
C1030 commonsourceibias.t187 gnd 0.17946f
C1031 commonsourceibias.n387 gnd 0.071604f
C1032 commonsourceibias.t96 gnd 0.17946f
C1033 commonsourceibias.n388 gnd 0.008375f
C1034 commonsourceibias.n389 gnd 0.009605f
C1035 commonsourceibias.t165 gnd 0.17946f
C1036 commonsourceibias.n390 gnd 0.011489f
C1037 commonsourceibias.n391 gnd 0.009605f
C1038 commonsourceibias.t175 gnd 0.17946f
C1039 commonsourceibias.n392 gnd 0.071604f
C1040 commonsourceibias.t199 gnd 0.17946f
C1041 commonsourceibias.n393 gnd 0.008208f
C1042 commonsourceibias.n394 gnd 0.009605f
C1043 commonsourceibias.t155 gnd 0.17946f
C1044 commonsourceibias.n395 gnd 0.011208f
C1045 commonsourceibias.t184 gnd 0.199526f
C1046 commonsourceibias.t150 gnd 0.17946f
C1047 commonsourceibias.n396 gnd 0.078221f
C1048 commonsourceibias.n397 gnd 0.085838f
C1049 commonsourceibias.n398 gnd 0.03983f
C1050 commonsourceibias.n399 gnd 0.009605f
C1051 commonsourceibias.n400 gnd 0.009349f
C1052 commonsourceibias.n401 gnd 0.013398f
C1053 commonsourceibias.n402 gnd 0.071604f
C1054 commonsourceibias.n403 gnd 0.013389f
C1055 commonsourceibias.n404 gnd 0.009605f
C1056 commonsourceibias.n405 gnd 0.009605f
C1057 commonsourceibias.n406 gnd 0.009605f
C1058 commonsourceibias.n407 gnd 0.012358f
C1059 commonsourceibias.n408 gnd 0.071604f
C1060 commonsourceibias.n409 gnd 0.012648f
C1061 commonsourceibias.n410 gnd 0.012288f
C1062 commonsourceibias.n411 gnd 0.009605f
C1063 commonsourceibias.n412 gnd 0.009605f
C1064 commonsourceibias.n413 gnd 0.009605f
C1065 commonsourceibias.n414 gnd 0.009057f
C1066 commonsourceibias.n415 gnd 0.01341f
C1067 commonsourceibias.n416 gnd 0.071604f
C1068 commonsourceibias.n417 gnd 0.013406f
C1069 commonsourceibias.n418 gnd 0.009605f
C1070 commonsourceibias.n419 gnd 0.009605f
C1071 commonsourceibias.n420 gnd 0.009605f
C1072 commonsourceibias.n421 gnd 0.012174f
C1073 commonsourceibias.n422 gnd 0.071604f
C1074 commonsourceibias.n423 gnd 0.012558f
C1075 commonsourceibias.n424 gnd 0.012378f
C1076 commonsourceibias.n425 gnd 0.009605f
C1077 commonsourceibias.n426 gnd 0.009605f
C1078 commonsourceibias.n427 gnd 0.009605f
C1079 commonsourceibias.n428 gnd 0.008798f
C1080 commonsourceibias.n429 gnd 0.013415f
C1081 commonsourceibias.n430 gnd 0.071604f
C1082 commonsourceibias.n431 gnd 0.013414f
C1083 commonsourceibias.n432 gnd 0.009605f
C1084 commonsourceibias.n433 gnd 0.009605f
C1085 commonsourceibias.n434 gnd 0.009605f
C1086 commonsourceibias.n435 gnd 0.01197f
C1087 commonsourceibias.n436 gnd 0.071604f
C1088 commonsourceibias.n437 gnd 0.012468f
C1089 commonsourceibias.n438 gnd 0.012468f
C1090 commonsourceibias.n439 gnd 0.009605f
C1091 commonsourceibias.n440 gnd 0.009605f
C1092 commonsourceibias.n441 gnd 0.009605f
C1093 commonsourceibias.n442 gnd 0.008571f
C1094 commonsourceibias.n443 gnd 0.013414f
C1095 commonsourceibias.n444 gnd 0.071604f
C1096 commonsourceibias.n445 gnd 0.013415f
C1097 commonsourceibias.n446 gnd 0.009605f
C1098 commonsourceibias.n447 gnd 0.009605f
C1099 commonsourceibias.n448 gnd 0.009605f
C1100 commonsourceibias.n449 gnd 0.011742f
C1101 commonsourceibias.n450 gnd 0.071604f
C1102 commonsourceibias.n451 gnd 0.012378f
C1103 commonsourceibias.n452 gnd 0.012558f
C1104 commonsourceibias.n453 gnd 0.009605f
C1105 commonsourceibias.n454 gnd 0.009605f
C1106 commonsourceibias.n455 gnd 0.009605f
C1107 commonsourceibias.n456 gnd 0.008375f
C1108 commonsourceibias.n457 gnd 0.013406f
C1109 commonsourceibias.n458 gnd 0.071604f
C1110 commonsourceibias.n459 gnd 0.01341f
C1111 commonsourceibias.n460 gnd 0.009605f
C1112 commonsourceibias.n461 gnd 0.009605f
C1113 commonsourceibias.n462 gnd 0.009605f
C1114 commonsourceibias.n463 gnd 0.011489f
C1115 commonsourceibias.n464 gnd 0.071604f
C1116 commonsourceibias.n465 gnd 0.012288f
C1117 commonsourceibias.n466 gnd 0.012648f
C1118 commonsourceibias.n467 gnd 0.009605f
C1119 commonsourceibias.n468 gnd 0.009605f
C1120 commonsourceibias.n469 gnd 0.009605f
C1121 commonsourceibias.n470 gnd 0.008208f
C1122 commonsourceibias.n471 gnd 0.013389f
C1123 commonsourceibias.n472 gnd 0.071604f
C1124 commonsourceibias.n473 gnd 0.013398f
C1125 commonsourceibias.n474 gnd 0.009605f
C1126 commonsourceibias.n475 gnd 0.009605f
C1127 commonsourceibias.n476 gnd 0.009605f
C1128 commonsourceibias.n477 gnd 0.011208f
C1129 commonsourceibias.n478 gnd 0.071604f
C1130 commonsourceibias.n479 gnd 0.011785f
C1131 commonsourceibias.t183 gnd 0.194086f
C1132 commonsourceibias.n480 gnd 0.085919f
C1133 commonsourceibias.n481 gnd 0.029883f
C1134 commonsourceibias.n482 gnd 0.456424f
C1135 commonsourceibias.n483 gnd 0.012817f
C1136 commonsourceibias.t112 gnd 0.194086f
C1137 commonsourceibias.t169 gnd 0.17946f
C1138 commonsourceibias.n484 gnd 0.009349f
C1139 commonsourceibias.n485 gnd 0.009605f
C1140 commonsourceibias.t142 gnd 0.17946f
C1141 commonsourceibias.n486 gnd 0.012358f
C1142 commonsourceibias.n487 gnd 0.009605f
C1143 commonsourceibias.t154 gnd 0.17946f
C1144 commonsourceibias.n488 gnd 0.009057f
C1145 commonsourceibias.n489 gnd 0.009605f
C1146 commonsourceibias.t108 gnd 0.17946f
C1147 commonsourceibias.n490 gnd 0.012174f
C1148 commonsourceibias.n491 gnd 0.009605f
C1149 commonsourceibias.t128 gnd 0.17946f
C1150 commonsourceibias.n492 gnd 0.008798f
C1151 commonsourceibias.n493 gnd 0.009605f
C1152 commonsourceibias.t109 gnd 0.17946f
C1153 commonsourceibias.n494 gnd 0.01197f
C1154 commonsourceibias.t69 gnd 0.020728f
C1155 commonsourceibias.t9 gnd 0.020728f
C1156 commonsourceibias.n495 gnd 0.18377f
C1157 commonsourceibias.t7 gnd 0.020728f
C1158 commonsourceibias.t67 gnd 0.020728f
C1159 commonsourceibias.n496 gnd 0.183157f
C1160 commonsourceibias.n497 gnd 0.170668f
C1161 commonsourceibias.t29 gnd 0.020728f
C1162 commonsourceibias.t79 gnd 0.020728f
C1163 commonsourceibias.n498 gnd 0.183157f
C1164 commonsourceibias.n499 gnd 0.084131f
C1165 commonsourceibias.t49 gnd 0.020728f
C1166 commonsourceibias.t3 gnd 0.020728f
C1167 commonsourceibias.n500 gnd 0.183157f
C1168 commonsourceibias.n501 gnd 0.084131f
C1169 commonsourceibias.t65 gnd 0.020728f
C1170 commonsourceibias.t51 gnd 0.020728f
C1171 commonsourceibias.n502 gnd 0.183157f
C1172 commonsourceibias.n503 gnd 0.070287f
C1173 commonsourceibias.n504 gnd 0.012817f
C1174 commonsourceibias.t76 gnd 0.17946f
C1175 commonsourceibias.n505 gnd 0.009349f
C1176 commonsourceibias.n506 gnd 0.009605f
C1177 commonsourceibias.t24 gnd 0.17946f
C1178 commonsourceibias.n507 gnd 0.012358f
C1179 commonsourceibias.n508 gnd 0.009605f
C1180 commonsourceibias.t12 gnd 0.17946f
C1181 commonsourceibias.n509 gnd 0.009057f
C1182 commonsourceibias.n510 gnd 0.009605f
C1183 commonsourceibias.t46 gnd 0.17946f
C1184 commonsourceibias.n511 gnd 0.012174f
C1185 commonsourceibias.n512 gnd 0.009605f
C1186 commonsourceibias.t32 gnd 0.17946f
C1187 commonsourceibias.n513 gnd 0.008798f
C1188 commonsourceibias.n514 gnd 0.009605f
C1189 commonsourceibias.t44 gnd 0.17946f
C1190 commonsourceibias.n515 gnd 0.01197f
C1191 commonsourceibias.n516 gnd 0.009605f
C1192 commonsourceibias.t50 gnd 0.17946f
C1193 commonsourceibias.n517 gnd 0.008571f
C1194 commonsourceibias.n518 gnd 0.009605f
C1195 commonsourceibias.t64 gnd 0.17946f
C1196 commonsourceibias.n519 gnd 0.011742f
C1197 commonsourceibias.n520 gnd 0.009605f
C1198 commonsourceibias.t48 gnd 0.17946f
C1199 commonsourceibias.n521 gnd 0.008375f
C1200 commonsourceibias.n522 gnd 0.009605f
C1201 commonsourceibias.t78 gnd 0.17946f
C1202 commonsourceibias.n523 gnd 0.011489f
C1203 commonsourceibias.n524 gnd 0.009605f
C1204 commonsourceibias.t66 gnd 0.17946f
C1205 commonsourceibias.n525 gnd 0.008208f
C1206 commonsourceibias.n526 gnd 0.009605f
C1207 commonsourceibias.t6 gnd 0.17946f
C1208 commonsourceibias.n527 gnd 0.011208f
C1209 commonsourceibias.t68 gnd 0.199526f
C1210 commonsourceibias.t8 gnd 0.17946f
C1211 commonsourceibias.n528 gnd 0.078221f
C1212 commonsourceibias.n529 gnd 0.085838f
C1213 commonsourceibias.n530 gnd 0.03983f
C1214 commonsourceibias.n531 gnd 0.009605f
C1215 commonsourceibias.n532 gnd 0.009349f
C1216 commonsourceibias.n533 gnd 0.013398f
C1217 commonsourceibias.n534 gnd 0.071604f
C1218 commonsourceibias.n535 gnd 0.013389f
C1219 commonsourceibias.n536 gnd 0.009605f
C1220 commonsourceibias.n537 gnd 0.009605f
C1221 commonsourceibias.n538 gnd 0.009605f
C1222 commonsourceibias.n539 gnd 0.012358f
C1223 commonsourceibias.n540 gnd 0.071604f
C1224 commonsourceibias.n541 gnd 0.012648f
C1225 commonsourceibias.t28 gnd 0.17946f
C1226 commonsourceibias.n542 gnd 0.071604f
C1227 commonsourceibias.n543 gnd 0.012288f
C1228 commonsourceibias.n544 gnd 0.009605f
C1229 commonsourceibias.n545 gnd 0.009605f
C1230 commonsourceibias.n546 gnd 0.009605f
C1231 commonsourceibias.n547 gnd 0.009057f
C1232 commonsourceibias.n548 gnd 0.01341f
C1233 commonsourceibias.n549 gnd 0.071604f
C1234 commonsourceibias.n550 gnd 0.013406f
C1235 commonsourceibias.n551 gnd 0.009605f
C1236 commonsourceibias.n552 gnd 0.009605f
C1237 commonsourceibias.n553 gnd 0.009605f
C1238 commonsourceibias.n554 gnd 0.012174f
C1239 commonsourceibias.n555 gnd 0.071604f
C1240 commonsourceibias.n556 gnd 0.012558f
C1241 commonsourceibias.t2 gnd 0.17946f
C1242 commonsourceibias.n557 gnd 0.071604f
C1243 commonsourceibias.n558 gnd 0.012378f
C1244 commonsourceibias.n559 gnd 0.009605f
C1245 commonsourceibias.n560 gnd 0.009605f
C1246 commonsourceibias.n561 gnd 0.009605f
C1247 commonsourceibias.n562 gnd 0.008798f
C1248 commonsourceibias.n563 gnd 0.013415f
C1249 commonsourceibias.n564 gnd 0.071604f
C1250 commonsourceibias.n565 gnd 0.013414f
C1251 commonsourceibias.n566 gnd 0.009605f
C1252 commonsourceibias.n567 gnd 0.009605f
C1253 commonsourceibias.n568 gnd 0.009605f
C1254 commonsourceibias.n569 gnd 0.01197f
C1255 commonsourceibias.n570 gnd 0.071604f
C1256 commonsourceibias.n571 gnd 0.012468f
C1257 commonsourceibias.t72 gnd 0.17946f
C1258 commonsourceibias.n572 gnd 0.071604f
C1259 commonsourceibias.n573 gnd 0.012468f
C1260 commonsourceibias.n574 gnd 0.009605f
C1261 commonsourceibias.n575 gnd 0.009605f
C1262 commonsourceibias.n576 gnd 0.009605f
C1263 commonsourceibias.n577 gnd 0.008571f
C1264 commonsourceibias.n578 gnd 0.013414f
C1265 commonsourceibias.n579 gnd 0.071604f
C1266 commonsourceibias.n580 gnd 0.013415f
C1267 commonsourceibias.n581 gnd 0.009605f
C1268 commonsourceibias.n582 gnd 0.009605f
C1269 commonsourceibias.n583 gnd 0.009605f
C1270 commonsourceibias.n584 gnd 0.011742f
C1271 commonsourceibias.n585 gnd 0.071604f
C1272 commonsourceibias.n586 gnd 0.012378f
C1273 commonsourceibias.t56 gnd 0.17946f
C1274 commonsourceibias.n587 gnd 0.071604f
C1275 commonsourceibias.n588 gnd 0.012558f
C1276 commonsourceibias.n589 gnd 0.009605f
C1277 commonsourceibias.n590 gnd 0.009605f
C1278 commonsourceibias.n591 gnd 0.009605f
C1279 commonsourceibias.n592 gnd 0.008375f
C1280 commonsourceibias.n593 gnd 0.013406f
C1281 commonsourceibias.n594 gnd 0.071604f
C1282 commonsourceibias.n595 gnd 0.01341f
C1283 commonsourceibias.n596 gnd 0.009605f
C1284 commonsourceibias.n597 gnd 0.009605f
C1285 commonsourceibias.n598 gnd 0.009605f
C1286 commonsourceibias.n599 gnd 0.011489f
C1287 commonsourceibias.n600 gnd 0.071604f
C1288 commonsourceibias.n601 gnd 0.012288f
C1289 commonsourceibias.t38 gnd 0.17946f
C1290 commonsourceibias.n602 gnd 0.071604f
C1291 commonsourceibias.n603 gnd 0.012648f
C1292 commonsourceibias.n604 gnd 0.009605f
C1293 commonsourceibias.n605 gnd 0.009605f
C1294 commonsourceibias.n606 gnd 0.009605f
C1295 commonsourceibias.n607 gnd 0.008208f
C1296 commonsourceibias.n608 gnd 0.013389f
C1297 commonsourceibias.n609 gnd 0.071604f
C1298 commonsourceibias.n610 gnd 0.013398f
C1299 commonsourceibias.n611 gnd 0.009605f
C1300 commonsourceibias.n612 gnd 0.009605f
C1301 commonsourceibias.n613 gnd 0.009605f
C1302 commonsourceibias.n614 gnd 0.011208f
C1303 commonsourceibias.n615 gnd 0.071604f
C1304 commonsourceibias.n616 gnd 0.011785f
C1305 commonsourceibias.t40 gnd 0.194086f
C1306 commonsourceibias.n617 gnd 0.085919f
C1307 commonsourceibias.n618 gnd 0.095702f
C1308 commonsourceibias.t77 gnd 0.020728f
C1309 commonsourceibias.t41 gnd 0.020728f
C1310 commonsourceibias.n619 gnd 0.183157f
C1311 commonsourceibias.n620 gnd 0.158432f
C1312 commonsourceibias.t39 gnd 0.020728f
C1313 commonsourceibias.t25 gnd 0.020728f
C1314 commonsourceibias.n621 gnd 0.183157f
C1315 commonsourceibias.n622 gnd 0.084131f
C1316 commonsourceibias.t47 gnd 0.020728f
C1317 commonsourceibias.t13 gnd 0.020728f
C1318 commonsourceibias.n623 gnd 0.183157f
C1319 commonsourceibias.n624 gnd 0.084131f
C1320 commonsourceibias.t33 gnd 0.020728f
C1321 commonsourceibias.t57 gnd 0.020728f
C1322 commonsourceibias.n625 gnd 0.183157f
C1323 commonsourceibias.n626 gnd 0.084131f
C1324 commonsourceibias.t73 gnd 0.020728f
C1325 commonsourceibias.t45 gnd 0.020728f
C1326 commonsourceibias.n627 gnd 0.183157f
C1327 commonsourceibias.n628 gnd 0.070287f
C1328 commonsourceibias.n629 gnd 0.085111f
C1329 commonsourceibias.n630 gnd 0.062167f
C1330 commonsourceibias.t102 gnd 0.17946f
C1331 commonsourceibias.n631 gnd 0.071604f
C1332 commonsourceibias.n632 gnd 0.009605f
C1333 commonsourceibias.t188 gnd 0.17946f
C1334 commonsourceibias.n633 gnd 0.071604f
C1335 commonsourceibias.n634 gnd 0.009605f
C1336 commonsourceibias.t162 gnd 0.17946f
C1337 commonsourceibias.n635 gnd 0.071604f
C1338 commonsourceibias.n636 gnd 0.009605f
C1339 commonsourceibias.t103 gnd 0.17946f
C1340 commonsourceibias.n637 gnd 0.008375f
C1341 commonsourceibias.n638 gnd 0.009605f
C1342 commonsourceibias.t166 gnd 0.17946f
C1343 commonsourceibias.n639 gnd 0.011489f
C1344 commonsourceibias.n640 gnd 0.009605f
C1345 commonsourceibias.t185 gnd 0.17946f
C1346 commonsourceibias.n641 gnd 0.008208f
C1347 commonsourceibias.n642 gnd 0.009605f
C1348 commonsourceibias.t160 gnd 0.17946f
C1349 commonsourceibias.n643 gnd 0.011208f
C1350 commonsourceibias.t177 gnd 0.199526f
C1351 commonsourceibias.t159 gnd 0.17946f
C1352 commonsourceibias.n644 gnd 0.078221f
C1353 commonsourceibias.n645 gnd 0.085838f
C1354 commonsourceibias.n646 gnd 0.03983f
C1355 commonsourceibias.n647 gnd 0.009605f
C1356 commonsourceibias.n648 gnd 0.009349f
C1357 commonsourceibias.n649 gnd 0.013398f
C1358 commonsourceibias.n650 gnd 0.071604f
C1359 commonsourceibias.n651 gnd 0.013389f
C1360 commonsourceibias.n652 gnd 0.009605f
C1361 commonsourceibias.n653 gnd 0.009605f
C1362 commonsourceibias.n654 gnd 0.009605f
C1363 commonsourceibias.n655 gnd 0.012358f
C1364 commonsourceibias.n656 gnd 0.071604f
C1365 commonsourceibias.n657 gnd 0.012648f
C1366 commonsourceibias.t135 gnd 0.17946f
C1367 commonsourceibias.n658 gnd 0.071604f
C1368 commonsourceibias.n659 gnd 0.012288f
C1369 commonsourceibias.n660 gnd 0.009605f
C1370 commonsourceibias.n661 gnd 0.009605f
C1371 commonsourceibias.n662 gnd 0.009605f
C1372 commonsourceibias.n663 gnd 0.009057f
C1373 commonsourceibias.n664 gnd 0.01341f
C1374 commonsourceibias.n665 gnd 0.071604f
C1375 commonsourceibias.n666 gnd 0.013406f
C1376 commonsourceibias.n667 gnd 0.009605f
C1377 commonsourceibias.n668 gnd 0.009605f
C1378 commonsourceibias.n669 gnd 0.009605f
C1379 commonsourceibias.n670 gnd 0.012174f
C1380 commonsourceibias.n671 gnd 0.071604f
C1381 commonsourceibias.n672 gnd 0.012558f
C1382 commonsourceibias.n673 gnd 0.012378f
C1383 commonsourceibias.n674 gnd 0.009605f
C1384 commonsourceibias.n675 gnd 0.009605f
C1385 commonsourceibias.n676 gnd 0.011742f
C1386 commonsourceibias.n677 gnd 0.008798f
C1387 commonsourceibias.n678 gnd 0.013415f
C1388 commonsourceibias.n679 gnd 0.009605f
C1389 commonsourceibias.n680 gnd 0.009605f
C1390 commonsourceibias.n681 gnd 0.013414f
C1391 commonsourceibias.n682 gnd 0.008571f
C1392 commonsourceibias.n683 gnd 0.01197f
C1393 commonsourceibias.n684 gnd 0.009605f
C1394 commonsourceibias.n685 gnd 0.008391f
C1395 commonsourceibias.n686 gnd 0.012468f
C1396 commonsourceibias.t174 gnd 0.17946f
C1397 commonsourceibias.n687 gnd 0.071604f
C1398 commonsourceibias.n688 gnd 0.012468f
C1399 commonsourceibias.n689 gnd 0.008391f
C1400 commonsourceibias.n690 gnd 0.009605f
C1401 commonsourceibias.n691 gnd 0.009605f
C1402 commonsourceibias.n692 gnd 0.008571f
C1403 commonsourceibias.n693 gnd 0.013414f
C1404 commonsourceibias.n694 gnd 0.071604f
C1405 commonsourceibias.n695 gnd 0.013415f
C1406 commonsourceibias.n696 gnd 0.009605f
C1407 commonsourceibias.n697 gnd 0.009605f
C1408 commonsourceibias.n698 gnd 0.009605f
C1409 commonsourceibias.n699 gnd 0.011742f
C1410 commonsourceibias.n700 gnd 0.071604f
C1411 commonsourceibias.n701 gnd 0.012378f
C1412 commonsourceibias.t90 gnd 0.17946f
C1413 commonsourceibias.n702 gnd 0.071604f
C1414 commonsourceibias.n703 gnd 0.012558f
C1415 commonsourceibias.n704 gnd 0.009605f
C1416 commonsourceibias.n705 gnd 0.009605f
C1417 commonsourceibias.n706 gnd 0.009605f
C1418 commonsourceibias.n707 gnd 0.008375f
C1419 commonsourceibias.n708 gnd 0.013406f
C1420 commonsourceibias.n709 gnd 0.071604f
C1421 commonsourceibias.n710 gnd 0.01341f
C1422 commonsourceibias.n711 gnd 0.009605f
C1423 commonsourceibias.n712 gnd 0.009605f
C1424 commonsourceibias.n713 gnd 0.009605f
C1425 commonsourceibias.n714 gnd 0.011489f
C1426 commonsourceibias.n715 gnd 0.071604f
C1427 commonsourceibias.n716 gnd 0.012288f
C1428 commonsourceibias.t116 gnd 0.17946f
C1429 commonsourceibias.n717 gnd 0.071604f
C1430 commonsourceibias.n718 gnd 0.012648f
C1431 commonsourceibias.n719 gnd 0.009605f
C1432 commonsourceibias.n720 gnd 0.009605f
C1433 commonsourceibias.n721 gnd 0.009605f
C1434 commonsourceibias.n722 gnd 0.008208f
C1435 commonsourceibias.n723 gnd 0.013389f
C1436 commonsourceibias.n724 gnd 0.071604f
C1437 commonsourceibias.n725 gnd 0.013398f
C1438 commonsourceibias.n726 gnd 0.009605f
C1439 commonsourceibias.n727 gnd 0.009605f
C1440 commonsourceibias.n728 gnd 0.009605f
C1441 commonsourceibias.n729 gnd 0.011208f
C1442 commonsourceibias.n730 gnd 0.071604f
C1443 commonsourceibias.n731 gnd 0.011785f
C1444 commonsourceibias.n732 gnd 0.085919f
C1445 commonsourceibias.n733 gnd 0.056156f
C1446 commonsourceibias.n734 gnd 0.012817f
C1447 commonsourceibias.t180 gnd 0.17946f
C1448 commonsourceibias.n735 gnd 0.009349f
C1449 commonsourceibias.n736 gnd 0.009605f
C1450 commonsourceibias.t82 gnd 0.17946f
C1451 commonsourceibias.n737 gnd 0.012358f
C1452 commonsourceibias.n738 gnd 0.009605f
C1453 commonsourceibias.t179 gnd 0.17946f
C1454 commonsourceibias.n739 gnd 0.009057f
C1455 commonsourceibias.n740 gnd 0.009605f
C1456 commonsourceibias.t81 gnd 0.17946f
C1457 commonsourceibias.n741 gnd 0.012174f
C1458 commonsourceibias.n742 gnd 0.009605f
C1459 commonsourceibias.t178 gnd 0.17946f
C1460 commonsourceibias.n743 gnd 0.008798f
C1461 commonsourceibias.n744 gnd 0.009605f
C1462 commonsourceibias.t89 gnd 0.17946f
C1463 commonsourceibias.n745 gnd 0.01197f
C1464 commonsourceibias.n746 gnd 0.009605f
C1465 commonsourceibias.t97 gnd 0.17946f
C1466 commonsourceibias.n747 gnd 0.008571f
C1467 commonsourceibias.n748 gnd 0.009605f
C1468 commonsourceibias.t86 gnd 0.17946f
C1469 commonsourceibias.n749 gnd 0.011742f
C1470 commonsourceibias.n750 gnd 0.009605f
C1471 commonsourceibias.t106 gnd 0.17946f
C1472 commonsourceibias.n751 gnd 0.008375f
C1473 commonsourceibias.n752 gnd 0.009605f
C1474 commonsourceibias.t85 gnd 0.17946f
C1475 commonsourceibias.n753 gnd 0.011489f
C1476 commonsourceibias.n754 gnd 0.009605f
C1477 commonsourceibias.t104 gnd 0.17946f
C1478 commonsourceibias.n755 gnd 0.008208f
C1479 commonsourceibias.n756 gnd 0.009605f
C1480 commonsourceibias.t132 gnd 0.17946f
C1481 commonsourceibias.n757 gnd 0.011208f
C1482 commonsourceibias.t98 gnd 0.199526f
C1483 commonsourceibias.t123 gnd 0.17946f
C1484 commonsourceibias.n758 gnd 0.078221f
C1485 commonsourceibias.n759 gnd 0.085838f
C1486 commonsourceibias.n760 gnd 0.03983f
C1487 commonsourceibias.n761 gnd 0.009605f
C1488 commonsourceibias.n762 gnd 0.009349f
C1489 commonsourceibias.n763 gnd 0.013398f
C1490 commonsourceibias.n764 gnd 0.071604f
C1491 commonsourceibias.n765 gnd 0.013389f
C1492 commonsourceibias.n766 gnd 0.009605f
C1493 commonsourceibias.n767 gnd 0.009605f
C1494 commonsourceibias.n768 gnd 0.009605f
C1495 commonsourceibias.n769 gnd 0.012358f
C1496 commonsourceibias.n770 gnd 0.071604f
C1497 commonsourceibias.n771 gnd 0.012648f
C1498 commonsourceibias.t118 gnd 0.17946f
C1499 commonsourceibias.n772 gnd 0.071604f
C1500 commonsourceibias.n773 gnd 0.012288f
C1501 commonsourceibias.n774 gnd 0.009605f
C1502 commonsourceibias.n775 gnd 0.009605f
C1503 commonsourceibias.n776 gnd 0.009605f
C1504 commonsourceibias.n777 gnd 0.009057f
C1505 commonsourceibias.n778 gnd 0.01341f
C1506 commonsourceibias.n779 gnd 0.071604f
C1507 commonsourceibias.n780 gnd 0.013406f
C1508 commonsourceibias.n781 gnd 0.009605f
C1509 commonsourceibias.n782 gnd 0.009605f
C1510 commonsourceibias.n783 gnd 0.009605f
C1511 commonsourceibias.n784 gnd 0.012174f
C1512 commonsourceibias.n785 gnd 0.071604f
C1513 commonsourceibias.n786 gnd 0.012558f
C1514 commonsourceibias.t119 gnd 0.17946f
C1515 commonsourceibias.n787 gnd 0.071604f
C1516 commonsourceibias.n788 gnd 0.012378f
C1517 commonsourceibias.n789 gnd 0.009605f
C1518 commonsourceibias.n790 gnd 0.009605f
C1519 commonsourceibias.n791 gnd 0.009605f
C1520 commonsourceibias.n792 gnd 0.008798f
C1521 commonsourceibias.n793 gnd 0.013415f
C1522 commonsourceibias.n794 gnd 0.071604f
C1523 commonsourceibias.n795 gnd 0.013414f
C1524 commonsourceibias.n796 gnd 0.009605f
C1525 commonsourceibias.n797 gnd 0.009605f
C1526 commonsourceibias.n798 gnd 0.009605f
C1527 commonsourceibias.n799 gnd 0.01197f
C1528 commonsourceibias.n800 gnd 0.071604f
C1529 commonsourceibias.n801 gnd 0.012468f
C1530 commonsourceibias.t120 gnd 0.17946f
C1531 commonsourceibias.n802 gnd 0.071604f
C1532 commonsourceibias.n803 gnd 0.012468f
C1533 commonsourceibias.n804 gnd 0.009605f
C1534 commonsourceibias.n805 gnd 0.009605f
C1535 commonsourceibias.n806 gnd 0.009605f
C1536 commonsourceibias.n807 gnd 0.008571f
C1537 commonsourceibias.n808 gnd 0.013414f
C1538 commonsourceibias.n809 gnd 0.071604f
C1539 commonsourceibias.n810 gnd 0.013415f
C1540 commonsourceibias.n811 gnd 0.009605f
C1541 commonsourceibias.n812 gnd 0.009605f
C1542 commonsourceibias.n813 gnd 0.009605f
C1543 commonsourceibias.n814 gnd 0.011742f
C1544 commonsourceibias.n815 gnd 0.071604f
C1545 commonsourceibias.n816 gnd 0.012378f
C1546 commonsourceibias.t121 gnd 0.17946f
C1547 commonsourceibias.n817 gnd 0.071604f
C1548 commonsourceibias.n818 gnd 0.012558f
C1549 commonsourceibias.n819 gnd 0.009605f
C1550 commonsourceibias.n820 gnd 0.009605f
C1551 commonsourceibias.n821 gnd 0.009605f
C1552 commonsourceibias.n822 gnd 0.008375f
C1553 commonsourceibias.n823 gnd 0.013406f
C1554 commonsourceibias.n824 gnd 0.071604f
C1555 commonsourceibias.n825 gnd 0.01341f
C1556 commonsourceibias.n826 gnd 0.009605f
C1557 commonsourceibias.n827 gnd 0.009605f
C1558 commonsourceibias.n828 gnd 0.009605f
C1559 commonsourceibias.n829 gnd 0.011489f
C1560 commonsourceibias.n830 gnd 0.071604f
C1561 commonsourceibias.n831 gnd 0.012288f
C1562 commonsourceibias.t193 gnd 0.17946f
C1563 commonsourceibias.n832 gnd 0.071604f
C1564 commonsourceibias.n833 gnd 0.012648f
C1565 commonsourceibias.n834 gnd 0.009605f
C1566 commonsourceibias.n835 gnd 0.009605f
C1567 commonsourceibias.n836 gnd 0.009605f
C1568 commonsourceibias.n837 gnd 0.008208f
C1569 commonsourceibias.n838 gnd 0.013389f
C1570 commonsourceibias.n839 gnd 0.071604f
C1571 commonsourceibias.n840 gnd 0.013398f
C1572 commonsourceibias.n841 gnd 0.009605f
C1573 commonsourceibias.n842 gnd 0.009605f
C1574 commonsourceibias.n843 gnd 0.009605f
C1575 commonsourceibias.n844 gnd 0.011208f
C1576 commonsourceibias.n845 gnd 0.071604f
C1577 commonsourceibias.n846 gnd 0.011785f
C1578 commonsourceibias.t189 gnd 0.194086f
C1579 commonsourceibias.n847 gnd 0.085919f
C1580 commonsourceibias.n848 gnd 0.029883f
C1581 commonsourceibias.n849 gnd 0.153509f
C1582 commonsourceibias.n850 gnd 0.012817f
C1583 commonsourceibias.t133 gnd 0.17946f
C1584 commonsourceibias.n851 gnd 0.009349f
C1585 commonsourceibias.n852 gnd 0.009605f
C1586 commonsourceibias.t153 gnd 0.17946f
C1587 commonsourceibias.n853 gnd 0.012358f
C1588 commonsourceibias.n854 gnd 0.009605f
C1589 commonsourceibias.t122 gnd 0.17946f
C1590 commonsourceibias.n855 gnd 0.009057f
C1591 commonsourceibias.n856 gnd 0.009605f
C1592 commonsourceibias.t143 gnd 0.17946f
C1593 commonsourceibias.n857 gnd 0.012174f
C1594 commonsourceibias.n858 gnd 0.009605f
C1595 commonsourceibias.t99 gnd 0.17946f
C1596 commonsourceibias.n859 gnd 0.008798f
C1597 commonsourceibias.n860 gnd 0.009605f
C1598 commonsourceibias.t87 gnd 0.17946f
C1599 commonsourceibias.n861 gnd 0.01197f
C1600 commonsourceibias.n862 gnd 0.009605f
C1601 commonsourceibias.t167 gnd 0.17946f
C1602 commonsourceibias.n863 gnd 0.008571f
C1603 commonsourceibias.n864 gnd 0.009605f
C1604 commonsourceibias.t192 gnd 0.17946f
C1605 commonsourceibias.n865 gnd 0.011742f
C1606 commonsourceibias.n866 gnd 0.009605f
C1607 commonsourceibias.t136 gnd 0.17946f
C1608 commonsourceibias.n867 gnd 0.008375f
C1609 commonsourceibias.n868 gnd 0.009605f
C1610 commonsourceibias.t181 gnd 0.17946f
C1611 commonsourceibias.n869 gnd 0.011489f
C1612 commonsourceibias.n870 gnd 0.009605f
C1613 commonsourceibias.t126 gnd 0.17946f
C1614 commonsourceibias.n871 gnd 0.008208f
C1615 commonsourceibias.n872 gnd 0.009605f
C1616 commonsourceibias.t146 gnd 0.17946f
C1617 commonsourceibias.n873 gnd 0.011208f
C1618 commonsourceibias.t191 gnd 0.199526f
C1619 commonsourceibias.t156 gnd 0.17946f
C1620 commonsourceibias.n874 gnd 0.078221f
C1621 commonsourceibias.n875 gnd 0.085838f
C1622 commonsourceibias.n876 gnd 0.03983f
C1623 commonsourceibias.n877 gnd 0.009605f
C1624 commonsourceibias.n878 gnd 0.009349f
C1625 commonsourceibias.n879 gnd 0.013398f
C1626 commonsourceibias.n880 gnd 0.071604f
C1627 commonsourceibias.n881 gnd 0.013389f
C1628 commonsourceibias.n882 gnd 0.009605f
C1629 commonsourceibias.n883 gnd 0.009605f
C1630 commonsourceibias.n884 gnd 0.009605f
C1631 commonsourceibias.n885 gnd 0.012358f
C1632 commonsourceibias.n886 gnd 0.071604f
C1633 commonsourceibias.n887 gnd 0.012648f
C1634 commonsourceibias.t91 gnd 0.17946f
C1635 commonsourceibias.n888 gnd 0.071604f
C1636 commonsourceibias.n889 gnd 0.012288f
C1637 commonsourceibias.n890 gnd 0.009605f
C1638 commonsourceibias.n891 gnd 0.009605f
C1639 commonsourceibias.n892 gnd 0.009605f
C1640 commonsourceibias.n893 gnd 0.009057f
C1641 commonsourceibias.n894 gnd 0.01341f
C1642 commonsourceibias.n895 gnd 0.071604f
C1643 commonsourceibias.n896 gnd 0.013406f
C1644 commonsourceibias.n897 gnd 0.009605f
C1645 commonsourceibias.n898 gnd 0.009605f
C1646 commonsourceibias.n899 gnd 0.009605f
C1647 commonsourceibias.n900 gnd 0.012174f
C1648 commonsourceibias.n901 gnd 0.071604f
C1649 commonsourceibias.n902 gnd 0.012558f
C1650 commonsourceibias.t107 gnd 0.17946f
C1651 commonsourceibias.n903 gnd 0.071604f
C1652 commonsourceibias.n904 gnd 0.012378f
C1653 commonsourceibias.n905 gnd 0.009605f
C1654 commonsourceibias.n906 gnd 0.009605f
C1655 commonsourceibias.n907 gnd 0.009605f
C1656 commonsourceibias.n908 gnd 0.008798f
C1657 commonsourceibias.n909 gnd 0.013415f
C1658 commonsourceibias.n910 gnd 0.071604f
C1659 commonsourceibias.n911 gnd 0.013414f
C1660 commonsourceibias.n912 gnd 0.009605f
C1661 commonsourceibias.n913 gnd 0.009605f
C1662 commonsourceibias.n914 gnd 0.009605f
C1663 commonsourceibias.n915 gnd 0.01197f
C1664 commonsourceibias.n916 gnd 0.071604f
C1665 commonsourceibias.n917 gnd 0.012468f
C1666 commonsourceibias.t127 gnd 0.17946f
C1667 commonsourceibias.n918 gnd 0.071604f
C1668 commonsourceibias.n919 gnd 0.012468f
C1669 commonsourceibias.n920 gnd 0.009605f
C1670 commonsourceibias.n921 gnd 0.009605f
C1671 commonsourceibias.n922 gnd 0.009605f
C1672 commonsourceibias.n923 gnd 0.008571f
C1673 commonsourceibias.n924 gnd 0.013414f
C1674 commonsourceibias.n925 gnd 0.071604f
C1675 commonsourceibias.n926 gnd 0.013415f
C1676 commonsourceibias.n927 gnd 0.009605f
C1677 commonsourceibias.n928 gnd 0.009605f
C1678 commonsourceibias.n929 gnd 0.009605f
C1679 commonsourceibias.n930 gnd 0.011742f
C1680 commonsourceibias.n931 gnd 0.071604f
C1681 commonsourceibias.n932 gnd 0.012378f
C1682 commonsourceibias.t137 gnd 0.17946f
C1683 commonsourceibias.n933 gnd 0.071604f
C1684 commonsourceibias.n934 gnd 0.012558f
C1685 commonsourceibias.n935 gnd 0.009605f
C1686 commonsourceibias.n936 gnd 0.009605f
C1687 commonsourceibias.n937 gnd 0.009605f
C1688 commonsourceibias.n938 gnd 0.008375f
C1689 commonsourceibias.n939 gnd 0.013406f
C1690 commonsourceibias.n940 gnd 0.071604f
C1691 commonsourceibias.n941 gnd 0.01341f
C1692 commonsourceibias.n942 gnd 0.009605f
C1693 commonsourceibias.n943 gnd 0.009605f
C1694 commonsourceibias.n944 gnd 0.009605f
C1695 commonsourceibias.n945 gnd 0.011489f
C1696 commonsourceibias.n946 gnd 0.071604f
C1697 commonsourceibias.n947 gnd 0.012288f
C1698 commonsourceibias.t170 gnd 0.17946f
C1699 commonsourceibias.n948 gnd 0.071604f
C1700 commonsourceibias.n949 gnd 0.012648f
C1701 commonsourceibias.n950 gnd 0.009605f
C1702 commonsourceibias.n951 gnd 0.009605f
C1703 commonsourceibias.n952 gnd 0.009605f
C1704 commonsourceibias.n953 gnd 0.008208f
C1705 commonsourceibias.n954 gnd 0.013389f
C1706 commonsourceibias.n955 gnd 0.071604f
C1707 commonsourceibias.n956 gnd 0.013398f
C1708 commonsourceibias.n957 gnd 0.009605f
C1709 commonsourceibias.n958 gnd 0.009605f
C1710 commonsourceibias.n959 gnd 0.009605f
C1711 commonsourceibias.n960 gnd 0.011208f
C1712 commonsourceibias.n961 gnd 0.071604f
C1713 commonsourceibias.n962 gnd 0.011785f
C1714 commonsourceibias.t101 gnd 0.194086f
C1715 commonsourceibias.n963 gnd 0.085919f
C1716 commonsourceibias.n964 gnd 0.029883f
C1717 commonsourceibias.n965 gnd 0.202572f
C1718 commonsourceibias.n966 gnd 5.28148f
C1719 a_n2140_13878.t11 gnd 0.186868f
C1720 a_n2140_13878.t10 gnd 0.186868f
C1721 a_n2140_13878.t5 gnd 0.186868f
C1722 a_n2140_13878.n0 gnd 1.47299f
C1723 a_n2140_13878.t2 gnd 0.186868f
C1724 a_n2140_13878.t4 gnd 0.186868f
C1725 a_n2140_13878.n1 gnd 1.47143f
C1726 a_n2140_13878.n2 gnd 2.05603f
C1727 a_n2140_13878.t12 gnd 0.186868f
C1728 a_n2140_13878.t3 gnd 0.186868f
C1729 a_n2140_13878.n3 gnd 1.47143f
C1730 a_n2140_13878.n4 gnd 1.00289f
C1731 a_n2140_13878.t9 gnd 0.186868f
C1732 a_n2140_13878.t1 gnd 0.186868f
C1733 a_n2140_13878.n5 gnd 1.47143f
C1734 a_n2140_13878.n6 gnd 4.06212f
C1735 a_n2140_13878.t17 gnd 1.74974f
C1736 a_n2140_13878.t20 gnd 0.186868f
C1737 a_n2140_13878.t21 gnd 0.186868f
C1738 a_n2140_13878.n7 gnd 1.3163f
C1739 a_n2140_13878.n8 gnd 1.47077f
C1740 a_n2140_13878.t16 gnd 1.74626f
C1741 a_n2140_13878.n9 gnd 0.740113f
C1742 a_n2140_13878.t19 gnd 1.74626f
C1743 a_n2140_13878.n10 gnd 0.740113f
C1744 a_n2140_13878.t22 gnd 0.186868f
C1745 a_n2140_13878.t23 gnd 0.186868f
C1746 a_n2140_13878.n11 gnd 1.3163f
C1747 a_n2140_13878.n12 gnd 0.74728f
C1748 a_n2140_13878.t18 gnd 1.74626f
C1749 a_n2140_13878.n13 gnd 2.09583f
C1750 a_n2140_13878.n14 gnd 2.85974f
C1751 a_n2140_13878.t6 gnd 0.186868f
C1752 a_n2140_13878.t7 gnd 0.186868f
C1753 a_n2140_13878.n15 gnd 1.47142f
C1754 a_n2140_13878.n16 gnd 2.01665f
C1755 a_n2140_13878.t13 gnd 0.186868f
C1756 a_n2140_13878.t14 gnd 0.186868f
C1757 a_n2140_13878.n17 gnd 1.47143f
C1758 a_n2140_13878.n18 gnd 0.651951f
C1759 a_n2140_13878.t0 gnd 0.186868f
C1760 a_n2140_13878.t8 gnd 0.186868f
C1761 a_n2140_13878.n19 gnd 1.47143f
C1762 a_n2140_13878.n20 gnd 1.32263f
C1763 a_n2140_13878.n21 gnd 1.47386f
C1764 a_n2140_13878.t15 gnd 0.186868f
C1765 a_n2408_n452.n0 gnd 3.95093f
C1766 a_n2408_n452.n1 gnd 2.90522f
C1767 a_n2408_n452.n2 gnd 3.88871f
C1768 a_n2408_n452.n3 gnd 0.820088f
C1769 a_n2408_n452.n4 gnd 0.82009f
C1770 a_n2408_n452.n5 gnd 0.668637f
C1771 a_n2408_n452.n6 gnd 0.204926f
C1772 a_n2408_n452.n7 gnd 0.150932f
C1773 a_n2408_n452.n8 gnd 0.237216f
C1774 a_n2408_n452.n9 gnd 0.183222f
C1775 a_n2408_n452.n10 gnd 0.204926f
C1776 a_n2408_n452.n11 gnd 1.1184f
C1777 a_n2408_n452.n12 gnd 0.150932f
C1778 a_n2408_n452.n13 gnd 0.722632f
C1779 a_n2408_n452.n14 gnd 0.512478f
C1780 a_n2408_n452.n15 gnd 0.215976f
C1781 a_n2408_n452.n16 gnd 0.215976f
C1782 a_n2408_n452.n17 gnd 0.44388f
C1783 a_n2408_n452.n18 gnd 0.215976f
C1784 a_n2408_n452.n19 gnd 0.215976f
C1785 a_n2408_n452.n20 gnd 0.215976f
C1786 a_n2408_n452.n21 gnd 0.747109f
C1787 a_n2408_n452.n22 gnd 0.215976f
C1788 a_n2408_n452.n23 gnd 0.44388f
C1789 a_n2408_n452.n24 gnd 3.3281f
C1790 a_n2408_n452.n25 gnd 0.668661f
C1791 a_n2408_n452.n26 gnd 0.215976f
C1792 a_n2408_n452.n27 gnd 1.7781f
C1793 a_n2408_n452.n28 gnd 2.07945f
C1794 a_n2408_n452.n29 gnd 1.89786f
C1795 a_n2408_n452.n30 gnd 1.7781f
C1796 a_n2408_n452.n31 gnd 0.285304f
C1797 a_n2408_n452.n32 gnd 0.004854f
C1798 a_n2408_n452.n33 gnd 0.010499f
C1799 a_n2408_n452.n34 gnd 0.010499f
C1800 a_n2408_n452.n35 gnd 0.285304f
C1801 a_n2408_n452.n36 gnd 0.285304f
C1802 a_n2408_n452.n37 gnd 0.004854f
C1803 a_n2408_n452.n38 gnd 0.010499f
C1804 a_n2408_n452.n39 gnd 0.010499f
C1805 a_n2408_n452.n40 gnd 0.004854f
C1806 a_n2408_n452.n41 gnd 0.285304f
C1807 a_n2408_n452.n42 gnd 0.285304f
C1808 a_n2408_n452.n43 gnd 0.76008f
C1809 a_n2408_n452.n44 gnd 0.004854f
C1810 a_n2408_n452.n45 gnd 0.010499f
C1811 a_n2408_n452.n46 gnd 0.010499f
C1812 a_n2408_n452.n47 gnd 0.004854f
C1813 a_n2408_n452.n48 gnd 0.285304f
C1814 a_n2408_n452.n49 gnd 0.285304f
C1815 a_n2408_n452.n50 gnd 0.44388f
C1816 a_n2408_n452.n51 gnd 0.004854f
C1817 a_n2408_n452.n52 gnd 0.010499f
C1818 a_n2408_n452.n53 gnd 0.010499f
C1819 a_n2408_n452.n54 gnd 0.004854f
C1820 a_n2408_n452.n55 gnd 0.285304f
C1821 a_n2408_n452.n56 gnd 0.008362f
C1822 a_n2408_n452.n57 gnd 0.285304f
C1823 a_n2408_n452.n58 gnd 0.008362f
C1824 a_n2408_n452.n59 gnd 0.285304f
C1825 a_n2408_n452.n60 gnd 0.008362f
C1826 a_n2408_n452.n61 gnd 0.285304f
C1827 a_n2408_n452.n62 gnd 0.008362f
C1828 a_n2408_n452.n63 gnd 0.285304f
C1829 a_n2408_n452.n64 gnd 0.004854f
C1830 a_n2408_n452.n65 gnd 0.304392f
C1831 a_n2408_n452.t15 gnd 0.149803f
C1832 a_n2408_n452.t8 gnd 0.708488f
C1833 a_n2408_n452.t16 gnd 0.696812f
C1834 a_n2408_n452.t6 gnd 0.696812f
C1835 a_n2408_n452.n66 gnd 0.304392f
C1836 a_n2408_n452.t14 gnd 0.696812f
C1837 a_n2408_n452.t2 gnd 0.696812f
C1838 a_n2408_n452.t22 gnd 0.696812f
C1839 a_n2408_n452.t12 gnd 0.708488f
C1840 a_n2408_n452.t86 gnd 0.708488f
C1841 a_n2408_n452.t67 gnd 0.696812f
C1842 a_n2408_n452.t71 gnd 0.696812f
C1843 a_n2408_n452.n67 gnd 0.304392f
C1844 a_n2408_n452.t61 gnd 0.696812f
C1845 a_n2408_n452.t76 gnd 0.696812f
C1846 a_n2408_n452.t83 gnd 0.696812f
C1847 a_n2408_n452.n68 gnd 0.304392f
C1848 a_n2408_n452.t84 gnd 0.696812f
C1849 a_n2408_n452.t58 gnd 0.708488f
C1850 a_n2408_n452.t19 gnd 1.40268f
C1851 a_n2408_n452.t25 gnd 0.149803f
C1852 a_n2408_n452.t31 gnd 0.149803f
C1853 a_n2408_n452.n69 gnd 1.05521f
C1854 a_n2408_n452.t33 gnd 0.149803f
C1855 a_n2408_n452.t21 gnd 0.149803f
C1856 a_n2408_n452.n70 gnd 1.05521f
C1857 a_n2408_n452.t11 gnd 0.149803f
C1858 a_n2408_n452.t29 gnd 0.149803f
C1859 a_n2408_n452.n71 gnd 1.05521f
C1860 a_n2408_n452.t27 gnd 1.39988f
C1861 a_n2408_n452.t10 gnd 0.696812f
C1862 a_n2408_n452.n72 gnd 0.304392f
C1863 a_n2408_n452.t32 gnd 0.696812f
C1864 a_n2408_n452.t18 gnd 0.708488f
C1865 a_n2408_n452.t24 gnd 0.696812f
C1866 a_n2408_n452.t66 gnd 0.696812f
C1867 a_n2408_n452.n73 gnd 0.304392f
C1868 a_n2408_n452.t80 gnd 0.696812f
C1869 a_n2408_n452.t82 gnd 0.708488f
C1870 a_n2408_n452.t60 gnd 0.696812f
C1871 a_n2408_n452.n74 gnd 0.306874f
C1872 a_n2408_n452.t79 gnd 0.696812f
C1873 a_n2408_n452.n75 gnd 0.304392f
C1874 a_n2408_n452.n76 gnd 0.299809f
C1875 a_n2408_n452.t57 gnd 0.696812f
C1876 a_n2408_n452.n77 gnd 0.299809f
C1877 a_n2408_n452.t74 gnd 0.696812f
C1878 a_n2408_n452.n78 gnd 0.306874f
C1879 a_n2408_n452.t59 gnd 0.708488f
C1880 a_n2408_n452.n79 gnd 0.306874f
C1881 a_n2408_n452.t30 gnd 0.696812f
C1882 a_n2408_n452.n80 gnd 0.304392f
C1883 a_n2408_n452.n81 gnd 0.299809f
C1884 a_n2408_n452.t20 gnd 0.696812f
C1885 a_n2408_n452.n82 gnd 0.299809f
C1886 a_n2408_n452.t28 gnd 0.696812f
C1887 a_n2408_n452.n83 gnd 0.306874f
C1888 a_n2408_n452.t26 gnd 0.708488f
C1889 a_n2408_n452.n84 gnd 1.19872f
C1890 a_n2408_n452.t64 gnd 0.696812f
C1891 a_n2408_n452.n85 gnd 0.302472f
C1892 a_n2408_n452.t70 gnd 0.696812f
C1893 a_n2408_n452.n86 gnd 0.302472f
C1894 a_n2408_n452.t62 gnd 0.696812f
C1895 a_n2408_n452.n87 gnd 0.302472f
C1896 a_n2408_n452.t75 gnd 0.696812f
C1897 a_n2408_n452.n88 gnd 0.302472f
C1898 a_n2408_n452.t65 gnd 0.696812f
C1899 a_n2408_n452.n89 gnd 0.296979f
C1900 a_n2408_n452.t87 gnd 0.696812f
C1901 a_n2408_n452.n90 gnd 0.306363f
C1902 a_n2408_n452.t68 gnd 0.708488f
C1903 a_n2408_n452.t77 gnd 0.696812f
C1904 a_n2408_n452.n91 gnd 0.296979f
C1905 a_n2408_n452.t63 gnd 0.696812f
C1906 a_n2408_n452.n92 gnd 0.306363f
C1907 a_n2408_n452.t72 gnd 0.708488f
C1908 a_n2408_n452.t81 gnd 0.696812f
C1909 a_n2408_n452.n93 gnd 0.296979f
C1910 a_n2408_n452.t69 gnd 0.696812f
C1911 a_n2408_n452.n94 gnd 0.306363f
C1912 a_n2408_n452.t85 gnd 0.708488f
C1913 a_n2408_n452.t73 gnd 0.696812f
C1914 a_n2408_n452.n95 gnd 0.296979f
C1915 a_n2408_n452.t56 gnd 0.696812f
C1916 a_n2408_n452.n96 gnd 0.306363f
C1917 a_n2408_n452.t78 gnd 0.708488f
C1918 a_n2408_n452.n97 gnd 1.45046f
C1919 a_n2408_n452.n98 gnd 0.306874f
C1920 a_n2408_n452.n99 gnd 0.299809f
C1921 a_n2408_n452.n100 gnd 0.299809f
C1922 a_n2408_n452.n101 gnd 0.306874f
C1923 a_n2408_n452.t4 gnd 0.696812f
C1924 a_n2408_n452.n102 gnd 0.306874f
C1925 a_n2408_n452.t49 gnd 0.116514f
C1926 a_n2408_n452.t52 gnd 0.116514f
C1927 a_n2408_n452.n103 gnd 1.03184f
C1928 a_n2408_n452.t0 gnd 0.116514f
C1929 a_n2408_n452.t38 gnd 0.116514f
C1930 a_n2408_n452.n104 gnd 1.02955f
C1931 a_n2408_n452.t1 gnd 0.116514f
C1932 a_n2408_n452.t50 gnd 0.116514f
C1933 a_n2408_n452.n105 gnd 1.02955f
C1934 a_n2408_n452.t41 gnd 0.116514f
C1935 a_n2408_n452.t46 gnd 0.116514f
C1936 a_n2408_n452.n106 gnd 1.03184f
C1937 a_n2408_n452.t37 gnd 0.116514f
C1938 a_n2408_n452.t43 gnd 0.116514f
C1939 a_n2408_n452.n107 gnd 1.02955f
C1940 a_n2408_n452.t48 gnd 0.116514f
C1941 a_n2408_n452.t55 gnd 0.116514f
C1942 a_n2408_n452.n108 gnd 1.02955f
C1943 a_n2408_n452.t53 gnd 0.116514f
C1944 a_n2408_n452.t39 gnd 0.116514f
C1945 a_n2408_n452.n109 gnd 1.02956f
C1946 a_n2408_n452.t44 gnd 0.116514f
C1947 a_n2408_n452.t47 gnd 0.116514f
C1948 a_n2408_n452.n110 gnd 1.02956f
C1949 a_n2408_n452.t54 gnd 0.116514f
C1950 a_n2408_n452.t34 gnd 0.116514f
C1951 a_n2408_n452.n111 gnd 1.02956f
C1952 a_n2408_n452.t36 gnd 0.116514f
C1953 a_n2408_n452.t45 gnd 0.116514f
C1954 a_n2408_n452.n112 gnd 1.03184f
C1955 a_n2408_n452.t42 gnd 0.116514f
C1956 a_n2408_n452.t40 gnd 0.116514f
C1957 a_n2408_n452.n113 gnd 1.02956f
C1958 a_n2408_n452.t35 gnd 0.116514f
C1959 a_n2408_n452.t51 gnd 0.116514f
C1960 a_n2408_n452.n114 gnd 1.02956f
C1961 a_n2408_n452.n115 gnd 0.299809f
C1962 a_n2408_n452.n116 gnd 0.299809f
C1963 a_n2408_n452.n117 gnd 0.306874f
C1964 a_n2408_n452.n118 gnd 0.859759f
C1965 a_n2408_n452.t9 gnd 1.39989f
C1966 a_n2408_n452.t17 gnd 0.149803f
C1967 a_n2408_n452.t7 gnd 0.149803f
C1968 a_n2408_n452.n119 gnd 1.05521f
C1969 a_n2408_n452.t13 gnd 1.40268f
C1970 a_n2408_n452.t23 gnd 0.149803f
C1971 a_n2408_n452.t5 gnd 0.149803f
C1972 a_n2408_n452.n120 gnd 1.05521f
C1973 a_n2408_n452.n121 gnd 1.05522f
C1974 a_n2408_n452.t3 gnd 0.149803f
C1975 a_n2903_n3924.t29 gnd 0.102925f
C1976 a_n2903_n3924.t35 gnd 0.102925f
C1977 a_n2903_n3924.n0 gnd 0.840607f
C1978 a_n2903_n3924.n1 gnd 0.382272f
C1979 a_n2903_n3924.t38 gnd 1.06972f
C1980 a_n2903_n3924.n2 gnd 0.962269f
C1981 a_n2903_n3924.t18 gnd 0.102925f
C1982 a_n2903_n3924.t36 gnd 0.102925f
C1983 a_n2903_n3924.n3 gnd 0.840608f
C1984 a_n2903_n3924.n4 gnd 0.382271f
C1985 a_n2903_n3924.t32 gnd 0.102925f
C1986 a_n2903_n3924.t34 gnd 0.102925f
C1987 a_n2903_n3924.n5 gnd 0.840608f
C1988 a_n2903_n3924.n6 gnd 0.382271f
C1989 a_n2903_n3924.t37 gnd 0.102925f
C1990 a_n2903_n3924.t39 gnd 0.102925f
C1991 a_n2903_n3924.n7 gnd 0.840608f
C1992 a_n2903_n3924.n8 gnd 0.382271f
C1993 a_n2903_n3924.t21 gnd 0.102925f
C1994 a_n2903_n3924.t19 gnd 0.102925f
C1995 a_n2903_n3924.n9 gnd 0.840608f
C1996 a_n2903_n3924.n10 gnd 0.382271f
C1997 a_n2903_n3924.t27 gnd 0.102925f
C1998 a_n2903_n3924.t20 gnd 0.102925f
C1999 a_n2903_n3924.n11 gnd 0.840608f
C2000 a_n2903_n3924.n12 gnd 0.382271f
C2001 a_n2903_n3924.t26 gnd 1.06972f
C2002 a_n2903_n3924.n13 gnd 0.383728f
C2003 a_n2903_n3924.t43 gnd 1.06972f
C2004 a_n2903_n3924.n14 gnd 0.383728f
C2005 a_n2903_n3924.t11 gnd 0.102925f
C2006 a_n2903_n3924.t6 gnd 0.102925f
C2007 a_n2903_n3924.n15 gnd 0.840608f
C2008 a_n2903_n3924.n16 gnd 0.382271f
C2009 a_n2903_n3924.t50 gnd 0.102925f
C2010 a_n2903_n3924.t14 gnd 0.102925f
C2011 a_n2903_n3924.n17 gnd 0.840608f
C2012 a_n2903_n3924.n18 gnd 0.382271f
C2013 a_n2903_n3924.t3 gnd 0.102925f
C2014 a_n2903_n3924.t4 gnd 0.102925f
C2015 a_n2903_n3924.n19 gnd 0.840608f
C2016 a_n2903_n3924.n20 gnd 0.382271f
C2017 a_n2903_n3924.t45 gnd 0.102925f
C2018 a_n2903_n3924.t54 gnd 0.102925f
C2019 a_n2903_n3924.n21 gnd 0.840608f
C2020 a_n2903_n3924.n22 gnd 0.382271f
C2021 a_n2903_n3924.t10 gnd 0.102925f
C2022 a_n2903_n3924.t17 gnd 0.102925f
C2023 a_n2903_n3924.n23 gnd 0.840608f
C2024 a_n2903_n3924.n24 gnd 0.382271f
C2025 a_n2903_n3924.t53 gnd 1.06972f
C2026 a_n2903_n3924.n25 gnd 0.962265f
C2027 a_n2903_n3924.t24 gnd 0.102925f
C2028 a_n2903_n3924.t30 gnd 0.102925f
C2029 a_n2903_n3924.n26 gnd 0.840607f
C2030 a_n2903_n3924.n27 gnd 0.382272f
C2031 a_n2903_n3924.t25 gnd 1.06972f
C2032 a_n2903_n3924.n28 gnd 0.625684f
C2033 a_n2903_n3924.n29 gnd 0.965474f
C2034 a_n2903_n3924.t2 gnd 1.32974f
C2035 a_n2903_n3924.n30 gnd 0.928343f
C2036 a_n2903_n3924.t12 gnd 1.3291f
C2037 a_n2903_n3924.n31 gnd 0.766359f
C2038 a_n2903_n3924.t48 gnd 1.3291f
C2039 a_n2903_n3924.n32 gnd 0.936111f
C2040 a_n2903_n3924.t15 gnd 1.3291f
C2041 a_n2903_n3924.n33 gnd 0.936111f
C2042 a_n2903_n3924.t9 gnd 1.3291f
C2043 a_n2903_n3924.n34 gnd 0.936111f
C2044 a_n2903_n3924.t42 gnd 1.3291f
C2045 a_n2903_n3924.n35 gnd 0.936111f
C2046 a_n2903_n3924.t5 gnd 1.3291f
C2047 a_n2903_n3924.n36 gnd 0.936111f
C2048 a_n2903_n3924.t52 gnd 1.3291f
C2049 a_n2903_n3924.n37 gnd 1.25723f
C2050 a_n2903_n3924.n38 gnd 1.02539f
C2051 a_n2903_n3924.t44 gnd 1.06972f
C2052 a_n2903_n3924.n39 gnd 0.625684f
C2053 a_n2903_n3924.t16 gnd 0.102925f
C2054 a_n2903_n3924.t13 gnd 0.102925f
C2055 a_n2903_n3924.n40 gnd 0.840607f
C2056 a_n2903_n3924.n41 gnd 0.382272f
C2057 a_n2903_n3924.t55 gnd 0.102925f
C2058 a_n2903_n3924.t7 gnd 0.102925f
C2059 a_n2903_n3924.n42 gnd 0.840607f
C2060 a_n2903_n3924.n43 gnd 0.382272f
C2061 a_n2903_n3924.t49 gnd 0.102925f
C2062 a_n2903_n3924.t46 gnd 0.102925f
C2063 a_n2903_n3924.n44 gnd 0.840607f
C2064 a_n2903_n3924.n45 gnd 0.382272f
C2065 a_n2903_n3924.t8 gnd 0.102925f
C2066 a_n2903_n3924.t1 gnd 0.102925f
C2067 a_n2903_n3924.n46 gnd 0.840607f
C2068 a_n2903_n3924.n47 gnd 0.382272f
C2069 a_n2903_n3924.t51 gnd 0.102925f
C2070 a_n2903_n3924.t0 gnd 0.102925f
C2071 a_n2903_n3924.n48 gnd 0.840607f
C2072 a_n2903_n3924.n49 gnd 0.382272f
C2073 a_n2903_n3924.t47 gnd 1.06972f
C2074 a_n2903_n3924.n50 gnd 0.383732f
C2075 a_n2903_n3924.t31 gnd 1.06972f
C2076 a_n2903_n3924.n51 gnd 0.383732f
C2077 a_n2903_n3924.t28 gnd 0.102925f
C2078 a_n2903_n3924.t33 gnd 0.102925f
C2079 a_n2903_n3924.n52 gnd 0.840607f
C2080 a_n2903_n3924.n53 gnd 0.382272f
C2081 a_n2903_n3924.t23 gnd 0.102925f
C2082 a_n2903_n3924.t22 gnd 0.102925f
C2083 a_n2903_n3924.n54 gnd 0.840607f
C2084 a_n2903_n3924.n55 gnd 0.382272f
C2085 a_n2903_n3924.n56 gnd 0.382275f
C2086 a_n2903_n3924.t40 gnd 0.102925f
C2087 a_n2903_n3924.n57 gnd 0.840604f
C2088 a_n2903_n3924.t41 gnd 0.102925f
C2089 plus.n0 gnd 0.023384f
C2090 plus.t21 gnd 0.330743f
C2091 plus.n1 gnd 0.023384f
C2092 plus.t22 gnd 0.330743f
C2093 plus.t16 gnd 0.330743f
C2094 plus.n2 gnd 0.146927f
C2095 plus.n3 gnd 0.023384f
C2096 plus.t17 gnd 0.330743f
C2097 plus.t11 gnd 0.330743f
C2098 plus.n4 gnd 0.146927f
C2099 plus.n5 gnd 0.023384f
C2100 plus.t5 gnd 0.330743f
C2101 plus.t6 gnd 0.330743f
C2102 plus.n6 gnd 0.146927f
C2103 plus.n7 gnd 0.023384f
C2104 plus.t23 gnd 0.330743f
C2105 plus.t24 gnd 0.330743f
C2106 plus.n8 gnd 0.146927f
C2107 plus.n9 gnd 0.023384f
C2108 plus.t18 gnd 0.330743f
C2109 plus.t13 gnd 0.330743f
C2110 plus.n10 gnd 0.151712f
C2111 plus.t15 gnd 0.342749f
C2112 plus.n11 gnd 0.136166f
C2113 plus.n12 gnd 0.100669f
C2114 plus.n13 gnd 0.005306f
C2115 plus.n14 gnd 0.146927f
C2116 plus.n15 gnd 0.005306f
C2117 plus.n16 gnd 0.023384f
C2118 plus.n17 gnd 0.023384f
C2119 plus.n18 gnd 0.023384f
C2120 plus.n19 gnd 0.005306f
C2121 plus.n20 gnd 0.146927f
C2122 plus.n21 gnd 0.005306f
C2123 plus.n22 gnd 0.023384f
C2124 plus.n23 gnd 0.023384f
C2125 plus.n24 gnd 0.023384f
C2126 plus.n25 gnd 0.005306f
C2127 plus.n26 gnd 0.146927f
C2128 plus.n27 gnd 0.005306f
C2129 plus.n28 gnd 0.023384f
C2130 plus.n29 gnd 0.023384f
C2131 plus.n30 gnd 0.023384f
C2132 plus.n31 gnd 0.005306f
C2133 plus.n32 gnd 0.146927f
C2134 plus.n33 gnd 0.005306f
C2135 plus.n34 gnd 0.023384f
C2136 plus.n35 gnd 0.023384f
C2137 plus.n36 gnd 0.023384f
C2138 plus.n37 gnd 0.005306f
C2139 plus.n38 gnd 0.146927f
C2140 plus.n39 gnd 0.005306f
C2141 plus.n40 gnd 0.147143f
C2142 plus.n41 gnd 0.264786f
C2143 plus.n42 gnd 0.023384f
C2144 plus.n43 gnd 0.005306f
C2145 plus.t10 gnd 0.330743f
C2146 plus.n44 gnd 0.023384f
C2147 plus.n45 gnd 0.005306f
C2148 plus.t12 gnd 0.330743f
C2149 plus.n46 gnd 0.023384f
C2150 plus.n47 gnd 0.005306f
C2151 plus.t7 gnd 0.330743f
C2152 plus.n48 gnd 0.023384f
C2153 plus.n49 gnd 0.005306f
C2154 plus.t27 gnd 0.330743f
C2155 plus.n50 gnd 0.023384f
C2156 plus.n51 gnd 0.005306f
C2157 plus.t26 gnd 0.330743f
C2158 plus.t20 gnd 0.342749f
C2159 plus.t19 gnd 0.330743f
C2160 plus.n52 gnd 0.151712f
C2161 plus.n53 gnd 0.136166f
C2162 plus.n54 gnd 0.100669f
C2163 plus.n55 gnd 0.023384f
C2164 plus.n56 gnd 0.146927f
C2165 plus.n57 gnd 0.005306f
C2166 plus.t25 gnd 0.330743f
C2167 plus.n58 gnd 0.146927f
C2168 plus.n59 gnd 0.023384f
C2169 plus.n60 gnd 0.023384f
C2170 plus.n61 gnd 0.023384f
C2171 plus.n62 gnd 0.146927f
C2172 plus.n63 gnd 0.005306f
C2173 plus.t9 gnd 0.330743f
C2174 plus.n64 gnd 0.146927f
C2175 plus.n65 gnd 0.023384f
C2176 plus.n66 gnd 0.023384f
C2177 plus.n67 gnd 0.023384f
C2178 plus.n68 gnd 0.146927f
C2179 plus.n69 gnd 0.005306f
C2180 plus.t14 gnd 0.330743f
C2181 plus.n70 gnd 0.146927f
C2182 plus.n71 gnd 0.023384f
C2183 plus.n72 gnd 0.023384f
C2184 plus.n73 gnd 0.023384f
C2185 plus.n74 gnd 0.146927f
C2186 plus.n75 gnd 0.005306f
C2187 plus.t28 gnd 0.330743f
C2188 plus.n76 gnd 0.146927f
C2189 plus.n77 gnd 0.023384f
C2190 plus.n78 gnd 0.023384f
C2191 plus.n79 gnd 0.023384f
C2192 plus.n80 gnd 0.146927f
C2193 plus.n81 gnd 0.005306f
C2194 plus.t8 gnd 0.330743f
C2195 plus.n82 gnd 0.147143f
C2196 plus.n83 gnd 0.774009f
C2197 plus.n84 gnd 1.15797f
C2198 plus.t3 gnd 0.040367f
C2199 plus.t4 gnd 0.007209f
C2200 plus.t1 gnd 0.007209f
C2201 plus.n85 gnd 0.023379f
C2202 plus.n86 gnd 0.18149f
C2203 plus.t2 gnd 0.007209f
C2204 plus.t0 gnd 0.007209f
C2205 plus.n87 gnd 0.023379f
C2206 plus.n88 gnd 0.136231f
C2207 plus.n89 gnd 2.97989f
C2208 CSoutput.n0 gnd 0.042211f
C2209 CSoutput.t202 gnd 0.27922f
C2210 CSoutput.n1 gnd 0.126082f
C2211 CSoutput.n2 gnd 0.042211f
C2212 CSoutput.t200 gnd 0.27922f
C2213 CSoutput.n3 gnd 0.033456f
C2214 CSoutput.n4 gnd 0.042211f
C2215 CSoutput.t193 gnd 0.27922f
C2216 CSoutput.n5 gnd 0.028849f
C2217 CSoutput.n6 gnd 0.042211f
C2218 CSoutput.t197 gnd 0.27922f
C2219 CSoutput.t207 gnd 0.27922f
C2220 CSoutput.n7 gnd 0.124708f
C2221 CSoutput.n8 gnd 0.042211f
C2222 CSoutput.t205 gnd 0.27922f
C2223 CSoutput.n9 gnd 0.027506f
C2224 CSoutput.n10 gnd 0.042211f
C2225 CSoutput.t194 gnd 0.27922f
C2226 CSoutput.t199 gnd 0.27922f
C2227 CSoutput.n11 gnd 0.124708f
C2228 CSoutput.n12 gnd 0.042211f
C2229 CSoutput.t204 gnd 0.27922f
C2230 CSoutput.n13 gnd 0.028849f
C2231 CSoutput.n14 gnd 0.042211f
C2232 CSoutput.t209 gnd 0.27922f
C2233 CSoutput.t196 gnd 0.27922f
C2234 CSoutput.n15 gnd 0.124708f
C2235 CSoutput.n16 gnd 0.042211f
C2236 CSoutput.t203 gnd 0.27922f
C2237 CSoutput.n17 gnd 0.030813f
C2238 CSoutput.t211 gnd 0.333675f
C2239 CSoutput.t201 gnd 0.27922f
C2240 CSoutput.n18 gnd 0.159203f
C2241 CSoutput.n19 gnd 0.154482f
C2242 CSoutput.n20 gnd 0.179218f
C2243 CSoutput.n21 gnd 0.042211f
C2244 CSoutput.n22 gnd 0.03523f
C2245 CSoutput.n23 gnd 0.124708f
C2246 CSoutput.n24 gnd 0.033961f
C2247 CSoutput.n25 gnd 0.033456f
C2248 CSoutput.n26 gnd 0.042211f
C2249 CSoutput.n27 gnd 0.042211f
C2250 CSoutput.n28 gnd 0.034959f
C2251 CSoutput.n29 gnd 0.029681f
C2252 CSoutput.n30 gnd 0.127484f
C2253 CSoutput.n31 gnd 0.03009f
C2254 CSoutput.n32 gnd 0.042211f
C2255 CSoutput.n33 gnd 0.042211f
C2256 CSoutput.n34 gnd 0.042211f
C2257 CSoutput.n35 gnd 0.034587f
C2258 CSoutput.n36 gnd 0.124708f
C2259 CSoutput.n37 gnd 0.033077f
C2260 CSoutput.n38 gnd 0.034339f
C2261 CSoutput.n39 gnd 0.042211f
C2262 CSoutput.n40 gnd 0.042211f
C2263 CSoutput.n41 gnd 0.035223f
C2264 CSoutput.n42 gnd 0.032194f
C2265 CSoutput.n43 gnd 0.124708f
C2266 CSoutput.n44 gnd 0.03301f
C2267 CSoutput.n45 gnd 0.042211f
C2268 CSoutput.n46 gnd 0.042211f
C2269 CSoutput.n47 gnd 0.042211f
C2270 CSoutput.n48 gnd 0.03301f
C2271 CSoutput.n49 gnd 0.124708f
C2272 CSoutput.n50 gnd 0.032194f
C2273 CSoutput.n51 gnd 0.035223f
C2274 CSoutput.n52 gnd 0.042211f
C2275 CSoutput.n53 gnd 0.042211f
C2276 CSoutput.n54 gnd 0.034339f
C2277 CSoutput.n55 gnd 0.033077f
C2278 CSoutput.n56 gnd 0.124708f
C2279 CSoutput.n57 gnd 0.034587f
C2280 CSoutput.n58 gnd 0.042211f
C2281 CSoutput.n59 gnd 0.042211f
C2282 CSoutput.n60 gnd 0.042211f
C2283 CSoutput.n61 gnd 0.03009f
C2284 CSoutput.n62 gnd 0.127484f
C2285 CSoutput.n63 gnd 0.029681f
C2286 CSoutput.t210 gnd 0.27922f
C2287 CSoutput.n64 gnd 0.124708f
C2288 CSoutput.n65 gnd 0.034959f
C2289 CSoutput.n66 gnd 0.042211f
C2290 CSoutput.n67 gnd 0.042211f
C2291 CSoutput.n68 gnd 0.042211f
C2292 CSoutput.n69 gnd 0.033961f
C2293 CSoutput.n70 gnd 0.124708f
C2294 CSoutput.n71 gnd 0.03523f
C2295 CSoutput.n72 gnd 0.030813f
C2296 CSoutput.n73 gnd 0.042211f
C2297 CSoutput.n74 gnd 0.042211f
C2298 CSoutput.n75 gnd 0.031955f
C2299 CSoutput.n76 gnd 0.018978f
C2300 CSoutput.t212 gnd 0.313724f
C2301 CSoutput.n77 gnd 0.155845f
C2302 CSoutput.n78 gnd 0.637555f
C2303 CSoutput.t143 gnd 0.052653f
C2304 CSoutput.t103 gnd 0.052653f
C2305 CSoutput.n79 gnd 0.407656f
C2306 CSoutput.t153 gnd 0.052653f
C2307 CSoutput.t117 gnd 0.052653f
C2308 CSoutput.n80 gnd 0.406929f
C2309 CSoutput.n81 gnd 0.413033f
C2310 CSoutput.t91 gnd 0.052653f
C2311 CSoutput.t127 gnd 0.052653f
C2312 CSoutput.n82 gnd 0.406929f
C2313 CSoutput.n83 gnd 0.203525f
C2314 CSoutput.t94 gnd 0.052653f
C2315 CSoutput.t111 gnd 0.052653f
C2316 CSoutput.n84 gnd 0.406929f
C2317 CSoutput.n85 gnd 0.203525f
C2318 CSoutput.t157 gnd 0.052653f
C2319 CSoutput.t123 gnd 0.052653f
C2320 CSoutput.n86 gnd 0.406929f
C2321 CSoutput.n87 gnd 0.203525f
C2322 CSoutput.t97 gnd 0.052653f
C2323 CSoutput.t146 gnd 0.052653f
C2324 CSoutput.n88 gnd 0.406929f
C2325 CSoutput.n89 gnd 0.373218f
C2326 CSoutput.t88 gnd 0.052653f
C2327 CSoutput.t141 gnd 0.052653f
C2328 CSoutput.n90 gnd 0.407656f
C2329 CSoutput.t133 gnd 0.052653f
C2330 CSoutput.t119 gnd 0.052653f
C2331 CSoutput.n91 gnd 0.406929f
C2332 CSoutput.n92 gnd 0.413033f
C2333 CSoutput.t104 gnd 0.052653f
C2334 CSoutput.t151 gnd 0.052653f
C2335 CSoutput.n93 gnd 0.406929f
C2336 CSoutput.n94 gnd 0.203525f
C2337 CSoutput.t132 gnd 0.052653f
C2338 CSoutput.t131 gnd 0.052653f
C2339 CSoutput.n95 gnd 0.406929f
C2340 CSoutput.n96 gnd 0.203525f
C2341 CSoutput.t124 gnd 0.052653f
C2342 CSoutput.t100 gnd 0.052653f
C2343 CSoutput.n97 gnd 0.406929f
C2344 CSoutput.n98 gnd 0.203525f
C2345 CSoutput.t90 gnd 0.052653f
C2346 CSoutput.t125 gnd 0.052653f
C2347 CSoutput.n99 gnd 0.406929f
C2348 CSoutput.n100 gnd 0.303507f
C2349 CSoutput.n101 gnd 0.382721f
C2350 CSoutput.t98 gnd 0.052653f
C2351 CSoutput.t150 gnd 0.052653f
C2352 CSoutput.n102 gnd 0.407656f
C2353 CSoutput.t138 gnd 0.052653f
C2354 CSoutput.t126 gnd 0.052653f
C2355 CSoutput.n103 gnd 0.406929f
C2356 CSoutput.n104 gnd 0.413033f
C2357 CSoutput.t113 gnd 0.052653f
C2358 CSoutput.t158 gnd 0.052653f
C2359 CSoutput.n105 gnd 0.406929f
C2360 CSoutput.n106 gnd 0.203525f
C2361 CSoutput.t137 gnd 0.052653f
C2362 CSoutput.t136 gnd 0.052653f
C2363 CSoutput.n107 gnd 0.406929f
C2364 CSoutput.n108 gnd 0.203525f
C2365 CSoutput.t129 gnd 0.052653f
C2366 CSoutput.t112 gnd 0.052653f
C2367 CSoutput.n109 gnd 0.406929f
C2368 CSoutput.n110 gnd 0.203525f
C2369 CSoutput.t99 gnd 0.052653f
C2370 CSoutput.t130 gnd 0.052653f
C2371 CSoutput.n111 gnd 0.406929f
C2372 CSoutput.n112 gnd 0.303507f
C2373 CSoutput.n113 gnd 0.427784f
C2374 CSoutput.n114 gnd 8.384171f
C2375 CSoutput.n116 gnd 0.746714f
C2376 CSoutput.n117 gnd 0.560036f
C2377 CSoutput.n118 gnd 0.746714f
C2378 CSoutput.n119 gnd 0.746714f
C2379 CSoutput.n120 gnd 2.01038f
C2380 CSoutput.n121 gnd 0.746714f
C2381 CSoutput.n122 gnd 0.746714f
C2382 CSoutput.t206 gnd 0.933393f
C2383 CSoutput.n123 gnd 0.746714f
C2384 CSoutput.n124 gnd 0.746714f
C2385 CSoutput.n128 gnd 0.746714f
C2386 CSoutput.n132 gnd 0.746714f
C2387 CSoutput.n133 gnd 0.746714f
C2388 CSoutput.n135 gnd 0.746714f
C2389 CSoutput.n140 gnd 0.746714f
C2390 CSoutput.n142 gnd 0.746714f
C2391 CSoutput.n143 gnd 0.746714f
C2392 CSoutput.n145 gnd 0.746714f
C2393 CSoutput.n146 gnd 0.746714f
C2394 CSoutput.n148 gnd 0.746714f
C2395 CSoutput.t195 gnd 12.4775f
C2396 CSoutput.n150 gnd 0.746714f
C2397 CSoutput.n151 gnd 0.560036f
C2398 CSoutput.n152 gnd 0.746714f
C2399 CSoutput.n153 gnd 0.746714f
C2400 CSoutput.n154 gnd 2.01038f
C2401 CSoutput.n155 gnd 0.746714f
C2402 CSoutput.n156 gnd 0.746714f
C2403 CSoutput.t213 gnd 0.933393f
C2404 CSoutput.n157 gnd 0.746714f
C2405 CSoutput.n158 gnd 0.746714f
C2406 CSoutput.n162 gnd 0.746714f
C2407 CSoutput.n166 gnd 0.746714f
C2408 CSoutput.n167 gnd 0.746714f
C2409 CSoutput.n169 gnd 0.746714f
C2410 CSoutput.n174 gnd 0.746714f
C2411 CSoutput.n176 gnd 0.746714f
C2412 CSoutput.n177 gnd 0.746714f
C2413 CSoutput.n179 gnd 0.746714f
C2414 CSoutput.n180 gnd 0.746714f
C2415 CSoutput.n182 gnd 0.746714f
C2416 CSoutput.n183 gnd 0.560036f
C2417 CSoutput.n185 gnd 0.746714f
C2418 CSoutput.n186 gnd 0.560036f
C2419 CSoutput.n187 gnd 0.746714f
C2420 CSoutput.n188 gnd 0.746714f
C2421 CSoutput.n189 gnd 2.01038f
C2422 CSoutput.n190 gnd 0.746714f
C2423 CSoutput.n191 gnd 0.746714f
C2424 CSoutput.t208 gnd 0.933393f
C2425 CSoutput.n192 gnd 0.746714f
C2426 CSoutput.n193 gnd 2.01038f
C2427 CSoutput.n195 gnd 0.746714f
C2428 CSoutput.n196 gnd 0.746714f
C2429 CSoutput.n198 gnd 0.746714f
C2430 CSoutput.n199 gnd 0.746714f
C2431 CSoutput.t192 gnd 12.2742f
C2432 CSoutput.t198 gnd 12.4775f
C2433 CSoutput.n205 gnd 2.34255f
C2434 CSoutput.n206 gnd 9.5427f
C2435 CSoutput.n207 gnd 9.942009f
C2436 CSoutput.n212 gnd 2.53761f
C2437 CSoutput.n218 gnd 0.746714f
C2438 CSoutput.n220 gnd 0.746714f
C2439 CSoutput.n222 gnd 0.746714f
C2440 CSoutput.n224 gnd 0.746714f
C2441 CSoutput.n226 gnd 0.746714f
C2442 CSoutput.n232 gnd 0.746714f
C2443 CSoutput.n239 gnd 1.36993f
C2444 CSoutput.n240 gnd 1.36993f
C2445 CSoutput.n241 gnd 0.746714f
C2446 CSoutput.n242 gnd 0.746714f
C2447 CSoutput.n244 gnd 0.560036f
C2448 CSoutput.n245 gnd 0.47962f
C2449 CSoutput.n247 gnd 0.560036f
C2450 CSoutput.n248 gnd 0.47962f
C2451 CSoutput.n249 gnd 0.560036f
C2452 CSoutput.n251 gnd 0.746714f
C2453 CSoutput.n253 gnd 2.01038f
C2454 CSoutput.n254 gnd 2.34255f
C2455 CSoutput.n255 gnd 8.77683f
C2456 CSoutput.n257 gnd 0.560036f
C2457 CSoutput.n258 gnd 1.44101f
C2458 CSoutput.n259 gnd 0.560036f
C2459 CSoutput.n261 gnd 0.746714f
C2460 CSoutput.n263 gnd 2.01038f
C2461 CSoutput.n264 gnd 4.37894f
C2462 CSoutput.t102 gnd 0.052653f
C2463 CSoutput.t142 gnd 0.052653f
C2464 CSoutput.n265 gnd 0.407656f
C2465 CSoutput.t116 gnd 0.052653f
C2466 CSoutput.t152 gnd 0.052653f
C2467 CSoutput.n266 gnd 0.406929f
C2468 CSoutput.n267 gnd 0.413033f
C2469 CSoutput.t139 gnd 0.052653f
C2470 CSoutput.t89 gnd 0.052653f
C2471 CSoutput.n268 gnd 0.406929f
C2472 CSoutput.n269 gnd 0.203525f
C2473 CSoutput.t110 gnd 0.052653f
C2474 CSoutput.t93 gnd 0.052653f
C2475 CSoutput.n270 gnd 0.406929f
C2476 CSoutput.n271 gnd 0.203525f
C2477 CSoutput.t122 gnd 0.052653f
C2478 CSoutput.t107 gnd 0.052653f
C2479 CSoutput.n272 gnd 0.406929f
C2480 CSoutput.n273 gnd 0.203525f
C2481 CSoutput.t145 gnd 0.052653f
C2482 CSoutput.t96 gnd 0.052653f
C2483 CSoutput.n274 gnd 0.406929f
C2484 CSoutput.n275 gnd 0.373218f
C2485 CSoutput.t121 gnd 0.052653f
C2486 CSoutput.t134 gnd 0.052653f
C2487 CSoutput.n276 gnd 0.407656f
C2488 CSoutput.t87 gnd 0.052653f
C2489 CSoutput.t108 gnd 0.052653f
C2490 CSoutput.n277 gnd 0.406929f
C2491 CSoutput.n278 gnd 0.413033f
C2492 CSoutput.t109 gnd 0.052653f
C2493 CSoutput.t149 gnd 0.052653f
C2494 CSoutput.n279 gnd 0.406929f
C2495 CSoutput.n280 gnd 0.203525f
C2496 CSoutput.t105 gnd 0.052653f
C2497 CSoutput.t106 gnd 0.052653f
C2498 CSoutput.n281 gnd 0.406929f
C2499 CSoutput.n282 gnd 0.203525f
C2500 CSoutput.t147 gnd 0.052653f
C2501 CSoutput.t148 gnd 0.052653f
C2502 CSoutput.n283 gnd 0.406929f
C2503 CSoutput.n284 gnd 0.203525f
C2504 CSoutput.t92 gnd 0.052653f
C2505 CSoutput.t135 gnd 0.052653f
C2506 CSoutput.n285 gnd 0.406929f
C2507 CSoutput.n286 gnd 0.303507f
C2508 CSoutput.n287 gnd 0.382721f
C2509 CSoutput.t128 gnd 0.052653f
C2510 CSoutput.t140 gnd 0.052653f
C2511 CSoutput.n288 gnd 0.407656f
C2512 CSoutput.t95 gnd 0.052653f
C2513 CSoutput.t118 gnd 0.052653f
C2514 CSoutput.n289 gnd 0.406929f
C2515 CSoutput.n290 gnd 0.413033f
C2516 CSoutput.t120 gnd 0.052653f
C2517 CSoutput.t156 gnd 0.052653f
C2518 CSoutput.n291 gnd 0.406929f
C2519 CSoutput.n292 gnd 0.203525f
C2520 CSoutput.t114 gnd 0.052653f
C2521 CSoutput.t115 gnd 0.052653f
C2522 CSoutput.n293 gnd 0.406929f
C2523 CSoutput.n294 gnd 0.203525f
C2524 CSoutput.t154 gnd 0.052653f
C2525 CSoutput.t155 gnd 0.052653f
C2526 CSoutput.n295 gnd 0.406929f
C2527 CSoutput.n296 gnd 0.203525f
C2528 CSoutput.t101 gnd 0.052653f
C2529 CSoutput.t144 gnd 0.052653f
C2530 CSoutput.n297 gnd 0.406928f
C2531 CSoutput.n298 gnd 0.303509f
C2532 CSoutput.n299 gnd 0.427784f
C2533 CSoutput.n300 gnd 11.741f
C2534 CSoutput.t191 gnd 0.046071f
C2535 CSoutput.t165 gnd 0.046071f
C2536 CSoutput.n301 gnd 0.408465f
C2537 CSoutput.t190 gnd 0.046071f
C2538 CSoutput.t28 gnd 0.046071f
C2539 CSoutput.n302 gnd 0.407102f
C2540 CSoutput.n303 gnd 0.379343f
C2541 CSoutput.t5 gnd 0.046071f
C2542 CSoutput.t17 gnd 0.046071f
C2543 CSoutput.n304 gnd 0.407102f
C2544 CSoutput.n305 gnd 0.186998f
C2545 CSoutput.t174 gnd 0.046071f
C2546 CSoutput.t166 gnd 0.046071f
C2547 CSoutput.n306 gnd 0.407102f
C2548 CSoutput.n307 gnd 0.186998f
C2549 CSoutput.t167 gnd 0.046071f
C2550 CSoutput.t178 gnd 0.046071f
C2551 CSoutput.n308 gnd 0.407102f
C2552 CSoutput.n309 gnd 0.186998f
C2553 CSoutput.t23 gnd 0.046071f
C2554 CSoutput.t84 gnd 0.046071f
C2555 CSoutput.n310 gnd 0.407102f
C2556 CSoutput.n311 gnd 0.186998f
C2557 CSoutput.t179 gnd 0.046071f
C2558 CSoutput.t82 gnd 0.046071f
C2559 CSoutput.n312 gnd 0.407102f
C2560 CSoutput.n313 gnd 0.186998f
C2561 CSoutput.t34 gnd 0.046071f
C2562 CSoutput.t186 gnd 0.046071f
C2563 CSoutput.n314 gnd 0.407102f
C2564 CSoutput.n315 gnd 0.186998f
C2565 CSoutput.t12 gnd 0.046071f
C2566 CSoutput.t176 gnd 0.046071f
C2567 CSoutput.n316 gnd 0.407102f
C2568 CSoutput.n317 gnd 0.186998f
C2569 CSoutput.t15 gnd 0.046071f
C2570 CSoutput.t161 gnd 0.046071f
C2571 CSoutput.n318 gnd 0.407102f
C2572 CSoutput.n319 gnd 0.344908f
C2573 CSoutput.t86 gnd 0.046071f
C2574 CSoutput.t183 gnd 0.046071f
C2575 CSoutput.n320 gnd 0.408465f
C2576 CSoutput.t170 gnd 0.046071f
C2577 CSoutput.t59 gnd 0.046071f
C2578 CSoutput.n321 gnd 0.407102f
C2579 CSoutput.n322 gnd 0.379343f
C2580 CSoutput.t75 gnd 0.046071f
C2581 CSoutput.t13 gnd 0.046071f
C2582 CSoutput.n323 gnd 0.407102f
C2583 CSoutput.n324 gnd 0.186998f
C2584 CSoutput.t189 gnd 0.046071f
C2585 CSoutput.t168 gnd 0.046071f
C2586 CSoutput.n325 gnd 0.407102f
C2587 CSoutput.n326 gnd 0.186998f
C2588 CSoutput.t24 gnd 0.046071f
C2589 CSoutput.t159 gnd 0.046071f
C2590 CSoutput.n327 gnd 0.407102f
C2591 CSoutput.n328 gnd 0.186998f
C2592 CSoutput.t80 gnd 0.046071f
C2593 CSoutput.t70 gnd 0.046071f
C2594 CSoutput.n329 gnd 0.407102f
C2595 CSoutput.n330 gnd 0.186998f
C2596 CSoutput.t67 gnd 0.046071f
C2597 CSoutput.t10 gnd 0.046071f
C2598 CSoutput.n331 gnd 0.407102f
C2599 CSoutput.n332 gnd 0.186998f
C2600 CSoutput.t163 gnd 0.046071f
C2601 CSoutput.t36 gnd 0.046071f
C2602 CSoutput.n333 gnd 0.407102f
C2603 CSoutput.n334 gnd 0.186998f
C2604 CSoutput.t160 gnd 0.046071f
C2605 CSoutput.t181 gnd 0.046071f
C2606 CSoutput.n335 gnd 0.407102f
C2607 CSoutput.n336 gnd 0.186998f
C2608 CSoutput.t33 gnd 0.046071f
C2609 CSoutput.t83 gnd 0.046071f
C2610 CSoutput.n337 gnd 0.407102f
C2611 CSoutput.n338 gnd 0.283904f
C2612 CSoutput.n339 gnd 0.358091f
C2613 CSoutput.t21 gnd 0.046071f
C2614 CSoutput.t73 gnd 0.046071f
C2615 CSoutput.n340 gnd 0.408465f
C2616 CSoutput.t173 gnd 0.046071f
C2617 CSoutput.t44 gnd 0.046071f
C2618 CSoutput.n341 gnd 0.407102f
C2619 CSoutput.n342 gnd 0.379343f
C2620 CSoutput.t50 gnd 0.046071f
C2621 CSoutput.t71 gnd 0.046071f
C2622 CSoutput.n343 gnd 0.407102f
C2623 CSoutput.n344 gnd 0.186998f
C2624 CSoutput.t79 gnd 0.046071f
C2625 CSoutput.t76 gnd 0.046071f
C2626 CSoutput.n345 gnd 0.407102f
C2627 CSoutput.n346 gnd 0.186998f
C2628 CSoutput.t18 gnd 0.046071f
C2629 CSoutput.t39 gnd 0.046071f
C2630 CSoutput.n347 gnd 0.407102f
C2631 CSoutput.n348 gnd 0.186998f
C2632 CSoutput.t52 gnd 0.046071f
C2633 CSoutput.t53 gnd 0.046071f
C2634 CSoutput.n349 gnd 0.407102f
C2635 CSoutput.n350 gnd 0.186998f
C2636 CSoutput.t184 gnd 0.046071f
C2637 CSoutput.t72 gnd 0.046071f
C2638 CSoutput.n351 gnd 0.407102f
C2639 CSoutput.n352 gnd 0.186998f
C2640 CSoutput.t54 gnd 0.046071f
C2641 CSoutput.t77 gnd 0.046071f
C2642 CSoutput.n353 gnd 0.407102f
C2643 CSoutput.n354 gnd 0.186998f
C2644 CSoutput.t49 gnd 0.046071f
C2645 CSoutput.t19 gnd 0.046071f
C2646 CSoutput.n355 gnd 0.407102f
C2647 CSoutput.n356 gnd 0.186998f
C2648 CSoutput.t30 gnd 0.046071f
C2649 CSoutput.t61 gnd 0.046071f
C2650 CSoutput.n357 gnd 0.407102f
C2651 CSoutput.n358 gnd 0.283904f
C2652 CSoutput.n359 gnd 0.384533f
C2653 CSoutput.n360 gnd 12.447599f
C2654 CSoutput.t43 gnd 0.046071f
C2655 CSoutput.t1 gnd 0.046071f
C2656 CSoutput.n361 gnd 0.408465f
C2657 CSoutput.t64 gnd 0.046071f
C2658 CSoutput.t22 gnd 0.046071f
C2659 CSoutput.n362 gnd 0.407102f
C2660 CSoutput.n363 gnd 0.379343f
C2661 CSoutput.t57 gnd 0.046071f
C2662 CSoutput.t7 gnd 0.046071f
C2663 CSoutput.n364 gnd 0.407102f
C2664 CSoutput.n365 gnd 0.186998f
C2665 CSoutput.t162 gnd 0.046071f
C2666 CSoutput.t14 gnd 0.046071f
C2667 CSoutput.n366 gnd 0.407102f
C2668 CSoutput.n367 gnd 0.186998f
C2669 CSoutput.t4 gnd 0.046071f
C2670 CSoutput.t85 gnd 0.046071f
C2671 CSoutput.n368 gnd 0.407102f
C2672 CSoutput.n369 gnd 0.186998f
C2673 CSoutput.t51 gnd 0.046071f
C2674 CSoutput.t38 gnd 0.046071f
C2675 CSoutput.n370 gnd 0.407102f
C2676 CSoutput.n371 gnd 0.186998f
C2677 CSoutput.t46 gnd 0.046071f
C2678 CSoutput.t16 gnd 0.046071f
C2679 CSoutput.n372 gnd 0.407102f
C2680 CSoutput.n373 gnd 0.186998f
C2681 CSoutput.t68 gnd 0.046071f
C2682 CSoutput.t172 gnd 0.046071f
C2683 CSoutput.n374 gnd 0.407102f
C2684 CSoutput.n375 gnd 0.186998f
C2685 CSoutput.t78 gnd 0.046071f
C2686 CSoutput.t81 gnd 0.046071f
C2687 CSoutput.n376 gnd 0.407102f
C2688 CSoutput.n377 gnd 0.186998f
C2689 CSoutput.t32 gnd 0.046071f
C2690 CSoutput.t6 gnd 0.046071f
C2691 CSoutput.n378 gnd 0.407102f
C2692 CSoutput.n379 gnd 0.344908f
C2693 CSoutput.t29 gnd 0.046071f
C2694 CSoutput.t31 gnd 0.046071f
C2695 CSoutput.n380 gnd 0.408465f
C2696 CSoutput.t3 gnd 0.046071f
C2697 CSoutput.t47 gnd 0.046071f
C2698 CSoutput.n381 gnd 0.407102f
C2699 CSoutput.n382 gnd 0.379343f
C2700 CSoutput.t41 gnd 0.046071f
C2701 CSoutput.t42 gnd 0.046071f
C2702 CSoutput.n383 gnd 0.407102f
C2703 CSoutput.n384 gnd 0.186998f
C2704 CSoutput.t35 gnd 0.046071f
C2705 CSoutput.t69 gnd 0.046071f
C2706 CSoutput.n385 gnd 0.407102f
C2707 CSoutput.n386 gnd 0.186998f
C2708 CSoutput.t56 gnd 0.046071f
C2709 CSoutput.t74 gnd 0.046071f
C2710 CSoutput.n387 gnd 0.407102f
C2711 CSoutput.n388 gnd 0.186998f
C2712 CSoutput.t66 gnd 0.046071f
C2713 CSoutput.t177 gnd 0.046071f
C2714 CSoutput.n389 gnd 0.407102f
C2715 CSoutput.n390 gnd 0.186998f
C2716 CSoutput.t25 gnd 0.046071f
C2717 CSoutput.t187 gnd 0.046071f
C2718 CSoutput.n391 gnd 0.407102f
C2719 CSoutput.n392 gnd 0.186998f
C2720 CSoutput.t175 gnd 0.046071f
C2721 CSoutput.t26 gnd 0.046071f
C2722 CSoutput.n393 gnd 0.407102f
C2723 CSoutput.n394 gnd 0.186998f
C2724 CSoutput.t63 gnd 0.046071f
C2725 CSoutput.t164 gnd 0.046071f
C2726 CSoutput.n395 gnd 0.407102f
C2727 CSoutput.n396 gnd 0.186998f
C2728 CSoutput.t188 gnd 0.046071f
C2729 CSoutput.t48 gnd 0.046071f
C2730 CSoutput.n397 gnd 0.407102f
C2731 CSoutput.n398 gnd 0.283904f
C2732 CSoutput.n399 gnd 0.358091f
C2733 CSoutput.t55 gnd 0.046071f
C2734 CSoutput.t182 gnd 0.046071f
C2735 CSoutput.n400 gnd 0.408465f
C2736 CSoutput.t171 gnd 0.046071f
C2737 CSoutput.t8 gnd 0.046071f
C2738 CSoutput.n401 gnd 0.407102f
C2739 CSoutput.n402 gnd 0.379343f
C2740 CSoutput.t62 gnd 0.046071f
C2741 CSoutput.t11 gnd 0.046071f
C2742 CSoutput.n403 gnd 0.407102f
C2743 CSoutput.n404 gnd 0.186998f
C2744 CSoutput.t58 gnd 0.046071f
C2745 CSoutput.t0 gnd 0.046071f
C2746 CSoutput.n405 gnd 0.407102f
C2747 CSoutput.n406 gnd 0.186998f
C2748 CSoutput.t45 gnd 0.046071f
C2749 CSoutput.t60 gnd 0.046071f
C2750 CSoutput.n407 gnd 0.407102f
C2751 CSoutput.n408 gnd 0.186998f
C2752 CSoutput.t169 gnd 0.046071f
C2753 CSoutput.t185 gnd 0.046071f
C2754 CSoutput.n409 gnd 0.407102f
C2755 CSoutput.n410 gnd 0.186998f
C2756 CSoutput.t9 gnd 0.046071f
C2757 CSoutput.t65 gnd 0.046071f
C2758 CSoutput.n411 gnd 0.407102f
C2759 CSoutput.n412 gnd 0.186998f
C2760 CSoutput.t2 gnd 0.046071f
C2761 CSoutput.t27 gnd 0.046071f
C2762 CSoutput.n413 gnd 0.407102f
C2763 CSoutput.n414 gnd 0.186998f
C2764 CSoutput.t180 gnd 0.046071f
C2765 CSoutput.t37 gnd 0.046071f
C2766 CSoutput.n415 gnd 0.407102f
C2767 CSoutput.n416 gnd 0.186998f
C2768 CSoutput.t20 gnd 0.046071f
C2769 CSoutput.t40 gnd 0.046071f
C2770 CSoutput.n417 gnd 0.407102f
C2771 CSoutput.n418 gnd 0.283904f
C2772 CSoutput.n419 gnd 0.384533f
C2773 CSoutput.n420 gnd 7.34439f
C2774 CSoutput.n421 gnd 12.9754f
C2775 vdd.t28 gnd 0.034663f
C2776 vdd.t121 gnd 0.034663f
C2777 vdd.n0 gnd 0.273395f
C2778 vdd.t137 gnd 0.034663f
C2779 vdd.t117 gnd 0.034663f
C2780 vdd.n1 gnd 0.272944f
C2781 vdd.n2 gnd 0.251706f
C2782 vdd.t113 gnd 0.034663f
C2783 vdd.t109 gnd 0.034663f
C2784 vdd.n3 gnd 0.272944f
C2785 vdd.n4 gnd 0.127297f
C2786 vdd.t111 gnd 0.034663f
C2787 vdd.t12 gnd 0.034663f
C2788 vdd.n5 gnd 0.272944f
C2789 vdd.n6 gnd 0.119445f
C2790 vdd.t235 gnd 0.034663f
C2791 vdd.t23 gnd 0.034663f
C2792 vdd.n7 gnd 0.273395f
C2793 vdd.t14 gnd 0.034663f
C2794 vdd.t26 gnd 0.034663f
C2795 vdd.n8 gnd 0.272944f
C2796 vdd.n9 gnd 0.251706f
C2797 vdd.t119 gnd 0.034663f
C2798 vdd.t115 gnd 0.034663f
C2799 vdd.n10 gnd 0.272944f
C2800 vdd.n11 gnd 0.127297f
C2801 vdd.t30 gnd 0.034663f
C2802 vdd.t8 gnd 0.034663f
C2803 vdd.n12 gnd 0.272944f
C2804 vdd.n13 gnd 0.119445f
C2805 vdd.n14 gnd 0.084445f
C2806 vdd.t127 gnd 0.019257f
C2807 vdd.t135 gnd 0.019257f
C2808 vdd.n15 gnd 0.177256f
C2809 vdd.t133 gnd 0.019257f
C2810 vdd.t125 gnd 0.019257f
C2811 vdd.n16 gnd 0.176737f
C2812 vdd.n17 gnd 0.307578f
C2813 vdd.t123 gnd 0.019257f
C2814 vdd.t4 gnd 0.019257f
C2815 vdd.n18 gnd 0.176737f
C2816 vdd.n19 gnd 0.127249f
C2817 vdd.t134 gnd 0.019257f
C2818 vdd.t126 gnd 0.019257f
C2819 vdd.n20 gnd 0.177256f
C2820 vdd.t128 gnd 0.019257f
C2821 vdd.t122 gnd 0.019257f
C2822 vdd.n21 gnd 0.176737f
C2823 vdd.n22 gnd 0.307578f
C2824 vdd.t132 gnd 0.019257f
C2825 vdd.t129 gnd 0.019257f
C2826 vdd.n23 gnd 0.176737f
C2827 vdd.n24 gnd 0.127249f
C2828 vdd.t124 gnd 0.019257f
C2829 vdd.t5 gnd 0.019257f
C2830 vdd.n25 gnd 0.176737f
C2831 vdd.t130 gnd 0.019257f
C2832 vdd.t131 gnd 0.019257f
C2833 vdd.n26 gnd 0.176737f
C2834 vdd.n27 gnd 19.5887f
C2835 vdd.n28 gnd 7.57335f
C2836 vdd.n29 gnd 0.005252f
C2837 vdd.n30 gnd 0.004874f
C2838 vdd.n31 gnd 0.002696f
C2839 vdd.n32 gnd 0.00619f
C2840 vdd.n33 gnd 0.002619f
C2841 vdd.n34 gnd 0.002773f
C2842 vdd.n35 gnd 0.004874f
C2843 vdd.n36 gnd 0.002619f
C2844 vdd.n37 gnd 0.00619f
C2845 vdd.n38 gnd 0.002773f
C2846 vdd.n39 gnd 0.004874f
C2847 vdd.n40 gnd 0.002619f
C2848 vdd.n41 gnd 0.004643f
C2849 vdd.n42 gnd 0.004657f
C2850 vdd.t167 gnd 0.0133f
C2851 vdd.n43 gnd 0.029591f
C2852 vdd.n44 gnd 0.153999f
C2853 vdd.n45 gnd 0.002619f
C2854 vdd.n46 gnd 0.002773f
C2855 vdd.n47 gnd 0.00619f
C2856 vdd.n48 gnd 0.00619f
C2857 vdd.n49 gnd 0.002773f
C2858 vdd.n50 gnd 0.002619f
C2859 vdd.n51 gnd 0.004874f
C2860 vdd.n52 gnd 0.004874f
C2861 vdd.n53 gnd 0.002619f
C2862 vdd.n54 gnd 0.002773f
C2863 vdd.n55 gnd 0.00619f
C2864 vdd.n56 gnd 0.00619f
C2865 vdd.n57 gnd 0.002773f
C2866 vdd.n58 gnd 0.002619f
C2867 vdd.n59 gnd 0.004874f
C2868 vdd.n60 gnd 0.004874f
C2869 vdd.n61 gnd 0.002619f
C2870 vdd.n62 gnd 0.002773f
C2871 vdd.n63 gnd 0.00619f
C2872 vdd.n64 gnd 0.00619f
C2873 vdd.n65 gnd 0.014635f
C2874 vdd.n66 gnd 0.002696f
C2875 vdd.n67 gnd 0.002619f
C2876 vdd.n68 gnd 0.012597f
C2877 vdd.n69 gnd 0.008795f
C2878 vdd.t217 gnd 0.030812f
C2879 vdd.t189 gnd 0.030812f
C2880 vdd.n70 gnd 0.21176f
C2881 vdd.n71 gnd 0.166517f
C2882 vdd.t227 gnd 0.030812f
C2883 vdd.t215 gnd 0.030812f
C2884 vdd.n72 gnd 0.21176f
C2885 vdd.n73 gnd 0.134378f
C2886 vdd.t147 gnd 0.030812f
C2887 vdd.t180 gnd 0.030812f
C2888 vdd.n74 gnd 0.21176f
C2889 vdd.n75 gnd 0.134378f
C2890 vdd.t155 gnd 0.030812f
C2891 vdd.t195 gnd 0.030812f
C2892 vdd.n76 gnd 0.21176f
C2893 vdd.n77 gnd 0.134378f
C2894 vdd.t175 gnd 0.030812f
C2895 vdd.t220 gnd 0.030812f
C2896 vdd.n78 gnd 0.21176f
C2897 vdd.n79 gnd 0.134378f
C2898 vdd.n80 gnd 0.005252f
C2899 vdd.n81 gnd 0.004874f
C2900 vdd.n82 gnd 0.002696f
C2901 vdd.n83 gnd 0.00619f
C2902 vdd.n84 gnd 0.002619f
C2903 vdd.n85 gnd 0.002773f
C2904 vdd.n86 gnd 0.004874f
C2905 vdd.n87 gnd 0.002619f
C2906 vdd.n88 gnd 0.00619f
C2907 vdd.n89 gnd 0.002773f
C2908 vdd.n90 gnd 0.004874f
C2909 vdd.n91 gnd 0.002619f
C2910 vdd.n92 gnd 0.004643f
C2911 vdd.n93 gnd 0.004657f
C2912 vdd.t160 gnd 0.0133f
C2913 vdd.n94 gnd 0.029591f
C2914 vdd.n95 gnd 0.153999f
C2915 vdd.n96 gnd 0.002619f
C2916 vdd.n97 gnd 0.002773f
C2917 vdd.n98 gnd 0.00619f
C2918 vdd.n99 gnd 0.00619f
C2919 vdd.n100 gnd 0.002773f
C2920 vdd.n101 gnd 0.002619f
C2921 vdd.n102 gnd 0.004874f
C2922 vdd.n103 gnd 0.004874f
C2923 vdd.n104 gnd 0.002619f
C2924 vdd.n105 gnd 0.002773f
C2925 vdd.n106 gnd 0.00619f
C2926 vdd.n107 gnd 0.00619f
C2927 vdd.n108 gnd 0.002773f
C2928 vdd.n109 gnd 0.002619f
C2929 vdd.n110 gnd 0.004874f
C2930 vdd.n111 gnd 0.004874f
C2931 vdd.n112 gnd 0.002619f
C2932 vdd.n113 gnd 0.002773f
C2933 vdd.n114 gnd 0.00619f
C2934 vdd.n115 gnd 0.00619f
C2935 vdd.n116 gnd 0.014635f
C2936 vdd.n117 gnd 0.002696f
C2937 vdd.n118 gnd 0.002619f
C2938 vdd.n119 gnd 0.012597f
C2939 vdd.n120 gnd 0.008519f
C2940 vdd.n121 gnd 0.099978f
C2941 vdd.n122 gnd 0.005252f
C2942 vdd.n123 gnd 0.004874f
C2943 vdd.n124 gnd 0.002696f
C2944 vdd.n125 gnd 0.00619f
C2945 vdd.n126 gnd 0.002619f
C2946 vdd.n127 gnd 0.002773f
C2947 vdd.n128 gnd 0.004874f
C2948 vdd.n129 gnd 0.002619f
C2949 vdd.n130 gnd 0.00619f
C2950 vdd.n131 gnd 0.002773f
C2951 vdd.n132 gnd 0.004874f
C2952 vdd.n133 gnd 0.002619f
C2953 vdd.n134 gnd 0.004643f
C2954 vdd.n135 gnd 0.004657f
C2955 vdd.t193 gnd 0.0133f
C2956 vdd.n136 gnd 0.029591f
C2957 vdd.n137 gnd 0.153999f
C2958 vdd.n138 gnd 0.002619f
C2959 vdd.n139 gnd 0.002773f
C2960 vdd.n140 gnd 0.00619f
C2961 vdd.n141 gnd 0.00619f
C2962 vdd.n142 gnd 0.002773f
C2963 vdd.n143 gnd 0.002619f
C2964 vdd.n144 gnd 0.004874f
C2965 vdd.n145 gnd 0.004874f
C2966 vdd.n146 gnd 0.002619f
C2967 vdd.n147 gnd 0.002773f
C2968 vdd.n148 gnd 0.00619f
C2969 vdd.n149 gnd 0.00619f
C2970 vdd.n150 gnd 0.002773f
C2971 vdd.n151 gnd 0.002619f
C2972 vdd.n152 gnd 0.004874f
C2973 vdd.n153 gnd 0.004874f
C2974 vdd.n154 gnd 0.002619f
C2975 vdd.n155 gnd 0.002773f
C2976 vdd.n156 gnd 0.00619f
C2977 vdd.n157 gnd 0.00619f
C2978 vdd.n158 gnd 0.014635f
C2979 vdd.n159 gnd 0.002696f
C2980 vdd.n160 gnd 0.002619f
C2981 vdd.n161 gnd 0.012597f
C2982 vdd.n162 gnd 0.008795f
C2983 vdd.t209 gnd 0.030812f
C2984 vdd.t139 gnd 0.030812f
C2985 vdd.n163 gnd 0.21176f
C2986 vdd.n164 gnd 0.166517f
C2987 vdd.t177 gnd 0.030812f
C2988 vdd.t179 gnd 0.030812f
C2989 vdd.n165 gnd 0.21176f
C2990 vdd.n166 gnd 0.134378f
C2991 vdd.t224 gnd 0.030812f
C2992 vdd.t172 gnd 0.030812f
C2993 vdd.n167 gnd 0.21176f
C2994 vdd.n168 gnd 0.134378f
C2995 vdd.t173 gnd 0.030812f
C2996 vdd.t222 gnd 0.030812f
C2997 vdd.n169 gnd 0.21176f
C2998 vdd.n170 gnd 0.134378f
C2999 vdd.t223 gnd 0.030812f
C3000 vdd.t153 gnd 0.030812f
C3001 vdd.n171 gnd 0.21176f
C3002 vdd.n172 gnd 0.134378f
C3003 vdd.n173 gnd 0.005252f
C3004 vdd.n174 gnd 0.004874f
C3005 vdd.n175 gnd 0.002696f
C3006 vdd.n176 gnd 0.00619f
C3007 vdd.n177 gnd 0.002619f
C3008 vdd.n178 gnd 0.002773f
C3009 vdd.n179 gnd 0.004874f
C3010 vdd.n180 gnd 0.002619f
C3011 vdd.n181 gnd 0.00619f
C3012 vdd.n182 gnd 0.002773f
C3013 vdd.n183 gnd 0.004874f
C3014 vdd.n184 gnd 0.002619f
C3015 vdd.n185 gnd 0.004643f
C3016 vdd.n186 gnd 0.004657f
C3017 vdd.t210 gnd 0.0133f
C3018 vdd.n187 gnd 0.029591f
C3019 vdd.n188 gnd 0.153999f
C3020 vdd.n189 gnd 0.002619f
C3021 vdd.n190 gnd 0.002773f
C3022 vdd.n191 gnd 0.00619f
C3023 vdd.n192 gnd 0.00619f
C3024 vdd.n193 gnd 0.002773f
C3025 vdd.n194 gnd 0.002619f
C3026 vdd.n195 gnd 0.004874f
C3027 vdd.n196 gnd 0.004874f
C3028 vdd.n197 gnd 0.002619f
C3029 vdd.n198 gnd 0.002773f
C3030 vdd.n199 gnd 0.00619f
C3031 vdd.n200 gnd 0.00619f
C3032 vdd.n201 gnd 0.002773f
C3033 vdd.n202 gnd 0.002619f
C3034 vdd.n203 gnd 0.004874f
C3035 vdd.n204 gnd 0.004874f
C3036 vdd.n205 gnd 0.002619f
C3037 vdd.n206 gnd 0.002773f
C3038 vdd.n207 gnd 0.00619f
C3039 vdd.n208 gnd 0.00619f
C3040 vdd.n209 gnd 0.014635f
C3041 vdd.n210 gnd 0.002696f
C3042 vdd.n211 gnd 0.002619f
C3043 vdd.n212 gnd 0.012597f
C3044 vdd.n213 gnd 0.008519f
C3045 vdd.n214 gnd 0.059477f
C3046 vdd.n215 gnd 0.214311f
C3047 vdd.n216 gnd 0.005252f
C3048 vdd.n217 gnd 0.004874f
C3049 vdd.n218 gnd 0.002696f
C3050 vdd.n219 gnd 0.00619f
C3051 vdd.n220 gnd 0.002619f
C3052 vdd.n221 gnd 0.002773f
C3053 vdd.n222 gnd 0.004874f
C3054 vdd.n223 gnd 0.002619f
C3055 vdd.n224 gnd 0.00619f
C3056 vdd.n225 gnd 0.002773f
C3057 vdd.n226 gnd 0.004874f
C3058 vdd.n227 gnd 0.002619f
C3059 vdd.n228 gnd 0.004643f
C3060 vdd.n229 gnd 0.004657f
C3061 vdd.t201 gnd 0.0133f
C3062 vdd.n230 gnd 0.029591f
C3063 vdd.n231 gnd 0.153999f
C3064 vdd.n232 gnd 0.002619f
C3065 vdd.n233 gnd 0.002773f
C3066 vdd.n234 gnd 0.00619f
C3067 vdd.n235 gnd 0.00619f
C3068 vdd.n236 gnd 0.002773f
C3069 vdd.n237 gnd 0.002619f
C3070 vdd.n238 gnd 0.004874f
C3071 vdd.n239 gnd 0.004874f
C3072 vdd.n240 gnd 0.002619f
C3073 vdd.n241 gnd 0.002773f
C3074 vdd.n242 gnd 0.00619f
C3075 vdd.n243 gnd 0.00619f
C3076 vdd.n244 gnd 0.002773f
C3077 vdd.n245 gnd 0.002619f
C3078 vdd.n246 gnd 0.004874f
C3079 vdd.n247 gnd 0.004874f
C3080 vdd.n248 gnd 0.002619f
C3081 vdd.n249 gnd 0.002773f
C3082 vdd.n250 gnd 0.00619f
C3083 vdd.n251 gnd 0.00619f
C3084 vdd.n252 gnd 0.014635f
C3085 vdd.n253 gnd 0.002696f
C3086 vdd.n254 gnd 0.002619f
C3087 vdd.n255 gnd 0.012597f
C3088 vdd.n256 gnd 0.008795f
C3089 vdd.t212 gnd 0.030812f
C3090 vdd.t158 gnd 0.030812f
C3091 vdd.n257 gnd 0.21176f
C3092 vdd.n258 gnd 0.166517f
C3093 vdd.t190 gnd 0.030812f
C3094 vdd.t192 gnd 0.030812f
C3095 vdd.n259 gnd 0.21176f
C3096 vdd.n260 gnd 0.134378f
C3097 vdd.t231 gnd 0.030812f
C3098 vdd.t187 gnd 0.030812f
C3099 vdd.n261 gnd 0.21176f
C3100 vdd.n262 gnd 0.134378f
C3101 vdd.t188 gnd 0.030812f
C3102 vdd.t229 gnd 0.030812f
C3103 vdd.n263 gnd 0.21176f
C3104 vdd.n264 gnd 0.134378f
C3105 vdd.t230 gnd 0.030812f
C3106 vdd.t165 gnd 0.030812f
C3107 vdd.n265 gnd 0.21176f
C3108 vdd.n266 gnd 0.134378f
C3109 vdd.n267 gnd 0.005252f
C3110 vdd.n268 gnd 0.004874f
C3111 vdd.n269 gnd 0.002696f
C3112 vdd.n270 gnd 0.00619f
C3113 vdd.n271 gnd 0.002619f
C3114 vdd.n272 gnd 0.002773f
C3115 vdd.n273 gnd 0.004874f
C3116 vdd.n274 gnd 0.002619f
C3117 vdd.n275 gnd 0.00619f
C3118 vdd.n276 gnd 0.002773f
C3119 vdd.n277 gnd 0.004874f
C3120 vdd.n278 gnd 0.002619f
C3121 vdd.n279 gnd 0.004643f
C3122 vdd.n280 gnd 0.004657f
C3123 vdd.t219 gnd 0.0133f
C3124 vdd.n281 gnd 0.029591f
C3125 vdd.n282 gnd 0.153999f
C3126 vdd.n283 gnd 0.002619f
C3127 vdd.n284 gnd 0.002773f
C3128 vdd.n285 gnd 0.00619f
C3129 vdd.n286 gnd 0.00619f
C3130 vdd.n287 gnd 0.002773f
C3131 vdd.n288 gnd 0.002619f
C3132 vdd.n289 gnd 0.004874f
C3133 vdd.n290 gnd 0.004874f
C3134 vdd.n291 gnd 0.002619f
C3135 vdd.n292 gnd 0.002773f
C3136 vdd.n293 gnd 0.00619f
C3137 vdd.n294 gnd 0.00619f
C3138 vdd.n295 gnd 0.002773f
C3139 vdd.n296 gnd 0.002619f
C3140 vdd.n297 gnd 0.004874f
C3141 vdd.n298 gnd 0.004874f
C3142 vdd.n299 gnd 0.002619f
C3143 vdd.n300 gnd 0.002773f
C3144 vdd.n301 gnd 0.00619f
C3145 vdd.n302 gnd 0.00619f
C3146 vdd.n303 gnd 0.014635f
C3147 vdd.n304 gnd 0.002696f
C3148 vdd.n305 gnd 0.002619f
C3149 vdd.n306 gnd 0.012597f
C3150 vdd.n307 gnd 0.008519f
C3151 vdd.n308 gnd 0.059477f
C3152 vdd.n309 gnd 0.235534f
C3153 vdd.n310 gnd 0.009537f
C3154 vdd.n311 gnd 0.009537f
C3155 vdd.n312 gnd 0.007703f
C3156 vdd.n313 gnd 0.007703f
C3157 vdd.n314 gnd 0.00957f
C3158 vdd.n315 gnd 0.00957f
C3159 vdd.t146 gnd 0.489021f
C3160 vdd.n316 gnd 0.00957f
C3161 vdd.n317 gnd 0.00957f
C3162 vdd.n318 gnd 0.00957f
C3163 vdd.t154 gnd 0.489021f
C3164 vdd.n319 gnd 0.00957f
C3165 vdd.n320 gnd 0.00957f
C3166 vdd.n321 gnd 0.00957f
C3167 vdd.n322 gnd 0.00957f
C3168 vdd.n323 gnd 0.007703f
C3169 vdd.n324 gnd 0.00957f
C3170 vdd.n325 gnd 0.787324f
C3171 vdd.n326 gnd 0.00957f
C3172 vdd.n327 gnd 0.00957f
C3173 vdd.n328 gnd 0.00957f
C3174 vdd.n329 gnd 0.669959f
C3175 vdd.n330 gnd 0.00957f
C3176 vdd.n331 gnd 0.00957f
C3177 vdd.n332 gnd 0.00957f
C3178 vdd.n333 gnd 0.00957f
C3179 vdd.n334 gnd 0.00957f
C3180 vdd.n335 gnd 0.007703f
C3181 vdd.n336 gnd 0.00957f
C3182 vdd.t152 gnd 0.489021f
C3183 vdd.n337 gnd 0.00957f
C3184 vdd.n338 gnd 0.00957f
C3185 vdd.n339 gnd 0.00957f
C3186 vdd.n340 gnd 0.978042f
C3187 vdd.n341 gnd 0.00957f
C3188 vdd.n342 gnd 0.00957f
C3189 vdd.n343 gnd 0.00957f
C3190 vdd.n344 gnd 0.00957f
C3191 vdd.n345 gnd 0.00957f
C3192 vdd.n346 gnd 0.007703f
C3193 vdd.n347 gnd 0.00957f
C3194 vdd.n348 gnd 0.00957f
C3195 vdd.n349 gnd 0.00957f
C3196 vdd.n350 gnd 0.022553f
C3197 vdd.n351 gnd 2.2495f
C3198 vdd.n352 gnd 0.022906f
C3199 vdd.n353 gnd 0.00957f
C3200 vdd.n354 gnd 0.00957f
C3201 vdd.n356 gnd 0.00957f
C3202 vdd.n357 gnd 0.00957f
C3203 vdd.n358 gnd 0.007703f
C3204 vdd.n359 gnd 0.007703f
C3205 vdd.n360 gnd 0.00957f
C3206 vdd.n361 gnd 0.00957f
C3207 vdd.n362 gnd 0.00957f
C3208 vdd.n363 gnd 0.00957f
C3209 vdd.n364 gnd 0.00957f
C3210 vdd.n365 gnd 0.00957f
C3211 vdd.n366 gnd 0.007703f
C3212 vdd.n368 gnd 0.00957f
C3213 vdd.n369 gnd 0.00957f
C3214 vdd.n370 gnd 0.00957f
C3215 vdd.n371 gnd 0.00957f
C3216 vdd.n372 gnd 0.00957f
C3217 vdd.n373 gnd 0.007703f
C3218 vdd.n375 gnd 0.00957f
C3219 vdd.n376 gnd 0.00957f
C3220 vdd.n377 gnd 0.00957f
C3221 vdd.n378 gnd 0.00957f
C3222 vdd.n379 gnd 0.00957f
C3223 vdd.n380 gnd 0.007703f
C3224 vdd.n382 gnd 0.00957f
C3225 vdd.n383 gnd 0.00957f
C3226 vdd.n384 gnd 0.00957f
C3227 vdd.n385 gnd 0.00957f
C3228 vdd.n386 gnd 0.006432f
C3229 vdd.t106 gnd 0.11774f
C3230 vdd.t105 gnd 0.125832f
C3231 vdd.t104 gnd 0.153767f
C3232 vdd.n387 gnd 0.197108f
C3233 vdd.n388 gnd 0.166376f
C3234 vdd.n390 gnd 0.00957f
C3235 vdd.n391 gnd 0.00957f
C3236 vdd.n392 gnd 0.007703f
C3237 vdd.n393 gnd 0.00957f
C3238 vdd.n395 gnd 0.00957f
C3239 vdd.n396 gnd 0.00957f
C3240 vdd.n397 gnd 0.00957f
C3241 vdd.n398 gnd 0.00957f
C3242 vdd.n399 gnd 0.007703f
C3243 vdd.n401 gnd 0.00957f
C3244 vdd.n402 gnd 0.00957f
C3245 vdd.n403 gnd 0.00957f
C3246 vdd.n404 gnd 0.00957f
C3247 vdd.n405 gnd 0.00957f
C3248 vdd.n406 gnd 0.007703f
C3249 vdd.n408 gnd 0.00957f
C3250 vdd.n409 gnd 0.00957f
C3251 vdd.n410 gnd 0.00957f
C3252 vdd.n411 gnd 0.00957f
C3253 vdd.n412 gnd 0.00957f
C3254 vdd.n413 gnd 0.007703f
C3255 vdd.n415 gnd 0.00957f
C3256 vdd.n416 gnd 0.00957f
C3257 vdd.n417 gnd 0.00957f
C3258 vdd.n418 gnd 0.00957f
C3259 vdd.n419 gnd 0.00957f
C3260 vdd.n420 gnd 0.007703f
C3261 vdd.n422 gnd 0.00957f
C3262 vdd.n423 gnd 0.00957f
C3263 vdd.n424 gnd 0.00957f
C3264 vdd.n425 gnd 0.00957f
C3265 vdd.n426 gnd 0.007626f
C3266 vdd.t100 gnd 0.11774f
C3267 vdd.t99 gnd 0.125832f
C3268 vdd.t98 gnd 0.153767f
C3269 vdd.n427 gnd 0.197108f
C3270 vdd.n428 gnd 0.166376f
C3271 vdd.n430 gnd 0.00957f
C3272 vdd.n431 gnd 0.00957f
C3273 vdd.n432 gnd 0.007703f
C3274 vdd.n433 gnd 0.00957f
C3275 vdd.n435 gnd 0.00957f
C3276 vdd.n436 gnd 0.00957f
C3277 vdd.n437 gnd 0.00957f
C3278 vdd.n438 gnd 0.00957f
C3279 vdd.n439 gnd 0.007703f
C3280 vdd.n441 gnd 0.00957f
C3281 vdd.n442 gnd 0.00957f
C3282 vdd.n443 gnd 0.00957f
C3283 vdd.n444 gnd 0.00957f
C3284 vdd.n445 gnd 0.00957f
C3285 vdd.n446 gnd 0.007703f
C3286 vdd.n448 gnd 0.00957f
C3287 vdd.n449 gnd 0.00957f
C3288 vdd.n450 gnd 0.00957f
C3289 vdd.n451 gnd 0.00957f
C3290 vdd.n452 gnd 0.00957f
C3291 vdd.n453 gnd 0.007703f
C3292 vdd.n455 gnd 0.00957f
C3293 vdd.n456 gnd 0.00957f
C3294 vdd.n457 gnd 0.00957f
C3295 vdd.n458 gnd 0.00957f
C3296 vdd.n459 gnd 0.00957f
C3297 vdd.n460 gnd 0.007703f
C3298 vdd.n462 gnd 0.00957f
C3299 vdd.n463 gnd 0.00957f
C3300 vdd.n464 gnd 0.00957f
C3301 vdd.n465 gnd 0.00957f
C3302 vdd.n466 gnd 0.00957f
C3303 vdd.n467 gnd 0.00957f
C3304 vdd.n468 gnd 0.007703f
C3305 vdd.n469 gnd 0.00957f
C3306 vdd.n470 gnd 0.00957f
C3307 vdd.n471 gnd 0.007703f
C3308 vdd.n472 gnd 0.00957f
C3309 vdd.n473 gnd 0.00957f
C3310 vdd.n474 gnd 0.007703f
C3311 vdd.n475 gnd 0.00957f
C3312 vdd.n476 gnd 0.007703f
C3313 vdd.n477 gnd 0.00957f
C3314 vdd.n478 gnd 0.007703f
C3315 vdd.n479 gnd 0.00957f
C3316 vdd.n480 gnd 0.00957f
C3317 vdd.t178 gnd 0.489021f
C3318 vdd.n481 gnd 0.523253f
C3319 vdd.n482 gnd 0.00957f
C3320 vdd.n483 gnd 0.007703f
C3321 vdd.n484 gnd 0.00957f
C3322 vdd.n485 gnd 0.007703f
C3323 vdd.n486 gnd 0.00957f
C3324 vdd.t176 gnd 0.489021f
C3325 vdd.n487 gnd 0.00957f
C3326 vdd.n488 gnd 0.007703f
C3327 vdd.n489 gnd 0.00957f
C3328 vdd.n490 gnd 0.007703f
C3329 vdd.n491 gnd 0.00957f
C3330 vdd.n492 gnd 0.767763f
C3331 vdd.n493 gnd 0.811775f
C3332 vdd.t138 gnd 0.489021f
C3333 vdd.n494 gnd 0.00957f
C3334 vdd.n495 gnd 0.007703f
C3335 vdd.n496 gnd 0.00957f
C3336 vdd.n497 gnd 0.007703f
C3337 vdd.n498 gnd 0.00957f
C3338 vdd.n499 gnd 0.601496f
C3339 vdd.n500 gnd 0.00957f
C3340 vdd.n501 gnd 0.007703f
C3341 vdd.n502 gnd 0.00957f
C3342 vdd.n503 gnd 0.007703f
C3343 vdd.n504 gnd 0.00957f
C3344 vdd.n505 gnd 0.978042f
C3345 vdd.t166 gnd 0.489021f
C3346 vdd.n506 gnd 0.00957f
C3347 vdd.n507 gnd 0.007703f
C3348 vdd.n508 gnd 0.00957f
C3349 vdd.n509 gnd 0.007703f
C3350 vdd.n510 gnd 0.00957f
C3351 vdd.n511 gnd 0.523253f
C3352 vdd.n512 gnd 0.00957f
C3353 vdd.n513 gnd 0.007703f
C3354 vdd.n514 gnd 0.022906f
C3355 vdd.n515 gnd 0.022906f
C3356 vdd.n516 gnd 8.62633f
C3357 vdd.t40 gnd 0.489021f
C3358 vdd.n517 gnd 0.022906f
C3359 vdd.n518 gnd 0.00823f
C3360 vdd.n519 gnd 0.007703f
C3361 vdd.n524 gnd 0.006125f
C3362 vdd.n525 gnd 0.007703f
C3363 vdd.n526 gnd 0.00957f
C3364 vdd.n527 gnd 0.00957f
C3365 vdd.n528 gnd 0.00957f
C3366 vdd.n529 gnd 0.00957f
C3367 vdd.n530 gnd 0.00957f
C3368 vdd.n531 gnd 0.007703f
C3369 vdd.n532 gnd 0.00957f
C3370 vdd.n533 gnd 0.00957f
C3371 vdd.n534 gnd 0.00957f
C3372 vdd.n535 gnd 0.00957f
C3373 vdd.n536 gnd 0.00957f
C3374 vdd.n537 gnd 0.007703f
C3375 vdd.n538 gnd 0.00957f
C3376 vdd.n539 gnd 0.00957f
C3377 vdd.n540 gnd 0.00957f
C3378 vdd.n541 gnd 0.00957f
C3379 vdd.n542 gnd 0.00957f
C3380 vdd.t69 gnd 0.11774f
C3381 vdd.t70 gnd 0.125832f
C3382 vdd.t68 gnd 0.153767f
C3383 vdd.n543 gnd 0.197108f
C3384 vdd.n544 gnd 0.165606f
C3385 vdd.n545 gnd 0.015714f
C3386 vdd.n546 gnd 0.00957f
C3387 vdd.n547 gnd 0.00957f
C3388 vdd.n548 gnd 0.00957f
C3389 vdd.n549 gnd 0.00957f
C3390 vdd.n550 gnd 0.00957f
C3391 vdd.n551 gnd 0.007703f
C3392 vdd.n552 gnd 0.00957f
C3393 vdd.n553 gnd 0.00957f
C3394 vdd.n554 gnd 0.00957f
C3395 vdd.n555 gnd 0.00957f
C3396 vdd.n556 gnd 0.00957f
C3397 vdd.n557 gnd 0.007703f
C3398 vdd.n558 gnd 0.00957f
C3399 vdd.n559 gnd 0.00957f
C3400 vdd.n560 gnd 0.00957f
C3401 vdd.n561 gnd 0.00957f
C3402 vdd.n562 gnd 0.00957f
C3403 vdd.n563 gnd 0.007703f
C3404 vdd.n564 gnd 0.00957f
C3405 vdd.n565 gnd 0.00957f
C3406 vdd.n566 gnd 0.00957f
C3407 vdd.n567 gnd 0.00957f
C3408 vdd.n568 gnd 0.00957f
C3409 vdd.n569 gnd 0.007703f
C3410 vdd.n570 gnd 0.00957f
C3411 vdd.n571 gnd 0.00957f
C3412 vdd.n572 gnd 0.00957f
C3413 vdd.n573 gnd 0.00957f
C3414 vdd.n574 gnd 0.00957f
C3415 vdd.n575 gnd 0.007703f
C3416 vdd.n576 gnd 0.00957f
C3417 vdd.n577 gnd 0.00957f
C3418 vdd.n578 gnd 0.00957f
C3419 vdd.n579 gnd 0.007626f
C3420 vdd.t56 gnd 0.11774f
C3421 vdd.t57 gnd 0.125832f
C3422 vdd.t55 gnd 0.153767f
C3423 vdd.n580 gnd 0.197108f
C3424 vdd.n581 gnd 0.165606f
C3425 vdd.n582 gnd 0.00957f
C3426 vdd.n583 gnd 0.007703f
C3427 vdd.n585 gnd 0.00957f
C3428 vdd.n587 gnd 0.00957f
C3429 vdd.n588 gnd 0.00957f
C3430 vdd.n589 gnd 0.007703f
C3431 vdd.n590 gnd 0.00957f
C3432 vdd.n591 gnd 0.00957f
C3433 vdd.n592 gnd 0.00957f
C3434 vdd.n593 gnd 0.00957f
C3435 vdd.n594 gnd 0.00957f
C3436 vdd.n595 gnd 0.007703f
C3437 vdd.n596 gnd 0.00957f
C3438 vdd.n597 gnd 0.00957f
C3439 vdd.n598 gnd 0.00957f
C3440 vdd.n599 gnd 0.00957f
C3441 vdd.n600 gnd 0.00957f
C3442 vdd.n601 gnd 0.007703f
C3443 vdd.n602 gnd 0.00957f
C3444 vdd.n603 gnd 0.00957f
C3445 vdd.n604 gnd 0.00957f
C3446 vdd.n605 gnd 0.006125f
C3447 vdd.n610 gnd 0.006508f
C3448 vdd.n611 gnd 0.006508f
C3449 vdd.n612 gnd 0.006508f
C3450 vdd.n613 gnd 8.3427f
C3451 vdd.n614 gnd 0.006508f
C3452 vdd.n615 gnd 0.006508f
C3453 vdd.n616 gnd 0.006508f
C3454 vdd.n618 gnd 0.006508f
C3455 vdd.n619 gnd 0.006508f
C3456 vdd.n621 gnd 0.006508f
C3457 vdd.n622 gnd 0.004737f
C3458 vdd.n624 gnd 0.006508f
C3459 vdd.t34 gnd 0.26298f
C3460 vdd.t33 gnd 0.269193f
C3461 vdd.t31 gnd 0.171684f
C3462 vdd.n625 gnd 0.092785f
C3463 vdd.n626 gnd 0.052631f
C3464 vdd.n627 gnd 0.009301f
C3465 vdd.n628 gnd 0.015064f
C3466 vdd.n630 gnd 0.006508f
C3467 vdd.n631 gnd 0.665069f
C3468 vdd.n632 gnd 0.014255f
C3469 vdd.n633 gnd 0.014255f
C3470 vdd.n634 gnd 0.006508f
C3471 vdd.n635 gnd 0.015221f
C3472 vdd.n636 gnd 0.006508f
C3473 vdd.n637 gnd 0.006508f
C3474 vdd.n638 gnd 0.006508f
C3475 vdd.n639 gnd 0.006508f
C3476 vdd.n640 gnd 0.006508f
C3477 vdd.n642 gnd 0.006508f
C3478 vdd.n643 gnd 0.006508f
C3479 vdd.n645 gnd 0.006508f
C3480 vdd.n646 gnd 0.006508f
C3481 vdd.n648 gnd 0.006508f
C3482 vdd.n649 gnd 0.006508f
C3483 vdd.n651 gnd 0.006508f
C3484 vdd.n652 gnd 0.006508f
C3485 vdd.n654 gnd 0.006508f
C3486 vdd.n655 gnd 0.006508f
C3487 vdd.n657 gnd 0.006508f
C3488 vdd.n658 gnd 0.004737f
C3489 vdd.n660 gnd 0.006508f
C3490 vdd.t103 gnd 0.26298f
C3491 vdd.t102 gnd 0.269193f
C3492 vdd.t101 gnd 0.171684f
C3493 vdd.n661 gnd 0.092785f
C3494 vdd.n662 gnd 0.052631f
C3495 vdd.n663 gnd 0.009301f
C3496 vdd.n664 gnd 0.006508f
C3497 vdd.n665 gnd 0.006508f
C3498 vdd.t32 gnd 0.332534f
C3499 vdd.n666 gnd 0.006508f
C3500 vdd.n667 gnd 0.006508f
C3501 vdd.n668 gnd 0.006508f
C3502 vdd.n669 gnd 0.006508f
C3503 vdd.n670 gnd 0.006508f
C3504 vdd.n671 gnd 0.665069f
C3505 vdd.n672 gnd 0.006508f
C3506 vdd.n673 gnd 0.006508f
C3507 vdd.n674 gnd 0.562374f
C3508 vdd.n675 gnd 0.006508f
C3509 vdd.n676 gnd 0.006508f
C3510 vdd.n677 gnd 0.006508f
C3511 vdd.n678 gnd 0.006508f
C3512 vdd.n679 gnd 0.650398f
C3513 vdd.n680 gnd 0.006508f
C3514 vdd.n681 gnd 0.006508f
C3515 vdd.n682 gnd 0.006508f
C3516 vdd.n683 gnd 0.006508f
C3517 vdd.n684 gnd 0.006508f
C3518 vdd.n685 gnd 0.665069f
C3519 vdd.n686 gnd 0.006508f
C3520 vdd.n687 gnd 0.006508f
C3521 vdd.t16 gnd 0.332534f
C3522 vdd.n688 gnd 0.006508f
C3523 vdd.n689 gnd 0.006508f
C3524 vdd.n690 gnd 0.006508f
C3525 vdd.t17 gnd 0.332534f
C3526 vdd.n691 gnd 0.006508f
C3527 vdd.n692 gnd 0.006508f
C3528 vdd.n693 gnd 0.006508f
C3529 vdd.n694 gnd 0.006508f
C3530 vdd.n695 gnd 0.006508f
C3531 vdd.t65 gnd 0.278742f
C3532 vdd.n696 gnd 0.006508f
C3533 vdd.n697 gnd 0.006508f
C3534 vdd.n698 gnd 0.533033f
C3535 vdd.n699 gnd 0.006508f
C3536 vdd.t66 gnd 0.269193f
C3537 vdd.t64 gnd 0.171684f
C3538 vdd.t67 gnd 0.269193f
C3539 vdd.n700 gnd 0.151297f
C3540 vdd.n701 gnd 0.006508f
C3541 vdd.n702 gnd 0.006508f
C3542 vdd.n703 gnd 0.425448f
C3543 vdd.n704 gnd 0.006508f
C3544 vdd.n705 gnd 0.006508f
C3545 vdd.t20 gnd 0.097804f
C3546 vdd.n706 gnd 0.386327f
C3547 vdd.n707 gnd 0.006508f
C3548 vdd.n708 gnd 0.006508f
C3549 vdd.n709 gnd 0.006508f
C3550 vdd.n710 gnd 0.572155f
C3551 vdd.n711 gnd 0.006508f
C3552 vdd.n712 gnd 0.006508f
C3553 vdd.t0 gnd 0.332534f
C3554 vdd.n713 gnd 0.006508f
C3555 vdd.n714 gnd 0.006508f
C3556 vdd.n715 gnd 0.006508f
C3557 vdd.t22 gnd 0.332534f
C3558 vdd.n716 gnd 0.006508f
C3559 vdd.n717 gnd 0.006508f
C3560 vdd.t19 gnd 0.332534f
C3561 vdd.n718 gnd 0.006508f
C3562 vdd.n719 gnd 0.006508f
C3563 vdd.n720 gnd 0.006508f
C3564 vdd.t9 gnd 0.264071f
C3565 vdd.n721 gnd 0.006508f
C3566 vdd.n722 gnd 0.006508f
C3567 vdd.n723 gnd 0.547704f
C3568 vdd.n724 gnd 0.006508f
C3569 vdd.n725 gnd 0.006508f
C3570 vdd.n726 gnd 0.006508f
C3571 vdd.t2 gnd 0.332534f
C3572 vdd.n727 gnd 0.006508f
C3573 vdd.n728 gnd 0.006508f
C3574 vdd.t234 gnd 0.278742f
C3575 vdd.n729 gnd 0.400997f
C3576 vdd.n730 gnd 0.006508f
C3577 vdd.n731 gnd 0.006508f
C3578 vdd.n732 gnd 0.006508f
C3579 vdd.n733 gnd 0.347205f
C3580 vdd.n734 gnd 0.006508f
C3581 vdd.n735 gnd 0.006508f
C3582 vdd.t25 gnd 0.332534f
C3583 vdd.n736 gnd 0.006508f
C3584 vdd.n737 gnd 0.006508f
C3585 vdd.n738 gnd 0.006508f
C3586 vdd.n739 gnd 0.665069f
C3587 vdd.n740 gnd 0.006508f
C3588 vdd.n741 gnd 0.006508f
C3589 vdd.t10 gnd 0.22495f
C3590 vdd.t13 gnd 0.317864f
C3591 vdd.n742 gnd 0.006508f
C3592 vdd.n743 gnd 0.006508f
C3593 vdd.n744 gnd 0.006508f
C3594 vdd.n745 gnd 0.498801f
C3595 vdd.n746 gnd 0.006508f
C3596 vdd.n747 gnd 0.006508f
C3597 vdd.n748 gnd 0.006508f
C3598 vdd.n749 gnd 0.006508f
C3599 vdd.n750 gnd 0.006508f
C3600 vdd.t82 gnd 0.332534f
C3601 vdd.n751 gnd 0.006508f
C3602 vdd.n752 gnd 0.006508f
C3603 vdd.t114 gnd 0.332534f
C3604 vdd.n753 gnd 0.006508f
C3605 vdd.n754 gnd 0.014255f
C3606 vdd.n755 gnd 0.014255f
C3607 vdd.n756 gnd 0.792214f
C3608 vdd.n757 gnd 0.006508f
C3609 vdd.n758 gnd 0.006508f
C3610 vdd.t118 gnd 0.332534f
C3611 vdd.n759 gnd 0.014255f
C3612 vdd.n760 gnd 0.006508f
C3613 vdd.n761 gnd 0.006508f
C3614 vdd.t110 gnd 0.606386f
C3615 vdd.n779 gnd 0.015221f
C3616 vdd.n797 gnd 0.014255f
C3617 vdd.n798 gnd 0.006508f
C3618 vdd.n799 gnd 0.014255f
C3619 vdd.t97 gnd 0.26298f
C3620 vdd.t96 gnd 0.269193f
C3621 vdd.t95 gnd 0.171684f
C3622 vdd.n800 gnd 0.092785f
C3623 vdd.n801 gnd 0.052631f
C3624 vdd.n802 gnd 0.015064f
C3625 vdd.n803 gnd 0.006508f
C3626 vdd.n804 gnd 0.352095f
C3627 vdd.n805 gnd 0.014255f
C3628 vdd.n806 gnd 0.006508f
C3629 vdd.n807 gnd 0.015221f
C3630 vdd.n808 gnd 0.006508f
C3631 vdd.t80 gnd 0.26298f
C3632 vdd.t79 gnd 0.269193f
C3633 vdd.t77 gnd 0.171684f
C3634 vdd.n809 gnd 0.092785f
C3635 vdd.n810 gnd 0.052631f
C3636 vdd.n811 gnd 0.009301f
C3637 vdd.n812 gnd 0.006508f
C3638 vdd.n813 gnd 0.006508f
C3639 vdd.t78 gnd 0.332534f
C3640 vdd.n814 gnd 0.006508f
C3641 vdd.t108 gnd 0.332534f
C3642 vdd.n815 gnd 0.006508f
C3643 vdd.n816 gnd 0.006508f
C3644 vdd.n817 gnd 0.006508f
C3645 vdd.n818 gnd 0.006508f
C3646 vdd.n819 gnd 0.006508f
C3647 vdd.n820 gnd 0.665069f
C3648 vdd.n821 gnd 0.006508f
C3649 vdd.n822 gnd 0.006508f
C3650 vdd.t112 gnd 0.332534f
C3651 vdd.n823 gnd 0.006508f
C3652 vdd.n824 gnd 0.006508f
C3653 vdd.n825 gnd 0.006508f
C3654 vdd.n826 gnd 0.006508f
C3655 vdd.n827 gnd 0.440119f
C3656 vdd.n828 gnd 0.006508f
C3657 vdd.n829 gnd 0.006508f
C3658 vdd.n830 gnd 0.006508f
C3659 vdd.n831 gnd 0.006508f
C3660 vdd.n832 gnd 0.006508f
C3661 vdd.n833 gnd 0.586825f
C3662 vdd.n834 gnd 0.006508f
C3663 vdd.n835 gnd 0.006508f
C3664 vdd.t116 gnd 0.317864f
C3665 vdd.t21 gnd 0.22495f
C3666 vdd.n836 gnd 0.006508f
C3667 vdd.n837 gnd 0.006508f
C3668 vdd.n838 gnd 0.006508f
C3669 vdd.t15 gnd 0.332534f
C3670 vdd.n839 gnd 0.006508f
C3671 vdd.n840 gnd 0.006508f
C3672 vdd.t136 gnd 0.332534f
C3673 vdd.n841 gnd 0.006508f
C3674 vdd.n842 gnd 0.006508f
C3675 vdd.n843 gnd 0.006508f
C3676 vdd.t120 gnd 0.278742f
C3677 vdd.n844 gnd 0.006508f
C3678 vdd.n845 gnd 0.006508f
C3679 vdd.n846 gnd 0.533033f
C3680 vdd.n847 gnd 0.006508f
C3681 vdd.n848 gnd 0.006508f
C3682 vdd.n849 gnd 0.006508f
C3683 vdd.t27 gnd 0.332534f
C3684 vdd.n850 gnd 0.006508f
C3685 vdd.n851 gnd 0.006508f
C3686 vdd.t3 gnd 0.264071f
C3687 vdd.n852 gnd 0.386327f
C3688 vdd.n853 gnd 0.006508f
C3689 vdd.n854 gnd 0.006508f
C3690 vdd.n855 gnd 0.006508f
C3691 vdd.n856 gnd 0.572155f
C3692 vdd.n857 gnd 0.006508f
C3693 vdd.n858 gnd 0.006508f
C3694 vdd.t107 gnd 0.332534f
C3695 vdd.n859 gnd 0.006508f
C3696 vdd.n860 gnd 0.006508f
C3697 vdd.n861 gnd 0.006508f
C3698 vdd.n862 gnd 0.665069f
C3699 vdd.n863 gnd 0.006508f
C3700 vdd.n864 gnd 0.006508f
C3701 vdd.t1 gnd 0.332534f
C3702 vdd.n865 gnd 0.006508f
C3703 vdd.n866 gnd 0.006508f
C3704 vdd.n867 gnd 0.006508f
C3705 vdd.t24 gnd 0.097804f
C3706 vdd.n868 gnd 0.006508f
C3707 vdd.n869 gnd 0.006508f
C3708 vdd.n870 gnd 0.006508f
C3709 vdd.t87 gnd 0.269193f
C3710 vdd.t85 gnd 0.171684f
C3711 vdd.t88 gnd 0.269193f
C3712 vdd.n871 gnd 0.151297f
C3713 vdd.n872 gnd 0.006508f
C3714 vdd.n873 gnd 0.006508f
C3715 vdd.t18 gnd 0.332534f
C3716 vdd.n874 gnd 0.006508f
C3717 vdd.n875 gnd 0.006508f
C3718 vdd.t86 gnd 0.278742f
C3719 vdd.n876 gnd 0.567264f
C3720 vdd.n877 gnd 0.006508f
C3721 vdd.n878 gnd 0.006508f
C3722 vdd.n879 gnd 0.006508f
C3723 vdd.n880 gnd 0.347205f
C3724 vdd.n881 gnd 0.006508f
C3725 vdd.n882 gnd 0.006508f
C3726 vdd.n883 gnd 0.46457f
C3727 vdd.n884 gnd 0.006508f
C3728 vdd.n885 gnd 0.006508f
C3729 vdd.n886 gnd 0.006508f
C3730 vdd.n887 gnd 0.665069f
C3731 vdd.n888 gnd 0.006508f
C3732 vdd.n889 gnd 0.006508f
C3733 vdd.t6 gnd 0.332534f
C3734 vdd.n890 gnd 0.006508f
C3735 vdd.n891 gnd 0.006508f
C3736 vdd.n892 gnd 0.006508f
C3737 vdd.n893 gnd 0.665069f
C3738 vdd.n894 gnd 0.006508f
C3739 vdd.n895 gnd 0.006508f
C3740 vdd.n896 gnd 0.006508f
C3741 vdd.n897 gnd 0.006508f
C3742 vdd.n898 gnd 0.006508f
C3743 vdd.t36 gnd 0.332534f
C3744 vdd.n899 gnd 0.006508f
C3745 vdd.n900 gnd 0.006508f
C3746 vdd.n901 gnd 0.006508f
C3747 vdd.n902 gnd 0.014255f
C3748 vdd.n903 gnd 0.014255f
C3749 vdd.n904 gnd 0.93892f
C3750 vdd.n905 gnd 0.006508f
C3751 vdd.n906 gnd 0.006508f
C3752 vdd.n907 gnd 0.435229f
C3753 vdd.n908 gnd 0.014255f
C3754 vdd.n909 gnd 0.006508f
C3755 vdd.n910 gnd 0.006508f
C3756 vdd.n911 gnd 8.62633f
C3757 vdd.n944 gnd 0.015221f
C3758 vdd.n945 gnd 0.006508f
C3759 vdd.n946 gnd 0.006508f
C3760 vdd.n947 gnd 0.006508f
C3761 vdd.n948 gnd 0.006125f
C3762 vdd.n951 gnd 0.022906f
C3763 vdd.n952 gnd 0.006393f
C3764 vdd.n953 gnd 0.007703f
C3765 vdd.n955 gnd 0.00957f
C3766 vdd.n956 gnd 0.00957f
C3767 vdd.n957 gnd 0.007703f
C3768 vdd.n959 gnd 0.00957f
C3769 vdd.n960 gnd 0.00957f
C3770 vdd.n961 gnd 0.00957f
C3771 vdd.n962 gnd 0.00957f
C3772 vdd.n963 gnd 0.00957f
C3773 vdd.n964 gnd 0.007703f
C3774 vdd.n966 gnd 0.00957f
C3775 vdd.n967 gnd 0.00957f
C3776 vdd.n968 gnd 0.00957f
C3777 vdd.n969 gnd 0.00957f
C3778 vdd.n970 gnd 0.00957f
C3779 vdd.n971 gnd 0.007703f
C3780 vdd.n973 gnd 0.00957f
C3781 vdd.n974 gnd 0.00957f
C3782 vdd.n975 gnd 0.00957f
C3783 vdd.n976 gnd 0.00957f
C3784 vdd.n977 gnd 0.006432f
C3785 vdd.t94 gnd 0.11774f
C3786 vdd.t93 gnd 0.125832f
C3787 vdd.t92 gnd 0.153767f
C3788 vdd.n978 gnd 0.197108f
C3789 vdd.n979 gnd 0.165606f
C3790 vdd.n981 gnd 0.00957f
C3791 vdd.n982 gnd 0.00957f
C3792 vdd.n983 gnd 0.007703f
C3793 vdd.n984 gnd 0.00957f
C3794 vdd.n986 gnd 0.00957f
C3795 vdd.n987 gnd 0.00957f
C3796 vdd.n988 gnd 0.00957f
C3797 vdd.n989 gnd 0.00957f
C3798 vdd.n990 gnd 0.007703f
C3799 vdd.n992 gnd 0.00957f
C3800 vdd.n993 gnd 0.00957f
C3801 vdd.n994 gnd 0.00957f
C3802 vdd.n995 gnd 0.00957f
C3803 vdd.n996 gnd 0.00957f
C3804 vdd.n997 gnd 0.007703f
C3805 vdd.n999 gnd 0.00957f
C3806 vdd.n1000 gnd 0.00957f
C3807 vdd.n1001 gnd 0.00957f
C3808 vdd.n1002 gnd 0.00957f
C3809 vdd.n1003 gnd 0.00957f
C3810 vdd.n1004 gnd 0.007703f
C3811 vdd.n1006 gnd 0.00957f
C3812 vdd.n1007 gnd 0.00957f
C3813 vdd.n1008 gnd 0.00957f
C3814 vdd.n1009 gnd 0.00957f
C3815 vdd.n1010 gnd 0.00957f
C3816 vdd.n1011 gnd 0.007703f
C3817 vdd.n1013 gnd 0.00957f
C3818 vdd.n1014 gnd 0.00957f
C3819 vdd.n1015 gnd 0.00957f
C3820 vdd.n1016 gnd 0.00957f
C3821 vdd.n1017 gnd 0.007626f
C3822 vdd.t76 gnd 0.11774f
C3823 vdd.t75 gnd 0.125832f
C3824 vdd.t74 gnd 0.153767f
C3825 vdd.n1018 gnd 0.197108f
C3826 vdd.n1019 gnd 0.165606f
C3827 vdd.n1021 gnd 0.00957f
C3828 vdd.n1022 gnd 0.00957f
C3829 vdd.n1023 gnd 0.007703f
C3830 vdd.n1024 gnd 0.00957f
C3831 vdd.n1026 gnd 0.00957f
C3832 vdd.n1027 gnd 0.00957f
C3833 vdd.n1028 gnd 0.00957f
C3834 vdd.n1029 gnd 0.00957f
C3835 vdd.n1030 gnd 0.007703f
C3836 vdd.n1032 gnd 0.00957f
C3837 vdd.n1033 gnd 0.00957f
C3838 vdd.n1034 gnd 0.00957f
C3839 vdd.n1035 gnd 0.00957f
C3840 vdd.n1036 gnd 0.00957f
C3841 vdd.n1037 gnd 0.007703f
C3842 vdd.n1039 gnd 0.00957f
C3843 vdd.n1040 gnd 0.00957f
C3844 vdd.n1041 gnd 0.00957f
C3845 vdd.n1042 gnd 0.00957f
C3846 vdd.n1043 gnd 0.00957f
C3847 vdd.n1044 gnd 0.007703f
C3848 vdd.n1046 gnd 0.00957f
C3849 vdd.n1047 gnd 0.00957f
C3850 vdd.n1048 gnd 0.006125f
C3851 vdd.n1049 gnd 0.007703f
C3852 vdd.n1050 gnd 0.006508f
C3853 vdd.n1051 gnd 0.006508f
C3854 vdd.n1052 gnd 0.006508f
C3855 vdd.n1053 gnd 0.006508f
C3856 vdd.n1054 gnd 0.006508f
C3857 vdd.n1055 gnd 0.006508f
C3858 vdd.n1056 gnd 0.006508f
C3859 vdd.n1057 gnd 0.006508f
C3860 vdd.n1058 gnd 0.006508f
C3861 vdd.n1059 gnd 0.006508f
C3862 vdd.n1060 gnd 0.006508f
C3863 vdd.n1061 gnd 0.006508f
C3864 vdd.n1062 gnd 0.006508f
C3865 vdd.n1063 gnd 0.006508f
C3866 vdd.n1064 gnd 0.006508f
C3867 vdd.n1065 gnd 0.006508f
C3868 vdd.n1066 gnd 0.006508f
C3869 vdd.n1067 gnd 0.006508f
C3870 vdd.n1068 gnd 0.006508f
C3871 vdd.n1069 gnd 0.006508f
C3872 vdd.n1070 gnd 0.006508f
C3873 vdd.n1071 gnd 0.006508f
C3874 vdd.n1072 gnd 0.006508f
C3875 vdd.n1073 gnd 0.006508f
C3876 vdd.n1074 gnd 0.006508f
C3877 vdd.n1075 gnd 0.006508f
C3878 vdd.n1076 gnd 0.006508f
C3879 vdd.n1077 gnd 0.006508f
C3880 vdd.n1078 gnd 0.006508f
C3881 vdd.n1079 gnd 0.006508f
C3882 vdd.n1080 gnd 0.006508f
C3883 vdd.t37 gnd 0.26298f
C3884 vdd.t38 gnd 0.269193f
C3885 vdd.t35 gnd 0.171684f
C3886 vdd.n1081 gnd 0.092785f
C3887 vdd.n1082 gnd 0.052631f
C3888 vdd.n1083 gnd 0.009301f
C3889 vdd.n1084 gnd 0.006508f
C3890 vdd.n1085 gnd 0.006508f
C3891 vdd.n1086 gnd 0.006508f
C3892 vdd.n1087 gnd 0.006508f
C3893 vdd.n1088 gnd 0.006508f
C3894 vdd.n1089 gnd 0.006508f
C3895 vdd.n1090 gnd 0.006508f
C3896 vdd.n1091 gnd 0.006508f
C3897 vdd.n1092 gnd 0.006508f
C3898 vdd.n1093 gnd 0.006508f
C3899 vdd.n1094 gnd 0.006508f
C3900 vdd.n1095 gnd 0.006508f
C3901 vdd.n1096 gnd 0.006508f
C3902 vdd.n1097 gnd 0.006508f
C3903 vdd.n1098 gnd 0.006508f
C3904 vdd.n1099 gnd 0.006508f
C3905 vdd.n1100 gnd 0.006508f
C3906 vdd.t62 gnd 0.26298f
C3907 vdd.t63 gnd 0.269193f
C3908 vdd.t61 gnd 0.171684f
C3909 vdd.n1101 gnd 0.092785f
C3910 vdd.n1102 gnd 0.052631f
C3911 vdd.n1103 gnd 0.006508f
C3912 vdd.n1104 gnd 0.006508f
C3913 vdd.n1105 gnd 0.006508f
C3914 vdd.n1106 gnd 0.006508f
C3915 vdd.n1107 gnd 0.006508f
C3916 vdd.n1108 gnd 0.006508f
C3917 vdd.n1109 gnd 0.006508f
C3918 vdd.n1110 gnd 0.006508f
C3919 vdd.n1111 gnd 0.006508f
C3920 vdd.n1112 gnd 0.006508f
C3921 vdd.n1113 gnd 0.006508f
C3922 vdd.n1114 gnd 0.006508f
C3923 vdd.n1115 gnd 0.006508f
C3924 vdd.n1116 gnd 0.006508f
C3925 vdd.n1117 gnd 0.006508f
C3926 vdd.n1118 gnd 0.006508f
C3927 vdd.n1119 gnd 0.006508f
C3928 vdd.n1120 gnd 0.006508f
C3929 vdd.n1121 gnd 0.006508f
C3930 vdd.n1122 gnd 0.006508f
C3931 vdd.n1123 gnd 0.006508f
C3932 vdd.n1124 gnd 0.006508f
C3933 vdd.n1125 gnd 0.006508f
C3934 vdd.n1126 gnd 0.006508f
C3935 vdd.n1127 gnd 0.006508f
C3936 vdd.n1128 gnd 0.006508f
C3937 vdd.n1129 gnd 0.004737f
C3938 vdd.n1130 gnd 0.009301f
C3939 vdd.n1131 gnd 0.005024f
C3940 vdd.n1132 gnd 0.006508f
C3941 vdd.n1133 gnd 0.006508f
C3942 vdd.n1134 gnd 0.006508f
C3943 vdd.n1135 gnd 0.015221f
C3944 vdd.n1136 gnd 0.015221f
C3945 vdd.n1137 gnd 0.014255f
C3946 vdd.n1138 gnd 0.014255f
C3947 vdd.n1139 gnd 0.006508f
C3948 vdd.n1140 gnd 0.006508f
C3949 vdd.n1141 gnd 0.006508f
C3950 vdd.n1142 gnd 0.006508f
C3951 vdd.n1143 gnd 0.006508f
C3952 vdd.n1144 gnd 0.006508f
C3953 vdd.n1145 gnd 0.006508f
C3954 vdd.n1146 gnd 0.006508f
C3955 vdd.n1147 gnd 0.006508f
C3956 vdd.n1148 gnd 0.006508f
C3957 vdd.n1149 gnd 0.006508f
C3958 vdd.n1150 gnd 0.006508f
C3959 vdd.n1151 gnd 0.006508f
C3960 vdd.n1152 gnd 0.006508f
C3961 vdd.n1153 gnd 0.006508f
C3962 vdd.n1154 gnd 0.006508f
C3963 vdd.n1155 gnd 0.006508f
C3964 vdd.n1156 gnd 0.006508f
C3965 vdd.n1157 gnd 0.006508f
C3966 vdd.n1158 gnd 0.006508f
C3967 vdd.n1159 gnd 0.006508f
C3968 vdd.n1160 gnd 0.006508f
C3969 vdd.n1161 gnd 0.006508f
C3970 vdd.n1162 gnd 0.006508f
C3971 vdd.n1163 gnd 0.006508f
C3972 vdd.n1164 gnd 0.006508f
C3973 vdd.n1165 gnd 0.006508f
C3974 vdd.n1166 gnd 0.396107f
C3975 vdd.n1167 gnd 0.006508f
C3976 vdd.n1168 gnd 0.006508f
C3977 vdd.n1169 gnd 0.006508f
C3978 vdd.n1170 gnd 0.006508f
C3979 vdd.n1171 gnd 0.006508f
C3980 vdd.n1172 gnd 0.006508f
C3981 vdd.n1173 gnd 0.006508f
C3982 vdd.n1174 gnd 0.006508f
C3983 vdd.n1175 gnd 0.006508f
C3984 vdd.n1176 gnd 0.006508f
C3985 vdd.n1177 gnd 0.006508f
C3986 vdd.n1178 gnd 0.006508f
C3987 vdd.n1179 gnd 0.006508f
C3988 vdd.n1180 gnd 0.006508f
C3989 vdd.n1181 gnd 0.006508f
C3990 vdd.n1182 gnd 0.006508f
C3991 vdd.n1183 gnd 0.006508f
C3992 vdd.n1184 gnd 0.006508f
C3993 vdd.n1185 gnd 0.006508f
C3994 vdd.n1186 gnd 0.006508f
C3995 vdd.n1187 gnd 0.210279f
C3996 vdd.n1188 gnd 0.006508f
C3997 vdd.n1189 gnd 0.006508f
C3998 vdd.n1190 gnd 0.006508f
C3999 vdd.n1191 gnd 0.006508f
C4000 vdd.n1192 gnd 0.006508f
C4001 vdd.n1193 gnd 0.006508f
C4002 vdd.n1194 gnd 0.006508f
C4003 vdd.n1195 gnd 0.006508f
C4004 vdd.n1196 gnd 0.006508f
C4005 vdd.n1197 gnd 0.006508f
C4006 vdd.n1198 gnd 0.006508f
C4007 vdd.n1199 gnd 0.006508f
C4008 vdd.n1200 gnd 0.006508f
C4009 vdd.n1201 gnd 0.006508f
C4010 vdd.n1202 gnd 0.006508f
C4011 vdd.n1203 gnd 0.006508f
C4012 vdd.n1204 gnd 0.006508f
C4013 vdd.n1205 gnd 0.006508f
C4014 vdd.n1206 gnd 0.006508f
C4015 vdd.n1207 gnd 0.006508f
C4016 vdd.n1208 gnd 0.006508f
C4017 vdd.n1209 gnd 0.006508f
C4018 vdd.n1210 gnd 0.006508f
C4019 vdd.n1211 gnd 0.006508f
C4020 vdd.n1212 gnd 0.006508f
C4021 vdd.n1213 gnd 0.006508f
C4022 vdd.n1214 gnd 0.006508f
C4023 vdd.n1215 gnd 0.014255f
C4024 vdd.n1216 gnd 0.014255f
C4025 vdd.n1217 gnd 0.015221f
C4026 vdd.n1218 gnd 0.006508f
C4027 vdd.n1219 gnd 0.006508f
C4028 vdd.n1220 gnd 0.005024f
C4029 vdd.n1221 gnd 0.006508f
C4030 vdd.n1222 gnd 0.006508f
C4031 vdd.n1223 gnd 0.004737f
C4032 vdd.n1224 gnd 0.006508f
C4033 vdd.n1225 gnd 0.006508f
C4034 vdd.n1226 gnd 0.006508f
C4035 vdd.n1227 gnd 0.006508f
C4036 vdd.n1228 gnd 0.006508f
C4037 vdd.n1229 gnd 0.006508f
C4038 vdd.n1230 gnd 0.006508f
C4039 vdd.n1231 gnd 0.006508f
C4040 vdd.n1232 gnd 0.006508f
C4041 vdd.n1233 gnd 0.006508f
C4042 vdd.n1234 gnd 0.006508f
C4043 vdd.n1235 gnd 0.006508f
C4044 vdd.n1236 gnd 0.006508f
C4045 vdd.n1237 gnd 0.006508f
C4046 vdd.n1238 gnd 0.006508f
C4047 vdd.n1239 gnd 0.006508f
C4048 vdd.n1240 gnd 0.006508f
C4049 vdd.n1241 gnd 0.006508f
C4050 vdd.n1242 gnd 0.006508f
C4051 vdd.n1243 gnd 0.006508f
C4052 vdd.n1244 gnd 0.006508f
C4053 vdd.n1245 gnd 0.006508f
C4054 vdd.n1246 gnd 0.006508f
C4055 vdd.n1247 gnd 0.006508f
C4056 vdd.n1248 gnd 0.006508f
C4057 vdd.n1249 gnd 0.006508f
C4058 vdd.n1250 gnd 0.026083f
C4059 vdd.n1252 gnd 0.022906f
C4060 vdd.n1253 gnd 0.007703f
C4061 vdd.n1255 gnd 0.00957f
C4062 vdd.n1256 gnd 0.007703f
C4063 vdd.n1257 gnd 0.00957f
C4064 vdd.n1259 gnd 0.00957f
C4065 vdd.n1260 gnd 0.00957f
C4066 vdd.n1262 gnd 0.00957f
C4067 vdd.n1263 gnd 0.006393f
C4068 vdd.t44 gnd 0.489021f
C4069 vdd.n1264 gnd 0.00957f
C4070 vdd.n1265 gnd 0.022906f
C4071 vdd.n1266 gnd 0.007703f
C4072 vdd.n1267 gnd 0.00957f
C4073 vdd.n1268 gnd 0.007703f
C4074 vdd.n1269 gnd 0.00957f
C4075 vdd.n1270 gnd 0.978042f
C4076 vdd.n1271 gnd 0.00957f
C4077 vdd.n1272 gnd 0.007703f
C4078 vdd.n1273 gnd 0.007703f
C4079 vdd.n1274 gnd 0.00957f
C4080 vdd.n1275 gnd 0.007703f
C4081 vdd.n1276 gnd 0.00957f
C4082 vdd.t168 gnd 0.489021f
C4083 vdd.n1277 gnd 0.00957f
C4084 vdd.n1278 gnd 0.007703f
C4085 vdd.n1279 gnd 0.00957f
C4086 vdd.n1280 gnd 0.007703f
C4087 vdd.n1281 gnd 0.00957f
C4088 vdd.t144 gnd 0.489021f
C4089 vdd.n1282 gnd 0.00957f
C4090 vdd.n1283 gnd 0.007703f
C4091 vdd.n1284 gnd 0.00957f
C4092 vdd.n1285 gnd 0.007703f
C4093 vdd.n1286 gnd 0.00957f
C4094 vdd.t185 gnd 0.489021f
C4095 vdd.n1287 gnd 0.767763f
C4096 vdd.n1288 gnd 0.00957f
C4097 vdd.n1289 gnd 0.007703f
C4098 vdd.n1290 gnd 0.00957f
C4099 vdd.n1291 gnd 0.007703f
C4100 vdd.n1292 gnd 0.00957f
C4101 vdd.n1293 gnd 0.68952f
C4102 vdd.n1294 gnd 0.00957f
C4103 vdd.n1295 gnd 0.007703f
C4104 vdd.n1296 gnd 0.00957f
C4105 vdd.n1297 gnd 0.007703f
C4106 vdd.n1298 gnd 0.00957f
C4107 vdd.n1299 gnd 0.523253f
C4108 vdd.t199 gnd 0.489021f
C4109 vdd.n1300 gnd 0.00957f
C4110 vdd.n1301 gnd 0.007703f
C4111 vdd.n1302 gnd 0.009537f
C4112 vdd.n1303 gnd 0.007703f
C4113 vdd.n1304 gnd 0.00957f
C4114 vdd.t181 gnd 0.489021f
C4115 vdd.n1305 gnd 0.00957f
C4116 vdd.n1306 gnd 0.007703f
C4117 vdd.n1307 gnd 0.00957f
C4118 vdd.n1308 gnd 0.007703f
C4119 vdd.n1309 gnd 0.00957f
C4120 vdd.t156 gnd 0.489021f
C4121 vdd.n1310 gnd 0.621057f
C4122 vdd.n1311 gnd 0.00957f
C4123 vdd.n1312 gnd 0.007703f
C4124 vdd.n1313 gnd 0.00957f
C4125 vdd.n1314 gnd 0.007703f
C4126 vdd.n1315 gnd 0.00957f
C4127 vdd.t142 gnd 0.489021f
C4128 vdd.n1316 gnd 0.00957f
C4129 vdd.n1317 gnd 0.007703f
C4130 vdd.n1318 gnd 0.00957f
C4131 vdd.n1319 gnd 0.007703f
C4132 vdd.n1320 gnd 0.00957f
C4133 vdd.n1321 gnd 0.669959f
C4134 vdd.n1322 gnd 0.811775f
C4135 vdd.t140 gnd 0.489021f
C4136 vdd.n1323 gnd 0.00957f
C4137 vdd.n1324 gnd 0.007703f
C4138 vdd.n1325 gnd 0.00957f
C4139 vdd.n1326 gnd 0.007703f
C4140 vdd.n1327 gnd 0.00957f
C4141 vdd.n1328 gnd 0.503692f
C4142 vdd.n1329 gnd 0.00957f
C4143 vdd.n1330 gnd 0.007703f
C4144 vdd.n1331 gnd 0.00957f
C4145 vdd.n1332 gnd 0.007703f
C4146 vdd.n1333 gnd 0.00957f
C4147 vdd.n1334 gnd 0.978042f
C4148 vdd.t148 gnd 0.489021f
C4149 vdd.n1335 gnd 0.00957f
C4150 vdd.n1336 gnd 0.007703f
C4151 vdd.n1337 gnd 0.00957f
C4152 vdd.n1338 gnd 0.007703f
C4153 vdd.n1339 gnd 0.00957f
C4154 vdd.t52 gnd 0.489021f
C4155 vdd.n1340 gnd 0.00957f
C4156 vdd.n1341 gnd 0.007703f
C4157 vdd.n1342 gnd 0.022906f
C4158 vdd.n1343 gnd 0.022906f
C4159 vdd.n1344 gnd 2.2495f
C4160 vdd.n1345 gnd 0.552594f
C4161 vdd.n1346 gnd 0.022906f
C4162 vdd.n1347 gnd 0.00957f
C4163 vdd.n1349 gnd 0.00957f
C4164 vdd.n1350 gnd 0.00957f
C4165 vdd.n1351 gnd 0.007703f
C4166 vdd.n1352 gnd 0.00957f
C4167 vdd.n1353 gnd 0.00957f
C4168 vdd.n1355 gnd 0.00957f
C4169 vdd.n1356 gnd 0.00957f
C4170 vdd.n1358 gnd 0.00957f
C4171 vdd.n1359 gnd 0.007703f
C4172 vdd.n1360 gnd 0.00957f
C4173 vdd.n1361 gnd 0.00957f
C4174 vdd.n1363 gnd 0.00957f
C4175 vdd.n1364 gnd 0.00957f
C4176 vdd.n1366 gnd 0.00957f
C4177 vdd.n1367 gnd 0.007703f
C4178 vdd.n1368 gnd 0.00957f
C4179 vdd.n1369 gnd 0.00957f
C4180 vdd.n1371 gnd 0.00957f
C4181 vdd.n1372 gnd 0.00957f
C4182 vdd.n1374 gnd 0.00957f
C4183 vdd.n1375 gnd 0.007703f
C4184 vdd.n1376 gnd 0.00957f
C4185 vdd.n1377 gnd 0.00957f
C4186 vdd.n1379 gnd 0.00957f
C4187 vdd.n1380 gnd 0.00957f
C4188 vdd.n1382 gnd 0.00957f
C4189 vdd.t72 gnd 0.11774f
C4190 vdd.t73 gnd 0.125832f
C4191 vdd.t71 gnd 0.153767f
C4192 vdd.n1383 gnd 0.197108f
C4193 vdd.n1384 gnd 0.166376f
C4194 vdd.n1385 gnd 0.016484f
C4195 vdd.n1386 gnd 0.00957f
C4196 vdd.n1387 gnd 0.00957f
C4197 vdd.n1389 gnd 0.00957f
C4198 vdd.n1390 gnd 0.00957f
C4199 vdd.n1392 gnd 0.00957f
C4200 vdd.n1393 gnd 0.007703f
C4201 vdd.n1394 gnd 0.00957f
C4202 vdd.n1395 gnd 0.00957f
C4203 vdd.n1397 gnd 0.00957f
C4204 vdd.n1398 gnd 0.00957f
C4205 vdd.n1400 gnd 0.00957f
C4206 vdd.n1401 gnd 0.007703f
C4207 vdd.n1402 gnd 0.00957f
C4208 vdd.n1403 gnd 0.00957f
C4209 vdd.n1405 gnd 0.00957f
C4210 vdd.n1406 gnd 0.00957f
C4211 vdd.n1408 gnd 0.00957f
C4212 vdd.n1409 gnd 0.007703f
C4213 vdd.n1410 gnd 0.00957f
C4214 vdd.n1411 gnd 0.00957f
C4215 vdd.n1413 gnd 0.00957f
C4216 vdd.n1414 gnd 0.00957f
C4217 vdd.n1416 gnd 0.00957f
C4218 vdd.n1417 gnd 0.007703f
C4219 vdd.n1418 gnd 0.00957f
C4220 vdd.n1419 gnd 0.00957f
C4221 vdd.n1421 gnd 0.00957f
C4222 vdd.n1422 gnd 0.00957f
C4223 vdd.n1424 gnd 0.00957f
C4224 vdd.n1425 gnd 0.007703f
C4225 vdd.n1426 gnd 0.00957f
C4226 vdd.n1427 gnd 0.00957f
C4227 vdd.n1429 gnd 0.00957f
C4228 vdd.n1430 gnd 0.007626f
C4229 vdd.n1432 gnd 0.007703f
C4230 vdd.n1433 gnd 0.00957f
C4231 vdd.n1434 gnd 0.00957f
C4232 vdd.n1435 gnd 0.00957f
C4233 vdd.n1436 gnd 0.00957f
C4234 vdd.n1438 gnd 0.00957f
C4235 vdd.n1439 gnd 0.00957f
C4236 vdd.n1440 gnd 0.007703f
C4237 vdd.n1441 gnd 0.00957f
C4238 vdd.n1443 gnd 0.00957f
C4239 vdd.n1444 gnd 0.00957f
C4240 vdd.n1446 gnd 0.00957f
C4241 vdd.n1447 gnd 0.00957f
C4242 vdd.n1448 gnd 0.007703f
C4243 vdd.n1449 gnd 0.00957f
C4244 vdd.n1451 gnd 0.00957f
C4245 vdd.n1452 gnd 0.00957f
C4246 vdd.n1454 gnd 0.00957f
C4247 vdd.n1455 gnd 0.00957f
C4248 vdd.n1456 gnd 0.007703f
C4249 vdd.n1457 gnd 0.00957f
C4250 vdd.n1459 gnd 0.00957f
C4251 vdd.n1460 gnd 0.00957f
C4252 vdd.n1462 gnd 0.00957f
C4253 vdd.n1463 gnd 0.00957f
C4254 vdd.n1464 gnd 0.007703f
C4255 vdd.n1465 gnd 0.00957f
C4256 vdd.n1467 gnd 0.00957f
C4257 vdd.n1468 gnd 0.00957f
C4258 vdd.n1470 gnd 0.00957f
C4259 vdd.n1471 gnd 0.003659f
C4260 vdd.t53 gnd 0.11774f
C4261 vdd.t54 gnd 0.125832f
C4262 vdd.t51 gnd 0.153767f
C4263 vdd.n1472 gnd 0.197108f
C4264 vdd.n1473 gnd 0.166376f
C4265 vdd.n1474 gnd 0.012633f
C4266 vdd.n1475 gnd 0.004044f
C4267 vdd.n1476 gnd 0.007703f
C4268 vdd.n1477 gnd 0.00957f
C4269 vdd.n1478 gnd 0.00957f
C4270 vdd.n1479 gnd 0.00957f
C4271 vdd.n1480 gnd 0.007703f
C4272 vdd.n1481 gnd 0.007703f
C4273 vdd.n1482 gnd 0.007703f
C4274 vdd.n1483 gnd 0.00957f
C4275 vdd.n1484 gnd 0.00957f
C4276 vdd.n1485 gnd 0.00957f
C4277 vdd.n1486 gnd 0.007703f
C4278 vdd.n1487 gnd 0.007703f
C4279 vdd.n1488 gnd 0.007703f
C4280 vdd.n1489 gnd 0.00957f
C4281 vdd.n1490 gnd 0.00957f
C4282 vdd.n1491 gnd 0.00957f
C4283 vdd.n1492 gnd 0.007703f
C4284 vdd.n1493 gnd 0.007703f
C4285 vdd.n1494 gnd 0.007703f
C4286 vdd.n1495 gnd 0.00957f
C4287 vdd.n1496 gnd 0.00957f
C4288 vdd.n1497 gnd 0.00957f
C4289 vdd.n1498 gnd 0.007703f
C4290 vdd.n1499 gnd 0.007703f
C4291 vdd.n1500 gnd 0.007703f
C4292 vdd.n1501 gnd 0.00957f
C4293 vdd.n1502 gnd 0.00957f
C4294 vdd.n1503 gnd 0.00957f
C4295 vdd.n1504 gnd 0.007703f
C4296 vdd.n1505 gnd 0.00957f
C4297 vdd.n1506 gnd 0.00957f
C4298 vdd.n1508 gnd 0.00957f
C4299 vdd.t59 gnd 0.11774f
C4300 vdd.t60 gnd 0.125832f
C4301 vdd.t58 gnd 0.153767f
C4302 vdd.n1509 gnd 0.197108f
C4303 vdd.n1510 gnd 0.166376f
C4304 vdd.n1511 gnd 0.016484f
C4305 vdd.n1512 gnd 0.005238f
C4306 vdd.n1513 gnd 0.00957f
C4307 vdd.n1514 gnd 0.00957f
C4308 vdd.n1515 gnd 0.00957f
C4309 vdd.n1516 gnd 0.007703f
C4310 vdd.n1517 gnd 0.007703f
C4311 vdd.n1518 gnd 0.007703f
C4312 vdd.n1519 gnd 0.00957f
C4313 vdd.n1520 gnd 0.00957f
C4314 vdd.n1521 gnd 0.00957f
C4315 vdd.n1522 gnd 0.007703f
C4316 vdd.n1523 gnd 0.007703f
C4317 vdd.n1524 gnd 0.007703f
C4318 vdd.n1525 gnd 0.00957f
C4319 vdd.n1526 gnd 0.00957f
C4320 vdd.n1527 gnd 0.00957f
C4321 vdd.n1528 gnd 0.007703f
C4322 vdd.n1529 gnd 0.007703f
C4323 vdd.n1530 gnd 0.007703f
C4324 vdd.n1531 gnd 0.00957f
C4325 vdd.n1532 gnd 0.00957f
C4326 vdd.n1533 gnd 0.00957f
C4327 vdd.n1534 gnd 0.007703f
C4328 vdd.n1535 gnd 0.007703f
C4329 vdd.n1536 gnd 0.007703f
C4330 vdd.n1537 gnd 0.00957f
C4331 vdd.n1538 gnd 0.00957f
C4332 vdd.n1539 gnd 0.00957f
C4333 vdd.n1540 gnd 0.007703f
C4334 vdd.n1541 gnd 0.007703f
C4335 vdd.n1542 gnd 0.006432f
C4336 vdd.n1543 gnd 0.00957f
C4337 vdd.n1544 gnd 0.00957f
C4338 vdd.n1545 gnd 0.00957f
C4339 vdd.n1546 gnd 0.006432f
C4340 vdd.n1547 gnd 0.007703f
C4341 vdd.n1548 gnd 0.007703f
C4342 vdd.n1549 gnd 0.00957f
C4343 vdd.n1550 gnd 0.00957f
C4344 vdd.n1551 gnd 0.00957f
C4345 vdd.n1552 gnd 0.007703f
C4346 vdd.n1553 gnd 0.007703f
C4347 vdd.n1554 gnd 0.007703f
C4348 vdd.n1555 gnd 0.00957f
C4349 vdd.n1556 gnd 0.00957f
C4350 vdd.n1557 gnd 0.00957f
C4351 vdd.n1558 gnd 0.007703f
C4352 vdd.n1559 gnd 0.007703f
C4353 vdd.n1560 gnd 0.007703f
C4354 vdd.n1561 gnd 0.00957f
C4355 vdd.n1562 gnd 0.00957f
C4356 vdd.n1563 gnd 0.00957f
C4357 vdd.n1564 gnd 0.007703f
C4358 vdd.n1565 gnd 0.007703f
C4359 vdd.n1566 gnd 0.007703f
C4360 vdd.n1567 gnd 0.00957f
C4361 vdd.n1568 gnd 0.00957f
C4362 vdd.n1569 gnd 0.00957f
C4363 vdd.n1570 gnd 0.007703f
C4364 vdd.n1571 gnd 0.007703f
C4365 vdd.n1572 gnd 0.006393f
C4366 vdd.n1573 gnd 0.022906f
C4367 vdd.n1574 gnd 0.022553f
C4368 vdd.n1575 gnd 0.006393f
C4369 vdd.n1576 gnd 0.022553f
C4370 vdd.n1577 gnd 1.37904f
C4371 vdd.n1578 gnd 0.022553f
C4372 vdd.n1579 gnd 0.006393f
C4373 vdd.n1580 gnd 0.022553f
C4374 vdd.n1581 gnd 0.00957f
C4375 vdd.n1582 gnd 0.00957f
C4376 vdd.n1583 gnd 0.007703f
C4377 vdd.n1584 gnd 0.00957f
C4378 vdd.n1585 gnd 0.914469f
C4379 vdd.n1586 gnd 0.00957f
C4380 vdd.n1587 gnd 0.007703f
C4381 vdd.n1588 gnd 0.00957f
C4382 vdd.n1589 gnd 0.00957f
C4383 vdd.n1590 gnd 0.00957f
C4384 vdd.n1591 gnd 0.007703f
C4385 vdd.n1592 gnd 0.00957f
C4386 vdd.n1593 gnd 0.963372f
C4387 vdd.n1594 gnd 0.00957f
C4388 vdd.n1595 gnd 0.007703f
C4389 vdd.n1596 gnd 0.00957f
C4390 vdd.n1597 gnd 0.00957f
C4391 vdd.n1598 gnd 0.00957f
C4392 vdd.n1599 gnd 0.007703f
C4393 vdd.n1600 gnd 0.00957f
C4394 vdd.t196 gnd 0.489021f
C4395 vdd.n1601 gnd 0.797104f
C4396 vdd.n1602 gnd 0.00957f
C4397 vdd.n1603 gnd 0.007703f
C4398 vdd.n1604 gnd 0.00957f
C4399 vdd.n1605 gnd 0.00957f
C4400 vdd.n1606 gnd 0.00957f
C4401 vdd.n1607 gnd 0.007703f
C4402 vdd.n1608 gnd 0.00957f
C4403 vdd.n1609 gnd 0.630837f
C4404 vdd.n1610 gnd 0.00957f
C4405 vdd.n1611 gnd 0.007703f
C4406 vdd.n1612 gnd 0.00957f
C4407 vdd.n1613 gnd 0.00957f
C4408 vdd.n1614 gnd 0.00957f
C4409 vdd.n1615 gnd 0.007703f
C4410 vdd.n1616 gnd 0.00957f
C4411 vdd.n1617 gnd 0.787324f
C4412 vdd.n1618 gnd 0.513472f
C4413 vdd.n1619 gnd 0.00957f
C4414 vdd.n1620 gnd 0.007703f
C4415 vdd.n1621 gnd 0.00957f
C4416 vdd.n1622 gnd 0.00957f
C4417 vdd.n1623 gnd 0.00957f
C4418 vdd.n1624 gnd 0.007703f
C4419 vdd.n1625 gnd 0.00957f
C4420 vdd.n1626 gnd 0.679739f
C4421 vdd.n1627 gnd 0.00957f
C4422 vdd.n1628 gnd 0.007703f
C4423 vdd.n1629 gnd 0.00957f
C4424 vdd.n1630 gnd 0.00957f
C4425 vdd.n1631 gnd 0.00957f
C4426 vdd.n1632 gnd 0.007703f
C4427 vdd.n1633 gnd 0.00957f
C4428 vdd.t150 gnd 0.489021f
C4429 vdd.n1634 gnd 0.811775f
C4430 vdd.n1635 gnd 0.00957f
C4431 vdd.n1636 gnd 0.007703f
C4432 vdd.n1637 gnd 0.005252f
C4433 vdd.n1638 gnd 0.004874f
C4434 vdd.n1639 gnd 0.002696f
C4435 vdd.n1640 gnd 0.00619f
C4436 vdd.n1641 gnd 0.002619f
C4437 vdd.n1642 gnd 0.002773f
C4438 vdd.n1643 gnd 0.004874f
C4439 vdd.n1644 gnd 0.002619f
C4440 vdd.n1645 gnd 0.00619f
C4441 vdd.n1646 gnd 0.002773f
C4442 vdd.n1647 gnd 0.004874f
C4443 vdd.n1648 gnd 0.002619f
C4444 vdd.n1649 gnd 0.004643f
C4445 vdd.n1650 gnd 0.004657f
C4446 vdd.t169 gnd 0.0133f
C4447 vdd.n1651 gnd 0.029591f
C4448 vdd.n1652 gnd 0.153999f
C4449 vdd.n1653 gnd 0.002619f
C4450 vdd.n1654 gnd 0.002773f
C4451 vdd.n1655 gnd 0.00619f
C4452 vdd.n1656 gnd 0.00619f
C4453 vdd.n1657 gnd 0.002773f
C4454 vdd.n1658 gnd 0.002619f
C4455 vdd.n1659 gnd 0.004874f
C4456 vdd.n1660 gnd 0.004874f
C4457 vdd.n1661 gnd 0.002619f
C4458 vdd.n1662 gnd 0.002773f
C4459 vdd.n1663 gnd 0.00619f
C4460 vdd.n1664 gnd 0.00619f
C4461 vdd.n1665 gnd 0.002773f
C4462 vdd.n1666 gnd 0.002619f
C4463 vdd.n1667 gnd 0.004874f
C4464 vdd.n1668 gnd 0.004874f
C4465 vdd.n1669 gnd 0.002619f
C4466 vdd.n1670 gnd 0.002773f
C4467 vdd.n1671 gnd 0.00619f
C4468 vdd.n1672 gnd 0.00619f
C4469 vdd.n1673 gnd 0.014635f
C4470 vdd.n1674 gnd 0.002696f
C4471 vdd.n1675 gnd 0.002619f
C4472 vdd.n1676 gnd 0.012597f
C4473 vdd.n1677 gnd 0.008795f
C4474 vdd.t186 gnd 0.030812f
C4475 vdd.t218 gnd 0.030812f
C4476 vdd.n1678 gnd 0.21176f
C4477 vdd.n1679 gnd 0.166517f
C4478 vdd.t200 gnd 0.030812f
C4479 vdd.t228 gnd 0.030812f
C4480 vdd.n1680 gnd 0.21176f
C4481 vdd.n1681 gnd 0.134378f
C4482 vdd.t182 gnd 0.030812f
C4483 vdd.t151 gnd 0.030812f
C4484 vdd.n1682 gnd 0.21176f
C4485 vdd.n1683 gnd 0.134378f
C4486 vdd.t143 gnd 0.030812f
C4487 vdd.t157 gnd 0.030812f
C4488 vdd.n1684 gnd 0.21176f
C4489 vdd.n1685 gnd 0.134378f
C4490 vdd.t221 gnd 0.030812f
C4491 vdd.t232 gnd 0.030812f
C4492 vdd.n1686 gnd 0.21176f
C4493 vdd.n1687 gnd 0.134378f
C4494 vdd.n1688 gnd 0.005252f
C4495 vdd.n1689 gnd 0.004874f
C4496 vdd.n1690 gnd 0.002696f
C4497 vdd.n1691 gnd 0.00619f
C4498 vdd.n1692 gnd 0.002619f
C4499 vdd.n1693 gnd 0.002773f
C4500 vdd.n1694 gnd 0.004874f
C4501 vdd.n1695 gnd 0.002619f
C4502 vdd.n1696 gnd 0.00619f
C4503 vdd.n1697 gnd 0.002773f
C4504 vdd.n1698 gnd 0.004874f
C4505 vdd.n1699 gnd 0.002619f
C4506 vdd.n1700 gnd 0.004643f
C4507 vdd.n1701 gnd 0.004657f
C4508 vdd.t161 gnd 0.0133f
C4509 vdd.n1702 gnd 0.029591f
C4510 vdd.n1703 gnd 0.153999f
C4511 vdd.n1704 gnd 0.002619f
C4512 vdd.n1705 gnd 0.002773f
C4513 vdd.n1706 gnd 0.00619f
C4514 vdd.n1707 gnd 0.00619f
C4515 vdd.n1708 gnd 0.002773f
C4516 vdd.n1709 gnd 0.002619f
C4517 vdd.n1710 gnd 0.004874f
C4518 vdd.n1711 gnd 0.004874f
C4519 vdd.n1712 gnd 0.002619f
C4520 vdd.n1713 gnd 0.002773f
C4521 vdd.n1714 gnd 0.00619f
C4522 vdd.n1715 gnd 0.00619f
C4523 vdd.n1716 gnd 0.002773f
C4524 vdd.n1717 gnd 0.002619f
C4525 vdd.n1718 gnd 0.004874f
C4526 vdd.n1719 gnd 0.004874f
C4527 vdd.n1720 gnd 0.002619f
C4528 vdd.n1721 gnd 0.002773f
C4529 vdd.n1722 gnd 0.00619f
C4530 vdd.n1723 gnd 0.00619f
C4531 vdd.n1724 gnd 0.014635f
C4532 vdd.n1725 gnd 0.002696f
C4533 vdd.n1726 gnd 0.002619f
C4534 vdd.n1727 gnd 0.012597f
C4535 vdd.n1728 gnd 0.008519f
C4536 vdd.n1729 gnd 0.099978f
C4537 vdd.n1730 gnd 0.005252f
C4538 vdd.n1731 gnd 0.004874f
C4539 vdd.n1732 gnd 0.002696f
C4540 vdd.n1733 gnd 0.00619f
C4541 vdd.n1734 gnd 0.002619f
C4542 vdd.n1735 gnd 0.002773f
C4543 vdd.n1736 gnd 0.004874f
C4544 vdd.n1737 gnd 0.002619f
C4545 vdd.n1738 gnd 0.00619f
C4546 vdd.n1739 gnd 0.002773f
C4547 vdd.n1740 gnd 0.004874f
C4548 vdd.n1741 gnd 0.002619f
C4549 vdd.n1742 gnd 0.004643f
C4550 vdd.n1743 gnd 0.004657f
C4551 vdd.t216 gnd 0.0133f
C4552 vdd.n1744 gnd 0.029591f
C4553 vdd.n1745 gnd 0.153999f
C4554 vdd.n1746 gnd 0.002619f
C4555 vdd.n1747 gnd 0.002773f
C4556 vdd.n1748 gnd 0.00619f
C4557 vdd.n1749 gnd 0.00619f
C4558 vdd.n1750 gnd 0.002773f
C4559 vdd.n1751 gnd 0.002619f
C4560 vdd.n1752 gnd 0.004874f
C4561 vdd.n1753 gnd 0.004874f
C4562 vdd.n1754 gnd 0.002619f
C4563 vdd.n1755 gnd 0.002773f
C4564 vdd.n1756 gnd 0.00619f
C4565 vdd.n1757 gnd 0.00619f
C4566 vdd.n1758 gnd 0.002773f
C4567 vdd.n1759 gnd 0.002619f
C4568 vdd.n1760 gnd 0.004874f
C4569 vdd.n1761 gnd 0.004874f
C4570 vdd.n1762 gnd 0.002619f
C4571 vdd.n1763 gnd 0.002773f
C4572 vdd.n1764 gnd 0.00619f
C4573 vdd.n1765 gnd 0.00619f
C4574 vdd.n1766 gnd 0.014635f
C4575 vdd.n1767 gnd 0.002696f
C4576 vdd.n1768 gnd 0.002619f
C4577 vdd.n1769 gnd 0.012597f
C4578 vdd.n1770 gnd 0.008795f
C4579 vdd.t191 gnd 0.030812f
C4580 vdd.t145 gnd 0.030812f
C4581 vdd.n1771 gnd 0.21176f
C4582 vdd.n1772 gnd 0.166517f
C4583 vdd.t226 gnd 0.030812f
C4584 vdd.t207 gnd 0.030812f
C4585 vdd.n1773 gnd 0.21176f
C4586 vdd.n1774 gnd 0.134378f
C4587 vdd.t204 gnd 0.030812f
C4588 vdd.t170 gnd 0.030812f
C4589 vdd.n1775 gnd 0.21176f
C4590 vdd.n1776 gnd 0.134378f
C4591 vdd.t164 gnd 0.030812f
C4592 vdd.t205 gnd 0.030812f
C4593 vdd.n1777 gnd 0.21176f
C4594 vdd.n1778 gnd 0.134378f
C4595 vdd.t197 gnd 0.030812f
C4596 vdd.t141 gnd 0.030812f
C4597 vdd.n1779 gnd 0.21176f
C4598 vdd.n1780 gnd 0.134378f
C4599 vdd.n1781 gnd 0.005252f
C4600 vdd.n1782 gnd 0.004874f
C4601 vdd.n1783 gnd 0.002696f
C4602 vdd.n1784 gnd 0.00619f
C4603 vdd.n1785 gnd 0.002619f
C4604 vdd.n1786 gnd 0.002773f
C4605 vdd.n1787 gnd 0.004874f
C4606 vdd.n1788 gnd 0.002619f
C4607 vdd.n1789 gnd 0.00619f
C4608 vdd.n1790 gnd 0.002773f
C4609 vdd.n1791 gnd 0.004874f
C4610 vdd.n1792 gnd 0.002619f
C4611 vdd.n1793 gnd 0.004643f
C4612 vdd.n1794 gnd 0.004657f
C4613 vdd.t149 gnd 0.0133f
C4614 vdd.n1795 gnd 0.029591f
C4615 vdd.n1796 gnd 0.153999f
C4616 vdd.n1797 gnd 0.002619f
C4617 vdd.n1798 gnd 0.002773f
C4618 vdd.n1799 gnd 0.00619f
C4619 vdd.n1800 gnd 0.00619f
C4620 vdd.n1801 gnd 0.002773f
C4621 vdd.n1802 gnd 0.002619f
C4622 vdd.n1803 gnd 0.004874f
C4623 vdd.n1804 gnd 0.004874f
C4624 vdd.n1805 gnd 0.002619f
C4625 vdd.n1806 gnd 0.002773f
C4626 vdd.n1807 gnd 0.00619f
C4627 vdd.n1808 gnd 0.00619f
C4628 vdd.n1809 gnd 0.002773f
C4629 vdd.n1810 gnd 0.002619f
C4630 vdd.n1811 gnd 0.004874f
C4631 vdd.n1812 gnd 0.004874f
C4632 vdd.n1813 gnd 0.002619f
C4633 vdd.n1814 gnd 0.002773f
C4634 vdd.n1815 gnd 0.00619f
C4635 vdd.n1816 gnd 0.00619f
C4636 vdd.n1817 gnd 0.014635f
C4637 vdd.n1818 gnd 0.002696f
C4638 vdd.n1819 gnd 0.002619f
C4639 vdd.n1820 gnd 0.012597f
C4640 vdd.n1821 gnd 0.008519f
C4641 vdd.n1822 gnd 0.059477f
C4642 vdd.n1823 gnd 0.214311f
C4643 vdd.n1824 gnd 0.005252f
C4644 vdd.n1825 gnd 0.004874f
C4645 vdd.n1826 gnd 0.002696f
C4646 vdd.n1827 gnd 0.00619f
C4647 vdd.n1828 gnd 0.002619f
C4648 vdd.n1829 gnd 0.002773f
C4649 vdd.n1830 gnd 0.004874f
C4650 vdd.n1831 gnd 0.002619f
C4651 vdd.n1832 gnd 0.00619f
C4652 vdd.n1833 gnd 0.002773f
C4653 vdd.n1834 gnd 0.004874f
C4654 vdd.n1835 gnd 0.002619f
C4655 vdd.n1836 gnd 0.004643f
C4656 vdd.n1837 gnd 0.004657f
C4657 vdd.t225 gnd 0.0133f
C4658 vdd.n1838 gnd 0.029591f
C4659 vdd.n1839 gnd 0.153999f
C4660 vdd.n1840 gnd 0.002619f
C4661 vdd.n1841 gnd 0.002773f
C4662 vdd.n1842 gnd 0.00619f
C4663 vdd.n1843 gnd 0.00619f
C4664 vdd.n1844 gnd 0.002773f
C4665 vdd.n1845 gnd 0.002619f
C4666 vdd.n1846 gnd 0.004874f
C4667 vdd.n1847 gnd 0.004874f
C4668 vdd.n1848 gnd 0.002619f
C4669 vdd.n1849 gnd 0.002773f
C4670 vdd.n1850 gnd 0.00619f
C4671 vdd.n1851 gnd 0.00619f
C4672 vdd.n1852 gnd 0.002773f
C4673 vdd.n1853 gnd 0.002619f
C4674 vdd.n1854 gnd 0.004874f
C4675 vdd.n1855 gnd 0.004874f
C4676 vdd.n1856 gnd 0.002619f
C4677 vdd.n1857 gnd 0.002773f
C4678 vdd.n1858 gnd 0.00619f
C4679 vdd.n1859 gnd 0.00619f
C4680 vdd.n1860 gnd 0.014635f
C4681 vdd.n1861 gnd 0.002696f
C4682 vdd.n1862 gnd 0.002619f
C4683 vdd.n1863 gnd 0.012597f
C4684 vdd.n1864 gnd 0.008795f
C4685 vdd.t198 gnd 0.030812f
C4686 vdd.t162 gnd 0.030812f
C4687 vdd.n1865 gnd 0.21176f
C4688 vdd.n1866 gnd 0.166517f
C4689 vdd.t233 gnd 0.030812f
C4690 vdd.t214 gnd 0.030812f
C4691 vdd.n1867 gnd 0.21176f
C4692 vdd.n1868 gnd 0.134378f
C4693 vdd.t211 gnd 0.030812f
C4694 vdd.t184 gnd 0.030812f
C4695 vdd.n1869 gnd 0.21176f
C4696 vdd.n1870 gnd 0.134378f
C4697 vdd.t183 gnd 0.030812f
C4698 vdd.t213 gnd 0.030812f
C4699 vdd.n1871 gnd 0.21176f
C4700 vdd.n1872 gnd 0.134378f
C4701 vdd.t203 gnd 0.030812f
C4702 vdd.t202 gnd 0.030812f
C4703 vdd.n1873 gnd 0.21176f
C4704 vdd.n1874 gnd 0.134378f
C4705 vdd.n1875 gnd 0.005252f
C4706 vdd.n1876 gnd 0.004874f
C4707 vdd.n1877 gnd 0.002696f
C4708 vdd.n1878 gnd 0.00619f
C4709 vdd.n1879 gnd 0.002619f
C4710 vdd.n1880 gnd 0.002773f
C4711 vdd.n1881 gnd 0.004874f
C4712 vdd.n1882 gnd 0.002619f
C4713 vdd.n1883 gnd 0.00619f
C4714 vdd.n1884 gnd 0.002773f
C4715 vdd.n1885 gnd 0.004874f
C4716 vdd.n1886 gnd 0.002619f
C4717 vdd.n1887 gnd 0.004643f
C4718 vdd.n1888 gnd 0.004657f
C4719 vdd.t163 gnd 0.0133f
C4720 vdd.n1889 gnd 0.029591f
C4721 vdd.n1890 gnd 0.153999f
C4722 vdd.n1891 gnd 0.002619f
C4723 vdd.n1892 gnd 0.002773f
C4724 vdd.n1893 gnd 0.00619f
C4725 vdd.n1894 gnd 0.00619f
C4726 vdd.n1895 gnd 0.002773f
C4727 vdd.n1896 gnd 0.002619f
C4728 vdd.n1897 gnd 0.004874f
C4729 vdd.n1898 gnd 0.004874f
C4730 vdd.n1899 gnd 0.002619f
C4731 vdd.n1900 gnd 0.002773f
C4732 vdd.n1901 gnd 0.00619f
C4733 vdd.n1902 gnd 0.00619f
C4734 vdd.n1903 gnd 0.002773f
C4735 vdd.n1904 gnd 0.002619f
C4736 vdd.n1905 gnd 0.004874f
C4737 vdd.n1906 gnd 0.004874f
C4738 vdd.n1907 gnd 0.002619f
C4739 vdd.n1908 gnd 0.002773f
C4740 vdd.n1909 gnd 0.00619f
C4741 vdd.n1910 gnd 0.00619f
C4742 vdd.n1911 gnd 0.014635f
C4743 vdd.n1912 gnd 0.002696f
C4744 vdd.n1913 gnd 0.002619f
C4745 vdd.n1914 gnd 0.012597f
C4746 vdd.n1915 gnd 0.008519f
C4747 vdd.n1916 gnd 0.059477f
C4748 vdd.n1917 gnd 0.235534f
C4749 vdd.n1918 gnd 2.23536f
C4750 vdd.n1919 gnd 0.5697f
C4751 vdd.n1920 gnd 0.009537f
C4752 vdd.n1921 gnd 0.00957f
C4753 vdd.n1922 gnd 0.007703f
C4754 vdd.n1923 gnd 0.00957f
C4755 vdd.n1924 gnd 0.777544f
C4756 vdd.n1925 gnd 0.00957f
C4757 vdd.n1926 gnd 0.007703f
C4758 vdd.n1927 gnd 0.00957f
C4759 vdd.n1928 gnd 0.00957f
C4760 vdd.n1929 gnd 0.00957f
C4761 vdd.n1930 gnd 0.007703f
C4762 vdd.n1931 gnd 0.00957f
C4763 vdd.n1932 gnd 0.811775f
C4764 vdd.t206 gnd 0.489021f
C4765 vdd.n1933 gnd 0.611276f
C4766 vdd.n1934 gnd 0.00957f
C4767 vdd.n1935 gnd 0.007703f
C4768 vdd.n1936 gnd 0.00957f
C4769 vdd.n1937 gnd 0.00957f
C4770 vdd.n1938 gnd 0.00957f
C4771 vdd.n1939 gnd 0.007703f
C4772 vdd.n1940 gnd 0.00957f
C4773 vdd.n1941 gnd 0.533033f
C4774 vdd.n1942 gnd 0.00957f
C4775 vdd.n1943 gnd 0.007703f
C4776 vdd.n1944 gnd 0.00957f
C4777 vdd.n1945 gnd 0.00957f
C4778 vdd.n1946 gnd 0.00957f
C4779 vdd.n1947 gnd 0.007703f
C4780 vdd.n1948 gnd 0.00957f
C4781 vdd.n1949 gnd 0.601496f
C4782 vdd.n1950 gnd 0.6993f
C4783 vdd.n1951 gnd 0.00957f
C4784 vdd.n1952 gnd 0.007703f
C4785 vdd.n1953 gnd 0.00957f
C4786 vdd.n1954 gnd 0.00957f
C4787 vdd.n1955 gnd 0.00957f
C4788 vdd.n1956 gnd 0.007703f
C4789 vdd.n1957 gnd 0.00957f
C4790 vdd.n1958 gnd 0.865567f
C4791 vdd.n1959 gnd 0.00957f
C4792 vdd.n1960 gnd 0.007703f
C4793 vdd.n1961 gnd 0.00957f
C4794 vdd.n1962 gnd 0.00957f
C4795 vdd.n1963 gnd 0.022553f
C4796 vdd.n1964 gnd 0.00957f
C4797 vdd.n1965 gnd 0.00957f
C4798 vdd.n1966 gnd 0.007703f
C4799 vdd.n1967 gnd 0.00957f
C4800 vdd.n1968 gnd 0.523253f
C4801 vdd.n1969 gnd 0.978042f
C4802 vdd.n1970 gnd 0.00957f
C4803 vdd.n1971 gnd 0.007703f
C4804 vdd.n1972 gnd 0.00957f
C4805 vdd.n1973 gnd 0.00957f
C4806 vdd.n1974 gnd 0.022553f
C4807 vdd.n1975 gnd 0.006393f
C4808 vdd.n1976 gnd 0.022553f
C4809 vdd.n1977 gnd 1.34481f
C4810 vdd.n1978 gnd 0.022553f
C4811 vdd.n1979 gnd 0.022906f
C4812 vdd.n1980 gnd 0.003659f
C4813 vdd.t46 gnd 0.11774f
C4814 vdd.t45 gnd 0.125832f
C4815 vdd.t43 gnd 0.153767f
C4816 vdd.n1981 gnd 0.197108f
C4817 vdd.n1982 gnd 0.165606f
C4818 vdd.n1983 gnd 0.011863f
C4819 vdd.n1984 gnd 0.004044f
C4820 vdd.n1985 gnd 0.00823f
C4821 vdd.n1986 gnd 0.72376f
C4822 vdd.n1988 gnd 0.007703f
C4823 vdd.n1989 gnd 0.007703f
C4824 vdd.n1990 gnd 0.00957f
C4825 vdd.n1992 gnd 0.00957f
C4826 vdd.n1993 gnd 0.00957f
C4827 vdd.n1994 gnd 0.007703f
C4828 vdd.n1995 gnd 0.007703f
C4829 vdd.n1996 gnd 0.007703f
C4830 vdd.n1997 gnd 0.00957f
C4831 vdd.n1999 gnd 0.00957f
C4832 vdd.n2000 gnd 0.00957f
C4833 vdd.n2001 gnd 0.007703f
C4834 vdd.n2002 gnd 0.007703f
C4835 vdd.n2003 gnd 0.007703f
C4836 vdd.n2004 gnd 0.00957f
C4837 vdd.n2006 gnd 0.00957f
C4838 vdd.n2007 gnd 0.00957f
C4839 vdd.n2008 gnd 0.007703f
C4840 vdd.n2009 gnd 0.007703f
C4841 vdd.n2010 gnd 0.007703f
C4842 vdd.n2011 gnd 0.00957f
C4843 vdd.n2013 gnd 0.00957f
C4844 vdd.n2014 gnd 0.00957f
C4845 vdd.n2015 gnd 0.007703f
C4846 vdd.n2016 gnd 0.00957f
C4847 vdd.n2017 gnd 0.00957f
C4848 vdd.n2018 gnd 0.00957f
C4849 vdd.n2019 gnd 0.015714f
C4850 vdd.n2020 gnd 0.005238f
C4851 vdd.n2021 gnd 0.007703f
C4852 vdd.n2022 gnd 0.00957f
C4853 vdd.n2024 gnd 0.00957f
C4854 vdd.n2025 gnd 0.00957f
C4855 vdd.n2026 gnd 0.007703f
C4856 vdd.n2027 gnd 0.007703f
C4857 vdd.n2028 gnd 0.007703f
C4858 vdd.n2029 gnd 0.00957f
C4859 vdd.n2031 gnd 0.00957f
C4860 vdd.n2032 gnd 0.00957f
C4861 vdd.n2033 gnd 0.007703f
C4862 vdd.n2034 gnd 0.007703f
C4863 vdd.n2035 gnd 0.007703f
C4864 vdd.n2036 gnd 0.00957f
C4865 vdd.n2038 gnd 0.00957f
C4866 vdd.n2039 gnd 0.00957f
C4867 vdd.n2040 gnd 0.007703f
C4868 vdd.n2041 gnd 0.007703f
C4869 vdd.n2042 gnd 0.007703f
C4870 vdd.n2043 gnd 0.00957f
C4871 vdd.n2045 gnd 0.00957f
C4872 vdd.n2046 gnd 0.00957f
C4873 vdd.n2047 gnd 0.007703f
C4874 vdd.n2048 gnd 0.007703f
C4875 vdd.n2049 gnd 0.007703f
C4876 vdd.n2050 gnd 0.00957f
C4877 vdd.n2052 gnd 0.00957f
C4878 vdd.n2053 gnd 0.00957f
C4879 vdd.n2054 gnd 0.007703f
C4880 vdd.n2055 gnd 0.00957f
C4881 vdd.n2056 gnd 0.00957f
C4882 vdd.n2057 gnd 0.00957f
C4883 vdd.n2058 gnd 0.015714f
C4884 vdd.n2059 gnd 0.006432f
C4885 vdd.n2060 gnd 0.007703f
C4886 vdd.n2061 gnd 0.00957f
C4887 vdd.n2063 gnd 0.00957f
C4888 vdd.n2064 gnd 0.00957f
C4889 vdd.n2065 gnd 0.007703f
C4890 vdd.n2066 gnd 0.007703f
C4891 vdd.n2067 gnd 0.007703f
C4892 vdd.n2068 gnd 0.00957f
C4893 vdd.n2070 gnd 0.00957f
C4894 vdd.n2071 gnd 0.00957f
C4895 vdd.n2072 gnd 0.007703f
C4896 vdd.n2073 gnd 0.007703f
C4897 vdd.n2074 gnd 0.007703f
C4898 vdd.n2075 gnd 0.00957f
C4899 vdd.n2077 gnd 0.00957f
C4900 vdd.n2078 gnd 0.00957f
C4901 vdd.n2079 gnd 0.007703f
C4902 vdd.n2080 gnd 0.007703f
C4903 vdd.n2081 gnd 0.007703f
C4904 vdd.n2082 gnd 0.00957f
C4905 vdd.n2084 gnd 0.00957f
C4906 vdd.n2085 gnd 0.007703f
C4907 vdd.n2086 gnd 0.007703f
C4908 vdd.n2087 gnd 0.00957f
C4909 vdd.n2089 gnd 0.00957f
C4910 vdd.n2090 gnd 0.00957f
C4911 vdd.n2091 gnd 0.007703f
C4912 vdd.n2092 gnd 0.00823f
C4913 vdd.n2093 gnd 0.72376f
C4914 vdd.n2094 gnd 0.026083f
C4915 vdd.n2095 gnd 0.006508f
C4916 vdd.n2096 gnd 0.006508f
C4917 vdd.n2097 gnd 0.006508f
C4918 vdd.n2098 gnd 0.006508f
C4919 vdd.n2099 gnd 0.006508f
C4920 vdd.n2100 gnd 0.006508f
C4921 vdd.n2101 gnd 0.006508f
C4922 vdd.n2102 gnd 0.006508f
C4923 vdd.n2103 gnd 0.006508f
C4924 vdd.n2104 gnd 0.006508f
C4925 vdd.n2105 gnd 0.006508f
C4926 vdd.n2106 gnd 0.006508f
C4927 vdd.n2107 gnd 0.006508f
C4928 vdd.n2108 gnd 0.006508f
C4929 vdd.n2109 gnd 0.006508f
C4930 vdd.n2110 gnd 0.006508f
C4931 vdd.n2111 gnd 0.006508f
C4932 vdd.n2112 gnd 0.006508f
C4933 vdd.n2113 gnd 0.006508f
C4934 vdd.n2114 gnd 0.006508f
C4935 vdd.n2115 gnd 0.006508f
C4936 vdd.n2116 gnd 0.006508f
C4937 vdd.n2117 gnd 0.006508f
C4938 vdd.n2118 gnd 0.006508f
C4939 vdd.n2119 gnd 0.006508f
C4940 vdd.n2120 gnd 0.006508f
C4941 vdd.n2121 gnd 0.006508f
C4942 vdd.n2122 gnd 0.006508f
C4943 vdd.n2123 gnd 0.006508f
C4944 vdd.n2124 gnd 0.006508f
C4945 vdd.n2125 gnd 0.006508f
C4946 vdd.n2126 gnd 0.015221f
C4947 vdd.n2127 gnd 0.015221f
C4948 vdd.n2129 gnd 8.3427f
C4949 vdd.n2131 gnd 0.015221f
C4950 vdd.n2132 gnd 0.015221f
C4951 vdd.n2133 gnd 0.014255f
C4952 vdd.n2134 gnd 0.006508f
C4953 vdd.n2135 gnd 0.006508f
C4954 vdd.n2136 gnd 0.665069f
C4955 vdd.n2137 gnd 0.006508f
C4956 vdd.n2138 gnd 0.006508f
C4957 vdd.n2139 gnd 0.006508f
C4958 vdd.n2140 gnd 0.006508f
C4959 vdd.n2141 gnd 0.006508f
C4960 vdd.n2142 gnd 0.562374f
C4961 vdd.n2143 gnd 0.006508f
C4962 vdd.n2144 gnd 0.006508f
C4963 vdd.n2145 gnd 0.006508f
C4964 vdd.n2146 gnd 0.006508f
C4965 vdd.n2147 gnd 0.006508f
C4966 vdd.n2148 gnd 0.665069f
C4967 vdd.n2149 gnd 0.006508f
C4968 vdd.n2150 gnd 0.006508f
C4969 vdd.n2151 gnd 0.006508f
C4970 vdd.n2152 gnd 0.006508f
C4971 vdd.n2153 gnd 0.006508f
C4972 vdd.n2154 gnd 0.650398f
C4973 vdd.n2155 gnd 0.006508f
C4974 vdd.n2156 gnd 0.006508f
C4975 vdd.n2157 gnd 0.006508f
C4976 vdd.n2158 gnd 0.006508f
C4977 vdd.n2159 gnd 0.006508f
C4978 vdd.n2160 gnd 0.665069f
C4979 vdd.n2161 gnd 0.006508f
C4980 vdd.n2162 gnd 0.006508f
C4981 vdd.n2163 gnd 0.006508f
C4982 vdd.n2164 gnd 0.006508f
C4983 vdd.n2165 gnd 0.006508f
C4984 vdd.n2166 gnd 0.533033f
C4985 vdd.n2167 gnd 0.006508f
C4986 vdd.n2168 gnd 0.006508f
C4987 vdd.n2169 gnd 0.005551f
C4988 vdd.n2170 gnd 0.018852f
C4989 vdd.n2171 gnd 0.004211f
C4990 vdd.n2172 gnd 0.006508f
C4991 vdd.n2173 gnd 0.386327f
C4992 vdd.n2174 gnd 0.006508f
C4993 vdd.n2175 gnd 0.006508f
C4994 vdd.n2176 gnd 0.006508f
C4995 vdd.n2177 gnd 0.006508f
C4996 vdd.n2178 gnd 0.006508f
C4997 vdd.n2179 gnd 0.425448f
C4998 vdd.n2180 gnd 0.006508f
C4999 vdd.n2181 gnd 0.006508f
C5000 vdd.n2182 gnd 0.006508f
C5001 vdd.n2183 gnd 0.006508f
C5002 vdd.n2184 gnd 0.006508f
C5003 vdd.n2185 gnd 0.572155f
C5004 vdd.n2186 gnd 0.006508f
C5005 vdd.n2187 gnd 0.006508f
C5006 vdd.n2188 gnd 0.006508f
C5007 vdd.n2189 gnd 0.006508f
C5008 vdd.n2190 gnd 0.006508f
C5009 vdd.n2191 gnd 0.547704f
C5010 vdd.n2192 gnd 0.006508f
C5011 vdd.n2193 gnd 0.006508f
C5012 vdd.n2194 gnd 0.006508f
C5013 vdd.n2195 gnd 0.006508f
C5014 vdd.n2196 gnd 0.006508f
C5015 vdd.n2197 gnd 0.400997f
C5016 vdd.n2198 gnd 0.006508f
C5017 vdd.n2199 gnd 0.006508f
C5018 vdd.n2200 gnd 0.006508f
C5019 vdd.n2201 gnd 0.006508f
C5020 vdd.n2202 gnd 0.006508f
C5021 vdd.n2203 gnd 0.210279f
C5022 vdd.n2204 gnd 0.006508f
C5023 vdd.n2205 gnd 0.006508f
C5024 vdd.n2206 gnd 0.006508f
C5025 vdd.n2207 gnd 0.006508f
C5026 vdd.n2208 gnd 0.006508f
C5027 vdd.n2209 gnd 0.347205f
C5028 vdd.n2210 gnd 0.006508f
C5029 vdd.n2211 gnd 0.006508f
C5030 vdd.n2212 gnd 0.006508f
C5031 vdd.n2213 gnd 0.006508f
C5032 vdd.n2214 gnd 0.006508f
C5033 vdd.n2215 gnd 0.665069f
C5034 vdd.n2216 gnd 0.006508f
C5035 vdd.n2217 gnd 0.006508f
C5036 vdd.n2218 gnd 0.006508f
C5037 vdd.n2219 gnd 0.006508f
C5038 vdd.n2220 gnd 0.006508f
C5039 vdd.n2221 gnd 0.006508f
C5040 vdd.n2222 gnd 0.006508f
C5041 vdd.n2223 gnd 0.498801f
C5042 vdd.n2224 gnd 0.006508f
C5043 vdd.n2225 gnd 0.006508f
C5044 vdd.n2226 gnd 0.006508f
C5045 vdd.n2227 gnd 0.006508f
C5046 vdd.n2228 gnd 0.006508f
C5047 vdd.n2229 gnd 0.006508f
C5048 vdd.n2230 gnd 0.415668f
C5049 vdd.n2231 gnd 0.006508f
C5050 vdd.n2232 gnd 0.006508f
C5051 vdd.n2233 gnd 0.006508f
C5052 vdd.n2234 gnd 0.015064f
C5053 vdd.n2235 gnd 0.014413f
C5054 vdd.n2236 gnd 0.006508f
C5055 vdd.n2237 gnd 0.006508f
C5056 vdd.n2238 gnd 0.005024f
C5057 vdd.n2239 gnd 0.006508f
C5058 vdd.n2240 gnd 0.006508f
C5059 vdd.n2241 gnd 0.004737f
C5060 vdd.n2242 gnd 0.006508f
C5061 vdd.n2243 gnd 0.006508f
C5062 vdd.n2244 gnd 0.006508f
C5063 vdd.n2245 gnd 0.006508f
C5064 vdd.n2246 gnd 0.006508f
C5065 vdd.n2247 gnd 0.006508f
C5066 vdd.n2248 gnd 0.006508f
C5067 vdd.n2249 gnd 0.006508f
C5068 vdd.n2250 gnd 0.006508f
C5069 vdd.n2251 gnd 0.006508f
C5070 vdd.n2252 gnd 0.006508f
C5071 vdd.n2253 gnd 0.006508f
C5072 vdd.n2254 gnd 0.006508f
C5073 vdd.n2255 gnd 0.006508f
C5074 vdd.n2256 gnd 0.006508f
C5075 vdd.n2257 gnd 0.006508f
C5076 vdd.n2258 gnd 0.006508f
C5077 vdd.n2259 gnd 0.006508f
C5078 vdd.n2260 gnd 0.006508f
C5079 vdd.n2261 gnd 0.006508f
C5080 vdd.n2262 gnd 0.006508f
C5081 vdd.n2263 gnd 0.006508f
C5082 vdd.n2264 gnd 0.006508f
C5083 vdd.n2265 gnd 0.006508f
C5084 vdd.n2266 gnd 0.006508f
C5085 vdd.n2267 gnd 0.006508f
C5086 vdd.n2268 gnd 0.006508f
C5087 vdd.n2269 gnd 0.006508f
C5088 vdd.n2270 gnd 0.006508f
C5089 vdd.n2271 gnd 0.006508f
C5090 vdd.n2272 gnd 0.006508f
C5091 vdd.n2273 gnd 0.006508f
C5092 vdd.n2274 gnd 0.006508f
C5093 vdd.n2275 gnd 0.006508f
C5094 vdd.n2276 gnd 0.006508f
C5095 vdd.n2277 gnd 0.006508f
C5096 vdd.n2278 gnd 0.006508f
C5097 vdd.n2279 gnd 0.006508f
C5098 vdd.n2280 gnd 0.006508f
C5099 vdd.n2281 gnd 0.006508f
C5100 vdd.n2282 gnd 0.006508f
C5101 vdd.n2283 gnd 0.006508f
C5102 vdd.n2284 gnd 0.006508f
C5103 vdd.n2285 gnd 0.006508f
C5104 vdd.n2286 gnd 0.006508f
C5105 vdd.n2287 gnd 0.006508f
C5106 vdd.n2288 gnd 0.006508f
C5107 vdd.n2289 gnd 0.006508f
C5108 vdd.n2290 gnd 0.006508f
C5109 vdd.n2291 gnd 0.006508f
C5110 vdd.n2292 gnd 0.006508f
C5111 vdd.n2293 gnd 0.006508f
C5112 vdd.n2294 gnd 0.006508f
C5113 vdd.n2295 gnd 0.006508f
C5114 vdd.n2296 gnd 0.006508f
C5115 vdd.n2297 gnd 0.006508f
C5116 vdd.n2298 gnd 0.006508f
C5117 vdd.n2299 gnd 0.006508f
C5118 vdd.n2300 gnd 0.006508f
C5119 vdd.n2301 gnd 0.006508f
C5120 vdd.n2302 gnd 0.015221f
C5121 vdd.n2303 gnd 0.014255f
C5122 vdd.n2304 gnd 0.014255f
C5123 vdd.n2305 gnd 0.792214f
C5124 vdd.n2306 gnd 0.014255f
C5125 vdd.n2307 gnd 0.015221f
C5126 vdd.n2308 gnd 0.014413f
C5127 vdd.n2309 gnd 0.006508f
C5128 vdd.n2310 gnd 0.006508f
C5129 vdd.n2311 gnd 0.006508f
C5130 vdd.n2312 gnd 0.005024f
C5131 vdd.n2313 gnd 0.009301f
C5132 vdd.n2314 gnd 0.004737f
C5133 vdd.n2315 gnd 0.006508f
C5134 vdd.n2316 gnd 0.006508f
C5135 vdd.n2317 gnd 0.006508f
C5136 vdd.n2318 gnd 0.006508f
C5137 vdd.n2319 gnd 0.006508f
C5138 vdd.n2320 gnd 0.006508f
C5139 vdd.n2321 gnd 0.006508f
C5140 vdd.n2322 gnd 0.006508f
C5141 vdd.n2323 gnd 0.006508f
C5142 vdd.n2324 gnd 0.006508f
C5143 vdd.n2325 gnd 0.006508f
C5144 vdd.n2326 gnd 0.006508f
C5145 vdd.n2327 gnd 0.006508f
C5146 vdd.n2328 gnd 0.006508f
C5147 vdd.n2329 gnd 0.006508f
C5148 vdd.n2330 gnd 0.006508f
C5149 vdd.n2331 gnd 0.006508f
C5150 vdd.n2332 gnd 0.006508f
C5151 vdd.n2333 gnd 0.006508f
C5152 vdd.n2334 gnd 0.006508f
C5153 vdd.n2335 gnd 0.006508f
C5154 vdd.n2336 gnd 0.006508f
C5155 vdd.n2337 gnd 0.006508f
C5156 vdd.n2338 gnd 0.006508f
C5157 vdd.n2339 gnd 0.006508f
C5158 vdd.n2340 gnd 0.006508f
C5159 vdd.n2341 gnd 0.006508f
C5160 vdd.n2342 gnd 0.006508f
C5161 vdd.n2343 gnd 0.006508f
C5162 vdd.n2344 gnd 0.006508f
C5163 vdd.n2345 gnd 0.006508f
C5164 vdd.n2346 gnd 0.006508f
C5165 vdd.n2347 gnd 0.006508f
C5166 vdd.n2348 gnd 0.006508f
C5167 vdd.n2349 gnd 0.006508f
C5168 vdd.n2350 gnd 0.006508f
C5169 vdd.n2351 gnd 0.006508f
C5170 vdd.n2352 gnd 0.006508f
C5171 vdd.n2353 gnd 0.006508f
C5172 vdd.n2354 gnd 0.006508f
C5173 vdd.n2355 gnd 0.006508f
C5174 vdd.n2356 gnd 0.006508f
C5175 vdd.n2357 gnd 0.006508f
C5176 vdd.n2358 gnd 0.006508f
C5177 vdd.n2359 gnd 0.006508f
C5178 vdd.n2360 gnd 0.006508f
C5179 vdd.n2361 gnd 0.006508f
C5180 vdd.n2362 gnd 0.006508f
C5181 vdd.n2363 gnd 0.006508f
C5182 vdd.n2364 gnd 0.006508f
C5183 vdd.n2365 gnd 0.006508f
C5184 vdd.n2366 gnd 0.006508f
C5185 vdd.n2367 gnd 0.006508f
C5186 vdd.n2368 gnd 0.006508f
C5187 vdd.n2369 gnd 0.006508f
C5188 vdd.n2370 gnd 0.006508f
C5189 vdd.n2371 gnd 0.006508f
C5190 vdd.n2372 gnd 0.006508f
C5191 vdd.n2373 gnd 0.006508f
C5192 vdd.n2374 gnd 0.006508f
C5193 vdd.n2375 gnd 0.015221f
C5194 vdd.n2376 gnd 0.015221f
C5195 vdd.n2377 gnd 0.811775f
C5196 vdd.t11 gnd 2.88522f
C5197 vdd.t29 gnd 2.88522f
C5198 vdd.n2410 gnd 0.015221f
C5199 vdd.t7 gnd 0.606386f
C5200 vdd.n2411 gnd 0.006508f
C5201 vdd.n2412 gnd 0.006508f
C5202 vdd.t83 gnd 0.26298f
C5203 vdd.t84 gnd 0.269193f
C5204 vdd.t81 gnd 0.171684f
C5205 vdd.n2413 gnd 0.092785f
C5206 vdd.n2414 gnd 0.052631f
C5207 vdd.n2415 gnd 0.006508f
C5208 vdd.t90 gnd 0.26298f
C5209 vdd.t91 gnd 0.269193f
C5210 vdd.t89 gnd 0.171684f
C5211 vdd.n2416 gnd 0.092785f
C5212 vdd.n2417 gnd 0.052631f
C5213 vdd.n2418 gnd 0.009301f
C5214 vdd.n2419 gnd 0.006508f
C5215 vdd.n2420 gnd 0.006508f
C5216 vdd.n2421 gnd 0.006508f
C5217 vdd.n2422 gnd 0.006508f
C5218 vdd.n2423 gnd 0.006508f
C5219 vdd.n2424 gnd 0.006508f
C5220 vdd.n2425 gnd 0.006508f
C5221 vdd.n2426 gnd 0.006508f
C5222 vdd.n2427 gnd 0.006508f
C5223 vdd.n2428 gnd 0.006508f
C5224 vdd.n2429 gnd 0.006508f
C5225 vdd.n2430 gnd 0.006508f
C5226 vdd.n2431 gnd 0.006508f
C5227 vdd.n2432 gnd 0.006508f
C5228 vdd.n2433 gnd 0.006508f
C5229 vdd.n2434 gnd 0.006508f
C5230 vdd.n2435 gnd 0.006508f
C5231 vdd.n2436 gnd 0.006508f
C5232 vdd.n2437 gnd 0.006508f
C5233 vdd.n2438 gnd 0.006508f
C5234 vdd.n2439 gnd 0.006508f
C5235 vdd.n2440 gnd 0.006508f
C5236 vdd.n2441 gnd 0.006508f
C5237 vdd.n2442 gnd 0.006508f
C5238 vdd.n2443 gnd 0.006508f
C5239 vdd.n2444 gnd 0.006508f
C5240 vdd.n2445 gnd 0.006508f
C5241 vdd.n2446 gnd 0.006508f
C5242 vdd.n2447 gnd 0.006508f
C5243 vdd.n2448 gnd 0.006508f
C5244 vdd.n2449 gnd 0.006508f
C5245 vdd.n2450 gnd 0.006508f
C5246 vdd.n2451 gnd 0.006508f
C5247 vdd.n2452 gnd 0.006508f
C5248 vdd.n2453 gnd 0.006508f
C5249 vdd.n2454 gnd 0.006508f
C5250 vdd.n2455 gnd 0.006508f
C5251 vdd.n2456 gnd 0.006508f
C5252 vdd.n2457 gnd 0.006508f
C5253 vdd.n2458 gnd 0.006508f
C5254 vdd.n2459 gnd 0.006508f
C5255 vdd.n2460 gnd 0.006508f
C5256 vdd.n2461 gnd 0.006508f
C5257 vdd.n2462 gnd 0.006508f
C5258 vdd.n2463 gnd 0.006508f
C5259 vdd.n2464 gnd 0.006508f
C5260 vdd.n2465 gnd 0.006508f
C5261 vdd.n2466 gnd 0.006508f
C5262 vdd.n2467 gnd 0.006508f
C5263 vdd.n2468 gnd 0.006508f
C5264 vdd.n2469 gnd 0.006508f
C5265 vdd.n2470 gnd 0.006508f
C5266 vdd.n2471 gnd 0.006508f
C5267 vdd.n2472 gnd 0.006508f
C5268 vdd.n2473 gnd 0.006508f
C5269 vdd.n2474 gnd 0.006508f
C5270 vdd.n2475 gnd 0.006508f
C5271 vdd.n2476 gnd 0.006508f
C5272 vdd.n2477 gnd 0.004737f
C5273 vdd.n2478 gnd 0.006508f
C5274 vdd.n2479 gnd 0.006508f
C5275 vdd.n2480 gnd 0.005024f
C5276 vdd.n2481 gnd 0.006508f
C5277 vdd.n2482 gnd 0.006508f
C5278 vdd.n2483 gnd 0.015221f
C5279 vdd.n2484 gnd 0.014255f
C5280 vdd.n2485 gnd 0.014255f
C5281 vdd.n2486 gnd 0.006508f
C5282 vdd.n2487 gnd 0.006508f
C5283 vdd.n2488 gnd 0.006508f
C5284 vdd.n2489 gnd 0.006508f
C5285 vdd.n2490 gnd 0.006508f
C5286 vdd.n2491 gnd 0.006508f
C5287 vdd.n2492 gnd 0.006508f
C5288 vdd.n2493 gnd 0.006508f
C5289 vdd.n2494 gnd 0.006508f
C5290 vdd.n2495 gnd 0.006508f
C5291 vdd.n2496 gnd 0.006508f
C5292 vdd.n2497 gnd 0.006508f
C5293 vdd.n2498 gnd 0.006508f
C5294 vdd.n2499 gnd 0.006508f
C5295 vdd.n2500 gnd 0.006508f
C5296 vdd.n2501 gnd 0.006508f
C5297 vdd.n2502 gnd 0.006508f
C5298 vdd.n2503 gnd 0.006508f
C5299 vdd.n2504 gnd 0.006508f
C5300 vdd.n2505 gnd 0.006508f
C5301 vdd.n2506 gnd 0.006508f
C5302 vdd.n2507 gnd 0.006508f
C5303 vdd.n2508 gnd 0.006508f
C5304 vdd.n2509 gnd 0.006508f
C5305 vdd.n2510 gnd 0.006508f
C5306 vdd.n2511 gnd 0.006508f
C5307 vdd.n2512 gnd 0.006508f
C5308 vdd.n2513 gnd 0.006508f
C5309 vdd.n2514 gnd 0.006508f
C5310 vdd.n2515 gnd 0.006508f
C5311 vdd.n2516 gnd 0.006508f
C5312 vdd.n2517 gnd 0.006508f
C5313 vdd.n2518 gnd 0.006508f
C5314 vdd.n2519 gnd 0.006508f
C5315 vdd.n2520 gnd 0.006508f
C5316 vdd.n2521 gnd 0.006508f
C5317 vdd.n2522 gnd 0.006508f
C5318 vdd.n2523 gnd 0.006508f
C5319 vdd.n2524 gnd 0.006508f
C5320 vdd.n2525 gnd 0.006508f
C5321 vdd.n2526 gnd 0.006508f
C5322 vdd.n2527 gnd 0.006508f
C5323 vdd.n2528 gnd 0.006508f
C5324 vdd.n2529 gnd 0.006508f
C5325 vdd.n2530 gnd 0.006508f
C5326 vdd.n2531 gnd 0.006508f
C5327 vdd.n2532 gnd 0.006508f
C5328 vdd.n2533 gnd 0.006508f
C5329 vdd.n2534 gnd 0.006508f
C5330 vdd.n2535 gnd 0.006508f
C5331 vdd.n2536 gnd 0.006508f
C5332 vdd.n2537 gnd 0.006508f
C5333 vdd.n2538 gnd 0.006508f
C5334 vdd.n2539 gnd 0.006508f
C5335 vdd.n2540 gnd 0.006508f
C5336 vdd.n2541 gnd 0.006508f
C5337 vdd.n2542 gnd 0.006508f
C5338 vdd.n2543 gnd 0.006508f
C5339 vdd.n2544 gnd 0.006508f
C5340 vdd.n2545 gnd 0.006508f
C5341 vdd.n2546 gnd 0.006508f
C5342 vdd.n2547 gnd 0.006508f
C5343 vdd.n2548 gnd 0.006508f
C5344 vdd.n2549 gnd 0.006508f
C5345 vdd.n2550 gnd 0.006508f
C5346 vdd.n2551 gnd 0.006508f
C5347 vdd.n2552 gnd 0.006508f
C5348 vdd.n2553 gnd 0.006508f
C5349 vdd.n2554 gnd 0.006508f
C5350 vdd.n2555 gnd 0.006508f
C5351 vdd.n2556 gnd 0.006508f
C5352 vdd.n2557 gnd 0.006508f
C5353 vdd.n2558 gnd 0.006508f
C5354 vdd.n2559 gnd 0.210279f
C5355 vdd.n2560 gnd 0.006508f
C5356 vdd.n2561 gnd 0.006508f
C5357 vdd.n2562 gnd 0.006508f
C5358 vdd.n2563 gnd 0.006508f
C5359 vdd.n2564 gnd 0.006508f
C5360 vdd.n2565 gnd 0.006508f
C5361 vdd.n2566 gnd 0.006508f
C5362 vdd.n2567 gnd 0.006508f
C5363 vdd.n2568 gnd 0.006508f
C5364 vdd.n2569 gnd 0.006508f
C5365 vdd.n2570 gnd 0.006508f
C5366 vdd.n2571 gnd 0.006508f
C5367 vdd.n2572 gnd 0.006508f
C5368 vdd.n2573 gnd 0.006508f
C5369 vdd.n2574 gnd 0.415668f
C5370 vdd.n2575 gnd 0.006508f
C5371 vdd.n2576 gnd 0.006508f
C5372 vdd.n2577 gnd 0.006508f
C5373 vdd.n2578 gnd 0.014255f
C5374 vdd.n2579 gnd 0.014255f
C5375 vdd.n2580 gnd 0.015221f
C5376 vdd.n2581 gnd 0.015221f
C5377 vdd.n2582 gnd 0.006508f
C5378 vdd.n2583 gnd 0.006508f
C5379 vdd.n2584 gnd 0.006508f
C5380 vdd.n2585 gnd 0.005024f
C5381 vdd.n2586 gnd 0.009301f
C5382 vdd.n2587 gnd 0.004737f
C5383 vdd.n2588 gnd 0.006508f
C5384 vdd.n2589 gnd 0.006508f
C5385 vdd.n2590 gnd 0.006508f
C5386 vdd.n2591 gnd 0.006508f
C5387 vdd.n2592 gnd 0.006508f
C5388 vdd.n2593 gnd 0.006508f
C5389 vdd.n2594 gnd 0.006508f
C5390 vdd.n2595 gnd 0.006508f
C5391 vdd.n2596 gnd 0.006508f
C5392 vdd.n2597 gnd 0.006508f
C5393 vdd.n2598 gnd 0.006508f
C5394 vdd.n2599 gnd 0.006508f
C5395 vdd.n2600 gnd 0.006508f
C5396 vdd.n2601 gnd 0.006508f
C5397 vdd.n2602 gnd 0.006508f
C5398 vdd.n2603 gnd 0.006508f
C5399 vdd.n2604 gnd 0.006508f
C5400 vdd.n2605 gnd 0.006508f
C5401 vdd.n2606 gnd 0.006508f
C5402 vdd.n2607 gnd 0.006508f
C5403 vdd.n2608 gnd 0.006508f
C5404 vdd.n2609 gnd 0.006508f
C5405 vdd.n2610 gnd 0.006508f
C5406 vdd.n2611 gnd 0.006508f
C5407 vdd.n2612 gnd 0.006508f
C5408 vdd.n2613 gnd 0.006508f
C5409 vdd.n2614 gnd 0.006508f
C5410 vdd.n2615 gnd 0.006508f
C5411 vdd.n2616 gnd 0.006508f
C5412 vdd.n2617 gnd 0.006508f
C5413 vdd.n2618 gnd 0.006508f
C5414 vdd.n2619 gnd 0.006508f
C5415 vdd.n2620 gnd 0.006508f
C5416 vdd.n2621 gnd 0.006508f
C5417 vdd.n2622 gnd 0.006508f
C5418 vdd.n2623 gnd 0.006508f
C5419 vdd.n2624 gnd 0.006508f
C5420 vdd.n2625 gnd 0.006508f
C5421 vdd.n2626 gnd 0.006508f
C5422 vdd.n2627 gnd 0.006508f
C5423 vdd.n2628 gnd 0.006508f
C5424 vdd.n2629 gnd 0.006508f
C5425 vdd.n2630 gnd 0.006508f
C5426 vdd.n2631 gnd 0.006508f
C5427 vdd.n2632 gnd 0.006508f
C5428 vdd.n2633 gnd 0.006508f
C5429 vdd.n2634 gnd 0.006508f
C5430 vdd.n2635 gnd 0.006508f
C5431 vdd.n2636 gnd 0.006508f
C5432 vdd.n2637 gnd 0.006508f
C5433 vdd.n2638 gnd 0.006508f
C5434 vdd.n2639 gnd 0.006508f
C5435 vdd.n2640 gnd 0.006508f
C5436 vdd.n2641 gnd 0.006508f
C5437 vdd.n2642 gnd 0.006508f
C5438 vdd.n2643 gnd 0.006508f
C5439 vdd.n2644 gnd 0.006508f
C5440 vdd.n2645 gnd 0.006508f
C5441 vdd.n2646 gnd 0.006508f
C5442 vdd.n2647 gnd 0.015221f
C5443 vdd.n2648 gnd 0.015221f
C5444 vdd.n2650 gnd 0.811775f
C5445 vdd.n2652 gnd 0.015221f
C5446 vdd.n2653 gnd 0.015221f
C5447 vdd.n2654 gnd 0.014255f
C5448 vdd.n2655 gnd 0.006508f
C5449 vdd.n2656 gnd 0.006508f
C5450 vdd.n2657 gnd 0.352095f
C5451 vdd.n2658 gnd 0.006508f
C5452 vdd.n2659 gnd 0.006508f
C5453 vdd.n2660 gnd 0.006508f
C5454 vdd.n2661 gnd 0.006508f
C5455 vdd.n2662 gnd 0.006508f
C5456 vdd.n2663 gnd 0.396107f
C5457 vdd.n2664 gnd 0.006508f
C5458 vdd.n2665 gnd 0.006508f
C5459 vdd.n2666 gnd 0.006508f
C5460 vdd.n2667 gnd 0.006508f
C5461 vdd.n2668 gnd 0.006508f
C5462 vdd.n2669 gnd 0.665069f
C5463 vdd.n2670 gnd 0.006508f
C5464 vdd.n2671 gnd 0.006508f
C5465 vdd.n2672 gnd 0.006508f
C5466 vdd.n2673 gnd 0.006508f
C5467 vdd.n2674 gnd 0.006508f
C5468 vdd.n2675 gnd 0.440119f
C5469 vdd.n2676 gnd 0.006508f
C5470 vdd.n2677 gnd 0.006508f
C5471 vdd.n2678 gnd 0.006508f
C5472 vdd.n2679 gnd 0.006508f
C5473 vdd.n2680 gnd 0.006508f
C5474 vdd.n2681 gnd 0.586825f
C5475 vdd.n2682 gnd 0.006508f
C5476 vdd.n2683 gnd 0.006508f
C5477 vdd.n2684 gnd 0.006508f
C5478 vdd.n2685 gnd 0.006508f
C5479 vdd.n2686 gnd 0.006508f
C5480 vdd.n2687 gnd 0.533033f
C5481 vdd.n2688 gnd 0.006508f
C5482 vdd.n2689 gnd 0.006508f
C5483 vdd.n2690 gnd 0.006508f
C5484 vdd.n2691 gnd 0.006508f
C5485 vdd.n2692 gnd 0.006508f
C5486 vdd.n2693 gnd 0.386327f
C5487 vdd.n2694 gnd 0.006508f
C5488 vdd.n2695 gnd 0.006508f
C5489 vdd.n2696 gnd 0.006508f
C5490 vdd.n2697 gnd 0.006508f
C5491 vdd.n2698 gnd 0.006508f
C5492 vdd.n2699 gnd 0.210279f
C5493 vdd.n2700 gnd 0.006508f
C5494 vdd.n2701 gnd 0.006508f
C5495 vdd.n2702 gnd 0.006508f
C5496 vdd.n2703 gnd 0.006508f
C5497 vdd.n2704 gnd 0.006508f
C5498 vdd.n2705 gnd 0.572155f
C5499 vdd.n2706 gnd 0.006508f
C5500 vdd.n2707 gnd 0.006508f
C5501 vdd.n2708 gnd 0.006508f
C5502 vdd.n2709 gnd 0.006508f
C5503 vdd.n2710 gnd 0.006508f
C5504 vdd.n2711 gnd 0.665069f
C5505 vdd.n2712 gnd 0.006508f
C5506 vdd.n2713 gnd 0.006508f
C5507 vdd.n2714 gnd 0.004211f
C5508 vdd.n2715 gnd 0.018852f
C5509 vdd.n2716 gnd 0.005551f
C5510 vdd.n2717 gnd 0.006508f
C5511 vdd.n2718 gnd 0.567264f
C5512 vdd.n2719 gnd 0.006508f
C5513 vdd.n2720 gnd 0.006508f
C5514 vdd.n2721 gnd 0.006508f
C5515 vdd.n2722 gnd 0.006508f
C5516 vdd.n2723 gnd 0.006508f
C5517 vdd.n2724 gnd 0.46457f
C5518 vdd.n2725 gnd 0.006508f
C5519 vdd.n2726 gnd 0.006508f
C5520 vdd.n2727 gnd 0.006508f
C5521 vdd.n2728 gnd 0.006508f
C5522 vdd.n2729 gnd 0.006508f
C5523 vdd.n2730 gnd 0.347205f
C5524 vdd.n2731 gnd 0.006508f
C5525 vdd.n2732 gnd 0.006508f
C5526 vdd.n2733 gnd 0.006508f
C5527 vdd.n2734 gnd 0.006508f
C5528 vdd.n2735 gnd 0.006508f
C5529 vdd.n2736 gnd 0.665069f
C5530 vdd.n2737 gnd 0.006508f
C5531 vdd.n2738 gnd 0.006508f
C5532 vdd.n2739 gnd 0.006508f
C5533 vdd.n2740 gnd 0.006508f
C5534 vdd.n2741 gnd 0.006508f
C5535 vdd.n2742 gnd 0.006508f
C5536 vdd.n2744 gnd 0.006508f
C5537 vdd.n2745 gnd 0.006508f
C5538 vdd.n2747 gnd 0.006508f
C5539 vdd.n2748 gnd 0.006508f
C5540 vdd.n2751 gnd 0.006508f
C5541 vdd.n2752 gnd 0.006508f
C5542 vdd.n2753 gnd 0.006508f
C5543 vdd.n2754 gnd 0.006508f
C5544 vdd.n2756 gnd 0.006508f
C5545 vdd.n2757 gnd 0.006508f
C5546 vdd.n2758 gnd 0.006508f
C5547 vdd.n2759 gnd 0.006508f
C5548 vdd.n2760 gnd 0.006508f
C5549 vdd.n2761 gnd 0.006508f
C5550 vdd.n2763 gnd 0.006508f
C5551 vdd.n2764 gnd 0.006508f
C5552 vdd.n2765 gnd 0.006508f
C5553 vdd.n2766 gnd 0.006508f
C5554 vdd.n2767 gnd 0.006508f
C5555 vdd.n2768 gnd 0.006508f
C5556 vdd.n2770 gnd 0.006508f
C5557 vdd.n2771 gnd 0.006508f
C5558 vdd.n2772 gnd 0.006508f
C5559 vdd.n2773 gnd 0.006508f
C5560 vdd.n2774 gnd 0.006508f
C5561 vdd.n2775 gnd 0.006508f
C5562 vdd.n2777 gnd 0.006508f
C5563 vdd.n2778 gnd 0.015221f
C5564 vdd.n2779 gnd 0.015221f
C5565 vdd.n2780 gnd 0.014255f
C5566 vdd.n2781 gnd 0.006508f
C5567 vdd.n2782 gnd 0.006508f
C5568 vdd.n2783 gnd 0.006508f
C5569 vdd.n2784 gnd 0.006508f
C5570 vdd.n2785 gnd 0.006508f
C5571 vdd.n2786 gnd 0.006508f
C5572 vdd.n2787 gnd 0.665069f
C5573 vdd.n2788 gnd 0.006508f
C5574 vdd.n2789 gnd 0.006508f
C5575 vdd.n2790 gnd 0.006508f
C5576 vdd.n2791 gnd 0.006508f
C5577 vdd.n2792 gnd 0.006508f
C5578 vdd.n2793 gnd 0.435229f
C5579 vdd.n2794 gnd 0.006508f
C5580 vdd.n2795 gnd 0.006508f
C5581 vdd.n2796 gnd 0.006508f
C5582 vdd.n2797 gnd 0.015064f
C5583 vdd.n2799 gnd 0.015221f
C5584 vdd.n2800 gnd 0.014413f
C5585 vdd.n2801 gnd 0.006508f
C5586 vdd.n2802 gnd 0.005024f
C5587 vdd.n2803 gnd 0.006508f
C5588 vdd.n2805 gnd 0.006508f
C5589 vdd.n2806 gnd 0.006508f
C5590 vdd.n2807 gnd 0.006508f
C5591 vdd.n2808 gnd 0.006508f
C5592 vdd.n2809 gnd 0.006508f
C5593 vdd.n2810 gnd 0.006508f
C5594 vdd.n2812 gnd 0.006508f
C5595 vdd.n2813 gnd 0.006508f
C5596 vdd.n2814 gnd 0.006508f
C5597 vdd.n2815 gnd 0.006508f
C5598 vdd.n2816 gnd 0.006508f
C5599 vdd.n2817 gnd 0.006508f
C5600 vdd.n2819 gnd 0.006508f
C5601 vdd.n2820 gnd 0.006508f
C5602 vdd.n2821 gnd 0.006508f
C5603 vdd.n2822 gnd 0.006508f
C5604 vdd.n2823 gnd 0.006508f
C5605 vdd.n2824 gnd 0.006508f
C5606 vdd.n2826 gnd 0.006508f
C5607 vdd.n2827 gnd 0.006508f
C5608 vdd.n2828 gnd 0.006508f
C5609 vdd.n2829 gnd 0.727493f
C5610 vdd.n2830 gnd 0.02235f
C5611 vdd.n2831 gnd 0.006508f
C5612 vdd.n2832 gnd 0.006508f
C5613 vdd.n2834 gnd 0.006508f
C5614 vdd.n2835 gnd 0.006508f
C5615 vdd.n2836 gnd 0.006508f
C5616 vdd.n2837 gnd 0.006508f
C5617 vdd.n2838 gnd 0.006508f
C5618 vdd.n2839 gnd 0.006508f
C5619 vdd.n2841 gnd 0.006508f
C5620 vdd.n2842 gnd 0.006508f
C5621 vdd.n2843 gnd 0.006508f
C5622 vdd.n2844 gnd 0.006508f
C5623 vdd.n2845 gnd 0.006508f
C5624 vdd.n2846 gnd 0.006508f
C5625 vdd.n2848 gnd 0.006508f
C5626 vdd.n2849 gnd 0.006508f
C5627 vdd.n2850 gnd 0.006508f
C5628 vdd.n2851 gnd 0.006508f
C5629 vdd.n2852 gnd 0.006508f
C5630 vdd.n2853 gnd 0.006508f
C5631 vdd.n2855 gnd 0.006508f
C5632 vdd.n2856 gnd 0.006508f
C5633 vdd.n2858 gnd 0.006508f
C5634 vdd.n2859 gnd 0.006508f
C5635 vdd.n2860 gnd 0.015221f
C5636 vdd.n2861 gnd 0.014255f
C5637 vdd.n2862 gnd 0.014255f
C5638 vdd.n2863 gnd 0.93892f
C5639 vdd.n2864 gnd 0.014255f
C5640 vdd.n2865 gnd 0.015221f
C5641 vdd.n2866 gnd 0.014413f
C5642 vdd.n2867 gnd 0.006508f
C5643 vdd.n2868 gnd 0.005024f
C5644 vdd.n2869 gnd 0.006508f
C5645 vdd.n2871 gnd 0.006508f
C5646 vdd.n2872 gnd 0.006508f
C5647 vdd.n2873 gnd 0.006508f
C5648 vdd.n2874 gnd 0.006508f
C5649 vdd.n2875 gnd 0.006508f
C5650 vdd.n2876 gnd 0.006508f
C5651 vdd.n2878 gnd 0.006508f
C5652 vdd.n2879 gnd 0.006508f
C5653 vdd.n2880 gnd 0.006508f
C5654 vdd.n2881 gnd 0.006508f
C5655 vdd.n2882 gnd 0.006508f
C5656 vdd.n2883 gnd 0.006508f
C5657 vdd.n2885 gnd 0.006508f
C5658 vdd.n2886 gnd 0.006508f
C5659 vdd.n2887 gnd 0.006508f
C5660 vdd.n2888 gnd 0.006508f
C5661 vdd.n2889 gnd 0.006508f
C5662 vdd.n2890 gnd 0.006508f
C5663 vdd.n2892 gnd 0.006508f
C5664 vdd.n2893 gnd 0.006508f
C5665 vdd.n2895 gnd 0.006508f
C5666 vdd.n2896 gnd 0.02235f
C5667 vdd.n2897 gnd 0.727493f
C5668 vdd.n2898 gnd 0.00823f
C5669 vdd.n2899 gnd 0.003659f
C5670 vdd.t41 gnd 0.11774f
C5671 vdd.t42 gnd 0.125832f
C5672 vdd.t39 gnd 0.153767f
C5673 vdd.n2900 gnd 0.197108f
C5674 vdd.n2901 gnd 0.165606f
C5675 vdd.n2902 gnd 0.011863f
C5676 vdd.n2903 gnd 0.00957f
C5677 vdd.n2904 gnd 0.004044f
C5678 vdd.n2905 gnd 0.007703f
C5679 vdd.n2906 gnd 0.00957f
C5680 vdd.n2907 gnd 0.00957f
C5681 vdd.n2908 gnd 0.007703f
C5682 vdd.n2909 gnd 0.007703f
C5683 vdd.n2910 gnd 0.00957f
C5684 vdd.n2912 gnd 0.00957f
C5685 vdd.n2913 gnd 0.007703f
C5686 vdd.n2914 gnd 0.007703f
C5687 vdd.n2915 gnd 0.007703f
C5688 vdd.n2916 gnd 0.00957f
C5689 vdd.n2918 gnd 0.00957f
C5690 vdd.n2920 gnd 0.00957f
C5691 vdd.n2921 gnd 0.007703f
C5692 vdd.n2922 gnd 0.007703f
C5693 vdd.n2923 gnd 0.007703f
C5694 vdd.n2924 gnd 0.00957f
C5695 vdd.n2926 gnd 0.00957f
C5696 vdd.n2928 gnd 0.00957f
C5697 vdd.n2929 gnd 0.007703f
C5698 vdd.n2930 gnd 0.007703f
C5699 vdd.n2931 gnd 0.007703f
C5700 vdd.n2932 gnd 0.00957f
C5701 vdd.n2934 gnd 0.00957f
C5702 vdd.n2935 gnd 0.00957f
C5703 vdd.n2936 gnd 0.007703f
C5704 vdd.n2937 gnd 0.007703f
C5705 vdd.n2938 gnd 0.00957f
C5706 vdd.n2939 gnd 0.00957f
C5707 vdd.n2941 gnd 0.00957f
C5708 vdd.n2942 gnd 0.007703f
C5709 vdd.n2943 gnd 0.00957f
C5710 vdd.n2944 gnd 0.00957f
C5711 vdd.n2945 gnd 0.00957f
C5712 vdd.n2946 gnd 0.015714f
C5713 vdd.n2947 gnd 0.005238f
C5714 vdd.n2948 gnd 0.00957f
C5715 vdd.n2950 gnd 0.00957f
C5716 vdd.n2952 gnd 0.00957f
C5717 vdd.n2953 gnd 0.007703f
C5718 vdd.n2954 gnd 0.007703f
C5719 vdd.n2955 gnd 0.007703f
C5720 vdd.n2956 gnd 0.00957f
C5721 vdd.n2958 gnd 0.00957f
C5722 vdd.n2960 gnd 0.00957f
C5723 vdd.n2961 gnd 0.007703f
C5724 vdd.n2962 gnd 0.007703f
C5725 vdd.n2963 gnd 0.007703f
C5726 vdd.n2964 gnd 0.00957f
C5727 vdd.n2966 gnd 0.00957f
C5728 vdd.n2968 gnd 0.00957f
C5729 vdd.n2969 gnd 0.007703f
C5730 vdd.n2970 gnd 0.007703f
C5731 vdd.n2971 gnd 0.007703f
C5732 vdd.n2972 gnd 0.00957f
C5733 vdd.n2974 gnd 0.00957f
C5734 vdd.n2976 gnd 0.00957f
C5735 vdd.n2977 gnd 0.007703f
C5736 vdd.n2978 gnd 0.007703f
C5737 vdd.n2979 gnd 0.007703f
C5738 vdd.n2980 gnd 0.00957f
C5739 vdd.n2982 gnd 0.00957f
C5740 vdd.n2984 gnd 0.00957f
C5741 vdd.n2985 gnd 0.007703f
C5742 vdd.n2986 gnd 0.007703f
C5743 vdd.n2987 gnd 0.006432f
C5744 vdd.n2988 gnd 0.00957f
C5745 vdd.n2990 gnd 0.00957f
C5746 vdd.n2992 gnd 0.00957f
C5747 vdd.n2993 gnd 0.006432f
C5748 vdd.n2994 gnd 0.007703f
C5749 vdd.n2995 gnd 0.007703f
C5750 vdd.n2996 gnd 0.00957f
C5751 vdd.n2998 gnd 0.00957f
C5752 vdd.n3000 gnd 0.00957f
C5753 vdd.n3001 gnd 0.007703f
C5754 vdd.n3002 gnd 0.007703f
C5755 vdd.n3003 gnd 0.007703f
C5756 vdd.n3004 gnd 0.00957f
C5757 vdd.n3006 gnd 0.00957f
C5758 vdd.n3008 gnd 0.00957f
C5759 vdd.n3009 gnd 0.007703f
C5760 vdd.n3010 gnd 0.007703f
C5761 vdd.n3011 gnd 0.007703f
C5762 vdd.n3012 gnd 0.00957f
C5763 vdd.n3014 gnd 0.00957f
C5764 vdd.n3015 gnd 0.00957f
C5765 vdd.n3016 gnd 0.007703f
C5766 vdd.n3017 gnd 0.007703f
C5767 vdd.n3018 gnd 0.00957f
C5768 vdd.n3019 gnd 0.00957f
C5769 vdd.n3020 gnd 0.007703f
C5770 vdd.n3021 gnd 0.007703f
C5771 vdd.n3022 gnd 0.00957f
C5772 vdd.n3023 gnd 0.00957f
C5773 vdd.n3025 gnd 0.00957f
C5774 vdd.n3026 gnd 0.007703f
C5775 vdd.n3027 gnd 0.006393f
C5776 vdd.n3028 gnd 0.022906f
C5777 vdd.n3029 gnd 0.022553f
C5778 vdd.n3030 gnd 0.006393f
C5779 vdd.n3031 gnd 0.022553f
C5780 vdd.n3032 gnd 1.34481f
C5781 vdd.n3033 gnd 0.022553f
C5782 vdd.n3034 gnd 0.006393f
C5783 vdd.n3035 gnd 0.022553f
C5784 vdd.n3036 gnd 0.00957f
C5785 vdd.n3037 gnd 0.00957f
C5786 vdd.n3038 gnd 0.007703f
C5787 vdd.n3039 gnd 0.00957f
C5788 vdd.n3040 gnd 0.978042f
C5789 vdd.n3041 gnd 0.00957f
C5790 vdd.n3042 gnd 0.007703f
C5791 vdd.n3043 gnd 0.00957f
C5792 vdd.n3044 gnd 0.00957f
C5793 vdd.n3045 gnd 0.00957f
C5794 vdd.n3046 gnd 0.007703f
C5795 vdd.n3047 gnd 0.00957f
C5796 vdd.n3048 gnd 0.865567f
C5797 vdd.n3049 gnd 0.00957f
C5798 vdd.n3050 gnd 0.007703f
C5799 vdd.n3051 gnd 0.00957f
C5800 vdd.n3052 gnd 0.00957f
C5801 vdd.n3053 gnd 0.00957f
C5802 vdd.n3054 gnd 0.007703f
C5803 vdd.n3055 gnd 0.00957f
C5804 vdd.t208 gnd 0.489021f
C5805 vdd.n3056 gnd 0.6993f
C5806 vdd.n3057 gnd 0.00957f
C5807 vdd.n3058 gnd 0.007703f
C5808 vdd.n3059 gnd 0.00957f
C5809 vdd.n3060 gnd 0.00957f
C5810 vdd.n3061 gnd 0.00957f
C5811 vdd.n3062 gnd 0.007703f
C5812 vdd.n3063 gnd 0.00957f
C5813 vdd.n3064 gnd 0.533033f
C5814 vdd.n3065 gnd 0.00957f
C5815 vdd.n3066 gnd 0.007703f
C5816 vdd.n3067 gnd 0.00957f
C5817 vdd.n3068 gnd 0.00957f
C5818 vdd.n3069 gnd 0.00957f
C5819 vdd.n3070 gnd 0.007703f
C5820 vdd.n3071 gnd 0.00957f
C5821 vdd.n3072 gnd 0.68952f
C5822 vdd.n3073 gnd 0.611276f
C5823 vdd.n3074 gnd 0.00957f
C5824 vdd.n3075 gnd 0.007703f
C5825 vdd.n3076 gnd 0.00957f
C5826 vdd.n3077 gnd 0.00957f
C5827 vdd.n3078 gnd 0.00957f
C5828 vdd.n3079 gnd 0.007703f
C5829 vdd.n3080 gnd 0.00957f
C5830 vdd.n3081 gnd 0.777544f
C5831 vdd.n3082 gnd 0.00957f
C5832 vdd.n3083 gnd 0.007703f
C5833 vdd.n3084 gnd 0.00957f
C5834 vdd.n3085 gnd 0.00957f
C5835 vdd.n3086 gnd 0.00957f
C5836 vdd.n3087 gnd 0.007703f
C5837 vdd.n3088 gnd 0.007703f
C5838 vdd.n3089 gnd 0.007703f
C5839 vdd.n3090 gnd 0.00957f
C5840 vdd.n3091 gnd 0.00957f
C5841 vdd.n3092 gnd 0.00957f
C5842 vdd.n3093 gnd 0.007703f
C5843 vdd.n3094 gnd 0.007703f
C5844 vdd.n3095 gnd 0.007703f
C5845 vdd.n3096 gnd 0.00957f
C5846 vdd.n3097 gnd 0.00957f
C5847 vdd.n3098 gnd 0.00957f
C5848 vdd.n3099 gnd 0.007703f
C5849 vdd.n3100 gnd 0.007703f
C5850 vdd.n3101 gnd 0.007703f
C5851 vdd.n3102 gnd 0.00957f
C5852 vdd.n3103 gnd 0.00957f
C5853 vdd.n3104 gnd 0.00957f
C5854 vdd.n3105 gnd 0.007703f
C5855 vdd.n3106 gnd 0.007703f
C5856 vdd.n3107 gnd 0.006393f
C5857 vdd.n3108 gnd 0.022553f
C5858 vdd.n3109 gnd 0.022906f
C5859 vdd.n3111 gnd 0.022906f
C5860 vdd.n3112 gnd 0.003659f
C5861 vdd.t50 gnd 0.11774f
C5862 vdd.t49 gnd 0.125832f
C5863 vdd.t47 gnd 0.153767f
C5864 vdd.n3113 gnd 0.197108f
C5865 vdd.n3114 gnd 0.166376f
C5866 vdd.n3115 gnd 0.012633f
C5867 vdd.n3116 gnd 0.004044f
C5868 vdd.n3117 gnd 0.007703f
C5869 vdd.n3118 gnd 0.00957f
C5870 vdd.n3120 gnd 0.00957f
C5871 vdd.n3121 gnd 0.00957f
C5872 vdd.n3122 gnd 0.007703f
C5873 vdd.n3123 gnd 0.007703f
C5874 vdd.n3124 gnd 0.007703f
C5875 vdd.n3125 gnd 0.00957f
C5876 vdd.n3127 gnd 0.00957f
C5877 vdd.n3128 gnd 0.00957f
C5878 vdd.n3129 gnd 0.007703f
C5879 vdd.n3130 gnd 0.007703f
C5880 vdd.n3131 gnd 0.007703f
C5881 vdd.n3132 gnd 0.00957f
C5882 vdd.n3134 gnd 0.00957f
C5883 vdd.n3135 gnd 0.00957f
C5884 vdd.n3136 gnd 0.007703f
C5885 vdd.n3137 gnd 0.007703f
C5886 vdd.n3138 gnd 0.007703f
C5887 vdd.n3139 gnd 0.00957f
C5888 vdd.n3141 gnd 0.00957f
C5889 vdd.n3142 gnd 0.00957f
C5890 vdd.n3143 gnd 0.007703f
C5891 vdd.n3144 gnd 0.007703f
C5892 vdd.n3145 gnd 0.007703f
C5893 vdd.n3146 gnd 0.00957f
C5894 vdd.n3148 gnd 0.00957f
C5895 vdd.n3149 gnd 0.00957f
C5896 vdd.n3150 gnd 0.007703f
C5897 vdd.n3151 gnd 0.00957f
C5898 vdd.n3152 gnd 0.00957f
C5899 vdd.n3153 gnd 0.00957f
C5900 vdd.n3154 gnd 0.016484f
C5901 vdd.n3155 gnd 0.005238f
C5902 vdd.n3156 gnd 0.007703f
C5903 vdd.n3157 gnd 0.00957f
C5904 vdd.n3159 gnd 0.00957f
C5905 vdd.n3160 gnd 0.00957f
C5906 vdd.n3161 gnd 0.007703f
C5907 vdd.n3162 gnd 0.007703f
C5908 vdd.n3163 gnd 0.007703f
C5909 vdd.n3164 gnd 0.00957f
C5910 vdd.n3166 gnd 0.00957f
C5911 vdd.n3167 gnd 0.00957f
C5912 vdd.n3168 gnd 0.007703f
C5913 vdd.n3169 gnd 0.007703f
C5914 vdd.n3170 gnd 0.007703f
C5915 vdd.n3171 gnd 0.00957f
C5916 vdd.n3173 gnd 0.00957f
C5917 vdd.n3174 gnd 0.00957f
C5918 vdd.n3175 gnd 0.007703f
C5919 vdd.n3176 gnd 0.007703f
C5920 vdd.n3177 gnd 0.007703f
C5921 vdd.n3178 gnd 0.00957f
C5922 vdd.n3180 gnd 0.00957f
C5923 vdd.n3181 gnd 0.00957f
C5924 vdd.n3182 gnd 0.007703f
C5925 vdd.n3183 gnd 0.007703f
C5926 vdd.n3184 gnd 0.007703f
C5927 vdd.n3185 gnd 0.00957f
C5928 vdd.n3187 gnd 0.00957f
C5929 vdd.n3188 gnd 0.00957f
C5930 vdd.n3189 gnd 0.007703f
C5931 vdd.n3190 gnd 0.00957f
C5932 vdd.n3191 gnd 0.00957f
C5933 vdd.n3192 gnd 0.00957f
C5934 vdd.n3193 gnd 0.016484f
C5935 vdd.n3194 gnd 0.006432f
C5936 vdd.n3195 gnd 0.007703f
C5937 vdd.n3196 gnd 0.00957f
C5938 vdd.n3198 gnd 0.00957f
C5939 vdd.n3199 gnd 0.00957f
C5940 vdd.n3200 gnd 0.007703f
C5941 vdd.n3201 gnd 0.007703f
C5942 vdd.n3202 gnd 0.007703f
C5943 vdd.n3203 gnd 0.00957f
C5944 vdd.n3205 gnd 0.00957f
C5945 vdd.n3206 gnd 0.00957f
C5946 vdd.n3207 gnd 0.007703f
C5947 vdd.n3208 gnd 0.007703f
C5948 vdd.n3209 gnd 0.007703f
C5949 vdd.n3210 gnd 0.00957f
C5950 vdd.n3212 gnd 0.00957f
C5951 vdd.n3213 gnd 0.00957f
C5952 vdd.n3214 gnd 0.007703f
C5953 vdd.n3215 gnd 0.007703f
C5954 vdd.n3216 gnd 0.007703f
C5955 vdd.n3217 gnd 0.00957f
C5956 vdd.n3219 gnd 0.00957f
C5957 vdd.n3220 gnd 0.00957f
C5958 vdd.n3222 gnd 0.00957f
C5959 vdd.n3223 gnd 0.007703f
C5960 vdd.n3224 gnd 0.007703f
C5961 vdd.n3225 gnd 0.006393f
C5962 vdd.n3226 gnd 0.022906f
C5963 vdd.n3227 gnd 0.022553f
C5964 vdd.n3228 gnd 0.006393f
C5965 vdd.n3229 gnd 0.022553f
C5966 vdd.n3230 gnd 1.37904f
C5967 vdd.n3231 gnd 0.552594f
C5968 vdd.t48 gnd 0.489021f
C5969 vdd.n3232 gnd 0.914469f
C5970 vdd.n3233 gnd 0.00957f
C5971 vdd.n3234 gnd 0.007703f
C5972 vdd.n3235 gnd 0.007703f
C5973 vdd.n3236 gnd 0.007703f
C5974 vdd.n3237 gnd 0.00957f
C5975 vdd.n3238 gnd 0.963372f
C5976 vdd.t159 gnd 0.489021f
C5977 vdd.n3239 gnd 0.503692f
C5978 vdd.n3240 gnd 0.797104f
C5979 vdd.n3241 gnd 0.00957f
C5980 vdd.n3242 gnd 0.007703f
C5981 vdd.n3243 gnd 0.007703f
C5982 vdd.n3244 gnd 0.007703f
C5983 vdd.n3245 gnd 0.00957f
C5984 vdd.n3246 gnd 0.630837f
C5985 vdd.t174 gnd 0.489021f
C5986 vdd.n3247 gnd 0.811775f
C5987 vdd.t194 gnd 0.489021f
C5988 vdd.n3248 gnd 0.513472f
C5989 vdd.n3249 gnd 0.00957f
C5990 vdd.n3250 gnd 0.007703f
C5991 vdd.n3251 gnd 0.007703f
C5992 vdd.n3252 gnd 0.007703f
C5993 vdd.n3253 gnd 0.00957f
C5994 vdd.n3254 gnd 0.679739f
C5995 vdd.n3255 gnd 0.621057f
C5996 vdd.t171 gnd 0.489021f
C5997 vdd.n3256 gnd 0.811775f
C5998 vdd.n3257 gnd 0.00957f
C5999 vdd.n3258 gnd 0.007703f
C6000 vdd.n3259 gnd 0.5697f
C6001 vdd.n3260 gnd 2.22459f
C6002 a_n6972_8799.n0 gnd 3.87083f
C6003 a_n6972_8799.n1 gnd 1.92936f
C6004 a_n6972_8799.n2 gnd 3.25853f
C6005 a_n6972_8799.n3 gnd 0.793559f
C6006 a_n6972_8799.n4 gnd 0.178461f
C6007 a_n6972_8799.n5 gnd 0.208989f
C6008 a_n6972_8799.n6 gnd 0.208989f
C6009 a_n6972_8799.n7 gnd 0.208989f
C6010 a_n6972_8799.n8 gnd 0.178461f
C6011 a_n6972_8799.n9 gnd 0.208989f
C6012 a_n6972_8799.n10 gnd 0.208989f
C6013 a_n6972_8799.n11 gnd 0.208989f
C6014 a_n6972_8799.n12 gnd 0.344724f
C6015 a_n6972_8799.n13 gnd 0.208989f
C6016 a_n6972_8799.n14 gnd 0.208989f
C6017 a_n6972_8799.n15 gnd 0.208989f
C6018 a_n6972_8799.n16 gnd 0.208989f
C6019 a_n6972_8799.n17 gnd 0.208989f
C6020 a_n6972_8799.n18 gnd 0.178461f
C6021 a_n6972_8799.n19 gnd 0.208989f
C6022 a_n6972_8799.n20 gnd 0.208989f
C6023 a_n6972_8799.n21 gnd 0.208989f
C6024 a_n6972_8799.n22 gnd 0.178461f
C6025 a_n6972_8799.n23 gnd 0.208989f
C6026 a_n6972_8799.n24 gnd 0.208989f
C6027 a_n6972_8799.n25 gnd 0.208989f
C6028 a_n6972_8799.n26 gnd 0.344724f
C6029 a_n6972_8799.n27 gnd 0.208989f
C6030 a_n6972_8799.n28 gnd 1.53172f
C6031 a_n6972_8799.n29 gnd 2.5338f
C6032 a_n6972_8799.n30 gnd 0.252736f
C6033 a_n6972_8799.n32 gnd 0.007784f
C6034 a_n6972_8799.n33 gnd 0.011766f
C6035 a_n6972_8799.n34 gnd 0.008091f
C6036 a_n6972_8799.n36 gnd 4.04e-19
C6037 a_n6972_8799.n37 gnd 0.008386f
C6038 a_n6972_8799.n38 gnd 0.264392f
C6039 a_n6972_8799.n39 gnd 0.252736f
C6040 a_n6972_8799.n41 gnd 0.007784f
C6041 a_n6972_8799.n42 gnd 0.011766f
C6042 a_n6972_8799.n43 gnd 0.008091f
C6043 a_n6972_8799.n45 gnd 4.04e-19
C6044 a_n6972_8799.n46 gnd 0.008386f
C6045 a_n6972_8799.n47 gnd 0.264392f
C6046 a_n6972_8799.n48 gnd 0.252736f
C6047 a_n6972_8799.n50 gnd 0.007784f
C6048 a_n6972_8799.n51 gnd 0.011766f
C6049 a_n6972_8799.n52 gnd 0.008091f
C6050 a_n6972_8799.n54 gnd 4.04e-19
C6051 a_n6972_8799.n55 gnd 0.008386f
C6052 a_n6972_8799.n56 gnd 0.264392f
C6053 a_n6972_8799.n57 gnd 0.008386f
C6054 a_n6972_8799.n58 gnd 0.264392f
C6055 a_n6972_8799.n59 gnd 4.04e-19
C6056 a_n6972_8799.n61 gnd 0.008091f
C6057 a_n6972_8799.n62 gnd 0.011766f
C6058 a_n6972_8799.n63 gnd 0.007784f
C6059 a_n6972_8799.n65 gnd 0.252736f
C6060 a_n6972_8799.n66 gnd 0.008386f
C6061 a_n6972_8799.n67 gnd 0.264392f
C6062 a_n6972_8799.n68 gnd 4.04e-19
C6063 a_n6972_8799.n70 gnd 0.008091f
C6064 a_n6972_8799.n71 gnd 0.011766f
C6065 a_n6972_8799.n72 gnd 0.007784f
C6066 a_n6972_8799.n74 gnd 0.252736f
C6067 a_n6972_8799.n75 gnd 0.008386f
C6068 a_n6972_8799.n76 gnd 0.264392f
C6069 a_n6972_8799.n77 gnd 4.04e-19
C6070 a_n6972_8799.n79 gnd 0.008091f
C6071 a_n6972_8799.n80 gnd 0.011766f
C6072 a_n6972_8799.n81 gnd 0.007784f
C6073 a_n6972_8799.n83 gnd 0.252736f
C6074 a_n6972_8799.t6 gnd 0.144957f
C6075 a_n6972_8799.t37 gnd 0.144957f
C6076 a_n6972_8799.t33 gnd 0.144957f
C6077 a_n6972_8799.n84 gnd 1.1433f
C6078 a_n6972_8799.t36 gnd 0.144957f
C6079 a_n6972_8799.t18 gnd 0.144957f
C6080 a_n6972_8799.n85 gnd 1.14329f
C6081 a_n6972_8799.t39 gnd 0.144957f
C6082 a_n6972_8799.t32 gnd 0.144957f
C6083 a_n6972_8799.n86 gnd 1.14141f
C6084 a_n6972_8799.t19 gnd 0.144957f
C6085 a_n6972_8799.t31 gnd 0.144957f
C6086 a_n6972_8799.n87 gnd 1.14141f
C6087 a_n6972_8799.t29 gnd 0.144957f
C6088 a_n6972_8799.t5 gnd 0.144957f
C6089 a_n6972_8799.n88 gnd 1.14141f
C6090 a_n6972_8799.n89 gnd 3.23927f
C6091 a_n6972_8799.t2 gnd 0.112744f
C6092 a_n6972_8799.t7 gnd 0.112744f
C6093 a_n6972_8799.n90 gnd 0.998463f
C6094 a_n6972_8799.t9 gnd 0.112744f
C6095 a_n6972_8799.t21 gnd 0.112744f
C6096 a_n6972_8799.n91 gnd 0.996248f
C6097 a_n6972_8799.t20 gnd 0.112744f
C6098 a_n6972_8799.t11 gnd 0.112744f
C6099 a_n6972_8799.n92 gnd 0.996248f
C6100 a_n6972_8799.t14 gnd 0.112744f
C6101 a_n6972_8799.t16 gnd 0.112744f
C6102 a_n6972_8799.n93 gnd 0.998462f
C6103 a_n6972_8799.t24 gnd 0.112744f
C6104 a_n6972_8799.t8 gnd 0.112744f
C6105 a_n6972_8799.n94 gnd 0.996247f
C6106 a_n6972_8799.t10 gnd 0.112744f
C6107 a_n6972_8799.t3 gnd 0.112744f
C6108 a_n6972_8799.n95 gnd 0.996247f
C6109 a_n6972_8799.t26 gnd 0.112744f
C6110 a_n6972_8799.t0 gnd 0.112744f
C6111 a_n6972_8799.n96 gnd 0.998462f
C6112 a_n6972_8799.t22 gnd 0.112744f
C6113 a_n6972_8799.t1 gnd 0.112744f
C6114 a_n6972_8799.n97 gnd 0.996247f
C6115 a_n6972_8799.t28 gnd 0.112744f
C6116 a_n6972_8799.t15 gnd 0.112744f
C6117 a_n6972_8799.n98 gnd 0.996247f
C6118 a_n6972_8799.t38 gnd 0.112744f
C6119 a_n6972_8799.t13 gnd 0.112744f
C6120 a_n6972_8799.n99 gnd 0.996248f
C6121 a_n6972_8799.t27 gnd 0.112744f
C6122 a_n6972_8799.t23 gnd 0.112744f
C6123 a_n6972_8799.n100 gnd 0.996248f
C6124 a_n6972_8799.t12 gnd 0.112744f
C6125 a_n6972_8799.t25 gnd 0.112744f
C6126 a_n6972_8799.n101 gnd 0.996248f
C6127 a_n6972_8799.t72 gnd 0.601059f
C6128 a_n6972_8799.n102 gnd 0.272033f
C6129 a_n6972_8799.t100 gnd 0.601059f
C6130 a_n6972_8799.t40 gnd 0.601059f
C6131 a_n6972_8799.n103 gnd 0.263129f
C6132 a_n6972_8799.t61 gnd 0.601059f
C6133 a_n6972_8799.n104 gnd 0.274581f
C6134 a_n6972_8799.t62 gnd 0.601059f
C6135 a_n6972_8799.t69 gnd 0.601059f
C6136 a_n6972_8799.n105 gnd 0.267961f
C6137 a_n6972_8799.t99 gnd 0.615185f
C6138 a_n6972_8799.t68 gnd 0.601059f
C6139 a_n6972_8799.n106 gnd 0.274143f
C6140 a_n6972_8799.n107 gnd 0.250554f
C6141 a_n6972_8799.t86 gnd 0.601059f
C6142 a_n6972_8799.n108 gnd 0.271915f
C6143 a_n6972_8799.n109 gnd 0.272048f
C6144 a_n6972_8799.t85 gnd 0.601059f
C6145 a_n6972_8799.n110 gnd 0.268283f
C6146 a_n6972_8799.t60 gnd 0.601059f
C6147 a_n6972_8799.n111 gnd 0.268535f
C6148 a_n6972_8799.n112 gnd 0.274144f
C6149 a_n6972_8799.t48 gnd 0.611971f
C6150 a_n6972_8799.t79 gnd 0.601059f
C6151 a_n6972_8799.n113 gnd 0.272033f
C6152 a_n6972_8799.t110 gnd 0.601059f
C6153 a_n6972_8799.t47 gnd 0.601059f
C6154 a_n6972_8799.n114 gnd 0.263129f
C6155 a_n6972_8799.t66 gnd 0.601059f
C6156 a_n6972_8799.n115 gnd 0.274581f
C6157 a_n6972_8799.t67 gnd 0.601059f
C6158 a_n6972_8799.t74 gnd 0.601059f
C6159 a_n6972_8799.n116 gnd 0.267961f
C6160 a_n6972_8799.t108 gnd 0.615185f
C6161 a_n6972_8799.t73 gnd 0.601059f
C6162 a_n6972_8799.n117 gnd 0.274143f
C6163 a_n6972_8799.n118 gnd 0.250554f
C6164 a_n6972_8799.t98 gnd 0.601059f
C6165 a_n6972_8799.n119 gnd 0.271915f
C6166 a_n6972_8799.n120 gnd 0.272048f
C6167 a_n6972_8799.t94 gnd 0.601059f
C6168 a_n6972_8799.n121 gnd 0.268283f
C6169 a_n6972_8799.t65 gnd 0.601059f
C6170 a_n6972_8799.n122 gnd 0.268535f
C6171 a_n6972_8799.n123 gnd 0.274144f
C6172 a_n6972_8799.t57 gnd 0.611971f
C6173 a_n6972_8799.n124 gnd 0.902354f
C6174 a_n6972_8799.t81 gnd 0.601059f
C6175 a_n6972_8799.n125 gnd 0.272033f
C6176 a_n6972_8799.t55 gnd 0.601059f
C6177 a_n6972_8799.t71 gnd 0.601059f
C6178 a_n6972_8799.n126 gnd 0.263129f
C6179 a_n6972_8799.t104 gnd 0.601059f
C6180 a_n6972_8799.n127 gnd 0.274581f
C6181 a_n6972_8799.t87 gnd 0.601059f
C6182 a_n6972_8799.t41 gnd 0.601059f
C6183 a_n6972_8799.n128 gnd 0.267961f
C6184 a_n6972_8799.t101 gnd 0.615185f
C6185 a_n6972_8799.t52 gnd 0.601059f
C6186 a_n6972_8799.n129 gnd 0.274143f
C6187 a_n6972_8799.n130 gnd 0.250554f
C6188 a_n6972_8799.t75 gnd 0.601059f
C6189 a_n6972_8799.n131 gnd 0.271915f
C6190 a_n6972_8799.n132 gnd 0.272048f
C6191 a_n6972_8799.t107 gnd 0.601059f
C6192 a_n6972_8799.n133 gnd 0.268283f
C6193 a_n6972_8799.t45 gnd 0.601059f
C6194 a_n6972_8799.n134 gnd 0.268535f
C6195 a_n6972_8799.n135 gnd 0.274144f
C6196 a_n6972_8799.t95 gnd 0.611971f
C6197 a_n6972_8799.n136 gnd 1.62811f
C6198 a_n6972_8799.t70 gnd 0.611971f
C6199 a_n6972_8799.t58 gnd 0.601059f
C6200 a_n6972_8799.t103 gnd 0.601059f
C6201 a_n6972_8799.t80 gnd 0.601059f
C6202 a_n6972_8799.n137 gnd 0.268535f
C6203 a_n6972_8799.t78 gnd 0.601059f
C6204 a_n6972_8799.t42 gnd 0.601059f
C6205 a_n6972_8799.t84 gnd 0.601059f
C6206 a_n6972_8799.n138 gnd 0.272048f
C6207 a_n6972_8799.t83 gnd 0.601059f
C6208 a_n6972_8799.t44 gnd 0.601059f
C6209 a_n6972_8799.t43 gnd 0.601059f
C6210 a_n6972_8799.n139 gnd 0.267961f
C6211 a_n6972_8799.t54 gnd 0.615185f
C6212 a_n6972_8799.t97 gnd 0.601059f
C6213 a_n6972_8799.n140 gnd 0.274143f
C6214 a_n6972_8799.n141 gnd 0.250554f
C6215 a_n6972_8799.n142 gnd 0.271915f
C6216 a_n6972_8799.n143 gnd 0.274581f
C6217 a_n6972_8799.n144 gnd 0.268283f
C6218 a_n6972_8799.n145 gnd 0.263129f
C6219 a_n6972_8799.n146 gnd 0.272033f
C6220 a_n6972_8799.n147 gnd 0.274144f
C6221 a_n6972_8799.t77 gnd 0.611971f
C6222 a_n6972_8799.t64 gnd 0.601059f
C6223 a_n6972_8799.t111 gnd 0.601059f
C6224 a_n6972_8799.t90 gnd 0.601059f
C6225 a_n6972_8799.n148 gnd 0.268535f
C6226 a_n6972_8799.t89 gnd 0.601059f
C6227 a_n6972_8799.t49 gnd 0.601059f
C6228 a_n6972_8799.t93 gnd 0.601059f
C6229 a_n6972_8799.n149 gnd 0.272048f
C6230 a_n6972_8799.t92 gnd 0.601059f
C6231 a_n6972_8799.t51 gnd 0.601059f
C6232 a_n6972_8799.t50 gnd 0.601059f
C6233 a_n6972_8799.n150 gnd 0.267961f
C6234 a_n6972_8799.t63 gnd 0.615185f
C6235 a_n6972_8799.t106 gnd 0.601059f
C6236 a_n6972_8799.n151 gnd 0.274143f
C6237 a_n6972_8799.n152 gnd 0.250554f
C6238 a_n6972_8799.n153 gnd 0.271915f
C6239 a_n6972_8799.n154 gnd 0.274581f
C6240 a_n6972_8799.n155 gnd 0.268283f
C6241 a_n6972_8799.n156 gnd 0.263129f
C6242 a_n6972_8799.n157 gnd 0.272033f
C6243 a_n6972_8799.n158 gnd 0.274144f
C6244 a_n6972_8799.n159 gnd 0.902354f
C6245 a_n6972_8799.t96 gnd 0.611971f
C6246 a_n6972_8799.t56 gnd 0.601059f
C6247 a_n6972_8799.t82 gnd 0.601059f
C6248 a_n6972_8799.t46 gnd 0.601059f
C6249 a_n6972_8799.n160 gnd 0.268535f
C6250 a_n6972_8799.t59 gnd 0.601059f
C6251 a_n6972_8799.t109 gnd 0.601059f
C6252 a_n6972_8799.t88 gnd 0.601059f
C6253 a_n6972_8799.n161 gnd 0.272048f
C6254 a_n6972_8799.t105 gnd 0.601059f
C6255 a_n6972_8799.t76 gnd 0.601059f
C6256 a_n6972_8799.t91 gnd 0.601059f
C6257 a_n6972_8799.n162 gnd 0.267961f
C6258 a_n6972_8799.t102 gnd 0.615185f
C6259 a_n6972_8799.t53 gnd 0.601059f
C6260 a_n6972_8799.n163 gnd 0.274143f
C6261 a_n6972_8799.n164 gnd 0.250554f
C6262 a_n6972_8799.n165 gnd 0.271915f
C6263 a_n6972_8799.n166 gnd 0.274581f
C6264 a_n6972_8799.n167 gnd 0.268283f
C6265 a_n6972_8799.n168 gnd 0.263129f
C6266 a_n6972_8799.n169 gnd 0.272033f
C6267 a_n6972_8799.n170 gnd 0.274144f
C6268 a_n6972_8799.n171 gnd 1.19276f
C6269 a_n6972_8799.n172 gnd 14.0386f
C6270 a_n6972_8799.n173 gnd 4.39888f
C6271 a_n6972_8799.n174 gnd 6.37523f
C6272 a_n6972_8799.t35 gnd 0.144957f
C6273 a_n6972_8799.t17 gnd 0.144957f
C6274 a_n6972_8799.n175 gnd 1.14141f
C6275 a_n6972_8799.t34 gnd 0.144957f
C6276 a_n6972_8799.t30 gnd 0.144957f
C6277 a_n6972_8799.n176 gnd 1.14141f
C6278 a_n6972_8799.n177 gnd 1.02599f
C6279 a_n6972_8799.n178 gnd 1.14141f
C6280 a_n6972_8799.t4 gnd 0.144957f
.ends

