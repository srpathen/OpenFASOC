* NGSPICE file created from opamp265.ext - technology: sky130A

.subckt opamp265 gnd CSoutput output vdd plus minus commonsourceibias outputibias
+ diffpairibias
X0 a_n2472_13878.t23 a_n2650_13878.t39 a_n2650_13878.t40 vdd.t213 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X1 CSoutput.t85 a_n7636_8799.t36 vdd.t5 vdd.t4 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=3.12 ps=16.78 w=8 l=0.5
X2 a_n2472_13878.t26 a_n2650_13878.t56 vdd.t225 vdd.t224 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X3 vdd.t7 a_n7636_8799.t37 CSoutput.t84 vdd.t6 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X4 gnd.t263 commonsourceibias.t20 commonsourceibias.t21 gnd.t201 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X5 a_n7636_8799.t35 plus.t5 a_n3827_n3924.t24 gnd.t310 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.9
X6 commonsourceibias.t19 commonsourceibias.t18 gnd.t262 gnd.t162 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X7 CSoutput.t83 a_n7636_8799.t38 vdd.t34 vdd.t33 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X8 a_n3827_n3924.t38 diffpairibias.t20 gnd.t318 gnd.t317 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=2.73 ps=14.78 w=7 l=1
X9 minus.t4 gnd.t139 gnd.t141 gnd.t140 sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.5
X10 vdd.t169 vdd.t167 vdd.t168 vdd.t125 sky130_fd_pr__pfet_01v8 ad=3.12 pd=16.78 as=0 ps=0 w=8 l=0.5
X11 a_n2650_8322.t25 a_n2650_13878.t57 a_n7636_8799.t14 vdd.t222 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X12 gnd.t261 commonsourceibias.t16 commonsourceibias.t17 gnd.t148 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X13 gnd.t260 commonsourceibias.t48 CSoutput.t131 gnd.t196 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X14 commonsourceibias.t15 commonsourceibias.t14 gnd.t259 gnd.t170 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X15 CSoutput.t82 a_n7636_8799.t39 vdd.t36 vdd.t35 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X16 vdd.t71 a_n7636_8799.t40 CSoutput.t81 vdd.t18 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X17 output.t19 outputibias.t8 gnd.t10 gnd.t9 sky130_fd_pr__nfet_01v8 ad=2.34 pd=12.78 as=2.34 ps=12.78 w=6 l=2
X18 gnd.t138 gnd.t136 gnd.t137 gnd.t60 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=0 ps=0 w=7 l=1
X19 a_n7636_8799.t20 a_n2650_13878.t58 a_n2650_8322.t24 vdd.t211 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X20 a_n2650_13878.t10 minus.t5 a_n3827_n3924.t34 gnd.t308 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.9
X21 a_n7636_8799.t8 plus.t6 a_n3827_n3924.t23 gnd.t314 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.9
X22 a_n2650_13878.t54 minus.t6 a_n3827_n3924.t40 gnd.t313 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.9
X23 vdd.t72 a_n7636_8799.t41 CSoutput.t80 vdd.t21 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X24 a_n7636_8799.t26 a_n2650_13878.t59 a_n2650_8322.t23 vdd.t175 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=3.51 ps=18.78 w=9 l=0.5
X25 commonsourceibias.t13 commonsourceibias.t12 gnd.t258 gnd.t199 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X26 gnd.t257 commonsourceibias.t49 CSoutput.t102 gnd.t156 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X27 CSoutput.t117 commonsourceibias.t50 gnd.t256 gnd.t168 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X28 gnd.t135 gnd.t132 gnd.t134 gnd.t133 sky130_fd_pr__nfet_01v8 ad=1.95 pd=10.78 as=0 ps=0 w=5 l=1
X29 gnd.t131 gnd.t128 gnd.t130 gnd.t129 sky130_fd_pr__nfet_01v8 ad=2.34 pd=12.78 as=0 ps=0 w=6 l=2
X30 CSoutput.t79 a_n7636_8799.t42 vdd.t75 vdd.t4 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=3.12 ps=16.78 w=8 l=0.5
X31 a_n3827_n3924.t22 plus.t7 a_n7636_8799.t1 gnd.t302 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=1.155 ps=7.33 w=7 l=0.9
X32 gnd.t254 commonsourceibias.t36 commonsourceibias.t37 gnd.t196 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X33 a_n3827_n3924.t1 minus.t7 a_n2650_13878.t1 gnd.t1 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.9
X34 a_n3827_n3924.t6 diffpairibias.t21 gnd.t15 gnd.t14 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=2.73 ps=14.78 w=7 l=1
X35 commonsourceibias.t39 commonsourceibias.t38 gnd.t255 gnd.t150 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=2.73 ps=14.78 w=7 l=1
X36 CSoutput.t78 a_n7636_8799.t43 vdd.t76 vdd.t33 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X37 vdd.t166 vdd.t164 vdd.t165 vdd.t103 sky130_fd_pr__pfet_01v8 ad=3.51 pd=18.78 as=0 ps=0 w=9 l=0.5
X38 CSoutput.t87 commonsourceibias.t51 gnd.t253 gnd.t158 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=2.73 ps=14.78 w=7 l=1
X39 gnd.t252 commonsourceibias.t34 commonsourceibias.t35 gnd.t188 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X40 a_n2472_13878.t22 a_n2650_13878.t23 a_n2650_13878.t24 vdd.t183 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X41 a_n2650_13878.t18 a_n2650_13878.t17 a_n2472_13878.t21 vdd.t194 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X42 vdd.t163 vdd.t161 vdd.t162 vdd.t125 sky130_fd_pr__pfet_01v8 ad=3.12 pd=16.78 as=0 ps=0 w=8 l=0.5
X43 CSoutput.t77 a_n7636_8799.t44 vdd.t234 vdd.t35 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X44 gnd.t127 gnd.t125 plus.t4 gnd.t126 sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.39 ps=2.78 w=1 l=0.5
X45 output.t18 outputibias.t9 gnd.t269 gnd.t268 sky130_fd_pr__nfet_01v8 ad=2.34 pd=12.78 as=2.34 ps=12.78 w=6 l=2
X46 vdd.t160 vdd.t158 vdd.t159 vdd.t141 sky130_fd_pr__pfet_01v8 ad=3.51 pd=18.78 as=0 ps=0 w=9 l=0.5
X47 vdd.t235 a_n7636_8799.t45 CSoutput.t76 vdd.t18 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X48 a_n3827_n3924.t21 plus.t8 a_n7636_8799.t34 gnd.t304 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.9
X49 diffpairibias.t19 diffpairibias.t18 gnd.t316 gnd.t315 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=2.73 ps=14.78 w=7 l=1
X50 a_n2650_13878.t22 a_n2650_13878.t21 a_n2472_13878.t20 vdd.t208 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X51 a_n7636_8799.t16 a_n2650_13878.t60 a_n2650_8322.t22 vdd.t203 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X52 vdd.t60 a_n7636_8799.t46 CSoutput.t75 vdd.t21 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X53 vdd.t61 a_n7636_8799.t47 CSoutput.t74 vdd.t10 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X54 a_n2650_13878.t28 a_n2650_13878.t27 a_n2472_13878.t19 vdd.t223 sky130_fd_pr__pfet_01v8 ad=3.51 pd=18.78 as=1.485 ps=9.33 w=9 l=0.5
X55 CSoutput.t73 a_n7636_8799.t48 vdd.t84 vdd.t49 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X56 CSoutput.t120 commonsourceibias.t52 gnd.t251 gnd.t190 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X57 gnd.t124 gnd.t122 gnd.t123 gnd.t31 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=0 ps=0 w=7 l=1
X58 CSoutput.t125 commonsourceibias.t53 gnd.t250 gnd.t211 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X59 a_n7636_8799.t24 a_n2650_13878.t61 a_n2650_8322.t21 vdd.t202 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=3.51 ps=18.78 w=9 l=0.5
X60 diffpairibias.t17 diffpairibias.t16 gnd.t323 gnd.t322 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=2.73 ps=14.78 w=7 l=1
X61 CSoutput.t72 a_n7636_8799.t49 vdd.t85 vdd.t27 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X62 gnd.t121 gnd.t119 gnd.t120 gnd.t31 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=0 ps=0 w=7 l=1
X63 CSoutput.t144 a_n2650_8322.t5 sky130_fd_pr__cap_mim_m3_1 l=12 w=12
X64 a_n2650_8322.t20 a_n2650_13878.t62 a_n7636_8799.t29 vdd.t223 sky130_fd_pr__pfet_01v8 ad=3.51 pd=18.78 as=1.485 ps=9.33 w=9 l=0.5
X65 CSoutput.t90 commonsourceibias.t54 gnd.t249 gnd.t190 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X66 CSoutput.t71 a_n7636_8799.t50 vdd.t1 vdd.t0 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=3.12 ps=16.78 w=8 l=0.5
X67 a_n3827_n3924.t5 minus.t8 a_n2650_13878.t3 gnd.t13 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.9
X68 a_n3827_n3924.t20 plus.t9 a_n7636_8799.t0 gnd.t4 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=1.155 ps=7.33 w=7 l=0.9
X69 gnd.t248 commonsourceibias.t55 CSoutput.t91 gnd.t176 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=1.155 ps=7.33 w=7 l=1
X70 output.t15 CSoutput.t145 vdd.t8 gnd.t287 sky130_fd_pr__nfet_01v8 ad=0.825 pd=5.33 as=0.825 ps=5.33 w=5 l=1
X71 gnd.t247 commonsourceibias.t56 CSoutput.t104 gnd.t164 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=1.155 ps=7.33 w=7 l=1
X72 CSoutput.t106 commonsourceibias.t57 gnd.t246 gnd.t185 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X73 CSoutput.t146 a_n2650_8322.t4 sky130_fd_pr__cap_mim_m3_1 l=12 w=12
X74 gnd.t118 gnd.t116 gnd.t117 gnd.t60 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=0 ps=0 w=7 l=1
X75 vdd.t3 a_n7636_8799.t51 CSoutput.t70 vdd.t2 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X76 a_n3827_n3924.t37 diffpairibias.t22 gnd.t312 gnd.t311 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=2.73 ps=14.78 w=7 l=1
X77 vdd.t15 a_n7636_8799.t52 CSoutput.t69 vdd.t14 sky130_fd_pr__pfet_01v8 ad=3.12 pd=16.78 as=1.32 ps=8.33 w=8 l=0.5
X78 a_n7636_8799.t15 a_n2650_13878.t63 a_n2650_8322.t19 vdd.t212 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X79 a_n2650_13878.t36 a_n2650_13878.t35 a_n2472_13878.t18 vdd.t222 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X80 a_n3827_n3924.t19 plus.t10 a_n7636_8799.t7 gnd.t299 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.9
X81 CSoutput.t133 commonsourceibias.t58 gnd.t245 gnd.t152 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X82 a_n2650_13878.t26 a_n2650_13878.t25 a_n2472_13878.t17 vdd.t178 sky130_fd_pr__pfet_01v8 ad=3.51 pd=18.78 as=1.485 ps=9.33 w=9 l=0.5
X83 outputibias.t7 outputibias.t6 gnd.t6 gnd.t5 sky130_fd_pr__nfet_01v8 ad=2.34 pd=12.78 as=2.34 ps=12.78 w=6 l=2
X84 CSoutput.t137 commonsourceibias.t59 gnd.t244 gnd.t162 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X85 gnd.t243 commonsourceibias.t60 CSoutput.t99 gnd.t174 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X86 commonsourceibias.t5 commonsourceibias.t4 gnd.t242 gnd.t168 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X87 CSoutput.t68 a_n7636_8799.t53 vdd.t17 vdd.t16 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X88 vdd.t73 a_n7636_8799.t54 CSoutput.t67 vdd.t47 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X89 gnd.t115 gnd.t113 gnd.t114 gnd.t56 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=0 ps=0 w=7 l=1
X90 diffpairibias.t15 diffpairibias.t14 gnd.t289 gnd.t288 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=2.73 ps=14.78 w=7 l=1
X91 outputibias.t5 outputibias.t4 gnd.t291 gnd.t290 sky130_fd_pr__nfet_01v8 ad=2.34 pd=12.78 as=2.34 ps=12.78 w=6 l=2
X92 CSoutput.t66 a_n7636_8799.t55 vdd.t74 vdd.t27 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X93 vdd.t157 vdd.t155 vdd.t156 vdd.t145 sky130_fd_pr__pfet_01v8 ad=3.51 pd=18.78 as=0 ps=0 w=9 l=0.5
X94 vdd.t154 vdd.t151 vdd.t153 vdd.t152 sky130_fd_pr__pfet_01v8 ad=3.51 pd=18.78 as=0 ps=0 w=9 l=0.5
X95 vdd.t150 vdd.t148 vdd.t149 vdd.t117 sky130_fd_pr__pfet_01v8 ad=3.12 pd=16.78 as=0 ps=0 w=8 l=0.5
X96 a_n2650_8322.t33 a_n2650_13878.t64 vdd.t221 vdd.t220 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X97 vdd.t219 a_n2650_13878.t65 a_n2650_8322.t32 vdd.t218 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X98 a_n2650_13878.t52 a_n2650_13878.t51 a_n2472_13878.t16 vdd.t186 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X99 gnd.t112 gnd.t110 minus.t3 gnd.t111 sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.39 ps=2.78 w=1 l=0.5
X100 CSoutput.t139 commonsourceibias.t61 gnd.t241 gnd.t199 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X101 output.t14 CSoutput.t147 vdd.t9 gnd.t286 sky130_fd_pr__nfet_01v8 ad=0.825 pd=5.33 as=0.825 ps=5.33 w=5 l=1
X102 gnd.t240 commonsourceibias.t10 commonsourceibias.t11 gnd.t160 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X103 CSoutput.t65 a_n7636_8799.t56 vdd.t46 vdd.t0 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=3.12 ps=16.78 w=8 l=0.5
X104 gnd.t239 commonsourceibias.t62 CSoutput.t86 gnd.t201 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X105 a_n3827_n3924.t29 diffpairibias.t23 gnd.t301 gnd.t300 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=2.73 ps=14.78 w=7 l=1
X106 gnd.t109 gnd.t107 gnd.t108 gnd.t52 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=0 ps=0 w=7 l=0.9
X107 vdd.t217 a_n2650_13878.t66 a_n2472_13878.t0 vdd.t216 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X108 commonsourceibias.t9 commonsourceibias.t8 gnd.t238 gnd.t158 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=2.73 ps=14.78 w=7 l=1
X109 gnd.t237 commonsourceibias.t63 CSoutput.t121 gnd.t146 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X110 vdd.t147 vdd.t144 vdd.t146 vdd.t145 sky130_fd_pr__pfet_01v8 ad=3.51 pd=18.78 as=0 ps=0 w=9 l=0.5
X111 gnd.t106 gnd.t104 gnd.t105 gnd.t27 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=0 ps=0 w=7 l=1
X112 gnd.t236 commonsourceibias.t6 commonsourceibias.t7 gnd.t156 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X113 gnd.t103 gnd.t101 gnd.t102 gnd.t56 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=0 ps=0 w=7 l=1
X114 CSoutput.t98 commonsourceibias.t64 gnd.t235 gnd.t185 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X115 a_n7636_8799.t32 a_n2650_13878.t67 a_n2650_8322.t18 vdd.t184 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X116 a_n2650_8322.t31 a_n2650_13878.t68 vdd.t215 vdd.t214 sky130_fd_pr__pfet_01v8 ad=3.51 pd=18.78 as=1.485 ps=9.33 w=9 l=0.5
X117 vdd.t143 vdd.t140 vdd.t142 vdd.t141 sky130_fd_pr__pfet_01v8 ad=3.51 pd=18.78 as=0 ps=0 w=9 l=0.5
X118 a_n7636_8799.t12 plus.t11 a_n3827_n3924.t18 gnd.t319 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=2.73 ps=14.78 w=7 l=0.9
X119 gnd.t234 commonsourceibias.t65 CSoutput.t141 gnd.t166 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X120 commonsourceibias.t41 commonsourceibias.t40 gnd.t233 gnd.t144 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X121 vdd.t48 a_n7636_8799.t57 CSoutput.t64 vdd.t47 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X122 vdd.t22 a_n7636_8799.t58 CSoutput.t63 vdd.t21 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X123 a_n2650_13878.t50 a_n2650_13878.t49 a_n2472_13878.t15 vdd.t197 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X124 CSoutput.t62 a_n7636_8799.t59 vdd.t24 vdd.t23 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X125 a_n7636_8799.t9 plus.t12 a_n3827_n3924.t17 gnd.t305 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=2.73 ps=14.78 w=7 l=0.9
X126 diffpairibias.t13 diffpairibias.t12 gnd.t19 gnd.t18 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=2.73 ps=14.78 w=7 l=1
X127 CSoutput.t61 a_n7636_8799.t60 vdd.t53 vdd.t16 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X128 a_n7636_8799.t19 a_n2650_13878.t69 a_n2650_8322.t17 vdd.t213 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X129 a_n2472_13878.t14 a_n2650_13878.t31 a_n2650_13878.t32 vdd.t212 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X130 gnd.t100 gnd.t98 gnd.t99 gnd.t23 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=0 ps=0 w=7 l=0.9
X131 gnd.t232 commonsourceibias.t66 CSoutput.t135 gnd.t172 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X132 gnd.t231 commonsourceibias.t67 CSoutput.t109 gnd.t160 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X133 vdd.t37 CSoutput.t148 output.t13 gnd.t285 sky130_fd_pr__nfet_01v8 ad=0.825 pd=5.33 as=0.825 ps=5.33 w=5 l=1
X134 output.t12 CSoutput.t149 vdd.t38 gnd.t284 sky130_fd_pr__nfet_01v8 ad=0.825 pd=5.33 as=0.825 ps=5.33 w=5 l=1
X135 a_n2472_13878.t13 a_n2650_13878.t45 a_n2650_13878.t46 vdd.t211 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X136 CSoutput.t60 a_n7636_8799.t61 vdd.t54 vdd.t49 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X137 vdd.t210 a_n2650_13878.t70 a_n2650_8322.t30 vdd.t209 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=3.51 ps=18.78 w=9 l=0.5
X138 a_n2650_13878.t30 a_n2650_13878.t29 a_n2472_13878.t12 vdd.t181 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X139 vdd.t55 a_n7636_8799.t62 CSoutput.t59 vdd.t6 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X140 vdd.t139 vdd.t137 vdd.t138 vdd.t117 sky130_fd_pr__pfet_01v8 ad=3.12 pd=16.78 as=0 ps=0 w=8 l=0.5
X141 a_n3827_n3924.t16 plus.t13 a_n7636_8799.t6 gnd.t309 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.9
X142 a_n2650_13878.t12 minus.t9 a_n3827_n3924.t36 gnd.t310 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.9
X143 gnd.t97 gnd.t95 gnd.t96 gnd.t60 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=0 ps=0 w=7 l=1
X144 plus.t3 gnd.t92 gnd.t94 gnd.t93 sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.5
X145 CSoutput.t108 commonsourceibias.t68 gnd.t230 gnd.t152 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X146 vdd.t39 CSoutput.t150 output.t11 gnd.t283 sky130_fd_pr__nfet_01v8 ad=0.825 pd=5.33 as=0.825 ps=5.33 w=5 l=1
X147 vdd.t56 a_n7636_8799.t63 CSoutput.t58 vdd.t51 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X148 gnd.t229 commonsourceibias.t69 CSoutput.t110 gnd.t174 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X149 gnd.t228 commonsourceibias.t70 CSoutput.t113 gnd.t176 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=1.155 ps=7.33 w=7 l=1
X150 gnd.t91 gnd.t89 minus.t2 gnd.t90 sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.5
X151 a_n3827_n3924.t7 diffpairibias.t24 gnd.t21 gnd.t20 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=2.73 ps=14.78 w=7 l=1
X152 a_n7636_8799.t5 plus.t14 a_n3827_n3924.t15 gnd.t296 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.9
X153 a_n3827_n3924.t8 diffpairibias.t25 gnd.t271 gnd.t270 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=2.73 ps=14.78 w=7 l=1
X154 vdd.t232 a_n7636_8799.t64 CSoutput.t57 vdd.t2 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X155 gnd.t88 gnd.t86 gnd.t87 gnd.t27 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=0 ps=0 w=7 l=1
X156 a_n2472_13878.t11 a_n2650_13878.t15 a_n2650_13878.t16 vdd.t185 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X157 a_n7636_8799.t4 plus.t15 a_n3827_n3924.t14 gnd.t313 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.9
X158 vdd.t136 vdd.t134 vdd.t135 vdd.t99 sky130_fd_pr__pfet_01v8 ad=3.51 pd=18.78 as=0 ps=0 w=9 l=0.5
X159 a_n2650_8322.t16 a_n2650_13878.t71 a_n7636_8799.t25 vdd.t208 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X160 CSoutput.t56 a_n7636_8799.t65 vdd.t233 vdd.t25 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X161 CSoutput.t55 a_n7636_8799.t66 vdd.t236 vdd.t4 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=3.12 ps=16.78 w=8 l=0.5
X162 CSoutput.t142 commonsourceibias.t71 gnd.t227 gnd.t211 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X163 vdd.t40 CSoutput.t151 output.t10 gnd.t282 sky130_fd_pr__nfet_01v8 ad=0.825 pd=5.33 as=0.825 ps=5.33 w=5 l=1
X164 a_n2472_13878.t25 a_n2650_13878.t72 vdd.t207 vdd.t206 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X165 gnd.t85 gnd.t83 gnd.t84 gnd.t31 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=0 ps=0 w=7 l=1
X166 gnd.t226 commonsourceibias.t72 CSoutput.t101 gnd.t146 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X167 output.t9 CSoutput.t152 vdd.t41 gnd.t281 sky130_fd_pr__nfet_01v8 ad=0.825 pd=5.33 as=0.825 ps=5.33 w=5 l=1
X168 diffpairibias.t11 diffpairibias.t10 gnd.t267 gnd.t266 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=2.73 ps=14.78 w=7 l=1
X169 vdd.t133 vdd.t131 vdd.t132 vdd.t121 sky130_fd_pr__pfet_01v8 ad=3.12 pd=16.78 as=0 ps=0 w=8 l=0.5
X170 vdd.t205 a_n2650_13878.t73 a_n2472_13878.t24 vdd.t204 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X171 a_n2650_13878.t0 minus.t10 a_n3827_n3924.t0 gnd.t0 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.9
X172 vdd.t237 a_n7636_8799.t67 CSoutput.t54 vdd.t6 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X173 CSoutput.t53 a_n7636_8799.t68 vdd.t50 vdd.t49 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X174 a_n3827_n3924.t13 plus.t16 a_n7636_8799.t3 gnd.t1 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.9
X175 gnd.t225 commonsourceibias.t73 CSoutput.t138 gnd.t196 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X176 CSoutput.t128 commonsourceibias.t74 gnd.t224 gnd.t158 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=2.73 ps=14.78 w=7 l=1
X177 vdd.t130 vdd.t128 vdd.t129 vdd.t121 sky130_fd_pr__pfet_01v8 ad=3.12 pd=16.78 as=0 ps=0 w=8 l=0.5
X178 output.t8 CSoutput.t153 vdd.t42 gnd.t280 sky130_fd_pr__nfet_01v8 ad=0.825 pd=5.33 as=0.825 ps=5.33 w=5 l=1
X179 a_n2472_13878.t10 a_n2650_13878.t13 a_n2650_13878.t14 vdd.t203 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X180 gnd.t223 commonsourceibias.t75 CSoutput.t118 gnd.t172 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X181 diffpairibias.t9 diffpairibias.t8 gnd.t325 gnd.t324 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=2.73 ps=14.78 w=7 l=1
X182 CSoutput.t154 a_n2650_8322.t3 sky130_fd_pr__cap_mim_m3_1 l=12 w=12
X183 vdd.t52 a_n7636_8799.t69 CSoutput.t52 vdd.t51 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X184 a_n2650_8322.t15 a_n2650_13878.t74 a_n7636_8799.t27 vdd.t174 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X185 gnd.t82 gnd.t80 gnd.t81 gnd.t27 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=0 ps=0 w=7 l=1
X186 a_n3827_n3924.t31 minus.t11 a_n2650_13878.t7 gnd.t303 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.9
X187 commonsourceibias.t25 commonsourceibias.t24 gnd.t222 gnd.t211 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X188 a_n2472_13878.t9 a_n2650_13878.t37 a_n2650_13878.t38 vdd.t202 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=3.51 ps=18.78 w=9 l=0.5
X189 vdd.t19 a_n7636_8799.t70 CSoutput.t51 vdd.t18 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X190 CSoutput.t50 a_n7636_8799.t71 vdd.t20 vdd.t12 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X191 diffpairibias.t7 diffpairibias.t6 gnd.t321 gnd.t320 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=2.73 ps=14.78 w=7 l=1
X192 vdd.t77 a_n7636_8799.t72 CSoutput.t49 vdd.t2 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X193 vdd.t201 a_n2650_13878.t75 a_n2650_8322.t29 vdd.t200 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=3.51 ps=18.78 w=9 l=0.5
X194 gnd.t79 gnd.t77 minus.t1 gnd.t78 sky130_fd_pr__nfet_01v8 ad=0.39 pd=2.78 as=0.165 ps=1.33 w=1 l=0.5
X195 plus.t2 gnd.t74 gnd.t76 gnd.t75 sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.5
X196 CSoutput.t155 a_n2650_8322.t2 sky130_fd_pr__cap_mim_m3_1 l=12 w=12
X197 output.t17 outputibias.t10 gnd.t293 gnd.t292 sky130_fd_pr__nfet_01v8 ad=2.34 pd=12.78 as=2.34 ps=12.78 w=6 l=2
X198 CSoutput.t136 commonsourceibias.t76 gnd.t221 gnd.t154 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X199 gnd.t73 gnd.t70 gnd.t72 gnd.t71 sky130_fd_pr__nfet_01v8 ad=1.95 pd=10.78 as=0 ps=0 w=5 l=1
X200 gnd.t69 gnd.t67 gnd.t68 gnd.t56 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=0 ps=0 w=7 l=1
X201 commonsourceibias.t23 commonsourceibias.t22 gnd.t220 gnd.t190 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X202 a_n2472_13878.t1 a_n2650_13878.t76 vdd.t199 vdd.t198 sky130_fd_pr__pfet_01v8 ad=3.51 pd=18.78 as=1.485 ps=9.33 w=9 l=0.5
X203 gnd.t66 gnd.t63 gnd.t65 gnd.t64 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=0 ps=0 w=7 l=1
X204 vdd.t78 a_n7636_8799.t73 CSoutput.t48 vdd.t14 sky130_fd_pr__pfet_01v8 ad=3.12 pd=16.78 as=1.32 ps=8.33 w=8 l=0.5
X205 CSoutput.t116 commonsourceibias.t77 gnd.t219 gnd.t154 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X206 vdd.t70 CSoutput.t156 output.t7 gnd.t279 sky130_fd_pr__nfet_01v8 ad=0.825 pd=5.33 as=0.825 ps=5.33 w=5 l=1
X207 output.t16 outputibias.t11 gnd.t143 gnd.t142 sky130_fd_pr__nfet_01v8 ad=2.34 pd=12.78 as=2.34 ps=12.78 w=6 l=2
X208 gnd.t218 commonsourceibias.t78 CSoutput.t112 gnd.t201 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X209 CSoutput.t111 commonsourceibias.t79 gnd.t217 gnd.t162 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X210 gnd.t216 commonsourceibias.t28 commonsourceibias.t29 gnd.t164 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=1.155 ps=7.33 w=7 l=1
X211 gnd.t215 commonsourceibias.t80 CSoutput.t4 gnd.t176 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=1.155 ps=7.33 w=7 l=1
X212 vdd.t127 vdd.t124 vdd.t126 vdd.t125 sky130_fd_pr__pfet_01v8 ad=3.12 pd=16.78 as=0 ps=0 w=8 l=0.5
X213 gnd.t62 gnd.t59 gnd.t61 gnd.t60 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=0 ps=0 w=7 l=1
X214 CSoutput.t126 commonsourceibias.t81 gnd.t214 gnd.t199 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X215 gnd.t213 commonsourceibias.t82 CSoutput.t1 gnd.t160 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X216 CSoutput.t2 commonsourceibias.t83 gnd.t212 gnd.t211 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X217 a_n2650_8322.t14 a_n2650_13878.t77 a_n7636_8799.t22 vdd.t197 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X218 vdd.t196 a_n2650_13878.t78 a_n2650_8322.t28 vdd.t195 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X219 vdd.t123 vdd.t120 vdd.t122 vdd.t121 sky130_fd_pr__pfet_01v8 ad=3.12 pd=16.78 as=0 ps=0 w=8 l=0.5
X220 commonsourceibias.t27 commonsourceibias.t26 gnd.t210 gnd.t152 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X221 a_n3827_n3924.t3 diffpairibias.t26 gnd.t8 gnd.t7 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=2.73 ps=14.78 w=7 l=1
X222 CSoutput.t47 a_n7636_8799.t74 vdd.t81 vdd.t64 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X223 vdd.t119 vdd.t116 vdd.t118 vdd.t117 sky130_fd_pr__pfet_01v8 ad=3.12 pd=16.78 as=0 ps=0 w=8 l=0.5
X224 CSoutput.t130 commonsourceibias.t84 gnd.t209 gnd.t170 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X225 gnd.t208 commonsourceibias.t85 CSoutput.t6 gnd.t148 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X226 a_n7636_8799.t2 plus.t17 a_n3827_n3924.t12 gnd.t308 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.9
X227 a_n2650_13878.t53 minus.t12 a_n3827_n3924.t39 gnd.t314 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.9
X228 vdd.t83 a_n7636_8799.t75 CSoutput.t46 vdd.t82 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X229 vdd.t30 a_n7636_8799.t76 CSoutput.t45 vdd.t29 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X230 vdd.t115 vdd.t113 vdd.t114 vdd.t95 sky130_fd_pr__pfet_01v8 ad=3.12 pd=16.78 as=0 ps=0 w=8 l=0.5
X231 a_n3827_n3924.t4 minus.t13 a_n2650_13878.t2 gnd.t4 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=1.155 ps=7.33 w=7 l=0.9
X232 gnd.t207 commonsourceibias.t86 CSoutput.t115 gnd.t188 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X233 CSoutput.t0 commonsourceibias.t87 gnd.t206 gnd.t170 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X234 CSoutput.t96 commonsourceibias.t88 gnd.t205 gnd.t144 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X235 gnd.t204 commonsourceibias.t89 CSoutput.t94 gnd.t164 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=1.155 ps=7.33 w=7 l=1
X236 vdd.t112 vdd.t109 vdd.t111 vdd.t110 sky130_fd_pr__pfet_01v8 ad=3.51 pd=18.78 as=0 ps=0 w=9 l=0.5
X237 vdd.t32 a_n7636_8799.t77 CSoutput.t44 vdd.t31 sky130_fd_pr__pfet_01v8 ad=3.12 pd=16.78 as=1.32 ps=8.33 w=8 l=0.5
X238 a_n3827_n3924.t28 minus.t14 a_n2650_13878.t5 gnd.t299 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.9
X239 gnd.t58 gnd.t55 gnd.t57 gnd.t56 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=0 ps=0 w=7 l=1
X240 CSoutput.t43 a_n7636_8799.t78 vdd.t172 vdd.t12 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X241 CSoutput.t42 a_n7636_8799.t79 vdd.t173 vdd.t0 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=3.12 ps=16.78 w=8 l=0.5
X242 a_n2472_13878.t8 a_n2650_13878.t47 a_n2650_13878.t48 vdd.t189 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X243 a_n3827_n3924.t30 minus.t15 a_n2650_13878.t6 gnd.t302 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=1.155 ps=7.33 w=7 l=0.9
X244 vdd.t108 vdd.t106 vdd.t107 vdd.t95 sky130_fd_pr__pfet_01v8 ad=3.12 pd=16.78 as=0 ps=0 w=8 l=0.5
X245 a_n2650_8322.t13 a_n2650_13878.t79 a_n7636_8799.t23 vdd.t194 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X246 diffpairibias.t5 diffpairibias.t4 gnd.t307 gnd.t306 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=2.73 ps=14.78 w=7 l=1
X247 CSoutput.t122 commonsourceibias.t90 gnd.t203 gnd.t185 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X248 gnd.t202 commonsourceibias.t91 CSoutput.t7 gnd.t201 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X249 output.t6 CSoutput.t157 vdd.t43 gnd.t278 sky130_fd_pr__nfet_01v8 ad=0.825 pd=5.33 as=0.825 ps=5.33 w=5 l=1
X250 CSoutput.t123 commonsourceibias.t92 gnd.t200 gnd.t199 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X251 CSoutput.t41 a_n7636_8799.t80 vdd.t230 vdd.t16 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X252 CSoutput.t40 a_n7636_8799.t81 vdd.t231 vdd.t23 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X253 vdd.t228 a_n7636_8799.t82 CSoutput.t39 vdd.t82 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X254 gnd.t198 commonsourceibias.t93 CSoutput.t129 gnd.t188 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X255 a_n3827_n3924.t25 diffpairibias.t27 gnd.t295 gnd.t294 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=2.73 ps=14.78 w=7 l=1
X256 vdd.t229 a_n7636_8799.t83 CSoutput.t38 vdd.t14 sky130_fd_pr__pfet_01v8 ad=3.12 pd=16.78 as=1.32 ps=8.33 w=8 l=0.5
X257 gnd.t197 commonsourceibias.t94 CSoutput.t11 gnd.t196 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X258 a_n2650_8322.t27 a_n2650_13878.t80 vdd.t193 vdd.t192 sky130_fd_pr__pfet_01v8 ad=3.51 pd=18.78 as=1.485 ps=9.33 w=9 l=0.5
X259 CSoutput.t143 commonsourceibias.t95 gnd.t195 gnd.t150 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=2.73 ps=14.78 w=7 l=1
X260 gnd.t147 commonsourceibias.t2 commonsourceibias.t3 gnd.t146 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X261 outputibias.t3 outputibias.t2 gnd.t327 gnd.t326 sky130_fd_pr__nfet_01v8 ad=2.34 pd=12.78 as=2.34 ps=12.78 w=6 l=2
X262 gnd.t194 commonsourceibias.t96 CSoutput.t5 gnd.t166 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X263 a_n3827_n3924.t32 minus.t16 a_n2650_13878.t8 gnd.t304 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.9
X264 vdd.t191 a_n2650_13878.t81 a_n2472_13878.t3 vdd.t190 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=3.51 ps=18.78 w=9 l=0.5
X265 CSoutput.t37 a_n7636_8799.t84 vdd.t66 vdd.t64 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X266 CSoutput.t36 a_n7636_8799.t85 vdd.t67 vdd.t35 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X267 CSoutput.t105 commonsourceibias.t97 gnd.t193 gnd.t150 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=2.73 ps=14.78 w=7 l=1
X268 gnd.t192 commonsourceibias.t98 CSoutput.t107 gnd.t156 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X269 CSoutput.t127 commonsourceibias.t99 gnd.t191 gnd.t190 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X270 gnd.t189 commonsourceibias.t100 CSoutput.t140 gnd.t188 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X271 vdd.t238 a_n7636_8799.t86 CSoutput.t35 vdd.t82 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X272 vdd.t239 a_n7636_8799.t87 CSoutput.t34 vdd.t29 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X273 gnd.t187 commonsourceibias.t101 CSoutput.t97 gnd.t174 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X274 gnd.t54 gnd.t51 gnd.t53 gnd.t52 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=0 ps=0 w=7 l=0.9
X275 commonsourceibias.t33 commonsourceibias.t32 gnd.t186 gnd.t185 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X276 gnd.t50 gnd.t48 plus.t1 gnd.t49 sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.5
X277 gnd.t184 commonsourceibias.t30 commonsourceibias.t31 gnd.t166 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X278 a_n7636_8799.t30 a_n2650_13878.t82 a_n2650_8322.t12 vdd.t189 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X279 a_n2650_8322.t11 a_n2650_13878.t83 a_n7636_8799.t18 vdd.t182 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X280 a_n2472_13878.t2 a_n2650_13878.t84 vdd.t188 vdd.t187 sky130_fd_pr__pfet_01v8 ad=3.51 pd=18.78 as=1.485 ps=9.33 w=9 l=0.5
X281 vdd.t105 vdd.t102 vdd.t104 vdd.t103 sky130_fd_pr__pfet_01v8 ad=3.51 pd=18.78 as=0 ps=0 w=9 l=0.5
X282 gnd.t183 commonsourceibias.t102 CSoutput.t103 gnd.t146 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X283 CSoutput.t93 commonsourceibias.t103 gnd.t182 gnd.t154 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X284 vdd.t11 a_n7636_8799.t88 CSoutput.t33 vdd.t10 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X285 CSoutput.t32 a_n7636_8799.t89 vdd.t13 vdd.t12 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X286 vdd.t101 vdd.t98 vdd.t100 vdd.t99 sky130_fd_pr__pfet_01v8 ad=3.51 pd=18.78 as=0 ps=0 w=9 l=0.5
X287 vdd.t44 CSoutput.t158 output.t5 gnd.t277 sky130_fd_pr__nfet_01v8 ad=0.825 pd=5.33 as=0.825 ps=5.33 w=5 l=1
X288 vdd.t97 vdd.t94 vdd.t96 vdd.t95 sky130_fd_pr__pfet_01v8 ad=3.12 pd=16.78 as=0 ps=0 w=8 l=0.5
X289 a_n3827_n3924.t11 plus.t18 a_n7636_8799.t10 gnd.t13 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.9
X290 gnd.t180 commonsourceibias.t46 commonsourceibias.t47 gnd.t172 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X291 a_n2650_8322.t10 a_n2650_13878.t85 a_n7636_8799.t21 vdd.t186 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X292 a_n7636_8799.t33 a_n2650_13878.t86 a_n2650_8322.t9 vdd.t185 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X293 CSoutput.t89 commonsourceibias.t104 gnd.t181 gnd.t144 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X294 a_n2650_13878.t9 minus.t17 a_n3827_n3924.t33 gnd.t305 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=2.73 ps=14.78 w=7 l=0.9
X295 CSoutput.t31 a_n7636_8799.t90 vdd.t79 vdd.t23 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X296 vdd.t80 a_n7636_8799.t91 CSoutput.t30 vdd.t51 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X297 CSoutput.t29 a_n7636_8799.t92 vdd.t88 vdd.t57 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X298 CSoutput.t28 a_n7636_8799.t93 vdd.t89 vdd.t57 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X299 a_n2472_13878.t7 a_n2650_13878.t33 a_n2650_13878.t34 vdd.t184 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X300 gnd.t179 commonsourceibias.t105 CSoutput.t124 gnd.t148 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X301 CSoutput.t88 commonsourceibias.t106 gnd.t178 gnd.t168 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X302 vdd.t86 a_n7636_8799.t94 CSoutput.t27 vdd.t62 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X303 gnd.t177 commonsourceibias.t44 commonsourceibias.t45 gnd.t176 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=1.155 ps=7.33 w=7 l=1
X304 gnd.t175 commonsourceibias.t42 commonsourceibias.t43 gnd.t174 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X305 vdd.t87 a_n7636_8799.t95 CSoutput.t26 vdd.t31 sky130_fd_pr__pfet_01v8 ad=3.12 pd=16.78 as=1.32 ps=8.33 w=8 l=0.5
X306 gnd.t173 commonsourceibias.t107 CSoutput.t95 gnd.t172 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X307 CSoutput.t3 commonsourceibias.t108 gnd.t171 gnd.t170 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X308 a_n3827_n3924.t35 minus.t18 a_n2650_13878.t11 gnd.t309 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.9
X309 a_n3827_n3924.t27 diffpairibias.t28 gnd.t298 gnd.t297 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=2.73 ps=14.78 w=7 l=1
X310 CSoutput.t25 a_n7636_8799.t96 vdd.t26 vdd.t25 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X311 a_n7636_8799.t28 a_n2650_13878.t87 a_n2650_8322.t8 vdd.t183 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X312 a_n2650_13878.t44 a_n2650_13878.t43 a_n2472_13878.t6 vdd.t182 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X313 output.t4 CSoutput.t159 vdd.t45 gnd.t276 sky130_fd_pr__nfet_01v8 ad=0.825 pd=5.33 as=0.825 ps=5.33 w=5 l=1
X314 CSoutput.t24 a_n7636_8799.t97 vdd.t28 vdd.t27 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X315 vdd.t63 a_n7636_8799.t98 CSoutput.t23 vdd.t62 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X316 gnd.t47 gnd.t44 gnd.t46 gnd.t45 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=0 ps=0 w=7 l=1
X317 CSoutput.t22 a_n7636_8799.t99 vdd.t65 vdd.t64 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X318 vdd.t170 a_n7636_8799.t100 CSoutput.t21 vdd.t47 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X319 minus.t0 gnd.t41 gnd.t43 gnd.t42 sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.5
X320 gnd.t40 gnd.t38 plus.t0 gnd.t39 sky130_fd_pr__nfet_01v8 ad=0.39 pd=2.78 as=0.165 ps=1.33 w=1 l=0.5
X321 CSoutput.t114 commonsourceibias.t109 gnd.t169 gnd.t168 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X322 gnd.t167 commonsourceibias.t110 CSoutput.t134 gnd.t166 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X323 diffpairibias.t3 diffpairibias.t2 gnd.t17 gnd.t16 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=2.73 ps=14.78 w=7 l=1
X324 gnd.t37 gnd.t34 gnd.t36 gnd.t35 sky130_fd_pr__nfet_01v8 ad=2.34 pd=12.78 as=0 ps=0 w=6 l=2
X325 a_n2650_8322.t7 a_n2650_13878.t88 a_n7636_8799.t17 vdd.t181 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X326 a_n2650_13878.t4 minus.t19 a_n3827_n3924.t26 gnd.t296 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.9
X327 vdd.t68 CSoutput.t160 output.t3 gnd.t275 sky130_fd_pr__nfet_01v8 ad=0.825 pd=5.33 as=0.825 ps=5.33 w=5 l=1
X328 output.t2 CSoutput.t161 vdd.t69 gnd.t274 sky130_fd_pr__nfet_01v8 ad=1.95 pd=10.78 as=0.825 ps=5.33 w=5 l=1
X329 vdd.t171 a_n7636_8799.t101 CSoutput.t20 vdd.t10 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X330 gnd.t165 commonsourceibias.t111 CSoutput.t92 gnd.t164 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=1.155 ps=7.33 w=7 l=1
X331 CSoutput.t162 a_n2650_8322.t1 sky130_fd_pr__cap_mim_m3_1 l=12 w=12
X332 gnd.t33 gnd.t30 gnd.t32 gnd.t31 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=0 ps=0 w=7 l=1
X333 CSoutput.t100 commonsourceibias.t112 gnd.t163 gnd.t162 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X334 diffpairibias.t1 diffpairibias.t0 gnd.t265 gnd.t264 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=2.73 ps=14.78 w=7 l=1
X335 outputibias.t1 outputibias.t0 gnd.t12 gnd.t11 sky130_fd_pr__nfet_01v8 ad=2.34 pd=12.78 as=2.34 ps=12.78 w=6 l=2
X336 CSoutput.t19 a_n7636_8799.t102 vdd.t58 vdd.t57 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X337 vdd.t180 a_n2650_13878.t89 a_n2472_13878.t27 vdd.t179 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=3.51 ps=18.78 w=9 l=0.5
X338 CSoutput.t163 a_n2650_8322.t0 sky130_fd_pr__cap_mim_m3_1 l=12 w=12
X339 vdd.t59 a_n7636_8799.t103 CSoutput.t18 vdd.t29 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X340 vdd.t226 a_n7636_8799.t104 CSoutput.t17 vdd.t62 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X341 CSoutput.t16 a_n7636_8799.t105 vdd.t227 vdd.t33 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X342 gnd.t161 commonsourceibias.t113 CSoutput.t13 gnd.t160 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X343 a_n7636_8799.t13 plus.t19 a_n3827_n3924.t10 gnd.t0 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.9
X344 gnd.t29 gnd.t26 gnd.t28 gnd.t27 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=0 ps=0 w=7 l=1
X345 a_n2650_8322.t6 a_n2650_13878.t90 a_n7636_8799.t31 vdd.t178 sky130_fd_pr__pfet_01v8 ad=3.51 pd=18.78 as=1.485 ps=9.33 w=9 l=0.5
X346 a_n2650_13878.t55 minus.t20 a_n3827_n3924.t41 gnd.t319 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=2.73 ps=14.78 w=7 l=0.9
X347 vdd.t92 CSoutput.t164 output.t1 gnd.t273 sky130_fd_pr__nfet_01v8 ad=0.825 pd=5.33 as=1.95 ps=10.78 w=5 l=1
X348 CSoutput.t15 a_n7636_8799.t106 vdd.t90 vdd.t25 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X349 vdd.t91 a_n7636_8799.t107 CSoutput.t14 vdd.t31 sky130_fd_pr__pfet_01v8 ad=3.12 pd=16.78 as=1.32 ps=8.33 w=8 l=0.5
X350 CSoutput.t9 commonsourceibias.t114 gnd.t159 gnd.t158 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=2.73 ps=14.78 w=7 l=1
X351 gnd.t157 commonsourceibias.t115 CSoutput.t10 gnd.t156 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X352 commonsourceibias.t1 commonsourceibias.t0 gnd.t155 gnd.t154 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X353 a_n2650_8322.t26 a_n2650_13878.t91 vdd.t177 vdd.t176 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X354 a_n2472_13878.t5 a_n2650_13878.t19 a_n2650_13878.t20 vdd.t175 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=3.51 ps=18.78 w=9 l=0.5
X355 gnd.t25 gnd.t22 gnd.t24 gnd.t23 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=0 ps=0 w=7 l=0.9
X356 CSoutput.t12 commonsourceibias.t116 gnd.t153 gnd.t152 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X357 a_n3827_n3924.t9 plus.t20 a_n7636_8799.t11 gnd.t303 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.9
X358 vdd.t93 CSoutput.t165 output.t0 gnd.t272 sky130_fd_pr__nfet_01v8 ad=0.825 pd=5.33 as=0.825 ps=5.33 w=5 l=1
X359 a_n2650_13878.t42 a_n2650_13878.t41 a_n2472_13878.t4 vdd.t174 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X360 CSoutput.t132 commonsourceibias.t117 gnd.t151 gnd.t150 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=2.73 ps=14.78 w=7 l=1
X361 gnd.t149 commonsourceibias.t118 CSoutput.t8 gnd.t148 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X362 CSoutput.t119 commonsourceibias.t119 gnd.t145 gnd.t144 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X363 a_n3827_n3924.t2 diffpairibias.t29 gnd.t3 gnd.t2 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=2.73 ps=14.78 w=7 l=1
R0 a_n2650_13878.n131 a_n2650_13878.t27 512.366
R1 a_n2650_13878.n130 a_n2650_13878.t15 512.366
R2 a_n2650_13878.n70 a_n2650_13878.t51 512.366
R3 a_n2650_13878.n129 a_n2650_13878.t13 512.366
R4 a_n2650_13878.n128 a_n2650_13878.t43 512.366
R5 a_n2650_13878.n71 a_n2650_13878.t47 512.366
R6 a_n2650_13878.n127 a_n2650_13878.t35 512.366
R7 a_n2650_13878.n126 a_n2650_13878.t33 512.366
R8 a_n2650_13878.n72 a_n2650_13878.t49 512.366
R9 a_n2650_13878.n117 a_n2650_13878.t90 512.366
R10 a_n2650_13878.n116 a_n2650_13878.t69 512.366
R11 a_n2650_13878.n73 a_n2650_13878.t74 512.366
R12 a_n2650_13878.n115 a_n2650_13878.t63 512.366
R13 a_n2650_13878.n114 a_n2650_13878.t79 512.366
R14 a_n2650_13878.n74 a_n2650_13878.t87 512.366
R15 a_n2650_13878.n113 a_n2650_13878.t88 512.366
R16 a_n2650_13878.n112 a_n2650_13878.t58 512.366
R17 a_n2650_13878.n75 a_n2650_13878.t71 512.366
R18 a_n2650_13878.n91 a_n2650_13878.t25 512.366
R19 a_n2650_13878.n92 a_n2650_13878.t39 512.366
R20 a_n2650_13878.n81 a_n2650_13878.t41 512.366
R21 a_n2650_13878.n93 a_n2650_13878.t31 512.366
R22 a_n2650_13878.n94 a_n2650_13878.t17 512.366
R23 a_n2650_13878.n95 a_n2650_13878.t23 512.366
R24 a_n2650_13878.n96 a_n2650_13878.t29 512.366
R25 a_n2650_13878.n80 a_n2650_13878.t45 512.366
R26 a_n2650_13878.n97 a_n2650_13878.t21 512.366
R27 a_n2650_13878.n84 a_n2650_13878.t62 512.366
R28 a_n2650_13878.n85 a_n2650_13878.t86 512.366
R29 a_n2650_13878.n83 a_n2650_13878.t85 512.366
R30 a_n2650_13878.n86 a_n2650_13878.t60 512.366
R31 a_n2650_13878.n87 a_n2650_13878.t83 512.366
R32 a_n2650_13878.n88 a_n2650_13878.t82 512.366
R33 a_n2650_13878.n89 a_n2650_13878.t57 512.366
R34 a_n2650_13878.n82 a_n2650_13878.t67 512.366
R35 a_n2650_13878.n90 a_n2650_13878.t77 512.366
R36 a_n2650_13878.n109 a_n2650_13878.t76 512.366
R37 a_n2650_13878.n99 a_n2650_13878.t66 512.366
R38 a_n2650_13878.n110 a_n2650_13878.t56 512.366
R39 a_n2650_13878.n107 a_n2650_13878.t84 512.366
R40 a_n2650_13878.n100 a_n2650_13878.t73 512.366
R41 a_n2650_13878.n108 a_n2650_13878.t72 512.366
R42 a_n2650_13878.n105 a_n2650_13878.t80 512.366
R43 a_n2650_13878.n101 a_n2650_13878.t65 512.366
R44 a_n2650_13878.n106 a_n2650_13878.t64 512.366
R45 a_n2650_13878.n103 a_n2650_13878.t68 512.366
R46 a_n2650_13878.n102 a_n2650_13878.t78 512.366
R47 a_n2650_13878.n104 a_n2650_13878.t91 512.366
R48 a_n2650_13878.n33 a_n2650_13878.n69 70.1674
R49 a_n2650_13878.n7 a_n2650_13878.n62 70.1674
R50 a_n2650_13878.n20 a_n2650_13878.n47 70.1674
R51 a_n2650_13878.n24 a_n2650_13878.n40 70.1674
R52 a_n2650_13878.n90 a_n2650_13878.n40 20.9683
R53 a_n2650_13878.n39 a_n2650_13878.n24 74.73
R54 a_n2650_13878.n39 a_n2650_13878.n82 11.843
R55 a_n2650_13878.n23 a_n2650_13878.n38 80.4688
R56 a_n2650_13878.n89 a_n2650_13878.n38 0.365327
R57 a_n2650_13878.n37 a_n2650_13878.n23 75.0448
R58 a_n2650_13878.n25 a_n2650_13878.n36 70.1674
R59 a_n2650_13878.n86 a_n2650_13878.n36 20.9683
R60 a_n2650_13878.n35 a_n2650_13878.n25 70.3058
R61 a_n2650_13878.n35 a_n2650_13878.n83 20.6913
R62 a_n2650_13878.n26 a_n2650_13878.n34 75.3623
R63 a_n2650_13878.n85 a_n2650_13878.n34 10.5784
R64 a_n2650_13878.n84 a_n2650_13878.n26 161.3
R65 a_n2650_13878.n97 a_n2650_13878.n47 20.9683
R66 a_n2650_13878.n46 a_n2650_13878.n20 74.73
R67 a_n2650_13878.n46 a_n2650_13878.n80 11.843
R68 a_n2650_13878.n19 a_n2650_13878.n45 80.4688
R69 a_n2650_13878.n96 a_n2650_13878.n45 0.365327
R70 a_n2650_13878.n44 a_n2650_13878.n19 75.0448
R71 a_n2650_13878.n21 a_n2650_13878.n43 70.1674
R72 a_n2650_13878.n93 a_n2650_13878.n43 20.9683
R73 a_n2650_13878.n42 a_n2650_13878.n21 70.3058
R74 a_n2650_13878.n42 a_n2650_13878.n81 20.6913
R75 a_n2650_13878.n22 a_n2650_13878.n41 75.3623
R76 a_n2650_13878.n92 a_n2650_13878.n41 10.5784
R77 a_n2650_13878.n91 a_n2650_13878.n22 161.3
R78 a_n2650_13878.n10 a_n2650_13878.n55 70.1674
R79 a_n2650_13878.n12 a_n2650_13878.n53 70.1674
R80 a_n2650_13878.n14 a_n2650_13878.n51 70.1674
R81 a_n2650_13878.n17 a_n2650_13878.n49 70.1674
R82 a_n2650_13878.n104 a_n2650_13878.n49 20.9683
R83 a_n2650_13878.n48 a_n2650_13878.n18 75.0448
R84 a_n2650_13878.n48 a_n2650_13878.n102 11.2134
R85 a_n2650_13878.n18 a_n2650_13878.n103 161.3
R86 a_n2650_13878.n106 a_n2650_13878.n51 20.9683
R87 a_n2650_13878.n50 a_n2650_13878.n15 75.0448
R88 a_n2650_13878.n50 a_n2650_13878.n101 11.2134
R89 a_n2650_13878.n15 a_n2650_13878.n105 161.3
R90 a_n2650_13878.n108 a_n2650_13878.n53 20.9683
R91 a_n2650_13878.n52 a_n2650_13878.n13 75.0448
R92 a_n2650_13878.n52 a_n2650_13878.n100 11.2134
R93 a_n2650_13878.n13 a_n2650_13878.n107 161.3
R94 a_n2650_13878.n110 a_n2650_13878.n55 20.9683
R95 a_n2650_13878.n54 a_n2650_13878.n11 75.0448
R96 a_n2650_13878.n54 a_n2650_13878.n99 11.2134
R97 a_n2650_13878.n11 a_n2650_13878.n109 161.3
R98 a_n2650_13878.n62 a_n2650_13878.n75 20.9683
R99 a_n2650_13878.n61 a_n2650_13878.n7 74.73
R100 a_n2650_13878.n112 a_n2650_13878.n61 11.843
R101 a_n2650_13878.n60 a_n2650_13878.n6 80.4688
R102 a_n2650_13878.n60 a_n2650_13878.n113 0.365327
R103 a_n2650_13878.n6 a_n2650_13878.n59 75.0448
R104 a_n2650_13878.n58 a_n2650_13878.n8 70.1674
R105 a_n2650_13878.n115 a_n2650_13878.n58 20.9683
R106 a_n2650_13878.n8 a_n2650_13878.n57 70.3058
R107 a_n2650_13878.n57 a_n2650_13878.n73 20.6913
R108 a_n2650_13878.n56 a_n2650_13878.n9 75.3623
R109 a_n2650_13878.n116 a_n2650_13878.n56 10.5784
R110 a_n2650_13878.n9 a_n2650_13878.n117 161.3
R111 a_n2650_13878.n69 a_n2650_13878.n72 20.9683
R112 a_n2650_13878.n68 a_n2650_13878.n33 74.73
R113 a_n2650_13878.n126 a_n2650_13878.n68 11.843
R114 a_n2650_13878.n67 a_n2650_13878.n4 80.4688
R115 a_n2650_13878.n67 a_n2650_13878.n127 0.365327
R116 a_n2650_13878.n4 a_n2650_13878.n66 75.0448
R117 a_n2650_13878.n65 a_n2650_13878.n3 70.1674
R118 a_n2650_13878.n129 a_n2650_13878.n65 20.9683
R119 a_n2650_13878.n3 a_n2650_13878.n64 70.3058
R120 a_n2650_13878.n64 a_n2650_13878.n70 20.6913
R121 a_n2650_13878.n63 a_n2650_13878.n5 75.3623
R122 a_n2650_13878.n130 a_n2650_13878.n63 10.5784
R123 a_n2650_13878.n5 a_n2650_13878.n131 161.3
R124 a_n2650_13878.n1 a_n2650_13878.n124 81.4626
R125 a_n2650_13878.n2 a_n2650_13878.n120 81.4626
R126 a_n2650_13878.n2 a_n2650_13878.n118 81.4626
R127 a_n2650_13878.n1 a_n2650_13878.n125 80.9324
R128 a_n2650_13878.n1 a_n2650_13878.n123 80.9324
R129 a_n2650_13878.n0 a_n2650_13878.n122 80.9324
R130 a_n2650_13878.n2 a_n2650_13878.n121 80.9324
R131 a_n2650_13878.n2 a_n2650_13878.n119 80.9324
R132 a_n2650_13878.n30 a_n2650_13878.t20 74.6477
R133 a_n2650_13878.n27 a_n2650_13878.t26 74.6477
R134 a_n2650_13878.n31 a_n2650_13878.t28 74.2899
R135 a_n2650_13878.n29 a_n2650_13878.t38 74.2897
R136 a_n2650_13878.n30 a_n2650_13878.n134 70.6783
R137 a_n2650_13878.n30 a_n2650_13878.n135 70.6783
R138 a_n2650_13878.n32 a_n2650_13878.n133 70.6783
R139 a_n2650_13878.n29 a_n2650_13878.n79 70.6783
R140 a_n2650_13878.n28 a_n2650_13878.n78 70.6783
R141 a_n2650_13878.n28 a_n2650_13878.n77 70.6783
R142 a_n2650_13878.n27 a_n2650_13878.n76 70.6783
R143 a_n2650_13878.n136 a_n2650_13878.n32 70.6782
R144 a_n2650_13878.n131 a_n2650_13878.n130 48.2005
R145 a_n2650_13878.n65 a_n2650_13878.n128 20.9683
R146 a_n2650_13878.n127 a_n2650_13878.n71 48.2005
R147 a_n2650_13878.t19 a_n2650_13878.n69 533.335
R148 a_n2650_13878.n117 a_n2650_13878.n116 48.2005
R149 a_n2650_13878.n58 a_n2650_13878.n114 20.9683
R150 a_n2650_13878.n113 a_n2650_13878.n74 48.2005
R151 a_n2650_13878.t61 a_n2650_13878.n62 533.335
R152 a_n2650_13878.n92 a_n2650_13878.n91 48.2005
R153 a_n2650_13878.n94 a_n2650_13878.n43 20.9683
R154 a_n2650_13878.n96 a_n2650_13878.n95 48.2005
R155 a_n2650_13878.t37 a_n2650_13878.n47 533.335
R156 a_n2650_13878.n85 a_n2650_13878.n84 48.2005
R157 a_n2650_13878.n87 a_n2650_13878.n36 20.9683
R158 a_n2650_13878.n89 a_n2650_13878.n88 48.2005
R159 a_n2650_13878.t59 a_n2650_13878.n40 533.335
R160 a_n2650_13878.n109 a_n2650_13878.n99 48.2005
R161 a_n2650_13878.t81 a_n2650_13878.n55 533.335
R162 a_n2650_13878.n107 a_n2650_13878.n100 48.2005
R163 a_n2650_13878.t89 a_n2650_13878.n53 533.335
R164 a_n2650_13878.n105 a_n2650_13878.n101 48.2005
R165 a_n2650_13878.t75 a_n2650_13878.n51 533.335
R166 a_n2650_13878.n103 a_n2650_13878.n102 48.2005
R167 a_n2650_13878.t70 a_n2650_13878.n49 533.335
R168 a_n2650_13878.n129 a_n2650_13878.n64 21.4216
R169 a_n2650_13878.n115 a_n2650_13878.n57 21.4216
R170 a_n2650_13878.n93 a_n2650_13878.n42 21.4216
R171 a_n2650_13878.n86 a_n2650_13878.n35 21.4216
R172 a_n2650_13878.n68 a_n2650_13878.n72 34.4824
R173 a_n2650_13878.n61 a_n2650_13878.n75 34.4824
R174 a_n2650_13878.n97 a_n2650_13878.n46 34.4824
R175 a_n2650_13878.n90 a_n2650_13878.n39 34.4824
R176 a_n2650_13878.n128 a_n2650_13878.n66 35.3134
R177 a_n2650_13878.n66 a_n2650_13878.n71 11.2134
R178 a_n2650_13878.n114 a_n2650_13878.n59 35.3134
R179 a_n2650_13878.n59 a_n2650_13878.n74 11.2134
R180 a_n2650_13878.n94 a_n2650_13878.n44 35.3134
R181 a_n2650_13878.n95 a_n2650_13878.n44 11.2134
R182 a_n2650_13878.n87 a_n2650_13878.n37 35.3134
R183 a_n2650_13878.n88 a_n2650_13878.n37 11.2134
R184 a_n2650_13878.n110 a_n2650_13878.n54 35.3134
R185 a_n2650_13878.n108 a_n2650_13878.n52 35.3134
R186 a_n2650_13878.n106 a_n2650_13878.n50 35.3134
R187 a_n2650_13878.n104 a_n2650_13878.n48 35.3134
R188 a_n2650_13878.n33 a_n2650_13878.n1 23.891
R189 a_n2650_13878.n63 a_n2650_13878.n70 36.139
R190 a_n2650_13878.n56 a_n2650_13878.n73 36.139
R191 a_n2650_13878.n81 a_n2650_13878.n41 36.139
R192 a_n2650_13878.n83 a_n2650_13878.n34 36.139
R193 a_n2650_13878.n26 a_n2650_13878.n16 13.3641
R194 a_n2650_13878.n7 a_n2650_13878.n111 13.1596
R195 a_n2650_13878.n132 a_n2650_13878.n5 11.8547
R196 a_n2650_13878.n98 a_n2650_13878.n29 10.2167
R197 a_n2650_13878.n18 a_n2650_13878.n16 9.99103
R198 a_n2650_13878.n111 a_n2650_13878.n10 9.99103
R199 a_n2650_13878.n98 a_n2650_13878.n20 8.01944
R200 a_n2650_13878.n31 a_n2650_13878.n132 6.37334
R201 a_n2650_13878.n111 a_n2650_13878.n98 5.3452
R202 a_n2650_13878.n22 a_n2650_13878.n24 4.07247
R203 a_n2650_13878.n33 a_n2650_13878.n9 4.06146
R204 a_n2650_13878.n134 a_n2650_13878.t34 3.61217
R205 a_n2650_13878.n134 a_n2650_13878.t50 3.61217
R206 a_n2650_13878.n135 a_n2650_13878.t48 3.61217
R207 a_n2650_13878.n135 a_n2650_13878.t36 3.61217
R208 a_n2650_13878.n133 a_n2650_13878.t16 3.61217
R209 a_n2650_13878.n133 a_n2650_13878.t52 3.61217
R210 a_n2650_13878.n79 a_n2650_13878.t46 3.61217
R211 a_n2650_13878.n79 a_n2650_13878.t22 3.61217
R212 a_n2650_13878.n78 a_n2650_13878.t24 3.61217
R213 a_n2650_13878.n78 a_n2650_13878.t30 3.61217
R214 a_n2650_13878.n77 a_n2650_13878.t32 3.61217
R215 a_n2650_13878.n77 a_n2650_13878.t18 3.61217
R216 a_n2650_13878.n76 a_n2650_13878.t40 3.61217
R217 a_n2650_13878.n76 a_n2650_13878.t42 3.61217
R218 a_n2650_13878.t14 a_n2650_13878.n136 3.61217
R219 a_n2650_13878.n136 a_n2650_13878.t44 3.61217
R220 a_n2650_13878.n124 a_n2650_13878.t8 2.82907
R221 a_n2650_13878.n124 a_n2650_13878.t55 2.82907
R222 a_n2650_13878.n125 a_n2650_13878.t7 2.82907
R223 a_n2650_13878.n125 a_n2650_13878.t0 2.82907
R224 a_n2650_13878.n123 a_n2650_13878.t1 2.82907
R225 a_n2650_13878.n123 a_n2650_13878.t54 2.82907
R226 a_n2650_13878.n122 a_n2650_13878.t6 2.82907
R227 a_n2650_13878.n122 a_n2650_13878.t53 2.82907
R228 a_n2650_13878.n120 a_n2650_13878.t5 2.82907
R229 a_n2650_13878.n120 a_n2650_13878.t9 2.82907
R230 a_n2650_13878.n121 a_n2650_13878.t11 2.82907
R231 a_n2650_13878.n121 a_n2650_13878.t4 2.82907
R232 a_n2650_13878.n119 a_n2650_13878.t3 2.82907
R233 a_n2650_13878.n119 a_n2650_13878.t10 2.82907
R234 a_n2650_13878.n118 a_n2650_13878.t2 2.82907
R235 a_n2650_13878.n118 a_n2650_13878.t12 2.82907
R236 a_n2650_13878.n132 a_n2650_13878.n16 1.30542
R237 a_n2650_13878.n13 a_n2650_13878.n14 1.04595
R238 a_n2650_13878.n67 a_n2650_13878.n126 47.835
R239 a_n2650_13878.n60 a_n2650_13878.n112 47.835
R240 a_n2650_13878.n80 a_n2650_13878.n45 47.835
R241 a_n2650_13878.n82 a_n2650_13878.n38 47.835
R242 a_n2650_13878.n0 a_n2650_13878.n2 32.5247
R243 a_n2650_13878.n24 a_n2650_13878.n23 1.13686
R244 a_n2650_13878.n20 a_n2650_13878.n19 1.13686
R245 a_n2650_13878.n7 a_n2650_13878.n6 1.13686
R246 a_n2650_13878.n33 a_n2650_13878.n4 1.11
R247 a_n2650_13878.n1 a_n2650_13878.n0 1.06084
R248 a_n2650_13878.n25 a_n2650_13878.n26 0.758076
R249 a_n2650_13878.n23 a_n2650_13878.n25 0.758076
R250 a_n2650_13878.n21 a_n2650_13878.n22 0.758076
R251 a_n2650_13878.n19 a_n2650_13878.n21 0.758076
R252 a_n2650_13878.n18 a_n2650_13878.n17 0.758076
R253 a_n2650_13878.n15 a_n2650_13878.n14 0.758076
R254 a_n2650_13878.n13 a_n2650_13878.n12 0.758076
R255 a_n2650_13878.n11 a_n2650_13878.n10 0.758076
R256 a_n2650_13878.n9 a_n2650_13878.n8 0.758076
R257 a_n2650_13878.n6 a_n2650_13878.n8 0.758076
R258 a_n2650_13878.n5 a_n2650_13878.n3 0.758076
R259 a_n2650_13878.n4 a_n2650_13878.n3 0.758076
R260 a_n2650_13878.n32 a_n2650_13878.n30 0.716017
R261 a_n2650_13878.n32 a_n2650_13878.n31 0.716017
R262 a_n2650_13878.n29 a_n2650_13878.n28 0.716017
R263 a_n2650_13878.n28 a_n2650_13878.n27 0.716017
R264 a_n2650_13878.n15 a_n2650_13878.n17 0.67853
R265 a_n2650_13878.n11 a_n2650_13878.n12 0.67853
R266 a_n2472_13878.n25 a_n2472_13878.n24 98.9632
R267 a_n2472_13878.n2 a_n2472_13878.n0 98.7517
R268 a_n2472_13878.n20 a_n2472_13878.n19 98.6055
R269 a_n2472_13878.n22 a_n2472_13878.n21 98.6055
R270 a_n2472_13878.n24 a_n2472_13878.n23 98.6055
R271 a_n2472_13878.n8 a_n2472_13878.n7 98.6055
R272 a_n2472_13878.n6 a_n2472_13878.n5 98.6055
R273 a_n2472_13878.n4 a_n2472_13878.n3 98.6055
R274 a_n2472_13878.n2 a_n2472_13878.n1 98.6055
R275 a_n2472_13878.n18 a_n2472_13878.n17 98.6054
R276 a_n2472_13878.n10 a_n2472_13878.t2 74.6477
R277 a_n2472_13878.n15 a_n2472_13878.t3 74.2899
R278 a_n2472_13878.n12 a_n2472_13878.t1 74.2899
R279 a_n2472_13878.n11 a_n2472_13878.t27 74.2899
R280 a_n2472_13878.n14 a_n2472_13878.n13 70.6783
R281 a_n2472_13878.n10 a_n2472_13878.n9 70.6783
R282 a_n2472_13878.n16 a_n2472_13878.n8 15.0004
R283 a_n2472_13878.n18 a_n2472_13878.n16 12.2917
R284 a_n2472_13878.n16 a_n2472_13878.n15 7.67184
R285 a_n2472_13878.n17 a_n2472_13878.t20 3.61217
R286 a_n2472_13878.n17 a_n2472_13878.t9 3.61217
R287 a_n2472_13878.n19 a_n2472_13878.t12 3.61217
R288 a_n2472_13878.n19 a_n2472_13878.t13 3.61217
R289 a_n2472_13878.n21 a_n2472_13878.t21 3.61217
R290 a_n2472_13878.n21 a_n2472_13878.t22 3.61217
R291 a_n2472_13878.n23 a_n2472_13878.t4 3.61217
R292 a_n2472_13878.n23 a_n2472_13878.t14 3.61217
R293 a_n2472_13878.n13 a_n2472_13878.t0 3.61217
R294 a_n2472_13878.n13 a_n2472_13878.t26 3.61217
R295 a_n2472_13878.n9 a_n2472_13878.t24 3.61217
R296 a_n2472_13878.n9 a_n2472_13878.t25 3.61217
R297 a_n2472_13878.n7 a_n2472_13878.t15 3.61217
R298 a_n2472_13878.n7 a_n2472_13878.t5 3.61217
R299 a_n2472_13878.n5 a_n2472_13878.t18 3.61217
R300 a_n2472_13878.n5 a_n2472_13878.t7 3.61217
R301 a_n2472_13878.n3 a_n2472_13878.t6 3.61217
R302 a_n2472_13878.n3 a_n2472_13878.t8 3.61217
R303 a_n2472_13878.n1 a_n2472_13878.t16 3.61217
R304 a_n2472_13878.n1 a_n2472_13878.t10 3.61217
R305 a_n2472_13878.n0 a_n2472_13878.t19 3.61217
R306 a_n2472_13878.n0 a_n2472_13878.t11 3.61217
R307 a_n2472_13878.n25 a_n2472_13878.t17 3.61217
R308 a_n2472_13878.t23 a_n2472_13878.n25 3.61217
R309 a_n2472_13878.n11 a_n2472_13878.n10 0.358259
R310 a_n2472_13878.n14 a_n2472_13878.n12 0.358259
R311 a_n2472_13878.n15 a_n2472_13878.n14 0.358259
R312 a_n2472_13878.n24 a_n2472_13878.n22 0.358259
R313 a_n2472_13878.n22 a_n2472_13878.n20 0.358259
R314 a_n2472_13878.n20 a_n2472_13878.n18 0.358259
R315 a_n2472_13878.n4 a_n2472_13878.n2 0.146627
R316 a_n2472_13878.n6 a_n2472_13878.n4 0.146627
R317 a_n2472_13878.n8 a_n2472_13878.n6 0.146627
R318 a_n2472_13878.n12 a_n2472_13878.n11 0.101793
R319 vdd.n303 vdd.n267 756.745
R320 vdd.n252 vdd.n216 756.745
R321 vdd.n209 vdd.n173 756.745
R322 vdd.n158 vdd.n122 756.745
R323 vdd.n116 vdd.n80 756.745
R324 vdd.n65 vdd.n29 756.745
R325 vdd.n1578 vdd.n1542 756.745
R326 vdd.n1629 vdd.n1593 756.745
R327 vdd.n1484 vdd.n1448 756.745
R328 vdd.n1535 vdd.n1499 756.745
R329 vdd.n1391 vdd.n1355 756.745
R330 vdd.n1442 vdd.n1406 756.745
R331 vdd.n964 vdd.t102 640.208
R332 vdd.n825 vdd.t140 640.208
R333 vdd.n958 vdd.t164 640.208
R334 vdd.n816 vdd.t158 640.208
R335 vdd.n713 vdd.t109 640.208
R336 vdd.n2473 vdd.t155 640.208
R337 vdd.n661 vdd.t134 640.208
R338 vdd.n2542 vdd.t144 640.208
R339 vdd.n625 vdd.t98 640.208
R340 vdd.n886 vdd.t151 640.208
R341 vdd.n1190 vdd.t128 592.009
R342 vdd.n1227 vdd.t120 592.009
R343 vdd.n1101 vdd.t131 592.009
R344 vdd.n1912 vdd.t116 592.009
R345 vdd.n1762 vdd.t137 592.009
R346 vdd.n1722 vdd.t148 592.009
R347 vdd.n3203 vdd.t124 592.009
R348 vdd.n427 vdd.t161 592.009
R349 vdd.n387 vdd.t167 592.009
R350 vdd.n580 vdd.t94 592.009
R351 vdd.n543 vdd.t106 592.009
R352 vdd.n2990 vdd.t113 592.009
R353 vdd.n304 vdd.n303 585
R354 vdd.n302 vdd.n269 585
R355 vdd.n301 vdd.n300 585
R356 vdd.n272 vdd.n270 585
R357 vdd.n295 vdd.n294 585
R358 vdd.n293 vdd.n292 585
R359 vdd.n276 vdd.n275 585
R360 vdd.n287 vdd.n286 585
R361 vdd.n285 vdd.n284 585
R362 vdd.n280 vdd.n279 585
R363 vdd.n253 vdd.n252 585
R364 vdd.n251 vdd.n218 585
R365 vdd.n250 vdd.n249 585
R366 vdd.n221 vdd.n219 585
R367 vdd.n244 vdd.n243 585
R368 vdd.n242 vdd.n241 585
R369 vdd.n225 vdd.n224 585
R370 vdd.n236 vdd.n235 585
R371 vdd.n234 vdd.n233 585
R372 vdd.n229 vdd.n228 585
R373 vdd.n210 vdd.n209 585
R374 vdd.n208 vdd.n175 585
R375 vdd.n207 vdd.n206 585
R376 vdd.n178 vdd.n176 585
R377 vdd.n201 vdd.n200 585
R378 vdd.n199 vdd.n198 585
R379 vdd.n182 vdd.n181 585
R380 vdd.n193 vdd.n192 585
R381 vdd.n191 vdd.n190 585
R382 vdd.n186 vdd.n185 585
R383 vdd.n159 vdd.n158 585
R384 vdd.n157 vdd.n124 585
R385 vdd.n156 vdd.n155 585
R386 vdd.n127 vdd.n125 585
R387 vdd.n150 vdd.n149 585
R388 vdd.n148 vdd.n147 585
R389 vdd.n131 vdd.n130 585
R390 vdd.n142 vdd.n141 585
R391 vdd.n140 vdd.n139 585
R392 vdd.n135 vdd.n134 585
R393 vdd.n117 vdd.n116 585
R394 vdd.n115 vdd.n82 585
R395 vdd.n114 vdd.n113 585
R396 vdd.n85 vdd.n83 585
R397 vdd.n108 vdd.n107 585
R398 vdd.n106 vdd.n105 585
R399 vdd.n89 vdd.n88 585
R400 vdd.n100 vdd.n99 585
R401 vdd.n98 vdd.n97 585
R402 vdd.n93 vdd.n92 585
R403 vdd.n66 vdd.n65 585
R404 vdd.n64 vdd.n31 585
R405 vdd.n63 vdd.n62 585
R406 vdd.n34 vdd.n32 585
R407 vdd.n57 vdd.n56 585
R408 vdd.n55 vdd.n54 585
R409 vdd.n38 vdd.n37 585
R410 vdd.n49 vdd.n48 585
R411 vdd.n47 vdd.n46 585
R412 vdd.n42 vdd.n41 585
R413 vdd.n1579 vdd.n1578 585
R414 vdd.n1577 vdd.n1544 585
R415 vdd.n1576 vdd.n1575 585
R416 vdd.n1547 vdd.n1545 585
R417 vdd.n1570 vdd.n1569 585
R418 vdd.n1568 vdd.n1567 585
R419 vdd.n1551 vdd.n1550 585
R420 vdd.n1562 vdd.n1561 585
R421 vdd.n1560 vdd.n1559 585
R422 vdd.n1555 vdd.n1554 585
R423 vdd.n1630 vdd.n1629 585
R424 vdd.n1628 vdd.n1595 585
R425 vdd.n1627 vdd.n1626 585
R426 vdd.n1598 vdd.n1596 585
R427 vdd.n1621 vdd.n1620 585
R428 vdd.n1619 vdd.n1618 585
R429 vdd.n1602 vdd.n1601 585
R430 vdd.n1613 vdd.n1612 585
R431 vdd.n1611 vdd.n1610 585
R432 vdd.n1606 vdd.n1605 585
R433 vdd.n1485 vdd.n1484 585
R434 vdd.n1483 vdd.n1450 585
R435 vdd.n1482 vdd.n1481 585
R436 vdd.n1453 vdd.n1451 585
R437 vdd.n1476 vdd.n1475 585
R438 vdd.n1474 vdd.n1473 585
R439 vdd.n1457 vdd.n1456 585
R440 vdd.n1468 vdd.n1467 585
R441 vdd.n1466 vdd.n1465 585
R442 vdd.n1461 vdd.n1460 585
R443 vdd.n1536 vdd.n1535 585
R444 vdd.n1534 vdd.n1501 585
R445 vdd.n1533 vdd.n1532 585
R446 vdd.n1504 vdd.n1502 585
R447 vdd.n1527 vdd.n1526 585
R448 vdd.n1525 vdd.n1524 585
R449 vdd.n1508 vdd.n1507 585
R450 vdd.n1519 vdd.n1518 585
R451 vdd.n1517 vdd.n1516 585
R452 vdd.n1512 vdd.n1511 585
R453 vdd.n1392 vdd.n1391 585
R454 vdd.n1390 vdd.n1357 585
R455 vdd.n1389 vdd.n1388 585
R456 vdd.n1360 vdd.n1358 585
R457 vdd.n1383 vdd.n1382 585
R458 vdd.n1381 vdd.n1380 585
R459 vdd.n1364 vdd.n1363 585
R460 vdd.n1375 vdd.n1374 585
R461 vdd.n1373 vdd.n1372 585
R462 vdd.n1368 vdd.n1367 585
R463 vdd.n1443 vdd.n1442 585
R464 vdd.n1441 vdd.n1408 585
R465 vdd.n1440 vdd.n1439 585
R466 vdd.n1411 vdd.n1409 585
R467 vdd.n1434 vdd.n1433 585
R468 vdd.n1432 vdd.n1431 585
R469 vdd.n1415 vdd.n1414 585
R470 vdd.n1426 vdd.n1425 585
R471 vdd.n1424 vdd.n1423 585
R472 vdd.n1419 vdd.n1418 585
R473 vdd.n3319 vdd.n352 488.781
R474 vdd.n3201 vdd.n350 488.781
R475 vdd.n3123 vdd.n515 488.781
R476 vdd.n3121 vdd.n517 488.781
R477 vdd.n1907 vdd.n983 488.781
R478 vdd.n1910 vdd.n1909 488.781
R479 vdd.n1296 vdd.n1061 488.781
R480 vdd.n1294 vdd.n1064 488.781
R481 vdd.n281 vdd.t1 329.043
R482 vdd.n230 vdd.t78 329.043
R483 vdd.n187 vdd.t46 329.043
R484 vdd.n136 vdd.t229 329.043
R485 vdd.n94 vdd.t173 329.043
R486 vdd.n43 vdd.t15 329.043
R487 vdd.n1556 vdd.t5 329.043
R488 vdd.n1607 vdd.t87 329.043
R489 vdd.n1462 vdd.t75 329.043
R490 vdd.n1513 vdd.t91 329.043
R491 vdd.n1369 vdd.t236 329.043
R492 vdd.n1420 vdd.t32 329.043
R493 vdd.n1190 vdd.t130 319.788
R494 vdd.n1227 vdd.t123 319.788
R495 vdd.n1101 vdd.t133 319.788
R496 vdd.n1912 vdd.t118 319.788
R497 vdd.n1762 vdd.t138 319.788
R498 vdd.n1722 vdd.t149 319.788
R499 vdd.n3203 vdd.t126 319.788
R500 vdd.n427 vdd.t162 319.788
R501 vdd.n387 vdd.t168 319.788
R502 vdd.n580 vdd.t97 319.788
R503 vdd.n543 vdd.t108 319.788
R504 vdd.n2990 vdd.t115 319.788
R505 vdd.n1191 vdd.t129 303.69
R506 vdd.n1228 vdd.t122 303.69
R507 vdd.n1102 vdd.t132 303.69
R508 vdd.n1913 vdd.t119 303.69
R509 vdd.n1763 vdd.t139 303.69
R510 vdd.n1723 vdd.t150 303.69
R511 vdd.n3204 vdd.t127 303.69
R512 vdd.n428 vdd.t163 303.69
R513 vdd.n388 vdd.t169 303.69
R514 vdd.n581 vdd.t96 303.69
R515 vdd.n544 vdd.t107 303.69
R516 vdd.n2991 vdd.t114 303.69
R517 vdd.n2728 vdd.n775 285.366
R518 vdd.n2952 vdd.n635 285.366
R519 vdd.n2889 vdd.n632 285.366
R520 vdd.n2607 vdd.n772 285.366
R521 vdd.n2437 vdd.n813 285.366
R522 vdd.n2368 vdd.n2367 285.366
R523 vdd.n2108 vdd.n939 285.366
R524 vdd.n2178 vdd.n941 285.366
R525 vdd.n2868 vdd.n633 285.366
R526 vdd.n2955 vdd.n2954 285.366
R527 vdd.n2721 vdd.n773 285.366
R528 vdd.n2730 vdd.n771 285.366
R529 vdd.n2365 vdd.n823 285.366
R530 vdd.n821 vdd.n795 285.366
R531 vdd.n1994 vdd.n940 285.366
R532 vdd.n2180 vdd.n937 285.366
R533 vdd.n981 vdd.n938 216.982
R534 vdd.n613 vdd.n516 216.982
R535 vdd.n2870 vdd.n633 185
R536 vdd.n2953 vdd.n633 185
R537 vdd.n2872 vdd.n2871 185
R538 vdd.n2871 vdd.n631 185
R539 vdd.n2873 vdd.n667 185
R540 vdd.n2883 vdd.n667 185
R541 vdd.n2874 vdd.n676 185
R542 vdd.n676 vdd.n674 185
R543 vdd.n2876 vdd.n2875 185
R544 vdd.n2877 vdd.n2876 185
R545 vdd.n2829 vdd.n675 185
R546 vdd.n675 vdd.n671 185
R547 vdd.n2828 vdd.n2827 185
R548 vdd.n2827 vdd.n2826 185
R549 vdd.n678 vdd.n677 185
R550 vdd.n679 vdd.n678 185
R551 vdd.n2819 vdd.n2818 185
R552 vdd.n2820 vdd.n2819 185
R553 vdd.n2817 vdd.n687 185
R554 vdd.n692 vdd.n687 185
R555 vdd.n2816 vdd.n2815 185
R556 vdd.n2815 vdd.n2814 185
R557 vdd.n689 vdd.n688 185
R558 vdd.n698 vdd.n689 185
R559 vdd.n2807 vdd.n2806 185
R560 vdd.n2808 vdd.n2807 185
R561 vdd.n2805 vdd.n699 185
R562 vdd.n705 vdd.n699 185
R563 vdd.n2804 vdd.n2803 185
R564 vdd.n2803 vdd.n2802 185
R565 vdd.n701 vdd.n700 185
R566 vdd.n702 vdd.n701 185
R567 vdd.n2795 vdd.n2794 185
R568 vdd.n2796 vdd.n2795 185
R569 vdd.n2793 vdd.n712 185
R570 vdd.n712 vdd.n709 185
R571 vdd.n2791 vdd.n2790 185
R572 vdd.n2790 vdd.n2789 185
R573 vdd.n715 vdd.n714 185
R574 vdd.n716 vdd.n715 185
R575 vdd.n2782 vdd.n2781 185
R576 vdd.n2783 vdd.n2782 185
R577 vdd.n2780 vdd.n724 185
R578 vdd.n729 vdd.n724 185
R579 vdd.n2779 vdd.n2778 185
R580 vdd.n2778 vdd.n2777 185
R581 vdd.n726 vdd.n725 185
R582 vdd.n2689 vdd.n726 185
R583 vdd.n2770 vdd.n2769 185
R584 vdd.n2771 vdd.n2770 185
R585 vdd.n2768 vdd.n736 185
R586 vdd.n736 vdd.n733 185
R587 vdd.n2767 vdd.n2766 185
R588 vdd.n2766 vdd.n2765 185
R589 vdd.n738 vdd.n737 185
R590 vdd.n739 vdd.n738 185
R591 vdd.n2758 vdd.n2757 185
R592 vdd.n2759 vdd.n2758 185
R593 vdd.n2756 vdd.n747 185
R594 vdd.n2701 vdd.n747 185
R595 vdd.n2755 vdd.n2754 185
R596 vdd.n2754 vdd.n2753 185
R597 vdd.n749 vdd.n748 185
R598 vdd.n758 vdd.n749 185
R599 vdd.n2746 vdd.n2745 185
R600 vdd.n2747 vdd.n2746 185
R601 vdd.n2744 vdd.n759 185
R602 vdd.n759 vdd.n755 185
R603 vdd.n2743 vdd.n2742 185
R604 vdd.n2742 vdd.n2741 185
R605 vdd.n761 vdd.n760 185
R606 vdd.n2713 vdd.n761 185
R607 vdd.n2734 vdd.n2733 185
R608 vdd.n2735 vdd.n2734 185
R609 vdd.n2732 vdd.n769 185
R610 vdd.n774 vdd.n769 185
R611 vdd.n2731 vdd.n2730 185
R612 vdd.n2730 vdd.n2729 185
R613 vdd.n771 vdd.n770 185
R614 vdd.n2477 vdd.n2476 185
R615 vdd.n2479 vdd.n2478 185
R616 vdd.n2481 vdd.n2480 185
R617 vdd.n2483 vdd.n2482 185
R618 vdd.n2485 vdd.n2484 185
R619 vdd.n2487 vdd.n2486 185
R620 vdd.n2489 vdd.n2488 185
R621 vdd.n2491 vdd.n2490 185
R622 vdd.n2493 vdd.n2492 185
R623 vdd.n2495 vdd.n2494 185
R624 vdd.n2497 vdd.n2496 185
R625 vdd.n2499 vdd.n2498 185
R626 vdd.n2501 vdd.n2500 185
R627 vdd.n2503 vdd.n2502 185
R628 vdd.n2505 vdd.n2504 185
R629 vdd.n2507 vdd.n2506 185
R630 vdd.n2509 vdd.n2508 185
R631 vdd.n2511 vdd.n2510 185
R632 vdd.n2513 vdd.n2512 185
R633 vdd.n2515 vdd.n2514 185
R634 vdd.n2517 vdd.n2516 185
R635 vdd.n2519 vdd.n2518 185
R636 vdd.n2521 vdd.n2520 185
R637 vdd.n2523 vdd.n2522 185
R638 vdd.n2525 vdd.n2524 185
R639 vdd.n2527 vdd.n2526 185
R640 vdd.n2529 vdd.n2528 185
R641 vdd.n2531 vdd.n2530 185
R642 vdd.n2533 vdd.n2532 185
R643 vdd.n2535 vdd.n2534 185
R644 vdd.n2537 vdd.n2536 185
R645 vdd.n2539 vdd.n2538 185
R646 vdd.n2540 vdd.n2472 185
R647 vdd.n2721 vdd.n2720 185
R648 vdd.n2722 vdd.n2721 185
R649 vdd.n2956 vdd.n2955 185
R650 vdd.n2957 vdd.n624 185
R651 vdd.n2959 vdd.n2958 185
R652 vdd.n2961 vdd.n622 185
R653 vdd.n2963 vdd.n2962 185
R654 vdd.n2964 vdd.n621 185
R655 vdd.n2966 vdd.n2965 185
R656 vdd.n2968 vdd.n619 185
R657 vdd.n2970 vdd.n2969 185
R658 vdd.n2971 vdd.n618 185
R659 vdd.n2973 vdd.n2972 185
R660 vdd.n2975 vdd.n616 185
R661 vdd.n2977 vdd.n2976 185
R662 vdd.n2978 vdd.n615 185
R663 vdd.n2980 vdd.n2979 185
R664 vdd.n2982 vdd.n614 185
R665 vdd.n2983 vdd.n611 185
R666 vdd.n2986 vdd.n2985 185
R667 vdd.n612 vdd.n610 185
R668 vdd.n2842 vdd.n2841 185
R669 vdd.n2844 vdd.n2843 185
R670 vdd.n2846 vdd.n2838 185
R671 vdd.n2848 vdd.n2847 185
R672 vdd.n2849 vdd.n2837 185
R673 vdd.n2851 vdd.n2850 185
R674 vdd.n2853 vdd.n2835 185
R675 vdd.n2855 vdd.n2854 185
R676 vdd.n2856 vdd.n2834 185
R677 vdd.n2858 vdd.n2857 185
R678 vdd.n2860 vdd.n2832 185
R679 vdd.n2862 vdd.n2861 185
R680 vdd.n2863 vdd.n2831 185
R681 vdd.n2865 vdd.n2864 185
R682 vdd.n2867 vdd.n2830 185
R683 vdd.n2869 vdd.n2868 185
R684 vdd.n2868 vdd.n613 185
R685 vdd.n2954 vdd.n628 185
R686 vdd.n2954 vdd.n2953 185
R687 vdd.n2620 vdd.n630 185
R688 vdd.n631 vdd.n630 185
R689 vdd.n2621 vdd.n666 185
R690 vdd.n2883 vdd.n666 185
R691 vdd.n2623 vdd.n2622 185
R692 vdd.n2622 vdd.n674 185
R693 vdd.n2624 vdd.n673 185
R694 vdd.n2877 vdd.n673 185
R695 vdd.n2626 vdd.n2625 185
R696 vdd.n2625 vdd.n671 185
R697 vdd.n2627 vdd.n681 185
R698 vdd.n2826 vdd.n681 185
R699 vdd.n2629 vdd.n2628 185
R700 vdd.n2628 vdd.n679 185
R701 vdd.n2630 vdd.n686 185
R702 vdd.n2820 vdd.n686 185
R703 vdd.n2632 vdd.n2631 185
R704 vdd.n2631 vdd.n692 185
R705 vdd.n2633 vdd.n691 185
R706 vdd.n2814 vdd.n691 185
R707 vdd.n2635 vdd.n2634 185
R708 vdd.n2634 vdd.n698 185
R709 vdd.n2636 vdd.n697 185
R710 vdd.n2808 vdd.n697 185
R711 vdd.n2638 vdd.n2637 185
R712 vdd.n2637 vdd.n705 185
R713 vdd.n2639 vdd.n704 185
R714 vdd.n2802 vdd.n704 185
R715 vdd.n2641 vdd.n2640 185
R716 vdd.n2640 vdd.n702 185
R717 vdd.n2642 vdd.n711 185
R718 vdd.n2796 vdd.n711 185
R719 vdd.n2644 vdd.n2643 185
R720 vdd.n2643 vdd.n709 185
R721 vdd.n2645 vdd.n718 185
R722 vdd.n2789 vdd.n718 185
R723 vdd.n2647 vdd.n2646 185
R724 vdd.n2646 vdd.n716 185
R725 vdd.n2648 vdd.n723 185
R726 vdd.n2783 vdd.n723 185
R727 vdd.n2650 vdd.n2649 185
R728 vdd.n2649 vdd.n729 185
R729 vdd.n2651 vdd.n728 185
R730 vdd.n2777 vdd.n728 185
R731 vdd.n2691 vdd.n2690 185
R732 vdd.n2690 vdd.n2689 185
R733 vdd.n2692 vdd.n735 185
R734 vdd.n2771 vdd.n735 185
R735 vdd.n2694 vdd.n2693 185
R736 vdd.n2693 vdd.n733 185
R737 vdd.n2695 vdd.n741 185
R738 vdd.n2765 vdd.n741 185
R739 vdd.n2697 vdd.n2696 185
R740 vdd.n2696 vdd.n739 185
R741 vdd.n2698 vdd.n746 185
R742 vdd.n2759 vdd.n746 185
R743 vdd.n2700 vdd.n2699 185
R744 vdd.n2701 vdd.n2700 185
R745 vdd.n2619 vdd.n751 185
R746 vdd.n2753 vdd.n751 185
R747 vdd.n2618 vdd.n2617 185
R748 vdd.n2617 vdd.n758 185
R749 vdd.n2616 vdd.n757 185
R750 vdd.n2747 vdd.n757 185
R751 vdd.n2615 vdd.n2614 185
R752 vdd.n2614 vdd.n755 185
R753 vdd.n2541 vdd.n763 185
R754 vdd.n2741 vdd.n763 185
R755 vdd.n2715 vdd.n2714 185
R756 vdd.n2714 vdd.n2713 185
R757 vdd.n2716 vdd.n768 185
R758 vdd.n2735 vdd.n768 185
R759 vdd.n2718 vdd.n2717 185
R760 vdd.n2717 vdd.n774 185
R761 vdd.n2719 vdd.n773 185
R762 vdd.n2729 vdd.n773 185
R763 vdd.n1907 vdd.n1906 185
R764 vdd.n1908 vdd.n1907 185
R765 vdd.n984 vdd.n982 185
R766 vdd.n1686 vdd.n982 185
R767 vdd.n1689 vdd.n1688 185
R768 vdd.n1688 vdd.n1687 185
R769 vdd.n987 vdd.n986 185
R770 vdd.n988 vdd.n987 185
R771 vdd.n1675 vdd.n1674 185
R772 vdd.n1676 vdd.n1675 185
R773 vdd.n996 vdd.n995 185
R774 vdd.n1667 vdd.n995 185
R775 vdd.n1670 vdd.n1669 185
R776 vdd.n1669 vdd.n1668 185
R777 vdd.n999 vdd.n998 185
R778 vdd.n1005 vdd.n999 185
R779 vdd.n1658 vdd.n1657 185
R780 vdd.n1659 vdd.n1658 185
R781 vdd.n1007 vdd.n1006 185
R782 vdd.n1650 vdd.n1006 185
R783 vdd.n1653 vdd.n1652 185
R784 vdd.n1652 vdd.n1651 185
R785 vdd.n1010 vdd.n1009 185
R786 vdd.n1011 vdd.n1010 185
R787 vdd.n1641 vdd.n1640 185
R788 vdd.n1642 vdd.n1641 185
R789 vdd.n1019 vdd.n1018 185
R790 vdd.n1018 vdd.n1017 185
R791 vdd.n1354 vdd.n1353 185
R792 vdd.n1353 vdd.n1352 185
R793 vdd.n1022 vdd.n1021 185
R794 vdd.n1028 vdd.n1022 185
R795 vdd.n1343 vdd.n1342 185
R796 vdd.n1344 vdd.n1343 185
R797 vdd.n1030 vdd.n1029 185
R798 vdd.n1335 vdd.n1029 185
R799 vdd.n1338 vdd.n1337 185
R800 vdd.n1337 vdd.n1336 185
R801 vdd.n1033 vdd.n1032 185
R802 vdd.n1040 vdd.n1033 185
R803 vdd.n1326 vdd.n1325 185
R804 vdd.n1327 vdd.n1326 185
R805 vdd.n1042 vdd.n1041 185
R806 vdd.n1041 vdd.n1039 185
R807 vdd.n1321 vdd.n1320 185
R808 vdd.n1320 vdd.n1319 185
R809 vdd.n1045 vdd.n1044 185
R810 vdd.n1046 vdd.n1045 185
R811 vdd.n1310 vdd.n1309 185
R812 vdd.n1311 vdd.n1310 185
R813 vdd.n1054 vdd.n1053 185
R814 vdd.n1053 vdd.n1052 185
R815 vdd.n1305 vdd.n1304 185
R816 vdd.n1304 vdd.n1303 185
R817 vdd.n1057 vdd.n1056 185
R818 vdd.n1063 vdd.n1057 185
R819 vdd.n1294 vdd.n1293 185
R820 vdd.n1295 vdd.n1294 185
R821 vdd.n1290 vdd.n1064 185
R822 vdd.n1289 vdd.n1067 185
R823 vdd.n1288 vdd.n1068 185
R824 vdd.n1068 vdd.n1062 185
R825 vdd.n1071 vdd.n1069 185
R826 vdd.n1284 vdd.n1073 185
R827 vdd.n1283 vdd.n1074 185
R828 vdd.n1282 vdd.n1076 185
R829 vdd.n1079 vdd.n1077 185
R830 vdd.n1278 vdd.n1081 185
R831 vdd.n1277 vdd.n1082 185
R832 vdd.n1276 vdd.n1084 185
R833 vdd.n1087 vdd.n1085 185
R834 vdd.n1272 vdd.n1089 185
R835 vdd.n1271 vdd.n1090 185
R836 vdd.n1270 vdd.n1092 185
R837 vdd.n1095 vdd.n1093 185
R838 vdd.n1266 vdd.n1097 185
R839 vdd.n1265 vdd.n1098 185
R840 vdd.n1264 vdd.n1100 185
R841 vdd.n1105 vdd.n1103 185
R842 vdd.n1260 vdd.n1107 185
R843 vdd.n1259 vdd.n1108 185
R844 vdd.n1258 vdd.n1110 185
R845 vdd.n1113 vdd.n1111 185
R846 vdd.n1254 vdd.n1115 185
R847 vdd.n1253 vdd.n1116 185
R848 vdd.n1252 vdd.n1118 185
R849 vdd.n1121 vdd.n1119 185
R850 vdd.n1248 vdd.n1123 185
R851 vdd.n1247 vdd.n1124 185
R852 vdd.n1246 vdd.n1126 185
R853 vdd.n1129 vdd.n1127 185
R854 vdd.n1242 vdd.n1131 185
R855 vdd.n1241 vdd.n1132 185
R856 vdd.n1240 vdd.n1134 185
R857 vdd.n1137 vdd.n1135 185
R858 vdd.n1236 vdd.n1139 185
R859 vdd.n1235 vdd.n1140 185
R860 vdd.n1234 vdd.n1142 185
R861 vdd.n1145 vdd.n1143 185
R862 vdd.n1230 vdd.n1147 185
R863 vdd.n1229 vdd.n1226 185
R864 vdd.n1224 vdd.n1148 185
R865 vdd.n1223 vdd.n1222 185
R866 vdd.n1153 vdd.n1150 185
R867 vdd.n1218 vdd.n1154 185
R868 vdd.n1217 vdd.n1156 185
R869 vdd.n1216 vdd.n1157 185
R870 vdd.n1161 vdd.n1158 185
R871 vdd.n1212 vdd.n1162 185
R872 vdd.n1211 vdd.n1164 185
R873 vdd.n1210 vdd.n1165 185
R874 vdd.n1169 vdd.n1166 185
R875 vdd.n1206 vdd.n1170 185
R876 vdd.n1205 vdd.n1172 185
R877 vdd.n1204 vdd.n1173 185
R878 vdd.n1177 vdd.n1174 185
R879 vdd.n1200 vdd.n1178 185
R880 vdd.n1199 vdd.n1180 185
R881 vdd.n1198 vdd.n1181 185
R882 vdd.n1185 vdd.n1182 185
R883 vdd.n1194 vdd.n1186 185
R884 vdd.n1193 vdd.n1188 185
R885 vdd.n1189 vdd.n1061 185
R886 vdd.n1062 vdd.n1061 185
R887 vdd.n1911 vdd.n1910 185
R888 vdd.n1915 vdd.n977 185
R889 vdd.n1791 vdd.n976 185
R890 vdd.n1794 vdd.n1793 185
R891 vdd.n1796 vdd.n1795 185
R892 vdd.n1799 vdd.n1798 185
R893 vdd.n1801 vdd.n1800 185
R894 vdd.n1803 vdd.n1789 185
R895 vdd.n1805 vdd.n1804 185
R896 vdd.n1806 vdd.n1783 185
R897 vdd.n1808 vdd.n1807 185
R898 vdd.n1810 vdd.n1781 185
R899 vdd.n1812 vdd.n1811 185
R900 vdd.n1813 vdd.n1776 185
R901 vdd.n1815 vdd.n1814 185
R902 vdd.n1817 vdd.n1774 185
R903 vdd.n1819 vdd.n1818 185
R904 vdd.n1820 vdd.n1770 185
R905 vdd.n1822 vdd.n1821 185
R906 vdd.n1824 vdd.n1767 185
R907 vdd.n1826 vdd.n1825 185
R908 vdd.n1768 vdd.n1761 185
R909 vdd.n1830 vdd.n1765 185
R910 vdd.n1831 vdd.n1757 185
R911 vdd.n1833 vdd.n1832 185
R912 vdd.n1835 vdd.n1755 185
R913 vdd.n1837 vdd.n1836 185
R914 vdd.n1838 vdd.n1750 185
R915 vdd.n1840 vdd.n1839 185
R916 vdd.n1842 vdd.n1748 185
R917 vdd.n1844 vdd.n1843 185
R918 vdd.n1845 vdd.n1743 185
R919 vdd.n1847 vdd.n1846 185
R920 vdd.n1849 vdd.n1741 185
R921 vdd.n1851 vdd.n1850 185
R922 vdd.n1852 vdd.n1736 185
R923 vdd.n1854 vdd.n1853 185
R924 vdd.n1856 vdd.n1734 185
R925 vdd.n1858 vdd.n1857 185
R926 vdd.n1859 vdd.n1730 185
R927 vdd.n1861 vdd.n1860 185
R928 vdd.n1863 vdd.n1727 185
R929 vdd.n1865 vdd.n1864 185
R930 vdd.n1728 vdd.n1721 185
R931 vdd.n1869 vdd.n1725 185
R932 vdd.n1870 vdd.n1717 185
R933 vdd.n1872 vdd.n1871 185
R934 vdd.n1874 vdd.n1715 185
R935 vdd.n1876 vdd.n1875 185
R936 vdd.n1877 vdd.n1710 185
R937 vdd.n1879 vdd.n1878 185
R938 vdd.n1881 vdd.n1708 185
R939 vdd.n1883 vdd.n1882 185
R940 vdd.n1884 vdd.n1703 185
R941 vdd.n1886 vdd.n1885 185
R942 vdd.n1888 vdd.n1702 185
R943 vdd.n1889 vdd.n1699 185
R944 vdd.n1892 vdd.n1891 185
R945 vdd.n1701 vdd.n1697 185
R946 vdd.n1896 vdd.n1695 185
R947 vdd.n1898 vdd.n1897 185
R948 vdd.n1900 vdd.n1693 185
R949 vdd.n1902 vdd.n1901 185
R950 vdd.n1903 vdd.n983 185
R951 vdd.n1909 vdd.n980 185
R952 vdd.n1909 vdd.n1908 185
R953 vdd.n991 vdd.n979 185
R954 vdd.n1686 vdd.n979 185
R955 vdd.n1685 vdd.n1684 185
R956 vdd.n1687 vdd.n1685 185
R957 vdd.n990 vdd.n989 185
R958 vdd.n989 vdd.n988 185
R959 vdd.n1678 vdd.n1677 185
R960 vdd.n1677 vdd.n1676 185
R961 vdd.n994 vdd.n993 185
R962 vdd.n1667 vdd.n994 185
R963 vdd.n1666 vdd.n1665 185
R964 vdd.n1668 vdd.n1666 185
R965 vdd.n1001 vdd.n1000 185
R966 vdd.n1005 vdd.n1000 185
R967 vdd.n1661 vdd.n1660 185
R968 vdd.n1660 vdd.n1659 185
R969 vdd.n1004 vdd.n1003 185
R970 vdd.n1650 vdd.n1004 185
R971 vdd.n1649 vdd.n1648 185
R972 vdd.n1651 vdd.n1649 185
R973 vdd.n1013 vdd.n1012 185
R974 vdd.n1012 vdd.n1011 185
R975 vdd.n1644 vdd.n1643 185
R976 vdd.n1643 vdd.n1642 185
R977 vdd.n1016 vdd.n1015 185
R978 vdd.n1017 vdd.n1016 185
R979 vdd.n1351 vdd.n1350 185
R980 vdd.n1352 vdd.n1351 185
R981 vdd.n1024 vdd.n1023 185
R982 vdd.n1028 vdd.n1023 185
R983 vdd.n1346 vdd.n1345 185
R984 vdd.n1345 vdd.n1344 185
R985 vdd.n1027 vdd.n1026 185
R986 vdd.n1335 vdd.n1027 185
R987 vdd.n1334 vdd.n1333 185
R988 vdd.n1336 vdd.n1334 185
R989 vdd.n1035 vdd.n1034 185
R990 vdd.n1040 vdd.n1034 185
R991 vdd.n1329 vdd.n1328 185
R992 vdd.n1328 vdd.n1327 185
R993 vdd.n1038 vdd.n1037 185
R994 vdd.n1039 vdd.n1038 185
R995 vdd.n1318 vdd.n1317 185
R996 vdd.n1319 vdd.n1318 185
R997 vdd.n1048 vdd.n1047 185
R998 vdd.n1047 vdd.n1046 185
R999 vdd.n1313 vdd.n1312 185
R1000 vdd.n1312 vdd.n1311 185
R1001 vdd.n1051 vdd.n1050 185
R1002 vdd.n1052 vdd.n1051 185
R1003 vdd.n1302 vdd.n1301 185
R1004 vdd.n1303 vdd.n1302 185
R1005 vdd.n1059 vdd.n1058 185
R1006 vdd.n1063 vdd.n1058 185
R1007 vdd.n1297 vdd.n1296 185
R1008 vdd.n1296 vdd.n1295 185
R1009 vdd.n815 vdd.n813 185
R1010 vdd.n2366 vdd.n813 185
R1011 vdd.n2288 vdd.n833 185
R1012 vdd.n833 vdd.n820 185
R1013 vdd.n2290 vdd.n2289 185
R1014 vdd.n2291 vdd.n2290 185
R1015 vdd.n2287 vdd.n832 185
R1016 vdd.n2046 vdd.n832 185
R1017 vdd.n2286 vdd.n2285 185
R1018 vdd.n2285 vdd.n2284 185
R1019 vdd.n835 vdd.n834 185
R1020 vdd.n836 vdd.n835 185
R1021 vdd.n2275 vdd.n2274 185
R1022 vdd.n2276 vdd.n2275 185
R1023 vdd.n2273 vdd.n846 185
R1024 vdd.n846 vdd.n843 185
R1025 vdd.n2272 vdd.n2271 185
R1026 vdd.n2271 vdd.n2270 185
R1027 vdd.n848 vdd.n847 185
R1028 vdd.n2058 vdd.n848 185
R1029 vdd.n2263 vdd.n2262 185
R1030 vdd.n2264 vdd.n2263 185
R1031 vdd.n2261 vdd.n856 185
R1032 vdd.n861 vdd.n856 185
R1033 vdd.n2260 vdd.n2259 185
R1034 vdd.n2259 vdd.n2258 185
R1035 vdd.n858 vdd.n857 185
R1036 vdd.n867 vdd.n858 185
R1037 vdd.n2251 vdd.n2250 185
R1038 vdd.n2252 vdd.n2251 185
R1039 vdd.n2249 vdd.n868 185
R1040 vdd.n2070 vdd.n868 185
R1041 vdd.n2248 vdd.n2247 185
R1042 vdd.n2247 vdd.n2246 185
R1043 vdd.n870 vdd.n869 185
R1044 vdd.n871 vdd.n870 185
R1045 vdd.n2239 vdd.n2238 185
R1046 vdd.n2240 vdd.n2239 185
R1047 vdd.n2237 vdd.n880 185
R1048 vdd.n880 vdd.n877 185
R1049 vdd.n2236 vdd.n2235 185
R1050 vdd.n2235 vdd.n2234 185
R1051 vdd.n882 vdd.n881 185
R1052 vdd.n891 vdd.n882 185
R1053 vdd.n2226 vdd.n2225 185
R1054 vdd.n2227 vdd.n2226 185
R1055 vdd.n2224 vdd.n892 185
R1056 vdd.n898 vdd.n892 185
R1057 vdd.n2223 vdd.n2222 185
R1058 vdd.n2222 vdd.n2221 185
R1059 vdd.n894 vdd.n893 185
R1060 vdd.n895 vdd.n894 185
R1061 vdd.n2214 vdd.n2213 185
R1062 vdd.n2215 vdd.n2214 185
R1063 vdd.n2212 vdd.n905 185
R1064 vdd.n905 vdd.n902 185
R1065 vdd.n2211 vdd.n2210 185
R1066 vdd.n2210 vdd.n2209 185
R1067 vdd.n907 vdd.n906 185
R1068 vdd.n908 vdd.n907 185
R1069 vdd.n2202 vdd.n2201 185
R1070 vdd.n2203 vdd.n2202 185
R1071 vdd.n2200 vdd.n917 185
R1072 vdd.n917 vdd.n914 185
R1073 vdd.n2199 vdd.n2198 185
R1074 vdd.n2198 vdd.n2197 185
R1075 vdd.n919 vdd.n918 185
R1076 vdd.n920 vdd.n919 185
R1077 vdd.n2190 vdd.n2189 185
R1078 vdd.n2191 vdd.n2190 185
R1079 vdd.n2188 vdd.n929 185
R1080 vdd.n929 vdd.n926 185
R1081 vdd.n2187 vdd.n2186 185
R1082 vdd.n2186 vdd.n2185 185
R1083 vdd.n931 vdd.n930 185
R1084 vdd.n932 vdd.n931 185
R1085 vdd.n2178 vdd.n2177 185
R1086 vdd.n2179 vdd.n2178 185
R1087 vdd.n2176 vdd.n941 185
R1088 vdd.n2175 vdd.n2174 185
R1089 vdd.n2172 vdd.n942 185
R1090 vdd.n2172 vdd.n938 185
R1091 vdd.n2171 vdd.n2170 185
R1092 vdd.n2169 vdd.n2168 185
R1093 vdd.n2167 vdd.n944 185
R1094 vdd.n2165 vdd.n2164 185
R1095 vdd.n2163 vdd.n945 185
R1096 vdd.n2162 vdd.n2161 185
R1097 vdd.n2159 vdd.n946 185
R1098 vdd.n2157 vdd.n2156 185
R1099 vdd.n2155 vdd.n947 185
R1100 vdd.n2154 vdd.n2153 185
R1101 vdd.n2151 vdd.n948 185
R1102 vdd.n2149 vdd.n2148 185
R1103 vdd.n2147 vdd.n949 185
R1104 vdd.n2146 vdd.n2145 185
R1105 vdd.n2143 vdd.n950 185
R1106 vdd.n2141 vdd.n2140 185
R1107 vdd.n2139 vdd.n951 185
R1108 vdd.n2138 vdd.n2137 185
R1109 vdd.n2135 vdd.n952 185
R1110 vdd.n2133 vdd.n2132 185
R1111 vdd.n2131 vdd.n953 185
R1112 vdd.n2130 vdd.n2129 185
R1113 vdd.n2127 vdd.n954 185
R1114 vdd.n2125 vdd.n2124 185
R1115 vdd.n2123 vdd.n955 185
R1116 vdd.n2122 vdd.n2121 185
R1117 vdd.n2119 vdd.n956 185
R1118 vdd.n2117 vdd.n2116 185
R1119 vdd.n2115 vdd.n957 185
R1120 vdd.n2113 vdd.n2112 185
R1121 vdd.n2110 vdd.n960 185
R1122 vdd.n2108 vdd.n2107 185
R1123 vdd.n2369 vdd.n2368 185
R1124 vdd.n2371 vdd.n2370 185
R1125 vdd.n2373 vdd.n2372 185
R1126 vdd.n2376 vdd.n2375 185
R1127 vdd.n2378 vdd.n2377 185
R1128 vdd.n2380 vdd.n2379 185
R1129 vdd.n2382 vdd.n2381 185
R1130 vdd.n2384 vdd.n2383 185
R1131 vdd.n2386 vdd.n2385 185
R1132 vdd.n2388 vdd.n2387 185
R1133 vdd.n2390 vdd.n2389 185
R1134 vdd.n2392 vdd.n2391 185
R1135 vdd.n2394 vdd.n2393 185
R1136 vdd.n2396 vdd.n2395 185
R1137 vdd.n2398 vdd.n2397 185
R1138 vdd.n2400 vdd.n2399 185
R1139 vdd.n2402 vdd.n2401 185
R1140 vdd.n2404 vdd.n2403 185
R1141 vdd.n2406 vdd.n2405 185
R1142 vdd.n2408 vdd.n2407 185
R1143 vdd.n2410 vdd.n2409 185
R1144 vdd.n2412 vdd.n2411 185
R1145 vdd.n2414 vdd.n2413 185
R1146 vdd.n2416 vdd.n2415 185
R1147 vdd.n2418 vdd.n2417 185
R1148 vdd.n2420 vdd.n2419 185
R1149 vdd.n2422 vdd.n2421 185
R1150 vdd.n2424 vdd.n2423 185
R1151 vdd.n2426 vdd.n2425 185
R1152 vdd.n2428 vdd.n2427 185
R1153 vdd.n2430 vdd.n2429 185
R1154 vdd.n2432 vdd.n2431 185
R1155 vdd.n2434 vdd.n2433 185
R1156 vdd.n2435 vdd.n814 185
R1157 vdd.n2437 vdd.n2436 185
R1158 vdd.n2438 vdd.n2437 185
R1159 vdd.n2367 vdd.n818 185
R1160 vdd.n2367 vdd.n2366 185
R1161 vdd.n2044 vdd.n819 185
R1162 vdd.n820 vdd.n819 185
R1163 vdd.n2045 vdd.n830 185
R1164 vdd.n2291 vdd.n830 185
R1165 vdd.n2048 vdd.n2047 185
R1166 vdd.n2047 vdd.n2046 185
R1167 vdd.n2049 vdd.n837 185
R1168 vdd.n2284 vdd.n837 185
R1169 vdd.n2051 vdd.n2050 185
R1170 vdd.n2050 vdd.n836 185
R1171 vdd.n2052 vdd.n844 185
R1172 vdd.n2276 vdd.n844 185
R1173 vdd.n2054 vdd.n2053 185
R1174 vdd.n2053 vdd.n843 185
R1175 vdd.n2055 vdd.n849 185
R1176 vdd.n2270 vdd.n849 185
R1177 vdd.n2057 vdd.n2056 185
R1178 vdd.n2058 vdd.n2057 185
R1179 vdd.n2043 vdd.n854 185
R1180 vdd.n2264 vdd.n854 185
R1181 vdd.n2042 vdd.n2041 185
R1182 vdd.n2041 vdd.n861 185
R1183 vdd.n2040 vdd.n859 185
R1184 vdd.n2258 vdd.n859 185
R1185 vdd.n2039 vdd.n2038 185
R1186 vdd.n2038 vdd.n867 185
R1187 vdd.n961 vdd.n865 185
R1188 vdd.n2252 vdd.n865 185
R1189 vdd.n2072 vdd.n2071 185
R1190 vdd.n2071 vdd.n2070 185
R1191 vdd.n2073 vdd.n872 185
R1192 vdd.n2246 vdd.n872 185
R1193 vdd.n2075 vdd.n2074 185
R1194 vdd.n2074 vdd.n871 185
R1195 vdd.n2076 vdd.n878 185
R1196 vdd.n2240 vdd.n878 185
R1197 vdd.n2078 vdd.n2077 185
R1198 vdd.n2077 vdd.n877 185
R1199 vdd.n2079 vdd.n883 185
R1200 vdd.n2234 vdd.n883 185
R1201 vdd.n2081 vdd.n2080 185
R1202 vdd.n2080 vdd.n891 185
R1203 vdd.n2082 vdd.n889 185
R1204 vdd.n2227 vdd.n889 185
R1205 vdd.n2084 vdd.n2083 185
R1206 vdd.n2083 vdd.n898 185
R1207 vdd.n2085 vdd.n896 185
R1208 vdd.n2221 vdd.n896 185
R1209 vdd.n2087 vdd.n2086 185
R1210 vdd.n2086 vdd.n895 185
R1211 vdd.n2088 vdd.n903 185
R1212 vdd.n2215 vdd.n903 185
R1213 vdd.n2090 vdd.n2089 185
R1214 vdd.n2089 vdd.n902 185
R1215 vdd.n2091 vdd.n909 185
R1216 vdd.n2209 vdd.n909 185
R1217 vdd.n2093 vdd.n2092 185
R1218 vdd.n2092 vdd.n908 185
R1219 vdd.n2094 vdd.n915 185
R1220 vdd.n2203 vdd.n915 185
R1221 vdd.n2096 vdd.n2095 185
R1222 vdd.n2095 vdd.n914 185
R1223 vdd.n2097 vdd.n921 185
R1224 vdd.n2197 vdd.n921 185
R1225 vdd.n2099 vdd.n2098 185
R1226 vdd.n2098 vdd.n920 185
R1227 vdd.n2100 vdd.n927 185
R1228 vdd.n2191 vdd.n927 185
R1229 vdd.n2102 vdd.n2101 185
R1230 vdd.n2101 vdd.n926 185
R1231 vdd.n2103 vdd.n933 185
R1232 vdd.n2185 vdd.n933 185
R1233 vdd.n2105 vdd.n2104 185
R1234 vdd.n2104 vdd.n932 185
R1235 vdd.n2106 vdd.n939 185
R1236 vdd.n2179 vdd.n939 185
R1237 vdd.n3319 vdd.n3318 185
R1238 vdd.n3320 vdd.n3319 185
R1239 vdd.n347 vdd.n346 185
R1240 vdd.n3321 vdd.n347 185
R1241 vdd.n3324 vdd.n3323 185
R1242 vdd.n3323 vdd.n3322 185
R1243 vdd.n3325 vdd.n341 185
R1244 vdd.n341 vdd.n340 185
R1245 vdd.n3327 vdd.n3326 185
R1246 vdd.n3328 vdd.n3327 185
R1247 vdd.n336 vdd.n335 185
R1248 vdd.n3329 vdd.n336 185
R1249 vdd.n3332 vdd.n3331 185
R1250 vdd.n3331 vdd.n3330 185
R1251 vdd.n3333 vdd.n330 185
R1252 vdd.n330 vdd.n329 185
R1253 vdd.n3335 vdd.n3334 185
R1254 vdd.n3336 vdd.n3335 185
R1255 vdd.n324 vdd.n323 185
R1256 vdd.n3337 vdd.n324 185
R1257 vdd.n3340 vdd.n3339 185
R1258 vdd.n3339 vdd.n3338 185
R1259 vdd.n3341 vdd.n319 185
R1260 vdd.n325 vdd.n319 185
R1261 vdd.n3343 vdd.n3342 185
R1262 vdd.n3344 vdd.n3343 185
R1263 vdd.n315 vdd.n313 185
R1264 vdd.n3345 vdd.n315 185
R1265 vdd.n3348 vdd.n3347 185
R1266 vdd.n3347 vdd.n3346 185
R1267 vdd.n314 vdd.n312 185
R1268 vdd.n481 vdd.n314 185
R1269 vdd.n3170 vdd.n3169 185
R1270 vdd.n3171 vdd.n3170 185
R1271 vdd.n483 vdd.n482 185
R1272 vdd.n3162 vdd.n482 185
R1273 vdd.n3165 vdd.n3164 185
R1274 vdd.n3164 vdd.n3163 185
R1275 vdd.n486 vdd.n485 185
R1276 vdd.n493 vdd.n486 185
R1277 vdd.n3153 vdd.n3152 185
R1278 vdd.n3154 vdd.n3153 185
R1279 vdd.n495 vdd.n494 185
R1280 vdd.n494 vdd.n492 185
R1281 vdd.n3148 vdd.n3147 185
R1282 vdd.n3147 vdd.n3146 185
R1283 vdd.n498 vdd.n497 185
R1284 vdd.n499 vdd.n498 185
R1285 vdd.n3137 vdd.n3136 185
R1286 vdd.n3138 vdd.n3137 185
R1287 vdd.n507 vdd.n506 185
R1288 vdd.n506 vdd.n505 185
R1289 vdd.n3132 vdd.n3131 185
R1290 vdd.n3131 vdd.n3130 185
R1291 vdd.n510 vdd.n509 185
R1292 vdd.n511 vdd.n510 185
R1293 vdd.n3121 vdd.n3120 185
R1294 vdd.n3122 vdd.n3121 185
R1295 vdd.n3117 vdd.n517 185
R1296 vdd.n3116 vdd.n3115 185
R1297 vdd.n3113 vdd.n519 185
R1298 vdd.n3113 vdd.n516 185
R1299 vdd.n3112 vdd.n3111 185
R1300 vdd.n3110 vdd.n3109 185
R1301 vdd.n3108 vdd.n3107 185
R1302 vdd.n3106 vdd.n3105 185
R1303 vdd.n3104 vdd.n525 185
R1304 vdd.n3102 vdd.n3101 185
R1305 vdd.n3100 vdd.n526 185
R1306 vdd.n3099 vdd.n3098 185
R1307 vdd.n3096 vdd.n531 185
R1308 vdd.n3094 vdd.n3093 185
R1309 vdd.n3092 vdd.n532 185
R1310 vdd.n3091 vdd.n3090 185
R1311 vdd.n3088 vdd.n537 185
R1312 vdd.n3086 vdd.n3085 185
R1313 vdd.n3084 vdd.n538 185
R1314 vdd.n3083 vdd.n3082 185
R1315 vdd.n3080 vdd.n545 185
R1316 vdd.n3078 vdd.n3077 185
R1317 vdd.n3076 vdd.n546 185
R1318 vdd.n3075 vdd.n3074 185
R1319 vdd.n3072 vdd.n551 185
R1320 vdd.n3070 vdd.n3069 185
R1321 vdd.n3068 vdd.n552 185
R1322 vdd.n3067 vdd.n3066 185
R1323 vdd.n3064 vdd.n557 185
R1324 vdd.n3062 vdd.n3061 185
R1325 vdd.n3060 vdd.n558 185
R1326 vdd.n3059 vdd.n3058 185
R1327 vdd.n3056 vdd.n563 185
R1328 vdd.n3054 vdd.n3053 185
R1329 vdd.n3052 vdd.n564 185
R1330 vdd.n3051 vdd.n3050 185
R1331 vdd.n3048 vdd.n569 185
R1332 vdd.n3046 vdd.n3045 185
R1333 vdd.n3044 vdd.n570 185
R1334 vdd.n3043 vdd.n3042 185
R1335 vdd.n3040 vdd.n575 185
R1336 vdd.n3038 vdd.n3037 185
R1337 vdd.n3036 vdd.n576 185
R1338 vdd.n585 vdd.n579 185
R1339 vdd.n3032 vdd.n3031 185
R1340 vdd.n3029 vdd.n583 185
R1341 vdd.n3028 vdd.n3027 185
R1342 vdd.n3026 vdd.n3025 185
R1343 vdd.n3024 vdd.n589 185
R1344 vdd.n3022 vdd.n3021 185
R1345 vdd.n3020 vdd.n590 185
R1346 vdd.n3019 vdd.n3018 185
R1347 vdd.n3016 vdd.n595 185
R1348 vdd.n3014 vdd.n3013 185
R1349 vdd.n3012 vdd.n596 185
R1350 vdd.n3011 vdd.n3010 185
R1351 vdd.n3008 vdd.n601 185
R1352 vdd.n3006 vdd.n3005 185
R1353 vdd.n3004 vdd.n602 185
R1354 vdd.n3003 vdd.n3002 185
R1355 vdd.n3000 vdd.n2999 185
R1356 vdd.n2998 vdd.n2997 185
R1357 vdd.n2996 vdd.n2995 185
R1358 vdd.n2994 vdd.n2993 185
R1359 vdd.n2989 vdd.n515 185
R1360 vdd.n516 vdd.n515 185
R1361 vdd.n3202 vdd.n3201 185
R1362 vdd.n3206 vdd.n462 185
R1363 vdd.n3208 vdd.n3207 185
R1364 vdd.n3210 vdd.n460 185
R1365 vdd.n3212 vdd.n3211 185
R1366 vdd.n3213 vdd.n455 185
R1367 vdd.n3215 vdd.n3214 185
R1368 vdd.n3217 vdd.n453 185
R1369 vdd.n3219 vdd.n3218 185
R1370 vdd.n3220 vdd.n448 185
R1371 vdd.n3222 vdd.n3221 185
R1372 vdd.n3224 vdd.n446 185
R1373 vdd.n3226 vdd.n3225 185
R1374 vdd.n3227 vdd.n441 185
R1375 vdd.n3229 vdd.n3228 185
R1376 vdd.n3231 vdd.n439 185
R1377 vdd.n3233 vdd.n3232 185
R1378 vdd.n3234 vdd.n435 185
R1379 vdd.n3236 vdd.n3235 185
R1380 vdd.n3238 vdd.n432 185
R1381 vdd.n3240 vdd.n3239 185
R1382 vdd.n433 vdd.n426 185
R1383 vdd.n3244 vdd.n430 185
R1384 vdd.n3245 vdd.n422 185
R1385 vdd.n3247 vdd.n3246 185
R1386 vdd.n3249 vdd.n420 185
R1387 vdd.n3251 vdd.n3250 185
R1388 vdd.n3252 vdd.n415 185
R1389 vdd.n3254 vdd.n3253 185
R1390 vdd.n3256 vdd.n413 185
R1391 vdd.n3258 vdd.n3257 185
R1392 vdd.n3259 vdd.n408 185
R1393 vdd.n3261 vdd.n3260 185
R1394 vdd.n3263 vdd.n406 185
R1395 vdd.n3265 vdd.n3264 185
R1396 vdd.n3266 vdd.n401 185
R1397 vdd.n3268 vdd.n3267 185
R1398 vdd.n3270 vdd.n399 185
R1399 vdd.n3272 vdd.n3271 185
R1400 vdd.n3273 vdd.n395 185
R1401 vdd.n3275 vdd.n3274 185
R1402 vdd.n3277 vdd.n392 185
R1403 vdd.n3279 vdd.n3278 185
R1404 vdd.n393 vdd.n386 185
R1405 vdd.n3283 vdd.n390 185
R1406 vdd.n3284 vdd.n382 185
R1407 vdd.n3286 vdd.n3285 185
R1408 vdd.n3288 vdd.n380 185
R1409 vdd.n3290 vdd.n3289 185
R1410 vdd.n3291 vdd.n375 185
R1411 vdd.n3293 vdd.n3292 185
R1412 vdd.n3295 vdd.n373 185
R1413 vdd.n3297 vdd.n3296 185
R1414 vdd.n3298 vdd.n368 185
R1415 vdd.n3300 vdd.n3299 185
R1416 vdd.n3302 vdd.n366 185
R1417 vdd.n3304 vdd.n3303 185
R1418 vdd.n3305 vdd.n360 185
R1419 vdd.n3307 vdd.n3306 185
R1420 vdd.n3309 vdd.n359 185
R1421 vdd.n3310 vdd.n358 185
R1422 vdd.n3313 vdd.n3312 185
R1423 vdd.n3314 vdd.n356 185
R1424 vdd.n3315 vdd.n352 185
R1425 vdd.n3197 vdd.n350 185
R1426 vdd.n3320 vdd.n350 185
R1427 vdd.n3196 vdd.n349 185
R1428 vdd.n3321 vdd.n349 185
R1429 vdd.n3195 vdd.n348 185
R1430 vdd.n3322 vdd.n348 185
R1431 vdd.n468 vdd.n467 185
R1432 vdd.n467 vdd.n340 185
R1433 vdd.n3191 vdd.n339 185
R1434 vdd.n3328 vdd.n339 185
R1435 vdd.n3190 vdd.n338 185
R1436 vdd.n3329 vdd.n338 185
R1437 vdd.n3189 vdd.n337 185
R1438 vdd.n3330 vdd.n337 185
R1439 vdd.n471 vdd.n470 185
R1440 vdd.n470 vdd.n329 185
R1441 vdd.n3185 vdd.n328 185
R1442 vdd.n3336 vdd.n328 185
R1443 vdd.n3184 vdd.n327 185
R1444 vdd.n3337 vdd.n327 185
R1445 vdd.n3183 vdd.n326 185
R1446 vdd.n3338 vdd.n326 185
R1447 vdd.n474 vdd.n473 185
R1448 vdd.n473 vdd.n325 185
R1449 vdd.n3179 vdd.n318 185
R1450 vdd.n3344 vdd.n318 185
R1451 vdd.n3178 vdd.n317 185
R1452 vdd.n3345 vdd.n317 185
R1453 vdd.n3177 vdd.n316 185
R1454 vdd.n3346 vdd.n316 185
R1455 vdd.n480 vdd.n476 185
R1456 vdd.n481 vdd.n480 185
R1457 vdd.n3173 vdd.n3172 185
R1458 vdd.n3172 vdd.n3171 185
R1459 vdd.n479 vdd.n478 185
R1460 vdd.n3162 vdd.n479 185
R1461 vdd.n3161 vdd.n3160 185
R1462 vdd.n3163 vdd.n3161 185
R1463 vdd.n488 vdd.n487 185
R1464 vdd.n493 vdd.n487 185
R1465 vdd.n3156 vdd.n3155 185
R1466 vdd.n3155 vdd.n3154 185
R1467 vdd.n491 vdd.n490 185
R1468 vdd.n492 vdd.n491 185
R1469 vdd.n3145 vdd.n3144 185
R1470 vdd.n3146 vdd.n3145 185
R1471 vdd.n501 vdd.n500 185
R1472 vdd.n500 vdd.n499 185
R1473 vdd.n3140 vdd.n3139 185
R1474 vdd.n3139 vdd.n3138 185
R1475 vdd.n504 vdd.n503 185
R1476 vdd.n505 vdd.n504 185
R1477 vdd.n3129 vdd.n3128 185
R1478 vdd.n3130 vdd.n3129 185
R1479 vdd.n513 vdd.n512 185
R1480 vdd.n512 vdd.n511 185
R1481 vdd.n3124 vdd.n3123 185
R1482 vdd.n3123 vdd.n3122 185
R1483 vdd.n2726 vdd.n775 185
R1484 vdd.n2725 vdd.n2724 185
R1485 vdd.n777 vdd.n776 185
R1486 vdd.n2722 vdd.n777 185
R1487 vdd.n2545 vdd.n2544 185
R1488 vdd.n2547 vdd.n2546 185
R1489 vdd.n2549 vdd.n2548 185
R1490 vdd.n2551 vdd.n2550 185
R1491 vdd.n2553 vdd.n2552 185
R1492 vdd.n2555 vdd.n2554 185
R1493 vdd.n2557 vdd.n2556 185
R1494 vdd.n2559 vdd.n2558 185
R1495 vdd.n2561 vdd.n2560 185
R1496 vdd.n2563 vdd.n2562 185
R1497 vdd.n2565 vdd.n2564 185
R1498 vdd.n2567 vdd.n2566 185
R1499 vdd.n2569 vdd.n2568 185
R1500 vdd.n2571 vdd.n2570 185
R1501 vdd.n2573 vdd.n2572 185
R1502 vdd.n2575 vdd.n2574 185
R1503 vdd.n2577 vdd.n2576 185
R1504 vdd.n2579 vdd.n2578 185
R1505 vdd.n2581 vdd.n2580 185
R1506 vdd.n2583 vdd.n2582 185
R1507 vdd.n2585 vdd.n2584 185
R1508 vdd.n2587 vdd.n2586 185
R1509 vdd.n2589 vdd.n2588 185
R1510 vdd.n2591 vdd.n2590 185
R1511 vdd.n2593 vdd.n2592 185
R1512 vdd.n2595 vdd.n2594 185
R1513 vdd.n2597 vdd.n2596 185
R1514 vdd.n2599 vdd.n2598 185
R1515 vdd.n2601 vdd.n2600 185
R1516 vdd.n2604 vdd.n2603 185
R1517 vdd.n2606 vdd.n2605 185
R1518 vdd.n2608 vdd.n2607 185
R1519 vdd.n2890 vdd.n2889 185
R1520 vdd.n2891 vdd.n660 185
R1521 vdd.n2893 vdd.n2892 185
R1522 vdd.n2895 vdd.n658 185
R1523 vdd.n2897 vdd.n2896 185
R1524 vdd.n2898 vdd.n657 185
R1525 vdd.n2900 vdd.n2899 185
R1526 vdd.n2902 vdd.n655 185
R1527 vdd.n2904 vdd.n2903 185
R1528 vdd.n2905 vdd.n654 185
R1529 vdd.n2907 vdd.n2906 185
R1530 vdd.n2909 vdd.n652 185
R1531 vdd.n2911 vdd.n2910 185
R1532 vdd.n2912 vdd.n651 185
R1533 vdd.n2914 vdd.n2913 185
R1534 vdd.n2916 vdd.n649 185
R1535 vdd.n2918 vdd.n2917 185
R1536 vdd.n2920 vdd.n648 185
R1537 vdd.n2922 vdd.n2921 185
R1538 vdd.n2924 vdd.n646 185
R1539 vdd.n2926 vdd.n2925 185
R1540 vdd.n2927 vdd.n645 185
R1541 vdd.n2929 vdd.n2928 185
R1542 vdd.n2931 vdd.n643 185
R1543 vdd.n2933 vdd.n2932 185
R1544 vdd.n2934 vdd.n642 185
R1545 vdd.n2936 vdd.n2935 185
R1546 vdd.n2938 vdd.n640 185
R1547 vdd.n2940 vdd.n2939 185
R1548 vdd.n2941 vdd.n639 185
R1549 vdd.n2943 vdd.n2942 185
R1550 vdd.n2945 vdd.n638 185
R1551 vdd.n2946 vdd.n637 185
R1552 vdd.n2949 vdd.n2948 185
R1553 vdd.n2950 vdd.n635 185
R1554 vdd.n635 vdd.n613 185
R1555 vdd.n2887 vdd.n632 185
R1556 vdd.n2953 vdd.n632 185
R1557 vdd.n2886 vdd.n2885 185
R1558 vdd.n2885 vdd.n631 185
R1559 vdd.n2884 vdd.n664 185
R1560 vdd.n2884 vdd.n2883 185
R1561 vdd.n2658 vdd.n665 185
R1562 vdd.n674 vdd.n665 185
R1563 vdd.n2659 vdd.n672 185
R1564 vdd.n2877 vdd.n672 185
R1565 vdd.n2661 vdd.n2660 185
R1566 vdd.n2660 vdd.n671 185
R1567 vdd.n2662 vdd.n680 185
R1568 vdd.n2826 vdd.n680 185
R1569 vdd.n2664 vdd.n2663 185
R1570 vdd.n2663 vdd.n679 185
R1571 vdd.n2665 vdd.n685 185
R1572 vdd.n2820 vdd.n685 185
R1573 vdd.n2667 vdd.n2666 185
R1574 vdd.n2666 vdd.n692 185
R1575 vdd.n2668 vdd.n690 185
R1576 vdd.n2814 vdd.n690 185
R1577 vdd.n2670 vdd.n2669 185
R1578 vdd.n2669 vdd.n698 185
R1579 vdd.n2671 vdd.n696 185
R1580 vdd.n2808 vdd.n696 185
R1581 vdd.n2673 vdd.n2672 185
R1582 vdd.n2672 vdd.n705 185
R1583 vdd.n2674 vdd.n703 185
R1584 vdd.n2802 vdd.n703 185
R1585 vdd.n2676 vdd.n2675 185
R1586 vdd.n2675 vdd.n702 185
R1587 vdd.n2677 vdd.n710 185
R1588 vdd.n2796 vdd.n710 185
R1589 vdd.n2679 vdd.n2678 185
R1590 vdd.n2678 vdd.n709 185
R1591 vdd.n2680 vdd.n717 185
R1592 vdd.n2789 vdd.n717 185
R1593 vdd.n2682 vdd.n2681 185
R1594 vdd.n2681 vdd.n716 185
R1595 vdd.n2683 vdd.n722 185
R1596 vdd.n2783 vdd.n722 185
R1597 vdd.n2685 vdd.n2684 185
R1598 vdd.n2684 vdd.n729 185
R1599 vdd.n2686 vdd.n727 185
R1600 vdd.n2777 vdd.n727 185
R1601 vdd.n2688 vdd.n2687 185
R1602 vdd.n2689 vdd.n2688 185
R1603 vdd.n2657 vdd.n734 185
R1604 vdd.n2771 vdd.n734 185
R1605 vdd.n2656 vdd.n2655 185
R1606 vdd.n2655 vdd.n733 185
R1607 vdd.n2654 vdd.n740 185
R1608 vdd.n2765 vdd.n740 185
R1609 vdd.n2653 vdd.n2652 185
R1610 vdd.n2652 vdd.n739 185
R1611 vdd.n2613 vdd.n745 185
R1612 vdd.n2759 vdd.n745 185
R1613 vdd.n2703 vdd.n2702 185
R1614 vdd.n2702 vdd.n2701 185
R1615 vdd.n2704 vdd.n750 185
R1616 vdd.n2753 vdd.n750 185
R1617 vdd.n2706 vdd.n2705 185
R1618 vdd.n2705 vdd.n758 185
R1619 vdd.n2707 vdd.n756 185
R1620 vdd.n2747 vdd.n756 185
R1621 vdd.n2709 vdd.n2708 185
R1622 vdd.n2708 vdd.n755 185
R1623 vdd.n2710 vdd.n762 185
R1624 vdd.n2741 vdd.n762 185
R1625 vdd.n2712 vdd.n2711 185
R1626 vdd.n2713 vdd.n2712 185
R1627 vdd.n2612 vdd.n767 185
R1628 vdd.n2735 vdd.n767 185
R1629 vdd.n2611 vdd.n2610 185
R1630 vdd.n2610 vdd.n774 185
R1631 vdd.n2609 vdd.n772 185
R1632 vdd.n2729 vdd.n772 185
R1633 vdd.n2728 vdd.n2727 185
R1634 vdd.n2729 vdd.n2728 185
R1635 vdd.n766 vdd.n765 185
R1636 vdd.n774 vdd.n766 185
R1637 vdd.n2737 vdd.n2736 185
R1638 vdd.n2736 vdd.n2735 185
R1639 vdd.n2738 vdd.n764 185
R1640 vdd.n2713 vdd.n764 185
R1641 vdd.n2740 vdd.n2739 185
R1642 vdd.n2741 vdd.n2740 185
R1643 vdd.n754 vdd.n753 185
R1644 vdd.n755 vdd.n754 185
R1645 vdd.n2749 vdd.n2748 185
R1646 vdd.n2748 vdd.n2747 185
R1647 vdd.n2750 vdd.n752 185
R1648 vdd.n758 vdd.n752 185
R1649 vdd.n2752 vdd.n2751 185
R1650 vdd.n2753 vdd.n2752 185
R1651 vdd.n744 vdd.n743 185
R1652 vdd.n2701 vdd.n744 185
R1653 vdd.n2761 vdd.n2760 185
R1654 vdd.n2760 vdd.n2759 185
R1655 vdd.n2762 vdd.n742 185
R1656 vdd.n742 vdd.n739 185
R1657 vdd.n2764 vdd.n2763 185
R1658 vdd.n2765 vdd.n2764 185
R1659 vdd.n732 vdd.n731 185
R1660 vdd.n733 vdd.n732 185
R1661 vdd.n2773 vdd.n2772 185
R1662 vdd.n2772 vdd.n2771 185
R1663 vdd.n2774 vdd.n730 185
R1664 vdd.n2689 vdd.n730 185
R1665 vdd.n2776 vdd.n2775 185
R1666 vdd.n2777 vdd.n2776 185
R1667 vdd.n721 vdd.n720 185
R1668 vdd.n729 vdd.n721 185
R1669 vdd.n2785 vdd.n2784 185
R1670 vdd.n2784 vdd.n2783 185
R1671 vdd.n2786 vdd.n719 185
R1672 vdd.n719 vdd.n716 185
R1673 vdd.n2788 vdd.n2787 185
R1674 vdd.n2789 vdd.n2788 185
R1675 vdd.n708 vdd.n707 185
R1676 vdd.n709 vdd.n708 185
R1677 vdd.n2798 vdd.n2797 185
R1678 vdd.n2797 vdd.n2796 185
R1679 vdd.n2799 vdd.n706 185
R1680 vdd.n706 vdd.n702 185
R1681 vdd.n2801 vdd.n2800 185
R1682 vdd.n2802 vdd.n2801 185
R1683 vdd.n695 vdd.n694 185
R1684 vdd.n705 vdd.n695 185
R1685 vdd.n2810 vdd.n2809 185
R1686 vdd.n2809 vdd.n2808 185
R1687 vdd.n2811 vdd.n693 185
R1688 vdd.n698 vdd.n693 185
R1689 vdd.n2813 vdd.n2812 185
R1690 vdd.n2814 vdd.n2813 185
R1691 vdd.n684 vdd.n683 185
R1692 vdd.n692 vdd.n684 185
R1693 vdd.n2822 vdd.n2821 185
R1694 vdd.n2821 vdd.n2820 185
R1695 vdd.n2823 vdd.n682 185
R1696 vdd.n682 vdd.n679 185
R1697 vdd.n2825 vdd.n2824 185
R1698 vdd.n2826 vdd.n2825 185
R1699 vdd.n670 vdd.n669 185
R1700 vdd.n671 vdd.n670 185
R1701 vdd.n2879 vdd.n2878 185
R1702 vdd.n2878 vdd.n2877 185
R1703 vdd.n2880 vdd.n668 185
R1704 vdd.n674 vdd.n668 185
R1705 vdd.n2882 vdd.n2881 185
R1706 vdd.n2883 vdd.n2882 185
R1707 vdd.n636 vdd.n634 185
R1708 vdd.n634 vdd.n631 185
R1709 vdd.n2952 vdd.n2951 185
R1710 vdd.n2953 vdd.n2952 185
R1711 vdd.n2365 vdd.n2364 185
R1712 vdd.n2366 vdd.n2365 185
R1713 vdd.n824 vdd.n822 185
R1714 vdd.n822 vdd.n820 185
R1715 vdd.n2280 vdd.n831 185
R1716 vdd.n2291 vdd.n831 185
R1717 vdd.n2281 vdd.n840 185
R1718 vdd.n2046 vdd.n840 185
R1719 vdd.n2283 vdd.n2282 185
R1720 vdd.n2284 vdd.n2283 185
R1721 vdd.n2279 vdd.n839 185
R1722 vdd.n839 vdd.n836 185
R1723 vdd.n2278 vdd.n2277 185
R1724 vdd.n2277 vdd.n2276 185
R1725 vdd.n842 vdd.n841 185
R1726 vdd.n843 vdd.n842 185
R1727 vdd.n2269 vdd.n2268 185
R1728 vdd.n2270 vdd.n2269 185
R1729 vdd.n2267 vdd.n851 185
R1730 vdd.n2058 vdd.n851 185
R1731 vdd.n2266 vdd.n2265 185
R1732 vdd.n2265 vdd.n2264 185
R1733 vdd.n853 vdd.n852 185
R1734 vdd.n861 vdd.n853 185
R1735 vdd.n2257 vdd.n2256 185
R1736 vdd.n2258 vdd.n2257 185
R1737 vdd.n2255 vdd.n862 185
R1738 vdd.n867 vdd.n862 185
R1739 vdd.n2254 vdd.n2253 185
R1740 vdd.n2253 vdd.n2252 185
R1741 vdd.n864 vdd.n863 185
R1742 vdd.n2070 vdd.n864 185
R1743 vdd.n2245 vdd.n2244 185
R1744 vdd.n2246 vdd.n2245 185
R1745 vdd.n2243 vdd.n874 185
R1746 vdd.n874 vdd.n871 185
R1747 vdd.n2242 vdd.n2241 185
R1748 vdd.n2241 vdd.n2240 185
R1749 vdd.n876 vdd.n875 185
R1750 vdd.n877 vdd.n876 185
R1751 vdd.n2233 vdd.n2232 185
R1752 vdd.n2234 vdd.n2233 185
R1753 vdd.n2230 vdd.n885 185
R1754 vdd.n891 vdd.n885 185
R1755 vdd.n2229 vdd.n2228 185
R1756 vdd.n2228 vdd.n2227 185
R1757 vdd.n888 vdd.n887 185
R1758 vdd.n898 vdd.n888 185
R1759 vdd.n2220 vdd.n2219 185
R1760 vdd.n2221 vdd.n2220 185
R1761 vdd.n2218 vdd.n899 185
R1762 vdd.n899 vdd.n895 185
R1763 vdd.n2217 vdd.n2216 185
R1764 vdd.n2216 vdd.n2215 185
R1765 vdd.n901 vdd.n900 185
R1766 vdd.n902 vdd.n901 185
R1767 vdd.n2208 vdd.n2207 185
R1768 vdd.n2209 vdd.n2208 185
R1769 vdd.n2206 vdd.n911 185
R1770 vdd.n911 vdd.n908 185
R1771 vdd.n2205 vdd.n2204 185
R1772 vdd.n2204 vdd.n2203 185
R1773 vdd.n913 vdd.n912 185
R1774 vdd.n914 vdd.n913 185
R1775 vdd.n2196 vdd.n2195 185
R1776 vdd.n2197 vdd.n2196 185
R1777 vdd.n2194 vdd.n923 185
R1778 vdd.n923 vdd.n920 185
R1779 vdd.n2193 vdd.n2192 185
R1780 vdd.n2192 vdd.n2191 185
R1781 vdd.n925 vdd.n924 185
R1782 vdd.n926 vdd.n925 185
R1783 vdd.n2184 vdd.n2183 185
R1784 vdd.n2185 vdd.n2184 185
R1785 vdd.n2182 vdd.n935 185
R1786 vdd.n935 vdd.n932 185
R1787 vdd.n2181 vdd.n2180 185
R1788 vdd.n2180 vdd.n2179 185
R1789 vdd.n2296 vdd.n795 185
R1790 vdd.n2438 vdd.n795 185
R1791 vdd.n2298 vdd.n2297 185
R1792 vdd.n2300 vdd.n2299 185
R1793 vdd.n2302 vdd.n2301 185
R1794 vdd.n2304 vdd.n2303 185
R1795 vdd.n2306 vdd.n2305 185
R1796 vdd.n2308 vdd.n2307 185
R1797 vdd.n2310 vdd.n2309 185
R1798 vdd.n2312 vdd.n2311 185
R1799 vdd.n2314 vdd.n2313 185
R1800 vdd.n2316 vdd.n2315 185
R1801 vdd.n2318 vdd.n2317 185
R1802 vdd.n2320 vdd.n2319 185
R1803 vdd.n2322 vdd.n2321 185
R1804 vdd.n2324 vdd.n2323 185
R1805 vdd.n2326 vdd.n2325 185
R1806 vdd.n2328 vdd.n2327 185
R1807 vdd.n2330 vdd.n2329 185
R1808 vdd.n2332 vdd.n2331 185
R1809 vdd.n2334 vdd.n2333 185
R1810 vdd.n2336 vdd.n2335 185
R1811 vdd.n2338 vdd.n2337 185
R1812 vdd.n2340 vdd.n2339 185
R1813 vdd.n2342 vdd.n2341 185
R1814 vdd.n2344 vdd.n2343 185
R1815 vdd.n2346 vdd.n2345 185
R1816 vdd.n2348 vdd.n2347 185
R1817 vdd.n2350 vdd.n2349 185
R1818 vdd.n2352 vdd.n2351 185
R1819 vdd.n2354 vdd.n2353 185
R1820 vdd.n2356 vdd.n2355 185
R1821 vdd.n2358 vdd.n2357 185
R1822 vdd.n2360 vdd.n2359 185
R1823 vdd.n2362 vdd.n2361 185
R1824 vdd.n2363 vdd.n823 185
R1825 vdd.n2295 vdd.n821 185
R1826 vdd.n2366 vdd.n821 185
R1827 vdd.n2294 vdd.n2293 185
R1828 vdd.n2293 vdd.n820 185
R1829 vdd.n2292 vdd.n828 185
R1830 vdd.n2292 vdd.n2291 185
R1831 vdd.n2030 vdd.n829 185
R1832 vdd.n2046 vdd.n829 185
R1833 vdd.n2031 vdd.n838 185
R1834 vdd.n2284 vdd.n838 185
R1835 vdd.n2033 vdd.n2032 185
R1836 vdd.n2032 vdd.n836 185
R1837 vdd.n2034 vdd.n845 185
R1838 vdd.n2276 vdd.n845 185
R1839 vdd.n2036 vdd.n2035 185
R1840 vdd.n2035 vdd.n843 185
R1841 vdd.n2037 vdd.n850 185
R1842 vdd.n2270 vdd.n850 185
R1843 vdd.n2060 vdd.n2059 185
R1844 vdd.n2059 vdd.n2058 185
R1845 vdd.n2061 vdd.n855 185
R1846 vdd.n2264 vdd.n855 185
R1847 vdd.n2063 vdd.n2062 185
R1848 vdd.n2062 vdd.n861 185
R1849 vdd.n2064 vdd.n860 185
R1850 vdd.n2258 vdd.n860 185
R1851 vdd.n2066 vdd.n2065 185
R1852 vdd.n2065 vdd.n867 185
R1853 vdd.n2067 vdd.n866 185
R1854 vdd.n2252 vdd.n866 185
R1855 vdd.n2069 vdd.n2068 185
R1856 vdd.n2070 vdd.n2069 185
R1857 vdd.n2029 vdd.n873 185
R1858 vdd.n2246 vdd.n873 185
R1859 vdd.n2028 vdd.n2027 185
R1860 vdd.n2027 vdd.n871 185
R1861 vdd.n2026 vdd.n879 185
R1862 vdd.n2240 vdd.n879 185
R1863 vdd.n2025 vdd.n2024 185
R1864 vdd.n2024 vdd.n877 185
R1865 vdd.n2023 vdd.n884 185
R1866 vdd.n2234 vdd.n884 185
R1867 vdd.n2022 vdd.n2021 185
R1868 vdd.n2021 vdd.n891 185
R1869 vdd.n2020 vdd.n890 185
R1870 vdd.n2227 vdd.n890 185
R1871 vdd.n2019 vdd.n2018 185
R1872 vdd.n2018 vdd.n898 185
R1873 vdd.n2017 vdd.n897 185
R1874 vdd.n2221 vdd.n897 185
R1875 vdd.n2016 vdd.n2015 185
R1876 vdd.n2015 vdd.n895 185
R1877 vdd.n2014 vdd.n904 185
R1878 vdd.n2215 vdd.n904 185
R1879 vdd.n2013 vdd.n2012 185
R1880 vdd.n2012 vdd.n902 185
R1881 vdd.n2011 vdd.n910 185
R1882 vdd.n2209 vdd.n910 185
R1883 vdd.n2010 vdd.n2009 185
R1884 vdd.n2009 vdd.n908 185
R1885 vdd.n2008 vdd.n916 185
R1886 vdd.n2203 vdd.n916 185
R1887 vdd.n2007 vdd.n2006 185
R1888 vdd.n2006 vdd.n914 185
R1889 vdd.n2005 vdd.n922 185
R1890 vdd.n2197 vdd.n922 185
R1891 vdd.n2004 vdd.n2003 185
R1892 vdd.n2003 vdd.n920 185
R1893 vdd.n2002 vdd.n928 185
R1894 vdd.n2191 vdd.n928 185
R1895 vdd.n2001 vdd.n2000 185
R1896 vdd.n2000 vdd.n926 185
R1897 vdd.n1999 vdd.n934 185
R1898 vdd.n2185 vdd.n934 185
R1899 vdd.n1998 vdd.n1997 185
R1900 vdd.n1997 vdd.n932 185
R1901 vdd.n1996 vdd.n940 185
R1902 vdd.n2179 vdd.n940 185
R1903 vdd.n937 vdd.n936 185
R1904 vdd.n1928 vdd.n1926 185
R1905 vdd.n1931 vdd.n1930 185
R1906 vdd.n1932 vdd.n1925 185
R1907 vdd.n1934 vdd.n1933 185
R1908 vdd.n1936 vdd.n1924 185
R1909 vdd.n1939 vdd.n1938 185
R1910 vdd.n1940 vdd.n1923 185
R1911 vdd.n1942 vdd.n1941 185
R1912 vdd.n1944 vdd.n1922 185
R1913 vdd.n1947 vdd.n1946 185
R1914 vdd.n1948 vdd.n1921 185
R1915 vdd.n1950 vdd.n1949 185
R1916 vdd.n1952 vdd.n1920 185
R1917 vdd.n1955 vdd.n1954 185
R1918 vdd.n1956 vdd.n1919 185
R1919 vdd.n1958 vdd.n1957 185
R1920 vdd.n1960 vdd.n1918 185
R1921 vdd.n1963 vdd.n1962 185
R1922 vdd.n1964 vdd.n971 185
R1923 vdd.n1966 vdd.n1965 185
R1924 vdd.n1968 vdd.n970 185
R1925 vdd.n1971 vdd.n1970 185
R1926 vdd.n1972 vdd.n969 185
R1927 vdd.n1974 vdd.n1973 185
R1928 vdd.n1976 vdd.n968 185
R1929 vdd.n1979 vdd.n1978 185
R1930 vdd.n1980 vdd.n967 185
R1931 vdd.n1982 vdd.n1981 185
R1932 vdd.n1984 vdd.n966 185
R1933 vdd.n1987 vdd.n1986 185
R1934 vdd.n1988 vdd.n963 185
R1935 vdd.n1991 vdd.n1990 185
R1936 vdd.n1993 vdd.n962 185
R1937 vdd.n1995 vdd.n1994 185
R1938 vdd.n1994 vdd.n938 185
R1939 vdd.n303 vdd.n302 171.744
R1940 vdd.n302 vdd.n301 171.744
R1941 vdd.n301 vdd.n270 171.744
R1942 vdd.n294 vdd.n270 171.744
R1943 vdd.n294 vdd.n293 171.744
R1944 vdd.n293 vdd.n275 171.744
R1945 vdd.n286 vdd.n275 171.744
R1946 vdd.n286 vdd.n285 171.744
R1947 vdd.n285 vdd.n279 171.744
R1948 vdd.n252 vdd.n251 171.744
R1949 vdd.n251 vdd.n250 171.744
R1950 vdd.n250 vdd.n219 171.744
R1951 vdd.n243 vdd.n219 171.744
R1952 vdd.n243 vdd.n242 171.744
R1953 vdd.n242 vdd.n224 171.744
R1954 vdd.n235 vdd.n224 171.744
R1955 vdd.n235 vdd.n234 171.744
R1956 vdd.n234 vdd.n228 171.744
R1957 vdd.n209 vdd.n208 171.744
R1958 vdd.n208 vdd.n207 171.744
R1959 vdd.n207 vdd.n176 171.744
R1960 vdd.n200 vdd.n176 171.744
R1961 vdd.n200 vdd.n199 171.744
R1962 vdd.n199 vdd.n181 171.744
R1963 vdd.n192 vdd.n181 171.744
R1964 vdd.n192 vdd.n191 171.744
R1965 vdd.n191 vdd.n185 171.744
R1966 vdd.n158 vdd.n157 171.744
R1967 vdd.n157 vdd.n156 171.744
R1968 vdd.n156 vdd.n125 171.744
R1969 vdd.n149 vdd.n125 171.744
R1970 vdd.n149 vdd.n148 171.744
R1971 vdd.n148 vdd.n130 171.744
R1972 vdd.n141 vdd.n130 171.744
R1973 vdd.n141 vdd.n140 171.744
R1974 vdd.n140 vdd.n134 171.744
R1975 vdd.n116 vdd.n115 171.744
R1976 vdd.n115 vdd.n114 171.744
R1977 vdd.n114 vdd.n83 171.744
R1978 vdd.n107 vdd.n83 171.744
R1979 vdd.n107 vdd.n106 171.744
R1980 vdd.n106 vdd.n88 171.744
R1981 vdd.n99 vdd.n88 171.744
R1982 vdd.n99 vdd.n98 171.744
R1983 vdd.n98 vdd.n92 171.744
R1984 vdd.n65 vdd.n64 171.744
R1985 vdd.n64 vdd.n63 171.744
R1986 vdd.n63 vdd.n32 171.744
R1987 vdd.n56 vdd.n32 171.744
R1988 vdd.n56 vdd.n55 171.744
R1989 vdd.n55 vdd.n37 171.744
R1990 vdd.n48 vdd.n37 171.744
R1991 vdd.n48 vdd.n47 171.744
R1992 vdd.n47 vdd.n41 171.744
R1993 vdd.n1578 vdd.n1577 171.744
R1994 vdd.n1577 vdd.n1576 171.744
R1995 vdd.n1576 vdd.n1545 171.744
R1996 vdd.n1569 vdd.n1545 171.744
R1997 vdd.n1569 vdd.n1568 171.744
R1998 vdd.n1568 vdd.n1550 171.744
R1999 vdd.n1561 vdd.n1550 171.744
R2000 vdd.n1561 vdd.n1560 171.744
R2001 vdd.n1560 vdd.n1554 171.744
R2002 vdd.n1629 vdd.n1628 171.744
R2003 vdd.n1628 vdd.n1627 171.744
R2004 vdd.n1627 vdd.n1596 171.744
R2005 vdd.n1620 vdd.n1596 171.744
R2006 vdd.n1620 vdd.n1619 171.744
R2007 vdd.n1619 vdd.n1601 171.744
R2008 vdd.n1612 vdd.n1601 171.744
R2009 vdd.n1612 vdd.n1611 171.744
R2010 vdd.n1611 vdd.n1605 171.744
R2011 vdd.n1484 vdd.n1483 171.744
R2012 vdd.n1483 vdd.n1482 171.744
R2013 vdd.n1482 vdd.n1451 171.744
R2014 vdd.n1475 vdd.n1451 171.744
R2015 vdd.n1475 vdd.n1474 171.744
R2016 vdd.n1474 vdd.n1456 171.744
R2017 vdd.n1467 vdd.n1456 171.744
R2018 vdd.n1467 vdd.n1466 171.744
R2019 vdd.n1466 vdd.n1460 171.744
R2020 vdd.n1535 vdd.n1534 171.744
R2021 vdd.n1534 vdd.n1533 171.744
R2022 vdd.n1533 vdd.n1502 171.744
R2023 vdd.n1526 vdd.n1502 171.744
R2024 vdd.n1526 vdd.n1525 171.744
R2025 vdd.n1525 vdd.n1507 171.744
R2026 vdd.n1518 vdd.n1507 171.744
R2027 vdd.n1518 vdd.n1517 171.744
R2028 vdd.n1517 vdd.n1511 171.744
R2029 vdd.n1391 vdd.n1390 171.744
R2030 vdd.n1390 vdd.n1389 171.744
R2031 vdd.n1389 vdd.n1358 171.744
R2032 vdd.n1382 vdd.n1358 171.744
R2033 vdd.n1382 vdd.n1381 171.744
R2034 vdd.n1381 vdd.n1363 171.744
R2035 vdd.n1374 vdd.n1363 171.744
R2036 vdd.n1374 vdd.n1373 171.744
R2037 vdd.n1373 vdd.n1367 171.744
R2038 vdd.n1442 vdd.n1441 171.744
R2039 vdd.n1441 vdd.n1440 171.744
R2040 vdd.n1440 vdd.n1409 171.744
R2041 vdd.n1433 vdd.n1409 171.744
R2042 vdd.n1433 vdd.n1432 171.744
R2043 vdd.n1432 vdd.n1414 171.744
R2044 vdd.n1425 vdd.n1414 171.744
R2045 vdd.n1425 vdd.n1424 171.744
R2046 vdd.n1424 vdd.n1418 171.744
R2047 vdd.n3312 vdd.n356 146.341
R2048 vdd.n3310 vdd.n3309 146.341
R2049 vdd.n3307 vdd.n360 146.341
R2050 vdd.n3303 vdd.n3302 146.341
R2051 vdd.n3300 vdd.n368 146.341
R2052 vdd.n3296 vdd.n3295 146.341
R2053 vdd.n3293 vdd.n375 146.341
R2054 vdd.n3289 vdd.n3288 146.341
R2055 vdd.n3286 vdd.n382 146.341
R2056 vdd.n393 vdd.n390 146.341
R2057 vdd.n3278 vdd.n3277 146.341
R2058 vdd.n3275 vdd.n395 146.341
R2059 vdd.n3271 vdd.n3270 146.341
R2060 vdd.n3268 vdd.n401 146.341
R2061 vdd.n3264 vdd.n3263 146.341
R2062 vdd.n3261 vdd.n408 146.341
R2063 vdd.n3257 vdd.n3256 146.341
R2064 vdd.n3254 vdd.n415 146.341
R2065 vdd.n3250 vdd.n3249 146.341
R2066 vdd.n3247 vdd.n422 146.341
R2067 vdd.n433 vdd.n430 146.341
R2068 vdd.n3239 vdd.n3238 146.341
R2069 vdd.n3236 vdd.n435 146.341
R2070 vdd.n3232 vdd.n3231 146.341
R2071 vdd.n3229 vdd.n441 146.341
R2072 vdd.n3225 vdd.n3224 146.341
R2073 vdd.n3222 vdd.n448 146.341
R2074 vdd.n3218 vdd.n3217 146.341
R2075 vdd.n3215 vdd.n455 146.341
R2076 vdd.n3211 vdd.n3210 146.341
R2077 vdd.n3208 vdd.n462 146.341
R2078 vdd.n3123 vdd.n512 146.341
R2079 vdd.n3129 vdd.n512 146.341
R2080 vdd.n3129 vdd.n504 146.341
R2081 vdd.n3139 vdd.n504 146.341
R2082 vdd.n3139 vdd.n500 146.341
R2083 vdd.n3145 vdd.n500 146.341
R2084 vdd.n3145 vdd.n491 146.341
R2085 vdd.n3155 vdd.n491 146.341
R2086 vdd.n3155 vdd.n487 146.341
R2087 vdd.n3161 vdd.n487 146.341
R2088 vdd.n3161 vdd.n479 146.341
R2089 vdd.n3172 vdd.n479 146.341
R2090 vdd.n3172 vdd.n480 146.341
R2091 vdd.n480 vdd.n316 146.341
R2092 vdd.n317 vdd.n316 146.341
R2093 vdd.n318 vdd.n317 146.341
R2094 vdd.n473 vdd.n318 146.341
R2095 vdd.n473 vdd.n326 146.341
R2096 vdd.n327 vdd.n326 146.341
R2097 vdd.n328 vdd.n327 146.341
R2098 vdd.n470 vdd.n328 146.341
R2099 vdd.n470 vdd.n337 146.341
R2100 vdd.n338 vdd.n337 146.341
R2101 vdd.n339 vdd.n338 146.341
R2102 vdd.n467 vdd.n339 146.341
R2103 vdd.n467 vdd.n348 146.341
R2104 vdd.n349 vdd.n348 146.341
R2105 vdd.n350 vdd.n349 146.341
R2106 vdd.n3115 vdd.n3113 146.341
R2107 vdd.n3113 vdd.n3112 146.341
R2108 vdd.n3109 vdd.n3108 146.341
R2109 vdd.n3105 vdd.n3104 146.341
R2110 vdd.n3102 vdd.n526 146.341
R2111 vdd.n3098 vdd.n3096 146.341
R2112 vdd.n3094 vdd.n532 146.341
R2113 vdd.n3090 vdd.n3088 146.341
R2114 vdd.n3086 vdd.n538 146.341
R2115 vdd.n3082 vdd.n3080 146.341
R2116 vdd.n3078 vdd.n546 146.341
R2117 vdd.n3074 vdd.n3072 146.341
R2118 vdd.n3070 vdd.n552 146.341
R2119 vdd.n3066 vdd.n3064 146.341
R2120 vdd.n3062 vdd.n558 146.341
R2121 vdd.n3058 vdd.n3056 146.341
R2122 vdd.n3054 vdd.n564 146.341
R2123 vdd.n3050 vdd.n3048 146.341
R2124 vdd.n3046 vdd.n570 146.341
R2125 vdd.n3042 vdd.n3040 146.341
R2126 vdd.n3038 vdd.n576 146.341
R2127 vdd.n3031 vdd.n585 146.341
R2128 vdd.n3029 vdd.n3028 146.341
R2129 vdd.n3025 vdd.n3024 146.341
R2130 vdd.n3022 vdd.n590 146.341
R2131 vdd.n3018 vdd.n3016 146.341
R2132 vdd.n3014 vdd.n596 146.341
R2133 vdd.n3010 vdd.n3008 146.341
R2134 vdd.n3006 vdd.n602 146.341
R2135 vdd.n3002 vdd.n3000 146.341
R2136 vdd.n2997 vdd.n2996 146.341
R2137 vdd.n2993 vdd.n515 146.341
R2138 vdd.n3121 vdd.n510 146.341
R2139 vdd.n3131 vdd.n510 146.341
R2140 vdd.n3131 vdd.n506 146.341
R2141 vdd.n3137 vdd.n506 146.341
R2142 vdd.n3137 vdd.n498 146.341
R2143 vdd.n3147 vdd.n498 146.341
R2144 vdd.n3147 vdd.n494 146.341
R2145 vdd.n3153 vdd.n494 146.341
R2146 vdd.n3153 vdd.n486 146.341
R2147 vdd.n3164 vdd.n486 146.341
R2148 vdd.n3164 vdd.n482 146.341
R2149 vdd.n3170 vdd.n482 146.341
R2150 vdd.n3170 vdd.n314 146.341
R2151 vdd.n3347 vdd.n314 146.341
R2152 vdd.n3347 vdd.n315 146.341
R2153 vdd.n3343 vdd.n315 146.341
R2154 vdd.n3343 vdd.n319 146.341
R2155 vdd.n3339 vdd.n319 146.341
R2156 vdd.n3339 vdd.n324 146.341
R2157 vdd.n3335 vdd.n324 146.341
R2158 vdd.n3335 vdd.n330 146.341
R2159 vdd.n3331 vdd.n330 146.341
R2160 vdd.n3331 vdd.n336 146.341
R2161 vdd.n3327 vdd.n336 146.341
R2162 vdd.n3327 vdd.n341 146.341
R2163 vdd.n3323 vdd.n341 146.341
R2164 vdd.n3323 vdd.n347 146.341
R2165 vdd.n3319 vdd.n347 146.341
R2166 vdd.n1901 vdd.n1900 146.341
R2167 vdd.n1898 vdd.n1695 146.341
R2168 vdd.n1891 vdd.n1701 146.341
R2169 vdd.n1889 vdd.n1888 146.341
R2170 vdd.n1886 vdd.n1703 146.341
R2171 vdd.n1882 vdd.n1881 146.341
R2172 vdd.n1879 vdd.n1710 146.341
R2173 vdd.n1875 vdd.n1874 146.341
R2174 vdd.n1872 vdd.n1717 146.341
R2175 vdd.n1728 vdd.n1725 146.341
R2176 vdd.n1864 vdd.n1863 146.341
R2177 vdd.n1861 vdd.n1730 146.341
R2178 vdd.n1857 vdd.n1856 146.341
R2179 vdd.n1854 vdd.n1736 146.341
R2180 vdd.n1850 vdd.n1849 146.341
R2181 vdd.n1847 vdd.n1743 146.341
R2182 vdd.n1843 vdd.n1842 146.341
R2183 vdd.n1840 vdd.n1750 146.341
R2184 vdd.n1836 vdd.n1835 146.341
R2185 vdd.n1833 vdd.n1757 146.341
R2186 vdd.n1768 vdd.n1765 146.341
R2187 vdd.n1825 vdd.n1824 146.341
R2188 vdd.n1822 vdd.n1770 146.341
R2189 vdd.n1818 vdd.n1817 146.341
R2190 vdd.n1815 vdd.n1776 146.341
R2191 vdd.n1811 vdd.n1810 146.341
R2192 vdd.n1808 vdd.n1783 146.341
R2193 vdd.n1804 vdd.n1803 146.341
R2194 vdd.n1801 vdd.n1798 146.341
R2195 vdd.n1796 vdd.n1793 146.341
R2196 vdd.n1791 vdd.n977 146.341
R2197 vdd.n1296 vdd.n1058 146.341
R2198 vdd.n1302 vdd.n1058 146.341
R2199 vdd.n1302 vdd.n1051 146.341
R2200 vdd.n1312 vdd.n1051 146.341
R2201 vdd.n1312 vdd.n1047 146.341
R2202 vdd.n1318 vdd.n1047 146.341
R2203 vdd.n1318 vdd.n1038 146.341
R2204 vdd.n1328 vdd.n1038 146.341
R2205 vdd.n1328 vdd.n1034 146.341
R2206 vdd.n1334 vdd.n1034 146.341
R2207 vdd.n1334 vdd.n1027 146.341
R2208 vdd.n1345 vdd.n1027 146.341
R2209 vdd.n1345 vdd.n1023 146.341
R2210 vdd.n1351 vdd.n1023 146.341
R2211 vdd.n1351 vdd.n1016 146.341
R2212 vdd.n1643 vdd.n1016 146.341
R2213 vdd.n1643 vdd.n1012 146.341
R2214 vdd.n1649 vdd.n1012 146.341
R2215 vdd.n1649 vdd.n1004 146.341
R2216 vdd.n1660 vdd.n1004 146.341
R2217 vdd.n1660 vdd.n1000 146.341
R2218 vdd.n1666 vdd.n1000 146.341
R2219 vdd.n1666 vdd.n994 146.341
R2220 vdd.n1677 vdd.n994 146.341
R2221 vdd.n1677 vdd.n989 146.341
R2222 vdd.n1685 vdd.n989 146.341
R2223 vdd.n1685 vdd.n979 146.341
R2224 vdd.n1909 vdd.n979 146.341
R2225 vdd.n1068 vdd.n1067 146.341
R2226 vdd.n1071 vdd.n1068 146.341
R2227 vdd.n1074 vdd.n1073 146.341
R2228 vdd.n1079 vdd.n1076 146.341
R2229 vdd.n1082 vdd.n1081 146.341
R2230 vdd.n1087 vdd.n1084 146.341
R2231 vdd.n1090 vdd.n1089 146.341
R2232 vdd.n1095 vdd.n1092 146.341
R2233 vdd.n1098 vdd.n1097 146.341
R2234 vdd.n1105 vdd.n1100 146.341
R2235 vdd.n1108 vdd.n1107 146.341
R2236 vdd.n1113 vdd.n1110 146.341
R2237 vdd.n1116 vdd.n1115 146.341
R2238 vdd.n1121 vdd.n1118 146.341
R2239 vdd.n1124 vdd.n1123 146.341
R2240 vdd.n1129 vdd.n1126 146.341
R2241 vdd.n1132 vdd.n1131 146.341
R2242 vdd.n1137 vdd.n1134 146.341
R2243 vdd.n1140 vdd.n1139 146.341
R2244 vdd.n1145 vdd.n1142 146.341
R2245 vdd.n1226 vdd.n1147 146.341
R2246 vdd.n1224 vdd.n1223 146.341
R2247 vdd.n1154 vdd.n1153 146.341
R2248 vdd.n1157 vdd.n1156 146.341
R2249 vdd.n1162 vdd.n1161 146.341
R2250 vdd.n1165 vdd.n1164 146.341
R2251 vdd.n1170 vdd.n1169 146.341
R2252 vdd.n1173 vdd.n1172 146.341
R2253 vdd.n1178 vdd.n1177 146.341
R2254 vdd.n1181 vdd.n1180 146.341
R2255 vdd.n1186 vdd.n1185 146.341
R2256 vdd.n1188 vdd.n1061 146.341
R2257 vdd.n1294 vdd.n1057 146.341
R2258 vdd.n1304 vdd.n1057 146.341
R2259 vdd.n1304 vdd.n1053 146.341
R2260 vdd.n1310 vdd.n1053 146.341
R2261 vdd.n1310 vdd.n1045 146.341
R2262 vdd.n1320 vdd.n1045 146.341
R2263 vdd.n1320 vdd.n1041 146.341
R2264 vdd.n1326 vdd.n1041 146.341
R2265 vdd.n1326 vdd.n1033 146.341
R2266 vdd.n1337 vdd.n1033 146.341
R2267 vdd.n1337 vdd.n1029 146.341
R2268 vdd.n1343 vdd.n1029 146.341
R2269 vdd.n1343 vdd.n1022 146.341
R2270 vdd.n1353 vdd.n1022 146.341
R2271 vdd.n1353 vdd.n1018 146.341
R2272 vdd.n1641 vdd.n1018 146.341
R2273 vdd.n1641 vdd.n1010 146.341
R2274 vdd.n1652 vdd.n1010 146.341
R2275 vdd.n1652 vdd.n1006 146.341
R2276 vdd.n1658 vdd.n1006 146.341
R2277 vdd.n1658 vdd.n999 146.341
R2278 vdd.n1669 vdd.n999 146.341
R2279 vdd.n1669 vdd.n995 146.341
R2280 vdd.n1675 vdd.n995 146.341
R2281 vdd.n1675 vdd.n987 146.341
R2282 vdd.n1688 vdd.n987 146.341
R2283 vdd.n1688 vdd.n982 146.341
R2284 vdd.n1907 vdd.n982 146.341
R2285 vdd.n964 vdd.t105 127.284
R2286 vdd.n825 vdd.t142 127.284
R2287 vdd.n958 vdd.t166 127.284
R2288 vdd.n816 vdd.t159 127.284
R2289 vdd.n713 vdd.t111 127.284
R2290 vdd.n713 vdd.t112 127.284
R2291 vdd.n2473 vdd.t157 127.284
R2292 vdd.n661 vdd.t135 127.284
R2293 vdd.n2542 vdd.t147 127.284
R2294 vdd.n625 vdd.t100 127.284
R2295 vdd.n886 vdd.t153 127.284
R2296 vdd.n886 vdd.t154 127.284
R2297 vdd.n22 vdd.n20 117.314
R2298 vdd.n17 vdd.n15 117.314
R2299 vdd.n27 vdd.n26 116.927
R2300 vdd.n24 vdd.n23 116.927
R2301 vdd.n22 vdd.n21 116.927
R2302 vdd.n17 vdd.n16 116.927
R2303 vdd.n19 vdd.n18 116.927
R2304 vdd.n27 vdd.n25 116.927
R2305 vdd.n965 vdd.t104 111.188
R2306 vdd.n826 vdd.t143 111.188
R2307 vdd.n959 vdd.t165 111.188
R2308 vdd.n817 vdd.t160 111.188
R2309 vdd.n2474 vdd.t156 111.188
R2310 vdd.n662 vdd.t136 111.188
R2311 vdd.n2543 vdd.t146 111.188
R2312 vdd.n626 vdd.t101 111.188
R2313 vdd.n2728 vdd.n766 99.5127
R2314 vdd.n2736 vdd.n766 99.5127
R2315 vdd.n2736 vdd.n764 99.5127
R2316 vdd.n2740 vdd.n764 99.5127
R2317 vdd.n2740 vdd.n754 99.5127
R2318 vdd.n2748 vdd.n754 99.5127
R2319 vdd.n2748 vdd.n752 99.5127
R2320 vdd.n2752 vdd.n752 99.5127
R2321 vdd.n2752 vdd.n744 99.5127
R2322 vdd.n2760 vdd.n744 99.5127
R2323 vdd.n2760 vdd.n742 99.5127
R2324 vdd.n2764 vdd.n742 99.5127
R2325 vdd.n2764 vdd.n732 99.5127
R2326 vdd.n2772 vdd.n732 99.5127
R2327 vdd.n2772 vdd.n730 99.5127
R2328 vdd.n2776 vdd.n730 99.5127
R2329 vdd.n2776 vdd.n721 99.5127
R2330 vdd.n2784 vdd.n721 99.5127
R2331 vdd.n2784 vdd.n719 99.5127
R2332 vdd.n2788 vdd.n719 99.5127
R2333 vdd.n2788 vdd.n708 99.5127
R2334 vdd.n2797 vdd.n708 99.5127
R2335 vdd.n2797 vdd.n706 99.5127
R2336 vdd.n2801 vdd.n706 99.5127
R2337 vdd.n2801 vdd.n695 99.5127
R2338 vdd.n2809 vdd.n695 99.5127
R2339 vdd.n2809 vdd.n693 99.5127
R2340 vdd.n2813 vdd.n693 99.5127
R2341 vdd.n2813 vdd.n684 99.5127
R2342 vdd.n2821 vdd.n684 99.5127
R2343 vdd.n2821 vdd.n682 99.5127
R2344 vdd.n2825 vdd.n682 99.5127
R2345 vdd.n2825 vdd.n670 99.5127
R2346 vdd.n2878 vdd.n670 99.5127
R2347 vdd.n2878 vdd.n668 99.5127
R2348 vdd.n2882 vdd.n668 99.5127
R2349 vdd.n2882 vdd.n634 99.5127
R2350 vdd.n2952 vdd.n634 99.5127
R2351 vdd.n2948 vdd.n635 99.5127
R2352 vdd.n2946 vdd.n2945 99.5127
R2353 vdd.n2943 vdd.n639 99.5127
R2354 vdd.n2939 vdd.n2938 99.5127
R2355 vdd.n2936 vdd.n642 99.5127
R2356 vdd.n2932 vdd.n2931 99.5127
R2357 vdd.n2929 vdd.n645 99.5127
R2358 vdd.n2925 vdd.n2924 99.5127
R2359 vdd.n2922 vdd.n648 99.5127
R2360 vdd.n2917 vdd.n2916 99.5127
R2361 vdd.n2914 vdd.n651 99.5127
R2362 vdd.n2910 vdd.n2909 99.5127
R2363 vdd.n2907 vdd.n654 99.5127
R2364 vdd.n2903 vdd.n2902 99.5127
R2365 vdd.n2900 vdd.n657 99.5127
R2366 vdd.n2896 vdd.n2895 99.5127
R2367 vdd.n2893 vdd.n660 99.5127
R2368 vdd.n2610 vdd.n772 99.5127
R2369 vdd.n2610 vdd.n767 99.5127
R2370 vdd.n2712 vdd.n767 99.5127
R2371 vdd.n2712 vdd.n762 99.5127
R2372 vdd.n2708 vdd.n762 99.5127
R2373 vdd.n2708 vdd.n756 99.5127
R2374 vdd.n2705 vdd.n756 99.5127
R2375 vdd.n2705 vdd.n750 99.5127
R2376 vdd.n2702 vdd.n750 99.5127
R2377 vdd.n2702 vdd.n745 99.5127
R2378 vdd.n2652 vdd.n745 99.5127
R2379 vdd.n2652 vdd.n740 99.5127
R2380 vdd.n2655 vdd.n740 99.5127
R2381 vdd.n2655 vdd.n734 99.5127
R2382 vdd.n2688 vdd.n734 99.5127
R2383 vdd.n2688 vdd.n727 99.5127
R2384 vdd.n2684 vdd.n727 99.5127
R2385 vdd.n2684 vdd.n722 99.5127
R2386 vdd.n2681 vdd.n722 99.5127
R2387 vdd.n2681 vdd.n717 99.5127
R2388 vdd.n2678 vdd.n717 99.5127
R2389 vdd.n2678 vdd.n710 99.5127
R2390 vdd.n2675 vdd.n710 99.5127
R2391 vdd.n2675 vdd.n703 99.5127
R2392 vdd.n2672 vdd.n703 99.5127
R2393 vdd.n2672 vdd.n696 99.5127
R2394 vdd.n2669 vdd.n696 99.5127
R2395 vdd.n2669 vdd.n690 99.5127
R2396 vdd.n2666 vdd.n690 99.5127
R2397 vdd.n2666 vdd.n685 99.5127
R2398 vdd.n2663 vdd.n685 99.5127
R2399 vdd.n2663 vdd.n680 99.5127
R2400 vdd.n2660 vdd.n680 99.5127
R2401 vdd.n2660 vdd.n672 99.5127
R2402 vdd.n672 vdd.n665 99.5127
R2403 vdd.n2884 vdd.n665 99.5127
R2404 vdd.n2885 vdd.n2884 99.5127
R2405 vdd.n2885 vdd.n632 99.5127
R2406 vdd.n2724 vdd.n777 99.5127
R2407 vdd.n2544 vdd.n777 99.5127
R2408 vdd.n2548 vdd.n2547 99.5127
R2409 vdd.n2552 vdd.n2551 99.5127
R2410 vdd.n2556 vdd.n2555 99.5127
R2411 vdd.n2560 vdd.n2559 99.5127
R2412 vdd.n2564 vdd.n2563 99.5127
R2413 vdd.n2568 vdd.n2567 99.5127
R2414 vdd.n2572 vdd.n2571 99.5127
R2415 vdd.n2576 vdd.n2575 99.5127
R2416 vdd.n2580 vdd.n2579 99.5127
R2417 vdd.n2584 vdd.n2583 99.5127
R2418 vdd.n2588 vdd.n2587 99.5127
R2419 vdd.n2592 vdd.n2591 99.5127
R2420 vdd.n2596 vdd.n2595 99.5127
R2421 vdd.n2600 vdd.n2599 99.5127
R2422 vdd.n2605 vdd.n2604 99.5127
R2423 vdd.n2437 vdd.n814 99.5127
R2424 vdd.n2433 vdd.n2432 99.5127
R2425 vdd.n2429 vdd.n2428 99.5127
R2426 vdd.n2425 vdd.n2424 99.5127
R2427 vdd.n2421 vdd.n2420 99.5127
R2428 vdd.n2417 vdd.n2416 99.5127
R2429 vdd.n2413 vdd.n2412 99.5127
R2430 vdd.n2409 vdd.n2408 99.5127
R2431 vdd.n2405 vdd.n2404 99.5127
R2432 vdd.n2401 vdd.n2400 99.5127
R2433 vdd.n2397 vdd.n2396 99.5127
R2434 vdd.n2393 vdd.n2392 99.5127
R2435 vdd.n2389 vdd.n2388 99.5127
R2436 vdd.n2385 vdd.n2384 99.5127
R2437 vdd.n2381 vdd.n2380 99.5127
R2438 vdd.n2377 vdd.n2376 99.5127
R2439 vdd.n2372 vdd.n2371 99.5127
R2440 vdd.n2104 vdd.n939 99.5127
R2441 vdd.n2104 vdd.n933 99.5127
R2442 vdd.n2101 vdd.n933 99.5127
R2443 vdd.n2101 vdd.n927 99.5127
R2444 vdd.n2098 vdd.n927 99.5127
R2445 vdd.n2098 vdd.n921 99.5127
R2446 vdd.n2095 vdd.n921 99.5127
R2447 vdd.n2095 vdd.n915 99.5127
R2448 vdd.n2092 vdd.n915 99.5127
R2449 vdd.n2092 vdd.n909 99.5127
R2450 vdd.n2089 vdd.n909 99.5127
R2451 vdd.n2089 vdd.n903 99.5127
R2452 vdd.n2086 vdd.n903 99.5127
R2453 vdd.n2086 vdd.n896 99.5127
R2454 vdd.n2083 vdd.n896 99.5127
R2455 vdd.n2083 vdd.n889 99.5127
R2456 vdd.n2080 vdd.n889 99.5127
R2457 vdd.n2080 vdd.n883 99.5127
R2458 vdd.n2077 vdd.n883 99.5127
R2459 vdd.n2077 vdd.n878 99.5127
R2460 vdd.n2074 vdd.n878 99.5127
R2461 vdd.n2074 vdd.n872 99.5127
R2462 vdd.n2071 vdd.n872 99.5127
R2463 vdd.n2071 vdd.n865 99.5127
R2464 vdd.n2038 vdd.n865 99.5127
R2465 vdd.n2038 vdd.n859 99.5127
R2466 vdd.n2041 vdd.n859 99.5127
R2467 vdd.n2041 vdd.n854 99.5127
R2468 vdd.n2057 vdd.n854 99.5127
R2469 vdd.n2057 vdd.n849 99.5127
R2470 vdd.n2053 vdd.n849 99.5127
R2471 vdd.n2053 vdd.n844 99.5127
R2472 vdd.n2050 vdd.n844 99.5127
R2473 vdd.n2050 vdd.n837 99.5127
R2474 vdd.n2047 vdd.n837 99.5127
R2475 vdd.n2047 vdd.n830 99.5127
R2476 vdd.n830 vdd.n819 99.5127
R2477 vdd.n2367 vdd.n819 99.5127
R2478 vdd.n2174 vdd.n2172 99.5127
R2479 vdd.n2172 vdd.n2171 99.5127
R2480 vdd.n2168 vdd.n2167 99.5127
R2481 vdd.n2165 vdd.n945 99.5127
R2482 vdd.n2161 vdd.n2159 99.5127
R2483 vdd.n2157 vdd.n947 99.5127
R2484 vdd.n2153 vdd.n2151 99.5127
R2485 vdd.n2149 vdd.n949 99.5127
R2486 vdd.n2145 vdd.n2143 99.5127
R2487 vdd.n2141 vdd.n951 99.5127
R2488 vdd.n2137 vdd.n2135 99.5127
R2489 vdd.n2133 vdd.n953 99.5127
R2490 vdd.n2129 vdd.n2127 99.5127
R2491 vdd.n2125 vdd.n955 99.5127
R2492 vdd.n2121 vdd.n2119 99.5127
R2493 vdd.n2117 vdd.n957 99.5127
R2494 vdd.n2112 vdd.n2110 99.5127
R2495 vdd.n2178 vdd.n931 99.5127
R2496 vdd.n2186 vdd.n931 99.5127
R2497 vdd.n2186 vdd.n929 99.5127
R2498 vdd.n2190 vdd.n929 99.5127
R2499 vdd.n2190 vdd.n919 99.5127
R2500 vdd.n2198 vdd.n919 99.5127
R2501 vdd.n2198 vdd.n917 99.5127
R2502 vdd.n2202 vdd.n917 99.5127
R2503 vdd.n2202 vdd.n907 99.5127
R2504 vdd.n2210 vdd.n907 99.5127
R2505 vdd.n2210 vdd.n905 99.5127
R2506 vdd.n2214 vdd.n905 99.5127
R2507 vdd.n2214 vdd.n894 99.5127
R2508 vdd.n2222 vdd.n894 99.5127
R2509 vdd.n2222 vdd.n892 99.5127
R2510 vdd.n2226 vdd.n892 99.5127
R2511 vdd.n2226 vdd.n882 99.5127
R2512 vdd.n2235 vdd.n882 99.5127
R2513 vdd.n2235 vdd.n880 99.5127
R2514 vdd.n2239 vdd.n880 99.5127
R2515 vdd.n2239 vdd.n870 99.5127
R2516 vdd.n2247 vdd.n870 99.5127
R2517 vdd.n2247 vdd.n868 99.5127
R2518 vdd.n2251 vdd.n868 99.5127
R2519 vdd.n2251 vdd.n858 99.5127
R2520 vdd.n2259 vdd.n858 99.5127
R2521 vdd.n2259 vdd.n856 99.5127
R2522 vdd.n2263 vdd.n856 99.5127
R2523 vdd.n2263 vdd.n848 99.5127
R2524 vdd.n2271 vdd.n848 99.5127
R2525 vdd.n2271 vdd.n846 99.5127
R2526 vdd.n2275 vdd.n846 99.5127
R2527 vdd.n2275 vdd.n835 99.5127
R2528 vdd.n2285 vdd.n835 99.5127
R2529 vdd.n2285 vdd.n832 99.5127
R2530 vdd.n2290 vdd.n832 99.5127
R2531 vdd.n2290 vdd.n833 99.5127
R2532 vdd.n833 vdd.n813 99.5127
R2533 vdd.n2868 vdd.n2867 99.5127
R2534 vdd.n2865 vdd.n2831 99.5127
R2535 vdd.n2861 vdd.n2860 99.5127
R2536 vdd.n2858 vdd.n2834 99.5127
R2537 vdd.n2854 vdd.n2853 99.5127
R2538 vdd.n2851 vdd.n2837 99.5127
R2539 vdd.n2847 vdd.n2846 99.5127
R2540 vdd.n2844 vdd.n2841 99.5127
R2541 vdd.n2985 vdd.n612 99.5127
R2542 vdd.n2983 vdd.n2982 99.5127
R2543 vdd.n2980 vdd.n615 99.5127
R2544 vdd.n2976 vdd.n2975 99.5127
R2545 vdd.n2973 vdd.n618 99.5127
R2546 vdd.n2969 vdd.n2968 99.5127
R2547 vdd.n2966 vdd.n621 99.5127
R2548 vdd.n2962 vdd.n2961 99.5127
R2549 vdd.n2959 vdd.n624 99.5127
R2550 vdd.n2717 vdd.n773 99.5127
R2551 vdd.n2717 vdd.n768 99.5127
R2552 vdd.n2714 vdd.n768 99.5127
R2553 vdd.n2714 vdd.n763 99.5127
R2554 vdd.n2614 vdd.n763 99.5127
R2555 vdd.n2614 vdd.n757 99.5127
R2556 vdd.n2617 vdd.n757 99.5127
R2557 vdd.n2617 vdd.n751 99.5127
R2558 vdd.n2700 vdd.n751 99.5127
R2559 vdd.n2700 vdd.n746 99.5127
R2560 vdd.n2696 vdd.n746 99.5127
R2561 vdd.n2696 vdd.n741 99.5127
R2562 vdd.n2693 vdd.n741 99.5127
R2563 vdd.n2693 vdd.n735 99.5127
R2564 vdd.n2690 vdd.n735 99.5127
R2565 vdd.n2690 vdd.n728 99.5127
R2566 vdd.n2649 vdd.n728 99.5127
R2567 vdd.n2649 vdd.n723 99.5127
R2568 vdd.n2646 vdd.n723 99.5127
R2569 vdd.n2646 vdd.n718 99.5127
R2570 vdd.n2643 vdd.n718 99.5127
R2571 vdd.n2643 vdd.n711 99.5127
R2572 vdd.n2640 vdd.n711 99.5127
R2573 vdd.n2640 vdd.n704 99.5127
R2574 vdd.n2637 vdd.n704 99.5127
R2575 vdd.n2637 vdd.n697 99.5127
R2576 vdd.n2634 vdd.n697 99.5127
R2577 vdd.n2634 vdd.n691 99.5127
R2578 vdd.n2631 vdd.n691 99.5127
R2579 vdd.n2631 vdd.n686 99.5127
R2580 vdd.n2628 vdd.n686 99.5127
R2581 vdd.n2628 vdd.n681 99.5127
R2582 vdd.n2625 vdd.n681 99.5127
R2583 vdd.n2625 vdd.n673 99.5127
R2584 vdd.n2622 vdd.n673 99.5127
R2585 vdd.n2622 vdd.n666 99.5127
R2586 vdd.n666 vdd.n630 99.5127
R2587 vdd.n2954 vdd.n630 99.5127
R2588 vdd.n2478 vdd.n2477 99.5127
R2589 vdd.n2482 vdd.n2481 99.5127
R2590 vdd.n2486 vdd.n2485 99.5127
R2591 vdd.n2490 vdd.n2489 99.5127
R2592 vdd.n2494 vdd.n2493 99.5127
R2593 vdd.n2498 vdd.n2497 99.5127
R2594 vdd.n2502 vdd.n2501 99.5127
R2595 vdd.n2506 vdd.n2505 99.5127
R2596 vdd.n2510 vdd.n2509 99.5127
R2597 vdd.n2514 vdd.n2513 99.5127
R2598 vdd.n2518 vdd.n2517 99.5127
R2599 vdd.n2522 vdd.n2521 99.5127
R2600 vdd.n2526 vdd.n2525 99.5127
R2601 vdd.n2530 vdd.n2529 99.5127
R2602 vdd.n2534 vdd.n2533 99.5127
R2603 vdd.n2538 vdd.n2537 99.5127
R2604 vdd.n2721 vdd.n2472 99.5127
R2605 vdd.n2730 vdd.n769 99.5127
R2606 vdd.n2734 vdd.n769 99.5127
R2607 vdd.n2734 vdd.n761 99.5127
R2608 vdd.n2742 vdd.n761 99.5127
R2609 vdd.n2742 vdd.n759 99.5127
R2610 vdd.n2746 vdd.n759 99.5127
R2611 vdd.n2746 vdd.n749 99.5127
R2612 vdd.n2754 vdd.n749 99.5127
R2613 vdd.n2754 vdd.n747 99.5127
R2614 vdd.n2758 vdd.n747 99.5127
R2615 vdd.n2758 vdd.n738 99.5127
R2616 vdd.n2766 vdd.n738 99.5127
R2617 vdd.n2766 vdd.n736 99.5127
R2618 vdd.n2770 vdd.n736 99.5127
R2619 vdd.n2770 vdd.n726 99.5127
R2620 vdd.n2778 vdd.n726 99.5127
R2621 vdd.n2778 vdd.n724 99.5127
R2622 vdd.n2782 vdd.n724 99.5127
R2623 vdd.n2782 vdd.n715 99.5127
R2624 vdd.n2790 vdd.n715 99.5127
R2625 vdd.n2790 vdd.n712 99.5127
R2626 vdd.n2795 vdd.n712 99.5127
R2627 vdd.n2795 vdd.n701 99.5127
R2628 vdd.n2803 vdd.n701 99.5127
R2629 vdd.n2803 vdd.n699 99.5127
R2630 vdd.n2807 vdd.n699 99.5127
R2631 vdd.n2807 vdd.n689 99.5127
R2632 vdd.n2815 vdd.n689 99.5127
R2633 vdd.n2815 vdd.n687 99.5127
R2634 vdd.n2819 vdd.n687 99.5127
R2635 vdd.n2819 vdd.n678 99.5127
R2636 vdd.n2827 vdd.n678 99.5127
R2637 vdd.n2827 vdd.n675 99.5127
R2638 vdd.n2876 vdd.n675 99.5127
R2639 vdd.n2876 vdd.n676 99.5127
R2640 vdd.n676 vdd.n667 99.5127
R2641 vdd.n2871 vdd.n667 99.5127
R2642 vdd.n2871 vdd.n633 99.5127
R2643 vdd.n2361 vdd.n2360 99.5127
R2644 vdd.n2357 vdd.n2356 99.5127
R2645 vdd.n2353 vdd.n2352 99.5127
R2646 vdd.n2349 vdd.n2348 99.5127
R2647 vdd.n2345 vdd.n2344 99.5127
R2648 vdd.n2341 vdd.n2340 99.5127
R2649 vdd.n2337 vdd.n2336 99.5127
R2650 vdd.n2333 vdd.n2332 99.5127
R2651 vdd.n2329 vdd.n2328 99.5127
R2652 vdd.n2325 vdd.n2324 99.5127
R2653 vdd.n2321 vdd.n2320 99.5127
R2654 vdd.n2317 vdd.n2316 99.5127
R2655 vdd.n2313 vdd.n2312 99.5127
R2656 vdd.n2309 vdd.n2308 99.5127
R2657 vdd.n2305 vdd.n2304 99.5127
R2658 vdd.n2301 vdd.n2300 99.5127
R2659 vdd.n2297 vdd.n795 99.5127
R2660 vdd.n1997 vdd.n940 99.5127
R2661 vdd.n1997 vdd.n934 99.5127
R2662 vdd.n2000 vdd.n934 99.5127
R2663 vdd.n2000 vdd.n928 99.5127
R2664 vdd.n2003 vdd.n928 99.5127
R2665 vdd.n2003 vdd.n922 99.5127
R2666 vdd.n2006 vdd.n922 99.5127
R2667 vdd.n2006 vdd.n916 99.5127
R2668 vdd.n2009 vdd.n916 99.5127
R2669 vdd.n2009 vdd.n910 99.5127
R2670 vdd.n2012 vdd.n910 99.5127
R2671 vdd.n2012 vdd.n904 99.5127
R2672 vdd.n2015 vdd.n904 99.5127
R2673 vdd.n2015 vdd.n897 99.5127
R2674 vdd.n2018 vdd.n897 99.5127
R2675 vdd.n2018 vdd.n890 99.5127
R2676 vdd.n2021 vdd.n890 99.5127
R2677 vdd.n2021 vdd.n884 99.5127
R2678 vdd.n2024 vdd.n884 99.5127
R2679 vdd.n2024 vdd.n879 99.5127
R2680 vdd.n2027 vdd.n879 99.5127
R2681 vdd.n2027 vdd.n873 99.5127
R2682 vdd.n2069 vdd.n873 99.5127
R2683 vdd.n2069 vdd.n866 99.5127
R2684 vdd.n2065 vdd.n866 99.5127
R2685 vdd.n2065 vdd.n860 99.5127
R2686 vdd.n2062 vdd.n860 99.5127
R2687 vdd.n2062 vdd.n855 99.5127
R2688 vdd.n2059 vdd.n855 99.5127
R2689 vdd.n2059 vdd.n850 99.5127
R2690 vdd.n2035 vdd.n850 99.5127
R2691 vdd.n2035 vdd.n845 99.5127
R2692 vdd.n2032 vdd.n845 99.5127
R2693 vdd.n2032 vdd.n838 99.5127
R2694 vdd.n838 vdd.n829 99.5127
R2695 vdd.n2292 vdd.n829 99.5127
R2696 vdd.n2293 vdd.n2292 99.5127
R2697 vdd.n2293 vdd.n821 99.5127
R2698 vdd.n1930 vdd.n1928 99.5127
R2699 vdd.n1934 vdd.n1925 99.5127
R2700 vdd.n1938 vdd.n1936 99.5127
R2701 vdd.n1942 vdd.n1923 99.5127
R2702 vdd.n1946 vdd.n1944 99.5127
R2703 vdd.n1950 vdd.n1921 99.5127
R2704 vdd.n1954 vdd.n1952 99.5127
R2705 vdd.n1958 vdd.n1919 99.5127
R2706 vdd.n1962 vdd.n1960 99.5127
R2707 vdd.n1966 vdd.n971 99.5127
R2708 vdd.n1970 vdd.n1968 99.5127
R2709 vdd.n1974 vdd.n969 99.5127
R2710 vdd.n1978 vdd.n1976 99.5127
R2711 vdd.n1982 vdd.n967 99.5127
R2712 vdd.n1986 vdd.n1984 99.5127
R2713 vdd.n1991 vdd.n963 99.5127
R2714 vdd.n1994 vdd.n1993 99.5127
R2715 vdd.n2180 vdd.n935 99.5127
R2716 vdd.n2184 vdd.n935 99.5127
R2717 vdd.n2184 vdd.n925 99.5127
R2718 vdd.n2192 vdd.n925 99.5127
R2719 vdd.n2192 vdd.n923 99.5127
R2720 vdd.n2196 vdd.n923 99.5127
R2721 vdd.n2196 vdd.n913 99.5127
R2722 vdd.n2204 vdd.n913 99.5127
R2723 vdd.n2204 vdd.n911 99.5127
R2724 vdd.n2208 vdd.n911 99.5127
R2725 vdd.n2208 vdd.n901 99.5127
R2726 vdd.n2216 vdd.n901 99.5127
R2727 vdd.n2216 vdd.n899 99.5127
R2728 vdd.n2220 vdd.n899 99.5127
R2729 vdd.n2220 vdd.n888 99.5127
R2730 vdd.n2228 vdd.n888 99.5127
R2731 vdd.n2228 vdd.n885 99.5127
R2732 vdd.n2233 vdd.n885 99.5127
R2733 vdd.n2233 vdd.n876 99.5127
R2734 vdd.n2241 vdd.n876 99.5127
R2735 vdd.n2241 vdd.n874 99.5127
R2736 vdd.n2245 vdd.n874 99.5127
R2737 vdd.n2245 vdd.n864 99.5127
R2738 vdd.n2253 vdd.n864 99.5127
R2739 vdd.n2253 vdd.n862 99.5127
R2740 vdd.n2257 vdd.n862 99.5127
R2741 vdd.n2257 vdd.n853 99.5127
R2742 vdd.n2265 vdd.n853 99.5127
R2743 vdd.n2265 vdd.n851 99.5127
R2744 vdd.n2269 vdd.n851 99.5127
R2745 vdd.n2269 vdd.n842 99.5127
R2746 vdd.n2277 vdd.n842 99.5127
R2747 vdd.n2277 vdd.n839 99.5127
R2748 vdd.n2283 vdd.n839 99.5127
R2749 vdd.n2283 vdd.n840 99.5127
R2750 vdd.n840 vdd.n831 99.5127
R2751 vdd.n831 vdd.n822 99.5127
R2752 vdd.n2365 vdd.n822 99.5127
R2753 vdd.n9 vdd.n7 98.9633
R2754 vdd.n2 vdd.n0 98.9633
R2755 vdd.n9 vdd.n8 98.6055
R2756 vdd.n11 vdd.n10 98.6055
R2757 vdd.n13 vdd.n12 98.6055
R2758 vdd.n6 vdd.n5 98.6055
R2759 vdd.n4 vdd.n3 98.6055
R2760 vdd.n2 vdd.n1 98.6055
R2761 vdd.t1 vdd.n279 85.8723
R2762 vdd.t78 vdd.n228 85.8723
R2763 vdd.t46 vdd.n185 85.8723
R2764 vdd.t229 vdd.n134 85.8723
R2765 vdd.t173 vdd.n92 85.8723
R2766 vdd.t15 vdd.n41 85.8723
R2767 vdd.t5 vdd.n1554 85.8723
R2768 vdd.t87 vdd.n1605 85.8723
R2769 vdd.t75 vdd.n1460 85.8723
R2770 vdd.t91 vdd.n1511 85.8723
R2771 vdd.t236 vdd.n1367 85.8723
R2772 vdd.t32 vdd.n1418 85.8723
R2773 vdd.n2792 vdd.n713 78.546
R2774 vdd.n2231 vdd.n886 78.546
R2775 vdd.n266 vdd.n265 75.1835
R2776 vdd.n264 vdd.n263 75.1835
R2777 vdd.n262 vdd.n261 75.1835
R2778 vdd.n260 vdd.n259 75.1835
R2779 vdd.n258 vdd.n257 75.1835
R2780 vdd.n172 vdd.n171 75.1835
R2781 vdd.n170 vdd.n169 75.1835
R2782 vdd.n168 vdd.n167 75.1835
R2783 vdd.n166 vdd.n165 75.1835
R2784 vdd.n164 vdd.n163 75.1835
R2785 vdd.n79 vdd.n78 75.1835
R2786 vdd.n77 vdd.n76 75.1835
R2787 vdd.n75 vdd.n74 75.1835
R2788 vdd.n73 vdd.n72 75.1835
R2789 vdd.n71 vdd.n70 75.1835
R2790 vdd.n1584 vdd.n1583 75.1835
R2791 vdd.n1586 vdd.n1585 75.1835
R2792 vdd.n1588 vdd.n1587 75.1835
R2793 vdd.n1590 vdd.n1589 75.1835
R2794 vdd.n1592 vdd.n1591 75.1835
R2795 vdd.n1490 vdd.n1489 75.1835
R2796 vdd.n1492 vdd.n1491 75.1835
R2797 vdd.n1494 vdd.n1493 75.1835
R2798 vdd.n1496 vdd.n1495 75.1835
R2799 vdd.n1498 vdd.n1497 75.1835
R2800 vdd.n1397 vdd.n1396 75.1835
R2801 vdd.n1399 vdd.n1398 75.1835
R2802 vdd.n1401 vdd.n1400 75.1835
R2803 vdd.n1403 vdd.n1402 75.1835
R2804 vdd.n1405 vdd.n1404 75.1835
R2805 vdd.n2722 vdd.n2455 72.8958
R2806 vdd.n2722 vdd.n2456 72.8958
R2807 vdd.n2722 vdd.n2457 72.8958
R2808 vdd.n2722 vdd.n2458 72.8958
R2809 vdd.n2722 vdd.n2459 72.8958
R2810 vdd.n2722 vdd.n2460 72.8958
R2811 vdd.n2722 vdd.n2461 72.8958
R2812 vdd.n2722 vdd.n2462 72.8958
R2813 vdd.n2722 vdd.n2463 72.8958
R2814 vdd.n2722 vdd.n2464 72.8958
R2815 vdd.n2722 vdd.n2465 72.8958
R2816 vdd.n2722 vdd.n2466 72.8958
R2817 vdd.n2722 vdd.n2467 72.8958
R2818 vdd.n2722 vdd.n2468 72.8958
R2819 vdd.n2722 vdd.n2469 72.8958
R2820 vdd.n2722 vdd.n2470 72.8958
R2821 vdd.n2722 vdd.n2471 72.8958
R2822 vdd.n629 vdd.n613 72.8958
R2823 vdd.n2960 vdd.n613 72.8958
R2824 vdd.n623 vdd.n613 72.8958
R2825 vdd.n2967 vdd.n613 72.8958
R2826 vdd.n620 vdd.n613 72.8958
R2827 vdd.n2974 vdd.n613 72.8958
R2828 vdd.n617 vdd.n613 72.8958
R2829 vdd.n2981 vdd.n613 72.8958
R2830 vdd.n2984 vdd.n613 72.8958
R2831 vdd.n2840 vdd.n613 72.8958
R2832 vdd.n2845 vdd.n613 72.8958
R2833 vdd.n2839 vdd.n613 72.8958
R2834 vdd.n2852 vdd.n613 72.8958
R2835 vdd.n2836 vdd.n613 72.8958
R2836 vdd.n2859 vdd.n613 72.8958
R2837 vdd.n2833 vdd.n613 72.8958
R2838 vdd.n2866 vdd.n613 72.8958
R2839 vdd.n2173 vdd.n938 72.8958
R2840 vdd.n943 vdd.n938 72.8958
R2841 vdd.n2166 vdd.n938 72.8958
R2842 vdd.n2160 vdd.n938 72.8958
R2843 vdd.n2158 vdd.n938 72.8958
R2844 vdd.n2152 vdd.n938 72.8958
R2845 vdd.n2150 vdd.n938 72.8958
R2846 vdd.n2144 vdd.n938 72.8958
R2847 vdd.n2142 vdd.n938 72.8958
R2848 vdd.n2136 vdd.n938 72.8958
R2849 vdd.n2134 vdd.n938 72.8958
R2850 vdd.n2128 vdd.n938 72.8958
R2851 vdd.n2126 vdd.n938 72.8958
R2852 vdd.n2120 vdd.n938 72.8958
R2853 vdd.n2118 vdd.n938 72.8958
R2854 vdd.n2111 vdd.n938 72.8958
R2855 vdd.n2109 vdd.n938 72.8958
R2856 vdd.n2438 vdd.n796 72.8958
R2857 vdd.n2438 vdd.n797 72.8958
R2858 vdd.n2438 vdd.n798 72.8958
R2859 vdd.n2438 vdd.n799 72.8958
R2860 vdd.n2438 vdd.n800 72.8958
R2861 vdd.n2438 vdd.n801 72.8958
R2862 vdd.n2438 vdd.n802 72.8958
R2863 vdd.n2438 vdd.n803 72.8958
R2864 vdd.n2438 vdd.n804 72.8958
R2865 vdd.n2438 vdd.n805 72.8958
R2866 vdd.n2438 vdd.n806 72.8958
R2867 vdd.n2438 vdd.n807 72.8958
R2868 vdd.n2438 vdd.n808 72.8958
R2869 vdd.n2438 vdd.n809 72.8958
R2870 vdd.n2438 vdd.n810 72.8958
R2871 vdd.n2438 vdd.n811 72.8958
R2872 vdd.n2438 vdd.n812 72.8958
R2873 vdd.n2723 vdd.n2722 72.8958
R2874 vdd.n2722 vdd.n2439 72.8958
R2875 vdd.n2722 vdd.n2440 72.8958
R2876 vdd.n2722 vdd.n2441 72.8958
R2877 vdd.n2722 vdd.n2442 72.8958
R2878 vdd.n2722 vdd.n2443 72.8958
R2879 vdd.n2722 vdd.n2444 72.8958
R2880 vdd.n2722 vdd.n2445 72.8958
R2881 vdd.n2722 vdd.n2446 72.8958
R2882 vdd.n2722 vdd.n2447 72.8958
R2883 vdd.n2722 vdd.n2448 72.8958
R2884 vdd.n2722 vdd.n2449 72.8958
R2885 vdd.n2722 vdd.n2450 72.8958
R2886 vdd.n2722 vdd.n2451 72.8958
R2887 vdd.n2722 vdd.n2452 72.8958
R2888 vdd.n2722 vdd.n2453 72.8958
R2889 vdd.n2722 vdd.n2454 72.8958
R2890 vdd.n2888 vdd.n613 72.8958
R2891 vdd.n2894 vdd.n613 72.8958
R2892 vdd.n659 vdd.n613 72.8958
R2893 vdd.n2901 vdd.n613 72.8958
R2894 vdd.n656 vdd.n613 72.8958
R2895 vdd.n2908 vdd.n613 72.8958
R2896 vdd.n653 vdd.n613 72.8958
R2897 vdd.n2915 vdd.n613 72.8958
R2898 vdd.n650 vdd.n613 72.8958
R2899 vdd.n2923 vdd.n613 72.8958
R2900 vdd.n647 vdd.n613 72.8958
R2901 vdd.n2930 vdd.n613 72.8958
R2902 vdd.n644 vdd.n613 72.8958
R2903 vdd.n2937 vdd.n613 72.8958
R2904 vdd.n641 vdd.n613 72.8958
R2905 vdd.n2944 vdd.n613 72.8958
R2906 vdd.n2947 vdd.n613 72.8958
R2907 vdd.n2438 vdd.n794 72.8958
R2908 vdd.n2438 vdd.n793 72.8958
R2909 vdd.n2438 vdd.n792 72.8958
R2910 vdd.n2438 vdd.n791 72.8958
R2911 vdd.n2438 vdd.n790 72.8958
R2912 vdd.n2438 vdd.n789 72.8958
R2913 vdd.n2438 vdd.n788 72.8958
R2914 vdd.n2438 vdd.n787 72.8958
R2915 vdd.n2438 vdd.n786 72.8958
R2916 vdd.n2438 vdd.n785 72.8958
R2917 vdd.n2438 vdd.n784 72.8958
R2918 vdd.n2438 vdd.n783 72.8958
R2919 vdd.n2438 vdd.n782 72.8958
R2920 vdd.n2438 vdd.n781 72.8958
R2921 vdd.n2438 vdd.n780 72.8958
R2922 vdd.n2438 vdd.n779 72.8958
R2923 vdd.n2438 vdd.n778 72.8958
R2924 vdd.n1927 vdd.n938 72.8958
R2925 vdd.n1929 vdd.n938 72.8958
R2926 vdd.n1935 vdd.n938 72.8958
R2927 vdd.n1937 vdd.n938 72.8958
R2928 vdd.n1943 vdd.n938 72.8958
R2929 vdd.n1945 vdd.n938 72.8958
R2930 vdd.n1951 vdd.n938 72.8958
R2931 vdd.n1953 vdd.n938 72.8958
R2932 vdd.n1959 vdd.n938 72.8958
R2933 vdd.n1961 vdd.n938 72.8958
R2934 vdd.n1967 vdd.n938 72.8958
R2935 vdd.n1969 vdd.n938 72.8958
R2936 vdd.n1975 vdd.n938 72.8958
R2937 vdd.n1977 vdd.n938 72.8958
R2938 vdd.n1983 vdd.n938 72.8958
R2939 vdd.n1985 vdd.n938 72.8958
R2940 vdd.n1992 vdd.n938 72.8958
R2941 vdd.n1066 vdd.n1062 66.2847
R2942 vdd.n1072 vdd.n1062 66.2847
R2943 vdd.n1075 vdd.n1062 66.2847
R2944 vdd.n1080 vdd.n1062 66.2847
R2945 vdd.n1083 vdd.n1062 66.2847
R2946 vdd.n1088 vdd.n1062 66.2847
R2947 vdd.n1091 vdd.n1062 66.2847
R2948 vdd.n1096 vdd.n1062 66.2847
R2949 vdd.n1099 vdd.n1062 66.2847
R2950 vdd.n1106 vdd.n1062 66.2847
R2951 vdd.n1109 vdd.n1062 66.2847
R2952 vdd.n1114 vdd.n1062 66.2847
R2953 vdd.n1117 vdd.n1062 66.2847
R2954 vdd.n1122 vdd.n1062 66.2847
R2955 vdd.n1125 vdd.n1062 66.2847
R2956 vdd.n1130 vdd.n1062 66.2847
R2957 vdd.n1133 vdd.n1062 66.2847
R2958 vdd.n1138 vdd.n1062 66.2847
R2959 vdd.n1141 vdd.n1062 66.2847
R2960 vdd.n1146 vdd.n1062 66.2847
R2961 vdd.n1225 vdd.n1062 66.2847
R2962 vdd.n1149 vdd.n1062 66.2847
R2963 vdd.n1155 vdd.n1062 66.2847
R2964 vdd.n1160 vdd.n1062 66.2847
R2965 vdd.n1163 vdd.n1062 66.2847
R2966 vdd.n1168 vdd.n1062 66.2847
R2967 vdd.n1171 vdd.n1062 66.2847
R2968 vdd.n1176 vdd.n1062 66.2847
R2969 vdd.n1179 vdd.n1062 66.2847
R2970 vdd.n1184 vdd.n1062 66.2847
R2971 vdd.n1187 vdd.n1062 66.2847
R2972 vdd.n981 vdd.n978 66.2847
R2973 vdd.n1792 vdd.n981 66.2847
R2974 vdd.n1797 vdd.n981 66.2847
R2975 vdd.n1802 vdd.n981 66.2847
R2976 vdd.n1790 vdd.n981 66.2847
R2977 vdd.n1809 vdd.n981 66.2847
R2978 vdd.n1782 vdd.n981 66.2847
R2979 vdd.n1816 vdd.n981 66.2847
R2980 vdd.n1775 vdd.n981 66.2847
R2981 vdd.n1823 vdd.n981 66.2847
R2982 vdd.n1769 vdd.n981 66.2847
R2983 vdd.n1764 vdd.n981 66.2847
R2984 vdd.n1834 vdd.n981 66.2847
R2985 vdd.n1756 vdd.n981 66.2847
R2986 vdd.n1841 vdd.n981 66.2847
R2987 vdd.n1749 vdd.n981 66.2847
R2988 vdd.n1848 vdd.n981 66.2847
R2989 vdd.n1742 vdd.n981 66.2847
R2990 vdd.n1855 vdd.n981 66.2847
R2991 vdd.n1735 vdd.n981 66.2847
R2992 vdd.n1862 vdd.n981 66.2847
R2993 vdd.n1729 vdd.n981 66.2847
R2994 vdd.n1724 vdd.n981 66.2847
R2995 vdd.n1873 vdd.n981 66.2847
R2996 vdd.n1716 vdd.n981 66.2847
R2997 vdd.n1880 vdd.n981 66.2847
R2998 vdd.n1709 vdd.n981 66.2847
R2999 vdd.n1887 vdd.n981 66.2847
R3000 vdd.n1890 vdd.n981 66.2847
R3001 vdd.n1700 vdd.n981 66.2847
R3002 vdd.n1899 vdd.n981 66.2847
R3003 vdd.n1694 vdd.n981 66.2847
R3004 vdd.n3114 vdd.n516 66.2847
R3005 vdd.n520 vdd.n516 66.2847
R3006 vdd.n523 vdd.n516 66.2847
R3007 vdd.n3103 vdd.n516 66.2847
R3008 vdd.n3097 vdd.n516 66.2847
R3009 vdd.n3095 vdd.n516 66.2847
R3010 vdd.n3089 vdd.n516 66.2847
R3011 vdd.n3087 vdd.n516 66.2847
R3012 vdd.n3081 vdd.n516 66.2847
R3013 vdd.n3079 vdd.n516 66.2847
R3014 vdd.n3073 vdd.n516 66.2847
R3015 vdd.n3071 vdd.n516 66.2847
R3016 vdd.n3065 vdd.n516 66.2847
R3017 vdd.n3063 vdd.n516 66.2847
R3018 vdd.n3057 vdd.n516 66.2847
R3019 vdd.n3055 vdd.n516 66.2847
R3020 vdd.n3049 vdd.n516 66.2847
R3021 vdd.n3047 vdd.n516 66.2847
R3022 vdd.n3041 vdd.n516 66.2847
R3023 vdd.n3039 vdd.n516 66.2847
R3024 vdd.n584 vdd.n516 66.2847
R3025 vdd.n3030 vdd.n516 66.2847
R3026 vdd.n586 vdd.n516 66.2847
R3027 vdd.n3023 vdd.n516 66.2847
R3028 vdd.n3017 vdd.n516 66.2847
R3029 vdd.n3015 vdd.n516 66.2847
R3030 vdd.n3009 vdd.n516 66.2847
R3031 vdd.n3007 vdd.n516 66.2847
R3032 vdd.n3001 vdd.n516 66.2847
R3033 vdd.n607 vdd.n516 66.2847
R3034 vdd.n609 vdd.n516 66.2847
R3035 vdd.n3200 vdd.n351 66.2847
R3036 vdd.n3209 vdd.n351 66.2847
R3037 vdd.n461 vdd.n351 66.2847
R3038 vdd.n3216 vdd.n351 66.2847
R3039 vdd.n454 vdd.n351 66.2847
R3040 vdd.n3223 vdd.n351 66.2847
R3041 vdd.n447 vdd.n351 66.2847
R3042 vdd.n3230 vdd.n351 66.2847
R3043 vdd.n440 vdd.n351 66.2847
R3044 vdd.n3237 vdd.n351 66.2847
R3045 vdd.n434 vdd.n351 66.2847
R3046 vdd.n429 vdd.n351 66.2847
R3047 vdd.n3248 vdd.n351 66.2847
R3048 vdd.n421 vdd.n351 66.2847
R3049 vdd.n3255 vdd.n351 66.2847
R3050 vdd.n414 vdd.n351 66.2847
R3051 vdd.n3262 vdd.n351 66.2847
R3052 vdd.n407 vdd.n351 66.2847
R3053 vdd.n3269 vdd.n351 66.2847
R3054 vdd.n400 vdd.n351 66.2847
R3055 vdd.n3276 vdd.n351 66.2847
R3056 vdd.n394 vdd.n351 66.2847
R3057 vdd.n389 vdd.n351 66.2847
R3058 vdd.n3287 vdd.n351 66.2847
R3059 vdd.n381 vdd.n351 66.2847
R3060 vdd.n3294 vdd.n351 66.2847
R3061 vdd.n374 vdd.n351 66.2847
R3062 vdd.n3301 vdd.n351 66.2847
R3063 vdd.n367 vdd.n351 66.2847
R3064 vdd.n3308 vdd.n351 66.2847
R3065 vdd.n3311 vdd.n351 66.2847
R3066 vdd.n355 vdd.n351 66.2847
R3067 vdd.n356 vdd.n355 52.4337
R3068 vdd.n3311 vdd.n3310 52.4337
R3069 vdd.n3308 vdd.n3307 52.4337
R3070 vdd.n3303 vdd.n367 52.4337
R3071 vdd.n3301 vdd.n3300 52.4337
R3072 vdd.n3296 vdd.n374 52.4337
R3073 vdd.n3294 vdd.n3293 52.4337
R3074 vdd.n3289 vdd.n381 52.4337
R3075 vdd.n3287 vdd.n3286 52.4337
R3076 vdd.n390 vdd.n389 52.4337
R3077 vdd.n3278 vdd.n394 52.4337
R3078 vdd.n3276 vdd.n3275 52.4337
R3079 vdd.n3271 vdd.n400 52.4337
R3080 vdd.n3269 vdd.n3268 52.4337
R3081 vdd.n3264 vdd.n407 52.4337
R3082 vdd.n3262 vdd.n3261 52.4337
R3083 vdd.n3257 vdd.n414 52.4337
R3084 vdd.n3255 vdd.n3254 52.4337
R3085 vdd.n3250 vdd.n421 52.4337
R3086 vdd.n3248 vdd.n3247 52.4337
R3087 vdd.n430 vdd.n429 52.4337
R3088 vdd.n3239 vdd.n434 52.4337
R3089 vdd.n3237 vdd.n3236 52.4337
R3090 vdd.n3232 vdd.n440 52.4337
R3091 vdd.n3230 vdd.n3229 52.4337
R3092 vdd.n3225 vdd.n447 52.4337
R3093 vdd.n3223 vdd.n3222 52.4337
R3094 vdd.n3218 vdd.n454 52.4337
R3095 vdd.n3216 vdd.n3215 52.4337
R3096 vdd.n3211 vdd.n461 52.4337
R3097 vdd.n3209 vdd.n3208 52.4337
R3098 vdd.n3201 vdd.n3200 52.4337
R3099 vdd.n3114 vdd.n517 52.4337
R3100 vdd.n3112 vdd.n520 52.4337
R3101 vdd.n3108 vdd.n523 52.4337
R3102 vdd.n3104 vdd.n3103 52.4337
R3103 vdd.n3097 vdd.n526 52.4337
R3104 vdd.n3096 vdd.n3095 52.4337
R3105 vdd.n3089 vdd.n532 52.4337
R3106 vdd.n3088 vdd.n3087 52.4337
R3107 vdd.n3081 vdd.n538 52.4337
R3108 vdd.n3080 vdd.n3079 52.4337
R3109 vdd.n3073 vdd.n546 52.4337
R3110 vdd.n3072 vdd.n3071 52.4337
R3111 vdd.n3065 vdd.n552 52.4337
R3112 vdd.n3064 vdd.n3063 52.4337
R3113 vdd.n3057 vdd.n558 52.4337
R3114 vdd.n3056 vdd.n3055 52.4337
R3115 vdd.n3049 vdd.n564 52.4337
R3116 vdd.n3048 vdd.n3047 52.4337
R3117 vdd.n3041 vdd.n570 52.4337
R3118 vdd.n3040 vdd.n3039 52.4337
R3119 vdd.n584 vdd.n576 52.4337
R3120 vdd.n3031 vdd.n3030 52.4337
R3121 vdd.n3028 vdd.n586 52.4337
R3122 vdd.n3024 vdd.n3023 52.4337
R3123 vdd.n3017 vdd.n590 52.4337
R3124 vdd.n3016 vdd.n3015 52.4337
R3125 vdd.n3009 vdd.n596 52.4337
R3126 vdd.n3008 vdd.n3007 52.4337
R3127 vdd.n3001 vdd.n602 52.4337
R3128 vdd.n3000 vdd.n607 52.4337
R3129 vdd.n2996 vdd.n609 52.4337
R3130 vdd.n1901 vdd.n1694 52.4337
R3131 vdd.n1899 vdd.n1898 52.4337
R3132 vdd.n1701 vdd.n1700 52.4337
R3133 vdd.n1890 vdd.n1889 52.4337
R3134 vdd.n1887 vdd.n1886 52.4337
R3135 vdd.n1882 vdd.n1709 52.4337
R3136 vdd.n1880 vdd.n1879 52.4337
R3137 vdd.n1875 vdd.n1716 52.4337
R3138 vdd.n1873 vdd.n1872 52.4337
R3139 vdd.n1725 vdd.n1724 52.4337
R3140 vdd.n1864 vdd.n1729 52.4337
R3141 vdd.n1862 vdd.n1861 52.4337
R3142 vdd.n1857 vdd.n1735 52.4337
R3143 vdd.n1855 vdd.n1854 52.4337
R3144 vdd.n1850 vdd.n1742 52.4337
R3145 vdd.n1848 vdd.n1847 52.4337
R3146 vdd.n1843 vdd.n1749 52.4337
R3147 vdd.n1841 vdd.n1840 52.4337
R3148 vdd.n1836 vdd.n1756 52.4337
R3149 vdd.n1834 vdd.n1833 52.4337
R3150 vdd.n1765 vdd.n1764 52.4337
R3151 vdd.n1825 vdd.n1769 52.4337
R3152 vdd.n1823 vdd.n1822 52.4337
R3153 vdd.n1818 vdd.n1775 52.4337
R3154 vdd.n1816 vdd.n1815 52.4337
R3155 vdd.n1811 vdd.n1782 52.4337
R3156 vdd.n1809 vdd.n1808 52.4337
R3157 vdd.n1804 vdd.n1790 52.4337
R3158 vdd.n1802 vdd.n1801 52.4337
R3159 vdd.n1797 vdd.n1796 52.4337
R3160 vdd.n1792 vdd.n1791 52.4337
R3161 vdd.n1910 vdd.n978 52.4337
R3162 vdd.n1066 vdd.n1064 52.4337
R3163 vdd.n1072 vdd.n1071 52.4337
R3164 vdd.n1075 vdd.n1074 52.4337
R3165 vdd.n1080 vdd.n1079 52.4337
R3166 vdd.n1083 vdd.n1082 52.4337
R3167 vdd.n1088 vdd.n1087 52.4337
R3168 vdd.n1091 vdd.n1090 52.4337
R3169 vdd.n1096 vdd.n1095 52.4337
R3170 vdd.n1099 vdd.n1098 52.4337
R3171 vdd.n1106 vdd.n1105 52.4337
R3172 vdd.n1109 vdd.n1108 52.4337
R3173 vdd.n1114 vdd.n1113 52.4337
R3174 vdd.n1117 vdd.n1116 52.4337
R3175 vdd.n1122 vdd.n1121 52.4337
R3176 vdd.n1125 vdd.n1124 52.4337
R3177 vdd.n1130 vdd.n1129 52.4337
R3178 vdd.n1133 vdd.n1132 52.4337
R3179 vdd.n1138 vdd.n1137 52.4337
R3180 vdd.n1141 vdd.n1140 52.4337
R3181 vdd.n1146 vdd.n1145 52.4337
R3182 vdd.n1226 vdd.n1225 52.4337
R3183 vdd.n1223 vdd.n1149 52.4337
R3184 vdd.n1155 vdd.n1154 52.4337
R3185 vdd.n1160 vdd.n1157 52.4337
R3186 vdd.n1163 vdd.n1162 52.4337
R3187 vdd.n1168 vdd.n1165 52.4337
R3188 vdd.n1171 vdd.n1170 52.4337
R3189 vdd.n1176 vdd.n1173 52.4337
R3190 vdd.n1179 vdd.n1178 52.4337
R3191 vdd.n1184 vdd.n1181 52.4337
R3192 vdd.n1187 vdd.n1186 52.4337
R3193 vdd.n1067 vdd.n1066 52.4337
R3194 vdd.n1073 vdd.n1072 52.4337
R3195 vdd.n1076 vdd.n1075 52.4337
R3196 vdd.n1081 vdd.n1080 52.4337
R3197 vdd.n1084 vdd.n1083 52.4337
R3198 vdd.n1089 vdd.n1088 52.4337
R3199 vdd.n1092 vdd.n1091 52.4337
R3200 vdd.n1097 vdd.n1096 52.4337
R3201 vdd.n1100 vdd.n1099 52.4337
R3202 vdd.n1107 vdd.n1106 52.4337
R3203 vdd.n1110 vdd.n1109 52.4337
R3204 vdd.n1115 vdd.n1114 52.4337
R3205 vdd.n1118 vdd.n1117 52.4337
R3206 vdd.n1123 vdd.n1122 52.4337
R3207 vdd.n1126 vdd.n1125 52.4337
R3208 vdd.n1131 vdd.n1130 52.4337
R3209 vdd.n1134 vdd.n1133 52.4337
R3210 vdd.n1139 vdd.n1138 52.4337
R3211 vdd.n1142 vdd.n1141 52.4337
R3212 vdd.n1147 vdd.n1146 52.4337
R3213 vdd.n1225 vdd.n1224 52.4337
R3214 vdd.n1153 vdd.n1149 52.4337
R3215 vdd.n1156 vdd.n1155 52.4337
R3216 vdd.n1161 vdd.n1160 52.4337
R3217 vdd.n1164 vdd.n1163 52.4337
R3218 vdd.n1169 vdd.n1168 52.4337
R3219 vdd.n1172 vdd.n1171 52.4337
R3220 vdd.n1177 vdd.n1176 52.4337
R3221 vdd.n1180 vdd.n1179 52.4337
R3222 vdd.n1185 vdd.n1184 52.4337
R3223 vdd.n1188 vdd.n1187 52.4337
R3224 vdd.n978 vdd.n977 52.4337
R3225 vdd.n1793 vdd.n1792 52.4337
R3226 vdd.n1798 vdd.n1797 52.4337
R3227 vdd.n1803 vdd.n1802 52.4337
R3228 vdd.n1790 vdd.n1783 52.4337
R3229 vdd.n1810 vdd.n1809 52.4337
R3230 vdd.n1782 vdd.n1776 52.4337
R3231 vdd.n1817 vdd.n1816 52.4337
R3232 vdd.n1775 vdd.n1770 52.4337
R3233 vdd.n1824 vdd.n1823 52.4337
R3234 vdd.n1769 vdd.n1768 52.4337
R3235 vdd.n1764 vdd.n1757 52.4337
R3236 vdd.n1835 vdd.n1834 52.4337
R3237 vdd.n1756 vdd.n1750 52.4337
R3238 vdd.n1842 vdd.n1841 52.4337
R3239 vdd.n1749 vdd.n1743 52.4337
R3240 vdd.n1849 vdd.n1848 52.4337
R3241 vdd.n1742 vdd.n1736 52.4337
R3242 vdd.n1856 vdd.n1855 52.4337
R3243 vdd.n1735 vdd.n1730 52.4337
R3244 vdd.n1863 vdd.n1862 52.4337
R3245 vdd.n1729 vdd.n1728 52.4337
R3246 vdd.n1724 vdd.n1717 52.4337
R3247 vdd.n1874 vdd.n1873 52.4337
R3248 vdd.n1716 vdd.n1710 52.4337
R3249 vdd.n1881 vdd.n1880 52.4337
R3250 vdd.n1709 vdd.n1703 52.4337
R3251 vdd.n1888 vdd.n1887 52.4337
R3252 vdd.n1891 vdd.n1890 52.4337
R3253 vdd.n1700 vdd.n1695 52.4337
R3254 vdd.n1900 vdd.n1899 52.4337
R3255 vdd.n1694 vdd.n983 52.4337
R3256 vdd.n3115 vdd.n3114 52.4337
R3257 vdd.n3109 vdd.n520 52.4337
R3258 vdd.n3105 vdd.n523 52.4337
R3259 vdd.n3103 vdd.n3102 52.4337
R3260 vdd.n3098 vdd.n3097 52.4337
R3261 vdd.n3095 vdd.n3094 52.4337
R3262 vdd.n3090 vdd.n3089 52.4337
R3263 vdd.n3087 vdd.n3086 52.4337
R3264 vdd.n3082 vdd.n3081 52.4337
R3265 vdd.n3079 vdd.n3078 52.4337
R3266 vdd.n3074 vdd.n3073 52.4337
R3267 vdd.n3071 vdd.n3070 52.4337
R3268 vdd.n3066 vdd.n3065 52.4337
R3269 vdd.n3063 vdd.n3062 52.4337
R3270 vdd.n3058 vdd.n3057 52.4337
R3271 vdd.n3055 vdd.n3054 52.4337
R3272 vdd.n3050 vdd.n3049 52.4337
R3273 vdd.n3047 vdd.n3046 52.4337
R3274 vdd.n3042 vdd.n3041 52.4337
R3275 vdd.n3039 vdd.n3038 52.4337
R3276 vdd.n585 vdd.n584 52.4337
R3277 vdd.n3030 vdd.n3029 52.4337
R3278 vdd.n3025 vdd.n586 52.4337
R3279 vdd.n3023 vdd.n3022 52.4337
R3280 vdd.n3018 vdd.n3017 52.4337
R3281 vdd.n3015 vdd.n3014 52.4337
R3282 vdd.n3010 vdd.n3009 52.4337
R3283 vdd.n3007 vdd.n3006 52.4337
R3284 vdd.n3002 vdd.n3001 52.4337
R3285 vdd.n2997 vdd.n607 52.4337
R3286 vdd.n2993 vdd.n609 52.4337
R3287 vdd.n3200 vdd.n462 52.4337
R3288 vdd.n3210 vdd.n3209 52.4337
R3289 vdd.n461 vdd.n455 52.4337
R3290 vdd.n3217 vdd.n3216 52.4337
R3291 vdd.n454 vdd.n448 52.4337
R3292 vdd.n3224 vdd.n3223 52.4337
R3293 vdd.n447 vdd.n441 52.4337
R3294 vdd.n3231 vdd.n3230 52.4337
R3295 vdd.n440 vdd.n435 52.4337
R3296 vdd.n3238 vdd.n3237 52.4337
R3297 vdd.n434 vdd.n433 52.4337
R3298 vdd.n429 vdd.n422 52.4337
R3299 vdd.n3249 vdd.n3248 52.4337
R3300 vdd.n421 vdd.n415 52.4337
R3301 vdd.n3256 vdd.n3255 52.4337
R3302 vdd.n414 vdd.n408 52.4337
R3303 vdd.n3263 vdd.n3262 52.4337
R3304 vdd.n407 vdd.n401 52.4337
R3305 vdd.n3270 vdd.n3269 52.4337
R3306 vdd.n400 vdd.n395 52.4337
R3307 vdd.n3277 vdd.n3276 52.4337
R3308 vdd.n394 vdd.n393 52.4337
R3309 vdd.n389 vdd.n382 52.4337
R3310 vdd.n3288 vdd.n3287 52.4337
R3311 vdd.n381 vdd.n375 52.4337
R3312 vdd.n3295 vdd.n3294 52.4337
R3313 vdd.n374 vdd.n368 52.4337
R3314 vdd.n3302 vdd.n3301 52.4337
R3315 vdd.n367 vdd.n360 52.4337
R3316 vdd.n3309 vdd.n3308 52.4337
R3317 vdd.n3312 vdd.n3311 52.4337
R3318 vdd.n355 vdd.n352 52.4337
R3319 vdd.t187 vdd.t200 51.4683
R3320 vdd.n258 vdd.n256 42.0461
R3321 vdd.n164 vdd.n162 42.0461
R3322 vdd.n71 vdd.n69 42.0461
R3323 vdd.n1584 vdd.n1582 42.0461
R3324 vdd.n1490 vdd.n1488 42.0461
R3325 vdd.n1397 vdd.n1395 42.0461
R3326 vdd.n308 vdd.n307 41.6884
R3327 vdd.n214 vdd.n213 41.6884
R3328 vdd.n121 vdd.n120 41.6884
R3329 vdd.n1634 vdd.n1633 41.6884
R3330 vdd.n1540 vdd.n1539 41.6884
R3331 vdd.n1447 vdd.n1446 41.6884
R3332 vdd.n1192 vdd.n1191 41.1157
R3333 vdd.n1229 vdd.n1228 41.1157
R3334 vdd.n1103 vdd.n1102 41.1157
R3335 vdd.n3205 vdd.n3204 41.1157
R3336 vdd.n3244 vdd.n428 41.1157
R3337 vdd.n3283 vdd.n388 41.1157
R3338 vdd.n2947 vdd.n2946 39.2114
R3339 vdd.n2944 vdd.n2943 39.2114
R3340 vdd.n2939 vdd.n641 39.2114
R3341 vdd.n2937 vdd.n2936 39.2114
R3342 vdd.n2932 vdd.n644 39.2114
R3343 vdd.n2930 vdd.n2929 39.2114
R3344 vdd.n2925 vdd.n647 39.2114
R3345 vdd.n2923 vdd.n2922 39.2114
R3346 vdd.n2917 vdd.n650 39.2114
R3347 vdd.n2915 vdd.n2914 39.2114
R3348 vdd.n2910 vdd.n653 39.2114
R3349 vdd.n2908 vdd.n2907 39.2114
R3350 vdd.n2903 vdd.n656 39.2114
R3351 vdd.n2901 vdd.n2900 39.2114
R3352 vdd.n2896 vdd.n659 39.2114
R3353 vdd.n2894 vdd.n2893 39.2114
R3354 vdd.n2889 vdd.n2888 39.2114
R3355 vdd.n2723 vdd.n775 39.2114
R3356 vdd.n2544 vdd.n2439 39.2114
R3357 vdd.n2548 vdd.n2440 39.2114
R3358 vdd.n2552 vdd.n2441 39.2114
R3359 vdd.n2556 vdd.n2442 39.2114
R3360 vdd.n2560 vdd.n2443 39.2114
R3361 vdd.n2564 vdd.n2444 39.2114
R3362 vdd.n2568 vdd.n2445 39.2114
R3363 vdd.n2572 vdd.n2446 39.2114
R3364 vdd.n2576 vdd.n2447 39.2114
R3365 vdd.n2580 vdd.n2448 39.2114
R3366 vdd.n2584 vdd.n2449 39.2114
R3367 vdd.n2588 vdd.n2450 39.2114
R3368 vdd.n2592 vdd.n2451 39.2114
R3369 vdd.n2596 vdd.n2452 39.2114
R3370 vdd.n2600 vdd.n2453 39.2114
R3371 vdd.n2605 vdd.n2454 39.2114
R3372 vdd.n2433 vdd.n812 39.2114
R3373 vdd.n2429 vdd.n811 39.2114
R3374 vdd.n2425 vdd.n810 39.2114
R3375 vdd.n2421 vdd.n809 39.2114
R3376 vdd.n2417 vdd.n808 39.2114
R3377 vdd.n2413 vdd.n807 39.2114
R3378 vdd.n2409 vdd.n806 39.2114
R3379 vdd.n2405 vdd.n805 39.2114
R3380 vdd.n2401 vdd.n804 39.2114
R3381 vdd.n2397 vdd.n803 39.2114
R3382 vdd.n2393 vdd.n802 39.2114
R3383 vdd.n2389 vdd.n801 39.2114
R3384 vdd.n2385 vdd.n800 39.2114
R3385 vdd.n2381 vdd.n799 39.2114
R3386 vdd.n2377 vdd.n798 39.2114
R3387 vdd.n2372 vdd.n797 39.2114
R3388 vdd.n2368 vdd.n796 39.2114
R3389 vdd.n2173 vdd.n941 39.2114
R3390 vdd.n2171 vdd.n943 39.2114
R3391 vdd.n2167 vdd.n2166 39.2114
R3392 vdd.n2160 vdd.n945 39.2114
R3393 vdd.n2159 vdd.n2158 39.2114
R3394 vdd.n2152 vdd.n947 39.2114
R3395 vdd.n2151 vdd.n2150 39.2114
R3396 vdd.n2144 vdd.n949 39.2114
R3397 vdd.n2143 vdd.n2142 39.2114
R3398 vdd.n2136 vdd.n951 39.2114
R3399 vdd.n2135 vdd.n2134 39.2114
R3400 vdd.n2128 vdd.n953 39.2114
R3401 vdd.n2127 vdd.n2126 39.2114
R3402 vdd.n2120 vdd.n955 39.2114
R3403 vdd.n2119 vdd.n2118 39.2114
R3404 vdd.n2111 vdd.n957 39.2114
R3405 vdd.n2110 vdd.n2109 39.2114
R3406 vdd.n2866 vdd.n2865 39.2114
R3407 vdd.n2861 vdd.n2833 39.2114
R3408 vdd.n2859 vdd.n2858 39.2114
R3409 vdd.n2854 vdd.n2836 39.2114
R3410 vdd.n2852 vdd.n2851 39.2114
R3411 vdd.n2847 vdd.n2839 39.2114
R3412 vdd.n2845 vdd.n2844 39.2114
R3413 vdd.n2840 vdd.n612 39.2114
R3414 vdd.n2984 vdd.n2983 39.2114
R3415 vdd.n2981 vdd.n2980 39.2114
R3416 vdd.n2976 vdd.n617 39.2114
R3417 vdd.n2974 vdd.n2973 39.2114
R3418 vdd.n2969 vdd.n620 39.2114
R3419 vdd.n2967 vdd.n2966 39.2114
R3420 vdd.n2962 vdd.n623 39.2114
R3421 vdd.n2960 vdd.n2959 39.2114
R3422 vdd.n2955 vdd.n629 39.2114
R3423 vdd.n2455 vdd.n771 39.2114
R3424 vdd.n2478 vdd.n2456 39.2114
R3425 vdd.n2482 vdd.n2457 39.2114
R3426 vdd.n2486 vdd.n2458 39.2114
R3427 vdd.n2490 vdd.n2459 39.2114
R3428 vdd.n2494 vdd.n2460 39.2114
R3429 vdd.n2498 vdd.n2461 39.2114
R3430 vdd.n2502 vdd.n2462 39.2114
R3431 vdd.n2506 vdd.n2463 39.2114
R3432 vdd.n2510 vdd.n2464 39.2114
R3433 vdd.n2514 vdd.n2465 39.2114
R3434 vdd.n2518 vdd.n2466 39.2114
R3435 vdd.n2522 vdd.n2467 39.2114
R3436 vdd.n2526 vdd.n2468 39.2114
R3437 vdd.n2530 vdd.n2469 39.2114
R3438 vdd.n2534 vdd.n2470 39.2114
R3439 vdd.n2538 vdd.n2471 39.2114
R3440 vdd.n2477 vdd.n2455 39.2114
R3441 vdd.n2481 vdd.n2456 39.2114
R3442 vdd.n2485 vdd.n2457 39.2114
R3443 vdd.n2489 vdd.n2458 39.2114
R3444 vdd.n2493 vdd.n2459 39.2114
R3445 vdd.n2497 vdd.n2460 39.2114
R3446 vdd.n2501 vdd.n2461 39.2114
R3447 vdd.n2505 vdd.n2462 39.2114
R3448 vdd.n2509 vdd.n2463 39.2114
R3449 vdd.n2513 vdd.n2464 39.2114
R3450 vdd.n2517 vdd.n2465 39.2114
R3451 vdd.n2521 vdd.n2466 39.2114
R3452 vdd.n2525 vdd.n2467 39.2114
R3453 vdd.n2529 vdd.n2468 39.2114
R3454 vdd.n2533 vdd.n2469 39.2114
R3455 vdd.n2537 vdd.n2470 39.2114
R3456 vdd.n2472 vdd.n2471 39.2114
R3457 vdd.n629 vdd.n624 39.2114
R3458 vdd.n2961 vdd.n2960 39.2114
R3459 vdd.n623 vdd.n621 39.2114
R3460 vdd.n2968 vdd.n2967 39.2114
R3461 vdd.n620 vdd.n618 39.2114
R3462 vdd.n2975 vdd.n2974 39.2114
R3463 vdd.n617 vdd.n615 39.2114
R3464 vdd.n2982 vdd.n2981 39.2114
R3465 vdd.n2985 vdd.n2984 39.2114
R3466 vdd.n2841 vdd.n2840 39.2114
R3467 vdd.n2846 vdd.n2845 39.2114
R3468 vdd.n2839 vdd.n2837 39.2114
R3469 vdd.n2853 vdd.n2852 39.2114
R3470 vdd.n2836 vdd.n2834 39.2114
R3471 vdd.n2860 vdd.n2859 39.2114
R3472 vdd.n2833 vdd.n2831 39.2114
R3473 vdd.n2867 vdd.n2866 39.2114
R3474 vdd.n2174 vdd.n2173 39.2114
R3475 vdd.n2168 vdd.n943 39.2114
R3476 vdd.n2166 vdd.n2165 39.2114
R3477 vdd.n2161 vdd.n2160 39.2114
R3478 vdd.n2158 vdd.n2157 39.2114
R3479 vdd.n2153 vdd.n2152 39.2114
R3480 vdd.n2150 vdd.n2149 39.2114
R3481 vdd.n2145 vdd.n2144 39.2114
R3482 vdd.n2142 vdd.n2141 39.2114
R3483 vdd.n2137 vdd.n2136 39.2114
R3484 vdd.n2134 vdd.n2133 39.2114
R3485 vdd.n2129 vdd.n2128 39.2114
R3486 vdd.n2126 vdd.n2125 39.2114
R3487 vdd.n2121 vdd.n2120 39.2114
R3488 vdd.n2118 vdd.n2117 39.2114
R3489 vdd.n2112 vdd.n2111 39.2114
R3490 vdd.n2109 vdd.n2108 39.2114
R3491 vdd.n2371 vdd.n796 39.2114
R3492 vdd.n2376 vdd.n797 39.2114
R3493 vdd.n2380 vdd.n798 39.2114
R3494 vdd.n2384 vdd.n799 39.2114
R3495 vdd.n2388 vdd.n800 39.2114
R3496 vdd.n2392 vdd.n801 39.2114
R3497 vdd.n2396 vdd.n802 39.2114
R3498 vdd.n2400 vdd.n803 39.2114
R3499 vdd.n2404 vdd.n804 39.2114
R3500 vdd.n2408 vdd.n805 39.2114
R3501 vdd.n2412 vdd.n806 39.2114
R3502 vdd.n2416 vdd.n807 39.2114
R3503 vdd.n2420 vdd.n808 39.2114
R3504 vdd.n2424 vdd.n809 39.2114
R3505 vdd.n2428 vdd.n810 39.2114
R3506 vdd.n2432 vdd.n811 39.2114
R3507 vdd.n814 vdd.n812 39.2114
R3508 vdd.n2724 vdd.n2723 39.2114
R3509 vdd.n2547 vdd.n2439 39.2114
R3510 vdd.n2551 vdd.n2440 39.2114
R3511 vdd.n2555 vdd.n2441 39.2114
R3512 vdd.n2559 vdd.n2442 39.2114
R3513 vdd.n2563 vdd.n2443 39.2114
R3514 vdd.n2567 vdd.n2444 39.2114
R3515 vdd.n2571 vdd.n2445 39.2114
R3516 vdd.n2575 vdd.n2446 39.2114
R3517 vdd.n2579 vdd.n2447 39.2114
R3518 vdd.n2583 vdd.n2448 39.2114
R3519 vdd.n2587 vdd.n2449 39.2114
R3520 vdd.n2591 vdd.n2450 39.2114
R3521 vdd.n2595 vdd.n2451 39.2114
R3522 vdd.n2599 vdd.n2452 39.2114
R3523 vdd.n2604 vdd.n2453 39.2114
R3524 vdd.n2607 vdd.n2454 39.2114
R3525 vdd.n2888 vdd.n660 39.2114
R3526 vdd.n2895 vdd.n2894 39.2114
R3527 vdd.n659 vdd.n657 39.2114
R3528 vdd.n2902 vdd.n2901 39.2114
R3529 vdd.n656 vdd.n654 39.2114
R3530 vdd.n2909 vdd.n2908 39.2114
R3531 vdd.n653 vdd.n651 39.2114
R3532 vdd.n2916 vdd.n2915 39.2114
R3533 vdd.n650 vdd.n648 39.2114
R3534 vdd.n2924 vdd.n2923 39.2114
R3535 vdd.n647 vdd.n645 39.2114
R3536 vdd.n2931 vdd.n2930 39.2114
R3537 vdd.n644 vdd.n642 39.2114
R3538 vdd.n2938 vdd.n2937 39.2114
R3539 vdd.n641 vdd.n639 39.2114
R3540 vdd.n2945 vdd.n2944 39.2114
R3541 vdd.n2948 vdd.n2947 39.2114
R3542 vdd.n823 vdd.n778 39.2114
R3543 vdd.n2360 vdd.n779 39.2114
R3544 vdd.n2356 vdd.n780 39.2114
R3545 vdd.n2352 vdd.n781 39.2114
R3546 vdd.n2348 vdd.n782 39.2114
R3547 vdd.n2344 vdd.n783 39.2114
R3548 vdd.n2340 vdd.n784 39.2114
R3549 vdd.n2336 vdd.n785 39.2114
R3550 vdd.n2332 vdd.n786 39.2114
R3551 vdd.n2328 vdd.n787 39.2114
R3552 vdd.n2324 vdd.n788 39.2114
R3553 vdd.n2320 vdd.n789 39.2114
R3554 vdd.n2316 vdd.n790 39.2114
R3555 vdd.n2312 vdd.n791 39.2114
R3556 vdd.n2308 vdd.n792 39.2114
R3557 vdd.n2304 vdd.n793 39.2114
R3558 vdd.n2300 vdd.n794 39.2114
R3559 vdd.n1927 vdd.n937 39.2114
R3560 vdd.n1930 vdd.n1929 39.2114
R3561 vdd.n1935 vdd.n1934 39.2114
R3562 vdd.n1938 vdd.n1937 39.2114
R3563 vdd.n1943 vdd.n1942 39.2114
R3564 vdd.n1946 vdd.n1945 39.2114
R3565 vdd.n1951 vdd.n1950 39.2114
R3566 vdd.n1954 vdd.n1953 39.2114
R3567 vdd.n1959 vdd.n1958 39.2114
R3568 vdd.n1962 vdd.n1961 39.2114
R3569 vdd.n1967 vdd.n1966 39.2114
R3570 vdd.n1970 vdd.n1969 39.2114
R3571 vdd.n1975 vdd.n1974 39.2114
R3572 vdd.n1978 vdd.n1977 39.2114
R3573 vdd.n1983 vdd.n1982 39.2114
R3574 vdd.n1986 vdd.n1985 39.2114
R3575 vdd.n1992 vdd.n1991 39.2114
R3576 vdd.n2297 vdd.n794 39.2114
R3577 vdd.n2301 vdd.n793 39.2114
R3578 vdd.n2305 vdd.n792 39.2114
R3579 vdd.n2309 vdd.n791 39.2114
R3580 vdd.n2313 vdd.n790 39.2114
R3581 vdd.n2317 vdd.n789 39.2114
R3582 vdd.n2321 vdd.n788 39.2114
R3583 vdd.n2325 vdd.n787 39.2114
R3584 vdd.n2329 vdd.n786 39.2114
R3585 vdd.n2333 vdd.n785 39.2114
R3586 vdd.n2337 vdd.n784 39.2114
R3587 vdd.n2341 vdd.n783 39.2114
R3588 vdd.n2345 vdd.n782 39.2114
R3589 vdd.n2349 vdd.n781 39.2114
R3590 vdd.n2353 vdd.n780 39.2114
R3591 vdd.n2357 vdd.n779 39.2114
R3592 vdd.n2361 vdd.n778 39.2114
R3593 vdd.n1928 vdd.n1927 39.2114
R3594 vdd.n1929 vdd.n1925 39.2114
R3595 vdd.n1936 vdd.n1935 39.2114
R3596 vdd.n1937 vdd.n1923 39.2114
R3597 vdd.n1944 vdd.n1943 39.2114
R3598 vdd.n1945 vdd.n1921 39.2114
R3599 vdd.n1952 vdd.n1951 39.2114
R3600 vdd.n1953 vdd.n1919 39.2114
R3601 vdd.n1960 vdd.n1959 39.2114
R3602 vdd.n1961 vdd.n971 39.2114
R3603 vdd.n1968 vdd.n1967 39.2114
R3604 vdd.n1969 vdd.n969 39.2114
R3605 vdd.n1976 vdd.n1975 39.2114
R3606 vdd.n1977 vdd.n967 39.2114
R3607 vdd.n1984 vdd.n1983 39.2114
R3608 vdd.n1985 vdd.n963 39.2114
R3609 vdd.n1993 vdd.n1992 39.2114
R3610 vdd.n1914 vdd.n1913 37.2369
R3611 vdd.n1830 vdd.n1763 37.2369
R3612 vdd.n1869 vdd.n1723 37.2369
R3613 vdd.n3036 vdd.n581 37.2369
R3614 vdd.n545 vdd.n544 37.2369
R3615 vdd.n2992 vdd.n2991 37.2369
R3616 vdd.n1989 vdd.n965 30.449
R3617 vdd.n827 vdd.n826 30.449
R3618 vdd.n2114 vdd.n959 30.449
R3619 vdd.n2374 vdd.n817 30.449
R3620 vdd.n2475 vdd.n2474 30.449
R3621 vdd.n663 vdd.n662 30.449
R3622 vdd.n2602 vdd.n2543 30.449
R3623 vdd.n627 vdd.n626 30.449
R3624 vdd.n2177 vdd.n2176 30.4395
R3625 vdd.n2436 vdd.n815 30.4395
R3626 vdd.n2369 vdd.n818 30.4395
R3627 vdd.n2107 vdd.n2106 30.4395
R3628 vdd.n2609 vdd.n2608 30.4395
R3629 vdd.n2890 vdd.n2887 30.4395
R3630 vdd.n2727 vdd.n2726 30.4395
R3631 vdd.n2951 vdd.n2950 30.4395
R3632 vdd.n2870 vdd.n2869 30.4395
R3633 vdd.n2956 vdd.n628 30.4395
R3634 vdd.n2720 vdd.n2719 30.4395
R3635 vdd.n2731 vdd.n770 30.4395
R3636 vdd.n2181 vdd.n936 30.4395
R3637 vdd.n2364 vdd.n2363 30.4395
R3638 vdd.n2296 vdd.n2295 30.4395
R3639 vdd.n1996 vdd.n1995 30.4395
R3640 vdd.n1295 vdd.n1062 20.633
R3641 vdd.n1908 vdd.n981 20.633
R3642 vdd.n3122 vdd.n516 20.633
R3643 vdd.n3320 vdd.n351 20.633
R3644 vdd.n1297 vdd.n1059 19.3944
R3645 vdd.n1301 vdd.n1059 19.3944
R3646 vdd.n1301 vdd.n1050 19.3944
R3647 vdd.n1313 vdd.n1050 19.3944
R3648 vdd.n1313 vdd.n1048 19.3944
R3649 vdd.n1317 vdd.n1048 19.3944
R3650 vdd.n1317 vdd.n1037 19.3944
R3651 vdd.n1329 vdd.n1037 19.3944
R3652 vdd.n1329 vdd.n1035 19.3944
R3653 vdd.n1333 vdd.n1035 19.3944
R3654 vdd.n1333 vdd.n1026 19.3944
R3655 vdd.n1346 vdd.n1026 19.3944
R3656 vdd.n1346 vdd.n1024 19.3944
R3657 vdd.n1350 vdd.n1024 19.3944
R3658 vdd.n1350 vdd.n1015 19.3944
R3659 vdd.n1644 vdd.n1015 19.3944
R3660 vdd.n1644 vdd.n1013 19.3944
R3661 vdd.n1648 vdd.n1013 19.3944
R3662 vdd.n1648 vdd.n1003 19.3944
R3663 vdd.n1661 vdd.n1003 19.3944
R3664 vdd.n1661 vdd.n1001 19.3944
R3665 vdd.n1665 vdd.n1001 19.3944
R3666 vdd.n1665 vdd.n993 19.3944
R3667 vdd.n1678 vdd.n993 19.3944
R3668 vdd.n1678 vdd.n990 19.3944
R3669 vdd.n1684 vdd.n990 19.3944
R3670 vdd.n1684 vdd.n991 19.3944
R3671 vdd.n991 vdd.n980 19.3944
R3672 vdd.n1222 vdd.n1148 19.3944
R3673 vdd.n1222 vdd.n1150 19.3944
R3674 vdd.n1218 vdd.n1150 19.3944
R3675 vdd.n1218 vdd.n1217 19.3944
R3676 vdd.n1217 vdd.n1216 19.3944
R3677 vdd.n1216 vdd.n1158 19.3944
R3678 vdd.n1212 vdd.n1158 19.3944
R3679 vdd.n1212 vdd.n1211 19.3944
R3680 vdd.n1211 vdd.n1210 19.3944
R3681 vdd.n1210 vdd.n1166 19.3944
R3682 vdd.n1206 vdd.n1166 19.3944
R3683 vdd.n1206 vdd.n1205 19.3944
R3684 vdd.n1205 vdd.n1204 19.3944
R3685 vdd.n1204 vdd.n1174 19.3944
R3686 vdd.n1200 vdd.n1174 19.3944
R3687 vdd.n1200 vdd.n1199 19.3944
R3688 vdd.n1199 vdd.n1198 19.3944
R3689 vdd.n1198 vdd.n1182 19.3944
R3690 vdd.n1194 vdd.n1182 19.3944
R3691 vdd.n1194 vdd.n1193 19.3944
R3692 vdd.n1260 vdd.n1259 19.3944
R3693 vdd.n1259 vdd.n1258 19.3944
R3694 vdd.n1258 vdd.n1111 19.3944
R3695 vdd.n1254 vdd.n1111 19.3944
R3696 vdd.n1254 vdd.n1253 19.3944
R3697 vdd.n1253 vdd.n1252 19.3944
R3698 vdd.n1252 vdd.n1119 19.3944
R3699 vdd.n1248 vdd.n1119 19.3944
R3700 vdd.n1248 vdd.n1247 19.3944
R3701 vdd.n1247 vdd.n1246 19.3944
R3702 vdd.n1246 vdd.n1127 19.3944
R3703 vdd.n1242 vdd.n1127 19.3944
R3704 vdd.n1242 vdd.n1241 19.3944
R3705 vdd.n1241 vdd.n1240 19.3944
R3706 vdd.n1240 vdd.n1135 19.3944
R3707 vdd.n1236 vdd.n1135 19.3944
R3708 vdd.n1236 vdd.n1235 19.3944
R3709 vdd.n1235 vdd.n1234 19.3944
R3710 vdd.n1234 vdd.n1143 19.3944
R3711 vdd.n1230 vdd.n1143 19.3944
R3712 vdd.n1290 vdd.n1289 19.3944
R3713 vdd.n1289 vdd.n1288 19.3944
R3714 vdd.n1288 vdd.n1069 19.3944
R3715 vdd.n1284 vdd.n1069 19.3944
R3716 vdd.n1284 vdd.n1283 19.3944
R3717 vdd.n1283 vdd.n1282 19.3944
R3718 vdd.n1282 vdd.n1077 19.3944
R3719 vdd.n1278 vdd.n1077 19.3944
R3720 vdd.n1278 vdd.n1277 19.3944
R3721 vdd.n1277 vdd.n1276 19.3944
R3722 vdd.n1276 vdd.n1085 19.3944
R3723 vdd.n1272 vdd.n1085 19.3944
R3724 vdd.n1272 vdd.n1271 19.3944
R3725 vdd.n1271 vdd.n1270 19.3944
R3726 vdd.n1270 vdd.n1093 19.3944
R3727 vdd.n1266 vdd.n1093 19.3944
R3728 vdd.n1266 vdd.n1265 19.3944
R3729 vdd.n1265 vdd.n1264 19.3944
R3730 vdd.n1826 vdd.n1761 19.3944
R3731 vdd.n1826 vdd.n1767 19.3944
R3732 vdd.n1821 vdd.n1767 19.3944
R3733 vdd.n1821 vdd.n1820 19.3944
R3734 vdd.n1820 vdd.n1819 19.3944
R3735 vdd.n1819 vdd.n1774 19.3944
R3736 vdd.n1814 vdd.n1774 19.3944
R3737 vdd.n1814 vdd.n1813 19.3944
R3738 vdd.n1813 vdd.n1812 19.3944
R3739 vdd.n1812 vdd.n1781 19.3944
R3740 vdd.n1807 vdd.n1781 19.3944
R3741 vdd.n1807 vdd.n1806 19.3944
R3742 vdd.n1806 vdd.n1805 19.3944
R3743 vdd.n1805 vdd.n1789 19.3944
R3744 vdd.n1800 vdd.n1789 19.3944
R3745 vdd.n1800 vdd.n1799 19.3944
R3746 vdd.n1795 vdd.n1794 19.3944
R3747 vdd.n1915 vdd.n976 19.3944
R3748 vdd.n1865 vdd.n1721 19.3944
R3749 vdd.n1865 vdd.n1727 19.3944
R3750 vdd.n1860 vdd.n1727 19.3944
R3751 vdd.n1860 vdd.n1859 19.3944
R3752 vdd.n1859 vdd.n1858 19.3944
R3753 vdd.n1858 vdd.n1734 19.3944
R3754 vdd.n1853 vdd.n1734 19.3944
R3755 vdd.n1853 vdd.n1852 19.3944
R3756 vdd.n1852 vdd.n1851 19.3944
R3757 vdd.n1851 vdd.n1741 19.3944
R3758 vdd.n1846 vdd.n1741 19.3944
R3759 vdd.n1846 vdd.n1845 19.3944
R3760 vdd.n1845 vdd.n1844 19.3944
R3761 vdd.n1844 vdd.n1748 19.3944
R3762 vdd.n1839 vdd.n1748 19.3944
R3763 vdd.n1839 vdd.n1838 19.3944
R3764 vdd.n1838 vdd.n1837 19.3944
R3765 vdd.n1837 vdd.n1755 19.3944
R3766 vdd.n1832 vdd.n1755 19.3944
R3767 vdd.n1832 vdd.n1831 19.3944
R3768 vdd.n1903 vdd.n1902 19.3944
R3769 vdd.n1902 vdd.n1693 19.3944
R3770 vdd.n1897 vdd.n1896 19.3944
R3771 vdd.n1892 vdd.n1697 19.3944
R3772 vdd.n1892 vdd.n1699 19.3944
R3773 vdd.n1702 vdd.n1699 19.3944
R3774 vdd.n1885 vdd.n1702 19.3944
R3775 vdd.n1885 vdd.n1884 19.3944
R3776 vdd.n1884 vdd.n1883 19.3944
R3777 vdd.n1883 vdd.n1708 19.3944
R3778 vdd.n1878 vdd.n1708 19.3944
R3779 vdd.n1878 vdd.n1877 19.3944
R3780 vdd.n1877 vdd.n1876 19.3944
R3781 vdd.n1876 vdd.n1715 19.3944
R3782 vdd.n1871 vdd.n1715 19.3944
R3783 vdd.n1871 vdd.n1870 19.3944
R3784 vdd.n1293 vdd.n1056 19.3944
R3785 vdd.n1305 vdd.n1056 19.3944
R3786 vdd.n1305 vdd.n1054 19.3944
R3787 vdd.n1309 vdd.n1054 19.3944
R3788 vdd.n1309 vdd.n1044 19.3944
R3789 vdd.n1321 vdd.n1044 19.3944
R3790 vdd.n1321 vdd.n1042 19.3944
R3791 vdd.n1325 vdd.n1042 19.3944
R3792 vdd.n1325 vdd.n1032 19.3944
R3793 vdd.n1338 vdd.n1032 19.3944
R3794 vdd.n1338 vdd.n1030 19.3944
R3795 vdd.n1342 vdd.n1030 19.3944
R3796 vdd.n1342 vdd.n1021 19.3944
R3797 vdd.n1354 vdd.n1021 19.3944
R3798 vdd.n1354 vdd.n1019 19.3944
R3799 vdd.n1640 vdd.n1019 19.3944
R3800 vdd.n1640 vdd.n1009 19.3944
R3801 vdd.n1653 vdd.n1009 19.3944
R3802 vdd.n1653 vdd.n1007 19.3944
R3803 vdd.n1657 vdd.n1007 19.3944
R3804 vdd.n1657 vdd.n998 19.3944
R3805 vdd.n1670 vdd.n998 19.3944
R3806 vdd.n1670 vdd.n996 19.3944
R3807 vdd.n1674 vdd.n996 19.3944
R3808 vdd.n1674 vdd.n986 19.3944
R3809 vdd.n1689 vdd.n986 19.3944
R3810 vdd.n1689 vdd.n984 19.3944
R3811 vdd.n1906 vdd.n984 19.3944
R3812 vdd.n3124 vdd.n513 19.3944
R3813 vdd.n3128 vdd.n513 19.3944
R3814 vdd.n3128 vdd.n503 19.3944
R3815 vdd.n3140 vdd.n503 19.3944
R3816 vdd.n3140 vdd.n501 19.3944
R3817 vdd.n3144 vdd.n501 19.3944
R3818 vdd.n3144 vdd.n490 19.3944
R3819 vdd.n3156 vdd.n490 19.3944
R3820 vdd.n3156 vdd.n488 19.3944
R3821 vdd.n3160 vdd.n488 19.3944
R3822 vdd.n3160 vdd.n478 19.3944
R3823 vdd.n3173 vdd.n478 19.3944
R3824 vdd.n3173 vdd.n476 19.3944
R3825 vdd.n3177 vdd.n476 19.3944
R3826 vdd.n3178 vdd.n3177 19.3944
R3827 vdd.n3179 vdd.n3178 19.3944
R3828 vdd.n3179 vdd.n474 19.3944
R3829 vdd.n3183 vdd.n474 19.3944
R3830 vdd.n3184 vdd.n3183 19.3944
R3831 vdd.n3185 vdd.n3184 19.3944
R3832 vdd.n3185 vdd.n471 19.3944
R3833 vdd.n3189 vdd.n471 19.3944
R3834 vdd.n3190 vdd.n3189 19.3944
R3835 vdd.n3191 vdd.n3190 19.3944
R3836 vdd.n3191 vdd.n468 19.3944
R3837 vdd.n3195 vdd.n468 19.3944
R3838 vdd.n3196 vdd.n3195 19.3944
R3839 vdd.n3197 vdd.n3196 19.3944
R3840 vdd.n3240 vdd.n426 19.3944
R3841 vdd.n3240 vdd.n432 19.3944
R3842 vdd.n3235 vdd.n432 19.3944
R3843 vdd.n3235 vdd.n3234 19.3944
R3844 vdd.n3234 vdd.n3233 19.3944
R3845 vdd.n3233 vdd.n439 19.3944
R3846 vdd.n3228 vdd.n439 19.3944
R3847 vdd.n3228 vdd.n3227 19.3944
R3848 vdd.n3227 vdd.n3226 19.3944
R3849 vdd.n3226 vdd.n446 19.3944
R3850 vdd.n3221 vdd.n446 19.3944
R3851 vdd.n3221 vdd.n3220 19.3944
R3852 vdd.n3220 vdd.n3219 19.3944
R3853 vdd.n3219 vdd.n453 19.3944
R3854 vdd.n3214 vdd.n453 19.3944
R3855 vdd.n3214 vdd.n3213 19.3944
R3856 vdd.n3213 vdd.n3212 19.3944
R3857 vdd.n3212 vdd.n460 19.3944
R3858 vdd.n3207 vdd.n460 19.3944
R3859 vdd.n3207 vdd.n3206 19.3944
R3860 vdd.n3279 vdd.n386 19.3944
R3861 vdd.n3279 vdd.n392 19.3944
R3862 vdd.n3274 vdd.n392 19.3944
R3863 vdd.n3274 vdd.n3273 19.3944
R3864 vdd.n3273 vdd.n3272 19.3944
R3865 vdd.n3272 vdd.n399 19.3944
R3866 vdd.n3267 vdd.n399 19.3944
R3867 vdd.n3267 vdd.n3266 19.3944
R3868 vdd.n3266 vdd.n3265 19.3944
R3869 vdd.n3265 vdd.n406 19.3944
R3870 vdd.n3260 vdd.n406 19.3944
R3871 vdd.n3260 vdd.n3259 19.3944
R3872 vdd.n3259 vdd.n3258 19.3944
R3873 vdd.n3258 vdd.n413 19.3944
R3874 vdd.n3253 vdd.n413 19.3944
R3875 vdd.n3253 vdd.n3252 19.3944
R3876 vdd.n3252 vdd.n3251 19.3944
R3877 vdd.n3251 vdd.n420 19.3944
R3878 vdd.n3246 vdd.n420 19.3944
R3879 vdd.n3246 vdd.n3245 19.3944
R3880 vdd.n3315 vdd.n3314 19.3944
R3881 vdd.n3314 vdd.n3313 19.3944
R3882 vdd.n3313 vdd.n358 19.3944
R3883 vdd.n359 vdd.n358 19.3944
R3884 vdd.n3306 vdd.n359 19.3944
R3885 vdd.n3306 vdd.n3305 19.3944
R3886 vdd.n3305 vdd.n3304 19.3944
R3887 vdd.n3304 vdd.n366 19.3944
R3888 vdd.n3299 vdd.n366 19.3944
R3889 vdd.n3299 vdd.n3298 19.3944
R3890 vdd.n3298 vdd.n3297 19.3944
R3891 vdd.n3297 vdd.n373 19.3944
R3892 vdd.n3292 vdd.n373 19.3944
R3893 vdd.n3292 vdd.n3291 19.3944
R3894 vdd.n3291 vdd.n3290 19.3944
R3895 vdd.n3290 vdd.n380 19.3944
R3896 vdd.n3285 vdd.n380 19.3944
R3897 vdd.n3285 vdd.n3284 19.3944
R3898 vdd.n3120 vdd.n509 19.3944
R3899 vdd.n3132 vdd.n509 19.3944
R3900 vdd.n3132 vdd.n507 19.3944
R3901 vdd.n3136 vdd.n507 19.3944
R3902 vdd.n3136 vdd.n497 19.3944
R3903 vdd.n3148 vdd.n497 19.3944
R3904 vdd.n3148 vdd.n495 19.3944
R3905 vdd.n3152 vdd.n495 19.3944
R3906 vdd.n3152 vdd.n485 19.3944
R3907 vdd.n3165 vdd.n485 19.3944
R3908 vdd.n3165 vdd.n483 19.3944
R3909 vdd.n3169 vdd.n483 19.3944
R3910 vdd.n3169 vdd.n312 19.3944
R3911 vdd.n3348 vdd.n312 19.3944
R3912 vdd.n3348 vdd.n313 19.3944
R3913 vdd.n3342 vdd.n313 19.3944
R3914 vdd.n3342 vdd.n3341 19.3944
R3915 vdd.n3341 vdd.n3340 19.3944
R3916 vdd.n3340 vdd.n323 19.3944
R3917 vdd.n3334 vdd.n323 19.3944
R3918 vdd.n3334 vdd.n3333 19.3944
R3919 vdd.n3333 vdd.n3332 19.3944
R3920 vdd.n3332 vdd.n335 19.3944
R3921 vdd.n3326 vdd.n335 19.3944
R3922 vdd.n3326 vdd.n3325 19.3944
R3923 vdd.n3325 vdd.n3324 19.3944
R3924 vdd.n3324 vdd.n346 19.3944
R3925 vdd.n3318 vdd.n346 19.3944
R3926 vdd.n3077 vdd.n3076 19.3944
R3927 vdd.n3076 vdd.n3075 19.3944
R3928 vdd.n3075 vdd.n551 19.3944
R3929 vdd.n3069 vdd.n551 19.3944
R3930 vdd.n3069 vdd.n3068 19.3944
R3931 vdd.n3068 vdd.n3067 19.3944
R3932 vdd.n3067 vdd.n557 19.3944
R3933 vdd.n3061 vdd.n557 19.3944
R3934 vdd.n3061 vdd.n3060 19.3944
R3935 vdd.n3060 vdd.n3059 19.3944
R3936 vdd.n3059 vdd.n563 19.3944
R3937 vdd.n3053 vdd.n563 19.3944
R3938 vdd.n3053 vdd.n3052 19.3944
R3939 vdd.n3052 vdd.n3051 19.3944
R3940 vdd.n3051 vdd.n569 19.3944
R3941 vdd.n3045 vdd.n569 19.3944
R3942 vdd.n3045 vdd.n3044 19.3944
R3943 vdd.n3044 vdd.n3043 19.3944
R3944 vdd.n3043 vdd.n575 19.3944
R3945 vdd.n3037 vdd.n575 19.3944
R3946 vdd.n3117 vdd.n3116 19.3944
R3947 vdd.n3116 vdd.n519 19.3944
R3948 vdd.n3111 vdd.n3110 19.3944
R3949 vdd.n3107 vdd.n3106 19.3944
R3950 vdd.n3106 vdd.n525 19.3944
R3951 vdd.n3101 vdd.n525 19.3944
R3952 vdd.n3101 vdd.n3100 19.3944
R3953 vdd.n3100 vdd.n3099 19.3944
R3954 vdd.n3099 vdd.n531 19.3944
R3955 vdd.n3093 vdd.n531 19.3944
R3956 vdd.n3093 vdd.n3092 19.3944
R3957 vdd.n3092 vdd.n3091 19.3944
R3958 vdd.n3091 vdd.n537 19.3944
R3959 vdd.n3085 vdd.n537 19.3944
R3960 vdd.n3085 vdd.n3084 19.3944
R3961 vdd.n3084 vdd.n3083 19.3944
R3962 vdd.n3032 vdd.n579 19.3944
R3963 vdd.n3032 vdd.n583 19.3944
R3964 vdd.n3027 vdd.n583 19.3944
R3965 vdd.n3027 vdd.n3026 19.3944
R3966 vdd.n3026 vdd.n589 19.3944
R3967 vdd.n3021 vdd.n589 19.3944
R3968 vdd.n3021 vdd.n3020 19.3944
R3969 vdd.n3020 vdd.n3019 19.3944
R3970 vdd.n3019 vdd.n595 19.3944
R3971 vdd.n3013 vdd.n595 19.3944
R3972 vdd.n3013 vdd.n3012 19.3944
R3973 vdd.n3012 vdd.n3011 19.3944
R3974 vdd.n3011 vdd.n601 19.3944
R3975 vdd.n3005 vdd.n601 19.3944
R3976 vdd.n3005 vdd.n3004 19.3944
R3977 vdd.n3004 vdd.n3003 19.3944
R3978 vdd.n2999 vdd.n2998 19.3944
R3979 vdd.n2995 vdd.n2994 19.3944
R3980 vdd.n1229 vdd.n1148 19.0066
R3981 vdd.n1830 vdd.n1761 19.0066
R3982 vdd.n3244 vdd.n426 19.0066
R3983 vdd.n3036 vdd.n579 19.0066
R3984 vdd.n965 vdd.n964 16.0975
R3985 vdd.n826 vdd.n825 16.0975
R3986 vdd.n1191 vdd.n1190 16.0975
R3987 vdd.n1228 vdd.n1227 16.0975
R3988 vdd.n1102 vdd.n1101 16.0975
R3989 vdd.n1913 vdd.n1912 16.0975
R3990 vdd.n1763 vdd.n1762 16.0975
R3991 vdd.n1723 vdd.n1722 16.0975
R3992 vdd.n959 vdd.n958 16.0975
R3993 vdd.n817 vdd.n816 16.0975
R3994 vdd.n2474 vdd.n2473 16.0975
R3995 vdd.n3204 vdd.n3203 16.0975
R3996 vdd.n428 vdd.n427 16.0975
R3997 vdd.n388 vdd.n387 16.0975
R3998 vdd.n581 vdd.n580 16.0975
R3999 vdd.n544 vdd.n543 16.0975
R4000 vdd.n662 vdd.n661 16.0975
R4001 vdd.n2543 vdd.n2542 16.0975
R4002 vdd.n2991 vdd.n2990 16.0975
R4003 vdd.n626 vdd.n625 16.0975
R4004 vdd.t200 vdd.n2438 15.4182
R4005 vdd.n2722 vdd.t187 15.4182
R4006 vdd.n28 vdd.n27 14.5458
R4007 vdd.n2179 vdd.n938 13.6043
R4008 vdd.n2953 vdd.n613 13.6043
R4009 vdd.n304 vdd.n269 13.1884
R4010 vdd.n253 vdd.n218 13.1884
R4011 vdd.n210 vdd.n175 13.1884
R4012 vdd.n159 vdd.n124 13.1884
R4013 vdd.n117 vdd.n82 13.1884
R4014 vdd.n66 vdd.n31 13.1884
R4015 vdd.n1579 vdd.n1544 13.1884
R4016 vdd.n1630 vdd.n1595 13.1884
R4017 vdd.n1485 vdd.n1450 13.1884
R4018 vdd.n1536 vdd.n1501 13.1884
R4019 vdd.n1392 vdd.n1357 13.1884
R4020 vdd.n1443 vdd.n1408 13.1884
R4021 vdd.n1260 vdd.n1103 12.9944
R4022 vdd.n1264 vdd.n1103 12.9944
R4023 vdd.n1869 vdd.n1721 12.9944
R4024 vdd.n1870 vdd.n1869 12.9944
R4025 vdd.n3283 vdd.n386 12.9944
R4026 vdd.n3284 vdd.n3283 12.9944
R4027 vdd.n3077 vdd.n545 12.9944
R4028 vdd.n3083 vdd.n545 12.9944
R4029 vdd.n305 vdd.n267 12.8005
R4030 vdd.n300 vdd.n271 12.8005
R4031 vdd.n254 vdd.n216 12.8005
R4032 vdd.n249 vdd.n220 12.8005
R4033 vdd.n211 vdd.n173 12.8005
R4034 vdd.n206 vdd.n177 12.8005
R4035 vdd.n160 vdd.n122 12.8005
R4036 vdd.n155 vdd.n126 12.8005
R4037 vdd.n118 vdd.n80 12.8005
R4038 vdd.n113 vdd.n84 12.8005
R4039 vdd.n67 vdd.n29 12.8005
R4040 vdd.n62 vdd.n33 12.8005
R4041 vdd.n1580 vdd.n1542 12.8005
R4042 vdd.n1575 vdd.n1546 12.8005
R4043 vdd.n1631 vdd.n1593 12.8005
R4044 vdd.n1626 vdd.n1597 12.8005
R4045 vdd.n1486 vdd.n1448 12.8005
R4046 vdd.n1481 vdd.n1452 12.8005
R4047 vdd.n1537 vdd.n1499 12.8005
R4048 vdd.n1532 vdd.n1503 12.8005
R4049 vdd.n1393 vdd.n1355 12.8005
R4050 vdd.n1388 vdd.n1359 12.8005
R4051 vdd.n1444 vdd.n1406 12.8005
R4052 vdd.n1439 vdd.n1410 12.8005
R4053 vdd.n299 vdd.n272 12.0247
R4054 vdd.n248 vdd.n221 12.0247
R4055 vdd.n205 vdd.n178 12.0247
R4056 vdd.n154 vdd.n127 12.0247
R4057 vdd.n112 vdd.n85 12.0247
R4058 vdd.n61 vdd.n34 12.0247
R4059 vdd.n1574 vdd.n1547 12.0247
R4060 vdd.n1625 vdd.n1598 12.0247
R4061 vdd.n1480 vdd.n1453 12.0247
R4062 vdd.n1531 vdd.n1504 12.0247
R4063 vdd.n1387 vdd.n1360 12.0247
R4064 vdd.n1438 vdd.n1411 12.0247
R4065 vdd.n1295 vdd.n1063 11.337
R4066 vdd.n1303 vdd.n1052 11.337
R4067 vdd.n1311 vdd.n1052 11.337
R4068 vdd.n1319 vdd.n1046 11.337
R4069 vdd.n1327 vdd.n1039 11.337
R4070 vdd.n1336 vdd.n1335 11.337
R4071 vdd.n1344 vdd.n1028 11.337
R4072 vdd.n1642 vdd.n1017 11.337
R4073 vdd.n1651 vdd.n1011 11.337
R4074 vdd.n1659 vdd.n1005 11.337
R4075 vdd.n1668 vdd.n1667 11.337
R4076 vdd.n1676 vdd.n988 11.337
R4077 vdd.n1687 vdd.n988 11.337
R4078 vdd.n1687 vdd.n1686 11.337
R4079 vdd.n3130 vdd.n511 11.337
R4080 vdd.n3130 vdd.n505 11.337
R4081 vdd.n3138 vdd.n505 11.337
R4082 vdd.n3146 vdd.n499 11.337
R4083 vdd.n3154 vdd.n492 11.337
R4084 vdd.n3163 vdd.n3162 11.337
R4085 vdd.n3171 vdd.n481 11.337
R4086 vdd.n3345 vdd.n3344 11.337
R4087 vdd.n3338 vdd.n325 11.337
R4088 vdd.n3336 vdd.n329 11.337
R4089 vdd.n3330 vdd.n3329 11.337
R4090 vdd.n3328 vdd.n340 11.337
R4091 vdd.n3322 vdd.n340 11.337
R4092 vdd.n3321 vdd.n3320 11.337
R4093 vdd.n296 vdd.n295 11.249
R4094 vdd.n245 vdd.n244 11.249
R4095 vdd.n202 vdd.n201 11.249
R4096 vdd.n151 vdd.n150 11.249
R4097 vdd.n109 vdd.n108 11.249
R4098 vdd.n58 vdd.n57 11.249
R4099 vdd.n1571 vdd.n1570 11.249
R4100 vdd.n1622 vdd.n1621 11.249
R4101 vdd.n1477 vdd.n1476 11.249
R4102 vdd.n1528 vdd.n1527 11.249
R4103 vdd.n1384 vdd.n1383 11.249
R4104 vdd.n1435 vdd.n1434 11.249
R4105 vdd.n1311 vdd.t31 10.9969
R4106 vdd.t0 vdd.n3328 10.9969
R4107 vdd.n1040 vdd.t23 10.7702
R4108 vdd.t21 vdd.n3337 10.7702
R4109 vdd.n281 vdd.n280 10.7238
R4110 vdd.n230 vdd.n229 10.7238
R4111 vdd.n187 vdd.n186 10.7238
R4112 vdd.n136 vdd.n135 10.7238
R4113 vdd.n94 vdd.n93 10.7238
R4114 vdd.n43 vdd.n42 10.7238
R4115 vdd.n1556 vdd.n1555 10.7238
R4116 vdd.n1607 vdd.n1606 10.7238
R4117 vdd.n1462 vdd.n1461 10.7238
R4118 vdd.n1513 vdd.n1512 10.7238
R4119 vdd.n1369 vdd.n1368 10.7238
R4120 vdd.n1420 vdd.n1419 10.7238
R4121 vdd.n2177 vdd.n930 10.6151
R4122 vdd.n2187 vdd.n930 10.6151
R4123 vdd.n2188 vdd.n2187 10.6151
R4124 vdd.n2189 vdd.n2188 10.6151
R4125 vdd.n2189 vdd.n918 10.6151
R4126 vdd.n2199 vdd.n918 10.6151
R4127 vdd.n2200 vdd.n2199 10.6151
R4128 vdd.n2201 vdd.n2200 10.6151
R4129 vdd.n2201 vdd.n906 10.6151
R4130 vdd.n2211 vdd.n906 10.6151
R4131 vdd.n2212 vdd.n2211 10.6151
R4132 vdd.n2213 vdd.n2212 10.6151
R4133 vdd.n2213 vdd.n893 10.6151
R4134 vdd.n2223 vdd.n893 10.6151
R4135 vdd.n2224 vdd.n2223 10.6151
R4136 vdd.n2225 vdd.n2224 10.6151
R4137 vdd.n2225 vdd.n881 10.6151
R4138 vdd.n2236 vdd.n881 10.6151
R4139 vdd.n2237 vdd.n2236 10.6151
R4140 vdd.n2238 vdd.n2237 10.6151
R4141 vdd.n2238 vdd.n869 10.6151
R4142 vdd.n2248 vdd.n869 10.6151
R4143 vdd.n2249 vdd.n2248 10.6151
R4144 vdd.n2250 vdd.n2249 10.6151
R4145 vdd.n2250 vdd.n857 10.6151
R4146 vdd.n2260 vdd.n857 10.6151
R4147 vdd.n2261 vdd.n2260 10.6151
R4148 vdd.n2262 vdd.n2261 10.6151
R4149 vdd.n2262 vdd.n847 10.6151
R4150 vdd.n2272 vdd.n847 10.6151
R4151 vdd.n2273 vdd.n2272 10.6151
R4152 vdd.n2274 vdd.n2273 10.6151
R4153 vdd.n2274 vdd.n834 10.6151
R4154 vdd.n2286 vdd.n834 10.6151
R4155 vdd.n2287 vdd.n2286 10.6151
R4156 vdd.n2289 vdd.n2287 10.6151
R4157 vdd.n2289 vdd.n2288 10.6151
R4158 vdd.n2288 vdd.n815 10.6151
R4159 vdd.n2436 vdd.n2435 10.6151
R4160 vdd.n2435 vdd.n2434 10.6151
R4161 vdd.n2434 vdd.n2431 10.6151
R4162 vdd.n2431 vdd.n2430 10.6151
R4163 vdd.n2430 vdd.n2427 10.6151
R4164 vdd.n2427 vdd.n2426 10.6151
R4165 vdd.n2426 vdd.n2423 10.6151
R4166 vdd.n2423 vdd.n2422 10.6151
R4167 vdd.n2422 vdd.n2419 10.6151
R4168 vdd.n2419 vdd.n2418 10.6151
R4169 vdd.n2418 vdd.n2415 10.6151
R4170 vdd.n2415 vdd.n2414 10.6151
R4171 vdd.n2414 vdd.n2411 10.6151
R4172 vdd.n2411 vdd.n2410 10.6151
R4173 vdd.n2410 vdd.n2407 10.6151
R4174 vdd.n2407 vdd.n2406 10.6151
R4175 vdd.n2406 vdd.n2403 10.6151
R4176 vdd.n2403 vdd.n2402 10.6151
R4177 vdd.n2402 vdd.n2399 10.6151
R4178 vdd.n2399 vdd.n2398 10.6151
R4179 vdd.n2398 vdd.n2395 10.6151
R4180 vdd.n2395 vdd.n2394 10.6151
R4181 vdd.n2394 vdd.n2391 10.6151
R4182 vdd.n2391 vdd.n2390 10.6151
R4183 vdd.n2390 vdd.n2387 10.6151
R4184 vdd.n2387 vdd.n2386 10.6151
R4185 vdd.n2386 vdd.n2383 10.6151
R4186 vdd.n2383 vdd.n2382 10.6151
R4187 vdd.n2382 vdd.n2379 10.6151
R4188 vdd.n2379 vdd.n2378 10.6151
R4189 vdd.n2378 vdd.n2375 10.6151
R4190 vdd.n2373 vdd.n2370 10.6151
R4191 vdd.n2370 vdd.n2369 10.6151
R4192 vdd.n2106 vdd.n2105 10.6151
R4193 vdd.n2105 vdd.n2103 10.6151
R4194 vdd.n2103 vdd.n2102 10.6151
R4195 vdd.n2102 vdd.n2100 10.6151
R4196 vdd.n2100 vdd.n2099 10.6151
R4197 vdd.n2099 vdd.n2097 10.6151
R4198 vdd.n2097 vdd.n2096 10.6151
R4199 vdd.n2096 vdd.n2094 10.6151
R4200 vdd.n2094 vdd.n2093 10.6151
R4201 vdd.n2093 vdd.n2091 10.6151
R4202 vdd.n2091 vdd.n2090 10.6151
R4203 vdd.n2090 vdd.n2088 10.6151
R4204 vdd.n2088 vdd.n2087 10.6151
R4205 vdd.n2087 vdd.n2085 10.6151
R4206 vdd.n2085 vdd.n2084 10.6151
R4207 vdd.n2084 vdd.n2082 10.6151
R4208 vdd.n2082 vdd.n2081 10.6151
R4209 vdd.n2081 vdd.n2079 10.6151
R4210 vdd.n2079 vdd.n2078 10.6151
R4211 vdd.n2078 vdd.n2076 10.6151
R4212 vdd.n2076 vdd.n2075 10.6151
R4213 vdd.n2075 vdd.n2073 10.6151
R4214 vdd.n2073 vdd.n2072 10.6151
R4215 vdd.n2072 vdd.n961 10.6151
R4216 vdd.n2039 vdd.n961 10.6151
R4217 vdd.n2040 vdd.n2039 10.6151
R4218 vdd.n2042 vdd.n2040 10.6151
R4219 vdd.n2043 vdd.n2042 10.6151
R4220 vdd.n2056 vdd.n2043 10.6151
R4221 vdd.n2056 vdd.n2055 10.6151
R4222 vdd.n2055 vdd.n2054 10.6151
R4223 vdd.n2054 vdd.n2052 10.6151
R4224 vdd.n2052 vdd.n2051 10.6151
R4225 vdd.n2051 vdd.n2049 10.6151
R4226 vdd.n2049 vdd.n2048 10.6151
R4227 vdd.n2048 vdd.n2045 10.6151
R4228 vdd.n2045 vdd.n2044 10.6151
R4229 vdd.n2044 vdd.n818 10.6151
R4230 vdd.n2176 vdd.n2175 10.6151
R4231 vdd.n2175 vdd.n942 10.6151
R4232 vdd.n2170 vdd.n942 10.6151
R4233 vdd.n2170 vdd.n2169 10.6151
R4234 vdd.n2169 vdd.n944 10.6151
R4235 vdd.n2164 vdd.n944 10.6151
R4236 vdd.n2164 vdd.n2163 10.6151
R4237 vdd.n2163 vdd.n2162 10.6151
R4238 vdd.n2162 vdd.n946 10.6151
R4239 vdd.n2156 vdd.n946 10.6151
R4240 vdd.n2156 vdd.n2155 10.6151
R4241 vdd.n2155 vdd.n2154 10.6151
R4242 vdd.n2154 vdd.n948 10.6151
R4243 vdd.n2148 vdd.n948 10.6151
R4244 vdd.n2148 vdd.n2147 10.6151
R4245 vdd.n2147 vdd.n2146 10.6151
R4246 vdd.n2146 vdd.n950 10.6151
R4247 vdd.n2140 vdd.n950 10.6151
R4248 vdd.n2140 vdd.n2139 10.6151
R4249 vdd.n2139 vdd.n2138 10.6151
R4250 vdd.n2138 vdd.n952 10.6151
R4251 vdd.n2132 vdd.n952 10.6151
R4252 vdd.n2132 vdd.n2131 10.6151
R4253 vdd.n2131 vdd.n2130 10.6151
R4254 vdd.n2130 vdd.n954 10.6151
R4255 vdd.n2124 vdd.n954 10.6151
R4256 vdd.n2124 vdd.n2123 10.6151
R4257 vdd.n2123 vdd.n2122 10.6151
R4258 vdd.n2122 vdd.n956 10.6151
R4259 vdd.n2116 vdd.n956 10.6151
R4260 vdd.n2116 vdd.n2115 10.6151
R4261 vdd.n2113 vdd.n960 10.6151
R4262 vdd.n2107 vdd.n960 10.6151
R4263 vdd.n2611 vdd.n2609 10.6151
R4264 vdd.n2612 vdd.n2611 10.6151
R4265 vdd.n2711 vdd.n2612 10.6151
R4266 vdd.n2711 vdd.n2710 10.6151
R4267 vdd.n2710 vdd.n2709 10.6151
R4268 vdd.n2709 vdd.n2707 10.6151
R4269 vdd.n2707 vdd.n2706 10.6151
R4270 vdd.n2706 vdd.n2704 10.6151
R4271 vdd.n2704 vdd.n2703 10.6151
R4272 vdd.n2703 vdd.n2613 10.6151
R4273 vdd.n2653 vdd.n2613 10.6151
R4274 vdd.n2654 vdd.n2653 10.6151
R4275 vdd.n2656 vdd.n2654 10.6151
R4276 vdd.n2657 vdd.n2656 10.6151
R4277 vdd.n2687 vdd.n2657 10.6151
R4278 vdd.n2687 vdd.n2686 10.6151
R4279 vdd.n2686 vdd.n2685 10.6151
R4280 vdd.n2685 vdd.n2683 10.6151
R4281 vdd.n2683 vdd.n2682 10.6151
R4282 vdd.n2682 vdd.n2680 10.6151
R4283 vdd.n2680 vdd.n2679 10.6151
R4284 vdd.n2679 vdd.n2677 10.6151
R4285 vdd.n2677 vdd.n2676 10.6151
R4286 vdd.n2676 vdd.n2674 10.6151
R4287 vdd.n2674 vdd.n2673 10.6151
R4288 vdd.n2673 vdd.n2671 10.6151
R4289 vdd.n2671 vdd.n2670 10.6151
R4290 vdd.n2670 vdd.n2668 10.6151
R4291 vdd.n2668 vdd.n2667 10.6151
R4292 vdd.n2667 vdd.n2665 10.6151
R4293 vdd.n2665 vdd.n2664 10.6151
R4294 vdd.n2664 vdd.n2662 10.6151
R4295 vdd.n2662 vdd.n2661 10.6151
R4296 vdd.n2661 vdd.n2659 10.6151
R4297 vdd.n2659 vdd.n2658 10.6151
R4298 vdd.n2658 vdd.n664 10.6151
R4299 vdd.n2886 vdd.n664 10.6151
R4300 vdd.n2887 vdd.n2886 10.6151
R4301 vdd.n2726 vdd.n2725 10.6151
R4302 vdd.n2725 vdd.n776 10.6151
R4303 vdd.n2545 vdd.n776 10.6151
R4304 vdd.n2546 vdd.n2545 10.6151
R4305 vdd.n2549 vdd.n2546 10.6151
R4306 vdd.n2550 vdd.n2549 10.6151
R4307 vdd.n2553 vdd.n2550 10.6151
R4308 vdd.n2554 vdd.n2553 10.6151
R4309 vdd.n2557 vdd.n2554 10.6151
R4310 vdd.n2558 vdd.n2557 10.6151
R4311 vdd.n2561 vdd.n2558 10.6151
R4312 vdd.n2562 vdd.n2561 10.6151
R4313 vdd.n2565 vdd.n2562 10.6151
R4314 vdd.n2566 vdd.n2565 10.6151
R4315 vdd.n2569 vdd.n2566 10.6151
R4316 vdd.n2570 vdd.n2569 10.6151
R4317 vdd.n2573 vdd.n2570 10.6151
R4318 vdd.n2574 vdd.n2573 10.6151
R4319 vdd.n2577 vdd.n2574 10.6151
R4320 vdd.n2578 vdd.n2577 10.6151
R4321 vdd.n2581 vdd.n2578 10.6151
R4322 vdd.n2582 vdd.n2581 10.6151
R4323 vdd.n2585 vdd.n2582 10.6151
R4324 vdd.n2586 vdd.n2585 10.6151
R4325 vdd.n2589 vdd.n2586 10.6151
R4326 vdd.n2590 vdd.n2589 10.6151
R4327 vdd.n2593 vdd.n2590 10.6151
R4328 vdd.n2594 vdd.n2593 10.6151
R4329 vdd.n2597 vdd.n2594 10.6151
R4330 vdd.n2598 vdd.n2597 10.6151
R4331 vdd.n2601 vdd.n2598 10.6151
R4332 vdd.n2606 vdd.n2603 10.6151
R4333 vdd.n2608 vdd.n2606 10.6151
R4334 vdd.n2727 vdd.n765 10.6151
R4335 vdd.n2737 vdd.n765 10.6151
R4336 vdd.n2738 vdd.n2737 10.6151
R4337 vdd.n2739 vdd.n2738 10.6151
R4338 vdd.n2739 vdd.n753 10.6151
R4339 vdd.n2749 vdd.n753 10.6151
R4340 vdd.n2750 vdd.n2749 10.6151
R4341 vdd.n2751 vdd.n2750 10.6151
R4342 vdd.n2751 vdd.n743 10.6151
R4343 vdd.n2761 vdd.n743 10.6151
R4344 vdd.n2762 vdd.n2761 10.6151
R4345 vdd.n2763 vdd.n2762 10.6151
R4346 vdd.n2763 vdd.n731 10.6151
R4347 vdd.n2773 vdd.n731 10.6151
R4348 vdd.n2774 vdd.n2773 10.6151
R4349 vdd.n2775 vdd.n2774 10.6151
R4350 vdd.n2775 vdd.n720 10.6151
R4351 vdd.n2785 vdd.n720 10.6151
R4352 vdd.n2786 vdd.n2785 10.6151
R4353 vdd.n2787 vdd.n2786 10.6151
R4354 vdd.n2787 vdd.n707 10.6151
R4355 vdd.n2798 vdd.n707 10.6151
R4356 vdd.n2799 vdd.n2798 10.6151
R4357 vdd.n2800 vdd.n2799 10.6151
R4358 vdd.n2800 vdd.n694 10.6151
R4359 vdd.n2810 vdd.n694 10.6151
R4360 vdd.n2811 vdd.n2810 10.6151
R4361 vdd.n2812 vdd.n2811 10.6151
R4362 vdd.n2812 vdd.n683 10.6151
R4363 vdd.n2822 vdd.n683 10.6151
R4364 vdd.n2823 vdd.n2822 10.6151
R4365 vdd.n2824 vdd.n2823 10.6151
R4366 vdd.n2824 vdd.n669 10.6151
R4367 vdd.n2879 vdd.n669 10.6151
R4368 vdd.n2880 vdd.n2879 10.6151
R4369 vdd.n2881 vdd.n2880 10.6151
R4370 vdd.n2881 vdd.n636 10.6151
R4371 vdd.n2951 vdd.n636 10.6151
R4372 vdd.n2950 vdd.n2949 10.6151
R4373 vdd.n2949 vdd.n637 10.6151
R4374 vdd.n638 vdd.n637 10.6151
R4375 vdd.n2942 vdd.n638 10.6151
R4376 vdd.n2942 vdd.n2941 10.6151
R4377 vdd.n2941 vdd.n2940 10.6151
R4378 vdd.n2940 vdd.n640 10.6151
R4379 vdd.n2935 vdd.n640 10.6151
R4380 vdd.n2935 vdd.n2934 10.6151
R4381 vdd.n2934 vdd.n2933 10.6151
R4382 vdd.n2933 vdd.n643 10.6151
R4383 vdd.n2928 vdd.n643 10.6151
R4384 vdd.n2928 vdd.n2927 10.6151
R4385 vdd.n2927 vdd.n2926 10.6151
R4386 vdd.n2926 vdd.n646 10.6151
R4387 vdd.n2921 vdd.n646 10.6151
R4388 vdd.n2921 vdd.n2920 10.6151
R4389 vdd.n2920 vdd.n2918 10.6151
R4390 vdd.n2918 vdd.n649 10.6151
R4391 vdd.n2913 vdd.n649 10.6151
R4392 vdd.n2913 vdd.n2912 10.6151
R4393 vdd.n2912 vdd.n2911 10.6151
R4394 vdd.n2911 vdd.n652 10.6151
R4395 vdd.n2906 vdd.n652 10.6151
R4396 vdd.n2906 vdd.n2905 10.6151
R4397 vdd.n2905 vdd.n2904 10.6151
R4398 vdd.n2904 vdd.n655 10.6151
R4399 vdd.n2899 vdd.n655 10.6151
R4400 vdd.n2899 vdd.n2898 10.6151
R4401 vdd.n2898 vdd.n2897 10.6151
R4402 vdd.n2897 vdd.n658 10.6151
R4403 vdd.n2892 vdd.n2891 10.6151
R4404 vdd.n2891 vdd.n2890 10.6151
R4405 vdd.n2869 vdd.n2830 10.6151
R4406 vdd.n2864 vdd.n2830 10.6151
R4407 vdd.n2864 vdd.n2863 10.6151
R4408 vdd.n2863 vdd.n2862 10.6151
R4409 vdd.n2862 vdd.n2832 10.6151
R4410 vdd.n2857 vdd.n2832 10.6151
R4411 vdd.n2857 vdd.n2856 10.6151
R4412 vdd.n2856 vdd.n2855 10.6151
R4413 vdd.n2855 vdd.n2835 10.6151
R4414 vdd.n2850 vdd.n2835 10.6151
R4415 vdd.n2850 vdd.n2849 10.6151
R4416 vdd.n2849 vdd.n2848 10.6151
R4417 vdd.n2848 vdd.n2838 10.6151
R4418 vdd.n2843 vdd.n2838 10.6151
R4419 vdd.n2843 vdd.n2842 10.6151
R4420 vdd.n2842 vdd.n610 10.6151
R4421 vdd.n2986 vdd.n610 10.6151
R4422 vdd.n2986 vdd.n611 10.6151
R4423 vdd.n614 vdd.n611 10.6151
R4424 vdd.n2979 vdd.n614 10.6151
R4425 vdd.n2979 vdd.n2978 10.6151
R4426 vdd.n2978 vdd.n2977 10.6151
R4427 vdd.n2977 vdd.n616 10.6151
R4428 vdd.n2972 vdd.n616 10.6151
R4429 vdd.n2972 vdd.n2971 10.6151
R4430 vdd.n2971 vdd.n2970 10.6151
R4431 vdd.n2970 vdd.n619 10.6151
R4432 vdd.n2965 vdd.n619 10.6151
R4433 vdd.n2965 vdd.n2964 10.6151
R4434 vdd.n2964 vdd.n2963 10.6151
R4435 vdd.n2963 vdd.n622 10.6151
R4436 vdd.n2958 vdd.n2957 10.6151
R4437 vdd.n2957 vdd.n2956 10.6151
R4438 vdd.n2719 vdd.n2718 10.6151
R4439 vdd.n2718 vdd.n2716 10.6151
R4440 vdd.n2716 vdd.n2715 10.6151
R4441 vdd.n2715 vdd.n2541 10.6151
R4442 vdd.n2615 vdd.n2541 10.6151
R4443 vdd.n2616 vdd.n2615 10.6151
R4444 vdd.n2618 vdd.n2616 10.6151
R4445 vdd.n2619 vdd.n2618 10.6151
R4446 vdd.n2699 vdd.n2619 10.6151
R4447 vdd.n2699 vdd.n2698 10.6151
R4448 vdd.n2698 vdd.n2697 10.6151
R4449 vdd.n2697 vdd.n2695 10.6151
R4450 vdd.n2695 vdd.n2694 10.6151
R4451 vdd.n2694 vdd.n2692 10.6151
R4452 vdd.n2692 vdd.n2691 10.6151
R4453 vdd.n2691 vdd.n2651 10.6151
R4454 vdd.n2651 vdd.n2650 10.6151
R4455 vdd.n2650 vdd.n2648 10.6151
R4456 vdd.n2648 vdd.n2647 10.6151
R4457 vdd.n2647 vdd.n2645 10.6151
R4458 vdd.n2645 vdd.n2644 10.6151
R4459 vdd.n2644 vdd.n2642 10.6151
R4460 vdd.n2642 vdd.n2641 10.6151
R4461 vdd.n2641 vdd.n2639 10.6151
R4462 vdd.n2639 vdd.n2638 10.6151
R4463 vdd.n2638 vdd.n2636 10.6151
R4464 vdd.n2636 vdd.n2635 10.6151
R4465 vdd.n2635 vdd.n2633 10.6151
R4466 vdd.n2633 vdd.n2632 10.6151
R4467 vdd.n2632 vdd.n2630 10.6151
R4468 vdd.n2630 vdd.n2629 10.6151
R4469 vdd.n2629 vdd.n2627 10.6151
R4470 vdd.n2627 vdd.n2626 10.6151
R4471 vdd.n2626 vdd.n2624 10.6151
R4472 vdd.n2624 vdd.n2623 10.6151
R4473 vdd.n2623 vdd.n2621 10.6151
R4474 vdd.n2621 vdd.n2620 10.6151
R4475 vdd.n2620 vdd.n628 10.6151
R4476 vdd.n2476 vdd.n770 10.6151
R4477 vdd.n2479 vdd.n2476 10.6151
R4478 vdd.n2480 vdd.n2479 10.6151
R4479 vdd.n2483 vdd.n2480 10.6151
R4480 vdd.n2484 vdd.n2483 10.6151
R4481 vdd.n2487 vdd.n2484 10.6151
R4482 vdd.n2488 vdd.n2487 10.6151
R4483 vdd.n2491 vdd.n2488 10.6151
R4484 vdd.n2492 vdd.n2491 10.6151
R4485 vdd.n2495 vdd.n2492 10.6151
R4486 vdd.n2496 vdd.n2495 10.6151
R4487 vdd.n2499 vdd.n2496 10.6151
R4488 vdd.n2500 vdd.n2499 10.6151
R4489 vdd.n2503 vdd.n2500 10.6151
R4490 vdd.n2504 vdd.n2503 10.6151
R4491 vdd.n2507 vdd.n2504 10.6151
R4492 vdd.n2508 vdd.n2507 10.6151
R4493 vdd.n2511 vdd.n2508 10.6151
R4494 vdd.n2512 vdd.n2511 10.6151
R4495 vdd.n2515 vdd.n2512 10.6151
R4496 vdd.n2516 vdd.n2515 10.6151
R4497 vdd.n2519 vdd.n2516 10.6151
R4498 vdd.n2520 vdd.n2519 10.6151
R4499 vdd.n2523 vdd.n2520 10.6151
R4500 vdd.n2524 vdd.n2523 10.6151
R4501 vdd.n2527 vdd.n2524 10.6151
R4502 vdd.n2528 vdd.n2527 10.6151
R4503 vdd.n2531 vdd.n2528 10.6151
R4504 vdd.n2532 vdd.n2531 10.6151
R4505 vdd.n2535 vdd.n2532 10.6151
R4506 vdd.n2536 vdd.n2535 10.6151
R4507 vdd.n2540 vdd.n2539 10.6151
R4508 vdd.n2720 vdd.n2540 10.6151
R4509 vdd.n2732 vdd.n2731 10.6151
R4510 vdd.n2733 vdd.n2732 10.6151
R4511 vdd.n2733 vdd.n760 10.6151
R4512 vdd.n2743 vdd.n760 10.6151
R4513 vdd.n2744 vdd.n2743 10.6151
R4514 vdd.n2745 vdd.n2744 10.6151
R4515 vdd.n2745 vdd.n748 10.6151
R4516 vdd.n2755 vdd.n748 10.6151
R4517 vdd.n2756 vdd.n2755 10.6151
R4518 vdd.n2757 vdd.n2756 10.6151
R4519 vdd.n2757 vdd.n737 10.6151
R4520 vdd.n2767 vdd.n737 10.6151
R4521 vdd.n2768 vdd.n2767 10.6151
R4522 vdd.n2769 vdd.n2768 10.6151
R4523 vdd.n2769 vdd.n725 10.6151
R4524 vdd.n2779 vdd.n725 10.6151
R4525 vdd.n2780 vdd.n2779 10.6151
R4526 vdd.n2781 vdd.n2780 10.6151
R4527 vdd.n2781 vdd.n714 10.6151
R4528 vdd.n2791 vdd.n714 10.6151
R4529 vdd.n2794 vdd.n2793 10.6151
R4530 vdd.n2794 vdd.n700 10.6151
R4531 vdd.n2804 vdd.n700 10.6151
R4532 vdd.n2805 vdd.n2804 10.6151
R4533 vdd.n2806 vdd.n2805 10.6151
R4534 vdd.n2806 vdd.n688 10.6151
R4535 vdd.n2816 vdd.n688 10.6151
R4536 vdd.n2817 vdd.n2816 10.6151
R4537 vdd.n2818 vdd.n2817 10.6151
R4538 vdd.n2818 vdd.n677 10.6151
R4539 vdd.n2828 vdd.n677 10.6151
R4540 vdd.n2829 vdd.n2828 10.6151
R4541 vdd.n2875 vdd.n2829 10.6151
R4542 vdd.n2875 vdd.n2874 10.6151
R4543 vdd.n2874 vdd.n2873 10.6151
R4544 vdd.n2873 vdd.n2872 10.6151
R4545 vdd.n2872 vdd.n2870 10.6151
R4546 vdd.n2182 vdd.n2181 10.6151
R4547 vdd.n2183 vdd.n2182 10.6151
R4548 vdd.n2183 vdd.n924 10.6151
R4549 vdd.n2193 vdd.n924 10.6151
R4550 vdd.n2194 vdd.n2193 10.6151
R4551 vdd.n2195 vdd.n2194 10.6151
R4552 vdd.n2195 vdd.n912 10.6151
R4553 vdd.n2205 vdd.n912 10.6151
R4554 vdd.n2206 vdd.n2205 10.6151
R4555 vdd.n2207 vdd.n2206 10.6151
R4556 vdd.n2207 vdd.n900 10.6151
R4557 vdd.n2217 vdd.n900 10.6151
R4558 vdd.n2218 vdd.n2217 10.6151
R4559 vdd.n2219 vdd.n2218 10.6151
R4560 vdd.n2219 vdd.n887 10.6151
R4561 vdd.n2229 vdd.n887 10.6151
R4562 vdd.n2230 vdd.n2229 10.6151
R4563 vdd.n2232 vdd.n875 10.6151
R4564 vdd.n2242 vdd.n875 10.6151
R4565 vdd.n2243 vdd.n2242 10.6151
R4566 vdd.n2244 vdd.n2243 10.6151
R4567 vdd.n2244 vdd.n863 10.6151
R4568 vdd.n2254 vdd.n863 10.6151
R4569 vdd.n2255 vdd.n2254 10.6151
R4570 vdd.n2256 vdd.n2255 10.6151
R4571 vdd.n2256 vdd.n852 10.6151
R4572 vdd.n2266 vdd.n852 10.6151
R4573 vdd.n2267 vdd.n2266 10.6151
R4574 vdd.n2268 vdd.n2267 10.6151
R4575 vdd.n2268 vdd.n841 10.6151
R4576 vdd.n2278 vdd.n841 10.6151
R4577 vdd.n2279 vdd.n2278 10.6151
R4578 vdd.n2282 vdd.n2279 10.6151
R4579 vdd.n2282 vdd.n2281 10.6151
R4580 vdd.n2281 vdd.n2280 10.6151
R4581 vdd.n2280 vdd.n824 10.6151
R4582 vdd.n2364 vdd.n824 10.6151
R4583 vdd.n2363 vdd.n2362 10.6151
R4584 vdd.n2362 vdd.n2359 10.6151
R4585 vdd.n2359 vdd.n2358 10.6151
R4586 vdd.n2358 vdd.n2355 10.6151
R4587 vdd.n2355 vdd.n2354 10.6151
R4588 vdd.n2354 vdd.n2351 10.6151
R4589 vdd.n2351 vdd.n2350 10.6151
R4590 vdd.n2350 vdd.n2347 10.6151
R4591 vdd.n2347 vdd.n2346 10.6151
R4592 vdd.n2346 vdd.n2343 10.6151
R4593 vdd.n2343 vdd.n2342 10.6151
R4594 vdd.n2342 vdd.n2339 10.6151
R4595 vdd.n2339 vdd.n2338 10.6151
R4596 vdd.n2338 vdd.n2335 10.6151
R4597 vdd.n2335 vdd.n2334 10.6151
R4598 vdd.n2334 vdd.n2331 10.6151
R4599 vdd.n2331 vdd.n2330 10.6151
R4600 vdd.n2330 vdd.n2327 10.6151
R4601 vdd.n2327 vdd.n2326 10.6151
R4602 vdd.n2326 vdd.n2323 10.6151
R4603 vdd.n2323 vdd.n2322 10.6151
R4604 vdd.n2322 vdd.n2319 10.6151
R4605 vdd.n2319 vdd.n2318 10.6151
R4606 vdd.n2318 vdd.n2315 10.6151
R4607 vdd.n2315 vdd.n2314 10.6151
R4608 vdd.n2314 vdd.n2311 10.6151
R4609 vdd.n2311 vdd.n2310 10.6151
R4610 vdd.n2310 vdd.n2307 10.6151
R4611 vdd.n2307 vdd.n2306 10.6151
R4612 vdd.n2306 vdd.n2303 10.6151
R4613 vdd.n2303 vdd.n2302 10.6151
R4614 vdd.n2299 vdd.n2298 10.6151
R4615 vdd.n2298 vdd.n2296 10.6151
R4616 vdd.n1998 vdd.n1996 10.6151
R4617 vdd.n1999 vdd.n1998 10.6151
R4618 vdd.n2001 vdd.n1999 10.6151
R4619 vdd.n2002 vdd.n2001 10.6151
R4620 vdd.n2004 vdd.n2002 10.6151
R4621 vdd.n2005 vdd.n2004 10.6151
R4622 vdd.n2007 vdd.n2005 10.6151
R4623 vdd.n2008 vdd.n2007 10.6151
R4624 vdd.n2010 vdd.n2008 10.6151
R4625 vdd.n2011 vdd.n2010 10.6151
R4626 vdd.n2013 vdd.n2011 10.6151
R4627 vdd.n2014 vdd.n2013 10.6151
R4628 vdd.n2016 vdd.n2014 10.6151
R4629 vdd.n2017 vdd.n2016 10.6151
R4630 vdd.n2019 vdd.n2017 10.6151
R4631 vdd.n2020 vdd.n2019 10.6151
R4632 vdd.n2022 vdd.n2020 10.6151
R4633 vdd.n2023 vdd.n2022 10.6151
R4634 vdd.n2025 vdd.n2023 10.6151
R4635 vdd.n2026 vdd.n2025 10.6151
R4636 vdd.n2028 vdd.n2026 10.6151
R4637 vdd.n2029 vdd.n2028 10.6151
R4638 vdd.n2068 vdd.n2029 10.6151
R4639 vdd.n2068 vdd.n2067 10.6151
R4640 vdd.n2067 vdd.n2066 10.6151
R4641 vdd.n2066 vdd.n2064 10.6151
R4642 vdd.n2064 vdd.n2063 10.6151
R4643 vdd.n2063 vdd.n2061 10.6151
R4644 vdd.n2061 vdd.n2060 10.6151
R4645 vdd.n2060 vdd.n2037 10.6151
R4646 vdd.n2037 vdd.n2036 10.6151
R4647 vdd.n2036 vdd.n2034 10.6151
R4648 vdd.n2034 vdd.n2033 10.6151
R4649 vdd.n2033 vdd.n2031 10.6151
R4650 vdd.n2031 vdd.n2030 10.6151
R4651 vdd.n2030 vdd.n828 10.6151
R4652 vdd.n2294 vdd.n828 10.6151
R4653 vdd.n2295 vdd.n2294 10.6151
R4654 vdd.n1926 vdd.n936 10.6151
R4655 vdd.n1931 vdd.n1926 10.6151
R4656 vdd.n1932 vdd.n1931 10.6151
R4657 vdd.n1933 vdd.n1932 10.6151
R4658 vdd.n1933 vdd.n1924 10.6151
R4659 vdd.n1939 vdd.n1924 10.6151
R4660 vdd.n1940 vdd.n1939 10.6151
R4661 vdd.n1941 vdd.n1940 10.6151
R4662 vdd.n1941 vdd.n1922 10.6151
R4663 vdd.n1947 vdd.n1922 10.6151
R4664 vdd.n1948 vdd.n1947 10.6151
R4665 vdd.n1949 vdd.n1948 10.6151
R4666 vdd.n1949 vdd.n1920 10.6151
R4667 vdd.n1955 vdd.n1920 10.6151
R4668 vdd.n1956 vdd.n1955 10.6151
R4669 vdd.n1957 vdd.n1956 10.6151
R4670 vdd.n1957 vdd.n1918 10.6151
R4671 vdd.n1963 vdd.n1918 10.6151
R4672 vdd.n1964 vdd.n1963 10.6151
R4673 vdd.n1965 vdd.n1964 10.6151
R4674 vdd.n1965 vdd.n970 10.6151
R4675 vdd.n1971 vdd.n970 10.6151
R4676 vdd.n1972 vdd.n1971 10.6151
R4677 vdd.n1973 vdd.n1972 10.6151
R4678 vdd.n1973 vdd.n968 10.6151
R4679 vdd.n1979 vdd.n968 10.6151
R4680 vdd.n1980 vdd.n1979 10.6151
R4681 vdd.n1981 vdd.n1980 10.6151
R4682 vdd.n1981 vdd.n966 10.6151
R4683 vdd.n1987 vdd.n966 10.6151
R4684 vdd.n1988 vdd.n1987 10.6151
R4685 vdd.n1990 vdd.n962 10.6151
R4686 vdd.n1995 vdd.n962 10.6151
R4687 vdd.n1352 vdd.t6 10.5435
R4688 vdd.n1908 vdd.t117 10.5435
R4689 vdd.n3122 vdd.t95 10.5435
R4690 vdd.n3346 vdd.t35 10.5435
R4691 vdd.n292 vdd.n274 10.4732
R4692 vdd.n241 vdd.n223 10.4732
R4693 vdd.n198 vdd.n180 10.4732
R4694 vdd.n147 vdd.n129 10.4732
R4695 vdd.n105 vdd.n87 10.4732
R4696 vdd.n54 vdd.n36 10.4732
R4697 vdd.n1567 vdd.n1549 10.4732
R4698 vdd.n1618 vdd.n1600 10.4732
R4699 vdd.n1473 vdd.n1455 10.4732
R4700 vdd.n1524 vdd.n1506 10.4732
R4701 vdd.n1380 vdd.n1362 10.4732
R4702 vdd.n1431 vdd.n1413 10.4732
R4703 vdd.n1650 vdd.t16 10.3167
R4704 vdd.t82 vdd.n493 10.3167
R4705 vdd.n2366 vdd.t220 10.2034
R4706 vdd.n2729 vdd.t204 10.2034
R4707 vdd.n1894 vdd.n950 9.88581
R4708 vdd.n2920 vdd.n2919 9.88581
R4709 vdd.n2987 vdd.n2986 9.88581
R4710 vdd.n1918 vdd.n1917 9.88581
R4711 vdd.n1303 vdd.t121 9.86327
R4712 vdd.n3322 vdd.t125 9.86327
R4713 vdd.n291 vdd.n276 9.69747
R4714 vdd.n240 vdd.n225 9.69747
R4715 vdd.n197 vdd.n182 9.69747
R4716 vdd.n146 vdd.n131 9.69747
R4717 vdd.n104 vdd.n89 9.69747
R4718 vdd.n53 vdd.n38 9.69747
R4719 vdd.n1566 vdd.n1551 9.69747
R4720 vdd.n1617 vdd.n1602 9.69747
R4721 vdd.n1472 vdd.n1457 9.69747
R4722 vdd.n1523 vdd.n1508 9.69747
R4723 vdd.n1379 vdd.n1364 9.69747
R4724 vdd.n1430 vdd.n1415 9.69747
R4725 vdd.n307 vdd.n306 9.45567
R4726 vdd.n256 vdd.n255 9.45567
R4727 vdd.n213 vdd.n212 9.45567
R4728 vdd.n162 vdd.n161 9.45567
R4729 vdd.n120 vdd.n119 9.45567
R4730 vdd.n69 vdd.n68 9.45567
R4731 vdd.n1582 vdd.n1581 9.45567
R4732 vdd.n1633 vdd.n1632 9.45567
R4733 vdd.n1488 vdd.n1487 9.45567
R4734 vdd.n1539 vdd.n1538 9.45567
R4735 vdd.n1395 vdd.n1394 9.45567
R4736 vdd.n1446 vdd.n1445 9.45567
R4737 vdd.n1867 vdd.n1721 9.3005
R4738 vdd.n1866 vdd.n1865 9.3005
R4739 vdd.n1727 vdd.n1726 9.3005
R4740 vdd.n1860 vdd.n1731 9.3005
R4741 vdd.n1859 vdd.n1732 9.3005
R4742 vdd.n1858 vdd.n1733 9.3005
R4743 vdd.n1737 vdd.n1734 9.3005
R4744 vdd.n1853 vdd.n1738 9.3005
R4745 vdd.n1852 vdd.n1739 9.3005
R4746 vdd.n1851 vdd.n1740 9.3005
R4747 vdd.n1744 vdd.n1741 9.3005
R4748 vdd.n1846 vdd.n1745 9.3005
R4749 vdd.n1845 vdd.n1746 9.3005
R4750 vdd.n1844 vdd.n1747 9.3005
R4751 vdd.n1751 vdd.n1748 9.3005
R4752 vdd.n1839 vdd.n1752 9.3005
R4753 vdd.n1838 vdd.n1753 9.3005
R4754 vdd.n1837 vdd.n1754 9.3005
R4755 vdd.n1758 vdd.n1755 9.3005
R4756 vdd.n1832 vdd.n1759 9.3005
R4757 vdd.n1831 vdd.n1760 9.3005
R4758 vdd.n1830 vdd.n1829 9.3005
R4759 vdd.n1828 vdd.n1761 9.3005
R4760 vdd.n1827 vdd.n1826 9.3005
R4761 vdd.n1767 vdd.n1766 9.3005
R4762 vdd.n1821 vdd.n1771 9.3005
R4763 vdd.n1820 vdd.n1772 9.3005
R4764 vdd.n1819 vdd.n1773 9.3005
R4765 vdd.n1777 vdd.n1774 9.3005
R4766 vdd.n1814 vdd.n1778 9.3005
R4767 vdd.n1813 vdd.n1779 9.3005
R4768 vdd.n1812 vdd.n1780 9.3005
R4769 vdd.n1784 vdd.n1781 9.3005
R4770 vdd.n1807 vdd.n1785 9.3005
R4771 vdd.n1806 vdd.n1786 9.3005
R4772 vdd.n1805 vdd.n1787 9.3005
R4773 vdd.n1789 vdd.n1788 9.3005
R4774 vdd.n1800 vdd.n972 9.3005
R4775 vdd.n1869 vdd.n1868 9.3005
R4776 vdd.n1893 vdd.n1892 9.3005
R4777 vdd.n1699 vdd.n1698 9.3005
R4778 vdd.n1704 vdd.n1702 9.3005
R4779 vdd.n1885 vdd.n1705 9.3005
R4780 vdd.n1884 vdd.n1706 9.3005
R4781 vdd.n1883 vdd.n1707 9.3005
R4782 vdd.n1711 vdd.n1708 9.3005
R4783 vdd.n1878 vdd.n1712 9.3005
R4784 vdd.n1877 vdd.n1713 9.3005
R4785 vdd.n1876 vdd.n1714 9.3005
R4786 vdd.n1718 vdd.n1715 9.3005
R4787 vdd.n1871 vdd.n1719 9.3005
R4788 vdd.n1870 vdd.n1720 9.3005
R4789 vdd.n1902 vdd.n1692 9.3005
R4790 vdd.n1904 vdd.n1903 9.3005
R4791 vdd.n1638 vdd.n1019 9.3005
R4792 vdd.n1640 vdd.n1639 9.3005
R4793 vdd.n1009 vdd.n1008 9.3005
R4794 vdd.n1654 vdd.n1653 9.3005
R4795 vdd.n1655 vdd.n1007 9.3005
R4796 vdd.n1657 vdd.n1656 9.3005
R4797 vdd.n998 vdd.n997 9.3005
R4798 vdd.n1671 vdd.n1670 9.3005
R4799 vdd.n1672 vdd.n996 9.3005
R4800 vdd.n1674 vdd.n1673 9.3005
R4801 vdd.n986 vdd.n985 9.3005
R4802 vdd.n1690 vdd.n1689 9.3005
R4803 vdd.n1691 vdd.n984 9.3005
R4804 vdd.n1906 vdd.n1905 9.3005
R4805 vdd.n283 vdd.n282 9.3005
R4806 vdd.n278 vdd.n277 9.3005
R4807 vdd.n289 vdd.n288 9.3005
R4808 vdd.n291 vdd.n290 9.3005
R4809 vdd.n274 vdd.n273 9.3005
R4810 vdd.n297 vdd.n296 9.3005
R4811 vdd.n299 vdd.n298 9.3005
R4812 vdd.n271 vdd.n268 9.3005
R4813 vdd.n306 vdd.n305 9.3005
R4814 vdd.n232 vdd.n231 9.3005
R4815 vdd.n227 vdd.n226 9.3005
R4816 vdd.n238 vdd.n237 9.3005
R4817 vdd.n240 vdd.n239 9.3005
R4818 vdd.n223 vdd.n222 9.3005
R4819 vdd.n246 vdd.n245 9.3005
R4820 vdd.n248 vdd.n247 9.3005
R4821 vdd.n220 vdd.n217 9.3005
R4822 vdd.n255 vdd.n254 9.3005
R4823 vdd.n189 vdd.n188 9.3005
R4824 vdd.n184 vdd.n183 9.3005
R4825 vdd.n195 vdd.n194 9.3005
R4826 vdd.n197 vdd.n196 9.3005
R4827 vdd.n180 vdd.n179 9.3005
R4828 vdd.n203 vdd.n202 9.3005
R4829 vdd.n205 vdd.n204 9.3005
R4830 vdd.n177 vdd.n174 9.3005
R4831 vdd.n212 vdd.n211 9.3005
R4832 vdd.n138 vdd.n137 9.3005
R4833 vdd.n133 vdd.n132 9.3005
R4834 vdd.n144 vdd.n143 9.3005
R4835 vdd.n146 vdd.n145 9.3005
R4836 vdd.n129 vdd.n128 9.3005
R4837 vdd.n152 vdd.n151 9.3005
R4838 vdd.n154 vdd.n153 9.3005
R4839 vdd.n126 vdd.n123 9.3005
R4840 vdd.n161 vdd.n160 9.3005
R4841 vdd.n96 vdd.n95 9.3005
R4842 vdd.n91 vdd.n90 9.3005
R4843 vdd.n102 vdd.n101 9.3005
R4844 vdd.n104 vdd.n103 9.3005
R4845 vdd.n87 vdd.n86 9.3005
R4846 vdd.n110 vdd.n109 9.3005
R4847 vdd.n112 vdd.n111 9.3005
R4848 vdd.n84 vdd.n81 9.3005
R4849 vdd.n119 vdd.n118 9.3005
R4850 vdd.n45 vdd.n44 9.3005
R4851 vdd.n40 vdd.n39 9.3005
R4852 vdd.n51 vdd.n50 9.3005
R4853 vdd.n53 vdd.n52 9.3005
R4854 vdd.n36 vdd.n35 9.3005
R4855 vdd.n59 vdd.n58 9.3005
R4856 vdd.n61 vdd.n60 9.3005
R4857 vdd.n33 vdd.n30 9.3005
R4858 vdd.n68 vdd.n67 9.3005
R4859 vdd.n3036 vdd.n3035 9.3005
R4860 vdd.n3037 vdd.n578 9.3005
R4861 vdd.n577 vdd.n575 9.3005
R4862 vdd.n3043 vdd.n574 9.3005
R4863 vdd.n3044 vdd.n573 9.3005
R4864 vdd.n3045 vdd.n572 9.3005
R4865 vdd.n571 vdd.n569 9.3005
R4866 vdd.n3051 vdd.n568 9.3005
R4867 vdd.n3052 vdd.n567 9.3005
R4868 vdd.n3053 vdd.n566 9.3005
R4869 vdd.n565 vdd.n563 9.3005
R4870 vdd.n3059 vdd.n562 9.3005
R4871 vdd.n3060 vdd.n561 9.3005
R4872 vdd.n3061 vdd.n560 9.3005
R4873 vdd.n559 vdd.n557 9.3005
R4874 vdd.n3067 vdd.n556 9.3005
R4875 vdd.n3068 vdd.n555 9.3005
R4876 vdd.n3069 vdd.n554 9.3005
R4877 vdd.n553 vdd.n551 9.3005
R4878 vdd.n3075 vdd.n550 9.3005
R4879 vdd.n3076 vdd.n549 9.3005
R4880 vdd.n3077 vdd.n548 9.3005
R4881 vdd.n547 vdd.n545 9.3005
R4882 vdd.n3083 vdd.n542 9.3005
R4883 vdd.n3084 vdd.n541 9.3005
R4884 vdd.n3085 vdd.n540 9.3005
R4885 vdd.n539 vdd.n537 9.3005
R4886 vdd.n3091 vdd.n536 9.3005
R4887 vdd.n3092 vdd.n535 9.3005
R4888 vdd.n3093 vdd.n534 9.3005
R4889 vdd.n533 vdd.n531 9.3005
R4890 vdd.n3099 vdd.n530 9.3005
R4891 vdd.n3100 vdd.n529 9.3005
R4892 vdd.n3101 vdd.n528 9.3005
R4893 vdd.n527 vdd.n525 9.3005
R4894 vdd.n3106 vdd.n524 9.3005
R4895 vdd.n3116 vdd.n518 9.3005
R4896 vdd.n3118 vdd.n3117 9.3005
R4897 vdd.n509 vdd.n508 9.3005
R4898 vdd.n3133 vdd.n3132 9.3005
R4899 vdd.n3134 vdd.n507 9.3005
R4900 vdd.n3136 vdd.n3135 9.3005
R4901 vdd.n497 vdd.n496 9.3005
R4902 vdd.n3149 vdd.n3148 9.3005
R4903 vdd.n3150 vdd.n495 9.3005
R4904 vdd.n3152 vdd.n3151 9.3005
R4905 vdd.n485 vdd.n484 9.3005
R4906 vdd.n3166 vdd.n3165 9.3005
R4907 vdd.n3167 vdd.n483 9.3005
R4908 vdd.n3169 vdd.n3168 9.3005
R4909 vdd.n312 vdd.n310 9.3005
R4910 vdd.n3120 vdd.n3119 9.3005
R4911 vdd.n3349 vdd.n3348 9.3005
R4912 vdd.n313 vdd.n311 9.3005
R4913 vdd.n3342 vdd.n320 9.3005
R4914 vdd.n3341 vdd.n321 9.3005
R4915 vdd.n3340 vdd.n322 9.3005
R4916 vdd.n331 vdd.n323 9.3005
R4917 vdd.n3334 vdd.n332 9.3005
R4918 vdd.n3333 vdd.n333 9.3005
R4919 vdd.n3332 vdd.n334 9.3005
R4920 vdd.n342 vdd.n335 9.3005
R4921 vdd.n3326 vdd.n343 9.3005
R4922 vdd.n3325 vdd.n344 9.3005
R4923 vdd.n3324 vdd.n345 9.3005
R4924 vdd.n353 vdd.n346 9.3005
R4925 vdd.n3318 vdd.n3317 9.3005
R4926 vdd.n3314 vdd.n354 9.3005
R4927 vdd.n3313 vdd.n357 9.3005
R4928 vdd.n361 vdd.n358 9.3005
R4929 vdd.n362 vdd.n359 9.3005
R4930 vdd.n3306 vdd.n363 9.3005
R4931 vdd.n3305 vdd.n364 9.3005
R4932 vdd.n3304 vdd.n365 9.3005
R4933 vdd.n369 vdd.n366 9.3005
R4934 vdd.n3299 vdd.n370 9.3005
R4935 vdd.n3298 vdd.n371 9.3005
R4936 vdd.n3297 vdd.n372 9.3005
R4937 vdd.n376 vdd.n373 9.3005
R4938 vdd.n3292 vdd.n377 9.3005
R4939 vdd.n3291 vdd.n378 9.3005
R4940 vdd.n3290 vdd.n379 9.3005
R4941 vdd.n383 vdd.n380 9.3005
R4942 vdd.n3285 vdd.n384 9.3005
R4943 vdd.n3284 vdd.n385 9.3005
R4944 vdd.n3283 vdd.n3282 9.3005
R4945 vdd.n3281 vdd.n386 9.3005
R4946 vdd.n3280 vdd.n3279 9.3005
R4947 vdd.n392 vdd.n391 9.3005
R4948 vdd.n3274 vdd.n396 9.3005
R4949 vdd.n3273 vdd.n397 9.3005
R4950 vdd.n3272 vdd.n398 9.3005
R4951 vdd.n402 vdd.n399 9.3005
R4952 vdd.n3267 vdd.n403 9.3005
R4953 vdd.n3266 vdd.n404 9.3005
R4954 vdd.n3265 vdd.n405 9.3005
R4955 vdd.n409 vdd.n406 9.3005
R4956 vdd.n3260 vdd.n410 9.3005
R4957 vdd.n3259 vdd.n411 9.3005
R4958 vdd.n3258 vdd.n412 9.3005
R4959 vdd.n416 vdd.n413 9.3005
R4960 vdd.n3253 vdd.n417 9.3005
R4961 vdd.n3252 vdd.n418 9.3005
R4962 vdd.n3251 vdd.n419 9.3005
R4963 vdd.n423 vdd.n420 9.3005
R4964 vdd.n3246 vdd.n424 9.3005
R4965 vdd.n3245 vdd.n425 9.3005
R4966 vdd.n3244 vdd.n3243 9.3005
R4967 vdd.n3242 vdd.n426 9.3005
R4968 vdd.n3241 vdd.n3240 9.3005
R4969 vdd.n432 vdd.n431 9.3005
R4970 vdd.n3235 vdd.n436 9.3005
R4971 vdd.n3234 vdd.n437 9.3005
R4972 vdd.n3233 vdd.n438 9.3005
R4973 vdd.n442 vdd.n439 9.3005
R4974 vdd.n3228 vdd.n443 9.3005
R4975 vdd.n3227 vdd.n444 9.3005
R4976 vdd.n3226 vdd.n445 9.3005
R4977 vdd.n449 vdd.n446 9.3005
R4978 vdd.n3221 vdd.n450 9.3005
R4979 vdd.n3220 vdd.n451 9.3005
R4980 vdd.n3219 vdd.n452 9.3005
R4981 vdd.n456 vdd.n453 9.3005
R4982 vdd.n3214 vdd.n457 9.3005
R4983 vdd.n3213 vdd.n458 9.3005
R4984 vdd.n3212 vdd.n459 9.3005
R4985 vdd.n463 vdd.n460 9.3005
R4986 vdd.n3207 vdd.n464 9.3005
R4987 vdd.n3206 vdd.n465 9.3005
R4988 vdd.n3202 vdd.n3199 9.3005
R4989 vdd.n3316 vdd.n3315 9.3005
R4990 vdd.n3126 vdd.n513 9.3005
R4991 vdd.n3128 vdd.n3127 9.3005
R4992 vdd.n503 vdd.n502 9.3005
R4993 vdd.n3141 vdd.n3140 9.3005
R4994 vdd.n3142 vdd.n501 9.3005
R4995 vdd.n3144 vdd.n3143 9.3005
R4996 vdd.n490 vdd.n489 9.3005
R4997 vdd.n3157 vdd.n3156 9.3005
R4998 vdd.n3158 vdd.n488 9.3005
R4999 vdd.n3160 vdd.n3159 9.3005
R5000 vdd.n478 vdd.n477 9.3005
R5001 vdd.n3174 vdd.n3173 9.3005
R5002 vdd.n3175 vdd.n476 9.3005
R5003 vdd.n3177 vdd.n3176 9.3005
R5004 vdd.n3178 vdd.n475 9.3005
R5005 vdd.n3180 vdd.n3179 9.3005
R5006 vdd.n3181 vdd.n474 9.3005
R5007 vdd.n3183 vdd.n3182 9.3005
R5008 vdd.n3184 vdd.n472 9.3005
R5009 vdd.n3186 vdd.n3185 9.3005
R5010 vdd.n3187 vdd.n471 9.3005
R5011 vdd.n3189 vdd.n3188 9.3005
R5012 vdd.n3190 vdd.n469 9.3005
R5013 vdd.n3192 vdd.n3191 9.3005
R5014 vdd.n3193 vdd.n468 9.3005
R5015 vdd.n3195 vdd.n3194 9.3005
R5016 vdd.n3196 vdd.n466 9.3005
R5017 vdd.n3198 vdd.n3197 9.3005
R5018 vdd.n3125 vdd.n3124 9.3005
R5019 vdd.n2989 vdd.n514 9.3005
R5020 vdd.n2994 vdd.n2988 9.3005
R5021 vdd.n3004 vdd.n605 9.3005
R5022 vdd.n3005 vdd.n604 9.3005
R5023 vdd.n603 vdd.n601 9.3005
R5024 vdd.n3011 vdd.n600 9.3005
R5025 vdd.n3012 vdd.n599 9.3005
R5026 vdd.n3013 vdd.n598 9.3005
R5027 vdd.n597 vdd.n595 9.3005
R5028 vdd.n3019 vdd.n594 9.3005
R5029 vdd.n3020 vdd.n593 9.3005
R5030 vdd.n3021 vdd.n592 9.3005
R5031 vdd.n591 vdd.n589 9.3005
R5032 vdd.n3026 vdd.n588 9.3005
R5033 vdd.n3027 vdd.n587 9.3005
R5034 vdd.n583 vdd.n582 9.3005
R5035 vdd.n3033 vdd.n3032 9.3005
R5036 vdd.n3034 vdd.n579 9.3005
R5037 vdd.n1916 vdd.n1915 9.3005
R5038 vdd.n1911 vdd.n975 9.3005
R5039 vdd.n1299 vdd.n1059 9.3005
R5040 vdd.n1301 vdd.n1300 9.3005
R5041 vdd.n1050 vdd.n1049 9.3005
R5042 vdd.n1314 vdd.n1313 9.3005
R5043 vdd.n1315 vdd.n1048 9.3005
R5044 vdd.n1317 vdd.n1316 9.3005
R5045 vdd.n1037 vdd.n1036 9.3005
R5046 vdd.n1330 vdd.n1329 9.3005
R5047 vdd.n1331 vdd.n1035 9.3005
R5048 vdd.n1333 vdd.n1332 9.3005
R5049 vdd.n1026 vdd.n1025 9.3005
R5050 vdd.n1347 vdd.n1346 9.3005
R5051 vdd.n1348 vdd.n1024 9.3005
R5052 vdd.n1350 vdd.n1349 9.3005
R5053 vdd.n1015 vdd.n1014 9.3005
R5054 vdd.n1645 vdd.n1644 9.3005
R5055 vdd.n1646 vdd.n1013 9.3005
R5056 vdd.n1648 vdd.n1647 9.3005
R5057 vdd.n1003 vdd.n1002 9.3005
R5058 vdd.n1662 vdd.n1661 9.3005
R5059 vdd.n1663 vdd.n1001 9.3005
R5060 vdd.n1665 vdd.n1664 9.3005
R5061 vdd.n993 vdd.n992 9.3005
R5062 vdd.n1679 vdd.n1678 9.3005
R5063 vdd.n1680 vdd.n990 9.3005
R5064 vdd.n1684 vdd.n1683 9.3005
R5065 vdd.n1682 vdd.n991 9.3005
R5066 vdd.n1681 vdd.n980 9.3005
R5067 vdd.n1298 vdd.n1297 9.3005
R5068 vdd.n1193 vdd.n1183 9.3005
R5069 vdd.n1195 vdd.n1194 9.3005
R5070 vdd.n1196 vdd.n1182 9.3005
R5071 vdd.n1198 vdd.n1197 9.3005
R5072 vdd.n1199 vdd.n1175 9.3005
R5073 vdd.n1201 vdd.n1200 9.3005
R5074 vdd.n1202 vdd.n1174 9.3005
R5075 vdd.n1204 vdd.n1203 9.3005
R5076 vdd.n1205 vdd.n1167 9.3005
R5077 vdd.n1207 vdd.n1206 9.3005
R5078 vdd.n1208 vdd.n1166 9.3005
R5079 vdd.n1210 vdd.n1209 9.3005
R5080 vdd.n1211 vdd.n1159 9.3005
R5081 vdd.n1213 vdd.n1212 9.3005
R5082 vdd.n1214 vdd.n1158 9.3005
R5083 vdd.n1216 vdd.n1215 9.3005
R5084 vdd.n1217 vdd.n1152 9.3005
R5085 vdd.n1219 vdd.n1218 9.3005
R5086 vdd.n1220 vdd.n1150 9.3005
R5087 vdd.n1222 vdd.n1221 9.3005
R5088 vdd.n1151 vdd.n1148 9.3005
R5089 vdd.n1229 vdd.n1144 9.3005
R5090 vdd.n1231 vdd.n1230 9.3005
R5091 vdd.n1232 vdd.n1143 9.3005
R5092 vdd.n1234 vdd.n1233 9.3005
R5093 vdd.n1235 vdd.n1136 9.3005
R5094 vdd.n1237 vdd.n1236 9.3005
R5095 vdd.n1238 vdd.n1135 9.3005
R5096 vdd.n1240 vdd.n1239 9.3005
R5097 vdd.n1241 vdd.n1128 9.3005
R5098 vdd.n1243 vdd.n1242 9.3005
R5099 vdd.n1244 vdd.n1127 9.3005
R5100 vdd.n1246 vdd.n1245 9.3005
R5101 vdd.n1247 vdd.n1120 9.3005
R5102 vdd.n1249 vdd.n1248 9.3005
R5103 vdd.n1250 vdd.n1119 9.3005
R5104 vdd.n1252 vdd.n1251 9.3005
R5105 vdd.n1253 vdd.n1112 9.3005
R5106 vdd.n1255 vdd.n1254 9.3005
R5107 vdd.n1256 vdd.n1111 9.3005
R5108 vdd.n1258 vdd.n1257 9.3005
R5109 vdd.n1259 vdd.n1104 9.3005
R5110 vdd.n1261 vdd.n1260 9.3005
R5111 vdd.n1262 vdd.n1103 9.3005
R5112 vdd.n1264 vdd.n1263 9.3005
R5113 vdd.n1265 vdd.n1094 9.3005
R5114 vdd.n1267 vdd.n1266 9.3005
R5115 vdd.n1268 vdd.n1093 9.3005
R5116 vdd.n1270 vdd.n1269 9.3005
R5117 vdd.n1271 vdd.n1086 9.3005
R5118 vdd.n1273 vdd.n1272 9.3005
R5119 vdd.n1274 vdd.n1085 9.3005
R5120 vdd.n1276 vdd.n1275 9.3005
R5121 vdd.n1277 vdd.n1078 9.3005
R5122 vdd.n1279 vdd.n1278 9.3005
R5123 vdd.n1280 vdd.n1077 9.3005
R5124 vdd.n1282 vdd.n1281 9.3005
R5125 vdd.n1283 vdd.n1070 9.3005
R5126 vdd.n1285 vdd.n1284 9.3005
R5127 vdd.n1286 vdd.n1069 9.3005
R5128 vdd.n1288 vdd.n1287 9.3005
R5129 vdd.n1289 vdd.n1065 9.3005
R5130 vdd.n1291 vdd.n1290 9.3005
R5131 vdd.n1189 vdd.n1060 9.3005
R5132 vdd.n1056 vdd.n1055 9.3005
R5133 vdd.n1306 vdd.n1305 9.3005
R5134 vdd.n1307 vdd.n1054 9.3005
R5135 vdd.n1309 vdd.n1308 9.3005
R5136 vdd.n1044 vdd.n1043 9.3005
R5137 vdd.n1322 vdd.n1321 9.3005
R5138 vdd.n1323 vdd.n1042 9.3005
R5139 vdd.n1325 vdd.n1324 9.3005
R5140 vdd.n1032 vdd.n1031 9.3005
R5141 vdd.n1339 vdd.n1338 9.3005
R5142 vdd.n1340 vdd.n1030 9.3005
R5143 vdd.n1342 vdd.n1341 9.3005
R5144 vdd.n1021 vdd.n1020 9.3005
R5145 vdd.n1293 vdd.n1292 9.3005
R5146 vdd.n1637 vdd.n1354 9.3005
R5147 vdd.n1558 vdd.n1557 9.3005
R5148 vdd.n1553 vdd.n1552 9.3005
R5149 vdd.n1564 vdd.n1563 9.3005
R5150 vdd.n1566 vdd.n1565 9.3005
R5151 vdd.n1549 vdd.n1548 9.3005
R5152 vdd.n1572 vdd.n1571 9.3005
R5153 vdd.n1574 vdd.n1573 9.3005
R5154 vdd.n1546 vdd.n1543 9.3005
R5155 vdd.n1581 vdd.n1580 9.3005
R5156 vdd.n1609 vdd.n1608 9.3005
R5157 vdd.n1604 vdd.n1603 9.3005
R5158 vdd.n1615 vdd.n1614 9.3005
R5159 vdd.n1617 vdd.n1616 9.3005
R5160 vdd.n1600 vdd.n1599 9.3005
R5161 vdd.n1623 vdd.n1622 9.3005
R5162 vdd.n1625 vdd.n1624 9.3005
R5163 vdd.n1597 vdd.n1594 9.3005
R5164 vdd.n1632 vdd.n1631 9.3005
R5165 vdd.n1464 vdd.n1463 9.3005
R5166 vdd.n1459 vdd.n1458 9.3005
R5167 vdd.n1470 vdd.n1469 9.3005
R5168 vdd.n1472 vdd.n1471 9.3005
R5169 vdd.n1455 vdd.n1454 9.3005
R5170 vdd.n1478 vdd.n1477 9.3005
R5171 vdd.n1480 vdd.n1479 9.3005
R5172 vdd.n1452 vdd.n1449 9.3005
R5173 vdd.n1487 vdd.n1486 9.3005
R5174 vdd.n1515 vdd.n1514 9.3005
R5175 vdd.n1510 vdd.n1509 9.3005
R5176 vdd.n1521 vdd.n1520 9.3005
R5177 vdd.n1523 vdd.n1522 9.3005
R5178 vdd.n1506 vdd.n1505 9.3005
R5179 vdd.n1529 vdd.n1528 9.3005
R5180 vdd.n1531 vdd.n1530 9.3005
R5181 vdd.n1503 vdd.n1500 9.3005
R5182 vdd.n1538 vdd.n1537 9.3005
R5183 vdd.n1371 vdd.n1370 9.3005
R5184 vdd.n1366 vdd.n1365 9.3005
R5185 vdd.n1377 vdd.n1376 9.3005
R5186 vdd.n1379 vdd.n1378 9.3005
R5187 vdd.n1362 vdd.n1361 9.3005
R5188 vdd.n1385 vdd.n1384 9.3005
R5189 vdd.n1387 vdd.n1386 9.3005
R5190 vdd.n1359 vdd.n1356 9.3005
R5191 vdd.n1394 vdd.n1393 9.3005
R5192 vdd.n1422 vdd.n1421 9.3005
R5193 vdd.n1417 vdd.n1416 9.3005
R5194 vdd.n1428 vdd.n1427 9.3005
R5195 vdd.n1430 vdd.n1429 9.3005
R5196 vdd.n1413 vdd.n1412 9.3005
R5197 vdd.n1436 vdd.n1435 9.3005
R5198 vdd.n1438 vdd.n1437 9.3005
R5199 vdd.n1410 vdd.n1407 9.3005
R5200 vdd.n1445 vdd.n1444 9.3005
R5201 vdd.n288 vdd.n287 8.92171
R5202 vdd.n237 vdd.n236 8.92171
R5203 vdd.n194 vdd.n193 8.92171
R5204 vdd.n143 vdd.n142 8.92171
R5205 vdd.n101 vdd.n100 8.92171
R5206 vdd.n50 vdd.n49 8.92171
R5207 vdd.n1563 vdd.n1562 8.92171
R5208 vdd.n1614 vdd.n1613 8.92171
R5209 vdd.n1469 vdd.n1468 8.92171
R5210 vdd.n1520 vdd.n1519 8.92171
R5211 vdd.n1376 vdd.n1375 8.92171
R5212 vdd.n1427 vdd.n1426 8.92171
R5213 vdd.n215 vdd.n121 8.81535
R5214 vdd.n1541 vdd.n1447 8.81535
R5215 vdd.n1676 vdd.t4 8.72962
R5216 vdd.n3138 vdd.t14 8.72962
R5217 vdd.t47 vdd.n1650 8.50289
R5218 vdd.n493 vdd.t64 8.50289
R5219 vdd.n28 vdd.n14 8.42249
R5220 vdd.n1352 vdd.t49 8.27616
R5221 vdd.n3346 vdd.t10 8.27616
R5222 vdd.n3350 vdd.n3349 8.16225
R5223 vdd.n1637 vdd.n1636 8.16225
R5224 vdd.n284 vdd.n278 8.14595
R5225 vdd.n233 vdd.n227 8.14595
R5226 vdd.n190 vdd.n184 8.14595
R5227 vdd.n139 vdd.n133 8.14595
R5228 vdd.n97 vdd.n91 8.14595
R5229 vdd.n46 vdd.n40 8.14595
R5230 vdd.n1559 vdd.n1553 8.14595
R5231 vdd.n1610 vdd.n1604 8.14595
R5232 vdd.n1465 vdd.n1459 8.14595
R5233 vdd.n1516 vdd.n1510 8.14595
R5234 vdd.n1372 vdd.n1366 8.14595
R5235 vdd.n1423 vdd.n1417 8.14595
R5236 vdd.t51 vdd.n1040 8.04943
R5237 vdd.n3337 vdd.t57 8.04943
R5238 vdd.n2179 vdd.n932 7.70933
R5239 vdd.n2185 vdd.n932 7.70933
R5240 vdd.n2191 vdd.n926 7.70933
R5241 vdd.n2191 vdd.n920 7.70933
R5242 vdd.n2197 vdd.n920 7.70933
R5243 vdd.n2197 vdd.n914 7.70933
R5244 vdd.n2203 vdd.n914 7.70933
R5245 vdd.n2209 vdd.n908 7.70933
R5246 vdd.n2215 vdd.n902 7.70933
R5247 vdd.n2221 vdd.n895 7.70933
R5248 vdd.n2221 vdd.n898 7.70933
R5249 vdd.n2227 vdd.n891 7.70933
R5250 vdd.n2234 vdd.n877 7.70933
R5251 vdd.n2240 vdd.n877 7.70933
R5252 vdd.n2246 vdd.n871 7.70933
R5253 vdd.n2252 vdd.n867 7.70933
R5254 vdd.n2258 vdd.n861 7.70933
R5255 vdd.n2276 vdd.n843 7.70933
R5256 vdd.n2276 vdd.n836 7.70933
R5257 vdd.n2284 vdd.n836 7.70933
R5258 vdd.n2366 vdd.n820 7.70933
R5259 vdd.n2729 vdd.n774 7.70933
R5260 vdd.n2741 vdd.n755 7.70933
R5261 vdd.n2747 vdd.n755 7.70933
R5262 vdd.n2747 vdd.n758 7.70933
R5263 vdd.n2765 vdd.n739 7.70933
R5264 vdd.n2771 vdd.n733 7.70933
R5265 vdd.n2777 vdd.n729 7.70933
R5266 vdd.n2783 vdd.n716 7.70933
R5267 vdd.n2789 vdd.n716 7.70933
R5268 vdd.n2796 vdd.n709 7.70933
R5269 vdd.n2802 vdd.n702 7.70933
R5270 vdd.n2802 vdd.n705 7.70933
R5271 vdd.n2808 vdd.n698 7.70933
R5272 vdd.n2814 vdd.n692 7.70933
R5273 vdd.n2820 vdd.n679 7.70933
R5274 vdd.n2826 vdd.n679 7.70933
R5275 vdd.n2826 vdd.n671 7.70933
R5276 vdd.n2877 vdd.n671 7.70933
R5277 vdd.n2877 vdd.n674 7.70933
R5278 vdd.n2883 vdd.n631 7.70933
R5279 vdd.n2953 vdd.n631 7.70933
R5280 vdd.t223 vdd.n908 7.59597
R5281 vdd.n2058 vdd.t175 7.59597
R5282 vdd.n2701 vdd.t178 7.59597
R5283 vdd.n692 vdd.t202 7.59597
R5284 vdd.n283 vdd.n280 7.3702
R5285 vdd.n232 vdd.n229 7.3702
R5286 vdd.n189 vdd.n186 7.3702
R5287 vdd.n138 vdd.n135 7.3702
R5288 vdd.n96 vdd.n93 7.3702
R5289 vdd.n45 vdd.n42 7.3702
R5290 vdd.n1558 vdd.n1555 7.3702
R5291 vdd.n1609 vdd.n1606 7.3702
R5292 vdd.n1464 vdd.n1461 7.3702
R5293 vdd.n1515 vdd.n1512 7.3702
R5294 vdd.n1371 vdd.n1368 7.3702
R5295 vdd.n1422 vdd.n1419 7.3702
R5296 vdd.n1319 vdd.t25 7.1425
R5297 vdd.n3330 vdd.t2 7.1425
R5298 vdd.n1230 vdd.n1229 6.98232
R5299 vdd.n1831 vdd.n1830 6.98232
R5300 vdd.n3245 vdd.n3244 6.98232
R5301 vdd.n3037 vdd.n3036 6.98232
R5302 vdd.n1335 vdd.t62 6.91577
R5303 vdd.n2215 vdd.t186 6.91577
R5304 vdd.n2808 vdd.t211 6.91577
R5305 vdd.n325 vdd.t27 6.91577
R5306 vdd.n2793 vdd.n2792 6.86879
R5307 vdd.n2231 vdd.n2230 6.86879
R5308 vdd.n2291 vdd.t218 6.80241
R5309 vdd.n2735 vdd.t206 6.80241
R5310 vdd.n1642 vdd.t12 6.68904
R5311 vdd.n3171 vdd.t18 6.68904
R5312 vdd.n1005 vdd.t29 6.46231
R5313 vdd.t33 vdd.n492 6.46231
R5314 vdd.n2058 vdd.t176 6.34895
R5315 vdd.n2701 vdd.t216 6.34895
R5316 vdd.n3350 vdd.n309 6.27748
R5317 vdd.n1636 vdd.n1635 6.27748
R5318 vdd.t189 vdd.n871 6.00885
R5319 vdd.n729 vdd.t194 6.00885
R5320 vdd.n284 vdd.n283 5.81868
R5321 vdd.n233 vdd.n232 5.81868
R5322 vdd.n190 vdd.n189 5.81868
R5323 vdd.n139 vdd.n138 5.81868
R5324 vdd.n97 vdd.n96 5.81868
R5325 vdd.n46 vdd.n45 5.81868
R5326 vdd.n1559 vdd.n1558 5.81868
R5327 vdd.n1610 vdd.n1609 5.81868
R5328 vdd.n1465 vdd.n1464 5.81868
R5329 vdd.n1516 vdd.n1515 5.81868
R5330 vdd.n1372 vdd.n1371 5.81868
R5331 vdd.n1423 vdd.n1422 5.81868
R5332 vdd.n2374 vdd.n2373 5.77611
R5333 vdd.n2114 vdd.n2113 5.77611
R5334 vdd.n2603 vdd.n2602 5.77611
R5335 vdd.n2892 vdd.n663 5.77611
R5336 vdd.n2958 vdd.n627 5.77611
R5337 vdd.n2539 vdd.n2475 5.77611
R5338 vdd.n2299 vdd.n827 5.77611
R5339 vdd.n1990 vdd.n1989 5.77611
R5340 vdd.n1192 vdd.n1189 5.62474
R5341 vdd.n1914 vdd.n1911 5.62474
R5342 vdd.n3205 vdd.n3202 5.62474
R5343 vdd.n2992 vdd.n2989 5.62474
R5344 vdd.n2252 vdd.t214 5.44203
R5345 vdd.n2771 vdd.t190 5.44203
R5346 vdd.n2227 vdd.t203 5.10193
R5347 vdd.n2246 vdd.t222 5.10193
R5348 vdd.n2777 vdd.t212 5.10193
R5349 vdd.n2796 vdd.t181 5.10193
R5350 vdd.n287 vdd.n278 5.04292
R5351 vdd.n236 vdd.n227 5.04292
R5352 vdd.n193 vdd.n184 5.04292
R5353 vdd.n142 vdd.n133 5.04292
R5354 vdd.n100 vdd.n91 5.04292
R5355 vdd.n49 vdd.n40 5.04292
R5356 vdd.n1562 vdd.n1553 5.04292
R5357 vdd.n1613 vdd.n1604 5.04292
R5358 vdd.n1468 vdd.n1459 5.04292
R5359 vdd.n1519 vdd.n1510 5.04292
R5360 vdd.n1375 vdd.n1366 5.04292
R5361 vdd.n1426 vdd.n1417 5.04292
R5362 vdd.n891 vdd.t152 4.98857
R5363 vdd.t110 vdd.n709 4.98857
R5364 vdd.n1668 vdd.t29 4.8752
R5365 vdd.t103 vdd.n926 4.8752
R5366 vdd.t184 vdd.t195 4.8752
R5367 vdd.n2046 vdd.t141 4.8752
R5368 vdd.n2713 vdd.t145 4.8752
R5369 vdd.t224 vdd.t174 4.8752
R5370 vdd.n674 vdd.t99 4.8752
R5371 vdd.n3146 vdd.t33 4.8752
R5372 vdd.n2375 vdd.n2374 4.83952
R5373 vdd.n2115 vdd.n2114 4.83952
R5374 vdd.n2602 vdd.n2601 4.83952
R5375 vdd.n663 vdd.n658 4.83952
R5376 vdd.n627 vdd.n622 4.83952
R5377 vdd.n2536 vdd.n2475 4.83952
R5378 vdd.n2302 vdd.n827 4.83952
R5379 vdd.n1989 vdd.n1988 4.83952
R5380 vdd.n2270 vdd.t209 4.76184
R5381 vdd.n2753 vdd.t198 4.76184
R5382 vdd.n1799 vdd.n973 4.74817
R5383 vdd.n1794 vdd.n974 4.74817
R5384 vdd.n1696 vdd.n1693 4.74817
R5385 vdd.n1895 vdd.n1697 4.74817
R5386 vdd.n1897 vdd.n1696 4.74817
R5387 vdd.n1896 vdd.n1895 4.74817
R5388 vdd.n521 vdd.n519 4.74817
R5389 vdd.n3107 vdd.n522 4.74817
R5390 vdd.n3110 vdd.n522 4.74817
R5391 vdd.n3111 vdd.n521 4.74817
R5392 vdd.n2999 vdd.n606 4.74817
R5393 vdd.n2995 vdd.n608 4.74817
R5394 vdd.n2998 vdd.n608 4.74817
R5395 vdd.n3003 vdd.n606 4.74817
R5396 vdd.n1795 vdd.n973 4.74817
R5397 vdd.n976 vdd.n974 4.74817
R5398 vdd.n309 vdd.n308 4.7074
R5399 vdd.n215 vdd.n214 4.7074
R5400 vdd.n1635 vdd.n1634 4.7074
R5401 vdd.n1541 vdd.n1540 4.7074
R5402 vdd.t12 vdd.n1011 4.64847
R5403 vdd.n3162 vdd.t18 4.64847
R5404 vdd.n1344 vdd.t62 4.42174
R5405 vdd.n3344 vdd.t27 4.42174
R5406 vdd.n2046 vdd.t192 4.30838
R5407 vdd.n2713 vdd.t179 4.30838
R5408 vdd.n288 vdd.n276 4.26717
R5409 vdd.n237 vdd.n225 4.26717
R5410 vdd.n194 vdd.n182 4.26717
R5411 vdd.n143 vdd.n131 4.26717
R5412 vdd.n101 vdd.n89 4.26717
R5413 vdd.n50 vdd.n38 4.26717
R5414 vdd.n1563 vdd.n1551 4.26717
R5415 vdd.n1614 vdd.n1602 4.26717
R5416 vdd.n1469 vdd.n1457 4.26717
R5417 vdd.n1520 vdd.n1508 4.26717
R5418 vdd.n1376 vdd.n1364 4.26717
R5419 vdd.n1427 vdd.n1415 4.26717
R5420 vdd.t25 vdd.n1039 4.19501
R5421 vdd.t185 vdd.n902 4.19501
R5422 vdd.n861 vdd.t197 4.19501
R5423 vdd.t213 vdd.n739 4.19501
R5424 vdd.n698 vdd.t208 4.19501
R5425 vdd.t2 vdd.n329 4.19501
R5426 vdd.n309 vdd.n215 4.10845
R5427 vdd.n1635 vdd.n1541 4.10845
R5428 vdd.n265 vdd.t88 4.06363
R5429 vdd.n265 vdd.t232 4.06363
R5430 vdd.n263 vdd.t85 4.06363
R5431 vdd.n263 vdd.t72 4.06363
R5432 vdd.n261 vdd.t36 4.06363
R5433 vdd.n261 vdd.t11 4.06363
R5434 vdd.n259 vdd.t81 4.06363
R5435 vdd.n259 vdd.t71 4.06363
R5436 vdd.n257 vdd.t34 4.06363
R5437 vdd.n257 vdd.t83 4.06363
R5438 vdd.n171 vdd.t58 4.06363
R5439 vdd.n171 vdd.t77 4.06363
R5440 vdd.n169 vdd.t74 4.06363
R5441 vdd.n169 vdd.t60 4.06363
R5442 vdd.n167 vdd.t234 4.06363
R5443 vdd.n167 vdd.t171 4.06363
R5444 vdd.n165 vdd.t66 4.06363
R5445 vdd.n165 vdd.t235 4.06363
R5446 vdd.n163 vdd.t76 4.06363
R5447 vdd.n163 vdd.t238 4.06363
R5448 vdd.n78 vdd.t89 4.06363
R5449 vdd.n78 vdd.t3 4.06363
R5450 vdd.n76 vdd.t28 4.06363
R5451 vdd.n76 vdd.t22 4.06363
R5452 vdd.n74 vdd.t67 4.06363
R5453 vdd.n74 vdd.t61 4.06363
R5454 vdd.n72 vdd.t65 4.06363
R5455 vdd.n72 vdd.t19 4.06363
R5456 vdd.n70 vdd.t227 4.06363
R5457 vdd.n70 vdd.t228 4.06363
R5458 vdd.n1583 vdd.t17 4.06363
R5459 vdd.n1583 vdd.t30 4.06363
R5460 vdd.n1585 vdd.t172 4.06363
R5461 vdd.n1585 vdd.t73 4.06363
R5462 vdd.n1587 vdd.t54 4.06363
R5463 vdd.n1587 vdd.t55 4.06363
R5464 vdd.n1589 vdd.t231 4.06363
R5465 vdd.n1589 vdd.t86 4.06363
R5466 vdd.n1591 vdd.t26 4.06363
R5467 vdd.n1591 vdd.t56 4.06363
R5468 vdd.n1489 vdd.t53 4.06363
R5469 vdd.n1489 vdd.t239 4.06363
R5470 vdd.n1491 vdd.t13 4.06363
R5471 vdd.n1491 vdd.t48 4.06363
R5472 vdd.n1493 vdd.t50 4.06363
R5473 vdd.n1493 vdd.t237 4.06363
R5474 vdd.n1495 vdd.t79 4.06363
R5475 vdd.n1495 vdd.t226 4.06363
R5476 vdd.n1497 vdd.t90 4.06363
R5477 vdd.n1497 vdd.t52 4.06363
R5478 vdd.n1396 vdd.t230 4.06363
R5479 vdd.n1396 vdd.t59 4.06363
R5480 vdd.n1398 vdd.t20 4.06363
R5481 vdd.n1398 vdd.t170 4.06363
R5482 vdd.n1400 vdd.t84 4.06363
R5483 vdd.n1400 vdd.t7 4.06363
R5484 vdd.n1402 vdd.t24 4.06363
R5485 vdd.n1402 vdd.t63 4.06363
R5486 vdd.n1404 vdd.t233 4.06363
R5487 vdd.n1404 vdd.t80 4.06363
R5488 vdd.n26 vdd.t43 3.9605
R5489 vdd.n26 vdd.t40 3.9605
R5490 vdd.n23 vdd.t42 3.9605
R5491 vdd.n23 vdd.t70 3.9605
R5492 vdd.n21 vdd.t41 3.9605
R5493 vdd.n21 vdd.t93 3.9605
R5494 vdd.n20 vdd.t69 3.9605
R5495 vdd.n20 vdd.t39 3.9605
R5496 vdd.n15 vdd.t8 3.9605
R5497 vdd.n15 vdd.t92 3.9605
R5498 vdd.n16 vdd.t45 3.9605
R5499 vdd.n16 vdd.t37 3.9605
R5500 vdd.n18 vdd.t9 3.9605
R5501 vdd.n18 vdd.t44 3.9605
R5502 vdd.n25 vdd.t38 3.9605
R5503 vdd.n25 vdd.t68 3.9605
R5504 vdd.n2792 vdd.n2791 3.74684
R5505 vdd.n2232 vdd.n2231 3.74684
R5506 vdd.n7 vdd.t225 3.61217
R5507 vdd.n7 vdd.t191 3.61217
R5508 vdd.n8 vdd.t199 3.61217
R5509 vdd.n8 vdd.t217 3.61217
R5510 vdd.n10 vdd.t207 3.61217
R5511 vdd.n10 vdd.t180 3.61217
R5512 vdd.n12 vdd.t188 3.61217
R5513 vdd.n12 vdd.t205 3.61217
R5514 vdd.n5 vdd.t221 3.61217
R5515 vdd.n5 vdd.t201 3.61217
R5516 vdd.n3 vdd.t193 3.61217
R5517 vdd.n3 vdd.t219 3.61217
R5518 vdd.n1 vdd.t177 3.61217
R5519 vdd.n1 vdd.t210 3.61217
R5520 vdd.n0 vdd.t215 3.61217
R5521 vdd.n0 vdd.t196 3.61217
R5522 vdd.n2209 vdd.t185 3.51482
R5523 vdd.n2264 vdd.t197 3.51482
R5524 vdd.n2759 vdd.t213 3.51482
R5525 vdd.n2814 vdd.t208 3.51482
R5526 vdd.n292 vdd.n291 3.49141
R5527 vdd.n241 vdd.n240 3.49141
R5528 vdd.n198 vdd.n197 3.49141
R5529 vdd.n147 vdd.n146 3.49141
R5530 vdd.n105 vdd.n104 3.49141
R5531 vdd.n54 vdd.n53 3.49141
R5532 vdd.n1567 vdd.n1566 3.49141
R5533 vdd.n1618 vdd.n1617 3.49141
R5534 vdd.n1473 vdd.n1472 3.49141
R5535 vdd.n1524 vdd.n1523 3.49141
R5536 vdd.n1380 vdd.n1379 3.49141
R5537 vdd.n1431 vdd.n1430 3.49141
R5538 vdd.n2284 vdd.t192 3.40145
R5539 vdd.n2438 vdd.t220 3.40145
R5540 vdd.n2722 vdd.t204 3.40145
R5541 vdd.n2741 vdd.t179 3.40145
R5542 vdd.n1327 vdd.t51 3.28809
R5543 vdd.t57 vdd.n3336 3.28809
R5544 vdd.n1028 vdd.t49 3.06136
R5545 vdd.t10 vdd.n3345 3.06136
R5546 vdd.t209 vdd.n843 2.94799
R5547 vdd.n758 vdd.t198 2.94799
R5548 vdd.n1651 vdd.t47 2.83463
R5549 vdd.n2185 vdd.t103 2.83463
R5550 vdd.n2291 vdd.t141 2.83463
R5551 vdd.n2735 vdd.t145 2.83463
R5552 vdd.n2883 vdd.t99 2.83463
R5553 vdd.n3163 vdd.t64 2.83463
R5554 vdd.n295 vdd.n274 2.71565
R5555 vdd.n244 vdd.n223 2.71565
R5556 vdd.n201 vdd.n180 2.71565
R5557 vdd.n150 vdd.n129 2.71565
R5558 vdd.n108 vdd.n87 2.71565
R5559 vdd.n57 vdd.n36 2.71565
R5560 vdd.n1570 vdd.n1549 2.71565
R5561 vdd.n1621 vdd.n1600 2.71565
R5562 vdd.n1476 vdd.n1455 2.71565
R5563 vdd.n1527 vdd.n1506 2.71565
R5564 vdd.n1383 vdd.n1362 2.71565
R5565 vdd.n1434 vdd.n1413 2.71565
R5566 vdd.n1667 vdd.t4 2.6079
R5567 vdd.n898 vdd.t203 2.6079
R5568 vdd.n2070 vdd.t222 2.6079
R5569 vdd.n2689 vdd.t212 2.6079
R5570 vdd.t181 vdd.n702 2.6079
R5571 vdd.t14 vdd.n499 2.6079
R5572 vdd.n282 vdd.n281 2.4129
R5573 vdd.n231 vdd.n230 2.4129
R5574 vdd.n188 vdd.n187 2.4129
R5575 vdd.n137 vdd.n136 2.4129
R5576 vdd.n95 vdd.n94 2.4129
R5577 vdd.n44 vdd.n43 2.4129
R5578 vdd.n1557 vdd.n1556 2.4129
R5579 vdd.n1608 vdd.n1607 2.4129
R5580 vdd.n1463 vdd.n1462 2.4129
R5581 vdd.n1514 vdd.n1513 2.4129
R5582 vdd.n1370 vdd.n1369 2.4129
R5583 vdd.n1421 vdd.n1420 2.4129
R5584 vdd.n1894 vdd.n1696 2.27742
R5585 vdd.n1895 vdd.n1894 2.27742
R5586 vdd.n2919 vdd.n522 2.27742
R5587 vdd.n2919 vdd.n521 2.27742
R5588 vdd.n2987 vdd.n608 2.27742
R5589 vdd.n2987 vdd.n606 2.27742
R5590 vdd.n1917 vdd.n973 2.27742
R5591 vdd.n1917 vdd.n974 2.27742
R5592 vdd.n2070 vdd.t214 2.2678
R5593 vdd.n2689 vdd.t190 2.2678
R5594 vdd.n2258 vdd.t195 2.04107
R5595 vdd.n2765 vdd.t224 2.04107
R5596 vdd.n296 vdd.n272 1.93989
R5597 vdd.n245 vdd.n221 1.93989
R5598 vdd.n202 vdd.n178 1.93989
R5599 vdd.n151 vdd.n127 1.93989
R5600 vdd.n109 vdd.n85 1.93989
R5601 vdd.n58 vdd.n34 1.93989
R5602 vdd.n1571 vdd.n1547 1.93989
R5603 vdd.n1622 vdd.n1598 1.93989
R5604 vdd.n1477 vdd.n1453 1.93989
R5605 vdd.n1528 vdd.n1504 1.93989
R5606 vdd.n1384 vdd.n1360 1.93989
R5607 vdd.n1435 vdd.n1411 1.93989
R5608 vdd.n2234 vdd.t182 1.70098
R5609 vdd.n2240 vdd.t189 1.70098
R5610 vdd.n2783 vdd.t194 1.70098
R5611 vdd.n2789 vdd.t183 1.70098
R5612 vdd.n1063 vdd.t121 1.47425
R5613 vdd.t125 vdd.n3321 1.47425
R5614 vdd.n2264 vdd.t176 1.36088
R5615 vdd.n2759 vdd.t216 1.36088
R5616 vdd.n307 vdd.n267 1.16414
R5617 vdd.n300 vdd.n299 1.16414
R5618 vdd.n256 vdd.n216 1.16414
R5619 vdd.n249 vdd.n248 1.16414
R5620 vdd.n213 vdd.n173 1.16414
R5621 vdd.n206 vdd.n205 1.16414
R5622 vdd.n162 vdd.n122 1.16414
R5623 vdd.n155 vdd.n154 1.16414
R5624 vdd.n120 vdd.n80 1.16414
R5625 vdd.n113 vdd.n112 1.16414
R5626 vdd.n69 vdd.n29 1.16414
R5627 vdd.n62 vdd.n61 1.16414
R5628 vdd.n1582 vdd.n1542 1.16414
R5629 vdd.n1575 vdd.n1574 1.16414
R5630 vdd.n1633 vdd.n1593 1.16414
R5631 vdd.n1626 vdd.n1625 1.16414
R5632 vdd.n1488 vdd.n1448 1.16414
R5633 vdd.n1481 vdd.n1480 1.16414
R5634 vdd.n1539 vdd.n1499 1.16414
R5635 vdd.n1532 vdd.n1531 1.16414
R5636 vdd.n1395 vdd.n1355 1.16414
R5637 vdd.n1388 vdd.n1387 1.16414
R5638 vdd.n1446 vdd.n1406 1.16414
R5639 vdd.n1439 vdd.n1438 1.16414
R5640 vdd.n1659 vdd.t16 1.02079
R5641 vdd.t152 vdd.t182 1.02079
R5642 vdd.t183 vdd.t110 1.02079
R5643 vdd.n3154 vdd.t82 1.02079
R5644 vdd.n1636 vdd.n28 1.00834
R5645 vdd vdd.n3350 1.0005
R5646 vdd.n1193 vdd.n1192 0.970197
R5647 vdd.n1915 vdd.n1914 0.970197
R5648 vdd.n3206 vdd.n3205 0.970197
R5649 vdd.n2994 vdd.n2992 0.970197
R5650 vdd.t218 vdd.n820 0.907421
R5651 vdd.n774 vdd.t206 0.907421
R5652 vdd.t6 vdd.n1017 0.794056
R5653 vdd.n1686 vdd.t117 0.794056
R5654 vdd.t186 vdd.n895 0.794056
R5655 vdd.n867 vdd.t184 0.794056
R5656 vdd.t174 vdd.n733 0.794056
R5657 vdd.n705 vdd.t211 0.794056
R5658 vdd.t95 vdd.n511 0.794056
R5659 vdd.n481 vdd.t35 0.794056
R5660 vdd.n1336 vdd.t23 0.567326
R5661 vdd.n3338 vdd.t21 0.567326
R5662 vdd.n1905 vdd.n1904 0.509646
R5663 vdd.n3119 vdd.n3118 0.509646
R5664 vdd.n3317 vdd.n3316 0.509646
R5665 vdd.n3199 vdd.n3198 0.509646
R5666 vdd.n3125 vdd.n514 0.509646
R5667 vdd.n1681 vdd.n975 0.509646
R5668 vdd.n1298 vdd.n1060 0.509646
R5669 vdd.n1292 vdd.n1291 0.509646
R5670 vdd.n4 vdd.n2 0.459552
R5671 vdd.n11 vdd.n9 0.459552
R5672 vdd.n305 vdd.n304 0.388379
R5673 vdd.n271 vdd.n269 0.388379
R5674 vdd.n254 vdd.n253 0.388379
R5675 vdd.n220 vdd.n218 0.388379
R5676 vdd.n211 vdd.n210 0.388379
R5677 vdd.n177 vdd.n175 0.388379
R5678 vdd.n160 vdd.n159 0.388379
R5679 vdd.n126 vdd.n124 0.388379
R5680 vdd.n118 vdd.n117 0.388379
R5681 vdd.n84 vdd.n82 0.388379
R5682 vdd.n67 vdd.n66 0.388379
R5683 vdd.n33 vdd.n31 0.388379
R5684 vdd.n1580 vdd.n1579 0.388379
R5685 vdd.n1546 vdd.n1544 0.388379
R5686 vdd.n1631 vdd.n1630 0.388379
R5687 vdd.n1597 vdd.n1595 0.388379
R5688 vdd.n1486 vdd.n1485 0.388379
R5689 vdd.n1452 vdd.n1450 0.388379
R5690 vdd.n1537 vdd.n1536 0.388379
R5691 vdd.n1503 vdd.n1501 0.388379
R5692 vdd.n1393 vdd.n1392 0.388379
R5693 vdd.n1359 vdd.n1357 0.388379
R5694 vdd.n1444 vdd.n1443 0.388379
R5695 vdd.n1410 vdd.n1408 0.388379
R5696 vdd.n19 vdd.n17 0.387128
R5697 vdd.n24 vdd.n22 0.387128
R5698 vdd.n6 vdd.n4 0.358259
R5699 vdd.n13 vdd.n11 0.358259
R5700 vdd.n260 vdd.n258 0.358259
R5701 vdd.n262 vdd.n260 0.358259
R5702 vdd.n264 vdd.n262 0.358259
R5703 vdd.n266 vdd.n264 0.358259
R5704 vdd.n308 vdd.n266 0.358259
R5705 vdd.n166 vdd.n164 0.358259
R5706 vdd.n168 vdd.n166 0.358259
R5707 vdd.n170 vdd.n168 0.358259
R5708 vdd.n172 vdd.n170 0.358259
R5709 vdd.n214 vdd.n172 0.358259
R5710 vdd.n73 vdd.n71 0.358259
R5711 vdd.n75 vdd.n73 0.358259
R5712 vdd.n77 vdd.n75 0.358259
R5713 vdd.n79 vdd.n77 0.358259
R5714 vdd.n121 vdd.n79 0.358259
R5715 vdd.n1634 vdd.n1592 0.358259
R5716 vdd.n1592 vdd.n1590 0.358259
R5717 vdd.n1590 vdd.n1588 0.358259
R5718 vdd.n1588 vdd.n1586 0.358259
R5719 vdd.n1586 vdd.n1584 0.358259
R5720 vdd.n1540 vdd.n1498 0.358259
R5721 vdd.n1498 vdd.n1496 0.358259
R5722 vdd.n1496 vdd.n1494 0.358259
R5723 vdd.n1494 vdd.n1492 0.358259
R5724 vdd.n1492 vdd.n1490 0.358259
R5725 vdd.n1447 vdd.n1405 0.358259
R5726 vdd.n1405 vdd.n1403 0.358259
R5727 vdd.n1403 vdd.n1401 0.358259
R5728 vdd.n1401 vdd.n1399 0.358259
R5729 vdd.n1399 vdd.n1397 0.358259
R5730 vdd.t31 vdd.n1046 0.340595
R5731 vdd.n3329 vdd.t0 0.340595
R5732 vdd.n14 vdd.n6 0.334552
R5733 vdd.n14 vdd.n13 0.334552
R5734 vdd.n27 vdd.n19 0.21707
R5735 vdd.n27 vdd.n24 0.21707
R5736 vdd.n306 vdd.n268 0.155672
R5737 vdd.n298 vdd.n268 0.155672
R5738 vdd.n298 vdd.n297 0.155672
R5739 vdd.n297 vdd.n273 0.155672
R5740 vdd.n290 vdd.n273 0.155672
R5741 vdd.n290 vdd.n289 0.155672
R5742 vdd.n289 vdd.n277 0.155672
R5743 vdd.n282 vdd.n277 0.155672
R5744 vdd.n255 vdd.n217 0.155672
R5745 vdd.n247 vdd.n217 0.155672
R5746 vdd.n247 vdd.n246 0.155672
R5747 vdd.n246 vdd.n222 0.155672
R5748 vdd.n239 vdd.n222 0.155672
R5749 vdd.n239 vdd.n238 0.155672
R5750 vdd.n238 vdd.n226 0.155672
R5751 vdd.n231 vdd.n226 0.155672
R5752 vdd.n212 vdd.n174 0.155672
R5753 vdd.n204 vdd.n174 0.155672
R5754 vdd.n204 vdd.n203 0.155672
R5755 vdd.n203 vdd.n179 0.155672
R5756 vdd.n196 vdd.n179 0.155672
R5757 vdd.n196 vdd.n195 0.155672
R5758 vdd.n195 vdd.n183 0.155672
R5759 vdd.n188 vdd.n183 0.155672
R5760 vdd.n161 vdd.n123 0.155672
R5761 vdd.n153 vdd.n123 0.155672
R5762 vdd.n153 vdd.n152 0.155672
R5763 vdd.n152 vdd.n128 0.155672
R5764 vdd.n145 vdd.n128 0.155672
R5765 vdd.n145 vdd.n144 0.155672
R5766 vdd.n144 vdd.n132 0.155672
R5767 vdd.n137 vdd.n132 0.155672
R5768 vdd.n119 vdd.n81 0.155672
R5769 vdd.n111 vdd.n81 0.155672
R5770 vdd.n111 vdd.n110 0.155672
R5771 vdd.n110 vdd.n86 0.155672
R5772 vdd.n103 vdd.n86 0.155672
R5773 vdd.n103 vdd.n102 0.155672
R5774 vdd.n102 vdd.n90 0.155672
R5775 vdd.n95 vdd.n90 0.155672
R5776 vdd.n68 vdd.n30 0.155672
R5777 vdd.n60 vdd.n30 0.155672
R5778 vdd.n60 vdd.n59 0.155672
R5779 vdd.n59 vdd.n35 0.155672
R5780 vdd.n52 vdd.n35 0.155672
R5781 vdd.n52 vdd.n51 0.155672
R5782 vdd.n51 vdd.n39 0.155672
R5783 vdd.n44 vdd.n39 0.155672
R5784 vdd.n1581 vdd.n1543 0.155672
R5785 vdd.n1573 vdd.n1543 0.155672
R5786 vdd.n1573 vdd.n1572 0.155672
R5787 vdd.n1572 vdd.n1548 0.155672
R5788 vdd.n1565 vdd.n1548 0.155672
R5789 vdd.n1565 vdd.n1564 0.155672
R5790 vdd.n1564 vdd.n1552 0.155672
R5791 vdd.n1557 vdd.n1552 0.155672
R5792 vdd.n1632 vdd.n1594 0.155672
R5793 vdd.n1624 vdd.n1594 0.155672
R5794 vdd.n1624 vdd.n1623 0.155672
R5795 vdd.n1623 vdd.n1599 0.155672
R5796 vdd.n1616 vdd.n1599 0.155672
R5797 vdd.n1616 vdd.n1615 0.155672
R5798 vdd.n1615 vdd.n1603 0.155672
R5799 vdd.n1608 vdd.n1603 0.155672
R5800 vdd.n1487 vdd.n1449 0.155672
R5801 vdd.n1479 vdd.n1449 0.155672
R5802 vdd.n1479 vdd.n1478 0.155672
R5803 vdd.n1478 vdd.n1454 0.155672
R5804 vdd.n1471 vdd.n1454 0.155672
R5805 vdd.n1471 vdd.n1470 0.155672
R5806 vdd.n1470 vdd.n1458 0.155672
R5807 vdd.n1463 vdd.n1458 0.155672
R5808 vdd.n1538 vdd.n1500 0.155672
R5809 vdd.n1530 vdd.n1500 0.155672
R5810 vdd.n1530 vdd.n1529 0.155672
R5811 vdd.n1529 vdd.n1505 0.155672
R5812 vdd.n1522 vdd.n1505 0.155672
R5813 vdd.n1522 vdd.n1521 0.155672
R5814 vdd.n1521 vdd.n1509 0.155672
R5815 vdd.n1514 vdd.n1509 0.155672
R5816 vdd.n1394 vdd.n1356 0.155672
R5817 vdd.n1386 vdd.n1356 0.155672
R5818 vdd.n1386 vdd.n1385 0.155672
R5819 vdd.n1385 vdd.n1361 0.155672
R5820 vdd.n1378 vdd.n1361 0.155672
R5821 vdd.n1378 vdd.n1377 0.155672
R5822 vdd.n1377 vdd.n1365 0.155672
R5823 vdd.n1370 vdd.n1365 0.155672
R5824 vdd.n1445 vdd.n1407 0.155672
R5825 vdd.n1437 vdd.n1407 0.155672
R5826 vdd.n1437 vdd.n1436 0.155672
R5827 vdd.n1436 vdd.n1412 0.155672
R5828 vdd.n1429 vdd.n1412 0.155672
R5829 vdd.n1429 vdd.n1428 0.155672
R5830 vdd.n1428 vdd.n1416 0.155672
R5831 vdd.n1421 vdd.n1416 0.155672
R5832 vdd.n1893 vdd.n1698 0.152939
R5833 vdd.n1704 vdd.n1698 0.152939
R5834 vdd.n1705 vdd.n1704 0.152939
R5835 vdd.n1706 vdd.n1705 0.152939
R5836 vdd.n1707 vdd.n1706 0.152939
R5837 vdd.n1711 vdd.n1707 0.152939
R5838 vdd.n1712 vdd.n1711 0.152939
R5839 vdd.n1713 vdd.n1712 0.152939
R5840 vdd.n1714 vdd.n1713 0.152939
R5841 vdd.n1718 vdd.n1714 0.152939
R5842 vdd.n1719 vdd.n1718 0.152939
R5843 vdd.n1720 vdd.n1719 0.152939
R5844 vdd.n1868 vdd.n1720 0.152939
R5845 vdd.n1868 vdd.n1867 0.152939
R5846 vdd.n1867 vdd.n1866 0.152939
R5847 vdd.n1866 vdd.n1726 0.152939
R5848 vdd.n1731 vdd.n1726 0.152939
R5849 vdd.n1732 vdd.n1731 0.152939
R5850 vdd.n1733 vdd.n1732 0.152939
R5851 vdd.n1737 vdd.n1733 0.152939
R5852 vdd.n1738 vdd.n1737 0.152939
R5853 vdd.n1739 vdd.n1738 0.152939
R5854 vdd.n1740 vdd.n1739 0.152939
R5855 vdd.n1744 vdd.n1740 0.152939
R5856 vdd.n1745 vdd.n1744 0.152939
R5857 vdd.n1746 vdd.n1745 0.152939
R5858 vdd.n1747 vdd.n1746 0.152939
R5859 vdd.n1751 vdd.n1747 0.152939
R5860 vdd.n1752 vdd.n1751 0.152939
R5861 vdd.n1753 vdd.n1752 0.152939
R5862 vdd.n1754 vdd.n1753 0.152939
R5863 vdd.n1758 vdd.n1754 0.152939
R5864 vdd.n1759 vdd.n1758 0.152939
R5865 vdd.n1760 vdd.n1759 0.152939
R5866 vdd.n1829 vdd.n1760 0.152939
R5867 vdd.n1829 vdd.n1828 0.152939
R5868 vdd.n1828 vdd.n1827 0.152939
R5869 vdd.n1827 vdd.n1766 0.152939
R5870 vdd.n1771 vdd.n1766 0.152939
R5871 vdd.n1772 vdd.n1771 0.152939
R5872 vdd.n1773 vdd.n1772 0.152939
R5873 vdd.n1777 vdd.n1773 0.152939
R5874 vdd.n1778 vdd.n1777 0.152939
R5875 vdd.n1779 vdd.n1778 0.152939
R5876 vdd.n1780 vdd.n1779 0.152939
R5877 vdd.n1784 vdd.n1780 0.152939
R5878 vdd.n1785 vdd.n1784 0.152939
R5879 vdd.n1786 vdd.n1785 0.152939
R5880 vdd.n1787 vdd.n1786 0.152939
R5881 vdd.n1788 vdd.n1787 0.152939
R5882 vdd.n1788 vdd.n972 0.152939
R5883 vdd.n1904 vdd.n1692 0.152939
R5884 vdd.n1639 vdd.n1638 0.152939
R5885 vdd.n1639 vdd.n1008 0.152939
R5886 vdd.n1654 vdd.n1008 0.152939
R5887 vdd.n1655 vdd.n1654 0.152939
R5888 vdd.n1656 vdd.n1655 0.152939
R5889 vdd.n1656 vdd.n997 0.152939
R5890 vdd.n1671 vdd.n997 0.152939
R5891 vdd.n1672 vdd.n1671 0.152939
R5892 vdd.n1673 vdd.n1672 0.152939
R5893 vdd.n1673 vdd.n985 0.152939
R5894 vdd.n1690 vdd.n985 0.152939
R5895 vdd.n1691 vdd.n1690 0.152939
R5896 vdd.n1905 vdd.n1691 0.152939
R5897 vdd.n527 vdd.n524 0.152939
R5898 vdd.n528 vdd.n527 0.152939
R5899 vdd.n529 vdd.n528 0.152939
R5900 vdd.n530 vdd.n529 0.152939
R5901 vdd.n533 vdd.n530 0.152939
R5902 vdd.n534 vdd.n533 0.152939
R5903 vdd.n535 vdd.n534 0.152939
R5904 vdd.n536 vdd.n535 0.152939
R5905 vdd.n539 vdd.n536 0.152939
R5906 vdd.n540 vdd.n539 0.152939
R5907 vdd.n541 vdd.n540 0.152939
R5908 vdd.n542 vdd.n541 0.152939
R5909 vdd.n547 vdd.n542 0.152939
R5910 vdd.n548 vdd.n547 0.152939
R5911 vdd.n549 vdd.n548 0.152939
R5912 vdd.n550 vdd.n549 0.152939
R5913 vdd.n553 vdd.n550 0.152939
R5914 vdd.n554 vdd.n553 0.152939
R5915 vdd.n555 vdd.n554 0.152939
R5916 vdd.n556 vdd.n555 0.152939
R5917 vdd.n559 vdd.n556 0.152939
R5918 vdd.n560 vdd.n559 0.152939
R5919 vdd.n561 vdd.n560 0.152939
R5920 vdd.n562 vdd.n561 0.152939
R5921 vdd.n565 vdd.n562 0.152939
R5922 vdd.n566 vdd.n565 0.152939
R5923 vdd.n567 vdd.n566 0.152939
R5924 vdd.n568 vdd.n567 0.152939
R5925 vdd.n571 vdd.n568 0.152939
R5926 vdd.n572 vdd.n571 0.152939
R5927 vdd.n573 vdd.n572 0.152939
R5928 vdd.n574 vdd.n573 0.152939
R5929 vdd.n577 vdd.n574 0.152939
R5930 vdd.n578 vdd.n577 0.152939
R5931 vdd.n3035 vdd.n578 0.152939
R5932 vdd.n3035 vdd.n3034 0.152939
R5933 vdd.n3034 vdd.n3033 0.152939
R5934 vdd.n3033 vdd.n582 0.152939
R5935 vdd.n587 vdd.n582 0.152939
R5936 vdd.n588 vdd.n587 0.152939
R5937 vdd.n591 vdd.n588 0.152939
R5938 vdd.n592 vdd.n591 0.152939
R5939 vdd.n593 vdd.n592 0.152939
R5940 vdd.n594 vdd.n593 0.152939
R5941 vdd.n597 vdd.n594 0.152939
R5942 vdd.n598 vdd.n597 0.152939
R5943 vdd.n599 vdd.n598 0.152939
R5944 vdd.n600 vdd.n599 0.152939
R5945 vdd.n603 vdd.n600 0.152939
R5946 vdd.n604 vdd.n603 0.152939
R5947 vdd.n605 vdd.n604 0.152939
R5948 vdd.n3118 vdd.n518 0.152939
R5949 vdd.n3119 vdd.n508 0.152939
R5950 vdd.n3133 vdd.n508 0.152939
R5951 vdd.n3134 vdd.n3133 0.152939
R5952 vdd.n3135 vdd.n3134 0.152939
R5953 vdd.n3135 vdd.n496 0.152939
R5954 vdd.n3149 vdd.n496 0.152939
R5955 vdd.n3150 vdd.n3149 0.152939
R5956 vdd.n3151 vdd.n3150 0.152939
R5957 vdd.n3151 vdd.n484 0.152939
R5958 vdd.n3166 vdd.n484 0.152939
R5959 vdd.n3167 vdd.n3166 0.152939
R5960 vdd.n3168 vdd.n3167 0.152939
R5961 vdd.n3168 vdd.n310 0.152939
R5962 vdd.n320 vdd.n311 0.152939
R5963 vdd.n321 vdd.n320 0.152939
R5964 vdd.n322 vdd.n321 0.152939
R5965 vdd.n331 vdd.n322 0.152939
R5966 vdd.n332 vdd.n331 0.152939
R5967 vdd.n333 vdd.n332 0.152939
R5968 vdd.n334 vdd.n333 0.152939
R5969 vdd.n342 vdd.n334 0.152939
R5970 vdd.n343 vdd.n342 0.152939
R5971 vdd.n344 vdd.n343 0.152939
R5972 vdd.n345 vdd.n344 0.152939
R5973 vdd.n353 vdd.n345 0.152939
R5974 vdd.n3317 vdd.n353 0.152939
R5975 vdd.n3316 vdd.n354 0.152939
R5976 vdd.n357 vdd.n354 0.152939
R5977 vdd.n361 vdd.n357 0.152939
R5978 vdd.n362 vdd.n361 0.152939
R5979 vdd.n363 vdd.n362 0.152939
R5980 vdd.n364 vdd.n363 0.152939
R5981 vdd.n365 vdd.n364 0.152939
R5982 vdd.n369 vdd.n365 0.152939
R5983 vdd.n370 vdd.n369 0.152939
R5984 vdd.n371 vdd.n370 0.152939
R5985 vdd.n372 vdd.n371 0.152939
R5986 vdd.n376 vdd.n372 0.152939
R5987 vdd.n377 vdd.n376 0.152939
R5988 vdd.n378 vdd.n377 0.152939
R5989 vdd.n379 vdd.n378 0.152939
R5990 vdd.n383 vdd.n379 0.152939
R5991 vdd.n384 vdd.n383 0.152939
R5992 vdd.n385 vdd.n384 0.152939
R5993 vdd.n3282 vdd.n385 0.152939
R5994 vdd.n3282 vdd.n3281 0.152939
R5995 vdd.n3281 vdd.n3280 0.152939
R5996 vdd.n3280 vdd.n391 0.152939
R5997 vdd.n396 vdd.n391 0.152939
R5998 vdd.n397 vdd.n396 0.152939
R5999 vdd.n398 vdd.n397 0.152939
R6000 vdd.n402 vdd.n398 0.152939
R6001 vdd.n403 vdd.n402 0.152939
R6002 vdd.n404 vdd.n403 0.152939
R6003 vdd.n405 vdd.n404 0.152939
R6004 vdd.n409 vdd.n405 0.152939
R6005 vdd.n410 vdd.n409 0.152939
R6006 vdd.n411 vdd.n410 0.152939
R6007 vdd.n412 vdd.n411 0.152939
R6008 vdd.n416 vdd.n412 0.152939
R6009 vdd.n417 vdd.n416 0.152939
R6010 vdd.n418 vdd.n417 0.152939
R6011 vdd.n419 vdd.n418 0.152939
R6012 vdd.n423 vdd.n419 0.152939
R6013 vdd.n424 vdd.n423 0.152939
R6014 vdd.n425 vdd.n424 0.152939
R6015 vdd.n3243 vdd.n425 0.152939
R6016 vdd.n3243 vdd.n3242 0.152939
R6017 vdd.n3242 vdd.n3241 0.152939
R6018 vdd.n3241 vdd.n431 0.152939
R6019 vdd.n436 vdd.n431 0.152939
R6020 vdd.n437 vdd.n436 0.152939
R6021 vdd.n438 vdd.n437 0.152939
R6022 vdd.n442 vdd.n438 0.152939
R6023 vdd.n443 vdd.n442 0.152939
R6024 vdd.n444 vdd.n443 0.152939
R6025 vdd.n445 vdd.n444 0.152939
R6026 vdd.n449 vdd.n445 0.152939
R6027 vdd.n450 vdd.n449 0.152939
R6028 vdd.n451 vdd.n450 0.152939
R6029 vdd.n452 vdd.n451 0.152939
R6030 vdd.n456 vdd.n452 0.152939
R6031 vdd.n457 vdd.n456 0.152939
R6032 vdd.n458 vdd.n457 0.152939
R6033 vdd.n459 vdd.n458 0.152939
R6034 vdd.n463 vdd.n459 0.152939
R6035 vdd.n464 vdd.n463 0.152939
R6036 vdd.n465 vdd.n464 0.152939
R6037 vdd.n3199 vdd.n465 0.152939
R6038 vdd.n3126 vdd.n3125 0.152939
R6039 vdd.n3127 vdd.n3126 0.152939
R6040 vdd.n3127 vdd.n502 0.152939
R6041 vdd.n3141 vdd.n502 0.152939
R6042 vdd.n3142 vdd.n3141 0.152939
R6043 vdd.n3143 vdd.n3142 0.152939
R6044 vdd.n3143 vdd.n489 0.152939
R6045 vdd.n3157 vdd.n489 0.152939
R6046 vdd.n3158 vdd.n3157 0.152939
R6047 vdd.n3159 vdd.n3158 0.152939
R6048 vdd.n3159 vdd.n477 0.152939
R6049 vdd.n3174 vdd.n477 0.152939
R6050 vdd.n3175 vdd.n3174 0.152939
R6051 vdd.n3176 vdd.n3175 0.152939
R6052 vdd.n3176 vdd.n475 0.152939
R6053 vdd.n3180 vdd.n475 0.152939
R6054 vdd.n3181 vdd.n3180 0.152939
R6055 vdd.n3182 vdd.n3181 0.152939
R6056 vdd.n3182 vdd.n472 0.152939
R6057 vdd.n3186 vdd.n472 0.152939
R6058 vdd.n3187 vdd.n3186 0.152939
R6059 vdd.n3188 vdd.n3187 0.152939
R6060 vdd.n3188 vdd.n469 0.152939
R6061 vdd.n3192 vdd.n469 0.152939
R6062 vdd.n3193 vdd.n3192 0.152939
R6063 vdd.n3194 vdd.n3193 0.152939
R6064 vdd.n3194 vdd.n466 0.152939
R6065 vdd.n3198 vdd.n466 0.152939
R6066 vdd.n2988 vdd.n514 0.152939
R6067 vdd.n1916 vdd.n975 0.152939
R6068 vdd.n1299 vdd.n1298 0.152939
R6069 vdd.n1300 vdd.n1299 0.152939
R6070 vdd.n1300 vdd.n1049 0.152939
R6071 vdd.n1314 vdd.n1049 0.152939
R6072 vdd.n1315 vdd.n1314 0.152939
R6073 vdd.n1316 vdd.n1315 0.152939
R6074 vdd.n1316 vdd.n1036 0.152939
R6075 vdd.n1330 vdd.n1036 0.152939
R6076 vdd.n1331 vdd.n1330 0.152939
R6077 vdd.n1332 vdd.n1331 0.152939
R6078 vdd.n1332 vdd.n1025 0.152939
R6079 vdd.n1347 vdd.n1025 0.152939
R6080 vdd.n1348 vdd.n1347 0.152939
R6081 vdd.n1349 vdd.n1348 0.152939
R6082 vdd.n1349 vdd.n1014 0.152939
R6083 vdd.n1645 vdd.n1014 0.152939
R6084 vdd.n1646 vdd.n1645 0.152939
R6085 vdd.n1647 vdd.n1646 0.152939
R6086 vdd.n1647 vdd.n1002 0.152939
R6087 vdd.n1662 vdd.n1002 0.152939
R6088 vdd.n1663 vdd.n1662 0.152939
R6089 vdd.n1664 vdd.n1663 0.152939
R6090 vdd.n1664 vdd.n992 0.152939
R6091 vdd.n1679 vdd.n992 0.152939
R6092 vdd.n1680 vdd.n1679 0.152939
R6093 vdd.n1683 vdd.n1680 0.152939
R6094 vdd.n1683 vdd.n1682 0.152939
R6095 vdd.n1682 vdd.n1681 0.152939
R6096 vdd.n1291 vdd.n1065 0.152939
R6097 vdd.n1287 vdd.n1065 0.152939
R6098 vdd.n1287 vdd.n1286 0.152939
R6099 vdd.n1286 vdd.n1285 0.152939
R6100 vdd.n1285 vdd.n1070 0.152939
R6101 vdd.n1281 vdd.n1070 0.152939
R6102 vdd.n1281 vdd.n1280 0.152939
R6103 vdd.n1280 vdd.n1279 0.152939
R6104 vdd.n1279 vdd.n1078 0.152939
R6105 vdd.n1275 vdd.n1078 0.152939
R6106 vdd.n1275 vdd.n1274 0.152939
R6107 vdd.n1274 vdd.n1273 0.152939
R6108 vdd.n1273 vdd.n1086 0.152939
R6109 vdd.n1269 vdd.n1086 0.152939
R6110 vdd.n1269 vdd.n1268 0.152939
R6111 vdd.n1268 vdd.n1267 0.152939
R6112 vdd.n1267 vdd.n1094 0.152939
R6113 vdd.n1263 vdd.n1094 0.152939
R6114 vdd.n1263 vdd.n1262 0.152939
R6115 vdd.n1262 vdd.n1261 0.152939
R6116 vdd.n1261 vdd.n1104 0.152939
R6117 vdd.n1257 vdd.n1104 0.152939
R6118 vdd.n1257 vdd.n1256 0.152939
R6119 vdd.n1256 vdd.n1255 0.152939
R6120 vdd.n1255 vdd.n1112 0.152939
R6121 vdd.n1251 vdd.n1112 0.152939
R6122 vdd.n1251 vdd.n1250 0.152939
R6123 vdd.n1250 vdd.n1249 0.152939
R6124 vdd.n1249 vdd.n1120 0.152939
R6125 vdd.n1245 vdd.n1120 0.152939
R6126 vdd.n1245 vdd.n1244 0.152939
R6127 vdd.n1244 vdd.n1243 0.152939
R6128 vdd.n1243 vdd.n1128 0.152939
R6129 vdd.n1239 vdd.n1128 0.152939
R6130 vdd.n1239 vdd.n1238 0.152939
R6131 vdd.n1238 vdd.n1237 0.152939
R6132 vdd.n1237 vdd.n1136 0.152939
R6133 vdd.n1233 vdd.n1136 0.152939
R6134 vdd.n1233 vdd.n1232 0.152939
R6135 vdd.n1232 vdd.n1231 0.152939
R6136 vdd.n1231 vdd.n1144 0.152939
R6137 vdd.n1151 vdd.n1144 0.152939
R6138 vdd.n1221 vdd.n1151 0.152939
R6139 vdd.n1221 vdd.n1220 0.152939
R6140 vdd.n1220 vdd.n1219 0.152939
R6141 vdd.n1219 vdd.n1152 0.152939
R6142 vdd.n1215 vdd.n1152 0.152939
R6143 vdd.n1215 vdd.n1214 0.152939
R6144 vdd.n1214 vdd.n1213 0.152939
R6145 vdd.n1213 vdd.n1159 0.152939
R6146 vdd.n1209 vdd.n1159 0.152939
R6147 vdd.n1209 vdd.n1208 0.152939
R6148 vdd.n1208 vdd.n1207 0.152939
R6149 vdd.n1207 vdd.n1167 0.152939
R6150 vdd.n1203 vdd.n1167 0.152939
R6151 vdd.n1203 vdd.n1202 0.152939
R6152 vdd.n1202 vdd.n1201 0.152939
R6153 vdd.n1201 vdd.n1175 0.152939
R6154 vdd.n1197 vdd.n1175 0.152939
R6155 vdd.n1197 vdd.n1196 0.152939
R6156 vdd.n1196 vdd.n1195 0.152939
R6157 vdd.n1195 vdd.n1183 0.152939
R6158 vdd.n1183 vdd.n1060 0.152939
R6159 vdd.n1292 vdd.n1055 0.152939
R6160 vdd.n1306 vdd.n1055 0.152939
R6161 vdd.n1307 vdd.n1306 0.152939
R6162 vdd.n1308 vdd.n1307 0.152939
R6163 vdd.n1308 vdd.n1043 0.152939
R6164 vdd.n1322 vdd.n1043 0.152939
R6165 vdd.n1323 vdd.n1322 0.152939
R6166 vdd.n1324 vdd.n1323 0.152939
R6167 vdd.n1324 vdd.n1031 0.152939
R6168 vdd.n1339 vdd.n1031 0.152939
R6169 vdd.n1340 vdd.n1339 0.152939
R6170 vdd.n1341 vdd.n1340 0.152939
R6171 vdd.n1341 vdd.n1020 0.152939
R6172 vdd.n1638 vdd.n1637 0.145814
R6173 vdd.n3349 vdd.n310 0.145814
R6174 vdd.n3349 vdd.n311 0.145814
R6175 vdd.n1637 vdd.n1020 0.145814
R6176 vdd.n2203 vdd.t223 0.113865
R6177 vdd.n2270 vdd.t175 0.113865
R6178 vdd.n2753 vdd.t178 0.113865
R6179 vdd.n2820 vdd.t202 0.113865
R6180 vdd.n1894 vdd.n1692 0.110256
R6181 vdd.n2919 vdd.n518 0.110256
R6182 vdd.n2988 vdd.n2987 0.110256
R6183 vdd.n1917 vdd.n1916 0.110256
R6184 vdd.n1894 vdd.n1893 0.0431829
R6185 vdd.n1917 vdd.n972 0.0431829
R6186 vdd.n2919 vdd.n524 0.0431829
R6187 vdd.n2987 vdd.n605 0.0431829
R6188 vdd vdd.n28 0.00833333
R6189 a_n7636_8799.n137 a_n7636_8799.t50 490.524
R6190 a_n7636_8799.n148 a_n7636_8799.t56 490.524
R6191 a_n7636_8799.n160 a_n7636_8799.t79 490.524
R6192 a_n7636_8799.n103 a_n7636_8799.t95 490.524
R6193 a_n7636_8799.n114 a_n7636_8799.t107 490.524
R6194 a_n7636_8799.n126 a_n7636_8799.t77 490.524
R6195 a_n7636_8799.n31 a_n7636_8799.t73 484.3
R6196 a_n7636_8799.n143 a_n7636_8799.t38 464.166
R6197 a_n7636_8799.n142 a_n7636_8799.t75 464.166
R6198 a_n7636_8799.n133 a_n7636_8799.t74 464.166
R6199 a_n7636_8799.n141 a_n7636_8799.t40 464.166
R6200 a_n7636_8799.n140 a_n7636_8799.t39 464.166
R6201 a_n7636_8799.n134 a_n7636_8799.t88 464.166
R6202 a_n7636_8799.n139 a_n7636_8799.t49 464.166
R6203 a_n7636_8799.n138 a_n7636_8799.t41 464.166
R6204 a_n7636_8799.n135 a_n7636_8799.t92 464.166
R6205 a_n7636_8799.n136 a_n7636_8799.t64 464.166
R6206 a_n7636_8799.n40 a_n7636_8799.t83 484.3
R6207 a_n7636_8799.n154 a_n7636_8799.t43 464.166
R6208 a_n7636_8799.n153 a_n7636_8799.t86 464.166
R6209 a_n7636_8799.n144 a_n7636_8799.t84 464.166
R6210 a_n7636_8799.n152 a_n7636_8799.t45 464.166
R6211 a_n7636_8799.n151 a_n7636_8799.t44 464.166
R6212 a_n7636_8799.n145 a_n7636_8799.t101 464.166
R6213 a_n7636_8799.n150 a_n7636_8799.t55 464.166
R6214 a_n7636_8799.n149 a_n7636_8799.t46 464.166
R6215 a_n7636_8799.n146 a_n7636_8799.t102 464.166
R6216 a_n7636_8799.n147 a_n7636_8799.t72 464.166
R6217 a_n7636_8799.n49 a_n7636_8799.t52 484.3
R6218 a_n7636_8799.n166 a_n7636_8799.t105 464.166
R6219 a_n7636_8799.n165 a_n7636_8799.t82 464.166
R6220 a_n7636_8799.n156 a_n7636_8799.t99 464.166
R6221 a_n7636_8799.n164 a_n7636_8799.t70 464.166
R6222 a_n7636_8799.n163 a_n7636_8799.t85 464.166
R6223 a_n7636_8799.n157 a_n7636_8799.t47 464.166
R6224 a_n7636_8799.n162 a_n7636_8799.t97 464.166
R6225 a_n7636_8799.n161 a_n7636_8799.t58 464.166
R6226 a_n7636_8799.n158 a_n7636_8799.t93 464.166
R6227 a_n7636_8799.n159 a_n7636_8799.t51 464.166
R6228 a_n7636_8799.n102 a_n7636_8799.t96 464.166
R6229 a_n7636_8799.n101 a_n7636_8799.t63 464.166
R6230 a_n7636_8799.n104 a_n7636_8799.t81 464.166
R6231 a_n7636_8799.n100 a_n7636_8799.t94 464.166
R6232 a_n7636_8799.n105 a_n7636_8799.t61 464.166
R6233 a_n7636_8799.n106 a_n7636_8799.t62 464.166
R6234 a_n7636_8799.n99 a_n7636_8799.t78 464.166
R6235 a_n7636_8799.n107 a_n7636_8799.t54 464.166
R6236 a_n7636_8799.n98 a_n7636_8799.t53 464.166
R6237 a_n7636_8799.n108 a_n7636_8799.t76 464.166
R6238 a_n7636_8799.n113 a_n7636_8799.t106 464.166
R6239 a_n7636_8799.n112 a_n7636_8799.t69 464.166
R6240 a_n7636_8799.n115 a_n7636_8799.t90 464.166
R6241 a_n7636_8799.n111 a_n7636_8799.t104 464.166
R6242 a_n7636_8799.n116 a_n7636_8799.t68 464.166
R6243 a_n7636_8799.n117 a_n7636_8799.t67 464.166
R6244 a_n7636_8799.n110 a_n7636_8799.t89 464.166
R6245 a_n7636_8799.n118 a_n7636_8799.t57 464.166
R6246 a_n7636_8799.n109 a_n7636_8799.t60 464.166
R6247 a_n7636_8799.n119 a_n7636_8799.t87 464.166
R6248 a_n7636_8799.n125 a_n7636_8799.t65 464.166
R6249 a_n7636_8799.n124 a_n7636_8799.t91 464.166
R6250 a_n7636_8799.n127 a_n7636_8799.t59 464.166
R6251 a_n7636_8799.n123 a_n7636_8799.t98 464.166
R6252 a_n7636_8799.n128 a_n7636_8799.t48 464.166
R6253 a_n7636_8799.n129 a_n7636_8799.t37 464.166
R6254 a_n7636_8799.n122 a_n7636_8799.t71 464.166
R6255 a_n7636_8799.n130 a_n7636_8799.t100 464.166
R6256 a_n7636_8799.n121 a_n7636_8799.t80 464.166
R6257 a_n7636_8799.n131 a_n7636_8799.t103 464.166
R6258 a_n7636_8799.n39 a_n7636_8799.n38 75.3623
R6259 a_n7636_8799.n37 a_n7636_8799.n23 70.3058
R6260 a_n7636_8799.n23 a_n7636_8799.n36 70.1674
R6261 a_n7636_8799.n36 a_n7636_8799.n134 20.9683
R6262 a_n7636_8799.n35 a_n7636_8799.n24 75.0448
R6263 a_n7636_8799.n140 a_n7636_8799.n35 11.2134
R6264 a_n7636_8799.n34 a_n7636_8799.n24 80.4688
R6265 a_n7636_8799.n26 a_n7636_8799.n33 74.73
R6266 a_n7636_8799.n32 a_n7636_8799.n26 70.1674
R6267 a_n7636_8799.n143 a_n7636_8799.n32 20.9683
R6268 a_n7636_8799.n25 a_n7636_8799.n31 70.5844
R6269 a_n7636_8799.n48 a_n7636_8799.n47 75.3623
R6270 a_n7636_8799.n46 a_n7636_8799.n19 70.3058
R6271 a_n7636_8799.n19 a_n7636_8799.n45 70.1674
R6272 a_n7636_8799.n45 a_n7636_8799.n145 20.9683
R6273 a_n7636_8799.n44 a_n7636_8799.n20 75.0448
R6274 a_n7636_8799.n151 a_n7636_8799.n44 11.2134
R6275 a_n7636_8799.n43 a_n7636_8799.n20 80.4688
R6276 a_n7636_8799.n22 a_n7636_8799.n42 74.73
R6277 a_n7636_8799.n41 a_n7636_8799.n22 70.1674
R6278 a_n7636_8799.n154 a_n7636_8799.n41 20.9683
R6279 a_n7636_8799.n21 a_n7636_8799.n40 70.5844
R6280 a_n7636_8799.n57 a_n7636_8799.n56 75.3623
R6281 a_n7636_8799.n55 a_n7636_8799.n15 70.3058
R6282 a_n7636_8799.n15 a_n7636_8799.n54 70.1674
R6283 a_n7636_8799.n54 a_n7636_8799.n157 20.9683
R6284 a_n7636_8799.n53 a_n7636_8799.n16 75.0448
R6285 a_n7636_8799.n163 a_n7636_8799.n53 11.2134
R6286 a_n7636_8799.n52 a_n7636_8799.n16 80.4688
R6287 a_n7636_8799.n18 a_n7636_8799.n51 74.73
R6288 a_n7636_8799.n50 a_n7636_8799.n18 70.1674
R6289 a_n7636_8799.n166 a_n7636_8799.n50 20.9683
R6290 a_n7636_8799.n17 a_n7636_8799.n49 70.5844
R6291 a_n7636_8799.n11 a_n7636_8799.n66 70.5844
R6292 a_n7636_8799.n65 a_n7636_8799.n12 70.1674
R6293 a_n7636_8799.n65 a_n7636_8799.n98 20.9683
R6294 a_n7636_8799.n12 a_n7636_8799.n64 74.73
R6295 a_n7636_8799.n107 a_n7636_8799.n64 11.843
R6296 a_n7636_8799.n63 a_n7636_8799.n13 80.4688
R6297 a_n7636_8799.n63 a_n7636_8799.n99 0.365327
R6298 a_n7636_8799.n13 a_n7636_8799.n62 75.0448
R6299 a_n7636_8799.n61 a_n7636_8799.n14 70.1674
R6300 a_n7636_8799.n61 a_n7636_8799.n100 20.9683
R6301 a_n7636_8799.n14 a_n7636_8799.n60 70.3058
R6302 a_n7636_8799.n104 a_n7636_8799.n60 20.6913
R6303 a_n7636_8799.n59 a_n7636_8799.n58 75.3623
R6304 a_n7636_8799.n7 a_n7636_8799.n75 70.5844
R6305 a_n7636_8799.n74 a_n7636_8799.n8 70.1674
R6306 a_n7636_8799.n74 a_n7636_8799.n109 20.9683
R6307 a_n7636_8799.n8 a_n7636_8799.n73 74.73
R6308 a_n7636_8799.n118 a_n7636_8799.n73 11.843
R6309 a_n7636_8799.n72 a_n7636_8799.n9 80.4688
R6310 a_n7636_8799.n72 a_n7636_8799.n110 0.365327
R6311 a_n7636_8799.n9 a_n7636_8799.n71 75.0448
R6312 a_n7636_8799.n70 a_n7636_8799.n10 70.1674
R6313 a_n7636_8799.n70 a_n7636_8799.n111 20.9683
R6314 a_n7636_8799.n10 a_n7636_8799.n69 70.3058
R6315 a_n7636_8799.n115 a_n7636_8799.n69 20.6913
R6316 a_n7636_8799.n68 a_n7636_8799.n67 75.3623
R6317 a_n7636_8799.n3 a_n7636_8799.n84 70.5844
R6318 a_n7636_8799.n83 a_n7636_8799.n4 70.1674
R6319 a_n7636_8799.n83 a_n7636_8799.n121 20.9683
R6320 a_n7636_8799.n4 a_n7636_8799.n82 74.73
R6321 a_n7636_8799.n130 a_n7636_8799.n82 11.843
R6322 a_n7636_8799.n81 a_n7636_8799.n5 80.4688
R6323 a_n7636_8799.n81 a_n7636_8799.n122 0.365327
R6324 a_n7636_8799.n5 a_n7636_8799.n80 75.0448
R6325 a_n7636_8799.n79 a_n7636_8799.n6 70.1674
R6326 a_n7636_8799.n79 a_n7636_8799.n123 20.9683
R6327 a_n7636_8799.n6 a_n7636_8799.n78 70.3058
R6328 a_n7636_8799.n127 a_n7636_8799.n78 20.6913
R6329 a_n7636_8799.n77 a_n7636_8799.n76 75.3623
R6330 a_n7636_8799.n27 a_n7636_8799.n85 98.9633
R6331 a_n7636_8799.n30 a_n7636_8799.n174 98.9631
R6332 a_n7636_8799.n30 a_n7636_8799.n173 98.6055
R6333 a_n7636_8799.n29 a_n7636_8799.n172 98.6055
R6334 a_n7636_8799.n29 a_n7636_8799.n171 98.6055
R6335 a_n7636_8799.n28 a_n7636_8799.n89 98.6055
R6336 a_n7636_8799.n28 a_n7636_8799.n88 98.6055
R6337 a_n7636_8799.n27 a_n7636_8799.n87 98.6055
R6338 a_n7636_8799.n27 a_n7636_8799.n86 98.6055
R6339 a_n7636_8799.n175 a_n7636_8799.n30 98.6054
R6340 a_n7636_8799.n1 a_n7636_8799.n90 81.4626
R6341 a_n7636_8799.n2 a_n7636_8799.n94 81.4626
R6342 a_n7636_8799.n2 a_n7636_8799.n92 81.4626
R6343 a_n7636_8799.n0 a_n7636_8799.n96 80.9324
R6344 a_n7636_8799.n1 a_n7636_8799.n97 80.9324
R6345 a_n7636_8799.n1 a_n7636_8799.n91 80.9324
R6346 a_n7636_8799.n2 a_n7636_8799.n95 80.9324
R6347 a_n7636_8799.n2 a_n7636_8799.n93 80.9324
R6348 a_n7636_8799.n32 a_n7636_8799.n142 20.9683
R6349 a_n7636_8799.n141 a_n7636_8799.n140 48.2005
R6350 a_n7636_8799.n139 a_n7636_8799.n36 20.9683
R6351 a_n7636_8799.n136 a_n7636_8799.n135 48.2005
R6352 a_n7636_8799.n41 a_n7636_8799.n153 20.9683
R6353 a_n7636_8799.n152 a_n7636_8799.n151 48.2005
R6354 a_n7636_8799.n150 a_n7636_8799.n45 20.9683
R6355 a_n7636_8799.n147 a_n7636_8799.n146 48.2005
R6356 a_n7636_8799.n50 a_n7636_8799.n165 20.9683
R6357 a_n7636_8799.n164 a_n7636_8799.n163 48.2005
R6358 a_n7636_8799.n162 a_n7636_8799.n54 20.9683
R6359 a_n7636_8799.n159 a_n7636_8799.n158 48.2005
R6360 a_n7636_8799.n102 a_n7636_8799.n101 48.2005
R6361 a_n7636_8799.n105 a_n7636_8799.n61 20.9683
R6362 a_n7636_8799.n106 a_n7636_8799.n99 48.2005
R6363 a_n7636_8799.n108 a_n7636_8799.n65 20.9683
R6364 a_n7636_8799.n113 a_n7636_8799.n112 48.2005
R6365 a_n7636_8799.n116 a_n7636_8799.n70 20.9683
R6366 a_n7636_8799.n117 a_n7636_8799.n110 48.2005
R6367 a_n7636_8799.n119 a_n7636_8799.n74 20.9683
R6368 a_n7636_8799.n125 a_n7636_8799.n124 48.2005
R6369 a_n7636_8799.n128 a_n7636_8799.n79 20.9683
R6370 a_n7636_8799.n129 a_n7636_8799.n122 48.2005
R6371 a_n7636_8799.n131 a_n7636_8799.n83 20.9683
R6372 a_n7636_8799.n34 a_n7636_8799.n133 47.835
R6373 a_n7636_8799.n37 a_n7636_8799.n138 20.6913
R6374 a_n7636_8799.n43 a_n7636_8799.n144 47.835
R6375 a_n7636_8799.n46 a_n7636_8799.n149 20.6913
R6376 a_n7636_8799.n52 a_n7636_8799.n156 47.835
R6377 a_n7636_8799.n55 a_n7636_8799.n161 20.6913
R6378 a_n7636_8799.n100 a_n7636_8799.n60 21.4216
R6379 a_n7636_8799.n111 a_n7636_8799.n69 21.4216
R6380 a_n7636_8799.n123 a_n7636_8799.n78 21.4216
R6381 a_n7636_8799.t36 a_n7636_8799.n66 484.3
R6382 a_n7636_8799.t42 a_n7636_8799.n75 484.3
R6383 a_n7636_8799.t66 a_n7636_8799.n84 484.3
R6384 a_n7636_8799.n59 a_n7636_8799.n103 45.0871
R6385 a_n7636_8799.n68 a_n7636_8799.n114 45.0871
R6386 a_n7636_8799.n77 a_n7636_8799.n126 45.0871
R6387 a_n7636_8799.n39 a_n7636_8799.n137 45.0871
R6388 a_n7636_8799.n48 a_n7636_8799.n148 45.0871
R6389 a_n7636_8799.n57 a_n7636_8799.n160 45.0871
R6390 a_n7636_8799.n29 a_n7636_8799.n170 32.8105
R6391 a_n7636_8799.n33 a_n7636_8799.n133 11.843
R6392 a_n7636_8799.n138 a_n7636_8799.n38 36.139
R6393 a_n7636_8799.n42 a_n7636_8799.n144 11.843
R6394 a_n7636_8799.n149 a_n7636_8799.n47 36.139
R6395 a_n7636_8799.n51 a_n7636_8799.n156 11.843
R6396 a_n7636_8799.n161 a_n7636_8799.n56 36.139
R6397 a_n7636_8799.n104 a_n7636_8799.n58 36.139
R6398 a_n7636_8799.n98 a_n7636_8799.n64 34.4824
R6399 a_n7636_8799.n115 a_n7636_8799.n67 36.139
R6400 a_n7636_8799.n109 a_n7636_8799.n73 34.4824
R6401 a_n7636_8799.n127 a_n7636_8799.n76 36.139
R6402 a_n7636_8799.n121 a_n7636_8799.n82 34.4824
R6403 a_n7636_8799.n35 a_n7636_8799.n134 35.3134
R6404 a_n7636_8799.n44 a_n7636_8799.n145 35.3134
R6405 a_n7636_8799.n53 a_n7636_8799.n157 35.3134
R6406 a_n7636_8799.n62 a_n7636_8799.n105 35.3134
R6407 a_n7636_8799.n106 a_n7636_8799.n62 11.2134
R6408 a_n7636_8799.n71 a_n7636_8799.n116 35.3134
R6409 a_n7636_8799.n117 a_n7636_8799.n71 11.2134
R6410 a_n7636_8799.n80 a_n7636_8799.n128 35.3134
R6411 a_n7636_8799.n129 a_n7636_8799.n80 11.2134
R6412 a_n7636_8799.n142 a_n7636_8799.n33 34.4824
R6413 a_n7636_8799.n38 a_n7636_8799.n135 10.5784
R6414 a_n7636_8799.n153 a_n7636_8799.n42 34.4824
R6415 a_n7636_8799.n47 a_n7636_8799.n146 10.5784
R6416 a_n7636_8799.n165 a_n7636_8799.n51 34.4824
R6417 a_n7636_8799.n56 a_n7636_8799.n158 10.5784
R6418 a_n7636_8799.n58 a_n7636_8799.n101 10.5784
R6419 a_n7636_8799.n67 a_n7636_8799.n112 10.5784
R6420 a_n7636_8799.n76 a_n7636_8799.n124 10.5784
R6421 a_n7636_8799.n170 a_n7636_8799.n28 19.9322
R6422 a_n7636_8799.n137 a_n7636_8799.n136 14.1472
R6423 a_n7636_8799.n148 a_n7636_8799.n147 14.1472
R6424 a_n7636_8799.n160 a_n7636_8799.n159 14.1472
R6425 a_n7636_8799.n103 a_n7636_8799.n102 14.1472
R6426 a_n7636_8799.n114 a_n7636_8799.n113 14.1472
R6427 a_n7636_8799.n126 a_n7636_8799.n125 14.1472
R6428 a_n7636_8799.n169 a_n7636_8799.n1 12.3339
R6429 a_n7636_8799.n170 a_n7636_8799.n169 11.4887
R6430 a_n7636_8799.n155 a_n7636_8799.n25 9.01755
R6431 a_n7636_8799.n120 a_n7636_8799.n11 9.01755
R6432 a_n7636_8799.n168 a_n7636_8799.n132 7.07069
R6433 a_n7636_8799.n168 a_n7636_8799.n167 6.72822
R6434 a_n7636_8799.n155 a_n7636_8799.n21 4.90959
R6435 a_n7636_8799.n167 a_n7636_8799.n17 4.90959
R6436 a_n7636_8799.n120 a_n7636_8799.n7 4.90959
R6437 a_n7636_8799.n132 a_n7636_8799.n3 4.90959
R6438 a_n7636_8799.n167 a_n7636_8799.n155 4.10845
R6439 a_n7636_8799.n132 a_n7636_8799.n120 4.10845
R6440 a_n7636_8799.n174 a_n7636_8799.t22 3.61217
R6441 a_n7636_8799.n174 a_n7636_8799.t26 3.61217
R6442 a_n7636_8799.n173 a_n7636_8799.t18 3.61217
R6443 a_n7636_8799.n173 a_n7636_8799.t30 3.61217
R6444 a_n7636_8799.n172 a_n7636_8799.t21 3.61217
R6445 a_n7636_8799.n172 a_n7636_8799.t16 3.61217
R6446 a_n7636_8799.n171 a_n7636_8799.t29 3.61217
R6447 a_n7636_8799.n171 a_n7636_8799.t33 3.61217
R6448 a_n7636_8799.n89 a_n7636_8799.t25 3.61217
R6449 a_n7636_8799.n89 a_n7636_8799.t24 3.61217
R6450 a_n7636_8799.n88 a_n7636_8799.t17 3.61217
R6451 a_n7636_8799.n88 a_n7636_8799.t20 3.61217
R6452 a_n7636_8799.n87 a_n7636_8799.t23 3.61217
R6453 a_n7636_8799.n87 a_n7636_8799.t28 3.61217
R6454 a_n7636_8799.n86 a_n7636_8799.t27 3.61217
R6455 a_n7636_8799.n86 a_n7636_8799.t15 3.61217
R6456 a_n7636_8799.n85 a_n7636_8799.t31 3.61217
R6457 a_n7636_8799.n85 a_n7636_8799.t19 3.61217
R6458 a_n7636_8799.t14 a_n7636_8799.n175 3.61217
R6459 a_n7636_8799.n175 a_n7636_8799.t32 3.61217
R6460 a_n7636_8799.n169 a_n7636_8799.n168 3.4105
R6461 a_n7636_8799.n96 a_n7636_8799.t7 2.82907
R6462 a_n7636_8799.n96 a_n7636_8799.t9 2.82907
R6463 a_n7636_8799.n97 a_n7636_8799.t6 2.82907
R6464 a_n7636_8799.n97 a_n7636_8799.t5 2.82907
R6465 a_n7636_8799.n91 a_n7636_8799.t10 2.82907
R6466 a_n7636_8799.n91 a_n7636_8799.t2 2.82907
R6467 a_n7636_8799.n90 a_n7636_8799.t0 2.82907
R6468 a_n7636_8799.n90 a_n7636_8799.t35 2.82907
R6469 a_n7636_8799.n94 a_n7636_8799.t34 2.82907
R6470 a_n7636_8799.n94 a_n7636_8799.t12 2.82907
R6471 a_n7636_8799.n95 a_n7636_8799.t11 2.82907
R6472 a_n7636_8799.n95 a_n7636_8799.t13 2.82907
R6473 a_n7636_8799.n93 a_n7636_8799.t3 2.82907
R6474 a_n7636_8799.n93 a_n7636_8799.t4 2.82907
R6475 a_n7636_8799.n92 a_n7636_8799.t1 2.82907
R6476 a_n7636_8799.n92 a_n7636_8799.t8 2.82907
R6477 a_n7636_8799.n31 a_n7636_8799.n143 22.3251
R6478 a_n7636_8799.n40 a_n7636_8799.n154 22.3251
R6479 a_n7636_8799.n49 a_n7636_8799.n166 22.3251
R6480 a_n7636_8799.n66 a_n7636_8799.n108 22.3251
R6481 a_n7636_8799.n75 a_n7636_8799.n119 22.3251
R6482 a_n7636_8799.n84 a_n7636_8799.n131 22.3251
R6483 a_n7636_8799.n34 a_n7636_8799.n141 0.365327
R6484 a_n7636_8799.n139 a_n7636_8799.n37 21.4216
R6485 a_n7636_8799.n43 a_n7636_8799.n152 0.365327
R6486 a_n7636_8799.n150 a_n7636_8799.n46 21.4216
R6487 a_n7636_8799.n52 a_n7636_8799.n164 0.365327
R6488 a_n7636_8799.n162 a_n7636_8799.n55 21.4216
R6489 a_n7636_8799.n107 a_n7636_8799.n63 47.835
R6490 a_n7636_8799.n118 a_n7636_8799.n72 47.835
R6491 a_n7636_8799.n130 a_n7636_8799.n81 47.835
R6492 a_n7636_8799.n0 a_n7636_8799.n2 33.2634
R6493 a_n7636_8799.n30 a_n7636_8799.n29 1.07378
R6494 a_n7636_8799.n28 a_n7636_8799.n27 1.07378
R6495 a_n7636_8799.n1 a_n7636_8799.n0 1.06084
R6496 a_n7636_8799.n26 a_n7636_8799.n24 0.758076
R6497 a_n7636_8799.n24 a_n7636_8799.n23 0.758076
R6498 a_n7636_8799.n39 a_n7636_8799.n23 0.758076
R6499 a_n7636_8799.n22 a_n7636_8799.n20 0.758076
R6500 a_n7636_8799.n20 a_n7636_8799.n19 0.758076
R6501 a_n7636_8799.n48 a_n7636_8799.n19 0.758076
R6502 a_n7636_8799.n18 a_n7636_8799.n16 0.758076
R6503 a_n7636_8799.n16 a_n7636_8799.n15 0.758076
R6504 a_n7636_8799.n57 a_n7636_8799.n15 0.758076
R6505 a_n7636_8799.n14 a_n7636_8799.n13 0.758076
R6506 a_n7636_8799.n13 a_n7636_8799.n12 0.758076
R6507 a_n7636_8799.n12 a_n7636_8799.n11 0.758076
R6508 a_n7636_8799.n10 a_n7636_8799.n9 0.758076
R6509 a_n7636_8799.n9 a_n7636_8799.n8 0.758076
R6510 a_n7636_8799.n8 a_n7636_8799.n7 0.758076
R6511 a_n7636_8799.n6 a_n7636_8799.n5 0.758076
R6512 a_n7636_8799.n5 a_n7636_8799.n4 0.758076
R6513 a_n7636_8799.n4 a_n7636_8799.n3 0.758076
R6514 a_n7636_8799.n77 a_n7636_8799.n6 0.568682
R6515 a_n7636_8799.n68 a_n7636_8799.n10 0.568682
R6516 a_n7636_8799.n59 a_n7636_8799.n14 0.568682
R6517 a_n7636_8799.n18 a_n7636_8799.n17 0.568682
R6518 a_n7636_8799.n22 a_n7636_8799.n21 0.568682
R6519 a_n7636_8799.n26 a_n7636_8799.n25 0.568682
R6520 CSoutput.n19 CSoutput.t161 184.661
R6521 CSoutput.n78 CSoutput.n77 165.8
R6522 CSoutput.n76 CSoutput.n0 165.8
R6523 CSoutput.n75 CSoutput.n74 165.8
R6524 CSoutput.n73 CSoutput.n72 165.8
R6525 CSoutput.n71 CSoutput.n2 165.8
R6526 CSoutput.n69 CSoutput.n68 165.8
R6527 CSoutput.n67 CSoutput.n3 165.8
R6528 CSoutput.n66 CSoutput.n65 165.8
R6529 CSoutput.n63 CSoutput.n4 165.8
R6530 CSoutput.n61 CSoutput.n60 165.8
R6531 CSoutput.n59 CSoutput.n5 165.8
R6532 CSoutput.n58 CSoutput.n57 165.8
R6533 CSoutput.n55 CSoutput.n6 165.8
R6534 CSoutput.n54 CSoutput.n53 165.8
R6535 CSoutput.n52 CSoutput.n51 165.8
R6536 CSoutput.n50 CSoutput.n8 165.8
R6537 CSoutput.n48 CSoutput.n47 165.8
R6538 CSoutput.n46 CSoutput.n9 165.8
R6539 CSoutput.n45 CSoutput.n44 165.8
R6540 CSoutput.n42 CSoutput.n10 165.8
R6541 CSoutput.n41 CSoutput.n40 165.8
R6542 CSoutput.n39 CSoutput.n38 165.8
R6543 CSoutput.n37 CSoutput.n12 165.8
R6544 CSoutput.n35 CSoutput.n34 165.8
R6545 CSoutput.n33 CSoutput.n13 165.8
R6546 CSoutput.n32 CSoutput.n31 165.8
R6547 CSoutput.n29 CSoutput.n14 165.8
R6548 CSoutput.n28 CSoutput.n27 165.8
R6549 CSoutput.n26 CSoutput.n25 165.8
R6550 CSoutput.n24 CSoutput.n16 165.8
R6551 CSoutput.n22 CSoutput.n21 165.8
R6552 CSoutput.n20 CSoutput.n17 165.8
R6553 CSoutput.n77 CSoutput.t164 162.194
R6554 CSoutput.n18 CSoutput.t150 120.501
R6555 CSoutput.n23 CSoutput.t152 120.501
R6556 CSoutput.n15 CSoutput.t165 120.501
R6557 CSoutput.n30 CSoutput.t153 120.501
R6558 CSoutput.n36 CSoutput.t156 120.501
R6559 CSoutput.n11 CSoutput.t149 120.501
R6560 CSoutput.n43 CSoutput.t160 120.501
R6561 CSoutput.n49 CSoutput.t157 120.501
R6562 CSoutput.n7 CSoutput.t151 120.501
R6563 CSoutput.n56 CSoutput.t147 120.501
R6564 CSoutput.n62 CSoutput.t158 120.501
R6565 CSoutput.n64 CSoutput.t159 120.501
R6566 CSoutput.n70 CSoutput.t148 120.501
R6567 CSoutput.n1 CSoutput.t145 120.501
R6568 CSoutput.n290 CSoutput.n288 103.469
R6569 CSoutput.n278 CSoutput.n276 103.469
R6570 CSoutput.n267 CSoutput.n265 103.469
R6571 CSoutput.n104 CSoutput.n102 103.469
R6572 CSoutput.n92 CSoutput.n90 103.469
R6573 CSoutput.n81 CSoutput.n79 103.469
R6574 CSoutput.n296 CSoutput.n295 103.111
R6575 CSoutput.n294 CSoutput.n293 103.111
R6576 CSoutput.n292 CSoutput.n291 103.111
R6577 CSoutput.n290 CSoutput.n289 103.111
R6578 CSoutput.n286 CSoutput.n285 103.111
R6579 CSoutput.n284 CSoutput.n283 103.111
R6580 CSoutput.n282 CSoutput.n281 103.111
R6581 CSoutput.n280 CSoutput.n279 103.111
R6582 CSoutput.n278 CSoutput.n277 103.111
R6583 CSoutput.n275 CSoutput.n274 103.111
R6584 CSoutput.n273 CSoutput.n272 103.111
R6585 CSoutput.n271 CSoutput.n270 103.111
R6586 CSoutput.n269 CSoutput.n268 103.111
R6587 CSoutput.n267 CSoutput.n266 103.111
R6588 CSoutput.n104 CSoutput.n103 103.111
R6589 CSoutput.n106 CSoutput.n105 103.111
R6590 CSoutput.n108 CSoutput.n107 103.111
R6591 CSoutput.n110 CSoutput.n109 103.111
R6592 CSoutput.n112 CSoutput.n111 103.111
R6593 CSoutput.n92 CSoutput.n91 103.111
R6594 CSoutput.n94 CSoutput.n93 103.111
R6595 CSoutput.n96 CSoutput.n95 103.111
R6596 CSoutput.n98 CSoutput.n97 103.111
R6597 CSoutput.n100 CSoutput.n99 103.111
R6598 CSoutput.n81 CSoutput.n80 103.111
R6599 CSoutput.n83 CSoutput.n82 103.111
R6600 CSoutput.n85 CSoutput.n84 103.111
R6601 CSoutput.n87 CSoutput.n86 103.111
R6602 CSoutput.n89 CSoutput.n88 103.111
R6603 CSoutput.n298 CSoutput.n297 103.111
R6604 CSoutput.n326 CSoutput.n324 81.5057
R6605 CSoutput.n314 CSoutput.n312 81.5057
R6606 CSoutput.n303 CSoutput.n301 81.5057
R6607 CSoutput.n362 CSoutput.n360 81.5057
R6608 CSoutput.n350 CSoutput.n348 81.5057
R6609 CSoutput.n339 CSoutput.n337 81.5057
R6610 CSoutput.n334 CSoutput.n333 80.9324
R6611 CSoutput.n332 CSoutput.n331 80.9324
R6612 CSoutput.n330 CSoutput.n329 80.9324
R6613 CSoutput.n328 CSoutput.n327 80.9324
R6614 CSoutput.n326 CSoutput.n325 80.9324
R6615 CSoutput.n322 CSoutput.n321 80.9324
R6616 CSoutput.n320 CSoutput.n319 80.9324
R6617 CSoutput.n318 CSoutput.n317 80.9324
R6618 CSoutput.n316 CSoutput.n315 80.9324
R6619 CSoutput.n314 CSoutput.n313 80.9324
R6620 CSoutput.n311 CSoutput.n310 80.9324
R6621 CSoutput.n309 CSoutput.n308 80.9324
R6622 CSoutput.n307 CSoutput.n306 80.9324
R6623 CSoutput.n305 CSoutput.n304 80.9324
R6624 CSoutput.n303 CSoutput.n302 80.9324
R6625 CSoutput.n362 CSoutput.n361 80.9324
R6626 CSoutput.n364 CSoutput.n363 80.9324
R6627 CSoutput.n366 CSoutput.n365 80.9324
R6628 CSoutput.n368 CSoutput.n367 80.9324
R6629 CSoutput.n370 CSoutput.n369 80.9324
R6630 CSoutput.n350 CSoutput.n349 80.9324
R6631 CSoutput.n352 CSoutput.n351 80.9324
R6632 CSoutput.n354 CSoutput.n353 80.9324
R6633 CSoutput.n356 CSoutput.n355 80.9324
R6634 CSoutput.n358 CSoutput.n357 80.9324
R6635 CSoutput.n339 CSoutput.n338 80.9324
R6636 CSoutput.n341 CSoutput.n340 80.9324
R6637 CSoutput.n343 CSoutput.n342 80.9324
R6638 CSoutput.n345 CSoutput.n344 80.9324
R6639 CSoutput.n347 CSoutput.n346 80.9324
R6640 CSoutput.n25 CSoutput.n24 48.1486
R6641 CSoutput.n69 CSoutput.n3 48.1486
R6642 CSoutput.n38 CSoutput.n37 48.1486
R6643 CSoutput.n42 CSoutput.n41 48.1486
R6644 CSoutput.n51 CSoutput.n50 48.1486
R6645 CSoutput.n55 CSoutput.n54 48.1486
R6646 CSoutput.n22 CSoutput.n17 46.462
R6647 CSoutput.n72 CSoutput.n71 46.462
R6648 CSoutput.n20 CSoutput.n19 44.9055
R6649 CSoutput.n29 CSoutput.n28 43.7635
R6650 CSoutput.n65 CSoutput.n63 43.7635
R6651 CSoutput.n35 CSoutput.n13 41.7396
R6652 CSoutput.n57 CSoutput.n5 41.7396
R6653 CSoutput.n44 CSoutput.n9 37.0171
R6654 CSoutput.n48 CSoutput.n9 37.0171
R6655 CSoutput.n76 CSoutput.n75 34.9932
R6656 CSoutput.n31 CSoutput.n13 32.2947
R6657 CSoutput.n61 CSoutput.n5 32.2947
R6658 CSoutput.n30 CSoutput.n29 29.6014
R6659 CSoutput.n63 CSoutput.n62 29.6014
R6660 CSoutput.n19 CSoutput.n18 28.4085
R6661 CSoutput.n18 CSoutput.n17 25.1176
R6662 CSoutput.n72 CSoutput.n1 25.1176
R6663 CSoutput.n43 CSoutput.n42 22.0922
R6664 CSoutput.n50 CSoutput.n49 22.0922
R6665 CSoutput.n77 CSoutput.n76 21.8586
R6666 CSoutput.n37 CSoutput.n36 18.9681
R6667 CSoutput.n56 CSoutput.n55 18.9681
R6668 CSoutput.n25 CSoutput.n15 17.6292
R6669 CSoutput.n64 CSoutput.n3 17.6292
R6670 CSoutput.n24 CSoutput.n23 15.844
R6671 CSoutput.n70 CSoutput.n69 15.844
R6672 CSoutput.n38 CSoutput.n11 14.5051
R6673 CSoutput.n54 CSoutput.n7 14.5051
R6674 CSoutput.n373 CSoutput.n78 11.4982
R6675 CSoutput.n41 CSoutput.n11 11.3811
R6676 CSoutput.n51 CSoutput.n7 11.3811
R6677 CSoutput.n23 CSoutput.n22 10.0422
R6678 CSoutput.n71 CSoutput.n70 10.0422
R6679 CSoutput.n287 CSoutput.n275 9.25285
R6680 CSoutput.n101 CSoutput.n89 9.25285
R6681 CSoutput.n323 CSoutput.n311 8.98182
R6682 CSoutput.n359 CSoutput.n347 8.98182
R6683 CSoutput.n336 CSoutput.n300 8.76129
R6684 CSoutput.n28 CSoutput.n15 8.25698
R6685 CSoutput.n65 CSoutput.n64 8.25698
R6686 CSoutput.n300 CSoutput.n299 7.12641
R6687 CSoutput.n114 CSoutput.n113 7.12641
R6688 CSoutput.n36 CSoutput.n35 6.91809
R6689 CSoutput.n57 CSoutput.n56 6.91809
R6690 CSoutput.n336 CSoutput.n335 6.02792
R6691 CSoutput.n372 CSoutput.n371 6.02792
R6692 CSoutput.n335 CSoutput.n334 5.25266
R6693 CSoutput.n323 CSoutput.n322 5.25266
R6694 CSoutput.n371 CSoutput.n370 5.25266
R6695 CSoutput.n359 CSoutput.n358 5.25266
R6696 CSoutput.n373 CSoutput.n114 5.16885
R6697 CSoutput.n299 CSoutput.n298 5.1449
R6698 CSoutput.n287 CSoutput.n286 5.1449
R6699 CSoutput.n113 CSoutput.n112 5.1449
R6700 CSoutput.n101 CSoutput.n100 5.1449
R6701 CSoutput.n205 CSoutput.n158 4.5005
R6702 CSoutput.n174 CSoutput.n158 4.5005
R6703 CSoutput.n169 CSoutput.n153 4.5005
R6704 CSoutput.n169 CSoutput.n155 4.5005
R6705 CSoutput.n169 CSoutput.n152 4.5005
R6706 CSoutput.n169 CSoutput.n156 4.5005
R6707 CSoutput.n169 CSoutput.n151 4.5005
R6708 CSoutput.n169 CSoutput.t162 4.5005
R6709 CSoutput.n169 CSoutput.n150 4.5005
R6710 CSoutput.n169 CSoutput.n157 4.5005
R6711 CSoutput.n169 CSoutput.n158 4.5005
R6712 CSoutput.n167 CSoutput.n153 4.5005
R6713 CSoutput.n167 CSoutput.n155 4.5005
R6714 CSoutput.n167 CSoutput.n152 4.5005
R6715 CSoutput.n167 CSoutput.n156 4.5005
R6716 CSoutput.n167 CSoutput.n151 4.5005
R6717 CSoutput.n167 CSoutput.t162 4.5005
R6718 CSoutput.n167 CSoutput.n150 4.5005
R6719 CSoutput.n167 CSoutput.n157 4.5005
R6720 CSoutput.n167 CSoutput.n158 4.5005
R6721 CSoutput.n166 CSoutput.n153 4.5005
R6722 CSoutput.n166 CSoutput.n155 4.5005
R6723 CSoutput.n166 CSoutput.n152 4.5005
R6724 CSoutput.n166 CSoutput.n156 4.5005
R6725 CSoutput.n166 CSoutput.n151 4.5005
R6726 CSoutput.n166 CSoutput.t162 4.5005
R6727 CSoutput.n166 CSoutput.n150 4.5005
R6728 CSoutput.n166 CSoutput.n157 4.5005
R6729 CSoutput.n166 CSoutput.n158 4.5005
R6730 CSoutput.n251 CSoutput.n153 4.5005
R6731 CSoutput.n251 CSoutput.n155 4.5005
R6732 CSoutput.n251 CSoutput.n152 4.5005
R6733 CSoutput.n251 CSoutput.n156 4.5005
R6734 CSoutput.n251 CSoutput.n151 4.5005
R6735 CSoutput.n251 CSoutput.t162 4.5005
R6736 CSoutput.n251 CSoutput.n150 4.5005
R6737 CSoutput.n251 CSoutput.n157 4.5005
R6738 CSoutput.n251 CSoutput.n158 4.5005
R6739 CSoutput.n249 CSoutput.n153 4.5005
R6740 CSoutput.n249 CSoutput.n155 4.5005
R6741 CSoutput.n249 CSoutput.n152 4.5005
R6742 CSoutput.n249 CSoutput.n156 4.5005
R6743 CSoutput.n249 CSoutput.n151 4.5005
R6744 CSoutput.n249 CSoutput.t162 4.5005
R6745 CSoutput.n249 CSoutput.n150 4.5005
R6746 CSoutput.n249 CSoutput.n157 4.5005
R6747 CSoutput.n247 CSoutput.n153 4.5005
R6748 CSoutput.n247 CSoutput.n155 4.5005
R6749 CSoutput.n247 CSoutput.n152 4.5005
R6750 CSoutput.n247 CSoutput.n156 4.5005
R6751 CSoutput.n247 CSoutput.n151 4.5005
R6752 CSoutput.n247 CSoutput.t162 4.5005
R6753 CSoutput.n247 CSoutput.n150 4.5005
R6754 CSoutput.n247 CSoutput.n157 4.5005
R6755 CSoutput.n177 CSoutput.n153 4.5005
R6756 CSoutput.n177 CSoutput.n155 4.5005
R6757 CSoutput.n177 CSoutput.n152 4.5005
R6758 CSoutput.n177 CSoutput.n156 4.5005
R6759 CSoutput.n177 CSoutput.n151 4.5005
R6760 CSoutput.n177 CSoutput.t162 4.5005
R6761 CSoutput.n177 CSoutput.n150 4.5005
R6762 CSoutput.n177 CSoutput.n157 4.5005
R6763 CSoutput.n177 CSoutput.n158 4.5005
R6764 CSoutput.n176 CSoutput.n153 4.5005
R6765 CSoutput.n176 CSoutput.n155 4.5005
R6766 CSoutput.n176 CSoutput.n152 4.5005
R6767 CSoutput.n176 CSoutput.n156 4.5005
R6768 CSoutput.n176 CSoutput.n151 4.5005
R6769 CSoutput.n176 CSoutput.t162 4.5005
R6770 CSoutput.n176 CSoutput.n150 4.5005
R6771 CSoutput.n176 CSoutput.n157 4.5005
R6772 CSoutput.n176 CSoutput.n158 4.5005
R6773 CSoutput.n180 CSoutput.n153 4.5005
R6774 CSoutput.n180 CSoutput.n155 4.5005
R6775 CSoutput.n180 CSoutput.n152 4.5005
R6776 CSoutput.n180 CSoutput.n156 4.5005
R6777 CSoutput.n180 CSoutput.n151 4.5005
R6778 CSoutput.n180 CSoutput.t162 4.5005
R6779 CSoutput.n180 CSoutput.n150 4.5005
R6780 CSoutput.n180 CSoutput.n157 4.5005
R6781 CSoutput.n180 CSoutput.n158 4.5005
R6782 CSoutput.n179 CSoutput.n153 4.5005
R6783 CSoutput.n179 CSoutput.n155 4.5005
R6784 CSoutput.n179 CSoutput.n152 4.5005
R6785 CSoutput.n179 CSoutput.n156 4.5005
R6786 CSoutput.n179 CSoutput.n151 4.5005
R6787 CSoutput.n179 CSoutput.t162 4.5005
R6788 CSoutput.n179 CSoutput.n150 4.5005
R6789 CSoutput.n179 CSoutput.n157 4.5005
R6790 CSoutput.n179 CSoutput.n158 4.5005
R6791 CSoutput.n162 CSoutput.n153 4.5005
R6792 CSoutput.n162 CSoutput.n155 4.5005
R6793 CSoutput.n162 CSoutput.n152 4.5005
R6794 CSoutput.n162 CSoutput.n156 4.5005
R6795 CSoutput.n162 CSoutput.n151 4.5005
R6796 CSoutput.n162 CSoutput.t162 4.5005
R6797 CSoutput.n162 CSoutput.n150 4.5005
R6798 CSoutput.n162 CSoutput.n157 4.5005
R6799 CSoutput.n162 CSoutput.n158 4.5005
R6800 CSoutput.n254 CSoutput.n153 4.5005
R6801 CSoutput.n254 CSoutput.n155 4.5005
R6802 CSoutput.n254 CSoutput.n152 4.5005
R6803 CSoutput.n254 CSoutput.n156 4.5005
R6804 CSoutput.n254 CSoutput.n151 4.5005
R6805 CSoutput.n254 CSoutput.t162 4.5005
R6806 CSoutput.n254 CSoutput.n150 4.5005
R6807 CSoutput.n254 CSoutput.n157 4.5005
R6808 CSoutput.n254 CSoutput.n158 4.5005
R6809 CSoutput.n241 CSoutput.n212 4.5005
R6810 CSoutput.n241 CSoutput.n218 4.5005
R6811 CSoutput.n199 CSoutput.n188 4.5005
R6812 CSoutput.n199 CSoutput.n190 4.5005
R6813 CSoutput.n199 CSoutput.n187 4.5005
R6814 CSoutput.n199 CSoutput.n191 4.5005
R6815 CSoutput.n199 CSoutput.n186 4.5005
R6816 CSoutput.n199 CSoutput.t155 4.5005
R6817 CSoutput.n199 CSoutput.n185 4.5005
R6818 CSoutput.n199 CSoutput.n192 4.5005
R6819 CSoutput.n241 CSoutput.n199 4.5005
R6820 CSoutput.n220 CSoutput.n188 4.5005
R6821 CSoutput.n220 CSoutput.n190 4.5005
R6822 CSoutput.n220 CSoutput.n187 4.5005
R6823 CSoutput.n220 CSoutput.n191 4.5005
R6824 CSoutput.n220 CSoutput.n186 4.5005
R6825 CSoutput.n220 CSoutput.t155 4.5005
R6826 CSoutput.n220 CSoutput.n185 4.5005
R6827 CSoutput.n220 CSoutput.n192 4.5005
R6828 CSoutput.n241 CSoutput.n220 4.5005
R6829 CSoutput.n198 CSoutput.n188 4.5005
R6830 CSoutput.n198 CSoutput.n190 4.5005
R6831 CSoutput.n198 CSoutput.n187 4.5005
R6832 CSoutput.n198 CSoutput.n191 4.5005
R6833 CSoutput.n198 CSoutput.n186 4.5005
R6834 CSoutput.n198 CSoutput.t155 4.5005
R6835 CSoutput.n198 CSoutput.n185 4.5005
R6836 CSoutput.n198 CSoutput.n192 4.5005
R6837 CSoutput.n241 CSoutput.n198 4.5005
R6838 CSoutput.n222 CSoutput.n188 4.5005
R6839 CSoutput.n222 CSoutput.n190 4.5005
R6840 CSoutput.n222 CSoutput.n187 4.5005
R6841 CSoutput.n222 CSoutput.n191 4.5005
R6842 CSoutput.n222 CSoutput.n186 4.5005
R6843 CSoutput.n222 CSoutput.t155 4.5005
R6844 CSoutput.n222 CSoutput.n185 4.5005
R6845 CSoutput.n222 CSoutput.n192 4.5005
R6846 CSoutput.n241 CSoutput.n222 4.5005
R6847 CSoutput.n188 CSoutput.n183 4.5005
R6848 CSoutput.n190 CSoutput.n183 4.5005
R6849 CSoutput.n187 CSoutput.n183 4.5005
R6850 CSoutput.n191 CSoutput.n183 4.5005
R6851 CSoutput.n186 CSoutput.n183 4.5005
R6852 CSoutput.t155 CSoutput.n183 4.5005
R6853 CSoutput.n185 CSoutput.n183 4.5005
R6854 CSoutput.n192 CSoutput.n183 4.5005
R6855 CSoutput.n244 CSoutput.n188 4.5005
R6856 CSoutput.n244 CSoutput.n190 4.5005
R6857 CSoutput.n244 CSoutput.n187 4.5005
R6858 CSoutput.n244 CSoutput.n191 4.5005
R6859 CSoutput.n244 CSoutput.n186 4.5005
R6860 CSoutput.n244 CSoutput.t155 4.5005
R6861 CSoutput.n244 CSoutput.n185 4.5005
R6862 CSoutput.n244 CSoutput.n192 4.5005
R6863 CSoutput.n242 CSoutput.n188 4.5005
R6864 CSoutput.n242 CSoutput.n190 4.5005
R6865 CSoutput.n242 CSoutput.n187 4.5005
R6866 CSoutput.n242 CSoutput.n191 4.5005
R6867 CSoutput.n242 CSoutput.n186 4.5005
R6868 CSoutput.n242 CSoutput.t155 4.5005
R6869 CSoutput.n242 CSoutput.n185 4.5005
R6870 CSoutput.n242 CSoutput.n192 4.5005
R6871 CSoutput.n242 CSoutput.n241 4.5005
R6872 CSoutput.n224 CSoutput.n188 4.5005
R6873 CSoutput.n224 CSoutput.n190 4.5005
R6874 CSoutput.n224 CSoutput.n187 4.5005
R6875 CSoutput.n224 CSoutput.n191 4.5005
R6876 CSoutput.n224 CSoutput.n186 4.5005
R6877 CSoutput.n224 CSoutput.t155 4.5005
R6878 CSoutput.n224 CSoutput.n185 4.5005
R6879 CSoutput.n224 CSoutput.n192 4.5005
R6880 CSoutput.n241 CSoutput.n224 4.5005
R6881 CSoutput.n196 CSoutput.n188 4.5005
R6882 CSoutput.n196 CSoutput.n190 4.5005
R6883 CSoutput.n196 CSoutput.n187 4.5005
R6884 CSoutput.n196 CSoutput.n191 4.5005
R6885 CSoutput.n196 CSoutput.n186 4.5005
R6886 CSoutput.n196 CSoutput.t155 4.5005
R6887 CSoutput.n196 CSoutput.n185 4.5005
R6888 CSoutput.n196 CSoutput.n192 4.5005
R6889 CSoutput.n241 CSoutput.n196 4.5005
R6890 CSoutput.n226 CSoutput.n188 4.5005
R6891 CSoutput.n226 CSoutput.n190 4.5005
R6892 CSoutput.n226 CSoutput.n187 4.5005
R6893 CSoutput.n226 CSoutput.n191 4.5005
R6894 CSoutput.n226 CSoutput.n186 4.5005
R6895 CSoutput.n226 CSoutput.t155 4.5005
R6896 CSoutput.n226 CSoutput.n185 4.5005
R6897 CSoutput.n226 CSoutput.n192 4.5005
R6898 CSoutput.n241 CSoutput.n226 4.5005
R6899 CSoutput.n195 CSoutput.n188 4.5005
R6900 CSoutput.n195 CSoutput.n190 4.5005
R6901 CSoutput.n195 CSoutput.n187 4.5005
R6902 CSoutput.n195 CSoutput.n191 4.5005
R6903 CSoutput.n195 CSoutput.n186 4.5005
R6904 CSoutput.n195 CSoutput.t155 4.5005
R6905 CSoutput.n195 CSoutput.n185 4.5005
R6906 CSoutput.n195 CSoutput.n192 4.5005
R6907 CSoutput.n241 CSoutput.n195 4.5005
R6908 CSoutput.n240 CSoutput.n188 4.5005
R6909 CSoutput.n240 CSoutput.n190 4.5005
R6910 CSoutput.n240 CSoutput.n187 4.5005
R6911 CSoutput.n240 CSoutput.n191 4.5005
R6912 CSoutput.n240 CSoutput.n186 4.5005
R6913 CSoutput.n240 CSoutput.t155 4.5005
R6914 CSoutput.n240 CSoutput.n185 4.5005
R6915 CSoutput.n240 CSoutput.n192 4.5005
R6916 CSoutput.n241 CSoutput.n240 4.5005
R6917 CSoutput.n239 CSoutput.n124 4.5005
R6918 CSoutput.n140 CSoutput.n124 4.5005
R6919 CSoutput.n135 CSoutput.n119 4.5005
R6920 CSoutput.n135 CSoutput.n121 4.5005
R6921 CSoutput.n135 CSoutput.n118 4.5005
R6922 CSoutput.n135 CSoutput.n122 4.5005
R6923 CSoutput.n135 CSoutput.n117 4.5005
R6924 CSoutput.n135 CSoutput.t154 4.5005
R6925 CSoutput.n135 CSoutput.n116 4.5005
R6926 CSoutput.n135 CSoutput.n123 4.5005
R6927 CSoutput.n135 CSoutput.n124 4.5005
R6928 CSoutput.n133 CSoutput.n119 4.5005
R6929 CSoutput.n133 CSoutput.n121 4.5005
R6930 CSoutput.n133 CSoutput.n118 4.5005
R6931 CSoutput.n133 CSoutput.n122 4.5005
R6932 CSoutput.n133 CSoutput.n117 4.5005
R6933 CSoutput.n133 CSoutput.t154 4.5005
R6934 CSoutput.n133 CSoutput.n116 4.5005
R6935 CSoutput.n133 CSoutput.n123 4.5005
R6936 CSoutput.n133 CSoutput.n124 4.5005
R6937 CSoutput.n132 CSoutput.n119 4.5005
R6938 CSoutput.n132 CSoutput.n121 4.5005
R6939 CSoutput.n132 CSoutput.n118 4.5005
R6940 CSoutput.n132 CSoutput.n122 4.5005
R6941 CSoutput.n132 CSoutput.n117 4.5005
R6942 CSoutput.n132 CSoutput.t154 4.5005
R6943 CSoutput.n132 CSoutput.n116 4.5005
R6944 CSoutput.n132 CSoutput.n123 4.5005
R6945 CSoutput.n132 CSoutput.n124 4.5005
R6946 CSoutput.n261 CSoutput.n119 4.5005
R6947 CSoutput.n261 CSoutput.n121 4.5005
R6948 CSoutput.n261 CSoutput.n118 4.5005
R6949 CSoutput.n261 CSoutput.n122 4.5005
R6950 CSoutput.n261 CSoutput.n117 4.5005
R6951 CSoutput.n261 CSoutput.t154 4.5005
R6952 CSoutput.n261 CSoutput.n116 4.5005
R6953 CSoutput.n261 CSoutput.n123 4.5005
R6954 CSoutput.n261 CSoutput.n124 4.5005
R6955 CSoutput.n259 CSoutput.n119 4.5005
R6956 CSoutput.n259 CSoutput.n121 4.5005
R6957 CSoutput.n259 CSoutput.n118 4.5005
R6958 CSoutput.n259 CSoutput.n122 4.5005
R6959 CSoutput.n259 CSoutput.n117 4.5005
R6960 CSoutput.n259 CSoutput.t154 4.5005
R6961 CSoutput.n259 CSoutput.n116 4.5005
R6962 CSoutput.n259 CSoutput.n123 4.5005
R6963 CSoutput.n257 CSoutput.n119 4.5005
R6964 CSoutput.n257 CSoutput.n121 4.5005
R6965 CSoutput.n257 CSoutput.n118 4.5005
R6966 CSoutput.n257 CSoutput.n122 4.5005
R6967 CSoutput.n257 CSoutput.n117 4.5005
R6968 CSoutput.n257 CSoutput.t154 4.5005
R6969 CSoutput.n257 CSoutput.n116 4.5005
R6970 CSoutput.n257 CSoutput.n123 4.5005
R6971 CSoutput.n143 CSoutput.n119 4.5005
R6972 CSoutput.n143 CSoutput.n121 4.5005
R6973 CSoutput.n143 CSoutput.n118 4.5005
R6974 CSoutput.n143 CSoutput.n122 4.5005
R6975 CSoutput.n143 CSoutput.n117 4.5005
R6976 CSoutput.n143 CSoutput.t154 4.5005
R6977 CSoutput.n143 CSoutput.n116 4.5005
R6978 CSoutput.n143 CSoutput.n123 4.5005
R6979 CSoutput.n143 CSoutput.n124 4.5005
R6980 CSoutput.n142 CSoutput.n119 4.5005
R6981 CSoutput.n142 CSoutput.n121 4.5005
R6982 CSoutput.n142 CSoutput.n118 4.5005
R6983 CSoutput.n142 CSoutput.n122 4.5005
R6984 CSoutput.n142 CSoutput.n117 4.5005
R6985 CSoutput.n142 CSoutput.t154 4.5005
R6986 CSoutput.n142 CSoutput.n116 4.5005
R6987 CSoutput.n142 CSoutput.n123 4.5005
R6988 CSoutput.n142 CSoutput.n124 4.5005
R6989 CSoutput.n146 CSoutput.n119 4.5005
R6990 CSoutput.n146 CSoutput.n121 4.5005
R6991 CSoutput.n146 CSoutput.n118 4.5005
R6992 CSoutput.n146 CSoutput.n122 4.5005
R6993 CSoutput.n146 CSoutput.n117 4.5005
R6994 CSoutput.n146 CSoutput.t154 4.5005
R6995 CSoutput.n146 CSoutput.n116 4.5005
R6996 CSoutput.n146 CSoutput.n123 4.5005
R6997 CSoutput.n146 CSoutput.n124 4.5005
R6998 CSoutput.n145 CSoutput.n119 4.5005
R6999 CSoutput.n145 CSoutput.n121 4.5005
R7000 CSoutput.n145 CSoutput.n118 4.5005
R7001 CSoutput.n145 CSoutput.n122 4.5005
R7002 CSoutput.n145 CSoutput.n117 4.5005
R7003 CSoutput.n145 CSoutput.t154 4.5005
R7004 CSoutput.n145 CSoutput.n116 4.5005
R7005 CSoutput.n145 CSoutput.n123 4.5005
R7006 CSoutput.n145 CSoutput.n124 4.5005
R7007 CSoutput.n128 CSoutput.n119 4.5005
R7008 CSoutput.n128 CSoutput.n121 4.5005
R7009 CSoutput.n128 CSoutput.n118 4.5005
R7010 CSoutput.n128 CSoutput.n122 4.5005
R7011 CSoutput.n128 CSoutput.n117 4.5005
R7012 CSoutput.n128 CSoutput.t154 4.5005
R7013 CSoutput.n128 CSoutput.n116 4.5005
R7014 CSoutput.n128 CSoutput.n123 4.5005
R7015 CSoutput.n128 CSoutput.n124 4.5005
R7016 CSoutput.n264 CSoutput.n119 4.5005
R7017 CSoutput.n264 CSoutput.n121 4.5005
R7018 CSoutput.n264 CSoutput.n118 4.5005
R7019 CSoutput.n264 CSoutput.n122 4.5005
R7020 CSoutput.n264 CSoutput.n117 4.5005
R7021 CSoutput.n264 CSoutput.t154 4.5005
R7022 CSoutput.n264 CSoutput.n116 4.5005
R7023 CSoutput.n264 CSoutput.n123 4.5005
R7024 CSoutput.n264 CSoutput.n124 4.5005
R7025 CSoutput.n299 CSoutput.n287 4.10845
R7026 CSoutput.n113 CSoutput.n101 4.10845
R7027 CSoutput.n297 CSoutput.t57 4.06363
R7028 CSoutput.n297 CSoutput.t71 4.06363
R7029 CSoutput.n295 CSoutput.t80 4.06363
R7030 CSoutput.n295 CSoutput.t29 4.06363
R7031 CSoutput.n293 CSoutput.t33 4.06363
R7032 CSoutput.n293 CSoutput.t72 4.06363
R7033 CSoutput.n291 CSoutput.t81 4.06363
R7034 CSoutput.n291 CSoutput.t82 4.06363
R7035 CSoutput.n289 CSoutput.t46 4.06363
R7036 CSoutput.n289 CSoutput.t47 4.06363
R7037 CSoutput.n288 CSoutput.t48 4.06363
R7038 CSoutput.n288 CSoutput.t83 4.06363
R7039 CSoutput.n285 CSoutput.t49 4.06363
R7040 CSoutput.n285 CSoutput.t65 4.06363
R7041 CSoutput.n283 CSoutput.t75 4.06363
R7042 CSoutput.n283 CSoutput.t19 4.06363
R7043 CSoutput.n281 CSoutput.t20 4.06363
R7044 CSoutput.n281 CSoutput.t66 4.06363
R7045 CSoutput.n279 CSoutput.t76 4.06363
R7046 CSoutput.n279 CSoutput.t77 4.06363
R7047 CSoutput.n277 CSoutput.t35 4.06363
R7048 CSoutput.n277 CSoutput.t37 4.06363
R7049 CSoutput.n276 CSoutput.t38 4.06363
R7050 CSoutput.n276 CSoutput.t78 4.06363
R7051 CSoutput.n274 CSoutput.t70 4.06363
R7052 CSoutput.n274 CSoutput.t42 4.06363
R7053 CSoutput.n272 CSoutput.t63 4.06363
R7054 CSoutput.n272 CSoutput.t28 4.06363
R7055 CSoutput.n270 CSoutput.t74 4.06363
R7056 CSoutput.n270 CSoutput.t24 4.06363
R7057 CSoutput.n268 CSoutput.t51 4.06363
R7058 CSoutput.n268 CSoutput.t36 4.06363
R7059 CSoutput.n266 CSoutput.t39 4.06363
R7060 CSoutput.n266 CSoutput.t22 4.06363
R7061 CSoutput.n265 CSoutput.t69 4.06363
R7062 CSoutput.n265 CSoutput.t16 4.06363
R7063 CSoutput.n102 CSoutput.t45 4.06363
R7064 CSoutput.n102 CSoutput.t85 4.06363
R7065 CSoutput.n103 CSoutput.t67 4.06363
R7066 CSoutput.n103 CSoutput.t68 4.06363
R7067 CSoutput.n105 CSoutput.t59 4.06363
R7068 CSoutput.n105 CSoutput.t43 4.06363
R7069 CSoutput.n107 CSoutput.t27 4.06363
R7070 CSoutput.n107 CSoutput.t60 4.06363
R7071 CSoutput.n109 CSoutput.t58 4.06363
R7072 CSoutput.n109 CSoutput.t40 4.06363
R7073 CSoutput.n111 CSoutput.t26 4.06363
R7074 CSoutput.n111 CSoutput.t25 4.06363
R7075 CSoutput.n90 CSoutput.t34 4.06363
R7076 CSoutput.n90 CSoutput.t79 4.06363
R7077 CSoutput.n91 CSoutput.t64 4.06363
R7078 CSoutput.n91 CSoutput.t61 4.06363
R7079 CSoutput.n93 CSoutput.t54 4.06363
R7080 CSoutput.n93 CSoutput.t32 4.06363
R7081 CSoutput.n95 CSoutput.t17 4.06363
R7082 CSoutput.n95 CSoutput.t53 4.06363
R7083 CSoutput.n97 CSoutput.t52 4.06363
R7084 CSoutput.n97 CSoutput.t31 4.06363
R7085 CSoutput.n99 CSoutput.t14 4.06363
R7086 CSoutput.n99 CSoutput.t15 4.06363
R7087 CSoutput.n79 CSoutput.t18 4.06363
R7088 CSoutput.n79 CSoutput.t55 4.06363
R7089 CSoutput.n80 CSoutput.t21 4.06363
R7090 CSoutput.n80 CSoutput.t41 4.06363
R7091 CSoutput.n82 CSoutput.t84 4.06363
R7092 CSoutput.n82 CSoutput.t50 4.06363
R7093 CSoutput.n84 CSoutput.t23 4.06363
R7094 CSoutput.n84 CSoutput.t73 4.06363
R7095 CSoutput.n86 CSoutput.t30 4.06363
R7096 CSoutput.n86 CSoutput.t62 4.06363
R7097 CSoutput.n88 CSoutput.t44 4.06363
R7098 CSoutput.n88 CSoutput.t56 4.06363
R7099 CSoutput.n44 CSoutput.n43 3.79402
R7100 CSoutput.n49 CSoutput.n48 3.79402
R7101 CSoutput.n335 CSoutput.n323 3.72967
R7102 CSoutput.n371 CSoutput.n359 3.72967
R7103 CSoutput.n373 CSoutput.n372 3.57343
R7104 CSoutput.n372 CSoutput.n336 3.04641
R7105 CSoutput.n333 CSoutput.t118 2.82907
R7106 CSoutput.n333 CSoutput.t132 2.82907
R7107 CSoutput.n331 CSoutput.t102 2.82907
R7108 CSoutput.n331 CSoutput.t137 2.82907
R7109 CSoutput.n329 CSoutput.t129 2.82907
R7110 CSoutput.n329 CSoutput.t130 2.82907
R7111 CSoutput.n327 CSoutput.t8 2.82907
R7112 CSoutput.n327 CSoutput.t120 2.82907
R7113 CSoutput.n325 CSoutput.t99 2.82907
R7114 CSoutput.n325 CSoutput.t89 2.82907
R7115 CSoutput.n324 CSoutput.t92 2.82907
R7116 CSoutput.n324 CSoutput.t117 2.82907
R7117 CSoutput.n321 CSoutput.t95 2.82907
R7118 CSoutput.n321 CSoutput.t105 2.82907
R7119 CSoutput.n319 CSoutput.t107 2.82907
R7120 CSoutput.n319 CSoutput.t100 2.82907
R7121 CSoutput.n317 CSoutput.t115 2.82907
R7122 CSoutput.n317 CSoutput.t3 2.82907
R7123 CSoutput.n315 CSoutput.t124 2.82907
R7124 CSoutput.n315 CSoutput.t127 2.82907
R7125 CSoutput.n313 CSoutput.t97 2.82907
R7126 CSoutput.n313 CSoutput.t96 2.82907
R7127 CSoutput.n312 CSoutput.t94 2.82907
R7128 CSoutput.n312 CSoutput.t88 2.82907
R7129 CSoutput.n310 CSoutput.t135 2.82907
R7130 CSoutput.n310 CSoutput.t143 2.82907
R7131 CSoutput.n308 CSoutput.t10 2.82907
R7132 CSoutput.n308 CSoutput.t111 2.82907
R7133 CSoutput.n306 CSoutput.t140 2.82907
R7134 CSoutput.n306 CSoutput.t0 2.82907
R7135 CSoutput.n304 CSoutput.t6 2.82907
R7136 CSoutput.n304 CSoutput.t90 2.82907
R7137 CSoutput.n302 CSoutput.t110 2.82907
R7138 CSoutput.n302 CSoutput.t119 2.82907
R7139 CSoutput.n301 CSoutput.t104 2.82907
R7140 CSoutput.n301 CSoutput.t114 2.82907
R7141 CSoutput.n360 CSoutput.t86 2.82907
R7142 CSoutput.n360 CSoutput.t87 2.82907
R7143 CSoutput.n361 CSoutput.t131 2.82907
R7144 CSoutput.n361 CSoutput.t142 2.82907
R7145 CSoutput.n363 CSoutput.t109 2.82907
R7146 CSoutput.n363 CSoutput.t106 2.82907
R7147 CSoutput.n365 CSoutput.t134 2.82907
R7148 CSoutput.n365 CSoutput.t116 2.82907
R7149 CSoutput.n367 CSoutput.t101 2.82907
R7150 CSoutput.n367 CSoutput.t139 2.82907
R7151 CSoutput.n369 CSoutput.t91 2.82907
R7152 CSoutput.n369 CSoutput.t108 2.82907
R7153 CSoutput.n348 CSoutput.t7 2.82907
R7154 CSoutput.n348 CSoutput.t128 2.82907
R7155 CSoutput.n349 CSoutput.t138 2.82907
R7156 CSoutput.n349 CSoutput.t2 2.82907
R7157 CSoutput.n351 CSoutput.t1 2.82907
R7158 CSoutput.n351 CSoutput.t122 2.82907
R7159 CSoutput.n353 CSoutput.t5 2.82907
R7160 CSoutput.n353 CSoutput.t93 2.82907
R7161 CSoutput.n355 CSoutput.t103 2.82907
R7162 CSoutput.n355 CSoutput.t126 2.82907
R7163 CSoutput.n357 CSoutput.t4 2.82907
R7164 CSoutput.n357 CSoutput.t12 2.82907
R7165 CSoutput.n337 CSoutput.t112 2.82907
R7166 CSoutput.n337 CSoutput.t9 2.82907
R7167 CSoutput.n338 CSoutput.t11 2.82907
R7168 CSoutput.n338 CSoutput.t125 2.82907
R7169 CSoutput.n340 CSoutput.t13 2.82907
R7170 CSoutput.n340 CSoutput.t98 2.82907
R7171 CSoutput.n342 CSoutput.t141 2.82907
R7172 CSoutput.n342 CSoutput.t136 2.82907
R7173 CSoutput.n344 CSoutput.t121 2.82907
R7174 CSoutput.n344 CSoutput.t123 2.82907
R7175 CSoutput.n346 CSoutput.t113 2.82907
R7176 CSoutput.n346 CSoutput.t133 2.82907
R7177 CSoutput.n300 CSoutput.n114 2.57547
R7178 CSoutput.n75 CSoutput.n1 2.45513
R7179 CSoutput.n205 CSoutput.n203 2.251
R7180 CSoutput.n205 CSoutput.n202 2.251
R7181 CSoutput.n205 CSoutput.n201 2.251
R7182 CSoutput.n205 CSoutput.n200 2.251
R7183 CSoutput.n174 CSoutput.n173 2.251
R7184 CSoutput.n174 CSoutput.n172 2.251
R7185 CSoutput.n174 CSoutput.n171 2.251
R7186 CSoutput.n174 CSoutput.n170 2.251
R7187 CSoutput.n247 CSoutput.n246 2.251
R7188 CSoutput.n212 CSoutput.n210 2.251
R7189 CSoutput.n212 CSoutput.n209 2.251
R7190 CSoutput.n212 CSoutput.n208 2.251
R7191 CSoutput.n230 CSoutput.n212 2.251
R7192 CSoutput.n218 CSoutput.n217 2.251
R7193 CSoutput.n218 CSoutput.n216 2.251
R7194 CSoutput.n218 CSoutput.n215 2.251
R7195 CSoutput.n218 CSoutput.n214 2.251
R7196 CSoutput.n244 CSoutput.n184 2.251
R7197 CSoutput.n239 CSoutput.n237 2.251
R7198 CSoutput.n239 CSoutput.n236 2.251
R7199 CSoutput.n239 CSoutput.n235 2.251
R7200 CSoutput.n239 CSoutput.n234 2.251
R7201 CSoutput.n140 CSoutput.n139 2.251
R7202 CSoutput.n140 CSoutput.n138 2.251
R7203 CSoutput.n140 CSoutput.n137 2.251
R7204 CSoutput.n140 CSoutput.n136 2.251
R7205 CSoutput.n257 CSoutput.n256 2.251
R7206 CSoutput.n174 CSoutput.n154 2.2505
R7207 CSoutput.n169 CSoutput.n154 2.2505
R7208 CSoutput.n167 CSoutput.n154 2.2505
R7209 CSoutput.n166 CSoutput.n154 2.2505
R7210 CSoutput.n251 CSoutput.n154 2.2505
R7211 CSoutput.n249 CSoutput.n154 2.2505
R7212 CSoutput.n247 CSoutput.n154 2.2505
R7213 CSoutput.n177 CSoutput.n154 2.2505
R7214 CSoutput.n176 CSoutput.n154 2.2505
R7215 CSoutput.n180 CSoutput.n154 2.2505
R7216 CSoutput.n179 CSoutput.n154 2.2505
R7217 CSoutput.n162 CSoutput.n154 2.2505
R7218 CSoutput.n254 CSoutput.n154 2.2505
R7219 CSoutput.n254 CSoutput.n253 2.2505
R7220 CSoutput.n218 CSoutput.n189 2.2505
R7221 CSoutput.n199 CSoutput.n189 2.2505
R7222 CSoutput.n220 CSoutput.n189 2.2505
R7223 CSoutput.n198 CSoutput.n189 2.2505
R7224 CSoutput.n222 CSoutput.n189 2.2505
R7225 CSoutput.n189 CSoutput.n183 2.2505
R7226 CSoutput.n244 CSoutput.n189 2.2505
R7227 CSoutput.n242 CSoutput.n189 2.2505
R7228 CSoutput.n224 CSoutput.n189 2.2505
R7229 CSoutput.n196 CSoutput.n189 2.2505
R7230 CSoutput.n226 CSoutput.n189 2.2505
R7231 CSoutput.n195 CSoutput.n189 2.2505
R7232 CSoutput.n240 CSoutput.n189 2.2505
R7233 CSoutput.n240 CSoutput.n193 2.2505
R7234 CSoutput.n140 CSoutput.n120 2.2505
R7235 CSoutput.n135 CSoutput.n120 2.2505
R7236 CSoutput.n133 CSoutput.n120 2.2505
R7237 CSoutput.n132 CSoutput.n120 2.2505
R7238 CSoutput.n261 CSoutput.n120 2.2505
R7239 CSoutput.n259 CSoutput.n120 2.2505
R7240 CSoutput.n257 CSoutput.n120 2.2505
R7241 CSoutput.n143 CSoutput.n120 2.2505
R7242 CSoutput.n142 CSoutput.n120 2.2505
R7243 CSoutput.n146 CSoutput.n120 2.2505
R7244 CSoutput.n145 CSoutput.n120 2.2505
R7245 CSoutput.n128 CSoutput.n120 2.2505
R7246 CSoutput.n264 CSoutput.n120 2.2505
R7247 CSoutput.n264 CSoutput.n263 2.2505
R7248 CSoutput.n182 CSoutput.n175 2.25024
R7249 CSoutput.n182 CSoutput.n168 2.25024
R7250 CSoutput.n250 CSoutput.n182 2.25024
R7251 CSoutput.n182 CSoutput.n178 2.25024
R7252 CSoutput.n182 CSoutput.n181 2.25024
R7253 CSoutput.n182 CSoutput.n149 2.25024
R7254 CSoutput.n232 CSoutput.n229 2.25024
R7255 CSoutput.n232 CSoutput.n228 2.25024
R7256 CSoutput.n232 CSoutput.n227 2.25024
R7257 CSoutput.n232 CSoutput.n194 2.25024
R7258 CSoutput.n232 CSoutput.n231 2.25024
R7259 CSoutput.n233 CSoutput.n232 2.25024
R7260 CSoutput.n148 CSoutput.n141 2.25024
R7261 CSoutput.n148 CSoutput.n134 2.25024
R7262 CSoutput.n260 CSoutput.n148 2.25024
R7263 CSoutput.n148 CSoutput.n144 2.25024
R7264 CSoutput.n148 CSoutput.n147 2.25024
R7265 CSoutput.n148 CSoutput.n115 2.25024
R7266 CSoutput.n249 CSoutput.n159 1.50111
R7267 CSoutput.n197 CSoutput.n183 1.50111
R7268 CSoutput.n259 CSoutput.n125 1.50111
R7269 CSoutput.n205 CSoutput.n204 1.501
R7270 CSoutput.n212 CSoutput.n211 1.501
R7271 CSoutput.n239 CSoutput.n238 1.501
R7272 CSoutput.n253 CSoutput.n164 1.12536
R7273 CSoutput.n253 CSoutput.n165 1.12536
R7274 CSoutput.n253 CSoutput.n252 1.12536
R7275 CSoutput.n213 CSoutput.n193 1.12536
R7276 CSoutput.n219 CSoutput.n193 1.12536
R7277 CSoutput.n221 CSoutput.n193 1.12536
R7278 CSoutput.n263 CSoutput.n130 1.12536
R7279 CSoutput.n263 CSoutput.n131 1.12536
R7280 CSoutput.n263 CSoutput.n262 1.12536
R7281 CSoutput.n253 CSoutput.n160 1.12536
R7282 CSoutput.n253 CSoutput.n161 1.12536
R7283 CSoutput.n253 CSoutput.n163 1.12536
R7284 CSoutput.n243 CSoutput.n193 1.12536
R7285 CSoutput.n223 CSoutput.n193 1.12536
R7286 CSoutput.n225 CSoutput.n193 1.12536
R7287 CSoutput.n263 CSoutput.n126 1.12536
R7288 CSoutput.n263 CSoutput.n127 1.12536
R7289 CSoutput.n263 CSoutput.n129 1.12536
R7290 CSoutput.n31 CSoutput.n30 0.669944
R7291 CSoutput.n62 CSoutput.n61 0.669944
R7292 CSoutput.n328 CSoutput.n326 0.573776
R7293 CSoutput.n330 CSoutput.n328 0.573776
R7294 CSoutput.n332 CSoutput.n330 0.573776
R7295 CSoutput.n334 CSoutput.n332 0.573776
R7296 CSoutput.n316 CSoutput.n314 0.573776
R7297 CSoutput.n318 CSoutput.n316 0.573776
R7298 CSoutput.n320 CSoutput.n318 0.573776
R7299 CSoutput.n322 CSoutput.n320 0.573776
R7300 CSoutput.n305 CSoutput.n303 0.573776
R7301 CSoutput.n307 CSoutput.n305 0.573776
R7302 CSoutput.n309 CSoutput.n307 0.573776
R7303 CSoutput.n311 CSoutput.n309 0.573776
R7304 CSoutput.n370 CSoutput.n368 0.573776
R7305 CSoutput.n368 CSoutput.n366 0.573776
R7306 CSoutput.n366 CSoutput.n364 0.573776
R7307 CSoutput.n364 CSoutput.n362 0.573776
R7308 CSoutput.n358 CSoutput.n356 0.573776
R7309 CSoutput.n356 CSoutput.n354 0.573776
R7310 CSoutput.n354 CSoutput.n352 0.573776
R7311 CSoutput.n352 CSoutput.n350 0.573776
R7312 CSoutput.n347 CSoutput.n345 0.573776
R7313 CSoutput.n345 CSoutput.n343 0.573776
R7314 CSoutput.n343 CSoutput.n341 0.573776
R7315 CSoutput.n341 CSoutput.n339 0.573776
R7316 CSoutput.n373 CSoutput.n264 0.53442
R7317 CSoutput.n292 CSoutput.n290 0.358259
R7318 CSoutput.n294 CSoutput.n292 0.358259
R7319 CSoutput.n296 CSoutput.n294 0.358259
R7320 CSoutput.n298 CSoutput.n296 0.358259
R7321 CSoutput.n280 CSoutput.n278 0.358259
R7322 CSoutput.n282 CSoutput.n280 0.358259
R7323 CSoutput.n284 CSoutput.n282 0.358259
R7324 CSoutput.n286 CSoutput.n284 0.358259
R7325 CSoutput.n269 CSoutput.n267 0.358259
R7326 CSoutput.n271 CSoutput.n269 0.358259
R7327 CSoutput.n273 CSoutput.n271 0.358259
R7328 CSoutput.n275 CSoutput.n273 0.358259
R7329 CSoutput.n112 CSoutput.n110 0.358259
R7330 CSoutput.n110 CSoutput.n108 0.358259
R7331 CSoutput.n108 CSoutput.n106 0.358259
R7332 CSoutput.n106 CSoutput.n104 0.358259
R7333 CSoutput.n100 CSoutput.n98 0.358259
R7334 CSoutput.n98 CSoutput.n96 0.358259
R7335 CSoutput.n96 CSoutput.n94 0.358259
R7336 CSoutput.n94 CSoutput.n92 0.358259
R7337 CSoutput.n89 CSoutput.n87 0.358259
R7338 CSoutput.n87 CSoutput.n85 0.358259
R7339 CSoutput.n85 CSoutput.n83 0.358259
R7340 CSoutput.n83 CSoutput.n81 0.358259
R7341 CSoutput.n21 CSoutput.n20 0.169105
R7342 CSoutput.n21 CSoutput.n16 0.169105
R7343 CSoutput.n26 CSoutput.n16 0.169105
R7344 CSoutput.n27 CSoutput.n26 0.169105
R7345 CSoutput.n27 CSoutput.n14 0.169105
R7346 CSoutput.n32 CSoutput.n14 0.169105
R7347 CSoutput.n33 CSoutput.n32 0.169105
R7348 CSoutput.n34 CSoutput.n33 0.169105
R7349 CSoutput.n34 CSoutput.n12 0.169105
R7350 CSoutput.n39 CSoutput.n12 0.169105
R7351 CSoutput.n40 CSoutput.n39 0.169105
R7352 CSoutput.n40 CSoutput.n10 0.169105
R7353 CSoutput.n45 CSoutput.n10 0.169105
R7354 CSoutput.n46 CSoutput.n45 0.169105
R7355 CSoutput.n47 CSoutput.n46 0.169105
R7356 CSoutput.n47 CSoutput.n8 0.169105
R7357 CSoutput.n52 CSoutput.n8 0.169105
R7358 CSoutput.n53 CSoutput.n52 0.169105
R7359 CSoutput.n53 CSoutput.n6 0.169105
R7360 CSoutput.n58 CSoutput.n6 0.169105
R7361 CSoutput.n59 CSoutput.n58 0.169105
R7362 CSoutput.n60 CSoutput.n59 0.169105
R7363 CSoutput.n60 CSoutput.n4 0.169105
R7364 CSoutput.n66 CSoutput.n4 0.169105
R7365 CSoutput.n67 CSoutput.n66 0.169105
R7366 CSoutput.n68 CSoutput.n67 0.169105
R7367 CSoutput.n68 CSoutput.n2 0.169105
R7368 CSoutput.n73 CSoutput.n2 0.169105
R7369 CSoutput.n74 CSoutput.n73 0.169105
R7370 CSoutput.n74 CSoutput.n0 0.169105
R7371 CSoutput.n78 CSoutput.n0 0.169105
R7372 CSoutput.n207 CSoutput.n206 0.0910737
R7373 CSoutput.n258 CSoutput.n255 0.0723685
R7374 CSoutput.n212 CSoutput.n207 0.0522944
R7375 CSoutput.n255 CSoutput.n254 0.0499135
R7376 CSoutput.n206 CSoutput.n205 0.0499135
R7377 CSoutput.n240 CSoutput.n239 0.0464294
R7378 CSoutput.n248 CSoutput.n245 0.0391444
R7379 CSoutput.n207 CSoutput.t163 0.023435
R7380 CSoutput.n255 CSoutput.t144 0.02262
R7381 CSoutput.n206 CSoutput.t146 0.02262
R7382 CSoutput CSoutput.n373 0.0052
R7383 CSoutput.n177 CSoutput.n160 0.00365111
R7384 CSoutput.n180 CSoutput.n161 0.00365111
R7385 CSoutput.n163 CSoutput.n162 0.00365111
R7386 CSoutput.n205 CSoutput.n164 0.00365111
R7387 CSoutput.n169 CSoutput.n165 0.00365111
R7388 CSoutput.n252 CSoutput.n166 0.00365111
R7389 CSoutput.n243 CSoutput.n242 0.00365111
R7390 CSoutput.n223 CSoutput.n196 0.00365111
R7391 CSoutput.n225 CSoutput.n195 0.00365111
R7392 CSoutput.n213 CSoutput.n212 0.00365111
R7393 CSoutput.n219 CSoutput.n199 0.00365111
R7394 CSoutput.n221 CSoutput.n198 0.00365111
R7395 CSoutput.n143 CSoutput.n126 0.00365111
R7396 CSoutput.n146 CSoutput.n127 0.00365111
R7397 CSoutput.n129 CSoutput.n128 0.00365111
R7398 CSoutput.n239 CSoutput.n130 0.00365111
R7399 CSoutput.n135 CSoutput.n131 0.00365111
R7400 CSoutput.n262 CSoutput.n132 0.00365111
R7401 CSoutput.n174 CSoutput.n164 0.00340054
R7402 CSoutput.n167 CSoutput.n165 0.00340054
R7403 CSoutput.n252 CSoutput.n251 0.00340054
R7404 CSoutput.n247 CSoutput.n160 0.00340054
R7405 CSoutput.n176 CSoutput.n161 0.00340054
R7406 CSoutput.n179 CSoutput.n163 0.00340054
R7407 CSoutput.n218 CSoutput.n213 0.00340054
R7408 CSoutput.n220 CSoutput.n219 0.00340054
R7409 CSoutput.n222 CSoutput.n221 0.00340054
R7410 CSoutput.n244 CSoutput.n243 0.00340054
R7411 CSoutput.n224 CSoutput.n223 0.00340054
R7412 CSoutput.n226 CSoutput.n225 0.00340054
R7413 CSoutput.n140 CSoutput.n130 0.00340054
R7414 CSoutput.n133 CSoutput.n131 0.00340054
R7415 CSoutput.n262 CSoutput.n261 0.00340054
R7416 CSoutput.n257 CSoutput.n126 0.00340054
R7417 CSoutput.n142 CSoutput.n127 0.00340054
R7418 CSoutput.n145 CSoutput.n129 0.00340054
R7419 CSoutput.n175 CSoutput.n169 0.00252698
R7420 CSoutput.n168 CSoutput.n166 0.00252698
R7421 CSoutput.n250 CSoutput.n249 0.00252698
R7422 CSoutput.n178 CSoutput.n176 0.00252698
R7423 CSoutput.n181 CSoutput.n179 0.00252698
R7424 CSoutput.n254 CSoutput.n149 0.00252698
R7425 CSoutput.n175 CSoutput.n174 0.00252698
R7426 CSoutput.n168 CSoutput.n167 0.00252698
R7427 CSoutput.n251 CSoutput.n250 0.00252698
R7428 CSoutput.n178 CSoutput.n177 0.00252698
R7429 CSoutput.n181 CSoutput.n180 0.00252698
R7430 CSoutput.n162 CSoutput.n149 0.00252698
R7431 CSoutput.n229 CSoutput.n199 0.00252698
R7432 CSoutput.n228 CSoutput.n198 0.00252698
R7433 CSoutput.n227 CSoutput.n183 0.00252698
R7434 CSoutput.n224 CSoutput.n194 0.00252698
R7435 CSoutput.n231 CSoutput.n226 0.00252698
R7436 CSoutput.n240 CSoutput.n233 0.00252698
R7437 CSoutput.n229 CSoutput.n218 0.00252698
R7438 CSoutput.n228 CSoutput.n220 0.00252698
R7439 CSoutput.n227 CSoutput.n222 0.00252698
R7440 CSoutput.n242 CSoutput.n194 0.00252698
R7441 CSoutput.n231 CSoutput.n196 0.00252698
R7442 CSoutput.n233 CSoutput.n195 0.00252698
R7443 CSoutput.n141 CSoutput.n135 0.00252698
R7444 CSoutput.n134 CSoutput.n132 0.00252698
R7445 CSoutput.n260 CSoutput.n259 0.00252698
R7446 CSoutput.n144 CSoutput.n142 0.00252698
R7447 CSoutput.n147 CSoutput.n145 0.00252698
R7448 CSoutput.n264 CSoutput.n115 0.00252698
R7449 CSoutput.n141 CSoutput.n140 0.00252698
R7450 CSoutput.n134 CSoutput.n133 0.00252698
R7451 CSoutput.n261 CSoutput.n260 0.00252698
R7452 CSoutput.n144 CSoutput.n143 0.00252698
R7453 CSoutput.n147 CSoutput.n146 0.00252698
R7454 CSoutput.n128 CSoutput.n115 0.00252698
R7455 CSoutput.n249 CSoutput.n248 0.0020275
R7456 CSoutput.n248 CSoutput.n247 0.0020275
R7457 CSoutput.n245 CSoutput.n183 0.0020275
R7458 CSoutput.n245 CSoutput.n244 0.0020275
R7459 CSoutput.n259 CSoutput.n258 0.0020275
R7460 CSoutput.n258 CSoutput.n257 0.0020275
R7461 CSoutput.n159 CSoutput.n158 0.00166668
R7462 CSoutput.n241 CSoutput.n197 0.00166668
R7463 CSoutput.n125 CSoutput.n124 0.00166668
R7464 CSoutput.n263 CSoutput.n125 0.00133328
R7465 CSoutput.n197 CSoutput.n193 0.00133328
R7466 CSoutput.n253 CSoutput.n159 0.00133328
R7467 CSoutput.n256 CSoutput.n148 0.001
R7468 CSoutput.n234 CSoutput.n148 0.001
R7469 CSoutput.n136 CSoutput.n116 0.001
R7470 CSoutput.n235 CSoutput.n116 0.001
R7471 CSoutput.n137 CSoutput.n117 0.001
R7472 CSoutput.n236 CSoutput.n117 0.001
R7473 CSoutput.n138 CSoutput.n118 0.001
R7474 CSoutput.n237 CSoutput.n118 0.001
R7475 CSoutput.n139 CSoutput.n119 0.001
R7476 CSoutput.n238 CSoutput.n119 0.001
R7477 CSoutput.n232 CSoutput.n184 0.001
R7478 CSoutput.n232 CSoutput.n230 0.001
R7479 CSoutput.n214 CSoutput.n185 0.001
R7480 CSoutput.n208 CSoutput.n185 0.001
R7481 CSoutput.n215 CSoutput.n186 0.001
R7482 CSoutput.n209 CSoutput.n186 0.001
R7483 CSoutput.n216 CSoutput.n187 0.001
R7484 CSoutput.n210 CSoutput.n187 0.001
R7485 CSoutput.n217 CSoutput.n188 0.001
R7486 CSoutput.n211 CSoutput.n188 0.001
R7487 CSoutput.n246 CSoutput.n182 0.001
R7488 CSoutput.n200 CSoutput.n182 0.001
R7489 CSoutput.n170 CSoutput.n150 0.001
R7490 CSoutput.n201 CSoutput.n150 0.001
R7491 CSoutput.n171 CSoutput.n151 0.001
R7492 CSoutput.n202 CSoutput.n151 0.001
R7493 CSoutput.n172 CSoutput.n152 0.001
R7494 CSoutput.n203 CSoutput.n152 0.001
R7495 CSoutput.n173 CSoutput.n153 0.001
R7496 CSoutput.n204 CSoutput.n153 0.001
R7497 CSoutput.n204 CSoutput.n154 0.001
R7498 CSoutput.n203 CSoutput.n155 0.001
R7499 CSoutput.n202 CSoutput.n156 0.001
R7500 CSoutput.n201 CSoutput.t162 0.001
R7501 CSoutput.n200 CSoutput.n157 0.001
R7502 CSoutput.n173 CSoutput.n155 0.001
R7503 CSoutput.n172 CSoutput.n156 0.001
R7504 CSoutput.n171 CSoutput.t162 0.001
R7505 CSoutput.n170 CSoutput.n157 0.001
R7506 CSoutput.n246 CSoutput.n158 0.001
R7507 CSoutput.n211 CSoutput.n189 0.001
R7508 CSoutput.n210 CSoutput.n190 0.001
R7509 CSoutput.n209 CSoutput.n191 0.001
R7510 CSoutput.n208 CSoutput.t155 0.001
R7511 CSoutput.n230 CSoutput.n192 0.001
R7512 CSoutput.n217 CSoutput.n190 0.001
R7513 CSoutput.n216 CSoutput.n191 0.001
R7514 CSoutput.n215 CSoutput.t155 0.001
R7515 CSoutput.n214 CSoutput.n192 0.001
R7516 CSoutput.n241 CSoutput.n184 0.001
R7517 CSoutput.n238 CSoutput.n120 0.001
R7518 CSoutput.n237 CSoutput.n121 0.001
R7519 CSoutput.n236 CSoutput.n122 0.001
R7520 CSoutput.n235 CSoutput.t154 0.001
R7521 CSoutput.n234 CSoutput.n123 0.001
R7522 CSoutput.n139 CSoutput.n121 0.001
R7523 CSoutput.n138 CSoutput.n122 0.001
R7524 CSoutput.n137 CSoutput.t154 0.001
R7525 CSoutput.n136 CSoutput.n123 0.001
R7526 CSoutput.n256 CSoutput.n124 0.001
R7527 commonsourceibias.n25 commonsourceibias.t38 230.006
R7528 commonsourceibias.n91 commonsourceibias.t95 230.006
R7529 commonsourceibias.n218 commonsourceibias.t117 230.006
R7530 commonsourceibias.n154 commonsourceibias.t97 230.006
R7531 commonsourceibias.n322 commonsourceibias.t44 230.006
R7532 commonsourceibias.n281 commonsourceibias.t70 230.006
R7533 commonsourceibias.n483 commonsourceibias.t55 230.006
R7534 commonsourceibias.n419 commonsourceibias.t80 230.006
R7535 commonsourceibias.n70 commonsourceibias.t28 207.983
R7536 commonsourceibias.n136 commonsourceibias.t56 207.983
R7537 commonsourceibias.n263 commonsourceibias.t111 207.983
R7538 commonsourceibias.n199 commonsourceibias.t89 207.983
R7539 commonsourceibias.n368 commonsourceibias.t8 207.983
R7540 commonsourceibias.n402 commonsourceibias.t114 207.983
R7541 commonsourceibias.n529 commonsourceibias.t51 207.983
R7542 commonsourceibias.n465 commonsourceibias.t74 207.983
R7543 commonsourceibias.n10 commonsourceibias.t4 168.701
R7544 commonsourceibias.n63 commonsourceibias.t42 168.701
R7545 commonsourceibias.n57 commonsourceibias.t40 168.701
R7546 commonsourceibias.n16 commonsourceibias.t16 168.701
R7547 commonsourceibias.n49 commonsourceibias.t22 168.701
R7548 commonsourceibias.n43 commonsourceibias.t34 168.701
R7549 commonsourceibias.n19 commonsourceibias.t14 168.701
R7550 commonsourceibias.n21 commonsourceibias.t6 168.701
R7551 commonsourceibias.n23 commonsourceibias.t18 168.701
R7552 commonsourceibias.n26 commonsourceibias.t46 168.701
R7553 commonsourceibias.n1 commonsourceibias.t109 168.701
R7554 commonsourceibias.n129 commonsourceibias.t69 168.701
R7555 commonsourceibias.n123 commonsourceibias.t119 168.701
R7556 commonsourceibias.n7 commonsourceibias.t85 168.701
R7557 commonsourceibias.n115 commonsourceibias.t54 168.701
R7558 commonsourceibias.n109 commonsourceibias.t100 168.701
R7559 commonsourceibias.n85 commonsourceibias.t87 168.701
R7560 commonsourceibias.n87 commonsourceibias.t115 168.701
R7561 commonsourceibias.n89 commonsourceibias.t79 168.701
R7562 commonsourceibias.n92 commonsourceibias.t66 168.701
R7563 commonsourceibias.n219 commonsourceibias.t75 168.701
R7564 commonsourceibias.n216 commonsourceibias.t59 168.701
R7565 commonsourceibias.n214 commonsourceibias.t49 168.701
R7566 commonsourceibias.n212 commonsourceibias.t84 168.701
R7567 commonsourceibias.n236 commonsourceibias.t93 168.701
R7568 commonsourceibias.n242 commonsourceibias.t52 168.701
R7569 commonsourceibias.n209 commonsourceibias.t118 168.701
R7570 commonsourceibias.n250 commonsourceibias.t104 168.701
R7571 commonsourceibias.n256 commonsourceibias.t60 168.701
R7572 commonsourceibias.n203 commonsourceibias.t50 168.701
R7573 commonsourceibias.n139 commonsourceibias.t106 168.701
R7574 commonsourceibias.n192 commonsourceibias.t101 168.701
R7575 commonsourceibias.n186 commonsourceibias.t88 168.701
R7576 commonsourceibias.n145 commonsourceibias.t105 168.701
R7577 commonsourceibias.n178 commonsourceibias.t99 168.701
R7578 commonsourceibias.n172 commonsourceibias.t86 168.701
R7579 commonsourceibias.n148 commonsourceibias.t108 168.701
R7580 commonsourceibias.n150 commonsourceibias.t98 168.701
R7581 commonsourceibias.n152 commonsourceibias.t112 168.701
R7582 commonsourceibias.n155 commonsourceibias.t107 168.701
R7583 commonsourceibias.n323 commonsourceibias.t26 168.701
R7584 commonsourceibias.n320 commonsourceibias.t2 168.701
R7585 commonsourceibias.n318 commonsourceibias.t12 168.701
R7586 commonsourceibias.n316 commonsourceibias.t30 168.701
R7587 commonsourceibias.n340 commonsourceibias.t0 168.701
R7588 commonsourceibias.n346 commonsourceibias.t10 168.701
R7589 commonsourceibias.n348 commonsourceibias.t32 168.701
R7590 commonsourceibias.n355 commonsourceibias.t36 168.701
R7591 commonsourceibias.n361 commonsourceibias.t24 168.701
R7592 commonsourceibias.n308 commonsourceibias.t20 168.701
R7593 commonsourceibias.n267 commonsourceibias.t78 168.701
R7594 commonsourceibias.n395 commonsourceibias.t53 168.701
R7595 commonsourceibias.n389 commonsourceibias.t94 168.701
R7596 commonsourceibias.n382 commonsourceibias.t64 168.701
R7597 commonsourceibias.n380 commonsourceibias.t113 168.701
R7598 commonsourceibias.n282 commonsourceibias.t58 168.701
R7599 commonsourceibias.n279 commonsourceibias.t63 168.701
R7600 commonsourceibias.n277 commonsourceibias.t92 168.701
R7601 commonsourceibias.n275 commonsourceibias.t65 168.701
R7602 commonsourceibias.n299 commonsourceibias.t76 168.701
R7603 commonsourceibias.n484 commonsourceibias.t68 168.701
R7604 commonsourceibias.n481 commonsourceibias.t72 168.701
R7605 commonsourceibias.n479 commonsourceibias.t61 168.701
R7606 commonsourceibias.n477 commonsourceibias.t110 168.701
R7607 commonsourceibias.n501 commonsourceibias.t77 168.701
R7608 commonsourceibias.n507 commonsourceibias.t67 168.701
R7609 commonsourceibias.n509 commonsourceibias.t57 168.701
R7610 commonsourceibias.n516 commonsourceibias.t48 168.701
R7611 commonsourceibias.n522 commonsourceibias.t71 168.701
R7612 commonsourceibias.n469 commonsourceibias.t62 168.701
R7613 commonsourceibias.n420 commonsourceibias.t116 168.701
R7614 commonsourceibias.n417 commonsourceibias.t102 168.701
R7615 commonsourceibias.n415 commonsourceibias.t81 168.701
R7616 commonsourceibias.n413 commonsourceibias.t96 168.701
R7617 commonsourceibias.n437 commonsourceibias.t103 168.701
R7618 commonsourceibias.n443 commonsourceibias.t82 168.701
R7619 commonsourceibias.n445 commonsourceibias.t90 168.701
R7620 commonsourceibias.n452 commonsourceibias.t73 168.701
R7621 commonsourceibias.n458 commonsourceibias.t83 168.701
R7622 commonsourceibias.n405 commonsourceibias.t91 168.701
R7623 commonsourceibias.n27 commonsourceibias.n24 161.3
R7624 commonsourceibias.n29 commonsourceibias.n28 161.3
R7625 commonsourceibias.n31 commonsourceibias.n30 161.3
R7626 commonsourceibias.n32 commonsourceibias.n22 161.3
R7627 commonsourceibias.n34 commonsourceibias.n33 161.3
R7628 commonsourceibias.n36 commonsourceibias.n35 161.3
R7629 commonsourceibias.n37 commonsourceibias.n20 161.3
R7630 commonsourceibias.n39 commonsourceibias.n38 161.3
R7631 commonsourceibias.n41 commonsourceibias.n40 161.3
R7632 commonsourceibias.n42 commonsourceibias.n18 161.3
R7633 commonsourceibias.n45 commonsourceibias.n44 161.3
R7634 commonsourceibias.n46 commonsourceibias.n17 161.3
R7635 commonsourceibias.n48 commonsourceibias.n47 161.3
R7636 commonsourceibias.n50 commonsourceibias.n15 161.3
R7637 commonsourceibias.n52 commonsourceibias.n51 161.3
R7638 commonsourceibias.n53 commonsourceibias.n14 161.3
R7639 commonsourceibias.n55 commonsourceibias.n54 161.3
R7640 commonsourceibias.n56 commonsourceibias.n13 161.3
R7641 commonsourceibias.n59 commonsourceibias.n58 161.3
R7642 commonsourceibias.n60 commonsourceibias.n12 161.3
R7643 commonsourceibias.n62 commonsourceibias.n61 161.3
R7644 commonsourceibias.n64 commonsourceibias.n11 161.3
R7645 commonsourceibias.n66 commonsourceibias.n65 161.3
R7646 commonsourceibias.n68 commonsourceibias.n67 161.3
R7647 commonsourceibias.n69 commonsourceibias.n9 161.3
R7648 commonsourceibias.n93 commonsourceibias.n90 161.3
R7649 commonsourceibias.n95 commonsourceibias.n94 161.3
R7650 commonsourceibias.n97 commonsourceibias.n96 161.3
R7651 commonsourceibias.n98 commonsourceibias.n88 161.3
R7652 commonsourceibias.n100 commonsourceibias.n99 161.3
R7653 commonsourceibias.n102 commonsourceibias.n101 161.3
R7654 commonsourceibias.n103 commonsourceibias.n86 161.3
R7655 commonsourceibias.n105 commonsourceibias.n104 161.3
R7656 commonsourceibias.n107 commonsourceibias.n106 161.3
R7657 commonsourceibias.n108 commonsourceibias.n84 161.3
R7658 commonsourceibias.n111 commonsourceibias.n110 161.3
R7659 commonsourceibias.n112 commonsourceibias.n8 161.3
R7660 commonsourceibias.n114 commonsourceibias.n113 161.3
R7661 commonsourceibias.n116 commonsourceibias.n6 161.3
R7662 commonsourceibias.n118 commonsourceibias.n117 161.3
R7663 commonsourceibias.n119 commonsourceibias.n5 161.3
R7664 commonsourceibias.n121 commonsourceibias.n120 161.3
R7665 commonsourceibias.n122 commonsourceibias.n4 161.3
R7666 commonsourceibias.n125 commonsourceibias.n124 161.3
R7667 commonsourceibias.n126 commonsourceibias.n3 161.3
R7668 commonsourceibias.n128 commonsourceibias.n127 161.3
R7669 commonsourceibias.n130 commonsourceibias.n2 161.3
R7670 commonsourceibias.n132 commonsourceibias.n131 161.3
R7671 commonsourceibias.n134 commonsourceibias.n133 161.3
R7672 commonsourceibias.n135 commonsourceibias.n0 161.3
R7673 commonsourceibias.n262 commonsourceibias.n202 161.3
R7674 commonsourceibias.n261 commonsourceibias.n260 161.3
R7675 commonsourceibias.n259 commonsourceibias.n258 161.3
R7676 commonsourceibias.n257 commonsourceibias.n204 161.3
R7677 commonsourceibias.n255 commonsourceibias.n254 161.3
R7678 commonsourceibias.n253 commonsourceibias.n205 161.3
R7679 commonsourceibias.n252 commonsourceibias.n251 161.3
R7680 commonsourceibias.n249 commonsourceibias.n206 161.3
R7681 commonsourceibias.n248 commonsourceibias.n247 161.3
R7682 commonsourceibias.n246 commonsourceibias.n207 161.3
R7683 commonsourceibias.n245 commonsourceibias.n244 161.3
R7684 commonsourceibias.n243 commonsourceibias.n208 161.3
R7685 commonsourceibias.n241 commonsourceibias.n240 161.3
R7686 commonsourceibias.n239 commonsourceibias.n210 161.3
R7687 commonsourceibias.n238 commonsourceibias.n237 161.3
R7688 commonsourceibias.n235 commonsourceibias.n211 161.3
R7689 commonsourceibias.n234 commonsourceibias.n233 161.3
R7690 commonsourceibias.n232 commonsourceibias.n231 161.3
R7691 commonsourceibias.n230 commonsourceibias.n213 161.3
R7692 commonsourceibias.n229 commonsourceibias.n228 161.3
R7693 commonsourceibias.n227 commonsourceibias.n226 161.3
R7694 commonsourceibias.n225 commonsourceibias.n215 161.3
R7695 commonsourceibias.n224 commonsourceibias.n223 161.3
R7696 commonsourceibias.n222 commonsourceibias.n221 161.3
R7697 commonsourceibias.n220 commonsourceibias.n217 161.3
R7698 commonsourceibias.n156 commonsourceibias.n153 161.3
R7699 commonsourceibias.n158 commonsourceibias.n157 161.3
R7700 commonsourceibias.n160 commonsourceibias.n159 161.3
R7701 commonsourceibias.n161 commonsourceibias.n151 161.3
R7702 commonsourceibias.n163 commonsourceibias.n162 161.3
R7703 commonsourceibias.n165 commonsourceibias.n164 161.3
R7704 commonsourceibias.n166 commonsourceibias.n149 161.3
R7705 commonsourceibias.n168 commonsourceibias.n167 161.3
R7706 commonsourceibias.n170 commonsourceibias.n169 161.3
R7707 commonsourceibias.n171 commonsourceibias.n147 161.3
R7708 commonsourceibias.n174 commonsourceibias.n173 161.3
R7709 commonsourceibias.n175 commonsourceibias.n146 161.3
R7710 commonsourceibias.n177 commonsourceibias.n176 161.3
R7711 commonsourceibias.n179 commonsourceibias.n144 161.3
R7712 commonsourceibias.n181 commonsourceibias.n180 161.3
R7713 commonsourceibias.n182 commonsourceibias.n143 161.3
R7714 commonsourceibias.n184 commonsourceibias.n183 161.3
R7715 commonsourceibias.n185 commonsourceibias.n142 161.3
R7716 commonsourceibias.n188 commonsourceibias.n187 161.3
R7717 commonsourceibias.n189 commonsourceibias.n141 161.3
R7718 commonsourceibias.n191 commonsourceibias.n190 161.3
R7719 commonsourceibias.n193 commonsourceibias.n140 161.3
R7720 commonsourceibias.n195 commonsourceibias.n194 161.3
R7721 commonsourceibias.n197 commonsourceibias.n196 161.3
R7722 commonsourceibias.n198 commonsourceibias.n138 161.3
R7723 commonsourceibias.n367 commonsourceibias.n307 161.3
R7724 commonsourceibias.n366 commonsourceibias.n365 161.3
R7725 commonsourceibias.n364 commonsourceibias.n363 161.3
R7726 commonsourceibias.n362 commonsourceibias.n309 161.3
R7727 commonsourceibias.n360 commonsourceibias.n359 161.3
R7728 commonsourceibias.n358 commonsourceibias.n310 161.3
R7729 commonsourceibias.n357 commonsourceibias.n356 161.3
R7730 commonsourceibias.n354 commonsourceibias.n311 161.3
R7731 commonsourceibias.n353 commonsourceibias.n352 161.3
R7732 commonsourceibias.n351 commonsourceibias.n312 161.3
R7733 commonsourceibias.n350 commonsourceibias.n349 161.3
R7734 commonsourceibias.n347 commonsourceibias.n313 161.3
R7735 commonsourceibias.n345 commonsourceibias.n344 161.3
R7736 commonsourceibias.n343 commonsourceibias.n314 161.3
R7737 commonsourceibias.n342 commonsourceibias.n341 161.3
R7738 commonsourceibias.n339 commonsourceibias.n315 161.3
R7739 commonsourceibias.n338 commonsourceibias.n337 161.3
R7740 commonsourceibias.n336 commonsourceibias.n335 161.3
R7741 commonsourceibias.n334 commonsourceibias.n317 161.3
R7742 commonsourceibias.n333 commonsourceibias.n332 161.3
R7743 commonsourceibias.n331 commonsourceibias.n330 161.3
R7744 commonsourceibias.n329 commonsourceibias.n319 161.3
R7745 commonsourceibias.n328 commonsourceibias.n327 161.3
R7746 commonsourceibias.n326 commonsourceibias.n325 161.3
R7747 commonsourceibias.n324 commonsourceibias.n321 161.3
R7748 commonsourceibias.n301 commonsourceibias.n300 161.3
R7749 commonsourceibias.n298 commonsourceibias.n274 161.3
R7750 commonsourceibias.n297 commonsourceibias.n296 161.3
R7751 commonsourceibias.n295 commonsourceibias.n294 161.3
R7752 commonsourceibias.n293 commonsourceibias.n276 161.3
R7753 commonsourceibias.n292 commonsourceibias.n291 161.3
R7754 commonsourceibias.n290 commonsourceibias.n289 161.3
R7755 commonsourceibias.n288 commonsourceibias.n278 161.3
R7756 commonsourceibias.n287 commonsourceibias.n286 161.3
R7757 commonsourceibias.n285 commonsourceibias.n284 161.3
R7758 commonsourceibias.n283 commonsourceibias.n280 161.3
R7759 commonsourceibias.n377 commonsourceibias.n273 161.3
R7760 commonsourceibias.n401 commonsourceibias.n266 161.3
R7761 commonsourceibias.n400 commonsourceibias.n399 161.3
R7762 commonsourceibias.n398 commonsourceibias.n397 161.3
R7763 commonsourceibias.n396 commonsourceibias.n268 161.3
R7764 commonsourceibias.n394 commonsourceibias.n393 161.3
R7765 commonsourceibias.n392 commonsourceibias.n269 161.3
R7766 commonsourceibias.n391 commonsourceibias.n390 161.3
R7767 commonsourceibias.n388 commonsourceibias.n270 161.3
R7768 commonsourceibias.n387 commonsourceibias.n386 161.3
R7769 commonsourceibias.n385 commonsourceibias.n271 161.3
R7770 commonsourceibias.n384 commonsourceibias.n383 161.3
R7771 commonsourceibias.n381 commonsourceibias.n272 161.3
R7772 commonsourceibias.n379 commonsourceibias.n378 161.3
R7773 commonsourceibias.n528 commonsourceibias.n468 161.3
R7774 commonsourceibias.n527 commonsourceibias.n526 161.3
R7775 commonsourceibias.n525 commonsourceibias.n524 161.3
R7776 commonsourceibias.n523 commonsourceibias.n470 161.3
R7777 commonsourceibias.n521 commonsourceibias.n520 161.3
R7778 commonsourceibias.n519 commonsourceibias.n471 161.3
R7779 commonsourceibias.n518 commonsourceibias.n517 161.3
R7780 commonsourceibias.n515 commonsourceibias.n472 161.3
R7781 commonsourceibias.n514 commonsourceibias.n513 161.3
R7782 commonsourceibias.n512 commonsourceibias.n473 161.3
R7783 commonsourceibias.n511 commonsourceibias.n510 161.3
R7784 commonsourceibias.n508 commonsourceibias.n474 161.3
R7785 commonsourceibias.n506 commonsourceibias.n505 161.3
R7786 commonsourceibias.n504 commonsourceibias.n475 161.3
R7787 commonsourceibias.n503 commonsourceibias.n502 161.3
R7788 commonsourceibias.n500 commonsourceibias.n476 161.3
R7789 commonsourceibias.n499 commonsourceibias.n498 161.3
R7790 commonsourceibias.n497 commonsourceibias.n496 161.3
R7791 commonsourceibias.n495 commonsourceibias.n478 161.3
R7792 commonsourceibias.n494 commonsourceibias.n493 161.3
R7793 commonsourceibias.n492 commonsourceibias.n491 161.3
R7794 commonsourceibias.n490 commonsourceibias.n480 161.3
R7795 commonsourceibias.n489 commonsourceibias.n488 161.3
R7796 commonsourceibias.n487 commonsourceibias.n486 161.3
R7797 commonsourceibias.n485 commonsourceibias.n482 161.3
R7798 commonsourceibias.n464 commonsourceibias.n404 161.3
R7799 commonsourceibias.n463 commonsourceibias.n462 161.3
R7800 commonsourceibias.n461 commonsourceibias.n460 161.3
R7801 commonsourceibias.n459 commonsourceibias.n406 161.3
R7802 commonsourceibias.n457 commonsourceibias.n456 161.3
R7803 commonsourceibias.n455 commonsourceibias.n407 161.3
R7804 commonsourceibias.n454 commonsourceibias.n453 161.3
R7805 commonsourceibias.n451 commonsourceibias.n408 161.3
R7806 commonsourceibias.n450 commonsourceibias.n449 161.3
R7807 commonsourceibias.n448 commonsourceibias.n409 161.3
R7808 commonsourceibias.n447 commonsourceibias.n446 161.3
R7809 commonsourceibias.n444 commonsourceibias.n410 161.3
R7810 commonsourceibias.n442 commonsourceibias.n441 161.3
R7811 commonsourceibias.n440 commonsourceibias.n411 161.3
R7812 commonsourceibias.n439 commonsourceibias.n438 161.3
R7813 commonsourceibias.n436 commonsourceibias.n412 161.3
R7814 commonsourceibias.n435 commonsourceibias.n434 161.3
R7815 commonsourceibias.n433 commonsourceibias.n432 161.3
R7816 commonsourceibias.n431 commonsourceibias.n414 161.3
R7817 commonsourceibias.n430 commonsourceibias.n429 161.3
R7818 commonsourceibias.n428 commonsourceibias.n427 161.3
R7819 commonsourceibias.n426 commonsourceibias.n416 161.3
R7820 commonsourceibias.n425 commonsourceibias.n424 161.3
R7821 commonsourceibias.n423 commonsourceibias.n422 161.3
R7822 commonsourceibias.n421 commonsourceibias.n418 161.3
R7823 commonsourceibias.n80 commonsourceibias.n78 81.5057
R7824 commonsourceibias.n304 commonsourceibias.n302 81.5057
R7825 commonsourceibias.n80 commonsourceibias.n79 80.9324
R7826 commonsourceibias.n82 commonsourceibias.n81 80.9324
R7827 commonsourceibias.n77 commonsourceibias.n76 80.9324
R7828 commonsourceibias.n75 commonsourceibias.n74 80.9324
R7829 commonsourceibias.n73 commonsourceibias.n72 80.9324
R7830 commonsourceibias.n371 commonsourceibias.n370 80.9324
R7831 commonsourceibias.n373 commonsourceibias.n372 80.9324
R7832 commonsourceibias.n375 commonsourceibias.n374 80.9324
R7833 commonsourceibias.n306 commonsourceibias.n305 80.9324
R7834 commonsourceibias.n304 commonsourceibias.n303 80.9324
R7835 commonsourceibias.n71 commonsourceibias.n70 80.6037
R7836 commonsourceibias.n137 commonsourceibias.n136 80.6037
R7837 commonsourceibias.n264 commonsourceibias.n263 80.6037
R7838 commonsourceibias.n200 commonsourceibias.n199 80.6037
R7839 commonsourceibias.n369 commonsourceibias.n368 80.6037
R7840 commonsourceibias.n403 commonsourceibias.n402 80.6037
R7841 commonsourceibias.n530 commonsourceibias.n529 80.6037
R7842 commonsourceibias.n466 commonsourceibias.n465 80.6037
R7843 commonsourceibias.n65 commonsourceibias.n64 56.5617
R7844 commonsourceibias.n51 commonsourceibias.n50 56.5617
R7845 commonsourceibias.n42 commonsourceibias.n41 56.5617
R7846 commonsourceibias.n28 commonsourceibias.n27 56.5617
R7847 commonsourceibias.n131 commonsourceibias.n130 56.5617
R7848 commonsourceibias.n117 commonsourceibias.n116 56.5617
R7849 commonsourceibias.n108 commonsourceibias.n107 56.5617
R7850 commonsourceibias.n94 commonsourceibias.n93 56.5617
R7851 commonsourceibias.n221 commonsourceibias.n220 56.5617
R7852 commonsourceibias.n235 commonsourceibias.n234 56.5617
R7853 commonsourceibias.n244 commonsourceibias.n243 56.5617
R7854 commonsourceibias.n258 commonsourceibias.n257 56.5617
R7855 commonsourceibias.n194 commonsourceibias.n193 56.5617
R7856 commonsourceibias.n180 commonsourceibias.n179 56.5617
R7857 commonsourceibias.n171 commonsourceibias.n170 56.5617
R7858 commonsourceibias.n157 commonsourceibias.n156 56.5617
R7859 commonsourceibias.n325 commonsourceibias.n324 56.5617
R7860 commonsourceibias.n339 commonsourceibias.n338 56.5617
R7861 commonsourceibias.n349 commonsourceibias.n347 56.5617
R7862 commonsourceibias.n363 commonsourceibias.n362 56.5617
R7863 commonsourceibias.n397 commonsourceibias.n396 56.5617
R7864 commonsourceibias.n383 commonsourceibias.n381 56.5617
R7865 commonsourceibias.n284 commonsourceibias.n283 56.5617
R7866 commonsourceibias.n298 commonsourceibias.n297 56.5617
R7867 commonsourceibias.n486 commonsourceibias.n485 56.5617
R7868 commonsourceibias.n500 commonsourceibias.n499 56.5617
R7869 commonsourceibias.n510 commonsourceibias.n508 56.5617
R7870 commonsourceibias.n524 commonsourceibias.n523 56.5617
R7871 commonsourceibias.n422 commonsourceibias.n421 56.5617
R7872 commonsourceibias.n436 commonsourceibias.n435 56.5617
R7873 commonsourceibias.n446 commonsourceibias.n444 56.5617
R7874 commonsourceibias.n460 commonsourceibias.n459 56.5617
R7875 commonsourceibias.n56 commonsourceibias.n55 56.0773
R7876 commonsourceibias.n37 commonsourceibias.n36 56.0773
R7877 commonsourceibias.n122 commonsourceibias.n121 56.0773
R7878 commonsourceibias.n103 commonsourceibias.n102 56.0773
R7879 commonsourceibias.n230 commonsourceibias.n229 56.0773
R7880 commonsourceibias.n249 commonsourceibias.n248 56.0773
R7881 commonsourceibias.n185 commonsourceibias.n184 56.0773
R7882 commonsourceibias.n166 commonsourceibias.n165 56.0773
R7883 commonsourceibias.n334 commonsourceibias.n333 56.0773
R7884 commonsourceibias.n354 commonsourceibias.n353 56.0773
R7885 commonsourceibias.n388 commonsourceibias.n387 56.0773
R7886 commonsourceibias.n293 commonsourceibias.n292 56.0773
R7887 commonsourceibias.n495 commonsourceibias.n494 56.0773
R7888 commonsourceibias.n515 commonsourceibias.n514 56.0773
R7889 commonsourceibias.n431 commonsourceibias.n430 56.0773
R7890 commonsourceibias.n451 commonsourceibias.n450 56.0773
R7891 commonsourceibias.n70 commonsourceibias.n69 46.0096
R7892 commonsourceibias.n136 commonsourceibias.n135 46.0096
R7893 commonsourceibias.n263 commonsourceibias.n262 46.0096
R7894 commonsourceibias.n199 commonsourceibias.n198 46.0096
R7895 commonsourceibias.n368 commonsourceibias.n367 46.0096
R7896 commonsourceibias.n402 commonsourceibias.n401 46.0096
R7897 commonsourceibias.n529 commonsourceibias.n528 46.0096
R7898 commonsourceibias.n465 commonsourceibias.n464 46.0096
R7899 commonsourceibias.n58 commonsourceibias.n12 41.5458
R7900 commonsourceibias.n33 commonsourceibias.n32 41.5458
R7901 commonsourceibias.n124 commonsourceibias.n3 41.5458
R7902 commonsourceibias.n99 commonsourceibias.n98 41.5458
R7903 commonsourceibias.n226 commonsourceibias.n225 41.5458
R7904 commonsourceibias.n251 commonsourceibias.n205 41.5458
R7905 commonsourceibias.n187 commonsourceibias.n141 41.5458
R7906 commonsourceibias.n162 commonsourceibias.n161 41.5458
R7907 commonsourceibias.n330 commonsourceibias.n329 41.5458
R7908 commonsourceibias.n356 commonsourceibias.n310 41.5458
R7909 commonsourceibias.n390 commonsourceibias.n269 41.5458
R7910 commonsourceibias.n289 commonsourceibias.n288 41.5458
R7911 commonsourceibias.n491 commonsourceibias.n490 41.5458
R7912 commonsourceibias.n517 commonsourceibias.n471 41.5458
R7913 commonsourceibias.n427 commonsourceibias.n426 41.5458
R7914 commonsourceibias.n453 commonsourceibias.n407 41.5458
R7915 commonsourceibias.n48 commonsourceibias.n17 40.577
R7916 commonsourceibias.n44 commonsourceibias.n17 40.577
R7917 commonsourceibias.n114 commonsourceibias.n8 40.577
R7918 commonsourceibias.n110 commonsourceibias.n8 40.577
R7919 commonsourceibias.n237 commonsourceibias.n210 40.577
R7920 commonsourceibias.n241 commonsourceibias.n210 40.577
R7921 commonsourceibias.n177 commonsourceibias.n146 40.577
R7922 commonsourceibias.n173 commonsourceibias.n146 40.577
R7923 commonsourceibias.n341 commonsourceibias.n314 40.577
R7924 commonsourceibias.n345 commonsourceibias.n314 40.577
R7925 commonsourceibias.n379 commonsourceibias.n273 40.577
R7926 commonsourceibias.n300 commonsourceibias.n273 40.577
R7927 commonsourceibias.n502 commonsourceibias.n475 40.577
R7928 commonsourceibias.n506 commonsourceibias.n475 40.577
R7929 commonsourceibias.n438 commonsourceibias.n411 40.577
R7930 commonsourceibias.n442 commonsourceibias.n411 40.577
R7931 commonsourceibias.n62 commonsourceibias.n12 39.6083
R7932 commonsourceibias.n32 commonsourceibias.n31 39.6083
R7933 commonsourceibias.n128 commonsourceibias.n3 39.6083
R7934 commonsourceibias.n98 commonsourceibias.n97 39.6083
R7935 commonsourceibias.n225 commonsourceibias.n224 39.6083
R7936 commonsourceibias.n255 commonsourceibias.n205 39.6083
R7937 commonsourceibias.n191 commonsourceibias.n141 39.6083
R7938 commonsourceibias.n161 commonsourceibias.n160 39.6083
R7939 commonsourceibias.n329 commonsourceibias.n328 39.6083
R7940 commonsourceibias.n360 commonsourceibias.n310 39.6083
R7941 commonsourceibias.n394 commonsourceibias.n269 39.6083
R7942 commonsourceibias.n288 commonsourceibias.n287 39.6083
R7943 commonsourceibias.n490 commonsourceibias.n489 39.6083
R7944 commonsourceibias.n521 commonsourceibias.n471 39.6083
R7945 commonsourceibias.n426 commonsourceibias.n425 39.6083
R7946 commonsourceibias.n457 commonsourceibias.n407 39.6083
R7947 commonsourceibias.n26 commonsourceibias.n25 33.0515
R7948 commonsourceibias.n92 commonsourceibias.n91 33.0515
R7949 commonsourceibias.n155 commonsourceibias.n154 33.0515
R7950 commonsourceibias.n219 commonsourceibias.n218 33.0515
R7951 commonsourceibias.n323 commonsourceibias.n322 33.0515
R7952 commonsourceibias.n282 commonsourceibias.n281 33.0515
R7953 commonsourceibias.n484 commonsourceibias.n483 33.0515
R7954 commonsourceibias.n420 commonsourceibias.n419 33.0515
R7955 commonsourceibias.n25 commonsourceibias.n24 28.5514
R7956 commonsourceibias.n91 commonsourceibias.n90 28.5514
R7957 commonsourceibias.n218 commonsourceibias.n217 28.5514
R7958 commonsourceibias.n154 commonsourceibias.n153 28.5514
R7959 commonsourceibias.n322 commonsourceibias.n321 28.5514
R7960 commonsourceibias.n281 commonsourceibias.n280 28.5514
R7961 commonsourceibias.n483 commonsourceibias.n482 28.5514
R7962 commonsourceibias.n419 commonsourceibias.n418 28.5514
R7963 commonsourceibias.n69 commonsourceibias.n68 26.0455
R7964 commonsourceibias.n135 commonsourceibias.n134 26.0455
R7965 commonsourceibias.n262 commonsourceibias.n261 26.0455
R7966 commonsourceibias.n198 commonsourceibias.n197 26.0455
R7967 commonsourceibias.n367 commonsourceibias.n366 26.0455
R7968 commonsourceibias.n401 commonsourceibias.n400 26.0455
R7969 commonsourceibias.n528 commonsourceibias.n527 26.0455
R7970 commonsourceibias.n464 commonsourceibias.n463 26.0455
R7971 commonsourceibias.n55 commonsourceibias.n14 25.0767
R7972 commonsourceibias.n38 commonsourceibias.n37 25.0767
R7973 commonsourceibias.n121 commonsourceibias.n5 25.0767
R7974 commonsourceibias.n104 commonsourceibias.n103 25.0767
R7975 commonsourceibias.n231 commonsourceibias.n230 25.0767
R7976 commonsourceibias.n248 commonsourceibias.n207 25.0767
R7977 commonsourceibias.n184 commonsourceibias.n143 25.0767
R7978 commonsourceibias.n167 commonsourceibias.n166 25.0767
R7979 commonsourceibias.n335 commonsourceibias.n334 25.0767
R7980 commonsourceibias.n353 commonsourceibias.n312 25.0767
R7981 commonsourceibias.n387 commonsourceibias.n271 25.0767
R7982 commonsourceibias.n294 commonsourceibias.n293 25.0767
R7983 commonsourceibias.n496 commonsourceibias.n495 25.0767
R7984 commonsourceibias.n514 commonsourceibias.n473 25.0767
R7985 commonsourceibias.n432 commonsourceibias.n431 25.0767
R7986 commonsourceibias.n450 commonsourceibias.n409 25.0767
R7987 commonsourceibias.n51 commonsourceibias.n16 24.3464
R7988 commonsourceibias.n41 commonsourceibias.n19 24.3464
R7989 commonsourceibias.n117 commonsourceibias.n7 24.3464
R7990 commonsourceibias.n107 commonsourceibias.n85 24.3464
R7991 commonsourceibias.n234 commonsourceibias.n212 24.3464
R7992 commonsourceibias.n244 commonsourceibias.n209 24.3464
R7993 commonsourceibias.n180 commonsourceibias.n145 24.3464
R7994 commonsourceibias.n170 commonsourceibias.n148 24.3464
R7995 commonsourceibias.n338 commonsourceibias.n316 24.3464
R7996 commonsourceibias.n349 commonsourceibias.n348 24.3464
R7997 commonsourceibias.n383 commonsourceibias.n382 24.3464
R7998 commonsourceibias.n297 commonsourceibias.n275 24.3464
R7999 commonsourceibias.n499 commonsourceibias.n477 24.3464
R8000 commonsourceibias.n510 commonsourceibias.n509 24.3464
R8001 commonsourceibias.n435 commonsourceibias.n413 24.3464
R8002 commonsourceibias.n446 commonsourceibias.n445 24.3464
R8003 commonsourceibias.n65 commonsourceibias.n10 23.8546
R8004 commonsourceibias.n27 commonsourceibias.n26 23.8546
R8005 commonsourceibias.n131 commonsourceibias.n1 23.8546
R8006 commonsourceibias.n93 commonsourceibias.n92 23.8546
R8007 commonsourceibias.n220 commonsourceibias.n219 23.8546
R8008 commonsourceibias.n258 commonsourceibias.n203 23.8546
R8009 commonsourceibias.n194 commonsourceibias.n139 23.8546
R8010 commonsourceibias.n156 commonsourceibias.n155 23.8546
R8011 commonsourceibias.n324 commonsourceibias.n323 23.8546
R8012 commonsourceibias.n363 commonsourceibias.n308 23.8546
R8013 commonsourceibias.n397 commonsourceibias.n267 23.8546
R8014 commonsourceibias.n283 commonsourceibias.n282 23.8546
R8015 commonsourceibias.n485 commonsourceibias.n484 23.8546
R8016 commonsourceibias.n524 commonsourceibias.n469 23.8546
R8017 commonsourceibias.n421 commonsourceibias.n420 23.8546
R8018 commonsourceibias.n460 commonsourceibias.n405 23.8546
R8019 commonsourceibias.n64 commonsourceibias.n63 16.9689
R8020 commonsourceibias.n28 commonsourceibias.n23 16.9689
R8021 commonsourceibias.n130 commonsourceibias.n129 16.9689
R8022 commonsourceibias.n94 commonsourceibias.n89 16.9689
R8023 commonsourceibias.n221 commonsourceibias.n216 16.9689
R8024 commonsourceibias.n257 commonsourceibias.n256 16.9689
R8025 commonsourceibias.n193 commonsourceibias.n192 16.9689
R8026 commonsourceibias.n157 commonsourceibias.n152 16.9689
R8027 commonsourceibias.n325 commonsourceibias.n320 16.9689
R8028 commonsourceibias.n362 commonsourceibias.n361 16.9689
R8029 commonsourceibias.n396 commonsourceibias.n395 16.9689
R8030 commonsourceibias.n284 commonsourceibias.n279 16.9689
R8031 commonsourceibias.n486 commonsourceibias.n481 16.9689
R8032 commonsourceibias.n523 commonsourceibias.n522 16.9689
R8033 commonsourceibias.n422 commonsourceibias.n417 16.9689
R8034 commonsourceibias.n459 commonsourceibias.n458 16.9689
R8035 commonsourceibias.n50 commonsourceibias.n49 16.477
R8036 commonsourceibias.n43 commonsourceibias.n42 16.477
R8037 commonsourceibias.n116 commonsourceibias.n115 16.477
R8038 commonsourceibias.n109 commonsourceibias.n108 16.477
R8039 commonsourceibias.n236 commonsourceibias.n235 16.477
R8040 commonsourceibias.n243 commonsourceibias.n242 16.477
R8041 commonsourceibias.n179 commonsourceibias.n178 16.477
R8042 commonsourceibias.n172 commonsourceibias.n171 16.477
R8043 commonsourceibias.n340 commonsourceibias.n339 16.477
R8044 commonsourceibias.n347 commonsourceibias.n346 16.477
R8045 commonsourceibias.n381 commonsourceibias.n380 16.477
R8046 commonsourceibias.n299 commonsourceibias.n298 16.477
R8047 commonsourceibias.n501 commonsourceibias.n500 16.477
R8048 commonsourceibias.n508 commonsourceibias.n507 16.477
R8049 commonsourceibias.n437 commonsourceibias.n436 16.477
R8050 commonsourceibias.n444 commonsourceibias.n443 16.477
R8051 commonsourceibias.n57 commonsourceibias.n56 15.9852
R8052 commonsourceibias.n36 commonsourceibias.n21 15.9852
R8053 commonsourceibias.n123 commonsourceibias.n122 15.9852
R8054 commonsourceibias.n102 commonsourceibias.n87 15.9852
R8055 commonsourceibias.n229 commonsourceibias.n214 15.9852
R8056 commonsourceibias.n250 commonsourceibias.n249 15.9852
R8057 commonsourceibias.n186 commonsourceibias.n185 15.9852
R8058 commonsourceibias.n165 commonsourceibias.n150 15.9852
R8059 commonsourceibias.n333 commonsourceibias.n318 15.9852
R8060 commonsourceibias.n355 commonsourceibias.n354 15.9852
R8061 commonsourceibias.n389 commonsourceibias.n388 15.9852
R8062 commonsourceibias.n292 commonsourceibias.n277 15.9852
R8063 commonsourceibias.n494 commonsourceibias.n479 15.9852
R8064 commonsourceibias.n516 commonsourceibias.n515 15.9852
R8065 commonsourceibias.n430 commonsourceibias.n415 15.9852
R8066 commonsourceibias.n452 commonsourceibias.n451 15.9852
R8067 commonsourceibias.n73 commonsourceibias.n71 13.2057
R8068 commonsourceibias.n371 commonsourceibias.n369 13.2057
R8069 commonsourceibias.n532 commonsourceibias.n265 10.4122
R8070 commonsourceibias.n112 commonsourceibias.n83 9.50363
R8071 commonsourceibias.n377 commonsourceibias.n376 9.50363
R8072 commonsourceibias.n201 commonsourceibias.n137 8.7339
R8073 commonsourceibias.n467 commonsourceibias.n403 8.7339
R8074 commonsourceibias.n58 commonsourceibias.n57 8.60764
R8075 commonsourceibias.n33 commonsourceibias.n21 8.60764
R8076 commonsourceibias.n124 commonsourceibias.n123 8.60764
R8077 commonsourceibias.n99 commonsourceibias.n87 8.60764
R8078 commonsourceibias.n226 commonsourceibias.n214 8.60764
R8079 commonsourceibias.n251 commonsourceibias.n250 8.60764
R8080 commonsourceibias.n187 commonsourceibias.n186 8.60764
R8081 commonsourceibias.n162 commonsourceibias.n150 8.60764
R8082 commonsourceibias.n330 commonsourceibias.n318 8.60764
R8083 commonsourceibias.n356 commonsourceibias.n355 8.60764
R8084 commonsourceibias.n390 commonsourceibias.n389 8.60764
R8085 commonsourceibias.n289 commonsourceibias.n277 8.60764
R8086 commonsourceibias.n491 commonsourceibias.n479 8.60764
R8087 commonsourceibias.n517 commonsourceibias.n516 8.60764
R8088 commonsourceibias.n427 commonsourceibias.n415 8.60764
R8089 commonsourceibias.n453 commonsourceibias.n452 8.60764
R8090 commonsourceibias.n532 commonsourceibias.n531 8.46921
R8091 commonsourceibias.n49 commonsourceibias.n48 8.11581
R8092 commonsourceibias.n44 commonsourceibias.n43 8.11581
R8093 commonsourceibias.n115 commonsourceibias.n114 8.11581
R8094 commonsourceibias.n110 commonsourceibias.n109 8.11581
R8095 commonsourceibias.n237 commonsourceibias.n236 8.11581
R8096 commonsourceibias.n242 commonsourceibias.n241 8.11581
R8097 commonsourceibias.n178 commonsourceibias.n177 8.11581
R8098 commonsourceibias.n173 commonsourceibias.n172 8.11581
R8099 commonsourceibias.n341 commonsourceibias.n340 8.11581
R8100 commonsourceibias.n346 commonsourceibias.n345 8.11581
R8101 commonsourceibias.n380 commonsourceibias.n379 8.11581
R8102 commonsourceibias.n300 commonsourceibias.n299 8.11581
R8103 commonsourceibias.n502 commonsourceibias.n501 8.11581
R8104 commonsourceibias.n507 commonsourceibias.n506 8.11581
R8105 commonsourceibias.n438 commonsourceibias.n437 8.11581
R8106 commonsourceibias.n443 commonsourceibias.n442 8.11581
R8107 commonsourceibias.n63 commonsourceibias.n62 7.62397
R8108 commonsourceibias.n31 commonsourceibias.n23 7.62397
R8109 commonsourceibias.n129 commonsourceibias.n128 7.62397
R8110 commonsourceibias.n97 commonsourceibias.n89 7.62397
R8111 commonsourceibias.n224 commonsourceibias.n216 7.62397
R8112 commonsourceibias.n256 commonsourceibias.n255 7.62397
R8113 commonsourceibias.n192 commonsourceibias.n191 7.62397
R8114 commonsourceibias.n160 commonsourceibias.n152 7.62397
R8115 commonsourceibias.n328 commonsourceibias.n320 7.62397
R8116 commonsourceibias.n361 commonsourceibias.n360 7.62397
R8117 commonsourceibias.n395 commonsourceibias.n394 7.62397
R8118 commonsourceibias.n287 commonsourceibias.n279 7.62397
R8119 commonsourceibias.n489 commonsourceibias.n481 7.62397
R8120 commonsourceibias.n522 commonsourceibias.n521 7.62397
R8121 commonsourceibias.n425 commonsourceibias.n417 7.62397
R8122 commonsourceibias.n458 commonsourceibias.n457 7.62397
R8123 commonsourceibias.n265 commonsourceibias.n264 5.00473
R8124 commonsourceibias.n201 commonsourceibias.n200 5.00473
R8125 commonsourceibias.n531 commonsourceibias.n530 5.00473
R8126 commonsourceibias.n467 commonsourceibias.n466 5.00473
R8127 commonsourceibias commonsourceibias.n532 3.87639
R8128 commonsourceibias.n265 commonsourceibias.n201 3.72967
R8129 commonsourceibias.n531 commonsourceibias.n467 3.72967
R8130 commonsourceibias.n78 commonsourceibias.t47 2.82907
R8131 commonsourceibias.n78 commonsourceibias.t39 2.82907
R8132 commonsourceibias.n79 commonsourceibias.t7 2.82907
R8133 commonsourceibias.n79 commonsourceibias.t19 2.82907
R8134 commonsourceibias.n81 commonsourceibias.t35 2.82907
R8135 commonsourceibias.n81 commonsourceibias.t15 2.82907
R8136 commonsourceibias.n76 commonsourceibias.t17 2.82907
R8137 commonsourceibias.n76 commonsourceibias.t23 2.82907
R8138 commonsourceibias.n74 commonsourceibias.t43 2.82907
R8139 commonsourceibias.n74 commonsourceibias.t41 2.82907
R8140 commonsourceibias.n72 commonsourceibias.t29 2.82907
R8141 commonsourceibias.n72 commonsourceibias.t5 2.82907
R8142 commonsourceibias.n370 commonsourceibias.t21 2.82907
R8143 commonsourceibias.n370 commonsourceibias.t9 2.82907
R8144 commonsourceibias.n372 commonsourceibias.t37 2.82907
R8145 commonsourceibias.n372 commonsourceibias.t25 2.82907
R8146 commonsourceibias.n374 commonsourceibias.t11 2.82907
R8147 commonsourceibias.n374 commonsourceibias.t33 2.82907
R8148 commonsourceibias.n305 commonsourceibias.t31 2.82907
R8149 commonsourceibias.n305 commonsourceibias.t1 2.82907
R8150 commonsourceibias.n303 commonsourceibias.t3 2.82907
R8151 commonsourceibias.n303 commonsourceibias.t13 2.82907
R8152 commonsourceibias.n302 commonsourceibias.t45 2.82907
R8153 commonsourceibias.n302 commonsourceibias.t27 2.82907
R8154 commonsourceibias.n68 commonsourceibias.n10 0.738255
R8155 commonsourceibias.n134 commonsourceibias.n1 0.738255
R8156 commonsourceibias.n261 commonsourceibias.n203 0.738255
R8157 commonsourceibias.n197 commonsourceibias.n139 0.738255
R8158 commonsourceibias.n366 commonsourceibias.n308 0.738255
R8159 commonsourceibias.n400 commonsourceibias.n267 0.738255
R8160 commonsourceibias.n527 commonsourceibias.n469 0.738255
R8161 commonsourceibias.n463 commonsourceibias.n405 0.738255
R8162 commonsourceibias.n75 commonsourceibias.n73 0.573776
R8163 commonsourceibias.n77 commonsourceibias.n75 0.573776
R8164 commonsourceibias.n82 commonsourceibias.n80 0.573776
R8165 commonsourceibias.n306 commonsourceibias.n304 0.573776
R8166 commonsourceibias.n375 commonsourceibias.n373 0.573776
R8167 commonsourceibias.n373 commonsourceibias.n371 0.573776
R8168 commonsourceibias.n83 commonsourceibias.n77 0.287138
R8169 commonsourceibias.n83 commonsourceibias.n82 0.287138
R8170 commonsourceibias.n376 commonsourceibias.n306 0.287138
R8171 commonsourceibias.n376 commonsourceibias.n375 0.287138
R8172 commonsourceibias.n71 commonsourceibias.n9 0.285035
R8173 commonsourceibias.n137 commonsourceibias.n0 0.285035
R8174 commonsourceibias.n264 commonsourceibias.n202 0.285035
R8175 commonsourceibias.n200 commonsourceibias.n138 0.285035
R8176 commonsourceibias.n369 commonsourceibias.n307 0.285035
R8177 commonsourceibias.n403 commonsourceibias.n266 0.285035
R8178 commonsourceibias.n530 commonsourceibias.n468 0.285035
R8179 commonsourceibias.n466 commonsourceibias.n404 0.285035
R8180 commonsourceibias.n16 commonsourceibias.n14 0.246418
R8181 commonsourceibias.n38 commonsourceibias.n19 0.246418
R8182 commonsourceibias.n7 commonsourceibias.n5 0.246418
R8183 commonsourceibias.n104 commonsourceibias.n85 0.246418
R8184 commonsourceibias.n231 commonsourceibias.n212 0.246418
R8185 commonsourceibias.n209 commonsourceibias.n207 0.246418
R8186 commonsourceibias.n145 commonsourceibias.n143 0.246418
R8187 commonsourceibias.n167 commonsourceibias.n148 0.246418
R8188 commonsourceibias.n335 commonsourceibias.n316 0.246418
R8189 commonsourceibias.n348 commonsourceibias.n312 0.246418
R8190 commonsourceibias.n382 commonsourceibias.n271 0.246418
R8191 commonsourceibias.n294 commonsourceibias.n275 0.246418
R8192 commonsourceibias.n496 commonsourceibias.n477 0.246418
R8193 commonsourceibias.n509 commonsourceibias.n473 0.246418
R8194 commonsourceibias.n432 commonsourceibias.n413 0.246418
R8195 commonsourceibias.n445 commonsourceibias.n409 0.246418
R8196 commonsourceibias.n67 commonsourceibias.n9 0.189894
R8197 commonsourceibias.n67 commonsourceibias.n66 0.189894
R8198 commonsourceibias.n66 commonsourceibias.n11 0.189894
R8199 commonsourceibias.n61 commonsourceibias.n11 0.189894
R8200 commonsourceibias.n61 commonsourceibias.n60 0.189894
R8201 commonsourceibias.n60 commonsourceibias.n59 0.189894
R8202 commonsourceibias.n59 commonsourceibias.n13 0.189894
R8203 commonsourceibias.n54 commonsourceibias.n13 0.189894
R8204 commonsourceibias.n54 commonsourceibias.n53 0.189894
R8205 commonsourceibias.n53 commonsourceibias.n52 0.189894
R8206 commonsourceibias.n52 commonsourceibias.n15 0.189894
R8207 commonsourceibias.n47 commonsourceibias.n15 0.189894
R8208 commonsourceibias.n47 commonsourceibias.n46 0.189894
R8209 commonsourceibias.n46 commonsourceibias.n45 0.189894
R8210 commonsourceibias.n45 commonsourceibias.n18 0.189894
R8211 commonsourceibias.n40 commonsourceibias.n18 0.189894
R8212 commonsourceibias.n40 commonsourceibias.n39 0.189894
R8213 commonsourceibias.n39 commonsourceibias.n20 0.189894
R8214 commonsourceibias.n35 commonsourceibias.n20 0.189894
R8215 commonsourceibias.n35 commonsourceibias.n34 0.189894
R8216 commonsourceibias.n34 commonsourceibias.n22 0.189894
R8217 commonsourceibias.n30 commonsourceibias.n22 0.189894
R8218 commonsourceibias.n30 commonsourceibias.n29 0.189894
R8219 commonsourceibias.n29 commonsourceibias.n24 0.189894
R8220 commonsourceibias.n111 commonsourceibias.n84 0.189894
R8221 commonsourceibias.n106 commonsourceibias.n84 0.189894
R8222 commonsourceibias.n106 commonsourceibias.n105 0.189894
R8223 commonsourceibias.n105 commonsourceibias.n86 0.189894
R8224 commonsourceibias.n101 commonsourceibias.n86 0.189894
R8225 commonsourceibias.n101 commonsourceibias.n100 0.189894
R8226 commonsourceibias.n100 commonsourceibias.n88 0.189894
R8227 commonsourceibias.n96 commonsourceibias.n88 0.189894
R8228 commonsourceibias.n96 commonsourceibias.n95 0.189894
R8229 commonsourceibias.n95 commonsourceibias.n90 0.189894
R8230 commonsourceibias.n133 commonsourceibias.n0 0.189894
R8231 commonsourceibias.n133 commonsourceibias.n132 0.189894
R8232 commonsourceibias.n132 commonsourceibias.n2 0.189894
R8233 commonsourceibias.n127 commonsourceibias.n2 0.189894
R8234 commonsourceibias.n127 commonsourceibias.n126 0.189894
R8235 commonsourceibias.n126 commonsourceibias.n125 0.189894
R8236 commonsourceibias.n125 commonsourceibias.n4 0.189894
R8237 commonsourceibias.n120 commonsourceibias.n4 0.189894
R8238 commonsourceibias.n120 commonsourceibias.n119 0.189894
R8239 commonsourceibias.n119 commonsourceibias.n118 0.189894
R8240 commonsourceibias.n118 commonsourceibias.n6 0.189894
R8241 commonsourceibias.n113 commonsourceibias.n6 0.189894
R8242 commonsourceibias.n260 commonsourceibias.n202 0.189894
R8243 commonsourceibias.n260 commonsourceibias.n259 0.189894
R8244 commonsourceibias.n259 commonsourceibias.n204 0.189894
R8245 commonsourceibias.n254 commonsourceibias.n204 0.189894
R8246 commonsourceibias.n254 commonsourceibias.n253 0.189894
R8247 commonsourceibias.n253 commonsourceibias.n252 0.189894
R8248 commonsourceibias.n252 commonsourceibias.n206 0.189894
R8249 commonsourceibias.n247 commonsourceibias.n206 0.189894
R8250 commonsourceibias.n247 commonsourceibias.n246 0.189894
R8251 commonsourceibias.n246 commonsourceibias.n245 0.189894
R8252 commonsourceibias.n245 commonsourceibias.n208 0.189894
R8253 commonsourceibias.n240 commonsourceibias.n208 0.189894
R8254 commonsourceibias.n240 commonsourceibias.n239 0.189894
R8255 commonsourceibias.n239 commonsourceibias.n238 0.189894
R8256 commonsourceibias.n238 commonsourceibias.n211 0.189894
R8257 commonsourceibias.n233 commonsourceibias.n211 0.189894
R8258 commonsourceibias.n233 commonsourceibias.n232 0.189894
R8259 commonsourceibias.n232 commonsourceibias.n213 0.189894
R8260 commonsourceibias.n228 commonsourceibias.n213 0.189894
R8261 commonsourceibias.n228 commonsourceibias.n227 0.189894
R8262 commonsourceibias.n227 commonsourceibias.n215 0.189894
R8263 commonsourceibias.n223 commonsourceibias.n215 0.189894
R8264 commonsourceibias.n223 commonsourceibias.n222 0.189894
R8265 commonsourceibias.n222 commonsourceibias.n217 0.189894
R8266 commonsourceibias.n196 commonsourceibias.n138 0.189894
R8267 commonsourceibias.n196 commonsourceibias.n195 0.189894
R8268 commonsourceibias.n195 commonsourceibias.n140 0.189894
R8269 commonsourceibias.n190 commonsourceibias.n140 0.189894
R8270 commonsourceibias.n190 commonsourceibias.n189 0.189894
R8271 commonsourceibias.n189 commonsourceibias.n188 0.189894
R8272 commonsourceibias.n188 commonsourceibias.n142 0.189894
R8273 commonsourceibias.n183 commonsourceibias.n142 0.189894
R8274 commonsourceibias.n183 commonsourceibias.n182 0.189894
R8275 commonsourceibias.n182 commonsourceibias.n181 0.189894
R8276 commonsourceibias.n181 commonsourceibias.n144 0.189894
R8277 commonsourceibias.n176 commonsourceibias.n144 0.189894
R8278 commonsourceibias.n176 commonsourceibias.n175 0.189894
R8279 commonsourceibias.n175 commonsourceibias.n174 0.189894
R8280 commonsourceibias.n174 commonsourceibias.n147 0.189894
R8281 commonsourceibias.n169 commonsourceibias.n147 0.189894
R8282 commonsourceibias.n169 commonsourceibias.n168 0.189894
R8283 commonsourceibias.n168 commonsourceibias.n149 0.189894
R8284 commonsourceibias.n164 commonsourceibias.n149 0.189894
R8285 commonsourceibias.n164 commonsourceibias.n163 0.189894
R8286 commonsourceibias.n163 commonsourceibias.n151 0.189894
R8287 commonsourceibias.n159 commonsourceibias.n151 0.189894
R8288 commonsourceibias.n159 commonsourceibias.n158 0.189894
R8289 commonsourceibias.n158 commonsourceibias.n153 0.189894
R8290 commonsourceibias.n326 commonsourceibias.n321 0.189894
R8291 commonsourceibias.n327 commonsourceibias.n326 0.189894
R8292 commonsourceibias.n327 commonsourceibias.n319 0.189894
R8293 commonsourceibias.n331 commonsourceibias.n319 0.189894
R8294 commonsourceibias.n332 commonsourceibias.n331 0.189894
R8295 commonsourceibias.n332 commonsourceibias.n317 0.189894
R8296 commonsourceibias.n336 commonsourceibias.n317 0.189894
R8297 commonsourceibias.n337 commonsourceibias.n336 0.189894
R8298 commonsourceibias.n337 commonsourceibias.n315 0.189894
R8299 commonsourceibias.n342 commonsourceibias.n315 0.189894
R8300 commonsourceibias.n343 commonsourceibias.n342 0.189894
R8301 commonsourceibias.n344 commonsourceibias.n343 0.189894
R8302 commonsourceibias.n344 commonsourceibias.n313 0.189894
R8303 commonsourceibias.n350 commonsourceibias.n313 0.189894
R8304 commonsourceibias.n351 commonsourceibias.n350 0.189894
R8305 commonsourceibias.n352 commonsourceibias.n351 0.189894
R8306 commonsourceibias.n352 commonsourceibias.n311 0.189894
R8307 commonsourceibias.n357 commonsourceibias.n311 0.189894
R8308 commonsourceibias.n358 commonsourceibias.n357 0.189894
R8309 commonsourceibias.n359 commonsourceibias.n358 0.189894
R8310 commonsourceibias.n359 commonsourceibias.n309 0.189894
R8311 commonsourceibias.n364 commonsourceibias.n309 0.189894
R8312 commonsourceibias.n365 commonsourceibias.n364 0.189894
R8313 commonsourceibias.n365 commonsourceibias.n307 0.189894
R8314 commonsourceibias.n285 commonsourceibias.n280 0.189894
R8315 commonsourceibias.n286 commonsourceibias.n285 0.189894
R8316 commonsourceibias.n286 commonsourceibias.n278 0.189894
R8317 commonsourceibias.n290 commonsourceibias.n278 0.189894
R8318 commonsourceibias.n291 commonsourceibias.n290 0.189894
R8319 commonsourceibias.n291 commonsourceibias.n276 0.189894
R8320 commonsourceibias.n295 commonsourceibias.n276 0.189894
R8321 commonsourceibias.n296 commonsourceibias.n295 0.189894
R8322 commonsourceibias.n296 commonsourceibias.n274 0.189894
R8323 commonsourceibias.n301 commonsourceibias.n274 0.189894
R8324 commonsourceibias.n378 commonsourceibias.n272 0.189894
R8325 commonsourceibias.n384 commonsourceibias.n272 0.189894
R8326 commonsourceibias.n385 commonsourceibias.n384 0.189894
R8327 commonsourceibias.n386 commonsourceibias.n385 0.189894
R8328 commonsourceibias.n386 commonsourceibias.n270 0.189894
R8329 commonsourceibias.n391 commonsourceibias.n270 0.189894
R8330 commonsourceibias.n392 commonsourceibias.n391 0.189894
R8331 commonsourceibias.n393 commonsourceibias.n392 0.189894
R8332 commonsourceibias.n393 commonsourceibias.n268 0.189894
R8333 commonsourceibias.n398 commonsourceibias.n268 0.189894
R8334 commonsourceibias.n399 commonsourceibias.n398 0.189894
R8335 commonsourceibias.n399 commonsourceibias.n266 0.189894
R8336 commonsourceibias.n487 commonsourceibias.n482 0.189894
R8337 commonsourceibias.n488 commonsourceibias.n487 0.189894
R8338 commonsourceibias.n488 commonsourceibias.n480 0.189894
R8339 commonsourceibias.n492 commonsourceibias.n480 0.189894
R8340 commonsourceibias.n493 commonsourceibias.n492 0.189894
R8341 commonsourceibias.n493 commonsourceibias.n478 0.189894
R8342 commonsourceibias.n497 commonsourceibias.n478 0.189894
R8343 commonsourceibias.n498 commonsourceibias.n497 0.189894
R8344 commonsourceibias.n498 commonsourceibias.n476 0.189894
R8345 commonsourceibias.n503 commonsourceibias.n476 0.189894
R8346 commonsourceibias.n504 commonsourceibias.n503 0.189894
R8347 commonsourceibias.n505 commonsourceibias.n504 0.189894
R8348 commonsourceibias.n505 commonsourceibias.n474 0.189894
R8349 commonsourceibias.n511 commonsourceibias.n474 0.189894
R8350 commonsourceibias.n512 commonsourceibias.n511 0.189894
R8351 commonsourceibias.n513 commonsourceibias.n512 0.189894
R8352 commonsourceibias.n513 commonsourceibias.n472 0.189894
R8353 commonsourceibias.n518 commonsourceibias.n472 0.189894
R8354 commonsourceibias.n519 commonsourceibias.n518 0.189894
R8355 commonsourceibias.n520 commonsourceibias.n519 0.189894
R8356 commonsourceibias.n520 commonsourceibias.n470 0.189894
R8357 commonsourceibias.n525 commonsourceibias.n470 0.189894
R8358 commonsourceibias.n526 commonsourceibias.n525 0.189894
R8359 commonsourceibias.n526 commonsourceibias.n468 0.189894
R8360 commonsourceibias.n423 commonsourceibias.n418 0.189894
R8361 commonsourceibias.n424 commonsourceibias.n423 0.189894
R8362 commonsourceibias.n424 commonsourceibias.n416 0.189894
R8363 commonsourceibias.n428 commonsourceibias.n416 0.189894
R8364 commonsourceibias.n429 commonsourceibias.n428 0.189894
R8365 commonsourceibias.n429 commonsourceibias.n414 0.189894
R8366 commonsourceibias.n433 commonsourceibias.n414 0.189894
R8367 commonsourceibias.n434 commonsourceibias.n433 0.189894
R8368 commonsourceibias.n434 commonsourceibias.n412 0.189894
R8369 commonsourceibias.n439 commonsourceibias.n412 0.189894
R8370 commonsourceibias.n440 commonsourceibias.n439 0.189894
R8371 commonsourceibias.n441 commonsourceibias.n440 0.189894
R8372 commonsourceibias.n441 commonsourceibias.n410 0.189894
R8373 commonsourceibias.n447 commonsourceibias.n410 0.189894
R8374 commonsourceibias.n448 commonsourceibias.n447 0.189894
R8375 commonsourceibias.n449 commonsourceibias.n448 0.189894
R8376 commonsourceibias.n449 commonsourceibias.n408 0.189894
R8377 commonsourceibias.n454 commonsourceibias.n408 0.189894
R8378 commonsourceibias.n455 commonsourceibias.n454 0.189894
R8379 commonsourceibias.n456 commonsourceibias.n455 0.189894
R8380 commonsourceibias.n456 commonsourceibias.n406 0.189894
R8381 commonsourceibias.n461 commonsourceibias.n406 0.189894
R8382 commonsourceibias.n462 commonsourceibias.n461 0.189894
R8383 commonsourceibias.n462 commonsourceibias.n404 0.189894
R8384 commonsourceibias.n112 commonsourceibias.n111 0.170955
R8385 commonsourceibias.n113 commonsourceibias.n112 0.170955
R8386 commonsourceibias.n377 commonsourceibias.n301 0.170955
R8387 commonsourceibias.n378 commonsourceibias.n377 0.170955
R8388 gnd.n6666 gnd.n310 1552.66
R8389 gnd.n3703 gnd.n3702 939.716
R8390 gnd.n7246 gnd.n171 838.452
R8391 gnd.n7188 gnd.n169 838.452
R8392 gnd.n1492 gnd.n1380 838.452
R8393 gnd.n5464 gnd.n1494 838.452
R8394 gnd.n5984 gnd.n863 838.452
R8395 gnd.n5904 gnd.n861 838.452
R8396 gnd.n3771 gnd.n3705 838.452
R8397 gnd.n3998 gnd.n2240 838.452
R8398 gnd.n7248 gnd.n166 783.196
R8399 gnd.n7063 gnd.n168 783.196
R8400 gnd.n5467 gnd.n5466 783.196
R8401 gnd.n5584 gnd.n1426 783.196
R8402 gnd.n5986 gnd.n858 783.196
R8403 gnd.n1069 gnd.n860 783.196
R8404 gnd.n3877 gnd.n3704 783.196
R8405 gnd.n3996 gnd.n3781 783.196
R8406 gnd.n3610 gnd.n2242 766.379
R8407 gnd.n3613 gnd.n3612 766.379
R8408 gnd.n2852 gnd.n2755 766.379
R8409 gnd.n2848 gnd.n2753 766.379
R8410 gnd.n3701 gnd.n2264 756.769
R8411 gnd.n3604 gnd.n3603 756.769
R8412 gnd.n2945 gnd.n2662 756.769
R8413 gnd.n2943 gnd.n2665 756.769
R8414 gnd.n6244 gnd.n562 756.769
R8415 gnd.n6665 gnd.n311 756.769
R8416 gnd.n6877 gnd.n6876 756.769
R8417 gnd.n6068 gnd.n727 756.769
R8418 gnd.n5965 gnd.n893 711.122
R8419 gnd.n5653 gnd.n1316 711.122
R8420 gnd.n5969 gnd.n875 711.122
R8421 gnd.n5655 gnd.n1311 711.122
R8422 gnd.n6240 gnd.n562 585
R8423 gnd.n562 gnd.n561 585
R8424 gnd.n6239 gnd.n6238 585
R8425 gnd.n6238 gnd.n6237 585
R8426 gnd.n565 gnd.n564 585
R8427 gnd.n6236 gnd.n565 585
R8428 gnd.n6234 gnd.n6233 585
R8429 gnd.n6235 gnd.n6234 585
R8430 gnd.n6232 gnd.n567 585
R8431 gnd.n567 gnd.n566 585
R8432 gnd.n6231 gnd.n6230 585
R8433 gnd.n6230 gnd.n6229 585
R8434 gnd.n573 gnd.n572 585
R8435 gnd.n6228 gnd.n573 585
R8436 gnd.n6226 gnd.n6225 585
R8437 gnd.n6227 gnd.n6226 585
R8438 gnd.n6224 gnd.n575 585
R8439 gnd.n575 gnd.n574 585
R8440 gnd.n6223 gnd.n6222 585
R8441 gnd.n6222 gnd.n6221 585
R8442 gnd.n581 gnd.n580 585
R8443 gnd.n6220 gnd.n581 585
R8444 gnd.n6218 gnd.n6217 585
R8445 gnd.n6219 gnd.n6218 585
R8446 gnd.n6216 gnd.n583 585
R8447 gnd.n583 gnd.n582 585
R8448 gnd.n6215 gnd.n6214 585
R8449 gnd.n6214 gnd.n6213 585
R8450 gnd.n589 gnd.n588 585
R8451 gnd.n6212 gnd.n589 585
R8452 gnd.n6210 gnd.n6209 585
R8453 gnd.n6211 gnd.n6210 585
R8454 gnd.n6208 gnd.n591 585
R8455 gnd.n591 gnd.n590 585
R8456 gnd.n6207 gnd.n6206 585
R8457 gnd.n6206 gnd.n6205 585
R8458 gnd.n597 gnd.n596 585
R8459 gnd.n6204 gnd.n597 585
R8460 gnd.n6202 gnd.n6201 585
R8461 gnd.n6203 gnd.n6202 585
R8462 gnd.n6200 gnd.n599 585
R8463 gnd.n599 gnd.n598 585
R8464 gnd.n6199 gnd.n6198 585
R8465 gnd.n6198 gnd.n6197 585
R8466 gnd.n605 gnd.n604 585
R8467 gnd.n6196 gnd.n605 585
R8468 gnd.n6194 gnd.n6193 585
R8469 gnd.n6195 gnd.n6194 585
R8470 gnd.n6192 gnd.n607 585
R8471 gnd.n607 gnd.n606 585
R8472 gnd.n6191 gnd.n6190 585
R8473 gnd.n6190 gnd.n6189 585
R8474 gnd.n613 gnd.n612 585
R8475 gnd.n6188 gnd.n613 585
R8476 gnd.n6186 gnd.n6185 585
R8477 gnd.n6187 gnd.n6186 585
R8478 gnd.n6184 gnd.n615 585
R8479 gnd.n615 gnd.n614 585
R8480 gnd.n6183 gnd.n6182 585
R8481 gnd.n6182 gnd.n6181 585
R8482 gnd.n621 gnd.n620 585
R8483 gnd.n6180 gnd.n621 585
R8484 gnd.n6178 gnd.n6177 585
R8485 gnd.n6179 gnd.n6178 585
R8486 gnd.n6176 gnd.n623 585
R8487 gnd.n623 gnd.n622 585
R8488 gnd.n6175 gnd.n6174 585
R8489 gnd.n6174 gnd.n6173 585
R8490 gnd.n629 gnd.n628 585
R8491 gnd.n6172 gnd.n629 585
R8492 gnd.n6170 gnd.n6169 585
R8493 gnd.n6171 gnd.n6170 585
R8494 gnd.n6168 gnd.n631 585
R8495 gnd.n631 gnd.n630 585
R8496 gnd.n6167 gnd.n6166 585
R8497 gnd.n6166 gnd.n6165 585
R8498 gnd.n637 gnd.n636 585
R8499 gnd.n6164 gnd.n637 585
R8500 gnd.n6162 gnd.n6161 585
R8501 gnd.n6163 gnd.n6162 585
R8502 gnd.n6160 gnd.n639 585
R8503 gnd.n639 gnd.n638 585
R8504 gnd.n6159 gnd.n6158 585
R8505 gnd.n6158 gnd.n6157 585
R8506 gnd.n645 gnd.n644 585
R8507 gnd.n6156 gnd.n645 585
R8508 gnd.n6154 gnd.n6153 585
R8509 gnd.n6155 gnd.n6154 585
R8510 gnd.n6152 gnd.n647 585
R8511 gnd.n647 gnd.n646 585
R8512 gnd.n6151 gnd.n6150 585
R8513 gnd.n6150 gnd.n6149 585
R8514 gnd.n653 gnd.n652 585
R8515 gnd.n6148 gnd.n653 585
R8516 gnd.n6146 gnd.n6145 585
R8517 gnd.n6147 gnd.n6146 585
R8518 gnd.n6144 gnd.n655 585
R8519 gnd.n655 gnd.n654 585
R8520 gnd.n6143 gnd.n6142 585
R8521 gnd.n6142 gnd.n6141 585
R8522 gnd.n661 gnd.n660 585
R8523 gnd.n6140 gnd.n661 585
R8524 gnd.n6138 gnd.n6137 585
R8525 gnd.n6139 gnd.n6138 585
R8526 gnd.n6136 gnd.n663 585
R8527 gnd.n663 gnd.n662 585
R8528 gnd.n6135 gnd.n6134 585
R8529 gnd.n6134 gnd.n6133 585
R8530 gnd.n669 gnd.n668 585
R8531 gnd.n6132 gnd.n669 585
R8532 gnd.n6130 gnd.n6129 585
R8533 gnd.n6131 gnd.n6130 585
R8534 gnd.n6128 gnd.n671 585
R8535 gnd.n671 gnd.n670 585
R8536 gnd.n6127 gnd.n6126 585
R8537 gnd.n6126 gnd.n6125 585
R8538 gnd.n677 gnd.n676 585
R8539 gnd.n6124 gnd.n677 585
R8540 gnd.n6122 gnd.n6121 585
R8541 gnd.n6123 gnd.n6122 585
R8542 gnd.n6120 gnd.n679 585
R8543 gnd.n679 gnd.n678 585
R8544 gnd.n6119 gnd.n6118 585
R8545 gnd.n6118 gnd.n6117 585
R8546 gnd.n685 gnd.n684 585
R8547 gnd.n6116 gnd.n685 585
R8548 gnd.n6114 gnd.n6113 585
R8549 gnd.n6115 gnd.n6114 585
R8550 gnd.n6112 gnd.n687 585
R8551 gnd.n687 gnd.n686 585
R8552 gnd.n6111 gnd.n6110 585
R8553 gnd.n6110 gnd.n6109 585
R8554 gnd.n693 gnd.n692 585
R8555 gnd.n6108 gnd.n693 585
R8556 gnd.n6106 gnd.n6105 585
R8557 gnd.n6107 gnd.n6106 585
R8558 gnd.n6104 gnd.n695 585
R8559 gnd.n695 gnd.n694 585
R8560 gnd.n6103 gnd.n6102 585
R8561 gnd.n6102 gnd.n6101 585
R8562 gnd.n701 gnd.n700 585
R8563 gnd.n6100 gnd.n701 585
R8564 gnd.n6098 gnd.n6097 585
R8565 gnd.n6099 gnd.n6098 585
R8566 gnd.n6096 gnd.n703 585
R8567 gnd.n703 gnd.n702 585
R8568 gnd.n6095 gnd.n6094 585
R8569 gnd.n6094 gnd.n6093 585
R8570 gnd.n709 gnd.n708 585
R8571 gnd.n6092 gnd.n709 585
R8572 gnd.n6090 gnd.n6089 585
R8573 gnd.n6091 gnd.n6090 585
R8574 gnd.n6088 gnd.n711 585
R8575 gnd.n711 gnd.n710 585
R8576 gnd.n6087 gnd.n6086 585
R8577 gnd.n6086 gnd.n6085 585
R8578 gnd.n717 gnd.n716 585
R8579 gnd.n6084 gnd.n717 585
R8580 gnd.n6082 gnd.n6081 585
R8581 gnd.n6083 gnd.n6082 585
R8582 gnd.n6080 gnd.n719 585
R8583 gnd.n719 gnd.n718 585
R8584 gnd.n6079 gnd.n6078 585
R8585 gnd.n6078 gnd.n6077 585
R8586 gnd.n725 gnd.n724 585
R8587 gnd.n6076 gnd.n725 585
R8588 gnd.n6074 gnd.n6073 585
R8589 gnd.n6075 gnd.n6074 585
R8590 gnd.n6244 gnd.n6243 585
R8591 gnd.n6245 gnd.n6244 585
R8592 gnd.n560 gnd.n559 585
R8593 gnd.n6246 gnd.n560 585
R8594 gnd.n6249 gnd.n6248 585
R8595 gnd.n6248 gnd.n6247 585
R8596 gnd.n557 gnd.n556 585
R8597 gnd.n556 gnd.n555 585
R8598 gnd.n6254 gnd.n6253 585
R8599 gnd.n6255 gnd.n6254 585
R8600 gnd.n554 gnd.n553 585
R8601 gnd.n6256 gnd.n554 585
R8602 gnd.n6259 gnd.n6258 585
R8603 gnd.n6258 gnd.n6257 585
R8604 gnd.n551 gnd.n550 585
R8605 gnd.n550 gnd.n549 585
R8606 gnd.n6264 gnd.n6263 585
R8607 gnd.n6265 gnd.n6264 585
R8608 gnd.n548 gnd.n547 585
R8609 gnd.n6266 gnd.n548 585
R8610 gnd.n6269 gnd.n6268 585
R8611 gnd.n6268 gnd.n6267 585
R8612 gnd.n545 gnd.n544 585
R8613 gnd.n544 gnd.n543 585
R8614 gnd.n6274 gnd.n6273 585
R8615 gnd.n6275 gnd.n6274 585
R8616 gnd.n542 gnd.n541 585
R8617 gnd.n6276 gnd.n542 585
R8618 gnd.n6279 gnd.n6278 585
R8619 gnd.n6278 gnd.n6277 585
R8620 gnd.n539 gnd.n538 585
R8621 gnd.n538 gnd.n537 585
R8622 gnd.n6284 gnd.n6283 585
R8623 gnd.n6285 gnd.n6284 585
R8624 gnd.n536 gnd.n535 585
R8625 gnd.n6286 gnd.n536 585
R8626 gnd.n6289 gnd.n6288 585
R8627 gnd.n6288 gnd.n6287 585
R8628 gnd.n533 gnd.n532 585
R8629 gnd.n532 gnd.n531 585
R8630 gnd.n6294 gnd.n6293 585
R8631 gnd.n6295 gnd.n6294 585
R8632 gnd.n530 gnd.n529 585
R8633 gnd.n6296 gnd.n530 585
R8634 gnd.n6299 gnd.n6298 585
R8635 gnd.n6298 gnd.n6297 585
R8636 gnd.n527 gnd.n526 585
R8637 gnd.n526 gnd.n525 585
R8638 gnd.n6304 gnd.n6303 585
R8639 gnd.n6305 gnd.n6304 585
R8640 gnd.n524 gnd.n523 585
R8641 gnd.n6306 gnd.n524 585
R8642 gnd.n6309 gnd.n6308 585
R8643 gnd.n6308 gnd.n6307 585
R8644 gnd.n521 gnd.n520 585
R8645 gnd.n520 gnd.n519 585
R8646 gnd.n6314 gnd.n6313 585
R8647 gnd.n6315 gnd.n6314 585
R8648 gnd.n518 gnd.n517 585
R8649 gnd.n6316 gnd.n518 585
R8650 gnd.n6319 gnd.n6318 585
R8651 gnd.n6318 gnd.n6317 585
R8652 gnd.n515 gnd.n514 585
R8653 gnd.n514 gnd.n513 585
R8654 gnd.n6324 gnd.n6323 585
R8655 gnd.n6325 gnd.n6324 585
R8656 gnd.n512 gnd.n511 585
R8657 gnd.n6326 gnd.n512 585
R8658 gnd.n6329 gnd.n6328 585
R8659 gnd.n6328 gnd.n6327 585
R8660 gnd.n509 gnd.n508 585
R8661 gnd.n508 gnd.n507 585
R8662 gnd.n6334 gnd.n6333 585
R8663 gnd.n6335 gnd.n6334 585
R8664 gnd.n506 gnd.n505 585
R8665 gnd.n6336 gnd.n506 585
R8666 gnd.n6339 gnd.n6338 585
R8667 gnd.n6338 gnd.n6337 585
R8668 gnd.n503 gnd.n502 585
R8669 gnd.n502 gnd.n501 585
R8670 gnd.n6344 gnd.n6343 585
R8671 gnd.n6345 gnd.n6344 585
R8672 gnd.n500 gnd.n499 585
R8673 gnd.n6346 gnd.n500 585
R8674 gnd.n6349 gnd.n6348 585
R8675 gnd.n6348 gnd.n6347 585
R8676 gnd.n497 gnd.n496 585
R8677 gnd.n496 gnd.n495 585
R8678 gnd.n6354 gnd.n6353 585
R8679 gnd.n6355 gnd.n6354 585
R8680 gnd.n494 gnd.n493 585
R8681 gnd.n6356 gnd.n494 585
R8682 gnd.n6359 gnd.n6358 585
R8683 gnd.n6358 gnd.n6357 585
R8684 gnd.n491 gnd.n490 585
R8685 gnd.n490 gnd.n489 585
R8686 gnd.n6364 gnd.n6363 585
R8687 gnd.n6365 gnd.n6364 585
R8688 gnd.n488 gnd.n487 585
R8689 gnd.n6366 gnd.n488 585
R8690 gnd.n6369 gnd.n6368 585
R8691 gnd.n6368 gnd.n6367 585
R8692 gnd.n485 gnd.n484 585
R8693 gnd.n484 gnd.n483 585
R8694 gnd.n6374 gnd.n6373 585
R8695 gnd.n6375 gnd.n6374 585
R8696 gnd.n482 gnd.n481 585
R8697 gnd.n6376 gnd.n482 585
R8698 gnd.n6379 gnd.n6378 585
R8699 gnd.n6378 gnd.n6377 585
R8700 gnd.n479 gnd.n478 585
R8701 gnd.n478 gnd.n477 585
R8702 gnd.n6384 gnd.n6383 585
R8703 gnd.n6385 gnd.n6384 585
R8704 gnd.n476 gnd.n475 585
R8705 gnd.n6386 gnd.n476 585
R8706 gnd.n6389 gnd.n6388 585
R8707 gnd.n6388 gnd.n6387 585
R8708 gnd.n473 gnd.n472 585
R8709 gnd.n472 gnd.n471 585
R8710 gnd.n6394 gnd.n6393 585
R8711 gnd.n6395 gnd.n6394 585
R8712 gnd.n470 gnd.n469 585
R8713 gnd.n6396 gnd.n470 585
R8714 gnd.n6399 gnd.n6398 585
R8715 gnd.n6398 gnd.n6397 585
R8716 gnd.n467 gnd.n466 585
R8717 gnd.n466 gnd.n465 585
R8718 gnd.n6404 gnd.n6403 585
R8719 gnd.n6405 gnd.n6404 585
R8720 gnd.n464 gnd.n463 585
R8721 gnd.n6406 gnd.n464 585
R8722 gnd.n6409 gnd.n6408 585
R8723 gnd.n6408 gnd.n6407 585
R8724 gnd.n461 gnd.n460 585
R8725 gnd.n460 gnd.n459 585
R8726 gnd.n6414 gnd.n6413 585
R8727 gnd.n6415 gnd.n6414 585
R8728 gnd.n458 gnd.n457 585
R8729 gnd.n6416 gnd.n458 585
R8730 gnd.n6419 gnd.n6418 585
R8731 gnd.n6418 gnd.n6417 585
R8732 gnd.n455 gnd.n454 585
R8733 gnd.n454 gnd.n453 585
R8734 gnd.n6424 gnd.n6423 585
R8735 gnd.n6425 gnd.n6424 585
R8736 gnd.n452 gnd.n451 585
R8737 gnd.n6426 gnd.n452 585
R8738 gnd.n6429 gnd.n6428 585
R8739 gnd.n6428 gnd.n6427 585
R8740 gnd.n449 gnd.n448 585
R8741 gnd.n448 gnd.n447 585
R8742 gnd.n6434 gnd.n6433 585
R8743 gnd.n6435 gnd.n6434 585
R8744 gnd.n446 gnd.n445 585
R8745 gnd.n6436 gnd.n446 585
R8746 gnd.n6439 gnd.n6438 585
R8747 gnd.n6438 gnd.n6437 585
R8748 gnd.n443 gnd.n442 585
R8749 gnd.n442 gnd.n441 585
R8750 gnd.n6444 gnd.n6443 585
R8751 gnd.n6445 gnd.n6444 585
R8752 gnd.n440 gnd.n439 585
R8753 gnd.n6446 gnd.n440 585
R8754 gnd.n6449 gnd.n6448 585
R8755 gnd.n6448 gnd.n6447 585
R8756 gnd.n437 gnd.n436 585
R8757 gnd.n436 gnd.n435 585
R8758 gnd.n6454 gnd.n6453 585
R8759 gnd.n6455 gnd.n6454 585
R8760 gnd.n434 gnd.n433 585
R8761 gnd.n6456 gnd.n434 585
R8762 gnd.n6459 gnd.n6458 585
R8763 gnd.n6458 gnd.n6457 585
R8764 gnd.n431 gnd.n430 585
R8765 gnd.n430 gnd.n429 585
R8766 gnd.n6464 gnd.n6463 585
R8767 gnd.n6465 gnd.n6464 585
R8768 gnd.n428 gnd.n427 585
R8769 gnd.n6466 gnd.n428 585
R8770 gnd.n6469 gnd.n6468 585
R8771 gnd.n6468 gnd.n6467 585
R8772 gnd.n425 gnd.n424 585
R8773 gnd.n424 gnd.n423 585
R8774 gnd.n6474 gnd.n6473 585
R8775 gnd.n6475 gnd.n6474 585
R8776 gnd.n422 gnd.n421 585
R8777 gnd.n6476 gnd.n422 585
R8778 gnd.n6479 gnd.n6478 585
R8779 gnd.n6478 gnd.n6477 585
R8780 gnd.n419 gnd.n418 585
R8781 gnd.n418 gnd.n417 585
R8782 gnd.n6484 gnd.n6483 585
R8783 gnd.n6485 gnd.n6484 585
R8784 gnd.n416 gnd.n415 585
R8785 gnd.n6486 gnd.n416 585
R8786 gnd.n6489 gnd.n6488 585
R8787 gnd.n6488 gnd.n6487 585
R8788 gnd.n413 gnd.n412 585
R8789 gnd.n412 gnd.n411 585
R8790 gnd.n6494 gnd.n6493 585
R8791 gnd.n6495 gnd.n6494 585
R8792 gnd.n410 gnd.n409 585
R8793 gnd.n6496 gnd.n410 585
R8794 gnd.n6499 gnd.n6498 585
R8795 gnd.n6498 gnd.n6497 585
R8796 gnd.n407 gnd.n406 585
R8797 gnd.n406 gnd.n405 585
R8798 gnd.n6504 gnd.n6503 585
R8799 gnd.n6505 gnd.n6504 585
R8800 gnd.n404 gnd.n403 585
R8801 gnd.n6506 gnd.n404 585
R8802 gnd.n6509 gnd.n6508 585
R8803 gnd.n6508 gnd.n6507 585
R8804 gnd.n401 gnd.n400 585
R8805 gnd.n400 gnd.n399 585
R8806 gnd.n6514 gnd.n6513 585
R8807 gnd.n6515 gnd.n6514 585
R8808 gnd.n398 gnd.n397 585
R8809 gnd.n6516 gnd.n398 585
R8810 gnd.n6519 gnd.n6518 585
R8811 gnd.n6518 gnd.n6517 585
R8812 gnd.n395 gnd.n394 585
R8813 gnd.n394 gnd.n393 585
R8814 gnd.n6524 gnd.n6523 585
R8815 gnd.n6525 gnd.n6524 585
R8816 gnd.n392 gnd.n391 585
R8817 gnd.n6526 gnd.n392 585
R8818 gnd.n6529 gnd.n6528 585
R8819 gnd.n6528 gnd.n6527 585
R8820 gnd.n389 gnd.n388 585
R8821 gnd.n388 gnd.n387 585
R8822 gnd.n6534 gnd.n6533 585
R8823 gnd.n6535 gnd.n6534 585
R8824 gnd.n386 gnd.n385 585
R8825 gnd.n6536 gnd.n386 585
R8826 gnd.n6539 gnd.n6538 585
R8827 gnd.n6538 gnd.n6537 585
R8828 gnd.n383 gnd.n382 585
R8829 gnd.n382 gnd.n381 585
R8830 gnd.n6544 gnd.n6543 585
R8831 gnd.n6545 gnd.n6544 585
R8832 gnd.n380 gnd.n379 585
R8833 gnd.n6546 gnd.n380 585
R8834 gnd.n6549 gnd.n6548 585
R8835 gnd.n6548 gnd.n6547 585
R8836 gnd.n377 gnd.n376 585
R8837 gnd.n376 gnd.n375 585
R8838 gnd.n6554 gnd.n6553 585
R8839 gnd.n6555 gnd.n6554 585
R8840 gnd.n374 gnd.n373 585
R8841 gnd.n6556 gnd.n374 585
R8842 gnd.n6559 gnd.n6558 585
R8843 gnd.n6558 gnd.n6557 585
R8844 gnd.n371 gnd.n370 585
R8845 gnd.n370 gnd.n369 585
R8846 gnd.n6564 gnd.n6563 585
R8847 gnd.n6565 gnd.n6564 585
R8848 gnd.n368 gnd.n367 585
R8849 gnd.n6566 gnd.n368 585
R8850 gnd.n6569 gnd.n6568 585
R8851 gnd.n6568 gnd.n6567 585
R8852 gnd.n365 gnd.n364 585
R8853 gnd.n364 gnd.n363 585
R8854 gnd.n6574 gnd.n6573 585
R8855 gnd.n6575 gnd.n6574 585
R8856 gnd.n362 gnd.n361 585
R8857 gnd.n6576 gnd.n362 585
R8858 gnd.n6579 gnd.n6578 585
R8859 gnd.n6578 gnd.n6577 585
R8860 gnd.n359 gnd.n358 585
R8861 gnd.n358 gnd.n357 585
R8862 gnd.n6584 gnd.n6583 585
R8863 gnd.n6585 gnd.n6584 585
R8864 gnd.n356 gnd.n355 585
R8865 gnd.n6586 gnd.n356 585
R8866 gnd.n6589 gnd.n6588 585
R8867 gnd.n6588 gnd.n6587 585
R8868 gnd.n353 gnd.n352 585
R8869 gnd.n352 gnd.n351 585
R8870 gnd.n6594 gnd.n6593 585
R8871 gnd.n6595 gnd.n6594 585
R8872 gnd.n350 gnd.n349 585
R8873 gnd.n6596 gnd.n350 585
R8874 gnd.n6599 gnd.n6598 585
R8875 gnd.n6598 gnd.n6597 585
R8876 gnd.n347 gnd.n346 585
R8877 gnd.n346 gnd.n345 585
R8878 gnd.n6604 gnd.n6603 585
R8879 gnd.n6605 gnd.n6604 585
R8880 gnd.n344 gnd.n343 585
R8881 gnd.n6606 gnd.n344 585
R8882 gnd.n6609 gnd.n6608 585
R8883 gnd.n6608 gnd.n6607 585
R8884 gnd.n341 gnd.n340 585
R8885 gnd.n340 gnd.n339 585
R8886 gnd.n6614 gnd.n6613 585
R8887 gnd.n6615 gnd.n6614 585
R8888 gnd.n338 gnd.n337 585
R8889 gnd.n6616 gnd.n338 585
R8890 gnd.n6619 gnd.n6618 585
R8891 gnd.n6618 gnd.n6617 585
R8892 gnd.n335 gnd.n334 585
R8893 gnd.n334 gnd.n333 585
R8894 gnd.n6624 gnd.n6623 585
R8895 gnd.n6625 gnd.n6624 585
R8896 gnd.n332 gnd.n331 585
R8897 gnd.n6626 gnd.n332 585
R8898 gnd.n6629 gnd.n6628 585
R8899 gnd.n6628 gnd.n6627 585
R8900 gnd.n329 gnd.n328 585
R8901 gnd.n328 gnd.n327 585
R8902 gnd.n6634 gnd.n6633 585
R8903 gnd.n6635 gnd.n6634 585
R8904 gnd.n326 gnd.n325 585
R8905 gnd.n6636 gnd.n326 585
R8906 gnd.n6639 gnd.n6638 585
R8907 gnd.n6638 gnd.n6637 585
R8908 gnd.n323 gnd.n322 585
R8909 gnd.n322 gnd.n321 585
R8910 gnd.n6644 gnd.n6643 585
R8911 gnd.n6645 gnd.n6644 585
R8912 gnd.n320 gnd.n319 585
R8913 gnd.n6646 gnd.n320 585
R8914 gnd.n6649 gnd.n6648 585
R8915 gnd.n6648 gnd.n6647 585
R8916 gnd.n317 gnd.n316 585
R8917 gnd.n316 gnd.n315 585
R8918 gnd.n6655 gnd.n6654 585
R8919 gnd.n6656 gnd.n6655 585
R8920 gnd.n314 gnd.n313 585
R8921 gnd.n6657 gnd.n314 585
R8922 gnd.n6660 gnd.n6659 585
R8923 gnd.n6659 gnd.n6658 585
R8924 gnd.n6661 gnd.n311 585
R8925 gnd.n311 gnd.n310 585
R8926 gnd.n186 gnd.n185 585
R8927 gnd.n6868 gnd.n185 585
R8928 gnd.n6871 gnd.n6870 585
R8929 gnd.n6870 gnd.n6869 585
R8930 gnd.n189 gnd.n188 585
R8931 gnd.n6867 gnd.n189 585
R8932 gnd.n6865 gnd.n6864 585
R8933 gnd.n6866 gnd.n6865 585
R8934 gnd.n192 gnd.n191 585
R8935 gnd.n191 gnd.n190 585
R8936 gnd.n6860 gnd.n6859 585
R8937 gnd.n6859 gnd.n6858 585
R8938 gnd.n195 gnd.n194 585
R8939 gnd.n6857 gnd.n195 585
R8940 gnd.n6855 gnd.n6854 585
R8941 gnd.n6856 gnd.n6855 585
R8942 gnd.n198 gnd.n197 585
R8943 gnd.n197 gnd.n196 585
R8944 gnd.n6850 gnd.n6849 585
R8945 gnd.n6849 gnd.n6848 585
R8946 gnd.n201 gnd.n200 585
R8947 gnd.n6847 gnd.n201 585
R8948 gnd.n6845 gnd.n6844 585
R8949 gnd.n6846 gnd.n6845 585
R8950 gnd.n204 gnd.n203 585
R8951 gnd.n203 gnd.n202 585
R8952 gnd.n6840 gnd.n6839 585
R8953 gnd.n6839 gnd.n6838 585
R8954 gnd.n207 gnd.n206 585
R8955 gnd.n6837 gnd.n207 585
R8956 gnd.n6835 gnd.n6834 585
R8957 gnd.n6836 gnd.n6835 585
R8958 gnd.n210 gnd.n209 585
R8959 gnd.n209 gnd.n208 585
R8960 gnd.n6830 gnd.n6829 585
R8961 gnd.n6829 gnd.n6828 585
R8962 gnd.n213 gnd.n212 585
R8963 gnd.n6827 gnd.n213 585
R8964 gnd.n6825 gnd.n6824 585
R8965 gnd.n6826 gnd.n6825 585
R8966 gnd.n216 gnd.n215 585
R8967 gnd.n215 gnd.n214 585
R8968 gnd.n6820 gnd.n6819 585
R8969 gnd.n6819 gnd.n6818 585
R8970 gnd.n219 gnd.n218 585
R8971 gnd.n6817 gnd.n219 585
R8972 gnd.n6815 gnd.n6814 585
R8973 gnd.n6816 gnd.n6815 585
R8974 gnd.n222 gnd.n221 585
R8975 gnd.n221 gnd.n220 585
R8976 gnd.n6810 gnd.n6809 585
R8977 gnd.n6809 gnd.n6808 585
R8978 gnd.n225 gnd.n224 585
R8979 gnd.n6807 gnd.n225 585
R8980 gnd.n6805 gnd.n6804 585
R8981 gnd.n6806 gnd.n6805 585
R8982 gnd.n228 gnd.n227 585
R8983 gnd.n227 gnd.n226 585
R8984 gnd.n6800 gnd.n6799 585
R8985 gnd.n6799 gnd.n6798 585
R8986 gnd.n231 gnd.n230 585
R8987 gnd.n6797 gnd.n231 585
R8988 gnd.n6795 gnd.n6794 585
R8989 gnd.n6796 gnd.n6795 585
R8990 gnd.n234 gnd.n233 585
R8991 gnd.n233 gnd.n232 585
R8992 gnd.n6790 gnd.n6789 585
R8993 gnd.n6789 gnd.n6788 585
R8994 gnd.n237 gnd.n236 585
R8995 gnd.n6787 gnd.n237 585
R8996 gnd.n6785 gnd.n6784 585
R8997 gnd.n6786 gnd.n6785 585
R8998 gnd.n240 gnd.n239 585
R8999 gnd.n239 gnd.n238 585
R9000 gnd.n6780 gnd.n6779 585
R9001 gnd.n6779 gnd.n6778 585
R9002 gnd.n243 gnd.n242 585
R9003 gnd.n6777 gnd.n243 585
R9004 gnd.n6775 gnd.n6774 585
R9005 gnd.n6776 gnd.n6775 585
R9006 gnd.n246 gnd.n245 585
R9007 gnd.n245 gnd.n244 585
R9008 gnd.n6770 gnd.n6769 585
R9009 gnd.n6769 gnd.n6768 585
R9010 gnd.n249 gnd.n248 585
R9011 gnd.n6767 gnd.n249 585
R9012 gnd.n6765 gnd.n6764 585
R9013 gnd.n6766 gnd.n6765 585
R9014 gnd.n252 gnd.n251 585
R9015 gnd.n251 gnd.n250 585
R9016 gnd.n6760 gnd.n6759 585
R9017 gnd.n6759 gnd.n6758 585
R9018 gnd.n255 gnd.n254 585
R9019 gnd.n6757 gnd.n255 585
R9020 gnd.n6755 gnd.n6754 585
R9021 gnd.n6756 gnd.n6755 585
R9022 gnd.n258 gnd.n257 585
R9023 gnd.n257 gnd.n256 585
R9024 gnd.n6750 gnd.n6749 585
R9025 gnd.n6749 gnd.n6748 585
R9026 gnd.n261 gnd.n260 585
R9027 gnd.n6747 gnd.n261 585
R9028 gnd.n6745 gnd.n6744 585
R9029 gnd.n6746 gnd.n6745 585
R9030 gnd.n264 gnd.n263 585
R9031 gnd.n263 gnd.n262 585
R9032 gnd.n6740 gnd.n6739 585
R9033 gnd.n6739 gnd.n6738 585
R9034 gnd.n267 gnd.n266 585
R9035 gnd.n6737 gnd.n267 585
R9036 gnd.n6735 gnd.n6734 585
R9037 gnd.n6736 gnd.n6735 585
R9038 gnd.n270 gnd.n269 585
R9039 gnd.n269 gnd.n268 585
R9040 gnd.n6730 gnd.n6729 585
R9041 gnd.n6729 gnd.n6728 585
R9042 gnd.n273 gnd.n272 585
R9043 gnd.n6727 gnd.n273 585
R9044 gnd.n6725 gnd.n6724 585
R9045 gnd.n6726 gnd.n6725 585
R9046 gnd.n276 gnd.n275 585
R9047 gnd.n275 gnd.n274 585
R9048 gnd.n6720 gnd.n6719 585
R9049 gnd.n6719 gnd.n6718 585
R9050 gnd.n279 gnd.n278 585
R9051 gnd.n6717 gnd.n279 585
R9052 gnd.n6715 gnd.n6714 585
R9053 gnd.n6716 gnd.n6715 585
R9054 gnd.n282 gnd.n281 585
R9055 gnd.n281 gnd.n280 585
R9056 gnd.n6710 gnd.n6709 585
R9057 gnd.n6709 gnd.n6708 585
R9058 gnd.n285 gnd.n284 585
R9059 gnd.n6707 gnd.n285 585
R9060 gnd.n6705 gnd.n6704 585
R9061 gnd.n6706 gnd.n6705 585
R9062 gnd.n288 gnd.n287 585
R9063 gnd.n287 gnd.n286 585
R9064 gnd.n6700 gnd.n6699 585
R9065 gnd.n6699 gnd.n6698 585
R9066 gnd.n291 gnd.n290 585
R9067 gnd.n6697 gnd.n291 585
R9068 gnd.n6695 gnd.n6694 585
R9069 gnd.n6696 gnd.n6695 585
R9070 gnd.n294 gnd.n293 585
R9071 gnd.n293 gnd.n292 585
R9072 gnd.n6690 gnd.n6689 585
R9073 gnd.n6689 gnd.n6688 585
R9074 gnd.n297 gnd.n296 585
R9075 gnd.n6687 gnd.n297 585
R9076 gnd.n6685 gnd.n6684 585
R9077 gnd.n6686 gnd.n6685 585
R9078 gnd.n300 gnd.n299 585
R9079 gnd.n299 gnd.n298 585
R9080 gnd.n6680 gnd.n6679 585
R9081 gnd.n6679 gnd.n6678 585
R9082 gnd.n303 gnd.n302 585
R9083 gnd.n6677 gnd.n303 585
R9084 gnd.n6675 gnd.n6674 585
R9085 gnd.n6676 gnd.n6675 585
R9086 gnd.n306 gnd.n305 585
R9087 gnd.n305 gnd.n304 585
R9088 gnd.n6670 gnd.n6669 585
R9089 gnd.n6669 gnd.n6668 585
R9090 gnd.n309 gnd.n308 585
R9091 gnd.n6667 gnd.n309 585
R9092 gnd.n6665 gnd.n6664 585
R9093 gnd.n6666 gnd.n6665 585
R9094 gnd.n5984 gnd.n5983 585
R9095 gnd.n5985 gnd.n5984 585
R9096 gnd.n849 gnd.n848 585
R9097 gnd.n5978 gnd.n849 585
R9098 gnd.n5993 gnd.n5992 585
R9099 gnd.n5992 gnd.n5991 585
R9100 gnd.n5994 gnd.n844 585
R9101 gnd.n4202 gnd.n844 585
R9102 gnd.n5996 gnd.n5995 585
R9103 gnd.n5997 gnd.n5996 585
R9104 gnd.n829 gnd.n828 585
R9105 gnd.n4196 gnd.n829 585
R9106 gnd.n6005 gnd.n6004 585
R9107 gnd.n6004 gnd.n6003 585
R9108 gnd.n6006 gnd.n824 585
R9109 gnd.n4191 gnd.n824 585
R9110 gnd.n6008 gnd.n6007 585
R9111 gnd.n6009 gnd.n6008 585
R9112 gnd.n808 gnd.n807 585
R9113 gnd.n4186 gnd.n808 585
R9114 gnd.n6017 gnd.n6016 585
R9115 gnd.n6016 gnd.n6015 585
R9116 gnd.n6018 gnd.n803 585
R9117 gnd.n4219 gnd.n803 585
R9118 gnd.n6020 gnd.n6019 585
R9119 gnd.n6021 gnd.n6020 585
R9120 gnd.n789 gnd.n788 585
R9121 gnd.n4179 gnd.n789 585
R9122 gnd.n6029 gnd.n6028 585
R9123 gnd.n6028 gnd.n6027 585
R9124 gnd.n6030 gnd.n784 585
R9125 gnd.n4171 gnd.n784 585
R9126 gnd.n6032 gnd.n6031 585
R9127 gnd.n6033 gnd.n6032 585
R9128 gnd.n771 gnd.n770 585
R9129 gnd.n4145 gnd.n771 585
R9130 gnd.n6042 gnd.n6041 585
R9131 gnd.n6041 gnd.n6040 585
R9132 gnd.n6043 gnd.n766 585
R9133 gnd.n4153 gnd.n766 585
R9134 gnd.n6045 gnd.n6044 585
R9135 gnd.n6046 gnd.n6045 585
R9136 gnd.n755 gnd.n754 585
R9137 gnd.n4134 gnd.n755 585
R9138 gnd.n6055 gnd.n6054 585
R9139 gnd.n6054 gnd.n6053 585
R9140 gnd.n6056 gnd.n749 585
R9141 gnd.n4126 gnd.n749 585
R9142 gnd.n6058 gnd.n6057 585
R9143 gnd.n6059 gnd.n6058 585
R9144 gnd.n750 gnd.n748 585
R9145 gnd.n4108 gnd.n748 585
R9146 gnd.n4083 gnd.n737 585
R9147 gnd.n6066 gnd.n737 585
R9148 gnd.n4085 gnd.n4084 585
R9149 gnd.n4084 gnd.n733 585
R9150 gnd.n4086 gnd.n2172 585
R9151 gnd.n4099 gnd.n2172 585
R9152 gnd.n4087 gnd.n2182 585
R9153 gnd.n2182 gnd.n2180 585
R9154 gnd.n4089 gnd.n4088 585
R9155 gnd.n4090 gnd.n4089 585
R9156 gnd.n2183 gnd.n2181 585
R9157 gnd.n4072 gnd.n2181 585
R9158 gnd.n4045 gnd.n4044 585
R9159 gnd.n4044 gnd.n2190 585
R9160 gnd.n4046 gnd.n2198 585
R9161 gnd.n4060 gnd.n2198 585
R9162 gnd.n4047 gnd.n2208 585
R9163 gnd.n2208 gnd.n2196 585
R9164 gnd.n4049 gnd.n4048 585
R9165 gnd.n4050 gnd.n4049 585
R9166 gnd.n2209 gnd.n2207 585
R9167 gnd.n4035 gnd.n2207 585
R9168 gnd.n4010 gnd.n4009 585
R9169 gnd.n4009 gnd.n2215 585
R9170 gnd.n4011 gnd.n2223 585
R9171 gnd.n4025 gnd.n2223 585
R9172 gnd.n4012 gnd.n2233 585
R9173 gnd.n2233 gnd.n2221 585
R9174 gnd.n4014 gnd.n4013 585
R9175 gnd.n4015 gnd.n4014 585
R9176 gnd.n2234 gnd.n2232 585
R9177 gnd.n3780 gnd.n2232 585
R9178 gnd.n3999 gnd.n3998 585
R9179 gnd.n3998 gnd.n3997 585
R9180 gnd.n3727 gnd.n2240 585
R9181 gnd.n3730 gnd.n3728 585
R9182 gnd.n3733 gnd.n3732 585
R9183 gnd.n3724 gnd.n3723 585
R9184 gnd.n3738 gnd.n3737 585
R9185 gnd.n3740 gnd.n3722 585
R9186 gnd.n3743 gnd.n3742 585
R9187 gnd.n3720 gnd.n3719 585
R9188 gnd.n3748 gnd.n3747 585
R9189 gnd.n3750 gnd.n3718 585
R9190 gnd.n3753 gnd.n3752 585
R9191 gnd.n3716 gnd.n3715 585
R9192 gnd.n3758 gnd.n3757 585
R9193 gnd.n3760 gnd.n3714 585
R9194 gnd.n3763 gnd.n3762 585
R9195 gnd.n3712 gnd.n3711 585
R9196 gnd.n3768 gnd.n3767 585
R9197 gnd.n3770 gnd.n3710 585
R9198 gnd.n3772 gnd.n3771 585
R9199 gnd.n3771 gnd.n3703 585
R9200 gnd.n5905 gnd.n5904 585
R9201 gnd.n5906 gnd.n964 585
R9202 gnd.n5907 gnd.n959 585
R9203 gnd.n977 gnd.n948 585
R9204 gnd.n5914 gnd.n947 585
R9205 gnd.n5915 gnd.n946 585
R9206 gnd.n974 gnd.n940 585
R9207 gnd.n5922 gnd.n939 585
R9208 gnd.n5923 gnd.n938 585
R9209 gnd.n972 gnd.n930 585
R9210 gnd.n5930 gnd.n929 585
R9211 gnd.n5931 gnd.n928 585
R9212 gnd.n969 gnd.n922 585
R9213 gnd.n5938 gnd.n921 585
R9214 gnd.n5939 gnd.n920 585
R9215 gnd.n967 gnd.n912 585
R9216 gnd.n5946 gnd.n911 585
R9217 gnd.n5947 gnd.n910 585
R9218 gnd.n909 gnd.n863 585
R9219 gnd.n5902 gnd.n863 585
R9220 gnd.n869 gnd.n861 585
R9221 gnd.n5985 gnd.n861 585
R9222 gnd.n5977 gnd.n5976 585
R9223 gnd.n5978 gnd.n5977 585
R9224 gnd.n868 gnd.n852 585
R9225 gnd.n5991 gnd.n852 585
R9226 gnd.n4205 gnd.n4203 585
R9227 gnd.n4203 gnd.n4202 585
R9228 gnd.n4206 gnd.n842 585
R9229 gnd.n5997 gnd.n842 585
R9230 gnd.n4207 gnd.n2142 585
R9231 gnd.n4196 gnd.n2142 585
R9232 gnd.n2140 gnd.n831 585
R9233 gnd.n6003 gnd.n831 585
R9234 gnd.n4211 gnd.n2139 585
R9235 gnd.n4191 gnd.n2139 585
R9236 gnd.n4212 gnd.n822 585
R9237 gnd.n6009 gnd.n822 585
R9238 gnd.n4213 gnd.n2138 585
R9239 gnd.n4186 gnd.n2138 585
R9240 gnd.n2135 gnd.n811 585
R9241 gnd.n6015 gnd.n811 585
R9242 gnd.n4218 gnd.n4217 585
R9243 gnd.n4219 gnd.n4218 585
R9244 gnd.n2134 gnd.n802 585
R9245 gnd.n6021 gnd.n802 585
R9246 gnd.n4178 gnd.n4177 585
R9247 gnd.n4179 gnd.n4178 585
R9248 gnd.n2145 gnd.n791 585
R9249 gnd.n6027 gnd.n791 585
R9250 gnd.n4173 gnd.n4172 585
R9251 gnd.n4172 gnd.n4171 585
R9252 gnd.n2147 gnd.n782 585
R9253 gnd.n6033 gnd.n782 585
R9254 gnd.n4147 gnd.n4146 585
R9255 gnd.n4146 gnd.n4145 585
R9256 gnd.n2157 gnd.n774 585
R9257 gnd.n6040 gnd.n774 585
R9258 gnd.n4152 gnd.n4151 585
R9259 gnd.n4153 gnd.n4152 585
R9260 gnd.n2156 gnd.n765 585
R9261 gnd.n6046 gnd.n765 585
R9262 gnd.n4133 gnd.n4132 585
R9263 gnd.n4134 gnd.n4133 585
R9264 gnd.n2161 gnd.n757 585
R9265 gnd.n6053 gnd.n757 585
R9266 gnd.n4128 gnd.n4127 585
R9267 gnd.n4127 gnd.n4126 585
R9268 gnd.n2163 gnd.n746 585
R9269 gnd.n6059 gnd.n746 585
R9270 gnd.n4107 gnd.n4106 585
R9271 gnd.n4108 gnd.n4107 585
R9272 gnd.n2166 gnd.n735 585
R9273 gnd.n6066 gnd.n735 585
R9274 gnd.n4102 gnd.n4101 585
R9275 gnd.n4101 gnd.n733 585
R9276 gnd.n4100 gnd.n2168 585
R9277 gnd.n4100 gnd.n4099 585
R9278 gnd.n4068 gnd.n2169 585
R9279 gnd.n2180 gnd.n2169 585
R9280 gnd.n4069 gnd.n2179 585
R9281 gnd.n4090 gnd.n2179 585
R9282 gnd.n4071 gnd.n4070 585
R9283 gnd.n4072 gnd.n4071 585
R9284 gnd.n2192 gnd.n2191 585
R9285 gnd.n2191 gnd.n2190 585
R9286 gnd.n4062 gnd.n4061 585
R9287 gnd.n4061 gnd.n4060 585
R9288 gnd.n2195 gnd.n2194 585
R9289 gnd.n2196 gnd.n2195 585
R9290 gnd.n4032 gnd.n2206 585
R9291 gnd.n4050 gnd.n2206 585
R9292 gnd.n4034 gnd.n4033 585
R9293 gnd.n4035 gnd.n4034 585
R9294 gnd.n2217 gnd.n2216 585
R9295 gnd.n2216 gnd.n2215 585
R9296 gnd.n4027 gnd.n4026 585
R9297 gnd.n4026 gnd.n4025 585
R9298 gnd.n2220 gnd.n2219 585
R9299 gnd.n2221 gnd.n2220 585
R9300 gnd.n3777 gnd.n2231 585
R9301 gnd.n4015 gnd.n2231 585
R9302 gnd.n3779 gnd.n3778 585
R9303 gnd.n3780 gnd.n3779 585
R9304 gnd.n3706 gnd.n3705 585
R9305 gnd.n3997 gnd.n3705 585
R9306 gnd.n3610 gnd.n3609 585
R9307 gnd.n3611 gnd.n3610 585
R9308 gnd.n2317 gnd.n2316 585
R9309 gnd.n2323 gnd.n2316 585
R9310 gnd.n3585 gnd.n2335 585
R9311 gnd.n2335 gnd.n2322 585
R9312 gnd.n3587 gnd.n3586 585
R9313 gnd.n3588 gnd.n3587 585
R9314 gnd.n2336 gnd.n2334 585
R9315 gnd.n2334 gnd.n2330 585
R9316 gnd.n3319 gnd.n3318 585
R9317 gnd.n3318 gnd.n3317 585
R9318 gnd.n2341 gnd.n2340 585
R9319 gnd.n3288 gnd.n2341 585
R9320 gnd.n3308 gnd.n3307 585
R9321 gnd.n3307 gnd.n3306 585
R9322 gnd.n2348 gnd.n2347 585
R9323 gnd.n3294 gnd.n2348 585
R9324 gnd.n3264 gnd.n2368 585
R9325 gnd.n2368 gnd.n2367 585
R9326 gnd.n3266 gnd.n3265 585
R9327 gnd.n3267 gnd.n3266 585
R9328 gnd.n2369 gnd.n2366 585
R9329 gnd.n2377 gnd.n2366 585
R9330 gnd.n3242 gnd.n2389 585
R9331 gnd.n2389 gnd.n2376 585
R9332 gnd.n3244 gnd.n3243 585
R9333 gnd.n3245 gnd.n3244 585
R9334 gnd.n2390 gnd.n2388 585
R9335 gnd.n2388 gnd.n2384 585
R9336 gnd.n3230 gnd.n3229 585
R9337 gnd.n3229 gnd.n3228 585
R9338 gnd.n2395 gnd.n2394 585
R9339 gnd.n2405 gnd.n2395 585
R9340 gnd.n3219 gnd.n3218 585
R9341 gnd.n3218 gnd.n3217 585
R9342 gnd.n2402 gnd.n2401 585
R9343 gnd.n3205 gnd.n2402 585
R9344 gnd.n3179 gnd.n2423 585
R9345 gnd.n2423 gnd.n2412 585
R9346 gnd.n3181 gnd.n3180 585
R9347 gnd.n3182 gnd.n3181 585
R9348 gnd.n2424 gnd.n2422 585
R9349 gnd.n2432 gnd.n2422 585
R9350 gnd.n3157 gnd.n2444 585
R9351 gnd.n2444 gnd.n2431 585
R9352 gnd.n3159 gnd.n3158 585
R9353 gnd.n3160 gnd.n3159 585
R9354 gnd.n2445 gnd.n2443 585
R9355 gnd.n2443 gnd.n2439 585
R9356 gnd.n3145 gnd.n3144 585
R9357 gnd.n3144 gnd.n3143 585
R9358 gnd.n2450 gnd.n2449 585
R9359 gnd.n2459 gnd.n2450 585
R9360 gnd.n3134 gnd.n3133 585
R9361 gnd.n3133 gnd.n3132 585
R9362 gnd.n2457 gnd.n2456 585
R9363 gnd.n3120 gnd.n2457 585
R9364 gnd.n2558 gnd.n2557 585
R9365 gnd.n2558 gnd.n2466 585
R9366 gnd.n3077 gnd.n3076 585
R9367 gnd.n3076 gnd.n3075 585
R9368 gnd.n3078 gnd.n2552 585
R9369 gnd.n2563 gnd.n2552 585
R9370 gnd.n3080 gnd.n3079 585
R9371 gnd.n3081 gnd.n3080 585
R9372 gnd.n2553 gnd.n2551 585
R9373 gnd.n2576 gnd.n2551 585
R9374 gnd.n2536 gnd.n2535 585
R9375 gnd.n2539 gnd.n2536 585
R9376 gnd.n3091 gnd.n3090 585
R9377 gnd.n3090 gnd.n3089 585
R9378 gnd.n3092 gnd.n2530 585
R9379 gnd.n3051 gnd.n2530 585
R9380 gnd.n3094 gnd.n3093 585
R9381 gnd.n3095 gnd.n3094 585
R9382 gnd.n2531 gnd.n2529 585
R9383 gnd.n2590 gnd.n2529 585
R9384 gnd.n3043 gnd.n3042 585
R9385 gnd.n3042 gnd.n3041 585
R9386 gnd.n2587 gnd.n2586 585
R9387 gnd.n3025 gnd.n2587 585
R9388 gnd.n3012 gnd.n2606 585
R9389 gnd.n2606 gnd.n2605 585
R9390 gnd.n3014 gnd.n3013 585
R9391 gnd.n3015 gnd.n3014 585
R9392 gnd.n2607 gnd.n2604 585
R9393 gnd.n2613 gnd.n2604 585
R9394 gnd.n2993 gnd.n2992 585
R9395 gnd.n2994 gnd.n2993 585
R9396 gnd.n2624 gnd.n2623 585
R9397 gnd.n2623 gnd.n2619 585
R9398 gnd.n2983 gnd.n2982 585
R9399 gnd.n2984 gnd.n2983 585
R9400 gnd.n2634 gnd.n2633 585
R9401 gnd.n2639 gnd.n2633 585
R9402 gnd.n2961 gnd.n2652 585
R9403 gnd.n2652 gnd.n2638 585
R9404 gnd.n2963 gnd.n2962 585
R9405 gnd.n2964 gnd.n2963 585
R9406 gnd.n2653 gnd.n2651 585
R9407 gnd.n2651 gnd.n2647 585
R9408 gnd.n2952 gnd.n2951 585
R9409 gnd.n2953 gnd.n2952 585
R9410 gnd.n2660 gnd.n2659 585
R9411 gnd.n2664 gnd.n2659 585
R9412 gnd.n2929 gnd.n2681 585
R9413 gnd.n2681 gnd.n2663 585
R9414 gnd.n2931 gnd.n2930 585
R9415 gnd.n2932 gnd.n2931 585
R9416 gnd.n2682 gnd.n2680 585
R9417 gnd.n2680 gnd.n2671 585
R9418 gnd.n2924 gnd.n2923 585
R9419 gnd.n2923 gnd.n2922 585
R9420 gnd.n2729 gnd.n2728 585
R9421 gnd.n2730 gnd.n2729 585
R9422 gnd.n2883 gnd.n2882 585
R9423 gnd.n2884 gnd.n2883 585
R9424 gnd.n2739 gnd.n2738 585
R9425 gnd.n2738 gnd.n2737 585
R9426 gnd.n2878 gnd.n2877 585
R9427 gnd.n2877 gnd.n2876 585
R9428 gnd.n2742 gnd.n2741 585
R9429 gnd.n2743 gnd.n2742 585
R9430 gnd.n2867 gnd.n2866 585
R9431 gnd.n2868 gnd.n2867 585
R9432 gnd.n2750 gnd.n2749 585
R9433 gnd.n2859 gnd.n2749 585
R9434 gnd.n2862 gnd.n2861 585
R9435 gnd.n2861 gnd.n2860 585
R9436 gnd.n2753 gnd.n2752 585
R9437 gnd.n2754 gnd.n2753 585
R9438 gnd.n2848 gnd.n2847 585
R9439 gnd.n2846 gnd.n2772 585
R9440 gnd.n2845 gnd.n2771 585
R9441 gnd.n2850 gnd.n2771 585
R9442 gnd.n2844 gnd.n2843 585
R9443 gnd.n2842 gnd.n2841 585
R9444 gnd.n2840 gnd.n2839 585
R9445 gnd.n2838 gnd.n2837 585
R9446 gnd.n2836 gnd.n2835 585
R9447 gnd.n2834 gnd.n2833 585
R9448 gnd.n2832 gnd.n2831 585
R9449 gnd.n2830 gnd.n2829 585
R9450 gnd.n2828 gnd.n2827 585
R9451 gnd.n2826 gnd.n2825 585
R9452 gnd.n2824 gnd.n2823 585
R9453 gnd.n2822 gnd.n2821 585
R9454 gnd.n2820 gnd.n2819 585
R9455 gnd.n2818 gnd.n2817 585
R9456 gnd.n2816 gnd.n2815 585
R9457 gnd.n2814 gnd.n2813 585
R9458 gnd.n2812 gnd.n2811 585
R9459 gnd.n2810 gnd.n2809 585
R9460 gnd.n2808 gnd.n2807 585
R9461 gnd.n2806 gnd.n2805 585
R9462 gnd.n2804 gnd.n2803 585
R9463 gnd.n2802 gnd.n2801 585
R9464 gnd.n2759 gnd.n2758 585
R9465 gnd.n2853 gnd.n2852 585
R9466 gnd.n3614 gnd.n3613 585
R9467 gnd.n3616 gnd.n3615 585
R9468 gnd.n3618 gnd.n3617 585
R9469 gnd.n3620 gnd.n3619 585
R9470 gnd.n3622 gnd.n3621 585
R9471 gnd.n3624 gnd.n3623 585
R9472 gnd.n3626 gnd.n3625 585
R9473 gnd.n3628 gnd.n3627 585
R9474 gnd.n3630 gnd.n3629 585
R9475 gnd.n3632 gnd.n3631 585
R9476 gnd.n3634 gnd.n3633 585
R9477 gnd.n3636 gnd.n3635 585
R9478 gnd.n3638 gnd.n3637 585
R9479 gnd.n3640 gnd.n3639 585
R9480 gnd.n3642 gnd.n3641 585
R9481 gnd.n3644 gnd.n3643 585
R9482 gnd.n3646 gnd.n3645 585
R9483 gnd.n3648 gnd.n3647 585
R9484 gnd.n3650 gnd.n3649 585
R9485 gnd.n3652 gnd.n3651 585
R9486 gnd.n3654 gnd.n3653 585
R9487 gnd.n3656 gnd.n3655 585
R9488 gnd.n3658 gnd.n3657 585
R9489 gnd.n3660 gnd.n3659 585
R9490 gnd.n3662 gnd.n3661 585
R9491 gnd.n3663 gnd.n2284 585
R9492 gnd.n3664 gnd.n2242 585
R9493 gnd.n3702 gnd.n2242 585
R9494 gnd.n3612 gnd.n2314 585
R9495 gnd.n3612 gnd.n3611 585
R9496 gnd.n3281 gnd.n2313 585
R9497 gnd.n2323 gnd.n2313 585
R9498 gnd.n3283 gnd.n3282 585
R9499 gnd.n3282 gnd.n2322 585
R9500 gnd.n3284 gnd.n2332 585
R9501 gnd.n3588 gnd.n2332 585
R9502 gnd.n3286 gnd.n3285 585
R9503 gnd.n3285 gnd.n2330 585
R9504 gnd.n3287 gnd.n2343 585
R9505 gnd.n3317 gnd.n2343 585
R9506 gnd.n3290 gnd.n3289 585
R9507 gnd.n3289 gnd.n3288 585
R9508 gnd.n3291 gnd.n2350 585
R9509 gnd.n3306 gnd.n2350 585
R9510 gnd.n3293 gnd.n3292 585
R9511 gnd.n3294 gnd.n3293 585
R9512 gnd.n2360 gnd.n2359 585
R9513 gnd.n2367 gnd.n2359 585
R9514 gnd.n3269 gnd.n3268 585
R9515 gnd.n3268 gnd.n3267 585
R9516 gnd.n2363 gnd.n2362 585
R9517 gnd.n2377 gnd.n2363 585
R9518 gnd.n3195 gnd.n3194 585
R9519 gnd.n3194 gnd.n2376 585
R9520 gnd.n3196 gnd.n2386 585
R9521 gnd.n3245 gnd.n2386 585
R9522 gnd.n3198 gnd.n3197 585
R9523 gnd.n3197 gnd.n2384 585
R9524 gnd.n3199 gnd.n2397 585
R9525 gnd.n3228 gnd.n2397 585
R9526 gnd.n3201 gnd.n3200 585
R9527 gnd.n3200 gnd.n2405 585
R9528 gnd.n3202 gnd.n2404 585
R9529 gnd.n3217 gnd.n2404 585
R9530 gnd.n3204 gnd.n3203 585
R9531 gnd.n3205 gnd.n3204 585
R9532 gnd.n2416 gnd.n2415 585
R9533 gnd.n2415 gnd.n2412 585
R9534 gnd.n3184 gnd.n3183 585
R9535 gnd.n3183 gnd.n3182 585
R9536 gnd.n2419 gnd.n2418 585
R9537 gnd.n2432 gnd.n2419 585
R9538 gnd.n3108 gnd.n3107 585
R9539 gnd.n3107 gnd.n2431 585
R9540 gnd.n3109 gnd.n2441 585
R9541 gnd.n3160 gnd.n2441 585
R9542 gnd.n3111 gnd.n3110 585
R9543 gnd.n3110 gnd.n2439 585
R9544 gnd.n3112 gnd.n2452 585
R9545 gnd.n3143 gnd.n2452 585
R9546 gnd.n3114 gnd.n3113 585
R9547 gnd.n3113 gnd.n2459 585
R9548 gnd.n3115 gnd.n2458 585
R9549 gnd.n3132 gnd.n2458 585
R9550 gnd.n3117 gnd.n3116 585
R9551 gnd.n3120 gnd.n3117 585
R9552 gnd.n2469 gnd.n2468 585
R9553 gnd.n2468 gnd.n2466 585
R9554 gnd.n2560 gnd.n2559 585
R9555 gnd.n3075 gnd.n2559 585
R9556 gnd.n2562 gnd.n2561 585
R9557 gnd.n2563 gnd.n2562 585
R9558 gnd.n2573 gnd.n2549 585
R9559 gnd.n3081 gnd.n2549 585
R9560 gnd.n2575 gnd.n2574 585
R9561 gnd.n2576 gnd.n2575 585
R9562 gnd.n2572 gnd.n2571 585
R9563 gnd.n2572 gnd.n2539 585
R9564 gnd.n2570 gnd.n2537 585
R9565 gnd.n3089 gnd.n2537 585
R9566 gnd.n2526 gnd.n2524 585
R9567 gnd.n3051 gnd.n2526 585
R9568 gnd.n3097 gnd.n3096 585
R9569 gnd.n3096 gnd.n3095 585
R9570 gnd.n2525 gnd.n2523 585
R9571 gnd.n2590 gnd.n2525 585
R9572 gnd.n3022 gnd.n2589 585
R9573 gnd.n3041 gnd.n2589 585
R9574 gnd.n3024 gnd.n3023 585
R9575 gnd.n3025 gnd.n3024 585
R9576 gnd.n2599 gnd.n2598 585
R9577 gnd.n2605 gnd.n2598 585
R9578 gnd.n3017 gnd.n3016 585
R9579 gnd.n3016 gnd.n3015 585
R9580 gnd.n2602 gnd.n2601 585
R9581 gnd.n2613 gnd.n2602 585
R9582 gnd.n2902 gnd.n2621 585
R9583 gnd.n2994 gnd.n2621 585
R9584 gnd.n2904 gnd.n2903 585
R9585 gnd.n2903 gnd.n2619 585
R9586 gnd.n2905 gnd.n2632 585
R9587 gnd.n2984 gnd.n2632 585
R9588 gnd.n2907 gnd.n2906 585
R9589 gnd.n2907 gnd.n2639 585
R9590 gnd.n2909 gnd.n2908 585
R9591 gnd.n2908 gnd.n2638 585
R9592 gnd.n2910 gnd.n2649 585
R9593 gnd.n2964 gnd.n2649 585
R9594 gnd.n2912 gnd.n2911 585
R9595 gnd.n2911 gnd.n2647 585
R9596 gnd.n2913 gnd.n2658 585
R9597 gnd.n2953 gnd.n2658 585
R9598 gnd.n2915 gnd.n2914 585
R9599 gnd.n2915 gnd.n2664 585
R9600 gnd.n2917 gnd.n2916 585
R9601 gnd.n2916 gnd.n2663 585
R9602 gnd.n2918 gnd.n2679 585
R9603 gnd.n2932 gnd.n2679 585
R9604 gnd.n2919 gnd.n2732 585
R9605 gnd.n2732 gnd.n2671 585
R9606 gnd.n2921 gnd.n2920 585
R9607 gnd.n2922 gnd.n2921 585
R9608 gnd.n2733 gnd.n2731 585
R9609 gnd.n2731 gnd.n2730 585
R9610 gnd.n2886 gnd.n2885 585
R9611 gnd.n2885 gnd.n2884 585
R9612 gnd.n2736 gnd.n2735 585
R9613 gnd.n2737 gnd.n2736 585
R9614 gnd.n2875 gnd.n2874 585
R9615 gnd.n2876 gnd.n2875 585
R9616 gnd.n2745 gnd.n2744 585
R9617 gnd.n2744 gnd.n2743 585
R9618 gnd.n2870 gnd.n2869 585
R9619 gnd.n2869 gnd.n2868 585
R9620 gnd.n2748 gnd.n2747 585
R9621 gnd.n2859 gnd.n2748 585
R9622 gnd.n2858 gnd.n2857 585
R9623 gnd.n2860 gnd.n2858 585
R9624 gnd.n2756 gnd.n2755 585
R9625 gnd.n2755 gnd.n2754 585
R9626 gnd.n7246 gnd.n7245 585
R9627 gnd.n7247 gnd.n7246 585
R9628 gnd.n158 gnd.n157 585
R9629 gnd.n167 gnd.n158 585
R9630 gnd.n7255 gnd.n7254 585
R9631 gnd.n7254 gnd.n7253 585
R9632 gnd.n7256 gnd.n153 585
R9633 gnd.n153 gnd.n152 585
R9634 gnd.n7258 gnd.n7257 585
R9635 gnd.n7259 gnd.n7258 585
R9636 gnd.n139 gnd.n138 585
R9637 gnd.n142 gnd.n139 585
R9638 gnd.n7267 gnd.n7266 585
R9639 gnd.n7266 gnd.n7265 585
R9640 gnd.n7268 gnd.n134 585
R9641 gnd.n134 gnd.n133 585
R9642 gnd.n7270 gnd.n7269 585
R9643 gnd.n7271 gnd.n7270 585
R9644 gnd.n119 gnd.n118 585
R9645 gnd.n130 gnd.n119 585
R9646 gnd.n7279 gnd.n7278 585
R9647 gnd.n7278 gnd.n7277 585
R9648 gnd.n7280 gnd.n114 585
R9649 gnd.n120 gnd.n114 585
R9650 gnd.n7282 gnd.n7281 585
R9651 gnd.n7283 gnd.n7282 585
R9652 gnd.n101 gnd.n100 585
R9653 gnd.n111 gnd.n101 585
R9654 gnd.n7291 gnd.n7290 585
R9655 gnd.n7290 gnd.n7289 585
R9656 gnd.n7292 gnd.n95 585
R9657 gnd.n7216 gnd.n95 585
R9658 gnd.n7294 gnd.n7293 585
R9659 gnd.n7295 gnd.n7294 585
R9660 gnd.n96 gnd.n94 585
R9661 gnd.n6891 gnd.n94 585
R9662 gnd.n6886 gnd.n6885 585
R9663 gnd.n6885 gnd.n6884 585
R9664 gnd.n180 gnd.n76 585
R9665 gnd.n7303 gnd.n76 585
R9666 gnd.n5394 gnd.n5393 585
R9667 gnd.n5395 gnd.n5394 585
R9668 gnd.n1606 gnd.n1605 585
R9669 gnd.n1605 gnd.n1603 585
R9670 gnd.n5385 gnd.n5384 585
R9671 gnd.n5386 gnd.n5385 585
R9672 gnd.n1584 gnd.n1583 585
R9673 gnd.n5404 gnd.n1584 585
R9674 gnd.n5411 gnd.n5410 585
R9675 gnd.n5410 gnd.n5409 585
R9676 gnd.n5412 gnd.n1579 585
R9677 gnd.n5377 gnd.n1579 585
R9678 gnd.n5414 gnd.n5413 585
R9679 gnd.n5415 gnd.n5414 585
R9680 gnd.n1567 gnd.n1566 585
R9681 gnd.n5365 gnd.n1567 585
R9682 gnd.n5423 gnd.n5422 585
R9683 gnd.n5422 gnd.n5421 585
R9684 gnd.n5424 gnd.n1562 585
R9685 gnd.n5358 gnd.n1562 585
R9686 gnd.n5426 gnd.n5425 585
R9687 gnd.n5427 gnd.n5426 585
R9688 gnd.n1547 gnd.n1546 585
R9689 gnd.n5350 gnd.n1547 585
R9690 gnd.n5435 gnd.n5434 585
R9691 gnd.n5434 gnd.n5433 585
R9692 gnd.n5436 gnd.n1542 585
R9693 gnd.n5290 gnd.n1542 585
R9694 gnd.n5438 gnd.n5437 585
R9695 gnd.n5439 gnd.n5438 585
R9696 gnd.n1527 gnd.n1526 585
R9697 gnd.n5281 gnd.n1527 585
R9698 gnd.n5447 gnd.n5446 585
R9699 gnd.n5446 gnd.n5445 585
R9700 gnd.n5448 gnd.n1520 585
R9701 gnd.n5275 gnd.n1520 585
R9702 gnd.n5450 gnd.n5449 585
R9703 gnd.n5451 gnd.n5450 585
R9704 gnd.n1521 gnd.n1519 585
R9705 gnd.n5268 gnd.n1519 585
R9706 gnd.n1503 gnd.n1497 585
R9707 gnd.n5457 gnd.n1503 585
R9708 gnd.n5462 gnd.n1495 585
R9709 gnd.n5307 gnd.n1495 585
R9710 gnd.n5464 gnd.n5463 585
R9711 gnd.n5465 gnd.n5464 585
R9712 gnd.n1494 gnd.n1334 585
R9713 gnd.n5632 gnd.n1335 585
R9714 gnd.n5631 gnd.n1336 585
R9715 gnd.n1411 gnd.n1337 585
R9716 gnd.n5624 gnd.n1343 585
R9717 gnd.n5623 gnd.n1344 585
R9718 gnd.n1414 gnd.n1345 585
R9719 gnd.n5616 gnd.n1351 585
R9720 gnd.n5615 gnd.n1352 585
R9721 gnd.n1416 gnd.n1353 585
R9722 gnd.n5608 gnd.n1359 585
R9723 gnd.n5607 gnd.n1360 585
R9724 gnd.n1419 gnd.n1361 585
R9725 gnd.n5600 gnd.n1367 585
R9726 gnd.n5599 gnd.n1368 585
R9727 gnd.n1421 gnd.n1369 585
R9728 gnd.n5592 gnd.n1377 585
R9729 gnd.n5591 gnd.n5588 585
R9730 gnd.n1380 gnd.n1378 585
R9731 gnd.n5586 gnd.n1380 585
R9732 gnd.n7189 gnd.n7188 585
R9733 gnd.n6915 gnd.n6914 585
R9734 gnd.n6972 gnd.n6971 585
R9735 gnd.n6924 gnd.n6923 585
R9736 gnd.n6967 gnd.n6966 585
R9737 gnd.n6965 gnd.n6964 585
R9738 gnd.n6963 gnd.n6962 585
R9739 gnd.n6956 gnd.n6926 585
R9740 gnd.n6958 gnd.n6957 585
R9741 gnd.n6955 gnd.n6954 585
R9742 gnd.n6953 gnd.n6952 585
R9743 gnd.n6946 gnd.n6928 585
R9744 gnd.n6948 gnd.n6947 585
R9745 gnd.n6945 gnd.n6944 585
R9746 gnd.n6943 gnd.n6942 585
R9747 gnd.n6936 gnd.n6930 585
R9748 gnd.n6938 gnd.n6937 585
R9749 gnd.n6935 gnd.n6934 585
R9750 gnd.n6933 gnd.n171 585
R9751 gnd.n7186 gnd.n171 585
R9752 gnd.n7192 gnd.n169 585
R9753 gnd.n7247 gnd.n169 585
R9754 gnd.n7194 gnd.n7193 585
R9755 gnd.n7193 gnd.n167 585
R9756 gnd.n7195 gnd.n160 585
R9757 gnd.n7253 gnd.n160 585
R9758 gnd.n7197 gnd.n7196 585
R9759 gnd.n7196 gnd.n152 585
R9760 gnd.n7198 gnd.n151 585
R9761 gnd.n7259 gnd.n151 585
R9762 gnd.n7200 gnd.n7199 585
R9763 gnd.n7199 gnd.n142 585
R9764 gnd.n7201 gnd.n141 585
R9765 gnd.n7265 gnd.n141 585
R9766 gnd.n7203 gnd.n7202 585
R9767 gnd.n7202 gnd.n133 585
R9768 gnd.n7204 gnd.n132 585
R9769 gnd.n7271 gnd.n132 585
R9770 gnd.n7206 gnd.n7205 585
R9771 gnd.n7205 gnd.n130 585
R9772 gnd.n7207 gnd.n122 585
R9773 gnd.n7277 gnd.n122 585
R9774 gnd.n7209 gnd.n7208 585
R9775 gnd.n7208 gnd.n120 585
R9776 gnd.n7210 gnd.n113 585
R9777 gnd.n7283 gnd.n113 585
R9778 gnd.n7212 gnd.n7211 585
R9779 gnd.n7211 gnd.n111 585
R9780 gnd.n7213 gnd.n103 585
R9781 gnd.n7289 gnd.n103 585
R9782 gnd.n7215 gnd.n7214 585
R9783 gnd.n7216 gnd.n7215 585
R9784 gnd.n175 gnd.n92 585
R9785 gnd.n7295 gnd.n92 585
R9786 gnd.n6893 gnd.n6892 585
R9787 gnd.n6892 gnd.n6891 585
R9788 gnd.n72 gnd.n71 585
R9789 gnd.n6884 gnd.n72 585
R9790 gnd.n7305 gnd.n7304 585
R9791 gnd.n7304 gnd.n7303 585
R9792 gnd.n7306 gnd.n70 585
R9793 gnd.n5395 gnd.n70 585
R9794 gnd.n1609 gnd.n68 585
R9795 gnd.n1609 gnd.n1603 585
R9796 gnd.n5370 gnd.n1610 585
R9797 gnd.n5386 gnd.n1610 585
R9798 gnd.n5371 gnd.n1593 585
R9799 gnd.n5404 gnd.n1593 585
R9800 gnd.n1614 gnd.n1587 585
R9801 gnd.n5409 gnd.n1587 585
R9802 gnd.n5376 gnd.n5375 585
R9803 gnd.n5377 gnd.n5376 585
R9804 gnd.n1613 gnd.n1577 585
R9805 gnd.n5415 gnd.n1577 585
R9806 gnd.n5367 gnd.n5366 585
R9807 gnd.n5366 gnd.n5365 585
R9808 gnd.n1616 gnd.n1570 585
R9809 gnd.n5421 gnd.n1570 585
R9810 gnd.n5357 gnd.n5356 585
R9811 gnd.n5358 gnd.n5357 585
R9812 gnd.n1619 gnd.n1560 585
R9813 gnd.n5427 gnd.n1560 585
R9814 gnd.n5352 gnd.n5351 585
R9815 gnd.n5351 gnd.n5350 585
R9816 gnd.n1621 gnd.n1550 585
R9817 gnd.n5433 gnd.n1550 585
R9818 gnd.n5293 gnd.n5291 585
R9819 gnd.n5291 gnd.n5290 585
R9820 gnd.n5294 gnd.n1540 585
R9821 gnd.n5439 gnd.n1540 585
R9822 gnd.n5295 gnd.n5273 585
R9823 gnd.n5281 gnd.n5273 585
R9824 gnd.n5271 gnd.n1530 585
R9825 gnd.n5445 gnd.n1530 585
R9826 gnd.n5299 gnd.n5270 585
R9827 gnd.n5275 gnd.n5270 585
R9828 gnd.n5300 gnd.n1517 585
R9829 gnd.n5451 gnd.n1517 585
R9830 gnd.n5301 gnd.n5269 585
R9831 gnd.n5269 gnd.n5268 585
R9832 gnd.n1638 gnd.n1501 585
R9833 gnd.n5457 gnd.n1501 585
R9834 gnd.n5306 gnd.n5305 585
R9835 gnd.n5307 gnd.n5306 585
R9836 gnd.n1637 gnd.n1492 585
R9837 gnd.n5465 gnd.n1492 585
R9838 gnd.n3597 gnd.n2264 585
R9839 gnd.n2264 gnd.n2241 585
R9840 gnd.n3598 gnd.n2325 585
R9841 gnd.n2325 gnd.n2315 585
R9842 gnd.n3600 gnd.n3599 585
R9843 gnd.n3601 gnd.n3600 585
R9844 gnd.n2326 gnd.n2324 585
R9845 gnd.n2333 gnd.n2324 585
R9846 gnd.n3591 gnd.n3590 585
R9847 gnd.n3590 gnd.n3589 585
R9848 gnd.n2329 gnd.n2328 585
R9849 gnd.n3316 gnd.n2329 585
R9850 gnd.n3302 gnd.n2352 585
R9851 gnd.n2352 gnd.n2342 585
R9852 gnd.n3304 gnd.n3303 585
R9853 gnd.n3305 gnd.n3304 585
R9854 gnd.n2353 gnd.n2351 585
R9855 gnd.n2351 gnd.n2349 585
R9856 gnd.n3297 gnd.n3296 585
R9857 gnd.n3296 gnd.n3295 585
R9858 gnd.n2356 gnd.n2355 585
R9859 gnd.n2365 gnd.n2356 585
R9860 gnd.n3253 gnd.n2379 585
R9861 gnd.n2379 gnd.n2364 585
R9862 gnd.n3255 gnd.n3254 585
R9863 gnd.n3256 gnd.n3255 585
R9864 gnd.n2380 gnd.n2378 585
R9865 gnd.n2387 gnd.n2378 585
R9866 gnd.n3248 gnd.n3247 585
R9867 gnd.n3247 gnd.n3246 585
R9868 gnd.n2383 gnd.n2382 585
R9869 gnd.n3227 gnd.n2383 585
R9870 gnd.n3213 gnd.n2407 585
R9871 gnd.n2407 gnd.n2396 585
R9872 gnd.n3215 gnd.n3214 585
R9873 gnd.n3216 gnd.n3215 585
R9874 gnd.n2408 gnd.n2406 585
R9875 gnd.n2406 gnd.n2403 585
R9876 gnd.n3208 gnd.n3207 585
R9877 gnd.n3207 gnd.n3206 585
R9878 gnd.n2411 gnd.n2410 585
R9879 gnd.n2421 gnd.n2411 585
R9880 gnd.n3168 gnd.n2434 585
R9881 gnd.n2434 gnd.n2420 585
R9882 gnd.n3170 gnd.n3169 585
R9883 gnd.n3171 gnd.n3170 585
R9884 gnd.n2435 gnd.n2433 585
R9885 gnd.n2442 gnd.n2433 585
R9886 gnd.n3163 gnd.n3162 585
R9887 gnd.n3162 gnd.n3161 585
R9888 gnd.n2438 gnd.n2437 585
R9889 gnd.n3142 gnd.n2438 585
R9890 gnd.n3128 gnd.n2461 585
R9891 gnd.n2461 gnd.n2451 585
R9892 gnd.n3130 gnd.n3129 585
R9893 gnd.n3131 gnd.n3130 585
R9894 gnd.n2462 gnd.n2460 585
R9895 gnd.n3119 gnd.n2460 585
R9896 gnd.n3123 gnd.n3122 585
R9897 gnd.n3122 gnd.n3121 585
R9898 gnd.n2465 gnd.n2464 585
R9899 gnd.n3074 gnd.n2465 585
R9900 gnd.n2567 gnd.n2566 585
R9901 gnd.n2568 gnd.n2567 585
R9902 gnd.n2547 gnd.n2546 585
R9903 gnd.n2550 gnd.n2547 585
R9904 gnd.n3084 gnd.n3083 585
R9905 gnd.n3083 gnd.n3082 585
R9906 gnd.n3085 gnd.n2541 585
R9907 gnd.n2577 gnd.n2541 585
R9908 gnd.n3087 gnd.n3086 585
R9909 gnd.n3088 gnd.n3087 585
R9910 gnd.n2542 gnd.n2540 585
R9911 gnd.n3052 gnd.n2540 585
R9912 gnd.n3036 gnd.n3035 585
R9913 gnd.n3035 gnd.n2528 585
R9914 gnd.n3037 gnd.n2592 585
R9915 gnd.n2592 gnd.n2527 585
R9916 gnd.n3039 gnd.n3038 585
R9917 gnd.n3040 gnd.n3039 585
R9918 gnd.n2593 gnd.n2591 585
R9919 gnd.n2591 gnd.n2588 585
R9920 gnd.n3028 gnd.n3027 585
R9921 gnd.n3027 gnd.n3026 585
R9922 gnd.n2596 gnd.n2595 585
R9923 gnd.n2603 gnd.n2596 585
R9924 gnd.n3002 gnd.n3001 585
R9925 gnd.n3003 gnd.n3002 585
R9926 gnd.n2615 gnd.n2614 585
R9927 gnd.n2622 gnd.n2614 585
R9928 gnd.n2997 gnd.n2996 585
R9929 gnd.n2996 gnd.n2995 585
R9930 gnd.n2618 gnd.n2617 585
R9931 gnd.n2985 gnd.n2618 585
R9932 gnd.n2972 gnd.n2642 585
R9933 gnd.n2642 gnd.n2641 585
R9934 gnd.n2974 gnd.n2973 585
R9935 gnd.n2975 gnd.n2974 585
R9936 gnd.n2643 gnd.n2640 585
R9937 gnd.n2650 gnd.n2640 585
R9938 gnd.n2967 gnd.n2966 585
R9939 gnd.n2966 gnd.n2965 585
R9940 gnd.n2646 gnd.n2645 585
R9941 gnd.n2954 gnd.n2646 585
R9942 gnd.n2941 gnd.n2667 585
R9943 gnd.n2667 gnd.n2666 585
R9944 gnd.n2943 gnd.n2942 585
R9945 gnd.n2944 gnd.n2943 585
R9946 gnd.n2937 gnd.n2665 585
R9947 gnd.n2936 gnd.n2935 585
R9948 gnd.n2670 gnd.n2669 585
R9949 gnd.n2933 gnd.n2670 585
R9950 gnd.n2692 gnd.n2691 585
R9951 gnd.n2695 gnd.n2694 585
R9952 gnd.n2693 gnd.n2688 585
R9953 gnd.n2700 gnd.n2699 585
R9954 gnd.n2702 gnd.n2701 585
R9955 gnd.n2705 gnd.n2704 585
R9956 gnd.n2703 gnd.n2686 585
R9957 gnd.n2710 gnd.n2709 585
R9958 gnd.n2712 gnd.n2711 585
R9959 gnd.n2715 gnd.n2714 585
R9960 gnd.n2713 gnd.n2684 585
R9961 gnd.n2720 gnd.n2719 585
R9962 gnd.n2724 gnd.n2721 585
R9963 gnd.n2725 gnd.n2662 585
R9964 gnd.n3603 gnd.n2279 585
R9965 gnd.n3670 gnd.n3669 585
R9966 gnd.n3672 gnd.n3671 585
R9967 gnd.n3674 gnd.n3673 585
R9968 gnd.n3676 gnd.n3675 585
R9969 gnd.n3678 gnd.n3677 585
R9970 gnd.n3680 gnd.n3679 585
R9971 gnd.n3682 gnd.n3681 585
R9972 gnd.n3684 gnd.n3683 585
R9973 gnd.n3686 gnd.n3685 585
R9974 gnd.n3688 gnd.n3687 585
R9975 gnd.n3690 gnd.n3689 585
R9976 gnd.n3692 gnd.n3691 585
R9977 gnd.n3695 gnd.n3694 585
R9978 gnd.n3693 gnd.n2267 585
R9979 gnd.n3699 gnd.n2265 585
R9980 gnd.n3701 gnd.n3700 585
R9981 gnd.n3702 gnd.n3701 585
R9982 gnd.n3604 gnd.n2320 585
R9983 gnd.n3604 gnd.n2241 585
R9984 gnd.n3606 gnd.n3605 585
R9985 gnd.n3605 gnd.n2315 585
R9986 gnd.n3602 gnd.n2319 585
R9987 gnd.n3602 gnd.n3601 585
R9988 gnd.n3581 gnd.n2321 585
R9989 gnd.n2333 gnd.n2321 585
R9990 gnd.n3580 gnd.n2331 585
R9991 gnd.n3589 gnd.n2331 585
R9992 gnd.n3315 gnd.n2338 585
R9993 gnd.n3316 gnd.n3315 585
R9994 gnd.n3314 gnd.n3313 585
R9995 gnd.n3314 gnd.n2342 585
R9996 gnd.n3312 gnd.n2344 585
R9997 gnd.n3305 gnd.n2344 585
R9998 gnd.n2357 gnd.n2345 585
R9999 gnd.n2357 gnd.n2349 585
R10000 gnd.n3261 gnd.n2358 585
R10001 gnd.n3295 gnd.n2358 585
R10002 gnd.n3260 gnd.n3259 585
R10003 gnd.n3259 gnd.n2365 585
R10004 gnd.n3258 gnd.n2373 585
R10005 gnd.n3258 gnd.n2364 585
R10006 gnd.n3257 gnd.n2375 585
R10007 gnd.n3257 gnd.n3256 585
R10008 gnd.n3236 gnd.n2374 585
R10009 gnd.n2387 gnd.n2374 585
R10010 gnd.n3235 gnd.n2385 585
R10011 gnd.n3246 gnd.n2385 585
R10012 gnd.n3226 gnd.n2392 585
R10013 gnd.n3227 gnd.n3226 585
R10014 gnd.n3225 gnd.n3224 585
R10015 gnd.n3225 gnd.n2396 585
R10016 gnd.n3223 gnd.n2398 585
R10017 gnd.n3216 gnd.n2398 585
R10018 gnd.n2413 gnd.n2399 585
R10019 gnd.n2413 gnd.n2403 585
R10020 gnd.n3176 gnd.n2414 585
R10021 gnd.n3206 gnd.n2414 585
R10022 gnd.n3175 gnd.n3174 585
R10023 gnd.n3174 gnd.n2421 585
R10024 gnd.n3173 gnd.n2428 585
R10025 gnd.n3173 gnd.n2420 585
R10026 gnd.n3172 gnd.n2430 585
R10027 gnd.n3172 gnd.n3171 585
R10028 gnd.n3151 gnd.n2429 585
R10029 gnd.n2442 gnd.n2429 585
R10030 gnd.n3150 gnd.n2440 585
R10031 gnd.n3161 gnd.n2440 585
R10032 gnd.n3141 gnd.n2447 585
R10033 gnd.n3142 gnd.n3141 585
R10034 gnd.n3140 gnd.n3139 585
R10035 gnd.n3140 gnd.n2451 585
R10036 gnd.n3138 gnd.n2453 585
R10037 gnd.n3131 gnd.n2453 585
R10038 gnd.n3118 gnd.n2454 585
R10039 gnd.n3119 gnd.n3118 585
R10040 gnd.n3071 gnd.n2467 585
R10041 gnd.n3121 gnd.n2467 585
R10042 gnd.n3073 gnd.n3072 585
R10043 gnd.n3074 gnd.n3073 585
R10044 gnd.n3066 gnd.n2569 585
R10045 gnd.n2569 gnd.n2568 585
R10046 gnd.n3064 gnd.n3063 585
R10047 gnd.n3063 gnd.n2550 585
R10048 gnd.n3061 gnd.n2548 585
R10049 gnd.n3082 gnd.n2548 585
R10050 gnd.n2579 gnd.n2578 585
R10051 gnd.n2578 gnd.n2577 585
R10052 gnd.n3055 gnd.n2538 585
R10053 gnd.n3088 gnd.n2538 585
R10054 gnd.n3054 gnd.n3053 585
R10055 gnd.n3053 gnd.n3052 585
R10056 gnd.n3050 gnd.n2581 585
R10057 gnd.n3050 gnd.n2528 585
R10058 gnd.n3049 gnd.n3048 585
R10059 gnd.n3049 gnd.n2527 585
R10060 gnd.n2584 gnd.n2583 585
R10061 gnd.n3040 gnd.n2583 585
R10062 gnd.n3008 gnd.n3007 585
R10063 gnd.n3007 gnd.n2588 585
R10064 gnd.n3009 gnd.n2597 585
R10065 gnd.n3026 gnd.n2597 585
R10066 gnd.n3006 gnd.n3005 585
R10067 gnd.n3005 gnd.n2603 585
R10068 gnd.n3004 gnd.n2611 585
R10069 gnd.n3004 gnd.n3003 585
R10070 gnd.n2989 gnd.n2612 585
R10071 gnd.n2622 gnd.n2612 585
R10072 gnd.n2988 gnd.n2620 585
R10073 gnd.n2995 gnd.n2620 585
R10074 gnd.n2987 gnd.n2986 585
R10075 gnd.n2986 gnd.n2985 585
R10076 gnd.n2631 gnd.n2628 585
R10077 gnd.n2641 gnd.n2631 585
R10078 gnd.n2977 gnd.n2976 585
R10079 gnd.n2976 gnd.n2975 585
R10080 gnd.n2637 gnd.n2636 585
R10081 gnd.n2650 gnd.n2637 585
R10082 gnd.n2957 gnd.n2648 585
R10083 gnd.n2965 gnd.n2648 585
R10084 gnd.n2956 gnd.n2955 585
R10085 gnd.n2955 gnd.n2954 585
R10086 gnd.n2657 gnd.n2655 585
R10087 gnd.n2666 gnd.n2657 585
R10088 gnd.n2946 gnd.n2945 585
R10089 gnd.n2945 gnd.n2944 585
R10090 gnd.n5075 gnd.n1776 585
R10091 gnd.n1776 gnd.n1732 585
R10092 gnd.n5077 gnd.n5076 585
R10093 gnd.n5078 gnd.n5077 585
R10094 gnd.n4986 gnd.n1775 585
R10095 gnd.n1780 gnd.n1775 585
R10096 gnd.n4985 gnd.n4984 585
R10097 gnd.n4984 gnd.n4983 585
R10098 gnd.n1778 gnd.n1777 585
R10099 gnd.n4959 gnd.n1778 585
R10100 gnd.n4971 gnd.n4970 585
R10101 gnd.n4972 gnd.n4971 585
R10102 gnd.n4969 gnd.n1791 585
R10103 gnd.n1791 gnd.n1788 585
R10104 gnd.n4968 gnd.n4967 585
R10105 gnd.n4967 gnd.n4966 585
R10106 gnd.n1793 gnd.n1792 585
R10107 gnd.n1806 gnd.n1793 585
R10108 gnd.n4925 gnd.n4924 585
R10109 gnd.n4924 gnd.n1805 585
R10110 gnd.n4926 gnd.n1818 585
R10111 gnd.n4913 gnd.n1818 585
R10112 gnd.n4928 gnd.n4927 585
R10113 gnd.n4929 gnd.n4928 585
R10114 gnd.n4923 gnd.n1817 585
R10115 gnd.n1817 gnd.n1812 585
R10116 gnd.n4922 gnd.n4921 585
R10117 gnd.n4921 gnd.n4920 585
R10118 gnd.n1820 gnd.n1819 585
R10119 gnd.n1826 gnd.n1820 585
R10120 gnd.n4906 gnd.n4905 585
R10121 gnd.n4907 gnd.n4906 585
R10122 gnd.n4904 gnd.n1828 585
R10123 gnd.n1834 gnd.n1828 585
R10124 gnd.n4903 gnd.n4902 585
R10125 gnd.n4902 gnd.n4901 585
R10126 gnd.n1830 gnd.n1829 585
R10127 gnd.n1845 gnd.n1830 585
R10128 gnd.n4889 gnd.n4888 585
R10129 gnd.t296 gnd.n4889 585
R10130 gnd.n4887 gnd.n1846 585
R10131 gnd.n1846 gnd.n1842 585
R10132 gnd.n4886 gnd.n4885 585
R10133 gnd.n4885 gnd.n4884 585
R10134 gnd.n1848 gnd.n1847 585
R10135 gnd.n1849 gnd.n1848 585
R10136 gnd.n4842 gnd.n1871 585
R10137 gnd.n4842 gnd.n4841 585
R10138 gnd.n4844 gnd.n4843 585
R10139 gnd.n4843 gnd.n1857 585
R10140 gnd.n4845 gnd.n1869 585
R10141 gnd.n4825 gnd.n1869 585
R10142 gnd.n4847 gnd.n4846 585
R10143 gnd.n4848 gnd.n4847 585
R10144 gnd.n1870 gnd.n1868 585
R10145 gnd.n1868 gnd.n1864 585
R10146 gnd.n1899 gnd.n1877 585
R10147 gnd.n4820 gnd.n1877 585
R10148 gnd.n1901 gnd.n1900 585
R10149 gnd.n1901 gnd.n1876 585
R10150 gnd.n4792 gnd.n1898 585
R10151 gnd.n4792 gnd.n4791 585
R10152 gnd.n4794 gnd.n4793 585
R10153 gnd.n4793 gnd.n1884 585
R10154 gnd.n4795 gnd.n1896 585
R10155 gnd.n4783 gnd.n1896 585
R10156 gnd.n4797 gnd.n4796 585
R10157 gnd.n4798 gnd.n4797 585
R10158 gnd.n1897 gnd.n1895 585
R10159 gnd.n1895 gnd.n1891 585
R10160 gnd.n4777 gnd.n4776 585
R10161 gnd.n4778 gnd.n4777 585
R10162 gnd.n4775 gnd.n1906 585
R10163 gnd.n1911 gnd.n1906 585
R10164 gnd.n4774 gnd.n4773 585
R10165 gnd.n4773 gnd.n4772 585
R10166 gnd.n1908 gnd.n1907 585
R10167 gnd.n4748 gnd.n1908 585
R10168 gnd.n4760 gnd.n4759 585
R10169 gnd.n4761 gnd.n4760 585
R10170 gnd.n4758 gnd.n1921 585
R10171 gnd.n1921 gnd.n1917 585
R10172 gnd.n4757 gnd.n4756 585
R10173 gnd.n4756 gnd.n4755 585
R10174 gnd.n1923 gnd.n1922 585
R10175 gnd.n1929 gnd.n1923 585
R10176 gnd.n4741 gnd.n4740 585
R10177 gnd.n4742 gnd.n4741 585
R10178 gnd.n4739 gnd.n1931 585
R10179 gnd.n1938 gnd.n1931 585
R10180 gnd.n4738 gnd.n4737 585
R10181 gnd.n4737 gnd.n4736 585
R10182 gnd.n1933 gnd.n1932 585
R10183 gnd.n1947 gnd.n1933 585
R10184 gnd.n4723 gnd.n4722 585
R10185 gnd.n4724 gnd.n4723 585
R10186 gnd.n4721 gnd.n1948 585
R10187 gnd.n4716 gnd.n1948 585
R10188 gnd.n4720 gnd.n4719 585
R10189 gnd.n4719 gnd.n4718 585
R10190 gnd.n1950 gnd.n1949 585
R10191 gnd.n1951 gnd.n1950 585
R10192 gnd.n4704 gnd.n4703 585
R10193 gnd.n4705 gnd.n4704 585
R10194 gnd.n4702 gnd.n1956 585
R10195 gnd.n1961 gnd.n1956 585
R10196 gnd.n4701 gnd.n4700 585
R10197 gnd.n4700 gnd.n4699 585
R10198 gnd.n1958 gnd.n1957 585
R10199 gnd.n1959 gnd.n1958 585
R10200 gnd.n4656 gnd.n4655 585
R10201 gnd.n4657 gnd.n4656 585
R10202 gnd.n4654 gnd.n1979 585
R10203 gnd.n4650 gnd.n1979 585
R10204 gnd.n4653 gnd.n4652 585
R10205 gnd.n4652 gnd.n4651 585
R10206 gnd.n1981 gnd.n1980 585
R10207 gnd.n4639 gnd.n1981 585
R10208 gnd.n4619 gnd.n4618 585
R10209 gnd.n4618 gnd.n1987 585
R10210 gnd.n4620 gnd.n1999 585
R10211 gnd.n4607 gnd.n1999 585
R10212 gnd.n4622 gnd.n4621 585
R10213 gnd.n4623 gnd.n4622 585
R10214 gnd.n4617 gnd.n1998 585
R10215 gnd.n1998 gnd.t1 585
R10216 gnd.n4616 gnd.n4615 585
R10217 gnd.n4615 gnd.n4614 585
R10218 gnd.n2001 gnd.n2000 585
R10219 gnd.n2008 gnd.n2001 585
R10220 gnd.n4602 gnd.n4601 585
R10221 gnd.n4603 gnd.n4602 585
R10222 gnd.n4600 gnd.n2010 585
R10223 gnd.n2016 gnd.n2010 585
R10224 gnd.n4599 gnd.n4598 585
R10225 gnd.n4598 gnd.n4597 585
R10226 gnd.n2012 gnd.n2011 585
R10227 gnd.n2025 gnd.n2012 585
R10228 gnd.n4583 gnd.n4582 585
R10229 gnd.n4584 gnd.n4583 585
R10230 gnd.n4581 gnd.n2026 585
R10231 gnd.n4576 gnd.n2026 585
R10232 gnd.n4580 gnd.n4579 585
R10233 gnd.n4579 gnd.n4578 585
R10234 gnd.n2028 gnd.n2027 585
R10235 gnd.n4566 gnd.n2028 585
R10236 gnd.n4509 gnd.n4508 585
R10237 gnd.n4509 gnd.n2033 585
R10238 gnd.n4511 gnd.n4510 585
R10239 gnd.n4510 gnd.n2035 585
R10240 gnd.n4512 gnd.n4505 585
R10241 gnd.n4505 gnd.n4504 585
R10242 gnd.n4514 gnd.n4513 585
R10243 gnd.n4515 gnd.n4514 585
R10244 gnd.n4507 gnd.n4503 585
R10245 gnd.n4503 gnd.n4502 585
R10246 gnd.n4506 gnd.n4424 585
R10247 gnd.n4521 gnd.n4424 585
R10248 gnd.n1200 gnd.n1199 585
R10249 gnd.n4423 gnd.n1200 585
R10250 gnd.n5780 gnd.n5779 585
R10251 gnd.n5779 gnd.n5778 585
R10252 gnd.n5781 gnd.n1178 585
R10253 gnd.n4492 gnd.n1178 585
R10254 gnd.n5846 gnd.n5845 585
R10255 gnd.n5844 gnd.n1177 585
R10256 gnd.n5843 gnd.n1176 585
R10257 gnd.n5848 gnd.n1176 585
R10258 gnd.n5842 gnd.n5841 585
R10259 gnd.n5840 gnd.n5839 585
R10260 gnd.n5838 gnd.n5837 585
R10261 gnd.n5836 gnd.n5835 585
R10262 gnd.n5834 gnd.n5833 585
R10263 gnd.n5832 gnd.n5831 585
R10264 gnd.n5830 gnd.n5829 585
R10265 gnd.n5828 gnd.n5827 585
R10266 gnd.n5826 gnd.n5825 585
R10267 gnd.n5824 gnd.n5823 585
R10268 gnd.n5822 gnd.n5821 585
R10269 gnd.n5820 gnd.n5819 585
R10270 gnd.n5818 gnd.n5817 585
R10271 gnd.n5816 gnd.n5815 585
R10272 gnd.n5814 gnd.n5813 585
R10273 gnd.n5812 gnd.n5811 585
R10274 gnd.n5810 gnd.n5809 585
R10275 gnd.n5808 gnd.n5807 585
R10276 gnd.n5806 gnd.n5805 585
R10277 gnd.n5804 gnd.n5803 585
R10278 gnd.n5802 gnd.n5801 585
R10279 gnd.n5800 gnd.n5799 585
R10280 gnd.n5798 gnd.n5797 585
R10281 gnd.n5796 gnd.n5795 585
R10282 gnd.n5794 gnd.n5793 585
R10283 gnd.n5792 gnd.n5791 585
R10284 gnd.n5790 gnd.n5789 585
R10285 gnd.n5788 gnd.n5787 585
R10286 gnd.n5786 gnd.n1140 585
R10287 gnd.n5851 gnd.n5850 585
R10288 gnd.n1142 gnd.n1139 585
R10289 gnd.n4430 gnd.n4429 585
R10290 gnd.n4432 gnd.n4431 585
R10291 gnd.n4435 gnd.n4434 585
R10292 gnd.n4437 gnd.n4436 585
R10293 gnd.n4439 gnd.n4438 585
R10294 gnd.n4441 gnd.n4440 585
R10295 gnd.n4443 gnd.n4442 585
R10296 gnd.n4445 gnd.n4444 585
R10297 gnd.n4447 gnd.n4446 585
R10298 gnd.n4449 gnd.n4448 585
R10299 gnd.n4451 gnd.n4450 585
R10300 gnd.n4453 gnd.n4452 585
R10301 gnd.n4455 gnd.n4454 585
R10302 gnd.n4457 gnd.n4456 585
R10303 gnd.n4459 gnd.n4458 585
R10304 gnd.n4461 gnd.n4460 585
R10305 gnd.n4463 gnd.n4462 585
R10306 gnd.n4465 gnd.n4464 585
R10307 gnd.n4467 gnd.n4466 585
R10308 gnd.n4469 gnd.n4468 585
R10309 gnd.n4471 gnd.n4470 585
R10310 gnd.n4473 gnd.n4472 585
R10311 gnd.n4475 gnd.n4474 585
R10312 gnd.n4477 gnd.n4476 585
R10313 gnd.n4479 gnd.n4478 585
R10314 gnd.n4481 gnd.n4480 585
R10315 gnd.n4483 gnd.n4482 585
R10316 gnd.n4485 gnd.n4484 585
R10317 gnd.n4487 gnd.n4486 585
R10318 gnd.n4489 gnd.n4488 585
R10319 gnd.n4491 gnd.n4490 585
R10320 gnd.n5082 gnd.n5081 585
R10321 gnd.n5084 gnd.n5083 585
R10322 gnd.n5086 gnd.n5085 585
R10323 gnd.n5088 gnd.n5087 585
R10324 gnd.n5090 gnd.n5089 585
R10325 gnd.n5092 gnd.n5091 585
R10326 gnd.n5094 gnd.n5093 585
R10327 gnd.n5096 gnd.n5095 585
R10328 gnd.n5098 gnd.n5097 585
R10329 gnd.n5100 gnd.n5099 585
R10330 gnd.n5102 gnd.n5101 585
R10331 gnd.n5104 gnd.n5103 585
R10332 gnd.n5106 gnd.n5105 585
R10333 gnd.n5108 gnd.n5107 585
R10334 gnd.n5110 gnd.n5109 585
R10335 gnd.n5112 gnd.n5111 585
R10336 gnd.n5114 gnd.n5113 585
R10337 gnd.n5116 gnd.n5115 585
R10338 gnd.n5118 gnd.n5117 585
R10339 gnd.n5120 gnd.n5119 585
R10340 gnd.n5122 gnd.n5121 585
R10341 gnd.n5124 gnd.n5123 585
R10342 gnd.n5126 gnd.n5125 585
R10343 gnd.n5128 gnd.n5127 585
R10344 gnd.n5130 gnd.n5129 585
R10345 gnd.n5132 gnd.n5131 585
R10346 gnd.n5134 gnd.n5133 585
R10347 gnd.n5136 gnd.n5135 585
R10348 gnd.n5138 gnd.n5137 585
R10349 gnd.n5141 gnd.n5140 585
R10350 gnd.n5143 gnd.n5142 585
R10351 gnd.n5145 gnd.n5144 585
R10352 gnd.n5147 gnd.n5146 585
R10353 gnd.n5008 gnd.n1455 585
R10354 gnd.n5010 gnd.n5009 585
R10355 gnd.n5012 gnd.n5011 585
R10356 gnd.n5014 gnd.n5013 585
R10357 gnd.n5017 gnd.n5016 585
R10358 gnd.n5019 gnd.n5018 585
R10359 gnd.n5021 gnd.n5020 585
R10360 gnd.n5023 gnd.n5022 585
R10361 gnd.n5025 gnd.n5024 585
R10362 gnd.n5027 gnd.n5026 585
R10363 gnd.n5029 gnd.n5028 585
R10364 gnd.n5031 gnd.n5030 585
R10365 gnd.n5033 gnd.n5032 585
R10366 gnd.n5035 gnd.n5034 585
R10367 gnd.n5037 gnd.n5036 585
R10368 gnd.n5039 gnd.n5038 585
R10369 gnd.n5041 gnd.n5040 585
R10370 gnd.n5043 gnd.n5042 585
R10371 gnd.n5045 gnd.n5044 585
R10372 gnd.n5047 gnd.n5046 585
R10373 gnd.n5049 gnd.n5048 585
R10374 gnd.n5051 gnd.n5050 585
R10375 gnd.n5053 gnd.n5052 585
R10376 gnd.n5055 gnd.n5054 585
R10377 gnd.n5057 gnd.n5056 585
R10378 gnd.n5059 gnd.n5058 585
R10379 gnd.n5061 gnd.n5060 585
R10380 gnd.n5063 gnd.n5062 585
R10381 gnd.n5065 gnd.n5064 585
R10382 gnd.n5067 gnd.n5066 585
R10383 gnd.n5069 gnd.n5068 585
R10384 gnd.n5071 gnd.n5070 585
R10385 gnd.n5073 gnd.n5072 585
R10386 gnd.n5080 gnd.n1771 585
R10387 gnd.n5080 gnd.n1732 585
R10388 gnd.n5079 gnd.n1773 585
R10389 gnd.n5079 gnd.n5078 585
R10390 gnd.n1798 gnd.n1772 585
R10391 gnd.n1780 gnd.n1772 585
R10392 gnd.n1799 gnd.n1781 585
R10393 gnd.n4983 gnd.n1781 585
R10394 gnd.n4961 gnd.n4960 585
R10395 gnd.n4960 gnd.n4959 585
R10396 gnd.n4962 gnd.n1790 585
R10397 gnd.n4972 gnd.n1790 585
R10398 gnd.n4963 gnd.n1796 585
R10399 gnd.n1796 gnd.n1788 585
R10400 gnd.n4965 gnd.n4964 585
R10401 gnd.n4966 gnd.n4965 585
R10402 gnd.n1797 gnd.n1795 585
R10403 gnd.n1806 gnd.n1795 585
R10404 gnd.n4912 gnd.n4911 585
R10405 gnd.n4912 gnd.n1805 585
R10406 gnd.n4915 gnd.n4914 585
R10407 gnd.n4914 gnd.n4913 585
R10408 gnd.n4916 gnd.n1814 585
R10409 gnd.n4929 gnd.n1814 585
R10410 gnd.n4917 gnd.n1823 585
R10411 gnd.n1823 gnd.n1812 585
R10412 gnd.n4919 gnd.n4918 585
R10413 gnd.n4920 gnd.n4919 585
R10414 gnd.n4910 gnd.n1822 585
R10415 gnd.n1826 gnd.n1822 585
R10416 gnd.n4909 gnd.n4908 585
R10417 gnd.n4908 gnd.n4907 585
R10418 gnd.n1825 gnd.n1824 585
R10419 gnd.n1834 gnd.n1825 585
R10420 gnd.n4829 gnd.n1832 585
R10421 gnd.n4901 gnd.n1832 585
R10422 gnd.n4831 gnd.n4830 585
R10423 gnd.n4830 gnd.n1845 585
R10424 gnd.n4832 gnd.n1844 585
R10425 gnd.t296 gnd.n1844 585
R10426 gnd.n4834 gnd.n4833 585
R10427 gnd.n4833 gnd.n1842 585
R10428 gnd.n4835 gnd.n1850 585
R10429 gnd.n4884 gnd.n1850 585
R10430 gnd.n4836 gnd.n1873 585
R10431 gnd.n1873 gnd.n1849 585
R10432 gnd.n4838 gnd.n4837 585
R10433 gnd.n4841 gnd.n4838 585
R10434 gnd.n4828 gnd.n1872 585
R10435 gnd.n1872 gnd.n1857 585
R10436 gnd.n4827 gnd.n4826 585
R10437 gnd.n4826 gnd.n4825 585
R10438 gnd.n4824 gnd.n1866 585
R10439 gnd.n4848 gnd.n1866 585
R10440 gnd.n4823 gnd.n4822 585
R10441 gnd.n4822 gnd.n1864 585
R10442 gnd.n4821 gnd.n1874 585
R10443 gnd.n4821 gnd.n4820 585
R10444 gnd.n4787 gnd.n1875 585
R10445 gnd.n1876 gnd.n1875 585
R10446 gnd.n4789 gnd.n4788 585
R10447 gnd.n4791 gnd.n4789 585
R10448 gnd.n4786 gnd.n1902 585
R10449 gnd.n1902 gnd.n1884 585
R10450 gnd.n4785 gnd.n4784 585
R10451 gnd.n4784 gnd.n4783 585
R10452 gnd.n4782 gnd.n1893 585
R10453 gnd.n4798 gnd.n1893 585
R10454 gnd.n4781 gnd.n4780 585
R10455 gnd.n4780 gnd.n1891 585
R10456 gnd.n4779 gnd.n1903 585
R10457 gnd.n4779 gnd.n4778 585
R10458 gnd.n4746 gnd.n1904 585
R10459 gnd.n1911 gnd.n1904 585
R10460 gnd.n4747 gnd.n1909 585
R10461 gnd.n4772 gnd.n1909 585
R10462 gnd.n4750 gnd.n4749 585
R10463 gnd.n4749 gnd.n4748 585
R10464 gnd.n4751 gnd.n1919 585
R10465 gnd.n4761 gnd.n1919 585
R10466 gnd.n4752 gnd.n1926 585
R10467 gnd.n1926 gnd.n1917 585
R10468 gnd.n4754 gnd.n4753 585
R10469 gnd.n4755 gnd.n4754 585
R10470 gnd.n4745 gnd.n1925 585
R10471 gnd.n1929 gnd.n1925 585
R10472 gnd.n4744 gnd.n4743 585
R10473 gnd.n4743 gnd.n4742 585
R10474 gnd.n1928 gnd.n1927 585
R10475 gnd.n1938 gnd.n1928 585
R10476 gnd.n4710 gnd.n1936 585
R10477 gnd.n4736 gnd.n1936 585
R10478 gnd.n4712 gnd.n4711 585
R10479 gnd.n4711 gnd.n1947 585
R10480 gnd.n4713 gnd.n1946 585
R10481 gnd.n4724 gnd.n1946 585
R10482 gnd.n4715 gnd.n4714 585
R10483 gnd.n4716 gnd.n4715 585
R10484 gnd.n4709 gnd.n1952 585
R10485 gnd.n4718 gnd.n1952 585
R10486 gnd.n4708 gnd.n4707 585
R10487 gnd.n4707 gnd.n1951 585
R10488 gnd.n4706 gnd.n1954 585
R10489 gnd.n4706 gnd.n4705 585
R10490 gnd.n4643 gnd.n1955 585
R10491 gnd.n1961 gnd.n1955 585
R10492 gnd.n4644 gnd.n1962 585
R10493 gnd.n4699 gnd.n1962 585
R10494 gnd.n4646 gnd.n4645 585
R10495 gnd.n4645 gnd.n1959 585
R10496 gnd.n4647 gnd.n1978 585
R10497 gnd.n4657 gnd.n1978 585
R10498 gnd.n4649 gnd.n4648 585
R10499 gnd.n4650 gnd.n4649 585
R10500 gnd.n4642 gnd.n1984 585
R10501 gnd.n4651 gnd.n1984 585
R10502 gnd.n4641 gnd.n4640 585
R10503 gnd.n4640 gnd.n4639 585
R10504 gnd.n1986 gnd.n1985 585
R10505 gnd.n1987 gnd.n1986 585
R10506 gnd.n4609 gnd.n4608 585
R10507 gnd.n4608 gnd.n4607 585
R10508 gnd.n4610 gnd.n1996 585
R10509 gnd.n4623 gnd.n1996 585
R10510 gnd.n4611 gnd.n2005 585
R10511 gnd.n2005 gnd.t1 585
R10512 gnd.n4613 gnd.n4612 585
R10513 gnd.n4614 gnd.n4613 585
R10514 gnd.n4606 gnd.n2004 585
R10515 gnd.n2008 gnd.n2004 585
R10516 gnd.n4605 gnd.n4604 585
R10517 gnd.n4604 gnd.n4603 585
R10518 gnd.n2007 gnd.n2006 585
R10519 gnd.n2016 gnd.n2007 585
R10520 gnd.n4570 gnd.n2014 585
R10521 gnd.n4597 gnd.n2014 585
R10522 gnd.n4572 gnd.n4571 585
R10523 gnd.n4571 gnd.n2025 585
R10524 gnd.n4573 gnd.n2024 585
R10525 gnd.n4584 gnd.n2024 585
R10526 gnd.n4575 gnd.n4574 585
R10527 gnd.n4576 gnd.n4575 585
R10528 gnd.n4569 gnd.n2029 585
R10529 gnd.n4578 gnd.n2029 585
R10530 gnd.n4568 gnd.n4567 585
R10531 gnd.n4567 gnd.n4566 585
R10532 gnd.n2032 gnd.n2031 585
R10533 gnd.n2033 gnd.n2032 585
R10534 gnd.n4499 gnd.n4498 585
R10535 gnd.n4499 gnd.n2035 585
R10536 gnd.n4500 gnd.n4497 585
R10537 gnd.n4504 gnd.n4500 585
R10538 gnd.n4517 gnd.n4516 585
R10539 gnd.n4516 gnd.n4515 585
R10540 gnd.n4518 gnd.n4426 585
R10541 gnd.n4502 gnd.n4426 585
R10542 gnd.n4520 gnd.n4519 585
R10543 gnd.n4521 gnd.n4520 585
R10544 gnd.n4496 gnd.n4425 585
R10545 gnd.n4425 gnd.n4423 585
R10546 gnd.n4495 gnd.n1202 585
R10547 gnd.n5778 gnd.n1202 585
R10548 gnd.n4494 gnd.n4493 585
R10549 gnd.n4493 gnd.n4492 585
R10550 gnd.n5987 gnd.n5986 585
R10551 gnd.n5986 gnd.n5985 585
R10552 gnd.n5988 gnd.n853 585
R10553 gnd.n5978 gnd.n853 585
R10554 gnd.n5990 gnd.n5989 585
R10555 gnd.n5991 gnd.n5990 585
R10556 gnd.n839 gnd.n838 585
R10557 gnd.n4202 gnd.n839 585
R10558 gnd.n5999 gnd.n5998 585
R10559 gnd.n5998 gnd.n5997 585
R10560 gnd.n6000 gnd.n833 585
R10561 gnd.n4196 gnd.n833 585
R10562 gnd.n6002 gnd.n6001 585
R10563 gnd.n6003 gnd.n6002 585
R10564 gnd.n819 gnd.n818 585
R10565 gnd.n4191 gnd.n819 585
R10566 gnd.n6011 gnd.n6010 585
R10567 gnd.n6010 gnd.n6009 585
R10568 gnd.n6012 gnd.n813 585
R10569 gnd.n4186 gnd.n813 585
R10570 gnd.n6014 gnd.n6013 585
R10571 gnd.n6015 gnd.n6014 585
R10572 gnd.n799 gnd.n798 585
R10573 gnd.n4219 gnd.n799 585
R10574 gnd.n6023 gnd.n6022 585
R10575 gnd.n6022 gnd.n6021 585
R10576 gnd.n6024 gnd.n793 585
R10577 gnd.n4179 gnd.n793 585
R10578 gnd.n6026 gnd.n6025 585
R10579 gnd.n6027 gnd.n6026 585
R10580 gnd.n779 gnd.n778 585
R10581 gnd.n4171 gnd.n779 585
R10582 gnd.n6035 gnd.n6034 585
R10583 gnd.n6034 gnd.n6033 585
R10584 gnd.n6036 gnd.n776 585
R10585 gnd.n4145 gnd.n776 585
R10586 gnd.n6039 gnd.n6038 585
R10587 gnd.n6040 gnd.n6039 585
R10588 gnd.n777 gnd.n762 585
R10589 gnd.n4153 gnd.n762 585
R10590 gnd.n6048 gnd.n6047 585
R10591 gnd.n6047 gnd.n6046 585
R10592 gnd.n6049 gnd.n759 585
R10593 gnd.n4134 gnd.n759 585
R10594 gnd.n6052 gnd.n6051 585
R10595 gnd.n6053 gnd.n6052 585
R10596 gnd.n760 gnd.n743 585
R10597 gnd.n4126 gnd.n743 585
R10598 gnd.n6061 gnd.n6060 585
R10599 gnd.n6060 gnd.n6059 585
R10600 gnd.n6062 gnd.n739 585
R10601 gnd.n4108 gnd.n739 585
R10602 gnd.n6065 gnd.n6064 585
R10603 gnd.n6066 gnd.n6065 585
R10604 gnd.n740 gnd.n738 585
R10605 gnd.n738 gnd.n733 585
R10606 gnd.n4098 gnd.n4097 585
R10607 gnd.n4099 gnd.n4098 585
R10608 gnd.n2174 gnd.n2173 585
R10609 gnd.n2180 gnd.n2173 585
R10610 gnd.n4092 gnd.n4091 585
R10611 gnd.n4091 gnd.n4090 585
R10612 gnd.n2177 gnd.n2176 585
R10613 gnd.n4072 gnd.n2177 585
R10614 gnd.n4057 gnd.n2200 585
R10615 gnd.n2200 gnd.n2190 585
R10616 gnd.n4059 gnd.n4058 585
R10617 gnd.n4060 gnd.n4059 585
R10618 gnd.n2201 gnd.n2199 585
R10619 gnd.n2199 gnd.n2196 585
R10620 gnd.n4052 gnd.n4051 585
R10621 gnd.n4051 gnd.n4050 585
R10622 gnd.n2204 gnd.n2203 585
R10623 gnd.n4035 gnd.n2204 585
R10624 gnd.n4022 gnd.n2225 585
R10625 gnd.n2225 gnd.n2215 585
R10626 gnd.n4024 gnd.n4023 585
R10627 gnd.n4025 gnd.n4024 585
R10628 gnd.n2226 gnd.n2224 585
R10629 gnd.n2224 gnd.n2221 585
R10630 gnd.n4017 gnd.n4016 585
R10631 gnd.n4016 gnd.n4015 585
R10632 gnd.n2229 gnd.n2228 585
R10633 gnd.n3780 gnd.n2229 585
R10634 gnd.n3996 gnd.n3995 585
R10635 gnd.n3997 gnd.n3996 585
R10636 gnd.n3992 gnd.n3781 585
R10637 gnd.n3991 gnd.n3990 585
R10638 gnd.n3988 gnd.n3783 585
R10639 gnd.n3988 gnd.n3703 585
R10640 gnd.n3987 gnd.n3986 585
R10641 gnd.n3985 gnd.n3984 585
R10642 gnd.n3983 gnd.n3788 585
R10643 gnd.n3981 gnd.n3980 585
R10644 gnd.n3979 gnd.n3789 585
R10645 gnd.n3978 gnd.n3977 585
R10646 gnd.n3975 gnd.n3794 585
R10647 gnd.n3973 gnd.n3972 585
R10648 gnd.n3971 gnd.n3795 585
R10649 gnd.n3970 gnd.n3969 585
R10650 gnd.n3967 gnd.n3800 585
R10651 gnd.n3965 gnd.n3964 585
R10652 gnd.n3963 gnd.n3801 585
R10653 gnd.n3962 gnd.n3961 585
R10654 gnd.n3959 gnd.n3806 585
R10655 gnd.n3957 gnd.n3956 585
R10656 gnd.n3955 gnd.n3807 585
R10657 gnd.n3954 gnd.n3953 585
R10658 gnd.n3951 gnd.n3815 585
R10659 gnd.n3949 gnd.n3948 585
R10660 gnd.n3947 gnd.n3816 585
R10661 gnd.n3946 gnd.n3945 585
R10662 gnd.n3943 gnd.n3821 585
R10663 gnd.n3941 gnd.n3940 585
R10664 gnd.n3939 gnd.n3822 585
R10665 gnd.n3938 gnd.n3937 585
R10666 gnd.n3935 gnd.n3827 585
R10667 gnd.n3933 gnd.n3932 585
R10668 gnd.n3931 gnd.n3828 585
R10669 gnd.n3930 gnd.n3929 585
R10670 gnd.n3927 gnd.n3833 585
R10671 gnd.n3925 gnd.n3924 585
R10672 gnd.n3923 gnd.n3834 585
R10673 gnd.n3922 gnd.n3921 585
R10674 gnd.n3919 gnd.n3841 585
R10675 gnd.n3917 gnd.n3916 585
R10676 gnd.n3915 gnd.n3842 585
R10677 gnd.n3914 gnd.n3913 585
R10678 gnd.n3911 gnd.n3847 585
R10679 gnd.n3909 gnd.n3908 585
R10680 gnd.n3907 gnd.n3848 585
R10681 gnd.n3906 gnd.n3905 585
R10682 gnd.n3903 gnd.n3853 585
R10683 gnd.n3901 gnd.n3900 585
R10684 gnd.n3899 gnd.n3854 585
R10685 gnd.n3898 gnd.n3897 585
R10686 gnd.n3895 gnd.n3859 585
R10687 gnd.n3893 gnd.n3892 585
R10688 gnd.n3891 gnd.n3860 585
R10689 gnd.n3890 gnd.n3889 585
R10690 gnd.n3887 gnd.n3865 585
R10691 gnd.n3885 gnd.n3884 585
R10692 gnd.n3883 gnd.n3866 585
R10693 gnd.n3882 gnd.n3881 585
R10694 gnd.n3879 gnd.n3873 585
R10695 gnd.n3877 gnd.n3876 585
R10696 gnd.n1070 gnd.n1069 585
R10697 gnd.n1076 gnd.n1075 585
R10698 gnd.n1078 gnd.n1077 585
R10699 gnd.n1080 gnd.n1079 585
R10700 gnd.n1082 gnd.n1081 585
R10701 gnd.n1084 gnd.n1083 585
R10702 gnd.n1086 gnd.n1085 585
R10703 gnd.n1088 gnd.n1087 585
R10704 gnd.n1090 gnd.n1089 585
R10705 gnd.n1092 gnd.n1091 585
R10706 gnd.n1094 gnd.n1093 585
R10707 gnd.n1096 gnd.n1095 585
R10708 gnd.n1098 gnd.n1097 585
R10709 gnd.n1100 gnd.n1099 585
R10710 gnd.n1102 gnd.n1101 585
R10711 gnd.n1104 gnd.n1103 585
R10712 gnd.n1106 gnd.n1105 585
R10713 gnd.n1108 gnd.n1107 585
R10714 gnd.n1110 gnd.n1109 585
R10715 gnd.n1113 gnd.n1112 585
R10716 gnd.n1111 gnd.n1049 585
R10717 gnd.n1118 gnd.n1117 585
R10718 gnd.n1120 gnd.n1119 585
R10719 gnd.n1122 gnd.n1121 585
R10720 gnd.n1124 gnd.n1123 585
R10721 gnd.n1126 gnd.n1125 585
R10722 gnd.n1128 gnd.n1127 585
R10723 gnd.n1130 gnd.n1129 585
R10724 gnd.n1132 gnd.n1131 585
R10725 gnd.n1135 gnd.n1134 585
R10726 gnd.n1133 gnd.n1040 585
R10727 gnd.n5854 gnd.n5853 585
R10728 gnd.n5856 gnd.n5855 585
R10729 gnd.n5858 gnd.n5857 585
R10730 gnd.n5860 gnd.n5859 585
R10731 gnd.n5862 gnd.n5861 585
R10732 gnd.n5864 gnd.n5863 585
R10733 gnd.n5866 gnd.n5865 585
R10734 gnd.n5868 gnd.n5867 585
R10735 gnd.n5871 gnd.n5870 585
R10736 gnd.n5873 gnd.n5872 585
R10737 gnd.n5875 gnd.n5874 585
R10738 gnd.n5877 gnd.n5876 585
R10739 gnd.n5879 gnd.n5878 585
R10740 gnd.n5881 gnd.n5880 585
R10741 gnd.n5883 gnd.n5882 585
R10742 gnd.n5885 gnd.n5884 585
R10743 gnd.n5887 gnd.n5886 585
R10744 gnd.n5889 gnd.n5888 585
R10745 gnd.n5891 gnd.n5890 585
R10746 gnd.n5893 gnd.n5892 585
R10747 gnd.n5895 gnd.n5894 585
R10748 gnd.n5897 gnd.n5896 585
R10749 gnd.n5898 gnd.n1009 585
R10750 gnd.n5900 gnd.n5899 585
R10751 gnd.n1010 gnd.n1008 585
R10752 gnd.n1011 gnd.n858 585
R10753 gnd.n5902 gnd.n858 585
R10754 gnd.n5981 gnd.n860 585
R10755 gnd.n5985 gnd.n860 585
R10756 gnd.n5980 gnd.n5979 585
R10757 gnd.n5979 gnd.n5978 585
R10758 gnd.n866 gnd.n851 585
R10759 gnd.n5991 gnd.n851 585
R10760 gnd.n4201 gnd.n4200 585
R10761 gnd.n4202 gnd.n4201 585
R10762 gnd.n4199 gnd.n841 585
R10763 gnd.n5997 gnd.n841 585
R10764 gnd.n4198 gnd.n4197 585
R10765 gnd.n4197 gnd.n4196 585
R10766 gnd.n4194 gnd.n830 585
R10767 gnd.n6003 gnd.n830 585
R10768 gnd.n4193 gnd.n4192 585
R10769 gnd.n4192 gnd.n4191 585
R10770 gnd.n4189 gnd.n821 585
R10771 gnd.n6009 gnd.n821 585
R10772 gnd.n4188 gnd.n4187 585
R10773 gnd.n4187 gnd.n4186 585
R10774 gnd.n4184 gnd.n810 585
R10775 gnd.n6015 gnd.n810 585
R10776 gnd.n4183 gnd.n2133 585
R10777 gnd.n4219 gnd.n2133 585
R10778 gnd.n4182 gnd.n801 585
R10779 gnd.n6021 gnd.n801 585
R10780 gnd.n4181 gnd.n4180 585
R10781 gnd.n4180 gnd.n4179 585
R10782 gnd.n2143 gnd.n790 585
R10783 gnd.n6027 gnd.n790 585
R10784 gnd.n4141 gnd.n2148 585
R10785 gnd.n4171 gnd.n2148 585
R10786 gnd.n4142 gnd.n781 585
R10787 gnd.n6033 gnd.n781 585
R10788 gnd.n4144 gnd.n4143 585
R10789 gnd.n4145 gnd.n4144 585
R10790 gnd.n4139 gnd.n773 585
R10791 gnd.n6040 gnd.n773 585
R10792 gnd.n4138 gnd.n2155 585
R10793 gnd.n4153 gnd.n2155 585
R10794 gnd.n4137 gnd.n764 585
R10795 gnd.n6046 gnd.n764 585
R10796 gnd.n4136 gnd.n4135 585
R10797 gnd.n4135 gnd.n4134 585
R10798 gnd.n2159 gnd.n756 585
R10799 gnd.n6053 gnd.n756 585
R10800 gnd.n4113 gnd.n4112 585
R10801 gnd.n4126 gnd.n4113 585
R10802 gnd.n4111 gnd.n745 585
R10803 gnd.n6059 gnd.n745 585
R10804 gnd.n4110 gnd.n4109 585
R10805 gnd.n4109 gnd.n4108 585
R10806 gnd.n2164 gnd.n734 585
R10807 gnd.n6066 gnd.n734 585
R10808 gnd.n4080 gnd.n4079 585
R10809 gnd.n4079 gnd.n733 585
R10810 gnd.n4078 gnd.n2171 585
R10811 gnd.n4099 gnd.n2171 585
R10812 gnd.n4077 gnd.n4076 585
R10813 gnd.n4076 gnd.n2180 585
R10814 gnd.n4075 gnd.n2178 585
R10815 gnd.n4090 gnd.n2178 585
R10816 gnd.n4074 gnd.n4073 585
R10817 gnd.n4073 gnd.n4072 585
R10818 gnd.n2189 gnd.n2187 585
R10819 gnd.n2190 gnd.n2189 585
R10820 gnd.n4041 gnd.n2197 585
R10821 gnd.n4060 gnd.n2197 585
R10822 gnd.n4040 gnd.n4039 585
R10823 gnd.n4039 gnd.n2196 585
R10824 gnd.n4038 gnd.n2205 585
R10825 gnd.n4050 gnd.n2205 585
R10826 gnd.n4037 gnd.n4036 585
R10827 gnd.n4036 gnd.n4035 585
R10828 gnd.n2214 gnd.n2212 585
R10829 gnd.n2215 gnd.n2214 585
R10830 gnd.n4006 gnd.n2222 585
R10831 gnd.n4025 gnd.n2222 585
R10832 gnd.n4005 gnd.n4004 585
R10833 gnd.n4004 gnd.n2221 585
R10834 gnd.n4003 gnd.n2230 585
R10835 gnd.n4015 gnd.n2230 585
R10836 gnd.n4002 gnd.n2238 585
R10837 gnd.n3780 gnd.n2238 585
R10838 gnd.n3704 gnd.n2237 585
R10839 gnd.n3997 gnd.n3704 585
R10840 gnd.n7249 gnd.n7248 585
R10841 gnd.n7248 gnd.n7247 585
R10842 gnd.n7250 gnd.n161 585
R10843 gnd.n167 gnd.n161 585
R10844 gnd.n7252 gnd.n7251 585
R10845 gnd.n7253 gnd.n7252 585
R10846 gnd.n149 gnd.n148 585
R10847 gnd.n152 gnd.n149 585
R10848 gnd.n7261 gnd.n7260 585
R10849 gnd.n7260 gnd.n7259 585
R10850 gnd.n7262 gnd.n143 585
R10851 gnd.n143 gnd.n142 585
R10852 gnd.n7264 gnd.n7263 585
R10853 gnd.n7265 gnd.n7264 585
R10854 gnd.n129 gnd.n128 585
R10855 gnd.n133 gnd.n129 585
R10856 gnd.n7273 gnd.n7272 585
R10857 gnd.n7272 gnd.n7271 585
R10858 gnd.n7274 gnd.n123 585
R10859 gnd.n130 gnd.n123 585
R10860 gnd.n7276 gnd.n7275 585
R10861 gnd.n7277 gnd.n7276 585
R10862 gnd.n110 gnd.n109 585
R10863 gnd.n120 gnd.n110 585
R10864 gnd.n7285 gnd.n7284 585
R10865 gnd.n7284 gnd.n7283 585
R10866 gnd.n7286 gnd.n105 585
R10867 gnd.n111 gnd.n105 585
R10868 gnd.n7288 gnd.n7287 585
R10869 gnd.n7289 gnd.n7288 585
R10870 gnd.n89 gnd.n87 585
R10871 gnd.n7216 gnd.n89 585
R10872 gnd.n7297 gnd.n7296 585
R10873 gnd.n7296 gnd.n7295 585
R10874 gnd.n88 gnd.n80 585
R10875 gnd.n6891 gnd.n88 585
R10876 gnd.n7300 gnd.n78 585
R10877 gnd.n6884 gnd.n78 585
R10878 gnd.n7302 gnd.n7301 585
R10879 gnd.n7303 gnd.n7302 585
R10880 gnd.n1600 gnd.n77 585
R10881 gnd.n5395 gnd.n77 585
R10882 gnd.n1602 gnd.n1601 585
R10883 gnd.n1603 gnd.n1602 585
R10884 gnd.n1590 gnd.n1589 585
R10885 gnd.n5386 gnd.n1589 585
R10886 gnd.n5405 gnd.n1591 585
R10887 gnd.n5405 gnd.n5404 585
R10888 gnd.n5408 gnd.n5407 585
R10889 gnd.n5409 gnd.n5408 585
R10890 gnd.n5406 gnd.n1574 585
R10891 gnd.n5377 gnd.n1574 585
R10892 gnd.n5417 gnd.n5416 585
R10893 gnd.n5416 gnd.n5415 585
R10894 gnd.n5418 gnd.n1571 585
R10895 gnd.n5365 gnd.n1571 585
R10896 gnd.n5420 gnd.n5419 585
R10897 gnd.n5421 gnd.n5420 585
R10898 gnd.n1558 gnd.n1557 585
R10899 gnd.n5358 gnd.n1558 585
R10900 gnd.n5429 gnd.n5428 585
R10901 gnd.n5428 gnd.n5427 585
R10902 gnd.n5430 gnd.n1552 585
R10903 gnd.n5350 gnd.n1552 585
R10904 gnd.n5432 gnd.n5431 585
R10905 gnd.n5433 gnd.n5432 585
R10906 gnd.n1537 gnd.n1536 585
R10907 gnd.n5290 gnd.n1537 585
R10908 gnd.n5441 gnd.n5440 585
R10909 gnd.n5440 gnd.n5439 585
R10910 gnd.n5442 gnd.n1531 585
R10911 gnd.n5281 gnd.n1531 585
R10912 gnd.n5444 gnd.n5443 585
R10913 gnd.n5445 gnd.n5444 585
R10914 gnd.n1514 gnd.n1513 585
R10915 gnd.n5275 gnd.n1514 585
R10916 gnd.n5453 gnd.n5452 585
R10917 gnd.n5452 gnd.n5451 585
R10918 gnd.n5454 gnd.n1505 585
R10919 gnd.n5268 gnd.n1505 585
R10920 gnd.n5456 gnd.n5455 585
R10921 gnd.n5457 gnd.n5456 585
R10922 gnd.n1506 gnd.n1504 585
R10923 gnd.n5307 gnd.n1504 585
R10924 gnd.n1507 gnd.n1426 585
R10925 gnd.n5465 gnd.n1426 585
R10926 gnd.n5584 gnd.n5583 585
R10927 gnd.n5582 gnd.n1425 585
R10928 gnd.n5581 gnd.n1424 585
R10929 gnd.n5586 gnd.n1424 585
R10930 gnd.n5580 gnd.n5579 585
R10931 gnd.n5578 gnd.n5577 585
R10932 gnd.n5576 gnd.n5575 585
R10933 gnd.n5574 gnd.n5573 585
R10934 gnd.n5572 gnd.n5571 585
R10935 gnd.n5570 gnd.n5569 585
R10936 gnd.n5568 gnd.n5567 585
R10937 gnd.n5566 gnd.n5565 585
R10938 gnd.n5564 gnd.n5563 585
R10939 gnd.n5562 gnd.n5561 585
R10940 gnd.n5560 gnd.n5559 585
R10941 gnd.n5558 gnd.n5557 585
R10942 gnd.n5556 gnd.n5555 585
R10943 gnd.n5554 gnd.n5553 585
R10944 gnd.n5552 gnd.n5551 585
R10945 gnd.n5549 gnd.n5548 585
R10946 gnd.n5547 gnd.n5546 585
R10947 gnd.n5545 gnd.n5544 585
R10948 gnd.n5543 gnd.n5542 585
R10949 gnd.n5541 gnd.n5540 585
R10950 gnd.n5539 gnd.n5538 585
R10951 gnd.n5537 gnd.n5536 585
R10952 gnd.n5535 gnd.n5534 585
R10953 gnd.n5532 gnd.n5531 585
R10954 gnd.n5530 gnd.n5529 585
R10955 gnd.n5528 gnd.n5527 585
R10956 gnd.n5526 gnd.n5525 585
R10957 gnd.n5524 gnd.n5523 585
R10958 gnd.n5522 gnd.n5521 585
R10959 gnd.n5520 gnd.n5519 585
R10960 gnd.n5518 gnd.n5517 585
R10961 gnd.n5516 gnd.n5515 585
R10962 gnd.n5514 gnd.n5513 585
R10963 gnd.n5512 gnd.n5511 585
R10964 gnd.n5510 gnd.n5509 585
R10965 gnd.n5508 gnd.n5507 585
R10966 gnd.n5506 gnd.n5505 585
R10967 gnd.n5504 gnd.n5503 585
R10968 gnd.n5502 gnd.n5501 585
R10969 gnd.n5500 gnd.n5499 585
R10970 gnd.n5498 gnd.n5497 585
R10971 gnd.n5496 gnd.n5495 585
R10972 gnd.n5494 gnd.n5493 585
R10973 gnd.n5492 gnd.n5491 585
R10974 gnd.n5490 gnd.n5489 585
R10975 gnd.n5488 gnd.n5487 585
R10976 gnd.n5486 gnd.n5485 585
R10977 gnd.n5484 gnd.n5483 585
R10978 gnd.n5482 gnd.n5481 585
R10979 gnd.n5480 gnd.n5479 585
R10980 gnd.n5478 gnd.n5477 585
R10981 gnd.n5476 gnd.n5475 585
R10982 gnd.n5474 gnd.n5473 585
R10983 gnd.n5468 gnd.n5467 585
R10984 gnd.n7064 gnd.n7063 585
R10985 gnd.n7070 gnd.n7069 585
R10986 gnd.n7072 gnd.n7071 585
R10987 gnd.n7074 gnd.n7073 585
R10988 gnd.n7076 gnd.n7075 585
R10989 gnd.n7078 gnd.n7077 585
R10990 gnd.n7080 gnd.n7079 585
R10991 gnd.n7082 gnd.n7081 585
R10992 gnd.n7084 gnd.n7083 585
R10993 gnd.n7086 gnd.n7085 585
R10994 gnd.n7088 gnd.n7087 585
R10995 gnd.n7090 gnd.n7089 585
R10996 gnd.n7092 gnd.n7091 585
R10997 gnd.n7094 gnd.n7093 585
R10998 gnd.n7096 gnd.n7095 585
R10999 gnd.n7098 gnd.n7097 585
R11000 gnd.n7100 gnd.n7099 585
R11001 gnd.n7102 gnd.n7101 585
R11002 gnd.n7104 gnd.n7103 585
R11003 gnd.n7107 gnd.n7106 585
R11004 gnd.n7105 gnd.n7043 585
R11005 gnd.n7112 gnd.n7111 585
R11006 gnd.n7114 gnd.n7113 585
R11007 gnd.n7116 gnd.n7115 585
R11008 gnd.n7118 gnd.n7117 585
R11009 gnd.n7120 gnd.n7119 585
R11010 gnd.n7122 gnd.n7121 585
R11011 gnd.n7124 gnd.n7123 585
R11012 gnd.n7126 gnd.n7125 585
R11013 gnd.n7128 gnd.n7127 585
R11014 gnd.n7130 gnd.n7129 585
R11015 gnd.n7132 gnd.n7131 585
R11016 gnd.n7134 gnd.n7133 585
R11017 gnd.n7136 gnd.n7135 585
R11018 gnd.n7138 gnd.n7137 585
R11019 gnd.n7140 gnd.n7139 585
R11020 gnd.n7142 gnd.n7141 585
R11021 gnd.n7144 gnd.n7143 585
R11022 gnd.n7146 gnd.n7145 585
R11023 gnd.n7148 gnd.n7147 585
R11024 gnd.n7150 gnd.n7149 585
R11025 gnd.n7155 gnd.n7154 585
R11026 gnd.n7157 gnd.n7156 585
R11027 gnd.n7159 gnd.n7158 585
R11028 gnd.n7161 gnd.n7160 585
R11029 gnd.n7163 gnd.n7162 585
R11030 gnd.n7165 gnd.n7164 585
R11031 gnd.n7167 gnd.n7166 585
R11032 gnd.n7169 gnd.n7168 585
R11033 gnd.n7171 gnd.n7170 585
R11034 gnd.n7173 gnd.n7172 585
R11035 gnd.n7175 gnd.n7174 585
R11036 gnd.n7177 gnd.n7176 585
R11037 gnd.n7179 gnd.n7178 585
R11038 gnd.n7181 gnd.n7180 585
R11039 gnd.n7182 gnd.n7003 585
R11040 gnd.n7184 gnd.n7183 585
R11041 gnd.n7004 gnd.n7002 585
R11042 gnd.n7005 gnd.n166 585
R11043 gnd.n7186 gnd.n166 585
R11044 gnd.n7243 gnd.n168 585
R11045 gnd.n7247 gnd.n168 585
R11046 gnd.n7242 gnd.n7241 585
R11047 gnd.n7241 gnd.n167 585
R11048 gnd.n7240 gnd.n159 585
R11049 gnd.n7253 gnd.n159 585
R11050 gnd.n7239 gnd.n7238 585
R11051 gnd.n7238 gnd.n152 585
R11052 gnd.n7237 gnd.n150 585
R11053 gnd.n7259 gnd.n150 585
R11054 gnd.n7236 gnd.n7235 585
R11055 gnd.n7235 gnd.n142 585
R11056 gnd.n7233 gnd.n140 585
R11057 gnd.n7265 gnd.n140 585
R11058 gnd.n7232 gnd.n7231 585
R11059 gnd.n7231 gnd.n133 585
R11060 gnd.n7230 gnd.n131 585
R11061 gnd.n7271 gnd.n131 585
R11062 gnd.n7229 gnd.n7228 585
R11063 gnd.n7228 gnd.n130 585
R11064 gnd.n7226 gnd.n121 585
R11065 gnd.n7277 gnd.n121 585
R11066 gnd.n7225 gnd.n7224 585
R11067 gnd.n7224 gnd.n120 585
R11068 gnd.n7223 gnd.n112 585
R11069 gnd.n7283 gnd.n112 585
R11070 gnd.n7222 gnd.n7221 585
R11071 gnd.n7221 gnd.n111 585
R11072 gnd.n7219 gnd.n102 585
R11073 gnd.n7289 gnd.n102 585
R11074 gnd.n7218 gnd.n7217 585
R11075 gnd.n7217 gnd.n7216 585
R11076 gnd.n174 gnd.n91 585
R11077 gnd.n7295 gnd.n91 585
R11078 gnd.n6890 gnd.n6889 585
R11079 gnd.n6891 gnd.n6890 585
R11080 gnd.n178 gnd.n177 585
R11081 gnd.n6884 gnd.n177 585
R11082 gnd.n5390 gnd.n74 585
R11083 gnd.n7303 gnd.n74 585
R11084 gnd.n5391 gnd.n1604 585
R11085 gnd.n5395 gnd.n1604 585
R11086 gnd.n5389 gnd.n5388 585
R11087 gnd.n5388 gnd.n1603 585
R11088 gnd.n5387 gnd.n1608 585
R11089 gnd.n5387 gnd.n5386 585
R11090 gnd.n5381 gnd.n1592 585
R11091 gnd.n5404 gnd.n1592 585
R11092 gnd.n5380 gnd.n1586 585
R11093 gnd.n5409 gnd.n1586 585
R11094 gnd.n5379 gnd.n5378 585
R11095 gnd.n5378 gnd.n5377 585
R11096 gnd.n1612 gnd.n1576 585
R11097 gnd.n5415 gnd.n1576 585
R11098 gnd.n5364 gnd.n5363 585
R11099 gnd.n5365 gnd.n5364 585
R11100 gnd.n5361 gnd.n1569 585
R11101 gnd.n5421 gnd.n1569 585
R11102 gnd.n5360 gnd.n5359 585
R11103 gnd.n5359 gnd.n5358 585
R11104 gnd.n1618 gnd.n1559 585
R11105 gnd.n5427 gnd.n1559 585
R11106 gnd.n5286 gnd.n1622 585
R11107 gnd.n5350 gnd.n1622 585
R11108 gnd.n5287 gnd.n1549 585
R11109 gnd.n5433 gnd.n1549 585
R11110 gnd.n5289 gnd.n5288 585
R11111 gnd.n5290 gnd.n5289 585
R11112 gnd.n5284 gnd.n1539 585
R11113 gnd.n5439 gnd.n1539 585
R11114 gnd.n5283 gnd.n5282 585
R11115 gnd.n5282 gnd.n5281 585
R11116 gnd.n5278 gnd.n1529 585
R11117 gnd.n5445 gnd.n1529 585
R11118 gnd.n5277 gnd.n5276 585
R11119 gnd.n5276 gnd.n5275 585
R11120 gnd.n5274 gnd.n1516 585
R11121 gnd.n5451 gnd.n1516 585
R11122 gnd.n1500 gnd.n1499 585
R11123 gnd.n5268 gnd.n1500 585
R11124 gnd.n5459 gnd.n5458 585
R11125 gnd.n5458 gnd.n5457 585
R11126 gnd.n5460 gnd.n1489 585
R11127 gnd.n5307 gnd.n1489 585
R11128 gnd.n5466 gnd.n1490 585
R11129 gnd.n5466 gnd.n5465 585
R11130 gnd.n6072 gnd.n727 585
R11131 gnd.n2170 gnd.n727 585
R11132 gnd.n6876 gnd.n6875 585
R11133 gnd.n6876 gnd.n104 585
R11134 gnd.n6878 gnd.n6877 585
R11135 gnd.n6877 gnd.n93 585
R11136 gnd.n6879 gnd.n182 585
R11137 gnd.n182 gnd.n90 585
R11138 gnd.n6882 gnd.n6881 585
R11139 gnd.n6883 gnd.n6882 585
R11140 gnd.n183 gnd.n181 585
R11141 gnd.n181 gnd.n75 585
R11142 gnd.n1599 gnd.n1598 585
R11143 gnd.n1599 gnd.n73 585
R11144 gnd.n5398 gnd.n5397 585
R11145 gnd.n5397 gnd.n5396 585
R11146 gnd.n5400 gnd.n1595 585
R11147 gnd.n1611 gnd.n1595 585
R11148 gnd.n5402 gnd.n5401 585
R11149 gnd.n5403 gnd.n5402 585
R11150 gnd.n5336 gnd.n1594 585
R11151 gnd.n1594 gnd.n1588 585
R11152 gnd.n5338 gnd.n5337 585
R11153 gnd.n5337 gnd.n1585 585
R11154 gnd.n5340 gnd.n5333 585
R11155 gnd.n5333 gnd.n1578 585
R11156 gnd.n5342 gnd.n5341 585
R11157 gnd.n5342 gnd.n1575 585
R11158 gnd.n5343 gnd.n5332 585
R11159 gnd.n5343 gnd.n1617 585
R11160 gnd.n5345 gnd.n5344 585
R11161 gnd.n5344 gnd.n1568 585
R11162 gnd.n5346 gnd.n1624 585
R11163 gnd.n1624 gnd.n1561 585
R11164 gnd.n5348 gnd.n5347 585
R11165 gnd.n5349 gnd.n5348 585
R11166 gnd.n1625 gnd.n1623 585
R11167 gnd.n1623 gnd.n1551 585
R11168 gnd.n5326 gnd.n5325 585
R11169 gnd.n5325 gnd.n1548 585
R11170 gnd.n5324 gnd.n1627 585
R11171 gnd.n5324 gnd.n1541 585
R11172 gnd.n5323 gnd.n5322 585
R11173 gnd.n5323 gnd.n1538 585
R11174 gnd.n1629 gnd.n1628 585
R11175 gnd.n5280 gnd.n1628 585
R11176 gnd.n5318 gnd.n5317 585
R11177 gnd.n5317 gnd.n1528 585
R11178 gnd.n5316 gnd.n1631 585
R11179 gnd.n5316 gnd.n1518 585
R11180 gnd.n5315 gnd.n5314 585
R11181 gnd.n5315 gnd.n1515 585
R11182 gnd.n1633 gnd.n1632 585
R11183 gnd.n1632 gnd.n1502 585
R11184 gnd.n5310 gnd.n5309 585
R11185 gnd.n5309 gnd.n5308 585
R11186 gnd.n1636 gnd.n1635 585
R11187 gnd.n1636 gnd.n1493 585
R11188 gnd.n5251 gnd.n5250 585
R11189 gnd.n5251 gnd.n1491 585
R11190 gnd.n5252 gnd.n5247 585
R11191 gnd.n5252 gnd.n1423 585
R11192 gnd.n5254 gnd.n5253 585
R11193 gnd.n5253 gnd.n1381 585
R11194 gnd.n5255 gnd.n1668 585
R11195 gnd.n1668 gnd.n1666 585
R11196 gnd.n5257 gnd.n5256 585
R11197 gnd.n5258 gnd.n5257 585
R11198 gnd.n1669 gnd.n1667 585
R11199 gnd.n1667 gnd.n1314 585
R11200 gnd.n5241 gnd.n1313 585
R11201 gnd.n5654 gnd.n1313 585
R11202 gnd.n5240 gnd.n5239 585
R11203 gnd.n5239 gnd.n1312 585
R11204 gnd.n5238 gnd.n1671 585
R11205 gnd.n5238 gnd.n5237 585
R11206 gnd.n5225 gnd.n1672 585
R11207 gnd.n1673 gnd.n1672 585
R11208 gnd.n5227 gnd.n5226 585
R11209 gnd.n5228 gnd.n5227 585
R11210 gnd.n1681 gnd.n1680 585
R11211 gnd.n1680 gnd.n1679 585
R11212 gnd.n5219 gnd.n5218 585
R11213 gnd.n5218 gnd.n5217 585
R11214 gnd.n1684 gnd.n1683 585
R11215 gnd.n1691 gnd.n1684 585
R11216 gnd.n5207 gnd.n5206 585
R11217 gnd.n5208 gnd.n5207 585
R11218 gnd.n1693 gnd.n1692 585
R11219 gnd.n1692 gnd.n1690 585
R11220 gnd.n5202 gnd.n5201 585
R11221 gnd.n5201 gnd.n5200 585
R11222 gnd.n1696 gnd.n1695 585
R11223 gnd.n1697 gnd.n1696 585
R11224 gnd.n5190 gnd.n5189 585
R11225 gnd.n5191 gnd.n5190 585
R11226 gnd.n1705 gnd.n1704 585
R11227 gnd.n1704 gnd.n1703 585
R11228 gnd.n5185 gnd.n5184 585
R11229 gnd.n5184 gnd.n5183 585
R11230 gnd.n1708 gnd.n1707 585
R11231 gnd.n1709 gnd.n1708 585
R11232 gnd.n5173 gnd.n5172 585
R11233 gnd.n5174 gnd.n5173 585
R11234 gnd.n1717 gnd.n1716 585
R11235 gnd.n1716 gnd.n1715 585
R11236 gnd.n5168 gnd.n5167 585
R11237 gnd.n5167 gnd.n5166 585
R11238 gnd.n1720 gnd.n1719 585
R11239 gnd.n1721 gnd.n1720 585
R11240 gnd.n5156 gnd.n5155 585
R11241 gnd.n5157 gnd.n5156 585
R11242 gnd.n1728 gnd.n1727 585
R11243 gnd.n1751 gnd.n1727 585
R11244 gnd.n5151 gnd.n5150 585
R11245 gnd.n5150 gnd.n5149 585
R11246 gnd.n1731 gnd.n1730 585
R11247 gnd.n4946 gnd.n1731 585
R11248 gnd.n4980 gnd.n1783 585
R11249 gnd.n1783 gnd.n1774 585
R11250 gnd.n4982 gnd.n4981 585
R11251 gnd.n4983 gnd.n4982 585
R11252 gnd.n1784 gnd.n1782 585
R11253 gnd.n4958 gnd.n1782 585
R11254 gnd.n4975 gnd.n4974 585
R11255 gnd.n4974 gnd.n4973 585
R11256 gnd.n1787 gnd.n1786 585
R11257 gnd.n1794 gnd.n1787 585
R11258 gnd.n4937 gnd.n4936 585
R11259 gnd.n4938 gnd.n4937 585
R11260 gnd.n1808 gnd.n1807 585
R11261 gnd.n1816 gnd.n1807 585
R11262 gnd.n4932 gnd.n4931 585
R11263 gnd.n4931 gnd.n4930 585
R11264 gnd.n1811 gnd.n1810 585
R11265 gnd.n1821 gnd.n1811 585
R11266 gnd.n4897 gnd.n1837 585
R11267 gnd.n1837 gnd.n1827 585
R11268 gnd.n4899 gnd.n4898 585
R11269 gnd.n4900 gnd.n4899 585
R11270 gnd.n1838 gnd.n1836 585
R11271 gnd.n1836 gnd.n1831 585
R11272 gnd.n4892 gnd.n4891 585
R11273 gnd.n4891 gnd.n4890 585
R11274 gnd.n1841 gnd.n1840 585
R11275 gnd.n4883 gnd.n1841 585
R11276 gnd.n4856 gnd.n1859 585
R11277 gnd.n4840 gnd.n1859 585
R11278 gnd.n4858 gnd.n4857 585
R11279 gnd.n4859 gnd.n4858 585
R11280 gnd.n1860 gnd.n1858 585
R11281 gnd.n1867 gnd.n1858 585
R11282 gnd.n4851 gnd.n4850 585
R11283 gnd.n4850 gnd.n4849 585
R11284 gnd.n1863 gnd.n1862 585
R11285 gnd.n4820 gnd.n1863 585
R11286 gnd.n4807 gnd.n1886 585
R11287 gnd.n4790 gnd.n1886 585
R11288 gnd.n4809 gnd.n4808 585
R11289 gnd.n4810 gnd.n4809 585
R11290 gnd.n1887 gnd.n1885 585
R11291 gnd.n1894 gnd.n1885 585
R11292 gnd.n4802 gnd.n4801 585
R11293 gnd.n4801 gnd.n4800 585
R11294 gnd.n1890 gnd.n1889 585
R11295 gnd.n1905 gnd.n1890 585
R11296 gnd.n4770 gnd.n4769 585
R11297 gnd.n4771 gnd.n4770 585
R11298 gnd.n1913 gnd.n1912 585
R11299 gnd.n1920 gnd.n1912 585
R11300 gnd.n4765 gnd.n4764 585
R11301 gnd.n4764 gnd.n4763 585
R11302 gnd.n1916 gnd.n1915 585
R11303 gnd.n1924 gnd.n1916 585
R11304 gnd.n4732 gnd.n1940 585
R11305 gnd.n1940 gnd.n1930 585
R11306 gnd.n4734 gnd.n4733 585
R11307 gnd.n4735 gnd.n4734 585
R11308 gnd.n1941 gnd.n1939 585
R11309 gnd.n1939 gnd.n1935 585
R11310 gnd.n4727 gnd.n4726 585
R11311 gnd.n4726 gnd.n4725 585
R11312 gnd.n1944 gnd.n1943 585
R11313 gnd.n4717 gnd.n1944 585
R11314 gnd.n4695 gnd.n4694 585
R11315 gnd.n4694 gnd.n4693 585
R11316 gnd.n4696 gnd.n1964 585
R11317 gnd.n1970 gnd.n1964 585
R11318 gnd.n4698 gnd.n4697 585
R11319 gnd.n4699 gnd.n4698 585
R11320 gnd.n1965 gnd.n1963 585
R11321 gnd.n4658 gnd.n1963 585
R11322 gnd.n4634 gnd.n4633 585
R11323 gnd.n4633 gnd.n1977 585
R11324 gnd.n4635 gnd.n1990 585
R11325 gnd.n1990 gnd.n1983 585
R11326 gnd.n4637 gnd.n4636 585
R11327 gnd.n4638 gnd.n4637 585
R11328 gnd.n1991 gnd.n1989 585
R11329 gnd.n1997 gnd.n1989 585
R11330 gnd.n4626 gnd.n4625 585
R11331 gnd.n4625 gnd.n4624 585
R11332 gnd.n1994 gnd.n1993 585
R11333 gnd.n2003 gnd.n1994 585
R11334 gnd.n4593 gnd.n2018 585
R11335 gnd.n2018 gnd.n2009 585
R11336 gnd.n4595 gnd.n4594 585
R11337 gnd.n4596 gnd.n4595 585
R11338 gnd.n2019 gnd.n2017 585
R11339 gnd.n2017 gnd.n2013 585
R11340 gnd.n4588 gnd.n4587 585
R11341 gnd.n4587 gnd.n4586 585
R11342 gnd.n2022 gnd.n2021 585
R11343 gnd.n4577 gnd.n2022 585
R11344 gnd.n4564 gnd.n4563 585
R11345 gnd.n4565 gnd.n4564 585
R11346 gnd.n4559 gnd.n4558 585
R11347 gnd.n4558 gnd.n4557 585
R11348 gnd.n1212 gnd.n1211 585
R11349 gnd.n4501 gnd.n1212 585
R11350 gnd.n5773 gnd.n5772 585
R11351 gnd.n5772 gnd.n5771 585
R11352 gnd.n5774 gnd.n1206 585
R11353 gnd.n4521 gnd.n1206 585
R11354 gnd.n5776 gnd.n5775 585
R11355 gnd.n5777 gnd.n5776 585
R11356 gnd.n1207 gnd.n1205 585
R11357 gnd.n1205 gnd.n1201 585
R11358 gnd.n4409 gnd.n4408 585
R11359 gnd.n4408 gnd.n1175 585
R11360 gnd.n4410 gnd.n2048 585
R11361 gnd.n2048 gnd.n1143 585
R11362 gnd.n4412 gnd.n4411 585
R11363 gnd.n4413 gnd.n4412 585
R11364 gnd.n2049 gnd.n2047 585
R11365 gnd.n2047 gnd.n2045 585
R11366 gnd.n4401 gnd.n4400 585
R11367 gnd.n4400 gnd.n4399 585
R11368 gnd.n2052 gnd.n2051 585
R11369 gnd.n2053 gnd.n2052 585
R11370 gnd.n4376 gnd.n4375 585
R11371 gnd.n4377 gnd.n4376 585
R11372 gnd.n2064 gnd.n2063 585
R11373 gnd.n2070 gnd.n2063 585
R11374 gnd.n4371 gnd.n4370 585
R11375 gnd.n4370 gnd.n4369 585
R11376 gnd.n2067 gnd.n2066 585
R11377 gnd.n2068 gnd.n2067 585
R11378 gnd.n4360 gnd.n4359 585
R11379 gnd.n4361 gnd.n4360 585
R11380 gnd.n2078 gnd.n2077 585
R11381 gnd.n2084 gnd.n2077 585
R11382 gnd.n4355 gnd.n4354 585
R11383 gnd.n4354 gnd.n4353 585
R11384 gnd.n2081 gnd.n2080 585
R11385 gnd.n2082 gnd.n2081 585
R11386 gnd.n4344 gnd.n4343 585
R11387 gnd.n4345 gnd.n4344 585
R11388 gnd.n2093 gnd.n2092 585
R11389 gnd.n2092 gnd.n2090 585
R11390 gnd.n4339 gnd.n4338 585
R11391 gnd.n4338 gnd.n4337 585
R11392 gnd.n2096 gnd.n2095 585
R11393 gnd.n2097 gnd.n2096 585
R11394 gnd.n4328 gnd.n4327 585
R11395 gnd.n4329 gnd.n4328 585
R11396 gnd.n2107 gnd.n2106 585
R11397 gnd.n2106 gnd.n2104 585
R11398 gnd.n4323 gnd.n4322 585
R11399 gnd.n4322 gnd.n4321 585
R11400 gnd.n2110 gnd.n2109 585
R11401 gnd.n4312 gnd.n2110 585
R11402 gnd.n4260 gnd.n4259 585
R11403 gnd.n4261 gnd.n4260 585
R11404 gnd.n2113 gnd.n2112 585
R11405 gnd.n2112 gnd.n890 585
R11406 gnd.n4255 gnd.n4254 585
R11407 gnd.n4254 gnd.n876 585
R11408 gnd.n4253 gnd.n2115 585
R11409 gnd.n4253 gnd.n4252 585
R11410 gnd.n4251 gnd.n4250 585
R11411 gnd.n4251 gnd.n979 585
R11412 gnd.n2117 gnd.n2116 585
R11413 gnd.n2116 gnd.n965 585
R11414 gnd.n4246 gnd.n4245 585
R11415 gnd.n4245 gnd.n862 585
R11416 gnd.n4244 gnd.n2119 585
R11417 gnd.n4244 gnd.n859 585
R11418 gnd.n4243 gnd.n4242 585
R11419 gnd.n4243 gnd.n867 585
R11420 gnd.n2121 gnd.n2120 585
R11421 gnd.n2120 gnd.n850 585
R11422 gnd.n4238 gnd.n4237 585
R11423 gnd.n4237 gnd.n843 585
R11424 gnd.n4236 gnd.n2123 585
R11425 gnd.n4236 gnd.n840 585
R11426 gnd.n4235 gnd.n4234 585
R11427 gnd.n4235 gnd.n832 585
R11428 gnd.n2125 gnd.n2124 585
R11429 gnd.n4190 gnd.n2124 585
R11430 gnd.n4230 gnd.n4229 585
R11431 gnd.n4229 gnd.n823 585
R11432 gnd.n4228 gnd.n2127 585
R11433 gnd.n4228 gnd.n820 585
R11434 gnd.n4227 gnd.n4226 585
R11435 gnd.n4227 gnd.n812 585
R11436 gnd.n2129 gnd.n2128 585
R11437 gnd.n2128 gnd.n809 585
R11438 gnd.n4222 gnd.n4221 585
R11439 gnd.n4221 gnd.n4220 585
R11440 gnd.n2132 gnd.n2131 585
R11441 gnd.n2132 gnd.n800 585
R11442 gnd.n4167 gnd.n2150 585
R11443 gnd.n2150 gnd.n792 585
R11444 gnd.n4169 gnd.n4168 585
R11445 gnd.n4170 gnd.n4169 585
R11446 gnd.n4163 gnd.n2149 585
R11447 gnd.n2149 gnd.n783 585
R11448 gnd.n4162 gnd.n4161 585
R11449 gnd.n4161 gnd.n780 585
R11450 gnd.n4160 gnd.n4159 585
R11451 gnd.n4160 gnd.n775 585
R11452 gnd.n4158 gnd.n2152 585
R11453 gnd.n2152 gnd.n772 585
R11454 gnd.n4156 gnd.n4155 585
R11455 gnd.n4155 gnd.n4154 585
R11456 gnd.n2154 gnd.n2153 585
R11457 gnd.n2154 gnd.n763 585
R11458 gnd.n4122 gnd.n4115 585
R11459 gnd.n4115 gnd.n758 585
R11460 gnd.n4124 gnd.n4123 585
R11461 gnd.n4125 gnd.n4124 585
R11462 gnd.n4119 gnd.n4114 585
R11463 gnd.n4114 gnd.n747 585
R11464 gnd.n4118 gnd.n4117 585
R11465 gnd.n4117 gnd.n744 585
R11466 gnd.n732 gnd.n731 585
R11467 gnd.n736 gnd.n732 585
R11468 gnd.n6069 gnd.n6068 585
R11469 gnd.n6068 gnd.n6067 585
R11470 gnd.n5653 gnd.n5652 585
R11471 gnd.n5654 gnd.n5653 585
R11472 gnd.n1317 gnd.n1315 585
R11473 gnd.n1315 gnd.n1312 585
R11474 gnd.n5235 gnd.n5234 585
R11475 gnd.n5237 gnd.n5235 585
R11476 gnd.n1675 gnd.n1674 585
R11477 gnd.n1674 gnd.n1673 585
R11478 gnd.n5230 gnd.n5229 585
R11479 gnd.n5229 gnd.n5228 585
R11480 gnd.n1678 gnd.n1677 585
R11481 gnd.n1679 gnd.n1678 585
R11482 gnd.n5215 gnd.n5214 585
R11483 gnd.n5217 gnd.n5215 585
R11484 gnd.n1686 gnd.n1685 585
R11485 gnd.n1691 gnd.n1685 585
R11486 gnd.n5210 gnd.n5209 585
R11487 gnd.n5209 gnd.n5208 585
R11488 gnd.n1689 gnd.n1688 585
R11489 gnd.n1690 gnd.n1689 585
R11490 gnd.n5198 gnd.n5197 585
R11491 gnd.n5200 gnd.n5198 585
R11492 gnd.n1699 gnd.n1698 585
R11493 gnd.n1698 gnd.n1697 585
R11494 gnd.n5193 gnd.n5192 585
R11495 gnd.n5192 gnd.n5191 585
R11496 gnd.n1702 gnd.n1701 585
R11497 gnd.n1703 gnd.n1702 585
R11498 gnd.n5181 gnd.n5180 585
R11499 gnd.n5183 gnd.n5181 585
R11500 gnd.n1711 gnd.n1710 585
R11501 gnd.n1710 gnd.n1709 585
R11502 gnd.n5176 gnd.n5175 585
R11503 gnd.n5175 gnd.n5174 585
R11504 gnd.n1714 gnd.n1713 585
R11505 gnd.n1715 gnd.n1714 585
R11506 gnd.n5164 gnd.n5163 585
R11507 gnd.n5166 gnd.n5164 585
R11508 gnd.n1723 gnd.n1722 585
R11509 gnd.n1722 gnd.n1721 585
R11510 gnd.n5159 gnd.n5158 585
R11511 gnd.n5158 gnd.n5157 585
R11512 gnd.n1726 gnd.n1725 585
R11513 gnd.n1751 gnd.n1726 585
R11514 gnd.n4949 gnd.n1733 585
R11515 gnd.n5149 gnd.n1733 585
R11516 gnd.n4950 gnd.n4947 585
R11517 gnd.n4947 gnd.n4946 585
R11518 gnd.n4951 gnd.n4945 585
R11519 gnd.n4945 gnd.n1774 585
R11520 gnd.n1801 gnd.n1779 585
R11521 gnd.n4983 gnd.n1779 585
R11522 gnd.n4956 gnd.n4955 585
R11523 gnd.n4958 gnd.n4956 585
R11524 gnd.n1800 gnd.n1789 585
R11525 gnd.n4973 gnd.n1789 585
R11526 gnd.n4941 gnd.n4940 585
R11527 gnd.n4940 gnd.n1794 585
R11528 gnd.n4939 gnd.n1803 585
R11529 gnd.n4939 gnd.n4938 585
R11530 gnd.n4870 gnd.n1804 585
R11531 gnd.n1816 gnd.n1804 585
R11532 gnd.n4871 gnd.n1813 585
R11533 gnd.n4930 gnd.n1813 585
R11534 gnd.n4868 gnd.n4867 585
R11535 gnd.n4867 gnd.n1821 585
R11536 gnd.n4875 gnd.n4866 585
R11537 gnd.n4866 gnd.n1827 585
R11538 gnd.n4876 gnd.n1833 585
R11539 gnd.n4900 gnd.n1833 585
R11540 gnd.n4877 gnd.n4865 585
R11541 gnd.n4865 gnd.n1831 585
R11542 gnd.n1853 gnd.n1843 585
R11543 gnd.n4890 gnd.n1843 585
R11544 gnd.n4882 gnd.n4881 585
R11545 gnd.n4883 gnd.n4882 585
R11546 gnd.n1852 gnd.n1851 585
R11547 gnd.n4840 gnd.n1851 585
R11548 gnd.n4861 gnd.n4860 585
R11549 gnd.n4860 gnd.n4859 585
R11550 gnd.n1856 gnd.n1855 585
R11551 gnd.n1867 gnd.n1856 585
R11552 gnd.n1880 gnd.n1865 585
R11553 gnd.n4849 gnd.n1865 585
R11554 gnd.n4818 gnd.n4817 585
R11555 gnd.n4820 gnd.n4818 585
R11556 gnd.n1879 gnd.n1878 585
R11557 gnd.n4790 gnd.n1878 585
R11558 gnd.n4812 gnd.n4811 585
R11559 gnd.n4811 gnd.n4810 585
R11560 gnd.n1883 gnd.n1882 585
R11561 gnd.n1894 gnd.n1883 585
R11562 gnd.n4674 gnd.n1892 585
R11563 gnd.n4800 gnd.n1892 585
R11564 gnd.n4675 gnd.n4673 585
R11565 gnd.n4673 gnd.n1905 585
R11566 gnd.n4671 gnd.n1910 585
R11567 gnd.n4771 gnd.n1910 585
R11568 gnd.n4679 gnd.n4670 585
R11569 gnd.n4670 gnd.n1920 585
R11570 gnd.n4680 gnd.n1918 585
R11571 gnd.n4763 gnd.n1918 585
R11572 gnd.n4681 gnd.n4669 585
R11573 gnd.n4669 gnd.n1924 585
R11574 gnd.n4668 gnd.n4666 585
R11575 gnd.n4668 gnd.n1930 585
R11576 gnd.n4685 gnd.n1937 585
R11577 gnd.n4735 gnd.n1937 585
R11578 gnd.n4686 gnd.n4665 585
R11579 gnd.n4665 gnd.n1935 585
R11580 gnd.n4687 gnd.n1945 585
R11581 gnd.n4725 gnd.n1945 585
R11582 gnd.n1973 gnd.n1953 585
R11583 gnd.n4717 gnd.n1953 585
R11584 gnd.n4692 gnd.n4691 585
R11585 gnd.n4693 gnd.n4692 585
R11586 gnd.n1972 gnd.n1971 585
R11587 gnd.n1971 gnd.n1970 585
R11588 gnd.n4661 gnd.n1960 585
R11589 gnd.n4699 gnd.n1960 585
R11590 gnd.n4660 gnd.n4659 585
R11591 gnd.n4659 gnd.n4658 585
R11592 gnd.n1976 gnd.n1975 585
R11593 gnd.n1977 gnd.n1976 585
R11594 gnd.n4538 gnd.n4537 585
R11595 gnd.n4537 gnd.n1983 585
R11596 gnd.n4539 gnd.n1988 585
R11597 gnd.n4638 gnd.n1988 585
R11598 gnd.n4534 gnd.n4533 585
R11599 gnd.n4533 gnd.n1997 585
R11600 gnd.n4543 gnd.n1995 585
R11601 gnd.n4624 gnd.n1995 585
R11602 gnd.n4544 gnd.n4532 585
R11603 gnd.n4532 gnd.n2003 585
R11604 gnd.n4545 gnd.n4531 585
R11605 gnd.n4531 gnd.n2009 585
R11606 gnd.n4529 gnd.n2015 585
R11607 gnd.n4596 gnd.n2015 585
R11608 gnd.n4549 gnd.n4528 585
R11609 gnd.n4528 gnd.n2013 585
R11610 gnd.n4550 gnd.n2023 585
R11611 gnd.n4586 gnd.n2023 585
R11612 gnd.n4551 gnd.n2030 585
R11613 gnd.n4577 gnd.n2030 585
R11614 gnd.n2038 gnd.n2034 585
R11615 gnd.n4565 gnd.n2034 585
R11616 gnd.n4556 gnd.n4555 585
R11617 gnd.n4557 gnd.n4556 585
R11618 gnd.n2037 gnd.n2036 585
R11619 gnd.n4501 gnd.n2036 585
R11620 gnd.n4524 gnd.n1213 585
R11621 gnd.n5771 gnd.n1213 585
R11622 gnd.n4523 gnd.n4522 585
R11623 gnd.n4522 gnd.n4521 585
R11624 gnd.n4422 gnd.n1203 585
R11625 gnd.n5777 gnd.n1203 585
R11626 gnd.n4416 gnd.n2040 585
R11627 gnd.n4416 gnd.n1201 585
R11628 gnd.n4418 gnd.n4417 585
R11629 gnd.n4417 gnd.n1175 585
R11630 gnd.n4415 gnd.n2042 585
R11631 gnd.n4415 gnd.n1143 585
R11632 gnd.n4414 gnd.n2044 585
R11633 gnd.n4414 gnd.n4413 585
R11634 gnd.n4282 gnd.n2043 585
R11635 gnd.n2045 gnd.n2043 585
R11636 gnd.n4280 gnd.n2054 585
R11637 gnd.n4399 gnd.n2054 585
R11638 gnd.n4286 gnd.n4279 585
R11639 gnd.n4279 gnd.n2053 585
R11640 gnd.n4287 gnd.n2062 585
R11641 gnd.n4377 gnd.n2062 585
R11642 gnd.n4288 gnd.n4278 585
R11643 gnd.n4278 gnd.n2070 585
R11644 gnd.n4276 gnd.n2069 585
R11645 gnd.n4369 gnd.n2069 585
R11646 gnd.n4292 gnd.n4275 585
R11647 gnd.n4275 gnd.n2068 585
R11648 gnd.n4293 gnd.n2076 585
R11649 gnd.n4361 gnd.n2076 585
R11650 gnd.n4294 gnd.n4274 585
R11651 gnd.n4274 gnd.n2084 585
R11652 gnd.n4272 gnd.n2083 585
R11653 gnd.n4353 gnd.n2083 585
R11654 gnd.n4298 gnd.n4271 585
R11655 gnd.n4271 gnd.n2082 585
R11656 gnd.n4299 gnd.n2091 585
R11657 gnd.n4345 gnd.n2091 585
R11658 gnd.n4300 gnd.n4270 585
R11659 gnd.n4270 gnd.n2090 585
R11660 gnd.n4268 gnd.n2098 585
R11661 gnd.n4337 gnd.n2098 585
R11662 gnd.n4304 gnd.n4267 585
R11663 gnd.n4267 gnd.n2097 585
R11664 gnd.n4305 gnd.n2105 585
R11665 gnd.n4329 gnd.n2105 585
R11666 gnd.n4306 gnd.n4266 585
R11667 gnd.n4266 gnd.n2104 585
R11668 gnd.n4263 gnd.n2111 585
R11669 gnd.n4321 gnd.n2111 585
R11670 gnd.n4311 gnd.n4310 585
R11671 gnd.n4312 gnd.n4311 585
R11672 gnd.n4262 gnd.n893 585
R11673 gnd.n4261 gnd.n893 585
R11674 gnd.n5965 gnd.n5964 585
R11675 gnd.n5963 gnd.n892 585
R11676 gnd.n895 gnd.n891 585
R11677 gnd.n5967 gnd.n891 585
R11678 gnd.n5959 gnd.n897 585
R11679 gnd.n5958 gnd.n898 585
R11680 gnd.n5957 gnd.n899 585
R11681 gnd.n902 gnd.n900 585
R11682 gnd.n5952 gnd.n903 585
R11683 gnd.n5951 gnd.n904 585
R11684 gnd.n5950 gnd.n905 585
R11685 gnd.n914 gnd.n906 585
R11686 gnd.n5943 gnd.n915 585
R11687 gnd.n5942 gnd.n916 585
R11688 gnd.n918 gnd.n917 585
R11689 gnd.n5935 gnd.n924 585
R11690 gnd.n5934 gnd.n925 585
R11691 gnd.n932 gnd.n926 585
R11692 gnd.n5927 gnd.n933 585
R11693 gnd.n5926 gnd.n934 585
R11694 gnd.n936 gnd.n935 585
R11695 gnd.n5919 gnd.n942 585
R11696 gnd.n5918 gnd.n943 585
R11697 gnd.n950 gnd.n944 585
R11698 gnd.n5911 gnd.n951 585
R11699 gnd.n5910 gnd.n952 585
R11700 gnd.n957 gnd.n956 585
R11701 gnd.n888 gnd.n873 585
R11702 gnd.n5971 gnd.n874 585
R11703 gnd.n5970 gnd.n5969 585
R11704 gnd.n5656 gnd.n5655 585
R11705 gnd.n5655 gnd.n5654 585
R11706 gnd.n5657 gnd.n1310 585
R11707 gnd.n1312 gnd.n1310 585
R11708 gnd.n5236 gnd.n1308 585
R11709 gnd.n5237 gnd.n5236 585
R11710 gnd.n5661 gnd.n1307 585
R11711 gnd.n1673 gnd.n1307 585
R11712 gnd.n5662 gnd.n1306 585
R11713 gnd.n5228 gnd.n1306 585
R11714 gnd.n5663 gnd.n1305 585
R11715 gnd.n1679 gnd.n1305 585
R11716 gnd.n5216 gnd.n1303 585
R11717 gnd.n5217 gnd.n5216 585
R11718 gnd.n5667 gnd.n1302 585
R11719 gnd.n1691 gnd.n1302 585
R11720 gnd.n5668 gnd.n1301 585
R11721 gnd.n5208 gnd.n1301 585
R11722 gnd.n5669 gnd.n1300 585
R11723 gnd.n1690 gnd.n1300 585
R11724 gnd.n5199 gnd.n1298 585
R11725 gnd.n5200 gnd.n5199 585
R11726 gnd.n5673 gnd.n1297 585
R11727 gnd.n1697 gnd.n1297 585
R11728 gnd.n5674 gnd.n1296 585
R11729 gnd.n5191 gnd.n1296 585
R11730 gnd.n5675 gnd.n1295 585
R11731 gnd.n1703 gnd.n1295 585
R11732 gnd.n5182 gnd.n1293 585
R11733 gnd.n5183 gnd.n5182 585
R11734 gnd.n5679 gnd.n1292 585
R11735 gnd.n1709 gnd.n1292 585
R11736 gnd.n5680 gnd.n1291 585
R11737 gnd.n5174 gnd.n1291 585
R11738 gnd.n5681 gnd.n1290 585
R11739 gnd.n1715 gnd.n1290 585
R11740 gnd.n5165 gnd.n1288 585
R11741 gnd.n5166 gnd.n5165 585
R11742 gnd.n5685 gnd.n1287 585
R11743 gnd.n1721 gnd.n1287 585
R11744 gnd.n5686 gnd.n1286 585
R11745 gnd.n5157 gnd.n1286 585
R11746 gnd.n5687 gnd.n1285 585
R11747 gnd.n1751 gnd.n1285 585
R11748 gnd.n5148 gnd.n1283 585
R11749 gnd.n5149 gnd.n5148 585
R11750 gnd.n5691 gnd.n1282 585
R11751 gnd.n4946 gnd.n1282 585
R11752 gnd.n5692 gnd.n1281 585
R11753 gnd.n1774 gnd.n1281 585
R11754 gnd.n5693 gnd.n1280 585
R11755 gnd.n4983 gnd.n1280 585
R11756 gnd.n4957 gnd.n1278 585
R11757 gnd.n4958 gnd.n4957 585
R11758 gnd.n5697 gnd.n1277 585
R11759 gnd.n4973 gnd.n1277 585
R11760 gnd.n5698 gnd.n1276 585
R11761 gnd.n1794 gnd.n1276 585
R11762 gnd.n5699 gnd.n1275 585
R11763 gnd.n4938 gnd.n1275 585
R11764 gnd.n1815 gnd.n1273 585
R11765 gnd.n1816 gnd.n1815 585
R11766 gnd.n5703 gnd.n1272 585
R11767 gnd.n4930 gnd.n1272 585
R11768 gnd.n5704 gnd.n1271 585
R11769 gnd.n1821 gnd.n1271 585
R11770 gnd.n5705 gnd.n1270 585
R11771 gnd.n1827 gnd.n1270 585
R11772 gnd.n1835 gnd.n1268 585
R11773 gnd.n4900 gnd.n1835 585
R11774 gnd.n5709 gnd.n1267 585
R11775 gnd.n1831 gnd.n1267 585
R11776 gnd.n5710 gnd.n1266 585
R11777 gnd.n4890 gnd.n1266 585
R11778 gnd.n5711 gnd.n1265 585
R11779 gnd.n4883 gnd.n1265 585
R11780 gnd.n4839 gnd.n1263 585
R11781 gnd.n4840 gnd.n4839 585
R11782 gnd.n5715 gnd.n1262 585
R11783 gnd.n4859 gnd.n1262 585
R11784 gnd.n5716 gnd.n1261 585
R11785 gnd.n1867 gnd.n1261 585
R11786 gnd.n5717 gnd.n1260 585
R11787 gnd.n4849 gnd.n1260 585
R11788 gnd.n4819 gnd.n1258 585
R11789 gnd.n4820 gnd.n4819 585
R11790 gnd.n5721 gnd.n1257 585
R11791 gnd.n4790 gnd.n1257 585
R11792 gnd.n5722 gnd.n1256 585
R11793 gnd.n4810 gnd.n1256 585
R11794 gnd.n5723 gnd.n1255 585
R11795 gnd.n1894 gnd.n1255 585
R11796 gnd.n4799 gnd.n1253 585
R11797 gnd.n4800 gnd.n4799 585
R11798 gnd.n5727 gnd.n1252 585
R11799 gnd.n1905 gnd.n1252 585
R11800 gnd.n5728 gnd.n1251 585
R11801 gnd.n4771 gnd.n1251 585
R11802 gnd.n5729 gnd.n1250 585
R11803 gnd.n1920 gnd.n1250 585
R11804 gnd.n4762 gnd.n1248 585
R11805 gnd.n4763 gnd.n4762 585
R11806 gnd.n5733 gnd.n1247 585
R11807 gnd.n1924 gnd.n1247 585
R11808 gnd.n5734 gnd.n1246 585
R11809 gnd.n1930 gnd.n1246 585
R11810 gnd.n5735 gnd.n1245 585
R11811 gnd.n4735 gnd.n1245 585
R11812 gnd.n1934 gnd.n1243 585
R11813 gnd.n1935 gnd.n1934 585
R11814 gnd.n5739 gnd.n1242 585
R11815 gnd.n4725 gnd.n1242 585
R11816 gnd.n5740 gnd.n1241 585
R11817 gnd.n4717 gnd.n1241 585
R11818 gnd.n5741 gnd.n1240 585
R11819 gnd.n4693 gnd.n1240 585
R11820 gnd.n1969 gnd.n1238 585
R11821 gnd.n1970 gnd.n1969 585
R11822 gnd.n5745 gnd.n1237 585
R11823 gnd.n4699 gnd.n1237 585
R11824 gnd.n5746 gnd.n1236 585
R11825 gnd.n4658 gnd.n1236 585
R11826 gnd.n5747 gnd.n1235 585
R11827 gnd.n1977 gnd.n1235 585
R11828 gnd.n1982 gnd.n1233 585
R11829 gnd.n1983 gnd.n1982 585
R11830 gnd.n5751 gnd.n1232 585
R11831 gnd.n4638 gnd.n1232 585
R11832 gnd.n5752 gnd.n1231 585
R11833 gnd.n1997 gnd.n1231 585
R11834 gnd.n5753 gnd.n1230 585
R11835 gnd.n4624 gnd.n1230 585
R11836 gnd.n2002 gnd.n1228 585
R11837 gnd.n2003 gnd.n2002 585
R11838 gnd.n5757 gnd.n1227 585
R11839 gnd.n2009 gnd.n1227 585
R11840 gnd.n5758 gnd.n1226 585
R11841 gnd.n4596 gnd.n1226 585
R11842 gnd.n5759 gnd.n1225 585
R11843 gnd.n2013 gnd.n1225 585
R11844 gnd.n4585 gnd.n1223 585
R11845 gnd.n4586 gnd.n4585 585
R11846 gnd.n5763 gnd.n1222 585
R11847 gnd.n4577 gnd.n1222 585
R11848 gnd.n5764 gnd.n1221 585
R11849 gnd.n4565 gnd.n1221 585
R11850 gnd.n5765 gnd.n1220 585
R11851 gnd.n4557 gnd.n1220 585
R11852 gnd.n1217 gnd.n1215 585
R11853 gnd.n4501 gnd.n1215 585
R11854 gnd.n5770 gnd.n5769 585
R11855 gnd.n5771 gnd.n5770 585
R11856 gnd.n1216 gnd.n1214 585
R11857 gnd.n4521 gnd.n1214 585
R11858 gnd.n4387 gnd.n1204 585
R11859 gnd.n5777 gnd.n1204 585
R11860 gnd.n4386 gnd.n4385 585
R11861 gnd.n4385 gnd.n1201 585
R11862 gnd.n4391 gnd.n4384 585
R11863 gnd.n4384 gnd.n1175 585
R11864 gnd.n4392 gnd.n4383 585
R11865 gnd.n4383 gnd.n1143 585
R11866 gnd.n4393 gnd.n2046 585
R11867 gnd.n4413 gnd.n2046 585
R11868 gnd.n2058 gnd.n2056 585
R11869 gnd.n2056 gnd.n2045 585
R11870 gnd.n4398 gnd.n4397 585
R11871 gnd.n4399 gnd.n4398 585
R11872 gnd.n2057 gnd.n2055 585
R11873 gnd.n2055 gnd.n2053 585
R11874 gnd.n4379 gnd.n4378 585
R11875 gnd.n4378 gnd.n4377 585
R11876 gnd.n2061 gnd.n2060 585
R11877 gnd.n2070 gnd.n2061 585
R11878 gnd.n4368 gnd.n4367 585
R11879 gnd.n4369 gnd.n4368 585
R11880 gnd.n2072 gnd.n2071 585
R11881 gnd.n2071 gnd.n2068 585
R11882 gnd.n4363 gnd.n4362 585
R11883 gnd.n4362 gnd.n4361 585
R11884 gnd.n2075 gnd.n2074 585
R11885 gnd.n2084 gnd.n2075 585
R11886 gnd.n4352 gnd.n4351 585
R11887 gnd.n4353 gnd.n4352 585
R11888 gnd.n2086 gnd.n2085 585
R11889 gnd.n2085 gnd.n2082 585
R11890 gnd.n4347 gnd.n4346 585
R11891 gnd.n4346 gnd.n4345 585
R11892 gnd.n2089 gnd.n2088 585
R11893 gnd.n2090 gnd.n2089 585
R11894 gnd.n4336 gnd.n4335 585
R11895 gnd.n4337 gnd.n4336 585
R11896 gnd.n2100 gnd.n2099 585
R11897 gnd.n2099 gnd.n2097 585
R11898 gnd.n4331 gnd.n4330 585
R11899 gnd.n4330 gnd.n4329 585
R11900 gnd.n2103 gnd.n2102 585
R11901 gnd.n2104 gnd.n2103 585
R11902 gnd.n4320 gnd.n4319 585
R11903 gnd.n4321 gnd.n4320 585
R11904 gnd.n4314 gnd.n4313 585
R11905 gnd.n4313 gnd.n4312 585
R11906 gnd.n4315 gnd.n875 585
R11907 gnd.n4261 gnd.n875 585
R11908 gnd.n5595 gnd.n1372 585
R11909 gnd.n5259 gnd.n1372 585
R11910 gnd.n5596 gnd.n1371 585
R11911 gnd.n1661 gnd.n1365 585
R11912 gnd.n5603 gnd.n1364 585
R11913 gnd.n5604 gnd.n1363 585
R11914 gnd.n1658 gnd.n1357 585
R11915 gnd.n5611 gnd.n1356 585
R11916 gnd.n5612 gnd.n1355 585
R11917 gnd.n1656 gnd.n1349 585
R11918 gnd.n5619 gnd.n1348 585
R11919 gnd.n5620 gnd.n1347 585
R11920 gnd.n1653 gnd.n1341 585
R11921 gnd.n5627 gnd.n1340 585
R11922 gnd.n5628 gnd.n1339 585
R11923 gnd.n1651 gnd.n1332 585
R11924 gnd.n5635 gnd.n1331 585
R11925 gnd.n5636 gnd.n1330 585
R11926 gnd.n1648 gnd.n1327 585
R11927 gnd.n5641 gnd.n1326 585
R11928 gnd.n5642 gnd.n1325 585
R11929 gnd.n5643 gnd.n1324 585
R11930 gnd.n1645 gnd.n1322 585
R11931 gnd.n5647 gnd.n1321 585
R11932 gnd.n5648 gnd.n1320 585
R11933 gnd.n5649 gnd.n1316 585
R11934 gnd.n5262 gnd.n1311 585
R11935 gnd.n5263 gnd.n5261 585
R11936 gnd.n1643 gnd.n1642 585
R11937 gnd.n1664 gnd.n1663 585
R11938 gnd.n5072 gnd.n1776 511.721
R11939 gnd.n5081 gnd.n5080 511.721
R11940 gnd.n4493 gnd.n4491 511.721
R11941 gnd.n5846 gnd.n1178 511.721
R11942 gnd.n6245 gnd.n561 498.228
R11943 gnd.n4427 gnd.t98 389.64
R11944 gnd.n1769 gnd.t51 389.64
R11945 gnd.n5783 gnd.t22 389.64
R11946 gnd.n5006 gnd.t107 389.64
R11947 gnd.n953 gnd.t63 371.625
R11948 gnd.n5589 gnd.t30 371.625
R11949 gnd.n960 gnd.t59 371.625
R11950 gnd.n1445 gnd.t119 371.625
R11951 gnd.n1468 gnd.t122 371.625
R11952 gnd.n5469 gnd.t83 371.625
R11953 gnd.n7065 gnd.t80 371.625
R11954 gnd.n7044 gnd.t86 371.625
R11955 gnd.n7151 gnd.t104 371.625
R11956 gnd.n6912 gnd.t26 371.625
R11957 gnd.n3808 gnd.t67 371.625
R11958 gnd.n3839 gnd.t101 371.625
R11959 gnd.n3871 gnd.t113 371.625
R11960 gnd.n3708 gnd.t55 371.625
R11961 gnd.n1030 gnd.t95 371.625
R11962 gnd.n1071 gnd.t116 371.625
R11963 gnd.n1050 gnd.t136 371.625
R11964 gnd.n1373 gnd.t44 371.625
R11965 gnd.n2722 gnd.t70 323.425
R11966 gnd.n2280 gnd.t132 323.425
R11967 gnd.n3570 gnd.n3544 289.615
R11968 gnd.n3538 gnd.n3512 289.615
R11969 gnd.n3506 gnd.n3480 289.615
R11970 gnd.n3475 gnd.n3449 289.615
R11971 gnd.n3443 gnd.n3417 289.615
R11972 gnd.n3411 gnd.n3385 289.615
R11973 gnd.n3379 gnd.n3353 289.615
R11974 gnd.n3348 gnd.n3322 289.615
R11975 gnd.n2796 gnd.t128 279.217
R11976 gnd.n2306 gnd.t34 279.217
R11977 gnd.n1185 gnd.t40 260.649
R11978 gnd.n4998 gnd.t79 260.649
R11979 gnd.n5848 gnd.n5847 256.663
R11980 gnd.n5848 gnd.n1144 256.663
R11981 gnd.n5848 gnd.n1145 256.663
R11982 gnd.n5848 gnd.n1146 256.663
R11983 gnd.n5848 gnd.n1147 256.663
R11984 gnd.n5848 gnd.n1148 256.663
R11985 gnd.n5848 gnd.n1149 256.663
R11986 gnd.n5848 gnd.n1150 256.663
R11987 gnd.n5848 gnd.n1151 256.663
R11988 gnd.n5848 gnd.n1152 256.663
R11989 gnd.n5848 gnd.n1153 256.663
R11990 gnd.n5848 gnd.n1154 256.663
R11991 gnd.n5848 gnd.n1155 256.663
R11992 gnd.n5848 gnd.n1156 256.663
R11993 gnd.n5848 gnd.n1157 256.663
R11994 gnd.n5848 gnd.n1158 256.663
R11995 gnd.n5851 gnd.n1141 256.663
R11996 gnd.n5849 gnd.n5848 256.663
R11997 gnd.n5848 gnd.n1159 256.663
R11998 gnd.n5848 gnd.n1160 256.663
R11999 gnd.n5848 gnd.n1161 256.663
R12000 gnd.n5848 gnd.n1162 256.663
R12001 gnd.n5848 gnd.n1163 256.663
R12002 gnd.n5848 gnd.n1164 256.663
R12003 gnd.n5848 gnd.n1165 256.663
R12004 gnd.n5848 gnd.n1166 256.663
R12005 gnd.n5848 gnd.n1167 256.663
R12006 gnd.n5848 gnd.n1168 256.663
R12007 gnd.n5848 gnd.n1169 256.663
R12008 gnd.n5848 gnd.n1170 256.663
R12009 gnd.n5848 gnd.n1171 256.663
R12010 gnd.n5848 gnd.n1172 256.663
R12011 gnd.n5848 gnd.n1173 256.663
R12012 gnd.n5848 gnd.n1174 256.663
R12013 gnd.n5147 gnd.n1752 256.663
R12014 gnd.n5147 gnd.n1753 256.663
R12015 gnd.n5147 gnd.n1754 256.663
R12016 gnd.n5147 gnd.n1755 256.663
R12017 gnd.n5147 gnd.n1756 256.663
R12018 gnd.n5147 gnd.n1757 256.663
R12019 gnd.n5147 gnd.n1758 256.663
R12020 gnd.n5147 gnd.n1759 256.663
R12021 gnd.n5147 gnd.n1760 256.663
R12022 gnd.n5147 gnd.n1761 256.663
R12023 gnd.n5147 gnd.n1762 256.663
R12024 gnd.n5147 gnd.n1763 256.663
R12025 gnd.n5147 gnd.n1764 256.663
R12026 gnd.n5147 gnd.n1765 256.663
R12027 gnd.n5147 gnd.n1766 256.663
R12028 gnd.n5147 gnd.n1767 256.663
R12029 gnd.n1768 gnd.n1455 256.663
R12030 gnd.n5147 gnd.n1750 256.663
R12031 gnd.n5147 gnd.n1749 256.663
R12032 gnd.n5147 gnd.n1748 256.663
R12033 gnd.n5147 gnd.n1747 256.663
R12034 gnd.n5147 gnd.n1746 256.663
R12035 gnd.n5147 gnd.n1745 256.663
R12036 gnd.n5147 gnd.n1744 256.663
R12037 gnd.n5147 gnd.n1743 256.663
R12038 gnd.n5147 gnd.n1742 256.663
R12039 gnd.n5147 gnd.n1741 256.663
R12040 gnd.n5147 gnd.n1740 256.663
R12041 gnd.n5147 gnd.n1739 256.663
R12042 gnd.n5147 gnd.n1738 256.663
R12043 gnd.n5147 gnd.n1737 256.663
R12044 gnd.n5147 gnd.n1736 256.663
R12045 gnd.n5147 gnd.n1735 256.663
R12046 gnd.n5147 gnd.n1734 256.663
R12047 gnd.n3729 gnd.n3703 242.672
R12048 gnd.n3731 gnd.n3703 242.672
R12049 gnd.n3739 gnd.n3703 242.672
R12050 gnd.n3741 gnd.n3703 242.672
R12051 gnd.n3749 gnd.n3703 242.672
R12052 gnd.n3751 gnd.n3703 242.672
R12053 gnd.n3759 gnd.n3703 242.672
R12054 gnd.n3761 gnd.n3703 242.672
R12055 gnd.n3769 gnd.n3703 242.672
R12056 gnd.n5903 gnd.n5902 242.672
R12057 gnd.n5902 gnd.n978 242.672
R12058 gnd.n5902 gnd.n976 242.672
R12059 gnd.n5902 gnd.n975 242.672
R12060 gnd.n5902 gnd.n973 242.672
R12061 gnd.n5902 gnd.n971 242.672
R12062 gnd.n5902 gnd.n970 242.672
R12063 gnd.n5902 gnd.n968 242.672
R12064 gnd.n5902 gnd.n966 242.672
R12065 gnd.n2850 gnd.n2849 242.672
R12066 gnd.n2850 gnd.n2760 242.672
R12067 gnd.n2850 gnd.n2761 242.672
R12068 gnd.n2850 gnd.n2762 242.672
R12069 gnd.n2850 gnd.n2763 242.672
R12070 gnd.n2850 gnd.n2764 242.672
R12071 gnd.n2850 gnd.n2765 242.672
R12072 gnd.n2850 gnd.n2766 242.672
R12073 gnd.n2850 gnd.n2767 242.672
R12074 gnd.n2850 gnd.n2768 242.672
R12075 gnd.n2850 gnd.n2769 242.672
R12076 gnd.n2850 gnd.n2770 242.672
R12077 gnd.n2851 gnd.n2850 242.672
R12078 gnd.n3702 gnd.n2255 242.672
R12079 gnd.n3702 gnd.n2254 242.672
R12080 gnd.n3702 gnd.n2253 242.672
R12081 gnd.n3702 gnd.n2252 242.672
R12082 gnd.n3702 gnd.n2251 242.672
R12083 gnd.n3702 gnd.n2250 242.672
R12084 gnd.n3702 gnd.n2249 242.672
R12085 gnd.n3702 gnd.n2248 242.672
R12086 gnd.n3702 gnd.n2247 242.672
R12087 gnd.n3702 gnd.n2246 242.672
R12088 gnd.n3702 gnd.n2245 242.672
R12089 gnd.n3702 gnd.n2244 242.672
R12090 gnd.n3702 gnd.n2243 242.672
R12091 gnd.n5586 gnd.n1410 242.672
R12092 gnd.n5586 gnd.n1412 242.672
R12093 gnd.n5586 gnd.n1413 242.672
R12094 gnd.n5586 gnd.n1415 242.672
R12095 gnd.n5586 gnd.n1417 242.672
R12096 gnd.n5586 gnd.n1418 242.672
R12097 gnd.n5586 gnd.n1420 242.672
R12098 gnd.n5586 gnd.n1422 242.672
R12099 gnd.n5587 gnd.n5586 242.672
R12100 gnd.n7187 gnd.n7186 242.672
R12101 gnd.n7186 gnd.n6973 242.672
R12102 gnd.n7186 gnd.n6922 242.672
R12103 gnd.n7186 gnd.n6921 242.672
R12104 gnd.n7186 gnd.n6920 242.672
R12105 gnd.n7186 gnd.n6919 242.672
R12106 gnd.n7186 gnd.n6918 242.672
R12107 gnd.n7186 gnd.n6917 242.672
R12108 gnd.n7186 gnd.n6916 242.672
R12109 gnd.n2934 gnd.n2933 242.672
R12110 gnd.n2933 gnd.n2672 242.672
R12111 gnd.n2933 gnd.n2673 242.672
R12112 gnd.n2933 gnd.n2674 242.672
R12113 gnd.n2933 gnd.n2675 242.672
R12114 gnd.n2933 gnd.n2676 242.672
R12115 gnd.n2933 gnd.n2677 242.672
R12116 gnd.n2933 gnd.n2678 242.672
R12117 gnd.n3702 gnd.n2256 242.672
R12118 gnd.n3702 gnd.n2257 242.672
R12119 gnd.n3702 gnd.n2258 242.672
R12120 gnd.n3702 gnd.n2259 242.672
R12121 gnd.n3702 gnd.n2260 242.672
R12122 gnd.n3702 gnd.n2261 242.672
R12123 gnd.n3702 gnd.n2262 242.672
R12124 gnd.n3702 gnd.n2263 242.672
R12125 gnd.n3989 gnd.n3703 242.672
R12126 gnd.n3784 gnd.n3703 242.672
R12127 gnd.n3982 gnd.n3703 242.672
R12128 gnd.n3976 gnd.n3703 242.672
R12129 gnd.n3974 gnd.n3703 242.672
R12130 gnd.n3968 gnd.n3703 242.672
R12131 gnd.n3966 gnd.n3703 242.672
R12132 gnd.n3960 gnd.n3703 242.672
R12133 gnd.n3958 gnd.n3703 242.672
R12134 gnd.n3952 gnd.n3703 242.672
R12135 gnd.n3950 gnd.n3703 242.672
R12136 gnd.n3944 gnd.n3703 242.672
R12137 gnd.n3942 gnd.n3703 242.672
R12138 gnd.n3936 gnd.n3703 242.672
R12139 gnd.n3934 gnd.n3703 242.672
R12140 gnd.n3928 gnd.n3703 242.672
R12141 gnd.n3926 gnd.n3703 242.672
R12142 gnd.n3920 gnd.n3703 242.672
R12143 gnd.n3918 gnd.n3703 242.672
R12144 gnd.n3912 gnd.n3703 242.672
R12145 gnd.n3910 gnd.n3703 242.672
R12146 gnd.n3904 gnd.n3703 242.672
R12147 gnd.n3902 gnd.n3703 242.672
R12148 gnd.n3896 gnd.n3703 242.672
R12149 gnd.n3894 gnd.n3703 242.672
R12150 gnd.n3888 gnd.n3703 242.672
R12151 gnd.n3886 gnd.n3703 242.672
R12152 gnd.n3880 gnd.n3703 242.672
R12153 gnd.n3878 gnd.n3703 242.672
R12154 gnd.n5902 gnd.n980 242.672
R12155 gnd.n5902 gnd.n981 242.672
R12156 gnd.n5902 gnd.n982 242.672
R12157 gnd.n5902 gnd.n983 242.672
R12158 gnd.n5902 gnd.n984 242.672
R12159 gnd.n5902 gnd.n985 242.672
R12160 gnd.n5902 gnd.n986 242.672
R12161 gnd.n5902 gnd.n987 242.672
R12162 gnd.n5902 gnd.n988 242.672
R12163 gnd.n5902 gnd.n989 242.672
R12164 gnd.n5902 gnd.n990 242.672
R12165 gnd.n5902 gnd.n991 242.672
R12166 gnd.n5902 gnd.n992 242.672
R12167 gnd.n5902 gnd.n993 242.672
R12168 gnd.n5902 gnd.n994 242.672
R12169 gnd.n5902 gnd.n995 242.672
R12170 gnd.n5852 gnd.n1041 242.672
R12171 gnd.n5902 gnd.n996 242.672
R12172 gnd.n5902 gnd.n997 242.672
R12173 gnd.n5902 gnd.n998 242.672
R12174 gnd.n5902 gnd.n999 242.672
R12175 gnd.n5902 gnd.n1000 242.672
R12176 gnd.n5902 gnd.n1001 242.672
R12177 gnd.n5902 gnd.n1002 242.672
R12178 gnd.n5902 gnd.n1003 242.672
R12179 gnd.n5902 gnd.n1004 242.672
R12180 gnd.n5902 gnd.n1005 242.672
R12181 gnd.n5902 gnd.n1006 242.672
R12182 gnd.n5902 gnd.n1007 242.672
R12183 gnd.n5902 gnd.n5901 242.672
R12184 gnd.n5586 gnd.n5585 242.672
R12185 gnd.n5586 gnd.n1382 242.672
R12186 gnd.n5586 gnd.n1383 242.672
R12187 gnd.n5586 gnd.n1384 242.672
R12188 gnd.n5586 gnd.n1385 242.672
R12189 gnd.n5586 gnd.n1386 242.672
R12190 gnd.n5586 gnd.n1387 242.672
R12191 gnd.n5586 gnd.n1388 242.672
R12192 gnd.n5586 gnd.n1389 242.672
R12193 gnd.n5586 gnd.n1390 242.672
R12194 gnd.n5586 gnd.n1391 242.672
R12195 gnd.n5586 gnd.n1392 242.672
R12196 gnd.n5586 gnd.n1393 242.672
R12197 gnd.n5533 gnd.n1456 242.672
R12198 gnd.n5586 gnd.n1394 242.672
R12199 gnd.n5586 gnd.n1395 242.672
R12200 gnd.n5586 gnd.n1396 242.672
R12201 gnd.n5586 gnd.n1397 242.672
R12202 gnd.n5586 gnd.n1398 242.672
R12203 gnd.n5586 gnd.n1399 242.672
R12204 gnd.n5586 gnd.n1400 242.672
R12205 gnd.n5586 gnd.n1401 242.672
R12206 gnd.n5586 gnd.n1402 242.672
R12207 gnd.n5586 gnd.n1403 242.672
R12208 gnd.n5586 gnd.n1404 242.672
R12209 gnd.n5586 gnd.n1405 242.672
R12210 gnd.n5586 gnd.n1406 242.672
R12211 gnd.n5586 gnd.n1407 242.672
R12212 gnd.n5586 gnd.n1408 242.672
R12213 gnd.n5586 gnd.n1409 242.672
R12214 gnd.n7186 gnd.n6974 242.672
R12215 gnd.n7186 gnd.n6975 242.672
R12216 gnd.n7186 gnd.n6976 242.672
R12217 gnd.n7186 gnd.n6977 242.672
R12218 gnd.n7186 gnd.n6978 242.672
R12219 gnd.n7186 gnd.n6979 242.672
R12220 gnd.n7186 gnd.n6980 242.672
R12221 gnd.n7186 gnd.n6981 242.672
R12222 gnd.n7186 gnd.n6982 242.672
R12223 gnd.n7186 gnd.n6983 242.672
R12224 gnd.n7186 gnd.n6984 242.672
R12225 gnd.n7186 gnd.n6985 242.672
R12226 gnd.n7186 gnd.n6986 242.672
R12227 gnd.n7186 gnd.n6987 242.672
R12228 gnd.n7186 gnd.n6988 242.672
R12229 gnd.n7186 gnd.n6989 242.672
R12230 gnd.n7186 gnd.n6990 242.672
R12231 gnd.n7186 gnd.n6991 242.672
R12232 gnd.n7186 gnd.n6992 242.672
R12233 gnd.n7186 gnd.n6993 242.672
R12234 gnd.n7186 gnd.n6994 242.672
R12235 gnd.n7186 gnd.n6995 242.672
R12236 gnd.n7186 gnd.n6996 242.672
R12237 gnd.n7186 gnd.n6997 242.672
R12238 gnd.n7186 gnd.n6998 242.672
R12239 gnd.n7186 gnd.n6999 242.672
R12240 gnd.n7186 gnd.n7000 242.672
R12241 gnd.n7186 gnd.n7001 242.672
R12242 gnd.n7186 gnd.n7185 242.672
R12243 gnd.n5967 gnd.n5966 242.672
R12244 gnd.n5967 gnd.n877 242.672
R12245 gnd.n5967 gnd.n878 242.672
R12246 gnd.n5967 gnd.n879 242.672
R12247 gnd.n5967 gnd.n880 242.672
R12248 gnd.n5967 gnd.n881 242.672
R12249 gnd.n5967 gnd.n882 242.672
R12250 gnd.n5967 gnd.n883 242.672
R12251 gnd.n5967 gnd.n884 242.672
R12252 gnd.n5967 gnd.n885 242.672
R12253 gnd.n5967 gnd.n886 242.672
R12254 gnd.n5967 gnd.n887 242.672
R12255 gnd.n5967 gnd.n889 242.672
R12256 gnd.n5968 gnd.n5967 242.672
R12257 gnd.n5259 gnd.n1662 242.672
R12258 gnd.n5259 gnd.n1660 242.672
R12259 gnd.n5259 gnd.n1659 242.672
R12260 gnd.n5259 gnd.n1657 242.672
R12261 gnd.n5259 gnd.n1655 242.672
R12262 gnd.n5259 gnd.n1654 242.672
R12263 gnd.n5259 gnd.n1652 242.672
R12264 gnd.n5259 gnd.n1650 242.672
R12265 gnd.n5259 gnd.n1649 242.672
R12266 gnd.n5259 gnd.n1647 242.672
R12267 gnd.n5259 gnd.n1646 242.672
R12268 gnd.n5259 gnd.n1644 242.672
R12269 gnd.n5260 gnd.n5259 242.672
R12270 gnd.n5259 gnd.n1665 242.672
R12271 gnd.n7002 gnd.n166 240.244
R12272 gnd.n7184 gnd.n7003 240.244
R12273 gnd.n7180 gnd.n7179 240.244
R12274 gnd.n7176 gnd.n7175 240.244
R12275 gnd.n7172 gnd.n7171 240.244
R12276 gnd.n7168 gnd.n7167 240.244
R12277 gnd.n7164 gnd.n7163 240.244
R12278 gnd.n7160 gnd.n7159 240.244
R12279 gnd.n7156 gnd.n7155 240.244
R12280 gnd.n7149 gnd.n7148 240.244
R12281 gnd.n7145 gnd.n7144 240.244
R12282 gnd.n7141 gnd.n7140 240.244
R12283 gnd.n7137 gnd.n7136 240.244
R12284 gnd.n7133 gnd.n7132 240.244
R12285 gnd.n7129 gnd.n7128 240.244
R12286 gnd.n7125 gnd.n7124 240.244
R12287 gnd.n7121 gnd.n7120 240.244
R12288 gnd.n7117 gnd.n7116 240.244
R12289 gnd.n7113 gnd.n7112 240.244
R12290 gnd.n7106 gnd.n7105 240.244
R12291 gnd.n7103 gnd.n7102 240.244
R12292 gnd.n7099 gnd.n7098 240.244
R12293 gnd.n7095 gnd.n7094 240.244
R12294 gnd.n7091 gnd.n7090 240.244
R12295 gnd.n7087 gnd.n7086 240.244
R12296 gnd.n7083 gnd.n7082 240.244
R12297 gnd.n7079 gnd.n7078 240.244
R12298 gnd.n7075 gnd.n7074 240.244
R12299 gnd.n7071 gnd.n7070 240.244
R12300 gnd.n5466 gnd.n1489 240.244
R12301 gnd.n5458 gnd.n1489 240.244
R12302 gnd.n5458 gnd.n1500 240.244
R12303 gnd.n1516 gnd.n1500 240.244
R12304 gnd.n5276 gnd.n1516 240.244
R12305 gnd.n5276 gnd.n1529 240.244
R12306 gnd.n5282 gnd.n1529 240.244
R12307 gnd.n5282 gnd.n1539 240.244
R12308 gnd.n5289 gnd.n1539 240.244
R12309 gnd.n5289 gnd.n1549 240.244
R12310 gnd.n1622 gnd.n1549 240.244
R12311 gnd.n1622 gnd.n1559 240.244
R12312 gnd.n5359 gnd.n1559 240.244
R12313 gnd.n5359 gnd.n1569 240.244
R12314 gnd.n5364 gnd.n1569 240.244
R12315 gnd.n5364 gnd.n1576 240.244
R12316 gnd.n5378 gnd.n1576 240.244
R12317 gnd.n5378 gnd.n1586 240.244
R12318 gnd.n1592 gnd.n1586 240.244
R12319 gnd.n5387 gnd.n1592 240.244
R12320 gnd.n5388 gnd.n5387 240.244
R12321 gnd.n5388 gnd.n1604 240.244
R12322 gnd.n1604 gnd.n74 240.244
R12323 gnd.n177 gnd.n74 240.244
R12324 gnd.n6890 gnd.n177 240.244
R12325 gnd.n6890 gnd.n91 240.244
R12326 gnd.n7217 gnd.n91 240.244
R12327 gnd.n7217 gnd.n102 240.244
R12328 gnd.n7221 gnd.n102 240.244
R12329 gnd.n7221 gnd.n112 240.244
R12330 gnd.n7224 gnd.n112 240.244
R12331 gnd.n7224 gnd.n121 240.244
R12332 gnd.n7228 gnd.n121 240.244
R12333 gnd.n7228 gnd.n131 240.244
R12334 gnd.n7231 gnd.n131 240.244
R12335 gnd.n7231 gnd.n140 240.244
R12336 gnd.n7235 gnd.n140 240.244
R12337 gnd.n7235 gnd.n150 240.244
R12338 gnd.n7238 gnd.n150 240.244
R12339 gnd.n7238 gnd.n159 240.244
R12340 gnd.n7241 gnd.n159 240.244
R12341 gnd.n7241 gnd.n168 240.244
R12342 gnd.n1425 gnd.n1424 240.244
R12343 gnd.n5579 gnd.n1424 240.244
R12344 gnd.n5577 gnd.n5576 240.244
R12345 gnd.n5573 gnd.n5572 240.244
R12346 gnd.n5569 gnd.n5568 240.244
R12347 gnd.n5565 gnd.n5564 240.244
R12348 gnd.n5561 gnd.n5560 240.244
R12349 gnd.n5557 gnd.n5556 240.244
R12350 gnd.n5553 gnd.n5552 240.244
R12351 gnd.n5548 gnd.n5547 240.244
R12352 gnd.n5544 gnd.n5543 240.244
R12353 gnd.n5540 gnd.n5539 240.244
R12354 gnd.n5536 gnd.n5535 240.244
R12355 gnd.n5531 gnd.n5530 240.244
R12356 gnd.n5527 gnd.n5526 240.244
R12357 gnd.n5523 gnd.n5522 240.244
R12358 gnd.n5519 gnd.n5518 240.244
R12359 gnd.n5515 gnd.n5514 240.244
R12360 gnd.n5511 gnd.n5510 240.244
R12361 gnd.n5507 gnd.n5506 240.244
R12362 gnd.n5503 gnd.n5502 240.244
R12363 gnd.n5499 gnd.n5498 240.244
R12364 gnd.n5495 gnd.n5494 240.244
R12365 gnd.n5491 gnd.n5490 240.244
R12366 gnd.n5487 gnd.n5486 240.244
R12367 gnd.n5483 gnd.n5482 240.244
R12368 gnd.n5479 gnd.n5478 240.244
R12369 gnd.n5475 gnd.n5474 240.244
R12370 gnd.n1504 gnd.n1426 240.244
R12371 gnd.n5456 gnd.n1504 240.244
R12372 gnd.n5456 gnd.n1505 240.244
R12373 gnd.n5452 gnd.n1505 240.244
R12374 gnd.n5452 gnd.n1514 240.244
R12375 gnd.n5444 gnd.n1514 240.244
R12376 gnd.n5444 gnd.n1531 240.244
R12377 gnd.n5440 gnd.n1531 240.244
R12378 gnd.n5440 gnd.n1537 240.244
R12379 gnd.n5432 gnd.n1537 240.244
R12380 gnd.n5432 gnd.n1552 240.244
R12381 gnd.n5428 gnd.n1552 240.244
R12382 gnd.n5428 gnd.n1558 240.244
R12383 gnd.n5420 gnd.n1558 240.244
R12384 gnd.n5420 gnd.n1571 240.244
R12385 gnd.n5416 gnd.n1571 240.244
R12386 gnd.n5416 gnd.n1574 240.244
R12387 gnd.n5408 gnd.n1574 240.244
R12388 gnd.n5408 gnd.n5405 240.244
R12389 gnd.n5405 gnd.n1589 240.244
R12390 gnd.n1602 gnd.n1589 240.244
R12391 gnd.n1602 gnd.n77 240.244
R12392 gnd.n7302 gnd.n77 240.244
R12393 gnd.n7302 gnd.n78 240.244
R12394 gnd.n88 gnd.n78 240.244
R12395 gnd.n7296 gnd.n88 240.244
R12396 gnd.n7296 gnd.n89 240.244
R12397 gnd.n7288 gnd.n89 240.244
R12398 gnd.n7288 gnd.n105 240.244
R12399 gnd.n7284 gnd.n105 240.244
R12400 gnd.n7284 gnd.n110 240.244
R12401 gnd.n7276 gnd.n110 240.244
R12402 gnd.n7276 gnd.n123 240.244
R12403 gnd.n7272 gnd.n123 240.244
R12404 gnd.n7272 gnd.n129 240.244
R12405 gnd.n7264 gnd.n129 240.244
R12406 gnd.n7264 gnd.n143 240.244
R12407 gnd.n7260 gnd.n143 240.244
R12408 gnd.n7260 gnd.n149 240.244
R12409 gnd.n7252 gnd.n149 240.244
R12410 gnd.n7252 gnd.n161 240.244
R12411 gnd.n7248 gnd.n161 240.244
R12412 gnd.n1008 gnd.n858 240.244
R12413 gnd.n5900 gnd.n1009 240.244
R12414 gnd.n5896 gnd.n5895 240.244
R12415 gnd.n5892 gnd.n5891 240.244
R12416 gnd.n5888 gnd.n5887 240.244
R12417 gnd.n5884 gnd.n5883 240.244
R12418 gnd.n5880 gnd.n5879 240.244
R12419 gnd.n5876 gnd.n5875 240.244
R12420 gnd.n5872 gnd.n5871 240.244
R12421 gnd.n5867 gnd.n5866 240.244
R12422 gnd.n5863 gnd.n5862 240.244
R12423 gnd.n5859 gnd.n5858 240.244
R12424 gnd.n5855 gnd.n5854 240.244
R12425 gnd.n1134 gnd.n1133 240.244
R12426 gnd.n1131 gnd.n1130 240.244
R12427 gnd.n1127 gnd.n1126 240.244
R12428 gnd.n1123 gnd.n1122 240.244
R12429 gnd.n1119 gnd.n1118 240.244
R12430 gnd.n1112 gnd.n1111 240.244
R12431 gnd.n1109 gnd.n1108 240.244
R12432 gnd.n1105 gnd.n1104 240.244
R12433 gnd.n1101 gnd.n1100 240.244
R12434 gnd.n1097 gnd.n1096 240.244
R12435 gnd.n1093 gnd.n1092 240.244
R12436 gnd.n1089 gnd.n1088 240.244
R12437 gnd.n1085 gnd.n1084 240.244
R12438 gnd.n1081 gnd.n1080 240.244
R12439 gnd.n1077 gnd.n1076 240.244
R12440 gnd.n3704 gnd.n2238 240.244
R12441 gnd.n2238 gnd.n2230 240.244
R12442 gnd.n4004 gnd.n2230 240.244
R12443 gnd.n4004 gnd.n2222 240.244
R12444 gnd.n2222 gnd.n2214 240.244
R12445 gnd.n4036 gnd.n2214 240.244
R12446 gnd.n4036 gnd.n2205 240.244
R12447 gnd.n4039 gnd.n2205 240.244
R12448 gnd.n4039 gnd.n2197 240.244
R12449 gnd.n2197 gnd.n2189 240.244
R12450 gnd.n4073 gnd.n2189 240.244
R12451 gnd.n4073 gnd.n2178 240.244
R12452 gnd.n4076 gnd.n2178 240.244
R12453 gnd.n4076 gnd.n2171 240.244
R12454 gnd.n4079 gnd.n2171 240.244
R12455 gnd.n4079 gnd.n734 240.244
R12456 gnd.n4109 gnd.n734 240.244
R12457 gnd.n4109 gnd.n745 240.244
R12458 gnd.n4113 gnd.n745 240.244
R12459 gnd.n4113 gnd.n756 240.244
R12460 gnd.n4135 gnd.n756 240.244
R12461 gnd.n4135 gnd.n764 240.244
R12462 gnd.n2155 gnd.n764 240.244
R12463 gnd.n2155 gnd.n773 240.244
R12464 gnd.n4144 gnd.n773 240.244
R12465 gnd.n4144 gnd.n781 240.244
R12466 gnd.n2148 gnd.n781 240.244
R12467 gnd.n2148 gnd.n790 240.244
R12468 gnd.n4180 gnd.n790 240.244
R12469 gnd.n4180 gnd.n801 240.244
R12470 gnd.n2133 gnd.n801 240.244
R12471 gnd.n2133 gnd.n810 240.244
R12472 gnd.n4187 gnd.n810 240.244
R12473 gnd.n4187 gnd.n821 240.244
R12474 gnd.n4192 gnd.n821 240.244
R12475 gnd.n4192 gnd.n830 240.244
R12476 gnd.n4197 gnd.n830 240.244
R12477 gnd.n4197 gnd.n841 240.244
R12478 gnd.n4201 gnd.n841 240.244
R12479 gnd.n4201 gnd.n851 240.244
R12480 gnd.n5979 gnd.n851 240.244
R12481 gnd.n5979 gnd.n860 240.244
R12482 gnd.n3990 gnd.n3988 240.244
R12483 gnd.n3988 gnd.n3987 240.244
R12484 gnd.n3984 gnd.n3983 240.244
R12485 gnd.n3981 gnd.n3789 240.244
R12486 gnd.n3977 gnd.n3975 240.244
R12487 gnd.n3973 gnd.n3795 240.244
R12488 gnd.n3969 gnd.n3967 240.244
R12489 gnd.n3965 gnd.n3801 240.244
R12490 gnd.n3961 gnd.n3959 240.244
R12491 gnd.n3957 gnd.n3807 240.244
R12492 gnd.n3953 gnd.n3951 240.244
R12493 gnd.n3949 gnd.n3816 240.244
R12494 gnd.n3945 gnd.n3943 240.244
R12495 gnd.n3941 gnd.n3822 240.244
R12496 gnd.n3937 gnd.n3935 240.244
R12497 gnd.n3933 gnd.n3828 240.244
R12498 gnd.n3929 gnd.n3927 240.244
R12499 gnd.n3925 gnd.n3834 240.244
R12500 gnd.n3921 gnd.n3919 240.244
R12501 gnd.n3917 gnd.n3842 240.244
R12502 gnd.n3913 gnd.n3911 240.244
R12503 gnd.n3909 gnd.n3848 240.244
R12504 gnd.n3905 gnd.n3903 240.244
R12505 gnd.n3901 gnd.n3854 240.244
R12506 gnd.n3897 gnd.n3895 240.244
R12507 gnd.n3893 gnd.n3860 240.244
R12508 gnd.n3889 gnd.n3887 240.244
R12509 gnd.n3885 gnd.n3866 240.244
R12510 gnd.n3881 gnd.n3879 240.244
R12511 gnd.n3996 gnd.n2229 240.244
R12512 gnd.n4016 gnd.n2229 240.244
R12513 gnd.n4016 gnd.n2224 240.244
R12514 gnd.n4024 gnd.n2224 240.244
R12515 gnd.n4024 gnd.n2225 240.244
R12516 gnd.n2225 gnd.n2204 240.244
R12517 gnd.n4051 gnd.n2204 240.244
R12518 gnd.n4051 gnd.n2199 240.244
R12519 gnd.n4059 gnd.n2199 240.244
R12520 gnd.n4059 gnd.n2200 240.244
R12521 gnd.n2200 gnd.n2177 240.244
R12522 gnd.n4091 gnd.n2177 240.244
R12523 gnd.n4091 gnd.n2173 240.244
R12524 gnd.n4098 gnd.n2173 240.244
R12525 gnd.n4098 gnd.n738 240.244
R12526 gnd.n6065 gnd.n738 240.244
R12527 gnd.n6065 gnd.n739 240.244
R12528 gnd.n6060 gnd.n739 240.244
R12529 gnd.n6060 gnd.n743 240.244
R12530 gnd.n6052 gnd.n743 240.244
R12531 gnd.n6052 gnd.n759 240.244
R12532 gnd.n6047 gnd.n759 240.244
R12533 gnd.n6047 gnd.n762 240.244
R12534 gnd.n6039 gnd.n762 240.244
R12535 gnd.n6039 gnd.n776 240.244
R12536 gnd.n6034 gnd.n776 240.244
R12537 gnd.n6034 gnd.n779 240.244
R12538 gnd.n6026 gnd.n779 240.244
R12539 gnd.n6026 gnd.n793 240.244
R12540 gnd.n6022 gnd.n793 240.244
R12541 gnd.n6022 gnd.n799 240.244
R12542 gnd.n6014 gnd.n799 240.244
R12543 gnd.n6014 gnd.n813 240.244
R12544 gnd.n6010 gnd.n813 240.244
R12545 gnd.n6010 gnd.n819 240.244
R12546 gnd.n6002 gnd.n819 240.244
R12547 gnd.n6002 gnd.n833 240.244
R12548 gnd.n5998 gnd.n833 240.244
R12549 gnd.n5998 gnd.n839 240.244
R12550 gnd.n5990 gnd.n839 240.244
R12551 gnd.n5990 gnd.n853 240.244
R12552 gnd.n5986 gnd.n853 240.244
R12553 gnd.n3701 gnd.n2265 240.244
R12554 gnd.n3694 gnd.n3693 240.244
R12555 gnd.n3691 gnd.n3690 240.244
R12556 gnd.n3687 gnd.n3686 240.244
R12557 gnd.n3683 gnd.n3682 240.244
R12558 gnd.n3679 gnd.n3678 240.244
R12559 gnd.n3675 gnd.n3674 240.244
R12560 gnd.n3671 gnd.n3670 240.244
R12561 gnd.n2945 gnd.n2657 240.244
R12562 gnd.n2955 gnd.n2657 240.244
R12563 gnd.n2955 gnd.n2648 240.244
R12564 gnd.n2648 gnd.n2637 240.244
R12565 gnd.n2976 gnd.n2637 240.244
R12566 gnd.n2976 gnd.n2631 240.244
R12567 gnd.n2986 gnd.n2631 240.244
R12568 gnd.n2986 gnd.n2620 240.244
R12569 gnd.n2620 gnd.n2612 240.244
R12570 gnd.n3004 gnd.n2612 240.244
R12571 gnd.n3005 gnd.n3004 240.244
R12572 gnd.n3005 gnd.n2597 240.244
R12573 gnd.n3007 gnd.n2597 240.244
R12574 gnd.n3007 gnd.n2583 240.244
R12575 gnd.n3049 gnd.n2583 240.244
R12576 gnd.n3050 gnd.n3049 240.244
R12577 gnd.n3053 gnd.n3050 240.244
R12578 gnd.n3053 gnd.n2538 240.244
R12579 gnd.n2578 gnd.n2538 240.244
R12580 gnd.n2578 gnd.n2548 240.244
R12581 gnd.n3063 gnd.n2548 240.244
R12582 gnd.n3063 gnd.n2569 240.244
R12583 gnd.n3073 gnd.n2569 240.244
R12584 gnd.n3073 gnd.n2467 240.244
R12585 gnd.n3118 gnd.n2467 240.244
R12586 gnd.n3118 gnd.n2453 240.244
R12587 gnd.n3140 gnd.n2453 240.244
R12588 gnd.n3141 gnd.n3140 240.244
R12589 gnd.n3141 gnd.n2440 240.244
R12590 gnd.n2440 gnd.n2429 240.244
R12591 gnd.n3172 gnd.n2429 240.244
R12592 gnd.n3173 gnd.n3172 240.244
R12593 gnd.n3174 gnd.n3173 240.244
R12594 gnd.n3174 gnd.n2414 240.244
R12595 gnd.n2414 gnd.n2413 240.244
R12596 gnd.n2413 gnd.n2398 240.244
R12597 gnd.n3225 gnd.n2398 240.244
R12598 gnd.n3226 gnd.n3225 240.244
R12599 gnd.n3226 gnd.n2385 240.244
R12600 gnd.n2385 gnd.n2374 240.244
R12601 gnd.n3257 gnd.n2374 240.244
R12602 gnd.n3258 gnd.n3257 240.244
R12603 gnd.n3259 gnd.n3258 240.244
R12604 gnd.n3259 gnd.n2358 240.244
R12605 gnd.n2358 gnd.n2357 240.244
R12606 gnd.n2357 gnd.n2344 240.244
R12607 gnd.n3314 gnd.n2344 240.244
R12608 gnd.n3315 gnd.n3314 240.244
R12609 gnd.n3315 gnd.n2331 240.244
R12610 gnd.n2331 gnd.n2321 240.244
R12611 gnd.n3602 gnd.n2321 240.244
R12612 gnd.n3605 gnd.n3602 240.244
R12613 gnd.n3605 gnd.n3604 240.244
R12614 gnd.n2935 gnd.n2670 240.244
R12615 gnd.n2691 gnd.n2670 240.244
R12616 gnd.n2694 gnd.n2693 240.244
R12617 gnd.n2701 gnd.n2700 240.244
R12618 gnd.n2704 gnd.n2703 240.244
R12619 gnd.n2711 gnd.n2710 240.244
R12620 gnd.n2714 gnd.n2713 240.244
R12621 gnd.n2721 gnd.n2720 240.244
R12622 gnd.n2943 gnd.n2667 240.244
R12623 gnd.n2667 gnd.n2646 240.244
R12624 gnd.n2966 gnd.n2646 240.244
R12625 gnd.n2966 gnd.n2640 240.244
R12626 gnd.n2974 gnd.n2640 240.244
R12627 gnd.n2974 gnd.n2642 240.244
R12628 gnd.n2642 gnd.n2618 240.244
R12629 gnd.n2996 gnd.n2618 240.244
R12630 gnd.n2996 gnd.n2614 240.244
R12631 gnd.n3002 gnd.n2614 240.244
R12632 gnd.n3002 gnd.n2596 240.244
R12633 gnd.n3027 gnd.n2596 240.244
R12634 gnd.n3027 gnd.n2591 240.244
R12635 gnd.n3039 gnd.n2591 240.244
R12636 gnd.n3039 gnd.n2592 240.244
R12637 gnd.n3035 gnd.n2592 240.244
R12638 gnd.n3035 gnd.n2540 240.244
R12639 gnd.n3087 gnd.n2540 240.244
R12640 gnd.n3087 gnd.n2541 240.244
R12641 gnd.n3083 gnd.n2541 240.244
R12642 gnd.n3083 gnd.n2547 240.244
R12643 gnd.n2567 gnd.n2547 240.244
R12644 gnd.n2567 gnd.n2465 240.244
R12645 gnd.n3122 gnd.n2465 240.244
R12646 gnd.n3122 gnd.n2460 240.244
R12647 gnd.n3130 gnd.n2460 240.244
R12648 gnd.n3130 gnd.n2461 240.244
R12649 gnd.n2461 gnd.n2438 240.244
R12650 gnd.n3162 gnd.n2438 240.244
R12651 gnd.n3162 gnd.n2433 240.244
R12652 gnd.n3170 gnd.n2433 240.244
R12653 gnd.n3170 gnd.n2434 240.244
R12654 gnd.n2434 gnd.n2411 240.244
R12655 gnd.n3207 gnd.n2411 240.244
R12656 gnd.n3207 gnd.n2406 240.244
R12657 gnd.n3215 gnd.n2406 240.244
R12658 gnd.n3215 gnd.n2407 240.244
R12659 gnd.n2407 gnd.n2383 240.244
R12660 gnd.n3247 gnd.n2383 240.244
R12661 gnd.n3247 gnd.n2378 240.244
R12662 gnd.n3255 gnd.n2378 240.244
R12663 gnd.n3255 gnd.n2379 240.244
R12664 gnd.n2379 gnd.n2356 240.244
R12665 gnd.n3296 gnd.n2356 240.244
R12666 gnd.n3296 gnd.n2351 240.244
R12667 gnd.n3304 gnd.n2351 240.244
R12668 gnd.n3304 gnd.n2352 240.244
R12669 gnd.n2352 gnd.n2329 240.244
R12670 gnd.n3590 gnd.n2329 240.244
R12671 gnd.n3590 gnd.n2324 240.244
R12672 gnd.n3600 gnd.n2324 240.244
R12673 gnd.n3600 gnd.n2325 240.244
R12674 gnd.n2325 gnd.n2264 240.244
R12675 gnd.n6934 gnd.n171 240.244
R12676 gnd.n6937 gnd.n6936 240.244
R12677 gnd.n6944 gnd.n6943 240.244
R12678 gnd.n6947 gnd.n6946 240.244
R12679 gnd.n6954 gnd.n6953 240.244
R12680 gnd.n6957 gnd.n6956 240.244
R12681 gnd.n6964 gnd.n6963 240.244
R12682 gnd.n6966 gnd.n6923 240.244
R12683 gnd.n6972 gnd.n6915 240.244
R12684 gnd.n5306 gnd.n1492 240.244
R12685 gnd.n5306 gnd.n1501 240.244
R12686 gnd.n5269 gnd.n1501 240.244
R12687 gnd.n5269 gnd.n1517 240.244
R12688 gnd.n5270 gnd.n1517 240.244
R12689 gnd.n5270 gnd.n1530 240.244
R12690 gnd.n5273 gnd.n1530 240.244
R12691 gnd.n5273 gnd.n1540 240.244
R12692 gnd.n5291 gnd.n1540 240.244
R12693 gnd.n5291 gnd.n1550 240.244
R12694 gnd.n5351 gnd.n1550 240.244
R12695 gnd.n5351 gnd.n1560 240.244
R12696 gnd.n5357 gnd.n1560 240.244
R12697 gnd.n5357 gnd.n1570 240.244
R12698 gnd.n5366 gnd.n1570 240.244
R12699 gnd.n5366 gnd.n1577 240.244
R12700 gnd.n5376 gnd.n1577 240.244
R12701 gnd.n5376 gnd.n1587 240.244
R12702 gnd.n1593 gnd.n1587 240.244
R12703 gnd.n1610 gnd.n1593 240.244
R12704 gnd.n1610 gnd.n1609 240.244
R12705 gnd.n1609 gnd.n70 240.244
R12706 gnd.n7304 gnd.n70 240.244
R12707 gnd.n7304 gnd.n72 240.244
R12708 gnd.n6892 gnd.n72 240.244
R12709 gnd.n6892 gnd.n92 240.244
R12710 gnd.n7215 gnd.n92 240.244
R12711 gnd.n7215 gnd.n103 240.244
R12712 gnd.n7211 gnd.n103 240.244
R12713 gnd.n7211 gnd.n113 240.244
R12714 gnd.n7208 gnd.n113 240.244
R12715 gnd.n7208 gnd.n122 240.244
R12716 gnd.n7205 gnd.n122 240.244
R12717 gnd.n7205 gnd.n132 240.244
R12718 gnd.n7202 gnd.n132 240.244
R12719 gnd.n7202 gnd.n141 240.244
R12720 gnd.n7199 gnd.n141 240.244
R12721 gnd.n7199 gnd.n151 240.244
R12722 gnd.n7196 gnd.n151 240.244
R12723 gnd.n7196 gnd.n160 240.244
R12724 gnd.n7193 gnd.n160 240.244
R12725 gnd.n7193 gnd.n169 240.244
R12726 gnd.n1336 gnd.n1335 240.244
R12727 gnd.n1411 gnd.n1343 240.244
R12728 gnd.n1414 gnd.n1344 240.244
R12729 gnd.n1352 gnd.n1351 240.244
R12730 gnd.n1416 gnd.n1359 240.244
R12731 gnd.n1419 gnd.n1360 240.244
R12732 gnd.n1368 gnd.n1367 240.244
R12733 gnd.n1421 gnd.n1377 240.244
R12734 gnd.n5588 gnd.n1380 240.244
R12735 gnd.n5464 gnd.n1495 240.244
R12736 gnd.n1503 gnd.n1495 240.244
R12737 gnd.n1519 gnd.n1503 240.244
R12738 gnd.n5450 gnd.n1519 240.244
R12739 gnd.n5450 gnd.n1520 240.244
R12740 gnd.n5446 gnd.n1520 240.244
R12741 gnd.n5446 gnd.n1527 240.244
R12742 gnd.n5438 gnd.n1527 240.244
R12743 gnd.n5438 gnd.n1542 240.244
R12744 gnd.n5434 gnd.n1542 240.244
R12745 gnd.n5434 gnd.n1547 240.244
R12746 gnd.n5426 gnd.n1547 240.244
R12747 gnd.n5426 gnd.n1562 240.244
R12748 gnd.n5422 gnd.n1562 240.244
R12749 gnd.n5422 gnd.n1567 240.244
R12750 gnd.n5414 gnd.n1567 240.244
R12751 gnd.n5414 gnd.n1579 240.244
R12752 gnd.n5410 gnd.n1579 240.244
R12753 gnd.n5410 gnd.n1584 240.244
R12754 gnd.n5385 gnd.n1584 240.244
R12755 gnd.n5385 gnd.n1605 240.244
R12756 gnd.n5394 gnd.n1605 240.244
R12757 gnd.n5394 gnd.n76 240.244
R12758 gnd.n6885 gnd.n76 240.244
R12759 gnd.n6885 gnd.n94 240.244
R12760 gnd.n7294 gnd.n94 240.244
R12761 gnd.n7294 gnd.n95 240.244
R12762 gnd.n7290 gnd.n95 240.244
R12763 gnd.n7290 gnd.n101 240.244
R12764 gnd.n7282 gnd.n101 240.244
R12765 gnd.n7282 gnd.n114 240.244
R12766 gnd.n7278 gnd.n114 240.244
R12767 gnd.n7278 gnd.n119 240.244
R12768 gnd.n7270 gnd.n119 240.244
R12769 gnd.n7270 gnd.n134 240.244
R12770 gnd.n7266 gnd.n134 240.244
R12771 gnd.n7266 gnd.n139 240.244
R12772 gnd.n7258 gnd.n139 240.244
R12773 gnd.n7258 gnd.n153 240.244
R12774 gnd.n7254 gnd.n153 240.244
R12775 gnd.n7254 gnd.n158 240.244
R12776 gnd.n7246 gnd.n158 240.244
R12777 gnd.n2284 gnd.n2242 240.244
R12778 gnd.n3661 gnd.n3660 240.244
R12779 gnd.n3657 gnd.n3656 240.244
R12780 gnd.n3653 gnd.n3652 240.244
R12781 gnd.n3649 gnd.n3648 240.244
R12782 gnd.n3645 gnd.n3644 240.244
R12783 gnd.n3641 gnd.n3640 240.244
R12784 gnd.n3637 gnd.n3636 240.244
R12785 gnd.n3633 gnd.n3632 240.244
R12786 gnd.n3629 gnd.n3628 240.244
R12787 gnd.n3625 gnd.n3624 240.244
R12788 gnd.n3621 gnd.n3620 240.244
R12789 gnd.n3617 gnd.n3616 240.244
R12790 gnd.n2858 gnd.n2755 240.244
R12791 gnd.n2858 gnd.n2748 240.244
R12792 gnd.n2869 gnd.n2748 240.244
R12793 gnd.n2869 gnd.n2744 240.244
R12794 gnd.n2875 gnd.n2744 240.244
R12795 gnd.n2875 gnd.n2736 240.244
R12796 gnd.n2885 gnd.n2736 240.244
R12797 gnd.n2885 gnd.n2731 240.244
R12798 gnd.n2921 gnd.n2731 240.244
R12799 gnd.n2921 gnd.n2732 240.244
R12800 gnd.n2732 gnd.n2679 240.244
R12801 gnd.n2916 gnd.n2679 240.244
R12802 gnd.n2916 gnd.n2915 240.244
R12803 gnd.n2915 gnd.n2658 240.244
R12804 gnd.n2911 gnd.n2658 240.244
R12805 gnd.n2911 gnd.n2649 240.244
R12806 gnd.n2908 gnd.n2649 240.244
R12807 gnd.n2908 gnd.n2907 240.244
R12808 gnd.n2907 gnd.n2632 240.244
R12809 gnd.n2903 gnd.n2632 240.244
R12810 gnd.n2903 gnd.n2621 240.244
R12811 gnd.n2621 gnd.n2602 240.244
R12812 gnd.n3016 gnd.n2602 240.244
R12813 gnd.n3016 gnd.n2598 240.244
R12814 gnd.n3024 gnd.n2598 240.244
R12815 gnd.n3024 gnd.n2589 240.244
R12816 gnd.n2589 gnd.n2525 240.244
R12817 gnd.n3096 gnd.n2525 240.244
R12818 gnd.n3096 gnd.n2526 240.244
R12819 gnd.n2537 gnd.n2526 240.244
R12820 gnd.n2572 gnd.n2537 240.244
R12821 gnd.n2575 gnd.n2572 240.244
R12822 gnd.n2575 gnd.n2549 240.244
R12823 gnd.n2562 gnd.n2549 240.244
R12824 gnd.n2562 gnd.n2559 240.244
R12825 gnd.n2559 gnd.n2468 240.244
R12826 gnd.n3117 gnd.n2468 240.244
R12827 gnd.n3117 gnd.n2458 240.244
R12828 gnd.n3113 gnd.n2458 240.244
R12829 gnd.n3113 gnd.n2452 240.244
R12830 gnd.n3110 gnd.n2452 240.244
R12831 gnd.n3110 gnd.n2441 240.244
R12832 gnd.n3107 gnd.n2441 240.244
R12833 gnd.n3107 gnd.n2419 240.244
R12834 gnd.n3183 gnd.n2419 240.244
R12835 gnd.n3183 gnd.n2415 240.244
R12836 gnd.n3204 gnd.n2415 240.244
R12837 gnd.n3204 gnd.n2404 240.244
R12838 gnd.n3200 gnd.n2404 240.244
R12839 gnd.n3200 gnd.n2397 240.244
R12840 gnd.n3197 gnd.n2397 240.244
R12841 gnd.n3197 gnd.n2386 240.244
R12842 gnd.n3194 gnd.n2386 240.244
R12843 gnd.n3194 gnd.n2363 240.244
R12844 gnd.n3268 gnd.n2363 240.244
R12845 gnd.n3268 gnd.n2359 240.244
R12846 gnd.n3293 gnd.n2359 240.244
R12847 gnd.n3293 gnd.n2350 240.244
R12848 gnd.n3289 gnd.n2350 240.244
R12849 gnd.n3289 gnd.n2343 240.244
R12850 gnd.n3285 gnd.n2343 240.244
R12851 gnd.n3285 gnd.n2332 240.244
R12852 gnd.n3282 gnd.n2332 240.244
R12853 gnd.n3282 gnd.n2313 240.244
R12854 gnd.n3612 gnd.n2313 240.244
R12855 gnd.n2772 gnd.n2771 240.244
R12856 gnd.n2843 gnd.n2771 240.244
R12857 gnd.n2841 gnd.n2840 240.244
R12858 gnd.n2837 gnd.n2836 240.244
R12859 gnd.n2833 gnd.n2832 240.244
R12860 gnd.n2829 gnd.n2828 240.244
R12861 gnd.n2825 gnd.n2824 240.244
R12862 gnd.n2821 gnd.n2820 240.244
R12863 gnd.n2817 gnd.n2816 240.244
R12864 gnd.n2813 gnd.n2812 240.244
R12865 gnd.n2809 gnd.n2808 240.244
R12866 gnd.n2805 gnd.n2804 240.244
R12867 gnd.n2801 gnd.n2759 240.244
R12868 gnd.n2861 gnd.n2753 240.244
R12869 gnd.n2861 gnd.n2749 240.244
R12870 gnd.n2867 gnd.n2749 240.244
R12871 gnd.n2867 gnd.n2742 240.244
R12872 gnd.n2877 gnd.n2742 240.244
R12873 gnd.n2877 gnd.n2738 240.244
R12874 gnd.n2883 gnd.n2738 240.244
R12875 gnd.n2883 gnd.n2729 240.244
R12876 gnd.n2923 gnd.n2729 240.244
R12877 gnd.n2923 gnd.n2680 240.244
R12878 gnd.n2931 gnd.n2680 240.244
R12879 gnd.n2931 gnd.n2681 240.244
R12880 gnd.n2681 gnd.n2659 240.244
R12881 gnd.n2952 gnd.n2659 240.244
R12882 gnd.n2952 gnd.n2651 240.244
R12883 gnd.n2963 gnd.n2651 240.244
R12884 gnd.n2963 gnd.n2652 240.244
R12885 gnd.n2652 gnd.n2633 240.244
R12886 gnd.n2983 gnd.n2633 240.244
R12887 gnd.n2983 gnd.n2623 240.244
R12888 gnd.n2993 gnd.n2623 240.244
R12889 gnd.n2993 gnd.n2604 240.244
R12890 gnd.n3014 gnd.n2604 240.244
R12891 gnd.n3014 gnd.n2606 240.244
R12892 gnd.n2606 gnd.n2587 240.244
R12893 gnd.n3042 gnd.n2587 240.244
R12894 gnd.n3042 gnd.n2529 240.244
R12895 gnd.n3094 gnd.n2529 240.244
R12896 gnd.n3094 gnd.n2530 240.244
R12897 gnd.n3090 gnd.n2530 240.244
R12898 gnd.n3090 gnd.n2536 240.244
R12899 gnd.n2551 gnd.n2536 240.244
R12900 gnd.n3080 gnd.n2551 240.244
R12901 gnd.n3080 gnd.n2552 240.244
R12902 gnd.n3076 gnd.n2552 240.244
R12903 gnd.n3076 gnd.n2558 240.244
R12904 gnd.n2558 gnd.n2457 240.244
R12905 gnd.n3133 gnd.n2457 240.244
R12906 gnd.n3133 gnd.n2450 240.244
R12907 gnd.n3144 gnd.n2450 240.244
R12908 gnd.n3144 gnd.n2443 240.244
R12909 gnd.n3159 gnd.n2443 240.244
R12910 gnd.n3159 gnd.n2444 240.244
R12911 gnd.n2444 gnd.n2422 240.244
R12912 gnd.n3181 gnd.n2422 240.244
R12913 gnd.n3181 gnd.n2423 240.244
R12914 gnd.n2423 gnd.n2402 240.244
R12915 gnd.n3218 gnd.n2402 240.244
R12916 gnd.n3218 gnd.n2395 240.244
R12917 gnd.n3229 gnd.n2395 240.244
R12918 gnd.n3229 gnd.n2388 240.244
R12919 gnd.n3244 gnd.n2388 240.244
R12920 gnd.n3244 gnd.n2389 240.244
R12921 gnd.n2389 gnd.n2366 240.244
R12922 gnd.n3266 gnd.n2366 240.244
R12923 gnd.n3266 gnd.n2368 240.244
R12924 gnd.n2368 gnd.n2348 240.244
R12925 gnd.n3307 gnd.n2348 240.244
R12926 gnd.n3307 gnd.n2341 240.244
R12927 gnd.n3318 gnd.n2341 240.244
R12928 gnd.n3318 gnd.n2334 240.244
R12929 gnd.n3587 gnd.n2334 240.244
R12930 gnd.n3587 gnd.n2335 240.244
R12931 gnd.n2335 gnd.n2316 240.244
R12932 gnd.n3610 gnd.n2316 240.244
R12933 gnd.n910 gnd.n863 240.244
R12934 gnd.n967 gnd.n911 240.244
R12935 gnd.n921 gnd.n920 240.244
R12936 gnd.n969 gnd.n928 240.244
R12937 gnd.n972 gnd.n929 240.244
R12938 gnd.n939 gnd.n938 240.244
R12939 gnd.n974 gnd.n946 240.244
R12940 gnd.n977 gnd.n947 240.244
R12941 gnd.n964 gnd.n959 240.244
R12942 gnd.n3779 gnd.n3705 240.244
R12943 gnd.n3779 gnd.n2231 240.244
R12944 gnd.n2231 gnd.n2220 240.244
R12945 gnd.n4026 gnd.n2220 240.244
R12946 gnd.n4026 gnd.n2216 240.244
R12947 gnd.n4034 gnd.n2216 240.244
R12948 gnd.n4034 gnd.n2206 240.244
R12949 gnd.n2206 gnd.n2195 240.244
R12950 gnd.n4061 gnd.n2195 240.244
R12951 gnd.n4061 gnd.n2191 240.244
R12952 gnd.n4071 gnd.n2191 240.244
R12953 gnd.n4071 gnd.n2179 240.244
R12954 gnd.n2179 gnd.n2169 240.244
R12955 gnd.n4100 gnd.n2169 240.244
R12956 gnd.n4101 gnd.n4100 240.244
R12957 gnd.n4101 gnd.n735 240.244
R12958 gnd.n4107 gnd.n735 240.244
R12959 gnd.n4107 gnd.n746 240.244
R12960 gnd.n4127 gnd.n746 240.244
R12961 gnd.n4127 gnd.n757 240.244
R12962 gnd.n4133 gnd.n757 240.244
R12963 gnd.n4133 gnd.n765 240.244
R12964 gnd.n4152 gnd.n765 240.244
R12965 gnd.n4152 gnd.n774 240.244
R12966 gnd.n4146 gnd.n774 240.244
R12967 gnd.n4146 gnd.n782 240.244
R12968 gnd.n4172 gnd.n782 240.244
R12969 gnd.n4172 gnd.n791 240.244
R12970 gnd.n4178 gnd.n791 240.244
R12971 gnd.n4178 gnd.n802 240.244
R12972 gnd.n4218 gnd.n802 240.244
R12973 gnd.n4218 gnd.n811 240.244
R12974 gnd.n2138 gnd.n811 240.244
R12975 gnd.n2138 gnd.n822 240.244
R12976 gnd.n2139 gnd.n822 240.244
R12977 gnd.n2139 gnd.n831 240.244
R12978 gnd.n2142 gnd.n831 240.244
R12979 gnd.n2142 gnd.n842 240.244
R12980 gnd.n4203 gnd.n842 240.244
R12981 gnd.n4203 gnd.n852 240.244
R12982 gnd.n5977 gnd.n852 240.244
R12983 gnd.n5977 gnd.n861 240.244
R12984 gnd.n3732 gnd.n3730 240.244
R12985 gnd.n3738 gnd.n3723 240.244
R12986 gnd.n3742 gnd.n3740 240.244
R12987 gnd.n3748 gnd.n3719 240.244
R12988 gnd.n3752 gnd.n3750 240.244
R12989 gnd.n3758 gnd.n3715 240.244
R12990 gnd.n3762 gnd.n3760 240.244
R12991 gnd.n3768 gnd.n3711 240.244
R12992 gnd.n3771 gnd.n3770 240.244
R12993 gnd.n3998 gnd.n2232 240.244
R12994 gnd.n4014 gnd.n2232 240.244
R12995 gnd.n4014 gnd.n2233 240.244
R12996 gnd.n2233 gnd.n2223 240.244
R12997 gnd.n4009 gnd.n2223 240.244
R12998 gnd.n4009 gnd.n2207 240.244
R12999 gnd.n4049 gnd.n2207 240.244
R13000 gnd.n4049 gnd.n2208 240.244
R13001 gnd.n2208 gnd.n2198 240.244
R13002 gnd.n4044 gnd.n2198 240.244
R13003 gnd.n4044 gnd.n2181 240.244
R13004 gnd.n4089 gnd.n2181 240.244
R13005 gnd.n4089 gnd.n2182 240.244
R13006 gnd.n2182 gnd.n2172 240.244
R13007 gnd.n4084 gnd.n2172 240.244
R13008 gnd.n4084 gnd.n737 240.244
R13009 gnd.n748 gnd.n737 240.244
R13010 gnd.n6058 gnd.n748 240.244
R13011 gnd.n6058 gnd.n749 240.244
R13012 gnd.n6054 gnd.n749 240.244
R13013 gnd.n6054 gnd.n755 240.244
R13014 gnd.n6045 gnd.n755 240.244
R13015 gnd.n6045 gnd.n766 240.244
R13016 gnd.n6041 gnd.n766 240.244
R13017 gnd.n6041 gnd.n771 240.244
R13018 gnd.n6032 gnd.n771 240.244
R13019 gnd.n6032 gnd.n784 240.244
R13020 gnd.n6028 gnd.n784 240.244
R13021 gnd.n6028 gnd.n789 240.244
R13022 gnd.n6020 gnd.n789 240.244
R13023 gnd.n6020 gnd.n803 240.244
R13024 gnd.n6016 gnd.n803 240.244
R13025 gnd.n6016 gnd.n808 240.244
R13026 gnd.n6008 gnd.n808 240.244
R13027 gnd.n6008 gnd.n824 240.244
R13028 gnd.n6004 gnd.n824 240.244
R13029 gnd.n6004 gnd.n829 240.244
R13030 gnd.n5996 gnd.n829 240.244
R13031 gnd.n5996 gnd.n844 240.244
R13032 gnd.n5992 gnd.n844 240.244
R13033 gnd.n5992 gnd.n849 240.244
R13034 gnd.n5984 gnd.n849 240.244
R13035 gnd.n6244 gnd.n560 240.244
R13036 gnd.n6248 gnd.n560 240.244
R13037 gnd.n6248 gnd.n556 240.244
R13038 gnd.n6254 gnd.n556 240.244
R13039 gnd.n6254 gnd.n554 240.244
R13040 gnd.n6258 gnd.n554 240.244
R13041 gnd.n6258 gnd.n550 240.244
R13042 gnd.n6264 gnd.n550 240.244
R13043 gnd.n6264 gnd.n548 240.244
R13044 gnd.n6268 gnd.n548 240.244
R13045 gnd.n6268 gnd.n544 240.244
R13046 gnd.n6274 gnd.n544 240.244
R13047 gnd.n6274 gnd.n542 240.244
R13048 gnd.n6278 gnd.n542 240.244
R13049 gnd.n6278 gnd.n538 240.244
R13050 gnd.n6284 gnd.n538 240.244
R13051 gnd.n6284 gnd.n536 240.244
R13052 gnd.n6288 gnd.n536 240.244
R13053 gnd.n6288 gnd.n532 240.244
R13054 gnd.n6294 gnd.n532 240.244
R13055 gnd.n6294 gnd.n530 240.244
R13056 gnd.n6298 gnd.n530 240.244
R13057 gnd.n6298 gnd.n526 240.244
R13058 gnd.n6304 gnd.n526 240.244
R13059 gnd.n6304 gnd.n524 240.244
R13060 gnd.n6308 gnd.n524 240.244
R13061 gnd.n6308 gnd.n520 240.244
R13062 gnd.n6314 gnd.n520 240.244
R13063 gnd.n6314 gnd.n518 240.244
R13064 gnd.n6318 gnd.n518 240.244
R13065 gnd.n6318 gnd.n514 240.244
R13066 gnd.n6324 gnd.n514 240.244
R13067 gnd.n6324 gnd.n512 240.244
R13068 gnd.n6328 gnd.n512 240.244
R13069 gnd.n6328 gnd.n508 240.244
R13070 gnd.n6334 gnd.n508 240.244
R13071 gnd.n6334 gnd.n506 240.244
R13072 gnd.n6338 gnd.n506 240.244
R13073 gnd.n6338 gnd.n502 240.244
R13074 gnd.n6344 gnd.n502 240.244
R13075 gnd.n6344 gnd.n500 240.244
R13076 gnd.n6348 gnd.n500 240.244
R13077 gnd.n6348 gnd.n496 240.244
R13078 gnd.n6354 gnd.n496 240.244
R13079 gnd.n6354 gnd.n494 240.244
R13080 gnd.n6358 gnd.n494 240.244
R13081 gnd.n6358 gnd.n490 240.244
R13082 gnd.n6364 gnd.n490 240.244
R13083 gnd.n6364 gnd.n488 240.244
R13084 gnd.n6368 gnd.n488 240.244
R13085 gnd.n6368 gnd.n484 240.244
R13086 gnd.n6374 gnd.n484 240.244
R13087 gnd.n6374 gnd.n482 240.244
R13088 gnd.n6378 gnd.n482 240.244
R13089 gnd.n6378 gnd.n478 240.244
R13090 gnd.n6384 gnd.n478 240.244
R13091 gnd.n6384 gnd.n476 240.244
R13092 gnd.n6388 gnd.n476 240.244
R13093 gnd.n6388 gnd.n472 240.244
R13094 gnd.n6394 gnd.n472 240.244
R13095 gnd.n6394 gnd.n470 240.244
R13096 gnd.n6398 gnd.n470 240.244
R13097 gnd.n6398 gnd.n466 240.244
R13098 gnd.n6404 gnd.n466 240.244
R13099 gnd.n6404 gnd.n464 240.244
R13100 gnd.n6408 gnd.n464 240.244
R13101 gnd.n6408 gnd.n460 240.244
R13102 gnd.n6414 gnd.n460 240.244
R13103 gnd.n6414 gnd.n458 240.244
R13104 gnd.n6418 gnd.n458 240.244
R13105 gnd.n6418 gnd.n454 240.244
R13106 gnd.n6424 gnd.n454 240.244
R13107 gnd.n6424 gnd.n452 240.244
R13108 gnd.n6428 gnd.n452 240.244
R13109 gnd.n6428 gnd.n448 240.244
R13110 gnd.n6434 gnd.n448 240.244
R13111 gnd.n6434 gnd.n446 240.244
R13112 gnd.n6438 gnd.n446 240.244
R13113 gnd.n6438 gnd.n442 240.244
R13114 gnd.n6444 gnd.n442 240.244
R13115 gnd.n6444 gnd.n440 240.244
R13116 gnd.n6448 gnd.n440 240.244
R13117 gnd.n6448 gnd.n436 240.244
R13118 gnd.n6454 gnd.n436 240.244
R13119 gnd.n6454 gnd.n434 240.244
R13120 gnd.n6458 gnd.n434 240.244
R13121 gnd.n6458 gnd.n430 240.244
R13122 gnd.n6464 gnd.n430 240.244
R13123 gnd.n6464 gnd.n428 240.244
R13124 gnd.n6468 gnd.n428 240.244
R13125 gnd.n6468 gnd.n424 240.244
R13126 gnd.n6474 gnd.n424 240.244
R13127 gnd.n6474 gnd.n422 240.244
R13128 gnd.n6478 gnd.n422 240.244
R13129 gnd.n6478 gnd.n418 240.244
R13130 gnd.n6484 gnd.n418 240.244
R13131 gnd.n6484 gnd.n416 240.244
R13132 gnd.n6488 gnd.n416 240.244
R13133 gnd.n6488 gnd.n412 240.244
R13134 gnd.n6494 gnd.n412 240.244
R13135 gnd.n6494 gnd.n410 240.244
R13136 gnd.n6498 gnd.n410 240.244
R13137 gnd.n6498 gnd.n406 240.244
R13138 gnd.n6504 gnd.n406 240.244
R13139 gnd.n6504 gnd.n404 240.244
R13140 gnd.n6508 gnd.n404 240.244
R13141 gnd.n6508 gnd.n400 240.244
R13142 gnd.n6514 gnd.n400 240.244
R13143 gnd.n6514 gnd.n398 240.244
R13144 gnd.n6518 gnd.n398 240.244
R13145 gnd.n6518 gnd.n394 240.244
R13146 gnd.n6524 gnd.n394 240.244
R13147 gnd.n6524 gnd.n392 240.244
R13148 gnd.n6528 gnd.n392 240.244
R13149 gnd.n6528 gnd.n388 240.244
R13150 gnd.n6534 gnd.n388 240.244
R13151 gnd.n6534 gnd.n386 240.244
R13152 gnd.n6538 gnd.n386 240.244
R13153 gnd.n6538 gnd.n382 240.244
R13154 gnd.n6544 gnd.n382 240.244
R13155 gnd.n6544 gnd.n380 240.244
R13156 gnd.n6548 gnd.n380 240.244
R13157 gnd.n6548 gnd.n376 240.244
R13158 gnd.n6554 gnd.n376 240.244
R13159 gnd.n6554 gnd.n374 240.244
R13160 gnd.n6558 gnd.n374 240.244
R13161 gnd.n6558 gnd.n370 240.244
R13162 gnd.n6564 gnd.n370 240.244
R13163 gnd.n6564 gnd.n368 240.244
R13164 gnd.n6568 gnd.n368 240.244
R13165 gnd.n6568 gnd.n364 240.244
R13166 gnd.n6574 gnd.n364 240.244
R13167 gnd.n6574 gnd.n362 240.244
R13168 gnd.n6578 gnd.n362 240.244
R13169 gnd.n6578 gnd.n358 240.244
R13170 gnd.n6584 gnd.n358 240.244
R13171 gnd.n6584 gnd.n356 240.244
R13172 gnd.n6588 gnd.n356 240.244
R13173 gnd.n6588 gnd.n352 240.244
R13174 gnd.n6594 gnd.n352 240.244
R13175 gnd.n6594 gnd.n350 240.244
R13176 gnd.n6598 gnd.n350 240.244
R13177 gnd.n6598 gnd.n346 240.244
R13178 gnd.n6604 gnd.n346 240.244
R13179 gnd.n6604 gnd.n344 240.244
R13180 gnd.n6608 gnd.n344 240.244
R13181 gnd.n6608 gnd.n340 240.244
R13182 gnd.n6614 gnd.n340 240.244
R13183 gnd.n6614 gnd.n338 240.244
R13184 gnd.n6618 gnd.n338 240.244
R13185 gnd.n6618 gnd.n334 240.244
R13186 gnd.n6624 gnd.n334 240.244
R13187 gnd.n6624 gnd.n332 240.244
R13188 gnd.n6628 gnd.n332 240.244
R13189 gnd.n6628 gnd.n328 240.244
R13190 gnd.n6634 gnd.n328 240.244
R13191 gnd.n6634 gnd.n326 240.244
R13192 gnd.n6638 gnd.n326 240.244
R13193 gnd.n6638 gnd.n322 240.244
R13194 gnd.n6644 gnd.n322 240.244
R13195 gnd.n6644 gnd.n320 240.244
R13196 gnd.n6648 gnd.n320 240.244
R13197 gnd.n6648 gnd.n316 240.244
R13198 gnd.n6655 gnd.n316 240.244
R13199 gnd.n6655 gnd.n314 240.244
R13200 gnd.n6659 gnd.n314 240.244
R13201 gnd.n6659 gnd.n311 240.244
R13202 gnd.n6665 gnd.n309 240.244
R13203 gnd.n6669 gnd.n309 240.244
R13204 gnd.n6669 gnd.n305 240.244
R13205 gnd.n6675 gnd.n305 240.244
R13206 gnd.n6675 gnd.n303 240.244
R13207 gnd.n6679 gnd.n303 240.244
R13208 gnd.n6679 gnd.n299 240.244
R13209 gnd.n6685 gnd.n299 240.244
R13210 gnd.n6685 gnd.n297 240.244
R13211 gnd.n6689 gnd.n297 240.244
R13212 gnd.n6689 gnd.n293 240.244
R13213 gnd.n6695 gnd.n293 240.244
R13214 gnd.n6695 gnd.n291 240.244
R13215 gnd.n6699 gnd.n291 240.244
R13216 gnd.n6699 gnd.n287 240.244
R13217 gnd.n6705 gnd.n287 240.244
R13218 gnd.n6705 gnd.n285 240.244
R13219 gnd.n6709 gnd.n285 240.244
R13220 gnd.n6709 gnd.n281 240.244
R13221 gnd.n6715 gnd.n281 240.244
R13222 gnd.n6715 gnd.n279 240.244
R13223 gnd.n6719 gnd.n279 240.244
R13224 gnd.n6719 gnd.n275 240.244
R13225 gnd.n6725 gnd.n275 240.244
R13226 gnd.n6725 gnd.n273 240.244
R13227 gnd.n6729 gnd.n273 240.244
R13228 gnd.n6729 gnd.n269 240.244
R13229 gnd.n6735 gnd.n269 240.244
R13230 gnd.n6735 gnd.n267 240.244
R13231 gnd.n6739 gnd.n267 240.244
R13232 gnd.n6739 gnd.n263 240.244
R13233 gnd.n6745 gnd.n263 240.244
R13234 gnd.n6745 gnd.n261 240.244
R13235 gnd.n6749 gnd.n261 240.244
R13236 gnd.n6749 gnd.n257 240.244
R13237 gnd.n6755 gnd.n257 240.244
R13238 gnd.n6755 gnd.n255 240.244
R13239 gnd.n6759 gnd.n255 240.244
R13240 gnd.n6759 gnd.n251 240.244
R13241 gnd.n6765 gnd.n251 240.244
R13242 gnd.n6765 gnd.n249 240.244
R13243 gnd.n6769 gnd.n249 240.244
R13244 gnd.n6769 gnd.n245 240.244
R13245 gnd.n6775 gnd.n245 240.244
R13246 gnd.n6775 gnd.n243 240.244
R13247 gnd.n6779 gnd.n243 240.244
R13248 gnd.n6779 gnd.n239 240.244
R13249 gnd.n6785 gnd.n239 240.244
R13250 gnd.n6785 gnd.n237 240.244
R13251 gnd.n6789 gnd.n237 240.244
R13252 gnd.n6789 gnd.n233 240.244
R13253 gnd.n6795 gnd.n233 240.244
R13254 gnd.n6795 gnd.n231 240.244
R13255 gnd.n6799 gnd.n231 240.244
R13256 gnd.n6799 gnd.n227 240.244
R13257 gnd.n6805 gnd.n227 240.244
R13258 gnd.n6805 gnd.n225 240.244
R13259 gnd.n6809 gnd.n225 240.244
R13260 gnd.n6809 gnd.n221 240.244
R13261 gnd.n6815 gnd.n221 240.244
R13262 gnd.n6815 gnd.n219 240.244
R13263 gnd.n6819 gnd.n219 240.244
R13264 gnd.n6819 gnd.n215 240.244
R13265 gnd.n6825 gnd.n215 240.244
R13266 gnd.n6825 gnd.n213 240.244
R13267 gnd.n6829 gnd.n213 240.244
R13268 gnd.n6829 gnd.n209 240.244
R13269 gnd.n6835 gnd.n209 240.244
R13270 gnd.n6835 gnd.n207 240.244
R13271 gnd.n6839 gnd.n207 240.244
R13272 gnd.n6839 gnd.n203 240.244
R13273 gnd.n6845 gnd.n203 240.244
R13274 gnd.n6845 gnd.n201 240.244
R13275 gnd.n6849 gnd.n201 240.244
R13276 gnd.n6849 gnd.n197 240.244
R13277 gnd.n6855 gnd.n197 240.244
R13278 gnd.n6855 gnd.n195 240.244
R13279 gnd.n6859 gnd.n195 240.244
R13280 gnd.n6859 gnd.n191 240.244
R13281 gnd.n6865 gnd.n191 240.244
R13282 gnd.n6865 gnd.n189 240.244
R13283 gnd.n6870 gnd.n189 240.244
R13284 gnd.n6870 gnd.n185 240.244
R13285 gnd.n6876 gnd.n185 240.244
R13286 gnd.n6068 gnd.n732 240.244
R13287 gnd.n4117 gnd.n732 240.244
R13288 gnd.n4117 gnd.n4114 240.244
R13289 gnd.n4124 gnd.n4114 240.244
R13290 gnd.n4124 gnd.n4115 240.244
R13291 gnd.n4115 gnd.n2154 240.244
R13292 gnd.n4155 gnd.n2154 240.244
R13293 gnd.n4155 gnd.n2152 240.244
R13294 gnd.n4160 gnd.n2152 240.244
R13295 gnd.n4161 gnd.n4160 240.244
R13296 gnd.n4161 gnd.n2149 240.244
R13297 gnd.n4169 gnd.n2149 240.244
R13298 gnd.n4169 gnd.n2150 240.244
R13299 gnd.n2150 gnd.n2132 240.244
R13300 gnd.n4221 gnd.n2132 240.244
R13301 gnd.n4221 gnd.n2128 240.244
R13302 gnd.n4227 gnd.n2128 240.244
R13303 gnd.n4228 gnd.n4227 240.244
R13304 gnd.n4229 gnd.n4228 240.244
R13305 gnd.n4229 gnd.n2124 240.244
R13306 gnd.n4235 gnd.n2124 240.244
R13307 gnd.n4236 gnd.n4235 240.244
R13308 gnd.n4237 gnd.n4236 240.244
R13309 gnd.n4237 gnd.n2120 240.244
R13310 gnd.n4243 gnd.n2120 240.244
R13311 gnd.n4244 gnd.n4243 240.244
R13312 gnd.n4245 gnd.n4244 240.244
R13313 gnd.n4245 gnd.n2116 240.244
R13314 gnd.n4251 gnd.n2116 240.244
R13315 gnd.n4253 gnd.n4251 240.244
R13316 gnd.n4254 gnd.n4253 240.244
R13317 gnd.n4254 gnd.n2112 240.244
R13318 gnd.n4260 gnd.n2112 240.244
R13319 gnd.n4260 gnd.n2110 240.244
R13320 gnd.n4322 gnd.n2110 240.244
R13321 gnd.n4322 gnd.n2106 240.244
R13322 gnd.n4328 gnd.n2106 240.244
R13323 gnd.n4328 gnd.n2096 240.244
R13324 gnd.n4338 gnd.n2096 240.244
R13325 gnd.n4338 gnd.n2092 240.244
R13326 gnd.n4344 gnd.n2092 240.244
R13327 gnd.n4344 gnd.n2081 240.244
R13328 gnd.n4354 gnd.n2081 240.244
R13329 gnd.n4354 gnd.n2077 240.244
R13330 gnd.n4360 gnd.n2077 240.244
R13331 gnd.n4360 gnd.n2067 240.244
R13332 gnd.n4370 gnd.n2067 240.244
R13333 gnd.n4370 gnd.n2063 240.244
R13334 gnd.n4376 gnd.n2063 240.244
R13335 gnd.n4376 gnd.n2052 240.244
R13336 gnd.n4400 gnd.n2052 240.244
R13337 gnd.n4400 gnd.n2047 240.244
R13338 gnd.n4412 gnd.n2047 240.244
R13339 gnd.n4412 gnd.n2048 240.244
R13340 gnd.n4408 gnd.n2048 240.244
R13341 gnd.n4408 gnd.n1205 240.244
R13342 gnd.n5776 gnd.n1205 240.244
R13343 gnd.n5776 gnd.n1206 240.244
R13344 gnd.n5772 gnd.n1206 240.244
R13345 gnd.n5772 gnd.n1212 240.244
R13346 gnd.n4558 gnd.n1212 240.244
R13347 gnd.n4564 gnd.n4558 240.244
R13348 gnd.n4564 gnd.n2022 240.244
R13349 gnd.n4587 gnd.n2022 240.244
R13350 gnd.n4587 gnd.n2017 240.244
R13351 gnd.n4595 gnd.n2017 240.244
R13352 gnd.n4595 gnd.n2018 240.244
R13353 gnd.n2018 gnd.n1994 240.244
R13354 gnd.n4625 gnd.n1994 240.244
R13355 gnd.n4625 gnd.n1989 240.244
R13356 gnd.n4637 gnd.n1989 240.244
R13357 gnd.n4637 gnd.n1990 240.244
R13358 gnd.n4633 gnd.n1990 240.244
R13359 gnd.n4633 gnd.n1963 240.244
R13360 gnd.n4698 gnd.n1963 240.244
R13361 gnd.n4698 gnd.n1964 240.244
R13362 gnd.n4694 gnd.n1964 240.244
R13363 gnd.n4694 gnd.n1944 240.244
R13364 gnd.n4726 gnd.n1944 240.244
R13365 gnd.n4726 gnd.n1939 240.244
R13366 gnd.n4734 gnd.n1939 240.244
R13367 gnd.n4734 gnd.n1940 240.244
R13368 gnd.n1940 gnd.n1916 240.244
R13369 gnd.n4764 gnd.n1916 240.244
R13370 gnd.n4764 gnd.n1912 240.244
R13371 gnd.n4770 gnd.n1912 240.244
R13372 gnd.n4770 gnd.n1890 240.244
R13373 gnd.n4801 gnd.n1890 240.244
R13374 gnd.n4801 gnd.n1885 240.244
R13375 gnd.n4809 gnd.n1885 240.244
R13376 gnd.n4809 gnd.n1886 240.244
R13377 gnd.n1886 gnd.n1863 240.244
R13378 gnd.n4850 gnd.n1863 240.244
R13379 gnd.n4850 gnd.n1858 240.244
R13380 gnd.n4858 gnd.n1858 240.244
R13381 gnd.n4858 gnd.n1859 240.244
R13382 gnd.n1859 gnd.n1841 240.244
R13383 gnd.n4891 gnd.n1841 240.244
R13384 gnd.n4891 gnd.n1836 240.244
R13385 gnd.n4899 gnd.n1836 240.244
R13386 gnd.n4899 gnd.n1837 240.244
R13387 gnd.n1837 gnd.n1811 240.244
R13388 gnd.n4931 gnd.n1811 240.244
R13389 gnd.n4931 gnd.n1807 240.244
R13390 gnd.n4937 gnd.n1807 240.244
R13391 gnd.n4937 gnd.n1787 240.244
R13392 gnd.n4974 gnd.n1787 240.244
R13393 gnd.n4974 gnd.n1782 240.244
R13394 gnd.n4982 gnd.n1782 240.244
R13395 gnd.n4982 gnd.n1783 240.244
R13396 gnd.n1783 gnd.n1731 240.244
R13397 gnd.n5150 gnd.n1731 240.244
R13398 gnd.n5150 gnd.n1727 240.244
R13399 gnd.n5156 gnd.n1727 240.244
R13400 gnd.n5156 gnd.n1720 240.244
R13401 gnd.n5167 gnd.n1720 240.244
R13402 gnd.n5167 gnd.n1716 240.244
R13403 gnd.n5173 gnd.n1716 240.244
R13404 gnd.n5173 gnd.n1708 240.244
R13405 gnd.n5184 gnd.n1708 240.244
R13406 gnd.n5184 gnd.n1704 240.244
R13407 gnd.n5190 gnd.n1704 240.244
R13408 gnd.n5190 gnd.n1696 240.244
R13409 gnd.n5201 gnd.n1696 240.244
R13410 gnd.n5201 gnd.n1692 240.244
R13411 gnd.n5207 gnd.n1692 240.244
R13412 gnd.n5207 gnd.n1684 240.244
R13413 gnd.n5218 gnd.n1684 240.244
R13414 gnd.n5218 gnd.n1680 240.244
R13415 gnd.n5227 gnd.n1680 240.244
R13416 gnd.n5227 gnd.n1672 240.244
R13417 gnd.n5238 gnd.n1672 240.244
R13418 gnd.n5239 gnd.n5238 240.244
R13419 gnd.n5239 gnd.n1313 240.244
R13420 gnd.n1667 gnd.n1313 240.244
R13421 gnd.n5257 gnd.n1667 240.244
R13422 gnd.n5257 gnd.n1668 240.244
R13423 gnd.n5253 gnd.n1668 240.244
R13424 gnd.n5253 gnd.n5252 240.244
R13425 gnd.n5252 gnd.n5251 240.244
R13426 gnd.n5251 gnd.n1636 240.244
R13427 gnd.n5309 gnd.n1636 240.244
R13428 gnd.n5309 gnd.n1632 240.244
R13429 gnd.n5315 gnd.n1632 240.244
R13430 gnd.n5316 gnd.n5315 240.244
R13431 gnd.n5317 gnd.n5316 240.244
R13432 gnd.n5317 gnd.n1628 240.244
R13433 gnd.n5323 gnd.n1628 240.244
R13434 gnd.n5324 gnd.n5323 240.244
R13435 gnd.n5325 gnd.n5324 240.244
R13436 gnd.n5325 gnd.n1623 240.244
R13437 gnd.n5348 gnd.n1623 240.244
R13438 gnd.n5348 gnd.n1624 240.244
R13439 gnd.n5344 gnd.n1624 240.244
R13440 gnd.n5344 gnd.n5343 240.244
R13441 gnd.n5343 gnd.n5342 240.244
R13442 gnd.n5342 gnd.n5333 240.244
R13443 gnd.n5337 gnd.n5333 240.244
R13444 gnd.n5337 gnd.n1594 240.244
R13445 gnd.n5402 gnd.n1594 240.244
R13446 gnd.n5402 gnd.n1595 240.244
R13447 gnd.n5397 gnd.n1595 240.244
R13448 gnd.n5397 gnd.n1599 240.244
R13449 gnd.n1599 gnd.n181 240.244
R13450 gnd.n6882 gnd.n181 240.244
R13451 gnd.n6882 gnd.n182 240.244
R13452 gnd.n6877 gnd.n182 240.244
R13453 gnd.n6238 gnd.n562 240.244
R13454 gnd.n6238 gnd.n565 240.244
R13455 gnd.n6234 gnd.n565 240.244
R13456 gnd.n6234 gnd.n567 240.244
R13457 gnd.n6230 gnd.n567 240.244
R13458 gnd.n6230 gnd.n573 240.244
R13459 gnd.n6226 gnd.n573 240.244
R13460 gnd.n6226 gnd.n575 240.244
R13461 gnd.n6222 gnd.n575 240.244
R13462 gnd.n6222 gnd.n581 240.244
R13463 gnd.n6218 gnd.n581 240.244
R13464 gnd.n6218 gnd.n583 240.244
R13465 gnd.n6214 gnd.n583 240.244
R13466 gnd.n6214 gnd.n589 240.244
R13467 gnd.n6210 gnd.n589 240.244
R13468 gnd.n6210 gnd.n591 240.244
R13469 gnd.n6206 gnd.n591 240.244
R13470 gnd.n6206 gnd.n597 240.244
R13471 gnd.n6202 gnd.n597 240.244
R13472 gnd.n6202 gnd.n599 240.244
R13473 gnd.n6198 gnd.n599 240.244
R13474 gnd.n6198 gnd.n605 240.244
R13475 gnd.n6194 gnd.n605 240.244
R13476 gnd.n6194 gnd.n607 240.244
R13477 gnd.n6190 gnd.n607 240.244
R13478 gnd.n6190 gnd.n613 240.244
R13479 gnd.n6186 gnd.n613 240.244
R13480 gnd.n6186 gnd.n615 240.244
R13481 gnd.n6182 gnd.n615 240.244
R13482 gnd.n6182 gnd.n621 240.244
R13483 gnd.n6178 gnd.n621 240.244
R13484 gnd.n6178 gnd.n623 240.244
R13485 gnd.n6174 gnd.n623 240.244
R13486 gnd.n6174 gnd.n629 240.244
R13487 gnd.n6170 gnd.n629 240.244
R13488 gnd.n6170 gnd.n631 240.244
R13489 gnd.n6166 gnd.n631 240.244
R13490 gnd.n6166 gnd.n637 240.244
R13491 gnd.n6162 gnd.n637 240.244
R13492 gnd.n6162 gnd.n639 240.244
R13493 gnd.n6158 gnd.n639 240.244
R13494 gnd.n6158 gnd.n645 240.244
R13495 gnd.n6154 gnd.n645 240.244
R13496 gnd.n6154 gnd.n647 240.244
R13497 gnd.n6150 gnd.n647 240.244
R13498 gnd.n6150 gnd.n653 240.244
R13499 gnd.n6146 gnd.n653 240.244
R13500 gnd.n6146 gnd.n655 240.244
R13501 gnd.n6142 gnd.n655 240.244
R13502 gnd.n6142 gnd.n661 240.244
R13503 gnd.n6138 gnd.n661 240.244
R13504 gnd.n6138 gnd.n663 240.244
R13505 gnd.n6134 gnd.n663 240.244
R13506 gnd.n6134 gnd.n669 240.244
R13507 gnd.n6130 gnd.n669 240.244
R13508 gnd.n6130 gnd.n671 240.244
R13509 gnd.n6126 gnd.n671 240.244
R13510 gnd.n6126 gnd.n677 240.244
R13511 gnd.n6122 gnd.n677 240.244
R13512 gnd.n6122 gnd.n679 240.244
R13513 gnd.n6118 gnd.n679 240.244
R13514 gnd.n6118 gnd.n685 240.244
R13515 gnd.n6114 gnd.n685 240.244
R13516 gnd.n6114 gnd.n687 240.244
R13517 gnd.n6110 gnd.n687 240.244
R13518 gnd.n6110 gnd.n693 240.244
R13519 gnd.n6106 gnd.n693 240.244
R13520 gnd.n6106 gnd.n695 240.244
R13521 gnd.n6102 gnd.n695 240.244
R13522 gnd.n6102 gnd.n701 240.244
R13523 gnd.n6098 gnd.n701 240.244
R13524 gnd.n6098 gnd.n703 240.244
R13525 gnd.n6094 gnd.n703 240.244
R13526 gnd.n6094 gnd.n709 240.244
R13527 gnd.n6090 gnd.n709 240.244
R13528 gnd.n6090 gnd.n711 240.244
R13529 gnd.n6086 gnd.n711 240.244
R13530 gnd.n6086 gnd.n717 240.244
R13531 gnd.n6082 gnd.n717 240.244
R13532 gnd.n6082 gnd.n719 240.244
R13533 gnd.n6078 gnd.n719 240.244
R13534 gnd.n6078 gnd.n725 240.244
R13535 gnd.n6074 gnd.n725 240.244
R13536 gnd.n6074 gnd.n727 240.244
R13537 gnd.n4311 gnd.n893 240.244
R13538 gnd.n4311 gnd.n2111 240.244
R13539 gnd.n4266 gnd.n2111 240.244
R13540 gnd.n4266 gnd.n2105 240.244
R13541 gnd.n4267 gnd.n2105 240.244
R13542 gnd.n4267 gnd.n2098 240.244
R13543 gnd.n4270 gnd.n2098 240.244
R13544 gnd.n4270 gnd.n2091 240.244
R13545 gnd.n4271 gnd.n2091 240.244
R13546 gnd.n4271 gnd.n2083 240.244
R13547 gnd.n4274 gnd.n2083 240.244
R13548 gnd.n4274 gnd.n2076 240.244
R13549 gnd.n4275 gnd.n2076 240.244
R13550 gnd.n4275 gnd.n2069 240.244
R13551 gnd.n4278 gnd.n2069 240.244
R13552 gnd.n4278 gnd.n2062 240.244
R13553 gnd.n4279 gnd.n2062 240.244
R13554 gnd.n4279 gnd.n2054 240.244
R13555 gnd.n2054 gnd.n2043 240.244
R13556 gnd.n4414 gnd.n2043 240.244
R13557 gnd.n4415 gnd.n4414 240.244
R13558 gnd.n4417 gnd.n4415 240.244
R13559 gnd.n4417 gnd.n4416 240.244
R13560 gnd.n4416 gnd.n1203 240.244
R13561 gnd.n4522 gnd.n1203 240.244
R13562 gnd.n4522 gnd.n1213 240.244
R13563 gnd.n2036 gnd.n1213 240.244
R13564 gnd.n4556 gnd.n2036 240.244
R13565 gnd.n4556 gnd.n2034 240.244
R13566 gnd.n2034 gnd.n2030 240.244
R13567 gnd.n2030 gnd.n2023 240.244
R13568 gnd.n4528 gnd.n2023 240.244
R13569 gnd.n4528 gnd.n2015 240.244
R13570 gnd.n4531 gnd.n2015 240.244
R13571 gnd.n4532 gnd.n4531 240.244
R13572 gnd.n4532 gnd.n1995 240.244
R13573 gnd.n4533 gnd.n1995 240.244
R13574 gnd.n4533 gnd.n1988 240.244
R13575 gnd.n4537 gnd.n1988 240.244
R13576 gnd.n4537 gnd.n1976 240.244
R13577 gnd.n4659 gnd.n1976 240.244
R13578 gnd.n4659 gnd.n1960 240.244
R13579 gnd.n1971 gnd.n1960 240.244
R13580 gnd.n4692 gnd.n1971 240.244
R13581 gnd.n4692 gnd.n1953 240.244
R13582 gnd.n1953 gnd.n1945 240.244
R13583 gnd.n4665 gnd.n1945 240.244
R13584 gnd.n4665 gnd.n1937 240.244
R13585 gnd.n4668 gnd.n1937 240.244
R13586 gnd.n4669 gnd.n4668 240.244
R13587 gnd.n4669 gnd.n1918 240.244
R13588 gnd.n4670 gnd.n1918 240.244
R13589 gnd.n4670 gnd.n1910 240.244
R13590 gnd.n4673 gnd.n1910 240.244
R13591 gnd.n4673 gnd.n1892 240.244
R13592 gnd.n1892 gnd.n1883 240.244
R13593 gnd.n4811 gnd.n1883 240.244
R13594 gnd.n4811 gnd.n1878 240.244
R13595 gnd.n4818 gnd.n1878 240.244
R13596 gnd.n4818 gnd.n1865 240.244
R13597 gnd.n1865 gnd.n1856 240.244
R13598 gnd.n4860 gnd.n1856 240.244
R13599 gnd.n4860 gnd.n1851 240.244
R13600 gnd.n4882 gnd.n1851 240.244
R13601 gnd.n4882 gnd.n1843 240.244
R13602 gnd.n4865 gnd.n1843 240.244
R13603 gnd.n4865 gnd.n1833 240.244
R13604 gnd.n4866 gnd.n1833 240.244
R13605 gnd.n4867 gnd.n4866 240.244
R13606 gnd.n4867 gnd.n1813 240.244
R13607 gnd.n1813 gnd.n1804 240.244
R13608 gnd.n4939 gnd.n1804 240.244
R13609 gnd.n4940 gnd.n4939 240.244
R13610 gnd.n4940 gnd.n1789 240.244
R13611 gnd.n4956 gnd.n1789 240.244
R13612 gnd.n4956 gnd.n1779 240.244
R13613 gnd.n4945 gnd.n1779 240.244
R13614 gnd.n4947 gnd.n4945 240.244
R13615 gnd.n4947 gnd.n1733 240.244
R13616 gnd.n1733 gnd.n1726 240.244
R13617 gnd.n5158 gnd.n1726 240.244
R13618 gnd.n5158 gnd.n1722 240.244
R13619 gnd.n5164 gnd.n1722 240.244
R13620 gnd.n5164 gnd.n1714 240.244
R13621 gnd.n5175 gnd.n1714 240.244
R13622 gnd.n5175 gnd.n1710 240.244
R13623 gnd.n5181 gnd.n1710 240.244
R13624 gnd.n5181 gnd.n1702 240.244
R13625 gnd.n5192 gnd.n1702 240.244
R13626 gnd.n5192 gnd.n1698 240.244
R13627 gnd.n5198 gnd.n1698 240.244
R13628 gnd.n5198 gnd.n1689 240.244
R13629 gnd.n5209 gnd.n1689 240.244
R13630 gnd.n5209 gnd.n1685 240.244
R13631 gnd.n5215 gnd.n1685 240.244
R13632 gnd.n5215 gnd.n1678 240.244
R13633 gnd.n5229 gnd.n1678 240.244
R13634 gnd.n5229 gnd.n1674 240.244
R13635 gnd.n5235 gnd.n1674 240.244
R13636 gnd.n5235 gnd.n1315 240.244
R13637 gnd.n5653 gnd.n1315 240.244
R13638 gnd.n892 gnd.n891 240.244
R13639 gnd.n897 gnd.n891 240.244
R13640 gnd.n899 gnd.n898 240.244
R13641 gnd.n903 gnd.n902 240.244
R13642 gnd.n905 gnd.n904 240.244
R13643 gnd.n915 gnd.n914 240.244
R13644 gnd.n917 gnd.n916 240.244
R13645 gnd.n925 gnd.n924 240.244
R13646 gnd.n933 gnd.n932 240.244
R13647 gnd.n935 gnd.n934 240.244
R13648 gnd.n943 gnd.n942 240.244
R13649 gnd.n951 gnd.n950 240.244
R13650 gnd.n956 gnd.n952 240.244
R13651 gnd.n888 gnd.n874 240.244
R13652 gnd.n4313 gnd.n875 240.244
R13653 gnd.n4320 gnd.n4313 240.244
R13654 gnd.n4320 gnd.n2103 240.244
R13655 gnd.n4330 gnd.n2103 240.244
R13656 gnd.n4330 gnd.n2099 240.244
R13657 gnd.n4336 gnd.n2099 240.244
R13658 gnd.n4336 gnd.n2089 240.244
R13659 gnd.n4346 gnd.n2089 240.244
R13660 gnd.n4346 gnd.n2085 240.244
R13661 gnd.n4352 gnd.n2085 240.244
R13662 gnd.n4352 gnd.n2075 240.244
R13663 gnd.n4362 gnd.n2075 240.244
R13664 gnd.n4362 gnd.n2071 240.244
R13665 gnd.n4368 gnd.n2071 240.244
R13666 gnd.n4368 gnd.n2061 240.244
R13667 gnd.n4378 gnd.n2061 240.244
R13668 gnd.n4378 gnd.n2055 240.244
R13669 gnd.n4398 gnd.n2055 240.244
R13670 gnd.n4398 gnd.n2056 240.244
R13671 gnd.n2056 gnd.n2046 240.244
R13672 gnd.n4383 gnd.n2046 240.244
R13673 gnd.n4384 gnd.n4383 240.244
R13674 gnd.n4385 gnd.n4384 240.244
R13675 gnd.n4385 gnd.n1204 240.244
R13676 gnd.n1214 gnd.n1204 240.244
R13677 gnd.n5770 gnd.n1214 240.244
R13678 gnd.n5770 gnd.n1215 240.244
R13679 gnd.n1220 gnd.n1215 240.244
R13680 gnd.n1221 gnd.n1220 240.244
R13681 gnd.n1222 gnd.n1221 240.244
R13682 gnd.n4585 gnd.n1222 240.244
R13683 gnd.n4585 gnd.n1225 240.244
R13684 gnd.n1226 gnd.n1225 240.244
R13685 gnd.n1227 gnd.n1226 240.244
R13686 gnd.n2002 gnd.n1227 240.244
R13687 gnd.n2002 gnd.n1230 240.244
R13688 gnd.n1231 gnd.n1230 240.244
R13689 gnd.n1232 gnd.n1231 240.244
R13690 gnd.n1982 gnd.n1232 240.244
R13691 gnd.n1982 gnd.n1235 240.244
R13692 gnd.n1236 gnd.n1235 240.244
R13693 gnd.n1237 gnd.n1236 240.244
R13694 gnd.n1969 gnd.n1237 240.244
R13695 gnd.n1969 gnd.n1240 240.244
R13696 gnd.n1241 gnd.n1240 240.244
R13697 gnd.n1242 gnd.n1241 240.244
R13698 gnd.n1934 gnd.n1242 240.244
R13699 gnd.n1934 gnd.n1245 240.244
R13700 gnd.n1246 gnd.n1245 240.244
R13701 gnd.n1247 gnd.n1246 240.244
R13702 gnd.n4762 gnd.n1247 240.244
R13703 gnd.n4762 gnd.n1250 240.244
R13704 gnd.n1251 gnd.n1250 240.244
R13705 gnd.n1252 gnd.n1251 240.244
R13706 gnd.n4799 gnd.n1252 240.244
R13707 gnd.n4799 gnd.n1255 240.244
R13708 gnd.n1256 gnd.n1255 240.244
R13709 gnd.n1257 gnd.n1256 240.244
R13710 gnd.n4819 gnd.n1257 240.244
R13711 gnd.n4819 gnd.n1260 240.244
R13712 gnd.n1261 gnd.n1260 240.244
R13713 gnd.n1262 gnd.n1261 240.244
R13714 gnd.n4839 gnd.n1262 240.244
R13715 gnd.n4839 gnd.n1265 240.244
R13716 gnd.n1266 gnd.n1265 240.244
R13717 gnd.n1267 gnd.n1266 240.244
R13718 gnd.n1835 gnd.n1267 240.244
R13719 gnd.n1835 gnd.n1270 240.244
R13720 gnd.n1271 gnd.n1270 240.244
R13721 gnd.n1272 gnd.n1271 240.244
R13722 gnd.n1815 gnd.n1272 240.244
R13723 gnd.n1815 gnd.n1275 240.244
R13724 gnd.n1276 gnd.n1275 240.244
R13725 gnd.n1277 gnd.n1276 240.244
R13726 gnd.n4957 gnd.n1277 240.244
R13727 gnd.n4957 gnd.n1280 240.244
R13728 gnd.n1281 gnd.n1280 240.244
R13729 gnd.n1282 gnd.n1281 240.244
R13730 gnd.n5148 gnd.n1282 240.244
R13731 gnd.n5148 gnd.n1285 240.244
R13732 gnd.n1286 gnd.n1285 240.244
R13733 gnd.n1287 gnd.n1286 240.244
R13734 gnd.n5165 gnd.n1287 240.244
R13735 gnd.n5165 gnd.n1290 240.244
R13736 gnd.n1291 gnd.n1290 240.244
R13737 gnd.n1292 gnd.n1291 240.244
R13738 gnd.n5182 gnd.n1292 240.244
R13739 gnd.n5182 gnd.n1295 240.244
R13740 gnd.n1296 gnd.n1295 240.244
R13741 gnd.n1297 gnd.n1296 240.244
R13742 gnd.n5199 gnd.n1297 240.244
R13743 gnd.n5199 gnd.n1300 240.244
R13744 gnd.n1301 gnd.n1300 240.244
R13745 gnd.n1302 gnd.n1301 240.244
R13746 gnd.n5216 gnd.n1302 240.244
R13747 gnd.n5216 gnd.n1305 240.244
R13748 gnd.n1306 gnd.n1305 240.244
R13749 gnd.n1307 gnd.n1306 240.244
R13750 gnd.n5236 gnd.n1307 240.244
R13751 gnd.n5236 gnd.n1310 240.244
R13752 gnd.n5655 gnd.n1310 240.244
R13753 gnd.n1321 gnd.n1320 240.244
R13754 gnd.n1645 gnd.n1324 240.244
R13755 gnd.n1326 gnd.n1325 240.244
R13756 gnd.n1648 gnd.n1330 240.244
R13757 gnd.n1651 gnd.n1331 240.244
R13758 gnd.n1340 gnd.n1339 240.244
R13759 gnd.n1653 gnd.n1347 240.244
R13760 gnd.n1656 gnd.n1348 240.244
R13761 gnd.n1356 gnd.n1355 240.244
R13762 gnd.n1658 gnd.n1363 240.244
R13763 gnd.n1661 gnd.n1364 240.244
R13764 gnd.n1372 gnd.n1371 240.244
R13765 gnd.n1664 gnd.n1372 240.244
R13766 gnd.n5261 gnd.n1643 240.244
R13767 gnd.n1185 gnd.n1184 240.132
R13768 gnd.n4998 gnd.n4997 240.132
R13769 gnd.n6246 gnd.n6245 225.874
R13770 gnd.n6247 gnd.n6246 225.874
R13771 gnd.n6247 gnd.n555 225.874
R13772 gnd.n6255 gnd.n555 225.874
R13773 gnd.n6256 gnd.n6255 225.874
R13774 gnd.n6257 gnd.n6256 225.874
R13775 gnd.n6257 gnd.n549 225.874
R13776 gnd.n6265 gnd.n549 225.874
R13777 gnd.n6266 gnd.n6265 225.874
R13778 gnd.n6267 gnd.n6266 225.874
R13779 gnd.n6267 gnd.n543 225.874
R13780 gnd.n6275 gnd.n543 225.874
R13781 gnd.n6276 gnd.n6275 225.874
R13782 gnd.n6277 gnd.n6276 225.874
R13783 gnd.n6277 gnd.n537 225.874
R13784 gnd.n6285 gnd.n537 225.874
R13785 gnd.n6286 gnd.n6285 225.874
R13786 gnd.n6287 gnd.n6286 225.874
R13787 gnd.n6287 gnd.n531 225.874
R13788 gnd.n6295 gnd.n531 225.874
R13789 gnd.n6296 gnd.n6295 225.874
R13790 gnd.n6297 gnd.n6296 225.874
R13791 gnd.n6297 gnd.n525 225.874
R13792 gnd.n6305 gnd.n525 225.874
R13793 gnd.n6306 gnd.n6305 225.874
R13794 gnd.n6307 gnd.n6306 225.874
R13795 gnd.n6307 gnd.n519 225.874
R13796 gnd.n6315 gnd.n519 225.874
R13797 gnd.n6316 gnd.n6315 225.874
R13798 gnd.n6317 gnd.n6316 225.874
R13799 gnd.n6317 gnd.n513 225.874
R13800 gnd.n6325 gnd.n513 225.874
R13801 gnd.n6326 gnd.n6325 225.874
R13802 gnd.n6327 gnd.n6326 225.874
R13803 gnd.n6327 gnd.n507 225.874
R13804 gnd.n6335 gnd.n507 225.874
R13805 gnd.n6336 gnd.n6335 225.874
R13806 gnd.n6337 gnd.n6336 225.874
R13807 gnd.n6337 gnd.n501 225.874
R13808 gnd.n6345 gnd.n501 225.874
R13809 gnd.n6346 gnd.n6345 225.874
R13810 gnd.n6347 gnd.n6346 225.874
R13811 gnd.n6347 gnd.n495 225.874
R13812 gnd.n6355 gnd.n495 225.874
R13813 gnd.n6356 gnd.n6355 225.874
R13814 gnd.n6357 gnd.n6356 225.874
R13815 gnd.n6357 gnd.n489 225.874
R13816 gnd.n6365 gnd.n489 225.874
R13817 gnd.n6366 gnd.n6365 225.874
R13818 gnd.n6367 gnd.n6366 225.874
R13819 gnd.n6367 gnd.n483 225.874
R13820 gnd.n6375 gnd.n483 225.874
R13821 gnd.n6376 gnd.n6375 225.874
R13822 gnd.n6377 gnd.n6376 225.874
R13823 gnd.n6377 gnd.n477 225.874
R13824 gnd.n6385 gnd.n477 225.874
R13825 gnd.n6386 gnd.n6385 225.874
R13826 gnd.n6387 gnd.n6386 225.874
R13827 gnd.n6387 gnd.n471 225.874
R13828 gnd.n6395 gnd.n471 225.874
R13829 gnd.n6396 gnd.n6395 225.874
R13830 gnd.n6397 gnd.n6396 225.874
R13831 gnd.n6397 gnd.n465 225.874
R13832 gnd.n6405 gnd.n465 225.874
R13833 gnd.n6406 gnd.n6405 225.874
R13834 gnd.n6407 gnd.n6406 225.874
R13835 gnd.n6407 gnd.n459 225.874
R13836 gnd.n6415 gnd.n459 225.874
R13837 gnd.n6416 gnd.n6415 225.874
R13838 gnd.n6417 gnd.n6416 225.874
R13839 gnd.n6417 gnd.n453 225.874
R13840 gnd.n6425 gnd.n453 225.874
R13841 gnd.n6426 gnd.n6425 225.874
R13842 gnd.n6427 gnd.n6426 225.874
R13843 gnd.n6427 gnd.n447 225.874
R13844 gnd.n6435 gnd.n447 225.874
R13845 gnd.n6436 gnd.n6435 225.874
R13846 gnd.n6437 gnd.n6436 225.874
R13847 gnd.n6437 gnd.n441 225.874
R13848 gnd.n6445 gnd.n441 225.874
R13849 gnd.n6446 gnd.n6445 225.874
R13850 gnd.n6447 gnd.n6446 225.874
R13851 gnd.n6447 gnd.n435 225.874
R13852 gnd.n6455 gnd.n435 225.874
R13853 gnd.n6456 gnd.n6455 225.874
R13854 gnd.n6457 gnd.n6456 225.874
R13855 gnd.n6457 gnd.n429 225.874
R13856 gnd.n6465 gnd.n429 225.874
R13857 gnd.n6466 gnd.n6465 225.874
R13858 gnd.n6467 gnd.n6466 225.874
R13859 gnd.n6467 gnd.n423 225.874
R13860 gnd.n6475 gnd.n423 225.874
R13861 gnd.n6476 gnd.n6475 225.874
R13862 gnd.n6477 gnd.n6476 225.874
R13863 gnd.n6477 gnd.n417 225.874
R13864 gnd.n6485 gnd.n417 225.874
R13865 gnd.n6486 gnd.n6485 225.874
R13866 gnd.n6487 gnd.n6486 225.874
R13867 gnd.n6487 gnd.n411 225.874
R13868 gnd.n6495 gnd.n411 225.874
R13869 gnd.n6496 gnd.n6495 225.874
R13870 gnd.n6497 gnd.n6496 225.874
R13871 gnd.n6497 gnd.n405 225.874
R13872 gnd.n6505 gnd.n405 225.874
R13873 gnd.n6506 gnd.n6505 225.874
R13874 gnd.n6507 gnd.n6506 225.874
R13875 gnd.n6507 gnd.n399 225.874
R13876 gnd.n6515 gnd.n399 225.874
R13877 gnd.n6516 gnd.n6515 225.874
R13878 gnd.n6517 gnd.n6516 225.874
R13879 gnd.n6517 gnd.n393 225.874
R13880 gnd.n6525 gnd.n393 225.874
R13881 gnd.n6526 gnd.n6525 225.874
R13882 gnd.n6527 gnd.n6526 225.874
R13883 gnd.n6527 gnd.n387 225.874
R13884 gnd.n6535 gnd.n387 225.874
R13885 gnd.n6536 gnd.n6535 225.874
R13886 gnd.n6537 gnd.n6536 225.874
R13887 gnd.n6537 gnd.n381 225.874
R13888 gnd.n6545 gnd.n381 225.874
R13889 gnd.n6546 gnd.n6545 225.874
R13890 gnd.n6547 gnd.n6546 225.874
R13891 gnd.n6547 gnd.n375 225.874
R13892 gnd.n6555 gnd.n375 225.874
R13893 gnd.n6556 gnd.n6555 225.874
R13894 gnd.n6557 gnd.n6556 225.874
R13895 gnd.n6557 gnd.n369 225.874
R13896 gnd.n6565 gnd.n369 225.874
R13897 gnd.n6566 gnd.n6565 225.874
R13898 gnd.n6567 gnd.n6566 225.874
R13899 gnd.n6567 gnd.n363 225.874
R13900 gnd.n6575 gnd.n363 225.874
R13901 gnd.n6576 gnd.n6575 225.874
R13902 gnd.n6577 gnd.n6576 225.874
R13903 gnd.n6577 gnd.n357 225.874
R13904 gnd.n6585 gnd.n357 225.874
R13905 gnd.n6586 gnd.n6585 225.874
R13906 gnd.n6587 gnd.n6586 225.874
R13907 gnd.n6587 gnd.n351 225.874
R13908 gnd.n6595 gnd.n351 225.874
R13909 gnd.n6596 gnd.n6595 225.874
R13910 gnd.n6597 gnd.n6596 225.874
R13911 gnd.n6597 gnd.n345 225.874
R13912 gnd.n6605 gnd.n345 225.874
R13913 gnd.n6606 gnd.n6605 225.874
R13914 gnd.n6607 gnd.n6606 225.874
R13915 gnd.n6607 gnd.n339 225.874
R13916 gnd.n6615 gnd.n339 225.874
R13917 gnd.n6616 gnd.n6615 225.874
R13918 gnd.n6617 gnd.n6616 225.874
R13919 gnd.n6617 gnd.n333 225.874
R13920 gnd.n6625 gnd.n333 225.874
R13921 gnd.n6626 gnd.n6625 225.874
R13922 gnd.n6627 gnd.n6626 225.874
R13923 gnd.n6627 gnd.n327 225.874
R13924 gnd.n6635 gnd.n327 225.874
R13925 gnd.n6636 gnd.n6635 225.874
R13926 gnd.n6637 gnd.n6636 225.874
R13927 gnd.n6637 gnd.n321 225.874
R13928 gnd.n6645 gnd.n321 225.874
R13929 gnd.n6646 gnd.n6645 225.874
R13930 gnd.n6647 gnd.n6646 225.874
R13931 gnd.n6647 gnd.n315 225.874
R13932 gnd.n6656 gnd.n315 225.874
R13933 gnd.n6657 gnd.n6656 225.874
R13934 gnd.n6658 gnd.n6657 225.874
R13935 gnd.n6658 gnd.n310 225.874
R13936 gnd.n2796 gnd.t131 224.174
R13937 gnd.n2306 gnd.t36 224.174
R13938 gnd.n1456 gnd.n1393 199.319
R13939 gnd.n1456 gnd.n1394 199.319
R13940 gnd.n1041 gnd.n996 199.319
R13941 gnd.n1041 gnd.n995 199.319
R13942 gnd.n1186 gnd.n1183 186.49
R13943 gnd.n4999 gnd.n4996 186.49
R13944 gnd.n3571 gnd.n3570 185
R13945 gnd.n3569 gnd.n3568 185
R13946 gnd.n3548 gnd.n3547 185
R13947 gnd.n3563 gnd.n3562 185
R13948 gnd.n3561 gnd.n3560 185
R13949 gnd.n3552 gnd.n3551 185
R13950 gnd.n3555 gnd.n3554 185
R13951 gnd.n3539 gnd.n3538 185
R13952 gnd.n3537 gnd.n3536 185
R13953 gnd.n3516 gnd.n3515 185
R13954 gnd.n3531 gnd.n3530 185
R13955 gnd.n3529 gnd.n3528 185
R13956 gnd.n3520 gnd.n3519 185
R13957 gnd.n3523 gnd.n3522 185
R13958 gnd.n3507 gnd.n3506 185
R13959 gnd.n3505 gnd.n3504 185
R13960 gnd.n3484 gnd.n3483 185
R13961 gnd.n3499 gnd.n3498 185
R13962 gnd.n3497 gnd.n3496 185
R13963 gnd.n3488 gnd.n3487 185
R13964 gnd.n3491 gnd.n3490 185
R13965 gnd.n3476 gnd.n3475 185
R13966 gnd.n3474 gnd.n3473 185
R13967 gnd.n3453 gnd.n3452 185
R13968 gnd.n3468 gnd.n3467 185
R13969 gnd.n3466 gnd.n3465 185
R13970 gnd.n3457 gnd.n3456 185
R13971 gnd.n3460 gnd.n3459 185
R13972 gnd.n3444 gnd.n3443 185
R13973 gnd.n3442 gnd.n3441 185
R13974 gnd.n3421 gnd.n3420 185
R13975 gnd.n3436 gnd.n3435 185
R13976 gnd.n3434 gnd.n3433 185
R13977 gnd.n3425 gnd.n3424 185
R13978 gnd.n3428 gnd.n3427 185
R13979 gnd.n3412 gnd.n3411 185
R13980 gnd.n3410 gnd.n3409 185
R13981 gnd.n3389 gnd.n3388 185
R13982 gnd.n3404 gnd.n3403 185
R13983 gnd.n3402 gnd.n3401 185
R13984 gnd.n3393 gnd.n3392 185
R13985 gnd.n3396 gnd.n3395 185
R13986 gnd.n3380 gnd.n3379 185
R13987 gnd.n3378 gnd.n3377 185
R13988 gnd.n3357 gnd.n3356 185
R13989 gnd.n3372 gnd.n3371 185
R13990 gnd.n3370 gnd.n3369 185
R13991 gnd.n3361 gnd.n3360 185
R13992 gnd.n3364 gnd.n3363 185
R13993 gnd.n3349 gnd.n3348 185
R13994 gnd.n3347 gnd.n3346 185
R13995 gnd.n3326 gnd.n3325 185
R13996 gnd.n3341 gnd.n3340 185
R13997 gnd.n3339 gnd.n3338 185
R13998 gnd.n3330 gnd.n3329 185
R13999 gnd.n3333 gnd.n3332 185
R14000 gnd.n2797 gnd.t130 178.987
R14001 gnd.n2307 gnd.t37 178.987
R14002 gnd.n1 gnd.t318 170.774
R14003 gnd.n9 gnd.t295 170.103
R14004 gnd.n8 gnd.t301 170.103
R14005 gnd.n7 gnd.t298 170.103
R14006 gnd.n6 gnd.t271 170.103
R14007 gnd.n5 gnd.t3 170.103
R14008 gnd.n4 gnd.t21 170.103
R14009 gnd.n3 gnd.t15 170.103
R14010 gnd.n2 gnd.t312 170.103
R14011 gnd.n1 gnd.t8 170.103
R14012 gnd.n5533 gnd.n1455 167.873
R14013 gnd.n5852 gnd.n5851 167.873
R14014 gnd.n5070 gnd.n5069 163.367
R14015 gnd.n5066 gnd.n5065 163.367
R14016 gnd.n5062 gnd.n5061 163.367
R14017 gnd.n5058 gnd.n5057 163.367
R14018 gnd.n5054 gnd.n5053 163.367
R14019 gnd.n5050 gnd.n5049 163.367
R14020 gnd.n5046 gnd.n5045 163.367
R14021 gnd.n5042 gnd.n5041 163.367
R14022 gnd.n5038 gnd.n5037 163.367
R14023 gnd.n5034 gnd.n5033 163.367
R14024 gnd.n5030 gnd.n5029 163.367
R14025 gnd.n5026 gnd.n5025 163.367
R14026 gnd.n5022 gnd.n5021 163.367
R14027 gnd.n5018 gnd.n5017 163.367
R14028 gnd.n5013 gnd.n5012 163.367
R14029 gnd.n5009 gnd.n5008 163.367
R14030 gnd.n5146 gnd.n5145 163.367
R14031 gnd.n5142 gnd.n5141 163.367
R14032 gnd.n5137 gnd.n5136 163.367
R14033 gnd.n5133 gnd.n5132 163.367
R14034 gnd.n5129 gnd.n5128 163.367
R14035 gnd.n5125 gnd.n5124 163.367
R14036 gnd.n5121 gnd.n5120 163.367
R14037 gnd.n5117 gnd.n5116 163.367
R14038 gnd.n5113 gnd.n5112 163.367
R14039 gnd.n5109 gnd.n5108 163.367
R14040 gnd.n5105 gnd.n5104 163.367
R14041 gnd.n5101 gnd.n5100 163.367
R14042 gnd.n5097 gnd.n5096 163.367
R14043 gnd.n5093 gnd.n5092 163.367
R14044 gnd.n5089 gnd.n5088 163.367
R14045 gnd.n5085 gnd.n5084 163.367
R14046 gnd.n4493 gnd.n1202 163.367
R14047 gnd.n4425 gnd.n1202 163.367
R14048 gnd.n4520 gnd.n4425 163.367
R14049 gnd.n4520 gnd.n4426 163.367
R14050 gnd.n4516 gnd.n4426 163.367
R14051 gnd.n4516 gnd.n4500 163.367
R14052 gnd.n4500 gnd.n4499 163.367
R14053 gnd.n4499 gnd.n2032 163.367
R14054 gnd.n4567 gnd.n2032 163.367
R14055 gnd.n4567 gnd.n2029 163.367
R14056 gnd.n4575 gnd.n2029 163.367
R14057 gnd.n4575 gnd.n2024 163.367
R14058 gnd.n4571 gnd.n2024 163.367
R14059 gnd.n4571 gnd.n2014 163.367
R14060 gnd.n2014 gnd.n2007 163.367
R14061 gnd.n4604 gnd.n2007 163.367
R14062 gnd.n4604 gnd.n2004 163.367
R14063 gnd.n4613 gnd.n2004 163.367
R14064 gnd.n4613 gnd.n2005 163.367
R14065 gnd.n2005 gnd.n1996 163.367
R14066 gnd.n4608 gnd.n1996 163.367
R14067 gnd.n4608 gnd.n1986 163.367
R14068 gnd.n4640 gnd.n1986 163.367
R14069 gnd.n4640 gnd.n1984 163.367
R14070 gnd.n4649 gnd.n1984 163.367
R14071 gnd.n4649 gnd.n1978 163.367
R14072 gnd.n4645 gnd.n1978 163.367
R14073 gnd.n4645 gnd.n1962 163.367
R14074 gnd.n1962 gnd.n1955 163.367
R14075 gnd.n4706 gnd.n1955 163.367
R14076 gnd.n4707 gnd.n4706 163.367
R14077 gnd.n4707 gnd.n1952 163.367
R14078 gnd.n4715 gnd.n1952 163.367
R14079 gnd.n4715 gnd.n1946 163.367
R14080 gnd.n4711 gnd.n1946 163.367
R14081 gnd.n4711 gnd.n1936 163.367
R14082 gnd.n1936 gnd.n1928 163.367
R14083 gnd.n4743 gnd.n1928 163.367
R14084 gnd.n4743 gnd.n1925 163.367
R14085 gnd.n4754 gnd.n1925 163.367
R14086 gnd.n4754 gnd.n1926 163.367
R14087 gnd.n1926 gnd.n1919 163.367
R14088 gnd.n4749 gnd.n1919 163.367
R14089 gnd.n4749 gnd.n1909 163.367
R14090 gnd.n1909 gnd.n1904 163.367
R14091 gnd.n4779 gnd.n1904 163.367
R14092 gnd.n4780 gnd.n4779 163.367
R14093 gnd.n4780 gnd.n1893 163.367
R14094 gnd.n4784 gnd.n1893 163.367
R14095 gnd.n4784 gnd.n1902 163.367
R14096 gnd.n4789 gnd.n1902 163.367
R14097 gnd.n4789 gnd.n1875 163.367
R14098 gnd.n4821 gnd.n1875 163.367
R14099 gnd.n4822 gnd.n4821 163.367
R14100 gnd.n4822 gnd.n1866 163.367
R14101 gnd.n4826 gnd.n1866 163.367
R14102 gnd.n4826 gnd.n1872 163.367
R14103 gnd.n4838 gnd.n1872 163.367
R14104 gnd.n4838 gnd.n1873 163.367
R14105 gnd.n1873 gnd.n1850 163.367
R14106 gnd.n4833 gnd.n1850 163.367
R14107 gnd.n4833 gnd.n1844 163.367
R14108 gnd.n4830 gnd.n1844 163.367
R14109 gnd.n4830 gnd.n1832 163.367
R14110 gnd.n1832 gnd.n1825 163.367
R14111 gnd.n4908 gnd.n1825 163.367
R14112 gnd.n4908 gnd.n1822 163.367
R14113 gnd.n4919 gnd.n1822 163.367
R14114 gnd.n4919 gnd.n1823 163.367
R14115 gnd.n1823 gnd.n1814 163.367
R14116 gnd.n4914 gnd.n1814 163.367
R14117 gnd.n4914 gnd.n4912 163.367
R14118 gnd.n4912 gnd.n1795 163.367
R14119 gnd.n4965 gnd.n1795 163.367
R14120 gnd.n4965 gnd.n1796 163.367
R14121 gnd.n1796 gnd.n1790 163.367
R14122 gnd.n4960 gnd.n1790 163.367
R14123 gnd.n4960 gnd.n1781 163.367
R14124 gnd.n1781 gnd.n1772 163.367
R14125 gnd.n5079 gnd.n1772 163.367
R14126 gnd.n5080 gnd.n5079 163.367
R14127 gnd.n1177 gnd.n1176 163.367
R14128 gnd.n5841 gnd.n1176 163.367
R14129 gnd.n5839 gnd.n5838 163.367
R14130 gnd.n5835 gnd.n5834 163.367
R14131 gnd.n5831 gnd.n5830 163.367
R14132 gnd.n5827 gnd.n5826 163.367
R14133 gnd.n5823 gnd.n5822 163.367
R14134 gnd.n5819 gnd.n5818 163.367
R14135 gnd.n5815 gnd.n5814 163.367
R14136 gnd.n5811 gnd.n5810 163.367
R14137 gnd.n5807 gnd.n5806 163.367
R14138 gnd.n5803 gnd.n5802 163.367
R14139 gnd.n5799 gnd.n5798 163.367
R14140 gnd.n5795 gnd.n5794 163.367
R14141 gnd.n5791 gnd.n5790 163.367
R14142 gnd.n5787 gnd.n5786 163.367
R14143 gnd.n5850 gnd.n1142 163.367
R14144 gnd.n4431 gnd.n4430 163.367
R14145 gnd.n4436 gnd.n4435 163.367
R14146 gnd.n4440 gnd.n4439 163.367
R14147 gnd.n4444 gnd.n4443 163.367
R14148 gnd.n4448 gnd.n4447 163.367
R14149 gnd.n4452 gnd.n4451 163.367
R14150 gnd.n4456 gnd.n4455 163.367
R14151 gnd.n4460 gnd.n4459 163.367
R14152 gnd.n4464 gnd.n4463 163.367
R14153 gnd.n4468 gnd.n4467 163.367
R14154 gnd.n4472 gnd.n4471 163.367
R14155 gnd.n4476 gnd.n4475 163.367
R14156 gnd.n4480 gnd.n4479 163.367
R14157 gnd.n4484 gnd.n4483 163.367
R14158 gnd.n4488 gnd.n4487 163.367
R14159 gnd.n5779 gnd.n1178 163.367
R14160 gnd.n5779 gnd.n1200 163.367
R14161 gnd.n4424 gnd.n1200 163.367
R14162 gnd.n4503 gnd.n4424 163.367
R14163 gnd.n4514 gnd.n4503 163.367
R14164 gnd.n4514 gnd.n4505 163.367
R14165 gnd.n4510 gnd.n4505 163.367
R14166 gnd.n4510 gnd.n4509 163.367
R14167 gnd.n4509 gnd.n2028 163.367
R14168 gnd.n4579 gnd.n2028 163.367
R14169 gnd.n4579 gnd.n2026 163.367
R14170 gnd.n4583 gnd.n2026 163.367
R14171 gnd.n4583 gnd.n2012 163.367
R14172 gnd.n4598 gnd.n2012 163.367
R14173 gnd.n4598 gnd.n2010 163.367
R14174 gnd.n4602 gnd.n2010 163.367
R14175 gnd.n4602 gnd.n2001 163.367
R14176 gnd.n4615 gnd.n2001 163.367
R14177 gnd.n4615 gnd.n1998 163.367
R14178 gnd.n4622 gnd.n1998 163.367
R14179 gnd.n4622 gnd.n1999 163.367
R14180 gnd.n4618 gnd.n1999 163.367
R14181 gnd.n4618 gnd.n1981 163.367
R14182 gnd.n4652 gnd.n1981 163.367
R14183 gnd.n4652 gnd.n1979 163.367
R14184 gnd.n4656 gnd.n1979 163.367
R14185 gnd.n4656 gnd.n1958 163.367
R14186 gnd.n4700 gnd.n1958 163.367
R14187 gnd.n4700 gnd.n1956 163.367
R14188 gnd.n4704 gnd.n1956 163.367
R14189 gnd.n4704 gnd.n1950 163.367
R14190 gnd.n4719 gnd.n1950 163.367
R14191 gnd.n4719 gnd.n1948 163.367
R14192 gnd.n4723 gnd.n1948 163.367
R14193 gnd.n4723 gnd.n1933 163.367
R14194 gnd.n4737 gnd.n1933 163.367
R14195 gnd.n4737 gnd.n1931 163.367
R14196 gnd.n4741 gnd.n1931 163.367
R14197 gnd.n4741 gnd.n1923 163.367
R14198 gnd.n4756 gnd.n1923 163.367
R14199 gnd.n4756 gnd.n1921 163.367
R14200 gnd.n4760 gnd.n1921 163.367
R14201 gnd.n4760 gnd.n1908 163.367
R14202 gnd.n4773 gnd.n1908 163.367
R14203 gnd.n4773 gnd.n1906 163.367
R14204 gnd.n4777 gnd.n1906 163.367
R14205 gnd.n4777 gnd.n1895 163.367
R14206 gnd.n4797 gnd.n1895 163.367
R14207 gnd.n4797 gnd.n1896 163.367
R14208 gnd.n4793 gnd.n1896 163.367
R14209 gnd.n4793 gnd.n4792 163.367
R14210 gnd.n4792 gnd.n1901 163.367
R14211 gnd.n1901 gnd.n1877 163.367
R14212 gnd.n1877 gnd.n1868 163.367
R14213 gnd.n4847 gnd.n1868 163.367
R14214 gnd.n4847 gnd.n1869 163.367
R14215 gnd.n4843 gnd.n1869 163.367
R14216 gnd.n4843 gnd.n4842 163.367
R14217 gnd.n4842 gnd.n1848 163.367
R14218 gnd.n4885 gnd.n1848 163.367
R14219 gnd.n4885 gnd.n1846 163.367
R14220 gnd.n4889 gnd.n1846 163.367
R14221 gnd.n4889 gnd.n1830 163.367
R14222 gnd.n4902 gnd.n1830 163.367
R14223 gnd.n4902 gnd.n1828 163.367
R14224 gnd.n4906 gnd.n1828 163.367
R14225 gnd.n4906 gnd.n1820 163.367
R14226 gnd.n4921 gnd.n1820 163.367
R14227 gnd.n4921 gnd.n1817 163.367
R14228 gnd.n4928 gnd.n1817 163.367
R14229 gnd.n4928 gnd.n1818 163.367
R14230 gnd.n4924 gnd.n1818 163.367
R14231 gnd.n4924 gnd.n1793 163.367
R14232 gnd.n4967 gnd.n1793 163.367
R14233 gnd.n4967 gnd.n1791 163.367
R14234 gnd.n4971 gnd.n1791 163.367
R14235 gnd.n4971 gnd.n1778 163.367
R14236 gnd.n4984 gnd.n1778 163.367
R14237 gnd.n4984 gnd.n1775 163.367
R14238 gnd.n5077 gnd.n1775 163.367
R14239 gnd.n5077 gnd.n1776 163.367
R14240 gnd.n5005 gnd.n5004 156.462
R14241 gnd.n3511 gnd.n3479 153.042
R14242 gnd.n3575 gnd.n3574 152.079
R14243 gnd.n3543 gnd.n3542 152.079
R14244 gnd.n3511 gnd.n3510 152.079
R14245 gnd.n1191 gnd.n1190 152
R14246 gnd.n1192 gnd.n1181 152
R14247 gnd.n1194 gnd.n1193 152
R14248 gnd.n1196 gnd.n1179 152
R14249 gnd.n1198 gnd.n1197 152
R14250 gnd.n5003 gnd.n4987 152
R14251 gnd.n4995 gnd.n4988 152
R14252 gnd.n4994 gnd.n4993 152
R14253 gnd.n4992 gnd.n4989 152
R14254 gnd.n4990 gnd.t77 150.546
R14255 gnd.t293 gnd.n3553 147.661
R14256 gnd.t269 gnd.n3521 147.661
R14257 gnd.t10 gnd.n3489 147.661
R14258 gnd.t143 gnd.n3458 147.661
R14259 gnd.t6 gnd.n3426 147.661
R14260 gnd.t12 gnd.n3394 147.661
R14261 gnd.t327 gnd.n3362 147.661
R14262 gnd.t291 gnd.n3331 147.661
R14263 gnd.n6667 gnd.n6666 143.933
R14264 gnd.n6668 gnd.n6667 143.933
R14265 gnd.n6668 gnd.n304 143.933
R14266 gnd.n6676 gnd.n304 143.933
R14267 gnd.n6677 gnd.n6676 143.933
R14268 gnd.n6678 gnd.n6677 143.933
R14269 gnd.n6678 gnd.n298 143.933
R14270 gnd.n6686 gnd.n298 143.933
R14271 gnd.n6687 gnd.n6686 143.933
R14272 gnd.n6688 gnd.n6687 143.933
R14273 gnd.n6688 gnd.n292 143.933
R14274 gnd.n6696 gnd.n292 143.933
R14275 gnd.n6697 gnd.n6696 143.933
R14276 gnd.n6698 gnd.n6697 143.933
R14277 gnd.n6698 gnd.n286 143.933
R14278 gnd.n6706 gnd.n286 143.933
R14279 gnd.n6707 gnd.n6706 143.933
R14280 gnd.n6708 gnd.n6707 143.933
R14281 gnd.n6708 gnd.n280 143.933
R14282 gnd.n6716 gnd.n280 143.933
R14283 gnd.n6717 gnd.n6716 143.933
R14284 gnd.n6718 gnd.n6717 143.933
R14285 gnd.n6718 gnd.n274 143.933
R14286 gnd.n6726 gnd.n274 143.933
R14287 gnd.n6727 gnd.n6726 143.933
R14288 gnd.n6728 gnd.n6727 143.933
R14289 gnd.n6728 gnd.n268 143.933
R14290 gnd.n6736 gnd.n268 143.933
R14291 gnd.n6737 gnd.n6736 143.933
R14292 gnd.n6738 gnd.n6737 143.933
R14293 gnd.n6738 gnd.n262 143.933
R14294 gnd.n6746 gnd.n262 143.933
R14295 gnd.n6747 gnd.n6746 143.933
R14296 gnd.n6748 gnd.n6747 143.933
R14297 gnd.n6748 gnd.n256 143.933
R14298 gnd.n6756 gnd.n256 143.933
R14299 gnd.n6757 gnd.n6756 143.933
R14300 gnd.n6758 gnd.n6757 143.933
R14301 gnd.n6758 gnd.n250 143.933
R14302 gnd.n6766 gnd.n250 143.933
R14303 gnd.n6767 gnd.n6766 143.933
R14304 gnd.n6768 gnd.n6767 143.933
R14305 gnd.n6768 gnd.n244 143.933
R14306 gnd.n6776 gnd.n244 143.933
R14307 gnd.n6777 gnd.n6776 143.933
R14308 gnd.n6778 gnd.n6777 143.933
R14309 gnd.n6778 gnd.n238 143.933
R14310 gnd.n6786 gnd.n238 143.933
R14311 gnd.n6787 gnd.n6786 143.933
R14312 gnd.n6788 gnd.n6787 143.933
R14313 gnd.n6788 gnd.n232 143.933
R14314 gnd.n6796 gnd.n232 143.933
R14315 gnd.n6797 gnd.n6796 143.933
R14316 gnd.n6798 gnd.n6797 143.933
R14317 gnd.n6798 gnd.n226 143.933
R14318 gnd.n6806 gnd.n226 143.933
R14319 gnd.n6807 gnd.n6806 143.933
R14320 gnd.n6808 gnd.n6807 143.933
R14321 gnd.n6808 gnd.n220 143.933
R14322 gnd.n6816 gnd.n220 143.933
R14323 gnd.n6817 gnd.n6816 143.933
R14324 gnd.n6818 gnd.n6817 143.933
R14325 gnd.n6818 gnd.n214 143.933
R14326 gnd.n6826 gnd.n214 143.933
R14327 gnd.n6827 gnd.n6826 143.933
R14328 gnd.n6828 gnd.n6827 143.933
R14329 gnd.n6828 gnd.n208 143.933
R14330 gnd.n6836 gnd.n208 143.933
R14331 gnd.n6837 gnd.n6836 143.933
R14332 gnd.n6838 gnd.n6837 143.933
R14333 gnd.n6838 gnd.n202 143.933
R14334 gnd.n6846 gnd.n202 143.933
R14335 gnd.n6847 gnd.n6846 143.933
R14336 gnd.n6848 gnd.n6847 143.933
R14337 gnd.n6848 gnd.n196 143.933
R14338 gnd.n6856 gnd.n196 143.933
R14339 gnd.n6857 gnd.n6856 143.933
R14340 gnd.n6858 gnd.n6857 143.933
R14341 gnd.n6858 gnd.n190 143.933
R14342 gnd.n6866 gnd.n190 143.933
R14343 gnd.n6867 gnd.n6866 143.933
R14344 gnd.n6869 gnd.n6867 143.933
R14345 gnd.n6869 gnd.n6868 143.933
R14346 gnd.n1768 gnd.n1750 143.351
R14347 gnd.n1158 gnd.n1141 143.351
R14348 gnd.n5849 gnd.n1141 143.351
R14349 gnd.n1188 gnd.t125 130.484
R14350 gnd.n1197 gnd.t38 126.766
R14351 gnd.n1195 gnd.t92 126.766
R14352 gnd.n1181 gnd.t48 126.766
R14353 gnd.n1189 gnd.t74 126.766
R14354 gnd.n4991 gnd.t139 126.766
R14355 gnd.n4993 gnd.t89 126.766
R14356 gnd.n5002 gnd.t41 126.766
R14357 gnd.n5004 gnd.t110 126.766
R14358 gnd.n3570 gnd.n3569 104.615
R14359 gnd.n3569 gnd.n3547 104.615
R14360 gnd.n3562 gnd.n3547 104.615
R14361 gnd.n3562 gnd.n3561 104.615
R14362 gnd.n3561 gnd.n3551 104.615
R14363 gnd.n3554 gnd.n3551 104.615
R14364 gnd.n3538 gnd.n3537 104.615
R14365 gnd.n3537 gnd.n3515 104.615
R14366 gnd.n3530 gnd.n3515 104.615
R14367 gnd.n3530 gnd.n3529 104.615
R14368 gnd.n3529 gnd.n3519 104.615
R14369 gnd.n3522 gnd.n3519 104.615
R14370 gnd.n3506 gnd.n3505 104.615
R14371 gnd.n3505 gnd.n3483 104.615
R14372 gnd.n3498 gnd.n3483 104.615
R14373 gnd.n3498 gnd.n3497 104.615
R14374 gnd.n3497 gnd.n3487 104.615
R14375 gnd.n3490 gnd.n3487 104.615
R14376 gnd.n3475 gnd.n3474 104.615
R14377 gnd.n3474 gnd.n3452 104.615
R14378 gnd.n3467 gnd.n3452 104.615
R14379 gnd.n3467 gnd.n3466 104.615
R14380 gnd.n3466 gnd.n3456 104.615
R14381 gnd.n3459 gnd.n3456 104.615
R14382 gnd.n3443 gnd.n3442 104.615
R14383 gnd.n3442 gnd.n3420 104.615
R14384 gnd.n3435 gnd.n3420 104.615
R14385 gnd.n3435 gnd.n3434 104.615
R14386 gnd.n3434 gnd.n3424 104.615
R14387 gnd.n3427 gnd.n3424 104.615
R14388 gnd.n3411 gnd.n3410 104.615
R14389 gnd.n3410 gnd.n3388 104.615
R14390 gnd.n3403 gnd.n3388 104.615
R14391 gnd.n3403 gnd.n3402 104.615
R14392 gnd.n3402 gnd.n3392 104.615
R14393 gnd.n3395 gnd.n3392 104.615
R14394 gnd.n3379 gnd.n3378 104.615
R14395 gnd.n3378 gnd.n3356 104.615
R14396 gnd.n3371 gnd.n3356 104.615
R14397 gnd.n3371 gnd.n3370 104.615
R14398 gnd.n3370 gnd.n3360 104.615
R14399 gnd.n3363 gnd.n3360 104.615
R14400 gnd.n3348 gnd.n3347 104.615
R14401 gnd.n3347 gnd.n3325 104.615
R14402 gnd.n3340 gnd.n3325 104.615
R14403 gnd.n3340 gnd.n3339 104.615
R14404 gnd.n3339 gnd.n3329 104.615
R14405 gnd.n3332 gnd.n3329 104.615
R14406 gnd.n2722 gnd.t73 100.632
R14407 gnd.n2280 gnd.t134 100.632
R14408 gnd.n7185 gnd.n7184 99.6594
R14409 gnd.n7180 gnd.n7001 99.6594
R14410 gnd.n7176 gnd.n7000 99.6594
R14411 gnd.n7172 gnd.n6999 99.6594
R14412 gnd.n7168 gnd.n6998 99.6594
R14413 gnd.n7164 gnd.n6997 99.6594
R14414 gnd.n7160 gnd.n6996 99.6594
R14415 gnd.n7156 gnd.n6995 99.6594
R14416 gnd.n7149 gnd.n6994 99.6594
R14417 gnd.n7145 gnd.n6993 99.6594
R14418 gnd.n7141 gnd.n6992 99.6594
R14419 gnd.n7137 gnd.n6991 99.6594
R14420 gnd.n7133 gnd.n6990 99.6594
R14421 gnd.n7129 gnd.n6989 99.6594
R14422 gnd.n7125 gnd.n6988 99.6594
R14423 gnd.n7121 gnd.n6987 99.6594
R14424 gnd.n7117 gnd.n6986 99.6594
R14425 gnd.n7113 gnd.n6985 99.6594
R14426 gnd.n7105 gnd.n6984 99.6594
R14427 gnd.n7103 gnd.n6983 99.6594
R14428 gnd.n7099 gnd.n6982 99.6594
R14429 gnd.n7095 gnd.n6981 99.6594
R14430 gnd.n7091 gnd.n6980 99.6594
R14431 gnd.n7087 gnd.n6979 99.6594
R14432 gnd.n7083 gnd.n6978 99.6594
R14433 gnd.n7079 gnd.n6977 99.6594
R14434 gnd.n7075 gnd.n6976 99.6594
R14435 gnd.n7071 gnd.n6975 99.6594
R14436 gnd.n7063 gnd.n6974 99.6594
R14437 gnd.n5585 gnd.n5584 99.6594
R14438 gnd.n5579 gnd.n1382 99.6594
R14439 gnd.n5576 gnd.n1383 99.6594
R14440 gnd.n5572 gnd.n1384 99.6594
R14441 gnd.n5568 gnd.n1385 99.6594
R14442 gnd.n5564 gnd.n1386 99.6594
R14443 gnd.n5560 gnd.n1387 99.6594
R14444 gnd.n5556 gnd.n1388 99.6594
R14445 gnd.n5552 gnd.n1389 99.6594
R14446 gnd.n5547 gnd.n1390 99.6594
R14447 gnd.n5543 gnd.n1391 99.6594
R14448 gnd.n5539 gnd.n1392 99.6594
R14449 gnd.n5535 gnd.n1393 99.6594
R14450 gnd.n5530 gnd.n1395 99.6594
R14451 gnd.n5526 gnd.n1396 99.6594
R14452 gnd.n5522 gnd.n1397 99.6594
R14453 gnd.n5518 gnd.n1398 99.6594
R14454 gnd.n5514 gnd.n1399 99.6594
R14455 gnd.n5510 gnd.n1400 99.6594
R14456 gnd.n5506 gnd.n1401 99.6594
R14457 gnd.n5502 gnd.n1402 99.6594
R14458 gnd.n5498 gnd.n1403 99.6594
R14459 gnd.n5494 gnd.n1404 99.6594
R14460 gnd.n5490 gnd.n1405 99.6594
R14461 gnd.n5486 gnd.n1406 99.6594
R14462 gnd.n5482 gnd.n1407 99.6594
R14463 gnd.n5478 gnd.n1408 99.6594
R14464 gnd.n5474 gnd.n1409 99.6594
R14465 gnd.n5901 gnd.n5900 99.6594
R14466 gnd.n5896 gnd.n1007 99.6594
R14467 gnd.n5892 gnd.n1006 99.6594
R14468 gnd.n5888 gnd.n1005 99.6594
R14469 gnd.n5884 gnd.n1004 99.6594
R14470 gnd.n5880 gnd.n1003 99.6594
R14471 gnd.n5876 gnd.n1002 99.6594
R14472 gnd.n5872 gnd.n1001 99.6594
R14473 gnd.n5867 gnd.n1000 99.6594
R14474 gnd.n5863 gnd.n999 99.6594
R14475 gnd.n5859 gnd.n998 99.6594
R14476 gnd.n5855 gnd.n997 99.6594
R14477 gnd.n1133 gnd.n995 99.6594
R14478 gnd.n1131 gnd.n994 99.6594
R14479 gnd.n1127 gnd.n993 99.6594
R14480 gnd.n1123 gnd.n992 99.6594
R14481 gnd.n1119 gnd.n991 99.6594
R14482 gnd.n1111 gnd.n990 99.6594
R14483 gnd.n1109 gnd.n989 99.6594
R14484 gnd.n1105 gnd.n988 99.6594
R14485 gnd.n1101 gnd.n987 99.6594
R14486 gnd.n1097 gnd.n986 99.6594
R14487 gnd.n1093 gnd.n985 99.6594
R14488 gnd.n1089 gnd.n984 99.6594
R14489 gnd.n1085 gnd.n983 99.6594
R14490 gnd.n1081 gnd.n982 99.6594
R14491 gnd.n1077 gnd.n981 99.6594
R14492 gnd.n1069 gnd.n980 99.6594
R14493 gnd.n3989 gnd.n3781 99.6594
R14494 gnd.n3987 gnd.n3784 99.6594
R14495 gnd.n3983 gnd.n3982 99.6594
R14496 gnd.n3976 gnd.n3789 99.6594
R14497 gnd.n3975 gnd.n3974 99.6594
R14498 gnd.n3968 gnd.n3795 99.6594
R14499 gnd.n3967 gnd.n3966 99.6594
R14500 gnd.n3960 gnd.n3801 99.6594
R14501 gnd.n3959 gnd.n3958 99.6594
R14502 gnd.n3952 gnd.n3807 99.6594
R14503 gnd.n3951 gnd.n3950 99.6594
R14504 gnd.n3944 gnd.n3816 99.6594
R14505 gnd.n3943 gnd.n3942 99.6594
R14506 gnd.n3936 gnd.n3822 99.6594
R14507 gnd.n3935 gnd.n3934 99.6594
R14508 gnd.n3928 gnd.n3828 99.6594
R14509 gnd.n3927 gnd.n3926 99.6594
R14510 gnd.n3920 gnd.n3834 99.6594
R14511 gnd.n3919 gnd.n3918 99.6594
R14512 gnd.n3912 gnd.n3842 99.6594
R14513 gnd.n3911 gnd.n3910 99.6594
R14514 gnd.n3904 gnd.n3848 99.6594
R14515 gnd.n3903 gnd.n3902 99.6594
R14516 gnd.n3896 gnd.n3854 99.6594
R14517 gnd.n3895 gnd.n3894 99.6594
R14518 gnd.n3888 gnd.n3860 99.6594
R14519 gnd.n3887 gnd.n3886 99.6594
R14520 gnd.n3880 gnd.n3866 99.6594
R14521 gnd.n3879 gnd.n3878 99.6594
R14522 gnd.n3693 gnd.n2263 99.6594
R14523 gnd.n3691 gnd.n2262 99.6594
R14524 gnd.n3687 gnd.n2261 99.6594
R14525 gnd.n3683 gnd.n2260 99.6594
R14526 gnd.n3679 gnd.n2259 99.6594
R14527 gnd.n3675 gnd.n2258 99.6594
R14528 gnd.n3671 gnd.n2257 99.6594
R14529 gnd.n3603 gnd.n2256 99.6594
R14530 gnd.n2934 gnd.n2665 99.6594
R14531 gnd.n2691 gnd.n2672 99.6594
R14532 gnd.n2693 gnd.n2673 99.6594
R14533 gnd.n2701 gnd.n2674 99.6594
R14534 gnd.n2703 gnd.n2675 99.6594
R14535 gnd.n2711 gnd.n2676 99.6594
R14536 gnd.n2713 gnd.n2677 99.6594
R14537 gnd.n2721 gnd.n2678 99.6594
R14538 gnd.n6937 gnd.n6916 99.6594
R14539 gnd.n6943 gnd.n6917 99.6594
R14540 gnd.n6947 gnd.n6918 99.6594
R14541 gnd.n6953 gnd.n6919 99.6594
R14542 gnd.n6957 gnd.n6920 99.6594
R14543 gnd.n6963 gnd.n6921 99.6594
R14544 gnd.n6966 gnd.n6922 99.6594
R14545 gnd.n6973 gnd.n6972 99.6594
R14546 gnd.n7188 gnd.n7187 99.6594
R14547 gnd.n1494 gnd.n1410 99.6594
R14548 gnd.n1412 gnd.n1336 99.6594
R14549 gnd.n1413 gnd.n1343 99.6594
R14550 gnd.n1415 gnd.n1414 99.6594
R14551 gnd.n1417 gnd.n1352 99.6594
R14552 gnd.n1418 gnd.n1359 99.6594
R14553 gnd.n1420 gnd.n1419 99.6594
R14554 gnd.n1422 gnd.n1368 99.6594
R14555 gnd.n5587 gnd.n1377 99.6594
R14556 gnd.n3661 gnd.n2243 99.6594
R14557 gnd.n3657 gnd.n2244 99.6594
R14558 gnd.n3653 gnd.n2245 99.6594
R14559 gnd.n3649 gnd.n2246 99.6594
R14560 gnd.n3645 gnd.n2247 99.6594
R14561 gnd.n3641 gnd.n2248 99.6594
R14562 gnd.n3637 gnd.n2249 99.6594
R14563 gnd.n3633 gnd.n2250 99.6594
R14564 gnd.n3629 gnd.n2251 99.6594
R14565 gnd.n3625 gnd.n2252 99.6594
R14566 gnd.n3621 gnd.n2253 99.6594
R14567 gnd.n3617 gnd.n2254 99.6594
R14568 gnd.n3613 gnd.n2255 99.6594
R14569 gnd.n2849 gnd.n2848 99.6594
R14570 gnd.n2843 gnd.n2760 99.6594
R14571 gnd.n2840 gnd.n2761 99.6594
R14572 gnd.n2836 gnd.n2762 99.6594
R14573 gnd.n2832 gnd.n2763 99.6594
R14574 gnd.n2828 gnd.n2764 99.6594
R14575 gnd.n2824 gnd.n2765 99.6594
R14576 gnd.n2820 gnd.n2766 99.6594
R14577 gnd.n2816 gnd.n2767 99.6594
R14578 gnd.n2812 gnd.n2768 99.6594
R14579 gnd.n2808 gnd.n2769 99.6594
R14580 gnd.n2804 gnd.n2770 99.6594
R14581 gnd.n2851 gnd.n2759 99.6594
R14582 gnd.n966 gnd.n911 99.6594
R14583 gnd.n968 gnd.n920 99.6594
R14584 gnd.n970 gnd.n969 99.6594
R14585 gnd.n971 gnd.n929 99.6594
R14586 gnd.n973 gnd.n938 99.6594
R14587 gnd.n975 gnd.n974 99.6594
R14588 gnd.n976 gnd.n947 99.6594
R14589 gnd.n978 gnd.n959 99.6594
R14590 gnd.n5904 gnd.n5903 99.6594
R14591 gnd.n3729 gnd.n2240 99.6594
R14592 gnd.n3732 gnd.n3731 99.6594
R14593 gnd.n3739 gnd.n3738 99.6594
R14594 gnd.n3742 gnd.n3741 99.6594
R14595 gnd.n3749 gnd.n3748 99.6594
R14596 gnd.n3752 gnd.n3751 99.6594
R14597 gnd.n3759 gnd.n3758 99.6594
R14598 gnd.n3762 gnd.n3761 99.6594
R14599 gnd.n3769 gnd.n3768 99.6594
R14600 gnd.n3730 gnd.n3729 99.6594
R14601 gnd.n3731 gnd.n3723 99.6594
R14602 gnd.n3740 gnd.n3739 99.6594
R14603 gnd.n3741 gnd.n3719 99.6594
R14604 gnd.n3750 gnd.n3749 99.6594
R14605 gnd.n3751 gnd.n3715 99.6594
R14606 gnd.n3760 gnd.n3759 99.6594
R14607 gnd.n3761 gnd.n3711 99.6594
R14608 gnd.n3770 gnd.n3769 99.6594
R14609 gnd.n5903 gnd.n964 99.6594
R14610 gnd.n978 gnd.n977 99.6594
R14611 gnd.n976 gnd.n946 99.6594
R14612 gnd.n975 gnd.n939 99.6594
R14613 gnd.n973 gnd.n972 99.6594
R14614 gnd.n971 gnd.n928 99.6594
R14615 gnd.n970 gnd.n921 99.6594
R14616 gnd.n968 gnd.n967 99.6594
R14617 gnd.n966 gnd.n910 99.6594
R14618 gnd.n2849 gnd.n2772 99.6594
R14619 gnd.n2841 gnd.n2760 99.6594
R14620 gnd.n2837 gnd.n2761 99.6594
R14621 gnd.n2833 gnd.n2762 99.6594
R14622 gnd.n2829 gnd.n2763 99.6594
R14623 gnd.n2825 gnd.n2764 99.6594
R14624 gnd.n2821 gnd.n2765 99.6594
R14625 gnd.n2817 gnd.n2766 99.6594
R14626 gnd.n2813 gnd.n2767 99.6594
R14627 gnd.n2809 gnd.n2768 99.6594
R14628 gnd.n2805 gnd.n2769 99.6594
R14629 gnd.n2801 gnd.n2770 99.6594
R14630 gnd.n2852 gnd.n2851 99.6594
R14631 gnd.n3616 gnd.n2255 99.6594
R14632 gnd.n3620 gnd.n2254 99.6594
R14633 gnd.n3624 gnd.n2253 99.6594
R14634 gnd.n3628 gnd.n2252 99.6594
R14635 gnd.n3632 gnd.n2251 99.6594
R14636 gnd.n3636 gnd.n2250 99.6594
R14637 gnd.n3640 gnd.n2249 99.6594
R14638 gnd.n3644 gnd.n2248 99.6594
R14639 gnd.n3648 gnd.n2247 99.6594
R14640 gnd.n3652 gnd.n2246 99.6594
R14641 gnd.n3656 gnd.n2245 99.6594
R14642 gnd.n3660 gnd.n2244 99.6594
R14643 gnd.n2284 gnd.n2243 99.6594
R14644 gnd.n1410 gnd.n1335 99.6594
R14645 gnd.n1412 gnd.n1411 99.6594
R14646 gnd.n1413 gnd.n1344 99.6594
R14647 gnd.n1415 gnd.n1351 99.6594
R14648 gnd.n1417 gnd.n1416 99.6594
R14649 gnd.n1418 gnd.n1360 99.6594
R14650 gnd.n1420 gnd.n1367 99.6594
R14651 gnd.n1422 gnd.n1421 99.6594
R14652 gnd.n5588 gnd.n5587 99.6594
R14653 gnd.n7187 gnd.n6915 99.6594
R14654 gnd.n6973 gnd.n6923 99.6594
R14655 gnd.n6964 gnd.n6922 99.6594
R14656 gnd.n6956 gnd.n6921 99.6594
R14657 gnd.n6954 gnd.n6920 99.6594
R14658 gnd.n6946 gnd.n6919 99.6594
R14659 gnd.n6944 gnd.n6918 99.6594
R14660 gnd.n6936 gnd.n6917 99.6594
R14661 gnd.n6934 gnd.n6916 99.6594
R14662 gnd.n2935 gnd.n2934 99.6594
R14663 gnd.n2694 gnd.n2672 99.6594
R14664 gnd.n2700 gnd.n2673 99.6594
R14665 gnd.n2704 gnd.n2674 99.6594
R14666 gnd.n2710 gnd.n2675 99.6594
R14667 gnd.n2714 gnd.n2676 99.6594
R14668 gnd.n2720 gnd.n2677 99.6594
R14669 gnd.n2678 gnd.n2662 99.6594
R14670 gnd.n3670 gnd.n2256 99.6594
R14671 gnd.n3674 gnd.n2257 99.6594
R14672 gnd.n3678 gnd.n2258 99.6594
R14673 gnd.n3682 gnd.n2259 99.6594
R14674 gnd.n3686 gnd.n2260 99.6594
R14675 gnd.n3690 gnd.n2261 99.6594
R14676 gnd.n3694 gnd.n2262 99.6594
R14677 gnd.n2265 gnd.n2263 99.6594
R14678 gnd.n3990 gnd.n3989 99.6594
R14679 gnd.n3984 gnd.n3784 99.6594
R14680 gnd.n3982 gnd.n3981 99.6594
R14681 gnd.n3977 gnd.n3976 99.6594
R14682 gnd.n3974 gnd.n3973 99.6594
R14683 gnd.n3969 gnd.n3968 99.6594
R14684 gnd.n3966 gnd.n3965 99.6594
R14685 gnd.n3961 gnd.n3960 99.6594
R14686 gnd.n3958 gnd.n3957 99.6594
R14687 gnd.n3953 gnd.n3952 99.6594
R14688 gnd.n3950 gnd.n3949 99.6594
R14689 gnd.n3945 gnd.n3944 99.6594
R14690 gnd.n3942 gnd.n3941 99.6594
R14691 gnd.n3937 gnd.n3936 99.6594
R14692 gnd.n3934 gnd.n3933 99.6594
R14693 gnd.n3929 gnd.n3928 99.6594
R14694 gnd.n3926 gnd.n3925 99.6594
R14695 gnd.n3921 gnd.n3920 99.6594
R14696 gnd.n3918 gnd.n3917 99.6594
R14697 gnd.n3913 gnd.n3912 99.6594
R14698 gnd.n3910 gnd.n3909 99.6594
R14699 gnd.n3905 gnd.n3904 99.6594
R14700 gnd.n3902 gnd.n3901 99.6594
R14701 gnd.n3897 gnd.n3896 99.6594
R14702 gnd.n3894 gnd.n3893 99.6594
R14703 gnd.n3889 gnd.n3888 99.6594
R14704 gnd.n3886 gnd.n3885 99.6594
R14705 gnd.n3881 gnd.n3880 99.6594
R14706 gnd.n3878 gnd.n3877 99.6594
R14707 gnd.n1076 gnd.n980 99.6594
R14708 gnd.n1080 gnd.n981 99.6594
R14709 gnd.n1084 gnd.n982 99.6594
R14710 gnd.n1088 gnd.n983 99.6594
R14711 gnd.n1092 gnd.n984 99.6594
R14712 gnd.n1096 gnd.n985 99.6594
R14713 gnd.n1100 gnd.n986 99.6594
R14714 gnd.n1104 gnd.n987 99.6594
R14715 gnd.n1108 gnd.n988 99.6594
R14716 gnd.n1112 gnd.n989 99.6594
R14717 gnd.n1118 gnd.n990 99.6594
R14718 gnd.n1122 gnd.n991 99.6594
R14719 gnd.n1126 gnd.n992 99.6594
R14720 gnd.n1130 gnd.n993 99.6594
R14721 gnd.n1134 gnd.n994 99.6594
R14722 gnd.n5854 gnd.n996 99.6594
R14723 gnd.n5858 gnd.n997 99.6594
R14724 gnd.n5862 gnd.n998 99.6594
R14725 gnd.n5866 gnd.n999 99.6594
R14726 gnd.n5871 gnd.n1000 99.6594
R14727 gnd.n5875 gnd.n1001 99.6594
R14728 gnd.n5879 gnd.n1002 99.6594
R14729 gnd.n5883 gnd.n1003 99.6594
R14730 gnd.n5887 gnd.n1004 99.6594
R14731 gnd.n5891 gnd.n1005 99.6594
R14732 gnd.n5895 gnd.n1006 99.6594
R14733 gnd.n1009 gnd.n1007 99.6594
R14734 gnd.n5901 gnd.n1008 99.6594
R14735 gnd.n5585 gnd.n1425 99.6594
R14736 gnd.n5577 gnd.n1382 99.6594
R14737 gnd.n5573 gnd.n1383 99.6594
R14738 gnd.n5569 gnd.n1384 99.6594
R14739 gnd.n5565 gnd.n1385 99.6594
R14740 gnd.n5561 gnd.n1386 99.6594
R14741 gnd.n5557 gnd.n1387 99.6594
R14742 gnd.n5553 gnd.n1388 99.6594
R14743 gnd.n5548 gnd.n1389 99.6594
R14744 gnd.n5544 gnd.n1390 99.6594
R14745 gnd.n5540 gnd.n1391 99.6594
R14746 gnd.n5536 gnd.n1392 99.6594
R14747 gnd.n5531 gnd.n1394 99.6594
R14748 gnd.n5527 gnd.n1395 99.6594
R14749 gnd.n5523 gnd.n1396 99.6594
R14750 gnd.n5519 gnd.n1397 99.6594
R14751 gnd.n5515 gnd.n1398 99.6594
R14752 gnd.n5511 gnd.n1399 99.6594
R14753 gnd.n5507 gnd.n1400 99.6594
R14754 gnd.n5503 gnd.n1401 99.6594
R14755 gnd.n5499 gnd.n1402 99.6594
R14756 gnd.n5495 gnd.n1403 99.6594
R14757 gnd.n5491 gnd.n1404 99.6594
R14758 gnd.n5487 gnd.n1405 99.6594
R14759 gnd.n5483 gnd.n1406 99.6594
R14760 gnd.n5479 gnd.n1407 99.6594
R14761 gnd.n5475 gnd.n1408 99.6594
R14762 gnd.n5467 gnd.n1409 99.6594
R14763 gnd.n7070 gnd.n6974 99.6594
R14764 gnd.n7074 gnd.n6975 99.6594
R14765 gnd.n7078 gnd.n6976 99.6594
R14766 gnd.n7082 gnd.n6977 99.6594
R14767 gnd.n7086 gnd.n6978 99.6594
R14768 gnd.n7090 gnd.n6979 99.6594
R14769 gnd.n7094 gnd.n6980 99.6594
R14770 gnd.n7098 gnd.n6981 99.6594
R14771 gnd.n7102 gnd.n6982 99.6594
R14772 gnd.n7106 gnd.n6983 99.6594
R14773 gnd.n7112 gnd.n6984 99.6594
R14774 gnd.n7116 gnd.n6985 99.6594
R14775 gnd.n7120 gnd.n6986 99.6594
R14776 gnd.n7124 gnd.n6987 99.6594
R14777 gnd.n7128 gnd.n6988 99.6594
R14778 gnd.n7132 gnd.n6989 99.6594
R14779 gnd.n7136 gnd.n6990 99.6594
R14780 gnd.n7140 gnd.n6991 99.6594
R14781 gnd.n7144 gnd.n6992 99.6594
R14782 gnd.n7148 gnd.n6993 99.6594
R14783 gnd.n7155 gnd.n6994 99.6594
R14784 gnd.n7159 gnd.n6995 99.6594
R14785 gnd.n7163 gnd.n6996 99.6594
R14786 gnd.n7167 gnd.n6997 99.6594
R14787 gnd.n7171 gnd.n6998 99.6594
R14788 gnd.n7175 gnd.n6999 99.6594
R14789 gnd.n7179 gnd.n7000 99.6594
R14790 gnd.n7003 gnd.n7001 99.6594
R14791 gnd.n7185 gnd.n7002 99.6594
R14792 gnd.n5966 gnd.n5965 99.6594
R14793 gnd.n897 gnd.n877 99.6594
R14794 gnd.n899 gnd.n878 99.6594
R14795 gnd.n903 gnd.n879 99.6594
R14796 gnd.n905 gnd.n880 99.6594
R14797 gnd.n915 gnd.n881 99.6594
R14798 gnd.n917 gnd.n882 99.6594
R14799 gnd.n925 gnd.n883 99.6594
R14800 gnd.n933 gnd.n884 99.6594
R14801 gnd.n935 gnd.n885 99.6594
R14802 gnd.n943 gnd.n886 99.6594
R14803 gnd.n951 gnd.n887 99.6594
R14804 gnd.n956 gnd.n889 99.6594
R14805 gnd.n5968 gnd.n874 99.6594
R14806 gnd.n5966 gnd.n892 99.6594
R14807 gnd.n898 gnd.n877 99.6594
R14808 gnd.n902 gnd.n878 99.6594
R14809 gnd.n904 gnd.n879 99.6594
R14810 gnd.n914 gnd.n880 99.6594
R14811 gnd.n916 gnd.n881 99.6594
R14812 gnd.n924 gnd.n882 99.6594
R14813 gnd.n932 gnd.n883 99.6594
R14814 gnd.n934 gnd.n884 99.6594
R14815 gnd.n942 gnd.n885 99.6594
R14816 gnd.n950 gnd.n886 99.6594
R14817 gnd.n952 gnd.n887 99.6594
R14818 gnd.n889 gnd.n888 99.6594
R14819 gnd.n5969 gnd.n5968 99.6594
R14820 gnd.n1644 gnd.n1320 99.6594
R14821 gnd.n1646 gnd.n1645 99.6594
R14822 gnd.n1647 gnd.n1325 99.6594
R14823 gnd.n1649 gnd.n1648 99.6594
R14824 gnd.n1650 gnd.n1331 99.6594
R14825 gnd.n1652 gnd.n1339 99.6594
R14826 gnd.n1654 gnd.n1653 99.6594
R14827 gnd.n1655 gnd.n1348 99.6594
R14828 gnd.n1657 gnd.n1355 99.6594
R14829 gnd.n1659 gnd.n1658 99.6594
R14830 gnd.n1660 gnd.n1364 99.6594
R14831 gnd.n1662 gnd.n1371 99.6594
R14832 gnd.n1665 gnd.n1664 99.6594
R14833 gnd.n5261 gnd.n5260 99.6594
R14834 gnd.n1662 gnd.n1661 99.6594
R14835 gnd.n1660 gnd.n1363 99.6594
R14836 gnd.n1659 gnd.n1356 99.6594
R14837 gnd.n1657 gnd.n1656 99.6594
R14838 gnd.n1655 gnd.n1347 99.6594
R14839 gnd.n1654 gnd.n1340 99.6594
R14840 gnd.n1652 gnd.n1651 99.6594
R14841 gnd.n1650 gnd.n1330 99.6594
R14842 gnd.n1649 gnd.n1326 99.6594
R14843 gnd.n1647 gnd.n1324 99.6594
R14844 gnd.n1646 gnd.n1321 99.6594
R14845 gnd.n1644 gnd.n1316 99.6594
R14846 gnd.n5260 gnd.n1311 99.6594
R14847 gnd.n1665 gnd.n1643 99.6594
R14848 gnd.n953 gnd.t66 98.63
R14849 gnd.n5589 gnd.t33 98.63
R14850 gnd.n960 gnd.t61 98.63
R14851 gnd.n1445 gnd.t121 98.63
R14852 gnd.n1468 gnd.t124 98.63
R14853 gnd.n5469 gnd.t85 98.63
R14854 gnd.n7065 gnd.t81 98.63
R14855 gnd.n7044 gnd.t87 98.63
R14856 gnd.n7151 gnd.t105 98.63
R14857 gnd.n6912 gnd.t28 98.63
R14858 gnd.n3808 gnd.t69 98.63
R14859 gnd.n3839 gnd.t103 98.63
R14860 gnd.n3871 gnd.t115 98.63
R14861 gnd.n3708 gnd.t58 98.63
R14862 gnd.n1030 gnd.t96 98.63
R14863 gnd.n1071 gnd.t117 98.63
R14864 gnd.n1050 gnd.t137 98.63
R14865 gnd.n1373 gnd.t46 98.63
R14866 gnd.n4427 gnd.t100 96.6984
R14867 gnd.n1769 gnd.t53 96.6984
R14868 gnd.n5783 gnd.t25 96.6906
R14869 gnd.n5006 gnd.t108 96.6906
R14870 gnd.n6868 gnd.n170 86.3597
R14871 gnd.n1188 gnd.n1187 81.8399
R14872 gnd.n2723 gnd.t72 74.8376
R14873 gnd.n2281 gnd.t135 74.8376
R14874 gnd.n4428 gnd.t99 72.8438
R14875 gnd.n1770 gnd.t54 72.8438
R14876 gnd.n1189 gnd.n1182 72.8411
R14877 gnd.n1195 gnd.n1180 72.8411
R14878 gnd.n5002 gnd.n5001 72.8411
R14879 gnd.n954 gnd.t65 72.836
R14880 gnd.n5784 gnd.t24 72.836
R14881 gnd.n5007 gnd.t109 72.836
R14882 gnd.n5590 gnd.t32 72.836
R14883 gnd.n961 gnd.t62 72.836
R14884 gnd.n1446 gnd.t120 72.836
R14885 gnd.n1469 gnd.t123 72.836
R14886 gnd.n5470 gnd.t84 72.836
R14887 gnd.n7066 gnd.t82 72.836
R14888 gnd.n7045 gnd.t88 72.836
R14889 gnd.n7152 gnd.t106 72.836
R14890 gnd.n6913 gnd.t29 72.836
R14891 gnd.n3809 gnd.t68 72.836
R14892 gnd.n3840 gnd.t102 72.836
R14893 gnd.n3872 gnd.t114 72.836
R14894 gnd.n3709 gnd.t57 72.836
R14895 gnd.n1031 gnd.t97 72.836
R14896 gnd.n1072 gnd.t118 72.836
R14897 gnd.n1051 gnd.t138 72.836
R14898 gnd.n1374 gnd.t47 72.836
R14899 gnd.n5070 gnd.n1734 71.676
R14900 gnd.n5066 gnd.n1735 71.676
R14901 gnd.n5062 gnd.n1736 71.676
R14902 gnd.n5058 gnd.n1737 71.676
R14903 gnd.n5054 gnd.n1738 71.676
R14904 gnd.n5050 gnd.n1739 71.676
R14905 gnd.n5046 gnd.n1740 71.676
R14906 gnd.n5042 gnd.n1741 71.676
R14907 gnd.n5038 gnd.n1742 71.676
R14908 gnd.n5034 gnd.n1743 71.676
R14909 gnd.n5030 gnd.n1744 71.676
R14910 gnd.n5026 gnd.n1745 71.676
R14911 gnd.n5022 gnd.n1746 71.676
R14912 gnd.n5018 gnd.n1747 71.676
R14913 gnd.n5013 gnd.n1748 71.676
R14914 gnd.n5009 gnd.n1749 71.676
R14915 gnd.n5146 gnd.n1768 71.676
R14916 gnd.n5142 gnd.n1767 71.676
R14917 gnd.n5137 gnd.n1766 71.676
R14918 gnd.n5133 gnd.n1765 71.676
R14919 gnd.n5129 gnd.n1764 71.676
R14920 gnd.n5125 gnd.n1763 71.676
R14921 gnd.n5121 gnd.n1762 71.676
R14922 gnd.n5117 gnd.n1761 71.676
R14923 gnd.n5113 gnd.n1760 71.676
R14924 gnd.n5109 gnd.n1759 71.676
R14925 gnd.n5105 gnd.n1758 71.676
R14926 gnd.n5101 gnd.n1757 71.676
R14927 gnd.n5097 gnd.n1756 71.676
R14928 gnd.n5093 gnd.n1755 71.676
R14929 gnd.n5089 gnd.n1754 71.676
R14930 gnd.n5085 gnd.n1753 71.676
R14931 gnd.n5081 gnd.n1752 71.676
R14932 gnd.n5847 gnd.n5846 71.676
R14933 gnd.n5841 gnd.n1144 71.676
R14934 gnd.n5838 gnd.n1145 71.676
R14935 gnd.n5834 gnd.n1146 71.676
R14936 gnd.n5830 gnd.n1147 71.676
R14937 gnd.n5826 gnd.n1148 71.676
R14938 gnd.n5822 gnd.n1149 71.676
R14939 gnd.n5818 gnd.n1150 71.676
R14940 gnd.n5814 gnd.n1151 71.676
R14941 gnd.n5810 gnd.n1152 71.676
R14942 gnd.n5806 gnd.n1153 71.676
R14943 gnd.n5802 gnd.n1154 71.676
R14944 gnd.n5798 gnd.n1155 71.676
R14945 gnd.n5794 gnd.n1156 71.676
R14946 gnd.n5790 gnd.n1157 71.676
R14947 gnd.n5786 gnd.n1158 71.676
R14948 gnd.n1159 gnd.n1142 71.676
R14949 gnd.n4431 gnd.n1160 71.676
R14950 gnd.n4436 gnd.n1161 71.676
R14951 gnd.n4440 gnd.n1162 71.676
R14952 gnd.n4444 gnd.n1163 71.676
R14953 gnd.n4448 gnd.n1164 71.676
R14954 gnd.n4452 gnd.n1165 71.676
R14955 gnd.n4456 gnd.n1166 71.676
R14956 gnd.n4460 gnd.n1167 71.676
R14957 gnd.n4464 gnd.n1168 71.676
R14958 gnd.n4468 gnd.n1169 71.676
R14959 gnd.n4472 gnd.n1170 71.676
R14960 gnd.n4476 gnd.n1171 71.676
R14961 gnd.n4480 gnd.n1172 71.676
R14962 gnd.n4484 gnd.n1173 71.676
R14963 gnd.n4488 gnd.n1174 71.676
R14964 gnd.n5847 gnd.n1177 71.676
R14965 gnd.n5839 gnd.n1144 71.676
R14966 gnd.n5835 gnd.n1145 71.676
R14967 gnd.n5831 gnd.n1146 71.676
R14968 gnd.n5827 gnd.n1147 71.676
R14969 gnd.n5823 gnd.n1148 71.676
R14970 gnd.n5819 gnd.n1149 71.676
R14971 gnd.n5815 gnd.n1150 71.676
R14972 gnd.n5811 gnd.n1151 71.676
R14973 gnd.n5807 gnd.n1152 71.676
R14974 gnd.n5803 gnd.n1153 71.676
R14975 gnd.n5799 gnd.n1154 71.676
R14976 gnd.n5795 gnd.n1155 71.676
R14977 gnd.n5791 gnd.n1156 71.676
R14978 gnd.n5787 gnd.n1157 71.676
R14979 gnd.n5850 gnd.n5849 71.676
R14980 gnd.n4430 gnd.n1159 71.676
R14981 gnd.n4435 gnd.n1160 71.676
R14982 gnd.n4439 gnd.n1161 71.676
R14983 gnd.n4443 gnd.n1162 71.676
R14984 gnd.n4447 gnd.n1163 71.676
R14985 gnd.n4451 gnd.n1164 71.676
R14986 gnd.n4455 gnd.n1165 71.676
R14987 gnd.n4459 gnd.n1166 71.676
R14988 gnd.n4463 gnd.n1167 71.676
R14989 gnd.n4467 gnd.n1168 71.676
R14990 gnd.n4471 gnd.n1169 71.676
R14991 gnd.n4475 gnd.n1170 71.676
R14992 gnd.n4479 gnd.n1171 71.676
R14993 gnd.n4483 gnd.n1172 71.676
R14994 gnd.n4487 gnd.n1173 71.676
R14995 gnd.n4491 gnd.n1174 71.676
R14996 gnd.n5084 gnd.n1752 71.676
R14997 gnd.n5088 gnd.n1753 71.676
R14998 gnd.n5092 gnd.n1754 71.676
R14999 gnd.n5096 gnd.n1755 71.676
R15000 gnd.n5100 gnd.n1756 71.676
R15001 gnd.n5104 gnd.n1757 71.676
R15002 gnd.n5108 gnd.n1758 71.676
R15003 gnd.n5112 gnd.n1759 71.676
R15004 gnd.n5116 gnd.n1760 71.676
R15005 gnd.n5120 gnd.n1761 71.676
R15006 gnd.n5124 gnd.n1762 71.676
R15007 gnd.n5128 gnd.n1763 71.676
R15008 gnd.n5132 gnd.n1764 71.676
R15009 gnd.n5136 gnd.n1765 71.676
R15010 gnd.n5141 gnd.n1766 71.676
R15011 gnd.n5145 gnd.n1767 71.676
R15012 gnd.n5008 gnd.n1750 71.676
R15013 gnd.n5012 gnd.n1749 71.676
R15014 gnd.n5017 gnd.n1748 71.676
R15015 gnd.n5021 gnd.n1747 71.676
R15016 gnd.n5025 gnd.n1746 71.676
R15017 gnd.n5029 gnd.n1745 71.676
R15018 gnd.n5033 gnd.n1744 71.676
R15019 gnd.n5037 gnd.n1743 71.676
R15020 gnd.n5041 gnd.n1742 71.676
R15021 gnd.n5045 gnd.n1741 71.676
R15022 gnd.n5049 gnd.n1740 71.676
R15023 gnd.n5053 gnd.n1739 71.676
R15024 gnd.n5057 gnd.n1738 71.676
R15025 gnd.n5061 gnd.n1737 71.676
R15026 gnd.n5065 gnd.n1736 71.676
R15027 gnd.n5069 gnd.n1735 71.676
R15028 gnd.n5072 gnd.n1734 71.676
R15029 gnd.n10 gnd.t325 69.1507
R15030 gnd.n18 gnd.t289 68.4792
R15031 gnd.n17 gnd.t265 68.4792
R15032 gnd.n16 gnd.t267 68.4792
R15033 gnd.n15 gnd.t19 68.4792
R15034 gnd.n14 gnd.t321 68.4792
R15035 gnd.n13 gnd.t17 68.4792
R15036 gnd.n12 gnd.t323 68.4792
R15037 gnd.n11 gnd.t307 68.4792
R15038 gnd.n10 gnd.t316 68.4792
R15039 gnd.n2850 gnd.n2754 64.369
R15040 gnd.n3997 gnd.n3703 63.0944
R15041 gnd.n4433 gnd.n4428 59.5399
R15042 gnd.n5139 gnd.n1770 59.5399
R15043 gnd.n5785 gnd.n5784 59.5399
R15044 gnd.n5015 gnd.n5007 59.5399
R15045 gnd.n5782 gnd.n1198 59.1804
R15046 gnd.n3702 gnd.n2241 57.3586
R15047 gnd.n2509 gnd.t238 56.407
R15048 gnd.n2474 gnd.t253 56.407
R15049 gnd.n2485 gnd.t224 56.407
R15050 gnd.n2497 gnd.t159 56.407
R15051 gnd.n56 gnd.t216 56.407
R15052 gnd.n21 gnd.t165 56.407
R15053 gnd.n32 gnd.t204 56.407
R15054 gnd.n44 gnd.t247 56.407
R15055 gnd.n2518 gnd.t177 55.8337
R15056 gnd.n2483 gnd.t248 55.8337
R15057 gnd.n2494 gnd.t215 55.8337
R15058 gnd.n2506 gnd.t228 55.8337
R15059 gnd.n65 gnd.t255 55.8337
R15060 gnd.n30 gnd.t151 55.8337
R15061 gnd.n41 gnd.t193 55.8337
R15062 gnd.n53 gnd.t195 55.8337
R15063 gnd.n7186 gnd.n170 55.7653
R15064 gnd.n1186 gnd.n1185 54.358
R15065 gnd.n4999 gnd.n4998 54.358
R15066 gnd.n2509 gnd.n2508 53.0052
R15067 gnd.n2511 gnd.n2510 53.0052
R15068 gnd.n2513 gnd.n2512 53.0052
R15069 gnd.n2515 gnd.n2514 53.0052
R15070 gnd.n2517 gnd.n2516 53.0052
R15071 gnd.n2474 gnd.n2473 53.0052
R15072 gnd.n2476 gnd.n2475 53.0052
R15073 gnd.n2478 gnd.n2477 53.0052
R15074 gnd.n2480 gnd.n2479 53.0052
R15075 gnd.n2482 gnd.n2481 53.0052
R15076 gnd.n2485 gnd.n2484 53.0052
R15077 gnd.n2487 gnd.n2486 53.0052
R15078 gnd.n2489 gnd.n2488 53.0052
R15079 gnd.n2491 gnd.n2490 53.0052
R15080 gnd.n2493 gnd.n2492 53.0052
R15081 gnd.n2497 gnd.n2496 53.0052
R15082 gnd.n2499 gnd.n2498 53.0052
R15083 gnd.n2501 gnd.n2500 53.0052
R15084 gnd.n2503 gnd.n2502 53.0052
R15085 gnd.n2505 gnd.n2504 53.0052
R15086 gnd.n64 gnd.n63 53.0052
R15087 gnd.n62 gnd.n61 53.0052
R15088 gnd.n60 gnd.n59 53.0052
R15089 gnd.n58 gnd.n57 53.0052
R15090 gnd.n56 gnd.n55 53.0052
R15091 gnd.n29 gnd.n28 53.0052
R15092 gnd.n27 gnd.n26 53.0052
R15093 gnd.n25 gnd.n24 53.0052
R15094 gnd.n23 gnd.n22 53.0052
R15095 gnd.n21 gnd.n20 53.0052
R15096 gnd.n40 gnd.n39 53.0052
R15097 gnd.n38 gnd.n37 53.0052
R15098 gnd.n36 gnd.n35 53.0052
R15099 gnd.n34 gnd.n33 53.0052
R15100 gnd.n32 gnd.n31 53.0052
R15101 gnd.n52 gnd.n51 53.0052
R15102 gnd.n50 gnd.n49 53.0052
R15103 gnd.n48 gnd.n47 53.0052
R15104 gnd.n46 gnd.n45 53.0052
R15105 gnd.n44 gnd.n43 53.0052
R15106 gnd.n4990 gnd.n4989 52.4801
R15107 gnd.n3554 gnd.t293 52.3082
R15108 gnd.n3522 gnd.t269 52.3082
R15109 gnd.n3490 gnd.t10 52.3082
R15110 gnd.n3459 gnd.t143 52.3082
R15111 gnd.n3427 gnd.t6 52.3082
R15112 gnd.n3395 gnd.t12 52.3082
R15113 gnd.n3363 gnd.t327 52.3082
R15114 gnd.n3332 gnd.t291 52.3082
R15115 gnd.n3384 gnd.n3352 51.4173
R15116 gnd.n3448 gnd.n3447 50.455
R15117 gnd.n3416 gnd.n3415 50.455
R15118 gnd.n3384 gnd.n3383 50.455
R15119 gnd.n2797 gnd.n2796 45.1884
R15120 gnd.n2307 gnd.n2306 45.1884
R15121 gnd.n5074 gnd.n5005 44.3322
R15122 gnd.n1189 gnd.n1188 44.3189
R15123 gnd.n955 gnd.n954 42.4732
R15124 gnd.n1375 gnd.n1374 42.4732
R15125 gnd.n5591 gnd.n5590 42.2793
R15126 gnd.n2798 gnd.n2797 42.2793
R15127 gnd.n2308 gnd.n2307 42.2793
R15128 gnd.n2724 gnd.n2723 42.2793
R15129 gnd.n3669 gnd.n2281 42.2793
R15130 gnd.n5906 gnd.n961 42.2793
R15131 gnd.n5550 gnd.n1446 42.2793
R15132 gnd.n5513 gnd.n1469 42.2793
R15133 gnd.n5473 gnd.n5470 42.2793
R15134 gnd.n7069 gnd.n7066 42.2793
R15135 gnd.n7111 gnd.n7045 42.2793
R15136 gnd.n7153 gnd.n7152 42.2793
R15137 gnd.n6914 gnd.n6913 42.2793
R15138 gnd.n3810 gnd.n3809 42.2793
R15139 gnd.n3841 gnd.n3840 42.2793
R15140 gnd.n3873 gnd.n3872 42.2793
R15141 gnd.n3710 gnd.n3709 42.2793
R15142 gnd.n5869 gnd.n1031 42.2793
R15143 gnd.n1075 gnd.n1072 42.2793
R15144 gnd.n1117 gnd.n1051 42.2793
R15145 gnd.n1187 gnd.n1186 41.6274
R15146 gnd.n5000 gnd.n4999 41.6274
R15147 gnd.n1196 gnd.n1195 40.8975
R15148 gnd.n5003 gnd.n5002 40.8975
R15149 gnd.n6237 gnd.n561 37.8532
R15150 gnd.n6237 gnd.n6236 37.8532
R15151 gnd.n6236 gnd.n6235 37.8532
R15152 gnd.n6235 gnd.n566 37.8532
R15153 gnd.n6229 gnd.n566 37.8532
R15154 gnd.n6229 gnd.n6228 37.8532
R15155 gnd.n6228 gnd.n6227 37.8532
R15156 gnd.n6227 gnd.n574 37.8532
R15157 gnd.n6221 gnd.n574 37.8532
R15158 gnd.n6221 gnd.n6220 37.8532
R15159 gnd.n6220 gnd.n6219 37.8532
R15160 gnd.n6219 gnd.n582 37.8532
R15161 gnd.n6213 gnd.n582 37.8532
R15162 gnd.n6213 gnd.n6212 37.8532
R15163 gnd.n6212 gnd.n6211 37.8532
R15164 gnd.n6211 gnd.n590 37.8532
R15165 gnd.n6205 gnd.n590 37.8532
R15166 gnd.n6205 gnd.n6204 37.8532
R15167 gnd.n6204 gnd.n6203 37.8532
R15168 gnd.n6203 gnd.n598 37.8532
R15169 gnd.n6197 gnd.n598 37.8532
R15170 gnd.n6197 gnd.n6196 37.8532
R15171 gnd.n6196 gnd.n6195 37.8532
R15172 gnd.n6195 gnd.n606 37.8532
R15173 gnd.n6189 gnd.n606 37.8532
R15174 gnd.n6189 gnd.n6188 37.8532
R15175 gnd.n6188 gnd.n6187 37.8532
R15176 gnd.n6187 gnd.n614 37.8532
R15177 gnd.n6181 gnd.n614 37.8532
R15178 gnd.n6181 gnd.n6180 37.8532
R15179 gnd.n6180 gnd.n6179 37.8532
R15180 gnd.n6179 gnd.n622 37.8532
R15181 gnd.n6173 gnd.n622 37.8532
R15182 gnd.n6173 gnd.n6172 37.8532
R15183 gnd.n6172 gnd.n6171 37.8532
R15184 gnd.n6171 gnd.n630 37.8532
R15185 gnd.n6165 gnd.n630 37.8532
R15186 gnd.n6165 gnd.n6164 37.8532
R15187 gnd.n6164 gnd.n6163 37.8532
R15188 gnd.n6163 gnd.n638 37.8532
R15189 gnd.n6157 gnd.n638 37.8532
R15190 gnd.n6157 gnd.n6156 37.8532
R15191 gnd.n6156 gnd.n6155 37.8532
R15192 gnd.n6155 gnd.n646 37.8532
R15193 gnd.n6149 gnd.n646 37.8532
R15194 gnd.n6149 gnd.n6148 37.8532
R15195 gnd.n6148 gnd.n6147 37.8532
R15196 gnd.n6147 gnd.n654 37.8532
R15197 gnd.n6141 gnd.n654 37.8532
R15198 gnd.n6141 gnd.n6140 37.8532
R15199 gnd.n6140 gnd.n6139 37.8532
R15200 gnd.n6139 gnd.n662 37.8532
R15201 gnd.n6133 gnd.n662 37.8532
R15202 gnd.n6133 gnd.n6132 37.8532
R15203 gnd.n6132 gnd.n6131 37.8532
R15204 gnd.n6131 gnd.n670 37.8532
R15205 gnd.n6125 gnd.n670 37.8532
R15206 gnd.n6125 gnd.n6124 37.8532
R15207 gnd.n6124 gnd.n6123 37.8532
R15208 gnd.n6123 gnd.n678 37.8532
R15209 gnd.n6117 gnd.n678 37.8532
R15210 gnd.n6117 gnd.n6116 37.8532
R15211 gnd.n6116 gnd.n6115 37.8532
R15212 gnd.n6115 gnd.n686 37.8532
R15213 gnd.n6109 gnd.n686 37.8532
R15214 gnd.n6109 gnd.n6108 37.8532
R15215 gnd.n6108 gnd.n6107 37.8532
R15216 gnd.n6107 gnd.n694 37.8532
R15217 gnd.n6101 gnd.n694 37.8532
R15218 gnd.n6101 gnd.n6100 37.8532
R15219 gnd.n6100 gnd.n6099 37.8532
R15220 gnd.n6099 gnd.n702 37.8532
R15221 gnd.n6093 gnd.n702 37.8532
R15222 gnd.n6093 gnd.n6092 37.8532
R15223 gnd.n6092 gnd.n6091 37.8532
R15224 gnd.n6091 gnd.n710 37.8532
R15225 gnd.n6085 gnd.n710 37.8532
R15226 gnd.n6085 gnd.n6084 37.8532
R15227 gnd.n6084 gnd.n6083 37.8532
R15228 gnd.n6083 gnd.n718 37.8532
R15229 gnd.n6077 gnd.n718 37.8532
R15230 gnd.n6077 gnd.n6076 37.8532
R15231 gnd.n6076 gnd.n6075 37.8532
R15232 gnd.n1195 gnd.n1194 35.055
R15233 gnd.n1190 gnd.n1189 35.055
R15234 gnd.n4992 gnd.n4991 35.055
R15235 gnd.n5002 gnd.n4988 35.055
R15236 gnd.n5082 gnd.n1771 33.2493
R15237 gnd.n4494 gnd.n4490 33.2493
R15238 gnd.n2860 gnd.n2754 31.8661
R15239 gnd.n2860 gnd.n2859 31.8661
R15240 gnd.n2868 gnd.n2743 31.8661
R15241 gnd.n2876 gnd.n2743 31.8661
R15242 gnd.n2876 gnd.n2737 31.8661
R15243 gnd.n2884 gnd.n2737 31.8661
R15244 gnd.n2884 gnd.n2730 31.8661
R15245 gnd.n2922 gnd.n2730 31.8661
R15246 gnd.n2932 gnd.n2663 31.8661
R15247 gnd.n3997 gnd.n3780 31.8661
R15248 gnd.n4015 gnd.n2221 31.8661
R15249 gnd.n4025 gnd.n2221 31.8661
R15250 gnd.n4025 gnd.n2215 31.8661
R15251 gnd.n4035 gnd.n2215 31.8661
R15252 gnd.n4050 gnd.n2196 31.8661
R15253 gnd.n4060 gnd.n2196 31.8661
R15254 gnd.n4072 gnd.n2190 31.8661
R15255 gnd.n4090 gnd.n2180 31.8661
R15256 gnd.n965 gnd.n862 31.8661
R15257 gnd.n4252 gnd.n979 31.8661
R15258 gnd.n4252 gnd.n876 31.8661
R15259 gnd.n4261 gnd.n890 31.8661
R15260 gnd.n4312 gnd.n4261 31.8661
R15261 gnd.n4321 gnd.n2104 31.8661
R15262 gnd.n4329 gnd.n2104 31.8661
R15263 gnd.n4329 gnd.n2097 31.8661
R15264 gnd.n4337 gnd.n2097 31.8661
R15265 gnd.n4345 gnd.n2090 31.8661
R15266 gnd.n4345 gnd.n2082 31.8661
R15267 gnd.n4353 gnd.n2082 31.8661
R15268 gnd.n4353 gnd.n2084 31.8661
R15269 gnd.n4361 gnd.n2068 31.8661
R15270 gnd.n4369 gnd.n2068 31.8661
R15271 gnd.n4369 gnd.n2070 31.8661
R15272 gnd.n4377 gnd.n2053 31.8661
R15273 gnd.n4399 gnd.n2053 31.8661
R15274 gnd.n4399 gnd.n2045 31.8661
R15275 gnd.n4413 gnd.n2045 31.8661
R15276 gnd.n5157 gnd.n1721 31.8661
R15277 gnd.n5166 gnd.n1721 31.8661
R15278 gnd.n5166 gnd.n1715 31.8661
R15279 gnd.n5174 gnd.n1715 31.8661
R15280 gnd.n5183 gnd.n1709 31.8661
R15281 gnd.n5183 gnd.n1703 31.8661
R15282 gnd.n5191 gnd.n1703 31.8661
R15283 gnd.n5200 gnd.n1697 31.8661
R15284 gnd.n5200 gnd.n1690 31.8661
R15285 gnd.n5208 gnd.n1690 31.8661
R15286 gnd.n5208 gnd.n1691 31.8661
R15287 gnd.n5217 gnd.n1679 31.8661
R15288 gnd.n5228 gnd.n1679 31.8661
R15289 gnd.n5228 gnd.n1673 31.8661
R15290 gnd.n5237 gnd.n1673 31.8661
R15291 gnd.n5654 gnd.n1312 31.8661
R15292 gnd.n5654 gnd.n1314 31.8661
R15293 gnd.n5258 gnd.n1666 31.8661
R15294 gnd.n1666 gnd.n1381 31.8661
R15295 gnd.n1491 gnd.n1423 31.8661
R15296 gnd.n7283 gnd.n111 31.8661
R15297 gnd.n7277 gnd.n120 31.8661
R15298 gnd.n7271 gnd.n130 31.8661
R15299 gnd.n7271 gnd.n133 31.8661
R15300 gnd.n7265 gnd.n142 31.8661
R15301 gnd.n7259 gnd.n142 31.8661
R15302 gnd.n7259 gnd.n152 31.8661
R15303 gnd.n7253 gnd.n152 31.8661
R15304 gnd.n7247 gnd.n167 31.8661
R15305 gnd.t152 gnd.n2190 30.9101
R15306 gnd.n7277 gnd.t172 30.9101
R15307 gnd.n5149 gnd.n1732 30.5915
R15308 gnd.n2070 gnd.t7 27.0862
R15309 gnd.t264 gnd.n1709 27.0862
R15310 gnd.n954 gnd.n953 25.7944
R15311 gnd.n5590 gnd.n5589 25.7944
R15312 gnd.n2723 gnd.n2722 25.7944
R15313 gnd.n2281 gnd.n2280 25.7944
R15314 gnd.n961 gnd.n960 25.7944
R15315 gnd.n1446 gnd.n1445 25.7944
R15316 gnd.n1469 gnd.n1468 25.7944
R15317 gnd.n5470 gnd.n5469 25.7944
R15318 gnd.n7066 gnd.n7065 25.7944
R15319 gnd.n7045 gnd.n7044 25.7944
R15320 gnd.n7152 gnd.n7151 25.7944
R15321 gnd.n6913 gnd.n6912 25.7944
R15322 gnd.n3809 gnd.n3808 25.7944
R15323 gnd.n3840 gnd.n3839 25.7944
R15324 gnd.n3872 gnd.n3871 25.7944
R15325 gnd.n3709 gnd.n3708 25.7944
R15326 gnd.n1031 gnd.n1030 25.7944
R15327 gnd.n1072 gnd.n1071 25.7944
R15328 gnd.n1051 gnd.n1050 25.7944
R15329 gnd.n1374 gnd.n1373 25.7944
R15330 gnd.n2944 gnd.n2664 24.8557
R15331 gnd.n2954 gnd.n2647 24.8557
R15332 gnd.n2650 gnd.n2638 24.8557
R15333 gnd.n2975 gnd.n2639 24.8557
R15334 gnd.n2985 gnd.n2619 24.8557
R15335 gnd.n2995 gnd.n2994 24.8557
R15336 gnd.n2605 gnd.n2603 24.8557
R15337 gnd.n3026 gnd.n3025 24.8557
R15338 gnd.n3041 gnd.n2588 24.8557
R15339 gnd.n3095 gnd.n2527 24.8557
R15340 gnd.n3051 gnd.n2528 24.8557
R15341 gnd.n3088 gnd.n2539 24.8557
R15342 gnd.n2577 gnd.n2576 24.8557
R15343 gnd.n3082 gnd.n3081 24.8557
R15344 gnd.n2563 gnd.n2550 24.8557
R15345 gnd.n3121 gnd.n3120 24.8557
R15346 gnd.n3131 gnd.n2459 24.8557
R15347 gnd.n3143 gnd.n2451 24.8557
R15348 gnd.n3142 gnd.n2439 24.8557
R15349 gnd.n3161 gnd.n3160 24.8557
R15350 gnd.n3171 gnd.n2432 24.8557
R15351 gnd.n3182 gnd.n2420 24.8557
R15352 gnd.n3206 gnd.n3205 24.8557
R15353 gnd.n3217 gnd.n2403 24.8557
R15354 gnd.n3216 gnd.n2405 24.8557
R15355 gnd.n3228 gnd.n2396 24.8557
R15356 gnd.n3246 gnd.n3245 24.8557
R15357 gnd.n2387 gnd.n2376 24.8557
R15358 gnd.n3267 gnd.n2364 24.8557
R15359 gnd.n3295 gnd.n3294 24.8557
R15360 gnd.n3306 gnd.n2349 24.8557
R15361 gnd.n3317 gnd.n2342 24.8557
R15362 gnd.n3316 gnd.n2330 24.8557
R15363 gnd.n3589 gnd.n3588 24.8557
R15364 gnd.n3611 gnd.n2315 24.8557
R15365 gnd.n4312 gnd.t64 24.537
R15366 gnd.n4361 gnd.t324 24.537
R15367 gnd.n5191 gnd.t294 24.537
R15368 gnd.t45 gnd.n1312 24.537
R15369 gnd.n5967 gnd.n890 23.8997
R15370 gnd.n5259 gnd.n1314 23.8997
R15371 gnd.n4428 gnd.n4427 23.855
R15372 gnd.n1770 gnd.n1769 23.855
R15373 gnd.n5784 gnd.n5783 23.855
R15374 gnd.n5007 gnd.n5006 23.855
R15375 gnd.n2965 gnd.t290 23.2624
R15376 gnd.n6075 gnd.n726 22.7121
R15377 gnd.n2666 gnd.t71 22.6251
R15378 gnd.n4072 gnd.t146 21.9878
R15379 gnd.n120 gnd.t162 21.9878
R15380 gnd.n4521 gnd.n4423 21.6691
R15381 gnd.n4584 gnd.n2025 21.6691
R15382 gnd.n4614 gnd.t1 21.6691
R15383 gnd.n4607 gnd.n1987 21.6691
R15384 gnd.n4651 gnd.n4650 21.6691
R15385 gnd.n4699 gnd.n1959 21.6691
R15386 gnd.n4699 gnd.n1961 21.6691
R15387 gnd.n4718 gnd.n1951 21.6691
R15388 gnd.n4724 gnd.n1947 21.6691
R15389 gnd.n4755 gnd.n1917 21.6691
R15390 gnd.n4778 gnd.n1891 21.6691
R15391 gnd.n4783 gnd.n1884 21.6691
R15392 gnd.n4820 gnd.n1876 21.6691
R15393 gnd.n4820 gnd.n1864 21.6691
R15394 gnd.n4825 gnd.n1857 21.6691
R15395 gnd.n4884 gnd.n1849 21.6691
R15396 gnd.t296 gnd.n1845 21.6691
R15397 gnd.n4920 gnd.n1812 21.6691
R15398 gnd.n4966 gnd.n1788 21.6691
R15399 gnd.t142 gnd.n2671 21.3504
R15400 gnd.n5782 gnd.n5781 21.0737
R15401 gnd.n5075 gnd.n5074 21.0737
R15402 gnd.t285 gnd.n2377 20.7131
R15403 gnd.n2180 gnd.n2170 20.7131
R15404 gnd.t199 gnd.n733 20.7131
R15405 gnd.n7216 gnd.t156 20.7131
R15406 gnd.n111 gnd.n104 20.7131
R15407 gnd.n5778 gnd.n1201 20.3945
R15408 gnd.n4515 gnd.n4501 20.3945
R15409 gnd.n4657 gnd.n1977 20.3945
R15410 gnd.n4848 gnd.n1867 20.3945
R15411 gnd.t286 gnd.n2412 20.0758
R15412 gnd.n4050 gnd.t176 20.0758
R15413 gnd.t297 gnd.n1805 20.0758
R15414 gnd.t150 gnd.n133 20.0758
R15415 gnd.n1184 gnd.t94 19.8005
R15416 gnd.n1184 gnd.t50 19.8005
R15417 gnd.n1183 gnd.t76 19.8005
R15418 gnd.n1183 gnd.t127 19.8005
R15419 gnd.n4997 gnd.t141 19.8005
R15420 gnd.n4997 gnd.t91 19.8005
R15421 gnd.n4996 gnd.t43 19.8005
R15422 gnd.n4996 gnd.t112 19.8005
R15423 gnd.n5902 gnd.n979 19.7572
R15424 gnd.n5586 gnd.n1381 19.7572
R15425 gnd.n1180 gnd.n1179 19.5087
R15426 gnd.n1193 gnd.n1180 19.5087
R15427 gnd.n1191 gnd.n1182 19.5087
R15428 gnd.n5001 gnd.n4995 19.5087
R15429 gnd.n3132 gnd.t275 19.4385
R15430 gnd.n4337 gnd.t317 19.4385
R15431 gnd.n5848 gnd.n1143 19.4385
R15432 gnd.n4742 gnd.t16 19.4385
R15433 gnd.n4748 gnd.t2 19.4385
R15434 gnd.n5217 gnd.t288 19.4385
R15435 gnd.n4315 gnd.n4314 19.3944
R15436 gnd.n4319 gnd.n4314 19.3944
R15437 gnd.n4319 gnd.n2102 19.3944
R15438 gnd.n4331 gnd.n2102 19.3944
R15439 gnd.n4331 gnd.n2100 19.3944
R15440 gnd.n4335 gnd.n2100 19.3944
R15441 gnd.n4335 gnd.n2088 19.3944
R15442 gnd.n4347 gnd.n2088 19.3944
R15443 gnd.n4347 gnd.n2086 19.3944
R15444 gnd.n4351 gnd.n2086 19.3944
R15445 gnd.n4351 gnd.n2074 19.3944
R15446 gnd.n4363 gnd.n2074 19.3944
R15447 gnd.n4363 gnd.n2072 19.3944
R15448 gnd.n4367 gnd.n2072 19.3944
R15449 gnd.n4367 gnd.n2060 19.3944
R15450 gnd.n4379 gnd.n2060 19.3944
R15451 gnd.n4379 gnd.n2057 19.3944
R15452 gnd.n4397 gnd.n2057 19.3944
R15453 gnd.n4397 gnd.n2058 19.3944
R15454 gnd.n4393 gnd.n2058 19.3944
R15455 gnd.n4393 gnd.n4392 19.3944
R15456 gnd.n4392 gnd.n4391 19.3944
R15457 gnd.n4391 gnd.n4386 19.3944
R15458 gnd.n4387 gnd.n4386 19.3944
R15459 gnd.n4387 gnd.n1216 19.3944
R15460 gnd.n5769 gnd.n1216 19.3944
R15461 gnd.n5769 gnd.n1217 19.3944
R15462 gnd.n5765 gnd.n1217 19.3944
R15463 gnd.n5765 gnd.n5764 19.3944
R15464 gnd.n5764 gnd.n5763 19.3944
R15465 gnd.n5763 gnd.n1223 19.3944
R15466 gnd.n5759 gnd.n1223 19.3944
R15467 gnd.n5759 gnd.n5758 19.3944
R15468 gnd.n5758 gnd.n5757 19.3944
R15469 gnd.n5757 gnd.n1228 19.3944
R15470 gnd.n5753 gnd.n1228 19.3944
R15471 gnd.n5753 gnd.n5752 19.3944
R15472 gnd.n5752 gnd.n5751 19.3944
R15473 gnd.n5751 gnd.n1233 19.3944
R15474 gnd.n5747 gnd.n1233 19.3944
R15475 gnd.n5747 gnd.n5746 19.3944
R15476 gnd.n5746 gnd.n5745 19.3944
R15477 gnd.n5745 gnd.n1238 19.3944
R15478 gnd.n5741 gnd.n1238 19.3944
R15479 gnd.n5741 gnd.n5740 19.3944
R15480 gnd.n5740 gnd.n5739 19.3944
R15481 gnd.n5739 gnd.n1243 19.3944
R15482 gnd.n5735 gnd.n1243 19.3944
R15483 gnd.n5735 gnd.n5734 19.3944
R15484 gnd.n5734 gnd.n5733 19.3944
R15485 gnd.n5733 gnd.n1248 19.3944
R15486 gnd.n5729 gnd.n1248 19.3944
R15487 gnd.n5729 gnd.n5728 19.3944
R15488 gnd.n5728 gnd.n5727 19.3944
R15489 gnd.n5727 gnd.n1253 19.3944
R15490 gnd.n5723 gnd.n1253 19.3944
R15491 gnd.n5723 gnd.n5722 19.3944
R15492 gnd.n5722 gnd.n5721 19.3944
R15493 gnd.n5721 gnd.n1258 19.3944
R15494 gnd.n5717 gnd.n1258 19.3944
R15495 gnd.n5717 gnd.n5716 19.3944
R15496 gnd.n5716 gnd.n5715 19.3944
R15497 gnd.n5715 gnd.n1263 19.3944
R15498 gnd.n5711 gnd.n1263 19.3944
R15499 gnd.n5711 gnd.n5710 19.3944
R15500 gnd.n5710 gnd.n5709 19.3944
R15501 gnd.n5709 gnd.n1268 19.3944
R15502 gnd.n5705 gnd.n1268 19.3944
R15503 gnd.n5705 gnd.n5704 19.3944
R15504 gnd.n5704 gnd.n5703 19.3944
R15505 gnd.n5703 gnd.n1273 19.3944
R15506 gnd.n5699 gnd.n1273 19.3944
R15507 gnd.n5699 gnd.n5698 19.3944
R15508 gnd.n5698 gnd.n5697 19.3944
R15509 gnd.n5697 gnd.n1278 19.3944
R15510 gnd.n5693 gnd.n1278 19.3944
R15511 gnd.n5693 gnd.n5692 19.3944
R15512 gnd.n5692 gnd.n5691 19.3944
R15513 gnd.n5691 gnd.n1283 19.3944
R15514 gnd.n5687 gnd.n1283 19.3944
R15515 gnd.n5687 gnd.n5686 19.3944
R15516 gnd.n5686 gnd.n5685 19.3944
R15517 gnd.n5685 gnd.n1288 19.3944
R15518 gnd.n5681 gnd.n1288 19.3944
R15519 gnd.n5681 gnd.n5680 19.3944
R15520 gnd.n5680 gnd.n5679 19.3944
R15521 gnd.n5679 gnd.n1293 19.3944
R15522 gnd.n5675 gnd.n1293 19.3944
R15523 gnd.n5675 gnd.n5674 19.3944
R15524 gnd.n5674 gnd.n5673 19.3944
R15525 gnd.n5673 gnd.n1298 19.3944
R15526 gnd.n5669 gnd.n1298 19.3944
R15527 gnd.n5669 gnd.n5668 19.3944
R15528 gnd.n5668 gnd.n5667 19.3944
R15529 gnd.n5667 gnd.n1303 19.3944
R15530 gnd.n5663 gnd.n1303 19.3944
R15531 gnd.n5663 gnd.n5662 19.3944
R15532 gnd.n5662 gnd.n5661 19.3944
R15533 gnd.n5661 gnd.n1308 19.3944
R15534 gnd.n5657 gnd.n1308 19.3944
R15535 gnd.n5657 gnd.n5656 19.3944
R15536 gnd.n957 gnd.n873 19.3944
R15537 gnd.n5971 gnd.n873 19.3944
R15538 gnd.n5971 gnd.n5970 19.3944
R15539 gnd.n5964 gnd.n5963 19.3944
R15540 gnd.n5963 gnd.n895 19.3944
R15541 gnd.n5959 gnd.n895 19.3944
R15542 gnd.n5959 gnd.n5958 19.3944
R15543 gnd.n5958 gnd.n5957 19.3944
R15544 gnd.n5957 gnd.n900 19.3944
R15545 gnd.n5952 gnd.n900 19.3944
R15546 gnd.n5952 gnd.n5951 19.3944
R15547 gnd.n5951 gnd.n5950 19.3944
R15548 gnd.n5950 gnd.n906 19.3944
R15549 gnd.n5943 gnd.n906 19.3944
R15550 gnd.n5943 gnd.n5942 19.3944
R15551 gnd.n5942 gnd.n918 19.3944
R15552 gnd.n5935 gnd.n918 19.3944
R15553 gnd.n5935 gnd.n5934 19.3944
R15554 gnd.n5934 gnd.n926 19.3944
R15555 gnd.n5927 gnd.n926 19.3944
R15556 gnd.n5927 gnd.n5926 19.3944
R15557 gnd.n5926 gnd.n936 19.3944
R15558 gnd.n5919 gnd.n936 19.3944
R15559 gnd.n5919 gnd.n5918 19.3944
R15560 gnd.n5918 gnd.n944 19.3944
R15561 gnd.n5911 gnd.n944 19.3944
R15562 gnd.n5911 gnd.n5910 19.3944
R15563 gnd.n5632 gnd.n1334 19.3944
R15564 gnd.n5632 gnd.n5631 19.3944
R15565 gnd.n5631 gnd.n1337 19.3944
R15566 gnd.n5624 gnd.n1337 19.3944
R15567 gnd.n5624 gnd.n5623 19.3944
R15568 gnd.n5623 gnd.n1345 19.3944
R15569 gnd.n5616 gnd.n1345 19.3944
R15570 gnd.n5616 gnd.n5615 19.3944
R15571 gnd.n5615 gnd.n1353 19.3944
R15572 gnd.n5608 gnd.n1353 19.3944
R15573 gnd.n5608 gnd.n5607 19.3944
R15574 gnd.n5607 gnd.n1361 19.3944
R15575 gnd.n5600 gnd.n1361 19.3944
R15576 gnd.n5600 gnd.n5599 19.3944
R15577 gnd.n5599 gnd.n1369 19.3944
R15578 gnd.n5592 gnd.n1369 19.3944
R15579 gnd.n2847 gnd.n2846 19.3944
R15580 gnd.n2846 gnd.n2845 19.3944
R15581 gnd.n2845 gnd.n2844 19.3944
R15582 gnd.n2844 gnd.n2842 19.3944
R15583 gnd.n2842 gnd.n2839 19.3944
R15584 gnd.n2839 gnd.n2838 19.3944
R15585 gnd.n2838 gnd.n2835 19.3944
R15586 gnd.n2835 gnd.n2834 19.3944
R15587 gnd.n2834 gnd.n2831 19.3944
R15588 gnd.n2831 gnd.n2830 19.3944
R15589 gnd.n2830 gnd.n2827 19.3944
R15590 gnd.n2827 gnd.n2826 19.3944
R15591 gnd.n2826 gnd.n2823 19.3944
R15592 gnd.n2823 gnd.n2822 19.3944
R15593 gnd.n2822 gnd.n2819 19.3944
R15594 gnd.n2819 gnd.n2818 19.3944
R15595 gnd.n2818 gnd.n2815 19.3944
R15596 gnd.n2815 gnd.n2814 19.3944
R15597 gnd.n2814 gnd.n2811 19.3944
R15598 gnd.n2811 gnd.n2810 19.3944
R15599 gnd.n2810 gnd.n2807 19.3944
R15600 gnd.n2807 gnd.n2806 19.3944
R15601 gnd.n2803 gnd.n2802 19.3944
R15602 gnd.n2802 gnd.n2758 19.3944
R15603 gnd.n2853 gnd.n2758 19.3944
R15604 gnd.n3619 gnd.n3618 19.3944
R15605 gnd.n3618 gnd.n3615 19.3944
R15606 gnd.n3615 gnd.n3614 19.3944
R15607 gnd.n3664 gnd.n3663 19.3944
R15608 gnd.n3663 gnd.n3662 19.3944
R15609 gnd.n3662 gnd.n3659 19.3944
R15610 gnd.n3659 gnd.n3658 19.3944
R15611 gnd.n3658 gnd.n3655 19.3944
R15612 gnd.n3655 gnd.n3654 19.3944
R15613 gnd.n3654 gnd.n3651 19.3944
R15614 gnd.n3651 gnd.n3650 19.3944
R15615 gnd.n3650 gnd.n3647 19.3944
R15616 gnd.n3647 gnd.n3646 19.3944
R15617 gnd.n3646 gnd.n3643 19.3944
R15618 gnd.n3643 gnd.n3642 19.3944
R15619 gnd.n3642 gnd.n3639 19.3944
R15620 gnd.n3639 gnd.n3638 19.3944
R15621 gnd.n3638 gnd.n3635 19.3944
R15622 gnd.n3635 gnd.n3634 19.3944
R15623 gnd.n3634 gnd.n3631 19.3944
R15624 gnd.n3631 gnd.n3630 19.3944
R15625 gnd.n3630 gnd.n3627 19.3944
R15626 gnd.n3627 gnd.n3626 19.3944
R15627 gnd.n3626 gnd.n3623 19.3944
R15628 gnd.n3623 gnd.n3622 19.3944
R15629 gnd.n2946 gnd.n2655 19.3944
R15630 gnd.n2956 gnd.n2655 19.3944
R15631 gnd.n2957 gnd.n2956 19.3944
R15632 gnd.n2957 gnd.n2636 19.3944
R15633 gnd.n2977 gnd.n2636 19.3944
R15634 gnd.n2977 gnd.n2628 19.3944
R15635 gnd.n2987 gnd.n2628 19.3944
R15636 gnd.n2988 gnd.n2987 19.3944
R15637 gnd.n2989 gnd.n2988 19.3944
R15638 gnd.n2989 gnd.n2611 19.3944
R15639 gnd.n3006 gnd.n2611 19.3944
R15640 gnd.n3009 gnd.n3006 19.3944
R15641 gnd.n3009 gnd.n3008 19.3944
R15642 gnd.n3008 gnd.n2584 19.3944
R15643 gnd.n3048 gnd.n2584 19.3944
R15644 gnd.n3048 gnd.n2581 19.3944
R15645 gnd.n3054 gnd.n2581 19.3944
R15646 gnd.n3055 gnd.n3054 19.3944
R15647 gnd.n3055 gnd.n2579 19.3944
R15648 gnd.n3061 gnd.n2579 19.3944
R15649 gnd.n3064 gnd.n3061 19.3944
R15650 gnd.n3066 gnd.n3064 19.3944
R15651 gnd.n3072 gnd.n3066 19.3944
R15652 gnd.n3072 gnd.n3071 19.3944
R15653 gnd.n3071 gnd.n2454 19.3944
R15654 gnd.n3138 gnd.n2454 19.3944
R15655 gnd.n3139 gnd.n3138 19.3944
R15656 gnd.n3139 gnd.n2447 19.3944
R15657 gnd.n3150 gnd.n2447 19.3944
R15658 gnd.n3151 gnd.n3150 19.3944
R15659 gnd.n3151 gnd.n2430 19.3944
R15660 gnd.n2430 gnd.n2428 19.3944
R15661 gnd.n3175 gnd.n2428 19.3944
R15662 gnd.n3176 gnd.n3175 19.3944
R15663 gnd.n3176 gnd.n2399 19.3944
R15664 gnd.n3223 gnd.n2399 19.3944
R15665 gnd.n3224 gnd.n3223 19.3944
R15666 gnd.n3224 gnd.n2392 19.3944
R15667 gnd.n3235 gnd.n2392 19.3944
R15668 gnd.n3236 gnd.n3235 19.3944
R15669 gnd.n3236 gnd.n2375 19.3944
R15670 gnd.n2375 gnd.n2373 19.3944
R15671 gnd.n3260 gnd.n2373 19.3944
R15672 gnd.n3261 gnd.n3260 19.3944
R15673 gnd.n3261 gnd.n2345 19.3944
R15674 gnd.n3312 gnd.n2345 19.3944
R15675 gnd.n3313 gnd.n3312 19.3944
R15676 gnd.n3313 gnd.n2338 19.3944
R15677 gnd.n3580 gnd.n2338 19.3944
R15678 gnd.n3581 gnd.n3580 19.3944
R15679 gnd.n3581 gnd.n2319 19.3944
R15680 gnd.n3606 gnd.n2319 19.3944
R15681 gnd.n3606 gnd.n2320 19.3944
R15682 gnd.n2937 gnd.n2936 19.3944
R15683 gnd.n2936 gnd.n2669 19.3944
R15684 gnd.n2692 gnd.n2669 19.3944
R15685 gnd.n2695 gnd.n2692 19.3944
R15686 gnd.n2695 gnd.n2688 19.3944
R15687 gnd.n2699 gnd.n2688 19.3944
R15688 gnd.n2702 gnd.n2699 19.3944
R15689 gnd.n2705 gnd.n2702 19.3944
R15690 gnd.n2705 gnd.n2686 19.3944
R15691 gnd.n2709 gnd.n2686 19.3944
R15692 gnd.n2712 gnd.n2709 19.3944
R15693 gnd.n2715 gnd.n2712 19.3944
R15694 gnd.n2715 gnd.n2684 19.3944
R15695 gnd.n2719 gnd.n2684 19.3944
R15696 gnd.n2942 gnd.n2941 19.3944
R15697 gnd.n2941 gnd.n2645 19.3944
R15698 gnd.n2967 gnd.n2645 19.3944
R15699 gnd.n2967 gnd.n2643 19.3944
R15700 gnd.n2973 gnd.n2643 19.3944
R15701 gnd.n2973 gnd.n2972 19.3944
R15702 gnd.n2972 gnd.n2617 19.3944
R15703 gnd.n2997 gnd.n2617 19.3944
R15704 gnd.n2997 gnd.n2615 19.3944
R15705 gnd.n3001 gnd.n2615 19.3944
R15706 gnd.n3001 gnd.n2595 19.3944
R15707 gnd.n3028 gnd.n2595 19.3944
R15708 gnd.n3028 gnd.n2593 19.3944
R15709 gnd.n3038 gnd.n2593 19.3944
R15710 gnd.n3038 gnd.n3037 19.3944
R15711 gnd.n3037 gnd.n3036 19.3944
R15712 gnd.n3036 gnd.n2542 19.3944
R15713 gnd.n3086 gnd.n2542 19.3944
R15714 gnd.n3086 gnd.n3085 19.3944
R15715 gnd.n3085 gnd.n3084 19.3944
R15716 gnd.n3084 gnd.n2546 19.3944
R15717 gnd.n2566 gnd.n2546 19.3944
R15718 gnd.n2566 gnd.n2464 19.3944
R15719 gnd.n3123 gnd.n2464 19.3944
R15720 gnd.n3123 gnd.n2462 19.3944
R15721 gnd.n3129 gnd.n2462 19.3944
R15722 gnd.n3129 gnd.n3128 19.3944
R15723 gnd.n3128 gnd.n2437 19.3944
R15724 gnd.n3163 gnd.n2437 19.3944
R15725 gnd.n3163 gnd.n2435 19.3944
R15726 gnd.n3169 gnd.n2435 19.3944
R15727 gnd.n3169 gnd.n3168 19.3944
R15728 gnd.n3168 gnd.n2410 19.3944
R15729 gnd.n3208 gnd.n2410 19.3944
R15730 gnd.n3208 gnd.n2408 19.3944
R15731 gnd.n3214 gnd.n2408 19.3944
R15732 gnd.n3214 gnd.n3213 19.3944
R15733 gnd.n3213 gnd.n2382 19.3944
R15734 gnd.n3248 gnd.n2382 19.3944
R15735 gnd.n3248 gnd.n2380 19.3944
R15736 gnd.n3254 gnd.n2380 19.3944
R15737 gnd.n3254 gnd.n3253 19.3944
R15738 gnd.n3253 gnd.n2355 19.3944
R15739 gnd.n3297 gnd.n2355 19.3944
R15740 gnd.n3297 gnd.n2353 19.3944
R15741 gnd.n3303 gnd.n2353 19.3944
R15742 gnd.n3303 gnd.n3302 19.3944
R15743 gnd.n3302 gnd.n2328 19.3944
R15744 gnd.n3591 gnd.n2328 19.3944
R15745 gnd.n3591 gnd.n2326 19.3944
R15746 gnd.n3599 gnd.n2326 19.3944
R15747 gnd.n3599 gnd.n3598 19.3944
R15748 gnd.n3598 gnd.n3597 19.3944
R15749 gnd.n3700 gnd.n3699 19.3944
R15750 gnd.n3699 gnd.n2267 19.3944
R15751 gnd.n3695 gnd.n2267 19.3944
R15752 gnd.n3695 gnd.n3692 19.3944
R15753 gnd.n3692 gnd.n3689 19.3944
R15754 gnd.n3689 gnd.n3688 19.3944
R15755 gnd.n3688 gnd.n3685 19.3944
R15756 gnd.n3685 gnd.n3684 19.3944
R15757 gnd.n3684 gnd.n3681 19.3944
R15758 gnd.n3681 gnd.n3680 19.3944
R15759 gnd.n3680 gnd.n3677 19.3944
R15760 gnd.n3677 gnd.n3676 19.3944
R15761 gnd.n3676 gnd.n3673 19.3944
R15762 gnd.n3673 gnd.n3672 19.3944
R15763 gnd.n2857 gnd.n2756 19.3944
R15764 gnd.n2857 gnd.n2747 19.3944
R15765 gnd.n2870 gnd.n2747 19.3944
R15766 gnd.n2870 gnd.n2745 19.3944
R15767 gnd.n2874 gnd.n2745 19.3944
R15768 gnd.n2874 gnd.n2735 19.3944
R15769 gnd.n2886 gnd.n2735 19.3944
R15770 gnd.n2886 gnd.n2733 19.3944
R15771 gnd.n2920 gnd.n2733 19.3944
R15772 gnd.n2920 gnd.n2919 19.3944
R15773 gnd.n2919 gnd.n2918 19.3944
R15774 gnd.n2918 gnd.n2917 19.3944
R15775 gnd.n2917 gnd.n2914 19.3944
R15776 gnd.n2914 gnd.n2913 19.3944
R15777 gnd.n2913 gnd.n2912 19.3944
R15778 gnd.n2912 gnd.n2910 19.3944
R15779 gnd.n2910 gnd.n2909 19.3944
R15780 gnd.n2909 gnd.n2906 19.3944
R15781 gnd.n2906 gnd.n2905 19.3944
R15782 gnd.n2905 gnd.n2904 19.3944
R15783 gnd.n2904 gnd.n2902 19.3944
R15784 gnd.n2902 gnd.n2601 19.3944
R15785 gnd.n3017 gnd.n2601 19.3944
R15786 gnd.n3017 gnd.n2599 19.3944
R15787 gnd.n3023 gnd.n2599 19.3944
R15788 gnd.n3023 gnd.n3022 19.3944
R15789 gnd.n3022 gnd.n2523 19.3944
R15790 gnd.n3097 gnd.n2523 19.3944
R15791 gnd.n3097 gnd.n2524 19.3944
R15792 gnd.n2571 gnd.n2570 19.3944
R15793 gnd.n2574 gnd.n2573 19.3944
R15794 gnd.n2561 gnd.n2560 19.3944
R15795 gnd.n3116 gnd.n2469 19.3944
R15796 gnd.n3116 gnd.n3115 19.3944
R15797 gnd.n3115 gnd.n3114 19.3944
R15798 gnd.n3114 gnd.n3112 19.3944
R15799 gnd.n3112 gnd.n3111 19.3944
R15800 gnd.n3111 gnd.n3109 19.3944
R15801 gnd.n3109 gnd.n3108 19.3944
R15802 gnd.n3108 gnd.n2418 19.3944
R15803 gnd.n3184 gnd.n2418 19.3944
R15804 gnd.n3184 gnd.n2416 19.3944
R15805 gnd.n3203 gnd.n2416 19.3944
R15806 gnd.n3203 gnd.n3202 19.3944
R15807 gnd.n3202 gnd.n3201 19.3944
R15808 gnd.n3201 gnd.n3199 19.3944
R15809 gnd.n3199 gnd.n3198 19.3944
R15810 gnd.n3198 gnd.n3196 19.3944
R15811 gnd.n3196 gnd.n3195 19.3944
R15812 gnd.n3195 gnd.n2362 19.3944
R15813 gnd.n3269 gnd.n2362 19.3944
R15814 gnd.n3269 gnd.n2360 19.3944
R15815 gnd.n3292 gnd.n2360 19.3944
R15816 gnd.n3292 gnd.n3291 19.3944
R15817 gnd.n3291 gnd.n3290 19.3944
R15818 gnd.n3290 gnd.n3287 19.3944
R15819 gnd.n3287 gnd.n3286 19.3944
R15820 gnd.n3286 gnd.n3284 19.3944
R15821 gnd.n3284 gnd.n3283 19.3944
R15822 gnd.n3283 gnd.n3281 19.3944
R15823 gnd.n3281 gnd.n2314 19.3944
R15824 gnd.n2862 gnd.n2752 19.3944
R15825 gnd.n2862 gnd.n2750 19.3944
R15826 gnd.n2866 gnd.n2750 19.3944
R15827 gnd.n2866 gnd.n2741 19.3944
R15828 gnd.n2878 gnd.n2741 19.3944
R15829 gnd.n2878 gnd.n2739 19.3944
R15830 gnd.n2882 gnd.n2739 19.3944
R15831 gnd.n2882 gnd.n2728 19.3944
R15832 gnd.n2924 gnd.n2728 19.3944
R15833 gnd.n2924 gnd.n2682 19.3944
R15834 gnd.n2930 gnd.n2682 19.3944
R15835 gnd.n2930 gnd.n2929 19.3944
R15836 gnd.n2929 gnd.n2660 19.3944
R15837 gnd.n2951 gnd.n2660 19.3944
R15838 gnd.n2951 gnd.n2653 19.3944
R15839 gnd.n2962 gnd.n2653 19.3944
R15840 gnd.n2962 gnd.n2961 19.3944
R15841 gnd.n2961 gnd.n2634 19.3944
R15842 gnd.n2982 gnd.n2634 19.3944
R15843 gnd.n2982 gnd.n2624 19.3944
R15844 gnd.n2992 gnd.n2624 19.3944
R15845 gnd.n2992 gnd.n2607 19.3944
R15846 gnd.n3013 gnd.n2607 19.3944
R15847 gnd.n3013 gnd.n3012 19.3944
R15848 gnd.n3012 gnd.n2586 19.3944
R15849 gnd.n3043 gnd.n2586 19.3944
R15850 gnd.n3043 gnd.n2531 19.3944
R15851 gnd.n3093 gnd.n2531 19.3944
R15852 gnd.n3093 gnd.n3092 19.3944
R15853 gnd.n3092 gnd.n3091 19.3944
R15854 gnd.n3091 gnd.n2535 19.3944
R15855 gnd.n2553 gnd.n2535 19.3944
R15856 gnd.n3079 gnd.n2553 19.3944
R15857 gnd.n3079 gnd.n3078 19.3944
R15858 gnd.n3078 gnd.n3077 19.3944
R15859 gnd.n3077 gnd.n2557 19.3944
R15860 gnd.n2557 gnd.n2456 19.3944
R15861 gnd.n3134 gnd.n2456 19.3944
R15862 gnd.n3134 gnd.n2449 19.3944
R15863 gnd.n3145 gnd.n2449 19.3944
R15864 gnd.n3145 gnd.n2445 19.3944
R15865 gnd.n3158 gnd.n2445 19.3944
R15866 gnd.n3158 gnd.n3157 19.3944
R15867 gnd.n3157 gnd.n2424 19.3944
R15868 gnd.n3180 gnd.n2424 19.3944
R15869 gnd.n3180 gnd.n3179 19.3944
R15870 gnd.n3179 gnd.n2401 19.3944
R15871 gnd.n3219 gnd.n2401 19.3944
R15872 gnd.n3219 gnd.n2394 19.3944
R15873 gnd.n3230 gnd.n2394 19.3944
R15874 gnd.n3230 gnd.n2390 19.3944
R15875 gnd.n3243 gnd.n2390 19.3944
R15876 gnd.n3243 gnd.n3242 19.3944
R15877 gnd.n3242 gnd.n2369 19.3944
R15878 gnd.n3265 gnd.n2369 19.3944
R15879 gnd.n3265 gnd.n3264 19.3944
R15880 gnd.n3264 gnd.n2347 19.3944
R15881 gnd.n3308 gnd.n2347 19.3944
R15882 gnd.n3308 gnd.n2340 19.3944
R15883 gnd.n3319 gnd.n2340 19.3944
R15884 gnd.n3319 gnd.n2336 19.3944
R15885 gnd.n3586 gnd.n2336 19.3944
R15886 gnd.n3586 gnd.n3585 19.3944
R15887 gnd.n3585 gnd.n2317 19.3944
R15888 gnd.n3609 gnd.n2317 19.3944
R15889 gnd.n5947 gnd.n909 19.3944
R15890 gnd.n5947 gnd.n5946 19.3944
R15891 gnd.n5946 gnd.n912 19.3944
R15892 gnd.n5939 gnd.n912 19.3944
R15893 gnd.n5939 gnd.n5938 19.3944
R15894 gnd.n5938 gnd.n922 19.3944
R15895 gnd.n5931 gnd.n922 19.3944
R15896 gnd.n5931 gnd.n5930 19.3944
R15897 gnd.n5930 gnd.n930 19.3944
R15898 gnd.n5923 gnd.n930 19.3944
R15899 gnd.n5923 gnd.n5922 19.3944
R15900 gnd.n5922 gnd.n940 19.3944
R15901 gnd.n5915 gnd.n940 19.3944
R15902 gnd.n5915 gnd.n5914 19.3944
R15903 gnd.n5914 gnd.n948 19.3944
R15904 gnd.n5907 gnd.n948 19.3944
R15905 gnd.n6664 gnd.n308 19.3944
R15906 gnd.n6670 gnd.n308 19.3944
R15907 gnd.n6670 gnd.n306 19.3944
R15908 gnd.n6674 gnd.n306 19.3944
R15909 gnd.n6674 gnd.n302 19.3944
R15910 gnd.n6680 gnd.n302 19.3944
R15911 gnd.n6680 gnd.n300 19.3944
R15912 gnd.n6684 gnd.n300 19.3944
R15913 gnd.n6684 gnd.n296 19.3944
R15914 gnd.n6690 gnd.n296 19.3944
R15915 gnd.n6690 gnd.n294 19.3944
R15916 gnd.n6694 gnd.n294 19.3944
R15917 gnd.n6694 gnd.n290 19.3944
R15918 gnd.n6700 gnd.n290 19.3944
R15919 gnd.n6700 gnd.n288 19.3944
R15920 gnd.n6704 gnd.n288 19.3944
R15921 gnd.n6704 gnd.n284 19.3944
R15922 gnd.n6710 gnd.n284 19.3944
R15923 gnd.n6710 gnd.n282 19.3944
R15924 gnd.n6714 gnd.n282 19.3944
R15925 gnd.n6714 gnd.n278 19.3944
R15926 gnd.n6720 gnd.n278 19.3944
R15927 gnd.n6720 gnd.n276 19.3944
R15928 gnd.n6724 gnd.n276 19.3944
R15929 gnd.n6724 gnd.n272 19.3944
R15930 gnd.n6730 gnd.n272 19.3944
R15931 gnd.n6730 gnd.n270 19.3944
R15932 gnd.n6734 gnd.n270 19.3944
R15933 gnd.n6734 gnd.n266 19.3944
R15934 gnd.n6740 gnd.n266 19.3944
R15935 gnd.n6740 gnd.n264 19.3944
R15936 gnd.n6744 gnd.n264 19.3944
R15937 gnd.n6744 gnd.n260 19.3944
R15938 gnd.n6750 gnd.n260 19.3944
R15939 gnd.n6750 gnd.n258 19.3944
R15940 gnd.n6754 gnd.n258 19.3944
R15941 gnd.n6754 gnd.n254 19.3944
R15942 gnd.n6760 gnd.n254 19.3944
R15943 gnd.n6760 gnd.n252 19.3944
R15944 gnd.n6764 gnd.n252 19.3944
R15945 gnd.n6764 gnd.n248 19.3944
R15946 gnd.n6770 gnd.n248 19.3944
R15947 gnd.n6770 gnd.n246 19.3944
R15948 gnd.n6774 gnd.n246 19.3944
R15949 gnd.n6774 gnd.n242 19.3944
R15950 gnd.n6780 gnd.n242 19.3944
R15951 gnd.n6780 gnd.n240 19.3944
R15952 gnd.n6784 gnd.n240 19.3944
R15953 gnd.n6784 gnd.n236 19.3944
R15954 gnd.n6790 gnd.n236 19.3944
R15955 gnd.n6790 gnd.n234 19.3944
R15956 gnd.n6794 gnd.n234 19.3944
R15957 gnd.n6794 gnd.n230 19.3944
R15958 gnd.n6800 gnd.n230 19.3944
R15959 gnd.n6800 gnd.n228 19.3944
R15960 gnd.n6804 gnd.n228 19.3944
R15961 gnd.n6804 gnd.n224 19.3944
R15962 gnd.n6810 gnd.n224 19.3944
R15963 gnd.n6810 gnd.n222 19.3944
R15964 gnd.n6814 gnd.n222 19.3944
R15965 gnd.n6814 gnd.n218 19.3944
R15966 gnd.n6820 gnd.n218 19.3944
R15967 gnd.n6820 gnd.n216 19.3944
R15968 gnd.n6824 gnd.n216 19.3944
R15969 gnd.n6824 gnd.n212 19.3944
R15970 gnd.n6830 gnd.n212 19.3944
R15971 gnd.n6830 gnd.n210 19.3944
R15972 gnd.n6834 gnd.n210 19.3944
R15973 gnd.n6834 gnd.n206 19.3944
R15974 gnd.n6840 gnd.n206 19.3944
R15975 gnd.n6840 gnd.n204 19.3944
R15976 gnd.n6844 gnd.n204 19.3944
R15977 gnd.n6844 gnd.n200 19.3944
R15978 gnd.n6850 gnd.n200 19.3944
R15979 gnd.n6850 gnd.n198 19.3944
R15980 gnd.n6854 gnd.n198 19.3944
R15981 gnd.n6854 gnd.n194 19.3944
R15982 gnd.n6860 gnd.n194 19.3944
R15983 gnd.n6860 gnd.n192 19.3944
R15984 gnd.n6864 gnd.n192 19.3944
R15985 gnd.n6864 gnd.n188 19.3944
R15986 gnd.n6871 gnd.n188 19.3944
R15987 gnd.n6871 gnd.n186 19.3944
R15988 gnd.n6875 gnd.n186 19.3944
R15989 gnd.n6243 gnd.n559 19.3944
R15990 gnd.n6249 gnd.n559 19.3944
R15991 gnd.n6249 gnd.n557 19.3944
R15992 gnd.n6253 gnd.n557 19.3944
R15993 gnd.n6253 gnd.n553 19.3944
R15994 gnd.n6259 gnd.n553 19.3944
R15995 gnd.n6259 gnd.n551 19.3944
R15996 gnd.n6263 gnd.n551 19.3944
R15997 gnd.n6263 gnd.n547 19.3944
R15998 gnd.n6269 gnd.n547 19.3944
R15999 gnd.n6269 gnd.n545 19.3944
R16000 gnd.n6273 gnd.n545 19.3944
R16001 gnd.n6273 gnd.n541 19.3944
R16002 gnd.n6279 gnd.n541 19.3944
R16003 gnd.n6279 gnd.n539 19.3944
R16004 gnd.n6283 gnd.n539 19.3944
R16005 gnd.n6283 gnd.n535 19.3944
R16006 gnd.n6289 gnd.n535 19.3944
R16007 gnd.n6289 gnd.n533 19.3944
R16008 gnd.n6293 gnd.n533 19.3944
R16009 gnd.n6293 gnd.n529 19.3944
R16010 gnd.n6299 gnd.n529 19.3944
R16011 gnd.n6299 gnd.n527 19.3944
R16012 gnd.n6303 gnd.n527 19.3944
R16013 gnd.n6303 gnd.n523 19.3944
R16014 gnd.n6309 gnd.n523 19.3944
R16015 gnd.n6309 gnd.n521 19.3944
R16016 gnd.n6313 gnd.n521 19.3944
R16017 gnd.n6313 gnd.n517 19.3944
R16018 gnd.n6319 gnd.n517 19.3944
R16019 gnd.n6319 gnd.n515 19.3944
R16020 gnd.n6323 gnd.n515 19.3944
R16021 gnd.n6323 gnd.n511 19.3944
R16022 gnd.n6329 gnd.n511 19.3944
R16023 gnd.n6329 gnd.n509 19.3944
R16024 gnd.n6333 gnd.n509 19.3944
R16025 gnd.n6333 gnd.n505 19.3944
R16026 gnd.n6339 gnd.n505 19.3944
R16027 gnd.n6339 gnd.n503 19.3944
R16028 gnd.n6343 gnd.n503 19.3944
R16029 gnd.n6343 gnd.n499 19.3944
R16030 gnd.n6349 gnd.n499 19.3944
R16031 gnd.n6349 gnd.n497 19.3944
R16032 gnd.n6353 gnd.n497 19.3944
R16033 gnd.n6353 gnd.n493 19.3944
R16034 gnd.n6359 gnd.n493 19.3944
R16035 gnd.n6359 gnd.n491 19.3944
R16036 gnd.n6363 gnd.n491 19.3944
R16037 gnd.n6363 gnd.n487 19.3944
R16038 gnd.n6369 gnd.n487 19.3944
R16039 gnd.n6369 gnd.n485 19.3944
R16040 gnd.n6373 gnd.n485 19.3944
R16041 gnd.n6373 gnd.n481 19.3944
R16042 gnd.n6379 gnd.n481 19.3944
R16043 gnd.n6379 gnd.n479 19.3944
R16044 gnd.n6383 gnd.n479 19.3944
R16045 gnd.n6383 gnd.n475 19.3944
R16046 gnd.n6389 gnd.n475 19.3944
R16047 gnd.n6389 gnd.n473 19.3944
R16048 gnd.n6393 gnd.n473 19.3944
R16049 gnd.n6393 gnd.n469 19.3944
R16050 gnd.n6399 gnd.n469 19.3944
R16051 gnd.n6399 gnd.n467 19.3944
R16052 gnd.n6403 gnd.n467 19.3944
R16053 gnd.n6403 gnd.n463 19.3944
R16054 gnd.n6409 gnd.n463 19.3944
R16055 gnd.n6409 gnd.n461 19.3944
R16056 gnd.n6413 gnd.n461 19.3944
R16057 gnd.n6413 gnd.n457 19.3944
R16058 gnd.n6419 gnd.n457 19.3944
R16059 gnd.n6419 gnd.n455 19.3944
R16060 gnd.n6423 gnd.n455 19.3944
R16061 gnd.n6423 gnd.n451 19.3944
R16062 gnd.n6429 gnd.n451 19.3944
R16063 gnd.n6429 gnd.n449 19.3944
R16064 gnd.n6433 gnd.n449 19.3944
R16065 gnd.n6433 gnd.n445 19.3944
R16066 gnd.n6439 gnd.n445 19.3944
R16067 gnd.n6439 gnd.n443 19.3944
R16068 gnd.n6443 gnd.n443 19.3944
R16069 gnd.n6443 gnd.n439 19.3944
R16070 gnd.n6449 gnd.n439 19.3944
R16071 gnd.n6449 gnd.n437 19.3944
R16072 gnd.n6453 gnd.n437 19.3944
R16073 gnd.n6453 gnd.n433 19.3944
R16074 gnd.n6459 gnd.n433 19.3944
R16075 gnd.n6459 gnd.n431 19.3944
R16076 gnd.n6463 gnd.n431 19.3944
R16077 gnd.n6463 gnd.n427 19.3944
R16078 gnd.n6469 gnd.n427 19.3944
R16079 gnd.n6469 gnd.n425 19.3944
R16080 gnd.n6473 gnd.n425 19.3944
R16081 gnd.n6473 gnd.n421 19.3944
R16082 gnd.n6479 gnd.n421 19.3944
R16083 gnd.n6479 gnd.n419 19.3944
R16084 gnd.n6483 gnd.n419 19.3944
R16085 gnd.n6483 gnd.n415 19.3944
R16086 gnd.n6489 gnd.n415 19.3944
R16087 gnd.n6489 gnd.n413 19.3944
R16088 gnd.n6493 gnd.n413 19.3944
R16089 gnd.n6493 gnd.n409 19.3944
R16090 gnd.n6499 gnd.n409 19.3944
R16091 gnd.n6499 gnd.n407 19.3944
R16092 gnd.n6503 gnd.n407 19.3944
R16093 gnd.n6503 gnd.n403 19.3944
R16094 gnd.n6509 gnd.n403 19.3944
R16095 gnd.n6509 gnd.n401 19.3944
R16096 gnd.n6513 gnd.n401 19.3944
R16097 gnd.n6513 gnd.n397 19.3944
R16098 gnd.n6519 gnd.n397 19.3944
R16099 gnd.n6519 gnd.n395 19.3944
R16100 gnd.n6523 gnd.n395 19.3944
R16101 gnd.n6523 gnd.n391 19.3944
R16102 gnd.n6529 gnd.n391 19.3944
R16103 gnd.n6529 gnd.n389 19.3944
R16104 gnd.n6533 gnd.n389 19.3944
R16105 gnd.n6533 gnd.n385 19.3944
R16106 gnd.n6539 gnd.n385 19.3944
R16107 gnd.n6539 gnd.n383 19.3944
R16108 gnd.n6543 gnd.n383 19.3944
R16109 gnd.n6543 gnd.n379 19.3944
R16110 gnd.n6549 gnd.n379 19.3944
R16111 gnd.n6549 gnd.n377 19.3944
R16112 gnd.n6553 gnd.n377 19.3944
R16113 gnd.n6553 gnd.n373 19.3944
R16114 gnd.n6559 gnd.n373 19.3944
R16115 gnd.n6559 gnd.n371 19.3944
R16116 gnd.n6563 gnd.n371 19.3944
R16117 gnd.n6563 gnd.n367 19.3944
R16118 gnd.n6569 gnd.n367 19.3944
R16119 gnd.n6569 gnd.n365 19.3944
R16120 gnd.n6573 gnd.n365 19.3944
R16121 gnd.n6573 gnd.n361 19.3944
R16122 gnd.n6579 gnd.n361 19.3944
R16123 gnd.n6579 gnd.n359 19.3944
R16124 gnd.n6583 gnd.n359 19.3944
R16125 gnd.n6583 gnd.n355 19.3944
R16126 gnd.n6589 gnd.n355 19.3944
R16127 gnd.n6589 gnd.n353 19.3944
R16128 gnd.n6593 gnd.n353 19.3944
R16129 gnd.n6593 gnd.n349 19.3944
R16130 gnd.n6599 gnd.n349 19.3944
R16131 gnd.n6599 gnd.n347 19.3944
R16132 gnd.n6603 gnd.n347 19.3944
R16133 gnd.n6603 gnd.n343 19.3944
R16134 gnd.n6609 gnd.n343 19.3944
R16135 gnd.n6609 gnd.n341 19.3944
R16136 gnd.n6613 gnd.n341 19.3944
R16137 gnd.n6613 gnd.n337 19.3944
R16138 gnd.n6619 gnd.n337 19.3944
R16139 gnd.n6619 gnd.n335 19.3944
R16140 gnd.n6623 gnd.n335 19.3944
R16141 gnd.n6623 gnd.n331 19.3944
R16142 gnd.n6629 gnd.n331 19.3944
R16143 gnd.n6629 gnd.n329 19.3944
R16144 gnd.n6633 gnd.n329 19.3944
R16145 gnd.n6633 gnd.n325 19.3944
R16146 gnd.n6639 gnd.n325 19.3944
R16147 gnd.n6639 gnd.n323 19.3944
R16148 gnd.n6643 gnd.n323 19.3944
R16149 gnd.n6643 gnd.n319 19.3944
R16150 gnd.n6649 gnd.n319 19.3944
R16151 gnd.n6649 gnd.n317 19.3944
R16152 gnd.n6654 gnd.n317 19.3944
R16153 gnd.n6654 gnd.n313 19.3944
R16154 gnd.n6660 gnd.n313 19.3944
R16155 gnd.n6661 gnd.n6660 19.3944
R16156 gnd.n5583 gnd.n5582 19.3944
R16157 gnd.n5582 gnd.n5581 19.3944
R16158 gnd.n5581 gnd.n5580 19.3944
R16159 gnd.n5580 gnd.n5578 19.3944
R16160 gnd.n5578 gnd.n5575 19.3944
R16161 gnd.n5575 gnd.n5574 19.3944
R16162 gnd.n5574 gnd.n5571 19.3944
R16163 gnd.n5571 gnd.n5570 19.3944
R16164 gnd.n5570 gnd.n5567 19.3944
R16165 gnd.n5567 gnd.n5566 19.3944
R16166 gnd.n5566 gnd.n5563 19.3944
R16167 gnd.n5563 gnd.n5562 19.3944
R16168 gnd.n5562 gnd.n5559 19.3944
R16169 gnd.n5559 gnd.n5558 19.3944
R16170 gnd.n5558 gnd.n5555 19.3944
R16171 gnd.n5555 gnd.n5554 19.3944
R16172 gnd.n5554 gnd.n5551 19.3944
R16173 gnd.n5549 gnd.n5546 19.3944
R16174 gnd.n5546 gnd.n5545 19.3944
R16175 gnd.n5545 gnd.n5542 19.3944
R16176 gnd.n5542 gnd.n5541 19.3944
R16177 gnd.n5541 gnd.n5538 19.3944
R16178 gnd.n5538 gnd.n5537 19.3944
R16179 gnd.n5537 gnd.n5534 19.3944
R16180 gnd.n5532 gnd.n5529 19.3944
R16181 gnd.n5529 gnd.n5528 19.3944
R16182 gnd.n5528 gnd.n5525 19.3944
R16183 gnd.n5525 gnd.n5524 19.3944
R16184 gnd.n5524 gnd.n5521 19.3944
R16185 gnd.n5521 gnd.n5520 19.3944
R16186 gnd.n5520 gnd.n5517 19.3944
R16187 gnd.n5517 gnd.n5516 19.3944
R16188 gnd.n5512 gnd.n5509 19.3944
R16189 gnd.n5509 gnd.n5508 19.3944
R16190 gnd.n5508 gnd.n5505 19.3944
R16191 gnd.n5505 gnd.n5504 19.3944
R16192 gnd.n5504 gnd.n5501 19.3944
R16193 gnd.n5501 gnd.n5500 19.3944
R16194 gnd.n5500 gnd.n5497 19.3944
R16195 gnd.n5497 gnd.n5496 19.3944
R16196 gnd.n5496 gnd.n5493 19.3944
R16197 gnd.n5493 gnd.n5492 19.3944
R16198 gnd.n5492 gnd.n5489 19.3944
R16199 gnd.n5489 gnd.n5488 19.3944
R16200 gnd.n5488 gnd.n5485 19.3944
R16201 gnd.n5485 gnd.n5484 19.3944
R16202 gnd.n5484 gnd.n5481 19.3944
R16203 gnd.n5481 gnd.n5480 19.3944
R16204 gnd.n5480 gnd.n5477 19.3944
R16205 gnd.n5477 gnd.n5476 19.3944
R16206 gnd.n5460 gnd.n1490 19.3944
R16207 gnd.n5460 gnd.n5459 19.3944
R16208 gnd.n5459 gnd.n1499 19.3944
R16209 gnd.n5274 gnd.n1499 19.3944
R16210 gnd.n5277 gnd.n5274 19.3944
R16211 gnd.n5278 gnd.n5277 19.3944
R16212 gnd.n5283 gnd.n5278 19.3944
R16213 gnd.n5284 gnd.n5283 19.3944
R16214 gnd.n5288 gnd.n5284 19.3944
R16215 gnd.n5288 gnd.n5287 19.3944
R16216 gnd.n5287 gnd.n5286 19.3944
R16217 gnd.n5286 gnd.n1618 19.3944
R16218 gnd.n5360 gnd.n1618 19.3944
R16219 gnd.n5361 gnd.n5360 19.3944
R16220 gnd.n5363 gnd.n5361 19.3944
R16221 gnd.n5363 gnd.n1612 19.3944
R16222 gnd.n5379 gnd.n1612 19.3944
R16223 gnd.n5380 gnd.n5379 19.3944
R16224 gnd.n5381 gnd.n5380 19.3944
R16225 gnd.n5381 gnd.n1608 19.3944
R16226 gnd.n5389 gnd.n1608 19.3944
R16227 gnd.n5391 gnd.n5389 19.3944
R16228 gnd.n5391 gnd.n5390 19.3944
R16229 gnd.n5390 gnd.n178 19.3944
R16230 gnd.n6889 gnd.n178 19.3944
R16231 gnd.n6889 gnd.n174 19.3944
R16232 gnd.n7218 gnd.n174 19.3944
R16233 gnd.n7219 gnd.n7218 19.3944
R16234 gnd.n7222 gnd.n7219 19.3944
R16235 gnd.n7223 gnd.n7222 19.3944
R16236 gnd.n7225 gnd.n7223 19.3944
R16237 gnd.n7226 gnd.n7225 19.3944
R16238 gnd.n7229 gnd.n7226 19.3944
R16239 gnd.n7230 gnd.n7229 19.3944
R16240 gnd.n7232 gnd.n7230 19.3944
R16241 gnd.n7233 gnd.n7232 19.3944
R16242 gnd.n7236 gnd.n7233 19.3944
R16243 gnd.n7237 gnd.n7236 19.3944
R16244 gnd.n7239 gnd.n7237 19.3944
R16245 gnd.n7240 gnd.n7239 19.3944
R16246 gnd.n7242 gnd.n7240 19.3944
R16247 gnd.n7243 gnd.n7242 19.3944
R16248 gnd.n5463 gnd.n5462 19.3944
R16249 gnd.n5462 gnd.n1497 19.3944
R16250 gnd.n1521 gnd.n1497 19.3944
R16251 gnd.n5449 gnd.n1521 19.3944
R16252 gnd.n5449 gnd.n5448 19.3944
R16253 gnd.n5448 gnd.n5447 19.3944
R16254 gnd.n5447 gnd.n1526 19.3944
R16255 gnd.n5437 gnd.n1526 19.3944
R16256 gnd.n5437 gnd.n5436 19.3944
R16257 gnd.n5436 gnd.n5435 19.3944
R16258 gnd.n5435 gnd.n1546 19.3944
R16259 gnd.n5425 gnd.n1546 19.3944
R16260 gnd.n5425 gnd.n5424 19.3944
R16261 gnd.n5424 gnd.n5423 19.3944
R16262 gnd.n5423 gnd.n1566 19.3944
R16263 gnd.n5413 gnd.n1566 19.3944
R16264 gnd.n5413 gnd.n5412 19.3944
R16265 gnd.n5412 gnd.n5411 19.3944
R16266 gnd.n5411 gnd.n1583 19.3944
R16267 gnd.n5384 gnd.n1583 19.3944
R16268 gnd.n5384 gnd.n1606 19.3944
R16269 gnd.n5393 gnd.n1606 19.3944
R16270 gnd.n5393 gnd.n180 19.3944
R16271 gnd.n6886 gnd.n180 19.3944
R16272 gnd.n6886 gnd.n96 19.3944
R16273 gnd.n7293 gnd.n96 19.3944
R16274 gnd.n7293 gnd.n7292 19.3944
R16275 gnd.n7292 gnd.n7291 19.3944
R16276 gnd.n7291 gnd.n100 19.3944
R16277 gnd.n7281 gnd.n100 19.3944
R16278 gnd.n7281 gnd.n7280 19.3944
R16279 gnd.n7280 gnd.n7279 19.3944
R16280 gnd.n7279 gnd.n118 19.3944
R16281 gnd.n7269 gnd.n118 19.3944
R16282 gnd.n7269 gnd.n7268 19.3944
R16283 gnd.n7268 gnd.n7267 19.3944
R16284 gnd.n7267 gnd.n138 19.3944
R16285 gnd.n7257 gnd.n138 19.3944
R16286 gnd.n7257 gnd.n7256 19.3944
R16287 gnd.n7256 gnd.n7255 19.3944
R16288 gnd.n7255 gnd.n157 19.3944
R16289 gnd.n7245 gnd.n157 19.3944
R16290 gnd.n7107 gnd.n7043 19.3944
R16291 gnd.n7107 gnd.n7104 19.3944
R16292 gnd.n7104 gnd.n7101 19.3944
R16293 gnd.n7101 gnd.n7100 19.3944
R16294 gnd.n7100 gnd.n7097 19.3944
R16295 gnd.n7097 gnd.n7096 19.3944
R16296 gnd.n7096 gnd.n7093 19.3944
R16297 gnd.n7093 gnd.n7092 19.3944
R16298 gnd.n7092 gnd.n7089 19.3944
R16299 gnd.n7089 gnd.n7088 19.3944
R16300 gnd.n7088 gnd.n7085 19.3944
R16301 gnd.n7085 gnd.n7084 19.3944
R16302 gnd.n7084 gnd.n7081 19.3944
R16303 gnd.n7081 gnd.n7080 19.3944
R16304 gnd.n7080 gnd.n7077 19.3944
R16305 gnd.n7077 gnd.n7076 19.3944
R16306 gnd.n7076 gnd.n7073 19.3944
R16307 gnd.n7073 gnd.n7072 19.3944
R16308 gnd.n7150 gnd.n7147 19.3944
R16309 gnd.n7147 gnd.n7146 19.3944
R16310 gnd.n7146 gnd.n7143 19.3944
R16311 gnd.n7143 gnd.n7142 19.3944
R16312 gnd.n7142 gnd.n7139 19.3944
R16313 gnd.n7139 gnd.n7138 19.3944
R16314 gnd.n7138 gnd.n7135 19.3944
R16315 gnd.n7135 gnd.n7134 19.3944
R16316 gnd.n7134 gnd.n7131 19.3944
R16317 gnd.n7131 gnd.n7130 19.3944
R16318 gnd.n7130 gnd.n7127 19.3944
R16319 gnd.n7127 gnd.n7126 19.3944
R16320 gnd.n7126 gnd.n7123 19.3944
R16321 gnd.n7123 gnd.n7122 19.3944
R16322 gnd.n7122 gnd.n7119 19.3944
R16323 gnd.n7119 gnd.n7118 19.3944
R16324 gnd.n7118 gnd.n7115 19.3944
R16325 gnd.n7115 gnd.n7114 19.3944
R16326 gnd.n7005 gnd.n7004 19.3944
R16327 gnd.n7183 gnd.n7004 19.3944
R16328 gnd.n7183 gnd.n7182 19.3944
R16329 gnd.n7182 gnd.n7181 19.3944
R16330 gnd.n7181 gnd.n7178 19.3944
R16331 gnd.n7178 gnd.n7177 19.3944
R16332 gnd.n7177 gnd.n7174 19.3944
R16333 gnd.n7174 gnd.n7173 19.3944
R16334 gnd.n7173 gnd.n7170 19.3944
R16335 gnd.n7170 gnd.n7169 19.3944
R16336 gnd.n7169 gnd.n7166 19.3944
R16337 gnd.n7166 gnd.n7165 19.3944
R16338 gnd.n7165 gnd.n7162 19.3944
R16339 gnd.n7162 gnd.n7161 19.3944
R16340 gnd.n7161 gnd.n7158 19.3944
R16341 gnd.n7158 gnd.n7157 19.3944
R16342 gnd.n7157 gnd.n7154 19.3944
R16343 gnd.n6935 gnd.n6933 19.3944
R16344 gnd.n6938 gnd.n6935 19.3944
R16345 gnd.n6938 gnd.n6930 19.3944
R16346 gnd.n6942 gnd.n6930 19.3944
R16347 gnd.n6945 gnd.n6942 19.3944
R16348 gnd.n6948 gnd.n6945 19.3944
R16349 gnd.n6948 gnd.n6928 19.3944
R16350 gnd.n6952 gnd.n6928 19.3944
R16351 gnd.n6955 gnd.n6952 19.3944
R16352 gnd.n6958 gnd.n6955 19.3944
R16353 gnd.n6958 gnd.n6926 19.3944
R16354 gnd.n6962 gnd.n6926 19.3944
R16355 gnd.n6965 gnd.n6962 19.3944
R16356 gnd.n6967 gnd.n6965 19.3944
R16357 gnd.n6967 gnd.n6924 19.3944
R16358 gnd.n6971 gnd.n6924 19.3944
R16359 gnd.n5305 gnd.n1637 19.3944
R16360 gnd.n5305 gnd.n1638 19.3944
R16361 gnd.n5301 gnd.n1638 19.3944
R16362 gnd.n5301 gnd.n5300 19.3944
R16363 gnd.n5300 gnd.n5299 19.3944
R16364 gnd.n5299 gnd.n5271 19.3944
R16365 gnd.n5295 gnd.n5271 19.3944
R16366 gnd.n5295 gnd.n5294 19.3944
R16367 gnd.n5294 gnd.n5293 19.3944
R16368 gnd.n5293 gnd.n1621 19.3944
R16369 gnd.n5352 gnd.n1621 19.3944
R16370 gnd.n5352 gnd.n1619 19.3944
R16371 gnd.n5356 gnd.n1619 19.3944
R16372 gnd.n5356 gnd.n1616 19.3944
R16373 gnd.n5367 gnd.n1616 19.3944
R16374 gnd.n5367 gnd.n1613 19.3944
R16375 gnd.n5375 gnd.n1613 19.3944
R16376 gnd.n5375 gnd.n1614 19.3944
R16377 gnd.n5371 gnd.n1614 19.3944
R16378 gnd.n5371 gnd.n5370 19.3944
R16379 gnd.n5370 gnd.n68 19.3944
R16380 gnd.n7306 gnd.n68 19.3944
R16381 gnd.n7306 gnd.n7305 19.3944
R16382 gnd.n7305 gnd.n71 19.3944
R16383 gnd.n6893 gnd.n71 19.3944
R16384 gnd.n6893 gnd.n175 19.3944
R16385 gnd.n7214 gnd.n175 19.3944
R16386 gnd.n7214 gnd.n7213 19.3944
R16387 gnd.n7213 gnd.n7212 19.3944
R16388 gnd.n7212 gnd.n7210 19.3944
R16389 gnd.n7210 gnd.n7209 19.3944
R16390 gnd.n7209 gnd.n7207 19.3944
R16391 gnd.n7207 gnd.n7206 19.3944
R16392 gnd.n7206 gnd.n7204 19.3944
R16393 gnd.n7204 gnd.n7203 19.3944
R16394 gnd.n7203 gnd.n7201 19.3944
R16395 gnd.n7201 gnd.n7200 19.3944
R16396 gnd.n7200 gnd.n7198 19.3944
R16397 gnd.n7198 gnd.n7197 19.3944
R16398 gnd.n7197 gnd.n7195 19.3944
R16399 gnd.n7195 gnd.n7194 19.3944
R16400 gnd.n7194 gnd.n7192 19.3944
R16401 gnd.n1507 gnd.n1506 19.3944
R16402 gnd.n5455 gnd.n1506 19.3944
R16403 gnd.n5455 gnd.n5454 19.3944
R16404 gnd.n5454 gnd.n5453 19.3944
R16405 gnd.n5453 gnd.n1513 19.3944
R16406 gnd.n5443 gnd.n1513 19.3944
R16407 gnd.n5443 gnd.n5442 19.3944
R16408 gnd.n5442 gnd.n5441 19.3944
R16409 gnd.n5441 gnd.n1536 19.3944
R16410 gnd.n5431 gnd.n1536 19.3944
R16411 gnd.n5431 gnd.n5430 19.3944
R16412 gnd.n5430 gnd.n5429 19.3944
R16413 gnd.n5429 gnd.n1557 19.3944
R16414 gnd.n5419 gnd.n1557 19.3944
R16415 gnd.n5419 gnd.n5418 19.3944
R16416 gnd.n5418 gnd.n5417 19.3944
R16417 gnd.n5407 gnd.n5406 19.3944
R16418 gnd.n1591 gnd.n1590 19.3944
R16419 gnd.n1601 gnd.n1600 19.3944
R16420 gnd.n7301 gnd.n7300 19.3944
R16421 gnd.n7297 gnd.n80 19.3944
R16422 gnd.n7297 gnd.n87 19.3944
R16423 gnd.n7287 gnd.n87 19.3944
R16424 gnd.n7287 gnd.n7286 19.3944
R16425 gnd.n7286 gnd.n7285 19.3944
R16426 gnd.n7285 gnd.n109 19.3944
R16427 gnd.n7275 gnd.n109 19.3944
R16428 gnd.n7275 gnd.n7274 19.3944
R16429 gnd.n7274 gnd.n7273 19.3944
R16430 gnd.n7273 gnd.n128 19.3944
R16431 gnd.n7263 gnd.n128 19.3944
R16432 gnd.n7263 gnd.n7262 19.3944
R16433 gnd.n7262 gnd.n7261 19.3944
R16434 gnd.n7261 gnd.n148 19.3944
R16435 gnd.n7251 gnd.n148 19.3944
R16436 gnd.n7251 gnd.n7250 19.3944
R16437 gnd.n7250 gnd.n7249 19.3944
R16438 gnd.n6069 gnd.n731 19.3944
R16439 gnd.n4119 gnd.n4118 19.3944
R16440 gnd.n4123 gnd.n4122 19.3944
R16441 gnd.n4156 gnd.n2153 19.3944
R16442 gnd.n4159 gnd.n4158 19.3944
R16443 gnd.n4163 gnd.n4162 19.3944
R16444 gnd.n4168 gnd.n4163 19.3944
R16445 gnd.n4168 gnd.n4167 19.3944
R16446 gnd.n4167 gnd.n2131 19.3944
R16447 gnd.n4222 gnd.n2131 19.3944
R16448 gnd.n4222 gnd.n2129 19.3944
R16449 gnd.n4226 gnd.n2129 19.3944
R16450 gnd.n4226 gnd.n2127 19.3944
R16451 gnd.n4230 gnd.n2127 19.3944
R16452 gnd.n4230 gnd.n2125 19.3944
R16453 gnd.n4234 gnd.n2125 19.3944
R16454 gnd.n4234 gnd.n2123 19.3944
R16455 gnd.n4238 gnd.n2123 19.3944
R16456 gnd.n4238 gnd.n2121 19.3944
R16457 gnd.n4242 gnd.n2121 19.3944
R16458 gnd.n4242 gnd.n2119 19.3944
R16459 gnd.n4246 gnd.n2119 19.3944
R16460 gnd.n4246 gnd.n2117 19.3944
R16461 gnd.n4250 gnd.n2117 19.3944
R16462 gnd.n4250 gnd.n2115 19.3944
R16463 gnd.n4255 gnd.n2115 19.3944
R16464 gnd.n4255 gnd.n2113 19.3944
R16465 gnd.n4259 gnd.n2113 19.3944
R16466 gnd.n4259 gnd.n2109 19.3944
R16467 gnd.n4323 gnd.n2109 19.3944
R16468 gnd.n4323 gnd.n2107 19.3944
R16469 gnd.n4327 gnd.n2107 19.3944
R16470 gnd.n4327 gnd.n2095 19.3944
R16471 gnd.n4339 gnd.n2095 19.3944
R16472 gnd.n4339 gnd.n2093 19.3944
R16473 gnd.n4343 gnd.n2093 19.3944
R16474 gnd.n4343 gnd.n2080 19.3944
R16475 gnd.n4355 gnd.n2080 19.3944
R16476 gnd.n4355 gnd.n2078 19.3944
R16477 gnd.n4359 gnd.n2078 19.3944
R16478 gnd.n4359 gnd.n2066 19.3944
R16479 gnd.n4371 gnd.n2066 19.3944
R16480 gnd.n4371 gnd.n2064 19.3944
R16481 gnd.n4375 gnd.n2064 19.3944
R16482 gnd.n4375 gnd.n2051 19.3944
R16483 gnd.n4401 gnd.n2051 19.3944
R16484 gnd.n4401 gnd.n2049 19.3944
R16485 gnd.n4411 gnd.n2049 19.3944
R16486 gnd.n4411 gnd.n4410 19.3944
R16487 gnd.n4410 gnd.n4409 19.3944
R16488 gnd.n4409 gnd.n1207 19.3944
R16489 gnd.n5775 gnd.n1207 19.3944
R16490 gnd.n5775 gnd.n5774 19.3944
R16491 gnd.n5774 gnd.n5773 19.3944
R16492 gnd.n5773 gnd.n1211 19.3944
R16493 gnd.n4559 gnd.n1211 19.3944
R16494 gnd.n4563 gnd.n4559 19.3944
R16495 gnd.n4563 gnd.n2021 19.3944
R16496 gnd.n4588 gnd.n2021 19.3944
R16497 gnd.n4588 gnd.n2019 19.3944
R16498 gnd.n4594 gnd.n2019 19.3944
R16499 gnd.n4594 gnd.n4593 19.3944
R16500 gnd.n4593 gnd.n1993 19.3944
R16501 gnd.n4626 gnd.n1993 19.3944
R16502 gnd.n4626 gnd.n1991 19.3944
R16503 gnd.n4636 gnd.n1991 19.3944
R16504 gnd.n4636 gnd.n4635 19.3944
R16505 gnd.n4635 gnd.n4634 19.3944
R16506 gnd.n4634 gnd.n1965 19.3944
R16507 gnd.n4697 gnd.n1965 19.3944
R16508 gnd.n4697 gnd.n4696 19.3944
R16509 gnd.n4696 gnd.n4695 19.3944
R16510 gnd.n4695 gnd.n1943 19.3944
R16511 gnd.n4727 gnd.n1943 19.3944
R16512 gnd.n4727 gnd.n1941 19.3944
R16513 gnd.n4733 gnd.n1941 19.3944
R16514 gnd.n4733 gnd.n4732 19.3944
R16515 gnd.n4732 gnd.n1915 19.3944
R16516 gnd.n4765 gnd.n1915 19.3944
R16517 gnd.n4765 gnd.n1913 19.3944
R16518 gnd.n4769 gnd.n1913 19.3944
R16519 gnd.n4769 gnd.n1889 19.3944
R16520 gnd.n4802 gnd.n1889 19.3944
R16521 gnd.n4802 gnd.n1887 19.3944
R16522 gnd.n4808 gnd.n1887 19.3944
R16523 gnd.n4808 gnd.n4807 19.3944
R16524 gnd.n4807 gnd.n1862 19.3944
R16525 gnd.n4851 gnd.n1862 19.3944
R16526 gnd.n4851 gnd.n1860 19.3944
R16527 gnd.n4857 gnd.n1860 19.3944
R16528 gnd.n4857 gnd.n4856 19.3944
R16529 gnd.n4856 gnd.n1840 19.3944
R16530 gnd.n4892 gnd.n1840 19.3944
R16531 gnd.n4892 gnd.n1838 19.3944
R16532 gnd.n4898 gnd.n1838 19.3944
R16533 gnd.n4898 gnd.n4897 19.3944
R16534 gnd.n4897 gnd.n1810 19.3944
R16535 gnd.n4932 gnd.n1810 19.3944
R16536 gnd.n4932 gnd.n1808 19.3944
R16537 gnd.n4936 gnd.n1808 19.3944
R16538 gnd.n4936 gnd.n1786 19.3944
R16539 gnd.n4975 gnd.n1786 19.3944
R16540 gnd.n4975 gnd.n1784 19.3944
R16541 gnd.n4981 gnd.n1784 19.3944
R16542 gnd.n4981 gnd.n4980 19.3944
R16543 gnd.n4980 gnd.n1730 19.3944
R16544 gnd.n5151 gnd.n1730 19.3944
R16545 gnd.n5151 gnd.n1728 19.3944
R16546 gnd.n5155 gnd.n1728 19.3944
R16547 gnd.n5155 gnd.n1719 19.3944
R16548 gnd.n5168 gnd.n1719 19.3944
R16549 gnd.n5168 gnd.n1717 19.3944
R16550 gnd.n5172 gnd.n1717 19.3944
R16551 gnd.n5172 gnd.n1707 19.3944
R16552 gnd.n5185 gnd.n1707 19.3944
R16553 gnd.n5185 gnd.n1705 19.3944
R16554 gnd.n5189 gnd.n1705 19.3944
R16555 gnd.n5189 gnd.n1695 19.3944
R16556 gnd.n5202 gnd.n1695 19.3944
R16557 gnd.n5202 gnd.n1693 19.3944
R16558 gnd.n5206 gnd.n1693 19.3944
R16559 gnd.n5206 gnd.n1683 19.3944
R16560 gnd.n5219 gnd.n1683 19.3944
R16561 gnd.n5219 gnd.n1681 19.3944
R16562 gnd.n5226 gnd.n1681 19.3944
R16563 gnd.n5226 gnd.n5225 19.3944
R16564 gnd.n5225 gnd.n1671 19.3944
R16565 gnd.n5240 gnd.n1671 19.3944
R16566 gnd.n5241 gnd.n5240 19.3944
R16567 gnd.n5241 gnd.n1669 19.3944
R16568 gnd.n5256 gnd.n1669 19.3944
R16569 gnd.n5256 gnd.n5255 19.3944
R16570 gnd.n5255 gnd.n5254 19.3944
R16571 gnd.n5254 gnd.n5247 19.3944
R16572 gnd.n5250 gnd.n5247 19.3944
R16573 gnd.n5250 gnd.n1635 19.3944
R16574 gnd.n5310 gnd.n1635 19.3944
R16575 gnd.n5310 gnd.n1633 19.3944
R16576 gnd.n5314 gnd.n1633 19.3944
R16577 gnd.n5314 gnd.n1631 19.3944
R16578 gnd.n5318 gnd.n1631 19.3944
R16579 gnd.n5318 gnd.n1629 19.3944
R16580 gnd.n5322 gnd.n1629 19.3944
R16581 gnd.n5322 gnd.n1627 19.3944
R16582 gnd.n5326 gnd.n1627 19.3944
R16583 gnd.n5326 gnd.n1625 19.3944
R16584 gnd.n5347 gnd.n1625 19.3944
R16585 gnd.n5347 gnd.n5346 19.3944
R16586 gnd.n5346 gnd.n5345 19.3944
R16587 gnd.n5345 gnd.n5332 19.3944
R16588 gnd.n5341 gnd.n5332 19.3944
R16589 gnd.n5341 gnd.n5340 19.3944
R16590 gnd.n5338 gnd.n5336 19.3944
R16591 gnd.n5401 gnd.n5400 19.3944
R16592 gnd.n5398 gnd.n1598 19.3944
R16593 gnd.n6881 gnd.n183 19.3944
R16594 gnd.n6879 gnd.n6878 19.3944
R16595 gnd.n3992 gnd.n3991 19.3944
R16596 gnd.n3991 gnd.n3783 19.3944
R16597 gnd.n3986 gnd.n3783 19.3944
R16598 gnd.n3986 gnd.n3985 19.3944
R16599 gnd.n3985 gnd.n3788 19.3944
R16600 gnd.n3980 gnd.n3788 19.3944
R16601 gnd.n3980 gnd.n3979 19.3944
R16602 gnd.n3979 gnd.n3978 19.3944
R16603 gnd.n3978 gnd.n3794 19.3944
R16604 gnd.n3972 gnd.n3794 19.3944
R16605 gnd.n3972 gnd.n3971 19.3944
R16606 gnd.n3971 gnd.n3970 19.3944
R16607 gnd.n3970 gnd.n3800 19.3944
R16608 gnd.n3964 gnd.n3800 19.3944
R16609 gnd.n3964 gnd.n3963 19.3944
R16610 gnd.n3963 gnd.n3962 19.3944
R16611 gnd.n3962 gnd.n3806 19.3944
R16612 gnd.n3956 gnd.n3955 19.3944
R16613 gnd.n3955 gnd.n3954 19.3944
R16614 gnd.n3954 gnd.n3815 19.3944
R16615 gnd.n3948 gnd.n3815 19.3944
R16616 gnd.n3948 gnd.n3947 19.3944
R16617 gnd.n3947 gnd.n3946 19.3944
R16618 gnd.n3946 gnd.n3821 19.3944
R16619 gnd.n3940 gnd.n3821 19.3944
R16620 gnd.n3940 gnd.n3939 19.3944
R16621 gnd.n3939 gnd.n3938 19.3944
R16622 gnd.n3938 gnd.n3827 19.3944
R16623 gnd.n3932 gnd.n3827 19.3944
R16624 gnd.n3932 gnd.n3931 19.3944
R16625 gnd.n3931 gnd.n3930 19.3944
R16626 gnd.n3930 gnd.n3833 19.3944
R16627 gnd.n3924 gnd.n3833 19.3944
R16628 gnd.n3924 gnd.n3923 19.3944
R16629 gnd.n3923 gnd.n3922 19.3944
R16630 gnd.n3916 gnd.n3915 19.3944
R16631 gnd.n3915 gnd.n3914 19.3944
R16632 gnd.n3914 gnd.n3847 19.3944
R16633 gnd.n3908 gnd.n3847 19.3944
R16634 gnd.n3908 gnd.n3907 19.3944
R16635 gnd.n3907 gnd.n3906 19.3944
R16636 gnd.n3906 gnd.n3853 19.3944
R16637 gnd.n3900 gnd.n3853 19.3944
R16638 gnd.n3900 gnd.n3899 19.3944
R16639 gnd.n3899 gnd.n3898 19.3944
R16640 gnd.n3898 gnd.n3859 19.3944
R16641 gnd.n3892 gnd.n3859 19.3944
R16642 gnd.n3892 gnd.n3891 19.3944
R16643 gnd.n3891 gnd.n3890 19.3944
R16644 gnd.n3890 gnd.n3865 19.3944
R16645 gnd.n3884 gnd.n3865 19.3944
R16646 gnd.n3884 gnd.n3883 19.3944
R16647 gnd.n3883 gnd.n3882 19.3944
R16648 gnd.n3728 gnd.n3727 19.3944
R16649 gnd.n3733 gnd.n3728 19.3944
R16650 gnd.n3733 gnd.n3724 19.3944
R16651 gnd.n3737 gnd.n3724 19.3944
R16652 gnd.n3737 gnd.n3722 19.3944
R16653 gnd.n3743 gnd.n3722 19.3944
R16654 gnd.n3743 gnd.n3720 19.3944
R16655 gnd.n3747 gnd.n3720 19.3944
R16656 gnd.n3747 gnd.n3718 19.3944
R16657 gnd.n3753 gnd.n3718 19.3944
R16658 gnd.n3753 gnd.n3716 19.3944
R16659 gnd.n3757 gnd.n3716 19.3944
R16660 gnd.n3757 gnd.n3714 19.3944
R16661 gnd.n3763 gnd.n3714 19.3944
R16662 gnd.n3763 gnd.n3712 19.3944
R16663 gnd.n3767 gnd.n3712 19.3944
R16664 gnd.n3778 gnd.n3706 19.3944
R16665 gnd.n3778 gnd.n3777 19.3944
R16666 gnd.n3777 gnd.n2219 19.3944
R16667 gnd.n4027 gnd.n2219 19.3944
R16668 gnd.n4027 gnd.n2217 19.3944
R16669 gnd.n4033 gnd.n2217 19.3944
R16670 gnd.n4033 gnd.n4032 19.3944
R16671 gnd.n4032 gnd.n2194 19.3944
R16672 gnd.n4062 gnd.n2194 19.3944
R16673 gnd.n4062 gnd.n2192 19.3944
R16674 gnd.n4070 gnd.n2192 19.3944
R16675 gnd.n4070 gnd.n4069 19.3944
R16676 gnd.n4069 gnd.n4068 19.3944
R16677 gnd.n4068 gnd.n2168 19.3944
R16678 gnd.n4102 gnd.n2168 19.3944
R16679 gnd.n4102 gnd.n2166 19.3944
R16680 gnd.n4106 gnd.n2166 19.3944
R16681 gnd.n4106 gnd.n2163 19.3944
R16682 gnd.n4128 gnd.n2163 19.3944
R16683 gnd.n4128 gnd.n2161 19.3944
R16684 gnd.n4132 gnd.n2161 19.3944
R16685 gnd.n4132 gnd.n2156 19.3944
R16686 gnd.n4151 gnd.n2156 19.3944
R16687 gnd.n4151 gnd.n2157 19.3944
R16688 gnd.n4147 gnd.n2157 19.3944
R16689 gnd.n4147 gnd.n2147 19.3944
R16690 gnd.n4173 gnd.n2147 19.3944
R16691 gnd.n4173 gnd.n2145 19.3944
R16692 gnd.n4177 gnd.n2145 19.3944
R16693 gnd.n4177 gnd.n2134 19.3944
R16694 gnd.n4217 gnd.n2134 19.3944
R16695 gnd.n4217 gnd.n2135 19.3944
R16696 gnd.n4213 gnd.n2135 19.3944
R16697 gnd.n4213 gnd.n4212 19.3944
R16698 gnd.n4212 gnd.n4211 19.3944
R16699 gnd.n4211 gnd.n2140 19.3944
R16700 gnd.n4207 gnd.n2140 19.3944
R16701 gnd.n4207 gnd.n4206 19.3944
R16702 gnd.n4206 gnd.n4205 19.3944
R16703 gnd.n4205 gnd.n868 19.3944
R16704 gnd.n5976 gnd.n868 19.3944
R16705 gnd.n5976 gnd.n869 19.3944
R16706 gnd.n4002 gnd.n2237 19.3944
R16707 gnd.n4003 gnd.n4002 19.3944
R16708 gnd.n4005 gnd.n4003 19.3944
R16709 gnd.n4006 gnd.n4005 19.3944
R16710 gnd.n4006 gnd.n2212 19.3944
R16711 gnd.n4037 gnd.n2212 19.3944
R16712 gnd.n4038 gnd.n4037 19.3944
R16713 gnd.n4040 gnd.n4038 19.3944
R16714 gnd.n4041 gnd.n4040 19.3944
R16715 gnd.n4041 gnd.n2187 19.3944
R16716 gnd.n4074 gnd.n2187 19.3944
R16717 gnd.n4075 gnd.n4074 19.3944
R16718 gnd.n4077 gnd.n4075 19.3944
R16719 gnd.n4078 gnd.n4077 19.3944
R16720 gnd.n4080 gnd.n4078 19.3944
R16721 gnd.n4080 gnd.n2164 19.3944
R16722 gnd.n4110 gnd.n2164 19.3944
R16723 gnd.n4111 gnd.n4110 19.3944
R16724 gnd.n4112 gnd.n4111 19.3944
R16725 gnd.n4112 gnd.n2159 19.3944
R16726 gnd.n4136 gnd.n2159 19.3944
R16727 gnd.n4137 gnd.n4136 19.3944
R16728 gnd.n4138 gnd.n4137 19.3944
R16729 gnd.n4139 gnd.n4138 19.3944
R16730 gnd.n4143 gnd.n4139 19.3944
R16731 gnd.n4143 gnd.n4142 19.3944
R16732 gnd.n4142 gnd.n4141 19.3944
R16733 gnd.n4141 gnd.n2143 19.3944
R16734 gnd.n4181 gnd.n2143 19.3944
R16735 gnd.n4182 gnd.n4181 19.3944
R16736 gnd.n4183 gnd.n4182 19.3944
R16737 gnd.n4184 gnd.n4183 19.3944
R16738 gnd.n4188 gnd.n4184 19.3944
R16739 gnd.n4189 gnd.n4188 19.3944
R16740 gnd.n4193 gnd.n4189 19.3944
R16741 gnd.n4194 gnd.n4193 19.3944
R16742 gnd.n4198 gnd.n4194 19.3944
R16743 gnd.n4199 gnd.n4198 19.3944
R16744 gnd.n4200 gnd.n4199 19.3944
R16745 gnd.n4200 gnd.n866 19.3944
R16746 gnd.n5980 gnd.n866 19.3944
R16747 gnd.n5981 gnd.n5980 19.3944
R16748 gnd.n3999 gnd.n2234 19.3944
R16749 gnd.n4013 gnd.n2234 19.3944
R16750 gnd.n4013 gnd.n4012 19.3944
R16751 gnd.n4012 gnd.n4011 19.3944
R16752 gnd.n4011 gnd.n4010 19.3944
R16753 gnd.n4010 gnd.n2209 19.3944
R16754 gnd.n4048 gnd.n2209 19.3944
R16755 gnd.n4048 gnd.n4047 19.3944
R16756 gnd.n4047 gnd.n4046 19.3944
R16757 gnd.n4046 gnd.n4045 19.3944
R16758 gnd.n4045 gnd.n2183 19.3944
R16759 gnd.n4088 gnd.n2183 19.3944
R16760 gnd.n4088 gnd.n4087 19.3944
R16761 gnd.n4087 gnd.n4086 19.3944
R16762 gnd.n4086 gnd.n4085 19.3944
R16763 gnd.n4085 gnd.n4083 19.3944
R16764 gnd.n4083 gnd.n750 19.3944
R16765 gnd.n6057 gnd.n750 19.3944
R16766 gnd.n6057 gnd.n6056 19.3944
R16767 gnd.n6056 gnd.n6055 19.3944
R16768 gnd.n6055 gnd.n754 19.3944
R16769 gnd.n6044 gnd.n754 19.3944
R16770 gnd.n6044 gnd.n6043 19.3944
R16771 gnd.n6043 gnd.n6042 19.3944
R16772 gnd.n6042 gnd.n770 19.3944
R16773 gnd.n6031 gnd.n770 19.3944
R16774 gnd.n6031 gnd.n6030 19.3944
R16775 gnd.n6030 gnd.n6029 19.3944
R16776 gnd.n6029 gnd.n788 19.3944
R16777 gnd.n6019 gnd.n788 19.3944
R16778 gnd.n6019 gnd.n6018 19.3944
R16779 gnd.n6018 gnd.n6017 19.3944
R16780 gnd.n6017 gnd.n807 19.3944
R16781 gnd.n6007 gnd.n807 19.3944
R16782 gnd.n6007 gnd.n6006 19.3944
R16783 gnd.n6006 gnd.n6005 19.3944
R16784 gnd.n6005 gnd.n828 19.3944
R16785 gnd.n5995 gnd.n828 19.3944
R16786 gnd.n5995 gnd.n5994 19.3944
R16787 gnd.n5994 gnd.n5993 19.3944
R16788 gnd.n5993 gnd.n848 19.3944
R16789 gnd.n5983 gnd.n848 19.3944
R16790 gnd.n1011 gnd.n1010 19.3944
R16791 gnd.n5899 gnd.n1010 19.3944
R16792 gnd.n5899 gnd.n5898 19.3944
R16793 gnd.n5898 gnd.n5897 19.3944
R16794 gnd.n5897 gnd.n5894 19.3944
R16795 gnd.n5894 gnd.n5893 19.3944
R16796 gnd.n5893 gnd.n5890 19.3944
R16797 gnd.n5890 gnd.n5889 19.3944
R16798 gnd.n5889 gnd.n5886 19.3944
R16799 gnd.n5886 gnd.n5885 19.3944
R16800 gnd.n5885 gnd.n5882 19.3944
R16801 gnd.n5882 gnd.n5881 19.3944
R16802 gnd.n5881 gnd.n5878 19.3944
R16803 gnd.n5878 gnd.n5877 19.3944
R16804 gnd.n5877 gnd.n5874 19.3944
R16805 gnd.n5874 gnd.n5873 19.3944
R16806 gnd.n5873 gnd.n5870 19.3944
R16807 gnd.n1113 gnd.n1049 19.3944
R16808 gnd.n1113 gnd.n1110 19.3944
R16809 gnd.n1110 gnd.n1107 19.3944
R16810 gnd.n1107 gnd.n1106 19.3944
R16811 gnd.n1106 gnd.n1103 19.3944
R16812 gnd.n1103 gnd.n1102 19.3944
R16813 gnd.n1102 gnd.n1099 19.3944
R16814 gnd.n1099 gnd.n1098 19.3944
R16815 gnd.n1098 gnd.n1095 19.3944
R16816 gnd.n1095 gnd.n1094 19.3944
R16817 gnd.n1094 gnd.n1091 19.3944
R16818 gnd.n1091 gnd.n1090 19.3944
R16819 gnd.n1090 gnd.n1087 19.3944
R16820 gnd.n1087 gnd.n1086 19.3944
R16821 gnd.n1086 gnd.n1083 19.3944
R16822 gnd.n1083 gnd.n1082 19.3944
R16823 gnd.n1082 gnd.n1079 19.3944
R16824 gnd.n1079 gnd.n1078 19.3944
R16825 gnd.n1135 gnd.n1040 19.3944
R16826 gnd.n1135 gnd.n1132 19.3944
R16827 gnd.n1132 gnd.n1129 19.3944
R16828 gnd.n1129 gnd.n1128 19.3944
R16829 gnd.n1128 gnd.n1125 19.3944
R16830 gnd.n1125 gnd.n1124 19.3944
R16831 gnd.n1124 gnd.n1121 19.3944
R16832 gnd.n1121 gnd.n1120 19.3944
R16833 gnd.n5868 gnd.n5865 19.3944
R16834 gnd.n5865 gnd.n5864 19.3944
R16835 gnd.n5864 gnd.n5861 19.3944
R16836 gnd.n5861 gnd.n5860 19.3944
R16837 gnd.n5860 gnd.n5857 19.3944
R16838 gnd.n5857 gnd.n5856 19.3944
R16839 gnd.n5856 gnd.n5853 19.3944
R16840 gnd.n3995 gnd.n2228 19.3944
R16841 gnd.n4017 gnd.n2228 19.3944
R16842 gnd.n4017 gnd.n2226 19.3944
R16843 gnd.n4023 gnd.n2226 19.3944
R16844 gnd.n4023 gnd.n4022 19.3944
R16845 gnd.n4022 gnd.n2203 19.3944
R16846 gnd.n4052 gnd.n2203 19.3944
R16847 gnd.n4052 gnd.n2201 19.3944
R16848 gnd.n4058 gnd.n2201 19.3944
R16849 gnd.n4058 gnd.n4057 19.3944
R16850 gnd.n4057 gnd.n2176 19.3944
R16851 gnd.n4092 gnd.n2176 19.3944
R16852 gnd.n4092 gnd.n2174 19.3944
R16853 gnd.n4097 gnd.n2174 19.3944
R16854 gnd.n4097 gnd.n740 19.3944
R16855 gnd.n6064 gnd.n740 19.3944
R16856 gnd.n6062 gnd.n6061 19.3944
R16857 gnd.n6051 gnd.n760 19.3944
R16858 gnd.n6049 gnd.n6048 19.3944
R16859 gnd.n6038 gnd.n777 19.3944
R16860 gnd.n6036 gnd.n6035 19.3944
R16861 gnd.n6035 gnd.n778 19.3944
R16862 gnd.n6025 gnd.n778 19.3944
R16863 gnd.n6025 gnd.n6024 19.3944
R16864 gnd.n6024 gnd.n6023 19.3944
R16865 gnd.n6023 gnd.n798 19.3944
R16866 gnd.n6013 gnd.n798 19.3944
R16867 gnd.n6013 gnd.n6012 19.3944
R16868 gnd.n6012 gnd.n6011 19.3944
R16869 gnd.n6011 gnd.n818 19.3944
R16870 gnd.n6001 gnd.n818 19.3944
R16871 gnd.n6001 gnd.n6000 19.3944
R16872 gnd.n6000 gnd.n5999 19.3944
R16873 gnd.n5999 gnd.n838 19.3944
R16874 gnd.n5989 gnd.n838 19.3944
R16875 gnd.n5989 gnd.n5988 19.3944
R16876 gnd.n5988 gnd.n5987 19.3944
R16877 gnd.n6240 gnd.n6239 19.3944
R16878 gnd.n6239 gnd.n564 19.3944
R16879 gnd.n6233 gnd.n564 19.3944
R16880 gnd.n6233 gnd.n6232 19.3944
R16881 gnd.n6232 gnd.n6231 19.3944
R16882 gnd.n6231 gnd.n572 19.3944
R16883 gnd.n6225 gnd.n572 19.3944
R16884 gnd.n6225 gnd.n6224 19.3944
R16885 gnd.n6224 gnd.n6223 19.3944
R16886 gnd.n6223 gnd.n580 19.3944
R16887 gnd.n6217 gnd.n580 19.3944
R16888 gnd.n6217 gnd.n6216 19.3944
R16889 gnd.n6216 gnd.n6215 19.3944
R16890 gnd.n6215 gnd.n588 19.3944
R16891 gnd.n6209 gnd.n588 19.3944
R16892 gnd.n6209 gnd.n6208 19.3944
R16893 gnd.n6208 gnd.n6207 19.3944
R16894 gnd.n6207 gnd.n596 19.3944
R16895 gnd.n6201 gnd.n596 19.3944
R16896 gnd.n6201 gnd.n6200 19.3944
R16897 gnd.n6200 gnd.n6199 19.3944
R16898 gnd.n6199 gnd.n604 19.3944
R16899 gnd.n6193 gnd.n604 19.3944
R16900 gnd.n6193 gnd.n6192 19.3944
R16901 gnd.n6192 gnd.n6191 19.3944
R16902 gnd.n6191 gnd.n612 19.3944
R16903 gnd.n6185 gnd.n612 19.3944
R16904 gnd.n6185 gnd.n6184 19.3944
R16905 gnd.n6184 gnd.n6183 19.3944
R16906 gnd.n6183 gnd.n620 19.3944
R16907 gnd.n6177 gnd.n620 19.3944
R16908 gnd.n6177 gnd.n6176 19.3944
R16909 gnd.n6176 gnd.n6175 19.3944
R16910 gnd.n6175 gnd.n628 19.3944
R16911 gnd.n6169 gnd.n628 19.3944
R16912 gnd.n6169 gnd.n6168 19.3944
R16913 gnd.n6168 gnd.n6167 19.3944
R16914 gnd.n6167 gnd.n636 19.3944
R16915 gnd.n6161 gnd.n636 19.3944
R16916 gnd.n6161 gnd.n6160 19.3944
R16917 gnd.n6160 gnd.n6159 19.3944
R16918 gnd.n6159 gnd.n644 19.3944
R16919 gnd.n6153 gnd.n644 19.3944
R16920 gnd.n6153 gnd.n6152 19.3944
R16921 gnd.n6152 gnd.n6151 19.3944
R16922 gnd.n6151 gnd.n652 19.3944
R16923 gnd.n6145 gnd.n652 19.3944
R16924 gnd.n6145 gnd.n6144 19.3944
R16925 gnd.n6144 gnd.n6143 19.3944
R16926 gnd.n6143 gnd.n660 19.3944
R16927 gnd.n6137 gnd.n660 19.3944
R16928 gnd.n6137 gnd.n6136 19.3944
R16929 gnd.n6136 gnd.n6135 19.3944
R16930 gnd.n6135 gnd.n668 19.3944
R16931 gnd.n6129 gnd.n668 19.3944
R16932 gnd.n6129 gnd.n6128 19.3944
R16933 gnd.n6128 gnd.n6127 19.3944
R16934 gnd.n6127 gnd.n676 19.3944
R16935 gnd.n6121 gnd.n676 19.3944
R16936 gnd.n6121 gnd.n6120 19.3944
R16937 gnd.n6120 gnd.n6119 19.3944
R16938 gnd.n6119 gnd.n684 19.3944
R16939 gnd.n6113 gnd.n684 19.3944
R16940 gnd.n6113 gnd.n6112 19.3944
R16941 gnd.n6112 gnd.n6111 19.3944
R16942 gnd.n6111 gnd.n692 19.3944
R16943 gnd.n6105 gnd.n692 19.3944
R16944 gnd.n6105 gnd.n6104 19.3944
R16945 gnd.n6104 gnd.n6103 19.3944
R16946 gnd.n6103 gnd.n700 19.3944
R16947 gnd.n6097 gnd.n700 19.3944
R16948 gnd.n6097 gnd.n6096 19.3944
R16949 gnd.n6096 gnd.n6095 19.3944
R16950 gnd.n6095 gnd.n708 19.3944
R16951 gnd.n6089 gnd.n708 19.3944
R16952 gnd.n6089 gnd.n6088 19.3944
R16953 gnd.n6088 gnd.n6087 19.3944
R16954 gnd.n6087 gnd.n716 19.3944
R16955 gnd.n6081 gnd.n716 19.3944
R16956 gnd.n6081 gnd.n6080 19.3944
R16957 gnd.n6080 gnd.n6079 19.3944
R16958 gnd.n6079 gnd.n724 19.3944
R16959 gnd.n6073 gnd.n724 19.3944
R16960 gnd.n6073 gnd.n6072 19.3944
R16961 gnd.n4310 gnd.n4262 19.3944
R16962 gnd.n4310 gnd.n4263 19.3944
R16963 gnd.n4306 gnd.n4263 19.3944
R16964 gnd.n4306 gnd.n4305 19.3944
R16965 gnd.n4305 gnd.n4304 19.3944
R16966 gnd.n4304 gnd.n4268 19.3944
R16967 gnd.n4300 gnd.n4268 19.3944
R16968 gnd.n4300 gnd.n4299 19.3944
R16969 gnd.n4299 gnd.n4298 19.3944
R16970 gnd.n4298 gnd.n4272 19.3944
R16971 gnd.n4294 gnd.n4272 19.3944
R16972 gnd.n4294 gnd.n4293 19.3944
R16973 gnd.n4293 gnd.n4292 19.3944
R16974 gnd.n4292 gnd.n4276 19.3944
R16975 gnd.n4288 gnd.n4276 19.3944
R16976 gnd.n4288 gnd.n4287 19.3944
R16977 gnd.n4287 gnd.n4286 19.3944
R16978 gnd.n4286 gnd.n4280 19.3944
R16979 gnd.n4282 gnd.n4280 19.3944
R16980 gnd.n4282 gnd.n2044 19.3944
R16981 gnd.n2044 gnd.n2042 19.3944
R16982 gnd.n4418 gnd.n2042 19.3944
R16983 gnd.n4418 gnd.n2040 19.3944
R16984 gnd.n4422 gnd.n2040 19.3944
R16985 gnd.n4523 gnd.n4422 19.3944
R16986 gnd.n4524 gnd.n4523 19.3944
R16987 gnd.n4524 gnd.n2037 19.3944
R16988 gnd.n4555 gnd.n2037 19.3944
R16989 gnd.n4555 gnd.n2038 19.3944
R16990 gnd.n4551 gnd.n2038 19.3944
R16991 gnd.n4551 gnd.n4550 19.3944
R16992 gnd.n4550 gnd.n4549 19.3944
R16993 gnd.n4549 gnd.n4529 19.3944
R16994 gnd.n4545 gnd.n4529 19.3944
R16995 gnd.n4545 gnd.n4544 19.3944
R16996 gnd.n4544 gnd.n4543 19.3944
R16997 gnd.n4543 gnd.n4534 19.3944
R16998 gnd.n4539 gnd.n4534 19.3944
R16999 gnd.n4539 gnd.n4538 19.3944
R17000 gnd.n4538 gnd.n1975 19.3944
R17001 gnd.n4660 gnd.n1975 19.3944
R17002 gnd.n4661 gnd.n4660 19.3944
R17003 gnd.n4661 gnd.n1972 19.3944
R17004 gnd.n4691 gnd.n1972 19.3944
R17005 gnd.n4691 gnd.n1973 19.3944
R17006 gnd.n4687 gnd.n1973 19.3944
R17007 gnd.n4687 gnd.n4686 19.3944
R17008 gnd.n4686 gnd.n4685 19.3944
R17009 gnd.n4685 gnd.n4666 19.3944
R17010 gnd.n4681 gnd.n4666 19.3944
R17011 gnd.n4681 gnd.n4680 19.3944
R17012 gnd.n4680 gnd.n4679 19.3944
R17013 gnd.n4679 gnd.n4671 19.3944
R17014 gnd.n4675 gnd.n4671 19.3944
R17015 gnd.n4675 gnd.n4674 19.3944
R17016 gnd.n4674 gnd.n1882 19.3944
R17017 gnd.n4812 gnd.n1882 19.3944
R17018 gnd.n4812 gnd.n1879 19.3944
R17019 gnd.n4817 gnd.n1879 19.3944
R17020 gnd.n4817 gnd.n1880 19.3944
R17021 gnd.n1880 gnd.n1855 19.3944
R17022 gnd.n4861 gnd.n1855 19.3944
R17023 gnd.n4861 gnd.n1852 19.3944
R17024 gnd.n4881 gnd.n1852 19.3944
R17025 gnd.n4881 gnd.n1853 19.3944
R17026 gnd.n4877 gnd.n1853 19.3944
R17027 gnd.n4877 gnd.n4876 19.3944
R17028 gnd.n4876 gnd.n4875 19.3944
R17029 gnd.n4875 gnd.n4868 19.3944
R17030 gnd.n4871 gnd.n4868 19.3944
R17031 gnd.n4871 gnd.n4870 19.3944
R17032 gnd.n4870 gnd.n1803 19.3944
R17033 gnd.n4941 gnd.n1803 19.3944
R17034 gnd.n4941 gnd.n1800 19.3944
R17035 gnd.n4955 gnd.n1800 19.3944
R17036 gnd.n4955 gnd.n1801 19.3944
R17037 gnd.n4951 gnd.n1801 19.3944
R17038 gnd.n4951 gnd.n4950 19.3944
R17039 gnd.n4950 gnd.n4949 19.3944
R17040 gnd.n4949 gnd.n1725 19.3944
R17041 gnd.n5159 gnd.n1725 19.3944
R17042 gnd.n5159 gnd.n1723 19.3944
R17043 gnd.n5163 gnd.n1723 19.3944
R17044 gnd.n5163 gnd.n1713 19.3944
R17045 gnd.n5176 gnd.n1713 19.3944
R17046 gnd.n5176 gnd.n1711 19.3944
R17047 gnd.n5180 gnd.n1711 19.3944
R17048 gnd.n5180 gnd.n1701 19.3944
R17049 gnd.n5193 gnd.n1701 19.3944
R17050 gnd.n5193 gnd.n1699 19.3944
R17051 gnd.n5197 gnd.n1699 19.3944
R17052 gnd.n5197 gnd.n1688 19.3944
R17053 gnd.n5210 gnd.n1688 19.3944
R17054 gnd.n5210 gnd.n1686 19.3944
R17055 gnd.n5214 gnd.n1686 19.3944
R17056 gnd.n5214 gnd.n1677 19.3944
R17057 gnd.n5230 gnd.n1677 19.3944
R17058 gnd.n5230 gnd.n1675 19.3944
R17059 gnd.n5234 gnd.n1675 19.3944
R17060 gnd.n5234 gnd.n1317 19.3944
R17061 gnd.n5652 gnd.n1317 19.3944
R17062 gnd.n5649 gnd.n5648 19.3944
R17063 gnd.n5648 gnd.n5647 19.3944
R17064 gnd.n5647 gnd.n1322 19.3944
R17065 gnd.n5643 gnd.n1322 19.3944
R17066 gnd.n5643 gnd.n5642 19.3944
R17067 gnd.n5642 gnd.n5641 19.3944
R17068 gnd.n5641 gnd.n1327 19.3944
R17069 gnd.n5636 gnd.n1327 19.3944
R17070 gnd.n5636 gnd.n5635 19.3944
R17071 gnd.n5635 gnd.n1332 19.3944
R17072 gnd.n5628 gnd.n1332 19.3944
R17073 gnd.n5628 gnd.n5627 19.3944
R17074 gnd.n5627 gnd.n1341 19.3944
R17075 gnd.n5620 gnd.n1341 19.3944
R17076 gnd.n5620 gnd.n5619 19.3944
R17077 gnd.n5619 gnd.n1349 19.3944
R17078 gnd.n5612 gnd.n1349 19.3944
R17079 gnd.n5612 gnd.n5611 19.3944
R17080 gnd.n5611 gnd.n1357 19.3944
R17081 gnd.n5604 gnd.n1357 19.3944
R17082 gnd.n5604 gnd.n5603 19.3944
R17083 gnd.n5603 gnd.n1365 19.3944
R17084 gnd.n5596 gnd.n1365 19.3944
R17085 gnd.n5596 gnd.n5595 19.3944
R17086 gnd.n1663 gnd.n1642 19.3944
R17087 gnd.n5263 gnd.n1642 19.3944
R17088 gnd.n5263 gnd.n5262 19.3944
R17089 gnd.n6067 gnd.n733 19.1199
R17090 gnd.n6066 gnd.n736 19.1199
R17091 gnd.n6059 gnd.n747 19.1199
R17092 gnd.n4126 gnd.n4125 19.1199
R17093 gnd.n6053 gnd.n758 19.1199
R17094 gnd.n4134 gnd.n763 19.1199
R17095 gnd.n4153 gnd.n772 19.1199
R17096 gnd.n6040 gnd.n775 19.1199
R17097 gnd.n4145 gnd.n780 19.1199
R17098 gnd.n6033 gnd.n783 19.1199
R17099 gnd.n4171 gnd.n4170 19.1199
R17100 gnd.n6027 gnd.n792 19.1199
R17101 gnd.n4179 gnd.n800 19.1199
R17102 gnd.n4219 gnd.n809 19.1199
R17103 gnd.n6015 gnd.n812 19.1199
R17104 gnd.n4186 gnd.n820 19.1199
R17105 gnd.n6009 gnd.n823 19.1199
R17106 gnd.n4191 gnd.n4190 19.1199
R17107 gnd.n6003 gnd.n832 19.1199
R17108 gnd.n4196 gnd.n840 19.1199
R17109 gnd.n5997 gnd.n843 19.1199
R17110 gnd.n4202 gnd.n850 19.1199
R17111 gnd.n5978 gnd.n859 19.1199
R17112 gnd.n5985 gnd.n862 19.1199
R17113 gnd.t39 gnd.n1175 19.1199
R17114 gnd.n4565 gnd.n2033 19.1199
R17115 gnd.n4938 gnd.n1806 19.1199
R17116 gnd.n5465 gnd.n1491 19.1199
R17117 gnd.n5307 gnd.n1493 19.1199
R17118 gnd.n5268 gnd.n1502 19.1199
R17119 gnd.n5451 gnd.n1515 19.1199
R17120 gnd.n5275 gnd.n1518 19.1199
R17121 gnd.n5445 gnd.n1528 19.1199
R17122 gnd.n5281 gnd.n5280 19.1199
R17123 gnd.n5439 gnd.n1538 19.1199
R17124 gnd.n5290 gnd.n1541 19.1199
R17125 gnd.n5433 gnd.n1548 19.1199
R17126 gnd.n5350 gnd.n1551 19.1199
R17127 gnd.n5358 gnd.n1561 19.1199
R17128 gnd.n5421 gnd.n1568 19.1199
R17129 gnd.n5365 gnd.n1617 19.1199
R17130 gnd.n5415 gnd.n1575 19.1199
R17131 gnd.n5377 gnd.n1578 19.1199
R17132 gnd.n5409 gnd.n1585 19.1199
R17133 gnd.n5404 gnd.n1588 19.1199
R17134 gnd.n1611 gnd.n1603 19.1199
R17135 gnd.n5396 gnd.n5395 19.1199
R17136 gnd.n7303 gnd.n73 19.1199
R17137 gnd.n6884 gnd.n75 19.1199
R17138 gnd.n7295 gnd.n90 19.1199
R17139 gnd.n7216 gnd.n93 19.1199
R17140 gnd.n3089 gnd.t280 18.8012
R17141 gnd.n3074 gnd.t268 18.8012
R17142 gnd.t166 gnd.n744 18.8012
R17143 gnd.n4502 gnd.t311 18.8012
R17144 gnd.n4959 gnd.t266 18.8012
R17145 gnd.n6883 gnd.t170 18.8012
R17146 gnd.n2933 gnd.n2932 18.4825
R17147 gnd.n5534 gnd.n5533 18.4247
R17148 gnd.n5853 gnd.n5852 18.4247
R17149 gnd.n5592 gnd.n5591 18.2308
R17150 gnd.n5907 gnd.n5906 18.2308
R17151 gnd.n6971 gnd.n6914 18.2308
R17152 gnd.n3767 gnd.n3710 18.2308
R17153 gnd.t283 gnd.n2613 18.1639
R17154 gnd.n4624 gnd.n4623 17.8452
R17155 gnd.n4736 gnd.n4735 17.8452
R17156 gnd.n4771 gnd.n1911 17.8452
R17157 gnd.n4890 gnd.n1842 17.8452
R17158 gnd.n4973 gnd.t140 17.8452
R17159 gnd.n2641 gnd.t274 17.5266
R17160 gnd.n4504 gnd.t75 17.2079
R17161 gnd.n3040 gnd.t272 16.8893
R17162 gnd.n3780 gnd.t56 16.8893
R17163 gnd.t315 gnd.n1143 16.8893
R17164 gnd.n1751 gnd.t300 16.8893
R17165 gnd.n167 gnd.t27 16.8893
R17166 gnd.n5516 gnd.n5513 16.6793
R17167 gnd.n7114 gnd.n7111 16.6793
R17168 gnd.n3922 gnd.n3841 16.6793
R17169 gnd.n1120 gnd.n1117 16.6793
R17170 gnd.n4576 gnd.t302 16.5706
R17171 gnd.n4597 gnd.n4596 16.5706
R17172 gnd.n1929 gnd.n1924 16.5706
R17173 gnd.n4763 gnd.n4761 16.5706
R17174 gnd.n1827 gnd.n1826 16.5706
R17175 gnd.t305 gnd.n4929 16.5706
R17176 gnd.n5078 gnd.t42 16.5706
R17177 gnd.n2868 gnd.t129 16.2519
R17178 gnd.n2568 gnd.t284 16.2519
R17179 gnd.n3555 gnd.n3553 15.6674
R17180 gnd.n3523 gnd.n3521 15.6674
R17181 gnd.n3491 gnd.n3489 15.6674
R17182 gnd.n3460 gnd.n3458 15.6674
R17183 gnd.n3428 gnd.n3426 15.6674
R17184 gnd.n3396 gnd.n3394 15.6674
R17185 gnd.n3364 gnd.n3362 15.6674
R17186 gnd.n3333 gnd.n3331 15.6674
R17187 gnd.n2859 gnd.t129 15.6146
R17188 gnd.t35 gnd.n2322 15.6146
R17189 gnd.t133 gnd.n2323 15.6146
R17190 gnd.n5473 gnd.n5468 15.3217
R17191 gnd.n7069 gnd.n7064 15.3217
R17192 gnd.n3876 gnd.n3873 15.3217
R17193 gnd.n1075 gnd.n1070 15.3217
R17194 gnd.n4597 gnd.n2013 15.296
R17195 gnd.n2008 gnd.n2003 15.296
R17196 gnd.n1930 gnd.n1929 15.296
R17197 gnd.n4761 gnd.n1920 15.296
R17198 gnd.n4901 gnd.n1831 15.296
R17199 gnd.n1826 gnd.n1821 15.296
R17200 gnd.n4991 gnd.n4990 15.0827
R17201 gnd.n1187 gnd.n1182 15.0481
R17202 gnd.n5001 gnd.n5000 15.0481
R17203 gnd.n3227 gnd.t276 14.9773
R17204 gnd.n4015 gnd.t56 14.9773
R17205 gnd.n5991 gnd.t60 14.9773
R17206 gnd.n4413 gnd.t315 14.9773
R17207 gnd.t126 gnd.t306 14.9773
R17208 gnd.n5157 gnd.t300 14.9773
R17209 gnd.n5457 gnd.t31 14.9773
R17210 gnd.n7253 gnd.t27 14.9773
R17211 gnd.t90 gnd.n1780 14.6587
R17212 gnd.t111 gnd.n1751 14.6587
R17213 gnd.n3305 gnd.t273 14.34
R17214 gnd.n4577 gnd.n4576 14.0214
R17215 gnd.n4623 gnd.n1997 14.0214
R17216 gnd.n4736 gnd.n1935 14.0214
R17217 gnd.n1911 gnd.n1905 14.0214
R17218 gnd.n4883 gnd.n1842 14.0214
R17219 gnd.n4929 gnd.n1816 14.0214
R17220 gnd.n3015 gnd.t9 13.7027
R17221 gnd.n4693 gnd.t20 13.7027
R17222 gnd.n4810 gnd.t320 13.7027
R17223 gnd.n2725 gnd.n2724 13.5763
R17224 gnd.n3669 gnd.n2279 13.5763
R17225 gnd.n2933 gnd.n2671 13.384
R17226 gnd.n4603 gnd.t314 13.384
R17227 gnd.n1834 gnd.t299 13.384
R17228 gnd.n1198 gnd.n1179 13.1884
R17229 gnd.n1193 gnd.n1192 13.1884
R17230 gnd.n1192 gnd.n1191 13.1884
R17231 gnd.n4994 gnd.n4989 13.1884
R17232 gnd.n4995 gnd.n4994 13.1884
R17233 gnd.n1194 gnd.n1181 13.146
R17234 gnd.n1190 gnd.n1181 13.146
R17235 gnd.n4993 gnd.n4992 13.146
R17236 gnd.n4993 gnd.n4988 13.146
R17237 gnd.n3556 gnd.n3552 12.8005
R17238 gnd.n3524 gnd.n3520 12.8005
R17239 gnd.n3492 gnd.n3488 12.8005
R17240 gnd.n3461 gnd.n3457 12.8005
R17241 gnd.n3429 gnd.n3425 12.8005
R17242 gnd.n3397 gnd.n3393 12.8005
R17243 gnd.n3365 gnd.n3361 12.8005
R17244 gnd.n3334 gnd.n3330 12.8005
R17245 gnd.n6067 gnd.n6066 12.7467
R17246 gnd.n4108 gnd.n736 12.7467
R17247 gnd.n6059 gnd.n744 12.7467
R17248 gnd.n4126 gnd.n747 12.7467
R17249 gnd.n4134 gnd.n758 12.7467
R17250 gnd.n6046 gnd.n763 12.7467
R17251 gnd.n4154 gnd.n4153 12.7467
R17252 gnd.n6040 gnd.n772 12.7467
R17253 gnd.n6033 gnd.n780 12.7467
R17254 gnd.n4171 gnd.n783 12.7467
R17255 gnd.n4179 gnd.n792 12.7467
R17256 gnd.n6021 gnd.n800 12.7467
R17257 gnd.n4220 gnd.n4219 12.7467
R17258 gnd.n6015 gnd.n809 12.7467
R17259 gnd.n6009 gnd.n820 12.7467
R17260 gnd.n4191 gnd.n823 12.7467
R17261 gnd.n4196 gnd.n832 12.7467
R17262 gnd.n5997 gnd.n840 12.7467
R17263 gnd.n4202 gnd.n843 12.7467
R17264 gnd.n5991 gnd.n850 12.7467
R17265 gnd.n5978 gnd.n867 12.7467
R17266 gnd.n5985 gnd.n859 12.7467
R17267 gnd.n4557 gnd.n2033 12.7467
R17268 gnd.n4717 gnd.n4716 12.7467
R17269 gnd.n4798 gnd.n1894 12.7467
R17270 gnd.n5465 gnd.n1493 12.7467
R17271 gnd.n5308 gnd.n5307 12.7467
R17272 gnd.n5457 gnd.n1502 12.7467
R17273 gnd.n5268 gnd.n1515 12.7467
R17274 gnd.n5451 gnd.n1518 12.7467
R17275 gnd.n5275 gnd.n1528 12.7467
R17276 gnd.n5281 gnd.n1538 12.7467
R17277 gnd.n5439 gnd.n1541 12.7467
R17278 gnd.n5433 gnd.n1551 12.7467
R17279 gnd.n5350 gnd.n5349 12.7467
R17280 gnd.n5427 gnd.n1561 12.7467
R17281 gnd.n5358 gnd.n1568 12.7467
R17282 gnd.n5365 gnd.n1575 12.7467
R17283 gnd.n5415 gnd.n1578 12.7467
R17284 gnd.n5409 gnd.n1588 12.7467
R17285 gnd.n5404 gnd.n5403 12.7467
R17286 gnd.n5386 gnd.n1611 12.7467
R17287 gnd.n5396 gnd.n1603 12.7467
R17288 gnd.n7303 gnd.n75 12.7467
R17289 gnd.n6884 gnd.n6883 12.7467
R17290 gnd.n6891 gnd.n90 12.7467
R17291 gnd.n7295 gnd.n93 12.7467
R17292 gnd.t185 gnd.n775 12.4281
R17293 gnd.t317 gnd.n2090 12.4281
R17294 gnd.n5848 gnd.n1175 12.4281
R17295 gnd.n5149 gnd.n5147 12.4281
R17296 gnd.n1691 gnd.t288 12.4281
R17297 gnd.t148 gnd.n1585 12.4281
R17298 gnd.n2724 gnd.n2719 12.4126
R17299 gnd.n3672 gnd.n3669 12.4126
R17300 gnd.n5845 gnd.n5782 12.1761
R17301 gnd.n5074 gnd.n5073 12.1761
R17302 gnd.n5902 gnd.n965 12.1094
R17303 gnd.n5586 gnd.n1423 12.1094
R17304 gnd.n3560 gnd.n3559 12.0247
R17305 gnd.n3528 gnd.n3527 12.0247
R17306 gnd.n3496 gnd.n3495 12.0247
R17307 gnd.n3465 gnd.n3464 12.0247
R17308 gnd.n3433 gnd.n3432 12.0247
R17309 gnd.n3401 gnd.n3400 12.0247
R17310 gnd.n3369 gnd.n3368 12.0247
R17311 gnd.n3338 gnd.n3337 12.0247
R17312 gnd.n4035 gnd.t176 11.7908
R17313 gnd.t201 gnd.n812 11.7908
R17314 gnd.n6003 gnd.t158 11.7908
R17315 gnd.n5445 gnd.t164 11.7908
R17316 gnd.t168 gnd.n1548 11.7908
R17317 gnd.n7265 gnd.t150 11.7908
R17318 gnd.n4492 gnd.t39 11.4721
R17319 gnd.n5778 gnd.n5777 11.4721
R17320 gnd.n5078 gnd.n1774 11.4721
R17321 gnd.n3563 gnd.n3550 11.249
R17322 gnd.n3531 gnd.n3518 11.249
R17323 gnd.n3499 gnd.n3486 11.249
R17324 gnd.n3468 gnd.n3455 11.249
R17325 gnd.n3436 gnd.n3423 11.249
R17326 gnd.n3404 gnd.n3391 11.249
R17327 gnd.n3372 gnd.n3359 11.249
R17328 gnd.n3341 gnd.n3328 11.249
R17329 gnd.n3003 gnd.t9 11.1535
R17330 gnd.n4099 gnd.n2170 11.1535
R17331 gnd.n4099 gnd.t199 11.1535
R17332 gnd.n6027 gnd.t196 11.1535
R17333 gnd.n4639 gnd.t322 11.1535
R17334 gnd.n4841 gnd.t270 11.1535
R17335 gnd.n5421 gnd.t144 11.1535
R17336 gnd.n7289 gnd.t156 11.1535
R17337 gnd.n7289 gnd.n104 11.1535
R17338 gnd.t313 gnd.n4638 10.8348
R17339 gnd.t309 gnd.n4840 10.8348
R17340 gnd.n5476 gnd.n5473 10.6672
R17341 gnd.n7072 gnd.n7069 10.6672
R17342 gnd.n3882 gnd.n3873 10.6672
R17343 gnd.n1078 gnd.n1075 10.6672
R17344 gnd.n5144 gnd.n5143 10.6151
R17345 gnd.n5143 gnd.n5140 10.6151
R17346 gnd.n5138 gnd.n5135 10.6151
R17347 gnd.n5135 gnd.n5134 10.6151
R17348 gnd.n5134 gnd.n5131 10.6151
R17349 gnd.n5131 gnd.n5130 10.6151
R17350 gnd.n5130 gnd.n5127 10.6151
R17351 gnd.n5127 gnd.n5126 10.6151
R17352 gnd.n5126 gnd.n5123 10.6151
R17353 gnd.n5123 gnd.n5122 10.6151
R17354 gnd.n5122 gnd.n5119 10.6151
R17355 gnd.n5119 gnd.n5118 10.6151
R17356 gnd.n5118 gnd.n5115 10.6151
R17357 gnd.n5115 gnd.n5114 10.6151
R17358 gnd.n5114 gnd.n5111 10.6151
R17359 gnd.n5111 gnd.n5110 10.6151
R17360 gnd.n5110 gnd.n5107 10.6151
R17361 gnd.n5107 gnd.n5106 10.6151
R17362 gnd.n5106 gnd.n5103 10.6151
R17363 gnd.n5103 gnd.n5102 10.6151
R17364 gnd.n5102 gnd.n5099 10.6151
R17365 gnd.n5099 gnd.n5098 10.6151
R17366 gnd.n5098 gnd.n5095 10.6151
R17367 gnd.n5095 gnd.n5094 10.6151
R17368 gnd.n5094 gnd.n5091 10.6151
R17369 gnd.n5091 gnd.n5090 10.6151
R17370 gnd.n5090 gnd.n5087 10.6151
R17371 gnd.n5087 gnd.n5086 10.6151
R17372 gnd.n5086 gnd.n5083 10.6151
R17373 gnd.n5083 gnd.n5082 10.6151
R17374 gnd.n4495 gnd.n4494 10.6151
R17375 gnd.n4496 gnd.n4495 10.6151
R17376 gnd.n4519 gnd.n4496 10.6151
R17377 gnd.n4519 gnd.n4518 10.6151
R17378 gnd.n4518 gnd.n4517 10.6151
R17379 gnd.n4517 gnd.n4497 10.6151
R17380 gnd.n4498 gnd.n4497 10.6151
R17381 gnd.n4498 gnd.n2031 10.6151
R17382 gnd.n4568 gnd.n2031 10.6151
R17383 gnd.n4569 gnd.n4568 10.6151
R17384 gnd.n4574 gnd.n4569 10.6151
R17385 gnd.n4574 gnd.n4573 10.6151
R17386 gnd.n4573 gnd.n4572 10.6151
R17387 gnd.n4572 gnd.n4570 10.6151
R17388 gnd.n4570 gnd.n2006 10.6151
R17389 gnd.n4605 gnd.n2006 10.6151
R17390 gnd.n4606 gnd.n4605 10.6151
R17391 gnd.n4612 gnd.n4606 10.6151
R17392 gnd.n4612 gnd.n4611 10.6151
R17393 gnd.n4611 gnd.n4610 10.6151
R17394 gnd.n4610 gnd.n4609 10.6151
R17395 gnd.n4609 gnd.n1985 10.6151
R17396 gnd.n4641 gnd.n1985 10.6151
R17397 gnd.n4642 gnd.n4641 10.6151
R17398 gnd.n4648 gnd.n4642 10.6151
R17399 gnd.n4648 gnd.n4647 10.6151
R17400 gnd.n4647 gnd.n4646 10.6151
R17401 gnd.n4646 gnd.n4644 10.6151
R17402 gnd.n4644 gnd.n4643 10.6151
R17403 gnd.n4643 gnd.n1954 10.6151
R17404 gnd.n4708 gnd.n1954 10.6151
R17405 gnd.n4709 gnd.n4708 10.6151
R17406 gnd.n4714 gnd.n4709 10.6151
R17407 gnd.n4714 gnd.n4713 10.6151
R17408 gnd.n4713 gnd.n4712 10.6151
R17409 gnd.n4712 gnd.n4710 10.6151
R17410 gnd.n4710 gnd.n1927 10.6151
R17411 gnd.n4744 gnd.n1927 10.6151
R17412 gnd.n4745 gnd.n4744 10.6151
R17413 gnd.n4753 gnd.n4745 10.6151
R17414 gnd.n4753 gnd.n4752 10.6151
R17415 gnd.n4752 gnd.n4751 10.6151
R17416 gnd.n4751 gnd.n4750 10.6151
R17417 gnd.n4750 gnd.n4747 10.6151
R17418 gnd.n4747 gnd.n4746 10.6151
R17419 gnd.n4746 gnd.n1903 10.6151
R17420 gnd.n4781 gnd.n1903 10.6151
R17421 gnd.n4782 gnd.n4781 10.6151
R17422 gnd.n4785 gnd.n4782 10.6151
R17423 gnd.n4786 gnd.n4785 10.6151
R17424 gnd.n4788 gnd.n4786 10.6151
R17425 gnd.n4788 gnd.n4787 10.6151
R17426 gnd.n4787 gnd.n1874 10.6151
R17427 gnd.n4823 gnd.n1874 10.6151
R17428 gnd.n4824 gnd.n4823 10.6151
R17429 gnd.n4827 gnd.n4824 10.6151
R17430 gnd.n4828 gnd.n4827 10.6151
R17431 gnd.n4837 gnd.n4828 10.6151
R17432 gnd.n4837 gnd.n4836 10.6151
R17433 gnd.n4836 gnd.n4835 10.6151
R17434 gnd.n4835 gnd.n4834 10.6151
R17435 gnd.n4834 gnd.n4832 10.6151
R17436 gnd.n4832 gnd.n4831 10.6151
R17437 gnd.n4831 gnd.n4829 10.6151
R17438 gnd.n4829 gnd.n1824 10.6151
R17439 gnd.n4909 gnd.n1824 10.6151
R17440 gnd.n4910 gnd.n4909 10.6151
R17441 gnd.n4918 gnd.n4910 10.6151
R17442 gnd.n4918 gnd.n4917 10.6151
R17443 gnd.n4917 gnd.n4916 10.6151
R17444 gnd.n4916 gnd.n4915 10.6151
R17445 gnd.n4915 gnd.n4911 10.6151
R17446 gnd.n4911 gnd.n1797 10.6151
R17447 gnd.n4964 gnd.n1797 10.6151
R17448 gnd.n4964 gnd.n4963 10.6151
R17449 gnd.n4963 gnd.n4962 10.6151
R17450 gnd.n4962 gnd.n4961 10.6151
R17451 gnd.n4961 gnd.n1799 10.6151
R17452 gnd.n1799 gnd.n1798 10.6151
R17453 gnd.n1798 gnd.n1773 10.6151
R17454 gnd.n1773 gnd.n1771 10.6151
R17455 gnd.n4429 gnd.n1139 10.6151
R17456 gnd.n4432 gnd.n4429 10.6151
R17457 gnd.n4437 gnd.n4434 10.6151
R17458 gnd.n4438 gnd.n4437 10.6151
R17459 gnd.n4441 gnd.n4438 10.6151
R17460 gnd.n4442 gnd.n4441 10.6151
R17461 gnd.n4445 gnd.n4442 10.6151
R17462 gnd.n4446 gnd.n4445 10.6151
R17463 gnd.n4449 gnd.n4446 10.6151
R17464 gnd.n4450 gnd.n4449 10.6151
R17465 gnd.n4453 gnd.n4450 10.6151
R17466 gnd.n4454 gnd.n4453 10.6151
R17467 gnd.n4457 gnd.n4454 10.6151
R17468 gnd.n4458 gnd.n4457 10.6151
R17469 gnd.n4461 gnd.n4458 10.6151
R17470 gnd.n4462 gnd.n4461 10.6151
R17471 gnd.n4465 gnd.n4462 10.6151
R17472 gnd.n4466 gnd.n4465 10.6151
R17473 gnd.n4469 gnd.n4466 10.6151
R17474 gnd.n4470 gnd.n4469 10.6151
R17475 gnd.n4473 gnd.n4470 10.6151
R17476 gnd.n4474 gnd.n4473 10.6151
R17477 gnd.n4477 gnd.n4474 10.6151
R17478 gnd.n4478 gnd.n4477 10.6151
R17479 gnd.n4481 gnd.n4478 10.6151
R17480 gnd.n4482 gnd.n4481 10.6151
R17481 gnd.n4485 gnd.n4482 10.6151
R17482 gnd.n4486 gnd.n4485 10.6151
R17483 gnd.n4489 gnd.n4486 10.6151
R17484 gnd.n4490 gnd.n4489 10.6151
R17485 gnd.n5845 gnd.n5844 10.6151
R17486 gnd.n5844 gnd.n5843 10.6151
R17487 gnd.n5843 gnd.n5842 10.6151
R17488 gnd.n5842 gnd.n5840 10.6151
R17489 gnd.n5840 gnd.n5837 10.6151
R17490 gnd.n5837 gnd.n5836 10.6151
R17491 gnd.n5836 gnd.n5833 10.6151
R17492 gnd.n5833 gnd.n5832 10.6151
R17493 gnd.n5832 gnd.n5829 10.6151
R17494 gnd.n5829 gnd.n5828 10.6151
R17495 gnd.n5828 gnd.n5825 10.6151
R17496 gnd.n5825 gnd.n5824 10.6151
R17497 gnd.n5824 gnd.n5821 10.6151
R17498 gnd.n5821 gnd.n5820 10.6151
R17499 gnd.n5820 gnd.n5817 10.6151
R17500 gnd.n5817 gnd.n5816 10.6151
R17501 gnd.n5816 gnd.n5813 10.6151
R17502 gnd.n5813 gnd.n5812 10.6151
R17503 gnd.n5812 gnd.n5809 10.6151
R17504 gnd.n5809 gnd.n5808 10.6151
R17505 gnd.n5808 gnd.n5805 10.6151
R17506 gnd.n5805 gnd.n5804 10.6151
R17507 gnd.n5804 gnd.n5801 10.6151
R17508 gnd.n5801 gnd.n5800 10.6151
R17509 gnd.n5800 gnd.n5797 10.6151
R17510 gnd.n5797 gnd.n5796 10.6151
R17511 gnd.n5796 gnd.n5793 10.6151
R17512 gnd.n5793 gnd.n5792 10.6151
R17513 gnd.n5789 gnd.n5788 10.6151
R17514 gnd.n5788 gnd.n1140 10.6151
R17515 gnd.n5073 gnd.n5071 10.6151
R17516 gnd.n5071 gnd.n5068 10.6151
R17517 gnd.n5068 gnd.n5067 10.6151
R17518 gnd.n5067 gnd.n5064 10.6151
R17519 gnd.n5064 gnd.n5063 10.6151
R17520 gnd.n5063 gnd.n5060 10.6151
R17521 gnd.n5060 gnd.n5059 10.6151
R17522 gnd.n5059 gnd.n5056 10.6151
R17523 gnd.n5056 gnd.n5055 10.6151
R17524 gnd.n5055 gnd.n5052 10.6151
R17525 gnd.n5052 gnd.n5051 10.6151
R17526 gnd.n5051 gnd.n5048 10.6151
R17527 gnd.n5048 gnd.n5047 10.6151
R17528 gnd.n5047 gnd.n5044 10.6151
R17529 gnd.n5044 gnd.n5043 10.6151
R17530 gnd.n5043 gnd.n5040 10.6151
R17531 gnd.n5040 gnd.n5039 10.6151
R17532 gnd.n5039 gnd.n5036 10.6151
R17533 gnd.n5036 gnd.n5035 10.6151
R17534 gnd.n5035 gnd.n5032 10.6151
R17535 gnd.n5032 gnd.n5031 10.6151
R17536 gnd.n5031 gnd.n5028 10.6151
R17537 gnd.n5028 gnd.n5027 10.6151
R17538 gnd.n5027 gnd.n5024 10.6151
R17539 gnd.n5024 gnd.n5023 10.6151
R17540 gnd.n5023 gnd.n5020 10.6151
R17541 gnd.n5020 gnd.n5019 10.6151
R17542 gnd.n5019 gnd.n5016 10.6151
R17543 gnd.n5014 gnd.n5011 10.6151
R17544 gnd.n5011 gnd.n5010 10.6151
R17545 gnd.n5781 gnd.n5780 10.6151
R17546 gnd.n5780 gnd.n1199 10.6151
R17547 gnd.n4506 gnd.n1199 10.6151
R17548 gnd.n4507 gnd.n4506 10.6151
R17549 gnd.n4513 gnd.n4507 10.6151
R17550 gnd.n4513 gnd.n4512 10.6151
R17551 gnd.n4512 gnd.n4511 10.6151
R17552 gnd.n4511 gnd.n4508 10.6151
R17553 gnd.n4508 gnd.n2027 10.6151
R17554 gnd.n4580 gnd.n2027 10.6151
R17555 gnd.n4581 gnd.n4580 10.6151
R17556 gnd.n4582 gnd.n4581 10.6151
R17557 gnd.n4582 gnd.n2011 10.6151
R17558 gnd.n4599 gnd.n2011 10.6151
R17559 gnd.n4600 gnd.n4599 10.6151
R17560 gnd.n4601 gnd.n4600 10.6151
R17561 gnd.n4601 gnd.n2000 10.6151
R17562 gnd.n4616 gnd.n2000 10.6151
R17563 gnd.n4617 gnd.n4616 10.6151
R17564 gnd.n4621 gnd.n4617 10.6151
R17565 gnd.n4621 gnd.n4620 10.6151
R17566 gnd.n4620 gnd.n4619 10.6151
R17567 gnd.n4619 gnd.n1980 10.6151
R17568 gnd.n4653 gnd.n1980 10.6151
R17569 gnd.n4654 gnd.n4653 10.6151
R17570 gnd.n4655 gnd.n4654 10.6151
R17571 gnd.n4655 gnd.n1957 10.6151
R17572 gnd.n4701 gnd.n1957 10.6151
R17573 gnd.n4702 gnd.n4701 10.6151
R17574 gnd.n4703 gnd.n4702 10.6151
R17575 gnd.n4703 gnd.n1949 10.6151
R17576 gnd.n4720 gnd.n1949 10.6151
R17577 gnd.n4721 gnd.n4720 10.6151
R17578 gnd.n4722 gnd.n4721 10.6151
R17579 gnd.n4722 gnd.n1932 10.6151
R17580 gnd.n4738 gnd.n1932 10.6151
R17581 gnd.n4739 gnd.n4738 10.6151
R17582 gnd.n4740 gnd.n4739 10.6151
R17583 gnd.n4740 gnd.n1922 10.6151
R17584 gnd.n4757 gnd.n1922 10.6151
R17585 gnd.n4758 gnd.n4757 10.6151
R17586 gnd.n4759 gnd.n4758 10.6151
R17587 gnd.n4759 gnd.n1907 10.6151
R17588 gnd.n4774 gnd.n1907 10.6151
R17589 gnd.n4775 gnd.n4774 10.6151
R17590 gnd.n4776 gnd.n4775 10.6151
R17591 gnd.n4776 gnd.n1897 10.6151
R17592 gnd.n4796 gnd.n1897 10.6151
R17593 gnd.n4796 gnd.n4795 10.6151
R17594 gnd.n4795 gnd.n4794 10.6151
R17595 gnd.n4794 gnd.n1898 10.6151
R17596 gnd.n1900 gnd.n1898 10.6151
R17597 gnd.n1900 gnd.n1899 10.6151
R17598 gnd.n1899 gnd.n1870 10.6151
R17599 gnd.n4846 gnd.n1870 10.6151
R17600 gnd.n4846 gnd.n4845 10.6151
R17601 gnd.n4845 gnd.n4844 10.6151
R17602 gnd.n4844 gnd.n1871 10.6151
R17603 gnd.n1871 gnd.n1847 10.6151
R17604 gnd.n4886 gnd.n1847 10.6151
R17605 gnd.n4887 gnd.n4886 10.6151
R17606 gnd.n4888 gnd.n4887 10.6151
R17607 gnd.n4888 gnd.n1829 10.6151
R17608 gnd.n4903 gnd.n1829 10.6151
R17609 gnd.n4904 gnd.n4903 10.6151
R17610 gnd.n4905 gnd.n4904 10.6151
R17611 gnd.n4905 gnd.n1819 10.6151
R17612 gnd.n4922 gnd.n1819 10.6151
R17613 gnd.n4923 gnd.n4922 10.6151
R17614 gnd.n4927 gnd.n4923 10.6151
R17615 gnd.n4927 gnd.n4926 10.6151
R17616 gnd.n4926 gnd.n4925 10.6151
R17617 gnd.n4925 gnd.n1792 10.6151
R17618 gnd.n4968 gnd.n1792 10.6151
R17619 gnd.n4969 gnd.n4968 10.6151
R17620 gnd.n4970 gnd.n4969 10.6151
R17621 gnd.n4970 gnd.n1777 10.6151
R17622 gnd.n4985 gnd.n1777 10.6151
R17623 gnd.n4986 gnd.n4985 10.6151
R17624 gnd.n5076 gnd.n4986 10.6151
R17625 gnd.n5076 gnd.n5075 10.6151
R17626 gnd.n2922 gnd.t142 10.5161
R17627 gnd.n2367 gnd.t5 10.5161
R17628 gnd.n3288 gnd.t273 10.5161
R17629 gnd.n6053 gnd.t154 10.5161
R17630 gnd.n6046 gnd.t160 10.5161
R17631 gnd.n2009 gnd.t14 10.5161
R17632 gnd.t18 gnd.n4900 10.5161
R17633 gnd.n5386 gnd.t190 10.5161
R17634 gnd.n5395 gnd.t188 10.5161
R17635 gnd.n3564 gnd.n3548 10.4732
R17636 gnd.n3532 gnd.n3516 10.4732
R17637 gnd.n3500 gnd.n3484 10.4732
R17638 gnd.n3469 gnd.n3453 10.4732
R17639 gnd.n3437 gnd.n3421 10.4732
R17640 gnd.n3405 gnd.n3389 10.4732
R17641 gnd.n3373 gnd.n3357 10.4732
R17642 gnd.n3342 gnd.n3326 10.4732
R17643 gnd.n5771 gnd.t23 10.1975
R17644 gnd.n4658 gnd.n1959 10.1975
R17645 gnd.n1970 gnd.n1961 10.1975
R17646 gnd.n4716 gnd.t304 10.1975
R17647 gnd.t310 gnd.n4798 10.1975
R17648 gnd.n4790 gnd.n1876 10.1975
R17649 gnd.n4849 gnd.n1864 10.1975
R17650 gnd.n4958 gnd.t52 10.1975
R17651 gnd.n4959 gnd.n4958 10.1975
R17652 gnd.n1780 gnd.n1774 10.1975
R17653 gnd.t276 gnd.n2384 9.87883
R17654 gnd.n4090 gnd.t146 9.87883
R17655 gnd.n6021 gnd.t211 9.87883
R17656 gnd.n5427 gnd.t174 9.87883
R17657 gnd.n7283 gnd.t162 9.87883
R17658 gnd.n3568 gnd.n3567 9.69747
R17659 gnd.n3536 gnd.n3535 9.69747
R17660 gnd.n3504 gnd.n3503 9.69747
R17661 gnd.n3473 gnd.n3472 9.69747
R17662 gnd.n3441 gnd.n3440 9.69747
R17663 gnd.n3409 gnd.n3408 9.69747
R17664 gnd.n3377 gnd.n3376 9.69747
R17665 gnd.n3346 gnd.n3345 9.69747
R17666 gnd.n1806 gnd.t78 9.56018
R17667 gnd.n3574 gnd.n3573 9.45567
R17668 gnd.n3542 gnd.n3541 9.45567
R17669 gnd.n3510 gnd.n3509 9.45567
R17670 gnd.n3479 gnd.n3478 9.45567
R17671 gnd.n3447 gnd.n3446 9.45567
R17672 gnd.n3415 gnd.n3414 9.45567
R17673 gnd.n3383 gnd.n3382 9.45567
R17674 gnd.n3352 gnd.n3351 9.45567
R17675 gnd.n5513 gnd.n5512 9.30959
R17676 gnd.n7111 gnd.n7043 9.30959
R17677 gnd.n3916 gnd.n3841 9.30959
R17678 gnd.n1117 gnd.n1049 9.30959
R17679 gnd.n3573 gnd.n3572 9.3005
R17680 gnd.n3546 gnd.n3545 9.3005
R17681 gnd.n3567 gnd.n3566 9.3005
R17682 gnd.n3565 gnd.n3564 9.3005
R17683 gnd.n3550 gnd.n3549 9.3005
R17684 gnd.n3559 gnd.n3558 9.3005
R17685 gnd.n3557 gnd.n3556 9.3005
R17686 gnd.n3541 gnd.n3540 9.3005
R17687 gnd.n3514 gnd.n3513 9.3005
R17688 gnd.n3535 gnd.n3534 9.3005
R17689 gnd.n3533 gnd.n3532 9.3005
R17690 gnd.n3518 gnd.n3517 9.3005
R17691 gnd.n3527 gnd.n3526 9.3005
R17692 gnd.n3525 gnd.n3524 9.3005
R17693 gnd.n3509 gnd.n3508 9.3005
R17694 gnd.n3482 gnd.n3481 9.3005
R17695 gnd.n3503 gnd.n3502 9.3005
R17696 gnd.n3501 gnd.n3500 9.3005
R17697 gnd.n3486 gnd.n3485 9.3005
R17698 gnd.n3495 gnd.n3494 9.3005
R17699 gnd.n3493 gnd.n3492 9.3005
R17700 gnd.n3478 gnd.n3477 9.3005
R17701 gnd.n3451 gnd.n3450 9.3005
R17702 gnd.n3472 gnd.n3471 9.3005
R17703 gnd.n3470 gnd.n3469 9.3005
R17704 gnd.n3455 gnd.n3454 9.3005
R17705 gnd.n3464 gnd.n3463 9.3005
R17706 gnd.n3462 gnd.n3461 9.3005
R17707 gnd.n3446 gnd.n3445 9.3005
R17708 gnd.n3419 gnd.n3418 9.3005
R17709 gnd.n3440 gnd.n3439 9.3005
R17710 gnd.n3438 gnd.n3437 9.3005
R17711 gnd.n3423 gnd.n3422 9.3005
R17712 gnd.n3432 gnd.n3431 9.3005
R17713 gnd.n3430 gnd.n3429 9.3005
R17714 gnd.n3414 gnd.n3413 9.3005
R17715 gnd.n3387 gnd.n3386 9.3005
R17716 gnd.n3408 gnd.n3407 9.3005
R17717 gnd.n3406 gnd.n3405 9.3005
R17718 gnd.n3391 gnd.n3390 9.3005
R17719 gnd.n3400 gnd.n3399 9.3005
R17720 gnd.n3398 gnd.n3397 9.3005
R17721 gnd.n3382 gnd.n3381 9.3005
R17722 gnd.n3355 gnd.n3354 9.3005
R17723 gnd.n3376 gnd.n3375 9.3005
R17724 gnd.n3374 gnd.n3373 9.3005
R17725 gnd.n3359 gnd.n3358 9.3005
R17726 gnd.n3368 gnd.n3367 9.3005
R17727 gnd.n3366 gnd.n3365 9.3005
R17728 gnd.n3351 gnd.n3350 9.3005
R17729 gnd.n3324 gnd.n3323 9.3005
R17730 gnd.n3345 gnd.n3344 9.3005
R17731 gnd.n3343 gnd.n3342 9.3005
R17732 gnd.n3328 gnd.n3327 9.3005
R17733 gnd.n3337 gnd.n3336 9.3005
R17734 gnd.n3335 gnd.n3334 9.3005
R17735 gnd.n3699 gnd.n3698 9.3005
R17736 gnd.n3697 gnd.n2267 9.3005
R17737 gnd.n3696 gnd.n3695 9.3005
R17738 gnd.n3692 gnd.n2268 9.3005
R17739 gnd.n3689 gnd.n2269 9.3005
R17740 gnd.n3688 gnd.n2270 9.3005
R17741 gnd.n3685 gnd.n2271 9.3005
R17742 gnd.n3684 gnd.n2272 9.3005
R17743 gnd.n3681 gnd.n2273 9.3005
R17744 gnd.n3680 gnd.n2274 9.3005
R17745 gnd.n3677 gnd.n2275 9.3005
R17746 gnd.n3676 gnd.n2276 9.3005
R17747 gnd.n3673 gnd.n2277 9.3005
R17748 gnd.n3672 gnd.n2278 9.3005
R17749 gnd.n3669 gnd.n3668 9.3005
R17750 gnd.n3667 gnd.n2279 9.3005
R17751 gnd.n3700 gnd.n2266 9.3005
R17752 gnd.n2941 gnd.n2940 9.3005
R17753 gnd.n2645 gnd.n2644 9.3005
R17754 gnd.n2968 gnd.n2967 9.3005
R17755 gnd.n2969 gnd.n2643 9.3005
R17756 gnd.n2973 gnd.n2970 9.3005
R17757 gnd.n2972 gnd.n2971 9.3005
R17758 gnd.n2617 gnd.n2616 9.3005
R17759 gnd.n2998 gnd.n2997 9.3005
R17760 gnd.n2999 gnd.n2615 9.3005
R17761 gnd.n3001 gnd.n3000 9.3005
R17762 gnd.n2595 gnd.n2594 9.3005
R17763 gnd.n3029 gnd.n3028 9.3005
R17764 gnd.n3030 gnd.n2593 9.3005
R17765 gnd.n3038 gnd.n3031 9.3005
R17766 gnd.n3037 gnd.n3032 9.3005
R17767 gnd.n3036 gnd.n3034 9.3005
R17768 gnd.n3033 gnd.n2542 9.3005
R17769 gnd.n3086 gnd.n2543 9.3005
R17770 gnd.n3085 gnd.n2544 9.3005
R17771 gnd.n3084 gnd.n2545 9.3005
R17772 gnd.n2564 gnd.n2546 9.3005
R17773 gnd.n2566 gnd.n2565 9.3005
R17774 gnd.n2464 gnd.n2463 9.3005
R17775 gnd.n3124 gnd.n3123 9.3005
R17776 gnd.n3125 gnd.n2462 9.3005
R17777 gnd.n3129 gnd.n3126 9.3005
R17778 gnd.n3128 gnd.n3127 9.3005
R17779 gnd.n2437 gnd.n2436 9.3005
R17780 gnd.n3164 gnd.n3163 9.3005
R17781 gnd.n3165 gnd.n2435 9.3005
R17782 gnd.n3169 gnd.n3166 9.3005
R17783 gnd.n3168 gnd.n3167 9.3005
R17784 gnd.n2410 gnd.n2409 9.3005
R17785 gnd.n3209 gnd.n3208 9.3005
R17786 gnd.n3210 gnd.n2408 9.3005
R17787 gnd.n3214 gnd.n3211 9.3005
R17788 gnd.n3213 gnd.n3212 9.3005
R17789 gnd.n2382 gnd.n2381 9.3005
R17790 gnd.n3249 gnd.n3248 9.3005
R17791 gnd.n3250 gnd.n2380 9.3005
R17792 gnd.n3254 gnd.n3251 9.3005
R17793 gnd.n3253 gnd.n3252 9.3005
R17794 gnd.n2355 gnd.n2354 9.3005
R17795 gnd.n3298 gnd.n3297 9.3005
R17796 gnd.n3299 gnd.n2353 9.3005
R17797 gnd.n3303 gnd.n3300 9.3005
R17798 gnd.n3302 gnd.n3301 9.3005
R17799 gnd.n2328 gnd.n2327 9.3005
R17800 gnd.n3592 gnd.n3591 9.3005
R17801 gnd.n3593 gnd.n2326 9.3005
R17802 gnd.n3599 gnd.n3594 9.3005
R17803 gnd.n3598 gnd.n3595 9.3005
R17804 gnd.n3597 gnd.n3596 9.3005
R17805 gnd.n2942 gnd.n2939 9.3005
R17806 gnd.n2724 gnd.n2683 9.3005
R17807 gnd.n2719 gnd.n2718 9.3005
R17808 gnd.n2717 gnd.n2684 9.3005
R17809 gnd.n2716 gnd.n2715 9.3005
R17810 gnd.n2712 gnd.n2685 9.3005
R17811 gnd.n2709 gnd.n2708 9.3005
R17812 gnd.n2707 gnd.n2686 9.3005
R17813 gnd.n2706 gnd.n2705 9.3005
R17814 gnd.n2702 gnd.n2687 9.3005
R17815 gnd.n2699 gnd.n2698 9.3005
R17816 gnd.n2697 gnd.n2688 9.3005
R17817 gnd.n2696 gnd.n2695 9.3005
R17818 gnd.n2692 gnd.n2690 9.3005
R17819 gnd.n2689 gnd.n2669 9.3005
R17820 gnd.n2936 gnd.n2668 9.3005
R17821 gnd.n2938 gnd.n2937 9.3005
R17822 gnd.n2726 gnd.n2725 9.3005
R17823 gnd.n2949 gnd.n2655 9.3005
R17824 gnd.n2956 gnd.n2656 9.3005
R17825 gnd.n2958 gnd.n2957 9.3005
R17826 gnd.n2959 gnd.n2636 9.3005
R17827 gnd.n2978 gnd.n2977 9.3005
R17828 gnd.n2980 gnd.n2628 9.3005
R17829 gnd.n2987 gnd.n2630 9.3005
R17830 gnd.n2988 gnd.n2625 9.3005
R17831 gnd.n2990 gnd.n2989 9.3005
R17832 gnd.n2626 gnd.n2611 9.3005
R17833 gnd.n3006 gnd.n2609 9.3005
R17834 gnd.n3010 gnd.n3009 9.3005
R17835 gnd.n3008 gnd.n2585 9.3005
R17836 gnd.n3045 gnd.n2584 9.3005
R17837 gnd.n3048 gnd.n3047 9.3005
R17838 gnd.n2581 gnd.n2580 9.3005
R17839 gnd.n3054 gnd.n2582 9.3005
R17840 gnd.n3056 gnd.n3055 9.3005
R17841 gnd.n3058 gnd.n2579 9.3005
R17842 gnd.n3061 gnd.n3060 9.3005
R17843 gnd.n3064 gnd.n3062 9.3005
R17844 gnd.n3066 gnd.n3065 9.3005
R17845 gnd.n3072 gnd.n3067 9.3005
R17846 gnd.n3071 gnd.n3070 9.3005
R17847 gnd.n2455 gnd.n2454 9.3005
R17848 gnd.n3138 gnd.n3137 9.3005
R17849 gnd.n3139 gnd.n2448 9.3005
R17850 gnd.n3147 gnd.n2447 9.3005
R17851 gnd.n3150 gnd.n3149 9.3005
R17852 gnd.n3152 gnd.n3151 9.3005
R17853 gnd.n3155 gnd.n2430 9.3005
R17854 gnd.n3153 gnd.n2428 9.3005
R17855 gnd.n3175 gnd.n2426 9.3005
R17856 gnd.n3177 gnd.n3176 9.3005
R17857 gnd.n2400 gnd.n2399 9.3005
R17858 gnd.n3223 gnd.n3222 9.3005
R17859 gnd.n3224 gnd.n2393 9.3005
R17860 gnd.n3232 gnd.n2392 9.3005
R17861 gnd.n3235 gnd.n3234 9.3005
R17862 gnd.n3237 gnd.n3236 9.3005
R17863 gnd.n3240 gnd.n2375 9.3005
R17864 gnd.n3238 gnd.n2373 9.3005
R17865 gnd.n3260 gnd.n2371 9.3005
R17866 gnd.n3262 gnd.n3261 9.3005
R17867 gnd.n2346 gnd.n2345 9.3005
R17868 gnd.n3312 gnd.n3311 9.3005
R17869 gnd.n3313 gnd.n2339 9.3005
R17870 gnd.n3321 gnd.n2338 9.3005
R17871 gnd.n3580 gnd.n3579 9.3005
R17872 gnd.n3582 gnd.n3581 9.3005
R17873 gnd.n3583 gnd.n2319 9.3005
R17874 gnd.n3607 gnd.n3606 9.3005
R17875 gnd.n2320 gnd.n2282 9.3005
R17876 gnd.n2947 gnd.n2946 9.3005
R17877 gnd.n3663 gnd.n2283 9.3005
R17878 gnd.n3662 gnd.n2285 9.3005
R17879 gnd.n3659 gnd.n2286 9.3005
R17880 gnd.n3658 gnd.n2287 9.3005
R17881 gnd.n3655 gnd.n2288 9.3005
R17882 gnd.n3654 gnd.n2289 9.3005
R17883 gnd.n3651 gnd.n2290 9.3005
R17884 gnd.n3650 gnd.n2291 9.3005
R17885 gnd.n3647 gnd.n2292 9.3005
R17886 gnd.n3646 gnd.n2293 9.3005
R17887 gnd.n3643 gnd.n2294 9.3005
R17888 gnd.n3642 gnd.n2295 9.3005
R17889 gnd.n3639 gnd.n2296 9.3005
R17890 gnd.n3638 gnd.n2297 9.3005
R17891 gnd.n3635 gnd.n2298 9.3005
R17892 gnd.n3634 gnd.n2299 9.3005
R17893 gnd.n3631 gnd.n2300 9.3005
R17894 gnd.n3630 gnd.n2301 9.3005
R17895 gnd.n3627 gnd.n2302 9.3005
R17896 gnd.n3626 gnd.n2303 9.3005
R17897 gnd.n3623 gnd.n2304 9.3005
R17898 gnd.n3622 gnd.n2305 9.3005
R17899 gnd.n3619 gnd.n2309 9.3005
R17900 gnd.n3618 gnd.n2310 9.3005
R17901 gnd.n3615 gnd.n2311 9.3005
R17902 gnd.n3614 gnd.n2312 9.3005
R17903 gnd.n3665 gnd.n3664 9.3005
R17904 gnd.n3116 gnd.n3100 9.3005
R17905 gnd.n3115 gnd.n3101 9.3005
R17906 gnd.n3114 gnd.n3102 9.3005
R17907 gnd.n3112 gnd.n3103 9.3005
R17908 gnd.n3111 gnd.n3104 9.3005
R17909 gnd.n3109 gnd.n3105 9.3005
R17910 gnd.n3108 gnd.n3106 9.3005
R17911 gnd.n2418 gnd.n2417 9.3005
R17912 gnd.n3185 gnd.n3184 9.3005
R17913 gnd.n3186 gnd.n2416 9.3005
R17914 gnd.n3203 gnd.n3187 9.3005
R17915 gnd.n3202 gnd.n3188 9.3005
R17916 gnd.n3201 gnd.n3189 9.3005
R17917 gnd.n3199 gnd.n3190 9.3005
R17918 gnd.n3198 gnd.n3191 9.3005
R17919 gnd.n3196 gnd.n3192 9.3005
R17920 gnd.n3195 gnd.n3193 9.3005
R17921 gnd.n2362 gnd.n2361 9.3005
R17922 gnd.n3270 gnd.n3269 9.3005
R17923 gnd.n3271 gnd.n2360 9.3005
R17924 gnd.n3292 gnd.n3272 9.3005
R17925 gnd.n3291 gnd.n3273 9.3005
R17926 gnd.n3290 gnd.n3274 9.3005
R17927 gnd.n3287 gnd.n3275 9.3005
R17928 gnd.n3286 gnd.n3276 9.3005
R17929 gnd.n3284 gnd.n3277 9.3005
R17930 gnd.n3283 gnd.n3278 9.3005
R17931 gnd.n3281 gnd.n3280 9.3005
R17932 gnd.n3279 gnd.n2314 9.3005
R17933 gnd.n2857 gnd.n2856 9.3005
R17934 gnd.n2747 gnd.n2746 9.3005
R17935 gnd.n2871 gnd.n2870 9.3005
R17936 gnd.n2872 gnd.n2745 9.3005
R17937 gnd.n2874 gnd.n2873 9.3005
R17938 gnd.n2735 gnd.n2734 9.3005
R17939 gnd.n2887 gnd.n2886 9.3005
R17940 gnd.n2888 gnd.n2733 9.3005
R17941 gnd.n2920 gnd.n2889 9.3005
R17942 gnd.n2919 gnd.n2890 9.3005
R17943 gnd.n2918 gnd.n2891 9.3005
R17944 gnd.n2917 gnd.n2892 9.3005
R17945 gnd.n2914 gnd.n2893 9.3005
R17946 gnd.n2913 gnd.n2894 9.3005
R17947 gnd.n2912 gnd.n2895 9.3005
R17948 gnd.n2910 gnd.n2896 9.3005
R17949 gnd.n2909 gnd.n2897 9.3005
R17950 gnd.n2906 gnd.n2898 9.3005
R17951 gnd.n2905 gnd.n2899 9.3005
R17952 gnd.n2904 gnd.n2900 9.3005
R17953 gnd.n2902 gnd.n2901 9.3005
R17954 gnd.n2601 gnd.n2600 9.3005
R17955 gnd.n3018 gnd.n3017 9.3005
R17956 gnd.n3019 gnd.n2599 9.3005
R17957 gnd.n3023 gnd.n3020 9.3005
R17958 gnd.n3022 gnd.n3021 9.3005
R17959 gnd.n2523 gnd.n2522 9.3005
R17960 gnd.n3098 gnd.n3097 9.3005
R17961 gnd.n2855 gnd.n2756 9.3005
R17962 gnd.n2758 gnd.n2757 9.3005
R17963 gnd.n2802 gnd.n2800 9.3005
R17964 gnd.n2803 gnd.n2799 9.3005
R17965 gnd.n2806 gnd.n2795 9.3005
R17966 gnd.n2807 gnd.n2794 9.3005
R17967 gnd.n2810 gnd.n2793 9.3005
R17968 gnd.n2811 gnd.n2792 9.3005
R17969 gnd.n2814 gnd.n2791 9.3005
R17970 gnd.n2815 gnd.n2790 9.3005
R17971 gnd.n2818 gnd.n2789 9.3005
R17972 gnd.n2819 gnd.n2788 9.3005
R17973 gnd.n2822 gnd.n2787 9.3005
R17974 gnd.n2823 gnd.n2786 9.3005
R17975 gnd.n2826 gnd.n2785 9.3005
R17976 gnd.n2827 gnd.n2784 9.3005
R17977 gnd.n2830 gnd.n2783 9.3005
R17978 gnd.n2831 gnd.n2782 9.3005
R17979 gnd.n2834 gnd.n2781 9.3005
R17980 gnd.n2835 gnd.n2780 9.3005
R17981 gnd.n2838 gnd.n2779 9.3005
R17982 gnd.n2839 gnd.n2778 9.3005
R17983 gnd.n2842 gnd.n2777 9.3005
R17984 gnd.n2844 gnd.n2776 9.3005
R17985 gnd.n2845 gnd.n2775 9.3005
R17986 gnd.n2846 gnd.n2774 9.3005
R17987 gnd.n2847 gnd.n2773 9.3005
R17988 gnd.n2854 gnd.n2853 9.3005
R17989 gnd.n2863 gnd.n2862 9.3005
R17990 gnd.n2864 gnd.n2750 9.3005
R17991 gnd.n2866 gnd.n2865 9.3005
R17992 gnd.n2741 gnd.n2740 9.3005
R17993 gnd.n2879 gnd.n2878 9.3005
R17994 gnd.n2880 gnd.n2739 9.3005
R17995 gnd.n2882 gnd.n2881 9.3005
R17996 gnd.n2728 gnd.n2727 9.3005
R17997 gnd.n2925 gnd.n2924 9.3005
R17998 gnd.n2926 gnd.n2682 9.3005
R17999 gnd.n2930 gnd.n2928 9.3005
R18000 gnd.n2929 gnd.n2661 9.3005
R18001 gnd.n2948 gnd.n2660 9.3005
R18002 gnd.n2951 gnd.n2950 9.3005
R18003 gnd.n2654 gnd.n2653 9.3005
R18004 gnd.n2962 gnd.n2960 9.3005
R18005 gnd.n2961 gnd.n2635 9.3005
R18006 gnd.n2979 gnd.n2634 9.3005
R18007 gnd.n2982 gnd.n2981 9.3005
R18008 gnd.n2629 gnd.n2624 9.3005
R18009 gnd.n2992 gnd.n2991 9.3005
R18010 gnd.n2627 gnd.n2607 9.3005
R18011 gnd.n3013 gnd.n2608 9.3005
R18012 gnd.n3012 gnd.n3011 9.3005
R18013 gnd.n2610 gnd.n2586 9.3005
R18014 gnd.n3044 gnd.n3043 9.3005
R18015 gnd.n3046 gnd.n2531 9.3005
R18016 gnd.n3093 gnd.n2532 9.3005
R18017 gnd.n3092 gnd.n2533 9.3005
R18018 gnd.n3091 gnd.n2534 9.3005
R18019 gnd.n3057 gnd.n2535 9.3005
R18020 gnd.n3059 gnd.n2553 9.3005
R18021 gnd.n3079 gnd.n2554 9.3005
R18022 gnd.n3078 gnd.n2555 9.3005
R18023 gnd.n3077 gnd.n2556 9.3005
R18024 gnd.n3068 gnd.n2557 9.3005
R18025 gnd.n3069 gnd.n2456 9.3005
R18026 gnd.n3135 gnd.n3134 9.3005
R18027 gnd.n3136 gnd.n2449 9.3005
R18028 gnd.n3146 gnd.n3145 9.3005
R18029 gnd.n3148 gnd.n2445 9.3005
R18030 gnd.n3158 gnd.n2446 9.3005
R18031 gnd.n3157 gnd.n3156 9.3005
R18032 gnd.n3154 gnd.n2424 9.3005
R18033 gnd.n3180 gnd.n2425 9.3005
R18034 gnd.n3179 gnd.n3178 9.3005
R18035 gnd.n2427 gnd.n2401 9.3005
R18036 gnd.n3220 gnd.n3219 9.3005
R18037 gnd.n3221 gnd.n2394 9.3005
R18038 gnd.n3231 gnd.n3230 9.3005
R18039 gnd.n3233 gnd.n2390 9.3005
R18040 gnd.n3243 gnd.n2391 9.3005
R18041 gnd.n3242 gnd.n3241 9.3005
R18042 gnd.n3239 gnd.n2369 9.3005
R18043 gnd.n3265 gnd.n2370 9.3005
R18044 gnd.n3264 gnd.n3263 9.3005
R18045 gnd.n2372 gnd.n2347 9.3005
R18046 gnd.n3309 gnd.n3308 9.3005
R18047 gnd.n3310 gnd.n2340 9.3005
R18048 gnd.n3320 gnd.n3319 9.3005
R18049 gnd.n3578 gnd.n2336 9.3005
R18050 gnd.n3586 gnd.n2337 9.3005
R18051 gnd.n3585 gnd.n3584 9.3005
R18052 gnd.n2318 gnd.n2317 9.3005
R18053 gnd.n3609 gnd.n3608 9.3005
R18054 gnd.n2752 gnd.n2751 9.3005
R18055 gnd.n6243 gnd.n6242 9.3005
R18056 gnd.n559 gnd.n558 9.3005
R18057 gnd.n6250 gnd.n6249 9.3005
R18058 gnd.n6251 gnd.n557 9.3005
R18059 gnd.n6253 gnd.n6252 9.3005
R18060 gnd.n553 gnd.n552 9.3005
R18061 gnd.n6260 gnd.n6259 9.3005
R18062 gnd.n6261 gnd.n551 9.3005
R18063 gnd.n6263 gnd.n6262 9.3005
R18064 gnd.n547 gnd.n546 9.3005
R18065 gnd.n6270 gnd.n6269 9.3005
R18066 gnd.n6271 gnd.n545 9.3005
R18067 gnd.n6273 gnd.n6272 9.3005
R18068 gnd.n541 gnd.n540 9.3005
R18069 gnd.n6280 gnd.n6279 9.3005
R18070 gnd.n6281 gnd.n539 9.3005
R18071 gnd.n6283 gnd.n6282 9.3005
R18072 gnd.n535 gnd.n534 9.3005
R18073 gnd.n6290 gnd.n6289 9.3005
R18074 gnd.n6291 gnd.n533 9.3005
R18075 gnd.n6293 gnd.n6292 9.3005
R18076 gnd.n529 gnd.n528 9.3005
R18077 gnd.n6300 gnd.n6299 9.3005
R18078 gnd.n6301 gnd.n527 9.3005
R18079 gnd.n6303 gnd.n6302 9.3005
R18080 gnd.n523 gnd.n522 9.3005
R18081 gnd.n6310 gnd.n6309 9.3005
R18082 gnd.n6311 gnd.n521 9.3005
R18083 gnd.n6313 gnd.n6312 9.3005
R18084 gnd.n517 gnd.n516 9.3005
R18085 gnd.n6320 gnd.n6319 9.3005
R18086 gnd.n6321 gnd.n515 9.3005
R18087 gnd.n6323 gnd.n6322 9.3005
R18088 gnd.n511 gnd.n510 9.3005
R18089 gnd.n6330 gnd.n6329 9.3005
R18090 gnd.n6331 gnd.n509 9.3005
R18091 gnd.n6333 gnd.n6332 9.3005
R18092 gnd.n505 gnd.n504 9.3005
R18093 gnd.n6340 gnd.n6339 9.3005
R18094 gnd.n6341 gnd.n503 9.3005
R18095 gnd.n6343 gnd.n6342 9.3005
R18096 gnd.n499 gnd.n498 9.3005
R18097 gnd.n6350 gnd.n6349 9.3005
R18098 gnd.n6351 gnd.n497 9.3005
R18099 gnd.n6353 gnd.n6352 9.3005
R18100 gnd.n493 gnd.n492 9.3005
R18101 gnd.n6360 gnd.n6359 9.3005
R18102 gnd.n6361 gnd.n491 9.3005
R18103 gnd.n6363 gnd.n6362 9.3005
R18104 gnd.n487 gnd.n486 9.3005
R18105 gnd.n6370 gnd.n6369 9.3005
R18106 gnd.n6371 gnd.n485 9.3005
R18107 gnd.n6373 gnd.n6372 9.3005
R18108 gnd.n481 gnd.n480 9.3005
R18109 gnd.n6380 gnd.n6379 9.3005
R18110 gnd.n6381 gnd.n479 9.3005
R18111 gnd.n6383 gnd.n6382 9.3005
R18112 gnd.n475 gnd.n474 9.3005
R18113 gnd.n6390 gnd.n6389 9.3005
R18114 gnd.n6391 gnd.n473 9.3005
R18115 gnd.n6393 gnd.n6392 9.3005
R18116 gnd.n469 gnd.n468 9.3005
R18117 gnd.n6400 gnd.n6399 9.3005
R18118 gnd.n6401 gnd.n467 9.3005
R18119 gnd.n6403 gnd.n6402 9.3005
R18120 gnd.n463 gnd.n462 9.3005
R18121 gnd.n6410 gnd.n6409 9.3005
R18122 gnd.n6411 gnd.n461 9.3005
R18123 gnd.n6413 gnd.n6412 9.3005
R18124 gnd.n457 gnd.n456 9.3005
R18125 gnd.n6420 gnd.n6419 9.3005
R18126 gnd.n6421 gnd.n455 9.3005
R18127 gnd.n6423 gnd.n6422 9.3005
R18128 gnd.n451 gnd.n450 9.3005
R18129 gnd.n6430 gnd.n6429 9.3005
R18130 gnd.n6431 gnd.n449 9.3005
R18131 gnd.n6433 gnd.n6432 9.3005
R18132 gnd.n445 gnd.n444 9.3005
R18133 gnd.n6440 gnd.n6439 9.3005
R18134 gnd.n6441 gnd.n443 9.3005
R18135 gnd.n6443 gnd.n6442 9.3005
R18136 gnd.n439 gnd.n438 9.3005
R18137 gnd.n6450 gnd.n6449 9.3005
R18138 gnd.n6451 gnd.n437 9.3005
R18139 gnd.n6453 gnd.n6452 9.3005
R18140 gnd.n433 gnd.n432 9.3005
R18141 gnd.n6460 gnd.n6459 9.3005
R18142 gnd.n6461 gnd.n431 9.3005
R18143 gnd.n6463 gnd.n6462 9.3005
R18144 gnd.n427 gnd.n426 9.3005
R18145 gnd.n6470 gnd.n6469 9.3005
R18146 gnd.n6471 gnd.n425 9.3005
R18147 gnd.n6473 gnd.n6472 9.3005
R18148 gnd.n421 gnd.n420 9.3005
R18149 gnd.n6480 gnd.n6479 9.3005
R18150 gnd.n6481 gnd.n419 9.3005
R18151 gnd.n6483 gnd.n6482 9.3005
R18152 gnd.n415 gnd.n414 9.3005
R18153 gnd.n6490 gnd.n6489 9.3005
R18154 gnd.n6491 gnd.n413 9.3005
R18155 gnd.n6493 gnd.n6492 9.3005
R18156 gnd.n409 gnd.n408 9.3005
R18157 gnd.n6500 gnd.n6499 9.3005
R18158 gnd.n6501 gnd.n407 9.3005
R18159 gnd.n6503 gnd.n6502 9.3005
R18160 gnd.n403 gnd.n402 9.3005
R18161 gnd.n6510 gnd.n6509 9.3005
R18162 gnd.n6511 gnd.n401 9.3005
R18163 gnd.n6513 gnd.n6512 9.3005
R18164 gnd.n397 gnd.n396 9.3005
R18165 gnd.n6520 gnd.n6519 9.3005
R18166 gnd.n6521 gnd.n395 9.3005
R18167 gnd.n6523 gnd.n6522 9.3005
R18168 gnd.n391 gnd.n390 9.3005
R18169 gnd.n6530 gnd.n6529 9.3005
R18170 gnd.n6531 gnd.n389 9.3005
R18171 gnd.n6533 gnd.n6532 9.3005
R18172 gnd.n385 gnd.n384 9.3005
R18173 gnd.n6540 gnd.n6539 9.3005
R18174 gnd.n6541 gnd.n383 9.3005
R18175 gnd.n6543 gnd.n6542 9.3005
R18176 gnd.n379 gnd.n378 9.3005
R18177 gnd.n6550 gnd.n6549 9.3005
R18178 gnd.n6551 gnd.n377 9.3005
R18179 gnd.n6553 gnd.n6552 9.3005
R18180 gnd.n373 gnd.n372 9.3005
R18181 gnd.n6560 gnd.n6559 9.3005
R18182 gnd.n6561 gnd.n371 9.3005
R18183 gnd.n6563 gnd.n6562 9.3005
R18184 gnd.n367 gnd.n366 9.3005
R18185 gnd.n6570 gnd.n6569 9.3005
R18186 gnd.n6571 gnd.n365 9.3005
R18187 gnd.n6573 gnd.n6572 9.3005
R18188 gnd.n361 gnd.n360 9.3005
R18189 gnd.n6580 gnd.n6579 9.3005
R18190 gnd.n6581 gnd.n359 9.3005
R18191 gnd.n6583 gnd.n6582 9.3005
R18192 gnd.n355 gnd.n354 9.3005
R18193 gnd.n6590 gnd.n6589 9.3005
R18194 gnd.n6591 gnd.n353 9.3005
R18195 gnd.n6593 gnd.n6592 9.3005
R18196 gnd.n349 gnd.n348 9.3005
R18197 gnd.n6600 gnd.n6599 9.3005
R18198 gnd.n6601 gnd.n347 9.3005
R18199 gnd.n6603 gnd.n6602 9.3005
R18200 gnd.n343 gnd.n342 9.3005
R18201 gnd.n6610 gnd.n6609 9.3005
R18202 gnd.n6611 gnd.n341 9.3005
R18203 gnd.n6613 gnd.n6612 9.3005
R18204 gnd.n337 gnd.n336 9.3005
R18205 gnd.n6620 gnd.n6619 9.3005
R18206 gnd.n6621 gnd.n335 9.3005
R18207 gnd.n6623 gnd.n6622 9.3005
R18208 gnd.n331 gnd.n330 9.3005
R18209 gnd.n6630 gnd.n6629 9.3005
R18210 gnd.n6631 gnd.n329 9.3005
R18211 gnd.n6633 gnd.n6632 9.3005
R18212 gnd.n325 gnd.n324 9.3005
R18213 gnd.n6640 gnd.n6639 9.3005
R18214 gnd.n6641 gnd.n323 9.3005
R18215 gnd.n6643 gnd.n6642 9.3005
R18216 gnd.n319 gnd.n318 9.3005
R18217 gnd.n6650 gnd.n6649 9.3005
R18218 gnd.n6651 gnd.n317 9.3005
R18219 gnd.n6654 gnd.n6653 9.3005
R18220 gnd.n6652 gnd.n313 9.3005
R18221 gnd.n6660 gnd.n312 9.3005
R18222 gnd.n6662 gnd.n6661 9.3005
R18223 gnd.n308 gnd.n307 9.3005
R18224 gnd.n6671 gnd.n6670 9.3005
R18225 gnd.n6672 gnd.n306 9.3005
R18226 gnd.n6674 gnd.n6673 9.3005
R18227 gnd.n302 gnd.n301 9.3005
R18228 gnd.n6681 gnd.n6680 9.3005
R18229 gnd.n6682 gnd.n300 9.3005
R18230 gnd.n6684 gnd.n6683 9.3005
R18231 gnd.n296 gnd.n295 9.3005
R18232 gnd.n6691 gnd.n6690 9.3005
R18233 gnd.n6692 gnd.n294 9.3005
R18234 gnd.n6694 gnd.n6693 9.3005
R18235 gnd.n290 gnd.n289 9.3005
R18236 gnd.n6701 gnd.n6700 9.3005
R18237 gnd.n6702 gnd.n288 9.3005
R18238 gnd.n6704 gnd.n6703 9.3005
R18239 gnd.n284 gnd.n283 9.3005
R18240 gnd.n6711 gnd.n6710 9.3005
R18241 gnd.n6712 gnd.n282 9.3005
R18242 gnd.n6714 gnd.n6713 9.3005
R18243 gnd.n278 gnd.n277 9.3005
R18244 gnd.n6721 gnd.n6720 9.3005
R18245 gnd.n6722 gnd.n276 9.3005
R18246 gnd.n6724 gnd.n6723 9.3005
R18247 gnd.n272 gnd.n271 9.3005
R18248 gnd.n6731 gnd.n6730 9.3005
R18249 gnd.n6732 gnd.n270 9.3005
R18250 gnd.n6734 gnd.n6733 9.3005
R18251 gnd.n266 gnd.n265 9.3005
R18252 gnd.n6741 gnd.n6740 9.3005
R18253 gnd.n6742 gnd.n264 9.3005
R18254 gnd.n6744 gnd.n6743 9.3005
R18255 gnd.n260 gnd.n259 9.3005
R18256 gnd.n6751 gnd.n6750 9.3005
R18257 gnd.n6752 gnd.n258 9.3005
R18258 gnd.n6754 gnd.n6753 9.3005
R18259 gnd.n254 gnd.n253 9.3005
R18260 gnd.n6761 gnd.n6760 9.3005
R18261 gnd.n6762 gnd.n252 9.3005
R18262 gnd.n6764 gnd.n6763 9.3005
R18263 gnd.n248 gnd.n247 9.3005
R18264 gnd.n6771 gnd.n6770 9.3005
R18265 gnd.n6772 gnd.n246 9.3005
R18266 gnd.n6774 gnd.n6773 9.3005
R18267 gnd.n242 gnd.n241 9.3005
R18268 gnd.n6781 gnd.n6780 9.3005
R18269 gnd.n6782 gnd.n240 9.3005
R18270 gnd.n6784 gnd.n6783 9.3005
R18271 gnd.n236 gnd.n235 9.3005
R18272 gnd.n6791 gnd.n6790 9.3005
R18273 gnd.n6792 gnd.n234 9.3005
R18274 gnd.n6794 gnd.n6793 9.3005
R18275 gnd.n230 gnd.n229 9.3005
R18276 gnd.n6801 gnd.n6800 9.3005
R18277 gnd.n6802 gnd.n228 9.3005
R18278 gnd.n6804 gnd.n6803 9.3005
R18279 gnd.n224 gnd.n223 9.3005
R18280 gnd.n6811 gnd.n6810 9.3005
R18281 gnd.n6812 gnd.n222 9.3005
R18282 gnd.n6814 gnd.n6813 9.3005
R18283 gnd.n218 gnd.n217 9.3005
R18284 gnd.n6821 gnd.n6820 9.3005
R18285 gnd.n6822 gnd.n216 9.3005
R18286 gnd.n6824 gnd.n6823 9.3005
R18287 gnd.n212 gnd.n211 9.3005
R18288 gnd.n6831 gnd.n6830 9.3005
R18289 gnd.n6832 gnd.n210 9.3005
R18290 gnd.n6834 gnd.n6833 9.3005
R18291 gnd.n206 gnd.n205 9.3005
R18292 gnd.n6841 gnd.n6840 9.3005
R18293 gnd.n6842 gnd.n204 9.3005
R18294 gnd.n6844 gnd.n6843 9.3005
R18295 gnd.n200 gnd.n199 9.3005
R18296 gnd.n6851 gnd.n6850 9.3005
R18297 gnd.n6852 gnd.n198 9.3005
R18298 gnd.n6854 gnd.n6853 9.3005
R18299 gnd.n194 gnd.n193 9.3005
R18300 gnd.n6861 gnd.n6860 9.3005
R18301 gnd.n6862 gnd.n192 9.3005
R18302 gnd.n6864 gnd.n6863 9.3005
R18303 gnd.n188 gnd.n187 9.3005
R18304 gnd.n6872 gnd.n6871 9.3005
R18305 gnd.n6873 gnd.n186 9.3005
R18306 gnd.n6875 gnd.n6874 9.3005
R18307 gnd.n6664 gnd.n6663 9.3005
R18308 gnd.n7307 gnd.n7306 9.3005
R18309 gnd.n7305 gnd.n69 9.3005
R18310 gnd.n176 gnd.n71 9.3005
R18311 gnd.n6894 gnd.n6893 9.3005
R18312 gnd.n6895 gnd.n175 9.3005
R18313 gnd.n7214 gnd.n6896 9.3005
R18314 gnd.n7213 gnd.n6897 9.3005
R18315 gnd.n7212 gnd.n6898 9.3005
R18316 gnd.n7210 gnd.n6899 9.3005
R18317 gnd.n7209 gnd.n6900 9.3005
R18318 gnd.n7207 gnd.n6901 9.3005
R18319 gnd.n7206 gnd.n6902 9.3005
R18320 gnd.n7204 gnd.n6903 9.3005
R18321 gnd.n7203 gnd.n6904 9.3005
R18322 gnd.n7201 gnd.n6905 9.3005
R18323 gnd.n7200 gnd.n6906 9.3005
R18324 gnd.n7198 gnd.n6907 9.3005
R18325 gnd.n7197 gnd.n6908 9.3005
R18326 gnd.n7195 gnd.n6909 9.3005
R18327 gnd.n7194 gnd.n6910 9.3005
R18328 gnd.n7192 gnd.n7191 9.3005
R18329 gnd.n6935 gnd.n6931 9.3005
R18330 gnd.n6939 gnd.n6938 9.3005
R18331 gnd.n6940 gnd.n6930 9.3005
R18332 gnd.n6942 gnd.n6941 9.3005
R18333 gnd.n6945 gnd.n6929 9.3005
R18334 gnd.n6949 gnd.n6948 9.3005
R18335 gnd.n6950 gnd.n6928 9.3005
R18336 gnd.n6952 gnd.n6951 9.3005
R18337 gnd.n6955 gnd.n6927 9.3005
R18338 gnd.n6959 gnd.n6958 9.3005
R18339 gnd.n6960 gnd.n6926 9.3005
R18340 gnd.n6962 gnd.n6961 9.3005
R18341 gnd.n6965 gnd.n6925 9.3005
R18342 gnd.n6968 gnd.n6967 9.3005
R18343 gnd.n6969 gnd.n6924 9.3005
R18344 gnd.n6971 gnd.n6970 9.3005
R18345 gnd.n6914 gnd.n6911 9.3005
R18346 gnd.n7190 gnd.n7189 9.3005
R18347 gnd.n6933 gnd.n6932 9.3005
R18348 gnd.n7007 gnd.n7004 9.3005
R18349 gnd.n7183 gnd.n7008 9.3005
R18350 gnd.n7182 gnd.n7009 9.3005
R18351 gnd.n7181 gnd.n7010 9.3005
R18352 gnd.n7178 gnd.n7011 9.3005
R18353 gnd.n7177 gnd.n7012 9.3005
R18354 gnd.n7174 gnd.n7013 9.3005
R18355 gnd.n7173 gnd.n7014 9.3005
R18356 gnd.n7170 gnd.n7015 9.3005
R18357 gnd.n7169 gnd.n7016 9.3005
R18358 gnd.n7166 gnd.n7017 9.3005
R18359 gnd.n7165 gnd.n7018 9.3005
R18360 gnd.n7162 gnd.n7019 9.3005
R18361 gnd.n7161 gnd.n7020 9.3005
R18362 gnd.n7158 gnd.n7021 9.3005
R18363 gnd.n7157 gnd.n7022 9.3005
R18364 gnd.n7154 gnd.n7023 9.3005
R18365 gnd.n7150 gnd.n7024 9.3005
R18366 gnd.n7147 gnd.n7025 9.3005
R18367 gnd.n7146 gnd.n7026 9.3005
R18368 gnd.n7143 gnd.n7027 9.3005
R18369 gnd.n7142 gnd.n7028 9.3005
R18370 gnd.n7139 gnd.n7029 9.3005
R18371 gnd.n7138 gnd.n7030 9.3005
R18372 gnd.n7135 gnd.n7031 9.3005
R18373 gnd.n7134 gnd.n7032 9.3005
R18374 gnd.n7131 gnd.n7033 9.3005
R18375 gnd.n7130 gnd.n7034 9.3005
R18376 gnd.n7127 gnd.n7035 9.3005
R18377 gnd.n7126 gnd.n7036 9.3005
R18378 gnd.n7123 gnd.n7037 9.3005
R18379 gnd.n7122 gnd.n7038 9.3005
R18380 gnd.n7119 gnd.n7039 9.3005
R18381 gnd.n7118 gnd.n7040 9.3005
R18382 gnd.n7115 gnd.n7041 9.3005
R18383 gnd.n7114 gnd.n7042 9.3005
R18384 gnd.n7111 gnd.n7110 9.3005
R18385 gnd.n7109 gnd.n7043 9.3005
R18386 gnd.n7108 gnd.n7107 9.3005
R18387 gnd.n7104 gnd.n7046 9.3005
R18388 gnd.n7101 gnd.n7047 9.3005
R18389 gnd.n7100 gnd.n7048 9.3005
R18390 gnd.n7097 gnd.n7049 9.3005
R18391 gnd.n7096 gnd.n7050 9.3005
R18392 gnd.n7093 gnd.n7051 9.3005
R18393 gnd.n7092 gnd.n7052 9.3005
R18394 gnd.n7089 gnd.n7053 9.3005
R18395 gnd.n7088 gnd.n7054 9.3005
R18396 gnd.n7085 gnd.n7055 9.3005
R18397 gnd.n7084 gnd.n7056 9.3005
R18398 gnd.n7081 gnd.n7057 9.3005
R18399 gnd.n7080 gnd.n7058 9.3005
R18400 gnd.n7077 gnd.n7059 9.3005
R18401 gnd.n7076 gnd.n7060 9.3005
R18402 gnd.n7073 gnd.n7061 9.3005
R18403 gnd.n7072 gnd.n7062 9.3005
R18404 gnd.n7069 gnd.n7068 9.3005
R18405 gnd.n7067 gnd.n7064 9.3005
R18406 gnd.n7006 gnd.n7005 9.3005
R18407 gnd.n5462 gnd.n5461 9.3005
R18408 gnd.n1498 gnd.n1497 9.3005
R18409 gnd.n1522 gnd.n1521 9.3005
R18410 gnd.n5449 gnd.n1523 9.3005
R18411 gnd.n5448 gnd.n1524 9.3005
R18412 gnd.n5447 gnd.n1525 9.3005
R18413 gnd.n5279 gnd.n1526 9.3005
R18414 gnd.n5437 gnd.n1543 9.3005
R18415 gnd.n5436 gnd.n1544 9.3005
R18416 gnd.n5435 gnd.n1545 9.3005
R18417 gnd.n5285 gnd.n1546 9.3005
R18418 gnd.n5425 gnd.n1563 9.3005
R18419 gnd.n5424 gnd.n1564 9.3005
R18420 gnd.n5423 gnd.n1565 9.3005
R18421 gnd.n5362 gnd.n1566 9.3005
R18422 gnd.n5413 gnd.n1580 9.3005
R18423 gnd.n5412 gnd.n1581 9.3005
R18424 gnd.n5411 gnd.n1582 9.3005
R18425 gnd.n5382 gnd.n1583 9.3005
R18426 gnd.n5384 gnd.n5383 9.3005
R18427 gnd.n1607 gnd.n1606 9.3005
R18428 gnd.n5393 gnd.n5392 9.3005
R18429 gnd.n180 gnd.n179 9.3005
R18430 gnd.n6887 gnd.n6886 9.3005
R18431 gnd.n6888 gnd.n96 9.3005
R18432 gnd.n7293 gnd.n97 9.3005
R18433 gnd.n7292 gnd.n98 9.3005
R18434 gnd.n7291 gnd.n99 9.3005
R18435 gnd.n7220 gnd.n100 9.3005
R18436 gnd.n7281 gnd.n115 9.3005
R18437 gnd.n7280 gnd.n116 9.3005
R18438 gnd.n7279 gnd.n117 9.3005
R18439 gnd.n7227 gnd.n118 9.3005
R18440 gnd.n7269 gnd.n135 9.3005
R18441 gnd.n7268 gnd.n136 9.3005
R18442 gnd.n7267 gnd.n137 9.3005
R18443 gnd.n7234 gnd.n138 9.3005
R18444 gnd.n7257 gnd.n154 9.3005
R18445 gnd.n7256 gnd.n155 9.3005
R18446 gnd.n7255 gnd.n156 9.3005
R18447 gnd.n172 gnd.n157 9.3005
R18448 gnd.n7245 gnd.n7244 9.3005
R18449 gnd.n5463 gnd.n1496 9.3005
R18450 gnd.n5461 gnd.n5460 9.3005
R18451 gnd.n5459 gnd.n1498 9.3005
R18452 gnd.n1522 gnd.n1499 9.3005
R18453 gnd.n5274 gnd.n1523 9.3005
R18454 gnd.n5277 gnd.n1524 9.3005
R18455 gnd.n5278 gnd.n1525 9.3005
R18456 gnd.n5283 gnd.n5279 9.3005
R18457 gnd.n5284 gnd.n1543 9.3005
R18458 gnd.n5288 gnd.n1544 9.3005
R18459 gnd.n5287 gnd.n1545 9.3005
R18460 gnd.n5286 gnd.n5285 9.3005
R18461 gnd.n1618 gnd.n1563 9.3005
R18462 gnd.n5360 gnd.n1564 9.3005
R18463 gnd.n5361 gnd.n1565 9.3005
R18464 gnd.n5363 gnd.n5362 9.3005
R18465 gnd.n1612 gnd.n1580 9.3005
R18466 gnd.n5379 gnd.n1581 9.3005
R18467 gnd.n5380 gnd.n1582 9.3005
R18468 gnd.n5382 gnd.n5381 9.3005
R18469 gnd.n5383 gnd.n1608 9.3005
R18470 gnd.n5389 gnd.n1607 9.3005
R18471 gnd.n5392 gnd.n5391 9.3005
R18472 gnd.n5390 gnd.n179 9.3005
R18473 gnd.n6887 gnd.n178 9.3005
R18474 gnd.n6889 gnd.n6888 9.3005
R18475 gnd.n174 gnd.n97 9.3005
R18476 gnd.n7218 gnd.n98 9.3005
R18477 gnd.n7219 gnd.n99 9.3005
R18478 gnd.n7222 gnd.n7220 9.3005
R18479 gnd.n7223 gnd.n115 9.3005
R18480 gnd.n7225 gnd.n116 9.3005
R18481 gnd.n7226 gnd.n117 9.3005
R18482 gnd.n7229 gnd.n7227 9.3005
R18483 gnd.n7230 gnd.n135 9.3005
R18484 gnd.n7232 gnd.n136 9.3005
R18485 gnd.n7233 gnd.n137 9.3005
R18486 gnd.n7236 gnd.n7234 9.3005
R18487 gnd.n7237 gnd.n154 9.3005
R18488 gnd.n7239 gnd.n155 9.3005
R18489 gnd.n7240 gnd.n156 9.3005
R18490 gnd.n7242 gnd.n172 9.3005
R18491 gnd.n7244 gnd.n7243 9.3005
R18492 gnd.n1496 gnd.n1490 9.3005
R18493 gnd.n5473 gnd.n5472 9.3005
R18494 gnd.n5476 gnd.n1488 9.3005
R18495 gnd.n5477 gnd.n1487 9.3005
R18496 gnd.n5480 gnd.n1486 9.3005
R18497 gnd.n5481 gnd.n1485 9.3005
R18498 gnd.n5484 gnd.n1484 9.3005
R18499 gnd.n5485 gnd.n1483 9.3005
R18500 gnd.n5488 gnd.n1482 9.3005
R18501 gnd.n5489 gnd.n1481 9.3005
R18502 gnd.n5492 gnd.n1480 9.3005
R18503 gnd.n5493 gnd.n1479 9.3005
R18504 gnd.n5496 gnd.n1478 9.3005
R18505 gnd.n5497 gnd.n1477 9.3005
R18506 gnd.n5500 gnd.n1476 9.3005
R18507 gnd.n5501 gnd.n1475 9.3005
R18508 gnd.n5504 gnd.n1474 9.3005
R18509 gnd.n5505 gnd.n1473 9.3005
R18510 gnd.n5508 gnd.n1472 9.3005
R18511 gnd.n5509 gnd.n1471 9.3005
R18512 gnd.n5512 gnd.n1470 9.3005
R18513 gnd.n5516 gnd.n1466 9.3005
R18514 gnd.n5517 gnd.n1465 9.3005
R18515 gnd.n5520 gnd.n1464 9.3005
R18516 gnd.n5521 gnd.n1463 9.3005
R18517 gnd.n5524 gnd.n1462 9.3005
R18518 gnd.n5525 gnd.n1461 9.3005
R18519 gnd.n5528 gnd.n1460 9.3005
R18520 gnd.n5529 gnd.n1459 9.3005
R18521 gnd.n5532 gnd.n1458 9.3005
R18522 gnd.n5534 gnd.n1454 9.3005
R18523 gnd.n5537 gnd.n1453 9.3005
R18524 gnd.n5538 gnd.n1452 9.3005
R18525 gnd.n5541 gnd.n1451 9.3005
R18526 gnd.n5542 gnd.n1450 9.3005
R18527 gnd.n5545 gnd.n1449 9.3005
R18528 gnd.n5546 gnd.n1448 9.3005
R18529 gnd.n5549 gnd.n1447 9.3005
R18530 gnd.n5551 gnd.n1444 9.3005
R18531 gnd.n5554 gnd.n1443 9.3005
R18532 gnd.n5555 gnd.n1442 9.3005
R18533 gnd.n5558 gnd.n1441 9.3005
R18534 gnd.n5559 gnd.n1440 9.3005
R18535 gnd.n5562 gnd.n1439 9.3005
R18536 gnd.n5563 gnd.n1438 9.3005
R18537 gnd.n5566 gnd.n1437 9.3005
R18538 gnd.n5567 gnd.n1436 9.3005
R18539 gnd.n5570 gnd.n1435 9.3005
R18540 gnd.n5571 gnd.n1434 9.3005
R18541 gnd.n5574 gnd.n1433 9.3005
R18542 gnd.n5575 gnd.n1432 9.3005
R18543 gnd.n5578 gnd.n1431 9.3005
R18544 gnd.n5580 gnd.n1430 9.3005
R18545 gnd.n5581 gnd.n1429 9.3005
R18546 gnd.n5582 gnd.n1428 9.3005
R18547 gnd.n5583 gnd.n1427 9.3005
R18548 gnd.n5513 gnd.n1467 9.3005
R18549 gnd.n5471 gnd.n5468 9.3005
R18550 gnd.n1509 gnd.n1506 9.3005
R18551 gnd.n5455 gnd.n1510 9.3005
R18552 gnd.n5454 gnd.n1511 9.3005
R18553 gnd.n5453 gnd.n1512 9.3005
R18554 gnd.n1532 gnd.n1513 9.3005
R18555 gnd.n5443 gnd.n1533 9.3005
R18556 gnd.n5442 gnd.n1534 9.3005
R18557 gnd.n5441 gnd.n1535 9.3005
R18558 gnd.n1553 gnd.n1536 9.3005
R18559 gnd.n5431 gnd.n1554 9.3005
R18560 gnd.n5430 gnd.n1555 9.3005
R18561 gnd.n5429 gnd.n1556 9.3005
R18562 gnd.n1572 gnd.n1557 9.3005
R18563 gnd.n5419 gnd.n1573 9.3005
R18564 gnd.n5418 gnd.n82 9.3005
R18565 gnd.n87 gnd.n81 9.3005
R18566 gnd.n7287 gnd.n106 9.3005
R18567 gnd.n7286 gnd.n107 9.3005
R18568 gnd.n7285 gnd.n108 9.3005
R18569 gnd.n124 gnd.n109 9.3005
R18570 gnd.n7275 gnd.n125 9.3005
R18571 gnd.n7274 gnd.n126 9.3005
R18572 gnd.n7273 gnd.n127 9.3005
R18573 gnd.n144 gnd.n128 9.3005
R18574 gnd.n7263 gnd.n145 9.3005
R18575 gnd.n7262 gnd.n146 9.3005
R18576 gnd.n7261 gnd.n147 9.3005
R18577 gnd.n162 gnd.n148 9.3005
R18578 gnd.n7251 gnd.n163 9.3005
R18579 gnd.n7250 gnd.n164 9.3005
R18580 gnd.n7249 gnd.n165 9.3005
R18581 gnd.n1508 gnd.n1507 9.3005
R18582 gnd.n7298 gnd.n7297 9.3005
R18583 gnd.n4164 gnd.n4163 9.3005
R18584 gnd.n4168 gnd.n4165 9.3005
R18585 gnd.n4167 gnd.n4166 9.3005
R18586 gnd.n2131 gnd.n2130 9.3005
R18587 gnd.n4223 gnd.n4222 9.3005
R18588 gnd.n4224 gnd.n2129 9.3005
R18589 gnd.n4226 gnd.n4225 9.3005
R18590 gnd.n2127 gnd.n2126 9.3005
R18591 gnd.n4231 gnd.n4230 9.3005
R18592 gnd.n4232 gnd.n2125 9.3005
R18593 gnd.n4234 gnd.n4233 9.3005
R18594 gnd.n2123 gnd.n2122 9.3005
R18595 gnd.n4239 gnd.n4238 9.3005
R18596 gnd.n4240 gnd.n2121 9.3005
R18597 gnd.n4242 gnd.n4241 9.3005
R18598 gnd.n2119 gnd.n2118 9.3005
R18599 gnd.n4247 gnd.n4246 9.3005
R18600 gnd.n4248 gnd.n2117 9.3005
R18601 gnd.n4250 gnd.n4249 9.3005
R18602 gnd.n2115 gnd.n2114 9.3005
R18603 gnd.n4256 gnd.n4255 9.3005
R18604 gnd.n4257 gnd.n2113 9.3005
R18605 gnd.n4259 gnd.n4258 9.3005
R18606 gnd.n2109 gnd.n2108 9.3005
R18607 gnd.n4324 gnd.n4323 9.3005
R18608 gnd.n4325 gnd.n2107 9.3005
R18609 gnd.n4327 gnd.n4326 9.3005
R18610 gnd.n2095 gnd.n2094 9.3005
R18611 gnd.n4340 gnd.n4339 9.3005
R18612 gnd.n4341 gnd.n2093 9.3005
R18613 gnd.n4343 gnd.n4342 9.3005
R18614 gnd.n2080 gnd.n2079 9.3005
R18615 gnd.n4356 gnd.n4355 9.3005
R18616 gnd.n4357 gnd.n2078 9.3005
R18617 gnd.n4359 gnd.n4358 9.3005
R18618 gnd.n2066 gnd.n2065 9.3005
R18619 gnd.n4372 gnd.n4371 9.3005
R18620 gnd.n4373 gnd.n2064 9.3005
R18621 gnd.n4375 gnd.n4374 9.3005
R18622 gnd.n2051 gnd.n2050 9.3005
R18623 gnd.n4402 gnd.n4401 9.3005
R18624 gnd.n4403 gnd.n2049 9.3005
R18625 gnd.n4411 gnd.n4404 9.3005
R18626 gnd.n4410 gnd.n4405 9.3005
R18627 gnd.n4409 gnd.n4407 9.3005
R18628 gnd.n4406 gnd.n1207 9.3005
R18629 gnd.n5775 gnd.n1208 9.3005
R18630 gnd.n5774 gnd.n1209 9.3005
R18631 gnd.n5773 gnd.n1210 9.3005
R18632 gnd.n4560 gnd.n1211 9.3005
R18633 gnd.n4561 gnd.n4559 9.3005
R18634 gnd.n4563 gnd.n4562 9.3005
R18635 gnd.n2021 gnd.n2020 9.3005
R18636 gnd.n4589 gnd.n4588 9.3005
R18637 gnd.n4590 gnd.n2019 9.3005
R18638 gnd.n4594 gnd.n4591 9.3005
R18639 gnd.n4593 gnd.n4592 9.3005
R18640 gnd.n1993 gnd.n1992 9.3005
R18641 gnd.n4627 gnd.n4626 9.3005
R18642 gnd.n4628 gnd.n1991 9.3005
R18643 gnd.n4636 gnd.n4629 9.3005
R18644 gnd.n4635 gnd.n4630 9.3005
R18645 gnd.n4634 gnd.n4632 9.3005
R18646 gnd.n4631 gnd.n1965 9.3005
R18647 gnd.n4697 gnd.n1966 9.3005
R18648 gnd.n4696 gnd.n1967 9.3005
R18649 gnd.n4695 gnd.n1968 9.3005
R18650 gnd.n1943 gnd.n1942 9.3005
R18651 gnd.n4728 gnd.n4727 9.3005
R18652 gnd.n4729 gnd.n1941 9.3005
R18653 gnd.n4733 gnd.n4730 9.3005
R18654 gnd.n4732 gnd.n4731 9.3005
R18655 gnd.n1915 gnd.n1914 9.3005
R18656 gnd.n4766 gnd.n4765 9.3005
R18657 gnd.n4767 gnd.n1913 9.3005
R18658 gnd.n4769 gnd.n4768 9.3005
R18659 gnd.n1889 gnd.n1888 9.3005
R18660 gnd.n4803 gnd.n4802 9.3005
R18661 gnd.n4804 gnd.n1887 9.3005
R18662 gnd.n4808 gnd.n4805 9.3005
R18663 gnd.n4807 gnd.n4806 9.3005
R18664 gnd.n1862 gnd.n1861 9.3005
R18665 gnd.n4852 gnd.n4851 9.3005
R18666 gnd.n4853 gnd.n1860 9.3005
R18667 gnd.n4857 gnd.n4854 9.3005
R18668 gnd.n4856 gnd.n4855 9.3005
R18669 gnd.n1840 gnd.n1839 9.3005
R18670 gnd.n4893 gnd.n4892 9.3005
R18671 gnd.n4894 gnd.n1838 9.3005
R18672 gnd.n4898 gnd.n4895 9.3005
R18673 gnd.n4897 gnd.n4896 9.3005
R18674 gnd.n1810 gnd.n1809 9.3005
R18675 gnd.n4933 gnd.n4932 9.3005
R18676 gnd.n4934 gnd.n1808 9.3005
R18677 gnd.n4936 gnd.n4935 9.3005
R18678 gnd.n1786 gnd.n1785 9.3005
R18679 gnd.n4976 gnd.n4975 9.3005
R18680 gnd.n4977 gnd.n1784 9.3005
R18681 gnd.n4981 gnd.n4978 9.3005
R18682 gnd.n4980 gnd.n4979 9.3005
R18683 gnd.n1730 gnd.n1729 9.3005
R18684 gnd.n5152 gnd.n5151 9.3005
R18685 gnd.n5153 gnd.n1728 9.3005
R18686 gnd.n5155 gnd.n5154 9.3005
R18687 gnd.n1719 gnd.n1718 9.3005
R18688 gnd.n5169 gnd.n5168 9.3005
R18689 gnd.n5170 gnd.n1717 9.3005
R18690 gnd.n5172 gnd.n5171 9.3005
R18691 gnd.n1707 gnd.n1706 9.3005
R18692 gnd.n5186 gnd.n5185 9.3005
R18693 gnd.n5187 gnd.n1705 9.3005
R18694 gnd.n5189 gnd.n5188 9.3005
R18695 gnd.n1695 gnd.n1694 9.3005
R18696 gnd.n5203 gnd.n5202 9.3005
R18697 gnd.n5204 gnd.n1693 9.3005
R18698 gnd.n5206 gnd.n5205 9.3005
R18699 gnd.n1683 gnd.n1682 9.3005
R18700 gnd.n5220 gnd.n5219 9.3005
R18701 gnd.n5221 gnd.n1681 9.3005
R18702 gnd.n5226 gnd.n5222 9.3005
R18703 gnd.n5225 gnd.n5224 9.3005
R18704 gnd.n5223 gnd.n1671 9.3005
R18705 gnd.n5240 gnd.n1670 9.3005
R18706 gnd.n5242 gnd.n5241 9.3005
R18707 gnd.n5243 gnd.n1669 9.3005
R18708 gnd.n5256 gnd.n5244 9.3005
R18709 gnd.n5255 gnd.n5245 9.3005
R18710 gnd.n5254 gnd.n5246 9.3005
R18711 gnd.n5248 gnd.n5247 9.3005
R18712 gnd.n5250 gnd.n5249 9.3005
R18713 gnd.n1635 gnd.n1634 9.3005
R18714 gnd.n5311 gnd.n5310 9.3005
R18715 gnd.n5312 gnd.n1633 9.3005
R18716 gnd.n5314 gnd.n5313 9.3005
R18717 gnd.n1631 gnd.n1630 9.3005
R18718 gnd.n5319 gnd.n5318 9.3005
R18719 gnd.n5320 gnd.n1629 9.3005
R18720 gnd.n5322 gnd.n5321 9.3005
R18721 gnd.n1627 gnd.n1626 9.3005
R18722 gnd.n5327 gnd.n5326 9.3005
R18723 gnd.n5328 gnd.n1625 9.3005
R18724 gnd.n5347 gnd.n5329 9.3005
R18725 gnd.n5346 gnd.n5330 9.3005
R18726 gnd.n5345 gnd.n5331 9.3005
R18727 gnd.n5334 gnd.n5332 9.3005
R18728 gnd.n5341 gnd.n5335 9.3005
R18729 gnd.n6878 gnd.n184 9.3005
R18730 gnd.n4132 gnd.n4131 9.3005
R18731 gnd.n3778 gnd.n3775 9.3005
R18732 gnd.n3777 gnd.n3776 9.3005
R18733 gnd.n2219 gnd.n2218 9.3005
R18734 gnd.n4028 gnd.n4027 9.3005
R18735 gnd.n4029 gnd.n2217 9.3005
R18736 gnd.n4033 gnd.n4030 9.3005
R18737 gnd.n4032 gnd.n4031 9.3005
R18738 gnd.n2194 gnd.n2193 9.3005
R18739 gnd.n4063 gnd.n4062 9.3005
R18740 gnd.n4064 gnd.n2192 9.3005
R18741 gnd.n4070 gnd.n4065 9.3005
R18742 gnd.n4069 gnd.n4066 9.3005
R18743 gnd.n4068 gnd.n4067 9.3005
R18744 gnd.n2168 gnd.n2167 9.3005
R18745 gnd.n4103 gnd.n4102 9.3005
R18746 gnd.n4104 gnd.n2166 9.3005
R18747 gnd.n4106 gnd.n4105 9.3005
R18748 gnd.n2163 gnd.n2162 9.3005
R18749 gnd.n4129 gnd.n4128 9.3005
R18750 gnd.n4130 gnd.n2161 9.3005
R18751 gnd.n3774 gnd.n3706 9.3005
R18752 gnd.n3767 gnd.n3766 9.3005
R18753 gnd.n3765 gnd.n3712 9.3005
R18754 gnd.n3764 gnd.n3763 9.3005
R18755 gnd.n3714 gnd.n3713 9.3005
R18756 gnd.n3757 gnd.n3756 9.3005
R18757 gnd.n3755 gnd.n3716 9.3005
R18758 gnd.n3754 gnd.n3753 9.3005
R18759 gnd.n3718 gnd.n3717 9.3005
R18760 gnd.n3747 gnd.n3746 9.3005
R18761 gnd.n3745 gnd.n3720 9.3005
R18762 gnd.n3744 gnd.n3743 9.3005
R18763 gnd.n3722 gnd.n3721 9.3005
R18764 gnd.n3737 gnd.n3736 9.3005
R18765 gnd.n3735 gnd.n3724 9.3005
R18766 gnd.n3734 gnd.n3733 9.3005
R18767 gnd.n3728 gnd.n3725 9.3005
R18768 gnd.n3727 gnd.n3726 9.3005
R18769 gnd.n3710 gnd.n3707 9.3005
R18770 gnd.n3773 gnd.n3772 9.3005
R18771 gnd.n5853 gnd.n1039 9.3005
R18772 gnd.n5856 gnd.n1038 9.3005
R18773 gnd.n5857 gnd.n1037 9.3005
R18774 gnd.n5860 gnd.n1036 9.3005
R18775 gnd.n5861 gnd.n1035 9.3005
R18776 gnd.n5864 gnd.n1034 9.3005
R18777 gnd.n5865 gnd.n1033 9.3005
R18778 gnd.n5868 gnd.n1032 9.3005
R18779 gnd.n5870 gnd.n1029 9.3005
R18780 gnd.n5873 gnd.n1028 9.3005
R18781 gnd.n5874 gnd.n1027 9.3005
R18782 gnd.n5877 gnd.n1026 9.3005
R18783 gnd.n5878 gnd.n1025 9.3005
R18784 gnd.n5881 gnd.n1024 9.3005
R18785 gnd.n5882 gnd.n1023 9.3005
R18786 gnd.n5885 gnd.n1022 9.3005
R18787 gnd.n5886 gnd.n1021 9.3005
R18788 gnd.n5889 gnd.n1020 9.3005
R18789 gnd.n5890 gnd.n1019 9.3005
R18790 gnd.n5893 gnd.n1018 9.3005
R18791 gnd.n5894 gnd.n1017 9.3005
R18792 gnd.n5897 gnd.n1016 9.3005
R18793 gnd.n5898 gnd.n1015 9.3005
R18794 gnd.n5899 gnd.n1014 9.3005
R18795 gnd.n1013 gnd.n1010 9.3005
R18796 gnd.n1012 gnd.n1011 9.3005
R18797 gnd.n1136 gnd.n1135 9.3005
R18798 gnd.n1132 gnd.n1042 9.3005
R18799 gnd.n1129 gnd.n1043 9.3005
R18800 gnd.n1128 gnd.n1044 9.3005
R18801 gnd.n1125 gnd.n1045 9.3005
R18802 gnd.n1124 gnd.n1046 9.3005
R18803 gnd.n1121 gnd.n1047 9.3005
R18804 gnd.n1120 gnd.n1048 9.3005
R18805 gnd.n1117 gnd.n1116 9.3005
R18806 gnd.n1115 gnd.n1049 9.3005
R18807 gnd.n1114 gnd.n1113 9.3005
R18808 gnd.n1110 gnd.n1052 9.3005
R18809 gnd.n1107 gnd.n1053 9.3005
R18810 gnd.n1106 gnd.n1054 9.3005
R18811 gnd.n1103 gnd.n1055 9.3005
R18812 gnd.n1102 gnd.n1056 9.3005
R18813 gnd.n1099 gnd.n1057 9.3005
R18814 gnd.n1098 gnd.n1058 9.3005
R18815 gnd.n1095 gnd.n1059 9.3005
R18816 gnd.n1094 gnd.n1060 9.3005
R18817 gnd.n1091 gnd.n1061 9.3005
R18818 gnd.n1090 gnd.n1062 9.3005
R18819 gnd.n1087 gnd.n1063 9.3005
R18820 gnd.n1086 gnd.n1064 9.3005
R18821 gnd.n1083 gnd.n1065 9.3005
R18822 gnd.n1082 gnd.n1066 9.3005
R18823 gnd.n1079 gnd.n1067 9.3005
R18824 gnd.n1078 gnd.n1068 9.3005
R18825 gnd.n1075 gnd.n1074 9.3005
R18826 gnd.n1073 gnd.n1070 9.3005
R18827 gnd.n1137 gnd.n1040 9.3005
R18828 gnd.n4001 gnd.n2234 9.3005
R18829 gnd.n4013 gnd.n2235 9.3005
R18830 gnd.n4012 gnd.n2236 9.3005
R18831 gnd.n4011 gnd.n4007 9.3005
R18832 gnd.n4010 gnd.n4008 9.3005
R18833 gnd.n2213 gnd.n2209 9.3005
R18834 gnd.n4048 gnd.n2210 9.3005
R18835 gnd.n4047 gnd.n2211 9.3005
R18836 gnd.n4046 gnd.n4042 9.3005
R18837 gnd.n4045 gnd.n4043 9.3005
R18838 gnd.n2188 gnd.n2183 9.3005
R18839 gnd.n4088 gnd.n2184 9.3005
R18840 gnd.n4087 gnd.n2185 9.3005
R18841 gnd.n4086 gnd.n2186 9.3005
R18842 gnd.n4085 gnd.n4081 9.3005
R18843 gnd.n4083 gnd.n4082 9.3005
R18844 gnd.n2165 gnd.n750 9.3005
R18845 gnd.n6057 gnd.n751 9.3005
R18846 gnd.n6056 gnd.n752 9.3005
R18847 gnd.n6055 gnd.n753 9.3005
R18848 gnd.n2160 gnd.n754 9.3005
R18849 gnd.n6044 gnd.n767 9.3005
R18850 gnd.n6043 gnd.n768 9.3005
R18851 gnd.n6042 gnd.n769 9.3005
R18852 gnd.n4140 gnd.n770 9.3005
R18853 gnd.n6031 gnd.n785 9.3005
R18854 gnd.n6030 gnd.n786 9.3005
R18855 gnd.n6029 gnd.n787 9.3005
R18856 gnd.n2144 gnd.n788 9.3005
R18857 gnd.n6019 gnd.n804 9.3005
R18858 gnd.n6018 gnd.n805 9.3005
R18859 gnd.n6017 gnd.n806 9.3005
R18860 gnd.n4185 gnd.n807 9.3005
R18861 gnd.n6007 gnd.n825 9.3005
R18862 gnd.n6006 gnd.n826 9.3005
R18863 gnd.n6005 gnd.n827 9.3005
R18864 gnd.n4195 gnd.n828 9.3005
R18865 gnd.n5995 gnd.n845 9.3005
R18866 gnd.n5994 gnd.n846 9.3005
R18867 gnd.n5993 gnd.n847 9.3005
R18868 gnd.n864 gnd.n848 9.3005
R18869 gnd.n5983 gnd.n5982 9.3005
R18870 gnd.n4000 gnd.n3999 9.3005
R18871 gnd.n4002 gnd.n4001 9.3005
R18872 gnd.n4003 gnd.n2235 9.3005
R18873 gnd.n4005 gnd.n2236 9.3005
R18874 gnd.n4007 gnd.n4006 9.3005
R18875 gnd.n4008 gnd.n2212 9.3005
R18876 gnd.n4037 gnd.n2213 9.3005
R18877 gnd.n4038 gnd.n2210 9.3005
R18878 gnd.n4040 gnd.n2211 9.3005
R18879 gnd.n4042 gnd.n4041 9.3005
R18880 gnd.n4043 gnd.n2187 9.3005
R18881 gnd.n4074 gnd.n2188 9.3005
R18882 gnd.n4075 gnd.n2184 9.3005
R18883 gnd.n4077 gnd.n2185 9.3005
R18884 gnd.n4078 gnd.n2186 9.3005
R18885 gnd.n4081 gnd.n4080 9.3005
R18886 gnd.n4082 gnd.n2164 9.3005
R18887 gnd.n4110 gnd.n2165 9.3005
R18888 gnd.n4111 gnd.n751 9.3005
R18889 gnd.n4112 gnd.n752 9.3005
R18890 gnd.n2159 gnd.n753 9.3005
R18891 gnd.n4136 gnd.n2160 9.3005
R18892 gnd.n4137 gnd.n767 9.3005
R18893 gnd.n4138 gnd.n768 9.3005
R18894 gnd.n4139 gnd.n769 9.3005
R18895 gnd.n4143 gnd.n4140 9.3005
R18896 gnd.n4142 gnd.n785 9.3005
R18897 gnd.n4141 gnd.n786 9.3005
R18898 gnd.n2143 gnd.n787 9.3005
R18899 gnd.n4181 gnd.n2144 9.3005
R18900 gnd.n4182 gnd.n804 9.3005
R18901 gnd.n4183 gnd.n805 9.3005
R18902 gnd.n4184 gnd.n806 9.3005
R18903 gnd.n4188 gnd.n4185 9.3005
R18904 gnd.n4189 gnd.n825 9.3005
R18905 gnd.n4193 gnd.n826 9.3005
R18906 gnd.n4194 gnd.n827 9.3005
R18907 gnd.n4198 gnd.n4195 9.3005
R18908 gnd.n4199 gnd.n845 9.3005
R18909 gnd.n4200 gnd.n846 9.3005
R18910 gnd.n866 gnd.n847 9.3005
R18911 gnd.n5980 gnd.n864 9.3005
R18912 gnd.n5982 gnd.n5981 9.3005
R18913 gnd.n4000 gnd.n2237 9.3005
R18914 gnd.n3874 gnd.n3873 9.3005
R18915 gnd.n3882 gnd.n3870 9.3005
R18916 gnd.n3883 gnd.n3869 9.3005
R18917 gnd.n3884 gnd.n3868 9.3005
R18918 gnd.n3867 gnd.n3865 9.3005
R18919 gnd.n3890 gnd.n3864 9.3005
R18920 gnd.n3891 gnd.n3863 9.3005
R18921 gnd.n3892 gnd.n3862 9.3005
R18922 gnd.n3861 gnd.n3859 9.3005
R18923 gnd.n3898 gnd.n3858 9.3005
R18924 gnd.n3899 gnd.n3857 9.3005
R18925 gnd.n3900 gnd.n3856 9.3005
R18926 gnd.n3855 gnd.n3853 9.3005
R18927 gnd.n3906 gnd.n3852 9.3005
R18928 gnd.n3907 gnd.n3851 9.3005
R18929 gnd.n3908 gnd.n3850 9.3005
R18930 gnd.n3849 gnd.n3847 9.3005
R18931 gnd.n3914 gnd.n3846 9.3005
R18932 gnd.n3915 gnd.n3845 9.3005
R18933 gnd.n3916 gnd.n3844 9.3005
R18934 gnd.n3922 gnd.n3838 9.3005
R18935 gnd.n3923 gnd.n3837 9.3005
R18936 gnd.n3924 gnd.n3836 9.3005
R18937 gnd.n3835 gnd.n3833 9.3005
R18938 gnd.n3930 gnd.n3832 9.3005
R18939 gnd.n3931 gnd.n3831 9.3005
R18940 gnd.n3932 gnd.n3830 9.3005
R18941 gnd.n3829 gnd.n3827 9.3005
R18942 gnd.n3938 gnd.n3826 9.3005
R18943 gnd.n3939 gnd.n3825 9.3005
R18944 gnd.n3940 gnd.n3824 9.3005
R18945 gnd.n3823 gnd.n3821 9.3005
R18946 gnd.n3946 gnd.n3820 9.3005
R18947 gnd.n3947 gnd.n3819 9.3005
R18948 gnd.n3948 gnd.n3818 9.3005
R18949 gnd.n3817 gnd.n3815 9.3005
R18950 gnd.n3954 gnd.n3814 9.3005
R18951 gnd.n3955 gnd.n3813 9.3005
R18952 gnd.n3956 gnd.n3812 9.3005
R18953 gnd.n3811 gnd.n3806 9.3005
R18954 gnd.n3962 gnd.n3805 9.3005
R18955 gnd.n3963 gnd.n3804 9.3005
R18956 gnd.n3964 gnd.n3803 9.3005
R18957 gnd.n3802 gnd.n3800 9.3005
R18958 gnd.n3970 gnd.n3799 9.3005
R18959 gnd.n3971 gnd.n3798 9.3005
R18960 gnd.n3972 gnd.n3797 9.3005
R18961 gnd.n3796 gnd.n3794 9.3005
R18962 gnd.n3978 gnd.n3793 9.3005
R18963 gnd.n3979 gnd.n3792 9.3005
R18964 gnd.n3980 gnd.n3791 9.3005
R18965 gnd.n3790 gnd.n3788 9.3005
R18966 gnd.n3985 gnd.n3787 9.3005
R18967 gnd.n3986 gnd.n3786 9.3005
R18968 gnd.n3785 gnd.n3783 9.3005
R18969 gnd.n3991 gnd.n3782 9.3005
R18970 gnd.n3993 gnd.n3992 9.3005
R18971 gnd.n3843 gnd.n3841 9.3005
R18972 gnd.n3876 gnd.n3875 9.3005
R18973 gnd.n2228 gnd.n2227 9.3005
R18974 gnd.n4018 gnd.n4017 9.3005
R18975 gnd.n4019 gnd.n2226 9.3005
R18976 gnd.n4023 gnd.n4020 9.3005
R18977 gnd.n4022 gnd.n4021 9.3005
R18978 gnd.n2203 gnd.n2202 9.3005
R18979 gnd.n4053 gnd.n4052 9.3005
R18980 gnd.n4054 gnd.n2201 9.3005
R18981 gnd.n4058 gnd.n4055 9.3005
R18982 gnd.n4057 gnd.n4056 9.3005
R18983 gnd.n2176 gnd.n2175 9.3005
R18984 gnd.n4093 gnd.n4092 9.3005
R18985 gnd.n4094 gnd.n2174 9.3005
R18986 gnd.n4097 gnd.n4096 9.3005
R18987 gnd.n4095 gnd.n740 9.3005
R18988 gnd.n794 gnd.n778 9.3005
R18989 gnd.n6025 gnd.n795 9.3005
R18990 gnd.n6024 gnd.n796 9.3005
R18991 gnd.n6023 gnd.n797 9.3005
R18992 gnd.n814 gnd.n798 9.3005
R18993 gnd.n6013 gnd.n815 9.3005
R18994 gnd.n6012 gnd.n816 9.3005
R18995 gnd.n6011 gnd.n817 9.3005
R18996 gnd.n834 gnd.n818 9.3005
R18997 gnd.n6001 gnd.n835 9.3005
R18998 gnd.n6000 gnd.n836 9.3005
R18999 gnd.n5999 gnd.n837 9.3005
R19000 gnd.n854 gnd.n838 9.3005
R19001 gnd.n5989 gnd.n855 9.3005
R19002 gnd.n5988 gnd.n856 9.3005
R19003 gnd.n5987 gnd.n857 9.3005
R19004 gnd.n3995 gnd.n3994 9.3005
R19005 gnd.n6035 gnd.n741 9.3005
R19006 gnd.n6070 gnd.n6069 9.3005
R19007 gnd.n6073 gnd.n729 9.3005
R19008 gnd.n728 gnd.n724 9.3005
R19009 gnd.n6079 gnd.n723 9.3005
R19010 gnd.n6080 gnd.n722 9.3005
R19011 gnd.n6081 gnd.n721 9.3005
R19012 gnd.n720 gnd.n716 9.3005
R19013 gnd.n6087 gnd.n715 9.3005
R19014 gnd.n6088 gnd.n714 9.3005
R19015 gnd.n6089 gnd.n713 9.3005
R19016 gnd.n712 gnd.n708 9.3005
R19017 gnd.n6095 gnd.n707 9.3005
R19018 gnd.n6096 gnd.n706 9.3005
R19019 gnd.n6097 gnd.n705 9.3005
R19020 gnd.n704 gnd.n700 9.3005
R19021 gnd.n6103 gnd.n699 9.3005
R19022 gnd.n6104 gnd.n698 9.3005
R19023 gnd.n6105 gnd.n697 9.3005
R19024 gnd.n696 gnd.n692 9.3005
R19025 gnd.n6111 gnd.n691 9.3005
R19026 gnd.n6112 gnd.n690 9.3005
R19027 gnd.n6113 gnd.n689 9.3005
R19028 gnd.n688 gnd.n684 9.3005
R19029 gnd.n6119 gnd.n683 9.3005
R19030 gnd.n6120 gnd.n682 9.3005
R19031 gnd.n6121 gnd.n681 9.3005
R19032 gnd.n680 gnd.n676 9.3005
R19033 gnd.n6127 gnd.n675 9.3005
R19034 gnd.n6128 gnd.n674 9.3005
R19035 gnd.n6129 gnd.n673 9.3005
R19036 gnd.n672 gnd.n668 9.3005
R19037 gnd.n6135 gnd.n667 9.3005
R19038 gnd.n6136 gnd.n666 9.3005
R19039 gnd.n6137 gnd.n665 9.3005
R19040 gnd.n664 gnd.n660 9.3005
R19041 gnd.n6143 gnd.n659 9.3005
R19042 gnd.n6144 gnd.n658 9.3005
R19043 gnd.n6145 gnd.n657 9.3005
R19044 gnd.n656 gnd.n652 9.3005
R19045 gnd.n6151 gnd.n651 9.3005
R19046 gnd.n6152 gnd.n650 9.3005
R19047 gnd.n6153 gnd.n649 9.3005
R19048 gnd.n648 gnd.n644 9.3005
R19049 gnd.n6159 gnd.n643 9.3005
R19050 gnd.n6160 gnd.n642 9.3005
R19051 gnd.n6161 gnd.n641 9.3005
R19052 gnd.n640 gnd.n636 9.3005
R19053 gnd.n6167 gnd.n635 9.3005
R19054 gnd.n6168 gnd.n634 9.3005
R19055 gnd.n6169 gnd.n633 9.3005
R19056 gnd.n632 gnd.n628 9.3005
R19057 gnd.n6175 gnd.n627 9.3005
R19058 gnd.n6176 gnd.n626 9.3005
R19059 gnd.n6177 gnd.n625 9.3005
R19060 gnd.n624 gnd.n620 9.3005
R19061 gnd.n6183 gnd.n619 9.3005
R19062 gnd.n6184 gnd.n618 9.3005
R19063 gnd.n6185 gnd.n617 9.3005
R19064 gnd.n616 gnd.n612 9.3005
R19065 gnd.n6191 gnd.n611 9.3005
R19066 gnd.n6192 gnd.n610 9.3005
R19067 gnd.n6193 gnd.n609 9.3005
R19068 gnd.n608 gnd.n604 9.3005
R19069 gnd.n6199 gnd.n603 9.3005
R19070 gnd.n6200 gnd.n602 9.3005
R19071 gnd.n6201 gnd.n601 9.3005
R19072 gnd.n600 gnd.n596 9.3005
R19073 gnd.n6207 gnd.n595 9.3005
R19074 gnd.n6208 gnd.n594 9.3005
R19075 gnd.n6209 gnd.n593 9.3005
R19076 gnd.n592 gnd.n588 9.3005
R19077 gnd.n6215 gnd.n587 9.3005
R19078 gnd.n6216 gnd.n586 9.3005
R19079 gnd.n6217 gnd.n585 9.3005
R19080 gnd.n584 gnd.n580 9.3005
R19081 gnd.n6223 gnd.n579 9.3005
R19082 gnd.n6224 gnd.n578 9.3005
R19083 gnd.n6225 gnd.n577 9.3005
R19084 gnd.n576 gnd.n572 9.3005
R19085 gnd.n6231 gnd.n571 9.3005
R19086 gnd.n6232 gnd.n570 9.3005
R19087 gnd.n6233 gnd.n569 9.3005
R19088 gnd.n568 gnd.n564 9.3005
R19089 gnd.n6239 gnd.n563 9.3005
R19090 gnd.n6241 gnd.n6240 9.3005
R19091 gnd.n6072 gnd.n6071 9.3005
R19092 gnd.n5262 gnd.n1639 9.3005
R19093 gnd.n4317 gnd.n4314 9.3005
R19094 gnd.n4319 gnd.n4318 9.3005
R19095 gnd.n2102 gnd.n2101 9.3005
R19096 gnd.n4332 gnd.n4331 9.3005
R19097 gnd.n4333 gnd.n2100 9.3005
R19098 gnd.n4335 gnd.n4334 9.3005
R19099 gnd.n2088 gnd.n2087 9.3005
R19100 gnd.n4348 gnd.n4347 9.3005
R19101 gnd.n4349 gnd.n2086 9.3005
R19102 gnd.n4351 gnd.n4350 9.3005
R19103 gnd.n2074 gnd.n2073 9.3005
R19104 gnd.n4364 gnd.n4363 9.3005
R19105 gnd.n4365 gnd.n2072 9.3005
R19106 gnd.n4367 gnd.n4366 9.3005
R19107 gnd.n2060 gnd.n2059 9.3005
R19108 gnd.n4380 gnd.n4379 9.3005
R19109 gnd.n4381 gnd.n2057 9.3005
R19110 gnd.n4397 gnd.n4396 9.3005
R19111 gnd.n4395 gnd.n2058 9.3005
R19112 gnd.n4394 gnd.n4393 9.3005
R19113 gnd.n4392 gnd.n4382 9.3005
R19114 gnd.n4391 gnd.n4390 9.3005
R19115 gnd.n4389 gnd.n4386 9.3005
R19116 gnd.n4388 gnd.n4387 9.3005
R19117 gnd.n1218 gnd.n1216 9.3005
R19118 gnd.n5769 gnd.n5768 9.3005
R19119 gnd.n5767 gnd.n1217 9.3005
R19120 gnd.n5766 gnd.n5765 9.3005
R19121 gnd.n5764 gnd.n1219 9.3005
R19122 gnd.n5763 gnd.n5762 9.3005
R19123 gnd.n5761 gnd.n1223 9.3005
R19124 gnd.n5760 gnd.n5759 9.3005
R19125 gnd.n5758 gnd.n1224 9.3005
R19126 gnd.n5757 gnd.n5756 9.3005
R19127 gnd.n5755 gnd.n1228 9.3005
R19128 gnd.n5754 gnd.n5753 9.3005
R19129 gnd.n5752 gnd.n1229 9.3005
R19130 gnd.n5751 gnd.n5750 9.3005
R19131 gnd.n5749 gnd.n1233 9.3005
R19132 gnd.n5748 gnd.n5747 9.3005
R19133 gnd.n5746 gnd.n1234 9.3005
R19134 gnd.n5745 gnd.n5744 9.3005
R19135 gnd.n5743 gnd.n1238 9.3005
R19136 gnd.n5742 gnd.n5741 9.3005
R19137 gnd.n5740 gnd.n1239 9.3005
R19138 gnd.n5739 gnd.n5738 9.3005
R19139 gnd.n5737 gnd.n1243 9.3005
R19140 gnd.n5736 gnd.n5735 9.3005
R19141 gnd.n5734 gnd.n1244 9.3005
R19142 gnd.n5733 gnd.n5732 9.3005
R19143 gnd.n5731 gnd.n1248 9.3005
R19144 gnd.n5730 gnd.n5729 9.3005
R19145 gnd.n5728 gnd.n1249 9.3005
R19146 gnd.n5727 gnd.n5726 9.3005
R19147 gnd.n5725 gnd.n1253 9.3005
R19148 gnd.n5724 gnd.n5723 9.3005
R19149 gnd.n5722 gnd.n1254 9.3005
R19150 gnd.n5721 gnd.n5720 9.3005
R19151 gnd.n5719 gnd.n1258 9.3005
R19152 gnd.n5718 gnd.n5717 9.3005
R19153 gnd.n5716 gnd.n1259 9.3005
R19154 gnd.n5715 gnd.n5714 9.3005
R19155 gnd.n5713 gnd.n1263 9.3005
R19156 gnd.n5712 gnd.n5711 9.3005
R19157 gnd.n5710 gnd.n1264 9.3005
R19158 gnd.n5709 gnd.n5708 9.3005
R19159 gnd.n5707 gnd.n1268 9.3005
R19160 gnd.n5706 gnd.n5705 9.3005
R19161 gnd.n5704 gnd.n1269 9.3005
R19162 gnd.n5703 gnd.n5702 9.3005
R19163 gnd.n5701 gnd.n1273 9.3005
R19164 gnd.n5700 gnd.n5699 9.3005
R19165 gnd.n5698 gnd.n1274 9.3005
R19166 gnd.n5697 gnd.n5696 9.3005
R19167 gnd.n5695 gnd.n1278 9.3005
R19168 gnd.n5694 gnd.n5693 9.3005
R19169 gnd.n5692 gnd.n1279 9.3005
R19170 gnd.n5691 gnd.n5690 9.3005
R19171 gnd.n5689 gnd.n1283 9.3005
R19172 gnd.n5688 gnd.n5687 9.3005
R19173 gnd.n5686 gnd.n1284 9.3005
R19174 gnd.n5685 gnd.n5684 9.3005
R19175 gnd.n5683 gnd.n1288 9.3005
R19176 gnd.n5682 gnd.n5681 9.3005
R19177 gnd.n5680 gnd.n1289 9.3005
R19178 gnd.n5679 gnd.n5678 9.3005
R19179 gnd.n5677 gnd.n1293 9.3005
R19180 gnd.n5676 gnd.n5675 9.3005
R19181 gnd.n5674 gnd.n1294 9.3005
R19182 gnd.n5673 gnd.n5672 9.3005
R19183 gnd.n5671 gnd.n1298 9.3005
R19184 gnd.n5670 gnd.n5669 9.3005
R19185 gnd.n5668 gnd.n1299 9.3005
R19186 gnd.n5667 gnd.n5666 9.3005
R19187 gnd.n5665 gnd.n1303 9.3005
R19188 gnd.n5664 gnd.n5663 9.3005
R19189 gnd.n5662 gnd.n1304 9.3005
R19190 gnd.n5661 gnd.n5660 9.3005
R19191 gnd.n5659 gnd.n1308 9.3005
R19192 gnd.n5658 gnd.n5657 9.3005
R19193 gnd.n5656 gnd.n1309 9.3005
R19194 gnd.n4316 gnd.n4315 9.3005
R19195 gnd.n5970 gnd.n871 9.3005
R19196 gnd.n2158 gnd.n2156 9.3005
R19197 gnd.n4151 gnd.n4150 9.3005
R19198 gnd.n4149 gnd.n2157 9.3005
R19199 gnd.n4148 gnd.n4147 9.3005
R19200 gnd.n2147 gnd.n2146 9.3005
R19201 gnd.n4174 gnd.n4173 9.3005
R19202 gnd.n4175 gnd.n2145 9.3005
R19203 gnd.n4177 gnd.n4176 9.3005
R19204 gnd.n2136 gnd.n2134 9.3005
R19205 gnd.n4217 gnd.n4216 9.3005
R19206 gnd.n4215 gnd.n2135 9.3005
R19207 gnd.n4214 gnd.n4213 9.3005
R19208 gnd.n4212 gnd.n2137 9.3005
R19209 gnd.n4211 gnd.n4210 9.3005
R19210 gnd.n4209 gnd.n2140 9.3005
R19211 gnd.n4208 gnd.n4207 9.3005
R19212 gnd.n4206 gnd.n2141 9.3005
R19213 gnd.n4205 gnd.n4204 9.3005
R19214 gnd.n870 gnd.n868 9.3005
R19215 gnd.n5976 gnd.n5975 9.3005
R19216 gnd.n5974 gnd.n869 9.3005
R19217 gnd.n5948 gnd.n5947 9.3005
R19218 gnd.n5946 gnd.n5945 9.3005
R19219 gnd.n913 gnd.n912 9.3005
R19220 gnd.n5940 gnd.n5939 9.3005
R19221 gnd.n5938 gnd.n5937 9.3005
R19222 gnd.n923 gnd.n922 9.3005
R19223 gnd.n5932 gnd.n5931 9.3005
R19224 gnd.n5930 gnd.n5929 9.3005
R19225 gnd.n931 gnd.n930 9.3005
R19226 gnd.n5924 gnd.n5923 9.3005
R19227 gnd.n5922 gnd.n5921 9.3005
R19228 gnd.n941 gnd.n940 9.3005
R19229 gnd.n5916 gnd.n5915 9.3005
R19230 gnd.n5914 gnd.n5913 9.3005
R19231 gnd.n949 gnd.n948 9.3005
R19232 gnd.n5908 gnd.n5907 9.3005
R19233 gnd.n5906 gnd.n963 9.3005
R19234 gnd.n5905 gnd.n872 9.3005
R19235 gnd.n909 gnd.n907 9.3005
R19236 gnd.n5972 gnd.n5971 9.3005
R19237 gnd.n962 gnd.n873 9.3005
R19238 gnd.n958 gnd.n957 9.3005
R19239 gnd.n5910 gnd.n5909 9.3005
R19240 gnd.n5912 gnd.n5911 9.3005
R19241 gnd.n945 gnd.n944 9.3005
R19242 gnd.n5918 gnd.n5917 9.3005
R19243 gnd.n5920 gnd.n5919 9.3005
R19244 gnd.n937 gnd.n936 9.3005
R19245 gnd.n5926 gnd.n5925 9.3005
R19246 gnd.n5928 gnd.n5927 9.3005
R19247 gnd.n927 gnd.n926 9.3005
R19248 gnd.n5934 gnd.n5933 9.3005
R19249 gnd.n5936 gnd.n5935 9.3005
R19250 gnd.n919 gnd.n918 9.3005
R19251 gnd.n5942 gnd.n5941 9.3005
R19252 gnd.n5944 gnd.n5943 9.3005
R19253 gnd.n908 gnd.n906 9.3005
R19254 gnd.n5950 gnd.n5949 9.3005
R19255 gnd.n5951 gnd.n901 9.3005
R19256 gnd.n5953 gnd.n5952 9.3005
R19257 gnd.n5955 gnd.n900 9.3005
R19258 gnd.n5957 gnd.n5956 9.3005
R19259 gnd.n5958 gnd.n896 9.3005
R19260 gnd.n5960 gnd.n5959 9.3005
R19261 gnd.n5961 gnd.n895 9.3005
R19262 gnd.n5963 gnd.n5962 9.3005
R19263 gnd.n5964 gnd.n894 9.3005
R19264 gnd.n4310 gnd.n4309 9.3005
R19265 gnd.n4308 gnd.n4263 9.3005
R19266 gnd.n4307 gnd.n4306 9.3005
R19267 gnd.n4305 gnd.n4265 9.3005
R19268 gnd.n4304 gnd.n4303 9.3005
R19269 gnd.n4302 gnd.n4268 9.3005
R19270 gnd.n4301 gnd.n4300 9.3005
R19271 gnd.n4299 gnd.n4269 9.3005
R19272 gnd.n4298 gnd.n4297 9.3005
R19273 gnd.n4296 gnd.n4272 9.3005
R19274 gnd.n4295 gnd.n4294 9.3005
R19275 gnd.n4293 gnd.n4273 9.3005
R19276 gnd.n4292 gnd.n4291 9.3005
R19277 gnd.n4290 gnd.n4276 9.3005
R19278 gnd.n4289 gnd.n4288 9.3005
R19279 gnd.n4287 gnd.n4277 9.3005
R19280 gnd.n4286 gnd.n4285 9.3005
R19281 gnd.n4284 gnd.n4280 9.3005
R19282 gnd.n4283 gnd.n4282 9.3005
R19283 gnd.n4281 gnd.n2044 9.3005
R19284 gnd.n2042 gnd.n2041 9.3005
R19285 gnd.n4419 gnd.n4418 9.3005
R19286 gnd.n4420 gnd.n2040 9.3005
R19287 gnd.n4422 gnd.n4421 9.3005
R19288 gnd.n4523 gnd.n2039 9.3005
R19289 gnd.n4525 gnd.n4524 9.3005
R19290 gnd.n4526 gnd.n2037 9.3005
R19291 gnd.n4555 gnd.n4554 9.3005
R19292 gnd.n4553 gnd.n2038 9.3005
R19293 gnd.n4552 gnd.n4551 9.3005
R19294 gnd.n4550 gnd.n4527 9.3005
R19295 gnd.n4549 gnd.n4548 9.3005
R19296 gnd.n4547 gnd.n4529 9.3005
R19297 gnd.n4546 gnd.n4545 9.3005
R19298 gnd.n4544 gnd.n4530 9.3005
R19299 gnd.n4543 gnd.n4542 9.3005
R19300 gnd.n4541 gnd.n4534 9.3005
R19301 gnd.n4540 gnd.n4539 9.3005
R19302 gnd.n4538 gnd.n4536 9.3005
R19303 gnd.n4535 gnd.n1975 9.3005
R19304 gnd.n4660 gnd.n1974 9.3005
R19305 gnd.n4662 gnd.n4661 9.3005
R19306 gnd.n4663 gnd.n1972 9.3005
R19307 gnd.n4691 gnd.n4690 9.3005
R19308 gnd.n4689 gnd.n1973 9.3005
R19309 gnd.n4688 gnd.n4687 9.3005
R19310 gnd.n4686 gnd.n4664 9.3005
R19311 gnd.n4685 gnd.n4684 9.3005
R19312 gnd.n4683 gnd.n4666 9.3005
R19313 gnd.n4682 gnd.n4681 9.3005
R19314 gnd.n4680 gnd.n4667 9.3005
R19315 gnd.n4679 gnd.n4678 9.3005
R19316 gnd.n4677 gnd.n4671 9.3005
R19317 gnd.n4676 gnd.n4675 9.3005
R19318 gnd.n4674 gnd.n4672 9.3005
R19319 gnd.n1882 gnd.n1881 9.3005
R19320 gnd.n4813 gnd.n4812 9.3005
R19321 gnd.n4814 gnd.n1879 9.3005
R19322 gnd.n4817 gnd.n4816 9.3005
R19323 gnd.n4815 gnd.n1880 9.3005
R19324 gnd.n1855 gnd.n1854 9.3005
R19325 gnd.n4862 gnd.n4861 9.3005
R19326 gnd.n4863 gnd.n1852 9.3005
R19327 gnd.n4881 gnd.n4880 9.3005
R19328 gnd.n4879 gnd.n1853 9.3005
R19329 gnd.n4878 gnd.n4877 9.3005
R19330 gnd.n4876 gnd.n4864 9.3005
R19331 gnd.n4875 gnd.n4874 9.3005
R19332 gnd.n4873 gnd.n4868 9.3005
R19333 gnd.n4872 gnd.n4871 9.3005
R19334 gnd.n4870 gnd.n4869 9.3005
R19335 gnd.n1803 gnd.n1802 9.3005
R19336 gnd.n4942 gnd.n4941 9.3005
R19337 gnd.n4943 gnd.n1800 9.3005
R19338 gnd.n4955 gnd.n4954 9.3005
R19339 gnd.n4953 gnd.n1801 9.3005
R19340 gnd.n4952 gnd.n4951 9.3005
R19341 gnd.n4950 gnd.n4944 9.3005
R19342 gnd.n4949 gnd.n4948 9.3005
R19343 gnd.n1725 gnd.n1724 9.3005
R19344 gnd.n5160 gnd.n5159 9.3005
R19345 gnd.n5161 gnd.n1723 9.3005
R19346 gnd.n5163 gnd.n5162 9.3005
R19347 gnd.n1713 gnd.n1712 9.3005
R19348 gnd.n5177 gnd.n5176 9.3005
R19349 gnd.n5178 gnd.n1711 9.3005
R19350 gnd.n5180 gnd.n5179 9.3005
R19351 gnd.n1701 gnd.n1700 9.3005
R19352 gnd.n5194 gnd.n5193 9.3005
R19353 gnd.n5195 gnd.n1699 9.3005
R19354 gnd.n5197 gnd.n5196 9.3005
R19355 gnd.n1688 gnd.n1687 9.3005
R19356 gnd.n5211 gnd.n5210 9.3005
R19357 gnd.n5212 gnd.n1686 9.3005
R19358 gnd.n5214 gnd.n5213 9.3005
R19359 gnd.n1677 gnd.n1676 9.3005
R19360 gnd.n5231 gnd.n5230 9.3005
R19361 gnd.n5232 gnd.n1675 9.3005
R19362 gnd.n5234 gnd.n5233 9.3005
R19363 gnd.n1318 gnd.n1317 9.3005
R19364 gnd.n5652 gnd.n5651 9.3005
R19365 gnd.n4264 gnd.n4262 9.3005
R19366 gnd.n5648 gnd.n1319 9.3005
R19367 gnd.n5647 gnd.n5646 9.3005
R19368 gnd.n5645 gnd.n1322 9.3005
R19369 gnd.n5644 gnd.n5643 9.3005
R19370 gnd.n5642 gnd.n1323 9.3005
R19371 gnd.n5641 gnd.n5640 9.3005
R19372 gnd.n5650 gnd.n5649 9.3005
R19373 gnd.n5593 gnd.n5592 9.3005
R19374 gnd.n1370 gnd.n1369 9.3005
R19375 gnd.n5599 gnd.n5598 9.3005
R19376 gnd.n5601 gnd.n5600 9.3005
R19377 gnd.n1362 gnd.n1361 9.3005
R19378 gnd.n5607 gnd.n5606 9.3005
R19379 gnd.n5609 gnd.n5608 9.3005
R19380 gnd.n1354 gnd.n1353 9.3005
R19381 gnd.n5615 gnd.n5614 9.3005
R19382 gnd.n5617 gnd.n5616 9.3005
R19383 gnd.n1346 gnd.n1345 9.3005
R19384 gnd.n5623 gnd.n5622 9.3005
R19385 gnd.n5625 gnd.n5624 9.3005
R19386 gnd.n1338 gnd.n1337 9.3005
R19387 gnd.n5631 gnd.n5630 9.3005
R19388 gnd.n5633 gnd.n5632 9.3005
R19389 gnd.n1334 gnd.n1329 9.3005
R19390 gnd.n5591 gnd.n1379 9.3005
R19391 gnd.n1640 gnd.n1378 9.3005
R19392 gnd.n5638 gnd.n1327 9.3005
R19393 gnd.n5637 gnd.n5636 9.3005
R19394 gnd.n5635 gnd.n5634 9.3005
R19395 gnd.n1333 gnd.n1332 9.3005
R19396 gnd.n5629 gnd.n5628 9.3005
R19397 gnd.n5627 gnd.n5626 9.3005
R19398 gnd.n1342 gnd.n1341 9.3005
R19399 gnd.n5621 gnd.n5620 9.3005
R19400 gnd.n5619 gnd.n5618 9.3005
R19401 gnd.n1350 gnd.n1349 9.3005
R19402 gnd.n5613 gnd.n5612 9.3005
R19403 gnd.n5611 gnd.n5610 9.3005
R19404 gnd.n1358 gnd.n1357 9.3005
R19405 gnd.n5605 gnd.n5604 9.3005
R19406 gnd.n5603 gnd.n5602 9.3005
R19407 gnd.n1366 gnd.n1365 9.3005
R19408 gnd.n5597 gnd.n5596 9.3005
R19409 gnd.n5595 gnd.n5594 9.3005
R19410 gnd.n1663 gnd.n1376 9.3005
R19411 gnd.n1642 gnd.n1641 9.3005
R19412 gnd.n5264 gnd.n5263 9.3005
R19413 gnd.n5305 gnd.n5304 9.3005
R19414 gnd.n5303 gnd.n1638 9.3005
R19415 gnd.n5302 gnd.n5301 9.3005
R19416 gnd.n5300 gnd.n5267 9.3005
R19417 gnd.n5299 gnd.n5298 9.3005
R19418 gnd.n5297 gnd.n5271 9.3005
R19419 gnd.n5296 gnd.n5295 9.3005
R19420 gnd.n5294 gnd.n5272 9.3005
R19421 gnd.n5293 gnd.n5292 9.3005
R19422 gnd.n1621 gnd.n1620 9.3005
R19423 gnd.n5353 gnd.n5352 9.3005
R19424 gnd.n5354 gnd.n1619 9.3005
R19425 gnd.n5356 gnd.n5355 9.3005
R19426 gnd.n1616 gnd.n1615 9.3005
R19427 gnd.n5368 gnd.n5367 9.3005
R19428 gnd.n5369 gnd.n1613 9.3005
R19429 gnd.n5375 gnd.n5374 9.3005
R19430 gnd.n5373 gnd.n1614 9.3005
R19431 gnd.n5372 gnd.n5371 9.3005
R19432 gnd.n5370 gnd.n67 9.3005
R19433 gnd.n5266 gnd.n1637 9.3005
R19434 gnd.n7308 gnd.n68 9.3005
R19435 gnd.t282 gnd.n2431 9.24152
R19436 gnd.n2333 gnd.t35 9.24152
R19437 gnd.n3601 gnd.t133 9.24152
R19438 gnd.n4220 gnd.t211 9.24152
R19439 gnd.n5349 gnd.t174 9.24152
R19440 gnd.t11 gnd.t282 8.92286
R19441 gnd.n4557 gnd.n2035 8.92286
R19442 gnd.n4651 gnd.n1983 8.92286
R19443 gnd.n4718 gnd.n4717 8.92286
R19444 gnd.n4725 gnd.t304 8.92286
R19445 gnd.n4800 gnd.t310 8.92286
R19446 gnd.n4783 gnd.n1894 8.92286
R19447 gnd.n4859 gnd.n1857 8.92286
R19448 gnd.n4966 gnd.n1794 8.92286
R19449 gnd.n3571 gnd.n3546 8.92171
R19450 gnd.n3539 gnd.n3514 8.92171
R19451 gnd.n3507 gnd.n3482 8.92171
R19452 gnd.n3476 gnd.n3451 8.92171
R19453 gnd.n3444 gnd.n3419 8.92171
R19454 gnd.n3412 gnd.n3387 8.92171
R19455 gnd.n3380 gnd.n3355 8.92171
R19456 gnd.n3349 gnd.n3324 8.92171
R19457 gnd.n5005 gnd.n4987 8.72777
R19458 gnd.n3075 gnd.t284 8.60421
R19459 gnd.n4154 gnd.t160 8.60421
R19460 gnd.n5403 gnd.t190 8.60421
R19461 gnd.n2495 gnd.n2483 8.43656
R19462 gnd.n42 gnd.n30 8.43656
R19463 gnd.n5777 gnd.t93 8.28555
R19464 gnd.n2016 gnd.t314 8.28555
R19465 gnd.n4639 gnd.t313 8.28555
R19466 gnd.n1970 gnd.t0 8.28555
R19467 gnd.t13 gnd.n4790 8.28555
R19468 gnd.n4841 gnd.t309 8.28555
R19469 gnd.n4907 gnd.t299 8.28555
R19470 gnd.n3572 gnd.n3544 8.14595
R19471 gnd.n3540 gnd.n3512 8.14595
R19472 gnd.n3508 gnd.n3480 8.14595
R19473 gnd.n3477 gnd.n3449 8.14595
R19474 gnd.n3445 gnd.n3417 8.14595
R19475 gnd.n3413 gnd.n3385 8.14595
R19476 gnd.n3381 gnd.n3353 8.14595
R19477 gnd.n3350 gnd.n3322 8.14595
R19478 gnd.n4131 gnd.n0 8.10675
R19479 gnd.n7309 gnd.n7308 8.10675
R19480 gnd.n3577 gnd.n3576 7.97301
R19481 gnd.t272 gnd.n2590 7.9669
R19482 gnd.n5967 gnd.n876 7.9669
R19483 gnd.n5259 gnd.n5258 7.9669
R19484 gnd.n7309 gnd.n66 7.78567
R19485 gnd.n5591 gnd.n1378 7.75808
R19486 gnd.n5906 gnd.n5905 7.75808
R19487 gnd.n7189 gnd.n6914 7.75808
R19488 gnd.n3772 gnd.n3710 7.75808
R19489 gnd.t5 gnd.n726 7.64824
R19490 gnd.n4502 gnd.t49 7.64824
R19491 gnd.n4578 gnd.n4577 7.64824
R19492 gnd.n4607 gnd.n1997 7.64824
R19493 gnd.n1947 gnd.n1935 7.64824
R19494 gnd.n4778 gnd.n1905 7.64824
R19495 gnd.n4884 gnd.n4883 7.64824
R19496 gnd.n4913 gnd.n1816 7.64824
R19497 gnd.n2520 gnd.n2519 7.53171
R19498 gnd.n2984 gnd.t274 7.32958
R19499 gnd.n4321 gnd.t64 7.32958
R19500 gnd.n2084 gnd.t324 7.32958
R19501 gnd.t294 gnd.n1697 7.32958
R19502 gnd.n5237 gnd.t45 7.32958
R19503 gnd.n7247 gnd.n170 7.32958
R19504 gnd.n1197 gnd.n1196 7.30353
R19505 gnd.n5004 gnd.n5003 7.30353
R19506 gnd.n2944 gnd.n2663 7.01093
R19507 gnd.n2666 gnd.n2664 7.01093
R19508 gnd.n2954 gnd.n2953 7.01093
R19509 gnd.n2965 gnd.n2647 7.01093
R19510 gnd.n2964 gnd.n2650 7.01093
R19511 gnd.n2975 gnd.n2638 7.01093
R19512 gnd.n2641 gnd.n2639 7.01093
R19513 gnd.n2985 gnd.n2984 7.01093
R19514 gnd.n2995 gnd.n2619 7.01093
R19515 gnd.n2994 gnd.n2622 7.01093
R19516 gnd.n3003 gnd.n2613 7.01093
R19517 gnd.n3015 gnd.n2603 7.01093
R19518 gnd.n3025 gnd.n2588 7.01093
R19519 gnd.n3041 gnd.n3040 7.01093
R19520 gnd.n2590 gnd.n2527 7.01093
R19521 gnd.n3095 gnd.n2528 7.01093
R19522 gnd.n3089 gnd.n3088 7.01093
R19523 gnd.n2577 gnd.n2539 7.01093
R19524 gnd.n3081 gnd.n2550 7.01093
R19525 gnd.n2568 gnd.n2563 7.01093
R19526 gnd.n3075 gnd.n3074 7.01093
R19527 gnd.n3121 gnd.n2466 7.01093
R19528 gnd.n3120 gnd.n3119 7.01093
R19529 gnd.n3132 gnd.n3131 7.01093
R19530 gnd.n2459 gnd.n2451 7.01093
R19531 gnd.n3161 gnd.n2439 7.01093
R19532 gnd.n3160 gnd.n2442 7.01093
R19533 gnd.n3171 gnd.n2431 7.01093
R19534 gnd.n2432 gnd.n2420 7.01093
R19535 gnd.n3182 gnd.n2421 7.01093
R19536 gnd.n3206 gnd.n2412 7.01093
R19537 gnd.n3205 gnd.n2403 7.01093
R19538 gnd.n3228 gnd.n3227 7.01093
R19539 gnd.n3246 gnd.n2384 7.01093
R19540 gnd.n3245 gnd.n2387 7.01093
R19541 gnd.n3256 gnd.n2376 7.01093
R19542 gnd.n2377 gnd.n2364 7.01093
R19543 gnd.n3267 gnd.n2365 7.01093
R19544 gnd.n3294 gnd.n2349 7.01093
R19545 gnd.n3306 gnd.n3305 7.01093
R19546 gnd.n3288 gnd.n2342 7.01093
R19547 gnd.n3317 gnd.n3316 7.01093
R19548 gnd.n3589 gnd.n2330 7.01093
R19549 gnd.n3588 gnd.n2333 7.01093
R19550 gnd.n3601 gnd.n2322 7.01093
R19551 gnd.n2323 gnd.n2315 7.01093
R19552 gnd.n3611 gnd.n2241 7.01093
R19553 gnd.n4983 gnd.t90 7.01093
R19554 gnd.n2622 gnd.t283 6.69227
R19555 gnd.n2442 gnd.t11 6.69227
R19556 gnd.n2365 gnd.n726 6.69227
R19557 gnd.n3295 gnd.t287 6.69227
R19558 gnd.n4705 gnd.t20 6.69227
R19559 gnd.n4791 gnd.t320 6.69227
R19560 gnd.n5140 gnd.n5139 6.5566
R19561 gnd.n4433 gnd.n4432 6.5566
R19562 gnd.n5789 gnd.n5785 6.5566
R19563 gnd.n5015 gnd.n5014 6.5566
R19564 gnd.n2025 gnd.n2013 6.37362
R19565 gnd.n4614 gnd.n2003 6.37362
R19566 gnd.n4658 gnd.t303 6.37362
R19567 gnd.n4742 gnd.n1930 6.37362
R19568 gnd.n4748 gnd.n1920 6.37362
R19569 gnd.n4849 gnd.t308 6.37362
R19570 gnd.n1845 gnd.n1831 6.37362
R19571 gnd.n4920 gnd.n1821 6.37362
R19572 gnd.n957 gnd.n955 6.20656
R19573 gnd.n1663 gnd.n1375 6.20656
R19574 gnd.t326 gnd.n3051 6.05496
R19575 gnd.n3052 gnd.t280 6.05496
R19576 gnd.t268 gnd.n2466 6.05496
R19577 gnd.t277 gnd.n3216 6.05496
R19578 gnd.t14 gnd.n2008 6.05496
R19579 gnd.n4901 gnd.t18 6.05496
R19580 gnd.n3574 gnd.n3544 5.81868
R19581 gnd.n3542 gnd.n3512 5.81868
R19582 gnd.n3510 gnd.n3480 5.81868
R19583 gnd.n3479 gnd.n3449 5.81868
R19584 gnd.n3447 gnd.n3417 5.81868
R19585 gnd.n3415 gnd.n3385 5.81868
R19586 gnd.n3383 gnd.n3353 5.81868
R19587 gnd.n3352 gnd.n3322 5.81868
R19588 gnd.n5144 gnd.n1455 5.62001
R19589 gnd.n5851 gnd.n1139 5.62001
R19590 gnd.n5851 gnd.n1140 5.62001
R19591 gnd.n5010 gnd.n1455 5.62001
R19592 gnd.n2803 gnd.n2798 5.4308
R19593 gnd.n3619 gnd.n2308 5.4308
R19594 gnd.n3119 gnd.t275 5.41765
R19595 gnd.t278 gnd.n3142 5.41765
R19596 gnd.t292 gnd.n2396 5.41765
R19597 gnd.n4566 gnd.t126 5.09899
R19598 gnd.n4596 gnd.n2016 5.09899
R19599 gnd.n4603 gnd.n2009 5.09899
R19600 gnd.t303 gnd.n4657 5.09899
R19601 gnd.n4755 gnd.n1924 5.09899
R19602 gnd.n4763 gnd.n1917 5.09899
R19603 gnd.t308 gnd.n4848 5.09899
R19604 gnd.n4900 gnd.n1834 5.09899
R19605 gnd.n4907 gnd.n1827 5.09899
R19606 gnd.n3572 gnd.n3571 5.04292
R19607 gnd.n3540 gnd.n3539 5.04292
R19608 gnd.n3508 gnd.n3507 5.04292
R19609 gnd.n3477 gnd.n3476 5.04292
R19610 gnd.n3445 gnd.n3444 5.04292
R19611 gnd.n3413 gnd.n3412 5.04292
R19612 gnd.n3381 gnd.n3380 5.04292
R19613 gnd.n3350 gnd.n3349 5.04292
R19614 gnd.n3082 gnd.t279 4.78034
R19615 gnd.n2421 gnd.t286 4.78034
R19616 gnd.n4377 gnd.t7 4.78034
R19617 gnd.n5147 gnd.t111 4.78034
R19618 gnd.n5174 gnd.t264 4.78034
R19619 gnd.n2524 gnd.n2521 4.74817
R19620 gnd.n2574 gnd.n2472 4.74817
R19621 gnd.n2561 gnd.n2471 4.74817
R19622 gnd.n2470 gnd.n2469 4.74817
R19623 gnd.n2570 gnd.n2521 4.74817
R19624 gnd.n2571 gnd.n2472 4.74817
R19625 gnd.n2573 gnd.n2471 4.74817
R19626 gnd.n2560 gnd.n2470 4.74817
R19627 gnd.n5406 gnd.n86 4.74817
R19628 gnd.n1591 gnd.n85 4.74817
R19629 gnd.n1601 gnd.n84 4.74817
R19630 gnd.n7301 gnd.n79 4.74817
R19631 gnd.n7299 gnd.n80 4.74817
R19632 gnd.n5417 gnd.n86 4.74817
R19633 gnd.n5407 gnd.n85 4.74817
R19634 gnd.n1590 gnd.n84 4.74817
R19635 gnd.n1600 gnd.n79 4.74817
R19636 gnd.n7300 gnd.n7299 4.74817
R19637 gnd.n4116 gnd.n731 4.74817
R19638 gnd.n4123 gnd.n4120 4.74817
R19639 gnd.n4121 gnd.n2153 4.74817
R19640 gnd.n4158 gnd.n4157 4.74817
R19641 gnd.n4162 gnd.n2151 4.74817
R19642 gnd.n5339 gnd.n5338 4.74817
R19643 gnd.n5401 gnd.n1596 4.74817
R19644 gnd.n5399 gnd.n5398 4.74817
R19645 gnd.n1597 gnd.n183 4.74817
R19646 gnd.n6880 gnd.n6879 4.74817
R19647 gnd.n5340 gnd.n5339 4.74817
R19648 gnd.n5336 gnd.n1596 4.74817
R19649 gnd.n5400 gnd.n5399 4.74817
R19650 gnd.n1598 gnd.n1597 4.74817
R19651 gnd.n6881 gnd.n6880 4.74817
R19652 gnd.n6063 gnd.n6062 4.74817
R19653 gnd.n760 gnd.n742 4.74817
R19654 gnd.n6050 gnd.n6049 4.74817
R19655 gnd.n777 gnd.n761 4.74817
R19656 gnd.n6037 gnd.n6036 4.74817
R19657 gnd.n6064 gnd.n6063 4.74817
R19658 gnd.n6061 gnd.n742 4.74817
R19659 gnd.n6051 gnd.n6050 4.74817
R19660 gnd.n6048 gnd.n761 4.74817
R19661 gnd.n6038 gnd.n6037 4.74817
R19662 gnd.n4118 gnd.n4116 4.74817
R19663 gnd.n4120 gnd.n4119 4.74817
R19664 gnd.n4122 gnd.n4121 4.74817
R19665 gnd.n4157 gnd.n4156 4.74817
R19666 gnd.n4159 gnd.n2151 4.74817
R19667 gnd.n2519 gnd.n2518 4.74296
R19668 gnd.n66 gnd.n65 4.74296
R19669 gnd.n2495 gnd.n2494 4.7074
R19670 gnd.n2507 gnd.n2506 4.7074
R19671 gnd.n42 gnd.n41 4.7074
R19672 gnd.n54 gnd.n53 4.7074
R19673 gnd.n2519 gnd.n2507 4.65959
R19674 gnd.n66 gnd.n54 4.65959
R19675 gnd.n5533 gnd.n1457 4.6132
R19676 gnd.n5852 gnd.n1138 4.6132
R19677 gnd.t75 gnd.n2035 4.46168
R19678 gnd.n5000 gnd.n4987 4.46111
R19679 gnd.n3557 gnd.n3553 4.38594
R19680 gnd.n3525 gnd.n3521 4.38594
R19681 gnd.n3493 gnd.n3489 4.38594
R19682 gnd.n3462 gnd.n3458 4.38594
R19683 gnd.n3430 gnd.n3426 4.38594
R19684 gnd.n3398 gnd.n3394 4.38594
R19685 gnd.n3366 gnd.n3362 4.38594
R19686 gnd.n3335 gnd.n3331 4.38594
R19687 gnd.n3568 gnd.n3546 4.26717
R19688 gnd.n3536 gnd.n3514 4.26717
R19689 gnd.n3504 gnd.n3482 4.26717
R19690 gnd.n3473 gnd.n3451 4.26717
R19691 gnd.n3441 gnd.n3419 4.26717
R19692 gnd.n3409 gnd.n3387 4.26717
R19693 gnd.n3377 gnd.n3355 4.26717
R19694 gnd.n3346 gnd.n3324 4.26717
R19695 gnd.n3026 gnd.t281 4.14303
R19696 gnd.n3256 gnd.t285 4.14303
R19697 gnd.n867 gnd.t60 4.14303
R19698 gnd.n5308 gnd.t31 4.14303
R19699 gnd.n3576 gnd.n3575 4.08274
R19700 gnd.n5139 gnd.n5138 4.05904
R19701 gnd.n4434 gnd.n4433 4.05904
R19702 gnd.n5792 gnd.n5785 4.05904
R19703 gnd.n5016 gnd.n5015 4.05904
R19704 gnd.n19 gnd.n9 3.99943
R19705 gnd.n4586 gnd.n4584 3.82437
R19706 gnd.n4624 gnd.t1 3.82437
R19707 gnd.n4735 gnd.n1938 3.82437
R19708 gnd.n4772 gnd.n4771 3.82437
R19709 gnd.n4890 gnd.t296 3.82437
R19710 gnd.n4930 gnd.n1812 3.82437
R19711 gnd.n4946 gnd.t42 3.82437
R19712 gnd.n3099 gnd.n2520 3.81325
R19713 gnd.n2507 gnd.n2495 3.72967
R19714 gnd.n54 gnd.n42 3.72967
R19715 gnd.n3576 gnd.n3448 3.70378
R19716 gnd.n19 gnd.n18 3.60163
R19717 gnd.n3567 gnd.n3548 3.49141
R19718 gnd.n3535 gnd.n3516 3.49141
R19719 gnd.n3503 gnd.n3484 3.49141
R19720 gnd.n3472 gnd.n3453 3.49141
R19721 gnd.n3440 gnd.n3421 3.49141
R19722 gnd.n3408 gnd.n3389 3.49141
R19723 gnd.n3376 gnd.n3357 3.49141
R19724 gnd.n3345 gnd.n3326 3.49141
R19725 gnd.n5551 gnd.n5550 3.29747
R19726 gnd.n5550 gnd.n5549 3.29747
R19727 gnd.n7153 gnd.n7150 3.29747
R19728 gnd.n7154 gnd.n7153 3.29747
R19729 gnd.n3810 gnd.n3806 3.29747
R19730 gnd.n3956 gnd.n3810 3.29747
R19731 gnd.n5870 gnd.n5869 3.29747
R19732 gnd.n5869 gnd.n5868 3.29747
R19733 gnd.n4705 gnd.t0 3.18706
R19734 gnd.n4791 gnd.t13 3.18706
R19735 gnd.t78 gnd.n1794 3.18706
R19736 gnd.n2605 gnd.t281 2.8684
R19737 gnd.n4521 gnd.t311 2.8684
R19738 gnd.n4983 gnd.t266 2.8684
R19739 gnd.n2508 gnd.t222 2.82907
R19740 gnd.n2508 gnd.t263 2.82907
R19741 gnd.n2510 gnd.t186 2.82907
R19742 gnd.n2510 gnd.t254 2.82907
R19743 gnd.n2512 gnd.t155 2.82907
R19744 gnd.n2512 gnd.t240 2.82907
R19745 gnd.n2514 gnd.t258 2.82907
R19746 gnd.n2514 gnd.t184 2.82907
R19747 gnd.n2516 gnd.t210 2.82907
R19748 gnd.n2516 gnd.t147 2.82907
R19749 gnd.n2473 gnd.t227 2.82907
R19750 gnd.n2473 gnd.t239 2.82907
R19751 gnd.n2475 gnd.t246 2.82907
R19752 gnd.n2475 gnd.t260 2.82907
R19753 gnd.n2477 gnd.t219 2.82907
R19754 gnd.n2477 gnd.t231 2.82907
R19755 gnd.n2479 gnd.t241 2.82907
R19756 gnd.n2479 gnd.t167 2.82907
R19757 gnd.n2481 gnd.t230 2.82907
R19758 gnd.n2481 gnd.t226 2.82907
R19759 gnd.n2484 gnd.t212 2.82907
R19760 gnd.n2484 gnd.t202 2.82907
R19761 gnd.n2486 gnd.t203 2.82907
R19762 gnd.n2486 gnd.t225 2.82907
R19763 gnd.n2488 gnd.t182 2.82907
R19764 gnd.n2488 gnd.t213 2.82907
R19765 gnd.n2490 gnd.t214 2.82907
R19766 gnd.n2490 gnd.t194 2.82907
R19767 gnd.n2492 gnd.t153 2.82907
R19768 gnd.n2492 gnd.t183 2.82907
R19769 gnd.n2496 gnd.t250 2.82907
R19770 gnd.n2496 gnd.t218 2.82907
R19771 gnd.n2498 gnd.t235 2.82907
R19772 gnd.n2498 gnd.t197 2.82907
R19773 gnd.n2500 gnd.t221 2.82907
R19774 gnd.n2500 gnd.t161 2.82907
R19775 gnd.n2502 gnd.t200 2.82907
R19776 gnd.n2502 gnd.t234 2.82907
R19777 gnd.n2504 gnd.t245 2.82907
R19778 gnd.n2504 gnd.t237 2.82907
R19779 gnd.n63 gnd.t262 2.82907
R19780 gnd.n63 gnd.t180 2.82907
R19781 gnd.n61 gnd.t259 2.82907
R19782 gnd.n61 gnd.t236 2.82907
R19783 gnd.n59 gnd.t220 2.82907
R19784 gnd.n59 gnd.t252 2.82907
R19785 gnd.n57 gnd.t233 2.82907
R19786 gnd.n57 gnd.t261 2.82907
R19787 gnd.n55 gnd.t242 2.82907
R19788 gnd.n55 gnd.t175 2.82907
R19789 gnd.n28 gnd.t244 2.82907
R19790 gnd.n28 gnd.t223 2.82907
R19791 gnd.n26 gnd.t209 2.82907
R19792 gnd.n26 gnd.t257 2.82907
R19793 gnd.n24 gnd.t251 2.82907
R19794 gnd.n24 gnd.t198 2.82907
R19795 gnd.n22 gnd.t181 2.82907
R19796 gnd.n22 gnd.t149 2.82907
R19797 gnd.n20 gnd.t256 2.82907
R19798 gnd.n20 gnd.t243 2.82907
R19799 gnd.n39 gnd.t163 2.82907
R19800 gnd.n39 gnd.t173 2.82907
R19801 gnd.n37 gnd.t171 2.82907
R19802 gnd.n37 gnd.t192 2.82907
R19803 gnd.n35 gnd.t191 2.82907
R19804 gnd.n35 gnd.t207 2.82907
R19805 gnd.n33 gnd.t205 2.82907
R19806 gnd.n33 gnd.t179 2.82907
R19807 gnd.n31 gnd.t178 2.82907
R19808 gnd.n31 gnd.t187 2.82907
R19809 gnd.n51 gnd.t217 2.82907
R19810 gnd.n51 gnd.t232 2.82907
R19811 gnd.n49 gnd.t206 2.82907
R19812 gnd.n49 gnd.t157 2.82907
R19813 gnd.n47 gnd.t249 2.82907
R19814 gnd.n47 gnd.t189 2.82907
R19815 gnd.n45 gnd.t145 2.82907
R19816 gnd.n45 gnd.t208 2.82907
R19817 gnd.n43 gnd.t169 2.82907
R19818 gnd.n43 gnd.t229 2.82907
R19819 gnd.n3564 gnd.n3563 2.71565
R19820 gnd.n3532 gnd.n3531 2.71565
R19821 gnd.n3500 gnd.n3499 2.71565
R19822 gnd.n3469 gnd.n3468 2.71565
R19823 gnd.n3437 gnd.n3436 2.71565
R19824 gnd.n3405 gnd.n3404 2.71565
R19825 gnd.n3373 gnd.n3372 2.71565
R19826 gnd.n3342 gnd.n3341 2.71565
R19827 gnd.n5771 gnd.t49 2.54975
R19828 gnd.n4566 gnd.n4565 2.54975
R19829 gnd.n4638 gnd.n1987 2.54975
R19830 gnd.n4725 gnd.n4724 2.54975
R19831 gnd.n4800 gnd.n1891 2.54975
R19832 gnd.n4840 gnd.n1849 2.54975
R19833 gnd.n4938 gnd.n1805 2.54975
R19834 gnd.t140 gnd.n4972 2.54975
R19835 gnd.n3099 gnd.n2521 2.27742
R19836 gnd.n3099 gnd.n2472 2.27742
R19837 gnd.n3099 gnd.n2471 2.27742
R19838 gnd.n3099 gnd.n2470 2.27742
R19839 gnd.n7298 gnd.n86 2.27742
R19840 gnd.n7298 gnd.n85 2.27742
R19841 gnd.n7298 gnd.n84 2.27742
R19842 gnd.n7298 gnd.n79 2.27742
R19843 gnd.n7299 gnd.n7298 2.27742
R19844 gnd.n5339 gnd.n83 2.27742
R19845 gnd.n1596 gnd.n83 2.27742
R19846 gnd.n5399 gnd.n83 2.27742
R19847 gnd.n1597 gnd.n83 2.27742
R19848 gnd.n6880 gnd.n83 2.27742
R19849 gnd.n6063 gnd.n741 2.27742
R19850 gnd.n742 gnd.n741 2.27742
R19851 gnd.n6050 gnd.n741 2.27742
R19852 gnd.n761 gnd.n741 2.27742
R19853 gnd.n6037 gnd.n741 2.27742
R19854 gnd.n4116 gnd.n730 2.27742
R19855 gnd.n4120 gnd.n730 2.27742
R19856 gnd.n4121 gnd.n730 2.27742
R19857 gnd.n4157 gnd.n730 2.27742
R19858 gnd.n2151 gnd.n730 2.27742
R19859 gnd.n2953 gnd.t71 2.23109
R19860 gnd.n2576 gnd.t279 2.23109
R19861 gnd.n4125 gnd.t154 2.23109
R19862 gnd.t188 gnd.n73 2.23109
R19863 gnd.n3560 gnd.n3550 1.93989
R19864 gnd.n3528 gnd.n3518 1.93989
R19865 gnd.n3496 gnd.n3486 1.93989
R19866 gnd.n3465 gnd.n3455 1.93989
R19867 gnd.n3433 gnd.n3423 1.93989
R19868 gnd.n3401 gnd.n3391 1.93989
R19869 gnd.n3369 gnd.n3359 1.93989
R19870 gnd.n3338 gnd.n3328 1.93989
R19871 gnd.n4423 gnd.t93 1.91244
R19872 gnd.n1938 gnd.t319 1.91244
R19873 gnd.n4772 gnd.t4 1.91244
R19874 gnd.t290 gnd.n2964 1.59378
R19875 gnd.n3143 gnd.t278 1.59378
R19876 gnd.n2405 gnd.t292 1.59378
R19877 gnd.n4170 gnd.t196 1.59378
R19878 gnd.n4578 gnd.t306 1.59378
R19879 gnd.t322 gnd.n1983 1.59378
R19880 gnd.n4859 gnd.t270 1.59378
R19881 gnd.n4913 gnd.t297 1.59378
R19882 gnd.n1617 gnd.t144 1.59378
R19883 gnd.n4492 gnd.n1201 1.27512
R19884 gnd.n4515 gnd.t23 1.27512
R19885 gnd.n4504 gnd.n4501 1.27512
R19886 gnd.n4586 gnd.t302 1.27512
R19887 gnd.n4650 gnd.n1977 1.27512
R19888 gnd.n4693 gnd.n1951 1.27512
R19889 gnd.n4810 gnd.n1884 1.27512
R19890 gnd.n4825 gnd.n1867 1.27512
R19891 gnd.n4930 gnd.t305 1.27512
R19892 gnd.n4973 gnd.n1788 1.27512
R19893 gnd.n4972 gnd.t52 1.27512
R19894 gnd.n4946 gnd.n1732 1.27512
R19895 gnd.n2806 gnd.n2798 1.16414
R19896 gnd.n3622 gnd.n2308 1.16414
R19897 gnd.n3559 gnd.n3552 1.16414
R19898 gnd.n3527 gnd.n3520 1.16414
R19899 gnd.n3495 gnd.n3488 1.16414
R19900 gnd.n3464 gnd.n3457 1.16414
R19901 gnd.n3432 gnd.n3425 1.16414
R19902 gnd.n3400 gnd.n3393 1.16414
R19903 gnd.n3368 gnd.n3361 1.16414
R19904 gnd.n3337 gnd.n3330 1.16414
R19905 gnd.n5533 gnd.n5532 0.970197
R19906 gnd.n5852 gnd.n1040 0.970197
R19907 gnd.n3543 gnd.n3511 0.962709
R19908 gnd.n3575 gnd.n3543 0.962709
R19909 gnd.n3416 gnd.n3384 0.962709
R19910 gnd.n3448 gnd.n3416 0.962709
R19911 gnd.n3052 gnd.t326 0.956468
R19912 gnd.n3217 gnd.t277 0.956468
R19913 gnd.n4060 gnd.t152 0.956468
R19914 gnd.n4186 gnd.t201 0.956468
R19915 gnd.n4190 gnd.t158 0.956468
R19916 gnd.n5280 gnd.t164 0.956468
R19917 gnd.n5290 gnd.t168 0.956468
R19918 gnd.n130 gnd.t172 0.956468
R19919 gnd.n2 gnd.n1 0.672012
R19920 gnd.n3 gnd.n2 0.672012
R19921 gnd.n4 gnd.n3 0.672012
R19922 gnd.n5 gnd.n4 0.672012
R19923 gnd.n6 gnd.n5 0.672012
R19924 gnd.n7 gnd.n6 0.672012
R19925 gnd.n8 gnd.n7 0.672012
R19926 gnd.n9 gnd.n8 0.672012
R19927 gnd.n11 gnd.n10 0.672012
R19928 gnd.n12 gnd.n11 0.672012
R19929 gnd.n13 gnd.n12 0.672012
R19930 gnd.n14 gnd.n13 0.672012
R19931 gnd.n15 gnd.n14 0.672012
R19932 gnd.n16 gnd.n15 0.672012
R19933 gnd.n17 gnd.n16 0.672012
R19934 gnd.n18 gnd.n17 0.672012
R19935 gnd gnd.n0 0.624033
R19936 gnd.n2518 gnd.n2517 0.573776
R19937 gnd.n2517 gnd.n2515 0.573776
R19938 gnd.n2515 gnd.n2513 0.573776
R19939 gnd.n2513 gnd.n2511 0.573776
R19940 gnd.n2511 gnd.n2509 0.573776
R19941 gnd.n2483 gnd.n2482 0.573776
R19942 gnd.n2482 gnd.n2480 0.573776
R19943 gnd.n2480 gnd.n2478 0.573776
R19944 gnd.n2478 gnd.n2476 0.573776
R19945 gnd.n2476 gnd.n2474 0.573776
R19946 gnd.n2494 gnd.n2493 0.573776
R19947 gnd.n2493 gnd.n2491 0.573776
R19948 gnd.n2491 gnd.n2489 0.573776
R19949 gnd.n2489 gnd.n2487 0.573776
R19950 gnd.n2487 gnd.n2485 0.573776
R19951 gnd.n2506 gnd.n2505 0.573776
R19952 gnd.n2505 gnd.n2503 0.573776
R19953 gnd.n2503 gnd.n2501 0.573776
R19954 gnd.n2501 gnd.n2499 0.573776
R19955 gnd.n2499 gnd.n2497 0.573776
R19956 gnd.n58 gnd.n56 0.573776
R19957 gnd.n60 gnd.n58 0.573776
R19958 gnd.n62 gnd.n60 0.573776
R19959 gnd.n64 gnd.n62 0.573776
R19960 gnd.n65 gnd.n64 0.573776
R19961 gnd.n23 gnd.n21 0.573776
R19962 gnd.n25 gnd.n23 0.573776
R19963 gnd.n27 gnd.n25 0.573776
R19964 gnd.n29 gnd.n27 0.573776
R19965 gnd.n30 gnd.n29 0.573776
R19966 gnd.n34 gnd.n32 0.573776
R19967 gnd.n36 gnd.n34 0.573776
R19968 gnd.n38 gnd.n36 0.573776
R19969 gnd.n40 gnd.n38 0.573776
R19970 gnd.n41 gnd.n40 0.573776
R19971 gnd.n46 gnd.n44 0.573776
R19972 gnd.n48 gnd.n46 0.573776
R19973 gnd.n50 gnd.n48 0.573776
R19974 gnd.n52 gnd.n50 0.573776
R19975 gnd.n53 gnd.n52 0.573776
R19976 gnd.n7191 gnd.n7190 0.532512
R19977 gnd.n3774 gnd.n3773 0.532512
R19978 gnd.n7006 gnd.n165 0.497451
R19979 gnd.n1012 gnd.n857 0.497451
R19980 gnd.n1508 gnd.n1427 0.497451
R19981 gnd.n3994 gnd.n3993 0.497451
R19982 gnd.n3279 gnd.n2312 0.486781
R19983 gnd.n2855 gnd.n2854 0.48678
R19984 gnd.n3596 gnd.n2266 0.480683
R19985 gnd.n2939 gnd.n2938 0.480683
R19986 gnd.n6242 gnd.n6241 0.480683
R19987 gnd.n6663 gnd.n6662 0.480683
R19988 gnd.n6874 gnd.n184 0.480683
R19989 gnd.n6071 gnd.n6070 0.480683
R19990 gnd.n7310 gnd.n7309 0.4705
R19991 gnd.n1639 gnd.n1309 0.451719
R19992 gnd.n4316 gnd.n871 0.451719
R19993 gnd.n4264 gnd.n894 0.451719
R19994 gnd.n5651 gnd.n5650 0.451719
R19995 gnd.n7298 gnd.n83 0.4255
R19996 gnd.n741 gnd.n730 0.4255
R19997 gnd.n5910 gnd.n955 0.388379
R19998 gnd.n3556 gnd.n3555 0.388379
R19999 gnd.n3524 gnd.n3523 0.388379
R20000 gnd.n3492 gnd.n3491 0.388379
R20001 gnd.n3461 gnd.n3460 0.388379
R20002 gnd.n3429 gnd.n3428 0.388379
R20003 gnd.n3397 gnd.n3396 0.388379
R20004 gnd.n3365 gnd.n3364 0.388379
R20005 gnd.n3334 gnd.n3333 0.388379
R20006 gnd.n5595 gnd.n1375 0.388379
R20007 gnd.n7310 gnd.n19 0.374463
R20008 gnd gnd.n7310 0.367492
R20009 gnd.n2367 gnd.t287 0.319156
R20010 gnd.n4108 gnd.t166 0.319156
R20011 gnd.n4145 gnd.t185 0.319156
R20012 gnd.t319 gnd.t16 0.319156
R20013 gnd.t2 gnd.t4 0.319156
R20014 gnd.n5377 gnd.t148 0.319156
R20015 gnd.n6891 gnd.t170 0.319156
R20016 gnd.n2773 gnd.n2751 0.311721
R20017 gnd.n5974 gnd.n5973 0.302329
R20018 gnd.n5266 gnd.n5265 0.302329
R20019 gnd.n6932 gnd.n173 0.293183
R20020 gnd.n3726 gnd.n2239 0.293183
R20021 gnd.n3667 gnd.n3666 0.268793
R20022 gnd.n7067 gnd.n173 0.258122
R20023 gnd.n5471 gnd.n1328 0.258122
R20024 gnd.n1073 gnd.n865 0.258122
R20025 gnd.n3875 gnd.n2239 0.258122
R20026 gnd.n3666 gnd.n3665 0.241354
R20027 gnd.n1457 gnd.n1454 0.229039
R20028 gnd.n1458 gnd.n1457 0.229039
R20029 gnd.n1138 gnd.n1039 0.229039
R20030 gnd.n1138 gnd.n1137 0.229039
R20031 gnd.n2927 gnd.n2726 0.206293
R20032 gnd.n3573 gnd.n3545 0.155672
R20033 gnd.n3566 gnd.n3545 0.155672
R20034 gnd.n3566 gnd.n3565 0.155672
R20035 gnd.n3565 gnd.n3549 0.155672
R20036 gnd.n3558 gnd.n3549 0.155672
R20037 gnd.n3558 gnd.n3557 0.155672
R20038 gnd.n3541 gnd.n3513 0.155672
R20039 gnd.n3534 gnd.n3513 0.155672
R20040 gnd.n3534 gnd.n3533 0.155672
R20041 gnd.n3533 gnd.n3517 0.155672
R20042 gnd.n3526 gnd.n3517 0.155672
R20043 gnd.n3526 gnd.n3525 0.155672
R20044 gnd.n3509 gnd.n3481 0.155672
R20045 gnd.n3502 gnd.n3481 0.155672
R20046 gnd.n3502 gnd.n3501 0.155672
R20047 gnd.n3501 gnd.n3485 0.155672
R20048 gnd.n3494 gnd.n3485 0.155672
R20049 gnd.n3494 gnd.n3493 0.155672
R20050 gnd.n3478 gnd.n3450 0.155672
R20051 gnd.n3471 gnd.n3450 0.155672
R20052 gnd.n3471 gnd.n3470 0.155672
R20053 gnd.n3470 gnd.n3454 0.155672
R20054 gnd.n3463 gnd.n3454 0.155672
R20055 gnd.n3463 gnd.n3462 0.155672
R20056 gnd.n3446 gnd.n3418 0.155672
R20057 gnd.n3439 gnd.n3418 0.155672
R20058 gnd.n3439 gnd.n3438 0.155672
R20059 gnd.n3438 gnd.n3422 0.155672
R20060 gnd.n3431 gnd.n3422 0.155672
R20061 gnd.n3431 gnd.n3430 0.155672
R20062 gnd.n3414 gnd.n3386 0.155672
R20063 gnd.n3407 gnd.n3386 0.155672
R20064 gnd.n3407 gnd.n3406 0.155672
R20065 gnd.n3406 gnd.n3390 0.155672
R20066 gnd.n3399 gnd.n3390 0.155672
R20067 gnd.n3399 gnd.n3398 0.155672
R20068 gnd.n3382 gnd.n3354 0.155672
R20069 gnd.n3375 gnd.n3354 0.155672
R20070 gnd.n3375 gnd.n3374 0.155672
R20071 gnd.n3374 gnd.n3358 0.155672
R20072 gnd.n3367 gnd.n3358 0.155672
R20073 gnd.n3367 gnd.n3366 0.155672
R20074 gnd.n3351 gnd.n3323 0.155672
R20075 gnd.n3344 gnd.n3323 0.155672
R20076 gnd.n3344 gnd.n3343 0.155672
R20077 gnd.n3343 gnd.n3327 0.155672
R20078 gnd.n3336 gnd.n3327 0.155672
R20079 gnd.n3336 gnd.n3335 0.155672
R20080 gnd.n3698 gnd.n2266 0.152939
R20081 gnd.n3698 gnd.n3697 0.152939
R20082 gnd.n3697 gnd.n3696 0.152939
R20083 gnd.n3696 gnd.n2268 0.152939
R20084 gnd.n2269 gnd.n2268 0.152939
R20085 gnd.n2270 gnd.n2269 0.152939
R20086 gnd.n2271 gnd.n2270 0.152939
R20087 gnd.n2272 gnd.n2271 0.152939
R20088 gnd.n2273 gnd.n2272 0.152939
R20089 gnd.n2274 gnd.n2273 0.152939
R20090 gnd.n2275 gnd.n2274 0.152939
R20091 gnd.n2276 gnd.n2275 0.152939
R20092 gnd.n2277 gnd.n2276 0.152939
R20093 gnd.n2278 gnd.n2277 0.152939
R20094 gnd.n3668 gnd.n2278 0.152939
R20095 gnd.n3668 gnd.n3667 0.152939
R20096 gnd.n2940 gnd.n2939 0.152939
R20097 gnd.n2940 gnd.n2644 0.152939
R20098 gnd.n2968 gnd.n2644 0.152939
R20099 gnd.n2969 gnd.n2968 0.152939
R20100 gnd.n2970 gnd.n2969 0.152939
R20101 gnd.n2971 gnd.n2970 0.152939
R20102 gnd.n2971 gnd.n2616 0.152939
R20103 gnd.n2998 gnd.n2616 0.152939
R20104 gnd.n2999 gnd.n2998 0.152939
R20105 gnd.n3000 gnd.n2999 0.152939
R20106 gnd.n3000 gnd.n2594 0.152939
R20107 gnd.n3029 gnd.n2594 0.152939
R20108 gnd.n3030 gnd.n3029 0.152939
R20109 gnd.n3031 gnd.n3030 0.152939
R20110 gnd.n3032 gnd.n3031 0.152939
R20111 gnd.n3034 gnd.n3032 0.152939
R20112 gnd.n3034 gnd.n3033 0.152939
R20113 gnd.n3033 gnd.n2543 0.152939
R20114 gnd.n2544 gnd.n2543 0.152939
R20115 gnd.n2545 gnd.n2544 0.152939
R20116 gnd.n2564 gnd.n2545 0.152939
R20117 gnd.n2565 gnd.n2564 0.152939
R20118 gnd.n2565 gnd.n2463 0.152939
R20119 gnd.n3124 gnd.n2463 0.152939
R20120 gnd.n3125 gnd.n3124 0.152939
R20121 gnd.n3126 gnd.n3125 0.152939
R20122 gnd.n3127 gnd.n3126 0.152939
R20123 gnd.n3127 gnd.n2436 0.152939
R20124 gnd.n3164 gnd.n2436 0.152939
R20125 gnd.n3165 gnd.n3164 0.152939
R20126 gnd.n3166 gnd.n3165 0.152939
R20127 gnd.n3167 gnd.n3166 0.152939
R20128 gnd.n3167 gnd.n2409 0.152939
R20129 gnd.n3209 gnd.n2409 0.152939
R20130 gnd.n3210 gnd.n3209 0.152939
R20131 gnd.n3211 gnd.n3210 0.152939
R20132 gnd.n3212 gnd.n3211 0.152939
R20133 gnd.n3212 gnd.n2381 0.152939
R20134 gnd.n3249 gnd.n2381 0.152939
R20135 gnd.n3250 gnd.n3249 0.152939
R20136 gnd.n3251 gnd.n3250 0.152939
R20137 gnd.n3252 gnd.n3251 0.152939
R20138 gnd.n3252 gnd.n2354 0.152939
R20139 gnd.n3298 gnd.n2354 0.152939
R20140 gnd.n3299 gnd.n3298 0.152939
R20141 gnd.n3300 gnd.n3299 0.152939
R20142 gnd.n3301 gnd.n3300 0.152939
R20143 gnd.n3301 gnd.n2327 0.152939
R20144 gnd.n3592 gnd.n2327 0.152939
R20145 gnd.n3593 gnd.n3592 0.152939
R20146 gnd.n3594 gnd.n3593 0.152939
R20147 gnd.n3595 gnd.n3594 0.152939
R20148 gnd.n3596 gnd.n3595 0.152939
R20149 gnd.n2938 gnd.n2668 0.152939
R20150 gnd.n2689 gnd.n2668 0.152939
R20151 gnd.n2690 gnd.n2689 0.152939
R20152 gnd.n2696 gnd.n2690 0.152939
R20153 gnd.n2697 gnd.n2696 0.152939
R20154 gnd.n2698 gnd.n2697 0.152939
R20155 gnd.n2698 gnd.n2687 0.152939
R20156 gnd.n2706 gnd.n2687 0.152939
R20157 gnd.n2707 gnd.n2706 0.152939
R20158 gnd.n2708 gnd.n2707 0.152939
R20159 gnd.n2708 gnd.n2685 0.152939
R20160 gnd.n2716 gnd.n2685 0.152939
R20161 gnd.n2717 gnd.n2716 0.152939
R20162 gnd.n2718 gnd.n2717 0.152939
R20163 gnd.n2718 gnd.n2683 0.152939
R20164 gnd.n2726 gnd.n2683 0.152939
R20165 gnd.n3665 gnd.n2283 0.152939
R20166 gnd.n2285 gnd.n2283 0.152939
R20167 gnd.n2286 gnd.n2285 0.152939
R20168 gnd.n2287 gnd.n2286 0.152939
R20169 gnd.n2288 gnd.n2287 0.152939
R20170 gnd.n2289 gnd.n2288 0.152939
R20171 gnd.n2290 gnd.n2289 0.152939
R20172 gnd.n2291 gnd.n2290 0.152939
R20173 gnd.n2292 gnd.n2291 0.152939
R20174 gnd.n2293 gnd.n2292 0.152939
R20175 gnd.n2294 gnd.n2293 0.152939
R20176 gnd.n2295 gnd.n2294 0.152939
R20177 gnd.n2296 gnd.n2295 0.152939
R20178 gnd.n2297 gnd.n2296 0.152939
R20179 gnd.n2298 gnd.n2297 0.152939
R20180 gnd.n2299 gnd.n2298 0.152939
R20181 gnd.n2300 gnd.n2299 0.152939
R20182 gnd.n2301 gnd.n2300 0.152939
R20183 gnd.n2302 gnd.n2301 0.152939
R20184 gnd.n2303 gnd.n2302 0.152939
R20185 gnd.n2304 gnd.n2303 0.152939
R20186 gnd.n2305 gnd.n2304 0.152939
R20187 gnd.n2309 gnd.n2305 0.152939
R20188 gnd.n2310 gnd.n2309 0.152939
R20189 gnd.n2311 gnd.n2310 0.152939
R20190 gnd.n2312 gnd.n2311 0.152939
R20191 gnd.n3101 gnd.n3100 0.152939
R20192 gnd.n3102 gnd.n3101 0.152939
R20193 gnd.n3103 gnd.n3102 0.152939
R20194 gnd.n3104 gnd.n3103 0.152939
R20195 gnd.n3105 gnd.n3104 0.152939
R20196 gnd.n3106 gnd.n3105 0.152939
R20197 gnd.n3106 gnd.n2417 0.152939
R20198 gnd.n3185 gnd.n2417 0.152939
R20199 gnd.n3186 gnd.n3185 0.152939
R20200 gnd.n3187 gnd.n3186 0.152939
R20201 gnd.n3188 gnd.n3187 0.152939
R20202 gnd.n3189 gnd.n3188 0.152939
R20203 gnd.n3190 gnd.n3189 0.152939
R20204 gnd.n3191 gnd.n3190 0.152939
R20205 gnd.n3192 gnd.n3191 0.152939
R20206 gnd.n3193 gnd.n3192 0.152939
R20207 gnd.n3193 gnd.n2361 0.152939
R20208 gnd.n3270 gnd.n2361 0.152939
R20209 gnd.n3271 gnd.n3270 0.152939
R20210 gnd.n3272 gnd.n3271 0.152939
R20211 gnd.n3273 gnd.n3272 0.152939
R20212 gnd.n3274 gnd.n3273 0.152939
R20213 gnd.n3275 gnd.n3274 0.152939
R20214 gnd.n3276 gnd.n3275 0.152939
R20215 gnd.n3277 gnd.n3276 0.152939
R20216 gnd.n3278 gnd.n3277 0.152939
R20217 gnd.n3280 gnd.n3278 0.152939
R20218 gnd.n3280 gnd.n3279 0.152939
R20219 gnd.n2856 gnd.n2855 0.152939
R20220 gnd.n2856 gnd.n2746 0.152939
R20221 gnd.n2871 gnd.n2746 0.152939
R20222 gnd.n2872 gnd.n2871 0.152939
R20223 gnd.n2873 gnd.n2872 0.152939
R20224 gnd.n2873 gnd.n2734 0.152939
R20225 gnd.n2887 gnd.n2734 0.152939
R20226 gnd.n2888 gnd.n2887 0.152939
R20227 gnd.n2889 gnd.n2888 0.152939
R20228 gnd.n2890 gnd.n2889 0.152939
R20229 gnd.n2891 gnd.n2890 0.152939
R20230 gnd.n2892 gnd.n2891 0.152939
R20231 gnd.n2893 gnd.n2892 0.152939
R20232 gnd.n2894 gnd.n2893 0.152939
R20233 gnd.n2895 gnd.n2894 0.152939
R20234 gnd.n2896 gnd.n2895 0.152939
R20235 gnd.n2897 gnd.n2896 0.152939
R20236 gnd.n2898 gnd.n2897 0.152939
R20237 gnd.n2899 gnd.n2898 0.152939
R20238 gnd.n2900 gnd.n2899 0.152939
R20239 gnd.n2901 gnd.n2900 0.152939
R20240 gnd.n2901 gnd.n2600 0.152939
R20241 gnd.n3018 gnd.n2600 0.152939
R20242 gnd.n3019 gnd.n3018 0.152939
R20243 gnd.n3020 gnd.n3019 0.152939
R20244 gnd.n3021 gnd.n3020 0.152939
R20245 gnd.n3021 gnd.n2522 0.152939
R20246 gnd.n3098 gnd.n2522 0.152939
R20247 gnd.n2774 gnd.n2773 0.152939
R20248 gnd.n2775 gnd.n2774 0.152939
R20249 gnd.n2776 gnd.n2775 0.152939
R20250 gnd.n2777 gnd.n2776 0.152939
R20251 gnd.n2778 gnd.n2777 0.152939
R20252 gnd.n2779 gnd.n2778 0.152939
R20253 gnd.n2780 gnd.n2779 0.152939
R20254 gnd.n2781 gnd.n2780 0.152939
R20255 gnd.n2782 gnd.n2781 0.152939
R20256 gnd.n2783 gnd.n2782 0.152939
R20257 gnd.n2784 gnd.n2783 0.152939
R20258 gnd.n2785 gnd.n2784 0.152939
R20259 gnd.n2786 gnd.n2785 0.152939
R20260 gnd.n2787 gnd.n2786 0.152939
R20261 gnd.n2788 gnd.n2787 0.152939
R20262 gnd.n2789 gnd.n2788 0.152939
R20263 gnd.n2790 gnd.n2789 0.152939
R20264 gnd.n2791 gnd.n2790 0.152939
R20265 gnd.n2792 gnd.n2791 0.152939
R20266 gnd.n2793 gnd.n2792 0.152939
R20267 gnd.n2794 gnd.n2793 0.152939
R20268 gnd.n2795 gnd.n2794 0.152939
R20269 gnd.n2799 gnd.n2795 0.152939
R20270 gnd.n2800 gnd.n2799 0.152939
R20271 gnd.n2800 gnd.n2757 0.152939
R20272 gnd.n2854 gnd.n2757 0.152939
R20273 gnd.n6242 gnd.n558 0.152939
R20274 gnd.n6250 gnd.n558 0.152939
R20275 gnd.n6251 gnd.n6250 0.152939
R20276 gnd.n6252 gnd.n6251 0.152939
R20277 gnd.n6252 gnd.n552 0.152939
R20278 gnd.n6260 gnd.n552 0.152939
R20279 gnd.n6261 gnd.n6260 0.152939
R20280 gnd.n6262 gnd.n6261 0.152939
R20281 gnd.n6262 gnd.n546 0.152939
R20282 gnd.n6270 gnd.n546 0.152939
R20283 gnd.n6271 gnd.n6270 0.152939
R20284 gnd.n6272 gnd.n6271 0.152939
R20285 gnd.n6272 gnd.n540 0.152939
R20286 gnd.n6280 gnd.n540 0.152939
R20287 gnd.n6281 gnd.n6280 0.152939
R20288 gnd.n6282 gnd.n6281 0.152939
R20289 gnd.n6282 gnd.n534 0.152939
R20290 gnd.n6290 gnd.n534 0.152939
R20291 gnd.n6291 gnd.n6290 0.152939
R20292 gnd.n6292 gnd.n6291 0.152939
R20293 gnd.n6292 gnd.n528 0.152939
R20294 gnd.n6300 gnd.n528 0.152939
R20295 gnd.n6301 gnd.n6300 0.152939
R20296 gnd.n6302 gnd.n6301 0.152939
R20297 gnd.n6302 gnd.n522 0.152939
R20298 gnd.n6310 gnd.n522 0.152939
R20299 gnd.n6311 gnd.n6310 0.152939
R20300 gnd.n6312 gnd.n6311 0.152939
R20301 gnd.n6312 gnd.n516 0.152939
R20302 gnd.n6320 gnd.n516 0.152939
R20303 gnd.n6321 gnd.n6320 0.152939
R20304 gnd.n6322 gnd.n6321 0.152939
R20305 gnd.n6322 gnd.n510 0.152939
R20306 gnd.n6330 gnd.n510 0.152939
R20307 gnd.n6331 gnd.n6330 0.152939
R20308 gnd.n6332 gnd.n6331 0.152939
R20309 gnd.n6332 gnd.n504 0.152939
R20310 gnd.n6340 gnd.n504 0.152939
R20311 gnd.n6341 gnd.n6340 0.152939
R20312 gnd.n6342 gnd.n6341 0.152939
R20313 gnd.n6342 gnd.n498 0.152939
R20314 gnd.n6350 gnd.n498 0.152939
R20315 gnd.n6351 gnd.n6350 0.152939
R20316 gnd.n6352 gnd.n6351 0.152939
R20317 gnd.n6352 gnd.n492 0.152939
R20318 gnd.n6360 gnd.n492 0.152939
R20319 gnd.n6361 gnd.n6360 0.152939
R20320 gnd.n6362 gnd.n6361 0.152939
R20321 gnd.n6362 gnd.n486 0.152939
R20322 gnd.n6370 gnd.n486 0.152939
R20323 gnd.n6371 gnd.n6370 0.152939
R20324 gnd.n6372 gnd.n6371 0.152939
R20325 gnd.n6372 gnd.n480 0.152939
R20326 gnd.n6380 gnd.n480 0.152939
R20327 gnd.n6381 gnd.n6380 0.152939
R20328 gnd.n6382 gnd.n6381 0.152939
R20329 gnd.n6382 gnd.n474 0.152939
R20330 gnd.n6390 gnd.n474 0.152939
R20331 gnd.n6391 gnd.n6390 0.152939
R20332 gnd.n6392 gnd.n6391 0.152939
R20333 gnd.n6392 gnd.n468 0.152939
R20334 gnd.n6400 gnd.n468 0.152939
R20335 gnd.n6401 gnd.n6400 0.152939
R20336 gnd.n6402 gnd.n6401 0.152939
R20337 gnd.n6402 gnd.n462 0.152939
R20338 gnd.n6410 gnd.n462 0.152939
R20339 gnd.n6411 gnd.n6410 0.152939
R20340 gnd.n6412 gnd.n6411 0.152939
R20341 gnd.n6412 gnd.n456 0.152939
R20342 gnd.n6420 gnd.n456 0.152939
R20343 gnd.n6421 gnd.n6420 0.152939
R20344 gnd.n6422 gnd.n6421 0.152939
R20345 gnd.n6422 gnd.n450 0.152939
R20346 gnd.n6430 gnd.n450 0.152939
R20347 gnd.n6431 gnd.n6430 0.152939
R20348 gnd.n6432 gnd.n6431 0.152939
R20349 gnd.n6432 gnd.n444 0.152939
R20350 gnd.n6440 gnd.n444 0.152939
R20351 gnd.n6441 gnd.n6440 0.152939
R20352 gnd.n6442 gnd.n6441 0.152939
R20353 gnd.n6442 gnd.n438 0.152939
R20354 gnd.n6450 gnd.n438 0.152939
R20355 gnd.n6451 gnd.n6450 0.152939
R20356 gnd.n6452 gnd.n6451 0.152939
R20357 gnd.n6452 gnd.n432 0.152939
R20358 gnd.n6460 gnd.n432 0.152939
R20359 gnd.n6461 gnd.n6460 0.152939
R20360 gnd.n6462 gnd.n6461 0.152939
R20361 gnd.n6462 gnd.n426 0.152939
R20362 gnd.n6470 gnd.n426 0.152939
R20363 gnd.n6471 gnd.n6470 0.152939
R20364 gnd.n6472 gnd.n6471 0.152939
R20365 gnd.n6472 gnd.n420 0.152939
R20366 gnd.n6480 gnd.n420 0.152939
R20367 gnd.n6481 gnd.n6480 0.152939
R20368 gnd.n6482 gnd.n6481 0.152939
R20369 gnd.n6482 gnd.n414 0.152939
R20370 gnd.n6490 gnd.n414 0.152939
R20371 gnd.n6491 gnd.n6490 0.152939
R20372 gnd.n6492 gnd.n6491 0.152939
R20373 gnd.n6492 gnd.n408 0.152939
R20374 gnd.n6500 gnd.n408 0.152939
R20375 gnd.n6501 gnd.n6500 0.152939
R20376 gnd.n6502 gnd.n6501 0.152939
R20377 gnd.n6502 gnd.n402 0.152939
R20378 gnd.n6510 gnd.n402 0.152939
R20379 gnd.n6511 gnd.n6510 0.152939
R20380 gnd.n6512 gnd.n6511 0.152939
R20381 gnd.n6512 gnd.n396 0.152939
R20382 gnd.n6520 gnd.n396 0.152939
R20383 gnd.n6521 gnd.n6520 0.152939
R20384 gnd.n6522 gnd.n6521 0.152939
R20385 gnd.n6522 gnd.n390 0.152939
R20386 gnd.n6530 gnd.n390 0.152939
R20387 gnd.n6531 gnd.n6530 0.152939
R20388 gnd.n6532 gnd.n6531 0.152939
R20389 gnd.n6532 gnd.n384 0.152939
R20390 gnd.n6540 gnd.n384 0.152939
R20391 gnd.n6541 gnd.n6540 0.152939
R20392 gnd.n6542 gnd.n6541 0.152939
R20393 gnd.n6542 gnd.n378 0.152939
R20394 gnd.n6550 gnd.n378 0.152939
R20395 gnd.n6551 gnd.n6550 0.152939
R20396 gnd.n6552 gnd.n6551 0.152939
R20397 gnd.n6552 gnd.n372 0.152939
R20398 gnd.n6560 gnd.n372 0.152939
R20399 gnd.n6561 gnd.n6560 0.152939
R20400 gnd.n6562 gnd.n6561 0.152939
R20401 gnd.n6562 gnd.n366 0.152939
R20402 gnd.n6570 gnd.n366 0.152939
R20403 gnd.n6571 gnd.n6570 0.152939
R20404 gnd.n6572 gnd.n6571 0.152939
R20405 gnd.n6572 gnd.n360 0.152939
R20406 gnd.n6580 gnd.n360 0.152939
R20407 gnd.n6581 gnd.n6580 0.152939
R20408 gnd.n6582 gnd.n6581 0.152939
R20409 gnd.n6582 gnd.n354 0.152939
R20410 gnd.n6590 gnd.n354 0.152939
R20411 gnd.n6591 gnd.n6590 0.152939
R20412 gnd.n6592 gnd.n6591 0.152939
R20413 gnd.n6592 gnd.n348 0.152939
R20414 gnd.n6600 gnd.n348 0.152939
R20415 gnd.n6601 gnd.n6600 0.152939
R20416 gnd.n6602 gnd.n6601 0.152939
R20417 gnd.n6602 gnd.n342 0.152939
R20418 gnd.n6610 gnd.n342 0.152939
R20419 gnd.n6611 gnd.n6610 0.152939
R20420 gnd.n6612 gnd.n6611 0.152939
R20421 gnd.n6612 gnd.n336 0.152939
R20422 gnd.n6620 gnd.n336 0.152939
R20423 gnd.n6621 gnd.n6620 0.152939
R20424 gnd.n6622 gnd.n6621 0.152939
R20425 gnd.n6622 gnd.n330 0.152939
R20426 gnd.n6630 gnd.n330 0.152939
R20427 gnd.n6631 gnd.n6630 0.152939
R20428 gnd.n6632 gnd.n6631 0.152939
R20429 gnd.n6632 gnd.n324 0.152939
R20430 gnd.n6640 gnd.n324 0.152939
R20431 gnd.n6641 gnd.n6640 0.152939
R20432 gnd.n6642 gnd.n6641 0.152939
R20433 gnd.n6642 gnd.n318 0.152939
R20434 gnd.n6650 gnd.n318 0.152939
R20435 gnd.n6651 gnd.n6650 0.152939
R20436 gnd.n6653 gnd.n6651 0.152939
R20437 gnd.n6653 gnd.n6652 0.152939
R20438 gnd.n6652 gnd.n312 0.152939
R20439 gnd.n6662 gnd.n312 0.152939
R20440 gnd.n6663 gnd.n307 0.152939
R20441 gnd.n6671 gnd.n307 0.152939
R20442 gnd.n6672 gnd.n6671 0.152939
R20443 gnd.n6673 gnd.n6672 0.152939
R20444 gnd.n6673 gnd.n301 0.152939
R20445 gnd.n6681 gnd.n301 0.152939
R20446 gnd.n6682 gnd.n6681 0.152939
R20447 gnd.n6683 gnd.n6682 0.152939
R20448 gnd.n6683 gnd.n295 0.152939
R20449 gnd.n6691 gnd.n295 0.152939
R20450 gnd.n6692 gnd.n6691 0.152939
R20451 gnd.n6693 gnd.n6692 0.152939
R20452 gnd.n6693 gnd.n289 0.152939
R20453 gnd.n6701 gnd.n289 0.152939
R20454 gnd.n6702 gnd.n6701 0.152939
R20455 gnd.n6703 gnd.n6702 0.152939
R20456 gnd.n6703 gnd.n283 0.152939
R20457 gnd.n6711 gnd.n283 0.152939
R20458 gnd.n6712 gnd.n6711 0.152939
R20459 gnd.n6713 gnd.n6712 0.152939
R20460 gnd.n6713 gnd.n277 0.152939
R20461 gnd.n6721 gnd.n277 0.152939
R20462 gnd.n6722 gnd.n6721 0.152939
R20463 gnd.n6723 gnd.n6722 0.152939
R20464 gnd.n6723 gnd.n271 0.152939
R20465 gnd.n6731 gnd.n271 0.152939
R20466 gnd.n6732 gnd.n6731 0.152939
R20467 gnd.n6733 gnd.n6732 0.152939
R20468 gnd.n6733 gnd.n265 0.152939
R20469 gnd.n6741 gnd.n265 0.152939
R20470 gnd.n6742 gnd.n6741 0.152939
R20471 gnd.n6743 gnd.n6742 0.152939
R20472 gnd.n6743 gnd.n259 0.152939
R20473 gnd.n6751 gnd.n259 0.152939
R20474 gnd.n6752 gnd.n6751 0.152939
R20475 gnd.n6753 gnd.n6752 0.152939
R20476 gnd.n6753 gnd.n253 0.152939
R20477 gnd.n6761 gnd.n253 0.152939
R20478 gnd.n6762 gnd.n6761 0.152939
R20479 gnd.n6763 gnd.n6762 0.152939
R20480 gnd.n6763 gnd.n247 0.152939
R20481 gnd.n6771 gnd.n247 0.152939
R20482 gnd.n6772 gnd.n6771 0.152939
R20483 gnd.n6773 gnd.n6772 0.152939
R20484 gnd.n6773 gnd.n241 0.152939
R20485 gnd.n6781 gnd.n241 0.152939
R20486 gnd.n6782 gnd.n6781 0.152939
R20487 gnd.n6783 gnd.n6782 0.152939
R20488 gnd.n6783 gnd.n235 0.152939
R20489 gnd.n6791 gnd.n235 0.152939
R20490 gnd.n6792 gnd.n6791 0.152939
R20491 gnd.n6793 gnd.n6792 0.152939
R20492 gnd.n6793 gnd.n229 0.152939
R20493 gnd.n6801 gnd.n229 0.152939
R20494 gnd.n6802 gnd.n6801 0.152939
R20495 gnd.n6803 gnd.n6802 0.152939
R20496 gnd.n6803 gnd.n223 0.152939
R20497 gnd.n6811 gnd.n223 0.152939
R20498 gnd.n6812 gnd.n6811 0.152939
R20499 gnd.n6813 gnd.n6812 0.152939
R20500 gnd.n6813 gnd.n217 0.152939
R20501 gnd.n6821 gnd.n217 0.152939
R20502 gnd.n6822 gnd.n6821 0.152939
R20503 gnd.n6823 gnd.n6822 0.152939
R20504 gnd.n6823 gnd.n211 0.152939
R20505 gnd.n6831 gnd.n211 0.152939
R20506 gnd.n6832 gnd.n6831 0.152939
R20507 gnd.n6833 gnd.n6832 0.152939
R20508 gnd.n6833 gnd.n205 0.152939
R20509 gnd.n6841 gnd.n205 0.152939
R20510 gnd.n6842 gnd.n6841 0.152939
R20511 gnd.n6843 gnd.n6842 0.152939
R20512 gnd.n6843 gnd.n199 0.152939
R20513 gnd.n6851 gnd.n199 0.152939
R20514 gnd.n6852 gnd.n6851 0.152939
R20515 gnd.n6853 gnd.n6852 0.152939
R20516 gnd.n6853 gnd.n193 0.152939
R20517 gnd.n6861 gnd.n193 0.152939
R20518 gnd.n6862 gnd.n6861 0.152939
R20519 gnd.n6863 gnd.n6862 0.152939
R20520 gnd.n6863 gnd.n187 0.152939
R20521 gnd.n6872 gnd.n187 0.152939
R20522 gnd.n6873 gnd.n6872 0.152939
R20523 gnd.n6874 gnd.n6873 0.152939
R20524 gnd.n7298 gnd.n81 0.152939
R20525 gnd.n106 gnd.n81 0.152939
R20526 gnd.n107 gnd.n106 0.152939
R20527 gnd.n108 gnd.n107 0.152939
R20528 gnd.n124 gnd.n108 0.152939
R20529 gnd.n125 gnd.n124 0.152939
R20530 gnd.n126 gnd.n125 0.152939
R20531 gnd.n127 gnd.n126 0.152939
R20532 gnd.n144 gnd.n127 0.152939
R20533 gnd.n145 gnd.n144 0.152939
R20534 gnd.n146 gnd.n145 0.152939
R20535 gnd.n147 gnd.n146 0.152939
R20536 gnd.n162 gnd.n147 0.152939
R20537 gnd.n163 gnd.n162 0.152939
R20538 gnd.n164 gnd.n163 0.152939
R20539 gnd.n165 gnd.n164 0.152939
R20540 gnd.n7307 gnd.n69 0.152939
R20541 gnd.n176 gnd.n69 0.152939
R20542 gnd.n6894 gnd.n176 0.152939
R20543 gnd.n6895 gnd.n6894 0.152939
R20544 gnd.n6896 gnd.n6895 0.152939
R20545 gnd.n6897 gnd.n6896 0.152939
R20546 gnd.n6898 gnd.n6897 0.152939
R20547 gnd.n6899 gnd.n6898 0.152939
R20548 gnd.n6900 gnd.n6899 0.152939
R20549 gnd.n6901 gnd.n6900 0.152939
R20550 gnd.n6902 gnd.n6901 0.152939
R20551 gnd.n6903 gnd.n6902 0.152939
R20552 gnd.n6904 gnd.n6903 0.152939
R20553 gnd.n6905 gnd.n6904 0.152939
R20554 gnd.n6906 gnd.n6905 0.152939
R20555 gnd.n6907 gnd.n6906 0.152939
R20556 gnd.n6908 gnd.n6907 0.152939
R20557 gnd.n6909 gnd.n6908 0.152939
R20558 gnd.n6910 gnd.n6909 0.152939
R20559 gnd.n7191 gnd.n6910 0.152939
R20560 gnd.n6932 gnd.n6931 0.152939
R20561 gnd.n6939 gnd.n6931 0.152939
R20562 gnd.n6940 gnd.n6939 0.152939
R20563 gnd.n6941 gnd.n6940 0.152939
R20564 gnd.n6941 gnd.n6929 0.152939
R20565 gnd.n6949 gnd.n6929 0.152939
R20566 gnd.n6950 gnd.n6949 0.152939
R20567 gnd.n6951 gnd.n6950 0.152939
R20568 gnd.n6951 gnd.n6927 0.152939
R20569 gnd.n6959 gnd.n6927 0.152939
R20570 gnd.n6960 gnd.n6959 0.152939
R20571 gnd.n6961 gnd.n6960 0.152939
R20572 gnd.n6961 gnd.n6925 0.152939
R20573 gnd.n6968 gnd.n6925 0.152939
R20574 gnd.n6969 gnd.n6968 0.152939
R20575 gnd.n6970 gnd.n6969 0.152939
R20576 gnd.n6970 gnd.n6911 0.152939
R20577 gnd.n7190 gnd.n6911 0.152939
R20578 gnd.n7007 gnd.n7006 0.152939
R20579 gnd.n7008 gnd.n7007 0.152939
R20580 gnd.n7009 gnd.n7008 0.152939
R20581 gnd.n7010 gnd.n7009 0.152939
R20582 gnd.n7011 gnd.n7010 0.152939
R20583 gnd.n7012 gnd.n7011 0.152939
R20584 gnd.n7013 gnd.n7012 0.152939
R20585 gnd.n7014 gnd.n7013 0.152939
R20586 gnd.n7015 gnd.n7014 0.152939
R20587 gnd.n7016 gnd.n7015 0.152939
R20588 gnd.n7017 gnd.n7016 0.152939
R20589 gnd.n7018 gnd.n7017 0.152939
R20590 gnd.n7019 gnd.n7018 0.152939
R20591 gnd.n7020 gnd.n7019 0.152939
R20592 gnd.n7021 gnd.n7020 0.152939
R20593 gnd.n7022 gnd.n7021 0.152939
R20594 gnd.n7023 gnd.n7022 0.152939
R20595 gnd.n7024 gnd.n7023 0.152939
R20596 gnd.n7025 gnd.n7024 0.152939
R20597 gnd.n7026 gnd.n7025 0.152939
R20598 gnd.n7027 gnd.n7026 0.152939
R20599 gnd.n7028 gnd.n7027 0.152939
R20600 gnd.n7029 gnd.n7028 0.152939
R20601 gnd.n7030 gnd.n7029 0.152939
R20602 gnd.n7031 gnd.n7030 0.152939
R20603 gnd.n7032 gnd.n7031 0.152939
R20604 gnd.n7033 gnd.n7032 0.152939
R20605 gnd.n7034 gnd.n7033 0.152939
R20606 gnd.n7035 gnd.n7034 0.152939
R20607 gnd.n7036 gnd.n7035 0.152939
R20608 gnd.n7037 gnd.n7036 0.152939
R20609 gnd.n7038 gnd.n7037 0.152939
R20610 gnd.n7039 gnd.n7038 0.152939
R20611 gnd.n7040 gnd.n7039 0.152939
R20612 gnd.n7041 gnd.n7040 0.152939
R20613 gnd.n7042 gnd.n7041 0.152939
R20614 gnd.n7110 gnd.n7042 0.152939
R20615 gnd.n7110 gnd.n7109 0.152939
R20616 gnd.n7109 gnd.n7108 0.152939
R20617 gnd.n7108 gnd.n7046 0.152939
R20618 gnd.n7047 gnd.n7046 0.152939
R20619 gnd.n7048 gnd.n7047 0.152939
R20620 gnd.n7049 gnd.n7048 0.152939
R20621 gnd.n7050 gnd.n7049 0.152939
R20622 gnd.n7051 gnd.n7050 0.152939
R20623 gnd.n7052 gnd.n7051 0.152939
R20624 gnd.n7053 gnd.n7052 0.152939
R20625 gnd.n7054 gnd.n7053 0.152939
R20626 gnd.n7055 gnd.n7054 0.152939
R20627 gnd.n7056 gnd.n7055 0.152939
R20628 gnd.n7057 gnd.n7056 0.152939
R20629 gnd.n7058 gnd.n7057 0.152939
R20630 gnd.n7059 gnd.n7058 0.152939
R20631 gnd.n7060 gnd.n7059 0.152939
R20632 gnd.n7061 gnd.n7060 0.152939
R20633 gnd.n7062 gnd.n7061 0.152939
R20634 gnd.n7068 gnd.n7062 0.152939
R20635 gnd.n7068 gnd.n7067 0.152939
R20636 gnd.n1428 gnd.n1427 0.152939
R20637 gnd.n1429 gnd.n1428 0.152939
R20638 gnd.n1430 gnd.n1429 0.152939
R20639 gnd.n1431 gnd.n1430 0.152939
R20640 gnd.n1432 gnd.n1431 0.152939
R20641 gnd.n1433 gnd.n1432 0.152939
R20642 gnd.n1434 gnd.n1433 0.152939
R20643 gnd.n1435 gnd.n1434 0.152939
R20644 gnd.n1436 gnd.n1435 0.152939
R20645 gnd.n1437 gnd.n1436 0.152939
R20646 gnd.n1438 gnd.n1437 0.152939
R20647 gnd.n1439 gnd.n1438 0.152939
R20648 gnd.n1440 gnd.n1439 0.152939
R20649 gnd.n1441 gnd.n1440 0.152939
R20650 gnd.n1442 gnd.n1441 0.152939
R20651 gnd.n1443 gnd.n1442 0.152939
R20652 gnd.n1444 gnd.n1443 0.152939
R20653 gnd.n1447 gnd.n1444 0.152939
R20654 gnd.n1448 gnd.n1447 0.152939
R20655 gnd.n1449 gnd.n1448 0.152939
R20656 gnd.n1450 gnd.n1449 0.152939
R20657 gnd.n1451 gnd.n1450 0.152939
R20658 gnd.n1452 gnd.n1451 0.152939
R20659 gnd.n1453 gnd.n1452 0.152939
R20660 gnd.n1454 gnd.n1453 0.152939
R20661 gnd.n1459 gnd.n1458 0.152939
R20662 gnd.n1460 gnd.n1459 0.152939
R20663 gnd.n1461 gnd.n1460 0.152939
R20664 gnd.n1462 gnd.n1461 0.152939
R20665 gnd.n1463 gnd.n1462 0.152939
R20666 gnd.n1464 gnd.n1463 0.152939
R20667 gnd.n1465 gnd.n1464 0.152939
R20668 gnd.n1466 gnd.n1465 0.152939
R20669 gnd.n1467 gnd.n1466 0.152939
R20670 gnd.n1470 gnd.n1467 0.152939
R20671 gnd.n1471 gnd.n1470 0.152939
R20672 gnd.n1472 gnd.n1471 0.152939
R20673 gnd.n1473 gnd.n1472 0.152939
R20674 gnd.n1474 gnd.n1473 0.152939
R20675 gnd.n1475 gnd.n1474 0.152939
R20676 gnd.n1476 gnd.n1475 0.152939
R20677 gnd.n1477 gnd.n1476 0.152939
R20678 gnd.n1478 gnd.n1477 0.152939
R20679 gnd.n1479 gnd.n1478 0.152939
R20680 gnd.n1480 gnd.n1479 0.152939
R20681 gnd.n1481 gnd.n1480 0.152939
R20682 gnd.n1482 gnd.n1481 0.152939
R20683 gnd.n1483 gnd.n1482 0.152939
R20684 gnd.n1484 gnd.n1483 0.152939
R20685 gnd.n1485 gnd.n1484 0.152939
R20686 gnd.n1486 gnd.n1485 0.152939
R20687 gnd.n1487 gnd.n1486 0.152939
R20688 gnd.n1488 gnd.n1487 0.152939
R20689 gnd.n5472 gnd.n1488 0.152939
R20690 gnd.n5472 gnd.n5471 0.152939
R20691 gnd.n1509 gnd.n1508 0.152939
R20692 gnd.n1510 gnd.n1509 0.152939
R20693 gnd.n1511 gnd.n1510 0.152939
R20694 gnd.n1512 gnd.n1511 0.152939
R20695 gnd.n1532 gnd.n1512 0.152939
R20696 gnd.n1533 gnd.n1532 0.152939
R20697 gnd.n1534 gnd.n1533 0.152939
R20698 gnd.n1535 gnd.n1534 0.152939
R20699 gnd.n1553 gnd.n1535 0.152939
R20700 gnd.n1554 gnd.n1553 0.152939
R20701 gnd.n1555 gnd.n1554 0.152939
R20702 gnd.n1556 gnd.n1555 0.152939
R20703 gnd.n1572 gnd.n1556 0.152939
R20704 gnd.n1573 gnd.n1572 0.152939
R20705 gnd.n1573 gnd.n82 0.152939
R20706 gnd.n7298 gnd.n82 0.152939
R20707 gnd.n4165 gnd.n4164 0.152939
R20708 gnd.n4166 gnd.n4165 0.152939
R20709 gnd.n4166 gnd.n2130 0.152939
R20710 gnd.n4223 gnd.n2130 0.152939
R20711 gnd.n4224 gnd.n4223 0.152939
R20712 gnd.n4225 gnd.n4224 0.152939
R20713 gnd.n4225 gnd.n2126 0.152939
R20714 gnd.n4231 gnd.n2126 0.152939
R20715 gnd.n4232 gnd.n4231 0.152939
R20716 gnd.n4233 gnd.n4232 0.152939
R20717 gnd.n4233 gnd.n2122 0.152939
R20718 gnd.n4239 gnd.n2122 0.152939
R20719 gnd.n4240 gnd.n4239 0.152939
R20720 gnd.n4241 gnd.n4240 0.152939
R20721 gnd.n4241 gnd.n2118 0.152939
R20722 gnd.n4247 gnd.n2118 0.152939
R20723 gnd.n4248 gnd.n4247 0.152939
R20724 gnd.n4249 gnd.n4248 0.152939
R20725 gnd.n4249 gnd.n2114 0.152939
R20726 gnd.n4256 gnd.n2114 0.152939
R20727 gnd.n4257 gnd.n4256 0.152939
R20728 gnd.n4258 gnd.n4257 0.152939
R20729 gnd.n4258 gnd.n2108 0.152939
R20730 gnd.n4324 gnd.n2108 0.152939
R20731 gnd.n4325 gnd.n4324 0.152939
R20732 gnd.n4326 gnd.n4325 0.152939
R20733 gnd.n4326 gnd.n2094 0.152939
R20734 gnd.n4340 gnd.n2094 0.152939
R20735 gnd.n4341 gnd.n4340 0.152939
R20736 gnd.n4342 gnd.n4341 0.152939
R20737 gnd.n4342 gnd.n2079 0.152939
R20738 gnd.n4356 gnd.n2079 0.152939
R20739 gnd.n4357 gnd.n4356 0.152939
R20740 gnd.n4358 gnd.n4357 0.152939
R20741 gnd.n4358 gnd.n2065 0.152939
R20742 gnd.n4372 gnd.n2065 0.152939
R20743 gnd.n4373 gnd.n4372 0.152939
R20744 gnd.n4374 gnd.n4373 0.152939
R20745 gnd.n4374 gnd.n2050 0.152939
R20746 gnd.n4402 gnd.n2050 0.152939
R20747 gnd.n4403 gnd.n4402 0.152939
R20748 gnd.n4404 gnd.n4403 0.152939
R20749 gnd.n4405 gnd.n4404 0.152939
R20750 gnd.n4407 gnd.n4405 0.152939
R20751 gnd.n4407 gnd.n4406 0.152939
R20752 gnd.n4406 gnd.n1208 0.152939
R20753 gnd.n1209 gnd.n1208 0.152939
R20754 gnd.n1210 gnd.n1209 0.152939
R20755 gnd.n4560 gnd.n1210 0.152939
R20756 gnd.n4561 gnd.n4560 0.152939
R20757 gnd.n4562 gnd.n4561 0.152939
R20758 gnd.n4562 gnd.n2020 0.152939
R20759 gnd.n4589 gnd.n2020 0.152939
R20760 gnd.n4590 gnd.n4589 0.152939
R20761 gnd.n4591 gnd.n4590 0.152939
R20762 gnd.n4592 gnd.n4591 0.152939
R20763 gnd.n4592 gnd.n1992 0.152939
R20764 gnd.n4627 gnd.n1992 0.152939
R20765 gnd.n4628 gnd.n4627 0.152939
R20766 gnd.n4629 gnd.n4628 0.152939
R20767 gnd.n4630 gnd.n4629 0.152939
R20768 gnd.n4632 gnd.n4630 0.152939
R20769 gnd.n4632 gnd.n4631 0.152939
R20770 gnd.n4631 gnd.n1966 0.152939
R20771 gnd.n1967 gnd.n1966 0.152939
R20772 gnd.n1968 gnd.n1967 0.152939
R20773 gnd.n1968 gnd.n1942 0.152939
R20774 gnd.n4728 gnd.n1942 0.152939
R20775 gnd.n4729 gnd.n4728 0.152939
R20776 gnd.n4730 gnd.n4729 0.152939
R20777 gnd.n4731 gnd.n4730 0.152939
R20778 gnd.n4731 gnd.n1914 0.152939
R20779 gnd.n4766 gnd.n1914 0.152939
R20780 gnd.n4767 gnd.n4766 0.152939
R20781 gnd.n4768 gnd.n4767 0.152939
R20782 gnd.n4768 gnd.n1888 0.152939
R20783 gnd.n4803 gnd.n1888 0.152939
R20784 gnd.n4804 gnd.n4803 0.152939
R20785 gnd.n4805 gnd.n4804 0.152939
R20786 gnd.n4806 gnd.n4805 0.152939
R20787 gnd.n4806 gnd.n1861 0.152939
R20788 gnd.n4852 gnd.n1861 0.152939
R20789 gnd.n4853 gnd.n4852 0.152939
R20790 gnd.n4854 gnd.n4853 0.152939
R20791 gnd.n4855 gnd.n4854 0.152939
R20792 gnd.n4855 gnd.n1839 0.152939
R20793 gnd.n4893 gnd.n1839 0.152939
R20794 gnd.n4894 gnd.n4893 0.152939
R20795 gnd.n4895 gnd.n4894 0.152939
R20796 gnd.n4896 gnd.n4895 0.152939
R20797 gnd.n4896 gnd.n1809 0.152939
R20798 gnd.n4933 gnd.n1809 0.152939
R20799 gnd.n4934 gnd.n4933 0.152939
R20800 gnd.n4935 gnd.n4934 0.152939
R20801 gnd.n4935 gnd.n1785 0.152939
R20802 gnd.n4976 gnd.n1785 0.152939
R20803 gnd.n4977 gnd.n4976 0.152939
R20804 gnd.n4978 gnd.n4977 0.152939
R20805 gnd.n4979 gnd.n4978 0.152939
R20806 gnd.n4979 gnd.n1729 0.152939
R20807 gnd.n5152 gnd.n1729 0.152939
R20808 gnd.n5153 gnd.n5152 0.152939
R20809 gnd.n5154 gnd.n5153 0.152939
R20810 gnd.n5154 gnd.n1718 0.152939
R20811 gnd.n5169 gnd.n1718 0.152939
R20812 gnd.n5170 gnd.n5169 0.152939
R20813 gnd.n5171 gnd.n5170 0.152939
R20814 gnd.n5171 gnd.n1706 0.152939
R20815 gnd.n5186 gnd.n1706 0.152939
R20816 gnd.n5187 gnd.n5186 0.152939
R20817 gnd.n5188 gnd.n5187 0.152939
R20818 gnd.n5188 gnd.n1694 0.152939
R20819 gnd.n5203 gnd.n1694 0.152939
R20820 gnd.n5204 gnd.n5203 0.152939
R20821 gnd.n5205 gnd.n5204 0.152939
R20822 gnd.n5205 gnd.n1682 0.152939
R20823 gnd.n5220 gnd.n1682 0.152939
R20824 gnd.n5221 gnd.n5220 0.152939
R20825 gnd.n5222 gnd.n5221 0.152939
R20826 gnd.n5224 gnd.n5222 0.152939
R20827 gnd.n5224 gnd.n5223 0.152939
R20828 gnd.n5223 gnd.n1670 0.152939
R20829 gnd.n5242 gnd.n1670 0.152939
R20830 gnd.n5243 gnd.n5242 0.152939
R20831 gnd.n5244 gnd.n5243 0.152939
R20832 gnd.n5245 gnd.n5244 0.152939
R20833 gnd.n5246 gnd.n5245 0.152939
R20834 gnd.n5248 gnd.n5246 0.152939
R20835 gnd.n5249 gnd.n5248 0.152939
R20836 gnd.n5249 gnd.n1634 0.152939
R20837 gnd.n5311 gnd.n1634 0.152939
R20838 gnd.n5312 gnd.n5311 0.152939
R20839 gnd.n5313 gnd.n5312 0.152939
R20840 gnd.n5313 gnd.n1630 0.152939
R20841 gnd.n5319 gnd.n1630 0.152939
R20842 gnd.n5320 gnd.n5319 0.152939
R20843 gnd.n5321 gnd.n5320 0.152939
R20844 gnd.n5321 gnd.n1626 0.152939
R20845 gnd.n5327 gnd.n1626 0.152939
R20846 gnd.n5328 gnd.n5327 0.152939
R20847 gnd.n5329 gnd.n5328 0.152939
R20848 gnd.n5330 gnd.n5329 0.152939
R20849 gnd.n5331 gnd.n5330 0.152939
R20850 gnd.n5334 gnd.n5331 0.152939
R20851 gnd.n5335 gnd.n5334 0.152939
R20852 gnd.n3775 gnd.n3774 0.152939
R20853 gnd.n3776 gnd.n3775 0.152939
R20854 gnd.n3776 gnd.n2218 0.152939
R20855 gnd.n4028 gnd.n2218 0.152939
R20856 gnd.n4029 gnd.n4028 0.152939
R20857 gnd.n4030 gnd.n4029 0.152939
R20858 gnd.n4031 gnd.n4030 0.152939
R20859 gnd.n4031 gnd.n2193 0.152939
R20860 gnd.n4063 gnd.n2193 0.152939
R20861 gnd.n4064 gnd.n4063 0.152939
R20862 gnd.n4065 gnd.n4064 0.152939
R20863 gnd.n4066 gnd.n4065 0.152939
R20864 gnd.n4067 gnd.n4066 0.152939
R20865 gnd.n4067 gnd.n2167 0.152939
R20866 gnd.n4103 gnd.n2167 0.152939
R20867 gnd.n4104 gnd.n4103 0.152939
R20868 gnd.n4105 gnd.n4104 0.152939
R20869 gnd.n4105 gnd.n2162 0.152939
R20870 gnd.n4129 gnd.n2162 0.152939
R20871 gnd.n4130 gnd.n4129 0.152939
R20872 gnd.n3726 gnd.n3725 0.152939
R20873 gnd.n3734 gnd.n3725 0.152939
R20874 gnd.n3735 gnd.n3734 0.152939
R20875 gnd.n3736 gnd.n3735 0.152939
R20876 gnd.n3736 gnd.n3721 0.152939
R20877 gnd.n3744 gnd.n3721 0.152939
R20878 gnd.n3745 gnd.n3744 0.152939
R20879 gnd.n3746 gnd.n3745 0.152939
R20880 gnd.n3746 gnd.n3717 0.152939
R20881 gnd.n3754 gnd.n3717 0.152939
R20882 gnd.n3755 gnd.n3754 0.152939
R20883 gnd.n3756 gnd.n3755 0.152939
R20884 gnd.n3756 gnd.n3713 0.152939
R20885 gnd.n3764 gnd.n3713 0.152939
R20886 gnd.n3765 gnd.n3764 0.152939
R20887 gnd.n3766 gnd.n3765 0.152939
R20888 gnd.n3766 gnd.n3707 0.152939
R20889 gnd.n3773 gnd.n3707 0.152939
R20890 gnd.n794 gnd.n741 0.152939
R20891 gnd.n795 gnd.n794 0.152939
R20892 gnd.n796 gnd.n795 0.152939
R20893 gnd.n797 gnd.n796 0.152939
R20894 gnd.n814 gnd.n797 0.152939
R20895 gnd.n815 gnd.n814 0.152939
R20896 gnd.n816 gnd.n815 0.152939
R20897 gnd.n817 gnd.n816 0.152939
R20898 gnd.n834 gnd.n817 0.152939
R20899 gnd.n835 gnd.n834 0.152939
R20900 gnd.n836 gnd.n835 0.152939
R20901 gnd.n837 gnd.n836 0.152939
R20902 gnd.n854 gnd.n837 0.152939
R20903 gnd.n855 gnd.n854 0.152939
R20904 gnd.n856 gnd.n855 0.152939
R20905 gnd.n857 gnd.n856 0.152939
R20906 gnd.n1013 gnd.n1012 0.152939
R20907 gnd.n1014 gnd.n1013 0.152939
R20908 gnd.n1015 gnd.n1014 0.152939
R20909 gnd.n1016 gnd.n1015 0.152939
R20910 gnd.n1017 gnd.n1016 0.152939
R20911 gnd.n1018 gnd.n1017 0.152939
R20912 gnd.n1019 gnd.n1018 0.152939
R20913 gnd.n1020 gnd.n1019 0.152939
R20914 gnd.n1021 gnd.n1020 0.152939
R20915 gnd.n1022 gnd.n1021 0.152939
R20916 gnd.n1023 gnd.n1022 0.152939
R20917 gnd.n1024 gnd.n1023 0.152939
R20918 gnd.n1025 gnd.n1024 0.152939
R20919 gnd.n1026 gnd.n1025 0.152939
R20920 gnd.n1027 gnd.n1026 0.152939
R20921 gnd.n1028 gnd.n1027 0.152939
R20922 gnd.n1029 gnd.n1028 0.152939
R20923 gnd.n1032 gnd.n1029 0.152939
R20924 gnd.n1033 gnd.n1032 0.152939
R20925 gnd.n1034 gnd.n1033 0.152939
R20926 gnd.n1035 gnd.n1034 0.152939
R20927 gnd.n1036 gnd.n1035 0.152939
R20928 gnd.n1037 gnd.n1036 0.152939
R20929 gnd.n1038 gnd.n1037 0.152939
R20930 gnd.n1039 gnd.n1038 0.152939
R20931 gnd.n1137 gnd.n1136 0.152939
R20932 gnd.n1136 gnd.n1042 0.152939
R20933 gnd.n1043 gnd.n1042 0.152939
R20934 gnd.n1044 gnd.n1043 0.152939
R20935 gnd.n1045 gnd.n1044 0.152939
R20936 gnd.n1046 gnd.n1045 0.152939
R20937 gnd.n1047 gnd.n1046 0.152939
R20938 gnd.n1048 gnd.n1047 0.152939
R20939 gnd.n1116 gnd.n1048 0.152939
R20940 gnd.n1116 gnd.n1115 0.152939
R20941 gnd.n1115 gnd.n1114 0.152939
R20942 gnd.n1114 gnd.n1052 0.152939
R20943 gnd.n1053 gnd.n1052 0.152939
R20944 gnd.n1054 gnd.n1053 0.152939
R20945 gnd.n1055 gnd.n1054 0.152939
R20946 gnd.n1056 gnd.n1055 0.152939
R20947 gnd.n1057 gnd.n1056 0.152939
R20948 gnd.n1058 gnd.n1057 0.152939
R20949 gnd.n1059 gnd.n1058 0.152939
R20950 gnd.n1060 gnd.n1059 0.152939
R20951 gnd.n1061 gnd.n1060 0.152939
R20952 gnd.n1062 gnd.n1061 0.152939
R20953 gnd.n1063 gnd.n1062 0.152939
R20954 gnd.n1064 gnd.n1063 0.152939
R20955 gnd.n1065 gnd.n1064 0.152939
R20956 gnd.n1066 gnd.n1065 0.152939
R20957 gnd.n1067 gnd.n1066 0.152939
R20958 gnd.n1068 gnd.n1067 0.152939
R20959 gnd.n1074 gnd.n1068 0.152939
R20960 gnd.n1074 gnd.n1073 0.152939
R20961 gnd.n3993 gnd.n3782 0.152939
R20962 gnd.n3785 gnd.n3782 0.152939
R20963 gnd.n3786 gnd.n3785 0.152939
R20964 gnd.n3787 gnd.n3786 0.152939
R20965 gnd.n3790 gnd.n3787 0.152939
R20966 gnd.n3791 gnd.n3790 0.152939
R20967 gnd.n3792 gnd.n3791 0.152939
R20968 gnd.n3793 gnd.n3792 0.152939
R20969 gnd.n3796 gnd.n3793 0.152939
R20970 gnd.n3797 gnd.n3796 0.152939
R20971 gnd.n3798 gnd.n3797 0.152939
R20972 gnd.n3799 gnd.n3798 0.152939
R20973 gnd.n3802 gnd.n3799 0.152939
R20974 gnd.n3803 gnd.n3802 0.152939
R20975 gnd.n3804 gnd.n3803 0.152939
R20976 gnd.n3805 gnd.n3804 0.152939
R20977 gnd.n3811 gnd.n3805 0.152939
R20978 gnd.n3812 gnd.n3811 0.152939
R20979 gnd.n3813 gnd.n3812 0.152939
R20980 gnd.n3814 gnd.n3813 0.152939
R20981 gnd.n3817 gnd.n3814 0.152939
R20982 gnd.n3818 gnd.n3817 0.152939
R20983 gnd.n3819 gnd.n3818 0.152939
R20984 gnd.n3820 gnd.n3819 0.152939
R20985 gnd.n3823 gnd.n3820 0.152939
R20986 gnd.n3824 gnd.n3823 0.152939
R20987 gnd.n3825 gnd.n3824 0.152939
R20988 gnd.n3826 gnd.n3825 0.152939
R20989 gnd.n3829 gnd.n3826 0.152939
R20990 gnd.n3830 gnd.n3829 0.152939
R20991 gnd.n3831 gnd.n3830 0.152939
R20992 gnd.n3832 gnd.n3831 0.152939
R20993 gnd.n3835 gnd.n3832 0.152939
R20994 gnd.n3836 gnd.n3835 0.152939
R20995 gnd.n3837 gnd.n3836 0.152939
R20996 gnd.n3838 gnd.n3837 0.152939
R20997 gnd.n3843 gnd.n3838 0.152939
R20998 gnd.n3844 gnd.n3843 0.152939
R20999 gnd.n3845 gnd.n3844 0.152939
R21000 gnd.n3846 gnd.n3845 0.152939
R21001 gnd.n3849 gnd.n3846 0.152939
R21002 gnd.n3850 gnd.n3849 0.152939
R21003 gnd.n3851 gnd.n3850 0.152939
R21004 gnd.n3852 gnd.n3851 0.152939
R21005 gnd.n3855 gnd.n3852 0.152939
R21006 gnd.n3856 gnd.n3855 0.152939
R21007 gnd.n3857 gnd.n3856 0.152939
R21008 gnd.n3858 gnd.n3857 0.152939
R21009 gnd.n3861 gnd.n3858 0.152939
R21010 gnd.n3862 gnd.n3861 0.152939
R21011 gnd.n3863 gnd.n3862 0.152939
R21012 gnd.n3864 gnd.n3863 0.152939
R21013 gnd.n3867 gnd.n3864 0.152939
R21014 gnd.n3868 gnd.n3867 0.152939
R21015 gnd.n3869 gnd.n3868 0.152939
R21016 gnd.n3870 gnd.n3869 0.152939
R21017 gnd.n3874 gnd.n3870 0.152939
R21018 gnd.n3875 gnd.n3874 0.152939
R21019 gnd.n3994 gnd.n2227 0.152939
R21020 gnd.n4018 gnd.n2227 0.152939
R21021 gnd.n4019 gnd.n4018 0.152939
R21022 gnd.n4020 gnd.n4019 0.152939
R21023 gnd.n4021 gnd.n4020 0.152939
R21024 gnd.n4021 gnd.n2202 0.152939
R21025 gnd.n4053 gnd.n2202 0.152939
R21026 gnd.n4054 gnd.n4053 0.152939
R21027 gnd.n4055 gnd.n4054 0.152939
R21028 gnd.n4056 gnd.n4055 0.152939
R21029 gnd.n4056 gnd.n2175 0.152939
R21030 gnd.n4093 gnd.n2175 0.152939
R21031 gnd.n4094 gnd.n4093 0.152939
R21032 gnd.n4096 gnd.n4094 0.152939
R21033 gnd.n4096 gnd.n4095 0.152939
R21034 gnd.n4095 gnd.n741 0.152939
R21035 gnd.n6241 gnd.n563 0.152939
R21036 gnd.n568 gnd.n563 0.152939
R21037 gnd.n569 gnd.n568 0.152939
R21038 gnd.n570 gnd.n569 0.152939
R21039 gnd.n571 gnd.n570 0.152939
R21040 gnd.n576 gnd.n571 0.152939
R21041 gnd.n577 gnd.n576 0.152939
R21042 gnd.n578 gnd.n577 0.152939
R21043 gnd.n579 gnd.n578 0.152939
R21044 gnd.n584 gnd.n579 0.152939
R21045 gnd.n585 gnd.n584 0.152939
R21046 gnd.n586 gnd.n585 0.152939
R21047 gnd.n587 gnd.n586 0.152939
R21048 gnd.n592 gnd.n587 0.152939
R21049 gnd.n593 gnd.n592 0.152939
R21050 gnd.n594 gnd.n593 0.152939
R21051 gnd.n595 gnd.n594 0.152939
R21052 gnd.n600 gnd.n595 0.152939
R21053 gnd.n601 gnd.n600 0.152939
R21054 gnd.n602 gnd.n601 0.152939
R21055 gnd.n603 gnd.n602 0.152939
R21056 gnd.n608 gnd.n603 0.152939
R21057 gnd.n609 gnd.n608 0.152939
R21058 gnd.n610 gnd.n609 0.152939
R21059 gnd.n611 gnd.n610 0.152939
R21060 gnd.n616 gnd.n611 0.152939
R21061 gnd.n617 gnd.n616 0.152939
R21062 gnd.n618 gnd.n617 0.152939
R21063 gnd.n619 gnd.n618 0.152939
R21064 gnd.n624 gnd.n619 0.152939
R21065 gnd.n625 gnd.n624 0.152939
R21066 gnd.n626 gnd.n625 0.152939
R21067 gnd.n627 gnd.n626 0.152939
R21068 gnd.n632 gnd.n627 0.152939
R21069 gnd.n633 gnd.n632 0.152939
R21070 gnd.n634 gnd.n633 0.152939
R21071 gnd.n635 gnd.n634 0.152939
R21072 gnd.n640 gnd.n635 0.152939
R21073 gnd.n641 gnd.n640 0.152939
R21074 gnd.n642 gnd.n641 0.152939
R21075 gnd.n643 gnd.n642 0.152939
R21076 gnd.n648 gnd.n643 0.152939
R21077 gnd.n649 gnd.n648 0.152939
R21078 gnd.n650 gnd.n649 0.152939
R21079 gnd.n651 gnd.n650 0.152939
R21080 gnd.n656 gnd.n651 0.152939
R21081 gnd.n657 gnd.n656 0.152939
R21082 gnd.n658 gnd.n657 0.152939
R21083 gnd.n659 gnd.n658 0.152939
R21084 gnd.n664 gnd.n659 0.152939
R21085 gnd.n665 gnd.n664 0.152939
R21086 gnd.n666 gnd.n665 0.152939
R21087 gnd.n667 gnd.n666 0.152939
R21088 gnd.n672 gnd.n667 0.152939
R21089 gnd.n673 gnd.n672 0.152939
R21090 gnd.n674 gnd.n673 0.152939
R21091 gnd.n675 gnd.n674 0.152939
R21092 gnd.n680 gnd.n675 0.152939
R21093 gnd.n681 gnd.n680 0.152939
R21094 gnd.n682 gnd.n681 0.152939
R21095 gnd.n683 gnd.n682 0.152939
R21096 gnd.n688 gnd.n683 0.152939
R21097 gnd.n689 gnd.n688 0.152939
R21098 gnd.n690 gnd.n689 0.152939
R21099 gnd.n691 gnd.n690 0.152939
R21100 gnd.n696 gnd.n691 0.152939
R21101 gnd.n697 gnd.n696 0.152939
R21102 gnd.n698 gnd.n697 0.152939
R21103 gnd.n699 gnd.n698 0.152939
R21104 gnd.n704 gnd.n699 0.152939
R21105 gnd.n705 gnd.n704 0.152939
R21106 gnd.n706 gnd.n705 0.152939
R21107 gnd.n707 gnd.n706 0.152939
R21108 gnd.n712 gnd.n707 0.152939
R21109 gnd.n713 gnd.n712 0.152939
R21110 gnd.n714 gnd.n713 0.152939
R21111 gnd.n715 gnd.n714 0.152939
R21112 gnd.n720 gnd.n715 0.152939
R21113 gnd.n721 gnd.n720 0.152939
R21114 gnd.n722 gnd.n721 0.152939
R21115 gnd.n723 gnd.n722 0.152939
R21116 gnd.n728 gnd.n723 0.152939
R21117 gnd.n729 gnd.n728 0.152939
R21118 gnd.n6071 gnd.n729 0.152939
R21119 gnd.n4317 gnd.n4316 0.152939
R21120 gnd.n4318 gnd.n4317 0.152939
R21121 gnd.n4318 gnd.n2101 0.152939
R21122 gnd.n4332 gnd.n2101 0.152939
R21123 gnd.n4333 gnd.n4332 0.152939
R21124 gnd.n4334 gnd.n4333 0.152939
R21125 gnd.n4334 gnd.n2087 0.152939
R21126 gnd.n4348 gnd.n2087 0.152939
R21127 gnd.n4349 gnd.n4348 0.152939
R21128 gnd.n4350 gnd.n4349 0.152939
R21129 gnd.n4350 gnd.n2073 0.152939
R21130 gnd.n4364 gnd.n2073 0.152939
R21131 gnd.n4365 gnd.n4364 0.152939
R21132 gnd.n4366 gnd.n4365 0.152939
R21133 gnd.n4366 gnd.n2059 0.152939
R21134 gnd.n4380 gnd.n2059 0.152939
R21135 gnd.n4381 gnd.n4380 0.152939
R21136 gnd.n4396 gnd.n4381 0.152939
R21137 gnd.n4396 gnd.n4395 0.152939
R21138 gnd.n4395 gnd.n4394 0.152939
R21139 gnd.n4394 gnd.n4382 0.152939
R21140 gnd.n4390 gnd.n4382 0.152939
R21141 gnd.n4390 gnd.n4389 0.152939
R21142 gnd.n4389 gnd.n4388 0.152939
R21143 gnd.n4388 gnd.n1218 0.152939
R21144 gnd.n5768 gnd.n1218 0.152939
R21145 gnd.n5768 gnd.n5767 0.152939
R21146 gnd.n5767 gnd.n5766 0.152939
R21147 gnd.n5766 gnd.n1219 0.152939
R21148 gnd.n5762 gnd.n1219 0.152939
R21149 gnd.n5762 gnd.n5761 0.152939
R21150 gnd.n5761 gnd.n5760 0.152939
R21151 gnd.n5760 gnd.n1224 0.152939
R21152 gnd.n5756 gnd.n1224 0.152939
R21153 gnd.n5756 gnd.n5755 0.152939
R21154 gnd.n5755 gnd.n5754 0.152939
R21155 gnd.n5754 gnd.n1229 0.152939
R21156 gnd.n5750 gnd.n1229 0.152939
R21157 gnd.n5750 gnd.n5749 0.152939
R21158 gnd.n5749 gnd.n5748 0.152939
R21159 gnd.n5748 gnd.n1234 0.152939
R21160 gnd.n5744 gnd.n1234 0.152939
R21161 gnd.n5744 gnd.n5743 0.152939
R21162 gnd.n5743 gnd.n5742 0.152939
R21163 gnd.n5742 gnd.n1239 0.152939
R21164 gnd.n5738 gnd.n1239 0.152939
R21165 gnd.n5738 gnd.n5737 0.152939
R21166 gnd.n5737 gnd.n5736 0.152939
R21167 gnd.n5736 gnd.n1244 0.152939
R21168 gnd.n5732 gnd.n1244 0.152939
R21169 gnd.n5732 gnd.n5731 0.152939
R21170 gnd.n5731 gnd.n5730 0.152939
R21171 gnd.n5730 gnd.n1249 0.152939
R21172 gnd.n5726 gnd.n1249 0.152939
R21173 gnd.n5726 gnd.n5725 0.152939
R21174 gnd.n5725 gnd.n5724 0.152939
R21175 gnd.n5724 gnd.n1254 0.152939
R21176 gnd.n5720 gnd.n1254 0.152939
R21177 gnd.n5720 gnd.n5719 0.152939
R21178 gnd.n5719 gnd.n5718 0.152939
R21179 gnd.n5718 gnd.n1259 0.152939
R21180 gnd.n5714 gnd.n1259 0.152939
R21181 gnd.n5714 gnd.n5713 0.152939
R21182 gnd.n5713 gnd.n5712 0.152939
R21183 gnd.n5712 gnd.n1264 0.152939
R21184 gnd.n5708 gnd.n1264 0.152939
R21185 gnd.n5708 gnd.n5707 0.152939
R21186 gnd.n5707 gnd.n5706 0.152939
R21187 gnd.n5706 gnd.n1269 0.152939
R21188 gnd.n5702 gnd.n1269 0.152939
R21189 gnd.n5702 gnd.n5701 0.152939
R21190 gnd.n5701 gnd.n5700 0.152939
R21191 gnd.n5700 gnd.n1274 0.152939
R21192 gnd.n5696 gnd.n1274 0.152939
R21193 gnd.n5696 gnd.n5695 0.152939
R21194 gnd.n5695 gnd.n5694 0.152939
R21195 gnd.n5694 gnd.n1279 0.152939
R21196 gnd.n5690 gnd.n1279 0.152939
R21197 gnd.n5690 gnd.n5689 0.152939
R21198 gnd.n5689 gnd.n5688 0.152939
R21199 gnd.n5688 gnd.n1284 0.152939
R21200 gnd.n5684 gnd.n1284 0.152939
R21201 gnd.n5684 gnd.n5683 0.152939
R21202 gnd.n5683 gnd.n5682 0.152939
R21203 gnd.n5682 gnd.n1289 0.152939
R21204 gnd.n5678 gnd.n1289 0.152939
R21205 gnd.n5678 gnd.n5677 0.152939
R21206 gnd.n5677 gnd.n5676 0.152939
R21207 gnd.n5676 gnd.n1294 0.152939
R21208 gnd.n5672 gnd.n1294 0.152939
R21209 gnd.n5672 gnd.n5671 0.152939
R21210 gnd.n5671 gnd.n5670 0.152939
R21211 gnd.n5670 gnd.n1299 0.152939
R21212 gnd.n5666 gnd.n1299 0.152939
R21213 gnd.n5666 gnd.n5665 0.152939
R21214 gnd.n5665 gnd.n5664 0.152939
R21215 gnd.n5664 gnd.n1304 0.152939
R21216 gnd.n5660 gnd.n1304 0.152939
R21217 gnd.n5660 gnd.n5659 0.152939
R21218 gnd.n5659 gnd.n5658 0.152939
R21219 gnd.n5658 gnd.n1309 0.152939
R21220 gnd.n4150 gnd.n2158 0.152939
R21221 gnd.n4150 gnd.n4149 0.152939
R21222 gnd.n4149 gnd.n4148 0.152939
R21223 gnd.n4148 gnd.n2146 0.152939
R21224 gnd.n4174 gnd.n2146 0.152939
R21225 gnd.n4175 gnd.n4174 0.152939
R21226 gnd.n4176 gnd.n4175 0.152939
R21227 gnd.n4176 gnd.n2136 0.152939
R21228 gnd.n4216 gnd.n2136 0.152939
R21229 gnd.n4216 gnd.n4215 0.152939
R21230 gnd.n4215 gnd.n4214 0.152939
R21231 gnd.n4214 gnd.n2137 0.152939
R21232 gnd.n4210 gnd.n2137 0.152939
R21233 gnd.n4210 gnd.n4209 0.152939
R21234 gnd.n4209 gnd.n4208 0.152939
R21235 gnd.n4208 gnd.n2141 0.152939
R21236 gnd.n4204 gnd.n2141 0.152939
R21237 gnd.n4204 gnd.n870 0.152939
R21238 gnd.n5975 gnd.n870 0.152939
R21239 gnd.n5975 gnd.n5974 0.152939
R21240 gnd.n5962 gnd.n894 0.152939
R21241 gnd.n5962 gnd.n5961 0.152939
R21242 gnd.n5961 gnd.n5960 0.152939
R21243 gnd.n5960 gnd.n896 0.152939
R21244 gnd.n5956 gnd.n896 0.152939
R21245 gnd.n5956 gnd.n5955 0.152939
R21246 gnd.n4309 gnd.n4264 0.152939
R21247 gnd.n4309 gnd.n4308 0.152939
R21248 gnd.n4308 gnd.n4307 0.152939
R21249 gnd.n4307 gnd.n4265 0.152939
R21250 gnd.n4303 gnd.n4265 0.152939
R21251 gnd.n4303 gnd.n4302 0.152939
R21252 gnd.n4302 gnd.n4301 0.152939
R21253 gnd.n4301 gnd.n4269 0.152939
R21254 gnd.n4297 gnd.n4269 0.152939
R21255 gnd.n4297 gnd.n4296 0.152939
R21256 gnd.n4296 gnd.n4295 0.152939
R21257 gnd.n4295 gnd.n4273 0.152939
R21258 gnd.n4291 gnd.n4273 0.152939
R21259 gnd.n4291 gnd.n4290 0.152939
R21260 gnd.n4290 gnd.n4289 0.152939
R21261 gnd.n4289 gnd.n4277 0.152939
R21262 gnd.n4285 gnd.n4277 0.152939
R21263 gnd.n4285 gnd.n4284 0.152939
R21264 gnd.n4284 gnd.n4283 0.152939
R21265 gnd.n4283 gnd.n4281 0.152939
R21266 gnd.n4281 gnd.n2041 0.152939
R21267 gnd.n4419 gnd.n2041 0.152939
R21268 gnd.n4420 gnd.n4419 0.152939
R21269 gnd.n4421 gnd.n4420 0.152939
R21270 gnd.n4421 gnd.n2039 0.152939
R21271 gnd.n4525 gnd.n2039 0.152939
R21272 gnd.n4526 gnd.n4525 0.152939
R21273 gnd.n4554 gnd.n4526 0.152939
R21274 gnd.n4554 gnd.n4553 0.152939
R21275 gnd.n4553 gnd.n4552 0.152939
R21276 gnd.n4552 gnd.n4527 0.152939
R21277 gnd.n4548 gnd.n4527 0.152939
R21278 gnd.n4548 gnd.n4547 0.152939
R21279 gnd.n4547 gnd.n4546 0.152939
R21280 gnd.n4546 gnd.n4530 0.152939
R21281 gnd.n4542 gnd.n4530 0.152939
R21282 gnd.n4542 gnd.n4541 0.152939
R21283 gnd.n4541 gnd.n4540 0.152939
R21284 gnd.n4540 gnd.n4536 0.152939
R21285 gnd.n4536 gnd.n4535 0.152939
R21286 gnd.n4535 gnd.n1974 0.152939
R21287 gnd.n4662 gnd.n1974 0.152939
R21288 gnd.n4663 gnd.n4662 0.152939
R21289 gnd.n4690 gnd.n4663 0.152939
R21290 gnd.n4690 gnd.n4689 0.152939
R21291 gnd.n4689 gnd.n4688 0.152939
R21292 gnd.n4688 gnd.n4664 0.152939
R21293 gnd.n4684 gnd.n4664 0.152939
R21294 gnd.n4684 gnd.n4683 0.152939
R21295 gnd.n4683 gnd.n4682 0.152939
R21296 gnd.n4682 gnd.n4667 0.152939
R21297 gnd.n4678 gnd.n4667 0.152939
R21298 gnd.n4678 gnd.n4677 0.152939
R21299 gnd.n4677 gnd.n4676 0.152939
R21300 gnd.n4676 gnd.n4672 0.152939
R21301 gnd.n4672 gnd.n1881 0.152939
R21302 gnd.n4813 gnd.n1881 0.152939
R21303 gnd.n4814 gnd.n4813 0.152939
R21304 gnd.n4816 gnd.n4814 0.152939
R21305 gnd.n4816 gnd.n4815 0.152939
R21306 gnd.n4815 gnd.n1854 0.152939
R21307 gnd.n4862 gnd.n1854 0.152939
R21308 gnd.n4863 gnd.n4862 0.152939
R21309 gnd.n4880 gnd.n4863 0.152939
R21310 gnd.n4880 gnd.n4879 0.152939
R21311 gnd.n4879 gnd.n4878 0.152939
R21312 gnd.n4878 gnd.n4864 0.152939
R21313 gnd.n4874 gnd.n4864 0.152939
R21314 gnd.n4874 gnd.n4873 0.152939
R21315 gnd.n4873 gnd.n4872 0.152939
R21316 gnd.n4872 gnd.n4869 0.152939
R21317 gnd.n4869 gnd.n1802 0.152939
R21318 gnd.n4942 gnd.n1802 0.152939
R21319 gnd.n4943 gnd.n4942 0.152939
R21320 gnd.n4954 gnd.n4943 0.152939
R21321 gnd.n4954 gnd.n4953 0.152939
R21322 gnd.n4953 gnd.n4952 0.152939
R21323 gnd.n4952 gnd.n4944 0.152939
R21324 gnd.n4948 gnd.n4944 0.152939
R21325 gnd.n4948 gnd.n1724 0.152939
R21326 gnd.n5160 gnd.n1724 0.152939
R21327 gnd.n5161 gnd.n5160 0.152939
R21328 gnd.n5162 gnd.n5161 0.152939
R21329 gnd.n5162 gnd.n1712 0.152939
R21330 gnd.n5177 gnd.n1712 0.152939
R21331 gnd.n5178 gnd.n5177 0.152939
R21332 gnd.n5179 gnd.n5178 0.152939
R21333 gnd.n5179 gnd.n1700 0.152939
R21334 gnd.n5194 gnd.n1700 0.152939
R21335 gnd.n5195 gnd.n5194 0.152939
R21336 gnd.n5196 gnd.n5195 0.152939
R21337 gnd.n5196 gnd.n1687 0.152939
R21338 gnd.n5211 gnd.n1687 0.152939
R21339 gnd.n5212 gnd.n5211 0.152939
R21340 gnd.n5213 gnd.n5212 0.152939
R21341 gnd.n5213 gnd.n1676 0.152939
R21342 gnd.n5231 gnd.n1676 0.152939
R21343 gnd.n5232 gnd.n5231 0.152939
R21344 gnd.n5233 gnd.n5232 0.152939
R21345 gnd.n5233 gnd.n1318 0.152939
R21346 gnd.n5651 gnd.n1318 0.152939
R21347 gnd.n5650 gnd.n1319 0.152939
R21348 gnd.n5646 gnd.n1319 0.152939
R21349 gnd.n5646 gnd.n5645 0.152939
R21350 gnd.n5645 gnd.n5644 0.152939
R21351 gnd.n5644 gnd.n1323 0.152939
R21352 gnd.n5640 gnd.n1323 0.152939
R21353 gnd.n5304 gnd.n5266 0.152939
R21354 gnd.n5304 gnd.n5303 0.152939
R21355 gnd.n5303 gnd.n5302 0.152939
R21356 gnd.n5302 gnd.n5267 0.152939
R21357 gnd.n5298 gnd.n5267 0.152939
R21358 gnd.n5298 gnd.n5297 0.152939
R21359 gnd.n5297 gnd.n5296 0.152939
R21360 gnd.n5296 gnd.n5272 0.152939
R21361 gnd.n5292 gnd.n5272 0.152939
R21362 gnd.n5292 gnd.n1620 0.152939
R21363 gnd.n5353 gnd.n1620 0.152939
R21364 gnd.n5354 gnd.n5353 0.152939
R21365 gnd.n5355 gnd.n5354 0.152939
R21366 gnd.n5355 gnd.n1615 0.152939
R21367 gnd.n5368 gnd.n1615 0.152939
R21368 gnd.n5369 gnd.n5368 0.152939
R21369 gnd.n5374 gnd.n5369 0.152939
R21370 gnd.n5374 gnd.n5373 0.152939
R21371 gnd.n5373 gnd.n5372 0.152939
R21372 gnd.n5372 gnd.n67 0.152939
R21373 gnd.n7308 gnd.n7307 0.145814
R21374 gnd.n4131 gnd.n4130 0.145814
R21375 gnd.n4131 gnd.n2158 0.145814
R21376 gnd.n7308 gnd.n67 0.145814
R21377 gnd.n5955 gnd.n5954 0.128549
R21378 gnd.n5640 gnd.n5639 0.128549
R21379 gnd.n2520 gnd.n0 0.127478
R21380 gnd.n4164 gnd.n730 0.0919634
R21381 gnd.n5335 gnd.n83 0.0919634
R21382 gnd.n3100 gnd.n3099 0.0767195
R21383 gnd.n3099 gnd.n3098 0.0767195
R21384 gnd.n5954 gnd.n865 0.063
R21385 gnd.n5639 gnd.n1328 0.063
R21386 gnd.n184 gnd.n83 0.0614756
R21387 gnd.n6070 gnd.n730 0.0614756
R21388 gnd.n1496 gnd.n1328 0.0538288
R21389 gnd.n7244 gnd.n173 0.0538288
R21390 gnd.n4000 gnd.n2239 0.0538288
R21391 gnd.n5982 gnd.n865 0.0538288
R21392 gnd.n3666 gnd.n2282 0.0477147
R21393 gnd.n2863 gnd.n2751 0.0442063
R21394 gnd.n2864 gnd.n2863 0.0442063
R21395 gnd.n2865 gnd.n2864 0.0442063
R21396 gnd.n2865 gnd.n2740 0.0442063
R21397 gnd.n2879 gnd.n2740 0.0442063
R21398 gnd.n2880 gnd.n2879 0.0442063
R21399 gnd.n2881 gnd.n2880 0.0442063
R21400 gnd.n2881 gnd.n2727 0.0442063
R21401 gnd.n2925 gnd.n2727 0.0442063
R21402 gnd.n2926 gnd.n2925 0.0442063
R21403 gnd.n2928 gnd.n2661 0.0344674
R21404 gnd.n5461 gnd.n1496 0.0344674
R21405 gnd.n5461 gnd.n1498 0.0344674
R21406 gnd.n1522 gnd.n1498 0.0344674
R21407 gnd.n1523 gnd.n1522 0.0344674
R21408 gnd.n1524 gnd.n1523 0.0344674
R21409 gnd.n1525 gnd.n1524 0.0344674
R21410 gnd.n5279 gnd.n1525 0.0344674
R21411 gnd.n5279 gnd.n1543 0.0344674
R21412 gnd.n1544 gnd.n1543 0.0344674
R21413 gnd.n1545 gnd.n1544 0.0344674
R21414 gnd.n5285 gnd.n1545 0.0344674
R21415 gnd.n5285 gnd.n1563 0.0344674
R21416 gnd.n1564 gnd.n1563 0.0344674
R21417 gnd.n1565 gnd.n1564 0.0344674
R21418 gnd.n5362 gnd.n1565 0.0344674
R21419 gnd.n5362 gnd.n1580 0.0344674
R21420 gnd.n1581 gnd.n1580 0.0344674
R21421 gnd.n1582 gnd.n1581 0.0344674
R21422 gnd.n5382 gnd.n1582 0.0344674
R21423 gnd.n5383 gnd.n5382 0.0344674
R21424 gnd.n5383 gnd.n1607 0.0344674
R21425 gnd.n5392 gnd.n1607 0.0344674
R21426 gnd.n5392 gnd.n179 0.0344674
R21427 gnd.n6887 gnd.n179 0.0344674
R21428 gnd.n6888 gnd.n6887 0.0344674
R21429 gnd.n6888 gnd.n97 0.0344674
R21430 gnd.n98 gnd.n97 0.0344674
R21431 gnd.n99 gnd.n98 0.0344674
R21432 gnd.n7220 gnd.n99 0.0344674
R21433 gnd.n7220 gnd.n115 0.0344674
R21434 gnd.n116 gnd.n115 0.0344674
R21435 gnd.n117 gnd.n116 0.0344674
R21436 gnd.n7227 gnd.n117 0.0344674
R21437 gnd.n7227 gnd.n135 0.0344674
R21438 gnd.n136 gnd.n135 0.0344674
R21439 gnd.n137 gnd.n136 0.0344674
R21440 gnd.n7234 gnd.n137 0.0344674
R21441 gnd.n7234 gnd.n154 0.0344674
R21442 gnd.n155 gnd.n154 0.0344674
R21443 gnd.n156 gnd.n155 0.0344674
R21444 gnd.n172 gnd.n156 0.0344674
R21445 gnd.n7244 gnd.n172 0.0344674
R21446 gnd.n4001 gnd.n4000 0.0344674
R21447 gnd.n4001 gnd.n2235 0.0344674
R21448 gnd.n2236 gnd.n2235 0.0344674
R21449 gnd.n4007 gnd.n2236 0.0344674
R21450 gnd.n4008 gnd.n4007 0.0344674
R21451 gnd.n4008 gnd.n2213 0.0344674
R21452 gnd.n2213 gnd.n2210 0.0344674
R21453 gnd.n2211 gnd.n2210 0.0344674
R21454 gnd.n4042 gnd.n2211 0.0344674
R21455 gnd.n4043 gnd.n4042 0.0344674
R21456 gnd.n4043 gnd.n2188 0.0344674
R21457 gnd.n2188 gnd.n2184 0.0344674
R21458 gnd.n2185 gnd.n2184 0.0344674
R21459 gnd.n2186 gnd.n2185 0.0344674
R21460 gnd.n4081 gnd.n2186 0.0344674
R21461 gnd.n4082 gnd.n4081 0.0344674
R21462 gnd.n4082 gnd.n2165 0.0344674
R21463 gnd.n2165 gnd.n751 0.0344674
R21464 gnd.n752 gnd.n751 0.0344674
R21465 gnd.n753 gnd.n752 0.0344674
R21466 gnd.n2160 gnd.n753 0.0344674
R21467 gnd.n2160 gnd.n767 0.0344674
R21468 gnd.n768 gnd.n767 0.0344674
R21469 gnd.n769 gnd.n768 0.0344674
R21470 gnd.n4140 gnd.n769 0.0344674
R21471 gnd.n4140 gnd.n785 0.0344674
R21472 gnd.n786 gnd.n785 0.0344674
R21473 gnd.n787 gnd.n786 0.0344674
R21474 gnd.n2144 gnd.n787 0.0344674
R21475 gnd.n2144 gnd.n804 0.0344674
R21476 gnd.n805 gnd.n804 0.0344674
R21477 gnd.n806 gnd.n805 0.0344674
R21478 gnd.n4185 gnd.n806 0.0344674
R21479 gnd.n4185 gnd.n825 0.0344674
R21480 gnd.n826 gnd.n825 0.0344674
R21481 gnd.n827 gnd.n826 0.0344674
R21482 gnd.n4195 gnd.n827 0.0344674
R21483 gnd.n4195 gnd.n845 0.0344674
R21484 gnd.n846 gnd.n845 0.0344674
R21485 gnd.n847 gnd.n846 0.0344674
R21486 gnd.n864 gnd.n847 0.0344674
R21487 gnd.n5982 gnd.n864 0.0344674
R21488 gnd.n5953 gnd.n901 0.0343753
R21489 gnd.n5638 gnd.n5637 0.0343753
R21490 gnd.n5973 gnd.n5972 0.0296328
R21491 gnd.n5265 gnd.n5264 0.0296328
R21492 gnd.n2948 gnd.n2947 0.0269946
R21493 gnd.n2950 gnd.n2949 0.0269946
R21494 gnd.n2656 gnd.n2654 0.0269946
R21495 gnd.n2960 gnd.n2958 0.0269946
R21496 gnd.n2959 gnd.n2635 0.0269946
R21497 gnd.n2979 gnd.n2978 0.0269946
R21498 gnd.n2981 gnd.n2980 0.0269946
R21499 gnd.n2630 gnd.n2629 0.0269946
R21500 gnd.n2991 gnd.n2625 0.0269946
R21501 gnd.n2990 gnd.n2627 0.0269946
R21502 gnd.n2626 gnd.n2608 0.0269946
R21503 gnd.n3011 gnd.n2609 0.0269946
R21504 gnd.n3010 gnd.n2610 0.0269946
R21505 gnd.n3044 gnd.n2585 0.0269946
R21506 gnd.n3046 gnd.n3045 0.0269946
R21507 gnd.n3047 gnd.n2532 0.0269946
R21508 gnd.n2580 gnd.n2533 0.0269946
R21509 gnd.n2582 gnd.n2534 0.0269946
R21510 gnd.n3057 gnd.n3056 0.0269946
R21511 gnd.n3059 gnd.n3058 0.0269946
R21512 gnd.n3060 gnd.n2554 0.0269946
R21513 gnd.n3062 gnd.n2555 0.0269946
R21514 gnd.n3065 gnd.n2556 0.0269946
R21515 gnd.n3068 gnd.n3067 0.0269946
R21516 gnd.n3070 gnd.n3069 0.0269946
R21517 gnd.n3135 gnd.n2455 0.0269946
R21518 gnd.n3137 gnd.n3136 0.0269946
R21519 gnd.n3146 gnd.n2448 0.0269946
R21520 gnd.n3148 gnd.n3147 0.0269946
R21521 gnd.n3149 gnd.n2446 0.0269946
R21522 gnd.n3156 gnd.n3152 0.0269946
R21523 gnd.n3155 gnd.n3154 0.0269946
R21524 gnd.n3153 gnd.n2425 0.0269946
R21525 gnd.n3178 gnd.n2426 0.0269946
R21526 gnd.n3177 gnd.n2427 0.0269946
R21527 gnd.n3220 gnd.n2400 0.0269946
R21528 gnd.n3222 gnd.n3221 0.0269946
R21529 gnd.n3231 gnd.n2393 0.0269946
R21530 gnd.n3233 gnd.n3232 0.0269946
R21531 gnd.n3234 gnd.n2391 0.0269946
R21532 gnd.n3241 gnd.n3237 0.0269946
R21533 gnd.n3240 gnd.n3239 0.0269946
R21534 gnd.n3238 gnd.n2370 0.0269946
R21535 gnd.n3263 gnd.n2371 0.0269946
R21536 gnd.n3262 gnd.n2372 0.0269946
R21537 gnd.n3309 gnd.n2346 0.0269946
R21538 gnd.n3311 gnd.n3310 0.0269946
R21539 gnd.n3320 gnd.n2339 0.0269946
R21540 gnd.n3579 gnd.n2337 0.0269946
R21541 gnd.n3584 gnd.n3582 0.0269946
R21542 gnd.n3583 gnd.n2318 0.0269946
R21543 gnd.n3608 gnd.n3607 0.0269946
R21544 gnd.n5949 gnd.n907 0.022519
R21545 gnd.n5948 gnd.n908 0.022519
R21546 gnd.n5945 gnd.n5944 0.022519
R21547 gnd.n5941 gnd.n913 0.022519
R21548 gnd.n5940 gnd.n919 0.022519
R21549 gnd.n5937 gnd.n5936 0.022519
R21550 gnd.n5933 gnd.n923 0.022519
R21551 gnd.n5932 gnd.n927 0.022519
R21552 gnd.n5929 gnd.n5928 0.022519
R21553 gnd.n5925 gnd.n931 0.022519
R21554 gnd.n5924 gnd.n937 0.022519
R21555 gnd.n5921 gnd.n5920 0.022519
R21556 gnd.n5917 gnd.n941 0.022519
R21557 gnd.n5916 gnd.n945 0.022519
R21558 gnd.n5913 gnd.n5912 0.022519
R21559 gnd.n5909 gnd.n949 0.022519
R21560 gnd.n5908 gnd.n958 0.022519
R21561 gnd.n963 gnd.n962 0.022519
R21562 gnd.n5972 gnd.n872 0.022519
R21563 gnd.n5634 gnd.n1329 0.022519
R21564 gnd.n5633 gnd.n1333 0.022519
R21565 gnd.n5630 gnd.n5629 0.022519
R21566 gnd.n5626 gnd.n1338 0.022519
R21567 gnd.n5625 gnd.n1342 0.022519
R21568 gnd.n5622 gnd.n5621 0.022519
R21569 gnd.n5618 gnd.n1346 0.022519
R21570 gnd.n5617 gnd.n1350 0.022519
R21571 gnd.n5614 gnd.n5613 0.022519
R21572 gnd.n5610 gnd.n1354 0.022519
R21573 gnd.n5609 gnd.n1358 0.022519
R21574 gnd.n5606 gnd.n5605 0.022519
R21575 gnd.n5602 gnd.n1362 0.022519
R21576 gnd.n5601 gnd.n1366 0.022519
R21577 gnd.n5598 gnd.n5597 0.022519
R21578 gnd.n5594 gnd.n1370 0.022519
R21579 gnd.n5593 gnd.n1376 0.022519
R21580 gnd.n1641 gnd.n1379 0.022519
R21581 gnd.n5264 gnd.n1640 0.022519
R21582 gnd.n5265 gnd.n1639 0.0218415
R21583 gnd.n5973 gnd.n871 0.0218415
R21584 gnd.n2928 gnd.n2927 0.0202011
R21585 gnd.n2927 gnd.n2926 0.0148637
R21586 gnd.n3577 gnd.n3321 0.0144266
R21587 gnd.n3578 gnd.n3577 0.0130679
R21588 gnd.n907 gnd.n901 0.0123564
R21589 gnd.n5949 gnd.n5948 0.0123564
R21590 gnd.n5945 gnd.n908 0.0123564
R21591 gnd.n5944 gnd.n913 0.0123564
R21592 gnd.n5941 gnd.n5940 0.0123564
R21593 gnd.n5937 gnd.n919 0.0123564
R21594 gnd.n5936 gnd.n923 0.0123564
R21595 gnd.n5933 gnd.n5932 0.0123564
R21596 gnd.n5929 gnd.n927 0.0123564
R21597 gnd.n5928 gnd.n931 0.0123564
R21598 gnd.n5925 gnd.n5924 0.0123564
R21599 gnd.n5921 gnd.n937 0.0123564
R21600 gnd.n5920 gnd.n941 0.0123564
R21601 gnd.n5917 gnd.n5916 0.0123564
R21602 gnd.n5913 gnd.n945 0.0123564
R21603 gnd.n5912 gnd.n949 0.0123564
R21604 gnd.n5909 gnd.n5908 0.0123564
R21605 gnd.n963 gnd.n958 0.0123564
R21606 gnd.n962 gnd.n872 0.0123564
R21607 gnd.n5637 gnd.n1329 0.0123564
R21608 gnd.n5634 gnd.n5633 0.0123564
R21609 gnd.n5630 gnd.n1333 0.0123564
R21610 gnd.n5629 gnd.n1338 0.0123564
R21611 gnd.n5626 gnd.n5625 0.0123564
R21612 gnd.n5622 gnd.n1342 0.0123564
R21613 gnd.n5621 gnd.n1346 0.0123564
R21614 gnd.n5618 gnd.n5617 0.0123564
R21615 gnd.n5614 gnd.n1350 0.0123564
R21616 gnd.n5613 gnd.n1354 0.0123564
R21617 gnd.n5610 gnd.n5609 0.0123564
R21618 gnd.n5606 gnd.n1358 0.0123564
R21619 gnd.n5605 gnd.n1362 0.0123564
R21620 gnd.n5602 gnd.n5601 0.0123564
R21621 gnd.n5598 gnd.n1366 0.0123564
R21622 gnd.n5597 gnd.n1370 0.0123564
R21623 gnd.n5594 gnd.n5593 0.0123564
R21624 gnd.n1379 gnd.n1376 0.0123564
R21625 gnd.n1641 gnd.n1640 0.0123564
R21626 gnd.n2947 gnd.n2661 0.00797283
R21627 gnd.n2949 gnd.n2948 0.00797283
R21628 gnd.n2950 gnd.n2656 0.00797283
R21629 gnd.n2958 gnd.n2654 0.00797283
R21630 gnd.n2960 gnd.n2959 0.00797283
R21631 gnd.n2978 gnd.n2635 0.00797283
R21632 gnd.n2980 gnd.n2979 0.00797283
R21633 gnd.n2981 gnd.n2630 0.00797283
R21634 gnd.n2629 gnd.n2625 0.00797283
R21635 gnd.n2991 gnd.n2990 0.00797283
R21636 gnd.n2627 gnd.n2626 0.00797283
R21637 gnd.n2609 gnd.n2608 0.00797283
R21638 gnd.n3011 gnd.n3010 0.00797283
R21639 gnd.n2610 gnd.n2585 0.00797283
R21640 gnd.n3045 gnd.n3044 0.00797283
R21641 gnd.n3047 gnd.n3046 0.00797283
R21642 gnd.n2580 gnd.n2532 0.00797283
R21643 gnd.n2582 gnd.n2533 0.00797283
R21644 gnd.n3056 gnd.n2534 0.00797283
R21645 gnd.n3058 gnd.n3057 0.00797283
R21646 gnd.n3060 gnd.n3059 0.00797283
R21647 gnd.n3062 gnd.n2554 0.00797283
R21648 gnd.n3065 gnd.n2555 0.00797283
R21649 gnd.n3067 gnd.n2556 0.00797283
R21650 gnd.n3070 gnd.n3068 0.00797283
R21651 gnd.n3069 gnd.n2455 0.00797283
R21652 gnd.n3137 gnd.n3135 0.00797283
R21653 gnd.n3136 gnd.n2448 0.00797283
R21654 gnd.n3147 gnd.n3146 0.00797283
R21655 gnd.n3149 gnd.n3148 0.00797283
R21656 gnd.n3152 gnd.n2446 0.00797283
R21657 gnd.n3156 gnd.n3155 0.00797283
R21658 gnd.n3154 gnd.n3153 0.00797283
R21659 gnd.n2426 gnd.n2425 0.00797283
R21660 gnd.n3178 gnd.n3177 0.00797283
R21661 gnd.n2427 gnd.n2400 0.00797283
R21662 gnd.n3222 gnd.n3220 0.00797283
R21663 gnd.n3221 gnd.n2393 0.00797283
R21664 gnd.n3232 gnd.n3231 0.00797283
R21665 gnd.n3234 gnd.n3233 0.00797283
R21666 gnd.n3237 gnd.n2391 0.00797283
R21667 gnd.n3241 gnd.n3240 0.00797283
R21668 gnd.n3239 gnd.n3238 0.00797283
R21669 gnd.n2371 gnd.n2370 0.00797283
R21670 gnd.n3263 gnd.n3262 0.00797283
R21671 gnd.n2372 gnd.n2346 0.00797283
R21672 gnd.n3311 gnd.n3309 0.00797283
R21673 gnd.n3310 gnd.n2339 0.00797283
R21674 gnd.n3321 gnd.n3320 0.00797283
R21675 gnd.n3579 gnd.n3578 0.00797283
R21676 gnd.n3582 gnd.n2337 0.00797283
R21677 gnd.n3584 gnd.n3583 0.00797283
R21678 gnd.n3607 gnd.n2318 0.00797283
R21679 gnd.n3608 gnd.n2282 0.00797283
R21680 gnd.n5954 gnd.n5953 0.00592005
R21681 gnd.n5639 gnd.n5638 0.00592005
R21682 plus.n46 plus.t9 252.611
R21683 plus.n9 plus.t11 252.611
R21684 plus.n76 plus.t4 243.97
R21685 plus.n72 plus.t12 231.093
R21686 plus.n35 plus.t7 231.093
R21687 plus.n76 plus.n75 223.454
R21688 plus.n78 plus.n77 223.454
R21689 plus.n47 plus.t5 187.445
R21690 plus.n44 plus.t18 187.445
R21691 plus.n42 plus.t17 187.445
R21692 plus.n59 plus.t13 187.445
R21693 plus.n65 plus.t14 187.445
R21694 plus.n38 plus.t10 187.445
R21695 plus.n1 plus.t6 187.445
R21696 plus.n28 plus.t16 187.445
R21697 plus.n22 plus.t15 187.445
R21698 plus.n5 plus.t20 187.445
R21699 plus.n7 plus.t19 187.445
R21700 plus.n10 plus.t8 187.445
R21701 plus.n73 plus.n72 161.3
R21702 plus.n71 plus.n37 161.3
R21703 plus.n70 plus.n69 161.3
R21704 plus.n68 plus.n67 161.3
R21705 plus.n66 plus.n39 161.3
R21706 plus.n64 plus.n63 161.3
R21707 plus.n62 plus.n40 161.3
R21708 plus.n61 plus.n60 161.3
R21709 plus.n58 plus.n41 161.3
R21710 plus.n57 plus.n56 161.3
R21711 plus.n55 plus.n54 161.3
R21712 plus.n53 plus.n43 161.3
R21713 plus.n52 plus.n51 161.3
R21714 plus.n50 plus.n49 161.3
R21715 plus.n48 plus.n45 161.3
R21716 plus.n11 plus.n8 161.3
R21717 plus.n13 plus.n12 161.3
R21718 plus.n15 plus.n14 161.3
R21719 plus.n16 plus.n6 161.3
R21720 plus.n18 plus.n17 161.3
R21721 plus.n20 plus.n19 161.3
R21722 plus.n21 plus.n4 161.3
R21723 plus.n24 plus.n23 161.3
R21724 plus.n25 plus.n3 161.3
R21725 plus.n27 plus.n26 161.3
R21726 plus.n29 plus.n2 161.3
R21727 plus.n31 plus.n30 161.3
R21728 plus.n33 plus.n32 161.3
R21729 plus.n34 plus.n0 161.3
R21730 plus.n36 plus.n35 161.3
R21731 plus.n49 plus.n48 56.5617
R21732 plus.n58 plus.n57 56.5617
R21733 plus.n67 plus.n66 56.5617
R21734 plus.n30 plus.n29 56.5617
R21735 plus.n21 plus.n20 56.5617
R21736 plus.n12 plus.n11 56.5617
R21737 plus.n71 plus.n70 46.3896
R21738 plus.n34 plus.n33 46.3896
R21739 plus.n46 plus.n45 42.8164
R21740 plus.n9 plus.n8 42.8164
R21741 plus.n54 plus.n53 42.5146
R21742 plus.n60 plus.n40 42.5146
R21743 plus.n23 plus.n3 42.5146
R21744 plus.n17 plus.n16 42.5146
R21745 plus.n53 plus.n52 38.6395
R21746 plus.n64 plus.n40 38.6395
R21747 plus.n27 plus.n3 38.6395
R21748 plus.n16 plus.n15 38.6395
R21749 plus.n47 plus.n46 38.2514
R21750 plus.n10 plus.n9 38.2514
R21751 plus.n74 plus.n73 31.491
R21752 plus.n49 plus.n44 19.9199
R21753 plus.n66 plus.n65 19.9199
R21754 plus.n29 plus.n28 19.9199
R21755 plus.n12 plus.n7 19.9199
R21756 plus.n75 plus.t1 19.8005
R21757 plus.n75 plus.t2 19.8005
R21758 plus.n77 plus.t0 19.8005
R21759 plus.n77 plus.t3 19.8005
R21760 plus.n57 plus.n42 17.9525
R21761 plus.n59 plus.n58 17.9525
R21762 plus.n22 plus.n21 17.9525
R21763 plus.n20 plus.n5 17.9525
R21764 plus.n48 plus.n47 15.9852
R21765 plus.n67 plus.n38 15.9852
R21766 plus.n30 plus.n1 15.9852
R21767 plus.n11 plus.n10 15.9852
R21768 plus.n72 plus.n71 15.3369
R21769 plus.n35 plus.n34 15.3369
R21770 plus plus.n79 14.3853
R21771 plus.n74 plus.n36 11.9494
R21772 plus.n70 plus.n38 8.60764
R21773 plus.n33 plus.n1 8.60764
R21774 plus.n54 plus.n42 6.6403
R21775 plus.n60 plus.n59 6.6403
R21776 plus.n23 plus.n22 6.6403
R21777 plus.n17 plus.n5 6.6403
R21778 plus.n79 plus.n78 5.40567
R21779 plus.n52 plus.n44 4.67295
R21780 plus.n65 plus.n64 4.67295
R21781 plus.n28 plus.n27 4.67295
R21782 plus.n15 plus.n7 4.67295
R21783 plus.n79 plus.n74 1.188
R21784 plus.n78 plus.n76 0.716017
R21785 plus.n50 plus.n45 0.189894
R21786 plus.n51 plus.n50 0.189894
R21787 plus.n51 plus.n43 0.189894
R21788 plus.n55 plus.n43 0.189894
R21789 plus.n56 plus.n55 0.189894
R21790 plus.n56 plus.n41 0.189894
R21791 plus.n61 plus.n41 0.189894
R21792 plus.n62 plus.n61 0.189894
R21793 plus.n63 plus.n62 0.189894
R21794 plus.n63 plus.n39 0.189894
R21795 plus.n68 plus.n39 0.189894
R21796 plus.n69 plus.n68 0.189894
R21797 plus.n69 plus.n37 0.189894
R21798 plus.n73 plus.n37 0.189894
R21799 plus.n36 plus.n0 0.189894
R21800 plus.n32 plus.n0 0.189894
R21801 plus.n32 plus.n31 0.189894
R21802 plus.n31 plus.n2 0.189894
R21803 plus.n26 plus.n2 0.189894
R21804 plus.n26 plus.n25 0.189894
R21805 plus.n25 plus.n24 0.189894
R21806 plus.n24 plus.n4 0.189894
R21807 plus.n19 plus.n4 0.189894
R21808 plus.n19 plus.n18 0.189894
R21809 plus.n18 plus.n6 0.189894
R21810 plus.n14 plus.n6 0.189894
R21811 plus.n14 plus.n13 0.189894
R21812 plus.n13 plus.n8 0.189894
R21813 a_n3827_n3924.n2 a_n3827_n3924.t25 214.994
R21814 a_n3827_n3924.n12 a_n3827_n3924.t38 214.994
R21815 a_n3827_n3924.n2 a_n3827_n3924.t29 214.321
R21816 a_n3827_n3924.n13 a_n3827_n3924.t27 214.321
R21817 a_n3827_n3924.n14 a_n3827_n3924.t8 214.321
R21818 a_n3827_n3924.n15 a_n3827_n3924.t2 214.321
R21819 a_n3827_n3924.n16 a_n3827_n3924.t7 214.321
R21820 a_n3827_n3924.n17 a_n3827_n3924.t6 214.321
R21821 a_n3827_n3924.n0 a_n3827_n3924.t37 214.321
R21822 a_n3827_n3924.n12 a_n3827_n3924.t3 214.321
R21823 a_n3827_n3924.n1 a_n3827_n3924.t20 55.8337
R21824 a_n3827_n3924.n4 a_n3827_n3924.t41 55.8337
R21825 a_n3827_n3924.n11 a_n3827_n3924.t30 55.8337
R21826 a_n3827_n3924.n36 a_n3827_n3924.t17 55.8335
R21827 a_n3827_n3924.n34 a_n3827_n3924.t33 55.8335
R21828 a_n3827_n3924.n27 a_n3827_n3924.t4 55.8335
R21829 a_n3827_n3924.n26 a_n3827_n3924.t18 55.8335
R21830 a_n3827_n3924.n19 a_n3827_n3924.t22 55.8335
R21831 a_n3827_n3924.n38 a_n3827_n3924.n37 53.0052
R21832 a_n3827_n3924.n40 a_n3827_n3924.n39 53.0052
R21833 a_n3827_n3924.n6 a_n3827_n3924.n5 53.0052
R21834 a_n3827_n3924.n8 a_n3827_n3924.n7 53.0052
R21835 a_n3827_n3924.n10 a_n3827_n3924.n9 53.0052
R21836 a_n3827_n3924.n33 a_n3827_n3924.n32 53.0051
R21837 a_n3827_n3924.n31 a_n3827_n3924.n30 53.0051
R21838 a_n3827_n3924.n29 a_n3827_n3924.n28 53.0051
R21839 a_n3827_n3924.n25 a_n3827_n3924.n24 53.0051
R21840 a_n3827_n3924.n23 a_n3827_n3924.n22 53.0051
R21841 a_n3827_n3924.n21 a_n3827_n3924.n20 53.0051
R21842 a_n3827_n3924.n42 a_n3827_n3924.n41 53.0051
R21843 a_n3827_n3924.n18 a_n3827_n3924.n11 12.2417
R21844 a_n3827_n3924.n36 a_n3827_n3924.n35 12.2417
R21845 a_n3827_n3924.n19 a_n3827_n3924.n18 5.16214
R21846 a_n3827_n3924.n35 a_n3827_n3924.n34 5.16214
R21847 a_n3827_n3924.n37 a_n3827_n3924.t15 2.82907
R21848 a_n3827_n3924.n37 a_n3827_n3924.t19 2.82907
R21849 a_n3827_n3924.n39 a_n3827_n3924.t12 2.82907
R21850 a_n3827_n3924.n39 a_n3827_n3924.t16 2.82907
R21851 a_n3827_n3924.n5 a_n3827_n3924.t0 2.82907
R21852 a_n3827_n3924.n5 a_n3827_n3924.t32 2.82907
R21853 a_n3827_n3924.n7 a_n3827_n3924.t40 2.82907
R21854 a_n3827_n3924.n7 a_n3827_n3924.t31 2.82907
R21855 a_n3827_n3924.n9 a_n3827_n3924.t39 2.82907
R21856 a_n3827_n3924.n9 a_n3827_n3924.t1 2.82907
R21857 a_n3827_n3924.n32 a_n3827_n3924.t26 2.82907
R21858 a_n3827_n3924.n32 a_n3827_n3924.t28 2.82907
R21859 a_n3827_n3924.n30 a_n3827_n3924.t34 2.82907
R21860 a_n3827_n3924.n30 a_n3827_n3924.t35 2.82907
R21861 a_n3827_n3924.n28 a_n3827_n3924.t36 2.82907
R21862 a_n3827_n3924.n28 a_n3827_n3924.t5 2.82907
R21863 a_n3827_n3924.n24 a_n3827_n3924.t10 2.82907
R21864 a_n3827_n3924.n24 a_n3827_n3924.t21 2.82907
R21865 a_n3827_n3924.n22 a_n3827_n3924.t14 2.82907
R21866 a_n3827_n3924.n22 a_n3827_n3924.t9 2.82907
R21867 a_n3827_n3924.n20 a_n3827_n3924.t23 2.82907
R21868 a_n3827_n3924.n20 a_n3827_n3924.t13 2.82907
R21869 a_n3827_n3924.t24 a_n3827_n3924.n42 2.82907
R21870 a_n3827_n3924.n42 a_n3827_n3924.t11 2.82907
R21871 a_n3827_n3924.n35 a_n3827_n3924.n3 1.95694
R21872 a_n3827_n3924.n18 a_n3827_n3924.n0 1.95694
R21873 a_n3827_n3924.n0 a_n3827_n3924.n17 0.672012
R21874 a_n3827_n3924.n17 a_n3827_n3924.n16 0.672012
R21875 a_n3827_n3924.n16 a_n3827_n3924.n15 0.672012
R21876 a_n3827_n3924.n15 a_n3827_n3924.n14 0.672012
R21877 a_n3827_n3924.n14 a_n3827_n3924.n13 0.672012
R21878 a_n3827_n3924.n0 a_n3827_n3924.n12 0.672012
R21879 a_n3827_n3924.n13 a_n3827_n3924.n3 0.541924
R21880 a_n3827_n3924.n21 a_n3827_n3924.n19 0.530672
R21881 a_n3827_n3924.n23 a_n3827_n3924.n21 0.530672
R21882 a_n3827_n3924.n25 a_n3827_n3924.n23 0.530672
R21883 a_n3827_n3924.n26 a_n3827_n3924.n25 0.530672
R21884 a_n3827_n3924.n29 a_n3827_n3924.n27 0.530672
R21885 a_n3827_n3924.n31 a_n3827_n3924.n29 0.530672
R21886 a_n3827_n3924.n33 a_n3827_n3924.n31 0.530672
R21887 a_n3827_n3924.n34 a_n3827_n3924.n33 0.530672
R21888 a_n3827_n3924.n11 a_n3827_n3924.n10 0.530672
R21889 a_n3827_n3924.n10 a_n3827_n3924.n8 0.530672
R21890 a_n3827_n3924.n8 a_n3827_n3924.n6 0.530672
R21891 a_n3827_n3924.n6 a_n3827_n3924.n4 0.530672
R21892 a_n3827_n3924.n41 a_n3827_n3924.n1 0.530672
R21893 a_n3827_n3924.n41 a_n3827_n3924.n40 0.530672
R21894 a_n3827_n3924.n40 a_n3827_n3924.n38 0.530672
R21895 a_n3827_n3924.n38 a_n3827_n3924.n36 0.530672
R21896 a_n3827_n3924.n27 a_n3827_n3924.n26 0.235414
R21897 a_n3827_n3924.n4 a_n3827_n3924.n1 0.235414
R21898 a_n3827_n3924.n3 a_n3827_n3924.n2 0.130587
R21899 diffpairibias.n0 diffpairibias.t27 436.822
R21900 diffpairibias.n27 diffpairibias.t24 435.479
R21901 diffpairibias.n26 diffpairibias.t21 435.479
R21902 diffpairibias.n25 diffpairibias.t22 435.479
R21903 diffpairibias.n24 diffpairibias.t26 435.479
R21904 diffpairibias.n23 diffpairibias.t20 435.479
R21905 diffpairibias.n0 diffpairibias.t23 435.479
R21906 diffpairibias.n1 diffpairibias.t28 435.479
R21907 diffpairibias.n2 diffpairibias.t25 435.479
R21908 diffpairibias.n3 diffpairibias.t29 435.479
R21909 diffpairibias.n13 diffpairibias.t14 377.536
R21910 diffpairibias.n13 diffpairibias.t0 376.193
R21911 diffpairibias.n14 diffpairibias.t10 376.193
R21912 diffpairibias.n15 diffpairibias.t12 376.193
R21913 diffpairibias.n16 diffpairibias.t6 376.193
R21914 diffpairibias.n17 diffpairibias.t2 376.193
R21915 diffpairibias.n18 diffpairibias.t16 376.193
R21916 diffpairibias.n19 diffpairibias.t4 376.193
R21917 diffpairibias.n20 diffpairibias.t18 376.193
R21918 diffpairibias.n21 diffpairibias.t8 376.193
R21919 diffpairibias.n4 diffpairibias.t15 113.368
R21920 diffpairibias.n4 diffpairibias.t1 112.698
R21921 diffpairibias.n5 diffpairibias.t11 112.698
R21922 diffpairibias.n6 diffpairibias.t13 112.698
R21923 diffpairibias.n7 diffpairibias.t7 112.698
R21924 diffpairibias.n8 diffpairibias.t3 112.698
R21925 diffpairibias.n9 diffpairibias.t17 112.698
R21926 diffpairibias.n10 diffpairibias.t5 112.698
R21927 diffpairibias.n11 diffpairibias.t19 112.698
R21928 diffpairibias.n12 diffpairibias.t9 112.698
R21929 diffpairibias.n22 diffpairibias.n21 4.77242
R21930 diffpairibias.n22 diffpairibias.n12 4.30807
R21931 diffpairibias.n23 diffpairibias.n22 4.13945
R21932 diffpairibias.n21 diffpairibias.n20 1.34352
R21933 diffpairibias.n20 diffpairibias.n19 1.34352
R21934 diffpairibias.n19 diffpairibias.n18 1.34352
R21935 diffpairibias.n18 diffpairibias.n17 1.34352
R21936 diffpairibias.n17 diffpairibias.n16 1.34352
R21937 diffpairibias.n16 diffpairibias.n15 1.34352
R21938 diffpairibias.n15 diffpairibias.n14 1.34352
R21939 diffpairibias.n14 diffpairibias.n13 1.34352
R21940 diffpairibias.n3 diffpairibias.n2 1.34352
R21941 diffpairibias.n2 diffpairibias.n1 1.34352
R21942 diffpairibias.n1 diffpairibias.n0 1.34352
R21943 diffpairibias.n24 diffpairibias.n23 1.34352
R21944 diffpairibias.n25 diffpairibias.n24 1.34352
R21945 diffpairibias.n26 diffpairibias.n25 1.34352
R21946 diffpairibias.n27 diffpairibias.n26 1.34352
R21947 diffpairibias.n28 diffpairibias.n27 0.862419
R21948 diffpairibias diffpairibias.n28 0.684875
R21949 diffpairibias.n12 diffpairibias.n11 0.672012
R21950 diffpairibias.n11 diffpairibias.n10 0.672012
R21951 diffpairibias.n10 diffpairibias.n9 0.672012
R21952 diffpairibias.n9 diffpairibias.n8 0.672012
R21953 diffpairibias.n8 diffpairibias.n7 0.672012
R21954 diffpairibias.n7 diffpairibias.n6 0.672012
R21955 diffpairibias.n6 diffpairibias.n5 0.672012
R21956 diffpairibias.n5 diffpairibias.n4 0.672012
R21957 diffpairibias.n28 diffpairibias.n3 0.190907
R21958 minus.n46 minus.t20 252.611
R21959 minus.n9 minus.t13 252.611
R21960 minus.n78 minus.t3 243.255
R21961 minus.n72 minus.t15 231.093
R21962 minus.n35 minus.t17 231.093
R21963 minus.n77 minus.n75 224.169
R21964 minus.n77 minus.n76 223.454
R21965 minus.n38 minus.t12 187.445
R21966 minus.n65 minus.t7 187.445
R21967 minus.n59 minus.t6 187.445
R21968 minus.n42 minus.t11 187.445
R21969 minus.n44 minus.t10 187.445
R21970 minus.n47 minus.t16 187.445
R21971 minus.n10 minus.t9 187.445
R21972 minus.n7 minus.t8 187.445
R21973 minus.n5 minus.t5 187.445
R21974 minus.n22 minus.t18 187.445
R21975 minus.n28 minus.t19 187.445
R21976 minus.n1 minus.t14 187.445
R21977 minus.n48 minus.n45 161.3
R21978 minus.n50 minus.n49 161.3
R21979 minus.n52 minus.n51 161.3
R21980 minus.n53 minus.n43 161.3
R21981 minus.n55 minus.n54 161.3
R21982 minus.n57 minus.n56 161.3
R21983 minus.n58 minus.n41 161.3
R21984 minus.n61 minus.n60 161.3
R21985 minus.n62 minus.n40 161.3
R21986 minus.n64 minus.n63 161.3
R21987 minus.n66 minus.n39 161.3
R21988 minus.n68 minus.n67 161.3
R21989 minus.n70 minus.n69 161.3
R21990 minus.n71 minus.n37 161.3
R21991 minus.n73 minus.n72 161.3
R21992 minus.n36 minus.n35 161.3
R21993 minus.n34 minus.n0 161.3
R21994 minus.n33 minus.n32 161.3
R21995 minus.n31 minus.n30 161.3
R21996 minus.n29 minus.n2 161.3
R21997 minus.n27 minus.n26 161.3
R21998 minus.n25 minus.n3 161.3
R21999 minus.n24 minus.n23 161.3
R22000 minus.n21 minus.n4 161.3
R22001 minus.n20 minus.n19 161.3
R22002 minus.n18 minus.n17 161.3
R22003 minus.n16 minus.n6 161.3
R22004 minus.n15 minus.n14 161.3
R22005 minus.n13 minus.n12 161.3
R22006 minus.n11 minus.n8 161.3
R22007 minus.n67 minus.n66 56.5617
R22008 minus.n58 minus.n57 56.5617
R22009 minus.n49 minus.n48 56.5617
R22010 minus.n12 minus.n11 56.5617
R22011 minus.n21 minus.n20 56.5617
R22012 minus.n30 minus.n29 56.5617
R22013 minus.n71 minus.n70 46.3896
R22014 minus.n34 minus.n33 46.3896
R22015 minus.n46 minus.n45 42.8164
R22016 minus.n9 minus.n8 42.8164
R22017 minus.n60 minus.n40 42.5146
R22018 minus.n54 minus.n53 42.5146
R22019 minus.n17 minus.n16 42.5146
R22020 minus.n23 minus.n3 42.5146
R22021 minus.n64 minus.n40 38.6395
R22022 minus.n53 minus.n52 38.6395
R22023 minus.n16 minus.n15 38.6395
R22024 minus.n27 minus.n3 38.6395
R22025 minus.n47 minus.n46 38.2514
R22026 minus.n10 minus.n9 38.2514
R22027 minus.n74 minus.n73 31.7069
R22028 minus.n66 minus.n65 19.9199
R22029 minus.n49 minus.n44 19.9199
R22030 minus.n12 minus.n7 19.9199
R22031 minus.n29 minus.n28 19.9199
R22032 minus.n76 minus.t2 19.8005
R22033 minus.n76 minus.t0 19.8005
R22034 minus.n75 minus.t1 19.8005
R22035 minus.n75 minus.t4 19.8005
R22036 minus.n59 minus.n58 17.9525
R22037 minus.n57 minus.n42 17.9525
R22038 minus.n20 minus.n5 17.9525
R22039 minus.n22 minus.n21 17.9525
R22040 minus.n67 minus.n38 15.9852
R22041 minus.n48 minus.n47 15.9852
R22042 minus.n11 minus.n10 15.9852
R22043 minus.n30 minus.n1 15.9852
R22044 minus.n72 minus.n71 15.3369
R22045 minus.n35 minus.n34 15.3369
R22046 minus.n74 minus.n36 12.1653
R22047 minus minus.n79 11.5131
R22048 minus.n70 minus.n38 8.60764
R22049 minus.n33 minus.n1 8.60764
R22050 minus.n60 minus.n59 6.6403
R22051 minus.n54 minus.n42 6.6403
R22052 minus.n17 minus.n5 6.6403
R22053 minus.n23 minus.n22 6.6403
R22054 minus.n79 minus.n78 4.80222
R22055 minus.n65 minus.n64 4.67295
R22056 minus.n52 minus.n44 4.67295
R22057 minus.n15 minus.n7 4.67295
R22058 minus.n28 minus.n27 4.67295
R22059 minus.n79 minus.n74 0.972091
R22060 minus.n78 minus.n77 0.716017
R22061 minus.n73 minus.n37 0.189894
R22062 minus.n69 minus.n37 0.189894
R22063 minus.n69 minus.n68 0.189894
R22064 minus.n68 minus.n39 0.189894
R22065 minus.n63 minus.n39 0.189894
R22066 minus.n63 minus.n62 0.189894
R22067 minus.n62 minus.n61 0.189894
R22068 minus.n61 minus.n41 0.189894
R22069 minus.n56 minus.n41 0.189894
R22070 minus.n56 minus.n55 0.189894
R22071 minus.n55 minus.n43 0.189894
R22072 minus.n51 minus.n43 0.189894
R22073 minus.n51 minus.n50 0.189894
R22074 minus.n50 minus.n45 0.189894
R22075 minus.n13 minus.n8 0.189894
R22076 minus.n14 minus.n13 0.189894
R22077 minus.n14 minus.n6 0.189894
R22078 minus.n18 minus.n6 0.189894
R22079 minus.n19 minus.n18 0.189894
R22080 minus.n19 minus.n4 0.189894
R22081 minus.n24 minus.n4 0.189894
R22082 minus.n25 minus.n24 0.189894
R22083 minus.n26 minus.n25 0.189894
R22084 minus.n26 minus.n2 0.189894
R22085 minus.n31 minus.n2 0.189894
R22086 minus.n32 minus.n31 0.189894
R22087 minus.n32 minus.n0 0.189894
R22088 minus.n36 minus.n0 0.189894
R22089 a_n2650_8322.n10 a_n2650_8322.t29 74.6477
R22090 a_n2650_8322.n1 a_n2650_8322.t21 74.6477
R22091 a_n2650_8322.n24 a_n2650_8322.t23 74.6474
R22092 a_n2650_8322.n18 a_n2650_8322.t20 74.2899
R22093 a_n2650_8322.n11 a_n2650_8322.t27 74.2899
R22094 a_n2650_8322.n12 a_n2650_8322.t30 74.2899
R22095 a_n2650_8322.n15 a_n2650_8322.t31 74.2899
R22096 a_n2650_8322.n8 a_n2650_8322.t6 74.2899
R22097 a_n2650_8322.n24 a_n2650_8322.n23 70.6783
R22098 a_n2650_8322.n22 a_n2650_8322.n21 70.6783
R22099 a_n2650_8322.n20 a_n2650_8322.n19 70.6783
R22100 a_n2650_8322.n10 a_n2650_8322.n9 70.6783
R22101 a_n2650_8322.n14 a_n2650_8322.n13 70.6783
R22102 a_n2650_8322.n1 a_n2650_8322.n0 70.6783
R22103 a_n2650_8322.n3 a_n2650_8322.n2 70.6783
R22104 a_n2650_8322.n5 a_n2650_8322.n4 70.6783
R22105 a_n2650_8322.n7 a_n2650_8322.n6 70.6783
R22106 a_n2650_8322.n26 a_n2650_8322.n25 70.6782
R22107 a_n2650_8322.n16 a_n2650_8322.n8 24.1867
R22108 a_n2650_8322.n17 a_n2650_8322.t0 9.73422
R22109 a_n2650_8322.n16 a_n2650_8322.n15 7.67184
R22110 a_n2650_8322.n18 a_n2650_8322.n17 6.55222
R22111 a_n2650_8322.n17 a_n2650_8322.n16 5.3452
R22112 a_n2650_8322.n23 a_n2650_8322.t18 3.61217
R22113 a_n2650_8322.n23 a_n2650_8322.t14 3.61217
R22114 a_n2650_8322.n21 a_n2650_8322.t22 3.61217
R22115 a_n2650_8322.n21 a_n2650_8322.t11 3.61217
R22116 a_n2650_8322.n19 a_n2650_8322.t9 3.61217
R22117 a_n2650_8322.n19 a_n2650_8322.t10 3.61217
R22118 a_n2650_8322.n9 a_n2650_8322.t32 3.61217
R22119 a_n2650_8322.n9 a_n2650_8322.t33 3.61217
R22120 a_n2650_8322.n13 a_n2650_8322.t28 3.61217
R22121 a_n2650_8322.n13 a_n2650_8322.t26 3.61217
R22122 a_n2650_8322.n0 a_n2650_8322.t24 3.61217
R22123 a_n2650_8322.n0 a_n2650_8322.t16 3.61217
R22124 a_n2650_8322.n2 a_n2650_8322.t8 3.61217
R22125 a_n2650_8322.n2 a_n2650_8322.t7 3.61217
R22126 a_n2650_8322.n4 a_n2650_8322.t19 3.61217
R22127 a_n2650_8322.n4 a_n2650_8322.t13 3.61217
R22128 a_n2650_8322.n6 a_n2650_8322.t17 3.61217
R22129 a_n2650_8322.n6 a_n2650_8322.t15 3.61217
R22130 a_n2650_8322.n26 a_n2650_8322.t12 3.61217
R22131 a_n2650_8322.t25 a_n2650_8322.n26 3.61217
R22132 a_n2650_8322.n15 a_n2650_8322.n14 0.358259
R22133 a_n2650_8322.n14 a_n2650_8322.n12 0.358259
R22134 a_n2650_8322.n11 a_n2650_8322.n10 0.358259
R22135 a_n2650_8322.n8 a_n2650_8322.n7 0.358259
R22136 a_n2650_8322.n7 a_n2650_8322.n5 0.358259
R22137 a_n2650_8322.n5 a_n2650_8322.n3 0.358259
R22138 a_n2650_8322.n3 a_n2650_8322.n1 0.358259
R22139 a_n2650_8322.n20 a_n2650_8322.n18 0.358259
R22140 a_n2650_8322.n22 a_n2650_8322.n20 0.358259
R22141 a_n2650_8322.n25 a_n2650_8322.n22 0.358259
R22142 a_n2650_8322.n25 a_n2650_8322.n24 0.358259
R22143 a_n2650_8322.n12 a_n2650_8322.n11 0.101793
R22144 a_n2650_8322.t5 a_n2650_8322.t3 0.0788333
R22145 a_n2650_8322.t1 a_n2650_8322.t2 0.0788333
R22146 a_n2650_8322.t0 a_n2650_8322.t4 0.0788333
R22147 a_n2650_8322.t1 a_n2650_8322.t5 0.0318333
R22148 a_n2650_8322.t0 a_n2650_8322.t2 0.0318333
R22149 a_n2650_8322.t3 a_n2650_8322.t2 0.0318333
R22150 a_n2650_8322.t4 a_n2650_8322.t1 0.0318333
R22151 outputibias.n27 outputibias.n1 289.615
R22152 outputibias.n58 outputibias.n32 289.615
R22153 outputibias.n90 outputibias.n64 289.615
R22154 outputibias.n122 outputibias.n96 289.615
R22155 outputibias.n28 outputibias.n27 185
R22156 outputibias.n26 outputibias.n25 185
R22157 outputibias.n5 outputibias.n4 185
R22158 outputibias.n20 outputibias.n19 185
R22159 outputibias.n18 outputibias.n17 185
R22160 outputibias.n9 outputibias.n8 185
R22161 outputibias.n12 outputibias.n11 185
R22162 outputibias.n59 outputibias.n58 185
R22163 outputibias.n57 outputibias.n56 185
R22164 outputibias.n36 outputibias.n35 185
R22165 outputibias.n51 outputibias.n50 185
R22166 outputibias.n49 outputibias.n48 185
R22167 outputibias.n40 outputibias.n39 185
R22168 outputibias.n43 outputibias.n42 185
R22169 outputibias.n91 outputibias.n90 185
R22170 outputibias.n89 outputibias.n88 185
R22171 outputibias.n68 outputibias.n67 185
R22172 outputibias.n83 outputibias.n82 185
R22173 outputibias.n81 outputibias.n80 185
R22174 outputibias.n72 outputibias.n71 185
R22175 outputibias.n75 outputibias.n74 185
R22176 outputibias.n123 outputibias.n122 185
R22177 outputibias.n121 outputibias.n120 185
R22178 outputibias.n100 outputibias.n99 185
R22179 outputibias.n115 outputibias.n114 185
R22180 outputibias.n113 outputibias.n112 185
R22181 outputibias.n104 outputibias.n103 185
R22182 outputibias.n107 outputibias.n106 185
R22183 outputibias.n0 outputibias.t10 178.945
R22184 outputibias.n133 outputibias.t8 177.018
R22185 outputibias.n132 outputibias.t11 177.018
R22186 outputibias.n0 outputibias.t9 177.018
R22187 outputibias.t7 outputibias.n10 147.661
R22188 outputibias.t1 outputibias.n41 147.661
R22189 outputibias.t3 outputibias.n73 147.661
R22190 outputibias.t5 outputibias.n105 147.661
R22191 outputibias.n128 outputibias.t6 132.363
R22192 outputibias.n128 outputibias.t0 130.436
R22193 outputibias.n129 outputibias.t2 130.436
R22194 outputibias.n130 outputibias.t4 130.436
R22195 outputibias.n27 outputibias.n26 104.615
R22196 outputibias.n26 outputibias.n4 104.615
R22197 outputibias.n19 outputibias.n4 104.615
R22198 outputibias.n19 outputibias.n18 104.615
R22199 outputibias.n18 outputibias.n8 104.615
R22200 outputibias.n11 outputibias.n8 104.615
R22201 outputibias.n58 outputibias.n57 104.615
R22202 outputibias.n57 outputibias.n35 104.615
R22203 outputibias.n50 outputibias.n35 104.615
R22204 outputibias.n50 outputibias.n49 104.615
R22205 outputibias.n49 outputibias.n39 104.615
R22206 outputibias.n42 outputibias.n39 104.615
R22207 outputibias.n90 outputibias.n89 104.615
R22208 outputibias.n89 outputibias.n67 104.615
R22209 outputibias.n82 outputibias.n67 104.615
R22210 outputibias.n82 outputibias.n81 104.615
R22211 outputibias.n81 outputibias.n71 104.615
R22212 outputibias.n74 outputibias.n71 104.615
R22213 outputibias.n122 outputibias.n121 104.615
R22214 outputibias.n121 outputibias.n99 104.615
R22215 outputibias.n114 outputibias.n99 104.615
R22216 outputibias.n114 outputibias.n113 104.615
R22217 outputibias.n113 outputibias.n103 104.615
R22218 outputibias.n106 outputibias.n103 104.615
R22219 outputibias.n63 outputibias.n31 95.6354
R22220 outputibias.n63 outputibias.n62 94.6732
R22221 outputibias.n95 outputibias.n94 94.6732
R22222 outputibias.n127 outputibias.n126 94.6732
R22223 outputibias.n11 outputibias.t7 52.3082
R22224 outputibias.n42 outputibias.t1 52.3082
R22225 outputibias.n74 outputibias.t3 52.3082
R22226 outputibias.n106 outputibias.t5 52.3082
R22227 outputibias.n12 outputibias.n10 15.6674
R22228 outputibias.n43 outputibias.n41 15.6674
R22229 outputibias.n75 outputibias.n73 15.6674
R22230 outputibias.n107 outputibias.n105 15.6674
R22231 outputibias.n13 outputibias.n9 12.8005
R22232 outputibias.n44 outputibias.n40 12.8005
R22233 outputibias.n76 outputibias.n72 12.8005
R22234 outputibias.n108 outputibias.n104 12.8005
R22235 outputibias.n17 outputibias.n16 12.0247
R22236 outputibias.n48 outputibias.n47 12.0247
R22237 outputibias.n80 outputibias.n79 12.0247
R22238 outputibias.n112 outputibias.n111 12.0247
R22239 outputibias.n20 outputibias.n7 11.249
R22240 outputibias.n51 outputibias.n38 11.249
R22241 outputibias.n83 outputibias.n70 11.249
R22242 outputibias.n115 outputibias.n102 11.249
R22243 outputibias.n21 outputibias.n5 10.4732
R22244 outputibias.n52 outputibias.n36 10.4732
R22245 outputibias.n84 outputibias.n68 10.4732
R22246 outputibias.n116 outputibias.n100 10.4732
R22247 outputibias.n25 outputibias.n24 9.69747
R22248 outputibias.n56 outputibias.n55 9.69747
R22249 outputibias.n88 outputibias.n87 9.69747
R22250 outputibias.n120 outputibias.n119 9.69747
R22251 outputibias.n31 outputibias.n30 9.45567
R22252 outputibias.n62 outputibias.n61 9.45567
R22253 outputibias.n94 outputibias.n93 9.45567
R22254 outputibias.n126 outputibias.n125 9.45567
R22255 outputibias.n30 outputibias.n29 9.3005
R22256 outputibias.n3 outputibias.n2 9.3005
R22257 outputibias.n24 outputibias.n23 9.3005
R22258 outputibias.n22 outputibias.n21 9.3005
R22259 outputibias.n7 outputibias.n6 9.3005
R22260 outputibias.n16 outputibias.n15 9.3005
R22261 outputibias.n14 outputibias.n13 9.3005
R22262 outputibias.n61 outputibias.n60 9.3005
R22263 outputibias.n34 outputibias.n33 9.3005
R22264 outputibias.n55 outputibias.n54 9.3005
R22265 outputibias.n53 outputibias.n52 9.3005
R22266 outputibias.n38 outputibias.n37 9.3005
R22267 outputibias.n47 outputibias.n46 9.3005
R22268 outputibias.n45 outputibias.n44 9.3005
R22269 outputibias.n93 outputibias.n92 9.3005
R22270 outputibias.n66 outputibias.n65 9.3005
R22271 outputibias.n87 outputibias.n86 9.3005
R22272 outputibias.n85 outputibias.n84 9.3005
R22273 outputibias.n70 outputibias.n69 9.3005
R22274 outputibias.n79 outputibias.n78 9.3005
R22275 outputibias.n77 outputibias.n76 9.3005
R22276 outputibias.n125 outputibias.n124 9.3005
R22277 outputibias.n98 outputibias.n97 9.3005
R22278 outputibias.n119 outputibias.n118 9.3005
R22279 outputibias.n117 outputibias.n116 9.3005
R22280 outputibias.n102 outputibias.n101 9.3005
R22281 outputibias.n111 outputibias.n110 9.3005
R22282 outputibias.n109 outputibias.n108 9.3005
R22283 outputibias.n28 outputibias.n3 8.92171
R22284 outputibias.n59 outputibias.n34 8.92171
R22285 outputibias.n91 outputibias.n66 8.92171
R22286 outputibias.n123 outputibias.n98 8.92171
R22287 outputibias.n29 outputibias.n1 8.14595
R22288 outputibias.n60 outputibias.n32 8.14595
R22289 outputibias.n92 outputibias.n64 8.14595
R22290 outputibias.n124 outputibias.n96 8.14595
R22291 outputibias.n31 outputibias.n1 5.81868
R22292 outputibias.n62 outputibias.n32 5.81868
R22293 outputibias.n94 outputibias.n64 5.81868
R22294 outputibias.n126 outputibias.n96 5.81868
R22295 outputibias.n131 outputibias.n130 5.20947
R22296 outputibias.n29 outputibias.n28 5.04292
R22297 outputibias.n60 outputibias.n59 5.04292
R22298 outputibias.n92 outputibias.n91 5.04292
R22299 outputibias.n124 outputibias.n123 5.04292
R22300 outputibias.n131 outputibias.n127 4.42209
R22301 outputibias.n14 outputibias.n10 4.38594
R22302 outputibias.n45 outputibias.n41 4.38594
R22303 outputibias.n77 outputibias.n73 4.38594
R22304 outputibias.n109 outputibias.n105 4.38594
R22305 outputibias.n132 outputibias.n131 4.28454
R22306 outputibias.n25 outputibias.n3 4.26717
R22307 outputibias.n56 outputibias.n34 4.26717
R22308 outputibias.n88 outputibias.n66 4.26717
R22309 outputibias.n120 outputibias.n98 4.26717
R22310 outputibias.n24 outputibias.n5 3.49141
R22311 outputibias.n55 outputibias.n36 3.49141
R22312 outputibias.n87 outputibias.n68 3.49141
R22313 outputibias.n119 outputibias.n100 3.49141
R22314 outputibias.n21 outputibias.n20 2.71565
R22315 outputibias.n52 outputibias.n51 2.71565
R22316 outputibias.n84 outputibias.n83 2.71565
R22317 outputibias.n116 outputibias.n115 2.71565
R22318 outputibias.n17 outputibias.n7 1.93989
R22319 outputibias.n48 outputibias.n38 1.93989
R22320 outputibias.n80 outputibias.n70 1.93989
R22321 outputibias.n112 outputibias.n102 1.93989
R22322 outputibias.n130 outputibias.n129 1.9266
R22323 outputibias.n129 outputibias.n128 1.9266
R22324 outputibias.n133 outputibias.n132 1.92658
R22325 outputibias.n134 outputibias.n133 1.29913
R22326 outputibias.n16 outputibias.n9 1.16414
R22327 outputibias.n47 outputibias.n40 1.16414
R22328 outputibias.n79 outputibias.n72 1.16414
R22329 outputibias.n111 outputibias.n104 1.16414
R22330 outputibias.n127 outputibias.n95 0.962709
R22331 outputibias.n95 outputibias.n63 0.962709
R22332 outputibias.n13 outputibias.n12 0.388379
R22333 outputibias.n44 outputibias.n43 0.388379
R22334 outputibias.n76 outputibias.n75 0.388379
R22335 outputibias.n108 outputibias.n107 0.388379
R22336 outputibias.n134 outputibias.n0 0.337251
R22337 outputibias outputibias.n134 0.302375
R22338 outputibias.n30 outputibias.n2 0.155672
R22339 outputibias.n23 outputibias.n2 0.155672
R22340 outputibias.n23 outputibias.n22 0.155672
R22341 outputibias.n22 outputibias.n6 0.155672
R22342 outputibias.n15 outputibias.n6 0.155672
R22343 outputibias.n15 outputibias.n14 0.155672
R22344 outputibias.n61 outputibias.n33 0.155672
R22345 outputibias.n54 outputibias.n33 0.155672
R22346 outputibias.n54 outputibias.n53 0.155672
R22347 outputibias.n53 outputibias.n37 0.155672
R22348 outputibias.n46 outputibias.n37 0.155672
R22349 outputibias.n46 outputibias.n45 0.155672
R22350 outputibias.n93 outputibias.n65 0.155672
R22351 outputibias.n86 outputibias.n65 0.155672
R22352 outputibias.n86 outputibias.n85 0.155672
R22353 outputibias.n85 outputibias.n69 0.155672
R22354 outputibias.n78 outputibias.n69 0.155672
R22355 outputibias.n78 outputibias.n77 0.155672
R22356 outputibias.n125 outputibias.n97 0.155672
R22357 outputibias.n118 outputibias.n97 0.155672
R22358 outputibias.n118 outputibias.n117 0.155672
R22359 outputibias.n117 outputibias.n101 0.155672
R22360 outputibias.n110 outputibias.n101 0.155672
R22361 outputibias.n110 outputibias.n109 0.155672
R22362 output.n41 output.n15 289.615
R22363 output.n72 output.n46 289.615
R22364 output.n104 output.n78 289.615
R22365 output.n136 output.n110 289.615
R22366 output.n77 output.n45 197.26
R22367 output.n77 output.n76 196.298
R22368 output.n109 output.n108 196.298
R22369 output.n141 output.n140 196.298
R22370 output.n42 output.n41 185
R22371 output.n40 output.n39 185
R22372 output.n19 output.n18 185
R22373 output.n34 output.n33 185
R22374 output.n32 output.n31 185
R22375 output.n23 output.n22 185
R22376 output.n26 output.n25 185
R22377 output.n73 output.n72 185
R22378 output.n71 output.n70 185
R22379 output.n50 output.n49 185
R22380 output.n65 output.n64 185
R22381 output.n63 output.n62 185
R22382 output.n54 output.n53 185
R22383 output.n57 output.n56 185
R22384 output.n105 output.n104 185
R22385 output.n103 output.n102 185
R22386 output.n82 output.n81 185
R22387 output.n97 output.n96 185
R22388 output.n95 output.n94 185
R22389 output.n86 output.n85 185
R22390 output.n89 output.n88 185
R22391 output.n137 output.n136 185
R22392 output.n135 output.n134 185
R22393 output.n114 output.n113 185
R22394 output.n129 output.n128 185
R22395 output.n127 output.n126 185
R22396 output.n118 output.n117 185
R22397 output.n121 output.n120 185
R22398 output.t17 output.n24 147.661
R22399 output.t18 output.n55 147.661
R22400 output.t19 output.n87 147.661
R22401 output.t16 output.n119 147.661
R22402 output.n41 output.n40 104.615
R22403 output.n40 output.n18 104.615
R22404 output.n33 output.n18 104.615
R22405 output.n33 output.n32 104.615
R22406 output.n32 output.n22 104.615
R22407 output.n25 output.n22 104.615
R22408 output.n72 output.n71 104.615
R22409 output.n71 output.n49 104.615
R22410 output.n64 output.n49 104.615
R22411 output.n64 output.n63 104.615
R22412 output.n63 output.n53 104.615
R22413 output.n56 output.n53 104.615
R22414 output.n104 output.n103 104.615
R22415 output.n103 output.n81 104.615
R22416 output.n96 output.n81 104.615
R22417 output.n96 output.n95 104.615
R22418 output.n95 output.n85 104.615
R22419 output.n88 output.n85 104.615
R22420 output.n136 output.n135 104.615
R22421 output.n135 output.n113 104.615
R22422 output.n128 output.n113 104.615
R22423 output.n128 output.n127 104.615
R22424 output.n127 output.n117 104.615
R22425 output.n120 output.n117 104.615
R22426 output.n1 output.t1 77.056
R22427 output.n14 output.t2 76.6694
R22428 output.n1 output.n0 72.7095
R22429 output.n3 output.n2 72.7095
R22430 output.n5 output.n4 72.7095
R22431 output.n7 output.n6 72.7095
R22432 output.n9 output.n8 72.7095
R22433 output.n11 output.n10 72.7095
R22434 output.n13 output.n12 72.7095
R22435 output.n25 output.t17 52.3082
R22436 output.n56 output.t18 52.3082
R22437 output.n88 output.t19 52.3082
R22438 output.n120 output.t16 52.3082
R22439 output.n26 output.n24 15.6674
R22440 output.n57 output.n55 15.6674
R22441 output.n89 output.n87 15.6674
R22442 output.n121 output.n119 15.6674
R22443 output.n27 output.n23 12.8005
R22444 output.n58 output.n54 12.8005
R22445 output.n90 output.n86 12.8005
R22446 output.n122 output.n118 12.8005
R22447 output.n31 output.n30 12.0247
R22448 output.n62 output.n61 12.0247
R22449 output.n94 output.n93 12.0247
R22450 output.n126 output.n125 12.0247
R22451 output.n34 output.n21 11.249
R22452 output.n65 output.n52 11.249
R22453 output.n97 output.n84 11.249
R22454 output.n129 output.n116 11.249
R22455 output.n35 output.n19 10.4732
R22456 output.n66 output.n50 10.4732
R22457 output.n98 output.n82 10.4732
R22458 output.n130 output.n114 10.4732
R22459 output.n39 output.n38 9.69747
R22460 output.n70 output.n69 9.69747
R22461 output.n102 output.n101 9.69747
R22462 output.n134 output.n133 9.69747
R22463 output.n45 output.n44 9.45567
R22464 output.n76 output.n75 9.45567
R22465 output.n108 output.n107 9.45567
R22466 output.n140 output.n139 9.45567
R22467 output.n44 output.n43 9.3005
R22468 output.n17 output.n16 9.3005
R22469 output.n38 output.n37 9.3005
R22470 output.n36 output.n35 9.3005
R22471 output.n21 output.n20 9.3005
R22472 output.n30 output.n29 9.3005
R22473 output.n28 output.n27 9.3005
R22474 output.n75 output.n74 9.3005
R22475 output.n48 output.n47 9.3005
R22476 output.n69 output.n68 9.3005
R22477 output.n67 output.n66 9.3005
R22478 output.n52 output.n51 9.3005
R22479 output.n61 output.n60 9.3005
R22480 output.n59 output.n58 9.3005
R22481 output.n107 output.n106 9.3005
R22482 output.n80 output.n79 9.3005
R22483 output.n101 output.n100 9.3005
R22484 output.n99 output.n98 9.3005
R22485 output.n84 output.n83 9.3005
R22486 output.n93 output.n92 9.3005
R22487 output.n91 output.n90 9.3005
R22488 output.n139 output.n138 9.3005
R22489 output.n112 output.n111 9.3005
R22490 output.n133 output.n132 9.3005
R22491 output.n131 output.n130 9.3005
R22492 output.n116 output.n115 9.3005
R22493 output.n125 output.n124 9.3005
R22494 output.n123 output.n122 9.3005
R22495 output.n42 output.n17 8.92171
R22496 output.n73 output.n48 8.92171
R22497 output.n105 output.n80 8.92171
R22498 output.n137 output.n112 8.92171
R22499 output output.n141 8.15037
R22500 output.n43 output.n15 8.14595
R22501 output.n74 output.n46 8.14595
R22502 output.n106 output.n78 8.14595
R22503 output.n138 output.n110 8.14595
R22504 output.n45 output.n15 5.81868
R22505 output.n76 output.n46 5.81868
R22506 output.n108 output.n78 5.81868
R22507 output.n140 output.n110 5.81868
R22508 output.n43 output.n42 5.04292
R22509 output.n74 output.n73 5.04292
R22510 output.n106 output.n105 5.04292
R22511 output.n138 output.n137 5.04292
R22512 output.n28 output.n24 4.38594
R22513 output.n59 output.n55 4.38594
R22514 output.n91 output.n87 4.38594
R22515 output.n123 output.n119 4.38594
R22516 output.n39 output.n17 4.26717
R22517 output.n70 output.n48 4.26717
R22518 output.n102 output.n80 4.26717
R22519 output.n134 output.n112 4.26717
R22520 output.n0 output.t13 3.9605
R22521 output.n0 output.t15 3.9605
R22522 output.n2 output.t5 3.9605
R22523 output.n2 output.t4 3.9605
R22524 output.n4 output.t10 3.9605
R22525 output.n4 output.t14 3.9605
R22526 output.n6 output.t3 3.9605
R22527 output.n6 output.t6 3.9605
R22528 output.n8 output.t7 3.9605
R22529 output.n8 output.t12 3.9605
R22530 output.n10 output.t0 3.9605
R22531 output.n10 output.t8 3.9605
R22532 output.n12 output.t11 3.9605
R22533 output.n12 output.t9 3.9605
R22534 output.n38 output.n19 3.49141
R22535 output.n69 output.n50 3.49141
R22536 output.n101 output.n82 3.49141
R22537 output.n133 output.n114 3.49141
R22538 output.n35 output.n34 2.71565
R22539 output.n66 output.n65 2.71565
R22540 output.n98 output.n97 2.71565
R22541 output.n130 output.n129 2.71565
R22542 output.n31 output.n21 1.93989
R22543 output.n62 output.n52 1.93989
R22544 output.n94 output.n84 1.93989
R22545 output.n126 output.n116 1.93989
R22546 output.n30 output.n23 1.16414
R22547 output.n61 output.n54 1.16414
R22548 output.n93 output.n86 1.16414
R22549 output.n125 output.n118 1.16414
R22550 output.n141 output.n109 0.962709
R22551 output.n109 output.n77 0.962709
R22552 output.n27 output.n26 0.388379
R22553 output.n58 output.n57 0.388379
R22554 output.n90 output.n89 0.388379
R22555 output.n122 output.n121 0.388379
R22556 output.n14 output.n13 0.387128
R22557 output.n13 output.n11 0.387128
R22558 output.n11 output.n9 0.387128
R22559 output.n9 output.n7 0.387128
R22560 output.n7 output.n5 0.387128
R22561 output.n5 output.n3 0.387128
R22562 output.n3 output.n1 0.387128
R22563 output.n44 output.n16 0.155672
R22564 output.n37 output.n16 0.155672
R22565 output.n37 output.n36 0.155672
R22566 output.n36 output.n20 0.155672
R22567 output.n29 output.n20 0.155672
R22568 output.n29 output.n28 0.155672
R22569 output.n75 output.n47 0.155672
R22570 output.n68 output.n47 0.155672
R22571 output.n68 output.n67 0.155672
R22572 output.n67 output.n51 0.155672
R22573 output.n60 output.n51 0.155672
R22574 output.n60 output.n59 0.155672
R22575 output.n107 output.n79 0.155672
R22576 output.n100 output.n79 0.155672
R22577 output.n100 output.n99 0.155672
R22578 output.n99 output.n83 0.155672
R22579 output.n92 output.n83 0.155672
R22580 output.n92 output.n91 0.155672
R22581 output.n139 output.n111 0.155672
R22582 output.n132 output.n111 0.155672
R22583 output.n132 output.n131 0.155672
R22584 output.n131 output.n115 0.155672
R22585 output.n124 output.n115 0.155672
R22586 output.n124 output.n123 0.155672
R22587 output output.n14 0.126227
C0 output outputibias 2.34152f
C1 vdd output 7.23429f
C2 CSoutput output 6.13881f
C3 CSoutput outputibias 0.032386f
C4 vdd CSoutput 92.5996f
C5 commonsourceibias output 0.006808f
C6 minus diffpairibias 3.46e-19
C7 CSoutput minus 2.73976f
C8 vdd plus 0.081257f
C9 plus diffpairibias 2.47e-19
C10 commonsourceibias outputibias 0.003832f
C11 vdd commonsourceibias 0.004218f
C12 CSoutput plus 0.854329f
C13 commonsourceibias diffpairibias 0.064336f
C14 CSoutput commonsourceibias 42.3358f
C15 minus plus 9.12235f
C16 minus commonsourceibias 0.331977f
C17 plus commonsourceibias 0.277692f
C18 diffpairibias gnd 60.00273f
C19 outputibias gnd 32.465668f
C20 output gnd 15.47879f
C21 commonsourceibias gnd 0.145029p
C22 plus gnd 32.580948f
C23 minus gnd 26.80269f
C24 CSoutput gnd 0.107678p
C25 vdd gnd 0.445486p
C26 output.t1 gnd 0.464308f
C27 output.t13 gnd 0.044422f
C28 output.t15 gnd 0.044422f
C29 output.n0 gnd 0.364624f
C30 output.n1 gnd 0.614102f
C31 output.t5 gnd 0.044422f
C32 output.t4 gnd 0.044422f
C33 output.n2 gnd 0.364624f
C34 output.n3 gnd 0.350265f
C35 output.t10 gnd 0.044422f
C36 output.t14 gnd 0.044422f
C37 output.n4 gnd 0.364624f
C38 output.n5 gnd 0.350265f
C39 output.t3 gnd 0.044422f
C40 output.t6 gnd 0.044422f
C41 output.n6 gnd 0.364624f
C42 output.n7 gnd 0.350265f
C43 output.t7 gnd 0.044422f
C44 output.t12 gnd 0.044422f
C45 output.n8 gnd 0.364624f
C46 output.n9 gnd 0.350265f
C47 output.t0 gnd 0.044422f
C48 output.t8 gnd 0.044422f
C49 output.n10 gnd 0.364624f
C50 output.n11 gnd 0.350265f
C51 output.t11 gnd 0.044422f
C52 output.t9 gnd 0.044422f
C53 output.n12 gnd 0.364624f
C54 output.n13 gnd 0.350265f
C55 output.t2 gnd 0.462979f
C56 output.n14 gnd 0.28994f
C57 output.n15 gnd 0.015803f
C58 output.n16 gnd 0.011243f
C59 output.n17 gnd 0.006041f
C60 output.n18 gnd 0.01428f
C61 output.n19 gnd 0.006397f
C62 output.n20 gnd 0.011243f
C63 output.n21 gnd 0.006041f
C64 output.n22 gnd 0.01428f
C65 output.n23 gnd 0.006397f
C66 output.n24 gnd 0.048111f
C67 output.t17 gnd 0.023274f
C68 output.n25 gnd 0.01071f
C69 output.n26 gnd 0.008435f
C70 output.n27 gnd 0.006041f
C71 output.n28 gnd 0.267512f
C72 output.n29 gnd 0.011243f
C73 output.n30 gnd 0.006041f
C74 output.n31 gnd 0.006397f
C75 output.n32 gnd 0.01428f
C76 output.n33 gnd 0.01428f
C77 output.n34 gnd 0.006397f
C78 output.n35 gnd 0.006041f
C79 output.n36 gnd 0.011243f
C80 output.n37 gnd 0.011243f
C81 output.n38 gnd 0.006041f
C82 output.n39 gnd 0.006397f
C83 output.n40 gnd 0.01428f
C84 output.n41 gnd 0.030913f
C85 output.n42 gnd 0.006397f
C86 output.n43 gnd 0.006041f
C87 output.n44 gnd 0.025987f
C88 output.n45 gnd 0.097665f
C89 output.n46 gnd 0.015803f
C90 output.n47 gnd 0.011243f
C91 output.n48 gnd 0.006041f
C92 output.n49 gnd 0.01428f
C93 output.n50 gnd 0.006397f
C94 output.n51 gnd 0.011243f
C95 output.n52 gnd 0.006041f
C96 output.n53 gnd 0.01428f
C97 output.n54 gnd 0.006397f
C98 output.n55 gnd 0.048111f
C99 output.t18 gnd 0.023274f
C100 output.n56 gnd 0.01071f
C101 output.n57 gnd 0.008435f
C102 output.n58 gnd 0.006041f
C103 output.n59 gnd 0.267512f
C104 output.n60 gnd 0.011243f
C105 output.n61 gnd 0.006041f
C106 output.n62 gnd 0.006397f
C107 output.n63 gnd 0.01428f
C108 output.n64 gnd 0.01428f
C109 output.n65 gnd 0.006397f
C110 output.n66 gnd 0.006041f
C111 output.n67 gnd 0.011243f
C112 output.n68 gnd 0.011243f
C113 output.n69 gnd 0.006041f
C114 output.n70 gnd 0.006397f
C115 output.n71 gnd 0.01428f
C116 output.n72 gnd 0.030913f
C117 output.n73 gnd 0.006397f
C118 output.n74 gnd 0.006041f
C119 output.n75 gnd 0.025987f
C120 output.n76 gnd 0.09306f
C121 output.n77 gnd 1.65264f
C122 output.n78 gnd 0.015803f
C123 output.n79 gnd 0.011243f
C124 output.n80 gnd 0.006041f
C125 output.n81 gnd 0.01428f
C126 output.n82 gnd 0.006397f
C127 output.n83 gnd 0.011243f
C128 output.n84 gnd 0.006041f
C129 output.n85 gnd 0.01428f
C130 output.n86 gnd 0.006397f
C131 output.n87 gnd 0.048111f
C132 output.t19 gnd 0.023274f
C133 output.n88 gnd 0.01071f
C134 output.n89 gnd 0.008435f
C135 output.n90 gnd 0.006041f
C136 output.n91 gnd 0.267512f
C137 output.n92 gnd 0.011243f
C138 output.n93 gnd 0.006041f
C139 output.n94 gnd 0.006397f
C140 output.n95 gnd 0.01428f
C141 output.n96 gnd 0.01428f
C142 output.n97 gnd 0.006397f
C143 output.n98 gnd 0.006041f
C144 output.n99 gnd 0.011243f
C145 output.n100 gnd 0.011243f
C146 output.n101 gnd 0.006041f
C147 output.n102 gnd 0.006397f
C148 output.n103 gnd 0.01428f
C149 output.n104 gnd 0.030913f
C150 output.n105 gnd 0.006397f
C151 output.n106 gnd 0.006041f
C152 output.n107 gnd 0.025987f
C153 output.n108 gnd 0.09306f
C154 output.n109 gnd 0.713089f
C155 output.n110 gnd 0.015803f
C156 output.n111 gnd 0.011243f
C157 output.n112 gnd 0.006041f
C158 output.n113 gnd 0.01428f
C159 output.n114 gnd 0.006397f
C160 output.n115 gnd 0.011243f
C161 output.n116 gnd 0.006041f
C162 output.n117 gnd 0.01428f
C163 output.n118 gnd 0.006397f
C164 output.n119 gnd 0.048111f
C165 output.t16 gnd 0.023274f
C166 output.n120 gnd 0.01071f
C167 output.n121 gnd 0.008435f
C168 output.n122 gnd 0.006041f
C169 output.n123 gnd 0.267512f
C170 output.n124 gnd 0.011243f
C171 output.n125 gnd 0.006041f
C172 output.n126 gnd 0.006397f
C173 output.n127 gnd 0.01428f
C174 output.n128 gnd 0.01428f
C175 output.n129 gnd 0.006397f
C176 output.n130 gnd 0.006041f
C177 output.n131 gnd 0.011243f
C178 output.n132 gnd 0.011243f
C179 output.n133 gnd 0.006041f
C180 output.n134 gnd 0.006397f
C181 output.n135 gnd 0.01428f
C182 output.n136 gnd 0.030913f
C183 output.n137 gnd 0.006397f
C184 output.n138 gnd 0.006041f
C185 output.n139 gnd 0.025987f
C186 output.n140 gnd 0.09306f
C187 output.n141 gnd 1.67353f
C188 outputibias.t9 gnd 0.11477f
C189 outputibias.t10 gnd 0.115567f
C190 outputibias.n0 gnd 0.130108f
C191 outputibias.n1 gnd 0.001372f
C192 outputibias.n2 gnd 9.76e-19
C193 outputibias.n3 gnd 5.24e-19
C194 outputibias.n4 gnd 0.001239f
C195 outputibias.n5 gnd 5.55e-19
C196 outputibias.n6 gnd 9.76e-19
C197 outputibias.n7 gnd 5.24e-19
C198 outputibias.n8 gnd 0.001239f
C199 outputibias.n9 gnd 5.55e-19
C200 outputibias.n10 gnd 0.004176f
C201 outputibias.t7 gnd 0.00202f
C202 outputibias.n11 gnd 9.3e-19
C203 outputibias.n12 gnd 7.32e-19
C204 outputibias.n13 gnd 5.24e-19
C205 outputibias.n14 gnd 0.02322f
C206 outputibias.n15 gnd 9.76e-19
C207 outputibias.n16 gnd 5.24e-19
C208 outputibias.n17 gnd 5.55e-19
C209 outputibias.n18 gnd 0.001239f
C210 outputibias.n19 gnd 0.001239f
C211 outputibias.n20 gnd 5.55e-19
C212 outputibias.n21 gnd 5.24e-19
C213 outputibias.n22 gnd 9.76e-19
C214 outputibias.n23 gnd 9.76e-19
C215 outputibias.n24 gnd 5.24e-19
C216 outputibias.n25 gnd 5.55e-19
C217 outputibias.n26 gnd 0.001239f
C218 outputibias.n27 gnd 0.002683f
C219 outputibias.n28 gnd 5.55e-19
C220 outputibias.n29 gnd 5.24e-19
C221 outputibias.n30 gnd 0.002256f
C222 outputibias.n31 gnd 0.005781f
C223 outputibias.n32 gnd 0.001372f
C224 outputibias.n33 gnd 9.76e-19
C225 outputibias.n34 gnd 5.24e-19
C226 outputibias.n35 gnd 0.001239f
C227 outputibias.n36 gnd 5.55e-19
C228 outputibias.n37 gnd 9.76e-19
C229 outputibias.n38 gnd 5.24e-19
C230 outputibias.n39 gnd 0.001239f
C231 outputibias.n40 gnd 5.55e-19
C232 outputibias.n41 gnd 0.004176f
C233 outputibias.t1 gnd 0.00202f
C234 outputibias.n42 gnd 9.3e-19
C235 outputibias.n43 gnd 7.32e-19
C236 outputibias.n44 gnd 5.24e-19
C237 outputibias.n45 gnd 0.02322f
C238 outputibias.n46 gnd 9.76e-19
C239 outputibias.n47 gnd 5.24e-19
C240 outputibias.n48 gnd 5.55e-19
C241 outputibias.n49 gnd 0.001239f
C242 outputibias.n50 gnd 0.001239f
C243 outputibias.n51 gnd 5.55e-19
C244 outputibias.n52 gnd 5.24e-19
C245 outputibias.n53 gnd 9.76e-19
C246 outputibias.n54 gnd 9.76e-19
C247 outputibias.n55 gnd 5.24e-19
C248 outputibias.n56 gnd 5.55e-19
C249 outputibias.n57 gnd 0.001239f
C250 outputibias.n58 gnd 0.002683f
C251 outputibias.n59 gnd 5.55e-19
C252 outputibias.n60 gnd 5.24e-19
C253 outputibias.n61 gnd 0.002256f
C254 outputibias.n62 gnd 0.005197f
C255 outputibias.n63 gnd 0.121892f
C256 outputibias.n64 gnd 0.001372f
C257 outputibias.n65 gnd 9.76e-19
C258 outputibias.n66 gnd 5.24e-19
C259 outputibias.n67 gnd 0.001239f
C260 outputibias.n68 gnd 5.55e-19
C261 outputibias.n69 gnd 9.76e-19
C262 outputibias.n70 gnd 5.24e-19
C263 outputibias.n71 gnd 0.001239f
C264 outputibias.n72 gnd 5.55e-19
C265 outputibias.n73 gnd 0.004176f
C266 outputibias.t3 gnd 0.00202f
C267 outputibias.n74 gnd 9.3e-19
C268 outputibias.n75 gnd 7.32e-19
C269 outputibias.n76 gnd 5.24e-19
C270 outputibias.n77 gnd 0.02322f
C271 outputibias.n78 gnd 9.76e-19
C272 outputibias.n79 gnd 5.24e-19
C273 outputibias.n80 gnd 5.55e-19
C274 outputibias.n81 gnd 0.001239f
C275 outputibias.n82 gnd 0.001239f
C276 outputibias.n83 gnd 5.55e-19
C277 outputibias.n84 gnd 5.24e-19
C278 outputibias.n85 gnd 9.76e-19
C279 outputibias.n86 gnd 9.76e-19
C280 outputibias.n87 gnd 5.24e-19
C281 outputibias.n88 gnd 5.55e-19
C282 outputibias.n89 gnd 0.001239f
C283 outputibias.n90 gnd 0.002683f
C284 outputibias.n91 gnd 5.55e-19
C285 outputibias.n92 gnd 5.24e-19
C286 outputibias.n93 gnd 0.002256f
C287 outputibias.n94 gnd 0.005197f
C288 outputibias.n95 gnd 0.064513f
C289 outputibias.n96 gnd 0.001372f
C290 outputibias.n97 gnd 9.76e-19
C291 outputibias.n98 gnd 5.24e-19
C292 outputibias.n99 gnd 0.001239f
C293 outputibias.n100 gnd 5.55e-19
C294 outputibias.n101 gnd 9.76e-19
C295 outputibias.n102 gnd 5.24e-19
C296 outputibias.n103 gnd 0.001239f
C297 outputibias.n104 gnd 5.55e-19
C298 outputibias.n105 gnd 0.004176f
C299 outputibias.t5 gnd 0.00202f
C300 outputibias.n106 gnd 9.3e-19
C301 outputibias.n107 gnd 7.32e-19
C302 outputibias.n108 gnd 5.24e-19
C303 outputibias.n109 gnd 0.02322f
C304 outputibias.n110 gnd 9.76e-19
C305 outputibias.n111 gnd 5.24e-19
C306 outputibias.n112 gnd 5.55e-19
C307 outputibias.n113 gnd 0.001239f
C308 outputibias.n114 gnd 0.001239f
C309 outputibias.n115 gnd 5.55e-19
C310 outputibias.n116 gnd 5.24e-19
C311 outputibias.n117 gnd 9.76e-19
C312 outputibias.n118 gnd 9.76e-19
C313 outputibias.n119 gnd 5.24e-19
C314 outputibias.n120 gnd 5.55e-19
C315 outputibias.n121 gnd 0.001239f
C316 outputibias.n122 gnd 0.002683f
C317 outputibias.n123 gnd 5.55e-19
C318 outputibias.n124 gnd 5.24e-19
C319 outputibias.n125 gnd 0.002256f
C320 outputibias.n126 gnd 0.005197f
C321 outputibias.n127 gnd 0.084814f
C322 outputibias.t4 gnd 0.108319f
C323 outputibias.t2 gnd 0.108319f
C324 outputibias.t0 gnd 0.108319f
C325 outputibias.t6 gnd 0.109238f
C326 outputibias.n128 gnd 0.134674f
C327 outputibias.n129 gnd 0.07244f
C328 outputibias.n130 gnd 0.079818f
C329 outputibias.n131 gnd 0.164901f
C330 outputibias.t11 gnd 0.11477f
C331 outputibias.n132 gnd 0.067481f
C332 outputibias.t8 gnd 0.11477f
C333 outputibias.n133 gnd 0.065115f
C334 outputibias.n134 gnd 0.029159f
C335 a_n2650_8322.t12 gnd 0.098025f
C336 a_n2650_8322.t2 gnd 20.3361f
C337 a_n2650_8322.t3 gnd 20.193499f
C338 a_n2650_8322.t5 gnd 20.193499f
C339 a_n2650_8322.t1 gnd 20.3361f
C340 a_n2650_8322.t4 gnd 20.193499f
C341 a_n2650_8322.t0 gnd 28.546698f
C342 a_n2650_8322.t21 gnd 0.917854f
C343 a_n2650_8322.t24 gnd 0.098025f
C344 a_n2650_8322.t16 gnd 0.098025f
C345 a_n2650_8322.n0 gnd 0.690486f
C346 a_n2650_8322.n1 gnd 0.771516f
C347 a_n2650_8322.t8 gnd 0.098025f
C348 a_n2650_8322.t7 gnd 0.098025f
C349 a_n2650_8322.n2 gnd 0.690486f
C350 a_n2650_8322.n3 gnd 0.391998f
C351 a_n2650_8322.t19 gnd 0.098025f
C352 a_n2650_8322.t13 gnd 0.098025f
C353 a_n2650_8322.n4 gnd 0.690486f
C354 a_n2650_8322.n5 gnd 0.391998f
C355 a_n2650_8322.t17 gnd 0.098025f
C356 a_n2650_8322.t15 gnd 0.098025f
C357 a_n2650_8322.n6 gnd 0.690486f
C358 a_n2650_8322.n7 gnd 0.391998f
C359 a_n2650_8322.t6 gnd 0.916026f
C360 a_n2650_8322.n8 gnd 1.7094f
C361 a_n2650_8322.t29 gnd 0.917854f
C362 a_n2650_8322.t32 gnd 0.098025f
C363 a_n2650_8322.t33 gnd 0.098025f
C364 a_n2650_8322.n9 gnd 0.690486f
C365 a_n2650_8322.n10 gnd 0.771516f
C366 a_n2650_8322.t27 gnd 0.916026f
C367 a_n2650_8322.n11 gnd 0.388238f
C368 a_n2650_8322.t30 gnd 0.916026f
C369 a_n2650_8322.n12 gnd 0.388238f
C370 a_n2650_8322.t28 gnd 0.098025f
C371 a_n2650_8322.t26 gnd 0.098025f
C372 a_n2650_8322.n13 gnd 0.690486f
C373 a_n2650_8322.n14 gnd 0.391998f
C374 a_n2650_8322.t31 gnd 0.916026f
C375 a_n2650_8322.n15 gnd 1.27375f
C376 a_n2650_8322.n16 gnd 2.08118f
C377 a_n2650_8322.n17 gnd 3.30568f
C378 a_n2650_8322.t20 gnd 0.916026f
C379 a_n2650_8322.n18 gnd 0.996372f
C380 a_n2650_8322.t9 gnd 0.098025f
C381 a_n2650_8322.t10 gnd 0.098025f
C382 a_n2650_8322.n19 gnd 0.690486f
C383 a_n2650_8322.n20 gnd 0.391998f
C384 a_n2650_8322.t22 gnd 0.098025f
C385 a_n2650_8322.t11 gnd 0.098025f
C386 a_n2650_8322.n21 gnd 0.690486f
C387 a_n2650_8322.n22 gnd 0.391998f
C388 a_n2650_8322.t23 gnd 0.917851f
C389 a_n2650_8322.t18 gnd 0.098025f
C390 a_n2650_8322.t14 gnd 0.098025f
C391 a_n2650_8322.n23 gnd 0.690486f
C392 a_n2650_8322.n24 gnd 0.771518f
C393 a_n2650_8322.n25 gnd 0.391996f
C394 a_n2650_8322.n26 gnd 0.690488f
C395 a_n2650_8322.t25 gnd 0.098025f
C396 minus.n0 gnd 0.030008f
C397 minus.t14 gnd 0.504578f
C398 minus.n1 gnd 0.204074f
C399 minus.n2 gnd 0.030008f
C400 minus.t19 gnd 0.504578f
C401 minus.n3 gnd 0.02439f
C402 minus.n4 gnd 0.030008f
C403 minus.t18 gnd 0.504578f
C404 minus.t5 gnd 0.504578f
C405 minus.n5 gnd 0.204074f
C406 minus.n6 gnd 0.030008f
C407 minus.t8 gnd 0.504578f
C408 minus.n7 gnd 0.204074f
C409 minus.n8 gnd 0.128812f
C410 minus.t9 gnd 0.504578f
C411 minus.t13 gnd 0.566509f
C412 minus.n9 gnd 0.236782f
C413 minus.n10 gnd 0.235673f
C414 minus.n11 gnd 0.037327f
C415 minus.n12 gnd 0.035081f
C416 minus.n13 gnd 0.030008f
C417 minus.n14 gnd 0.030008f
C418 minus.n15 gnd 0.03759f
C419 minus.n16 gnd 0.02439f
C420 minus.n17 gnd 0.038604f
C421 minus.n18 gnd 0.030008f
C422 minus.n19 gnd 0.030008f
C423 minus.n20 gnd 0.036204f
C424 minus.n21 gnd 0.036204f
C425 minus.n22 gnd 0.204074f
C426 minus.n23 gnd 0.038604f
C427 minus.n24 gnd 0.030008f
C428 minus.n25 gnd 0.030008f
C429 minus.n26 gnd 0.030008f
C430 minus.n27 gnd 0.03759f
C431 minus.n28 gnd 0.204074f
C432 minus.n29 gnd 0.035081f
C433 minus.n30 gnd 0.037327f
C434 minus.n31 gnd 0.030008f
C435 minus.n32 gnd 0.030008f
C436 minus.n33 gnd 0.039081f
C437 minus.n34 gnd 0.012429f
C438 minus.t17 gnd 0.545701f
C439 minus.n35 gnd 0.237023f
C440 minus.n36 gnd 0.352598f
C441 minus.n37 gnd 0.030008f
C442 minus.t15 gnd 0.545701f
C443 minus.t12 gnd 0.504578f
C444 minus.n38 gnd 0.204074f
C445 minus.n39 gnd 0.030008f
C446 minus.t7 gnd 0.504578f
C447 minus.n40 gnd 0.02439f
C448 minus.n41 gnd 0.030008f
C449 minus.t6 gnd 0.504578f
C450 minus.t11 gnd 0.504578f
C451 minus.n42 gnd 0.204074f
C452 minus.n43 gnd 0.030008f
C453 minus.t10 gnd 0.504578f
C454 minus.n44 gnd 0.204074f
C455 minus.n45 gnd 0.128812f
C456 minus.t16 gnd 0.504578f
C457 minus.t20 gnd 0.566509f
C458 minus.n46 gnd 0.236782f
C459 minus.n47 gnd 0.235673f
C460 minus.n48 gnd 0.037327f
C461 minus.n49 gnd 0.035081f
C462 minus.n50 gnd 0.030008f
C463 minus.n51 gnd 0.030008f
C464 minus.n52 gnd 0.03759f
C465 minus.n53 gnd 0.02439f
C466 minus.n54 gnd 0.038604f
C467 minus.n55 gnd 0.030008f
C468 minus.n56 gnd 0.030008f
C469 minus.n57 gnd 0.036204f
C470 minus.n58 gnd 0.036204f
C471 minus.n59 gnd 0.204074f
C472 minus.n60 gnd 0.038604f
C473 minus.n61 gnd 0.030008f
C474 minus.n62 gnd 0.030008f
C475 minus.n63 gnd 0.030008f
C476 minus.n64 gnd 0.03759f
C477 minus.n65 gnd 0.204074f
C478 minus.n66 gnd 0.035081f
C479 minus.n67 gnd 0.037327f
C480 minus.n68 gnd 0.030008f
C481 minus.n69 gnd 0.030008f
C482 minus.n70 gnd 0.039081f
C483 minus.n71 gnd 0.012429f
C484 minus.n72 gnd 0.237023f
C485 minus.n73 gnd 0.935033f
C486 minus.n74 gnd 1.40543f
C487 minus.t1 gnd 0.009251f
C488 minus.t4 gnd 0.009251f
C489 minus.n75 gnd 0.030418f
C490 minus.t2 gnd 0.009251f
C491 minus.t0 gnd 0.009251f
C492 minus.n76 gnd 0.030001f
C493 minus.n77 gnd 0.256047f
C494 minus.t3 gnd 0.051488f
C495 minus.n78 gnd 0.139722f
C496 minus.n79 gnd 1.86779f
C497 diffpairibias.t27 gnd 0.090128f
C498 diffpairibias.t23 gnd 0.08996f
C499 diffpairibias.n0 gnd 0.105991f
C500 diffpairibias.t28 gnd 0.08996f
C501 diffpairibias.n1 gnd 0.051736f
C502 diffpairibias.t25 gnd 0.08996f
C503 diffpairibias.n2 gnd 0.051736f
C504 diffpairibias.t29 gnd 0.08996f
C505 diffpairibias.n3 gnd 0.041084f
C506 diffpairibias.t15 gnd 0.086371f
C507 diffpairibias.t1 gnd 0.085993f
C508 diffpairibias.n4 gnd 0.13579f
C509 diffpairibias.t11 gnd 0.085993f
C510 diffpairibias.n5 gnd 0.072463f
C511 diffpairibias.t13 gnd 0.085993f
C512 diffpairibias.n6 gnd 0.072463f
C513 diffpairibias.t7 gnd 0.085993f
C514 diffpairibias.n7 gnd 0.072463f
C515 diffpairibias.t3 gnd 0.085993f
C516 diffpairibias.n8 gnd 0.072463f
C517 diffpairibias.t17 gnd 0.085993f
C518 diffpairibias.n9 gnd 0.072463f
C519 diffpairibias.t5 gnd 0.085993f
C520 diffpairibias.n10 gnd 0.072463f
C521 diffpairibias.t19 gnd 0.085993f
C522 diffpairibias.n11 gnd 0.072463f
C523 diffpairibias.t9 gnd 0.085993f
C524 diffpairibias.n12 gnd 0.102883f
C525 diffpairibias.t14 gnd 0.086899f
C526 diffpairibias.t0 gnd 0.086748f
C527 diffpairibias.n13 gnd 0.094648f
C528 diffpairibias.t10 gnd 0.086748f
C529 diffpairibias.n14 gnd 0.052262f
C530 diffpairibias.t12 gnd 0.086748f
C531 diffpairibias.n15 gnd 0.052262f
C532 diffpairibias.t6 gnd 0.086748f
C533 diffpairibias.n16 gnd 0.052262f
C534 diffpairibias.t2 gnd 0.086748f
C535 diffpairibias.n17 gnd 0.052262f
C536 diffpairibias.t16 gnd 0.086748f
C537 diffpairibias.n18 gnd 0.052262f
C538 diffpairibias.t4 gnd 0.086748f
C539 diffpairibias.n19 gnd 0.052262f
C540 diffpairibias.t18 gnd 0.086748f
C541 diffpairibias.n20 gnd 0.052262f
C542 diffpairibias.t8 gnd 0.086748f
C543 diffpairibias.n21 gnd 0.061849f
C544 diffpairibias.n22 gnd 0.233513f
C545 diffpairibias.t20 gnd 0.08996f
C546 diffpairibias.n23 gnd 0.051747f
C547 diffpairibias.t26 gnd 0.08996f
C548 diffpairibias.n24 gnd 0.051736f
C549 diffpairibias.t22 gnd 0.08996f
C550 diffpairibias.n25 gnd 0.051736f
C551 diffpairibias.t21 gnd 0.08996f
C552 diffpairibias.n26 gnd 0.051736f
C553 diffpairibias.t24 gnd 0.08996f
C554 diffpairibias.n27 gnd 0.04729f
C555 diffpairibias.n28 gnd 0.047711f
C556 a_n3827_n3924.n0 gnd 0.8843f
C557 a_n3827_n3924.t11 gnd 0.083157f
C558 a_n3827_n3924.t20 gnd 0.864269f
C559 a_n3827_n3924.n1 gnd 0.326732f
C560 a_n3827_n3924.t25 gnd 1.07678f
C561 a_n3827_n3924.t29 gnd 1.07383f
C562 a_n3827_n3924.n2 gnd 1.46419f
C563 a_n3827_n3924.n3 gnd 0.408778f
C564 a_n3827_n3924.t41 gnd 0.864269f
C565 a_n3827_n3924.n4 gnd 0.326732f
C566 a_n3827_n3924.t0 gnd 0.083157f
C567 a_n3827_n3924.t32 gnd 0.083157f
C568 a_n3827_n3924.n5 gnd 0.67916f
C569 a_n3827_n3924.n6 gnd 0.342258f
C570 a_n3827_n3924.t40 gnd 0.083157f
C571 a_n3827_n3924.t31 gnd 0.083157f
C572 a_n3827_n3924.n7 gnd 0.67916f
C573 a_n3827_n3924.n8 gnd 0.342258f
C574 a_n3827_n3924.t39 gnd 0.083157f
C575 a_n3827_n3924.t1 gnd 0.083157f
C576 a_n3827_n3924.n9 gnd 0.67916f
C577 a_n3827_n3924.n10 gnd 0.342258f
C578 a_n3827_n3924.t30 gnd 0.864269f
C579 a_n3827_n3924.n11 gnd 0.809022f
C580 a_n3827_n3924.t38 gnd 1.07537f
C581 a_n3827_n3924.t3 gnd 1.07383f
C582 a_n3827_n3924.n12 gnd 1.24022f
C583 a_n3827_n3924.t27 gnd 1.07383f
C584 a_n3827_n3924.n13 gnd 0.700903f
C585 a_n3827_n3924.t8 gnd 1.07383f
C586 a_n3827_n3924.n14 gnd 0.75632f
C587 a_n3827_n3924.t2 gnd 1.07383f
C588 a_n3827_n3924.n15 gnd 0.75632f
C589 a_n3827_n3924.t7 gnd 1.07383f
C590 a_n3827_n3924.n16 gnd 0.75632f
C591 a_n3827_n3924.t6 gnd 1.07383f
C592 a_n3827_n3924.n17 gnd 0.75632f
C593 a_n3827_n3924.t37 gnd 1.07383f
C594 a_n3827_n3924.n18 gnd 0.783961f
C595 a_n3827_n3924.t22 gnd 0.864266f
C596 a_n3827_n3924.n19 gnd 0.536839f
C597 a_n3827_n3924.t23 gnd 0.083157f
C598 a_n3827_n3924.t13 gnd 0.083157f
C599 a_n3827_n3924.n20 gnd 0.679159f
C600 a_n3827_n3924.n21 gnd 0.342259f
C601 a_n3827_n3924.t14 gnd 0.083157f
C602 a_n3827_n3924.t9 gnd 0.083157f
C603 a_n3827_n3924.n22 gnd 0.679159f
C604 a_n3827_n3924.n23 gnd 0.342259f
C605 a_n3827_n3924.t10 gnd 0.083157f
C606 a_n3827_n3924.t21 gnd 0.083157f
C607 a_n3827_n3924.n24 gnd 0.679159f
C608 a_n3827_n3924.n25 gnd 0.342259f
C609 a_n3827_n3924.t18 gnd 0.864266f
C610 a_n3827_n3924.n26 gnd 0.326736f
C611 a_n3827_n3924.t4 gnd 0.864266f
C612 a_n3827_n3924.n27 gnd 0.326736f
C613 a_n3827_n3924.t36 gnd 0.083157f
C614 a_n3827_n3924.t5 gnd 0.083157f
C615 a_n3827_n3924.n28 gnd 0.679159f
C616 a_n3827_n3924.n29 gnd 0.342259f
C617 a_n3827_n3924.t34 gnd 0.083157f
C618 a_n3827_n3924.t35 gnd 0.083157f
C619 a_n3827_n3924.n30 gnd 0.679159f
C620 a_n3827_n3924.n31 gnd 0.342259f
C621 a_n3827_n3924.t26 gnd 0.083157f
C622 a_n3827_n3924.t28 gnd 0.083157f
C623 a_n3827_n3924.n32 gnd 0.679159f
C624 a_n3827_n3924.n33 gnd 0.342259f
C625 a_n3827_n3924.t33 gnd 0.864266f
C626 a_n3827_n3924.n34 gnd 0.536839f
C627 a_n3827_n3924.n35 gnd 0.783961f
C628 a_n3827_n3924.t17 gnd 0.864266f
C629 a_n3827_n3924.n36 gnd 0.809025f
C630 a_n3827_n3924.t15 gnd 0.083157f
C631 a_n3827_n3924.t19 gnd 0.083157f
C632 a_n3827_n3924.n37 gnd 0.67916f
C633 a_n3827_n3924.n38 gnd 0.342258f
C634 a_n3827_n3924.t12 gnd 0.083157f
C635 a_n3827_n3924.t16 gnd 0.083157f
C636 a_n3827_n3924.n39 gnd 0.67916f
C637 a_n3827_n3924.n40 gnd 0.342258f
C638 a_n3827_n3924.n41 gnd 0.342257f
C639 a_n3827_n3924.n42 gnd 0.679161f
C640 a_n3827_n3924.t24 gnd 0.083157f
C641 plus.n0 gnd 0.022063f
C642 plus.t7 gnd 0.401225f
C643 plus.t6 gnd 0.37099f
C644 plus.n1 gnd 0.150045f
C645 plus.n2 gnd 0.022063f
C646 plus.t16 gnd 0.37099f
C647 plus.n3 gnd 0.017933f
C648 plus.n4 gnd 0.022063f
C649 plus.t15 gnd 0.37099f
C650 plus.t20 gnd 0.37099f
C651 plus.n5 gnd 0.150045f
C652 plus.n6 gnd 0.022063f
C653 plus.t19 gnd 0.37099f
C654 plus.n7 gnd 0.150045f
C655 plus.n8 gnd 0.094709f
C656 plus.t8 gnd 0.37099f
C657 plus.t11 gnd 0.416524f
C658 plus.n9 gnd 0.174093f
C659 plus.n10 gnd 0.173278f
C660 plus.n11 gnd 0.027445f
C661 plus.n12 gnd 0.025793f
C662 plus.n13 gnd 0.022063f
C663 plus.n14 gnd 0.022063f
C664 plus.n15 gnd 0.027638f
C665 plus.n16 gnd 0.017933f
C666 plus.n17 gnd 0.028383f
C667 plus.n18 gnd 0.022063f
C668 plus.n19 gnd 0.022063f
C669 plus.n20 gnd 0.026619f
C670 plus.n21 gnd 0.026619f
C671 plus.n22 gnd 0.150045f
C672 plus.n23 gnd 0.028383f
C673 plus.n24 gnd 0.022063f
C674 plus.n25 gnd 0.022063f
C675 plus.n26 gnd 0.022063f
C676 plus.n27 gnd 0.027638f
C677 plus.n28 gnd 0.150045f
C678 plus.n29 gnd 0.025793f
C679 plus.n30 gnd 0.027445f
C680 plus.n31 gnd 0.022063f
C681 plus.n32 gnd 0.022063f
C682 plus.n33 gnd 0.028734f
C683 plus.n34 gnd 0.009138f
C684 plus.n35 gnd 0.174271f
C685 plus.n36 gnd 0.253573f
C686 plus.n37 gnd 0.022063f
C687 plus.t10 gnd 0.37099f
C688 plus.n38 gnd 0.150045f
C689 plus.n39 gnd 0.022063f
C690 plus.t14 gnd 0.37099f
C691 plus.n40 gnd 0.017933f
C692 plus.n41 gnd 0.022063f
C693 plus.t13 gnd 0.37099f
C694 plus.t17 gnd 0.37099f
C695 plus.n42 gnd 0.150045f
C696 plus.n43 gnd 0.022063f
C697 plus.t18 gnd 0.37099f
C698 plus.n44 gnd 0.150045f
C699 plus.n45 gnd 0.094709f
C700 plus.t5 gnd 0.37099f
C701 plus.t9 gnd 0.416524f
C702 plus.n46 gnd 0.174093f
C703 plus.n47 gnd 0.173278f
C704 plus.n48 gnd 0.027445f
C705 plus.n49 gnd 0.025793f
C706 plus.n50 gnd 0.022063f
C707 plus.n51 gnd 0.022063f
C708 plus.n52 gnd 0.027638f
C709 plus.n53 gnd 0.017933f
C710 plus.n54 gnd 0.028383f
C711 plus.n55 gnd 0.022063f
C712 plus.n56 gnd 0.022063f
C713 plus.n57 gnd 0.026619f
C714 plus.n58 gnd 0.026619f
C715 plus.n59 gnd 0.150045f
C716 plus.n60 gnd 0.028383f
C717 plus.n61 gnd 0.022063f
C718 plus.n62 gnd 0.022063f
C719 plus.n63 gnd 0.022063f
C720 plus.n64 gnd 0.027638f
C721 plus.n65 gnd 0.150045f
C722 plus.n66 gnd 0.025793f
C723 plus.n67 gnd 0.027445f
C724 plus.n68 gnd 0.022063f
C725 plus.n69 gnd 0.022063f
C726 plus.n70 gnd 0.028734f
C727 plus.n71 gnd 0.009138f
C728 plus.t12 gnd 0.401225f
C729 plus.n72 gnd 0.174271f
C730 plus.n73 gnd 0.67864f
C731 plus.n74 gnd 1.02459f
C732 plus.t4 gnd 0.038088f
C733 plus.t1 gnd 0.006801f
C734 plus.t2 gnd 0.006801f
C735 plus.n75 gnd 0.022058f
C736 plus.n76 gnd 0.17124f
C737 plus.t0 gnd 0.006801f
C738 plus.t3 gnd 0.006801f
C739 plus.n77 gnd 0.022058f
C740 plus.n78 gnd 0.128537f
C741 plus.n79 gnd 2.4535f
C742 commonsourceibias.n0 gnd 0.012299f
C743 commonsourceibias.t56 gnd 0.18623f
C744 commonsourceibias.t109 gnd 0.172196f
C745 commonsourceibias.n1 gnd 0.068706f
C746 commonsourceibias.n2 gnd 0.009217f
C747 commonsourceibias.t69 gnd 0.172196f
C748 commonsourceibias.n3 gnd 0.007456f
C749 commonsourceibias.n4 gnd 0.009217f
C750 commonsourceibias.t119 gnd 0.172196f
C751 commonsourceibias.n5 gnd 0.008898f
C752 commonsourceibias.n6 gnd 0.009217f
C753 commonsourceibias.t85 gnd 0.172196f
C754 commonsourceibias.n7 gnd 0.068706f
C755 commonsourceibias.t54 gnd 0.172196f
C756 commonsourceibias.n8 gnd 0.007444f
C757 commonsourceibias.n9 gnd 0.012299f
C758 commonsourceibias.t28 gnd 0.18623f
C759 commonsourceibias.t4 gnd 0.172196f
C760 commonsourceibias.n10 gnd 0.068706f
C761 commonsourceibias.n11 gnd 0.009217f
C762 commonsourceibias.t42 gnd 0.172196f
C763 commonsourceibias.n12 gnd 0.007456f
C764 commonsourceibias.n13 gnd 0.009217f
C765 commonsourceibias.t40 gnd 0.172196f
C766 commonsourceibias.n14 gnd 0.008898f
C767 commonsourceibias.n15 gnd 0.009217f
C768 commonsourceibias.t16 gnd 0.172196f
C769 commonsourceibias.n16 gnd 0.068706f
C770 commonsourceibias.t22 gnd 0.172196f
C771 commonsourceibias.n17 gnd 0.007444f
C772 commonsourceibias.n18 gnd 0.009217f
C773 commonsourceibias.t34 gnd 0.172196f
C774 commonsourceibias.t14 gnd 0.172196f
C775 commonsourceibias.n19 gnd 0.068706f
C776 commonsourceibias.n20 gnd 0.009217f
C777 commonsourceibias.t6 gnd 0.172196f
C778 commonsourceibias.n21 gnd 0.068706f
C779 commonsourceibias.n22 gnd 0.009217f
C780 commonsourceibias.t18 gnd 0.172196f
C781 commonsourceibias.n23 gnd 0.068706f
C782 commonsourceibias.n24 gnd 0.046399f
C783 commonsourceibias.t46 gnd 0.172196f
C784 commonsourceibias.t38 gnd 0.194303f
C785 commonsourceibias.n25 gnd 0.079733f
C786 commonsourceibias.n26 gnd 0.082545f
C787 commonsourceibias.n27 gnd 0.01136f
C788 commonsourceibias.n28 gnd 0.012567f
C789 commonsourceibias.n29 gnd 0.009217f
C790 commonsourceibias.n30 gnd 0.009217f
C791 commonsourceibias.n31 gnd 0.012485f
C792 commonsourceibias.n32 gnd 0.007456f
C793 commonsourceibias.n33 gnd 0.01264f
C794 commonsourceibias.n34 gnd 0.009217f
C795 commonsourceibias.n35 gnd 0.009217f
C796 commonsourceibias.n36 gnd 0.012717f
C797 commonsourceibias.n37 gnd 0.010966f
C798 commonsourceibias.n38 gnd 0.008898f
C799 commonsourceibias.n39 gnd 0.009217f
C800 commonsourceibias.n40 gnd 0.009217f
C801 commonsourceibias.n41 gnd 0.011274f
C802 commonsourceibias.n42 gnd 0.012653f
C803 commonsourceibias.n43 gnd 0.068706f
C804 commonsourceibias.n44 gnd 0.012568f
C805 commonsourceibias.n45 gnd 0.009217f
C806 commonsourceibias.n46 gnd 0.009217f
C807 commonsourceibias.n47 gnd 0.009217f
C808 commonsourceibias.n48 gnd 0.012568f
C809 commonsourceibias.n49 gnd 0.068706f
C810 commonsourceibias.n50 gnd 0.012653f
C811 commonsourceibias.n51 gnd 0.011274f
C812 commonsourceibias.n52 gnd 0.009217f
C813 commonsourceibias.n53 gnd 0.009217f
C814 commonsourceibias.n54 gnd 0.009217f
C815 commonsourceibias.n55 gnd 0.010966f
C816 commonsourceibias.n56 gnd 0.012717f
C817 commonsourceibias.n57 gnd 0.068706f
C818 commonsourceibias.n58 gnd 0.01264f
C819 commonsourceibias.n59 gnd 0.009217f
C820 commonsourceibias.n60 gnd 0.009217f
C821 commonsourceibias.n61 gnd 0.009217f
C822 commonsourceibias.n62 gnd 0.012485f
C823 commonsourceibias.n63 gnd 0.068706f
C824 commonsourceibias.n64 gnd 0.012567f
C825 commonsourceibias.n65 gnd 0.01136f
C826 commonsourceibias.n66 gnd 0.009217f
C827 commonsourceibias.n67 gnd 0.009217f
C828 commonsourceibias.n68 gnd 0.009349f
C829 commonsourceibias.n69 gnd 0.009666f
C830 commonsourceibias.n70 gnd 0.082208f
C831 commonsourceibias.n71 gnd 0.091197f
C832 commonsourceibias.t29 gnd 0.019889f
C833 commonsourceibias.t5 gnd 0.019889f
C834 commonsourceibias.n72 gnd 0.175743f
C835 commonsourceibias.n73 gnd 0.151855f
C836 commonsourceibias.t43 gnd 0.019889f
C837 commonsourceibias.t41 gnd 0.019889f
C838 commonsourceibias.n74 gnd 0.175743f
C839 commonsourceibias.n75 gnd 0.080726f
C840 commonsourceibias.t17 gnd 0.019889f
C841 commonsourceibias.t23 gnd 0.019889f
C842 commonsourceibias.n76 gnd 0.175743f
C843 commonsourceibias.n77 gnd 0.067443f
C844 commonsourceibias.t47 gnd 0.019889f
C845 commonsourceibias.t39 gnd 0.019889f
C846 commonsourceibias.n78 gnd 0.176331f
C847 commonsourceibias.t7 gnd 0.019889f
C848 commonsourceibias.t19 gnd 0.019889f
C849 commonsourceibias.n79 gnd 0.175743f
C850 commonsourceibias.n80 gnd 0.16376f
C851 commonsourceibias.t35 gnd 0.019889f
C852 commonsourceibias.t15 gnd 0.019889f
C853 commonsourceibias.n81 gnd 0.175743f
C854 commonsourceibias.n82 gnd 0.067443f
C855 commonsourceibias.n83 gnd 0.081666f
C856 commonsourceibias.n84 gnd 0.009217f
C857 commonsourceibias.t100 gnd 0.172196f
C858 commonsourceibias.t87 gnd 0.172196f
C859 commonsourceibias.n85 gnd 0.068706f
C860 commonsourceibias.n86 gnd 0.009217f
C861 commonsourceibias.t115 gnd 0.172196f
C862 commonsourceibias.n87 gnd 0.068706f
C863 commonsourceibias.n88 gnd 0.009217f
C864 commonsourceibias.t79 gnd 0.172196f
C865 commonsourceibias.n89 gnd 0.068706f
C866 commonsourceibias.n90 gnd 0.046399f
C867 commonsourceibias.t66 gnd 0.172196f
C868 commonsourceibias.t95 gnd 0.194303f
C869 commonsourceibias.n91 gnd 0.079733f
C870 commonsourceibias.n92 gnd 0.082545f
C871 commonsourceibias.n93 gnd 0.01136f
C872 commonsourceibias.n94 gnd 0.012567f
C873 commonsourceibias.n95 gnd 0.009217f
C874 commonsourceibias.n96 gnd 0.009217f
C875 commonsourceibias.n97 gnd 0.012485f
C876 commonsourceibias.n98 gnd 0.007456f
C877 commonsourceibias.n99 gnd 0.01264f
C878 commonsourceibias.n100 gnd 0.009217f
C879 commonsourceibias.n101 gnd 0.009217f
C880 commonsourceibias.n102 gnd 0.012717f
C881 commonsourceibias.n103 gnd 0.010966f
C882 commonsourceibias.n104 gnd 0.008898f
C883 commonsourceibias.n105 gnd 0.009217f
C884 commonsourceibias.n106 gnd 0.009217f
C885 commonsourceibias.n107 gnd 0.011274f
C886 commonsourceibias.n108 gnd 0.012653f
C887 commonsourceibias.n109 gnd 0.068706f
C888 commonsourceibias.n110 gnd 0.012568f
C889 commonsourceibias.n111 gnd 0.009172f
C890 commonsourceibias.n112 gnd 0.066626f
C891 commonsourceibias.n113 gnd 0.009172f
C892 commonsourceibias.n114 gnd 0.012568f
C893 commonsourceibias.n115 gnd 0.068706f
C894 commonsourceibias.n116 gnd 0.012653f
C895 commonsourceibias.n117 gnd 0.011274f
C896 commonsourceibias.n118 gnd 0.009217f
C897 commonsourceibias.n119 gnd 0.009217f
C898 commonsourceibias.n120 gnd 0.009217f
C899 commonsourceibias.n121 gnd 0.010966f
C900 commonsourceibias.n122 gnd 0.012717f
C901 commonsourceibias.n123 gnd 0.068706f
C902 commonsourceibias.n124 gnd 0.01264f
C903 commonsourceibias.n125 gnd 0.009217f
C904 commonsourceibias.n126 gnd 0.009217f
C905 commonsourceibias.n127 gnd 0.009217f
C906 commonsourceibias.n128 gnd 0.012485f
C907 commonsourceibias.n129 gnd 0.068706f
C908 commonsourceibias.n130 gnd 0.012567f
C909 commonsourceibias.n131 gnd 0.01136f
C910 commonsourceibias.n132 gnd 0.009217f
C911 commonsourceibias.n133 gnd 0.009217f
C912 commonsourceibias.n134 gnd 0.009349f
C913 commonsourceibias.n135 gnd 0.009666f
C914 commonsourceibias.n136 gnd 0.082208f
C915 commonsourceibias.n137 gnd 0.05322f
C916 commonsourceibias.n138 gnd 0.012299f
C917 commonsourceibias.t89 gnd 0.18623f
C918 commonsourceibias.t106 gnd 0.172196f
C919 commonsourceibias.n139 gnd 0.068706f
C920 commonsourceibias.n140 gnd 0.009217f
C921 commonsourceibias.t101 gnd 0.172196f
C922 commonsourceibias.n141 gnd 0.007456f
C923 commonsourceibias.n142 gnd 0.009217f
C924 commonsourceibias.t88 gnd 0.172196f
C925 commonsourceibias.n143 gnd 0.008898f
C926 commonsourceibias.n144 gnd 0.009217f
C927 commonsourceibias.t105 gnd 0.172196f
C928 commonsourceibias.n145 gnd 0.068706f
C929 commonsourceibias.t99 gnd 0.172196f
C930 commonsourceibias.n146 gnd 0.007444f
C931 commonsourceibias.n147 gnd 0.009217f
C932 commonsourceibias.t86 gnd 0.172196f
C933 commonsourceibias.t108 gnd 0.172196f
C934 commonsourceibias.n148 gnd 0.068706f
C935 commonsourceibias.n149 gnd 0.009217f
C936 commonsourceibias.t98 gnd 0.172196f
C937 commonsourceibias.n150 gnd 0.068706f
C938 commonsourceibias.n151 gnd 0.009217f
C939 commonsourceibias.t112 gnd 0.172196f
C940 commonsourceibias.n152 gnd 0.068706f
C941 commonsourceibias.n153 gnd 0.046399f
C942 commonsourceibias.t107 gnd 0.172196f
C943 commonsourceibias.t97 gnd 0.194303f
C944 commonsourceibias.n154 gnd 0.079733f
C945 commonsourceibias.n155 gnd 0.082545f
C946 commonsourceibias.n156 gnd 0.01136f
C947 commonsourceibias.n157 gnd 0.012567f
C948 commonsourceibias.n158 gnd 0.009217f
C949 commonsourceibias.n159 gnd 0.009217f
C950 commonsourceibias.n160 gnd 0.012485f
C951 commonsourceibias.n161 gnd 0.007456f
C952 commonsourceibias.n162 gnd 0.01264f
C953 commonsourceibias.n163 gnd 0.009217f
C954 commonsourceibias.n164 gnd 0.009217f
C955 commonsourceibias.n165 gnd 0.012717f
C956 commonsourceibias.n166 gnd 0.010966f
C957 commonsourceibias.n167 gnd 0.008898f
C958 commonsourceibias.n168 gnd 0.009217f
C959 commonsourceibias.n169 gnd 0.009217f
C960 commonsourceibias.n170 gnd 0.011274f
C961 commonsourceibias.n171 gnd 0.012653f
C962 commonsourceibias.n172 gnd 0.068706f
C963 commonsourceibias.n173 gnd 0.012568f
C964 commonsourceibias.n174 gnd 0.009217f
C965 commonsourceibias.n175 gnd 0.009217f
C966 commonsourceibias.n176 gnd 0.009217f
C967 commonsourceibias.n177 gnd 0.012568f
C968 commonsourceibias.n178 gnd 0.068706f
C969 commonsourceibias.n179 gnd 0.012653f
C970 commonsourceibias.n180 gnd 0.011274f
C971 commonsourceibias.n181 gnd 0.009217f
C972 commonsourceibias.n182 gnd 0.009217f
C973 commonsourceibias.n183 gnd 0.009217f
C974 commonsourceibias.n184 gnd 0.010966f
C975 commonsourceibias.n185 gnd 0.012717f
C976 commonsourceibias.n186 gnd 0.068706f
C977 commonsourceibias.n187 gnd 0.01264f
C978 commonsourceibias.n188 gnd 0.009217f
C979 commonsourceibias.n189 gnd 0.009217f
C980 commonsourceibias.n190 gnd 0.009217f
C981 commonsourceibias.n191 gnd 0.012485f
C982 commonsourceibias.n192 gnd 0.068706f
C983 commonsourceibias.n193 gnd 0.012567f
C984 commonsourceibias.n194 gnd 0.01136f
C985 commonsourceibias.n195 gnd 0.009217f
C986 commonsourceibias.n196 gnd 0.009217f
C987 commonsourceibias.n197 gnd 0.009349f
C988 commonsourceibias.n198 gnd 0.009666f
C989 commonsourceibias.n199 gnd 0.082208f
C990 commonsourceibias.n200 gnd 0.027976f
C991 commonsourceibias.n201 gnd 0.147064f
C992 commonsourceibias.n202 gnd 0.012299f
C993 commonsourceibias.t50 gnd 0.172196f
C994 commonsourceibias.n203 gnd 0.068706f
C995 commonsourceibias.n204 gnd 0.009217f
C996 commonsourceibias.t60 gnd 0.172196f
C997 commonsourceibias.n205 gnd 0.007456f
C998 commonsourceibias.n206 gnd 0.009217f
C999 commonsourceibias.t104 gnd 0.172196f
C1000 commonsourceibias.n207 gnd 0.008898f
C1001 commonsourceibias.n208 gnd 0.009217f
C1002 commonsourceibias.t118 gnd 0.172196f
C1003 commonsourceibias.n209 gnd 0.068706f
C1004 commonsourceibias.t52 gnd 0.172196f
C1005 commonsourceibias.n210 gnd 0.007444f
C1006 commonsourceibias.n211 gnd 0.009217f
C1007 commonsourceibias.t93 gnd 0.172196f
C1008 commonsourceibias.t84 gnd 0.172196f
C1009 commonsourceibias.n212 gnd 0.068706f
C1010 commonsourceibias.n213 gnd 0.009217f
C1011 commonsourceibias.t49 gnd 0.172196f
C1012 commonsourceibias.n214 gnd 0.068706f
C1013 commonsourceibias.n215 gnd 0.009217f
C1014 commonsourceibias.t59 gnd 0.172196f
C1015 commonsourceibias.n216 gnd 0.068706f
C1016 commonsourceibias.n217 gnd 0.046399f
C1017 commonsourceibias.t75 gnd 0.172196f
C1018 commonsourceibias.t117 gnd 0.194303f
C1019 commonsourceibias.n218 gnd 0.079733f
C1020 commonsourceibias.n219 gnd 0.082545f
C1021 commonsourceibias.n220 gnd 0.01136f
C1022 commonsourceibias.n221 gnd 0.012567f
C1023 commonsourceibias.n222 gnd 0.009217f
C1024 commonsourceibias.n223 gnd 0.009217f
C1025 commonsourceibias.n224 gnd 0.012485f
C1026 commonsourceibias.n225 gnd 0.007456f
C1027 commonsourceibias.n226 gnd 0.01264f
C1028 commonsourceibias.n227 gnd 0.009217f
C1029 commonsourceibias.n228 gnd 0.009217f
C1030 commonsourceibias.n229 gnd 0.012717f
C1031 commonsourceibias.n230 gnd 0.010966f
C1032 commonsourceibias.n231 gnd 0.008898f
C1033 commonsourceibias.n232 gnd 0.009217f
C1034 commonsourceibias.n233 gnd 0.009217f
C1035 commonsourceibias.n234 gnd 0.011274f
C1036 commonsourceibias.n235 gnd 0.012653f
C1037 commonsourceibias.n236 gnd 0.068706f
C1038 commonsourceibias.n237 gnd 0.012568f
C1039 commonsourceibias.n238 gnd 0.009217f
C1040 commonsourceibias.n239 gnd 0.009217f
C1041 commonsourceibias.n240 gnd 0.009217f
C1042 commonsourceibias.n241 gnd 0.012568f
C1043 commonsourceibias.n242 gnd 0.068706f
C1044 commonsourceibias.n243 gnd 0.012653f
C1045 commonsourceibias.n244 gnd 0.011274f
C1046 commonsourceibias.n245 gnd 0.009217f
C1047 commonsourceibias.n246 gnd 0.009217f
C1048 commonsourceibias.n247 gnd 0.009217f
C1049 commonsourceibias.n248 gnd 0.010966f
C1050 commonsourceibias.n249 gnd 0.012717f
C1051 commonsourceibias.n250 gnd 0.068706f
C1052 commonsourceibias.n251 gnd 0.01264f
C1053 commonsourceibias.n252 gnd 0.009217f
C1054 commonsourceibias.n253 gnd 0.009217f
C1055 commonsourceibias.n254 gnd 0.009217f
C1056 commonsourceibias.n255 gnd 0.012485f
C1057 commonsourceibias.n256 gnd 0.068706f
C1058 commonsourceibias.n257 gnd 0.012567f
C1059 commonsourceibias.n258 gnd 0.01136f
C1060 commonsourceibias.n259 gnd 0.009217f
C1061 commonsourceibias.n260 gnd 0.009217f
C1062 commonsourceibias.n261 gnd 0.009349f
C1063 commonsourceibias.n262 gnd 0.009666f
C1064 commonsourceibias.t111 gnd 0.18623f
C1065 commonsourceibias.n263 gnd 0.082208f
C1066 commonsourceibias.n264 gnd 0.027976f
C1067 commonsourceibias.n265 gnd 0.517265f
C1068 commonsourceibias.n266 gnd 0.012299f
C1069 commonsourceibias.t114 gnd 0.18623f
C1070 commonsourceibias.t78 gnd 0.172196f
C1071 commonsourceibias.n267 gnd 0.068706f
C1072 commonsourceibias.n268 gnd 0.009217f
C1073 commonsourceibias.t53 gnd 0.172196f
C1074 commonsourceibias.n269 gnd 0.007456f
C1075 commonsourceibias.n270 gnd 0.009217f
C1076 commonsourceibias.t94 gnd 0.172196f
C1077 commonsourceibias.n271 gnd 0.008898f
C1078 commonsourceibias.n272 gnd 0.009217f
C1079 commonsourceibias.t113 gnd 0.172196f
C1080 commonsourceibias.n273 gnd 0.007444f
C1081 commonsourceibias.n274 gnd 0.009217f
C1082 commonsourceibias.t76 gnd 0.172196f
C1083 commonsourceibias.t65 gnd 0.172196f
C1084 commonsourceibias.n275 gnd 0.068706f
C1085 commonsourceibias.n276 gnd 0.009217f
C1086 commonsourceibias.t92 gnd 0.172196f
C1087 commonsourceibias.n277 gnd 0.068706f
C1088 commonsourceibias.n278 gnd 0.009217f
C1089 commonsourceibias.t63 gnd 0.172196f
C1090 commonsourceibias.n279 gnd 0.068706f
C1091 commonsourceibias.n280 gnd 0.046399f
C1092 commonsourceibias.t58 gnd 0.172196f
C1093 commonsourceibias.t70 gnd 0.194303f
C1094 commonsourceibias.n281 gnd 0.079733f
C1095 commonsourceibias.n282 gnd 0.082545f
C1096 commonsourceibias.n283 gnd 0.01136f
C1097 commonsourceibias.n284 gnd 0.012567f
C1098 commonsourceibias.n285 gnd 0.009217f
C1099 commonsourceibias.n286 gnd 0.009217f
C1100 commonsourceibias.n287 gnd 0.012485f
C1101 commonsourceibias.n288 gnd 0.007456f
C1102 commonsourceibias.n289 gnd 0.01264f
C1103 commonsourceibias.n290 gnd 0.009217f
C1104 commonsourceibias.n291 gnd 0.009217f
C1105 commonsourceibias.n292 gnd 0.012717f
C1106 commonsourceibias.n293 gnd 0.010966f
C1107 commonsourceibias.n294 gnd 0.008898f
C1108 commonsourceibias.n295 gnd 0.009217f
C1109 commonsourceibias.n296 gnd 0.009217f
C1110 commonsourceibias.n297 gnd 0.011274f
C1111 commonsourceibias.n298 gnd 0.012653f
C1112 commonsourceibias.n299 gnd 0.068706f
C1113 commonsourceibias.n300 gnd 0.012568f
C1114 commonsourceibias.n301 gnd 0.009172f
C1115 commonsourceibias.t45 gnd 0.019889f
C1116 commonsourceibias.t27 gnd 0.019889f
C1117 commonsourceibias.n302 gnd 0.176331f
C1118 commonsourceibias.t3 gnd 0.019889f
C1119 commonsourceibias.t13 gnd 0.019889f
C1120 commonsourceibias.n303 gnd 0.175743f
C1121 commonsourceibias.n304 gnd 0.16376f
C1122 commonsourceibias.t31 gnd 0.019889f
C1123 commonsourceibias.t1 gnd 0.019889f
C1124 commonsourceibias.n305 gnd 0.175743f
C1125 commonsourceibias.n306 gnd 0.067443f
C1126 commonsourceibias.n307 gnd 0.012299f
C1127 commonsourceibias.t20 gnd 0.172196f
C1128 commonsourceibias.n308 gnd 0.068706f
C1129 commonsourceibias.n309 gnd 0.009217f
C1130 commonsourceibias.t24 gnd 0.172196f
C1131 commonsourceibias.n310 gnd 0.007456f
C1132 commonsourceibias.n311 gnd 0.009217f
C1133 commonsourceibias.t36 gnd 0.172196f
C1134 commonsourceibias.n312 gnd 0.008898f
C1135 commonsourceibias.n313 gnd 0.009217f
C1136 commonsourceibias.t10 gnd 0.172196f
C1137 commonsourceibias.n314 gnd 0.007444f
C1138 commonsourceibias.n315 gnd 0.009217f
C1139 commonsourceibias.t0 gnd 0.172196f
C1140 commonsourceibias.t30 gnd 0.172196f
C1141 commonsourceibias.n316 gnd 0.068706f
C1142 commonsourceibias.n317 gnd 0.009217f
C1143 commonsourceibias.t12 gnd 0.172196f
C1144 commonsourceibias.n318 gnd 0.068706f
C1145 commonsourceibias.n319 gnd 0.009217f
C1146 commonsourceibias.t2 gnd 0.172196f
C1147 commonsourceibias.n320 gnd 0.068706f
C1148 commonsourceibias.n321 gnd 0.046399f
C1149 commonsourceibias.t26 gnd 0.172196f
C1150 commonsourceibias.t44 gnd 0.194303f
C1151 commonsourceibias.n322 gnd 0.079733f
C1152 commonsourceibias.n323 gnd 0.082545f
C1153 commonsourceibias.n324 gnd 0.01136f
C1154 commonsourceibias.n325 gnd 0.012567f
C1155 commonsourceibias.n326 gnd 0.009217f
C1156 commonsourceibias.n327 gnd 0.009217f
C1157 commonsourceibias.n328 gnd 0.012485f
C1158 commonsourceibias.n329 gnd 0.007456f
C1159 commonsourceibias.n330 gnd 0.01264f
C1160 commonsourceibias.n331 gnd 0.009217f
C1161 commonsourceibias.n332 gnd 0.009217f
C1162 commonsourceibias.n333 gnd 0.012717f
C1163 commonsourceibias.n334 gnd 0.010966f
C1164 commonsourceibias.n335 gnd 0.008898f
C1165 commonsourceibias.n336 gnd 0.009217f
C1166 commonsourceibias.n337 gnd 0.009217f
C1167 commonsourceibias.n338 gnd 0.011274f
C1168 commonsourceibias.n339 gnd 0.012653f
C1169 commonsourceibias.n340 gnd 0.068706f
C1170 commonsourceibias.n341 gnd 0.012568f
C1171 commonsourceibias.n342 gnd 0.009217f
C1172 commonsourceibias.n343 gnd 0.009217f
C1173 commonsourceibias.n344 gnd 0.009217f
C1174 commonsourceibias.n345 gnd 0.012568f
C1175 commonsourceibias.n346 gnd 0.068706f
C1176 commonsourceibias.n347 gnd 0.012653f
C1177 commonsourceibias.t32 gnd 0.172196f
C1178 commonsourceibias.n348 gnd 0.068706f
C1179 commonsourceibias.n349 gnd 0.011274f
C1180 commonsourceibias.n350 gnd 0.009217f
C1181 commonsourceibias.n351 gnd 0.009217f
C1182 commonsourceibias.n352 gnd 0.009217f
C1183 commonsourceibias.n353 gnd 0.010966f
C1184 commonsourceibias.n354 gnd 0.012717f
C1185 commonsourceibias.n355 gnd 0.068706f
C1186 commonsourceibias.n356 gnd 0.01264f
C1187 commonsourceibias.n357 gnd 0.009217f
C1188 commonsourceibias.n358 gnd 0.009217f
C1189 commonsourceibias.n359 gnd 0.009217f
C1190 commonsourceibias.n360 gnd 0.012485f
C1191 commonsourceibias.n361 gnd 0.068706f
C1192 commonsourceibias.n362 gnd 0.012567f
C1193 commonsourceibias.n363 gnd 0.01136f
C1194 commonsourceibias.n364 gnd 0.009217f
C1195 commonsourceibias.n365 gnd 0.009217f
C1196 commonsourceibias.n366 gnd 0.009349f
C1197 commonsourceibias.n367 gnd 0.009666f
C1198 commonsourceibias.t8 gnd 0.18623f
C1199 commonsourceibias.n368 gnd 0.082208f
C1200 commonsourceibias.n369 gnd 0.091197f
C1201 commonsourceibias.t21 gnd 0.019889f
C1202 commonsourceibias.t9 gnd 0.019889f
C1203 commonsourceibias.n370 gnd 0.175743f
C1204 commonsourceibias.n371 gnd 0.151855f
C1205 commonsourceibias.t37 gnd 0.019889f
C1206 commonsourceibias.t25 gnd 0.019889f
C1207 commonsourceibias.n372 gnd 0.175743f
C1208 commonsourceibias.n373 gnd 0.080726f
C1209 commonsourceibias.t11 gnd 0.019889f
C1210 commonsourceibias.t33 gnd 0.019889f
C1211 commonsourceibias.n374 gnd 0.175743f
C1212 commonsourceibias.n375 gnd 0.067443f
C1213 commonsourceibias.n376 gnd 0.081666f
C1214 commonsourceibias.n377 gnd 0.066626f
C1215 commonsourceibias.n378 gnd 0.009172f
C1216 commonsourceibias.n379 gnd 0.012568f
C1217 commonsourceibias.n380 gnd 0.068706f
C1218 commonsourceibias.n381 gnd 0.012653f
C1219 commonsourceibias.t64 gnd 0.172196f
C1220 commonsourceibias.n382 gnd 0.068706f
C1221 commonsourceibias.n383 gnd 0.011274f
C1222 commonsourceibias.n384 gnd 0.009217f
C1223 commonsourceibias.n385 gnd 0.009217f
C1224 commonsourceibias.n386 gnd 0.009217f
C1225 commonsourceibias.n387 gnd 0.010966f
C1226 commonsourceibias.n388 gnd 0.012717f
C1227 commonsourceibias.n389 gnd 0.068706f
C1228 commonsourceibias.n390 gnd 0.01264f
C1229 commonsourceibias.n391 gnd 0.009217f
C1230 commonsourceibias.n392 gnd 0.009217f
C1231 commonsourceibias.n393 gnd 0.009217f
C1232 commonsourceibias.n394 gnd 0.012485f
C1233 commonsourceibias.n395 gnd 0.068706f
C1234 commonsourceibias.n396 gnd 0.012567f
C1235 commonsourceibias.n397 gnd 0.01136f
C1236 commonsourceibias.n398 gnd 0.009217f
C1237 commonsourceibias.n399 gnd 0.009217f
C1238 commonsourceibias.n400 gnd 0.009349f
C1239 commonsourceibias.n401 gnd 0.009666f
C1240 commonsourceibias.n402 gnd 0.082208f
C1241 commonsourceibias.n403 gnd 0.05322f
C1242 commonsourceibias.n404 gnd 0.012299f
C1243 commonsourceibias.t91 gnd 0.172196f
C1244 commonsourceibias.n405 gnd 0.068706f
C1245 commonsourceibias.n406 gnd 0.009217f
C1246 commonsourceibias.t83 gnd 0.172196f
C1247 commonsourceibias.n407 gnd 0.007456f
C1248 commonsourceibias.n408 gnd 0.009217f
C1249 commonsourceibias.t73 gnd 0.172196f
C1250 commonsourceibias.n409 gnd 0.008898f
C1251 commonsourceibias.n410 gnd 0.009217f
C1252 commonsourceibias.t82 gnd 0.172196f
C1253 commonsourceibias.n411 gnd 0.007444f
C1254 commonsourceibias.n412 gnd 0.009217f
C1255 commonsourceibias.t103 gnd 0.172196f
C1256 commonsourceibias.t96 gnd 0.172196f
C1257 commonsourceibias.n413 gnd 0.068706f
C1258 commonsourceibias.n414 gnd 0.009217f
C1259 commonsourceibias.t81 gnd 0.172196f
C1260 commonsourceibias.n415 gnd 0.068706f
C1261 commonsourceibias.n416 gnd 0.009217f
C1262 commonsourceibias.t102 gnd 0.172196f
C1263 commonsourceibias.n417 gnd 0.068706f
C1264 commonsourceibias.n418 gnd 0.046399f
C1265 commonsourceibias.t116 gnd 0.172196f
C1266 commonsourceibias.t80 gnd 0.194303f
C1267 commonsourceibias.n419 gnd 0.079733f
C1268 commonsourceibias.n420 gnd 0.082545f
C1269 commonsourceibias.n421 gnd 0.01136f
C1270 commonsourceibias.n422 gnd 0.012567f
C1271 commonsourceibias.n423 gnd 0.009217f
C1272 commonsourceibias.n424 gnd 0.009217f
C1273 commonsourceibias.n425 gnd 0.012485f
C1274 commonsourceibias.n426 gnd 0.007456f
C1275 commonsourceibias.n427 gnd 0.01264f
C1276 commonsourceibias.n428 gnd 0.009217f
C1277 commonsourceibias.n429 gnd 0.009217f
C1278 commonsourceibias.n430 gnd 0.012717f
C1279 commonsourceibias.n431 gnd 0.010966f
C1280 commonsourceibias.n432 gnd 0.008898f
C1281 commonsourceibias.n433 gnd 0.009217f
C1282 commonsourceibias.n434 gnd 0.009217f
C1283 commonsourceibias.n435 gnd 0.011274f
C1284 commonsourceibias.n436 gnd 0.012653f
C1285 commonsourceibias.n437 gnd 0.068706f
C1286 commonsourceibias.n438 gnd 0.012568f
C1287 commonsourceibias.n439 gnd 0.009217f
C1288 commonsourceibias.n440 gnd 0.009217f
C1289 commonsourceibias.n441 gnd 0.009217f
C1290 commonsourceibias.n442 gnd 0.012568f
C1291 commonsourceibias.n443 gnd 0.068706f
C1292 commonsourceibias.n444 gnd 0.012653f
C1293 commonsourceibias.t90 gnd 0.172196f
C1294 commonsourceibias.n445 gnd 0.068706f
C1295 commonsourceibias.n446 gnd 0.011274f
C1296 commonsourceibias.n447 gnd 0.009217f
C1297 commonsourceibias.n448 gnd 0.009217f
C1298 commonsourceibias.n449 gnd 0.009217f
C1299 commonsourceibias.n450 gnd 0.010966f
C1300 commonsourceibias.n451 gnd 0.012717f
C1301 commonsourceibias.n452 gnd 0.068706f
C1302 commonsourceibias.n453 gnd 0.01264f
C1303 commonsourceibias.n454 gnd 0.009217f
C1304 commonsourceibias.n455 gnd 0.009217f
C1305 commonsourceibias.n456 gnd 0.009217f
C1306 commonsourceibias.n457 gnd 0.012485f
C1307 commonsourceibias.n458 gnd 0.068706f
C1308 commonsourceibias.n459 gnd 0.012567f
C1309 commonsourceibias.n460 gnd 0.01136f
C1310 commonsourceibias.n461 gnd 0.009217f
C1311 commonsourceibias.n462 gnd 0.009217f
C1312 commonsourceibias.n463 gnd 0.009349f
C1313 commonsourceibias.n464 gnd 0.009666f
C1314 commonsourceibias.t74 gnd 0.18623f
C1315 commonsourceibias.n465 gnd 0.082208f
C1316 commonsourceibias.n466 gnd 0.027976f
C1317 commonsourceibias.n467 gnd 0.147064f
C1318 commonsourceibias.n468 gnd 0.012299f
C1319 commonsourceibias.t62 gnd 0.172196f
C1320 commonsourceibias.n469 gnd 0.068706f
C1321 commonsourceibias.n470 gnd 0.009217f
C1322 commonsourceibias.t71 gnd 0.172196f
C1323 commonsourceibias.n471 gnd 0.007456f
C1324 commonsourceibias.n472 gnd 0.009217f
C1325 commonsourceibias.t48 gnd 0.172196f
C1326 commonsourceibias.n473 gnd 0.008898f
C1327 commonsourceibias.n474 gnd 0.009217f
C1328 commonsourceibias.t67 gnd 0.172196f
C1329 commonsourceibias.n475 gnd 0.007444f
C1330 commonsourceibias.n476 gnd 0.009217f
C1331 commonsourceibias.t77 gnd 0.172196f
C1332 commonsourceibias.t110 gnd 0.172196f
C1333 commonsourceibias.n477 gnd 0.068706f
C1334 commonsourceibias.n478 gnd 0.009217f
C1335 commonsourceibias.t61 gnd 0.172196f
C1336 commonsourceibias.n479 gnd 0.068706f
C1337 commonsourceibias.n480 gnd 0.009217f
C1338 commonsourceibias.t72 gnd 0.172196f
C1339 commonsourceibias.n481 gnd 0.068706f
C1340 commonsourceibias.n482 gnd 0.046399f
C1341 commonsourceibias.t68 gnd 0.172196f
C1342 commonsourceibias.t55 gnd 0.194303f
C1343 commonsourceibias.n483 gnd 0.079733f
C1344 commonsourceibias.n484 gnd 0.082545f
C1345 commonsourceibias.n485 gnd 0.01136f
C1346 commonsourceibias.n486 gnd 0.012567f
C1347 commonsourceibias.n487 gnd 0.009217f
C1348 commonsourceibias.n488 gnd 0.009217f
C1349 commonsourceibias.n489 gnd 0.012485f
C1350 commonsourceibias.n490 gnd 0.007456f
C1351 commonsourceibias.n491 gnd 0.01264f
C1352 commonsourceibias.n492 gnd 0.009217f
C1353 commonsourceibias.n493 gnd 0.009217f
C1354 commonsourceibias.n494 gnd 0.012717f
C1355 commonsourceibias.n495 gnd 0.010966f
C1356 commonsourceibias.n496 gnd 0.008898f
C1357 commonsourceibias.n497 gnd 0.009217f
C1358 commonsourceibias.n498 gnd 0.009217f
C1359 commonsourceibias.n499 gnd 0.011274f
C1360 commonsourceibias.n500 gnd 0.012653f
C1361 commonsourceibias.n501 gnd 0.068706f
C1362 commonsourceibias.n502 gnd 0.012568f
C1363 commonsourceibias.n503 gnd 0.009217f
C1364 commonsourceibias.n504 gnd 0.009217f
C1365 commonsourceibias.n505 gnd 0.009217f
C1366 commonsourceibias.n506 gnd 0.012568f
C1367 commonsourceibias.n507 gnd 0.068706f
C1368 commonsourceibias.n508 gnd 0.012653f
C1369 commonsourceibias.t57 gnd 0.172196f
C1370 commonsourceibias.n509 gnd 0.068706f
C1371 commonsourceibias.n510 gnd 0.011274f
C1372 commonsourceibias.n511 gnd 0.009217f
C1373 commonsourceibias.n512 gnd 0.009217f
C1374 commonsourceibias.n513 gnd 0.009217f
C1375 commonsourceibias.n514 gnd 0.010966f
C1376 commonsourceibias.n515 gnd 0.012717f
C1377 commonsourceibias.n516 gnd 0.068706f
C1378 commonsourceibias.n517 gnd 0.01264f
C1379 commonsourceibias.n518 gnd 0.009217f
C1380 commonsourceibias.n519 gnd 0.009217f
C1381 commonsourceibias.n520 gnd 0.009217f
C1382 commonsourceibias.n521 gnd 0.012485f
C1383 commonsourceibias.n522 gnd 0.068706f
C1384 commonsourceibias.n523 gnd 0.012567f
C1385 commonsourceibias.n524 gnd 0.01136f
C1386 commonsourceibias.n525 gnd 0.009217f
C1387 commonsourceibias.n526 gnd 0.009217f
C1388 commonsourceibias.n527 gnd 0.009349f
C1389 commonsourceibias.n528 gnd 0.009666f
C1390 commonsourceibias.t51 gnd 0.18623f
C1391 commonsourceibias.n529 gnd 0.082208f
C1392 commonsourceibias.n530 gnd 0.027976f
C1393 commonsourceibias.n531 gnd 0.194274f
C1394 commonsourceibias.n532 gnd 5.09694f
C1395 CSoutput.n0 gnd 0.041334f
C1396 CSoutput.t145 gnd 0.273414f
C1397 CSoutput.n1 gnd 0.12346f
C1398 CSoutput.n2 gnd 0.041334f
C1399 CSoutput.t148 gnd 0.273414f
C1400 CSoutput.n3 gnd 0.03276f
C1401 CSoutput.n4 gnd 0.041334f
C1402 CSoutput.t158 gnd 0.273414f
C1403 CSoutput.n5 gnd 0.02825f
C1404 CSoutput.n6 gnd 0.041334f
C1405 CSoutput.t147 gnd 0.273414f
C1406 CSoutput.t151 gnd 0.273414f
C1407 CSoutput.n7 gnd 0.122114f
C1408 CSoutput.n8 gnd 0.041334f
C1409 CSoutput.t157 gnd 0.273414f
C1410 CSoutput.n9 gnd 0.026934f
C1411 CSoutput.n10 gnd 0.041334f
C1412 CSoutput.t160 gnd 0.273414f
C1413 CSoutput.t149 gnd 0.273414f
C1414 CSoutput.n11 gnd 0.122114f
C1415 CSoutput.n12 gnd 0.041334f
C1416 CSoutput.t156 gnd 0.273414f
C1417 CSoutput.n13 gnd 0.02825f
C1418 CSoutput.n14 gnd 0.041334f
C1419 CSoutput.t153 gnd 0.273414f
C1420 CSoutput.t165 gnd 0.273414f
C1421 CSoutput.n15 gnd 0.122114f
C1422 CSoutput.n16 gnd 0.041334f
C1423 CSoutput.t152 gnd 0.273414f
C1424 CSoutput.n17 gnd 0.030172f
C1425 CSoutput.t161 gnd 0.326737f
C1426 CSoutput.t150 gnd 0.273414f
C1427 CSoutput.n18 gnd 0.155893f
C1428 CSoutput.n19 gnd 0.15127f
C1429 CSoutput.n20 gnd 0.175491f
C1430 CSoutput.n21 gnd 0.041334f
C1431 CSoutput.n22 gnd 0.034498f
C1432 CSoutput.n23 gnd 0.122114f
C1433 CSoutput.n24 gnd 0.033255f
C1434 CSoutput.n25 gnd 0.03276f
C1435 CSoutput.n26 gnd 0.041334f
C1436 CSoutput.n27 gnd 0.041334f
C1437 CSoutput.n28 gnd 0.034232f
C1438 CSoutput.n29 gnd 0.029064f
C1439 CSoutput.n30 gnd 0.124833f
C1440 CSoutput.n31 gnd 0.029465f
C1441 CSoutput.n32 gnd 0.041334f
C1442 CSoutput.n33 gnd 0.041334f
C1443 CSoutput.n34 gnd 0.041334f
C1444 CSoutput.n35 gnd 0.033868f
C1445 CSoutput.n36 gnd 0.122114f
C1446 CSoutput.n37 gnd 0.03239f
C1447 CSoutput.n38 gnd 0.033625f
C1448 CSoutput.n39 gnd 0.041334f
C1449 CSoutput.n40 gnd 0.041334f
C1450 CSoutput.n41 gnd 0.03449f
C1451 CSoutput.n42 gnd 0.031524f
C1452 CSoutput.n43 gnd 0.122114f
C1453 CSoutput.n44 gnd 0.032324f
C1454 CSoutput.n45 gnd 0.041334f
C1455 CSoutput.n46 gnd 0.041334f
C1456 CSoutput.n47 gnd 0.041334f
C1457 CSoutput.n48 gnd 0.032324f
C1458 CSoutput.n49 gnd 0.122114f
C1459 CSoutput.n50 gnd 0.031524f
C1460 CSoutput.n51 gnd 0.03449f
C1461 CSoutput.n52 gnd 0.041334f
C1462 CSoutput.n53 gnd 0.041334f
C1463 CSoutput.n54 gnd 0.033625f
C1464 CSoutput.n55 gnd 0.03239f
C1465 CSoutput.n56 gnd 0.122114f
C1466 CSoutput.n57 gnd 0.033868f
C1467 CSoutput.n58 gnd 0.041334f
C1468 CSoutput.n59 gnd 0.041334f
C1469 CSoutput.n60 gnd 0.041334f
C1470 CSoutput.n61 gnd 0.029465f
C1471 CSoutput.n62 gnd 0.124833f
C1472 CSoutput.n63 gnd 0.029064f
C1473 CSoutput.t159 gnd 0.273414f
C1474 CSoutput.n64 gnd 0.122114f
C1475 CSoutput.n65 gnd 0.034232f
C1476 CSoutput.n66 gnd 0.041334f
C1477 CSoutput.n67 gnd 0.041334f
C1478 CSoutput.n68 gnd 0.041334f
C1479 CSoutput.n69 gnd 0.033255f
C1480 CSoutput.n70 gnd 0.122114f
C1481 CSoutput.n71 gnd 0.034498f
C1482 CSoutput.n72 gnd 0.030172f
C1483 CSoutput.n73 gnd 0.041334f
C1484 CSoutput.n74 gnd 0.041334f
C1485 CSoutput.n75 gnd 0.03129f
C1486 CSoutput.n76 gnd 0.018583f
C1487 CSoutput.t164 gnd 0.3072f
C1488 CSoutput.n77 gnd 0.152605f
C1489 CSoutput.n78 gnd 0.624298f
C1490 CSoutput.t18 gnd 0.051558f
C1491 CSoutput.t55 gnd 0.051558f
C1492 CSoutput.n79 gnd 0.39918f
C1493 CSoutput.t21 gnd 0.051558f
C1494 CSoutput.t41 gnd 0.051558f
C1495 CSoutput.n80 gnd 0.398468f
C1496 CSoutput.n81 gnd 0.404444f
C1497 CSoutput.t84 gnd 0.051558f
C1498 CSoutput.t50 gnd 0.051558f
C1499 CSoutput.n82 gnd 0.398468f
C1500 CSoutput.n83 gnd 0.199293f
C1501 CSoutput.t23 gnd 0.051558f
C1502 CSoutput.t73 gnd 0.051558f
C1503 CSoutput.n84 gnd 0.398468f
C1504 CSoutput.n85 gnd 0.199293f
C1505 CSoutput.t30 gnd 0.051558f
C1506 CSoutput.t62 gnd 0.051558f
C1507 CSoutput.n86 gnd 0.398468f
C1508 CSoutput.n87 gnd 0.199293f
C1509 CSoutput.t44 gnd 0.051558f
C1510 CSoutput.t56 gnd 0.051558f
C1511 CSoutput.n88 gnd 0.398468f
C1512 CSoutput.n89 gnd 0.365458f
C1513 CSoutput.t34 gnd 0.051558f
C1514 CSoutput.t79 gnd 0.051558f
C1515 CSoutput.n90 gnd 0.39918f
C1516 CSoutput.t64 gnd 0.051558f
C1517 CSoutput.t61 gnd 0.051558f
C1518 CSoutput.n91 gnd 0.398468f
C1519 CSoutput.n92 gnd 0.404444f
C1520 CSoutput.t54 gnd 0.051558f
C1521 CSoutput.t32 gnd 0.051558f
C1522 CSoutput.n93 gnd 0.398468f
C1523 CSoutput.n94 gnd 0.199293f
C1524 CSoutput.t17 gnd 0.051558f
C1525 CSoutput.t53 gnd 0.051558f
C1526 CSoutput.n95 gnd 0.398468f
C1527 CSoutput.n96 gnd 0.199293f
C1528 CSoutput.t52 gnd 0.051558f
C1529 CSoutput.t31 gnd 0.051558f
C1530 CSoutput.n97 gnd 0.398468f
C1531 CSoutput.n98 gnd 0.199293f
C1532 CSoutput.t14 gnd 0.051558f
C1533 CSoutput.t15 gnd 0.051558f
C1534 CSoutput.n99 gnd 0.398468f
C1535 CSoutput.n100 gnd 0.297196f
C1536 CSoutput.n101 gnd 0.374762f
C1537 CSoutput.t45 gnd 0.051558f
C1538 CSoutput.t85 gnd 0.051558f
C1539 CSoutput.n102 gnd 0.39918f
C1540 CSoutput.t67 gnd 0.051558f
C1541 CSoutput.t68 gnd 0.051558f
C1542 CSoutput.n103 gnd 0.398468f
C1543 CSoutput.n104 gnd 0.404444f
C1544 CSoutput.t59 gnd 0.051558f
C1545 CSoutput.t43 gnd 0.051558f
C1546 CSoutput.n105 gnd 0.398468f
C1547 CSoutput.n106 gnd 0.199293f
C1548 CSoutput.t27 gnd 0.051558f
C1549 CSoutput.t60 gnd 0.051558f
C1550 CSoutput.n107 gnd 0.398468f
C1551 CSoutput.n108 gnd 0.199293f
C1552 CSoutput.t58 gnd 0.051558f
C1553 CSoutput.t40 gnd 0.051558f
C1554 CSoutput.n109 gnd 0.398468f
C1555 CSoutput.n110 gnd 0.199293f
C1556 CSoutput.t26 gnd 0.051558f
C1557 CSoutput.t25 gnd 0.051558f
C1558 CSoutput.n111 gnd 0.398468f
C1559 CSoutput.n112 gnd 0.297196f
C1560 CSoutput.n113 gnd 0.418889f
C1561 CSoutput.n114 gnd 7.67994f
C1562 CSoutput.n116 gnd 0.731187f
C1563 CSoutput.n117 gnd 0.54839f
C1564 CSoutput.n118 gnd 0.731187f
C1565 CSoutput.n119 gnd 0.731187f
C1566 CSoutput.n120 gnd 1.96858f
C1567 CSoutput.n121 gnd 0.731187f
C1568 CSoutput.n122 gnd 0.731187f
C1569 CSoutput.t154 gnd 0.913984f
C1570 CSoutput.n123 gnd 0.731187f
C1571 CSoutput.n124 gnd 0.731187f
C1572 CSoutput.n128 gnd 0.731187f
C1573 CSoutput.n132 gnd 0.731187f
C1574 CSoutput.n133 gnd 0.731187f
C1575 CSoutput.n135 gnd 0.731187f
C1576 CSoutput.n140 gnd 0.731187f
C1577 CSoutput.n142 gnd 0.731187f
C1578 CSoutput.n143 gnd 0.731187f
C1579 CSoutput.n145 gnd 0.731187f
C1580 CSoutput.n146 gnd 0.731187f
C1581 CSoutput.n148 gnd 0.731187f
C1582 CSoutput.t144 gnd 12.2181f
C1583 CSoutput.n150 gnd 0.731187f
C1584 CSoutput.n151 gnd 0.54839f
C1585 CSoutput.n152 gnd 0.731187f
C1586 CSoutput.n153 gnd 0.731187f
C1587 CSoutput.n154 gnd 1.96858f
C1588 CSoutput.n155 gnd 0.731187f
C1589 CSoutput.n156 gnd 0.731187f
C1590 CSoutput.t162 gnd 0.913984f
C1591 CSoutput.n157 gnd 0.731187f
C1592 CSoutput.n158 gnd 0.731187f
C1593 CSoutput.n162 gnd 0.731187f
C1594 CSoutput.n166 gnd 0.731187f
C1595 CSoutput.n167 gnd 0.731187f
C1596 CSoutput.n169 gnd 0.731187f
C1597 CSoutput.n174 gnd 0.731187f
C1598 CSoutput.n176 gnd 0.731187f
C1599 CSoutput.n177 gnd 0.731187f
C1600 CSoutput.n179 gnd 0.731187f
C1601 CSoutput.n180 gnd 0.731187f
C1602 CSoutput.n182 gnd 0.731187f
C1603 CSoutput.n183 gnd 0.54839f
C1604 CSoutput.n185 gnd 0.731187f
C1605 CSoutput.n186 gnd 0.54839f
C1606 CSoutput.n187 gnd 0.731187f
C1607 CSoutput.n188 gnd 0.731187f
C1608 CSoutput.n189 gnd 1.96858f
C1609 CSoutput.n190 gnd 0.731187f
C1610 CSoutput.n191 gnd 0.731187f
C1611 CSoutput.t155 gnd 0.913984f
C1612 CSoutput.n192 gnd 0.731187f
C1613 CSoutput.n193 gnd 1.96858f
C1614 CSoutput.n195 gnd 0.731187f
C1615 CSoutput.n196 gnd 0.731187f
C1616 CSoutput.n198 gnd 0.731187f
C1617 CSoutput.n199 gnd 0.731187f
C1618 CSoutput.t163 gnd 12.0189f
C1619 CSoutput.t146 gnd 12.2181f
C1620 CSoutput.n205 gnd 2.29384f
C1621 CSoutput.n206 gnd 9.344269f
C1622 CSoutput.n207 gnd 9.73528f
C1623 CSoutput.n212 gnd 2.48485f
C1624 CSoutput.n218 gnd 0.731187f
C1625 CSoutput.n220 gnd 0.731187f
C1626 CSoutput.n222 gnd 0.731187f
C1627 CSoutput.n224 gnd 0.731187f
C1628 CSoutput.n226 gnd 0.731187f
C1629 CSoutput.n232 gnd 0.731187f
C1630 CSoutput.n239 gnd 1.34145f
C1631 CSoutput.n240 gnd 1.34145f
C1632 CSoutput.n241 gnd 0.731187f
C1633 CSoutput.n242 gnd 0.731187f
C1634 CSoutput.n244 gnd 0.54839f
C1635 CSoutput.n245 gnd 0.469647f
C1636 CSoutput.n247 gnd 0.54839f
C1637 CSoutput.n248 gnd 0.469647f
C1638 CSoutput.n249 gnd 0.54839f
C1639 CSoutput.n251 gnd 0.731187f
C1640 CSoutput.n253 gnd 1.96858f
C1641 CSoutput.n254 gnd 2.29384f
C1642 CSoutput.n255 gnd 8.59433f
C1643 CSoutput.n257 gnd 0.54839f
C1644 CSoutput.n258 gnd 1.41104f
C1645 CSoutput.n259 gnd 0.54839f
C1646 CSoutput.n261 gnd 0.731187f
C1647 CSoutput.n263 gnd 1.96858f
C1648 CSoutput.n264 gnd 4.28789f
C1649 CSoutput.t69 gnd 0.051558f
C1650 CSoutput.t16 gnd 0.051558f
C1651 CSoutput.n265 gnd 0.39918f
C1652 CSoutput.t39 gnd 0.051558f
C1653 CSoutput.t22 gnd 0.051558f
C1654 CSoutput.n266 gnd 0.398468f
C1655 CSoutput.n267 gnd 0.404444f
C1656 CSoutput.t51 gnd 0.051558f
C1657 CSoutput.t36 gnd 0.051558f
C1658 CSoutput.n268 gnd 0.398468f
C1659 CSoutput.n269 gnd 0.199293f
C1660 CSoutput.t74 gnd 0.051558f
C1661 CSoutput.t24 gnd 0.051558f
C1662 CSoutput.n270 gnd 0.398468f
C1663 CSoutput.n271 gnd 0.199293f
C1664 CSoutput.t63 gnd 0.051558f
C1665 CSoutput.t28 gnd 0.051558f
C1666 CSoutput.n272 gnd 0.398468f
C1667 CSoutput.n273 gnd 0.199293f
C1668 CSoutput.t70 gnd 0.051558f
C1669 CSoutput.t42 gnd 0.051558f
C1670 CSoutput.n274 gnd 0.398468f
C1671 CSoutput.n275 gnd 0.365458f
C1672 CSoutput.t38 gnd 0.051558f
C1673 CSoutput.t78 gnd 0.051558f
C1674 CSoutput.n276 gnd 0.39918f
C1675 CSoutput.t35 gnd 0.051558f
C1676 CSoutput.t37 gnd 0.051558f
C1677 CSoutput.n277 gnd 0.398468f
C1678 CSoutput.n278 gnd 0.404444f
C1679 CSoutput.t76 gnd 0.051558f
C1680 CSoutput.t77 gnd 0.051558f
C1681 CSoutput.n279 gnd 0.398468f
C1682 CSoutput.n280 gnd 0.199293f
C1683 CSoutput.t20 gnd 0.051558f
C1684 CSoutput.t66 gnd 0.051558f
C1685 CSoutput.n281 gnd 0.398468f
C1686 CSoutput.n282 gnd 0.199293f
C1687 CSoutput.t75 gnd 0.051558f
C1688 CSoutput.t19 gnd 0.051558f
C1689 CSoutput.n283 gnd 0.398468f
C1690 CSoutput.n284 gnd 0.199293f
C1691 CSoutput.t49 gnd 0.051558f
C1692 CSoutput.t65 gnd 0.051558f
C1693 CSoutput.n285 gnd 0.398468f
C1694 CSoutput.n286 gnd 0.297196f
C1695 CSoutput.n287 gnd 0.374762f
C1696 CSoutput.t48 gnd 0.051558f
C1697 CSoutput.t83 gnd 0.051558f
C1698 CSoutput.n288 gnd 0.39918f
C1699 CSoutput.t46 gnd 0.051558f
C1700 CSoutput.t47 gnd 0.051558f
C1701 CSoutput.n289 gnd 0.398468f
C1702 CSoutput.n290 gnd 0.404444f
C1703 CSoutput.t81 gnd 0.051558f
C1704 CSoutput.t82 gnd 0.051558f
C1705 CSoutput.n291 gnd 0.398468f
C1706 CSoutput.n292 gnd 0.199293f
C1707 CSoutput.t33 gnd 0.051558f
C1708 CSoutput.t72 gnd 0.051558f
C1709 CSoutput.n293 gnd 0.398468f
C1710 CSoutput.n294 gnd 0.199293f
C1711 CSoutput.t80 gnd 0.051558f
C1712 CSoutput.t29 gnd 0.051558f
C1713 CSoutput.n295 gnd 0.398468f
C1714 CSoutput.n296 gnd 0.199293f
C1715 CSoutput.t57 gnd 0.051558f
C1716 CSoutput.t71 gnd 0.051558f
C1717 CSoutput.n297 gnd 0.398466f
C1718 CSoutput.n298 gnd 0.297198f
C1719 CSoutput.n299 gnd 0.418889f
C1720 CSoutput.n300 gnd 11.0052f
C1721 CSoutput.t104 gnd 0.045113f
C1722 CSoutput.t114 gnd 0.045113f
C1723 CSoutput.n301 gnd 0.399971f
C1724 CSoutput.t110 gnd 0.045113f
C1725 CSoutput.t119 gnd 0.045113f
C1726 CSoutput.n302 gnd 0.398637f
C1727 CSoutput.n303 gnd 0.371455f
C1728 CSoutput.t6 gnd 0.045113f
C1729 CSoutput.t90 gnd 0.045113f
C1730 CSoutput.n304 gnd 0.398637f
C1731 CSoutput.n305 gnd 0.18311f
C1732 CSoutput.t140 gnd 0.045113f
C1733 CSoutput.t0 gnd 0.045113f
C1734 CSoutput.n306 gnd 0.398637f
C1735 CSoutput.n307 gnd 0.18311f
C1736 CSoutput.t10 gnd 0.045113f
C1737 CSoutput.t111 gnd 0.045113f
C1738 CSoutput.n308 gnd 0.398637f
C1739 CSoutput.n309 gnd 0.18311f
C1740 CSoutput.t135 gnd 0.045113f
C1741 CSoutput.t143 gnd 0.045113f
C1742 CSoutput.n310 gnd 0.398637f
C1743 CSoutput.n311 gnd 0.337736f
C1744 CSoutput.t94 gnd 0.045113f
C1745 CSoutput.t88 gnd 0.045113f
C1746 CSoutput.n312 gnd 0.399971f
C1747 CSoutput.t97 gnd 0.045113f
C1748 CSoutput.t96 gnd 0.045113f
C1749 CSoutput.n313 gnd 0.398637f
C1750 CSoutput.n314 gnd 0.371455f
C1751 CSoutput.t124 gnd 0.045113f
C1752 CSoutput.t127 gnd 0.045113f
C1753 CSoutput.n315 gnd 0.398637f
C1754 CSoutput.n316 gnd 0.18311f
C1755 CSoutput.t115 gnd 0.045113f
C1756 CSoutput.t3 gnd 0.045113f
C1757 CSoutput.n317 gnd 0.398637f
C1758 CSoutput.n318 gnd 0.18311f
C1759 CSoutput.t107 gnd 0.045113f
C1760 CSoutput.t100 gnd 0.045113f
C1761 CSoutput.n319 gnd 0.398637f
C1762 CSoutput.n320 gnd 0.18311f
C1763 CSoutput.t95 gnd 0.045113f
C1764 CSoutput.t105 gnd 0.045113f
C1765 CSoutput.n321 gnd 0.398637f
C1766 CSoutput.n322 gnd 0.278f
C1767 CSoutput.n323 gnd 0.350645f
C1768 CSoutput.t92 gnd 0.045113f
C1769 CSoutput.t117 gnd 0.045113f
C1770 CSoutput.n324 gnd 0.399971f
C1771 CSoutput.t99 gnd 0.045113f
C1772 CSoutput.t89 gnd 0.045113f
C1773 CSoutput.n325 gnd 0.398637f
C1774 CSoutput.n326 gnd 0.371455f
C1775 CSoutput.t8 gnd 0.045113f
C1776 CSoutput.t120 gnd 0.045113f
C1777 CSoutput.n327 gnd 0.398637f
C1778 CSoutput.n328 gnd 0.18311f
C1779 CSoutput.t129 gnd 0.045113f
C1780 CSoutput.t130 gnd 0.045113f
C1781 CSoutput.n329 gnd 0.398637f
C1782 CSoutput.n330 gnd 0.18311f
C1783 CSoutput.t102 gnd 0.045113f
C1784 CSoutput.t137 gnd 0.045113f
C1785 CSoutput.n331 gnd 0.398637f
C1786 CSoutput.n332 gnd 0.18311f
C1787 CSoutput.t118 gnd 0.045113f
C1788 CSoutput.t132 gnd 0.045113f
C1789 CSoutput.n333 gnd 0.398637f
C1790 CSoutput.n334 gnd 0.278f
C1791 CSoutput.n335 gnd 0.376537f
C1792 CSoutput.n336 gnd 11.272f
C1793 CSoutput.t112 gnd 0.045113f
C1794 CSoutput.t9 gnd 0.045113f
C1795 CSoutput.n337 gnd 0.399971f
C1796 CSoutput.t11 gnd 0.045113f
C1797 CSoutput.t125 gnd 0.045113f
C1798 CSoutput.n338 gnd 0.398637f
C1799 CSoutput.n339 gnd 0.371455f
C1800 CSoutput.t13 gnd 0.045113f
C1801 CSoutput.t98 gnd 0.045113f
C1802 CSoutput.n340 gnd 0.398637f
C1803 CSoutput.n341 gnd 0.18311f
C1804 CSoutput.t141 gnd 0.045113f
C1805 CSoutput.t136 gnd 0.045113f
C1806 CSoutput.n342 gnd 0.398637f
C1807 CSoutput.n343 gnd 0.18311f
C1808 CSoutput.t121 gnd 0.045113f
C1809 CSoutput.t123 gnd 0.045113f
C1810 CSoutput.n344 gnd 0.398637f
C1811 CSoutput.n345 gnd 0.18311f
C1812 CSoutput.t113 gnd 0.045113f
C1813 CSoutput.t133 gnd 0.045113f
C1814 CSoutput.n346 gnd 0.398637f
C1815 CSoutput.n347 gnd 0.337736f
C1816 CSoutput.t7 gnd 0.045113f
C1817 CSoutput.t128 gnd 0.045113f
C1818 CSoutput.n348 gnd 0.399971f
C1819 CSoutput.t138 gnd 0.045113f
C1820 CSoutput.t2 gnd 0.045113f
C1821 CSoutput.n349 gnd 0.398637f
C1822 CSoutput.n350 gnd 0.371455f
C1823 CSoutput.t1 gnd 0.045113f
C1824 CSoutput.t122 gnd 0.045113f
C1825 CSoutput.n351 gnd 0.398637f
C1826 CSoutput.n352 gnd 0.18311f
C1827 CSoutput.t5 gnd 0.045113f
C1828 CSoutput.t93 gnd 0.045113f
C1829 CSoutput.n353 gnd 0.398637f
C1830 CSoutput.n354 gnd 0.18311f
C1831 CSoutput.t103 gnd 0.045113f
C1832 CSoutput.t126 gnd 0.045113f
C1833 CSoutput.n355 gnd 0.398637f
C1834 CSoutput.n356 gnd 0.18311f
C1835 CSoutput.t4 gnd 0.045113f
C1836 CSoutput.t12 gnd 0.045113f
C1837 CSoutput.n357 gnd 0.398637f
C1838 CSoutput.n358 gnd 0.278f
C1839 CSoutput.n359 gnd 0.350645f
C1840 CSoutput.t86 gnd 0.045113f
C1841 CSoutput.t87 gnd 0.045113f
C1842 CSoutput.n360 gnd 0.399971f
C1843 CSoutput.t131 gnd 0.045113f
C1844 CSoutput.t142 gnd 0.045113f
C1845 CSoutput.n361 gnd 0.398637f
C1846 CSoutput.n362 gnd 0.371455f
C1847 CSoutput.t109 gnd 0.045113f
C1848 CSoutput.t106 gnd 0.045113f
C1849 CSoutput.n363 gnd 0.398637f
C1850 CSoutput.n364 gnd 0.18311f
C1851 CSoutput.t134 gnd 0.045113f
C1852 CSoutput.t116 gnd 0.045113f
C1853 CSoutput.n365 gnd 0.398637f
C1854 CSoutput.n366 gnd 0.18311f
C1855 CSoutput.t101 gnd 0.045113f
C1856 CSoutput.t139 gnd 0.045113f
C1857 CSoutput.n367 gnd 0.398637f
C1858 CSoutput.n368 gnd 0.18311f
C1859 CSoutput.t91 gnd 0.045113f
C1860 CSoutput.t108 gnd 0.045113f
C1861 CSoutput.n369 gnd 0.398637f
C1862 CSoutput.n370 gnd 0.278f
C1863 CSoutput.n371 gnd 0.376537f
C1864 CSoutput.n372 gnd 6.48744f
C1865 CSoutput.n373 gnd 12.5312f
C1866 a_n7636_8799.n0 gnd 2.71476f
C1867 a_n7636_8799.n1 gnd 1.6448f
C1868 a_n7636_8799.n2 gnd 3.76313f
C1869 a_n7636_8799.n3 gnd 0.17526f
C1870 a_n7636_8799.n4 gnd 0.205241f
C1871 a_n7636_8799.n5 gnd 0.205241f
C1872 a_n7636_8799.n6 gnd 0.205241f
C1873 a_n7636_8799.n7 gnd 0.17526f
C1874 a_n7636_8799.n8 gnd 0.205241f
C1875 a_n7636_8799.n9 gnd 0.205241f
C1876 a_n7636_8799.n10 gnd 0.205241f
C1877 a_n7636_8799.n11 gnd 0.338541f
C1878 a_n7636_8799.n12 gnd 0.205241f
C1879 a_n7636_8799.n13 gnd 0.205241f
C1880 a_n7636_8799.n14 gnd 0.205241f
C1881 a_n7636_8799.n15 gnd 0.205241f
C1882 a_n7636_8799.n16 gnd 0.205241f
C1883 a_n7636_8799.n17 gnd 0.17526f
C1884 a_n7636_8799.n18 gnd 0.205241f
C1885 a_n7636_8799.n19 gnd 0.205241f
C1886 a_n7636_8799.n20 gnd 0.205241f
C1887 a_n7636_8799.n21 gnd 0.17526f
C1888 a_n7636_8799.n22 gnd 0.205241f
C1889 a_n7636_8799.n23 gnd 0.205241f
C1890 a_n7636_8799.n24 gnd 0.205241f
C1891 a_n7636_8799.n25 gnd 0.338541f
C1892 a_n7636_8799.n26 gnd 0.205241f
C1893 a_n7636_8799.n27 gnd 1.50425f
C1894 a_n7636_8799.n28 gnd 2.74588f
C1895 a_n7636_8799.n29 gnd 3.88534f
C1896 a_n7636_8799.n30 gnd 1.50425f
C1897 a_n7636_8799.n31 gnd 0.248204f
C1898 a_n7636_8799.n33 gnd 0.007645f
C1899 a_n7636_8799.n34 gnd 0.011555f
C1900 a_n7636_8799.n35 gnd 0.007946f
C1901 a_n7636_8799.n37 gnd 3.97e-19
C1902 a_n7636_8799.n38 gnd 0.008235f
C1903 a_n7636_8799.n39 gnd 0.259651f
C1904 a_n7636_8799.n40 gnd 0.248204f
C1905 a_n7636_8799.n42 gnd 0.007645f
C1906 a_n7636_8799.n43 gnd 0.011555f
C1907 a_n7636_8799.n44 gnd 0.007946f
C1908 a_n7636_8799.n46 gnd 3.97e-19
C1909 a_n7636_8799.n47 gnd 0.008235f
C1910 a_n7636_8799.n48 gnd 0.259651f
C1911 a_n7636_8799.n49 gnd 0.248204f
C1912 a_n7636_8799.n51 gnd 0.007645f
C1913 a_n7636_8799.n52 gnd 0.011555f
C1914 a_n7636_8799.n53 gnd 0.007946f
C1915 a_n7636_8799.n55 gnd 3.97e-19
C1916 a_n7636_8799.n56 gnd 0.008235f
C1917 a_n7636_8799.n57 gnd 0.259651f
C1918 a_n7636_8799.n58 gnd 0.008235f
C1919 a_n7636_8799.n59 gnd 0.259651f
C1920 a_n7636_8799.n60 gnd 3.97e-19
C1921 a_n7636_8799.n62 gnd 0.007946f
C1922 a_n7636_8799.n63 gnd 0.011555f
C1923 a_n7636_8799.n64 gnd 0.007645f
C1924 a_n7636_8799.n66 gnd 0.248204f
C1925 a_n7636_8799.n67 gnd 0.008235f
C1926 a_n7636_8799.n68 gnd 0.259651f
C1927 a_n7636_8799.n69 gnd 3.97e-19
C1928 a_n7636_8799.n71 gnd 0.007946f
C1929 a_n7636_8799.n72 gnd 0.011555f
C1930 a_n7636_8799.n73 gnd 0.007645f
C1931 a_n7636_8799.n75 gnd 0.248204f
C1932 a_n7636_8799.n76 gnd 0.008235f
C1933 a_n7636_8799.n77 gnd 0.259651f
C1934 a_n7636_8799.n78 gnd 3.97e-19
C1935 a_n7636_8799.n80 gnd 0.007946f
C1936 a_n7636_8799.n81 gnd 0.011555f
C1937 a_n7636_8799.n82 gnd 0.007645f
C1938 a_n7636_8799.n84 gnd 0.248204f
C1939 a_n7636_8799.t32 gnd 0.142357f
C1940 a_n7636_8799.t31 gnd 0.142357f
C1941 a_n7636_8799.t19 gnd 0.142357f
C1942 a_n7636_8799.n85 gnd 1.12279f
C1943 a_n7636_8799.t27 gnd 0.142357f
C1944 a_n7636_8799.t15 gnd 0.142357f
C1945 a_n7636_8799.n86 gnd 1.12094f
C1946 a_n7636_8799.t23 gnd 0.142357f
C1947 a_n7636_8799.t28 gnd 0.142357f
C1948 a_n7636_8799.n87 gnd 1.12094f
C1949 a_n7636_8799.t17 gnd 0.142357f
C1950 a_n7636_8799.t20 gnd 0.142357f
C1951 a_n7636_8799.n88 gnd 1.12094f
C1952 a_n7636_8799.t25 gnd 0.142357f
C1953 a_n7636_8799.t24 gnd 0.142357f
C1954 a_n7636_8799.n89 gnd 1.12094f
C1955 a_n7636_8799.t0 gnd 0.110722f
C1956 a_n7636_8799.t35 gnd 0.110722f
C1957 a_n7636_8799.n90 gnd 0.981266f
C1958 a_n7636_8799.t10 gnd 0.110722f
C1959 a_n7636_8799.t2 gnd 0.110722f
C1960 a_n7636_8799.n91 gnd 0.978381f
C1961 a_n7636_8799.t1 gnd 0.110722f
C1962 a_n7636_8799.t8 gnd 0.110722f
C1963 a_n7636_8799.n92 gnd 0.981265f
C1964 a_n7636_8799.t3 gnd 0.110722f
C1965 a_n7636_8799.t4 gnd 0.110722f
C1966 a_n7636_8799.n93 gnd 0.97838f
C1967 a_n7636_8799.t34 gnd 0.110722f
C1968 a_n7636_8799.t12 gnd 0.110722f
C1969 a_n7636_8799.n94 gnd 0.981265f
C1970 a_n7636_8799.t11 gnd 0.110722f
C1971 a_n7636_8799.t13 gnd 0.110722f
C1972 a_n7636_8799.n95 gnd 0.97838f
C1973 a_n7636_8799.t7 gnd 0.110722f
C1974 a_n7636_8799.t9 gnd 0.110722f
C1975 a_n7636_8799.n96 gnd 0.978381f
C1976 a_n7636_8799.t6 gnd 0.110722f
C1977 a_n7636_8799.t5 gnd 0.110722f
C1978 a_n7636_8799.n97 gnd 0.978381f
C1979 a_n7636_8799.t53 gnd 0.590279f
C1980 a_n7636_8799.n98 gnd 0.267154f
C1981 a_n7636_8799.t76 gnd 0.590279f
C1982 a_n7636_8799.t78 gnd 0.590279f
C1983 a_n7636_8799.n99 gnd 0.25841f
C1984 a_n7636_8799.t94 gnd 0.590279f
C1985 a_n7636_8799.n100 gnd 0.269657f
C1986 a_n7636_8799.t61 gnd 0.590279f
C1987 a_n7636_8799.t63 gnd 0.590279f
C1988 a_n7636_8799.n101 gnd 0.263156f
C1989 a_n7636_8799.t95 gnd 0.604153f
C1990 a_n7636_8799.t96 gnd 0.590279f
C1991 a_n7636_8799.n102 gnd 0.269227f
C1992 a_n7636_8799.n103 gnd 0.24606f
C1993 a_n7636_8799.t81 gnd 0.590279f
C1994 a_n7636_8799.n104 gnd 0.267038f
C1995 a_n7636_8799.n105 gnd 0.267169f
C1996 a_n7636_8799.t62 gnd 0.590279f
C1997 a_n7636_8799.n106 gnd 0.263472f
C1998 a_n7636_8799.t54 gnd 0.590279f
C1999 a_n7636_8799.n107 gnd 0.263719f
C2000 a_n7636_8799.n108 gnd 0.269227f
C2001 a_n7636_8799.t36 gnd 0.600996f
C2002 a_n7636_8799.t60 gnd 0.590279f
C2003 a_n7636_8799.n109 gnd 0.267154f
C2004 a_n7636_8799.t87 gnd 0.590279f
C2005 a_n7636_8799.t89 gnd 0.590279f
C2006 a_n7636_8799.n110 gnd 0.25841f
C2007 a_n7636_8799.t104 gnd 0.590279f
C2008 a_n7636_8799.n111 gnd 0.269657f
C2009 a_n7636_8799.t68 gnd 0.590279f
C2010 a_n7636_8799.t69 gnd 0.590279f
C2011 a_n7636_8799.n112 gnd 0.263156f
C2012 a_n7636_8799.t107 gnd 0.604153f
C2013 a_n7636_8799.t106 gnd 0.590279f
C2014 a_n7636_8799.n113 gnd 0.269227f
C2015 a_n7636_8799.n114 gnd 0.24606f
C2016 a_n7636_8799.t90 gnd 0.590279f
C2017 a_n7636_8799.n115 gnd 0.267038f
C2018 a_n7636_8799.n116 gnd 0.267169f
C2019 a_n7636_8799.t67 gnd 0.590279f
C2020 a_n7636_8799.n117 gnd 0.263472f
C2021 a_n7636_8799.t57 gnd 0.590279f
C2022 a_n7636_8799.n118 gnd 0.263719f
C2023 a_n7636_8799.n119 gnd 0.269227f
C2024 a_n7636_8799.t42 gnd 0.600996f
C2025 a_n7636_8799.n120 gnd 0.886171f
C2026 a_n7636_8799.t80 gnd 0.590279f
C2027 a_n7636_8799.n121 gnd 0.267154f
C2028 a_n7636_8799.t103 gnd 0.590279f
C2029 a_n7636_8799.t71 gnd 0.590279f
C2030 a_n7636_8799.n122 gnd 0.25841f
C2031 a_n7636_8799.t98 gnd 0.590279f
C2032 a_n7636_8799.n123 gnd 0.269657f
C2033 a_n7636_8799.t48 gnd 0.590279f
C2034 a_n7636_8799.t91 gnd 0.590279f
C2035 a_n7636_8799.n124 gnd 0.263156f
C2036 a_n7636_8799.t77 gnd 0.604153f
C2037 a_n7636_8799.t65 gnd 0.590279f
C2038 a_n7636_8799.n125 gnd 0.269227f
C2039 a_n7636_8799.n126 gnd 0.24606f
C2040 a_n7636_8799.t59 gnd 0.590279f
C2041 a_n7636_8799.n127 gnd 0.267038f
C2042 a_n7636_8799.n128 gnd 0.267169f
C2043 a_n7636_8799.t37 gnd 0.590279f
C2044 a_n7636_8799.n129 gnd 0.263472f
C2045 a_n7636_8799.t100 gnd 0.590279f
C2046 a_n7636_8799.n130 gnd 0.263719f
C2047 a_n7636_8799.n131 gnd 0.269227f
C2048 a_n7636_8799.t66 gnd 0.600996f
C2049 a_n7636_8799.n132 gnd 1.68026f
C2050 a_n7636_8799.t73 gnd 0.600996f
C2051 a_n7636_8799.t38 gnd 0.590279f
C2052 a_n7636_8799.t75 gnd 0.590279f
C2053 a_n7636_8799.t74 gnd 0.590279f
C2054 a_n7636_8799.n133 gnd 0.263719f
C2055 a_n7636_8799.t40 gnd 0.590279f
C2056 a_n7636_8799.t39 gnd 0.590279f
C2057 a_n7636_8799.t88 gnd 0.590279f
C2058 a_n7636_8799.n134 gnd 0.267169f
C2059 a_n7636_8799.t49 gnd 0.590279f
C2060 a_n7636_8799.t41 gnd 0.590279f
C2061 a_n7636_8799.t92 gnd 0.590279f
C2062 a_n7636_8799.n135 gnd 0.263156f
C2063 a_n7636_8799.t50 gnd 0.604153f
C2064 a_n7636_8799.t64 gnd 0.590279f
C2065 a_n7636_8799.n136 gnd 0.269227f
C2066 a_n7636_8799.n137 gnd 0.24606f
C2067 a_n7636_8799.n138 gnd 0.267038f
C2068 a_n7636_8799.n139 gnd 0.269657f
C2069 a_n7636_8799.n140 gnd 0.263472f
C2070 a_n7636_8799.n141 gnd 0.25841f
C2071 a_n7636_8799.n142 gnd 0.267154f
C2072 a_n7636_8799.n143 gnd 0.269227f
C2073 a_n7636_8799.t83 gnd 0.600996f
C2074 a_n7636_8799.t43 gnd 0.590279f
C2075 a_n7636_8799.t86 gnd 0.590279f
C2076 a_n7636_8799.t84 gnd 0.590279f
C2077 a_n7636_8799.n144 gnd 0.263719f
C2078 a_n7636_8799.t45 gnd 0.590279f
C2079 a_n7636_8799.t44 gnd 0.590279f
C2080 a_n7636_8799.t101 gnd 0.590279f
C2081 a_n7636_8799.n145 gnd 0.267169f
C2082 a_n7636_8799.t55 gnd 0.590279f
C2083 a_n7636_8799.t46 gnd 0.590279f
C2084 a_n7636_8799.t102 gnd 0.590279f
C2085 a_n7636_8799.n146 gnd 0.263156f
C2086 a_n7636_8799.t56 gnd 0.604153f
C2087 a_n7636_8799.t72 gnd 0.590279f
C2088 a_n7636_8799.n147 gnd 0.269227f
C2089 a_n7636_8799.n148 gnd 0.24606f
C2090 a_n7636_8799.n149 gnd 0.267038f
C2091 a_n7636_8799.n150 gnd 0.269657f
C2092 a_n7636_8799.n151 gnd 0.263472f
C2093 a_n7636_8799.n152 gnd 0.25841f
C2094 a_n7636_8799.n153 gnd 0.267154f
C2095 a_n7636_8799.n154 gnd 0.269227f
C2096 a_n7636_8799.n155 gnd 0.886171f
C2097 a_n7636_8799.t52 gnd 0.600996f
C2098 a_n7636_8799.t105 gnd 0.590279f
C2099 a_n7636_8799.t82 gnd 0.590279f
C2100 a_n7636_8799.t99 gnd 0.590279f
C2101 a_n7636_8799.n156 gnd 0.263719f
C2102 a_n7636_8799.t70 gnd 0.590279f
C2103 a_n7636_8799.t85 gnd 0.590279f
C2104 a_n7636_8799.t47 gnd 0.590279f
C2105 a_n7636_8799.n157 gnd 0.267169f
C2106 a_n7636_8799.t97 gnd 0.590279f
C2107 a_n7636_8799.t58 gnd 0.590279f
C2108 a_n7636_8799.t93 gnd 0.590279f
C2109 a_n7636_8799.n158 gnd 0.263156f
C2110 a_n7636_8799.t79 gnd 0.604153f
C2111 a_n7636_8799.t51 gnd 0.590279f
C2112 a_n7636_8799.n159 gnd 0.269227f
C2113 a_n7636_8799.n160 gnd 0.24606f
C2114 a_n7636_8799.n161 gnd 0.267038f
C2115 a_n7636_8799.n162 gnd 0.269657f
C2116 a_n7636_8799.n163 gnd 0.263472f
C2117 a_n7636_8799.n164 gnd 0.25841f
C2118 a_n7636_8799.n165 gnd 0.267154f
C2119 a_n7636_8799.n166 gnd 0.269227f
C2120 a_n7636_8799.n167 gnd 1.29577f
C2121 a_n7636_8799.n168 gnd 15.4907f
C2122 a_n7636_8799.n169 gnd 4.319991f
C2123 a_n7636_8799.n170 gnd 6.90345f
C2124 a_n7636_8799.t29 gnd 0.142357f
C2125 a_n7636_8799.t33 gnd 0.142357f
C2126 a_n7636_8799.n171 gnd 1.12094f
C2127 a_n7636_8799.t21 gnd 0.142357f
C2128 a_n7636_8799.t16 gnd 0.142357f
C2129 a_n7636_8799.n172 gnd 1.12094f
C2130 a_n7636_8799.t18 gnd 0.142357f
C2131 a_n7636_8799.t30 gnd 0.142357f
C2132 a_n7636_8799.n173 gnd 1.12094f
C2133 a_n7636_8799.t22 gnd 0.142357f
C2134 a_n7636_8799.t26 gnd 0.142357f
C2135 a_n7636_8799.n174 gnd 1.12279f
C2136 a_n7636_8799.n175 gnd 1.12094f
C2137 a_n7636_8799.t14 gnd 0.142357f
C2138 vdd.t215 gnd 0.033456f
C2139 vdd.t196 gnd 0.033456f
C2140 vdd.n0 gnd 0.263872f
C2141 vdd.t177 gnd 0.033456f
C2142 vdd.t210 gnd 0.033456f
C2143 vdd.n1 gnd 0.263437f
C2144 vdd.n2 gnd 0.242939f
C2145 vdd.t193 gnd 0.033456f
C2146 vdd.t219 gnd 0.033456f
C2147 vdd.n3 gnd 0.263437f
C2148 vdd.n4 gnd 0.122863f
C2149 vdd.t221 gnd 0.033456f
C2150 vdd.t201 gnd 0.033456f
C2151 vdd.n5 gnd 0.263437f
C2152 vdd.n6 gnd 0.115284f
C2153 vdd.t225 gnd 0.033456f
C2154 vdd.t191 gnd 0.033456f
C2155 vdd.n7 gnd 0.263872f
C2156 vdd.t199 gnd 0.033456f
C2157 vdd.t217 gnd 0.033456f
C2158 vdd.n8 gnd 0.263437f
C2159 vdd.n9 gnd 0.242939f
C2160 vdd.t207 gnd 0.033456f
C2161 vdd.t180 gnd 0.033456f
C2162 vdd.n10 gnd 0.263437f
C2163 vdd.n11 gnd 0.122863f
C2164 vdd.t188 gnd 0.033456f
C2165 vdd.t205 gnd 0.033456f
C2166 vdd.n12 gnd 0.263437f
C2167 vdd.n13 gnd 0.115284f
C2168 vdd.n14 gnd 0.081504f
C2169 vdd.t8 gnd 0.018587f
C2170 vdd.t92 gnd 0.018587f
C2171 vdd.n15 gnd 0.171082f
C2172 vdd.t45 gnd 0.018587f
C2173 vdd.t37 gnd 0.018587f
C2174 vdd.n16 gnd 0.170581f
C2175 vdd.n17 gnd 0.296865f
C2176 vdd.t9 gnd 0.018587f
C2177 vdd.t44 gnd 0.018587f
C2178 vdd.n18 gnd 0.170581f
C2179 vdd.n19 gnd 0.122817f
C2180 vdd.t69 gnd 0.018587f
C2181 vdd.t39 gnd 0.018587f
C2182 vdd.n20 gnd 0.171082f
C2183 vdd.t41 gnd 0.018587f
C2184 vdd.t93 gnd 0.018587f
C2185 vdd.n21 gnd 0.170581f
C2186 vdd.n22 gnd 0.296865f
C2187 vdd.t42 gnd 0.018587f
C2188 vdd.t70 gnd 0.018587f
C2189 vdd.n23 gnd 0.170581f
C2190 vdd.n24 gnd 0.122817f
C2191 vdd.t38 gnd 0.018587f
C2192 vdd.t68 gnd 0.018587f
C2193 vdd.n25 gnd 0.170581f
C2194 vdd.t43 gnd 0.018587f
C2195 vdd.t40 gnd 0.018587f
C2196 vdd.n26 gnd 0.170581f
C2197 vdd.n27 gnd 18.6758f
C2198 vdd.n28 gnd 7.24673f
C2199 vdd.n29 gnd 0.005069f
C2200 vdd.n30 gnd 0.004704f
C2201 vdd.n31 gnd 0.002602f
C2202 vdd.n32 gnd 0.005975f
C2203 vdd.n33 gnd 0.002528f
C2204 vdd.n34 gnd 0.002676f
C2205 vdd.n35 gnd 0.004704f
C2206 vdd.n36 gnd 0.002528f
C2207 vdd.n37 gnd 0.005975f
C2208 vdd.n38 gnd 0.002676f
C2209 vdd.n39 gnd 0.004704f
C2210 vdd.n40 gnd 0.002528f
C2211 vdd.n41 gnd 0.004481f
C2212 vdd.n42 gnd 0.004494f
C2213 vdd.t15 gnd 0.012836f
C2214 vdd.n43 gnd 0.02856f
C2215 vdd.n44 gnd 0.148635f
C2216 vdd.n45 gnd 0.002528f
C2217 vdd.n46 gnd 0.002676f
C2218 vdd.n47 gnd 0.005975f
C2219 vdd.n48 gnd 0.005975f
C2220 vdd.n49 gnd 0.002676f
C2221 vdd.n50 gnd 0.002528f
C2222 vdd.n51 gnd 0.004704f
C2223 vdd.n52 gnd 0.004704f
C2224 vdd.n53 gnd 0.002528f
C2225 vdd.n54 gnd 0.002676f
C2226 vdd.n55 gnd 0.005975f
C2227 vdd.n56 gnd 0.005975f
C2228 vdd.n57 gnd 0.002676f
C2229 vdd.n58 gnd 0.002528f
C2230 vdd.n59 gnd 0.004704f
C2231 vdd.n60 gnd 0.004704f
C2232 vdd.n61 gnd 0.002528f
C2233 vdd.n62 gnd 0.002676f
C2234 vdd.n63 gnd 0.005975f
C2235 vdd.n64 gnd 0.005975f
C2236 vdd.n65 gnd 0.014125f
C2237 vdd.n66 gnd 0.002602f
C2238 vdd.n67 gnd 0.002528f
C2239 vdd.n68 gnd 0.012159f
C2240 vdd.n69 gnd 0.008488f
C2241 vdd.t227 gnd 0.029739f
C2242 vdd.t228 gnd 0.029739f
C2243 vdd.n70 gnd 0.204384f
C2244 vdd.n71 gnd 0.160717f
C2245 vdd.t65 gnd 0.029739f
C2246 vdd.t19 gnd 0.029739f
C2247 vdd.n72 gnd 0.204384f
C2248 vdd.n73 gnd 0.129698f
C2249 vdd.t67 gnd 0.029739f
C2250 vdd.t61 gnd 0.029739f
C2251 vdd.n74 gnd 0.204384f
C2252 vdd.n75 gnd 0.129698f
C2253 vdd.t28 gnd 0.029739f
C2254 vdd.t22 gnd 0.029739f
C2255 vdd.n76 gnd 0.204384f
C2256 vdd.n77 gnd 0.129698f
C2257 vdd.t89 gnd 0.029739f
C2258 vdd.t3 gnd 0.029739f
C2259 vdd.n78 gnd 0.204384f
C2260 vdd.n79 gnd 0.129698f
C2261 vdd.n80 gnd 0.005069f
C2262 vdd.n81 gnd 0.004704f
C2263 vdd.n82 gnd 0.002602f
C2264 vdd.n83 gnd 0.005975f
C2265 vdd.n84 gnd 0.002528f
C2266 vdd.n85 gnd 0.002676f
C2267 vdd.n86 gnd 0.004704f
C2268 vdd.n87 gnd 0.002528f
C2269 vdd.n88 gnd 0.005975f
C2270 vdd.n89 gnd 0.002676f
C2271 vdd.n90 gnd 0.004704f
C2272 vdd.n91 gnd 0.002528f
C2273 vdd.n92 gnd 0.004481f
C2274 vdd.n93 gnd 0.004494f
C2275 vdd.t173 gnd 0.012836f
C2276 vdd.n94 gnd 0.02856f
C2277 vdd.n95 gnd 0.148635f
C2278 vdd.n96 gnd 0.002528f
C2279 vdd.n97 gnd 0.002676f
C2280 vdd.n98 gnd 0.005975f
C2281 vdd.n99 gnd 0.005975f
C2282 vdd.n100 gnd 0.002676f
C2283 vdd.n101 gnd 0.002528f
C2284 vdd.n102 gnd 0.004704f
C2285 vdd.n103 gnd 0.004704f
C2286 vdd.n104 gnd 0.002528f
C2287 vdd.n105 gnd 0.002676f
C2288 vdd.n106 gnd 0.005975f
C2289 vdd.n107 gnd 0.005975f
C2290 vdd.n108 gnd 0.002676f
C2291 vdd.n109 gnd 0.002528f
C2292 vdd.n110 gnd 0.004704f
C2293 vdd.n111 gnd 0.004704f
C2294 vdd.n112 gnd 0.002528f
C2295 vdd.n113 gnd 0.002676f
C2296 vdd.n114 gnd 0.005975f
C2297 vdd.n115 gnd 0.005975f
C2298 vdd.n116 gnd 0.014125f
C2299 vdd.n117 gnd 0.002602f
C2300 vdd.n118 gnd 0.002528f
C2301 vdd.n119 gnd 0.012159f
C2302 vdd.n120 gnd 0.008222f
C2303 vdd.n121 gnd 0.096496f
C2304 vdd.n122 gnd 0.005069f
C2305 vdd.n123 gnd 0.004704f
C2306 vdd.n124 gnd 0.002602f
C2307 vdd.n125 gnd 0.005975f
C2308 vdd.n126 gnd 0.002528f
C2309 vdd.n127 gnd 0.002676f
C2310 vdd.n128 gnd 0.004704f
C2311 vdd.n129 gnd 0.002528f
C2312 vdd.n130 gnd 0.005975f
C2313 vdd.n131 gnd 0.002676f
C2314 vdd.n132 gnd 0.004704f
C2315 vdd.n133 gnd 0.002528f
C2316 vdd.n134 gnd 0.004481f
C2317 vdd.n135 gnd 0.004494f
C2318 vdd.t229 gnd 0.012836f
C2319 vdd.n136 gnd 0.02856f
C2320 vdd.n137 gnd 0.148635f
C2321 vdd.n138 gnd 0.002528f
C2322 vdd.n139 gnd 0.002676f
C2323 vdd.n140 gnd 0.005975f
C2324 vdd.n141 gnd 0.005975f
C2325 vdd.n142 gnd 0.002676f
C2326 vdd.n143 gnd 0.002528f
C2327 vdd.n144 gnd 0.004704f
C2328 vdd.n145 gnd 0.004704f
C2329 vdd.n146 gnd 0.002528f
C2330 vdd.n147 gnd 0.002676f
C2331 vdd.n148 gnd 0.005975f
C2332 vdd.n149 gnd 0.005975f
C2333 vdd.n150 gnd 0.002676f
C2334 vdd.n151 gnd 0.002528f
C2335 vdd.n152 gnd 0.004704f
C2336 vdd.n153 gnd 0.004704f
C2337 vdd.n154 gnd 0.002528f
C2338 vdd.n155 gnd 0.002676f
C2339 vdd.n156 gnd 0.005975f
C2340 vdd.n157 gnd 0.005975f
C2341 vdd.n158 gnd 0.014125f
C2342 vdd.n159 gnd 0.002602f
C2343 vdd.n160 gnd 0.002528f
C2344 vdd.n161 gnd 0.012159f
C2345 vdd.n162 gnd 0.008488f
C2346 vdd.t76 gnd 0.029739f
C2347 vdd.t238 gnd 0.029739f
C2348 vdd.n163 gnd 0.204384f
C2349 vdd.n164 gnd 0.160717f
C2350 vdd.t66 gnd 0.029739f
C2351 vdd.t235 gnd 0.029739f
C2352 vdd.n165 gnd 0.204384f
C2353 vdd.n166 gnd 0.129698f
C2354 vdd.t234 gnd 0.029739f
C2355 vdd.t171 gnd 0.029739f
C2356 vdd.n167 gnd 0.204384f
C2357 vdd.n168 gnd 0.129698f
C2358 vdd.t74 gnd 0.029739f
C2359 vdd.t60 gnd 0.029739f
C2360 vdd.n169 gnd 0.204384f
C2361 vdd.n170 gnd 0.129698f
C2362 vdd.t58 gnd 0.029739f
C2363 vdd.t77 gnd 0.029739f
C2364 vdd.n171 gnd 0.204384f
C2365 vdd.n172 gnd 0.129698f
C2366 vdd.n173 gnd 0.005069f
C2367 vdd.n174 gnd 0.004704f
C2368 vdd.n175 gnd 0.002602f
C2369 vdd.n176 gnd 0.005975f
C2370 vdd.n177 gnd 0.002528f
C2371 vdd.n178 gnd 0.002676f
C2372 vdd.n179 gnd 0.004704f
C2373 vdd.n180 gnd 0.002528f
C2374 vdd.n181 gnd 0.005975f
C2375 vdd.n182 gnd 0.002676f
C2376 vdd.n183 gnd 0.004704f
C2377 vdd.n184 gnd 0.002528f
C2378 vdd.n185 gnd 0.004481f
C2379 vdd.n186 gnd 0.004494f
C2380 vdd.t46 gnd 0.012836f
C2381 vdd.n187 gnd 0.02856f
C2382 vdd.n188 gnd 0.148635f
C2383 vdd.n189 gnd 0.002528f
C2384 vdd.n190 gnd 0.002676f
C2385 vdd.n191 gnd 0.005975f
C2386 vdd.n192 gnd 0.005975f
C2387 vdd.n193 gnd 0.002676f
C2388 vdd.n194 gnd 0.002528f
C2389 vdd.n195 gnd 0.004704f
C2390 vdd.n196 gnd 0.004704f
C2391 vdd.n197 gnd 0.002528f
C2392 vdd.n198 gnd 0.002676f
C2393 vdd.n199 gnd 0.005975f
C2394 vdd.n200 gnd 0.005975f
C2395 vdd.n201 gnd 0.002676f
C2396 vdd.n202 gnd 0.002528f
C2397 vdd.n203 gnd 0.004704f
C2398 vdd.n204 gnd 0.004704f
C2399 vdd.n205 gnd 0.002528f
C2400 vdd.n206 gnd 0.002676f
C2401 vdd.n207 gnd 0.005975f
C2402 vdd.n208 gnd 0.005975f
C2403 vdd.n209 gnd 0.014125f
C2404 vdd.n210 gnd 0.002602f
C2405 vdd.n211 gnd 0.002528f
C2406 vdd.n212 gnd 0.012159f
C2407 vdd.n213 gnd 0.008222f
C2408 vdd.n214 gnd 0.057405f
C2409 vdd.n215 gnd 0.206846f
C2410 vdd.n216 gnd 0.005069f
C2411 vdd.n217 gnd 0.004704f
C2412 vdd.n218 gnd 0.002602f
C2413 vdd.n219 gnd 0.005975f
C2414 vdd.n220 gnd 0.002528f
C2415 vdd.n221 gnd 0.002676f
C2416 vdd.n222 gnd 0.004704f
C2417 vdd.n223 gnd 0.002528f
C2418 vdd.n224 gnd 0.005975f
C2419 vdd.n225 gnd 0.002676f
C2420 vdd.n226 gnd 0.004704f
C2421 vdd.n227 gnd 0.002528f
C2422 vdd.n228 gnd 0.004481f
C2423 vdd.n229 gnd 0.004494f
C2424 vdd.t78 gnd 0.012836f
C2425 vdd.n230 gnd 0.02856f
C2426 vdd.n231 gnd 0.148635f
C2427 vdd.n232 gnd 0.002528f
C2428 vdd.n233 gnd 0.002676f
C2429 vdd.n234 gnd 0.005975f
C2430 vdd.n235 gnd 0.005975f
C2431 vdd.n236 gnd 0.002676f
C2432 vdd.n237 gnd 0.002528f
C2433 vdd.n238 gnd 0.004704f
C2434 vdd.n239 gnd 0.004704f
C2435 vdd.n240 gnd 0.002528f
C2436 vdd.n241 gnd 0.002676f
C2437 vdd.n242 gnd 0.005975f
C2438 vdd.n243 gnd 0.005975f
C2439 vdd.n244 gnd 0.002676f
C2440 vdd.n245 gnd 0.002528f
C2441 vdd.n246 gnd 0.004704f
C2442 vdd.n247 gnd 0.004704f
C2443 vdd.n248 gnd 0.002528f
C2444 vdd.n249 gnd 0.002676f
C2445 vdd.n250 gnd 0.005975f
C2446 vdd.n251 gnd 0.005975f
C2447 vdd.n252 gnd 0.014125f
C2448 vdd.n253 gnd 0.002602f
C2449 vdd.n254 gnd 0.002528f
C2450 vdd.n255 gnd 0.012159f
C2451 vdd.n256 gnd 0.008488f
C2452 vdd.t34 gnd 0.029739f
C2453 vdd.t83 gnd 0.029739f
C2454 vdd.n257 gnd 0.204384f
C2455 vdd.n258 gnd 0.160717f
C2456 vdd.t81 gnd 0.029739f
C2457 vdd.t71 gnd 0.029739f
C2458 vdd.n259 gnd 0.204384f
C2459 vdd.n260 gnd 0.129698f
C2460 vdd.t36 gnd 0.029739f
C2461 vdd.t11 gnd 0.029739f
C2462 vdd.n261 gnd 0.204384f
C2463 vdd.n262 gnd 0.129698f
C2464 vdd.t85 gnd 0.029739f
C2465 vdd.t72 gnd 0.029739f
C2466 vdd.n263 gnd 0.204384f
C2467 vdd.n264 gnd 0.129698f
C2468 vdd.t88 gnd 0.029739f
C2469 vdd.t232 gnd 0.029739f
C2470 vdd.n265 gnd 0.204384f
C2471 vdd.n266 gnd 0.129698f
C2472 vdd.n267 gnd 0.005069f
C2473 vdd.n268 gnd 0.004704f
C2474 vdd.n269 gnd 0.002602f
C2475 vdd.n270 gnd 0.005975f
C2476 vdd.n271 gnd 0.002528f
C2477 vdd.n272 gnd 0.002676f
C2478 vdd.n273 gnd 0.004704f
C2479 vdd.n274 gnd 0.002528f
C2480 vdd.n275 gnd 0.005975f
C2481 vdd.n276 gnd 0.002676f
C2482 vdd.n277 gnd 0.004704f
C2483 vdd.n278 gnd 0.002528f
C2484 vdd.n279 gnd 0.004481f
C2485 vdd.n280 gnd 0.004494f
C2486 vdd.t1 gnd 0.012836f
C2487 vdd.n281 gnd 0.02856f
C2488 vdd.n282 gnd 0.148635f
C2489 vdd.n283 gnd 0.002528f
C2490 vdd.n284 gnd 0.002676f
C2491 vdd.n285 gnd 0.005975f
C2492 vdd.n286 gnd 0.005975f
C2493 vdd.n287 gnd 0.002676f
C2494 vdd.n288 gnd 0.002528f
C2495 vdd.n289 gnd 0.004704f
C2496 vdd.n290 gnd 0.004704f
C2497 vdd.n291 gnd 0.002528f
C2498 vdd.n292 gnd 0.002676f
C2499 vdd.n293 gnd 0.005975f
C2500 vdd.n294 gnd 0.005975f
C2501 vdd.n295 gnd 0.002676f
C2502 vdd.n296 gnd 0.002528f
C2503 vdd.n297 gnd 0.004704f
C2504 vdd.n298 gnd 0.004704f
C2505 vdd.n299 gnd 0.002528f
C2506 vdd.n300 gnd 0.002676f
C2507 vdd.n301 gnd 0.005975f
C2508 vdd.n302 gnd 0.005975f
C2509 vdd.n303 gnd 0.014125f
C2510 vdd.n304 gnd 0.002602f
C2511 vdd.n305 gnd 0.002528f
C2512 vdd.n306 gnd 0.012159f
C2513 vdd.n307 gnd 0.008222f
C2514 vdd.n308 gnd 0.057405f
C2515 vdd.n309 gnd 0.22733f
C2516 vdd.n310 gnd 0.009205f
C2517 vdd.n311 gnd 0.009205f
C2518 vdd.n312 gnd 0.007435f
C2519 vdd.n313 gnd 0.007435f
C2520 vdd.n314 gnd 0.009237f
C2521 vdd.n315 gnd 0.009237f
C2522 vdd.t35 gnd 0.471988f
C2523 vdd.n316 gnd 0.009237f
C2524 vdd.n317 gnd 0.009237f
C2525 vdd.n318 gnd 0.009237f
C2526 vdd.t27 gnd 0.471988f
C2527 vdd.n319 gnd 0.009237f
C2528 vdd.n320 gnd 0.009237f
C2529 vdd.n321 gnd 0.009237f
C2530 vdd.n322 gnd 0.009237f
C2531 vdd.n323 gnd 0.007435f
C2532 vdd.n324 gnd 0.009237f
C2533 vdd.n325 gnd 0.7599f
C2534 vdd.n326 gnd 0.009237f
C2535 vdd.n327 gnd 0.009237f
C2536 vdd.n328 gnd 0.009237f
C2537 vdd.n329 gnd 0.646623f
C2538 vdd.n330 gnd 0.009237f
C2539 vdd.n331 gnd 0.009237f
C2540 vdd.n332 gnd 0.009237f
C2541 vdd.n333 gnd 0.009237f
C2542 vdd.n334 gnd 0.009237f
C2543 vdd.n335 gnd 0.007435f
C2544 vdd.n336 gnd 0.009237f
C2545 vdd.t2 gnd 0.471988f
C2546 vdd.n337 gnd 0.009237f
C2547 vdd.n338 gnd 0.009237f
C2548 vdd.n339 gnd 0.009237f
C2549 vdd.n340 gnd 0.943976f
C2550 vdd.n341 gnd 0.009237f
C2551 vdd.n342 gnd 0.009237f
C2552 vdd.n343 gnd 0.009237f
C2553 vdd.n344 gnd 0.009237f
C2554 vdd.n345 gnd 0.009237f
C2555 vdd.n346 gnd 0.007435f
C2556 vdd.n347 gnd 0.009237f
C2557 vdd.n348 gnd 0.009237f
C2558 vdd.n349 gnd 0.009237f
C2559 vdd.n350 gnd 0.021768f
C2560 vdd.n351 gnd 2.17114f
C2561 vdd.n352 gnd 0.022108f
C2562 vdd.n353 gnd 0.009237f
C2563 vdd.n354 gnd 0.009237f
C2564 vdd.n356 gnd 0.009237f
C2565 vdd.n357 gnd 0.009237f
C2566 vdd.n358 gnd 0.007435f
C2567 vdd.n359 gnd 0.007435f
C2568 vdd.n360 gnd 0.009237f
C2569 vdd.n361 gnd 0.009237f
C2570 vdd.n362 gnd 0.009237f
C2571 vdd.n363 gnd 0.009237f
C2572 vdd.n364 gnd 0.009237f
C2573 vdd.n365 gnd 0.009237f
C2574 vdd.n366 gnd 0.007435f
C2575 vdd.n368 gnd 0.009237f
C2576 vdd.n369 gnd 0.009237f
C2577 vdd.n370 gnd 0.009237f
C2578 vdd.n371 gnd 0.009237f
C2579 vdd.n372 gnd 0.009237f
C2580 vdd.n373 gnd 0.007435f
C2581 vdd.n375 gnd 0.009237f
C2582 vdd.n376 gnd 0.009237f
C2583 vdd.n377 gnd 0.009237f
C2584 vdd.n378 gnd 0.009237f
C2585 vdd.n379 gnd 0.009237f
C2586 vdd.n380 gnd 0.007435f
C2587 vdd.n382 gnd 0.009237f
C2588 vdd.n383 gnd 0.009237f
C2589 vdd.n384 gnd 0.009237f
C2590 vdd.n385 gnd 0.009237f
C2591 vdd.n386 gnd 0.006208f
C2592 vdd.t169 gnd 0.113639f
C2593 vdd.t168 gnd 0.121449f
C2594 vdd.t167 gnd 0.148411f
C2595 vdd.n387 gnd 0.190242f
C2596 vdd.n388 gnd 0.160581f
C2597 vdd.n390 gnd 0.009237f
C2598 vdd.n391 gnd 0.009237f
C2599 vdd.n392 gnd 0.007435f
C2600 vdd.n393 gnd 0.009237f
C2601 vdd.n395 gnd 0.009237f
C2602 vdd.n396 gnd 0.009237f
C2603 vdd.n397 gnd 0.009237f
C2604 vdd.n398 gnd 0.009237f
C2605 vdd.n399 gnd 0.007435f
C2606 vdd.n401 gnd 0.009237f
C2607 vdd.n402 gnd 0.009237f
C2608 vdd.n403 gnd 0.009237f
C2609 vdd.n404 gnd 0.009237f
C2610 vdd.n405 gnd 0.009237f
C2611 vdd.n406 gnd 0.007435f
C2612 vdd.n408 gnd 0.009237f
C2613 vdd.n409 gnd 0.009237f
C2614 vdd.n410 gnd 0.009237f
C2615 vdd.n411 gnd 0.009237f
C2616 vdd.n412 gnd 0.009237f
C2617 vdd.n413 gnd 0.007435f
C2618 vdd.n415 gnd 0.009237f
C2619 vdd.n416 gnd 0.009237f
C2620 vdd.n417 gnd 0.009237f
C2621 vdd.n418 gnd 0.009237f
C2622 vdd.n419 gnd 0.009237f
C2623 vdd.n420 gnd 0.007435f
C2624 vdd.n422 gnd 0.009237f
C2625 vdd.n423 gnd 0.009237f
C2626 vdd.n424 gnd 0.009237f
C2627 vdd.n425 gnd 0.009237f
C2628 vdd.n426 gnd 0.00736f
C2629 vdd.t163 gnd 0.113639f
C2630 vdd.t162 gnd 0.121449f
C2631 vdd.t161 gnd 0.148411f
C2632 vdd.n427 gnd 0.190242f
C2633 vdd.n428 gnd 0.160581f
C2634 vdd.n430 gnd 0.009237f
C2635 vdd.n431 gnd 0.009237f
C2636 vdd.n432 gnd 0.007435f
C2637 vdd.n433 gnd 0.009237f
C2638 vdd.n435 gnd 0.009237f
C2639 vdd.n436 gnd 0.009237f
C2640 vdd.n437 gnd 0.009237f
C2641 vdd.n438 gnd 0.009237f
C2642 vdd.n439 gnd 0.007435f
C2643 vdd.n441 gnd 0.009237f
C2644 vdd.n442 gnd 0.009237f
C2645 vdd.n443 gnd 0.009237f
C2646 vdd.n444 gnd 0.009237f
C2647 vdd.n445 gnd 0.009237f
C2648 vdd.n446 gnd 0.007435f
C2649 vdd.n448 gnd 0.009237f
C2650 vdd.n449 gnd 0.009237f
C2651 vdd.n450 gnd 0.009237f
C2652 vdd.n451 gnd 0.009237f
C2653 vdd.n452 gnd 0.009237f
C2654 vdd.n453 gnd 0.007435f
C2655 vdd.n455 gnd 0.009237f
C2656 vdd.n456 gnd 0.009237f
C2657 vdd.n457 gnd 0.009237f
C2658 vdd.n458 gnd 0.009237f
C2659 vdd.n459 gnd 0.009237f
C2660 vdd.n460 gnd 0.007435f
C2661 vdd.n462 gnd 0.009237f
C2662 vdd.n463 gnd 0.009237f
C2663 vdd.n464 gnd 0.009237f
C2664 vdd.n465 gnd 0.009237f
C2665 vdd.n466 gnd 0.009237f
C2666 vdd.n467 gnd 0.009237f
C2667 vdd.n468 gnd 0.007435f
C2668 vdd.n469 gnd 0.009237f
C2669 vdd.n470 gnd 0.009237f
C2670 vdd.n471 gnd 0.007435f
C2671 vdd.n472 gnd 0.009237f
C2672 vdd.n473 gnd 0.009237f
C2673 vdd.n474 gnd 0.007435f
C2674 vdd.n475 gnd 0.009237f
C2675 vdd.n476 gnd 0.007435f
C2676 vdd.n477 gnd 0.009237f
C2677 vdd.n478 gnd 0.007435f
C2678 vdd.n479 gnd 0.009237f
C2679 vdd.n480 gnd 0.009237f
C2680 vdd.t18 gnd 0.471988f
C2681 vdd.n481 gnd 0.505027f
C2682 vdd.n482 gnd 0.009237f
C2683 vdd.n483 gnd 0.007435f
C2684 vdd.n484 gnd 0.009237f
C2685 vdd.n485 gnd 0.007435f
C2686 vdd.n486 gnd 0.009237f
C2687 vdd.t64 gnd 0.471988f
C2688 vdd.n487 gnd 0.009237f
C2689 vdd.n488 gnd 0.007435f
C2690 vdd.n489 gnd 0.009237f
C2691 vdd.n490 gnd 0.007435f
C2692 vdd.n491 gnd 0.009237f
C2693 vdd.n492 gnd 0.741021f
C2694 vdd.n493 gnd 0.7835f
C2695 vdd.t82 gnd 0.471988f
C2696 vdd.n494 gnd 0.009237f
C2697 vdd.n495 gnd 0.007435f
C2698 vdd.n496 gnd 0.009237f
C2699 vdd.n497 gnd 0.007435f
C2700 vdd.n498 gnd 0.009237f
C2701 vdd.n499 gnd 0.580545f
C2702 vdd.n500 gnd 0.009237f
C2703 vdd.n501 gnd 0.007435f
C2704 vdd.n502 gnd 0.009237f
C2705 vdd.n503 gnd 0.007435f
C2706 vdd.n504 gnd 0.009237f
C2707 vdd.n505 gnd 0.943976f
C2708 vdd.t14 gnd 0.471988f
C2709 vdd.n506 gnd 0.009237f
C2710 vdd.n507 gnd 0.007435f
C2711 vdd.n508 gnd 0.009237f
C2712 vdd.n509 gnd 0.007435f
C2713 vdd.n510 gnd 0.009237f
C2714 vdd.n511 gnd 0.505027f
C2715 vdd.n512 gnd 0.009237f
C2716 vdd.n513 gnd 0.007435f
C2717 vdd.n514 gnd 0.022108f
C2718 vdd.n515 gnd 0.022108f
C2719 vdd.n516 gnd 9.892871f
C2720 vdd.t95 gnd 0.471988f
C2721 vdd.n517 gnd 0.022108f
C2722 vdd.n518 gnd 0.007944f
C2723 vdd.n519 gnd 0.007435f
C2724 vdd.n524 gnd 0.005912f
C2725 vdd.n525 gnd 0.007435f
C2726 vdd.n526 gnd 0.009237f
C2727 vdd.n527 gnd 0.009237f
C2728 vdd.n528 gnd 0.009237f
C2729 vdd.n529 gnd 0.009237f
C2730 vdd.n530 gnd 0.009237f
C2731 vdd.n531 gnd 0.007435f
C2732 vdd.n532 gnd 0.009237f
C2733 vdd.n533 gnd 0.009237f
C2734 vdd.n534 gnd 0.009237f
C2735 vdd.n535 gnd 0.009237f
C2736 vdd.n536 gnd 0.009237f
C2737 vdd.n537 gnd 0.007435f
C2738 vdd.n538 gnd 0.009237f
C2739 vdd.n539 gnd 0.009237f
C2740 vdd.n540 gnd 0.009237f
C2741 vdd.n541 gnd 0.009237f
C2742 vdd.n542 gnd 0.009237f
C2743 vdd.t107 gnd 0.113639f
C2744 vdd.t108 gnd 0.121449f
C2745 vdd.t106 gnd 0.148411f
C2746 vdd.n543 gnd 0.190242f
C2747 vdd.n544 gnd 0.159838f
C2748 vdd.n545 gnd 0.015167f
C2749 vdd.n546 gnd 0.009237f
C2750 vdd.n547 gnd 0.009237f
C2751 vdd.n548 gnd 0.009237f
C2752 vdd.n549 gnd 0.009237f
C2753 vdd.n550 gnd 0.009237f
C2754 vdd.n551 gnd 0.007435f
C2755 vdd.n552 gnd 0.009237f
C2756 vdd.n553 gnd 0.009237f
C2757 vdd.n554 gnd 0.009237f
C2758 vdd.n555 gnd 0.009237f
C2759 vdd.n556 gnd 0.009237f
C2760 vdd.n557 gnd 0.007435f
C2761 vdd.n558 gnd 0.009237f
C2762 vdd.n559 gnd 0.009237f
C2763 vdd.n560 gnd 0.009237f
C2764 vdd.n561 gnd 0.009237f
C2765 vdd.n562 gnd 0.009237f
C2766 vdd.n563 gnd 0.007435f
C2767 vdd.n564 gnd 0.009237f
C2768 vdd.n565 gnd 0.009237f
C2769 vdd.n566 gnd 0.009237f
C2770 vdd.n567 gnd 0.009237f
C2771 vdd.n568 gnd 0.009237f
C2772 vdd.n569 gnd 0.007435f
C2773 vdd.n570 gnd 0.009237f
C2774 vdd.n571 gnd 0.009237f
C2775 vdd.n572 gnd 0.009237f
C2776 vdd.n573 gnd 0.009237f
C2777 vdd.n574 gnd 0.009237f
C2778 vdd.n575 gnd 0.007435f
C2779 vdd.n576 gnd 0.009237f
C2780 vdd.n577 gnd 0.009237f
C2781 vdd.n578 gnd 0.009237f
C2782 vdd.n579 gnd 0.00736f
C2783 vdd.t96 gnd 0.113639f
C2784 vdd.t97 gnd 0.121449f
C2785 vdd.t94 gnd 0.148411f
C2786 vdd.n580 gnd 0.190242f
C2787 vdd.n581 gnd 0.159838f
C2788 vdd.n582 gnd 0.009237f
C2789 vdd.n583 gnd 0.007435f
C2790 vdd.n585 gnd 0.009237f
C2791 vdd.n587 gnd 0.009237f
C2792 vdd.n588 gnd 0.009237f
C2793 vdd.n589 gnd 0.007435f
C2794 vdd.n590 gnd 0.009237f
C2795 vdd.n591 gnd 0.009237f
C2796 vdd.n592 gnd 0.009237f
C2797 vdd.n593 gnd 0.009237f
C2798 vdd.n594 gnd 0.009237f
C2799 vdd.n595 gnd 0.007435f
C2800 vdd.n596 gnd 0.009237f
C2801 vdd.n597 gnd 0.009237f
C2802 vdd.n598 gnd 0.009237f
C2803 vdd.n599 gnd 0.009237f
C2804 vdd.n600 gnd 0.009237f
C2805 vdd.n601 gnd 0.007435f
C2806 vdd.n602 gnd 0.009237f
C2807 vdd.n603 gnd 0.009237f
C2808 vdd.n604 gnd 0.009237f
C2809 vdd.n605 gnd 0.005912f
C2810 vdd.n610 gnd 0.006281f
C2811 vdd.n611 gnd 0.006281f
C2812 vdd.n612 gnd 0.006281f
C2813 vdd.n613 gnd 9.600231f
C2814 vdd.n614 gnd 0.006281f
C2815 vdd.n615 gnd 0.006281f
C2816 vdd.n616 gnd 0.006281f
C2817 vdd.n618 gnd 0.006281f
C2818 vdd.n619 gnd 0.006281f
C2819 vdd.n621 gnd 0.006281f
C2820 vdd.n622 gnd 0.004572f
C2821 vdd.n624 gnd 0.006281f
C2822 vdd.t101 gnd 0.25382f
C2823 vdd.t100 gnd 0.259817f
C2824 vdd.t98 gnd 0.165704f
C2825 vdd.n625 gnd 0.089554f
C2826 vdd.n626 gnd 0.050798f
C2827 vdd.n627 gnd 0.008977f
C2828 vdd.n628 gnd 0.0144f
C2829 vdd.n630 gnd 0.006281f
C2830 vdd.n631 gnd 0.641903f
C2831 vdd.n632 gnd 0.013603f
C2832 vdd.n633 gnd 0.013603f
C2833 vdd.n634 gnd 0.006281f
C2834 vdd.n635 gnd 0.014477f
C2835 vdd.n636 gnd 0.006281f
C2836 vdd.n637 gnd 0.006281f
C2837 vdd.n638 gnd 0.006281f
C2838 vdd.n639 gnd 0.006281f
C2839 vdd.n640 gnd 0.006281f
C2840 vdd.n642 gnd 0.006281f
C2841 vdd.n643 gnd 0.006281f
C2842 vdd.n645 gnd 0.006281f
C2843 vdd.n646 gnd 0.006281f
C2844 vdd.n648 gnd 0.006281f
C2845 vdd.n649 gnd 0.006281f
C2846 vdd.n651 gnd 0.006281f
C2847 vdd.n652 gnd 0.006281f
C2848 vdd.n654 gnd 0.006281f
C2849 vdd.n655 gnd 0.006281f
C2850 vdd.n657 gnd 0.006281f
C2851 vdd.n658 gnd 0.004572f
C2852 vdd.n660 gnd 0.006281f
C2853 vdd.t136 gnd 0.25382f
C2854 vdd.t135 gnd 0.259817f
C2855 vdd.t134 gnd 0.165704f
C2856 vdd.n661 gnd 0.089554f
C2857 vdd.n662 gnd 0.050798f
C2858 vdd.n663 gnd 0.008977f
C2859 vdd.n664 gnd 0.006281f
C2860 vdd.n665 gnd 0.006281f
C2861 vdd.t99 gnd 0.320952f
C2862 vdd.n666 gnd 0.006281f
C2863 vdd.n667 gnd 0.006281f
C2864 vdd.n668 gnd 0.006281f
C2865 vdd.n669 gnd 0.006281f
C2866 vdd.n670 gnd 0.006281f
C2867 vdd.n671 gnd 0.641903f
C2868 vdd.n672 gnd 0.006281f
C2869 vdd.n673 gnd 0.006281f
C2870 vdd.n674 gnd 0.523906f
C2871 vdd.n675 gnd 0.006281f
C2872 vdd.n676 gnd 0.006281f
C2873 vdd.n677 gnd 0.006281f
C2874 vdd.n678 gnd 0.006281f
C2875 vdd.n679 gnd 0.641903f
C2876 vdd.n680 gnd 0.006281f
C2877 vdd.n681 gnd 0.006281f
C2878 vdd.n682 gnd 0.006281f
C2879 vdd.n683 gnd 0.006281f
C2880 vdd.n684 gnd 0.006281f
C2881 vdd.t202 gnd 0.320952f
C2882 vdd.n685 gnd 0.006281f
C2883 vdd.n686 gnd 0.006281f
C2884 vdd.n687 gnd 0.006281f
C2885 vdd.n688 gnd 0.006281f
C2886 vdd.n689 gnd 0.006281f
C2887 vdd.t208 gnd 0.320952f
C2888 vdd.n690 gnd 0.006281f
C2889 vdd.n691 gnd 0.006281f
C2890 vdd.n692 gnd 0.637184f
C2891 vdd.n693 gnd 0.006281f
C2892 vdd.n694 gnd 0.006281f
C2893 vdd.n695 gnd 0.006281f
C2894 vdd.t211 gnd 0.320952f
C2895 vdd.n696 gnd 0.006281f
C2896 vdd.n697 gnd 0.006281f
C2897 vdd.n698 gnd 0.495587f
C2898 vdd.n699 gnd 0.006281f
C2899 vdd.n700 gnd 0.006281f
C2900 vdd.n701 gnd 0.006281f
C2901 vdd.n702 gnd 0.429509f
C2902 vdd.n703 gnd 0.006281f
C2903 vdd.n704 gnd 0.006281f
C2904 vdd.n705 gnd 0.353991f
C2905 vdd.n706 gnd 0.006281f
C2906 vdd.n707 gnd 0.006281f
C2907 vdd.n708 gnd 0.006281f
C2908 vdd.n709 gnd 0.528626f
C2909 vdd.n710 gnd 0.006281f
C2910 vdd.n711 gnd 0.006281f
C2911 vdd.t181 gnd 0.320952f
C2912 vdd.n712 gnd 0.006281f
C2913 vdd.t111 gnd 0.259817f
C2914 vdd.t109 gnd 0.165704f
C2915 vdd.t112 gnd 0.259817f
C2916 vdd.n713 gnd 0.146028f
C2917 vdd.n714 gnd 0.006281f
C2918 vdd.n715 gnd 0.006281f
C2919 vdd.n716 gnd 0.641903f
C2920 vdd.n717 gnd 0.006281f
C2921 vdd.n718 gnd 0.006281f
C2922 vdd.t110 gnd 0.250154f
C2923 vdd.t183 gnd 0.113277f
C2924 vdd.n719 gnd 0.006281f
C2925 vdd.n720 gnd 0.006281f
C2926 vdd.n721 gnd 0.006281f
C2927 vdd.t194 gnd 0.320952f
C2928 vdd.n722 gnd 0.006281f
C2929 vdd.n723 gnd 0.006281f
C2930 vdd.n724 gnd 0.006281f
C2931 vdd.n725 gnd 0.006281f
C2932 vdd.n726 gnd 0.006281f
C2933 vdd.t212 gnd 0.320952f
C2934 vdd.n727 gnd 0.006281f
C2935 vdd.n728 gnd 0.006281f
C2936 vdd.n729 gnd 0.571105f
C2937 vdd.n730 gnd 0.006281f
C2938 vdd.n731 gnd 0.006281f
C2939 vdd.n732 gnd 0.006281f
C2940 vdd.n733 gnd 0.353991f
C2941 vdd.n734 gnd 0.006281f
C2942 vdd.n735 gnd 0.006281f
C2943 vdd.t190 gnd 0.320952f
C2944 vdd.n736 gnd 0.006281f
C2945 vdd.n737 gnd 0.006281f
C2946 vdd.n738 gnd 0.006281f
C2947 vdd.n739 gnd 0.495587f
C2948 vdd.n740 gnd 0.006281f
C2949 vdd.n741 gnd 0.006281f
C2950 vdd.t174 gnd 0.235994f
C2951 vdd.t224 gnd 0.287913f
C2952 vdd.n742 gnd 0.006281f
C2953 vdd.n743 gnd 0.006281f
C2954 vdd.n744 gnd 0.006281f
C2955 vdd.t216 gnd 0.320952f
C2956 vdd.n745 gnd 0.006281f
C2957 vdd.n746 gnd 0.006281f
C2958 vdd.t213 gnd 0.320952f
C2959 vdd.n747 gnd 0.006281f
C2960 vdd.n748 gnd 0.006281f
C2961 vdd.n749 gnd 0.006281f
C2962 vdd.t198 gnd 0.320952f
C2963 vdd.n750 gnd 0.006281f
C2964 vdd.n751 gnd 0.006281f
C2965 vdd.t178 gnd 0.320952f
C2966 vdd.n752 gnd 0.006281f
C2967 vdd.n753 gnd 0.006281f
C2968 vdd.n754 gnd 0.006281f
C2969 vdd.n755 gnd 0.641903f
C2970 vdd.n756 gnd 0.006281f
C2971 vdd.n757 gnd 0.006281f
C2972 vdd.n758 gnd 0.443669f
C2973 vdd.n759 gnd 0.006281f
C2974 vdd.n760 gnd 0.006281f
C2975 vdd.n761 gnd 0.006281f
C2976 vdd.t179 gnd 0.320952f
C2977 vdd.n762 gnd 0.006281f
C2978 vdd.n763 gnd 0.006281f
C2979 vdd.n764 gnd 0.006281f
C2980 vdd.n765 gnd 0.006281f
C2981 vdd.n766 gnd 0.006281f
C2982 vdd.t206 gnd 0.320952f
C2983 vdd.n767 gnd 0.006281f
C2984 vdd.n768 gnd 0.006281f
C2985 vdd.t145 gnd 0.320952f
C2986 vdd.n769 gnd 0.006281f
C2987 vdd.n770 gnd 0.014477f
C2988 vdd.n771 gnd 0.014477f
C2989 vdd.t204 gnd 0.566385f
C2990 vdd.n772 gnd 0.013603f
C2991 vdd.n773 gnd 0.013603f
C2992 vdd.n774 gnd 0.358711f
C2993 vdd.n775 gnd 0.014477f
C2994 vdd.n776 gnd 0.006281f
C2995 vdd.n777 gnd 0.006281f
C2996 vdd.t220 gnd 0.566385f
C2997 vdd.n795 gnd 0.014477f
C2998 vdd.n813 gnd 0.013603f
C2999 vdd.n814 gnd 0.006281f
C3000 vdd.n815 gnd 0.013603f
C3001 vdd.t160 gnd 0.25382f
C3002 vdd.t159 gnd 0.259817f
C3003 vdd.t158 gnd 0.165704f
C3004 vdd.n816 gnd 0.089554f
C3005 vdd.n817 gnd 0.050798f
C3006 vdd.n818 gnd 0.0144f
C3007 vdd.n819 gnd 0.006281f
C3008 vdd.n820 gnd 0.358711f
C3009 vdd.n821 gnd 0.013603f
C3010 vdd.n822 gnd 0.006281f
C3011 vdd.n823 gnd 0.014477f
C3012 vdd.n824 gnd 0.006281f
C3013 vdd.t143 gnd 0.25382f
C3014 vdd.t142 gnd 0.259817f
C3015 vdd.t140 gnd 0.165704f
C3016 vdd.n825 gnd 0.089554f
C3017 vdd.n826 gnd 0.050798f
C3018 vdd.n827 gnd 0.008977f
C3019 vdd.n828 gnd 0.006281f
C3020 vdd.n829 gnd 0.006281f
C3021 vdd.t141 gnd 0.320952f
C3022 vdd.n830 gnd 0.006281f
C3023 vdd.t218 gnd 0.320952f
C3024 vdd.n831 gnd 0.006281f
C3025 vdd.n832 gnd 0.006281f
C3026 vdd.n833 gnd 0.006281f
C3027 vdd.n834 gnd 0.006281f
C3028 vdd.n835 gnd 0.006281f
C3029 vdd.n836 gnd 0.641903f
C3030 vdd.n837 gnd 0.006281f
C3031 vdd.n838 gnd 0.006281f
C3032 vdd.t192 gnd 0.320952f
C3033 vdd.n839 gnd 0.006281f
C3034 vdd.n840 gnd 0.006281f
C3035 vdd.n841 gnd 0.006281f
C3036 vdd.n842 gnd 0.006281f
C3037 vdd.n843 gnd 0.443669f
C3038 vdd.n844 gnd 0.006281f
C3039 vdd.n845 gnd 0.006281f
C3040 vdd.n846 gnd 0.006281f
C3041 vdd.n847 gnd 0.006281f
C3042 vdd.n848 gnd 0.006281f
C3043 vdd.t175 gnd 0.320952f
C3044 vdd.n849 gnd 0.006281f
C3045 vdd.n850 gnd 0.006281f
C3046 vdd.t209 gnd 0.320952f
C3047 vdd.n851 gnd 0.006281f
C3048 vdd.n852 gnd 0.006281f
C3049 vdd.n853 gnd 0.006281f
C3050 vdd.t197 gnd 0.320952f
C3051 vdd.n854 gnd 0.006281f
C3052 vdd.n855 gnd 0.006281f
C3053 vdd.t176 gnd 0.320952f
C3054 vdd.n856 gnd 0.006281f
C3055 vdd.n857 gnd 0.006281f
C3056 vdd.n858 gnd 0.006281f
C3057 vdd.t195 gnd 0.287913f
C3058 vdd.n859 gnd 0.006281f
C3059 vdd.n860 gnd 0.006281f
C3060 vdd.n861 gnd 0.495587f
C3061 vdd.n862 gnd 0.006281f
C3062 vdd.n863 gnd 0.006281f
C3063 vdd.n864 gnd 0.006281f
C3064 vdd.t214 gnd 0.320952f
C3065 vdd.n865 gnd 0.006281f
C3066 vdd.n866 gnd 0.006281f
C3067 vdd.t184 gnd 0.235994f
C3068 vdd.n867 gnd 0.353991f
C3069 vdd.n868 gnd 0.006281f
C3070 vdd.n869 gnd 0.006281f
C3071 vdd.n870 gnd 0.006281f
C3072 vdd.n871 gnd 0.571105f
C3073 vdd.n872 gnd 0.006281f
C3074 vdd.n873 gnd 0.006281f
C3075 vdd.t222 gnd 0.320952f
C3076 vdd.n874 gnd 0.006281f
C3077 vdd.n875 gnd 0.006281f
C3078 vdd.n876 gnd 0.006281f
C3079 vdd.n877 gnd 0.641903f
C3080 vdd.n878 gnd 0.006281f
C3081 vdd.n879 gnd 0.006281f
C3082 vdd.t189 gnd 0.320952f
C3083 vdd.n880 gnd 0.006281f
C3084 vdd.n881 gnd 0.006281f
C3085 vdd.n882 gnd 0.006281f
C3086 vdd.t182 gnd 0.113277f
C3087 vdd.n883 gnd 0.006281f
C3088 vdd.n884 gnd 0.006281f
C3089 vdd.n885 gnd 0.006281f
C3090 vdd.t153 gnd 0.259817f
C3091 vdd.t151 gnd 0.165704f
C3092 vdd.t154 gnd 0.259817f
C3093 vdd.n886 gnd 0.146028f
C3094 vdd.n887 gnd 0.006281f
C3095 vdd.n888 gnd 0.006281f
C3096 vdd.t203 gnd 0.320952f
C3097 vdd.n889 gnd 0.006281f
C3098 vdd.n890 gnd 0.006281f
C3099 vdd.t152 gnd 0.250154f
C3100 vdd.n891 gnd 0.528626f
C3101 vdd.n892 gnd 0.006281f
C3102 vdd.n893 gnd 0.006281f
C3103 vdd.n894 gnd 0.006281f
C3104 vdd.n895 gnd 0.353991f
C3105 vdd.n896 gnd 0.006281f
C3106 vdd.n897 gnd 0.006281f
C3107 vdd.n898 gnd 0.429509f
C3108 vdd.n899 gnd 0.006281f
C3109 vdd.n900 gnd 0.006281f
C3110 vdd.n901 gnd 0.006281f
C3111 vdd.n902 gnd 0.495587f
C3112 vdd.n903 gnd 0.006281f
C3113 vdd.n904 gnd 0.006281f
C3114 vdd.t186 gnd 0.320952f
C3115 vdd.n905 gnd 0.006281f
C3116 vdd.n906 gnd 0.006281f
C3117 vdd.n907 gnd 0.006281f
C3118 vdd.n908 gnd 0.637184f
C3119 vdd.n909 gnd 0.006281f
C3120 vdd.n910 gnd 0.006281f
C3121 vdd.t185 gnd 0.320952f
C3122 vdd.n911 gnd 0.006281f
C3123 vdd.n912 gnd 0.006281f
C3124 vdd.n913 gnd 0.006281f
C3125 vdd.n914 gnd 0.641903f
C3126 vdd.n915 gnd 0.006281f
C3127 vdd.n916 gnd 0.006281f
C3128 vdd.t223 gnd 0.320952f
C3129 vdd.n917 gnd 0.006281f
C3130 vdd.n918 gnd 0.006281f
C3131 vdd.n919 gnd 0.006281f
C3132 vdd.n920 gnd 0.641903f
C3133 vdd.n921 gnd 0.006281f
C3134 vdd.n922 gnd 0.006281f
C3135 vdd.n923 gnd 0.006281f
C3136 vdd.n924 gnd 0.006281f
C3137 vdd.n925 gnd 0.006281f
C3138 vdd.n926 gnd 0.523906f
C3139 vdd.n927 gnd 0.006281f
C3140 vdd.n928 gnd 0.006281f
C3141 vdd.n929 gnd 0.006281f
C3142 vdd.n930 gnd 0.006281f
C3143 vdd.n931 gnd 0.006281f
C3144 vdd.n932 gnd 0.641903f
C3145 vdd.n933 gnd 0.006281f
C3146 vdd.n934 gnd 0.006281f
C3147 vdd.t103 gnd 0.320952f
C3148 vdd.n935 gnd 0.006281f
C3149 vdd.n936 gnd 0.014477f
C3150 vdd.n937 gnd 0.014477f
C3151 vdd.n938 gnd 9.600231f
C3152 vdd.n939 gnd 0.013603f
C3153 vdd.n940 gnd 0.013603f
C3154 vdd.n941 gnd 0.014477f
C3155 vdd.n942 gnd 0.006281f
C3156 vdd.n944 gnd 0.006281f
C3157 vdd.n945 gnd 0.006281f
C3158 vdd.n946 gnd 0.006281f
C3159 vdd.n947 gnd 0.006281f
C3160 vdd.n948 gnd 0.006281f
C3161 vdd.n949 gnd 0.006281f
C3162 vdd.n950 gnd 0.033049f
C3163 vdd.n951 gnd 0.006281f
C3164 vdd.n952 gnd 0.006281f
C3165 vdd.n953 gnd 0.006281f
C3166 vdd.n954 gnd 0.006281f
C3167 vdd.n955 gnd 0.006281f
C3168 vdd.n956 gnd 0.006281f
C3169 vdd.n957 gnd 0.006281f
C3170 vdd.t165 gnd 0.25382f
C3171 vdd.t166 gnd 0.259817f
C3172 vdd.t164 gnd 0.165704f
C3173 vdd.n958 gnd 0.089554f
C3174 vdd.n959 gnd 0.050798f
C3175 vdd.n960 gnd 0.006281f
C3176 vdd.n961 gnd 0.006281f
C3177 vdd.n962 gnd 0.006281f
C3178 vdd.n963 gnd 0.006281f
C3179 vdd.t104 gnd 0.25382f
C3180 vdd.t105 gnd 0.259817f
C3181 vdd.t102 gnd 0.165704f
C3182 vdd.n964 gnd 0.089554f
C3183 vdd.n965 gnd 0.050798f
C3184 vdd.n966 gnd 0.006281f
C3185 vdd.n967 gnd 0.006281f
C3186 vdd.n968 gnd 0.006281f
C3187 vdd.n969 gnd 0.006281f
C3188 vdd.n970 gnd 0.006281f
C3189 vdd.n971 gnd 0.006281f
C3190 vdd.n972 gnd 0.005912f
C3191 vdd.n975 gnd 0.022108f
C3192 vdd.n976 gnd 0.007435f
C3193 vdd.n977 gnd 0.009237f
C3194 vdd.n979 gnd 0.009237f
C3195 vdd.n980 gnd 0.006171f
C3196 vdd.t117 gnd 0.471988f
C3197 vdd.n981 gnd 9.892871f
C3198 vdd.n982 gnd 0.009237f
C3199 vdd.n983 gnd 0.022108f
C3200 vdd.n984 gnd 0.007435f
C3201 vdd.n985 gnd 0.009237f
C3202 vdd.n986 gnd 0.007435f
C3203 vdd.n987 gnd 0.009237f
C3204 vdd.n988 gnd 0.943976f
C3205 vdd.n989 gnd 0.009237f
C3206 vdd.n990 gnd 0.007435f
C3207 vdd.n991 gnd 0.007435f
C3208 vdd.n992 gnd 0.009237f
C3209 vdd.n993 gnd 0.007435f
C3210 vdd.n994 gnd 0.009237f
C3211 vdd.t4 gnd 0.471988f
C3212 vdd.n995 gnd 0.009237f
C3213 vdd.n996 gnd 0.007435f
C3214 vdd.n997 gnd 0.009237f
C3215 vdd.n998 gnd 0.007435f
C3216 vdd.n999 gnd 0.009237f
C3217 vdd.t29 gnd 0.471988f
C3218 vdd.n1000 gnd 0.009237f
C3219 vdd.n1001 gnd 0.007435f
C3220 vdd.n1002 gnd 0.009237f
C3221 vdd.n1003 gnd 0.007435f
C3222 vdd.n1004 gnd 0.009237f
C3223 vdd.t16 gnd 0.471988f
C3224 vdd.n1005 gnd 0.741021f
C3225 vdd.n1006 gnd 0.009237f
C3226 vdd.n1007 gnd 0.007435f
C3227 vdd.n1008 gnd 0.009237f
C3228 vdd.n1009 gnd 0.007435f
C3229 vdd.n1010 gnd 0.009237f
C3230 vdd.n1011 gnd 0.665503f
C3231 vdd.n1012 gnd 0.009237f
C3232 vdd.n1013 gnd 0.007435f
C3233 vdd.n1014 gnd 0.009237f
C3234 vdd.n1015 gnd 0.007435f
C3235 vdd.n1016 gnd 0.009237f
C3236 vdd.n1017 gnd 0.505027f
C3237 vdd.t12 gnd 0.471988f
C3238 vdd.n1018 gnd 0.009237f
C3239 vdd.n1019 gnd 0.007435f
C3240 vdd.n1020 gnd 0.009205f
C3241 vdd.n1021 gnd 0.007435f
C3242 vdd.n1022 gnd 0.009237f
C3243 vdd.t49 gnd 0.471988f
C3244 vdd.n1023 gnd 0.009237f
C3245 vdd.n1024 gnd 0.007435f
C3246 vdd.n1025 gnd 0.009237f
C3247 vdd.n1026 gnd 0.007435f
C3248 vdd.n1027 gnd 0.009237f
C3249 vdd.t62 gnd 0.471988f
C3250 vdd.n1028 gnd 0.599425f
C3251 vdd.n1029 gnd 0.009237f
C3252 vdd.n1030 gnd 0.007435f
C3253 vdd.n1031 gnd 0.009237f
C3254 vdd.n1032 gnd 0.007435f
C3255 vdd.n1033 gnd 0.009237f
C3256 vdd.t23 gnd 0.471988f
C3257 vdd.n1034 gnd 0.009237f
C3258 vdd.n1035 gnd 0.007435f
C3259 vdd.n1036 gnd 0.009237f
C3260 vdd.n1037 gnd 0.007435f
C3261 vdd.n1038 gnd 0.009237f
C3262 vdd.n1039 gnd 0.646623f
C3263 vdd.n1040 gnd 0.7835f
C3264 vdd.t51 gnd 0.471988f
C3265 vdd.n1041 gnd 0.009237f
C3266 vdd.n1042 gnd 0.007435f
C3267 vdd.n1043 gnd 0.009237f
C3268 vdd.n1044 gnd 0.007435f
C3269 vdd.n1045 gnd 0.009237f
C3270 vdd.n1046 gnd 0.486147f
C3271 vdd.n1047 gnd 0.009237f
C3272 vdd.n1048 gnd 0.007435f
C3273 vdd.n1049 gnd 0.009237f
C3274 vdd.n1050 gnd 0.007435f
C3275 vdd.n1051 gnd 0.009237f
C3276 vdd.n1052 gnd 0.943976f
C3277 vdd.t31 gnd 0.471988f
C3278 vdd.n1053 gnd 0.009237f
C3279 vdd.n1054 gnd 0.007435f
C3280 vdd.n1055 gnd 0.009237f
C3281 vdd.n1056 gnd 0.007435f
C3282 vdd.n1057 gnd 0.009237f
C3283 vdd.t121 gnd 0.471988f
C3284 vdd.n1058 gnd 0.009237f
C3285 vdd.n1059 gnd 0.007435f
C3286 vdd.n1060 gnd 0.022108f
C3287 vdd.n1061 gnd 0.022108f
C3288 vdd.n1062 gnd 2.17114f
C3289 vdd.n1063 gnd 0.533346f
C3290 vdd.n1064 gnd 0.022108f
C3291 vdd.n1065 gnd 0.009237f
C3292 vdd.n1067 gnd 0.009237f
C3293 vdd.n1068 gnd 0.009237f
C3294 vdd.n1069 gnd 0.007435f
C3295 vdd.n1070 gnd 0.009237f
C3296 vdd.n1071 gnd 0.009237f
C3297 vdd.n1073 gnd 0.009237f
C3298 vdd.n1074 gnd 0.009237f
C3299 vdd.n1076 gnd 0.009237f
C3300 vdd.n1077 gnd 0.007435f
C3301 vdd.n1078 gnd 0.009237f
C3302 vdd.n1079 gnd 0.009237f
C3303 vdd.n1081 gnd 0.009237f
C3304 vdd.n1082 gnd 0.009237f
C3305 vdd.n1084 gnd 0.009237f
C3306 vdd.n1085 gnd 0.007435f
C3307 vdd.n1086 gnd 0.009237f
C3308 vdd.n1087 gnd 0.009237f
C3309 vdd.n1089 gnd 0.009237f
C3310 vdd.n1090 gnd 0.009237f
C3311 vdd.n1092 gnd 0.009237f
C3312 vdd.n1093 gnd 0.007435f
C3313 vdd.n1094 gnd 0.009237f
C3314 vdd.n1095 gnd 0.009237f
C3315 vdd.n1097 gnd 0.009237f
C3316 vdd.n1098 gnd 0.009237f
C3317 vdd.n1100 gnd 0.009237f
C3318 vdd.t132 gnd 0.113639f
C3319 vdd.t133 gnd 0.121449f
C3320 vdd.t131 gnd 0.148411f
C3321 vdd.n1101 gnd 0.190242f
C3322 vdd.n1102 gnd 0.160581f
C3323 vdd.n1103 gnd 0.01591f
C3324 vdd.n1104 gnd 0.009237f
C3325 vdd.n1105 gnd 0.009237f
C3326 vdd.n1107 gnd 0.009237f
C3327 vdd.n1108 gnd 0.009237f
C3328 vdd.n1110 gnd 0.009237f
C3329 vdd.n1111 gnd 0.007435f
C3330 vdd.n1112 gnd 0.009237f
C3331 vdd.n1113 gnd 0.009237f
C3332 vdd.n1115 gnd 0.009237f
C3333 vdd.n1116 gnd 0.009237f
C3334 vdd.n1118 gnd 0.009237f
C3335 vdd.n1119 gnd 0.007435f
C3336 vdd.n1120 gnd 0.009237f
C3337 vdd.n1121 gnd 0.009237f
C3338 vdd.n1123 gnd 0.009237f
C3339 vdd.n1124 gnd 0.009237f
C3340 vdd.n1126 gnd 0.009237f
C3341 vdd.n1127 gnd 0.007435f
C3342 vdd.n1128 gnd 0.009237f
C3343 vdd.n1129 gnd 0.009237f
C3344 vdd.n1131 gnd 0.009237f
C3345 vdd.n1132 gnd 0.009237f
C3346 vdd.n1134 gnd 0.009237f
C3347 vdd.n1135 gnd 0.007435f
C3348 vdd.n1136 gnd 0.009237f
C3349 vdd.n1137 gnd 0.009237f
C3350 vdd.n1139 gnd 0.009237f
C3351 vdd.n1140 gnd 0.009237f
C3352 vdd.n1142 gnd 0.009237f
C3353 vdd.n1143 gnd 0.007435f
C3354 vdd.n1144 gnd 0.009237f
C3355 vdd.n1145 gnd 0.009237f
C3356 vdd.n1147 gnd 0.009237f
C3357 vdd.n1148 gnd 0.00736f
C3358 vdd.n1150 gnd 0.007435f
C3359 vdd.n1151 gnd 0.009237f
C3360 vdd.n1152 gnd 0.009237f
C3361 vdd.n1153 gnd 0.009237f
C3362 vdd.n1154 gnd 0.009237f
C3363 vdd.n1156 gnd 0.009237f
C3364 vdd.n1157 gnd 0.009237f
C3365 vdd.n1158 gnd 0.007435f
C3366 vdd.n1159 gnd 0.009237f
C3367 vdd.n1161 gnd 0.009237f
C3368 vdd.n1162 gnd 0.009237f
C3369 vdd.n1164 gnd 0.009237f
C3370 vdd.n1165 gnd 0.009237f
C3371 vdd.n1166 gnd 0.007435f
C3372 vdd.n1167 gnd 0.009237f
C3373 vdd.n1169 gnd 0.009237f
C3374 vdd.n1170 gnd 0.009237f
C3375 vdd.n1172 gnd 0.009237f
C3376 vdd.n1173 gnd 0.009237f
C3377 vdd.n1174 gnd 0.007435f
C3378 vdd.n1175 gnd 0.009237f
C3379 vdd.n1177 gnd 0.009237f
C3380 vdd.n1178 gnd 0.009237f
C3381 vdd.n1180 gnd 0.009237f
C3382 vdd.n1181 gnd 0.009237f
C3383 vdd.n1182 gnd 0.007435f
C3384 vdd.n1183 gnd 0.009237f
C3385 vdd.n1185 gnd 0.009237f
C3386 vdd.n1186 gnd 0.009237f
C3387 vdd.n1188 gnd 0.009237f
C3388 vdd.n1189 gnd 0.003531f
C3389 vdd.t129 gnd 0.113639f
C3390 vdd.t130 gnd 0.121449f
C3391 vdd.t128 gnd 0.148411f
C3392 vdd.n1190 gnd 0.190242f
C3393 vdd.n1191 gnd 0.160581f
C3394 vdd.n1192 gnd 0.012193f
C3395 vdd.n1193 gnd 0.003903f
C3396 vdd.n1194 gnd 0.007435f
C3397 vdd.n1195 gnd 0.009237f
C3398 vdd.n1196 gnd 0.009237f
C3399 vdd.n1197 gnd 0.009237f
C3400 vdd.n1198 gnd 0.007435f
C3401 vdd.n1199 gnd 0.007435f
C3402 vdd.n1200 gnd 0.007435f
C3403 vdd.n1201 gnd 0.009237f
C3404 vdd.n1202 gnd 0.009237f
C3405 vdd.n1203 gnd 0.009237f
C3406 vdd.n1204 gnd 0.007435f
C3407 vdd.n1205 gnd 0.007435f
C3408 vdd.n1206 gnd 0.007435f
C3409 vdd.n1207 gnd 0.009237f
C3410 vdd.n1208 gnd 0.009237f
C3411 vdd.n1209 gnd 0.009237f
C3412 vdd.n1210 gnd 0.007435f
C3413 vdd.n1211 gnd 0.007435f
C3414 vdd.n1212 gnd 0.007435f
C3415 vdd.n1213 gnd 0.009237f
C3416 vdd.n1214 gnd 0.009237f
C3417 vdd.n1215 gnd 0.009237f
C3418 vdd.n1216 gnd 0.007435f
C3419 vdd.n1217 gnd 0.007435f
C3420 vdd.n1218 gnd 0.007435f
C3421 vdd.n1219 gnd 0.009237f
C3422 vdd.n1220 gnd 0.009237f
C3423 vdd.n1221 gnd 0.009237f
C3424 vdd.n1222 gnd 0.007435f
C3425 vdd.n1223 gnd 0.009237f
C3426 vdd.n1224 gnd 0.009237f
C3427 vdd.n1226 gnd 0.009237f
C3428 vdd.t122 gnd 0.113639f
C3429 vdd.t123 gnd 0.121449f
C3430 vdd.t120 gnd 0.148411f
C3431 vdd.n1227 gnd 0.190242f
C3432 vdd.n1228 gnd 0.160581f
C3433 vdd.n1229 gnd 0.01591f
C3434 vdd.n1230 gnd 0.005056f
C3435 vdd.n1231 gnd 0.009237f
C3436 vdd.n1232 gnd 0.009237f
C3437 vdd.n1233 gnd 0.009237f
C3438 vdd.n1234 gnd 0.007435f
C3439 vdd.n1235 gnd 0.007435f
C3440 vdd.n1236 gnd 0.007435f
C3441 vdd.n1237 gnd 0.009237f
C3442 vdd.n1238 gnd 0.009237f
C3443 vdd.n1239 gnd 0.009237f
C3444 vdd.n1240 gnd 0.007435f
C3445 vdd.n1241 gnd 0.007435f
C3446 vdd.n1242 gnd 0.007435f
C3447 vdd.n1243 gnd 0.009237f
C3448 vdd.n1244 gnd 0.009237f
C3449 vdd.n1245 gnd 0.009237f
C3450 vdd.n1246 gnd 0.007435f
C3451 vdd.n1247 gnd 0.007435f
C3452 vdd.n1248 gnd 0.007435f
C3453 vdd.n1249 gnd 0.009237f
C3454 vdd.n1250 gnd 0.009237f
C3455 vdd.n1251 gnd 0.009237f
C3456 vdd.n1252 gnd 0.007435f
C3457 vdd.n1253 gnd 0.007435f
C3458 vdd.n1254 gnd 0.007435f
C3459 vdd.n1255 gnd 0.009237f
C3460 vdd.n1256 gnd 0.009237f
C3461 vdd.n1257 gnd 0.009237f
C3462 vdd.n1258 gnd 0.007435f
C3463 vdd.n1259 gnd 0.007435f
C3464 vdd.n1260 gnd 0.006208f
C3465 vdd.n1261 gnd 0.009237f
C3466 vdd.n1262 gnd 0.009237f
C3467 vdd.n1263 gnd 0.009237f
C3468 vdd.n1264 gnd 0.006208f
C3469 vdd.n1265 gnd 0.007435f
C3470 vdd.n1266 gnd 0.007435f
C3471 vdd.n1267 gnd 0.009237f
C3472 vdd.n1268 gnd 0.009237f
C3473 vdd.n1269 gnd 0.009237f
C3474 vdd.n1270 gnd 0.007435f
C3475 vdd.n1271 gnd 0.007435f
C3476 vdd.n1272 gnd 0.007435f
C3477 vdd.n1273 gnd 0.009237f
C3478 vdd.n1274 gnd 0.009237f
C3479 vdd.n1275 gnd 0.009237f
C3480 vdd.n1276 gnd 0.007435f
C3481 vdd.n1277 gnd 0.007435f
C3482 vdd.n1278 gnd 0.007435f
C3483 vdd.n1279 gnd 0.009237f
C3484 vdd.n1280 gnd 0.009237f
C3485 vdd.n1281 gnd 0.009237f
C3486 vdd.n1282 gnd 0.007435f
C3487 vdd.n1283 gnd 0.007435f
C3488 vdd.n1284 gnd 0.007435f
C3489 vdd.n1285 gnd 0.009237f
C3490 vdd.n1286 gnd 0.009237f
C3491 vdd.n1287 gnd 0.009237f
C3492 vdd.n1288 gnd 0.007435f
C3493 vdd.n1289 gnd 0.007435f
C3494 vdd.n1290 gnd 0.006171f
C3495 vdd.n1291 gnd 0.022108f
C3496 vdd.n1292 gnd 0.021768f
C3497 vdd.n1293 gnd 0.006171f
C3498 vdd.n1294 gnd 0.021768f
C3499 vdd.n1295 gnd 1.33101f
C3500 vdd.n1296 gnd 0.021768f
C3501 vdd.n1297 gnd 0.006171f
C3502 vdd.n1298 gnd 0.021768f
C3503 vdd.n1299 gnd 0.009237f
C3504 vdd.n1300 gnd 0.009237f
C3505 vdd.n1301 gnd 0.007435f
C3506 vdd.n1302 gnd 0.009237f
C3507 vdd.n1303 gnd 0.882617f
C3508 vdd.n1304 gnd 0.009237f
C3509 vdd.n1305 gnd 0.007435f
C3510 vdd.n1306 gnd 0.009237f
C3511 vdd.n1307 gnd 0.009237f
C3512 vdd.n1308 gnd 0.009237f
C3513 vdd.n1309 gnd 0.007435f
C3514 vdd.n1310 gnd 0.009237f
C3515 vdd.n1311 gnd 0.929816f
C3516 vdd.n1312 gnd 0.009237f
C3517 vdd.n1313 gnd 0.007435f
C3518 vdd.n1314 gnd 0.009237f
C3519 vdd.n1315 gnd 0.009237f
C3520 vdd.n1316 gnd 0.009237f
C3521 vdd.n1317 gnd 0.007435f
C3522 vdd.n1318 gnd 0.009237f
C3523 vdd.t25 gnd 0.471988f
C3524 vdd.n1319 gnd 0.76934f
C3525 vdd.n1320 gnd 0.009237f
C3526 vdd.n1321 gnd 0.007435f
C3527 vdd.n1322 gnd 0.009237f
C3528 vdd.n1323 gnd 0.009237f
C3529 vdd.n1324 gnd 0.009237f
C3530 vdd.n1325 gnd 0.007435f
C3531 vdd.n1326 gnd 0.009237f
C3532 vdd.n1327 gnd 0.608864f
C3533 vdd.n1328 gnd 0.009237f
C3534 vdd.n1329 gnd 0.007435f
C3535 vdd.n1330 gnd 0.009237f
C3536 vdd.n1331 gnd 0.009237f
C3537 vdd.n1332 gnd 0.009237f
C3538 vdd.n1333 gnd 0.007435f
C3539 vdd.n1334 gnd 0.009237f
C3540 vdd.n1335 gnd 0.7599f
C3541 vdd.n1336 gnd 0.495587f
C3542 vdd.n1337 gnd 0.009237f
C3543 vdd.n1338 gnd 0.007435f
C3544 vdd.n1339 gnd 0.009237f
C3545 vdd.n1340 gnd 0.009237f
C3546 vdd.n1341 gnd 0.009237f
C3547 vdd.n1342 gnd 0.007435f
C3548 vdd.n1343 gnd 0.009237f
C3549 vdd.n1344 gnd 0.656063f
C3550 vdd.n1345 gnd 0.009237f
C3551 vdd.n1346 gnd 0.007435f
C3552 vdd.n1347 gnd 0.009237f
C3553 vdd.n1348 gnd 0.009237f
C3554 vdd.n1349 gnd 0.009237f
C3555 vdd.n1350 gnd 0.007435f
C3556 vdd.n1351 gnd 0.009237f
C3557 vdd.t6 gnd 0.471988f
C3558 vdd.n1352 gnd 0.7835f
C3559 vdd.n1353 gnd 0.009237f
C3560 vdd.n1354 gnd 0.007435f
C3561 vdd.n1355 gnd 0.005069f
C3562 vdd.n1356 gnd 0.004704f
C3563 vdd.n1357 gnd 0.002602f
C3564 vdd.n1358 gnd 0.005975f
C3565 vdd.n1359 gnd 0.002528f
C3566 vdd.n1360 gnd 0.002676f
C3567 vdd.n1361 gnd 0.004704f
C3568 vdd.n1362 gnd 0.002528f
C3569 vdd.n1363 gnd 0.005975f
C3570 vdd.n1364 gnd 0.002676f
C3571 vdd.n1365 gnd 0.004704f
C3572 vdd.n1366 gnd 0.002528f
C3573 vdd.n1367 gnd 0.004481f
C3574 vdd.n1368 gnd 0.004494f
C3575 vdd.t236 gnd 0.012836f
C3576 vdd.n1369 gnd 0.02856f
C3577 vdd.n1370 gnd 0.148635f
C3578 vdd.n1371 gnd 0.002528f
C3579 vdd.n1372 gnd 0.002676f
C3580 vdd.n1373 gnd 0.005975f
C3581 vdd.n1374 gnd 0.005975f
C3582 vdd.n1375 gnd 0.002676f
C3583 vdd.n1376 gnd 0.002528f
C3584 vdd.n1377 gnd 0.004704f
C3585 vdd.n1378 gnd 0.004704f
C3586 vdd.n1379 gnd 0.002528f
C3587 vdd.n1380 gnd 0.002676f
C3588 vdd.n1381 gnd 0.005975f
C3589 vdd.n1382 gnd 0.005975f
C3590 vdd.n1383 gnd 0.002676f
C3591 vdd.n1384 gnd 0.002528f
C3592 vdd.n1385 gnd 0.004704f
C3593 vdd.n1386 gnd 0.004704f
C3594 vdd.n1387 gnd 0.002528f
C3595 vdd.n1388 gnd 0.002676f
C3596 vdd.n1389 gnd 0.005975f
C3597 vdd.n1390 gnd 0.005975f
C3598 vdd.n1391 gnd 0.014125f
C3599 vdd.n1392 gnd 0.002602f
C3600 vdd.n1393 gnd 0.002528f
C3601 vdd.n1394 gnd 0.012159f
C3602 vdd.n1395 gnd 0.008488f
C3603 vdd.t230 gnd 0.029739f
C3604 vdd.t59 gnd 0.029739f
C3605 vdd.n1396 gnd 0.204384f
C3606 vdd.n1397 gnd 0.160717f
C3607 vdd.t20 gnd 0.029739f
C3608 vdd.t170 gnd 0.029739f
C3609 vdd.n1398 gnd 0.204384f
C3610 vdd.n1399 gnd 0.129698f
C3611 vdd.t84 gnd 0.029739f
C3612 vdd.t7 gnd 0.029739f
C3613 vdd.n1400 gnd 0.204384f
C3614 vdd.n1401 gnd 0.129698f
C3615 vdd.t24 gnd 0.029739f
C3616 vdd.t63 gnd 0.029739f
C3617 vdd.n1402 gnd 0.204384f
C3618 vdd.n1403 gnd 0.129698f
C3619 vdd.t233 gnd 0.029739f
C3620 vdd.t80 gnd 0.029739f
C3621 vdd.n1404 gnd 0.204384f
C3622 vdd.n1405 gnd 0.129698f
C3623 vdd.n1406 gnd 0.005069f
C3624 vdd.n1407 gnd 0.004704f
C3625 vdd.n1408 gnd 0.002602f
C3626 vdd.n1409 gnd 0.005975f
C3627 vdd.n1410 gnd 0.002528f
C3628 vdd.n1411 gnd 0.002676f
C3629 vdd.n1412 gnd 0.004704f
C3630 vdd.n1413 gnd 0.002528f
C3631 vdd.n1414 gnd 0.005975f
C3632 vdd.n1415 gnd 0.002676f
C3633 vdd.n1416 gnd 0.004704f
C3634 vdd.n1417 gnd 0.002528f
C3635 vdd.n1418 gnd 0.004481f
C3636 vdd.n1419 gnd 0.004494f
C3637 vdd.t32 gnd 0.012836f
C3638 vdd.n1420 gnd 0.02856f
C3639 vdd.n1421 gnd 0.148635f
C3640 vdd.n1422 gnd 0.002528f
C3641 vdd.n1423 gnd 0.002676f
C3642 vdd.n1424 gnd 0.005975f
C3643 vdd.n1425 gnd 0.005975f
C3644 vdd.n1426 gnd 0.002676f
C3645 vdd.n1427 gnd 0.002528f
C3646 vdd.n1428 gnd 0.004704f
C3647 vdd.n1429 gnd 0.004704f
C3648 vdd.n1430 gnd 0.002528f
C3649 vdd.n1431 gnd 0.002676f
C3650 vdd.n1432 gnd 0.005975f
C3651 vdd.n1433 gnd 0.005975f
C3652 vdd.n1434 gnd 0.002676f
C3653 vdd.n1435 gnd 0.002528f
C3654 vdd.n1436 gnd 0.004704f
C3655 vdd.n1437 gnd 0.004704f
C3656 vdd.n1438 gnd 0.002528f
C3657 vdd.n1439 gnd 0.002676f
C3658 vdd.n1440 gnd 0.005975f
C3659 vdd.n1441 gnd 0.005975f
C3660 vdd.n1442 gnd 0.014125f
C3661 vdd.n1443 gnd 0.002602f
C3662 vdd.n1444 gnd 0.002528f
C3663 vdd.n1445 gnd 0.012159f
C3664 vdd.n1446 gnd 0.008222f
C3665 vdd.n1447 gnd 0.096496f
C3666 vdd.n1448 gnd 0.005069f
C3667 vdd.n1449 gnd 0.004704f
C3668 vdd.n1450 gnd 0.002602f
C3669 vdd.n1451 gnd 0.005975f
C3670 vdd.n1452 gnd 0.002528f
C3671 vdd.n1453 gnd 0.002676f
C3672 vdd.n1454 gnd 0.004704f
C3673 vdd.n1455 gnd 0.002528f
C3674 vdd.n1456 gnd 0.005975f
C3675 vdd.n1457 gnd 0.002676f
C3676 vdd.n1458 gnd 0.004704f
C3677 vdd.n1459 gnd 0.002528f
C3678 vdd.n1460 gnd 0.004481f
C3679 vdd.n1461 gnd 0.004494f
C3680 vdd.t75 gnd 0.012836f
C3681 vdd.n1462 gnd 0.02856f
C3682 vdd.n1463 gnd 0.148635f
C3683 vdd.n1464 gnd 0.002528f
C3684 vdd.n1465 gnd 0.002676f
C3685 vdd.n1466 gnd 0.005975f
C3686 vdd.n1467 gnd 0.005975f
C3687 vdd.n1468 gnd 0.002676f
C3688 vdd.n1469 gnd 0.002528f
C3689 vdd.n1470 gnd 0.004704f
C3690 vdd.n1471 gnd 0.004704f
C3691 vdd.n1472 gnd 0.002528f
C3692 vdd.n1473 gnd 0.002676f
C3693 vdd.n1474 gnd 0.005975f
C3694 vdd.n1475 gnd 0.005975f
C3695 vdd.n1476 gnd 0.002676f
C3696 vdd.n1477 gnd 0.002528f
C3697 vdd.n1478 gnd 0.004704f
C3698 vdd.n1479 gnd 0.004704f
C3699 vdd.n1480 gnd 0.002528f
C3700 vdd.n1481 gnd 0.002676f
C3701 vdd.n1482 gnd 0.005975f
C3702 vdd.n1483 gnd 0.005975f
C3703 vdd.n1484 gnd 0.014125f
C3704 vdd.n1485 gnd 0.002602f
C3705 vdd.n1486 gnd 0.002528f
C3706 vdd.n1487 gnd 0.012159f
C3707 vdd.n1488 gnd 0.008488f
C3708 vdd.t53 gnd 0.029739f
C3709 vdd.t239 gnd 0.029739f
C3710 vdd.n1489 gnd 0.204384f
C3711 vdd.n1490 gnd 0.160717f
C3712 vdd.t13 gnd 0.029739f
C3713 vdd.t48 gnd 0.029739f
C3714 vdd.n1491 gnd 0.204384f
C3715 vdd.n1492 gnd 0.129698f
C3716 vdd.t50 gnd 0.029739f
C3717 vdd.t237 gnd 0.029739f
C3718 vdd.n1493 gnd 0.204384f
C3719 vdd.n1494 gnd 0.129698f
C3720 vdd.t79 gnd 0.029739f
C3721 vdd.t226 gnd 0.029739f
C3722 vdd.n1495 gnd 0.204384f
C3723 vdd.n1496 gnd 0.129698f
C3724 vdd.t90 gnd 0.029739f
C3725 vdd.t52 gnd 0.029739f
C3726 vdd.n1497 gnd 0.204384f
C3727 vdd.n1498 gnd 0.129698f
C3728 vdd.n1499 gnd 0.005069f
C3729 vdd.n1500 gnd 0.004704f
C3730 vdd.n1501 gnd 0.002602f
C3731 vdd.n1502 gnd 0.005975f
C3732 vdd.n1503 gnd 0.002528f
C3733 vdd.n1504 gnd 0.002676f
C3734 vdd.n1505 gnd 0.004704f
C3735 vdd.n1506 gnd 0.002528f
C3736 vdd.n1507 gnd 0.005975f
C3737 vdd.n1508 gnd 0.002676f
C3738 vdd.n1509 gnd 0.004704f
C3739 vdd.n1510 gnd 0.002528f
C3740 vdd.n1511 gnd 0.004481f
C3741 vdd.n1512 gnd 0.004494f
C3742 vdd.t91 gnd 0.012836f
C3743 vdd.n1513 gnd 0.02856f
C3744 vdd.n1514 gnd 0.148635f
C3745 vdd.n1515 gnd 0.002528f
C3746 vdd.n1516 gnd 0.002676f
C3747 vdd.n1517 gnd 0.005975f
C3748 vdd.n1518 gnd 0.005975f
C3749 vdd.n1519 gnd 0.002676f
C3750 vdd.n1520 gnd 0.002528f
C3751 vdd.n1521 gnd 0.004704f
C3752 vdd.n1522 gnd 0.004704f
C3753 vdd.n1523 gnd 0.002528f
C3754 vdd.n1524 gnd 0.002676f
C3755 vdd.n1525 gnd 0.005975f
C3756 vdd.n1526 gnd 0.005975f
C3757 vdd.n1527 gnd 0.002676f
C3758 vdd.n1528 gnd 0.002528f
C3759 vdd.n1529 gnd 0.004704f
C3760 vdd.n1530 gnd 0.004704f
C3761 vdd.n1531 gnd 0.002528f
C3762 vdd.n1532 gnd 0.002676f
C3763 vdd.n1533 gnd 0.005975f
C3764 vdd.n1534 gnd 0.005975f
C3765 vdd.n1535 gnd 0.014125f
C3766 vdd.n1536 gnd 0.002602f
C3767 vdd.n1537 gnd 0.002528f
C3768 vdd.n1538 gnd 0.012159f
C3769 vdd.n1539 gnd 0.008222f
C3770 vdd.n1540 gnd 0.057405f
C3771 vdd.n1541 gnd 0.206846f
C3772 vdd.n1542 gnd 0.005069f
C3773 vdd.n1543 gnd 0.004704f
C3774 vdd.n1544 gnd 0.002602f
C3775 vdd.n1545 gnd 0.005975f
C3776 vdd.n1546 gnd 0.002528f
C3777 vdd.n1547 gnd 0.002676f
C3778 vdd.n1548 gnd 0.004704f
C3779 vdd.n1549 gnd 0.002528f
C3780 vdd.n1550 gnd 0.005975f
C3781 vdd.n1551 gnd 0.002676f
C3782 vdd.n1552 gnd 0.004704f
C3783 vdd.n1553 gnd 0.002528f
C3784 vdd.n1554 gnd 0.004481f
C3785 vdd.n1555 gnd 0.004494f
C3786 vdd.t5 gnd 0.012836f
C3787 vdd.n1556 gnd 0.02856f
C3788 vdd.n1557 gnd 0.148635f
C3789 vdd.n1558 gnd 0.002528f
C3790 vdd.n1559 gnd 0.002676f
C3791 vdd.n1560 gnd 0.005975f
C3792 vdd.n1561 gnd 0.005975f
C3793 vdd.n1562 gnd 0.002676f
C3794 vdd.n1563 gnd 0.002528f
C3795 vdd.n1564 gnd 0.004704f
C3796 vdd.n1565 gnd 0.004704f
C3797 vdd.n1566 gnd 0.002528f
C3798 vdd.n1567 gnd 0.002676f
C3799 vdd.n1568 gnd 0.005975f
C3800 vdd.n1569 gnd 0.005975f
C3801 vdd.n1570 gnd 0.002676f
C3802 vdd.n1571 gnd 0.002528f
C3803 vdd.n1572 gnd 0.004704f
C3804 vdd.n1573 gnd 0.004704f
C3805 vdd.n1574 gnd 0.002528f
C3806 vdd.n1575 gnd 0.002676f
C3807 vdd.n1576 gnd 0.005975f
C3808 vdd.n1577 gnd 0.005975f
C3809 vdd.n1578 gnd 0.014125f
C3810 vdd.n1579 gnd 0.002602f
C3811 vdd.n1580 gnd 0.002528f
C3812 vdd.n1581 gnd 0.012159f
C3813 vdd.n1582 gnd 0.008488f
C3814 vdd.t17 gnd 0.029739f
C3815 vdd.t30 gnd 0.029739f
C3816 vdd.n1583 gnd 0.204384f
C3817 vdd.n1584 gnd 0.160717f
C3818 vdd.t172 gnd 0.029739f
C3819 vdd.t73 gnd 0.029739f
C3820 vdd.n1585 gnd 0.204384f
C3821 vdd.n1586 gnd 0.129698f
C3822 vdd.t54 gnd 0.029739f
C3823 vdd.t55 gnd 0.029739f
C3824 vdd.n1587 gnd 0.204384f
C3825 vdd.n1588 gnd 0.129698f
C3826 vdd.t231 gnd 0.029739f
C3827 vdd.t86 gnd 0.029739f
C3828 vdd.n1589 gnd 0.204384f
C3829 vdd.n1590 gnd 0.129698f
C3830 vdd.t26 gnd 0.029739f
C3831 vdd.t56 gnd 0.029739f
C3832 vdd.n1591 gnd 0.204384f
C3833 vdd.n1592 gnd 0.129698f
C3834 vdd.n1593 gnd 0.005069f
C3835 vdd.n1594 gnd 0.004704f
C3836 vdd.n1595 gnd 0.002602f
C3837 vdd.n1596 gnd 0.005975f
C3838 vdd.n1597 gnd 0.002528f
C3839 vdd.n1598 gnd 0.002676f
C3840 vdd.n1599 gnd 0.004704f
C3841 vdd.n1600 gnd 0.002528f
C3842 vdd.n1601 gnd 0.005975f
C3843 vdd.n1602 gnd 0.002676f
C3844 vdd.n1603 gnd 0.004704f
C3845 vdd.n1604 gnd 0.002528f
C3846 vdd.n1605 gnd 0.004481f
C3847 vdd.n1606 gnd 0.004494f
C3848 vdd.t87 gnd 0.012836f
C3849 vdd.n1607 gnd 0.02856f
C3850 vdd.n1608 gnd 0.148635f
C3851 vdd.n1609 gnd 0.002528f
C3852 vdd.n1610 gnd 0.002676f
C3853 vdd.n1611 gnd 0.005975f
C3854 vdd.n1612 gnd 0.005975f
C3855 vdd.n1613 gnd 0.002676f
C3856 vdd.n1614 gnd 0.002528f
C3857 vdd.n1615 gnd 0.004704f
C3858 vdd.n1616 gnd 0.004704f
C3859 vdd.n1617 gnd 0.002528f
C3860 vdd.n1618 gnd 0.002676f
C3861 vdd.n1619 gnd 0.005975f
C3862 vdd.n1620 gnd 0.005975f
C3863 vdd.n1621 gnd 0.002676f
C3864 vdd.n1622 gnd 0.002528f
C3865 vdd.n1623 gnd 0.004704f
C3866 vdd.n1624 gnd 0.004704f
C3867 vdd.n1625 gnd 0.002528f
C3868 vdd.n1626 gnd 0.002676f
C3869 vdd.n1627 gnd 0.005975f
C3870 vdd.n1628 gnd 0.005975f
C3871 vdd.n1629 gnd 0.014125f
C3872 vdd.n1630 gnd 0.002602f
C3873 vdd.n1631 gnd 0.002528f
C3874 vdd.n1632 gnd 0.012159f
C3875 vdd.n1633 gnd 0.008222f
C3876 vdd.n1634 gnd 0.057405f
C3877 vdd.n1635 gnd 0.22733f
C3878 vdd.n1636 gnd 2.26913f
C3879 vdd.n1637 gnd 0.549857f
C3880 vdd.n1638 gnd 0.009205f
C3881 vdd.n1639 gnd 0.009237f
C3882 vdd.n1640 gnd 0.007435f
C3883 vdd.n1641 gnd 0.009237f
C3884 vdd.n1642 gnd 0.750461f
C3885 vdd.n1643 gnd 0.009237f
C3886 vdd.n1644 gnd 0.007435f
C3887 vdd.n1645 gnd 0.009237f
C3888 vdd.n1646 gnd 0.009237f
C3889 vdd.n1647 gnd 0.009237f
C3890 vdd.n1648 gnd 0.007435f
C3891 vdd.n1649 gnd 0.009237f
C3892 vdd.n1650 gnd 0.7835f
C3893 vdd.t47 gnd 0.471988f
C3894 vdd.n1651 gnd 0.589985f
C3895 vdd.n1652 gnd 0.009237f
C3896 vdd.n1653 gnd 0.007435f
C3897 vdd.n1654 gnd 0.009237f
C3898 vdd.n1655 gnd 0.009237f
C3899 vdd.n1656 gnd 0.009237f
C3900 vdd.n1657 gnd 0.007435f
C3901 vdd.n1658 gnd 0.009237f
C3902 vdd.n1659 gnd 0.514467f
C3903 vdd.n1660 gnd 0.009237f
C3904 vdd.n1661 gnd 0.007435f
C3905 vdd.n1662 gnd 0.009237f
C3906 vdd.n1663 gnd 0.009237f
C3907 vdd.n1664 gnd 0.009237f
C3908 vdd.n1665 gnd 0.007435f
C3909 vdd.n1666 gnd 0.009237f
C3910 vdd.n1667 gnd 0.580545f
C3911 vdd.n1668 gnd 0.674943f
C3912 vdd.n1669 gnd 0.009237f
C3913 vdd.n1670 gnd 0.007435f
C3914 vdd.n1671 gnd 0.009237f
C3915 vdd.n1672 gnd 0.009237f
C3916 vdd.n1673 gnd 0.009237f
C3917 vdd.n1674 gnd 0.007435f
C3918 vdd.n1675 gnd 0.009237f
C3919 vdd.n1676 gnd 0.835418f
C3920 vdd.n1677 gnd 0.009237f
C3921 vdd.n1678 gnd 0.007435f
C3922 vdd.n1679 gnd 0.009237f
C3923 vdd.n1680 gnd 0.009237f
C3924 vdd.n1681 gnd 0.021768f
C3925 vdd.n1682 gnd 0.009237f
C3926 vdd.n1683 gnd 0.009237f
C3927 vdd.n1684 gnd 0.007435f
C3928 vdd.n1685 gnd 0.009237f
C3929 vdd.n1686 gnd 0.505027f
C3930 vdd.n1687 gnd 0.943976f
C3931 vdd.n1688 gnd 0.009237f
C3932 vdd.n1689 gnd 0.007435f
C3933 vdd.n1690 gnd 0.009237f
C3934 vdd.n1691 gnd 0.009237f
C3935 vdd.n1692 gnd 0.007944f
C3936 vdd.n1693 gnd 0.007435f
C3937 vdd.n1695 gnd 0.009237f
C3938 vdd.n1697 gnd 0.007435f
C3939 vdd.n1698 gnd 0.009237f
C3940 vdd.n1699 gnd 0.007435f
C3941 vdd.n1701 gnd 0.009237f
C3942 vdd.n1702 gnd 0.007435f
C3943 vdd.n1703 gnd 0.009237f
C3944 vdd.n1704 gnd 0.009237f
C3945 vdd.n1705 gnd 0.009237f
C3946 vdd.n1706 gnd 0.009237f
C3947 vdd.n1707 gnd 0.009237f
C3948 vdd.n1708 gnd 0.007435f
C3949 vdd.n1710 gnd 0.009237f
C3950 vdd.n1711 gnd 0.009237f
C3951 vdd.n1712 gnd 0.009237f
C3952 vdd.n1713 gnd 0.009237f
C3953 vdd.n1714 gnd 0.009237f
C3954 vdd.n1715 gnd 0.007435f
C3955 vdd.n1717 gnd 0.009237f
C3956 vdd.n1718 gnd 0.009237f
C3957 vdd.n1719 gnd 0.009237f
C3958 vdd.n1720 gnd 0.009237f
C3959 vdd.n1721 gnd 0.006208f
C3960 vdd.t150 gnd 0.113639f
C3961 vdd.t149 gnd 0.121449f
C3962 vdd.t148 gnd 0.148411f
C3963 vdd.n1722 gnd 0.190242f
C3964 vdd.n1723 gnd 0.159838f
C3965 vdd.n1725 gnd 0.009237f
C3966 vdd.n1726 gnd 0.009237f
C3967 vdd.n1727 gnd 0.007435f
C3968 vdd.n1728 gnd 0.009237f
C3969 vdd.n1730 gnd 0.009237f
C3970 vdd.n1731 gnd 0.009237f
C3971 vdd.n1732 gnd 0.009237f
C3972 vdd.n1733 gnd 0.009237f
C3973 vdd.n1734 gnd 0.007435f
C3974 vdd.n1736 gnd 0.009237f
C3975 vdd.n1737 gnd 0.009237f
C3976 vdd.n1738 gnd 0.009237f
C3977 vdd.n1739 gnd 0.009237f
C3978 vdd.n1740 gnd 0.009237f
C3979 vdd.n1741 gnd 0.007435f
C3980 vdd.n1743 gnd 0.009237f
C3981 vdd.n1744 gnd 0.009237f
C3982 vdd.n1745 gnd 0.009237f
C3983 vdd.n1746 gnd 0.009237f
C3984 vdd.n1747 gnd 0.009237f
C3985 vdd.n1748 gnd 0.007435f
C3986 vdd.n1750 gnd 0.009237f
C3987 vdd.n1751 gnd 0.009237f
C3988 vdd.n1752 gnd 0.009237f
C3989 vdd.n1753 gnd 0.009237f
C3990 vdd.n1754 gnd 0.009237f
C3991 vdd.n1755 gnd 0.007435f
C3992 vdd.n1757 gnd 0.009237f
C3993 vdd.n1758 gnd 0.009237f
C3994 vdd.n1759 gnd 0.009237f
C3995 vdd.n1760 gnd 0.009237f
C3996 vdd.n1761 gnd 0.00736f
C3997 vdd.t139 gnd 0.113639f
C3998 vdd.t138 gnd 0.121449f
C3999 vdd.t137 gnd 0.148411f
C4000 vdd.n1762 gnd 0.190242f
C4001 vdd.n1763 gnd 0.159838f
C4002 vdd.n1765 gnd 0.009237f
C4003 vdd.n1766 gnd 0.009237f
C4004 vdd.n1767 gnd 0.007435f
C4005 vdd.n1768 gnd 0.009237f
C4006 vdd.n1770 gnd 0.009237f
C4007 vdd.n1771 gnd 0.009237f
C4008 vdd.n1772 gnd 0.009237f
C4009 vdd.n1773 gnd 0.009237f
C4010 vdd.n1774 gnd 0.007435f
C4011 vdd.n1776 gnd 0.009237f
C4012 vdd.n1777 gnd 0.009237f
C4013 vdd.n1778 gnd 0.009237f
C4014 vdd.n1779 gnd 0.009237f
C4015 vdd.n1780 gnd 0.009237f
C4016 vdd.n1781 gnd 0.007435f
C4017 vdd.n1783 gnd 0.009237f
C4018 vdd.n1784 gnd 0.009237f
C4019 vdd.n1785 gnd 0.009237f
C4020 vdd.n1786 gnd 0.009237f
C4021 vdd.n1787 gnd 0.009237f
C4022 vdd.n1788 gnd 0.009237f
C4023 vdd.n1789 gnd 0.007435f
C4024 vdd.n1791 gnd 0.009237f
C4025 vdd.n1793 gnd 0.009237f
C4026 vdd.n1794 gnd 0.007435f
C4027 vdd.n1795 gnd 0.007435f
C4028 vdd.n1796 gnd 0.009237f
C4029 vdd.n1798 gnd 0.009237f
C4030 vdd.n1799 gnd 0.007435f
C4031 vdd.n1800 gnd 0.007435f
C4032 vdd.n1801 gnd 0.009237f
C4033 vdd.n1803 gnd 0.009237f
C4034 vdd.n1804 gnd 0.009237f
C4035 vdd.n1805 gnd 0.007435f
C4036 vdd.n1806 gnd 0.007435f
C4037 vdd.n1807 gnd 0.007435f
C4038 vdd.n1808 gnd 0.009237f
C4039 vdd.n1810 gnd 0.009237f
C4040 vdd.n1811 gnd 0.009237f
C4041 vdd.n1812 gnd 0.007435f
C4042 vdd.n1813 gnd 0.007435f
C4043 vdd.n1814 gnd 0.007435f
C4044 vdd.n1815 gnd 0.009237f
C4045 vdd.n1817 gnd 0.009237f
C4046 vdd.n1818 gnd 0.009237f
C4047 vdd.n1819 gnd 0.007435f
C4048 vdd.n1820 gnd 0.007435f
C4049 vdd.n1821 gnd 0.007435f
C4050 vdd.n1822 gnd 0.009237f
C4051 vdd.n1824 gnd 0.009237f
C4052 vdd.n1825 gnd 0.009237f
C4053 vdd.n1826 gnd 0.007435f
C4054 vdd.n1827 gnd 0.009237f
C4055 vdd.n1828 gnd 0.009237f
C4056 vdd.n1829 gnd 0.009237f
C4057 vdd.n1830 gnd 0.015167f
C4058 vdd.n1831 gnd 0.005056f
C4059 vdd.n1832 gnd 0.007435f
C4060 vdd.n1833 gnd 0.009237f
C4061 vdd.n1835 gnd 0.009237f
C4062 vdd.n1836 gnd 0.009237f
C4063 vdd.n1837 gnd 0.007435f
C4064 vdd.n1838 gnd 0.007435f
C4065 vdd.n1839 gnd 0.007435f
C4066 vdd.n1840 gnd 0.009237f
C4067 vdd.n1842 gnd 0.009237f
C4068 vdd.n1843 gnd 0.009237f
C4069 vdd.n1844 gnd 0.007435f
C4070 vdd.n1845 gnd 0.007435f
C4071 vdd.n1846 gnd 0.007435f
C4072 vdd.n1847 gnd 0.009237f
C4073 vdd.n1849 gnd 0.009237f
C4074 vdd.n1850 gnd 0.009237f
C4075 vdd.n1851 gnd 0.007435f
C4076 vdd.n1852 gnd 0.007435f
C4077 vdd.n1853 gnd 0.007435f
C4078 vdd.n1854 gnd 0.009237f
C4079 vdd.n1856 gnd 0.009237f
C4080 vdd.n1857 gnd 0.009237f
C4081 vdd.n1858 gnd 0.007435f
C4082 vdd.n1859 gnd 0.007435f
C4083 vdd.n1860 gnd 0.007435f
C4084 vdd.n1861 gnd 0.009237f
C4085 vdd.n1863 gnd 0.009237f
C4086 vdd.n1864 gnd 0.009237f
C4087 vdd.n1865 gnd 0.007435f
C4088 vdd.n1866 gnd 0.009237f
C4089 vdd.n1867 gnd 0.009237f
C4090 vdd.n1868 gnd 0.009237f
C4091 vdd.n1869 gnd 0.015167f
C4092 vdd.n1870 gnd 0.006208f
C4093 vdd.n1871 gnd 0.007435f
C4094 vdd.n1872 gnd 0.009237f
C4095 vdd.n1874 gnd 0.009237f
C4096 vdd.n1875 gnd 0.009237f
C4097 vdd.n1876 gnd 0.007435f
C4098 vdd.n1877 gnd 0.007435f
C4099 vdd.n1878 gnd 0.007435f
C4100 vdd.n1879 gnd 0.009237f
C4101 vdd.n1881 gnd 0.009237f
C4102 vdd.n1882 gnd 0.009237f
C4103 vdd.n1883 gnd 0.007435f
C4104 vdd.n1884 gnd 0.007435f
C4105 vdd.n1885 gnd 0.007435f
C4106 vdd.n1886 gnd 0.009237f
C4107 vdd.n1888 gnd 0.009237f
C4108 vdd.n1889 gnd 0.009237f
C4109 vdd.n1891 gnd 0.009237f
C4110 vdd.n1892 gnd 0.007435f
C4111 vdd.n1893 gnd 0.005912f
C4112 vdd.n1894 gnd 0.840271f
C4113 vdd.n1896 gnd 0.007435f
C4114 vdd.n1897 gnd 0.007435f
C4115 vdd.n1898 gnd 0.009237f
C4116 vdd.n1900 gnd 0.009237f
C4117 vdd.n1901 gnd 0.009237f
C4118 vdd.n1902 gnd 0.007435f
C4119 vdd.n1903 gnd 0.006171f
C4120 vdd.n1904 gnd 0.022108f
C4121 vdd.n1905 gnd 0.021768f
C4122 vdd.n1906 gnd 0.006171f
C4123 vdd.n1907 gnd 0.021768f
C4124 vdd.n1908 gnd 1.29797f
C4125 vdd.n1909 gnd 0.021768f
C4126 vdd.n1910 gnd 0.022108f
C4127 vdd.n1911 gnd 0.003531f
C4128 vdd.t119 gnd 0.113639f
C4129 vdd.t118 gnd 0.121449f
C4130 vdd.t116 gnd 0.148411f
C4131 vdd.n1912 gnd 0.190242f
C4132 vdd.n1913 gnd 0.159838f
C4133 vdd.n1914 gnd 0.011449f
C4134 vdd.n1915 gnd 0.003903f
C4135 vdd.n1916 gnd 0.007944f
C4136 vdd.n1917 gnd 0.840271f
C4137 vdd.n1918 gnd 0.033049f
C4138 vdd.n1919 gnd 0.006281f
C4139 vdd.n1920 gnd 0.006281f
C4140 vdd.n1921 gnd 0.006281f
C4141 vdd.n1922 gnd 0.006281f
C4142 vdd.n1923 gnd 0.006281f
C4143 vdd.n1924 gnd 0.006281f
C4144 vdd.n1925 gnd 0.006281f
C4145 vdd.n1926 gnd 0.006281f
C4146 vdd.n1928 gnd 0.006281f
C4147 vdd.n1930 gnd 0.006281f
C4148 vdd.n1931 gnd 0.006281f
C4149 vdd.n1932 gnd 0.006281f
C4150 vdd.n1933 gnd 0.006281f
C4151 vdd.n1934 gnd 0.006281f
C4152 vdd.n1936 gnd 0.006281f
C4153 vdd.n1938 gnd 0.006281f
C4154 vdd.n1939 gnd 0.006281f
C4155 vdd.n1940 gnd 0.006281f
C4156 vdd.n1941 gnd 0.006281f
C4157 vdd.n1942 gnd 0.006281f
C4158 vdd.n1944 gnd 0.006281f
C4159 vdd.n1946 gnd 0.006281f
C4160 vdd.n1947 gnd 0.006281f
C4161 vdd.n1948 gnd 0.006281f
C4162 vdd.n1949 gnd 0.006281f
C4163 vdd.n1950 gnd 0.006281f
C4164 vdd.n1952 gnd 0.006281f
C4165 vdd.n1954 gnd 0.006281f
C4166 vdd.n1955 gnd 0.006281f
C4167 vdd.n1956 gnd 0.006281f
C4168 vdd.n1957 gnd 0.006281f
C4169 vdd.n1958 gnd 0.006281f
C4170 vdd.n1960 gnd 0.006281f
C4171 vdd.n1962 gnd 0.006281f
C4172 vdd.n1963 gnd 0.006281f
C4173 vdd.n1964 gnd 0.006281f
C4174 vdd.n1965 gnd 0.006281f
C4175 vdd.n1966 gnd 0.006281f
C4176 vdd.n1968 gnd 0.006281f
C4177 vdd.n1970 gnd 0.006281f
C4178 vdd.n1971 gnd 0.006281f
C4179 vdd.n1972 gnd 0.006281f
C4180 vdd.n1973 gnd 0.006281f
C4181 vdd.n1974 gnd 0.006281f
C4182 vdd.n1976 gnd 0.006281f
C4183 vdd.n1978 gnd 0.006281f
C4184 vdd.n1979 gnd 0.006281f
C4185 vdd.n1980 gnd 0.006281f
C4186 vdd.n1981 gnd 0.006281f
C4187 vdd.n1982 gnd 0.006281f
C4188 vdd.n1984 gnd 0.006281f
C4189 vdd.n1986 gnd 0.006281f
C4190 vdd.n1987 gnd 0.006281f
C4191 vdd.n1988 gnd 0.004572f
C4192 vdd.n1989 gnd 0.008977f
C4193 vdd.n1990 gnd 0.004849f
C4194 vdd.n1991 gnd 0.006281f
C4195 vdd.n1993 gnd 0.006281f
C4196 vdd.n1994 gnd 0.014477f
C4197 vdd.n1995 gnd 0.014477f
C4198 vdd.n1996 gnd 0.013603f
C4199 vdd.n1997 gnd 0.006281f
C4200 vdd.n1998 gnd 0.006281f
C4201 vdd.n1999 gnd 0.006281f
C4202 vdd.n2000 gnd 0.006281f
C4203 vdd.n2001 gnd 0.006281f
C4204 vdd.n2002 gnd 0.006281f
C4205 vdd.n2003 gnd 0.006281f
C4206 vdd.n2004 gnd 0.006281f
C4207 vdd.n2005 gnd 0.006281f
C4208 vdd.n2006 gnd 0.006281f
C4209 vdd.n2007 gnd 0.006281f
C4210 vdd.n2008 gnd 0.006281f
C4211 vdd.n2009 gnd 0.006281f
C4212 vdd.n2010 gnd 0.006281f
C4213 vdd.n2011 gnd 0.006281f
C4214 vdd.n2012 gnd 0.006281f
C4215 vdd.n2013 gnd 0.006281f
C4216 vdd.n2014 gnd 0.006281f
C4217 vdd.n2015 gnd 0.006281f
C4218 vdd.n2016 gnd 0.006281f
C4219 vdd.n2017 gnd 0.006281f
C4220 vdd.n2018 gnd 0.006281f
C4221 vdd.n2019 gnd 0.006281f
C4222 vdd.n2020 gnd 0.006281f
C4223 vdd.n2021 gnd 0.006281f
C4224 vdd.n2022 gnd 0.006281f
C4225 vdd.n2023 gnd 0.006281f
C4226 vdd.n2024 gnd 0.006281f
C4227 vdd.n2025 gnd 0.006281f
C4228 vdd.n2026 gnd 0.006281f
C4229 vdd.n2027 gnd 0.006281f
C4230 vdd.n2028 gnd 0.006281f
C4231 vdd.n2029 gnd 0.006281f
C4232 vdd.n2030 gnd 0.006281f
C4233 vdd.n2031 gnd 0.006281f
C4234 vdd.n2032 gnd 0.006281f
C4235 vdd.n2033 gnd 0.006281f
C4236 vdd.n2034 gnd 0.006281f
C4237 vdd.n2035 gnd 0.006281f
C4238 vdd.n2036 gnd 0.006281f
C4239 vdd.n2037 gnd 0.006281f
C4240 vdd.n2038 gnd 0.006281f
C4241 vdd.n2039 gnd 0.006281f
C4242 vdd.n2040 gnd 0.006281f
C4243 vdd.n2041 gnd 0.006281f
C4244 vdd.n2042 gnd 0.006281f
C4245 vdd.n2043 gnd 0.006281f
C4246 vdd.n2044 gnd 0.006281f
C4247 vdd.n2045 gnd 0.006281f
C4248 vdd.n2046 gnd 0.38231f
C4249 vdd.n2047 gnd 0.006281f
C4250 vdd.n2048 gnd 0.006281f
C4251 vdd.n2049 gnd 0.006281f
C4252 vdd.n2050 gnd 0.006281f
C4253 vdd.n2051 gnd 0.006281f
C4254 vdd.n2052 gnd 0.006281f
C4255 vdd.n2053 gnd 0.006281f
C4256 vdd.n2054 gnd 0.006281f
C4257 vdd.n2055 gnd 0.006281f
C4258 vdd.n2056 gnd 0.006281f
C4259 vdd.n2057 gnd 0.006281f
C4260 vdd.n2058 gnd 0.580545f
C4261 vdd.n2059 gnd 0.006281f
C4262 vdd.n2060 gnd 0.006281f
C4263 vdd.n2061 gnd 0.006281f
C4264 vdd.n2062 gnd 0.006281f
C4265 vdd.n2063 gnd 0.006281f
C4266 vdd.n2064 gnd 0.006281f
C4267 vdd.n2065 gnd 0.006281f
C4268 vdd.n2066 gnd 0.006281f
C4269 vdd.n2067 gnd 0.006281f
C4270 vdd.n2068 gnd 0.006281f
C4271 vdd.n2069 gnd 0.006281f
C4272 vdd.n2070 gnd 0.202955f
C4273 vdd.n2071 gnd 0.006281f
C4274 vdd.n2072 gnd 0.006281f
C4275 vdd.n2073 gnd 0.006281f
C4276 vdd.n2074 gnd 0.006281f
C4277 vdd.n2075 gnd 0.006281f
C4278 vdd.n2076 gnd 0.006281f
C4279 vdd.n2077 gnd 0.006281f
C4280 vdd.n2078 gnd 0.006281f
C4281 vdd.n2079 gnd 0.006281f
C4282 vdd.n2080 gnd 0.006281f
C4283 vdd.n2081 gnd 0.006281f
C4284 vdd.n2082 gnd 0.006281f
C4285 vdd.n2083 gnd 0.006281f
C4286 vdd.n2084 gnd 0.006281f
C4287 vdd.n2085 gnd 0.006281f
C4288 vdd.n2086 gnd 0.006281f
C4289 vdd.n2087 gnd 0.006281f
C4290 vdd.n2088 gnd 0.006281f
C4291 vdd.n2089 gnd 0.006281f
C4292 vdd.n2090 gnd 0.006281f
C4293 vdd.n2091 gnd 0.006281f
C4294 vdd.n2092 gnd 0.006281f
C4295 vdd.n2093 gnd 0.006281f
C4296 vdd.n2094 gnd 0.006281f
C4297 vdd.n2095 gnd 0.006281f
C4298 vdd.n2096 gnd 0.006281f
C4299 vdd.n2097 gnd 0.006281f
C4300 vdd.n2098 gnd 0.006281f
C4301 vdd.n2099 gnd 0.006281f
C4302 vdd.n2100 gnd 0.006281f
C4303 vdd.n2101 gnd 0.006281f
C4304 vdd.n2102 gnd 0.006281f
C4305 vdd.n2103 gnd 0.006281f
C4306 vdd.n2104 gnd 0.006281f
C4307 vdd.n2105 gnd 0.006281f
C4308 vdd.n2106 gnd 0.013603f
C4309 vdd.n2107 gnd 0.014477f
C4310 vdd.n2108 gnd 0.014477f
C4311 vdd.n2110 gnd 0.006281f
C4312 vdd.n2112 gnd 0.006281f
C4313 vdd.n2113 gnd 0.004849f
C4314 vdd.n2114 gnd 0.008977f
C4315 vdd.n2115 gnd 0.004572f
C4316 vdd.n2116 gnd 0.006281f
C4317 vdd.n2117 gnd 0.006281f
C4318 vdd.n2119 gnd 0.006281f
C4319 vdd.n2121 gnd 0.006281f
C4320 vdd.n2122 gnd 0.006281f
C4321 vdd.n2123 gnd 0.006281f
C4322 vdd.n2124 gnd 0.006281f
C4323 vdd.n2125 gnd 0.006281f
C4324 vdd.n2127 gnd 0.006281f
C4325 vdd.n2129 gnd 0.006281f
C4326 vdd.n2130 gnd 0.006281f
C4327 vdd.n2131 gnd 0.006281f
C4328 vdd.n2132 gnd 0.006281f
C4329 vdd.n2133 gnd 0.006281f
C4330 vdd.n2135 gnd 0.006281f
C4331 vdd.n2137 gnd 0.006281f
C4332 vdd.n2138 gnd 0.006281f
C4333 vdd.n2139 gnd 0.006281f
C4334 vdd.n2140 gnd 0.006281f
C4335 vdd.n2141 gnd 0.006281f
C4336 vdd.n2143 gnd 0.006281f
C4337 vdd.n2145 gnd 0.006281f
C4338 vdd.n2146 gnd 0.006281f
C4339 vdd.n2147 gnd 0.006281f
C4340 vdd.n2148 gnd 0.006281f
C4341 vdd.n2149 gnd 0.006281f
C4342 vdd.n2151 gnd 0.006281f
C4343 vdd.n2153 gnd 0.006281f
C4344 vdd.n2154 gnd 0.006281f
C4345 vdd.n2155 gnd 0.006281f
C4346 vdd.n2156 gnd 0.006281f
C4347 vdd.n2157 gnd 0.006281f
C4348 vdd.n2159 gnd 0.006281f
C4349 vdd.n2161 gnd 0.006281f
C4350 vdd.n2162 gnd 0.006281f
C4351 vdd.n2163 gnd 0.006281f
C4352 vdd.n2164 gnd 0.006281f
C4353 vdd.n2165 gnd 0.006281f
C4354 vdd.n2167 gnd 0.006281f
C4355 vdd.n2168 gnd 0.006281f
C4356 vdd.n2169 gnd 0.006281f
C4357 vdd.n2170 gnd 0.006281f
C4358 vdd.n2171 gnd 0.006281f
C4359 vdd.n2172 gnd 0.006281f
C4360 vdd.n2174 gnd 0.006281f
C4361 vdd.n2175 gnd 0.006281f
C4362 vdd.n2176 gnd 0.014477f
C4363 vdd.n2177 gnd 0.013603f
C4364 vdd.n2178 gnd 0.013603f
C4365 vdd.n2179 gnd 0.887337f
C4366 vdd.n2180 gnd 0.013603f
C4367 vdd.n2181 gnd 0.013603f
C4368 vdd.n2182 gnd 0.006281f
C4369 vdd.n2183 gnd 0.006281f
C4370 vdd.n2184 gnd 0.006281f
C4371 vdd.n2185 gnd 0.438949f
C4372 vdd.n2186 gnd 0.006281f
C4373 vdd.n2187 gnd 0.006281f
C4374 vdd.n2188 gnd 0.006281f
C4375 vdd.n2189 gnd 0.006281f
C4376 vdd.n2190 gnd 0.006281f
C4377 vdd.n2191 gnd 0.641903f
C4378 vdd.n2192 gnd 0.006281f
C4379 vdd.n2193 gnd 0.006281f
C4380 vdd.n2194 gnd 0.006281f
C4381 vdd.n2195 gnd 0.006281f
C4382 vdd.n2196 gnd 0.006281f
C4383 vdd.n2197 gnd 0.641903f
C4384 vdd.n2198 gnd 0.006281f
C4385 vdd.n2199 gnd 0.006281f
C4386 vdd.n2200 gnd 0.006281f
C4387 vdd.n2201 gnd 0.006281f
C4388 vdd.n2202 gnd 0.006281f
C4389 vdd.n2203 gnd 0.325672f
C4390 vdd.n2204 gnd 0.006281f
C4391 vdd.n2205 gnd 0.006281f
C4392 vdd.n2206 gnd 0.006281f
C4393 vdd.n2207 gnd 0.006281f
C4394 vdd.n2208 gnd 0.006281f
C4395 vdd.n2209 gnd 0.467268f
C4396 vdd.n2210 gnd 0.006281f
C4397 vdd.n2211 gnd 0.006281f
C4398 vdd.n2212 gnd 0.006281f
C4399 vdd.n2213 gnd 0.006281f
C4400 vdd.n2214 gnd 0.006281f
C4401 vdd.n2215 gnd 0.608864f
C4402 vdd.n2216 gnd 0.006281f
C4403 vdd.n2217 gnd 0.006281f
C4404 vdd.n2218 gnd 0.006281f
C4405 vdd.n2219 gnd 0.006281f
C4406 vdd.n2220 gnd 0.006281f
C4407 vdd.n2221 gnd 0.641903f
C4408 vdd.n2222 gnd 0.006281f
C4409 vdd.n2223 gnd 0.006281f
C4410 vdd.n2224 gnd 0.006281f
C4411 vdd.n2225 gnd 0.006281f
C4412 vdd.n2226 gnd 0.006281f
C4413 vdd.n2227 gnd 0.533346f
C4414 vdd.n2228 gnd 0.006281f
C4415 vdd.n2229 gnd 0.006281f
C4416 vdd.n2230 gnd 0.005173f
C4417 vdd.n2231 gnd 0.018196f
C4418 vdd.n2232 gnd 0.004249f
C4419 vdd.n2233 gnd 0.006281f
C4420 vdd.n2234 gnd 0.39175f
C4421 vdd.n2235 gnd 0.006281f
C4422 vdd.n2236 gnd 0.006281f
C4423 vdd.n2237 gnd 0.006281f
C4424 vdd.n2238 gnd 0.006281f
C4425 vdd.n2239 gnd 0.006281f
C4426 vdd.n2240 gnd 0.39175f
C4427 vdd.n2241 gnd 0.006281f
C4428 vdd.n2242 gnd 0.006281f
C4429 vdd.n2243 gnd 0.006281f
C4430 vdd.n2244 gnd 0.006281f
C4431 vdd.n2245 gnd 0.006281f
C4432 vdd.n2246 gnd 0.533346f
C4433 vdd.n2247 gnd 0.006281f
C4434 vdd.n2248 gnd 0.006281f
C4435 vdd.n2249 gnd 0.006281f
C4436 vdd.n2250 gnd 0.006281f
C4437 vdd.n2251 gnd 0.006281f
C4438 vdd.n2252 gnd 0.547506f
C4439 vdd.n2253 gnd 0.006281f
C4440 vdd.n2254 gnd 0.006281f
C4441 vdd.n2255 gnd 0.006281f
C4442 vdd.n2256 gnd 0.006281f
C4443 vdd.n2257 gnd 0.006281f
C4444 vdd.n2258 gnd 0.40591f
C4445 vdd.n2259 gnd 0.006281f
C4446 vdd.n2260 gnd 0.006281f
C4447 vdd.n2261 gnd 0.006281f
C4448 vdd.n2262 gnd 0.006281f
C4449 vdd.n2263 gnd 0.006281f
C4450 vdd.n2264 gnd 0.202955f
C4451 vdd.n2265 gnd 0.006281f
C4452 vdd.n2266 gnd 0.006281f
C4453 vdd.n2267 gnd 0.006281f
C4454 vdd.n2268 gnd 0.006281f
C4455 vdd.n2269 gnd 0.006281f
C4456 vdd.n2270 gnd 0.202955f
C4457 vdd.n2271 gnd 0.006281f
C4458 vdd.n2272 gnd 0.006281f
C4459 vdd.n2273 gnd 0.006281f
C4460 vdd.n2274 gnd 0.006281f
C4461 vdd.n2275 gnd 0.006281f
C4462 vdd.n2276 gnd 0.641903f
C4463 vdd.n2277 gnd 0.006281f
C4464 vdd.n2278 gnd 0.006281f
C4465 vdd.n2279 gnd 0.006281f
C4466 vdd.n2280 gnd 0.006281f
C4467 vdd.n2281 gnd 0.006281f
C4468 vdd.n2282 gnd 0.006281f
C4469 vdd.n2283 gnd 0.006281f
C4470 vdd.n2284 gnd 0.462548f
C4471 vdd.n2285 gnd 0.006281f
C4472 vdd.n2286 gnd 0.006281f
C4473 vdd.n2287 gnd 0.006281f
C4474 vdd.n2288 gnd 0.006281f
C4475 vdd.n2289 gnd 0.006281f
C4476 vdd.n2290 gnd 0.006281f
C4477 vdd.n2291 gnd 0.40119f
C4478 vdd.n2292 gnd 0.006281f
C4479 vdd.n2293 gnd 0.006281f
C4480 vdd.n2294 gnd 0.006281f
C4481 vdd.n2295 gnd 0.0144f
C4482 vdd.n2296 gnd 0.013681f
C4483 vdd.n2297 gnd 0.006281f
C4484 vdd.n2298 gnd 0.006281f
C4485 vdd.n2299 gnd 0.004849f
C4486 vdd.n2300 gnd 0.006281f
C4487 vdd.n2301 gnd 0.006281f
C4488 vdd.n2302 gnd 0.004572f
C4489 vdd.n2303 gnd 0.006281f
C4490 vdd.n2304 gnd 0.006281f
C4491 vdd.n2305 gnd 0.006281f
C4492 vdd.n2306 gnd 0.006281f
C4493 vdd.n2307 gnd 0.006281f
C4494 vdd.n2308 gnd 0.006281f
C4495 vdd.n2309 gnd 0.006281f
C4496 vdd.n2310 gnd 0.006281f
C4497 vdd.n2311 gnd 0.006281f
C4498 vdd.n2312 gnd 0.006281f
C4499 vdd.n2313 gnd 0.006281f
C4500 vdd.n2314 gnd 0.006281f
C4501 vdd.n2315 gnd 0.006281f
C4502 vdd.n2316 gnd 0.006281f
C4503 vdd.n2317 gnd 0.006281f
C4504 vdd.n2318 gnd 0.006281f
C4505 vdd.n2319 gnd 0.006281f
C4506 vdd.n2320 gnd 0.006281f
C4507 vdd.n2321 gnd 0.006281f
C4508 vdd.n2322 gnd 0.006281f
C4509 vdd.n2323 gnd 0.006281f
C4510 vdd.n2324 gnd 0.006281f
C4511 vdd.n2325 gnd 0.006281f
C4512 vdd.n2326 gnd 0.006281f
C4513 vdd.n2327 gnd 0.006281f
C4514 vdd.n2328 gnd 0.006281f
C4515 vdd.n2329 gnd 0.006281f
C4516 vdd.n2330 gnd 0.006281f
C4517 vdd.n2331 gnd 0.006281f
C4518 vdd.n2332 gnd 0.006281f
C4519 vdd.n2333 gnd 0.006281f
C4520 vdd.n2334 gnd 0.006281f
C4521 vdd.n2335 gnd 0.006281f
C4522 vdd.n2336 gnd 0.006281f
C4523 vdd.n2337 gnd 0.006281f
C4524 vdd.n2338 gnd 0.006281f
C4525 vdd.n2339 gnd 0.006281f
C4526 vdd.n2340 gnd 0.006281f
C4527 vdd.n2341 gnd 0.006281f
C4528 vdd.n2342 gnd 0.006281f
C4529 vdd.n2343 gnd 0.006281f
C4530 vdd.n2344 gnd 0.006281f
C4531 vdd.n2345 gnd 0.006281f
C4532 vdd.n2346 gnd 0.006281f
C4533 vdd.n2347 gnd 0.006281f
C4534 vdd.n2348 gnd 0.006281f
C4535 vdd.n2349 gnd 0.006281f
C4536 vdd.n2350 gnd 0.006281f
C4537 vdd.n2351 gnd 0.006281f
C4538 vdd.n2352 gnd 0.006281f
C4539 vdd.n2353 gnd 0.006281f
C4540 vdd.n2354 gnd 0.006281f
C4541 vdd.n2355 gnd 0.006281f
C4542 vdd.n2356 gnd 0.006281f
C4543 vdd.n2357 gnd 0.006281f
C4544 vdd.n2358 gnd 0.006281f
C4545 vdd.n2359 gnd 0.006281f
C4546 vdd.n2360 gnd 0.006281f
C4547 vdd.n2361 gnd 0.006281f
C4548 vdd.n2362 gnd 0.006281f
C4549 vdd.n2363 gnd 0.014477f
C4550 vdd.n2364 gnd 0.013603f
C4551 vdd.n2365 gnd 0.013603f
C4552 vdd.n2366 gnd 0.745741f
C4553 vdd.n2367 gnd 0.013603f
C4554 vdd.n2368 gnd 0.014477f
C4555 vdd.n2369 gnd 0.013681f
C4556 vdd.n2370 gnd 0.006281f
C4557 vdd.n2371 gnd 0.006281f
C4558 vdd.n2372 gnd 0.006281f
C4559 vdd.n2373 gnd 0.004849f
C4560 vdd.n2374 gnd 0.008977f
C4561 vdd.n2375 gnd 0.004572f
C4562 vdd.n2376 gnd 0.006281f
C4563 vdd.n2377 gnd 0.006281f
C4564 vdd.n2378 gnd 0.006281f
C4565 vdd.n2379 gnd 0.006281f
C4566 vdd.n2380 gnd 0.006281f
C4567 vdd.n2381 gnd 0.006281f
C4568 vdd.n2382 gnd 0.006281f
C4569 vdd.n2383 gnd 0.006281f
C4570 vdd.n2384 gnd 0.006281f
C4571 vdd.n2385 gnd 0.006281f
C4572 vdd.n2386 gnd 0.006281f
C4573 vdd.n2387 gnd 0.006281f
C4574 vdd.n2388 gnd 0.006281f
C4575 vdd.n2389 gnd 0.006281f
C4576 vdd.n2390 gnd 0.006281f
C4577 vdd.n2391 gnd 0.006281f
C4578 vdd.n2392 gnd 0.006281f
C4579 vdd.n2393 gnd 0.006281f
C4580 vdd.n2394 gnd 0.006281f
C4581 vdd.n2395 gnd 0.006281f
C4582 vdd.n2396 gnd 0.006281f
C4583 vdd.n2397 gnd 0.006281f
C4584 vdd.n2398 gnd 0.006281f
C4585 vdd.n2399 gnd 0.006281f
C4586 vdd.n2400 gnd 0.006281f
C4587 vdd.n2401 gnd 0.006281f
C4588 vdd.n2402 gnd 0.006281f
C4589 vdd.n2403 gnd 0.006281f
C4590 vdd.n2404 gnd 0.006281f
C4591 vdd.n2405 gnd 0.006281f
C4592 vdd.n2406 gnd 0.006281f
C4593 vdd.n2407 gnd 0.006281f
C4594 vdd.n2408 gnd 0.006281f
C4595 vdd.n2409 gnd 0.006281f
C4596 vdd.n2410 gnd 0.006281f
C4597 vdd.n2411 gnd 0.006281f
C4598 vdd.n2412 gnd 0.006281f
C4599 vdd.n2413 gnd 0.006281f
C4600 vdd.n2414 gnd 0.006281f
C4601 vdd.n2415 gnd 0.006281f
C4602 vdd.n2416 gnd 0.006281f
C4603 vdd.n2417 gnd 0.006281f
C4604 vdd.n2418 gnd 0.006281f
C4605 vdd.n2419 gnd 0.006281f
C4606 vdd.n2420 gnd 0.006281f
C4607 vdd.n2421 gnd 0.006281f
C4608 vdd.n2422 gnd 0.006281f
C4609 vdd.n2423 gnd 0.006281f
C4610 vdd.n2424 gnd 0.006281f
C4611 vdd.n2425 gnd 0.006281f
C4612 vdd.n2426 gnd 0.006281f
C4613 vdd.n2427 gnd 0.006281f
C4614 vdd.n2428 gnd 0.006281f
C4615 vdd.n2429 gnd 0.006281f
C4616 vdd.n2430 gnd 0.006281f
C4617 vdd.n2431 gnd 0.006281f
C4618 vdd.n2432 gnd 0.006281f
C4619 vdd.n2433 gnd 0.006281f
C4620 vdd.n2434 gnd 0.006281f
C4621 vdd.n2435 gnd 0.006281f
C4622 vdd.n2436 gnd 0.014477f
C4623 vdd.n2437 gnd 0.014477f
C4624 vdd.n2438 gnd 0.7835f
C4625 vdd.t200 gnd 2.78473f
C4626 vdd.t187 gnd 2.78473f
C4627 vdd.n2472 gnd 0.006281f
C4628 vdd.t156 gnd 0.25382f
C4629 vdd.t157 gnd 0.259817f
C4630 vdd.t155 gnd 0.165704f
C4631 vdd.n2473 gnd 0.089554f
C4632 vdd.n2474 gnd 0.050798f
C4633 vdd.n2475 gnd 0.008977f
C4634 vdd.n2476 gnd 0.006281f
C4635 vdd.n2477 gnd 0.006281f
C4636 vdd.n2478 gnd 0.006281f
C4637 vdd.n2479 gnd 0.006281f
C4638 vdd.n2480 gnd 0.006281f
C4639 vdd.n2481 gnd 0.006281f
C4640 vdd.n2482 gnd 0.006281f
C4641 vdd.n2483 gnd 0.006281f
C4642 vdd.n2484 gnd 0.006281f
C4643 vdd.n2485 gnd 0.006281f
C4644 vdd.n2486 gnd 0.006281f
C4645 vdd.n2487 gnd 0.006281f
C4646 vdd.n2488 gnd 0.006281f
C4647 vdd.n2489 gnd 0.006281f
C4648 vdd.n2490 gnd 0.006281f
C4649 vdd.n2491 gnd 0.006281f
C4650 vdd.n2492 gnd 0.006281f
C4651 vdd.n2493 gnd 0.006281f
C4652 vdd.n2494 gnd 0.006281f
C4653 vdd.n2495 gnd 0.006281f
C4654 vdd.n2496 gnd 0.006281f
C4655 vdd.n2497 gnd 0.006281f
C4656 vdd.n2498 gnd 0.006281f
C4657 vdd.n2499 gnd 0.006281f
C4658 vdd.n2500 gnd 0.006281f
C4659 vdd.n2501 gnd 0.006281f
C4660 vdd.n2502 gnd 0.006281f
C4661 vdd.n2503 gnd 0.006281f
C4662 vdd.n2504 gnd 0.006281f
C4663 vdd.n2505 gnd 0.006281f
C4664 vdd.n2506 gnd 0.006281f
C4665 vdd.n2507 gnd 0.006281f
C4666 vdd.n2508 gnd 0.006281f
C4667 vdd.n2509 gnd 0.006281f
C4668 vdd.n2510 gnd 0.006281f
C4669 vdd.n2511 gnd 0.006281f
C4670 vdd.n2512 gnd 0.006281f
C4671 vdd.n2513 gnd 0.006281f
C4672 vdd.n2514 gnd 0.006281f
C4673 vdd.n2515 gnd 0.006281f
C4674 vdd.n2516 gnd 0.006281f
C4675 vdd.n2517 gnd 0.006281f
C4676 vdd.n2518 gnd 0.006281f
C4677 vdd.n2519 gnd 0.006281f
C4678 vdd.n2520 gnd 0.006281f
C4679 vdd.n2521 gnd 0.006281f
C4680 vdd.n2522 gnd 0.006281f
C4681 vdd.n2523 gnd 0.006281f
C4682 vdd.n2524 gnd 0.006281f
C4683 vdd.n2525 gnd 0.006281f
C4684 vdd.n2526 gnd 0.006281f
C4685 vdd.n2527 gnd 0.006281f
C4686 vdd.n2528 gnd 0.006281f
C4687 vdd.n2529 gnd 0.006281f
C4688 vdd.n2530 gnd 0.006281f
C4689 vdd.n2531 gnd 0.006281f
C4690 vdd.n2532 gnd 0.006281f
C4691 vdd.n2533 gnd 0.006281f
C4692 vdd.n2534 gnd 0.006281f
C4693 vdd.n2535 gnd 0.006281f
C4694 vdd.n2536 gnd 0.004572f
C4695 vdd.n2537 gnd 0.006281f
C4696 vdd.n2538 gnd 0.006281f
C4697 vdd.n2539 gnd 0.004849f
C4698 vdd.n2540 gnd 0.006281f
C4699 vdd.n2541 gnd 0.006281f
C4700 vdd.t146 gnd 0.25382f
C4701 vdd.t147 gnd 0.259817f
C4702 vdd.t144 gnd 0.165704f
C4703 vdd.n2542 gnd 0.089554f
C4704 vdd.n2543 gnd 0.050798f
C4705 vdd.n2544 gnd 0.006281f
C4706 vdd.n2545 gnd 0.006281f
C4707 vdd.n2546 gnd 0.006281f
C4708 vdd.n2547 gnd 0.006281f
C4709 vdd.n2548 gnd 0.006281f
C4710 vdd.n2549 gnd 0.006281f
C4711 vdd.n2550 gnd 0.006281f
C4712 vdd.n2551 gnd 0.006281f
C4713 vdd.n2552 gnd 0.006281f
C4714 vdd.n2553 gnd 0.006281f
C4715 vdd.n2554 gnd 0.006281f
C4716 vdd.n2555 gnd 0.006281f
C4717 vdd.n2556 gnd 0.006281f
C4718 vdd.n2557 gnd 0.006281f
C4719 vdd.n2558 gnd 0.006281f
C4720 vdd.n2559 gnd 0.006281f
C4721 vdd.n2560 gnd 0.006281f
C4722 vdd.n2561 gnd 0.006281f
C4723 vdd.n2562 gnd 0.006281f
C4724 vdd.n2563 gnd 0.006281f
C4725 vdd.n2564 gnd 0.006281f
C4726 vdd.n2565 gnd 0.006281f
C4727 vdd.n2566 gnd 0.006281f
C4728 vdd.n2567 gnd 0.006281f
C4729 vdd.n2568 gnd 0.006281f
C4730 vdd.n2569 gnd 0.006281f
C4731 vdd.n2570 gnd 0.006281f
C4732 vdd.n2571 gnd 0.006281f
C4733 vdd.n2572 gnd 0.006281f
C4734 vdd.n2573 gnd 0.006281f
C4735 vdd.n2574 gnd 0.006281f
C4736 vdd.n2575 gnd 0.006281f
C4737 vdd.n2576 gnd 0.006281f
C4738 vdd.n2577 gnd 0.006281f
C4739 vdd.n2578 gnd 0.006281f
C4740 vdd.n2579 gnd 0.006281f
C4741 vdd.n2580 gnd 0.006281f
C4742 vdd.n2581 gnd 0.006281f
C4743 vdd.n2582 gnd 0.006281f
C4744 vdd.n2583 gnd 0.006281f
C4745 vdd.n2584 gnd 0.006281f
C4746 vdd.n2585 gnd 0.006281f
C4747 vdd.n2586 gnd 0.006281f
C4748 vdd.n2587 gnd 0.006281f
C4749 vdd.n2588 gnd 0.006281f
C4750 vdd.n2589 gnd 0.006281f
C4751 vdd.n2590 gnd 0.006281f
C4752 vdd.n2591 gnd 0.006281f
C4753 vdd.n2592 gnd 0.006281f
C4754 vdd.n2593 gnd 0.006281f
C4755 vdd.n2594 gnd 0.006281f
C4756 vdd.n2595 gnd 0.006281f
C4757 vdd.n2596 gnd 0.006281f
C4758 vdd.n2597 gnd 0.006281f
C4759 vdd.n2598 gnd 0.006281f
C4760 vdd.n2599 gnd 0.006281f
C4761 vdd.n2600 gnd 0.006281f
C4762 vdd.n2601 gnd 0.004572f
C4763 vdd.n2602 gnd 0.008977f
C4764 vdd.n2603 gnd 0.004849f
C4765 vdd.n2604 gnd 0.006281f
C4766 vdd.n2605 gnd 0.006281f
C4767 vdd.n2606 gnd 0.006281f
C4768 vdd.n2607 gnd 0.014477f
C4769 vdd.n2608 gnd 0.014477f
C4770 vdd.n2609 gnd 0.013603f
C4771 vdd.n2610 gnd 0.006281f
C4772 vdd.n2611 gnd 0.006281f
C4773 vdd.n2612 gnd 0.006281f
C4774 vdd.n2613 gnd 0.006281f
C4775 vdd.n2614 gnd 0.006281f
C4776 vdd.n2615 gnd 0.006281f
C4777 vdd.n2616 gnd 0.006281f
C4778 vdd.n2617 gnd 0.006281f
C4779 vdd.n2618 gnd 0.006281f
C4780 vdd.n2619 gnd 0.006281f
C4781 vdd.n2620 gnd 0.006281f
C4782 vdd.n2621 gnd 0.006281f
C4783 vdd.n2622 gnd 0.006281f
C4784 vdd.n2623 gnd 0.006281f
C4785 vdd.n2624 gnd 0.006281f
C4786 vdd.n2625 gnd 0.006281f
C4787 vdd.n2626 gnd 0.006281f
C4788 vdd.n2627 gnd 0.006281f
C4789 vdd.n2628 gnd 0.006281f
C4790 vdd.n2629 gnd 0.006281f
C4791 vdd.n2630 gnd 0.006281f
C4792 vdd.n2631 gnd 0.006281f
C4793 vdd.n2632 gnd 0.006281f
C4794 vdd.n2633 gnd 0.006281f
C4795 vdd.n2634 gnd 0.006281f
C4796 vdd.n2635 gnd 0.006281f
C4797 vdd.n2636 gnd 0.006281f
C4798 vdd.n2637 gnd 0.006281f
C4799 vdd.n2638 gnd 0.006281f
C4800 vdd.n2639 gnd 0.006281f
C4801 vdd.n2640 gnd 0.006281f
C4802 vdd.n2641 gnd 0.006281f
C4803 vdd.n2642 gnd 0.006281f
C4804 vdd.n2643 gnd 0.006281f
C4805 vdd.n2644 gnd 0.006281f
C4806 vdd.n2645 gnd 0.006281f
C4807 vdd.n2646 gnd 0.006281f
C4808 vdd.n2647 gnd 0.006281f
C4809 vdd.n2648 gnd 0.006281f
C4810 vdd.n2649 gnd 0.006281f
C4811 vdd.n2650 gnd 0.006281f
C4812 vdd.n2651 gnd 0.006281f
C4813 vdd.n2652 gnd 0.006281f
C4814 vdd.n2653 gnd 0.006281f
C4815 vdd.n2654 gnd 0.006281f
C4816 vdd.n2655 gnd 0.006281f
C4817 vdd.n2656 gnd 0.006281f
C4818 vdd.n2657 gnd 0.006281f
C4819 vdd.n2658 gnd 0.006281f
C4820 vdd.n2659 gnd 0.006281f
C4821 vdd.n2660 gnd 0.006281f
C4822 vdd.n2661 gnd 0.006281f
C4823 vdd.n2662 gnd 0.006281f
C4824 vdd.n2663 gnd 0.006281f
C4825 vdd.n2664 gnd 0.006281f
C4826 vdd.n2665 gnd 0.006281f
C4827 vdd.n2666 gnd 0.006281f
C4828 vdd.n2667 gnd 0.006281f
C4829 vdd.n2668 gnd 0.006281f
C4830 vdd.n2669 gnd 0.006281f
C4831 vdd.n2670 gnd 0.006281f
C4832 vdd.n2671 gnd 0.006281f
C4833 vdd.n2672 gnd 0.006281f
C4834 vdd.n2673 gnd 0.006281f
C4835 vdd.n2674 gnd 0.006281f
C4836 vdd.n2675 gnd 0.006281f
C4837 vdd.n2676 gnd 0.006281f
C4838 vdd.n2677 gnd 0.006281f
C4839 vdd.n2678 gnd 0.006281f
C4840 vdd.n2679 gnd 0.006281f
C4841 vdd.n2680 gnd 0.006281f
C4842 vdd.n2681 gnd 0.006281f
C4843 vdd.n2682 gnd 0.006281f
C4844 vdd.n2683 gnd 0.006281f
C4845 vdd.n2684 gnd 0.006281f
C4846 vdd.n2685 gnd 0.006281f
C4847 vdd.n2686 gnd 0.006281f
C4848 vdd.n2687 gnd 0.006281f
C4849 vdd.n2688 gnd 0.006281f
C4850 vdd.n2689 gnd 0.202955f
C4851 vdd.n2690 gnd 0.006281f
C4852 vdd.n2691 gnd 0.006281f
C4853 vdd.n2692 gnd 0.006281f
C4854 vdd.n2693 gnd 0.006281f
C4855 vdd.n2694 gnd 0.006281f
C4856 vdd.n2695 gnd 0.006281f
C4857 vdd.n2696 gnd 0.006281f
C4858 vdd.n2697 gnd 0.006281f
C4859 vdd.n2698 gnd 0.006281f
C4860 vdd.n2699 gnd 0.006281f
C4861 vdd.n2700 gnd 0.006281f
C4862 vdd.n2701 gnd 0.580545f
C4863 vdd.n2702 gnd 0.006281f
C4864 vdd.n2703 gnd 0.006281f
C4865 vdd.n2704 gnd 0.006281f
C4866 vdd.n2705 gnd 0.006281f
C4867 vdd.n2706 gnd 0.006281f
C4868 vdd.n2707 gnd 0.006281f
C4869 vdd.n2708 gnd 0.006281f
C4870 vdd.n2709 gnd 0.006281f
C4871 vdd.n2710 gnd 0.006281f
C4872 vdd.n2711 gnd 0.006281f
C4873 vdd.n2712 gnd 0.006281f
C4874 vdd.n2713 gnd 0.38231f
C4875 vdd.n2714 gnd 0.006281f
C4876 vdd.n2715 gnd 0.006281f
C4877 vdd.n2716 gnd 0.006281f
C4878 vdd.n2717 gnd 0.006281f
C4879 vdd.n2718 gnd 0.006281f
C4880 vdd.n2719 gnd 0.013603f
C4881 vdd.n2720 gnd 0.014477f
C4882 vdd.n2721 gnd 0.014477f
C4883 vdd.n2722 gnd 0.7835f
C4884 vdd.n2724 gnd 0.006281f
C4885 vdd.n2725 gnd 0.006281f
C4886 vdd.n2726 gnd 0.014477f
C4887 vdd.n2727 gnd 0.013603f
C4888 vdd.n2728 gnd 0.013603f
C4889 vdd.n2729 gnd 0.745741f
C4890 vdd.n2730 gnd 0.013603f
C4891 vdd.n2731 gnd 0.013603f
C4892 vdd.n2732 gnd 0.006281f
C4893 vdd.n2733 gnd 0.006281f
C4894 vdd.n2734 gnd 0.006281f
C4895 vdd.n2735 gnd 0.40119f
C4896 vdd.n2736 gnd 0.006281f
C4897 vdd.n2737 gnd 0.006281f
C4898 vdd.n2738 gnd 0.006281f
C4899 vdd.n2739 gnd 0.006281f
C4900 vdd.n2740 gnd 0.006281f
C4901 vdd.n2741 gnd 0.462548f
C4902 vdd.n2742 gnd 0.006281f
C4903 vdd.n2743 gnd 0.006281f
C4904 vdd.n2744 gnd 0.006281f
C4905 vdd.n2745 gnd 0.006281f
C4906 vdd.n2746 gnd 0.006281f
C4907 vdd.n2747 gnd 0.641903f
C4908 vdd.n2748 gnd 0.006281f
C4909 vdd.n2749 gnd 0.006281f
C4910 vdd.n2750 gnd 0.006281f
C4911 vdd.n2751 gnd 0.006281f
C4912 vdd.n2752 gnd 0.006281f
C4913 vdd.n2753 gnd 0.202955f
C4914 vdd.n2754 gnd 0.006281f
C4915 vdd.n2755 gnd 0.006281f
C4916 vdd.n2756 gnd 0.006281f
C4917 vdd.n2757 gnd 0.006281f
C4918 vdd.n2758 gnd 0.006281f
C4919 vdd.n2759 gnd 0.202955f
C4920 vdd.n2760 gnd 0.006281f
C4921 vdd.n2761 gnd 0.006281f
C4922 vdd.n2762 gnd 0.006281f
C4923 vdd.n2763 gnd 0.006281f
C4924 vdd.n2764 gnd 0.006281f
C4925 vdd.n2765 gnd 0.40591f
C4926 vdd.n2766 gnd 0.006281f
C4927 vdd.n2767 gnd 0.006281f
C4928 vdd.n2768 gnd 0.006281f
C4929 vdd.n2769 gnd 0.006281f
C4930 vdd.n2770 gnd 0.006281f
C4931 vdd.n2771 gnd 0.547506f
C4932 vdd.n2772 gnd 0.006281f
C4933 vdd.n2773 gnd 0.006281f
C4934 vdd.n2774 gnd 0.006281f
C4935 vdd.n2775 gnd 0.006281f
C4936 vdd.n2776 gnd 0.006281f
C4937 vdd.n2777 gnd 0.533346f
C4938 vdd.n2778 gnd 0.006281f
C4939 vdd.n2779 gnd 0.006281f
C4940 vdd.n2780 gnd 0.006281f
C4941 vdd.n2781 gnd 0.006281f
C4942 vdd.n2782 gnd 0.006281f
C4943 vdd.n2783 gnd 0.39175f
C4944 vdd.n2784 gnd 0.006281f
C4945 vdd.n2785 gnd 0.006281f
C4946 vdd.n2786 gnd 0.006281f
C4947 vdd.n2787 gnd 0.006281f
C4948 vdd.n2788 gnd 0.006281f
C4949 vdd.n2789 gnd 0.39175f
C4950 vdd.n2790 gnd 0.006281f
C4951 vdd.n2791 gnd 0.004249f
C4952 vdd.n2792 gnd 0.018196f
C4953 vdd.n2793 gnd 0.005173f
C4954 vdd.n2794 gnd 0.006281f
C4955 vdd.n2795 gnd 0.006281f
C4956 vdd.n2796 gnd 0.533346f
C4957 vdd.n2797 gnd 0.006281f
C4958 vdd.n2798 gnd 0.006281f
C4959 vdd.n2799 gnd 0.006281f
C4960 vdd.n2800 gnd 0.006281f
C4961 vdd.n2801 gnd 0.006281f
C4962 vdd.n2802 gnd 0.641903f
C4963 vdd.n2803 gnd 0.006281f
C4964 vdd.n2804 gnd 0.006281f
C4965 vdd.n2805 gnd 0.006281f
C4966 vdd.n2806 gnd 0.006281f
C4967 vdd.n2807 gnd 0.006281f
C4968 vdd.n2808 gnd 0.608864f
C4969 vdd.n2809 gnd 0.006281f
C4970 vdd.n2810 gnd 0.006281f
C4971 vdd.n2811 gnd 0.006281f
C4972 vdd.n2812 gnd 0.006281f
C4973 vdd.n2813 gnd 0.006281f
C4974 vdd.n2814 gnd 0.467268f
C4975 vdd.n2815 gnd 0.006281f
C4976 vdd.n2816 gnd 0.006281f
C4977 vdd.n2817 gnd 0.006281f
C4978 vdd.n2818 gnd 0.006281f
C4979 vdd.n2819 gnd 0.006281f
C4980 vdd.n2820 gnd 0.325672f
C4981 vdd.n2821 gnd 0.006281f
C4982 vdd.n2822 gnd 0.006281f
C4983 vdd.n2823 gnd 0.006281f
C4984 vdd.n2824 gnd 0.006281f
C4985 vdd.n2825 gnd 0.006281f
C4986 vdd.n2826 gnd 0.641903f
C4987 vdd.n2827 gnd 0.006281f
C4988 vdd.n2828 gnd 0.006281f
C4989 vdd.n2829 gnd 0.006281f
C4990 vdd.n2830 gnd 0.006281f
C4991 vdd.n2831 gnd 0.006281f
C4992 vdd.n2832 gnd 0.006281f
C4993 vdd.n2834 gnd 0.006281f
C4994 vdd.n2835 gnd 0.006281f
C4995 vdd.n2837 gnd 0.006281f
C4996 vdd.n2838 gnd 0.006281f
C4997 vdd.n2841 gnd 0.006281f
C4998 vdd.n2842 gnd 0.006281f
C4999 vdd.n2843 gnd 0.006281f
C5000 vdd.n2844 gnd 0.006281f
C5001 vdd.n2846 gnd 0.006281f
C5002 vdd.n2847 gnd 0.006281f
C5003 vdd.n2848 gnd 0.006281f
C5004 vdd.n2849 gnd 0.006281f
C5005 vdd.n2850 gnd 0.006281f
C5006 vdd.n2851 gnd 0.006281f
C5007 vdd.n2853 gnd 0.006281f
C5008 vdd.n2854 gnd 0.006281f
C5009 vdd.n2855 gnd 0.006281f
C5010 vdd.n2856 gnd 0.006281f
C5011 vdd.n2857 gnd 0.006281f
C5012 vdd.n2858 gnd 0.006281f
C5013 vdd.n2860 gnd 0.006281f
C5014 vdd.n2861 gnd 0.006281f
C5015 vdd.n2862 gnd 0.006281f
C5016 vdd.n2863 gnd 0.006281f
C5017 vdd.n2864 gnd 0.006281f
C5018 vdd.n2865 gnd 0.006281f
C5019 vdd.n2867 gnd 0.006281f
C5020 vdd.n2868 gnd 0.014477f
C5021 vdd.n2869 gnd 0.014477f
C5022 vdd.n2870 gnd 0.013603f
C5023 vdd.n2871 gnd 0.006281f
C5024 vdd.n2872 gnd 0.006281f
C5025 vdd.n2873 gnd 0.006281f
C5026 vdd.n2874 gnd 0.006281f
C5027 vdd.n2875 gnd 0.006281f
C5028 vdd.n2876 gnd 0.006281f
C5029 vdd.n2877 gnd 0.641903f
C5030 vdd.n2878 gnd 0.006281f
C5031 vdd.n2879 gnd 0.006281f
C5032 vdd.n2880 gnd 0.006281f
C5033 vdd.n2881 gnd 0.006281f
C5034 vdd.n2882 gnd 0.006281f
C5035 vdd.n2883 gnd 0.438949f
C5036 vdd.n2884 gnd 0.006281f
C5037 vdd.n2885 gnd 0.006281f
C5038 vdd.n2886 gnd 0.006281f
C5039 vdd.n2887 gnd 0.0144f
C5040 vdd.n2889 gnd 0.014477f
C5041 vdd.n2890 gnd 0.013681f
C5042 vdd.n2891 gnd 0.006281f
C5043 vdd.n2892 gnd 0.004849f
C5044 vdd.n2893 gnd 0.006281f
C5045 vdd.n2895 gnd 0.006281f
C5046 vdd.n2896 gnd 0.006281f
C5047 vdd.n2897 gnd 0.006281f
C5048 vdd.n2898 gnd 0.006281f
C5049 vdd.n2899 gnd 0.006281f
C5050 vdd.n2900 gnd 0.006281f
C5051 vdd.n2902 gnd 0.006281f
C5052 vdd.n2903 gnd 0.006281f
C5053 vdd.n2904 gnd 0.006281f
C5054 vdd.n2905 gnd 0.006281f
C5055 vdd.n2906 gnd 0.006281f
C5056 vdd.n2907 gnd 0.006281f
C5057 vdd.n2909 gnd 0.006281f
C5058 vdd.n2910 gnd 0.006281f
C5059 vdd.n2911 gnd 0.006281f
C5060 vdd.n2912 gnd 0.006281f
C5061 vdd.n2913 gnd 0.006281f
C5062 vdd.n2914 gnd 0.006281f
C5063 vdd.n2916 gnd 0.006281f
C5064 vdd.n2917 gnd 0.006281f
C5065 vdd.n2918 gnd 0.006281f
C5066 vdd.n2919 gnd 0.843836f
C5067 vdd.n2920 gnd 0.029484f
C5068 vdd.n2921 gnd 0.006281f
C5069 vdd.n2922 gnd 0.006281f
C5070 vdd.n2924 gnd 0.006281f
C5071 vdd.n2925 gnd 0.006281f
C5072 vdd.n2926 gnd 0.006281f
C5073 vdd.n2927 gnd 0.006281f
C5074 vdd.n2928 gnd 0.006281f
C5075 vdd.n2929 gnd 0.006281f
C5076 vdd.n2931 gnd 0.006281f
C5077 vdd.n2932 gnd 0.006281f
C5078 vdd.n2933 gnd 0.006281f
C5079 vdd.n2934 gnd 0.006281f
C5080 vdd.n2935 gnd 0.006281f
C5081 vdd.n2936 gnd 0.006281f
C5082 vdd.n2938 gnd 0.006281f
C5083 vdd.n2939 gnd 0.006281f
C5084 vdd.n2940 gnd 0.006281f
C5085 vdd.n2941 gnd 0.006281f
C5086 vdd.n2942 gnd 0.006281f
C5087 vdd.n2943 gnd 0.006281f
C5088 vdd.n2945 gnd 0.006281f
C5089 vdd.n2946 gnd 0.006281f
C5090 vdd.n2948 gnd 0.006281f
C5091 vdd.n2949 gnd 0.006281f
C5092 vdd.n2950 gnd 0.014477f
C5093 vdd.n2951 gnd 0.013603f
C5094 vdd.n2952 gnd 0.013603f
C5095 vdd.n2953 gnd 0.887337f
C5096 vdd.n2954 gnd 0.013603f
C5097 vdd.n2955 gnd 0.014477f
C5098 vdd.n2956 gnd 0.013681f
C5099 vdd.n2957 gnd 0.006281f
C5100 vdd.n2958 gnd 0.004849f
C5101 vdd.n2959 gnd 0.006281f
C5102 vdd.n2961 gnd 0.006281f
C5103 vdd.n2962 gnd 0.006281f
C5104 vdd.n2963 gnd 0.006281f
C5105 vdd.n2964 gnd 0.006281f
C5106 vdd.n2965 gnd 0.006281f
C5107 vdd.n2966 gnd 0.006281f
C5108 vdd.n2968 gnd 0.006281f
C5109 vdd.n2969 gnd 0.006281f
C5110 vdd.n2970 gnd 0.006281f
C5111 vdd.n2971 gnd 0.006281f
C5112 vdd.n2972 gnd 0.006281f
C5113 vdd.n2973 gnd 0.006281f
C5114 vdd.n2975 gnd 0.006281f
C5115 vdd.n2976 gnd 0.006281f
C5116 vdd.n2977 gnd 0.006281f
C5117 vdd.n2978 gnd 0.006281f
C5118 vdd.n2979 gnd 0.006281f
C5119 vdd.n2980 gnd 0.006281f
C5120 vdd.n2982 gnd 0.006281f
C5121 vdd.n2983 gnd 0.006281f
C5122 vdd.n2985 gnd 0.006281f
C5123 vdd.n2986 gnd 0.029484f
C5124 vdd.n2987 gnd 0.843836f
C5125 vdd.n2988 gnd 0.007944f
C5126 vdd.n2989 gnd 0.003531f
C5127 vdd.t114 gnd 0.113639f
C5128 vdd.t115 gnd 0.121449f
C5129 vdd.t113 gnd 0.148411f
C5130 vdd.n2990 gnd 0.190242f
C5131 vdd.n2991 gnd 0.159838f
C5132 vdd.n2992 gnd 0.011449f
C5133 vdd.n2993 gnd 0.009237f
C5134 vdd.n2994 gnd 0.003903f
C5135 vdd.n2995 gnd 0.007435f
C5136 vdd.n2996 gnd 0.009237f
C5137 vdd.n2997 gnd 0.009237f
C5138 vdd.n2998 gnd 0.007435f
C5139 vdd.n2999 gnd 0.007435f
C5140 vdd.n3000 gnd 0.009237f
C5141 vdd.n3002 gnd 0.009237f
C5142 vdd.n3003 gnd 0.007435f
C5143 vdd.n3004 gnd 0.007435f
C5144 vdd.n3005 gnd 0.007435f
C5145 vdd.n3006 gnd 0.009237f
C5146 vdd.n3008 gnd 0.009237f
C5147 vdd.n3010 gnd 0.009237f
C5148 vdd.n3011 gnd 0.007435f
C5149 vdd.n3012 gnd 0.007435f
C5150 vdd.n3013 gnd 0.007435f
C5151 vdd.n3014 gnd 0.009237f
C5152 vdd.n3016 gnd 0.009237f
C5153 vdd.n3018 gnd 0.009237f
C5154 vdd.n3019 gnd 0.007435f
C5155 vdd.n3020 gnd 0.007435f
C5156 vdd.n3021 gnd 0.007435f
C5157 vdd.n3022 gnd 0.009237f
C5158 vdd.n3024 gnd 0.009237f
C5159 vdd.n3025 gnd 0.009237f
C5160 vdd.n3026 gnd 0.007435f
C5161 vdd.n3027 gnd 0.007435f
C5162 vdd.n3028 gnd 0.009237f
C5163 vdd.n3029 gnd 0.009237f
C5164 vdd.n3031 gnd 0.009237f
C5165 vdd.n3032 gnd 0.007435f
C5166 vdd.n3033 gnd 0.009237f
C5167 vdd.n3034 gnd 0.009237f
C5168 vdd.n3035 gnd 0.009237f
C5169 vdd.n3036 gnd 0.015167f
C5170 vdd.n3037 gnd 0.005056f
C5171 vdd.n3038 gnd 0.009237f
C5172 vdd.n3040 gnd 0.009237f
C5173 vdd.n3042 gnd 0.009237f
C5174 vdd.n3043 gnd 0.007435f
C5175 vdd.n3044 gnd 0.007435f
C5176 vdd.n3045 gnd 0.007435f
C5177 vdd.n3046 gnd 0.009237f
C5178 vdd.n3048 gnd 0.009237f
C5179 vdd.n3050 gnd 0.009237f
C5180 vdd.n3051 gnd 0.007435f
C5181 vdd.n3052 gnd 0.007435f
C5182 vdd.n3053 gnd 0.007435f
C5183 vdd.n3054 gnd 0.009237f
C5184 vdd.n3056 gnd 0.009237f
C5185 vdd.n3058 gnd 0.009237f
C5186 vdd.n3059 gnd 0.007435f
C5187 vdd.n3060 gnd 0.007435f
C5188 vdd.n3061 gnd 0.007435f
C5189 vdd.n3062 gnd 0.009237f
C5190 vdd.n3064 gnd 0.009237f
C5191 vdd.n3066 gnd 0.009237f
C5192 vdd.n3067 gnd 0.007435f
C5193 vdd.n3068 gnd 0.007435f
C5194 vdd.n3069 gnd 0.007435f
C5195 vdd.n3070 gnd 0.009237f
C5196 vdd.n3072 gnd 0.009237f
C5197 vdd.n3074 gnd 0.009237f
C5198 vdd.n3075 gnd 0.007435f
C5199 vdd.n3076 gnd 0.007435f
C5200 vdd.n3077 gnd 0.006208f
C5201 vdd.n3078 gnd 0.009237f
C5202 vdd.n3080 gnd 0.009237f
C5203 vdd.n3082 gnd 0.009237f
C5204 vdd.n3083 gnd 0.006208f
C5205 vdd.n3084 gnd 0.007435f
C5206 vdd.n3085 gnd 0.007435f
C5207 vdd.n3086 gnd 0.009237f
C5208 vdd.n3088 gnd 0.009237f
C5209 vdd.n3090 gnd 0.009237f
C5210 vdd.n3091 gnd 0.007435f
C5211 vdd.n3092 gnd 0.007435f
C5212 vdd.n3093 gnd 0.007435f
C5213 vdd.n3094 gnd 0.009237f
C5214 vdd.n3096 gnd 0.009237f
C5215 vdd.n3098 gnd 0.009237f
C5216 vdd.n3099 gnd 0.007435f
C5217 vdd.n3100 gnd 0.007435f
C5218 vdd.n3101 gnd 0.007435f
C5219 vdd.n3102 gnd 0.009237f
C5220 vdd.n3104 gnd 0.009237f
C5221 vdd.n3105 gnd 0.009237f
C5222 vdd.n3106 gnd 0.007435f
C5223 vdd.n3107 gnd 0.007435f
C5224 vdd.n3108 gnd 0.009237f
C5225 vdd.n3109 gnd 0.009237f
C5226 vdd.n3110 gnd 0.007435f
C5227 vdd.n3111 gnd 0.007435f
C5228 vdd.n3112 gnd 0.009237f
C5229 vdd.n3113 gnd 0.009237f
C5230 vdd.n3115 gnd 0.009237f
C5231 vdd.n3116 gnd 0.007435f
C5232 vdd.n3117 gnd 0.006171f
C5233 vdd.n3118 gnd 0.022108f
C5234 vdd.n3119 gnd 0.021768f
C5235 vdd.n3120 gnd 0.006171f
C5236 vdd.n3121 gnd 0.021768f
C5237 vdd.n3122 gnd 1.29797f
C5238 vdd.n3123 gnd 0.021768f
C5239 vdd.n3124 gnd 0.006171f
C5240 vdd.n3125 gnd 0.021768f
C5241 vdd.n3126 gnd 0.009237f
C5242 vdd.n3127 gnd 0.009237f
C5243 vdd.n3128 gnd 0.007435f
C5244 vdd.n3129 gnd 0.009237f
C5245 vdd.n3130 gnd 0.943976f
C5246 vdd.n3131 gnd 0.009237f
C5247 vdd.n3132 gnd 0.007435f
C5248 vdd.n3133 gnd 0.009237f
C5249 vdd.n3134 gnd 0.009237f
C5250 vdd.n3135 gnd 0.009237f
C5251 vdd.n3136 gnd 0.007435f
C5252 vdd.n3137 gnd 0.009237f
C5253 vdd.n3138 gnd 0.835418f
C5254 vdd.n3139 gnd 0.009237f
C5255 vdd.n3140 gnd 0.007435f
C5256 vdd.n3141 gnd 0.009237f
C5257 vdd.n3142 gnd 0.009237f
C5258 vdd.n3143 gnd 0.009237f
C5259 vdd.n3144 gnd 0.007435f
C5260 vdd.n3145 gnd 0.009237f
C5261 vdd.t33 gnd 0.471988f
C5262 vdd.n3146 gnd 0.674943f
C5263 vdd.n3147 gnd 0.009237f
C5264 vdd.n3148 gnd 0.007435f
C5265 vdd.n3149 gnd 0.009237f
C5266 vdd.n3150 gnd 0.009237f
C5267 vdd.n3151 gnd 0.009237f
C5268 vdd.n3152 gnd 0.007435f
C5269 vdd.n3153 gnd 0.009237f
C5270 vdd.n3154 gnd 0.514467f
C5271 vdd.n3155 gnd 0.009237f
C5272 vdd.n3156 gnd 0.007435f
C5273 vdd.n3157 gnd 0.009237f
C5274 vdd.n3158 gnd 0.009237f
C5275 vdd.n3159 gnd 0.009237f
C5276 vdd.n3160 gnd 0.007435f
C5277 vdd.n3161 gnd 0.009237f
C5278 vdd.n3162 gnd 0.665503f
C5279 vdd.n3163 gnd 0.589985f
C5280 vdd.n3164 gnd 0.009237f
C5281 vdd.n3165 gnd 0.007435f
C5282 vdd.n3166 gnd 0.009237f
C5283 vdd.n3167 gnd 0.009237f
C5284 vdd.n3168 gnd 0.009237f
C5285 vdd.n3169 gnd 0.007435f
C5286 vdd.n3170 gnd 0.009237f
C5287 vdd.n3171 gnd 0.750461f
C5288 vdd.n3172 gnd 0.009237f
C5289 vdd.n3173 gnd 0.007435f
C5290 vdd.n3174 gnd 0.009237f
C5291 vdd.n3175 gnd 0.009237f
C5292 vdd.n3176 gnd 0.009237f
C5293 vdd.n3177 gnd 0.007435f
C5294 vdd.n3178 gnd 0.007435f
C5295 vdd.n3179 gnd 0.007435f
C5296 vdd.n3180 gnd 0.009237f
C5297 vdd.n3181 gnd 0.009237f
C5298 vdd.n3182 gnd 0.009237f
C5299 vdd.n3183 gnd 0.007435f
C5300 vdd.n3184 gnd 0.007435f
C5301 vdd.n3185 gnd 0.007435f
C5302 vdd.n3186 gnd 0.009237f
C5303 vdd.n3187 gnd 0.009237f
C5304 vdd.n3188 gnd 0.009237f
C5305 vdd.n3189 gnd 0.007435f
C5306 vdd.n3190 gnd 0.007435f
C5307 vdd.n3191 gnd 0.007435f
C5308 vdd.n3192 gnd 0.009237f
C5309 vdd.n3193 gnd 0.009237f
C5310 vdd.n3194 gnd 0.009237f
C5311 vdd.n3195 gnd 0.007435f
C5312 vdd.n3196 gnd 0.007435f
C5313 vdd.n3197 gnd 0.006171f
C5314 vdd.n3198 gnd 0.021768f
C5315 vdd.n3199 gnd 0.022108f
C5316 vdd.n3201 gnd 0.022108f
C5317 vdd.n3202 gnd 0.003531f
C5318 vdd.t127 gnd 0.113639f
C5319 vdd.t126 gnd 0.121449f
C5320 vdd.t124 gnd 0.148411f
C5321 vdd.n3203 gnd 0.190242f
C5322 vdd.n3204 gnd 0.160581f
C5323 vdd.n3205 gnd 0.012193f
C5324 vdd.n3206 gnd 0.003903f
C5325 vdd.n3207 gnd 0.007435f
C5326 vdd.n3208 gnd 0.009237f
C5327 vdd.n3210 gnd 0.009237f
C5328 vdd.n3211 gnd 0.009237f
C5329 vdd.n3212 gnd 0.007435f
C5330 vdd.n3213 gnd 0.007435f
C5331 vdd.n3214 gnd 0.007435f
C5332 vdd.n3215 gnd 0.009237f
C5333 vdd.n3217 gnd 0.009237f
C5334 vdd.n3218 gnd 0.009237f
C5335 vdd.n3219 gnd 0.007435f
C5336 vdd.n3220 gnd 0.007435f
C5337 vdd.n3221 gnd 0.007435f
C5338 vdd.n3222 gnd 0.009237f
C5339 vdd.n3224 gnd 0.009237f
C5340 vdd.n3225 gnd 0.009237f
C5341 vdd.n3226 gnd 0.007435f
C5342 vdd.n3227 gnd 0.007435f
C5343 vdd.n3228 gnd 0.007435f
C5344 vdd.n3229 gnd 0.009237f
C5345 vdd.n3231 gnd 0.009237f
C5346 vdd.n3232 gnd 0.009237f
C5347 vdd.n3233 gnd 0.007435f
C5348 vdd.n3234 gnd 0.007435f
C5349 vdd.n3235 gnd 0.007435f
C5350 vdd.n3236 gnd 0.009237f
C5351 vdd.n3238 gnd 0.009237f
C5352 vdd.n3239 gnd 0.009237f
C5353 vdd.n3240 gnd 0.007435f
C5354 vdd.n3241 gnd 0.009237f
C5355 vdd.n3242 gnd 0.009237f
C5356 vdd.n3243 gnd 0.009237f
C5357 vdd.n3244 gnd 0.01591f
C5358 vdd.n3245 gnd 0.005056f
C5359 vdd.n3246 gnd 0.007435f
C5360 vdd.n3247 gnd 0.009237f
C5361 vdd.n3249 gnd 0.009237f
C5362 vdd.n3250 gnd 0.009237f
C5363 vdd.n3251 gnd 0.007435f
C5364 vdd.n3252 gnd 0.007435f
C5365 vdd.n3253 gnd 0.007435f
C5366 vdd.n3254 gnd 0.009237f
C5367 vdd.n3256 gnd 0.009237f
C5368 vdd.n3257 gnd 0.009237f
C5369 vdd.n3258 gnd 0.007435f
C5370 vdd.n3259 gnd 0.007435f
C5371 vdd.n3260 gnd 0.007435f
C5372 vdd.n3261 gnd 0.009237f
C5373 vdd.n3263 gnd 0.009237f
C5374 vdd.n3264 gnd 0.009237f
C5375 vdd.n3265 gnd 0.007435f
C5376 vdd.n3266 gnd 0.007435f
C5377 vdd.n3267 gnd 0.007435f
C5378 vdd.n3268 gnd 0.009237f
C5379 vdd.n3270 gnd 0.009237f
C5380 vdd.n3271 gnd 0.009237f
C5381 vdd.n3272 gnd 0.007435f
C5382 vdd.n3273 gnd 0.007435f
C5383 vdd.n3274 gnd 0.007435f
C5384 vdd.n3275 gnd 0.009237f
C5385 vdd.n3277 gnd 0.009237f
C5386 vdd.n3278 gnd 0.009237f
C5387 vdd.n3279 gnd 0.007435f
C5388 vdd.n3280 gnd 0.009237f
C5389 vdd.n3281 gnd 0.009237f
C5390 vdd.n3282 gnd 0.009237f
C5391 vdd.n3283 gnd 0.01591f
C5392 vdd.n3284 gnd 0.006208f
C5393 vdd.n3285 gnd 0.007435f
C5394 vdd.n3286 gnd 0.009237f
C5395 vdd.n3288 gnd 0.009237f
C5396 vdd.n3289 gnd 0.009237f
C5397 vdd.n3290 gnd 0.007435f
C5398 vdd.n3291 gnd 0.007435f
C5399 vdd.n3292 gnd 0.007435f
C5400 vdd.n3293 gnd 0.009237f
C5401 vdd.n3295 gnd 0.009237f
C5402 vdd.n3296 gnd 0.009237f
C5403 vdd.n3297 gnd 0.007435f
C5404 vdd.n3298 gnd 0.007435f
C5405 vdd.n3299 gnd 0.007435f
C5406 vdd.n3300 gnd 0.009237f
C5407 vdd.n3302 gnd 0.009237f
C5408 vdd.n3303 gnd 0.009237f
C5409 vdd.n3304 gnd 0.007435f
C5410 vdd.n3305 gnd 0.007435f
C5411 vdd.n3306 gnd 0.007435f
C5412 vdd.n3307 gnd 0.009237f
C5413 vdd.n3309 gnd 0.009237f
C5414 vdd.n3310 gnd 0.009237f
C5415 vdd.n3312 gnd 0.009237f
C5416 vdd.n3313 gnd 0.007435f
C5417 vdd.n3314 gnd 0.007435f
C5418 vdd.n3315 gnd 0.006171f
C5419 vdd.n3316 gnd 0.022108f
C5420 vdd.n3317 gnd 0.021768f
C5421 vdd.n3318 gnd 0.006171f
C5422 vdd.n3319 gnd 0.021768f
C5423 vdd.n3320 gnd 1.33101f
C5424 vdd.n3321 gnd 0.533346f
C5425 vdd.t125 gnd 0.471988f
C5426 vdd.n3322 gnd 0.882617f
C5427 vdd.n3323 gnd 0.009237f
C5428 vdd.n3324 gnd 0.007435f
C5429 vdd.n3325 gnd 0.007435f
C5430 vdd.n3326 gnd 0.007435f
C5431 vdd.n3327 gnd 0.009237f
C5432 vdd.n3328 gnd 0.929816f
C5433 vdd.t0 gnd 0.471988f
C5434 vdd.n3329 gnd 0.486147f
C5435 vdd.n3330 gnd 0.76934f
C5436 vdd.n3331 gnd 0.009237f
C5437 vdd.n3332 gnd 0.007435f
C5438 vdd.n3333 gnd 0.007435f
C5439 vdd.n3334 gnd 0.007435f
C5440 vdd.n3335 gnd 0.009237f
C5441 vdd.n3336 gnd 0.608864f
C5442 vdd.t57 gnd 0.471988f
C5443 vdd.n3337 gnd 0.7835f
C5444 vdd.t21 gnd 0.471988f
C5445 vdd.n3338 gnd 0.495587f
C5446 vdd.n3339 gnd 0.009237f
C5447 vdd.n3340 gnd 0.007435f
C5448 vdd.n3341 gnd 0.007435f
C5449 vdd.n3342 gnd 0.007435f
C5450 vdd.n3343 gnd 0.009237f
C5451 vdd.n3344 gnd 0.656063f
C5452 vdd.n3345 gnd 0.599425f
C5453 vdd.t10 gnd 0.471988f
C5454 vdd.n3346 gnd 0.7835f
C5455 vdd.n3347 gnd 0.009237f
C5456 vdd.n3348 gnd 0.007435f
C5457 vdd.n3349 gnd 0.549857f
C5458 vdd.n3350 gnd 2.25893f
C5459 a_n2472_13878.t17 gnd 0.187752f
C5460 a_n2472_13878.t19 gnd 0.187752f
C5461 a_n2472_13878.t11 gnd 0.187752f
C5462 a_n2472_13878.n0 gnd 1.47995f
C5463 a_n2472_13878.t16 gnd 0.187752f
C5464 a_n2472_13878.t10 gnd 0.187752f
C5465 a_n2472_13878.n1 gnd 1.47838f
C5466 a_n2472_13878.n2 gnd 2.06575f
C5467 a_n2472_13878.t6 gnd 0.187752f
C5468 a_n2472_13878.t8 gnd 0.187752f
C5469 a_n2472_13878.n3 gnd 1.47838f
C5470 a_n2472_13878.n4 gnd 1.00763f
C5471 a_n2472_13878.t18 gnd 0.187752f
C5472 a_n2472_13878.t7 gnd 0.187752f
C5473 a_n2472_13878.n5 gnd 1.47838f
C5474 a_n2472_13878.n6 gnd 1.00763f
C5475 a_n2472_13878.t15 gnd 0.187752f
C5476 a_n2472_13878.t5 gnd 0.187752f
C5477 a_n2472_13878.n7 gnd 1.47838f
C5478 a_n2472_13878.n8 gnd 4.40971f
C5479 a_n2472_13878.t2 gnd 1.75801f
C5480 a_n2472_13878.t24 gnd 0.187752f
C5481 a_n2472_13878.t25 gnd 0.187752f
C5482 a_n2472_13878.n9 gnd 1.32252f
C5483 a_n2472_13878.n10 gnd 1.47772f
C5484 a_n2472_13878.t27 gnd 1.75451f
C5485 a_n2472_13878.n11 gnd 0.743612f
C5486 a_n2472_13878.t1 gnd 1.75451f
C5487 a_n2472_13878.n12 gnd 0.743612f
C5488 a_n2472_13878.t0 gnd 0.187752f
C5489 a_n2472_13878.t26 gnd 0.187752f
C5490 a_n2472_13878.n13 gnd 1.32252f
C5491 a_n2472_13878.n14 gnd 0.750813f
C5492 a_n2472_13878.t3 gnd 1.75451f
C5493 a_n2472_13878.n15 gnd 2.43968f
C5494 a_n2472_13878.n16 gnd 3.23176f
C5495 a_n2472_13878.t20 gnd 0.187752f
C5496 a_n2472_13878.t9 gnd 0.187752f
C5497 a_n2472_13878.n17 gnd 1.47838f
C5498 a_n2472_13878.n18 gnd 2.22265f
C5499 a_n2472_13878.t12 gnd 0.187752f
C5500 a_n2472_13878.t13 gnd 0.187752f
C5501 a_n2472_13878.n19 gnd 1.47838f
C5502 a_n2472_13878.n20 gnd 0.655033f
C5503 a_n2472_13878.t21 gnd 0.187752f
C5504 a_n2472_13878.t22 gnd 0.187752f
C5505 a_n2472_13878.n21 gnd 1.47838f
C5506 a_n2472_13878.n22 gnd 0.655033f
C5507 a_n2472_13878.t4 gnd 0.187752f
C5508 a_n2472_13878.t14 gnd 0.187752f
C5509 a_n2472_13878.n23 gnd 1.47838f
C5510 a_n2472_13878.n24 gnd 1.32888f
C5511 a_n2472_13878.n25 gnd 1.48083f
C5512 a_n2472_13878.t23 gnd 0.187752f
C5513 a_n2650_13878.n0 gnd 2.71632f
C5514 a_n2650_13878.n1 gnd 3.9242f
C5515 a_n2650_13878.n2 gnd 3.79431f
C5516 a_n2650_13878.n3 gnd 0.209626f
C5517 a_n2650_13878.n4 gnd 0.209626f
C5518 a_n2650_13878.n5 gnd 0.779569f
C5519 a_n2650_13878.n6 gnd 0.209626f
C5520 a_n2650_13878.n7 gnd 0.907703f
C5521 a_n2650_13878.n8 gnd 0.209626f
C5522 a_n2650_13878.n9 gnd 0.487486f
C5523 a_n2650_13878.n10 gnd 0.779488f
C5524 a_n2650_13878.n11 gnd 0.198901f
C5525 a_n2650_13878.n12 gnd 0.146494f
C5526 a_n2650_13878.n13 gnd 0.230242f
C5527 a_n2650_13878.n14 gnd 0.177836f
C5528 a_n2650_13878.n15 gnd 0.198901f
C5529 a_n2650_13878.n16 gnd 1.20434f
C5530 a_n2650_13878.n17 gnd 0.146494f
C5531 a_n2650_13878.n18 gnd 0.831895f
C5532 a_n2650_13878.n19 gnd 0.209626f
C5533 a_n2650_13878.n20 gnd 0.676448f
C5534 a_n2650_13878.n21 gnd 0.209626f
C5535 a_n2650_13878.n22 gnd 0.488406f
C5536 a_n2650_13878.n23 gnd 0.209626f
C5537 a_n2650_13878.n24 gnd 0.540812f
C5538 a_n2650_13878.n25 gnd 0.209626f
C5539 a_n2650_13878.n26 gnd 0.867796f
C5540 a_n2650_13878.n27 gnd 1.14438f
C5541 a_n2650_13878.n28 gnd 1.16289f
C5542 a_n2650_13878.n29 gnd 2.17246f
C5543 a_n2650_13878.n30 gnd 1.72583f
C5544 a_n2650_13878.n31 gnd 1.40392f
C5545 a_n2650_13878.n32 gnd 1.16289f
C5546 a_n2650_13878.n33 gnd 3.13153f
C5547 a_n2650_13878.n34 gnd 0.008411f
C5548 a_n2650_13878.n35 gnd 4.05e-19
C5549 a_n2650_13878.n37 gnd 0.008116f
C5550 a_n2650_13878.n38 gnd 0.011801f
C5551 a_n2650_13878.n39 gnd 0.007808f
C5552 a_n2650_13878.n40 gnd 0.276916f
C5553 a_n2650_13878.n41 gnd 0.008411f
C5554 a_n2650_13878.n42 gnd 4.05e-19
C5555 a_n2650_13878.n44 gnd 0.008116f
C5556 a_n2650_13878.n45 gnd 0.011801f
C5557 a_n2650_13878.n46 gnd 0.007808f
C5558 a_n2650_13878.n47 gnd 0.276916f
C5559 a_n2650_13878.n48 gnd 0.008116f
C5560 a_n2650_13878.n49 gnd 0.276916f
C5561 a_n2650_13878.n50 gnd 0.008116f
C5562 a_n2650_13878.n51 gnd 0.276916f
C5563 a_n2650_13878.n52 gnd 0.008116f
C5564 a_n2650_13878.n53 gnd 0.276916f
C5565 a_n2650_13878.n54 gnd 0.008116f
C5566 a_n2650_13878.n55 gnd 0.276916f
C5567 a_n2650_13878.n56 gnd 0.008411f
C5568 a_n2650_13878.n57 gnd 4.05e-19
C5569 a_n2650_13878.n59 gnd 0.008116f
C5570 a_n2650_13878.n60 gnd 0.011801f
C5571 a_n2650_13878.n61 gnd 0.007808f
C5572 a_n2650_13878.n62 gnd 0.276916f
C5573 a_n2650_13878.n63 gnd 0.008411f
C5574 a_n2650_13878.n64 gnd 4.05e-19
C5575 a_n2650_13878.n66 gnd 0.008116f
C5576 a_n2650_13878.n67 gnd 0.011801f
C5577 a_n2650_13878.n68 gnd 0.007808f
C5578 a_n2650_13878.n69 gnd 0.276916f
C5579 a_n2650_13878.t44 gnd 0.145399f
C5580 a_n2650_13878.t27 gnd 0.676325f
C5581 a_n2650_13878.t15 gnd 0.676325f
C5582 a_n2650_13878.t51 gnd 0.676325f
C5583 a_n2650_13878.n70 gnd 0.297222f
C5584 a_n2650_13878.t13 gnd 0.676325f
C5585 a_n2650_13878.t43 gnd 0.676325f
C5586 a_n2650_13878.t47 gnd 0.676325f
C5587 a_n2650_13878.n71 gnd 0.293579f
C5588 a_n2650_13878.t35 gnd 0.676325f
C5589 a_n2650_13878.t33 gnd 0.676325f
C5590 a_n2650_13878.t49 gnd 0.676325f
C5591 a_n2650_13878.n72 gnd 0.29734f
C5592 a_n2650_13878.t90 gnd 0.676325f
C5593 a_n2650_13878.t69 gnd 0.676325f
C5594 a_n2650_13878.t74 gnd 0.676325f
C5595 a_n2650_13878.n73 gnd 0.297222f
C5596 a_n2650_13878.t63 gnd 0.676325f
C5597 a_n2650_13878.t79 gnd 0.676325f
C5598 a_n2650_13878.t87 gnd 0.676325f
C5599 a_n2650_13878.n74 gnd 0.293579f
C5600 a_n2650_13878.t88 gnd 0.676325f
C5601 a_n2650_13878.t58 gnd 0.676325f
C5602 a_n2650_13878.t71 gnd 0.676325f
C5603 a_n2650_13878.n75 gnd 0.29734f
C5604 a_n2650_13878.t26 gnd 1.36144f
C5605 a_n2650_13878.t40 gnd 0.145399f
C5606 a_n2650_13878.t42 gnd 0.145399f
C5607 a_n2650_13878.n76 gnd 1.02419f
C5608 a_n2650_13878.t32 gnd 0.145399f
C5609 a_n2650_13878.t18 gnd 0.145399f
C5610 a_n2650_13878.n77 gnd 1.02419f
C5611 a_n2650_13878.t24 gnd 0.145399f
C5612 a_n2650_13878.t30 gnd 0.145399f
C5613 a_n2650_13878.n78 gnd 1.02419f
C5614 a_n2650_13878.t46 gnd 0.145399f
C5615 a_n2650_13878.t22 gnd 0.145399f
C5616 a_n2650_13878.n79 gnd 1.02419f
C5617 a_n2650_13878.t38 gnd 1.35873f
C5618 a_n2650_13878.t45 gnd 0.676325f
C5619 a_n2650_13878.n80 gnd 0.293831f
C5620 a_n2650_13878.t23 gnd 0.676325f
C5621 a_n2650_13878.t41 gnd 0.676325f
C5622 a_n2650_13878.n81 gnd 0.297222f
C5623 a_n2650_13878.t25 gnd 0.676325f
C5624 a_n2650_13878.t67 gnd 0.676325f
C5625 a_n2650_13878.n82 gnd 0.293831f
C5626 a_n2650_13878.t82 gnd 0.676325f
C5627 a_n2650_13878.t85 gnd 0.676325f
C5628 a_n2650_13878.n83 gnd 0.297222f
C5629 a_n2650_13878.t62 gnd 0.676325f
C5630 a_n2650_13878.n84 gnd 0.288248f
C5631 a_n2650_13878.t86 gnd 0.676325f
C5632 a_n2650_13878.n85 gnd 0.293256f
C5633 a_n2650_13878.t60 gnd 0.676325f
C5634 a_n2650_13878.n86 gnd 0.299896f
C5635 a_n2650_13878.t83 gnd 0.676325f
C5636 a_n2650_13878.n87 gnd 0.297355f
C5637 a_n2650_13878.n88 gnd 0.293579f
C5638 a_n2650_13878.t57 gnd 0.676325f
C5639 a_n2650_13878.n89 gnd 0.288409f
C5640 a_n2650_13878.t77 gnd 0.676325f
C5641 a_n2650_13878.n90 gnd 0.29734f
C5642 a_n2650_13878.t59 gnd 0.687657f
C5643 a_n2650_13878.n91 gnd 0.288248f
C5644 a_n2650_13878.t39 gnd 0.676325f
C5645 a_n2650_13878.n92 gnd 0.293256f
C5646 a_n2650_13878.t31 gnd 0.676325f
C5647 a_n2650_13878.n93 gnd 0.299896f
C5648 a_n2650_13878.t17 gnd 0.676325f
C5649 a_n2650_13878.n94 gnd 0.297355f
C5650 a_n2650_13878.n95 gnd 0.293579f
C5651 a_n2650_13878.t29 gnd 0.676325f
C5652 a_n2650_13878.n96 gnd 0.288409f
C5653 a_n2650_13878.t21 gnd 0.676325f
C5654 a_n2650_13878.n97 gnd 0.29734f
C5655 a_n2650_13878.t37 gnd 0.687657f
C5656 a_n2650_13878.n98 gnd 1.23608f
C5657 a_n2650_13878.t66 gnd 0.676325f
C5658 a_n2650_13878.n99 gnd 0.293579f
C5659 a_n2650_13878.t73 gnd 0.676325f
C5660 a_n2650_13878.n100 gnd 0.293579f
C5661 a_n2650_13878.t65 gnd 0.676325f
C5662 a_n2650_13878.n101 gnd 0.293579f
C5663 a_n2650_13878.t78 gnd 0.676325f
C5664 a_n2650_13878.n102 gnd 0.293579f
C5665 a_n2650_13878.t68 gnd 0.676325f
C5666 a_n2650_13878.n103 gnd 0.288248f
C5667 a_n2650_13878.t91 gnd 0.676325f
C5668 a_n2650_13878.n104 gnd 0.297355f
C5669 a_n2650_13878.t70 gnd 0.687657f
C5670 a_n2650_13878.t80 gnd 0.676325f
C5671 a_n2650_13878.n105 gnd 0.288248f
C5672 a_n2650_13878.t64 gnd 0.676325f
C5673 a_n2650_13878.n106 gnd 0.297355f
C5674 a_n2650_13878.t75 gnd 0.687657f
C5675 a_n2650_13878.t84 gnd 0.676325f
C5676 a_n2650_13878.n107 gnd 0.288248f
C5677 a_n2650_13878.t72 gnd 0.676325f
C5678 a_n2650_13878.n108 gnd 0.297355f
C5679 a_n2650_13878.t89 gnd 0.687657f
C5680 a_n2650_13878.t76 gnd 0.676325f
C5681 a_n2650_13878.n109 gnd 0.288248f
C5682 a_n2650_13878.t56 gnd 0.676325f
C5683 a_n2650_13878.n110 gnd 0.297355f
C5684 a_n2650_13878.t81 gnd 0.687657f
C5685 a_n2650_13878.n111 gnd 1.52654f
C5686 a_n2650_13878.t61 gnd 0.687657f
C5687 a_n2650_13878.n112 gnd 0.293831f
C5688 a_n2650_13878.n113 gnd 0.288409f
C5689 a_n2650_13878.n114 gnd 0.297355f
C5690 a_n2650_13878.n115 gnd 0.299896f
C5691 a_n2650_13878.n116 gnd 0.293256f
C5692 a_n2650_13878.n117 gnd 0.288248f
C5693 a_n2650_13878.t19 gnd 0.687657f
C5694 a_n2650_13878.t2 gnd 0.113088f
C5695 a_n2650_13878.t12 gnd 0.113088f
C5696 a_n2650_13878.n118 gnd 1.00223f
C5697 a_n2650_13878.t3 gnd 0.113088f
C5698 a_n2650_13878.t10 gnd 0.113088f
C5699 a_n2650_13878.n119 gnd 0.999285f
C5700 a_n2650_13878.t5 gnd 0.113088f
C5701 a_n2650_13878.t9 gnd 0.113088f
C5702 a_n2650_13878.n120 gnd 1.00223f
C5703 a_n2650_13878.t11 gnd 0.113088f
C5704 a_n2650_13878.t4 gnd 0.113088f
C5705 a_n2650_13878.n121 gnd 0.999285f
C5706 a_n2650_13878.t6 gnd 0.113088f
C5707 a_n2650_13878.t53 gnd 0.113088f
C5708 a_n2650_13878.n122 gnd 0.999285f
C5709 a_n2650_13878.t1 gnd 0.113088f
C5710 a_n2650_13878.t54 gnd 0.113088f
C5711 a_n2650_13878.n123 gnd 0.999285f
C5712 a_n2650_13878.t8 gnd 0.113088f
C5713 a_n2650_13878.t55 gnd 0.113088f
C5714 a_n2650_13878.n124 gnd 1.00223f
C5715 a_n2650_13878.t7 gnd 0.113088f
C5716 a_n2650_13878.t0 gnd 0.113088f
C5717 a_n2650_13878.n125 gnd 0.999285f
C5718 a_n2650_13878.n126 gnd 0.293831f
C5719 a_n2650_13878.n127 gnd 0.288409f
C5720 a_n2650_13878.n128 gnd 0.297355f
C5721 a_n2650_13878.n129 gnd 0.299896f
C5722 a_n2650_13878.n130 gnd 0.293256f
C5723 a_n2650_13878.n131 gnd 0.288248f
C5724 a_n2650_13878.n132 gnd 0.913993f
C5725 a_n2650_13878.t28 gnd 1.35873f
C5726 a_n2650_13878.t16 gnd 0.145399f
C5727 a_n2650_13878.t52 gnd 0.145399f
C5728 a_n2650_13878.n133 gnd 1.02419f
C5729 a_n2650_13878.t20 gnd 1.36144f
C5730 a_n2650_13878.t34 gnd 0.145399f
C5731 a_n2650_13878.t50 gnd 0.145399f
C5732 a_n2650_13878.n134 gnd 1.02419f
C5733 a_n2650_13878.t48 gnd 0.145399f
C5734 a_n2650_13878.t36 gnd 0.145399f
C5735 a_n2650_13878.n135 gnd 1.02419f
C5736 a_n2650_13878.n136 gnd 1.02419f
C5737 a_n2650_13878.t14 gnd 0.145399f
.ends

