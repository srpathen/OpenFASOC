* NGSPICE file created from diffpair.ext - technology: sky130A

.subckt diffpair minus drain_right drain_left source plus
X0 source.t30 plus.t0 drain_left.t3 a_n3110_n2688# sky130_fd_pr__nfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=1
X1 source.t3 minus.t0 drain_right.t15 a_n3110_n2688# sky130_fd_pr__nfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=1
X2 source.t4 minus.t1 drain_right.t14 a_n3110_n2688# sky130_fd_pr__nfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=1
X3 source.t29 plus.t1 drain_left.t8 a_n3110_n2688# sky130_fd_pr__nfet_01v8 ad=3.51 pd=18.78 as=1.485 ps=9.33 w=9 l=1
X4 drain_left.t6 plus.t2 source.t28 a_n3110_n2688# sky130_fd_pr__nfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=1
X5 drain_left.t13 plus.t3 source.t27 a_n3110_n2688# sky130_fd_pr__nfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=1
X6 drain_right.t13 minus.t2 source.t1 a_n3110_n2688# sky130_fd_pr__nfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=1
X7 source.t14 minus.t3 drain_right.t12 a_n3110_n2688# sky130_fd_pr__nfet_01v8 ad=3.51 pd=18.78 as=1.485 ps=9.33 w=9 l=1
X8 drain_left.t2 plus.t4 source.t26 a_n3110_n2688# sky130_fd_pr__nfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=1
X9 drain_right.t11 minus.t4 source.t10 a_n3110_n2688# sky130_fd_pr__nfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=1
X10 drain_left.t9 plus.t5 source.t25 a_n3110_n2688# sky130_fd_pr__nfet_01v8 ad=1.485 pd=9.33 as=3.51 ps=18.78 w=9 l=1
X11 source.t24 plus.t6 drain_left.t15 a_n3110_n2688# sky130_fd_pr__nfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=1
X12 drain_left.t4 plus.t7 source.t23 a_n3110_n2688# sky130_fd_pr__nfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=1
X13 drain_right.t10 minus.t5 source.t11 a_n3110_n2688# sky130_fd_pr__nfet_01v8 ad=1.485 pd=9.33 as=3.51 ps=18.78 w=9 l=1
X14 source.t22 plus.t8 drain_left.t0 a_n3110_n2688# sky130_fd_pr__nfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=1
X15 drain_left.t7 plus.t9 source.t21 a_n3110_n2688# sky130_fd_pr__nfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=1
X16 a_n3110_n2688# a_n3110_n2688# a_n3110_n2688# a_n3110_n2688# sky130_fd_pr__nfet_01v8 ad=3.51 pd=18.78 as=28.08 ps=150.24 w=9 l=1
X17 source.t2 minus.t6 drain_right.t9 a_n3110_n2688# sky130_fd_pr__nfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=1
X18 source.t20 plus.t10 drain_left.t5 a_n3110_n2688# sky130_fd_pr__nfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=1
X19 source.t19 plus.t11 drain_left.t1 a_n3110_n2688# sky130_fd_pr__nfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=1
X20 source.t18 plus.t12 drain_left.t11 a_n3110_n2688# sky130_fd_pr__nfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=1
X21 drain_right.t8 minus.t7 source.t31 a_n3110_n2688# sky130_fd_pr__nfet_01v8 ad=1.485 pd=9.33 as=3.51 ps=18.78 w=9 l=1
X22 a_n3110_n2688# a_n3110_n2688# a_n3110_n2688# a_n3110_n2688# sky130_fd_pr__nfet_01v8 ad=3.51 pd=18.78 as=0 ps=0 w=9 l=1
X23 drain_left.t10 plus.t13 source.t17 a_n3110_n2688# sky130_fd_pr__nfet_01v8 ad=1.485 pd=9.33 as=3.51 ps=18.78 w=9 l=1
X24 drain_right.t7 minus.t8 source.t6 a_n3110_n2688# sky130_fd_pr__nfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=1
X25 drain_right.t6 minus.t9 source.t7 a_n3110_n2688# sky130_fd_pr__nfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=1
X26 a_n3110_n2688# a_n3110_n2688# a_n3110_n2688# a_n3110_n2688# sky130_fd_pr__nfet_01v8 ad=3.51 pd=18.78 as=0 ps=0 w=9 l=1
X27 source.t8 minus.t10 drain_right.t5 a_n3110_n2688# sky130_fd_pr__nfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=1
X28 source.t9 minus.t11 drain_right.t4 a_n3110_n2688# sky130_fd_pr__nfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=1
X29 a_n3110_n2688# a_n3110_n2688# a_n3110_n2688# a_n3110_n2688# sky130_fd_pr__nfet_01v8 ad=3.51 pd=18.78 as=0 ps=0 w=9 l=1
X30 source.t13 minus.t12 drain_right.t3 a_n3110_n2688# sky130_fd_pr__nfet_01v8 ad=3.51 pd=18.78 as=1.485 ps=9.33 w=9 l=1
X31 source.t12 minus.t13 drain_right.t2 a_n3110_n2688# sky130_fd_pr__nfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=1
X32 drain_right.t1 minus.t14 source.t0 a_n3110_n2688# sky130_fd_pr__nfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=1
X33 source.t16 plus.t14 drain_left.t14 a_n3110_n2688# sky130_fd_pr__nfet_01v8 ad=3.51 pd=18.78 as=1.485 ps=9.33 w=9 l=1
X34 drain_right.t0 minus.t15 source.t5 a_n3110_n2688# sky130_fd_pr__nfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=1
X35 drain_left.t12 plus.t15 source.t15 a_n3110_n2688# sky130_fd_pr__nfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=1
R0 plus.n9 plus.t14 270.457
R1 plus.n49 plus.t13 270.457
R2 plus.n37 plus.t5 256.183
R3 plus.n76 plus.t1 256.183
R4 plus.n35 plus.t8 216.9
R5 plus.n29 plus.t4 216.9
R6 plus.n22 plus.t6 216.9
R7 plus.n20 plus.t3 216.9
R8 plus.n14 plus.t0 216.9
R9 plus.n8 plus.t2 216.9
R10 plus.n74 plus.t9 216.9
R11 plus.n68 plus.t12 216.9
R12 plus.n44 plus.t7 216.9
R13 plus.n60 plus.t10 216.9
R14 plus.n54 plus.t15 216.9
R15 plus.n48 plus.t11 216.9
R16 plus.n10 plus.n7 161.3
R17 plus.n12 plus.n11 161.3
R18 plus.n13 plus.n6 161.3
R19 plus.n16 plus.n15 161.3
R20 plus.n17 plus.n5 161.3
R21 plus.n19 plus.n18 161.3
R22 plus.n21 plus.n4 161.3
R23 plus.n24 plus.n23 161.3
R24 plus.n25 plus.n3 161.3
R25 plus.n27 plus.n26 161.3
R26 plus.n28 plus.n2 161.3
R27 plus.n31 plus.n30 161.3
R28 plus.n32 plus.n1 161.3
R29 plus.n34 plus.n33 161.3
R30 plus.n36 plus.n0 161.3
R31 plus.n50 plus.n47 161.3
R32 plus.n52 plus.n51 161.3
R33 plus.n53 plus.n46 161.3
R34 plus.n56 plus.n55 161.3
R35 plus.n57 plus.n45 161.3
R36 plus.n59 plus.n58 161.3
R37 plus.n61 plus.n43 161.3
R38 plus.n63 plus.n62 161.3
R39 plus.n64 plus.n42 161.3
R40 plus.n66 plus.n65 161.3
R41 plus.n67 plus.n41 161.3
R42 plus.n70 plus.n69 161.3
R43 plus.n71 plus.n40 161.3
R44 plus.n73 plus.n72 161.3
R45 plus.n75 plus.n39 161.3
R46 plus.n38 plus.n37 80.6037
R47 plus.n77 plus.n76 80.6037
R48 plus.n23 plus.n21 56.5617
R49 plus.n62 plus.n61 56.5617
R50 plus.n37 plus.n36 51.8893
R51 plus.n76 plus.n75 51.8893
R52 plus.n9 plus.n8 49.3649
R53 plus.n49 plus.n48 49.3649
R54 plus.n30 plus.n1 49.296
R55 plus.n13 plus.n12 49.296
R56 plus.n69 plus.n40 49.296
R57 plus.n53 plus.n52 49.296
R58 plus.n28 plus.n27 48.3272
R59 plus.n15 plus.n5 48.3272
R60 plus.n67 plus.n66 48.3272
R61 plus.n55 plus.n45 48.3272
R62 plus.n10 plus.n9 44.557
R63 plus.n50 plus.n49 44.557
R64 plus plus.n77 33.9919
R65 plus.n27 plus.n3 32.8269
R66 plus.n19 plus.n5 32.8269
R67 plus.n66 plus.n42 32.8269
R68 plus.n59 plus.n45 32.8269
R69 plus.n34 plus.n1 31.8581
R70 plus.n12 plus.n7 31.8581
R71 plus.n73 plus.n40 31.8581
R72 plus.n52 plus.n47 31.8581
R73 plus.n36 plus.n35 20.9036
R74 plus.n75 plus.n74 20.9036
R75 plus.n23 plus.n22 20.4117
R76 plus.n21 plus.n20 20.4117
R77 plus.n62 plus.n44 20.4117
R78 plus.n61 plus.n60 20.4117
R79 plus.n30 plus.n29 12.5423
R80 plus.n14 plus.n13 12.5423
R81 plus.n69 plus.n68 12.5423
R82 plus.n54 plus.n53 12.5423
R83 plus.n29 plus.n28 12.0505
R84 plus.n15 plus.n14 12.0505
R85 plus.n68 plus.n67 12.0505
R86 plus.n55 plus.n54 12.0505
R87 plus plus.n38 11.3532
R88 plus.n22 plus.n3 4.18111
R89 plus.n20 plus.n19 4.18111
R90 plus.n44 plus.n42 4.18111
R91 plus.n60 plus.n59 4.18111
R92 plus.n35 plus.n34 3.68928
R93 plus.n8 plus.n7 3.68928
R94 plus.n74 plus.n73 3.68928
R95 plus.n48 plus.n47 3.68928
R96 plus.n38 plus.n0 0.285035
R97 plus.n77 plus.n39 0.285035
R98 plus.n11 plus.n10 0.189894
R99 plus.n11 plus.n6 0.189894
R100 plus.n16 plus.n6 0.189894
R101 plus.n17 plus.n16 0.189894
R102 plus.n18 plus.n17 0.189894
R103 plus.n18 plus.n4 0.189894
R104 plus.n24 plus.n4 0.189894
R105 plus.n25 plus.n24 0.189894
R106 plus.n26 plus.n25 0.189894
R107 plus.n26 plus.n2 0.189894
R108 plus.n31 plus.n2 0.189894
R109 plus.n32 plus.n31 0.189894
R110 plus.n33 plus.n32 0.189894
R111 plus.n33 plus.n0 0.189894
R112 plus.n72 plus.n39 0.189894
R113 plus.n72 plus.n71 0.189894
R114 plus.n71 plus.n70 0.189894
R115 plus.n70 plus.n41 0.189894
R116 plus.n65 plus.n41 0.189894
R117 plus.n65 plus.n64 0.189894
R118 plus.n64 plus.n63 0.189894
R119 plus.n63 plus.n43 0.189894
R120 plus.n58 plus.n43 0.189894
R121 plus.n58 plus.n57 0.189894
R122 plus.n57 plus.n56 0.189894
R123 plus.n56 plus.n46 0.189894
R124 plus.n51 plus.n46 0.189894
R125 plus.n51 plus.n50 0.189894
R126 drain_left.n9 drain_left.n7 66.6841
R127 drain_left.n5 drain_left.n3 66.6839
R128 drain_left.n2 drain_left.n0 66.6839
R129 drain_left.n11 drain_left.n10 65.5376
R130 drain_left.n9 drain_left.n8 65.5376
R131 drain_left.n13 drain_left.n12 65.5374
R132 drain_left.n5 drain_left.n4 65.5373
R133 drain_left.n2 drain_left.n1 65.5373
R134 drain_left drain_left.n6 32.5469
R135 drain_left drain_left.n13 6.79977
R136 drain_left.n3 drain_left.t1 2.2005
R137 drain_left.n3 drain_left.t10 2.2005
R138 drain_left.n4 drain_left.t5 2.2005
R139 drain_left.n4 drain_left.t12 2.2005
R140 drain_left.n1 drain_left.t11 2.2005
R141 drain_left.n1 drain_left.t4 2.2005
R142 drain_left.n0 drain_left.t8 2.2005
R143 drain_left.n0 drain_left.t7 2.2005
R144 drain_left.n12 drain_left.t0 2.2005
R145 drain_left.n12 drain_left.t9 2.2005
R146 drain_left.n10 drain_left.t15 2.2005
R147 drain_left.n10 drain_left.t2 2.2005
R148 drain_left.n8 drain_left.t3 2.2005
R149 drain_left.n8 drain_left.t13 2.2005
R150 drain_left.n7 drain_left.t14 2.2005
R151 drain_left.n7 drain_left.t6 2.2005
R152 drain_left.n11 drain_left.n9 1.14705
R153 drain_left.n13 drain_left.n11 1.14705
R154 drain_left.n6 drain_left.n5 0.51843
R155 drain_left.n6 drain_left.n2 0.51843
R156 source.n7 source.t16 51.0588
R157 source.n8 source.t31 51.0588
R158 source.n15 source.t14 51.0588
R159 source.n31 source.t11 51.0586
R160 source.n24 source.t13 51.0586
R161 source.n23 source.t17 51.0586
R162 source.n16 source.t29 51.0586
R163 source.n0 source.t25 51.0586
R164 source.n2 source.n1 48.8588
R165 source.n4 source.n3 48.8588
R166 source.n6 source.n5 48.8588
R167 source.n10 source.n9 48.8588
R168 source.n12 source.n11 48.8588
R169 source.n14 source.n13 48.8588
R170 source.n30 source.n29 48.8586
R171 source.n28 source.n27 48.8586
R172 source.n26 source.n25 48.8586
R173 source.n22 source.n21 48.8586
R174 source.n20 source.n19 48.8586
R175 source.n18 source.n17 48.8586
R176 source.n16 source.n15 20.1616
R177 source.n32 source.n0 14.3253
R178 source.n32 source.n31 5.83671
R179 source.n29 source.t0 2.2005
R180 source.n29 source.t8 2.2005
R181 source.n27 source.t5 2.2005
R182 source.n27 source.t2 2.2005
R183 source.n25 source.t7 2.2005
R184 source.n25 source.t4 2.2005
R185 source.n21 source.t15 2.2005
R186 source.n21 source.t19 2.2005
R187 source.n19 source.t23 2.2005
R188 source.n19 source.t20 2.2005
R189 source.n17 source.t21 2.2005
R190 source.n17 source.t18 2.2005
R191 source.n1 source.t26 2.2005
R192 source.n1 source.t22 2.2005
R193 source.n3 source.t27 2.2005
R194 source.n3 source.t24 2.2005
R195 source.n5 source.t28 2.2005
R196 source.n5 source.t30 2.2005
R197 source.n9 source.t6 2.2005
R198 source.n9 source.t9 2.2005
R199 source.n11 source.t1 2.2005
R200 source.n11 source.t12 2.2005
R201 source.n13 source.t10 2.2005
R202 source.n13 source.t3 2.2005
R203 source.n15 source.n14 1.14705
R204 source.n14 source.n12 1.14705
R205 source.n12 source.n10 1.14705
R206 source.n10 source.n8 1.14705
R207 source.n7 source.n6 1.14705
R208 source.n6 source.n4 1.14705
R209 source.n4 source.n2 1.14705
R210 source.n2 source.n0 1.14705
R211 source.n18 source.n16 1.14705
R212 source.n20 source.n18 1.14705
R213 source.n22 source.n20 1.14705
R214 source.n23 source.n22 1.14705
R215 source.n26 source.n24 1.14705
R216 source.n28 source.n26 1.14705
R217 source.n30 source.n28 1.14705
R218 source.n31 source.n30 1.14705
R219 source.n8 source.n7 0.470328
R220 source.n24 source.n23 0.470328
R221 source source.n32 0.188
R222 minus.n10 minus.t7 270.457
R223 minus.n48 minus.t12 270.457
R224 minus.n37 minus.t3 256.183
R225 minus.n76 minus.t5 256.183
R226 minus.n9 minus.t11 216.9
R227 minus.n15 minus.t8 216.9
R228 minus.n21 minus.t13 216.9
R229 minus.n5 minus.t2 216.9
R230 minus.n29 minus.t0 216.9
R231 minus.n35 minus.t4 216.9
R232 minus.n47 minus.t9 216.9
R233 minus.n53 minus.t1 216.9
R234 minus.n59 minus.t15 216.9
R235 minus.n61 minus.t6 216.9
R236 minus.n68 minus.t14 216.9
R237 minus.n74 minus.t10 216.9
R238 minus.n36 minus.n0 161.3
R239 minus.n34 minus.n33 161.3
R240 minus.n32 minus.n1 161.3
R241 minus.n31 minus.n30 161.3
R242 minus.n28 minus.n2 161.3
R243 minus.n27 minus.n26 161.3
R244 minus.n25 minus.n3 161.3
R245 minus.n24 minus.n23 161.3
R246 minus.n22 minus.n4 161.3
R247 minus.n20 minus.n19 161.3
R248 minus.n18 minus.n6 161.3
R249 minus.n17 minus.n16 161.3
R250 minus.n14 minus.n7 161.3
R251 minus.n13 minus.n12 161.3
R252 minus.n11 minus.n8 161.3
R253 minus.n75 minus.n39 161.3
R254 minus.n73 minus.n72 161.3
R255 minus.n71 minus.n40 161.3
R256 minus.n70 minus.n69 161.3
R257 minus.n67 minus.n41 161.3
R258 minus.n66 minus.n65 161.3
R259 minus.n64 minus.n42 161.3
R260 minus.n63 minus.n62 161.3
R261 minus.n60 minus.n43 161.3
R262 minus.n58 minus.n57 161.3
R263 minus.n56 minus.n44 161.3
R264 minus.n55 minus.n54 161.3
R265 minus.n52 minus.n45 161.3
R266 minus.n51 minus.n50 161.3
R267 minus.n49 minus.n46 161.3
R268 minus.n38 minus.n37 80.6037
R269 minus.n77 minus.n76 80.6037
R270 minus.n23 minus.n22 56.5617
R271 minus.n62 minus.n60 56.5617
R272 minus.n37 minus.n36 51.8893
R273 minus.n76 minus.n75 51.8893
R274 minus.n10 minus.n9 49.3649
R275 minus.n48 minus.n47 49.3649
R276 minus.n14 minus.n13 49.296
R277 minus.n30 minus.n1 49.296
R278 minus.n52 minus.n51 49.296
R279 minus.n69 minus.n40 49.296
R280 minus.n16 minus.n6 48.3272
R281 minus.n28 minus.n27 48.3272
R282 minus.n54 minus.n44 48.3272
R283 minus.n67 minus.n66 48.3272
R284 minus.n11 minus.n10 44.557
R285 minus.n49 minus.n48 44.557
R286 minus.n78 minus.n38 38.9744
R287 minus.n20 minus.n6 32.8269
R288 minus.n27 minus.n3 32.8269
R289 minus.n58 minus.n44 32.8269
R290 minus.n66 minus.n42 32.8269
R291 minus.n13 minus.n8 31.8581
R292 minus.n34 minus.n1 31.8581
R293 minus.n51 minus.n46 31.8581
R294 minus.n73 minus.n40 31.8581
R295 minus.n36 minus.n35 20.9036
R296 minus.n75 minus.n74 20.9036
R297 minus.n22 minus.n21 20.4117
R298 minus.n23 minus.n5 20.4117
R299 minus.n60 minus.n59 20.4117
R300 minus.n62 minus.n61 20.4117
R301 minus.n15 minus.n14 12.5423
R302 minus.n30 minus.n29 12.5423
R303 minus.n53 minus.n52 12.5423
R304 minus.n69 minus.n68 12.5423
R305 minus.n16 minus.n15 12.0505
R306 minus.n29 minus.n28 12.0505
R307 minus.n54 minus.n53 12.0505
R308 minus.n68 minus.n67 12.0505
R309 minus.n78 minus.n77 6.84564
R310 minus.n21 minus.n20 4.18111
R311 minus.n5 minus.n3 4.18111
R312 minus.n59 minus.n58 4.18111
R313 minus.n61 minus.n42 4.18111
R314 minus.n9 minus.n8 3.68928
R315 minus.n35 minus.n34 3.68928
R316 minus.n47 minus.n46 3.68928
R317 minus.n74 minus.n73 3.68928
R318 minus.n38 minus.n0 0.285035
R319 minus.n77 minus.n39 0.285035
R320 minus.n33 minus.n0 0.189894
R321 minus.n33 minus.n32 0.189894
R322 minus.n32 minus.n31 0.189894
R323 minus.n31 minus.n2 0.189894
R324 minus.n26 minus.n2 0.189894
R325 minus.n26 minus.n25 0.189894
R326 minus.n25 minus.n24 0.189894
R327 minus.n24 minus.n4 0.189894
R328 minus.n19 minus.n4 0.189894
R329 minus.n19 minus.n18 0.189894
R330 minus.n18 minus.n17 0.189894
R331 minus.n17 minus.n7 0.189894
R332 minus.n12 minus.n7 0.189894
R333 minus.n12 minus.n11 0.189894
R334 minus.n50 minus.n49 0.189894
R335 minus.n50 minus.n45 0.189894
R336 minus.n55 minus.n45 0.189894
R337 minus.n56 minus.n55 0.189894
R338 minus.n57 minus.n56 0.189894
R339 minus.n57 minus.n43 0.189894
R340 minus.n63 minus.n43 0.189894
R341 minus.n64 minus.n63 0.189894
R342 minus.n65 minus.n64 0.189894
R343 minus.n65 minus.n41 0.189894
R344 minus.n70 minus.n41 0.189894
R345 minus.n71 minus.n70 0.189894
R346 minus.n72 minus.n71 0.189894
R347 minus.n72 minus.n39 0.189894
R348 minus minus.n78 0.188
R349 drain_right.n9 drain_right.n7 66.684
R350 drain_right.n5 drain_right.n3 66.6839
R351 drain_right.n2 drain_right.n0 66.6839
R352 drain_right.n9 drain_right.n8 65.5376
R353 drain_right.n11 drain_right.n10 65.5376
R354 drain_right.n13 drain_right.n12 65.5376
R355 drain_right.n5 drain_right.n4 65.5373
R356 drain_right.n2 drain_right.n1 65.5373
R357 drain_right drain_right.n6 31.9937
R358 drain_right drain_right.n13 6.79977
R359 drain_right.n3 drain_right.t5 2.2005
R360 drain_right.n3 drain_right.t10 2.2005
R361 drain_right.n4 drain_right.t9 2.2005
R362 drain_right.n4 drain_right.t1 2.2005
R363 drain_right.n1 drain_right.t14 2.2005
R364 drain_right.n1 drain_right.t0 2.2005
R365 drain_right.n0 drain_right.t3 2.2005
R366 drain_right.n0 drain_right.t6 2.2005
R367 drain_right.n7 drain_right.t4 2.2005
R368 drain_right.n7 drain_right.t8 2.2005
R369 drain_right.n8 drain_right.t2 2.2005
R370 drain_right.n8 drain_right.t7 2.2005
R371 drain_right.n10 drain_right.t15 2.2005
R372 drain_right.n10 drain_right.t13 2.2005
R373 drain_right.n12 drain_right.t12 2.2005
R374 drain_right.n12 drain_right.t11 2.2005
R375 drain_right.n13 drain_right.n11 1.14705
R376 drain_right.n11 drain_right.n9 1.14705
R377 drain_right.n6 drain_right.n5 0.51843
R378 drain_right.n6 drain_right.n2 0.51843
C0 source drain_right 13.562201f
C1 source minus 9.695651f
C2 plus drain_right 0.468824f
C3 plus minus 6.46402f
C4 drain_right minus 9.32971f
C5 source drain_left 13.5583f
C6 drain_left plus 9.64056f
C7 drain_left drain_right 1.64323f
C8 drain_left minus 0.174261f
C9 source plus 9.70969f
C10 drain_right a_n3110_n2688# 6.72435f
C11 drain_left a_n3110_n2688# 7.15598f
C12 source a_n3110_n2688# 7.928731f
C13 minus a_n3110_n2688# 12.321501f
C14 plus a_n3110_n2688# 13.8221f
C15 drain_right.t3 a_n3110_n2688# 0.182123f
C16 drain_right.t6 a_n3110_n2688# 0.182123f
C17 drain_right.n0 a_n3110_n2688# 1.59993f
C18 drain_right.t14 a_n3110_n2688# 0.182123f
C19 drain_right.t0 a_n3110_n2688# 0.182123f
C20 drain_right.n1 a_n3110_n2688# 1.59297f
C21 drain_right.n2 a_n3110_n2688# 0.741297f
C22 drain_right.t5 a_n3110_n2688# 0.182123f
C23 drain_right.t10 a_n3110_n2688# 0.182123f
C24 drain_right.n3 a_n3110_n2688# 1.59993f
C25 drain_right.t9 a_n3110_n2688# 0.182123f
C26 drain_right.t1 a_n3110_n2688# 0.182123f
C27 drain_right.n4 a_n3110_n2688# 1.59297f
C28 drain_right.n5 a_n3110_n2688# 0.741297f
C29 drain_right.n6 a_n3110_n2688# 1.40462f
C30 drain_right.t4 a_n3110_n2688# 0.182123f
C31 drain_right.t8 a_n3110_n2688# 0.182123f
C32 drain_right.n7 a_n3110_n2688# 1.59992f
C33 drain_right.t2 a_n3110_n2688# 0.182123f
C34 drain_right.t7 a_n3110_n2688# 0.182123f
C35 drain_right.n8 a_n3110_n2688# 1.59297f
C36 drain_right.n9 a_n3110_n2688# 0.792021f
C37 drain_right.t15 a_n3110_n2688# 0.182123f
C38 drain_right.t13 a_n3110_n2688# 0.182123f
C39 drain_right.n10 a_n3110_n2688# 1.59297f
C40 drain_right.n11 a_n3110_n2688# 0.394329f
C41 drain_right.t12 a_n3110_n2688# 0.182123f
C42 drain_right.t11 a_n3110_n2688# 0.182123f
C43 drain_right.n12 a_n3110_n2688# 1.59297f
C44 drain_right.n13 a_n3110_n2688# 0.629956f
C45 minus.n0 a_n3110_n2688# 0.047144f
C46 minus.t4 a_n3110_n2688# 0.858107f
C47 minus.n1 a_n3110_n2688# 0.03236f
C48 minus.n2 a_n3110_n2688# 0.03533f
C49 minus.t0 a_n3110_n2688# 0.858107f
C50 minus.n3 a_n3110_n2688# 0.044026f
C51 minus.n4 a_n3110_n2688# 0.03533f
C52 minus.t2 a_n3110_n2688# 0.858107f
C53 minus.n5 a_n3110_n2688# 0.329381f
C54 minus.t13 a_n3110_n2688# 0.858107f
C55 minus.n6 a_n3110_n2688# 0.031527f
C56 minus.n7 a_n3110_n2688# 0.03533f
C57 minus.t8 a_n3110_n2688# 0.858107f
C58 minus.n8 a_n3110_n2688# 0.043188f
C59 minus.t7 a_n3110_n2688# 0.932092f
C60 minus.t11 a_n3110_n2688# 0.858107f
C61 minus.n9 a_n3110_n2688# 0.354955f
C62 minus.n10 a_n3110_n2688# 0.381622f
C63 minus.n11 a_n3110_n2688# 0.147365f
C64 minus.n12 a_n3110_n2688# 0.03533f
C65 minus.n13 a_n3110_n2688# 0.03236f
C66 minus.n14 a_n3110_n2688# 0.049344f
C67 minus.n15 a_n3110_n2688# 0.329381f
C68 minus.n16 a_n3110_n2688# 0.049339f
C69 minus.n17 a_n3110_n2688# 0.03533f
C70 minus.n18 a_n3110_n2688# 0.03533f
C71 minus.n19 a_n3110_n2688# 0.03533f
C72 minus.n20 a_n3110_n2688# 0.044026f
C73 minus.n21 a_n3110_n2688# 0.329381f
C74 minus.n22 a_n3110_n2688# 0.04586f
C75 minus.n23 a_n3110_n2688# 0.04586f
C76 minus.n24 a_n3110_n2688# 0.03533f
C77 minus.n25 a_n3110_n2688# 0.03533f
C78 minus.n26 a_n3110_n2688# 0.03533f
C79 minus.n27 a_n3110_n2688# 0.031527f
C80 minus.n28 a_n3110_n2688# 0.049339f
C81 minus.n29 a_n3110_n2688# 0.329381f
C82 minus.n30 a_n3110_n2688# 0.049344f
C83 minus.n31 a_n3110_n2688# 0.03533f
C84 minus.n32 a_n3110_n2688# 0.03533f
C85 minus.n33 a_n3110_n2688# 0.03533f
C86 minus.n34 a_n3110_n2688# 0.043188f
C87 minus.n35 a_n3110_n2688# 0.329381f
C88 minus.n36 a_n3110_n2688# 0.044357f
C89 minus.t3 a_n3110_n2688# 0.911904f
C90 minus.n37 a_n3110_n2688# 0.382319f
C91 minus.n38 a_n3110_n2688# 1.42058f
C92 minus.n39 a_n3110_n2688# 0.047144f
C93 minus.t10 a_n3110_n2688# 0.858107f
C94 minus.n40 a_n3110_n2688# 0.03236f
C95 minus.n41 a_n3110_n2688# 0.03533f
C96 minus.t14 a_n3110_n2688# 0.858107f
C97 minus.n42 a_n3110_n2688# 0.044026f
C98 minus.n43 a_n3110_n2688# 0.03533f
C99 minus.t15 a_n3110_n2688# 0.858107f
C100 minus.n44 a_n3110_n2688# 0.031527f
C101 minus.n45 a_n3110_n2688# 0.03533f
C102 minus.t1 a_n3110_n2688# 0.858107f
C103 minus.n46 a_n3110_n2688# 0.043188f
C104 minus.t12 a_n3110_n2688# 0.932092f
C105 minus.t9 a_n3110_n2688# 0.858107f
C106 minus.n47 a_n3110_n2688# 0.354955f
C107 minus.n48 a_n3110_n2688# 0.381622f
C108 minus.n49 a_n3110_n2688# 0.147365f
C109 minus.n50 a_n3110_n2688# 0.03533f
C110 minus.n51 a_n3110_n2688# 0.03236f
C111 minus.n52 a_n3110_n2688# 0.049344f
C112 minus.n53 a_n3110_n2688# 0.329381f
C113 minus.n54 a_n3110_n2688# 0.049339f
C114 minus.n55 a_n3110_n2688# 0.03533f
C115 minus.n56 a_n3110_n2688# 0.03533f
C116 minus.n57 a_n3110_n2688# 0.03533f
C117 minus.n58 a_n3110_n2688# 0.044026f
C118 minus.n59 a_n3110_n2688# 0.329381f
C119 minus.n60 a_n3110_n2688# 0.04586f
C120 minus.t6 a_n3110_n2688# 0.858107f
C121 minus.n61 a_n3110_n2688# 0.329381f
C122 minus.n62 a_n3110_n2688# 0.04586f
C123 minus.n63 a_n3110_n2688# 0.03533f
C124 minus.n64 a_n3110_n2688# 0.03533f
C125 minus.n65 a_n3110_n2688# 0.03533f
C126 minus.n66 a_n3110_n2688# 0.031527f
C127 minus.n67 a_n3110_n2688# 0.049339f
C128 minus.n68 a_n3110_n2688# 0.329381f
C129 minus.n69 a_n3110_n2688# 0.049344f
C130 minus.n70 a_n3110_n2688# 0.03533f
C131 minus.n71 a_n3110_n2688# 0.03533f
C132 minus.n72 a_n3110_n2688# 0.03533f
C133 minus.n73 a_n3110_n2688# 0.043188f
C134 minus.n74 a_n3110_n2688# 0.329381f
C135 minus.n75 a_n3110_n2688# 0.044357f
C136 minus.t5 a_n3110_n2688# 0.911904f
C137 minus.n76 a_n3110_n2688# 0.382319f
C138 minus.n77 a_n3110_n2688# 0.271612f
C139 minus.n78 a_n3110_n2688# 1.68882f
C140 source.t25 a_n3110_n2688# 1.75532f
C141 source.n0 a_n3110_n2688# 1.08454f
C142 source.t26 a_n3110_n2688# 0.164611f
C143 source.t22 a_n3110_n2688# 0.164611f
C144 source.n1 a_n3110_n2688# 1.37802f
C145 source.n2 a_n3110_n2688# 0.386736f
C146 source.t27 a_n3110_n2688# 0.164611f
C147 source.t24 a_n3110_n2688# 0.164611f
C148 source.n3 a_n3110_n2688# 1.37802f
C149 source.n4 a_n3110_n2688# 0.386736f
C150 source.t28 a_n3110_n2688# 0.164611f
C151 source.t30 a_n3110_n2688# 0.164611f
C152 source.n5 a_n3110_n2688# 1.37802f
C153 source.n6 a_n3110_n2688# 0.386736f
C154 source.t16 a_n3110_n2688# 1.75533f
C155 source.n7 a_n3110_n2688# 0.407894f
C156 source.t31 a_n3110_n2688# 1.75533f
C157 source.n8 a_n3110_n2688# 0.407894f
C158 source.t6 a_n3110_n2688# 0.164611f
C159 source.t9 a_n3110_n2688# 0.164611f
C160 source.n9 a_n3110_n2688# 1.37802f
C161 source.n10 a_n3110_n2688# 0.386736f
C162 source.t1 a_n3110_n2688# 0.164611f
C163 source.t12 a_n3110_n2688# 0.164611f
C164 source.n11 a_n3110_n2688# 1.37802f
C165 source.n12 a_n3110_n2688# 0.386736f
C166 source.t10 a_n3110_n2688# 0.164611f
C167 source.t3 a_n3110_n2688# 0.164611f
C168 source.n13 a_n3110_n2688# 1.37802f
C169 source.n14 a_n3110_n2688# 0.386736f
C170 source.t14 a_n3110_n2688# 1.75533f
C171 source.n15 a_n3110_n2688# 1.43567f
C172 source.t29 a_n3110_n2688# 1.75532f
C173 source.n16 a_n3110_n2688# 1.43567f
C174 source.t21 a_n3110_n2688# 0.164611f
C175 source.t18 a_n3110_n2688# 0.164611f
C176 source.n17 a_n3110_n2688# 1.37801f
C177 source.n18 a_n3110_n2688# 0.386741f
C178 source.t23 a_n3110_n2688# 0.164611f
C179 source.t20 a_n3110_n2688# 0.164611f
C180 source.n19 a_n3110_n2688# 1.37801f
C181 source.n20 a_n3110_n2688# 0.386741f
C182 source.t15 a_n3110_n2688# 0.164611f
C183 source.t19 a_n3110_n2688# 0.164611f
C184 source.n21 a_n3110_n2688# 1.37801f
C185 source.n22 a_n3110_n2688# 0.386741f
C186 source.t17 a_n3110_n2688# 1.75532f
C187 source.n23 a_n3110_n2688# 0.407898f
C188 source.t13 a_n3110_n2688# 1.75532f
C189 source.n24 a_n3110_n2688# 0.407898f
C190 source.t7 a_n3110_n2688# 0.164611f
C191 source.t4 a_n3110_n2688# 0.164611f
C192 source.n25 a_n3110_n2688# 1.37801f
C193 source.n26 a_n3110_n2688# 0.386741f
C194 source.t5 a_n3110_n2688# 0.164611f
C195 source.t2 a_n3110_n2688# 0.164611f
C196 source.n27 a_n3110_n2688# 1.37801f
C197 source.n28 a_n3110_n2688# 0.386741f
C198 source.t0 a_n3110_n2688# 0.164611f
C199 source.t8 a_n3110_n2688# 0.164611f
C200 source.n29 a_n3110_n2688# 1.37801f
C201 source.n30 a_n3110_n2688# 0.386741f
C202 source.t11 a_n3110_n2688# 1.75532f
C203 source.n31 a_n3110_n2688# 0.573828f
C204 source.n32 a_n3110_n2688# 1.22943f
C205 drain_left.t8 a_n3110_n2688# 0.183706f
C206 drain_left.t7 a_n3110_n2688# 0.183706f
C207 drain_left.n0 a_n3110_n2688# 1.61383f
C208 drain_left.t11 a_n3110_n2688# 0.183706f
C209 drain_left.t4 a_n3110_n2688# 0.183706f
C210 drain_left.n1 a_n3110_n2688# 1.60681f
C211 drain_left.n2 a_n3110_n2688# 0.747737f
C212 drain_left.t1 a_n3110_n2688# 0.183706f
C213 drain_left.t10 a_n3110_n2688# 0.183706f
C214 drain_left.n3 a_n3110_n2688# 1.61383f
C215 drain_left.t5 a_n3110_n2688# 0.183706f
C216 drain_left.t12 a_n3110_n2688# 0.183706f
C217 drain_left.n4 a_n3110_n2688# 1.60681f
C218 drain_left.n5 a_n3110_n2688# 0.747737f
C219 drain_left.n6 a_n3110_n2688# 1.46896f
C220 drain_left.t14 a_n3110_n2688# 0.183706f
C221 drain_left.t6 a_n3110_n2688# 0.183706f
C222 drain_left.n7 a_n3110_n2688# 1.61383f
C223 drain_left.t3 a_n3110_n2688# 0.183706f
C224 drain_left.t13 a_n3110_n2688# 0.183706f
C225 drain_left.n8 a_n3110_n2688# 1.60681f
C226 drain_left.n9 a_n3110_n2688# 0.798895f
C227 drain_left.t15 a_n3110_n2688# 0.183706f
C228 drain_left.t2 a_n3110_n2688# 0.183706f
C229 drain_left.n10 a_n3110_n2688# 1.60681f
C230 drain_left.n11 a_n3110_n2688# 0.397755f
C231 drain_left.t0 a_n3110_n2688# 0.183706f
C232 drain_left.t9 a_n3110_n2688# 0.183706f
C233 drain_left.n12 a_n3110_n2688# 1.60681f
C234 drain_left.n13 a_n3110_n2688# 0.635435f
C235 plus.n0 a_n3110_n2688# 0.047833f
C236 plus.t5 a_n3110_n2688# 0.925225f
C237 plus.t8 a_n3110_n2688# 0.870642f
C238 plus.n1 a_n3110_n2688# 0.032833f
C239 plus.n2 a_n3110_n2688# 0.035847f
C240 plus.t4 a_n3110_n2688# 0.870642f
C241 plus.n3 a_n3110_n2688# 0.04467f
C242 plus.n4 a_n3110_n2688# 0.035847f
C243 plus.t3 a_n3110_n2688# 0.870642f
C244 plus.n5 a_n3110_n2688# 0.031987f
C245 plus.n6 a_n3110_n2688# 0.035847f
C246 plus.t0 a_n3110_n2688# 0.870642f
C247 plus.n7 a_n3110_n2688# 0.043819f
C248 plus.t2 a_n3110_n2688# 0.870642f
C249 plus.n8 a_n3110_n2688# 0.36014f
C250 plus.t14 a_n3110_n2688# 0.945708f
C251 plus.n9 a_n3110_n2688# 0.387196f
C252 plus.n10 a_n3110_n2688# 0.149518f
C253 plus.n11 a_n3110_n2688# 0.035847f
C254 plus.n12 a_n3110_n2688# 0.032833f
C255 plus.n13 a_n3110_n2688# 0.050065f
C256 plus.n14 a_n3110_n2688# 0.334193f
C257 plus.n15 a_n3110_n2688# 0.05006f
C258 plus.n16 a_n3110_n2688# 0.035847f
C259 plus.n17 a_n3110_n2688# 0.035847f
C260 plus.n18 a_n3110_n2688# 0.035847f
C261 plus.n19 a_n3110_n2688# 0.04467f
C262 plus.n20 a_n3110_n2688# 0.334193f
C263 plus.n21 a_n3110_n2688# 0.04653f
C264 plus.t6 a_n3110_n2688# 0.870642f
C265 plus.n22 a_n3110_n2688# 0.334193f
C266 plus.n23 a_n3110_n2688# 0.04653f
C267 plus.n24 a_n3110_n2688# 0.035847f
C268 plus.n25 a_n3110_n2688# 0.035847f
C269 plus.n26 a_n3110_n2688# 0.035847f
C270 plus.n27 a_n3110_n2688# 0.031987f
C271 plus.n28 a_n3110_n2688# 0.05006f
C272 plus.n29 a_n3110_n2688# 0.334193f
C273 plus.n30 a_n3110_n2688# 0.050065f
C274 plus.n31 a_n3110_n2688# 0.035847f
C275 plus.n32 a_n3110_n2688# 0.035847f
C276 plus.n33 a_n3110_n2688# 0.035847f
C277 plus.n34 a_n3110_n2688# 0.043819f
C278 plus.n35 a_n3110_n2688# 0.334193f
C279 plus.n36 a_n3110_n2688# 0.045005f
C280 plus.n37 a_n3110_n2688# 0.387903f
C281 plus.n38 a_n3110_n2688# 0.39447f
C282 plus.n39 a_n3110_n2688# 0.047833f
C283 plus.t1 a_n3110_n2688# 0.925225f
C284 plus.t9 a_n3110_n2688# 0.870642f
C285 plus.n40 a_n3110_n2688# 0.032833f
C286 plus.n41 a_n3110_n2688# 0.035847f
C287 plus.t12 a_n3110_n2688# 0.870642f
C288 plus.n42 a_n3110_n2688# 0.04467f
C289 plus.n43 a_n3110_n2688# 0.035847f
C290 plus.t7 a_n3110_n2688# 0.870642f
C291 plus.n44 a_n3110_n2688# 0.334193f
C292 plus.t10 a_n3110_n2688# 0.870642f
C293 plus.n45 a_n3110_n2688# 0.031987f
C294 plus.n46 a_n3110_n2688# 0.035847f
C295 plus.t15 a_n3110_n2688# 0.870642f
C296 plus.n47 a_n3110_n2688# 0.043819f
C297 plus.t13 a_n3110_n2688# 0.945708f
C298 plus.t11 a_n3110_n2688# 0.870642f
C299 plus.n48 a_n3110_n2688# 0.36014f
C300 plus.n49 a_n3110_n2688# 0.387196f
C301 plus.n50 a_n3110_n2688# 0.149518f
C302 plus.n51 a_n3110_n2688# 0.035847f
C303 plus.n52 a_n3110_n2688# 0.032833f
C304 plus.n53 a_n3110_n2688# 0.050065f
C305 plus.n54 a_n3110_n2688# 0.334193f
C306 plus.n55 a_n3110_n2688# 0.05006f
C307 plus.n56 a_n3110_n2688# 0.035847f
C308 plus.n57 a_n3110_n2688# 0.035847f
C309 plus.n58 a_n3110_n2688# 0.035847f
C310 plus.n59 a_n3110_n2688# 0.04467f
C311 plus.n60 a_n3110_n2688# 0.334193f
C312 plus.n61 a_n3110_n2688# 0.04653f
C313 plus.n62 a_n3110_n2688# 0.04653f
C314 plus.n63 a_n3110_n2688# 0.035847f
C315 plus.n64 a_n3110_n2688# 0.035847f
C316 plus.n65 a_n3110_n2688# 0.035847f
C317 plus.n66 a_n3110_n2688# 0.031987f
C318 plus.n67 a_n3110_n2688# 0.05006f
C319 plus.n68 a_n3110_n2688# 0.334193f
C320 plus.n69 a_n3110_n2688# 0.050065f
C321 plus.n70 a_n3110_n2688# 0.035847f
C322 plus.n71 a_n3110_n2688# 0.035847f
C323 plus.n72 a_n3110_n2688# 0.035847f
C324 plus.n73 a_n3110_n2688# 0.043819f
C325 plus.n74 a_n3110_n2688# 0.334193f
C326 plus.n75 a_n3110_n2688# 0.045005f
C327 plus.n76 a_n3110_n2688# 0.387903f
C328 plus.n77 a_n3110_n2688# 1.27239f
.ends

