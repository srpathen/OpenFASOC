* NGSPICE file created from opamp614.ext - technology: sky130A

.subckt opamp614 gnd CSoutput output vdd plus minus commonsourceibias outputibias
+ diffpairibias
X0 gnd.t307 commonsourceibias.t64 CSoutput.t102 gnd.t190 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X1 a_n7636_8799.t22 plus.t5 a_n2903_n3924.t23 gnd.t136 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.7
X2 CSoutput.t4 a_n7636_8799.t32 vdd.t170 vdd.t109 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X3 commonsourceibias.t7 commonsourceibias.t6 gnd.t306 gnd.t277 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X4 a_n1808_13878.t19 a_n1996_n452.t44 vdd.t291 vdd.t290 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X5 a_n1808_13878.t11 a_n1996_n452.t15 a_n1996_n452.t16 vdd.t171 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X6 CSoutput.t184 a_n1986_8322.t21 sky130_fd_pr__cap_mim_m3_1 l=12 w=12
X7 vdd.t169 a_n7636_8799.t33 CSoutput.t6 vdd.t104 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X8 CSoutput.t23 a_n7636_8799.t34 vdd.t168 vdd.t23 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X9 gnd.t124 gnd.t122 plus.t4 gnd.t123 sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.5
X10 CSoutput.t43 a_n7636_8799.t35 vdd.t167 vdd.t25 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X11 a_n2903_n3924.t12 plus.t6 a_n7636_8799.t21 gnd.t128 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.7
X12 gnd.t305 commonsourceibias.t65 CSoutput.t101 gnd.t272 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X13 gnd.t121 gnd.t119 gnd.t120 gnd.t18 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=0 ps=0 w=7 l=1
X14 gnd.t304 commonsourceibias.t4 commonsourceibias.t5 gnd.t184 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X15 gnd.t303 commonsourceibias.t66 CSoutput.t100 gnd.t184 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X16 vdd.t281 vdd.t279 vdd.t280 vdd.t233 sky130_fd_pr__pfet_01v8 ad=3.12 pd=16.78 as=0 ps=0 w=8 l=0.5
X17 a_n2903_n3924.t45 minus.t5 a_n1996_n452.t43 gnd.t4 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=1.155 ps=7.33 w=7 l=0.7
X18 a_n1986_8322.t11 a_n1996_n452.t45 a_n7636_8799.t2 vdd.t6 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X19 output.t17 CSoutput.t185 vdd.t183 gnd.t165 sky130_fd_pr__nfet_01v8 ad=0.825 pd=5.33 as=0.825 ps=5.33 w=5 l=1
X20 CSoutput.t60 a_n7636_8799.t36 vdd.t166 vdd.t68 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X21 gnd.t302 commonsourceibias.t67 CSoutput.t99 gnd.t213 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X22 vdd.t165 a_n7636_8799.t37 CSoutput.t67 vdd.t97 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X23 a_n1996_n452.t5 minus.t6 a_n2903_n3924.t7 gnd.t6 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.7
X24 gnd.t301 commonsourceibias.t2 commonsourceibias.t3 gnd.t226 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X25 vdd.t164 a_n7636_8799.t38 CSoutput.t18 vdd.t124 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X26 a_n1996_n452.t1 minus.t7 a_n2903_n3924.t3 gnd.t13 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.7
X27 CSoutput.t75 a_n7636_8799.t39 vdd.t163 vdd.t70 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X28 vdd.t162 a_n7636_8799.t40 CSoutput.t73 vdd.t121 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X29 vdd.t161 a_n7636_8799.t41 CSoutput.t55 vdd.t148 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X30 output.t0 outputibias.t8 gnd.t140 gnd.t139 sky130_fd_pr__nfet_01v8 ad=2.34 pd=12.78 as=2.34 ps=12.78 w=6 l=2
X31 CSoutput.t186 a_n1986_8322.t20 sky130_fd_pr__cap_mim_m3_1 l=12 w=12
X32 a_n7636_8799.t24 a_n1996_n452.t46 a_n1986_8322.t10 vdd.t178 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=3.51 ps=18.78 w=9 l=0.5
X33 CSoutput.t1 a_n7636_8799.t42 vdd.t160 vdd.t17 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=3.12 ps=16.78 w=8 l=0.5
X34 CSoutput.t98 commonsourceibias.t68 gnd.t300 gnd.t182 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X35 gnd.t118 gnd.t116 gnd.t117 gnd.t64 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=0 ps=0 w=7 l=1
X36 a_n2903_n3924.t32 minus.t8 a_n1996_n452.t32 gnd.t7 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=1.155 ps=7.33 w=7 l=0.7
X37 gnd.t299 commonsourceibias.t0 commonsourceibias.t1 gnd.t268 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X38 output.t1 outputibias.t9 gnd.t145 gnd.t144 sky130_fd_pr__nfet_01v8 ad=2.34 pd=12.78 as=2.34 ps=12.78 w=6 l=2
X39 CSoutput.t93 a_n7636_8799.t43 vdd.t159 vdd.t109 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X40 vdd.t184 CSoutput.t187 output.t16 gnd.t164 sky130_fd_pr__nfet_01v8 ad=0.825 pd=5.33 as=0.825 ps=5.33 w=5 l=1
X41 vdd.t278 vdd.t276 vdd.t277 vdd.t211 sky130_fd_pr__pfet_01v8 ad=3.12 pd=16.78 as=0 ps=0 w=8 l=0.5
X42 CSoutput.t111 commonsourceibias.t69 gnd.t298 gnd.t196 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X43 a_n2903_n3924.t37 diffpairibias.t16 gnd.t175 gnd.t174 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=2.73 ps=14.78 w=7 l=1
X44 CSoutput.t175 a_n7636_8799.t44 vdd.t158 vdd.t62 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X45 output.t19 outputibias.t10 gnd.t311 gnd.t310 sky130_fd_pr__nfet_01v8 ad=2.34 pd=12.78 as=2.34 ps=12.78 w=6 l=2
X46 CSoutput.t110 commonsourceibias.t70 gnd.t297 gnd.t192 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X47 CSoutput.t16 a_n7636_8799.t45 vdd.t157 vdd.t25 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X48 a_n2903_n3924.t26 plus.t7 a_n7636_8799.t20 gnd.t143 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.7
X49 output.t15 CSoutput.t188 vdd.t185 gnd.t163 sky130_fd_pr__nfet_01v8 ad=1.95 pd=10.78 as=0.825 ps=5.33 w=5 l=1
X50 gnd.t296 commonsourceibias.t14 commonsourceibias.t15 gnd.t234 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=1.155 ps=7.33 w=7 l=1
X51 vdd.t156 a_n7636_8799.t46 CSoutput.t25 vdd.t148 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X52 vdd.t275 vdd.t273 vdd.t274 vdd.t233 sky130_fd_pr__pfet_01v8 ad=3.12 pd=16.78 as=0 ps=0 w=8 l=0.5
X53 a_n1808_13878.t10 a_n1996_n452.t29 a_n1996_n452.t30 vdd.t176 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=3.51 ps=18.78 w=9 l=0.5
X54 CSoutput.t109 commonsourceibias.t71 gnd.t295 gnd.t277 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X55 CSoutput.t33 a_n7636_8799.t47 vdd.t155 vdd.t102 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X56 a_n1996_n452.t26 a_n1996_n452.t25 a_n1808_13878.t9 vdd.t1 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X57 a_n7636_8799.t19 plus.t8 a_n2903_n3924.t28 gnd.t130 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.7
X58 CSoutput.t179 a_n7636_8799.t48 vdd.t154 vdd.t68 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X59 vdd.t272 vdd.t270 vdd.t271 vdd.t246 sky130_fd_pr__pfet_01v8 ad=3.51 pd=18.78 as=0 ps=0 w=9 l=0.5
X60 vdd.t153 a_n7636_8799.t49 CSoutput.t183 vdd.t97 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X61 diffpairibias.t15 diffpairibias.t14 gnd.t177 gnd.t176 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=2.73 ps=14.78 w=7 l=1
X62 a_n1996_n452.t0 minus.t9 a_n2903_n3924.t1 gnd.t3 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.7
X63 CSoutput.t27 a_n7636_8799.t50 vdd.t152 vdd.t106 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X64 vdd.t151 a_n7636_8799.t51 CSoutput.t20 vdd.t35 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X65 vdd.t150 a_n7636_8799.t52 CSoutput.t85 vdd.t121 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X66 vdd.t149 a_n7636_8799.t53 CSoutput.t182 vdd.t148 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X67 gnd.t294 commonsourceibias.t72 CSoutput.t108 gnd.t272 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X68 plus.t3 gnd.t113 gnd.t115 gnd.t114 sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.5
X69 vdd.t147 a_n7636_8799.t54 CSoutput.t10 vdd.t94 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X70 diffpairibias.t13 diffpairibias.t12 gnd.t168 gnd.t167 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=2.73 ps=14.78 w=7 l=1
X71 gnd.t293 commonsourceibias.t73 CSoutput.t107 gnd.t180 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X72 CSoutput.t56 a_n7636_8799.t55 vdd.t146 vdd.t17 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=3.12 ps=16.78 w=8 l=0.5
X73 CSoutput.t58 a_n7636_8799.t56 vdd.t145 vdd.t42 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X74 output.t14 CSoutput.t189 vdd.t193 gnd.t162 sky130_fd_pr__nfet_01v8 ad=0.825 pd=5.33 as=0.825 ps=5.33 w=5 l=1
X75 commonsourceibias.t13 commonsourceibias.t12 gnd.t292 gnd.t182 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X76 vdd.t197 CSoutput.t190 output.t13 gnd.t161 sky130_fd_pr__nfet_01v8 ad=0.825 pd=5.33 as=1.95 ps=10.78 w=5 l=1
X77 gnd.t112 gnd.t110 gnd.t111 gnd.t43 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=0 ps=0 w=7 l=0.7
X78 gnd.t291 commonsourceibias.t74 CSoutput.t106 gnd.t268 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X79 vdd.t144 a_n7636_8799.t57 CSoutput.t168 vdd.t19 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X80 CSoutput.t51 a_n7636_8799.t58 vdd.t143 vdd.t129 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X81 CSoutput.t170 a_n7636_8799.t59 vdd.t142 vdd.t62 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X82 CSoutput.t14 a_n7636_8799.t60 vdd.t141 vdd.t79 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=3.12 ps=16.78 w=8 l=0.5
X83 commonsourceibias.t11 commonsourceibias.t10 gnd.t290 gnd.t228 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X84 gnd.t289 commonsourceibias.t75 CSoutput.t105 gnd.t213 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X85 CSoutput.t65 a_n7636_8799.t61 vdd.t140 vdd.t129 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X86 CSoutput.t191 a_n1986_8322.t20 sky130_fd_pr__cap_mim_m3_1 l=12 w=12
X87 vdd.t139 a_n7636_8799.t62 CSoutput.t78 vdd.t126 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X88 commonsourceibias.t9 commonsourceibias.t8 gnd.t288 gnd.t215 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X89 gnd.t287 commonsourceibias.t76 CSoutput.t104 gnd.t265 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X90 a_n2903_n3924.t25 plus.t9 a_n7636_8799.t18 gnd.t125 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.7
X91 CSoutput.t103 commonsourceibias.t77 gnd.t286 gnd.t262 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=2.73 ps=14.78 w=7 l=1
X92 gnd.t285 commonsourceibias.t36 commonsourceibias.t37 gnd.t265 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X93 a_n2903_n3924.t8 diffpairibias.t17 gnd.t127 gnd.t126 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=2.73 ps=14.78 w=7 l=1
X94 vdd.t138 a_n7636_8799.t63 CSoutput.t17 vdd.t91 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X95 a_n1996_n452.t18 a_n1996_n452.t17 a_n1808_13878.t8 vdd.t6 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X96 vdd.t137 a_n7636_8799.t64 CSoutput.t35 vdd.t72 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X97 a_n7636_8799.t26 a_n1996_n452.t47 a_n1986_8322.t9 vdd.t199 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X98 vdd.t136 a_n7636_8799.t65 CSoutput.t47 vdd.t124 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X99 a_n1996_n452.t20 a_n1996_n452.t19 a_n1808_13878.t7 vdd.t177 sky130_fd_pr__pfet_01v8 ad=3.51 pd=18.78 as=1.485 ps=9.33 w=9 l=0.5
X100 gnd.t284 commonsourceibias.t34 commonsourceibias.t35 gnd.t255 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=1.155 ps=7.33 w=7 l=1
X101 vdd.t135 a_n7636_8799.t66 CSoutput.t90 vdd.t126 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X102 gnd.t109 gnd.t107 gnd.t108 gnd.t64 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=0 ps=0 w=7 l=1
X103 commonsourceibias.t33 commonsourceibias.t32 gnd.t283 gnd.t192 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X104 CSoutput.t120 commonsourceibias.t78 gnd.t282 gnd.t196 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X105 vdd.t134 a_n7636_8799.t67 CSoutput.t24 vdd.t39 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X106 CSoutput.t48 a_n7636_8799.t68 vdd.t133 vdd.t76 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X107 CSoutput.t149 commonsourceibias.t79 gnd.t253 gnd.t251 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X108 vdd.t196 CSoutput.t192 output.t12 gnd.t160 sky130_fd_pr__nfet_01v8 ad=0.825 pd=5.33 as=0.825 ps=5.33 w=5 l=1
X109 a_n1996_n452.t2 minus.t10 a_n2903_n3924.t4 gnd.t14 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.7
X110 vdd.t269 vdd.t267 vdd.t268 vdd.t254 sky130_fd_pr__pfet_01v8 ad=3.51 pd=18.78 as=0 ps=0 w=9 l=0.5
X111 vdd.t132 a_n7636_8799.t69 CSoutput.t165 vdd.t94 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X112 CSoutput.t119 commonsourceibias.t80 gnd.t281 gnd.t257 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X113 CSoutput.t181 a_n7636_8799.t70 vdd.t131 vdd.t42 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X114 vdd.t266 vdd.t263 vdd.t265 vdd.t264 sky130_fd_pr__pfet_01v8 ad=3.51 pd=18.78 as=0 ps=0 w=9 l=0.5
X115 gnd.t280 commonsourceibias.t81 CSoutput.t118 gnd.t255 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=1.155 ps=7.33 w=7 l=1
X116 commonsourceibias.t31 commonsourceibias.t30 gnd.t279 gnd.t211 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X117 a_n2903_n3924.t6 minus.t11 a_n1996_n452.t4 gnd.t5 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.7
X118 CSoutput.t117 commonsourceibias.t82 gnd.t278 gnd.t277 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X119 vdd.t262 vdd.t260 vdd.t261 vdd.t207 sky130_fd_pr__pfet_01v8 ad=3.51 pd=18.78 as=0 ps=0 w=9 l=0.5
X120 CSoutput.t193 a_n1986_8322.t21 sky130_fd_pr__cap_mim_m3_1 l=12 w=12
X121 vdd.t259 vdd.t257 vdd.t258 vdd.t250 sky130_fd_pr__pfet_01v8 ad=3.51 pd=18.78 as=0 ps=0 w=9 l=0.5
X122 vdd.t173 a_n1996_n452.t48 a_n1986_8322.t19 vdd.t172 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X123 a_n1986_8322.t18 a_n1996_n452.t49 vdd.t295 vdd.t294 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X124 a_n2903_n3924.t2 diffpairibias.t18 gnd.t10 gnd.t9 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=2.73 ps=14.78 w=7 l=1
X125 CSoutput.t42 a_n7636_8799.t71 vdd.t130 vdd.t129 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X126 CSoutput.t3 a_n7636_8799.t72 vdd.t128 vdd.t79 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=3.12 ps=16.78 w=8 l=0.5
X127 output.t18 outputibias.t11 gnd.t173 gnd.t172 sky130_fd_pr__nfet_01v8 ad=2.34 pd=12.78 as=2.34 ps=12.78 w=6 l=2
X128 gnd.t106 gnd.t104 gnd.t105 gnd.t25 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=0 ps=0 w=7 l=0.7
X129 gnd.t276 commonsourceibias.t83 CSoutput.t116 gnd.t232 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X130 vdd.t127 a_n7636_8799.t73 CSoutput.t72 vdd.t126 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X131 a_n2903_n3924.t39 minus.t12 a_n1996_n452.t37 gnd.t166 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.7
X132 CSoutput.t194 a_n1986_8322.t21 sky130_fd_pr__cap_mim_m3_1 l=12 w=12
X133 commonsourceibias.t29 commonsourceibias.t28 gnd.t275 gnd.t257 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X134 vdd.t8 a_n1996_n452.t50 a_n1808_13878.t18 vdd.t7 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X135 a_n1996_n452.t3 minus.t13 a_n2903_n3924.t5 gnd.t2 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=2.73 ps=14.78 w=7 l=0.7
X136 a_n2903_n3924.t24 plus.t10 a_n7636_8799.t17 gnd.t8 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.7
X137 a_n2903_n3924.t27 plus.t11 a_n7636_8799.t16 gnd.t169 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.7
X138 vdd.t256 vdd.t253 vdd.t255 vdd.t254 sky130_fd_pr__pfet_01v8 ad=3.51 pd=18.78 as=0 ps=0 w=9 l=0.5
X139 gnd.t274 commonsourceibias.t84 CSoutput.t115 gnd.t180 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X140 vdd.t125 a_n7636_8799.t74 CSoutput.t9 vdd.t124 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X141 vdd.t252 vdd.t249 vdd.t251 vdd.t250 sky130_fd_pr__pfet_01v8 ad=3.51 pd=18.78 as=0 ps=0 w=9 l=0.5
X142 gnd.t273 commonsourceibias.t26 commonsourceibias.t27 gnd.t272 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X143 a_n7636_8799.t15 plus.t12 a_n2903_n3924.t18 gnd.t129 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.7
X144 a_n7636_8799.t14 plus.t13 a_n2903_n3924.t16 gnd.t131 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=2.73 ps=14.78 w=7 l=0.7
X145 vdd.t248 vdd.t245 vdd.t247 vdd.t246 sky130_fd_pr__pfet_01v8 ad=3.51 pd=18.78 as=0 ps=0 w=9 l=0.5
X146 a_n1986_8322.t17 a_n1996_n452.t51 vdd.t203 vdd.t202 sky130_fd_pr__pfet_01v8 ad=3.51 pd=18.78 as=1.485 ps=9.33 w=9 l=0.5
X147 commonsourceibias.t41 commonsourceibias.t40 gnd.t271 gnd.t219 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X148 gnd.t270 commonsourceibias.t85 CSoutput.t128 gnd.t222 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X149 gnd.t269 commonsourceibias.t86 CSoutput.t127 gnd.t268 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X150 a_n7636_8799.t29 a_n1996_n452.t52 a_n1986_8322.t8 vdd.t3 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X151 CSoutput.t41 a_n7636_8799.t75 vdd.t123 vdd.t53 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X152 diffpairibias.t11 diffpairibias.t10 gnd.t12 gnd.t11 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=2.73 ps=14.78 w=7 l=1
X153 vdd.t122 a_n7636_8799.t76 CSoutput.t79 vdd.t121 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X154 a_n1996_n452.t35 minus.t14 a_n2903_n3924.t36 gnd.t135 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.7
X155 a_n1996_n452.t8 a_n1996_n452.t7 a_n1808_13878.t6 vdd.t0 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X156 vdd.t120 a_n7636_8799.t77 CSoutput.t87 vdd.t39 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X157 a_n7636_8799.t25 a_n1996_n452.t53 a_n1986_8322.t7 vdd.t171 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X158 CSoutput.t62 a_n7636_8799.t78 vdd.t119 vdd.t76 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X159 gnd.t103 gnd.t100 gnd.t102 gnd.t101 sky130_fd_pr__nfet_01v8 ad=2.34 pd=12.78 as=0 ps=0 w=6 l=2
X160 gnd.t267 commonsourceibias.t87 CSoutput.t126 gnd.t240 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X161 a_n1808_13878.t5 a_n1996_n452.t11 a_n1996_n452.t12 vdd.t199 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X162 gnd.t99 gnd.t97 minus.t4 gnd.t98 sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.39 ps=2.78 w=1 l=0.5
X163 a_n2903_n3924.t42 minus.t15 a_n1996_n452.t40 gnd.t132 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.7
X164 gnd.t266 commonsourceibias.t88 CSoutput.t125 gnd.t265 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X165 CSoutput.t124 commonsourceibias.t89 gnd.t264 gnd.t262 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=2.73 ps=14.78 w=7 l=1
X166 commonsourceibias.t39 commonsourceibias.t38 gnd.t263 gnd.t262 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=2.73 ps=14.78 w=7 l=1
X167 CSoutput.t12 a_n7636_8799.t79 vdd.t118 vdd.t106 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X168 vdd.t175 a_n1996_n452.t54 a_n1986_8322.t16 vdd.t174 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=3.51 ps=18.78 w=9 l=0.5
X169 CSoutput.t123 commonsourceibias.t90 gnd.t261 gnd.t203 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X170 vdd.t117 a_n7636_8799.t80 CSoutput.t68 vdd.t104 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X171 CSoutput.t94 a_n7636_8799.t81 vdd.t116 vdd.t102 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X172 vdd.t115 a_n7636_8799.t82 CSoutput.t44 vdd.t13 sky130_fd_pr__pfet_01v8 ad=3.12 pd=16.78 as=1.32 ps=8.33 w=8 l=0.5
X173 a_n2903_n3924.t22 plus.t14 a_n7636_8799.t13 gnd.t4 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=1.155 ps=7.33 w=7 l=0.7
X174 gnd.t96 gnd.t94 minus.t3 gnd.t95 sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.5
X175 vdd.t114 a_n7636_8799.t83 CSoutput.t36 vdd.t55 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X176 CSoutput.t122 commonsourceibias.t91 gnd.t260 gnd.t251 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X177 a_n2903_n3924.t35 diffpairibias.t19 gnd.t171 gnd.t170 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=2.73 ps=14.78 w=7 l=1
X178 gnd.t93 gnd.t90 gnd.t92 gnd.t91 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=0 ps=0 w=7 l=1
X179 a_n2903_n3924.t0 diffpairibias.t20 gnd.t1 gnd.t0 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=2.73 ps=14.78 w=7 l=1
X180 vdd.t195 CSoutput.t195 output.t11 gnd.t159 sky130_fd_pr__nfet_01v8 ad=0.825 pd=5.33 as=0.825 ps=5.33 w=5 l=1
X181 CSoutput.t121 commonsourceibias.t92 gnd.t259 gnd.t188 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X182 CSoutput.t152 commonsourceibias.t93 gnd.t258 gnd.t257 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X183 vdd.t113 a_n7636_8799.t84 CSoutput.t84 vdd.t91 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X184 a_n7636_8799.t12 plus.t15 a_n2903_n3924.t13 gnd.t6 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.7
X185 vdd.t112 a_n7636_8799.t85 CSoutput.t39 vdd.t60 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X186 gnd.t256 commonsourceibias.t94 CSoutput.t151 gnd.t255 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=1.155 ps=7.33 w=7 l=1
X187 gnd.t254 commonsourceibias.t95 CSoutput.t150 gnd.t234 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=1.155 ps=7.33 w=7 l=1
X188 commonsourceibias.t61 commonsourceibias.t60 gnd.t252 gnd.t251 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X189 CSoutput.t148 commonsourceibias.t96 gnd.t250 gnd.t209 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X190 CSoutput.t22 a_n7636_8799.t86 vdd.t111 vdd.t15 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X191 gnd.t249 commonsourceibias.t97 CSoutput.t147 gnd.t232 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X192 CSoutput.t7 a_n7636_8799.t87 vdd.t110 vdd.t109 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X193 CSoutput.t30 a_n7636_8799.t88 vdd.t108 vdd.t86 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X194 gnd.t89 gnd.t87 gnd.t88 gnd.t50 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=0 ps=0 w=7 l=1
X195 CSoutput.t146 commonsourceibias.t98 gnd.t248 gnd.t228 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X196 diffpairibias.t9 diffpairibias.t8 gnd.t309 gnd.t308 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=2.73 ps=14.78 w=7 l=1
X197 a_n1808_13878.t17 a_n1996_n452.t55 vdd.t5 vdd.t4 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X198 vdd.t287 a_n1996_n452.t56 a_n1808_13878.t16 vdd.t286 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X199 vdd.t244 vdd.t242 vdd.t243 vdd.t218 sky130_fd_pr__pfet_01v8 ad=3.12 pd=16.78 as=0 ps=0 w=8 l=0.5
X200 vdd.t241 vdd.t239 vdd.t240 vdd.t226 sky130_fd_pr__pfet_01v8 ad=3.12 pd=16.78 as=0 ps=0 w=8 l=0.5
X201 CSoutput.t26 a_n7636_8799.t89 vdd.t107 vdd.t106 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X202 vdd.t105 a_n7636_8799.t90 CSoutput.t166 vdd.t104 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X203 vdd.t238 vdd.t236 vdd.t237 vdd.t226 sky130_fd_pr__pfet_01v8 ad=3.12 pd=16.78 as=0 ps=0 w=8 l=0.5
X204 gnd.t247 commonsourceibias.t99 CSoutput.t145 gnd.t226 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X205 CSoutput.t144 commonsourceibias.t100 gnd.t246 gnd.t186 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=2.73 ps=14.78 w=7 l=1
X206 gnd.t245 commonsourceibias.t58 commonsourceibias.t59 gnd.t201 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X207 gnd.t244 commonsourceibias.t101 CSoutput.t136 gnd.t222 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X208 a_n2903_n3924.t33 minus.t16 a_n1996_n452.t33 gnd.t143 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.7
X209 CSoutput.t53 a_n7636_8799.t91 vdd.t103 vdd.t102 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X210 vdd.t101 a_n7636_8799.t92 CSoutput.t64 vdd.t13 sky130_fd_pr__pfet_01v8 ad=3.12 pd=16.78 as=1.32 ps=8.33 w=8 l=0.5
X211 vdd.t100 a_n7636_8799.t93 CSoutput.t163 vdd.t55 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X212 gnd.t243 commonsourceibias.t102 CSoutput.t135 gnd.t240 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X213 a_n1986_8322.t6 a_n1996_n452.t57 a_n7636_8799.t30 vdd.t204 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X214 vdd.t191 CSoutput.t196 output.t10 gnd.t158 sky130_fd_pr__nfet_01v8 ad=0.825 pd=5.33 as=0.825 ps=5.33 w=5 l=1
X215 CSoutput.t34 a_n7636_8799.t94 vdd.t99 vdd.t57 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X216 diffpairibias.t7 diffpairibias.t6 gnd.t142 gnd.t141 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=2.73 ps=14.78 w=7 l=1
X217 CSoutput.t134 commonsourceibias.t103 gnd.t242 gnd.t219 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X218 vdd.t98 a_n7636_8799.t95 CSoutput.t82 vdd.t97 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X219 a_n1996_n452.t36 minus.t17 a_n2903_n3924.t38 gnd.t130 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.7
X220 CSoutput.t50 a_n7636_8799.t96 vdd.t96 vdd.t31 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X221 a_n1996_n452.t34 minus.t18 a_n2903_n3924.t34 gnd.t136 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.7
X222 vdd.t95 a_n7636_8799.t97 CSoutput.t45 vdd.t94 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X223 plus.t2 gnd.t84 gnd.t86 gnd.t85 sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.5
X224 vdd.t182 a_n1996_n452.t58 a_n1986_8322.t15 vdd.t181 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=3.51 ps=18.78 w=9 l=0.5
X225 gnd.t241 commonsourceibias.t46 commonsourceibias.t47 gnd.t240 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X226 gnd.t83 gnd.t80 gnd.t82 gnd.t81 sky130_fd_pr__nfet_01v8 ad=1.95 pd=10.78 as=0 ps=0 w=5 l=1
X227 vdd.t93 a_n7636_8799.t98 CSoutput.t88 vdd.t60 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X228 vdd.t92 a_n7636_8799.t99 CSoutput.t63 vdd.t91 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X229 gnd.t72 gnd.t70 gnd.t71 gnd.t50 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=0 ps=0 w=7 l=1
X230 CSoutput.t133 commonsourceibias.t104 gnd.t239 gnd.t215 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X231 a_n7636_8799.t11 plus.t16 a_n2903_n3924.t30 gnd.t3 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.7
X232 gnd.t79 gnd.t77 minus.t2 gnd.t78 sky130_fd_pr__nfet_01v8 ad=0.39 pd=2.78 as=0.165 ps=1.33 w=1 l=0.5
X233 a_n2903_n3924.t10 minus.t19 a_n1996_n452.t31 gnd.t128 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.7
X234 CSoutput.t132 commonsourceibias.t105 gnd.t238 gnd.t203 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X235 a_n1808_13878.t15 a_n1996_n452.t59 vdd.t10 vdd.t9 sky130_fd_pr__pfet_01v8 ad=3.51 pd=18.78 as=1.485 ps=9.33 w=9 l=0.5
X236 vdd.t90 a_n7636_8799.t100 CSoutput.t32 vdd.t72 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X237 CSoutput.t74 a_n7636_8799.t101 vdd.t89 vdd.t86 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X238 CSoutput.t29 a_n7636_8799.t102 vdd.t88 vdd.t70 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X239 gnd.t237 commonsourceibias.t44 commonsourceibias.t45 gnd.t206 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X240 vdd.t235 vdd.t232 vdd.t234 vdd.t233 sky130_fd_pr__pfet_01v8 ad=3.12 pd=16.78 as=0 ps=0 w=8 l=0.5
X241 gnd.t76 gnd.t73 gnd.t75 gnd.t74 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=0 ps=0 w=7 l=1
X242 minus.t1 gnd.t67 gnd.t69 gnd.t68 sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.5
X243 vdd.t231 vdd.t229 vdd.t230 vdd.t218 sky130_fd_pr__pfet_01v8 ad=3.12 pd=16.78 as=0 ps=0 w=8 l=0.5
X244 a_n2903_n3924.t31 diffpairibias.t21 gnd.t138 gnd.t137 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=2.73 ps=14.78 w=7 l=1
X245 gnd.t66 gnd.t63 gnd.t65 gnd.t64 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=0 ps=0 w=7 l=1
X246 CSoutput.t157 commonsourceibias.t106 gnd.t224 gnd.t211 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X247 vdd.t228 vdd.t225 vdd.t227 vdd.t226 sky130_fd_pr__pfet_01v8 ad=3.12 pd=16.78 as=0 ps=0 w=8 l=0.5
X248 vdd.t283 a_n1996_n452.t60 a_n1986_8322.t14 vdd.t282 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X249 a_n1986_8322.t5 a_n1996_n452.t61 a_n7636_8799.t28 vdd.t0 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X250 CSoutput.t164 a_n7636_8799.t103 vdd.t87 vdd.t86 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X251 vdd.t85 a_n7636_8799.t104 CSoutput.t40 vdd.t11 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X252 CSoutput.t52 a_n7636_8799.t105 vdd.t84 vdd.t37 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X253 CSoutput.t131 commonsourceibias.t107 gnd.t236 gnd.t188 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X254 vdd.t83 a_n7636_8799.t106 CSoutput.t86 vdd.t65 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X255 gnd.t235 commonsourceibias.t108 CSoutput.t130 gnd.t234 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=1.155 ps=7.33 w=7 l=1
X256 vdd.t82 a_n7636_8799.t107 CSoutput.t169 vdd.t29 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X257 gnd.t233 commonsourceibias.t42 commonsourceibias.t43 gnd.t232 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X258 a_n7636_8799.t10 plus.t17 a_n2903_n3924.t11 gnd.t13 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.7
X259 gnd.t62 gnd.t59 gnd.t61 gnd.t60 sky130_fd_pr__nfet_01v8 ad=2.34 pd=12.78 as=0 ps=0 w=6 l=2
X260 CSoutput.t129 commonsourceibias.t109 gnd.t231 gnd.t209 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X261 output.t9 CSoutput.t197 vdd.t192 gnd.t157 sky130_fd_pr__nfet_01v8 ad=0.825 pd=5.33 as=0.825 ps=5.33 w=5 l=1
X262 gnd.t230 commonsourceibias.t110 CSoutput.t161 gnd.t206 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X263 vdd.t224 vdd.t221 vdd.t223 vdd.t222 sky130_fd_pr__pfet_01v8 ad=3.51 pd=18.78 as=0 ps=0 w=9 l=0.5
X264 a_n2903_n3924.t14 plus.t18 a_n7636_8799.t9 gnd.t7 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=1.155 ps=7.33 w=7 l=0.7
X265 gnd.t58 gnd.t56 gnd.t57 gnd.t32 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=0 ps=0 w=7 l=1
X266 vdd.t81 a_n7636_8799.t108 CSoutput.t37 vdd.t21 sky130_fd_pr__pfet_01v8 ad=3.12 pd=16.78 as=1.32 ps=8.33 w=8 l=0.5
X267 CSoutput.t80 a_n7636_8799.t109 vdd.t80 vdd.t79 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=3.12 ps=16.78 w=8 l=0.5
X268 outputibias.t7 outputibias.t6 gnd.t16 gnd.t15 sky130_fd_pr__nfet_01v8 ad=2.34 pd=12.78 as=2.34 ps=12.78 w=6 l=2
X269 a_n1808_13878.t4 a_n1996_n452.t13 a_n1996_n452.t14 vdd.t205 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X270 CSoutput.t19 a_n7636_8799.t110 vdd.t78 vdd.t57 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X271 gnd.t55 gnd.t53 gnd.t54 gnd.t32 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=0 ps=0 w=7 l=1
X272 CSoutput.t160 commonsourceibias.t111 gnd.t229 gnd.t228 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X273 a_n1986_8322.t4 a_n1996_n452.t62 a_n7636_8799.t1 vdd.t1 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X274 diffpairibias.t5 diffpairibias.t4 gnd.t315 gnd.t314 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=2.73 ps=14.78 w=7 l=1
X275 outputibias.t5 outputibias.t4 gnd.t147 gnd.t146 sky130_fd_pr__nfet_01v8 ad=2.34 pd=12.78 as=2.34 ps=12.78 w=6 l=2
X276 CSoutput.t13 a_n7636_8799.t111 vdd.t77 vdd.t76 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X277 CSoutput.t97 a_n7636_8799.t112 vdd.t75 vdd.t53 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X278 vdd.t74 a_n7636_8799.t113 CSoutput.t76 vdd.t65 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X279 gnd.t227 commonsourceibias.t112 CSoutput.t159 gnd.t226 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X280 CSoutput.t158 commonsourceibias.t113 gnd.t225 gnd.t186 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=2.73 ps=14.78 w=7 l=1
X281 vdd.t73 a_n7636_8799.t114 CSoutput.t66 vdd.t72 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X282 outputibias.t3 outputibias.t2 gnd.t134 gnd.t133 sky130_fd_pr__nfet_01v8 ad=2.34 pd=12.78 as=2.34 ps=12.78 w=6 l=2
X283 output.t8 CSoutput.t198 vdd.t198 gnd.t156 sky130_fd_pr__nfet_01v8 ad=0.825 pd=5.33 as=0.825 ps=5.33 w=5 l=1
X284 a_n1986_8322.t13 a_n1996_n452.t63 vdd.t289 vdd.t288 sky130_fd_pr__pfet_01v8 ad=3.51 pd=18.78 as=1.485 ps=9.33 w=9 l=0.5
X285 gnd.t223 commonsourceibias.t62 commonsourceibias.t63 gnd.t222 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X286 outputibias.t1 outputibias.t0 gnd.t149 gnd.t148 sky130_fd_pr__nfet_01v8 ad=2.34 pd=12.78 as=2.34 ps=12.78 w=6 l=2
X287 gnd.t221 commonsourceibias.t114 CSoutput.t156 gnd.t201 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X288 CSoutput.t176 a_n7636_8799.t115 vdd.t71 vdd.t70 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X289 CSoutput.t155 commonsourceibias.t115 gnd.t220 gnd.t219 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X290 vdd.t285 a_n1996_n452.t64 a_n1808_13878.t14 vdd.t284 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=3.51 ps=18.78 w=9 l=0.5
X291 CSoutput.t61 a_n7636_8799.t116 vdd.t69 vdd.t68 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X292 output.t7 CSoutput.t199 vdd.t186 gnd.t155 sky130_fd_pr__nfet_01v8 ad=0.825 pd=5.33 as=0.825 ps=5.33 w=5 l=1
X293 CSoutput.t2 a_n7636_8799.t117 vdd.t67 vdd.t37 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X294 gnd.t27 gnd.t24 gnd.t26 gnd.t25 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=0 ps=0 w=7 l=0.7
X295 gnd.t52 gnd.t49 gnd.t51 gnd.t50 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=0 ps=0 w=7 l=1
X296 vdd.t188 CSoutput.t200 output.t6 gnd.t154 sky130_fd_pr__nfet_01v8 ad=0.825 pd=5.33 as=0.825 ps=5.33 w=5 l=1
X297 gnd.t218 commonsourceibias.t116 CSoutput.t154 gnd.t194 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X298 CSoutput.t153 commonsourceibias.t117 gnd.t217 gnd.t198 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X299 CSoutput.t141 commonsourceibias.t118 gnd.t216 gnd.t215 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X300 vdd.t66 a_n7636_8799.t118 CSoutput.t167 vdd.t65 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X301 gnd.t214 commonsourceibias.t54 commonsourceibias.t55 gnd.t213 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X302 vdd.t64 a_n7636_8799.t119 CSoutput.t83 vdd.t29 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X303 vdd.t220 vdd.t217 vdd.t219 vdd.t218 sky130_fd_pr__pfet_01v8 ad=3.12 pd=16.78 as=0 ps=0 w=8 l=0.5
X304 minus.t0 gnd.t46 gnd.t48 gnd.t47 sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.5
X305 a_n2903_n3924.t43 minus.t20 a_n1996_n452.t41 gnd.t8 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.7
X306 a_n1986_8322.t3 a_n1996_n452.t65 a_n7636_8799.t0 vdd.t2 sky130_fd_pr__pfet_01v8 ad=3.51 pd=18.78 as=1.485 ps=9.33 w=9 l=0.5
X307 CSoutput.t5 a_n7636_8799.t120 vdd.t63 vdd.t62 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X308 vdd.t216 vdd.t214 vdd.t215 vdd.t211 sky130_fd_pr__pfet_01v8 ad=3.12 pd=16.78 as=0 ps=0 w=8 l=0.5
X309 a_n7636_8799.t31 a_n1996_n452.t66 a_n1986_8322.t2 vdd.t205 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X310 vdd.t61 a_n7636_8799.t121 CSoutput.t89 vdd.t60 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X311 a_n1808_13878.t13 a_n1996_n452.t67 vdd.t293 vdd.t292 sky130_fd_pr__pfet_01v8 ad=3.51 pd=18.78 as=1.485 ps=9.33 w=9 l=0.5
X312 gnd.t45 gnd.t42 gnd.t44 gnd.t43 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=0 ps=0 w=7 l=0.7
X313 vdd.t59 a_n7636_8799.t122 CSoutput.t28 vdd.t35 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X314 a_n1996_n452.t42 minus.t21 a_n2903_n3924.t44 gnd.t129 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.7
X315 CSoutput.t77 a_n7636_8799.t123 vdd.t58 vdd.t57 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X316 CSoutput.t140 commonsourceibias.t119 gnd.t212 gnd.t211 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X317 a_n7636_8799.t8 plus.t19 a_n2903_n3924.t21 gnd.t135 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.7
X318 a_n2903_n3924.t9 minus.t22 a_n1996_n452.t6 gnd.t125 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.7
X319 vdd.t56 a_n7636_8799.t124 CSoutput.t69 vdd.t55 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X320 CSoutput.t70 a_n7636_8799.t125 vdd.t54 vdd.t53 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X321 CSoutput.t96 a_n7636_8799.t126 vdd.t52 vdd.t33 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X322 CSoutput.t8 a_n7636_8799.t127 vdd.t51 vdd.t33 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X323 output.t5 CSoutput.t201 vdd.t190 gnd.t153 sky130_fd_pr__nfet_01v8 ad=0.825 pd=5.33 as=0.825 ps=5.33 w=5 l=1
X324 a_n1808_13878.t3 a_n1996_n452.t21 a_n1996_n452.t22 vdd.t3 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X325 CSoutput.t38 a_n7636_8799.t128 vdd.t50 vdd.t31 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X326 commonsourceibias.t53 commonsourceibias.t52 gnd.t210 gnd.t209 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X327 gnd.t208 commonsourceibias.t120 CSoutput.t139 gnd.t190 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X328 a_n2903_n3924.t20 plus.t20 a_n7636_8799.t7 gnd.t132 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.7
X329 vdd.t49 a_n7636_8799.t129 CSoutput.t171 vdd.t27 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X330 gnd.t41 gnd.t38 gnd.t40 gnd.t39 sky130_fd_pr__nfet_01v8 ad=1.95 pd=10.78 as=0 ps=0 w=5 l=1
X331 gnd.t207 commonsourceibias.t121 CSoutput.t138 gnd.t206 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X332 CSoutput.t11 a_n7636_8799.t130 vdd.t48 vdd.t23 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X333 output.t4 CSoutput.t202 vdd.t194 gnd.t152 sky130_fd_pr__nfet_01v8 ad=0.825 pd=5.33 as=0.825 ps=5.33 w=5 l=1
X334 gnd.t37 gnd.t35 gnd.t36 gnd.t18 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=0 ps=0 w=7 l=1
X335 a_n2903_n3924.t46 diffpairibias.t22 gnd.t313 gnd.t312 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=2.73 ps=14.78 w=7 l=1
X336 vdd.t47 a_n7636_8799.t131 CSoutput.t162 vdd.t21 sky130_fd_pr__pfet_01v8 ad=3.12 pd=16.78 as=1.32 ps=8.33 w=8 l=0.5
X337 vdd.t46 a_n7636_8799.t132 CSoutput.t91 vdd.t19 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X338 gnd.t34 gnd.t31 gnd.t33 gnd.t32 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=0 ps=0 w=7 l=1
X339 gnd.t185 commonsourceibias.t122 CSoutput.t143 gnd.t184 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X340 CSoutput.t177 a_n7636_8799.t133 vdd.t45 vdd.t15 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X341 a_n1996_n452.t28 a_n1996_n452.t27 a_n1808_13878.t2 vdd.t2 sky130_fd_pr__pfet_01v8 ad=3.51 pd=18.78 as=1.485 ps=9.33 w=9 l=0.5
X342 commonsourceibias.t51 commonsourceibias.t50 gnd.t205 gnd.t198 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X343 a_n7636_8799.t27 a_n1996_n452.t68 a_n1986_8322.t1 vdd.t176 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=3.51 ps=18.78 w=9 l=0.5
X344 vdd.t44 a_n7636_8799.t134 CSoutput.t95 vdd.t27 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X345 CSoutput.t49 a_n7636_8799.t135 vdd.t43 vdd.t42 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X346 a_n7636_8799.t6 plus.t21 a_n2903_n3924.t17 gnd.t14 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.7
X347 vdd.t41 a_n7636_8799.t136 CSoutput.t57 vdd.t11 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X348 gnd.t30 gnd.t28 plus.t1 gnd.t29 sky130_fd_pr__nfet_01v8 ad=0.39 pd=2.78 as=0.165 ps=1.33 w=1 l=0.5
X349 diffpairibias.t3 diffpairibias.t2 gnd.t319 gnd.t318 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=2.73 ps=14.78 w=7 l=1
X350 vdd.t40 a_n7636_8799.t137 CSoutput.t59 vdd.t39 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X351 vdd.t213 vdd.t210 vdd.t212 vdd.t211 sky130_fd_pr__pfet_01v8 ad=3.12 pd=16.78 as=0 ps=0 w=8 l=0.5
X352 CSoutput.t203 a_n1986_8322.t20 sky130_fd_pr__cap_mim_m3_1 l=12 w=12
X353 CSoutput.t172 a_n7636_8799.t138 vdd.t38 vdd.t37 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X354 a_n2903_n3924.t15 plus.t22 a_n7636_8799.t5 gnd.t5 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.7
X355 gnd.t23 gnd.t21 plus.t0 gnd.t22 sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.39 ps=2.78 w=1 l=0.5
X356 commonsourceibias.t49 commonsourceibias.t48 gnd.t204 gnd.t203 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X357 vdd.t36 a_n7636_8799.t139 CSoutput.t46 vdd.t35 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X358 gnd.t202 commonsourceibias.t123 CSoutput.t137 gnd.t201 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X359 gnd.t20 gnd.t17 gnd.t19 gnd.t18 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=0 ps=0 w=7 l=1
X360 diffpairibias.t1 diffpairibias.t0 gnd.t179 gnd.t178 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=2.73 ps=14.78 w=7 l=1
X361 a_n2903_n3924.t19 plus.t23 a_n7636_8799.t4 gnd.t166 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.7
X362 vdd.t187 CSoutput.t204 output.t3 gnd.t151 sky130_fd_pr__nfet_01v8 ad=0.825 pd=5.33 as=0.825 ps=5.33 w=5 l=1
X363 CSoutput.t142 commonsourceibias.t124 gnd.t183 gnd.t182 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X364 vdd.t201 a_n1996_n452.t69 a_n1808_13878.t12 vdd.t200 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=3.51 ps=18.78 w=9 l=0.5
X365 a_n7636_8799.t3 plus.t24 a_n2903_n3924.t29 gnd.t2 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=2.73 ps=14.78 w=7 l=0.7
X366 CSoutput.t21 a_n7636_8799.t140 vdd.t34 vdd.t33 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X367 gnd.t200 commonsourceibias.t125 CSoutput.t114 gnd.t194 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X368 CSoutput.t113 commonsourceibias.t126 gnd.t199 gnd.t198 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X369 a_n2903_n3924.t41 minus.t23 a_n1996_n452.t39 gnd.t169 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.7
X370 CSoutput.t178 a_n7636_8799.t141 vdd.t32 vdd.t31 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X371 vdd.t30 a_n7636_8799.t142 CSoutput.t174 vdd.t29 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X372 commonsourceibias.t25 commonsourceibias.t24 gnd.t197 gnd.t196 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X373 vdd.t28 a_n7636_8799.t143 CSoutput.t92 vdd.t27 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X374 CSoutput.t173 a_n7636_8799.t144 vdd.t26 vdd.t25 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X375 gnd.t195 commonsourceibias.t22 commonsourceibias.t23 gnd.t194 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X376 vdd.t189 CSoutput.t205 output.t2 gnd.t150 sky130_fd_pr__nfet_01v8 ad=0.825 pd=5.33 as=0.825 ps=5.33 w=5 l=1
X377 a_n1996_n452.t38 minus.t24 a_n2903_n3924.t40 gnd.t131 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=2.73 ps=14.78 w=7 l=0.7
X378 CSoutput.t112 commonsourceibias.t127 gnd.t193 gnd.t192 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X379 CSoutput.t54 a_n7636_8799.t145 vdd.t24 vdd.t23 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X380 a_n1986_8322.t0 a_n1996_n452.t70 a_n7636_8799.t23 vdd.t177 sky130_fd_pr__pfet_01v8 ad=3.51 pd=18.78 as=1.485 ps=9.33 w=9 l=0.5
X381 gnd.t191 commonsourceibias.t20 commonsourceibias.t21 gnd.t190 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X382 vdd.t22 a_n7636_8799.t146 CSoutput.t15 vdd.t21 sky130_fd_pr__pfet_01v8 ad=3.12 pd=16.78 as=1.32 ps=8.33 w=8 l=0.5
X383 vdd.t20 a_n7636_8799.t147 CSoutput.t71 vdd.t19 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X384 CSoutput.t81 a_n7636_8799.t148 vdd.t18 vdd.t17 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=3.12 ps=16.78 w=8 l=0.5
X385 CSoutput.t31 a_n7636_8799.t149 vdd.t16 vdd.t15 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X386 vdd.t14 a_n7636_8799.t150 CSoutput.t180 vdd.t13 sky130_fd_pr__pfet_01v8 ad=3.12 pd=16.78 as=1.32 ps=8.33 w=8 l=0.5
X387 commonsourceibias.t19 commonsourceibias.t18 gnd.t189 gnd.t188 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X388 a_n1986_8322.t12 a_n1996_n452.t71 vdd.t180 vdd.t179 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X389 a_n1808_13878.t1 a_n1996_n452.t23 a_n1996_n452.t24 vdd.t178 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=3.51 ps=18.78 w=9 l=0.5
X390 vdd.t12 a_n7636_8799.t151 CSoutput.t0 vdd.t11 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X391 commonsourceibias.t17 commonsourceibias.t16 gnd.t187 gnd.t186 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=2.73 ps=14.78 w=7 l=1
X392 a_n2903_n3924.t47 diffpairibias.t23 gnd.t317 gnd.t316 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=2.73 ps=14.78 w=7 l=1
X393 gnd.t181 commonsourceibias.t56 commonsourceibias.t57 gnd.t180 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X394 a_n1996_n452.t10 a_n1996_n452.t9 a_n1808_13878.t0 vdd.t204 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X395 vdd.t209 vdd.t206 vdd.t208 vdd.t207 sky130_fd_pr__pfet_01v8 ad=3.51 pd=18.78 as=0 ps=0 w=9 l=0.5
R0 commonsourceibias.n35 commonsourceibias.t38 223.028
R1 commonsourceibias.n128 commonsourceibias.t89 223.028
R2 commonsourceibias.n217 commonsourceibias.t77 223.028
R3 commonsourceibias.n364 commonsourceibias.t14 223.028
R4 commonsourceibias.n305 commonsourceibias.t108 223.028
R5 commonsourceibias.n499 commonsourceibias.t95 223.028
R6 commonsourceibias.n99 commonsourceibias.t34 207.983
R7 commonsourceibias.n192 commonsourceibias.t94 207.983
R8 commonsourceibias.n281 commonsourceibias.t81 207.983
R9 commonsourceibias.n430 commonsourceibias.t16 207.983
R10 commonsourceibias.n476 commonsourceibias.t113 207.983
R11 commonsourceibias.n565 commonsourceibias.t100 207.983
R12 commonsourceibias.n97 commonsourceibias.t52 168.701
R13 commonsourceibias.n91 commonsourceibias.t26 168.701
R14 commonsourceibias.n17 commonsourceibias.t32 168.701
R15 commonsourceibias.n83 commonsourceibias.t46 168.701
R16 commonsourceibias.n77 commonsourceibias.t8 168.701
R17 commonsourceibias.n22 commonsourceibias.t4 168.701
R18 commonsourceibias.n69 commonsourceibias.t28 168.701
R19 commonsourceibias.n63 commonsourceibias.t36 168.701
R20 commonsourceibias.n25 commonsourceibias.t48 168.701
R21 commonsourceibias.n27 commonsourceibias.t0 168.701
R22 commonsourceibias.n29 commonsourceibias.t6 168.701
R23 commonsourceibias.n46 commonsourceibias.t42 168.701
R24 commonsourceibias.n40 commonsourceibias.t10 168.701
R25 commonsourceibias.n34 commonsourceibias.t54 168.701
R26 commonsourceibias.n190 commonsourceibias.t109 168.701
R27 commonsourceibias.n184 commonsourceibias.t72 168.701
R28 commonsourceibias.n5 commonsourceibias.t70 168.701
R29 commonsourceibias.n176 commonsourceibias.t102 168.701
R30 commonsourceibias.n170 commonsourceibias.t118 168.701
R31 commonsourceibias.n10 commonsourceibias.t66 168.701
R32 commonsourceibias.n162 commonsourceibias.t93 168.701
R33 commonsourceibias.n156 commonsourceibias.t88 168.701
R34 commonsourceibias.n118 commonsourceibias.t105 168.701
R35 commonsourceibias.n120 commonsourceibias.t86 168.701
R36 commonsourceibias.n122 commonsourceibias.t82 168.701
R37 commonsourceibias.n139 commonsourceibias.t97 168.701
R38 commonsourceibias.n133 commonsourceibias.t111 168.701
R39 commonsourceibias.n127 commonsourceibias.t75 168.701
R40 commonsourceibias.n216 commonsourceibias.t67 168.701
R41 commonsourceibias.n222 commonsourceibias.t98 168.701
R42 commonsourceibias.n228 commonsourceibias.t83 168.701
R43 commonsourceibias.n211 commonsourceibias.t71 168.701
R44 commonsourceibias.n209 commonsourceibias.t74 168.701
R45 commonsourceibias.n207 commonsourceibias.t90 168.701
R46 commonsourceibias.n245 commonsourceibias.t76 168.701
R47 commonsourceibias.n251 commonsourceibias.t80 168.701
R48 commonsourceibias.n204 commonsourceibias.t122 168.701
R49 commonsourceibias.n259 commonsourceibias.t104 168.701
R50 commonsourceibias.n265 commonsourceibias.t87 168.701
R51 commonsourceibias.n199 commonsourceibias.t127 168.701
R52 commonsourceibias.n273 commonsourceibias.t65 168.701
R53 commonsourceibias.n279 commonsourceibias.t96 168.701
R54 commonsourceibias.n363 commonsourceibias.t60 168.701
R55 commonsourceibias.n369 commonsourceibias.t22 168.701
R56 commonsourceibias.n375 commonsourceibias.t40 168.701
R57 commonsourceibias.n358 commonsourceibias.t62 168.701
R58 commonsourceibias.n356 commonsourceibias.t24 168.701
R59 commonsourceibias.n354 commonsourceibias.t44 168.701
R60 commonsourceibias.n392 commonsourceibias.t18 168.701
R61 commonsourceibias.n398 commonsourceibias.t2 168.701
R62 commonsourceibias.n400 commonsourceibias.t50 168.701
R63 commonsourceibias.n407 commonsourceibias.t20 168.701
R64 commonsourceibias.n413 commonsourceibias.t30 168.701
R65 commonsourceibias.n415 commonsourceibias.t56 168.701
R66 commonsourceibias.n422 commonsourceibias.t12 168.701
R67 commonsourceibias.n428 commonsourceibias.t58 168.701
R68 commonsourceibias.n474 commonsourceibias.t123 168.701
R69 commonsourceibias.n468 commonsourceibias.t68 168.701
R70 commonsourceibias.n461 commonsourceibias.t84 168.701
R71 commonsourceibias.n459 commonsourceibias.t119 168.701
R72 commonsourceibias.n453 commonsourceibias.t64 168.701
R73 commonsourceibias.n446 commonsourceibias.t126 168.701
R74 commonsourceibias.n444 commonsourceibias.t112 168.701
R75 commonsourceibias.n304 commonsourceibias.t91 168.701
R76 commonsourceibias.n310 commonsourceibias.t125 168.701
R77 commonsourceibias.n316 commonsourceibias.t115 168.701
R78 commonsourceibias.n299 commonsourceibias.t101 168.701
R79 commonsourceibias.n297 commonsourceibias.t78 168.701
R80 commonsourceibias.n295 commonsourceibias.t121 168.701
R81 commonsourceibias.n333 commonsourceibias.t107 168.701
R82 commonsourceibias.n498 commonsourceibias.t79 168.701
R83 commonsourceibias.n504 commonsourceibias.t116 168.701
R84 commonsourceibias.n510 commonsourceibias.t103 168.701
R85 commonsourceibias.n493 commonsourceibias.t85 168.701
R86 commonsourceibias.n491 commonsourceibias.t69 168.701
R87 commonsourceibias.n489 commonsourceibias.t110 168.701
R88 commonsourceibias.n527 commonsourceibias.t92 168.701
R89 commonsourceibias.n533 commonsourceibias.t99 168.701
R90 commonsourceibias.n535 commonsourceibias.t117 168.701
R91 commonsourceibias.n542 commonsourceibias.t120 168.701
R92 commonsourceibias.n548 commonsourceibias.t106 168.701
R93 commonsourceibias.n550 commonsourceibias.t73 168.701
R94 commonsourceibias.n557 commonsourceibias.t124 168.701
R95 commonsourceibias.n563 commonsourceibias.t114 168.701
R96 commonsourceibias.n36 commonsourceibias.n33 161.3
R97 commonsourceibias.n38 commonsourceibias.n37 161.3
R98 commonsourceibias.n39 commonsourceibias.n32 161.3
R99 commonsourceibias.n42 commonsourceibias.n41 161.3
R100 commonsourceibias.n43 commonsourceibias.n31 161.3
R101 commonsourceibias.n45 commonsourceibias.n44 161.3
R102 commonsourceibias.n47 commonsourceibias.n30 161.3
R103 commonsourceibias.n49 commonsourceibias.n48 161.3
R104 commonsourceibias.n51 commonsourceibias.n50 161.3
R105 commonsourceibias.n52 commonsourceibias.n28 161.3
R106 commonsourceibias.n54 commonsourceibias.n53 161.3
R107 commonsourceibias.n56 commonsourceibias.n55 161.3
R108 commonsourceibias.n57 commonsourceibias.n26 161.3
R109 commonsourceibias.n59 commonsourceibias.n58 161.3
R110 commonsourceibias.n61 commonsourceibias.n60 161.3
R111 commonsourceibias.n62 commonsourceibias.n24 161.3
R112 commonsourceibias.n65 commonsourceibias.n64 161.3
R113 commonsourceibias.n66 commonsourceibias.n23 161.3
R114 commonsourceibias.n68 commonsourceibias.n67 161.3
R115 commonsourceibias.n70 commonsourceibias.n21 161.3
R116 commonsourceibias.n72 commonsourceibias.n71 161.3
R117 commonsourceibias.n73 commonsourceibias.n20 161.3
R118 commonsourceibias.n75 commonsourceibias.n74 161.3
R119 commonsourceibias.n76 commonsourceibias.n19 161.3
R120 commonsourceibias.n79 commonsourceibias.n78 161.3
R121 commonsourceibias.n80 commonsourceibias.n18 161.3
R122 commonsourceibias.n82 commonsourceibias.n81 161.3
R123 commonsourceibias.n84 commonsourceibias.n16 161.3
R124 commonsourceibias.n86 commonsourceibias.n85 161.3
R125 commonsourceibias.n87 commonsourceibias.n15 161.3
R126 commonsourceibias.n89 commonsourceibias.n88 161.3
R127 commonsourceibias.n90 commonsourceibias.n14 161.3
R128 commonsourceibias.n93 commonsourceibias.n92 161.3
R129 commonsourceibias.n94 commonsourceibias.n13 161.3
R130 commonsourceibias.n96 commonsourceibias.n95 161.3
R131 commonsourceibias.n98 commonsourceibias.n12 161.3
R132 commonsourceibias.n129 commonsourceibias.n126 161.3
R133 commonsourceibias.n131 commonsourceibias.n130 161.3
R134 commonsourceibias.n132 commonsourceibias.n125 161.3
R135 commonsourceibias.n135 commonsourceibias.n134 161.3
R136 commonsourceibias.n136 commonsourceibias.n124 161.3
R137 commonsourceibias.n138 commonsourceibias.n137 161.3
R138 commonsourceibias.n140 commonsourceibias.n123 161.3
R139 commonsourceibias.n142 commonsourceibias.n141 161.3
R140 commonsourceibias.n144 commonsourceibias.n143 161.3
R141 commonsourceibias.n145 commonsourceibias.n121 161.3
R142 commonsourceibias.n147 commonsourceibias.n146 161.3
R143 commonsourceibias.n149 commonsourceibias.n148 161.3
R144 commonsourceibias.n150 commonsourceibias.n119 161.3
R145 commonsourceibias.n152 commonsourceibias.n151 161.3
R146 commonsourceibias.n154 commonsourceibias.n153 161.3
R147 commonsourceibias.n155 commonsourceibias.n117 161.3
R148 commonsourceibias.n158 commonsourceibias.n157 161.3
R149 commonsourceibias.n159 commonsourceibias.n11 161.3
R150 commonsourceibias.n161 commonsourceibias.n160 161.3
R151 commonsourceibias.n163 commonsourceibias.n9 161.3
R152 commonsourceibias.n165 commonsourceibias.n164 161.3
R153 commonsourceibias.n166 commonsourceibias.n8 161.3
R154 commonsourceibias.n168 commonsourceibias.n167 161.3
R155 commonsourceibias.n169 commonsourceibias.n7 161.3
R156 commonsourceibias.n172 commonsourceibias.n171 161.3
R157 commonsourceibias.n173 commonsourceibias.n6 161.3
R158 commonsourceibias.n175 commonsourceibias.n174 161.3
R159 commonsourceibias.n177 commonsourceibias.n4 161.3
R160 commonsourceibias.n179 commonsourceibias.n178 161.3
R161 commonsourceibias.n180 commonsourceibias.n3 161.3
R162 commonsourceibias.n182 commonsourceibias.n181 161.3
R163 commonsourceibias.n183 commonsourceibias.n2 161.3
R164 commonsourceibias.n186 commonsourceibias.n185 161.3
R165 commonsourceibias.n187 commonsourceibias.n1 161.3
R166 commonsourceibias.n189 commonsourceibias.n188 161.3
R167 commonsourceibias.n191 commonsourceibias.n0 161.3
R168 commonsourceibias.n280 commonsourceibias.n194 161.3
R169 commonsourceibias.n278 commonsourceibias.n277 161.3
R170 commonsourceibias.n276 commonsourceibias.n195 161.3
R171 commonsourceibias.n275 commonsourceibias.n274 161.3
R172 commonsourceibias.n272 commonsourceibias.n196 161.3
R173 commonsourceibias.n271 commonsourceibias.n270 161.3
R174 commonsourceibias.n269 commonsourceibias.n197 161.3
R175 commonsourceibias.n268 commonsourceibias.n267 161.3
R176 commonsourceibias.n266 commonsourceibias.n198 161.3
R177 commonsourceibias.n264 commonsourceibias.n263 161.3
R178 commonsourceibias.n262 commonsourceibias.n200 161.3
R179 commonsourceibias.n261 commonsourceibias.n260 161.3
R180 commonsourceibias.n258 commonsourceibias.n201 161.3
R181 commonsourceibias.n257 commonsourceibias.n256 161.3
R182 commonsourceibias.n255 commonsourceibias.n202 161.3
R183 commonsourceibias.n254 commonsourceibias.n253 161.3
R184 commonsourceibias.n252 commonsourceibias.n203 161.3
R185 commonsourceibias.n250 commonsourceibias.n249 161.3
R186 commonsourceibias.n248 commonsourceibias.n205 161.3
R187 commonsourceibias.n247 commonsourceibias.n246 161.3
R188 commonsourceibias.n244 commonsourceibias.n206 161.3
R189 commonsourceibias.n243 commonsourceibias.n242 161.3
R190 commonsourceibias.n241 commonsourceibias.n240 161.3
R191 commonsourceibias.n239 commonsourceibias.n208 161.3
R192 commonsourceibias.n238 commonsourceibias.n237 161.3
R193 commonsourceibias.n236 commonsourceibias.n235 161.3
R194 commonsourceibias.n234 commonsourceibias.n210 161.3
R195 commonsourceibias.n233 commonsourceibias.n232 161.3
R196 commonsourceibias.n231 commonsourceibias.n230 161.3
R197 commonsourceibias.n229 commonsourceibias.n212 161.3
R198 commonsourceibias.n227 commonsourceibias.n226 161.3
R199 commonsourceibias.n225 commonsourceibias.n213 161.3
R200 commonsourceibias.n224 commonsourceibias.n223 161.3
R201 commonsourceibias.n221 commonsourceibias.n214 161.3
R202 commonsourceibias.n220 commonsourceibias.n219 161.3
R203 commonsourceibias.n218 commonsourceibias.n215 161.3
R204 commonsourceibias.n429 commonsourceibias.n343 161.3
R205 commonsourceibias.n427 commonsourceibias.n426 161.3
R206 commonsourceibias.n425 commonsourceibias.n344 161.3
R207 commonsourceibias.n424 commonsourceibias.n423 161.3
R208 commonsourceibias.n421 commonsourceibias.n345 161.3
R209 commonsourceibias.n420 commonsourceibias.n419 161.3
R210 commonsourceibias.n418 commonsourceibias.n346 161.3
R211 commonsourceibias.n417 commonsourceibias.n416 161.3
R212 commonsourceibias.n414 commonsourceibias.n347 161.3
R213 commonsourceibias.n412 commonsourceibias.n411 161.3
R214 commonsourceibias.n410 commonsourceibias.n348 161.3
R215 commonsourceibias.n409 commonsourceibias.n408 161.3
R216 commonsourceibias.n406 commonsourceibias.n349 161.3
R217 commonsourceibias.n405 commonsourceibias.n404 161.3
R218 commonsourceibias.n403 commonsourceibias.n350 161.3
R219 commonsourceibias.n402 commonsourceibias.n401 161.3
R220 commonsourceibias.n399 commonsourceibias.n351 161.3
R221 commonsourceibias.n397 commonsourceibias.n396 161.3
R222 commonsourceibias.n395 commonsourceibias.n352 161.3
R223 commonsourceibias.n394 commonsourceibias.n393 161.3
R224 commonsourceibias.n391 commonsourceibias.n353 161.3
R225 commonsourceibias.n390 commonsourceibias.n389 161.3
R226 commonsourceibias.n388 commonsourceibias.n387 161.3
R227 commonsourceibias.n386 commonsourceibias.n355 161.3
R228 commonsourceibias.n385 commonsourceibias.n384 161.3
R229 commonsourceibias.n383 commonsourceibias.n382 161.3
R230 commonsourceibias.n381 commonsourceibias.n357 161.3
R231 commonsourceibias.n380 commonsourceibias.n379 161.3
R232 commonsourceibias.n378 commonsourceibias.n377 161.3
R233 commonsourceibias.n376 commonsourceibias.n359 161.3
R234 commonsourceibias.n374 commonsourceibias.n373 161.3
R235 commonsourceibias.n372 commonsourceibias.n360 161.3
R236 commonsourceibias.n371 commonsourceibias.n370 161.3
R237 commonsourceibias.n368 commonsourceibias.n361 161.3
R238 commonsourceibias.n367 commonsourceibias.n366 161.3
R239 commonsourceibias.n365 commonsourceibias.n362 161.3
R240 commonsourceibias.n335 commonsourceibias.n334 161.3
R241 commonsourceibias.n332 commonsourceibias.n294 161.3
R242 commonsourceibias.n331 commonsourceibias.n330 161.3
R243 commonsourceibias.n329 commonsourceibias.n328 161.3
R244 commonsourceibias.n327 commonsourceibias.n296 161.3
R245 commonsourceibias.n326 commonsourceibias.n325 161.3
R246 commonsourceibias.n324 commonsourceibias.n323 161.3
R247 commonsourceibias.n322 commonsourceibias.n298 161.3
R248 commonsourceibias.n321 commonsourceibias.n320 161.3
R249 commonsourceibias.n319 commonsourceibias.n318 161.3
R250 commonsourceibias.n317 commonsourceibias.n300 161.3
R251 commonsourceibias.n315 commonsourceibias.n314 161.3
R252 commonsourceibias.n313 commonsourceibias.n301 161.3
R253 commonsourceibias.n312 commonsourceibias.n311 161.3
R254 commonsourceibias.n309 commonsourceibias.n302 161.3
R255 commonsourceibias.n308 commonsourceibias.n307 161.3
R256 commonsourceibias.n306 commonsourceibias.n303 161.3
R257 commonsourceibias.n441 commonsourceibias.n293 161.3
R258 commonsourceibias.n475 commonsourceibias.n284 161.3
R259 commonsourceibias.n473 commonsourceibias.n472 161.3
R260 commonsourceibias.n471 commonsourceibias.n285 161.3
R261 commonsourceibias.n470 commonsourceibias.n469 161.3
R262 commonsourceibias.n467 commonsourceibias.n286 161.3
R263 commonsourceibias.n466 commonsourceibias.n465 161.3
R264 commonsourceibias.n464 commonsourceibias.n287 161.3
R265 commonsourceibias.n463 commonsourceibias.n462 161.3
R266 commonsourceibias.n460 commonsourceibias.n288 161.3
R267 commonsourceibias.n458 commonsourceibias.n457 161.3
R268 commonsourceibias.n456 commonsourceibias.n289 161.3
R269 commonsourceibias.n455 commonsourceibias.n454 161.3
R270 commonsourceibias.n452 commonsourceibias.n290 161.3
R271 commonsourceibias.n451 commonsourceibias.n450 161.3
R272 commonsourceibias.n449 commonsourceibias.n291 161.3
R273 commonsourceibias.n448 commonsourceibias.n447 161.3
R274 commonsourceibias.n445 commonsourceibias.n292 161.3
R275 commonsourceibias.n443 commonsourceibias.n442 161.3
R276 commonsourceibias.n564 commonsourceibias.n478 161.3
R277 commonsourceibias.n562 commonsourceibias.n561 161.3
R278 commonsourceibias.n560 commonsourceibias.n479 161.3
R279 commonsourceibias.n559 commonsourceibias.n558 161.3
R280 commonsourceibias.n556 commonsourceibias.n480 161.3
R281 commonsourceibias.n555 commonsourceibias.n554 161.3
R282 commonsourceibias.n553 commonsourceibias.n481 161.3
R283 commonsourceibias.n552 commonsourceibias.n551 161.3
R284 commonsourceibias.n549 commonsourceibias.n482 161.3
R285 commonsourceibias.n547 commonsourceibias.n546 161.3
R286 commonsourceibias.n545 commonsourceibias.n483 161.3
R287 commonsourceibias.n544 commonsourceibias.n543 161.3
R288 commonsourceibias.n541 commonsourceibias.n484 161.3
R289 commonsourceibias.n540 commonsourceibias.n539 161.3
R290 commonsourceibias.n538 commonsourceibias.n485 161.3
R291 commonsourceibias.n537 commonsourceibias.n536 161.3
R292 commonsourceibias.n534 commonsourceibias.n486 161.3
R293 commonsourceibias.n532 commonsourceibias.n531 161.3
R294 commonsourceibias.n530 commonsourceibias.n487 161.3
R295 commonsourceibias.n529 commonsourceibias.n528 161.3
R296 commonsourceibias.n526 commonsourceibias.n488 161.3
R297 commonsourceibias.n525 commonsourceibias.n524 161.3
R298 commonsourceibias.n523 commonsourceibias.n522 161.3
R299 commonsourceibias.n521 commonsourceibias.n490 161.3
R300 commonsourceibias.n520 commonsourceibias.n519 161.3
R301 commonsourceibias.n518 commonsourceibias.n517 161.3
R302 commonsourceibias.n516 commonsourceibias.n492 161.3
R303 commonsourceibias.n515 commonsourceibias.n514 161.3
R304 commonsourceibias.n513 commonsourceibias.n512 161.3
R305 commonsourceibias.n511 commonsourceibias.n494 161.3
R306 commonsourceibias.n509 commonsourceibias.n508 161.3
R307 commonsourceibias.n507 commonsourceibias.n495 161.3
R308 commonsourceibias.n506 commonsourceibias.n505 161.3
R309 commonsourceibias.n503 commonsourceibias.n496 161.3
R310 commonsourceibias.n502 commonsourceibias.n501 161.3
R311 commonsourceibias.n500 commonsourceibias.n497 161.3
R312 commonsourceibias.n111 commonsourceibias.n109 81.5057
R313 commonsourceibias.n338 commonsourceibias.n336 81.5057
R314 commonsourceibias.n111 commonsourceibias.n110 80.9324
R315 commonsourceibias.n113 commonsourceibias.n112 80.9324
R316 commonsourceibias.n115 commonsourceibias.n114 80.9324
R317 commonsourceibias.n108 commonsourceibias.n107 80.9324
R318 commonsourceibias.n106 commonsourceibias.n105 80.9324
R319 commonsourceibias.n104 commonsourceibias.n103 80.9324
R320 commonsourceibias.n102 commonsourceibias.n101 80.9324
R321 commonsourceibias.n433 commonsourceibias.n432 80.9324
R322 commonsourceibias.n435 commonsourceibias.n434 80.9324
R323 commonsourceibias.n437 commonsourceibias.n436 80.9324
R324 commonsourceibias.n439 commonsourceibias.n438 80.9324
R325 commonsourceibias.n342 commonsourceibias.n341 80.9324
R326 commonsourceibias.n340 commonsourceibias.n339 80.9324
R327 commonsourceibias.n338 commonsourceibias.n337 80.9324
R328 commonsourceibias.n100 commonsourceibias.n99 80.6037
R329 commonsourceibias.n193 commonsourceibias.n192 80.6037
R330 commonsourceibias.n282 commonsourceibias.n281 80.6037
R331 commonsourceibias.n431 commonsourceibias.n430 80.6037
R332 commonsourceibias.n477 commonsourceibias.n476 80.6037
R333 commonsourceibias.n566 commonsourceibias.n565 80.6037
R334 commonsourceibias.n85 commonsourceibias.n84 56.5617
R335 commonsourceibias.n71 commonsourceibias.n70 56.5617
R336 commonsourceibias.n62 commonsourceibias.n61 56.5617
R337 commonsourceibias.n48 commonsourceibias.n47 56.5617
R338 commonsourceibias.n178 commonsourceibias.n177 56.5617
R339 commonsourceibias.n164 commonsourceibias.n163 56.5617
R340 commonsourceibias.n155 commonsourceibias.n154 56.5617
R341 commonsourceibias.n141 commonsourceibias.n140 56.5617
R342 commonsourceibias.n230 commonsourceibias.n229 56.5617
R343 commonsourceibias.n244 commonsourceibias.n243 56.5617
R344 commonsourceibias.n253 commonsourceibias.n252 56.5617
R345 commonsourceibias.n267 commonsourceibias.n266 56.5617
R346 commonsourceibias.n377 commonsourceibias.n376 56.5617
R347 commonsourceibias.n391 commonsourceibias.n390 56.5617
R348 commonsourceibias.n401 commonsourceibias.n399 56.5617
R349 commonsourceibias.n416 commonsourceibias.n414 56.5617
R350 commonsourceibias.n462 commonsourceibias.n460 56.5617
R351 commonsourceibias.n447 commonsourceibias.n445 56.5617
R352 commonsourceibias.n318 commonsourceibias.n317 56.5617
R353 commonsourceibias.n332 commonsourceibias.n331 56.5617
R354 commonsourceibias.n512 commonsourceibias.n511 56.5617
R355 commonsourceibias.n526 commonsourceibias.n525 56.5617
R356 commonsourceibias.n536 commonsourceibias.n534 56.5617
R357 commonsourceibias.n551 commonsourceibias.n549 56.5617
R358 commonsourceibias.n76 commonsourceibias.n75 56.0773
R359 commonsourceibias.n57 commonsourceibias.n56 56.0773
R360 commonsourceibias.n169 commonsourceibias.n168 56.0773
R361 commonsourceibias.n150 commonsourceibias.n149 56.0773
R362 commonsourceibias.n239 commonsourceibias.n238 56.0773
R363 commonsourceibias.n258 commonsourceibias.n257 56.0773
R364 commonsourceibias.n386 commonsourceibias.n385 56.0773
R365 commonsourceibias.n406 commonsourceibias.n405 56.0773
R366 commonsourceibias.n452 commonsourceibias.n451 56.0773
R367 commonsourceibias.n327 commonsourceibias.n326 56.0773
R368 commonsourceibias.n521 commonsourceibias.n520 56.0773
R369 commonsourceibias.n541 commonsourceibias.n540 56.0773
R370 commonsourceibias.n99 commonsourceibias.n98 55.3321
R371 commonsourceibias.n192 commonsourceibias.n191 55.3321
R372 commonsourceibias.n281 commonsourceibias.n280 55.3321
R373 commonsourceibias.n430 commonsourceibias.n429 55.3321
R374 commonsourceibias.n476 commonsourceibias.n475 55.3321
R375 commonsourceibias.n565 commonsourceibias.n564 55.3321
R376 commonsourceibias.n90 commonsourceibias.n89 55.1086
R377 commonsourceibias.n41 commonsourceibias.n31 55.1086
R378 commonsourceibias.n183 commonsourceibias.n182 55.1086
R379 commonsourceibias.n134 commonsourceibias.n124 55.1086
R380 commonsourceibias.n223 commonsourceibias.n213 55.1086
R381 commonsourceibias.n272 commonsourceibias.n271 55.1086
R382 commonsourceibias.n370 commonsourceibias.n360 55.1086
R383 commonsourceibias.n421 commonsourceibias.n420 55.1086
R384 commonsourceibias.n467 commonsourceibias.n466 55.1086
R385 commonsourceibias.n311 commonsourceibias.n301 55.1086
R386 commonsourceibias.n505 commonsourceibias.n495 55.1086
R387 commonsourceibias.n556 commonsourceibias.n555 55.1086
R388 commonsourceibias.n35 commonsourceibias.n34 47.4592
R389 commonsourceibias.n128 commonsourceibias.n127 47.4592
R390 commonsourceibias.n217 commonsourceibias.n216 47.4592
R391 commonsourceibias.n364 commonsourceibias.n363 47.4592
R392 commonsourceibias.n305 commonsourceibias.n304 47.4592
R393 commonsourceibias.n499 commonsourceibias.n498 47.4592
R394 commonsourceibias.n218 commonsourceibias.n217 44.0436
R395 commonsourceibias.n365 commonsourceibias.n364 44.0436
R396 commonsourceibias.n306 commonsourceibias.n305 44.0436
R397 commonsourceibias.n500 commonsourceibias.n499 44.0436
R398 commonsourceibias.n36 commonsourceibias.n35 44.0436
R399 commonsourceibias.n129 commonsourceibias.n128 44.0436
R400 commonsourceibias.n92 commonsourceibias.n13 42.5146
R401 commonsourceibias.n39 commonsourceibias.n38 42.5146
R402 commonsourceibias.n185 commonsourceibias.n1 42.5146
R403 commonsourceibias.n132 commonsourceibias.n131 42.5146
R404 commonsourceibias.n221 commonsourceibias.n220 42.5146
R405 commonsourceibias.n274 commonsourceibias.n195 42.5146
R406 commonsourceibias.n368 commonsourceibias.n367 42.5146
R407 commonsourceibias.n423 commonsourceibias.n344 42.5146
R408 commonsourceibias.n469 commonsourceibias.n285 42.5146
R409 commonsourceibias.n309 commonsourceibias.n308 42.5146
R410 commonsourceibias.n503 commonsourceibias.n502 42.5146
R411 commonsourceibias.n558 commonsourceibias.n479 42.5146
R412 commonsourceibias.n78 commonsourceibias.n18 41.5458
R413 commonsourceibias.n53 commonsourceibias.n52 41.5458
R414 commonsourceibias.n171 commonsourceibias.n6 41.5458
R415 commonsourceibias.n146 commonsourceibias.n145 41.5458
R416 commonsourceibias.n235 commonsourceibias.n234 41.5458
R417 commonsourceibias.n260 commonsourceibias.n200 41.5458
R418 commonsourceibias.n382 commonsourceibias.n381 41.5458
R419 commonsourceibias.n408 commonsourceibias.n348 41.5458
R420 commonsourceibias.n454 commonsourceibias.n289 41.5458
R421 commonsourceibias.n323 commonsourceibias.n322 41.5458
R422 commonsourceibias.n517 commonsourceibias.n516 41.5458
R423 commonsourceibias.n543 commonsourceibias.n483 41.5458
R424 commonsourceibias.n68 commonsourceibias.n23 40.577
R425 commonsourceibias.n64 commonsourceibias.n23 40.577
R426 commonsourceibias.n161 commonsourceibias.n11 40.577
R427 commonsourceibias.n157 commonsourceibias.n11 40.577
R428 commonsourceibias.n246 commonsourceibias.n205 40.577
R429 commonsourceibias.n250 commonsourceibias.n205 40.577
R430 commonsourceibias.n393 commonsourceibias.n352 40.577
R431 commonsourceibias.n397 commonsourceibias.n352 40.577
R432 commonsourceibias.n443 commonsourceibias.n293 40.577
R433 commonsourceibias.n334 commonsourceibias.n293 40.577
R434 commonsourceibias.n528 commonsourceibias.n487 40.577
R435 commonsourceibias.n532 commonsourceibias.n487 40.577
R436 commonsourceibias.n82 commonsourceibias.n18 39.6083
R437 commonsourceibias.n52 commonsourceibias.n51 39.6083
R438 commonsourceibias.n175 commonsourceibias.n6 39.6083
R439 commonsourceibias.n145 commonsourceibias.n144 39.6083
R440 commonsourceibias.n234 commonsourceibias.n233 39.6083
R441 commonsourceibias.n264 commonsourceibias.n200 39.6083
R442 commonsourceibias.n381 commonsourceibias.n380 39.6083
R443 commonsourceibias.n412 commonsourceibias.n348 39.6083
R444 commonsourceibias.n458 commonsourceibias.n289 39.6083
R445 commonsourceibias.n322 commonsourceibias.n321 39.6083
R446 commonsourceibias.n516 commonsourceibias.n515 39.6083
R447 commonsourceibias.n547 commonsourceibias.n483 39.6083
R448 commonsourceibias.n96 commonsourceibias.n13 38.6395
R449 commonsourceibias.n38 commonsourceibias.n33 38.6395
R450 commonsourceibias.n189 commonsourceibias.n1 38.6395
R451 commonsourceibias.n131 commonsourceibias.n126 38.6395
R452 commonsourceibias.n220 commonsourceibias.n215 38.6395
R453 commonsourceibias.n278 commonsourceibias.n195 38.6395
R454 commonsourceibias.n367 commonsourceibias.n362 38.6395
R455 commonsourceibias.n427 commonsourceibias.n344 38.6395
R456 commonsourceibias.n473 commonsourceibias.n285 38.6395
R457 commonsourceibias.n308 commonsourceibias.n303 38.6395
R458 commonsourceibias.n502 commonsourceibias.n497 38.6395
R459 commonsourceibias.n562 commonsourceibias.n479 38.6395
R460 commonsourceibias.n89 commonsourceibias.n15 26.0455
R461 commonsourceibias.n45 commonsourceibias.n31 26.0455
R462 commonsourceibias.n182 commonsourceibias.n3 26.0455
R463 commonsourceibias.n138 commonsourceibias.n124 26.0455
R464 commonsourceibias.n227 commonsourceibias.n213 26.0455
R465 commonsourceibias.n271 commonsourceibias.n197 26.0455
R466 commonsourceibias.n374 commonsourceibias.n360 26.0455
R467 commonsourceibias.n420 commonsourceibias.n346 26.0455
R468 commonsourceibias.n466 commonsourceibias.n287 26.0455
R469 commonsourceibias.n315 commonsourceibias.n301 26.0455
R470 commonsourceibias.n509 commonsourceibias.n495 26.0455
R471 commonsourceibias.n555 commonsourceibias.n481 26.0455
R472 commonsourceibias.n75 commonsourceibias.n20 25.0767
R473 commonsourceibias.n58 commonsourceibias.n57 25.0767
R474 commonsourceibias.n168 commonsourceibias.n8 25.0767
R475 commonsourceibias.n151 commonsourceibias.n150 25.0767
R476 commonsourceibias.n240 commonsourceibias.n239 25.0767
R477 commonsourceibias.n257 commonsourceibias.n202 25.0767
R478 commonsourceibias.n387 commonsourceibias.n386 25.0767
R479 commonsourceibias.n405 commonsourceibias.n350 25.0767
R480 commonsourceibias.n451 commonsourceibias.n291 25.0767
R481 commonsourceibias.n328 commonsourceibias.n327 25.0767
R482 commonsourceibias.n522 commonsourceibias.n521 25.0767
R483 commonsourceibias.n540 commonsourceibias.n485 25.0767
R484 commonsourceibias.n71 commonsourceibias.n22 24.3464
R485 commonsourceibias.n61 commonsourceibias.n25 24.3464
R486 commonsourceibias.n164 commonsourceibias.n10 24.3464
R487 commonsourceibias.n154 commonsourceibias.n118 24.3464
R488 commonsourceibias.n243 commonsourceibias.n207 24.3464
R489 commonsourceibias.n253 commonsourceibias.n204 24.3464
R490 commonsourceibias.n390 commonsourceibias.n354 24.3464
R491 commonsourceibias.n401 commonsourceibias.n400 24.3464
R492 commonsourceibias.n447 commonsourceibias.n446 24.3464
R493 commonsourceibias.n331 commonsourceibias.n295 24.3464
R494 commonsourceibias.n525 commonsourceibias.n489 24.3464
R495 commonsourceibias.n536 commonsourceibias.n535 24.3464
R496 commonsourceibias.n85 commonsourceibias.n17 23.8546
R497 commonsourceibias.n47 commonsourceibias.n46 23.8546
R498 commonsourceibias.n178 commonsourceibias.n5 23.8546
R499 commonsourceibias.n140 commonsourceibias.n139 23.8546
R500 commonsourceibias.n229 commonsourceibias.n228 23.8546
R501 commonsourceibias.n267 commonsourceibias.n199 23.8546
R502 commonsourceibias.n376 commonsourceibias.n375 23.8546
R503 commonsourceibias.n416 commonsourceibias.n415 23.8546
R504 commonsourceibias.n462 commonsourceibias.n461 23.8546
R505 commonsourceibias.n317 commonsourceibias.n316 23.8546
R506 commonsourceibias.n511 commonsourceibias.n510 23.8546
R507 commonsourceibias.n551 commonsourceibias.n550 23.8546
R508 commonsourceibias.n98 commonsourceibias.n97 17.4607
R509 commonsourceibias.n191 commonsourceibias.n190 17.4607
R510 commonsourceibias.n280 commonsourceibias.n279 17.4607
R511 commonsourceibias.n429 commonsourceibias.n428 17.4607
R512 commonsourceibias.n475 commonsourceibias.n474 17.4607
R513 commonsourceibias.n564 commonsourceibias.n563 17.4607
R514 commonsourceibias.n84 commonsourceibias.n83 16.9689
R515 commonsourceibias.n48 commonsourceibias.n29 16.9689
R516 commonsourceibias.n177 commonsourceibias.n176 16.9689
R517 commonsourceibias.n141 commonsourceibias.n122 16.9689
R518 commonsourceibias.n230 commonsourceibias.n211 16.9689
R519 commonsourceibias.n266 commonsourceibias.n265 16.9689
R520 commonsourceibias.n377 commonsourceibias.n358 16.9689
R521 commonsourceibias.n414 commonsourceibias.n413 16.9689
R522 commonsourceibias.n460 commonsourceibias.n459 16.9689
R523 commonsourceibias.n318 commonsourceibias.n299 16.9689
R524 commonsourceibias.n512 commonsourceibias.n493 16.9689
R525 commonsourceibias.n549 commonsourceibias.n548 16.9689
R526 commonsourceibias.n70 commonsourceibias.n69 16.477
R527 commonsourceibias.n63 commonsourceibias.n62 16.477
R528 commonsourceibias.n163 commonsourceibias.n162 16.477
R529 commonsourceibias.n156 commonsourceibias.n155 16.477
R530 commonsourceibias.n245 commonsourceibias.n244 16.477
R531 commonsourceibias.n252 commonsourceibias.n251 16.477
R532 commonsourceibias.n392 commonsourceibias.n391 16.477
R533 commonsourceibias.n399 commonsourceibias.n398 16.477
R534 commonsourceibias.n445 commonsourceibias.n444 16.477
R535 commonsourceibias.n333 commonsourceibias.n332 16.477
R536 commonsourceibias.n527 commonsourceibias.n526 16.477
R537 commonsourceibias.n534 commonsourceibias.n533 16.477
R538 commonsourceibias.n77 commonsourceibias.n76 15.9852
R539 commonsourceibias.n56 commonsourceibias.n27 15.9852
R540 commonsourceibias.n170 commonsourceibias.n169 15.9852
R541 commonsourceibias.n149 commonsourceibias.n120 15.9852
R542 commonsourceibias.n238 commonsourceibias.n209 15.9852
R543 commonsourceibias.n259 commonsourceibias.n258 15.9852
R544 commonsourceibias.n385 commonsourceibias.n356 15.9852
R545 commonsourceibias.n407 commonsourceibias.n406 15.9852
R546 commonsourceibias.n453 commonsourceibias.n452 15.9852
R547 commonsourceibias.n326 commonsourceibias.n297 15.9852
R548 commonsourceibias.n520 commonsourceibias.n491 15.9852
R549 commonsourceibias.n542 commonsourceibias.n541 15.9852
R550 commonsourceibias.n91 commonsourceibias.n90 15.4934
R551 commonsourceibias.n41 commonsourceibias.n40 15.4934
R552 commonsourceibias.n184 commonsourceibias.n183 15.4934
R553 commonsourceibias.n134 commonsourceibias.n133 15.4934
R554 commonsourceibias.n223 commonsourceibias.n222 15.4934
R555 commonsourceibias.n273 commonsourceibias.n272 15.4934
R556 commonsourceibias.n370 commonsourceibias.n369 15.4934
R557 commonsourceibias.n422 commonsourceibias.n421 15.4934
R558 commonsourceibias.n468 commonsourceibias.n467 15.4934
R559 commonsourceibias.n311 commonsourceibias.n310 15.4934
R560 commonsourceibias.n505 commonsourceibias.n504 15.4934
R561 commonsourceibias.n557 commonsourceibias.n556 15.4934
R562 commonsourceibias.n102 commonsourceibias.n100 13.2663
R563 commonsourceibias.n433 commonsourceibias.n431 13.2663
R564 commonsourceibias.n568 commonsourceibias.n283 11.9876
R565 commonsourceibias.n568 commonsourceibias.n567 10.3347
R566 commonsourceibias.n159 commonsourceibias.n116 9.50363
R567 commonsourceibias.n441 commonsourceibias.n440 9.50363
R568 commonsourceibias.n92 commonsourceibias.n91 9.09948
R569 commonsourceibias.n40 commonsourceibias.n39 9.09948
R570 commonsourceibias.n185 commonsourceibias.n184 9.09948
R571 commonsourceibias.n133 commonsourceibias.n132 9.09948
R572 commonsourceibias.n222 commonsourceibias.n221 9.09948
R573 commonsourceibias.n274 commonsourceibias.n273 9.09948
R574 commonsourceibias.n369 commonsourceibias.n368 9.09948
R575 commonsourceibias.n423 commonsourceibias.n422 9.09948
R576 commonsourceibias.n469 commonsourceibias.n468 9.09948
R577 commonsourceibias.n310 commonsourceibias.n309 9.09948
R578 commonsourceibias.n504 commonsourceibias.n503 9.09948
R579 commonsourceibias.n558 commonsourceibias.n557 9.09948
R580 commonsourceibias.n283 commonsourceibias.n193 8.79261
R581 commonsourceibias.n567 commonsourceibias.n477 8.79261
R582 commonsourceibias.n78 commonsourceibias.n77 8.60764
R583 commonsourceibias.n53 commonsourceibias.n27 8.60764
R584 commonsourceibias.n171 commonsourceibias.n170 8.60764
R585 commonsourceibias.n146 commonsourceibias.n120 8.60764
R586 commonsourceibias.n235 commonsourceibias.n209 8.60764
R587 commonsourceibias.n260 commonsourceibias.n259 8.60764
R588 commonsourceibias.n382 commonsourceibias.n356 8.60764
R589 commonsourceibias.n408 commonsourceibias.n407 8.60764
R590 commonsourceibias.n454 commonsourceibias.n453 8.60764
R591 commonsourceibias.n323 commonsourceibias.n297 8.60764
R592 commonsourceibias.n517 commonsourceibias.n491 8.60764
R593 commonsourceibias.n543 commonsourceibias.n542 8.60764
R594 commonsourceibias.n69 commonsourceibias.n68 8.11581
R595 commonsourceibias.n64 commonsourceibias.n63 8.11581
R596 commonsourceibias.n162 commonsourceibias.n161 8.11581
R597 commonsourceibias.n157 commonsourceibias.n156 8.11581
R598 commonsourceibias.n246 commonsourceibias.n245 8.11581
R599 commonsourceibias.n251 commonsourceibias.n250 8.11581
R600 commonsourceibias.n393 commonsourceibias.n392 8.11581
R601 commonsourceibias.n398 commonsourceibias.n397 8.11581
R602 commonsourceibias.n444 commonsourceibias.n443 8.11581
R603 commonsourceibias.n334 commonsourceibias.n333 8.11581
R604 commonsourceibias.n528 commonsourceibias.n527 8.11581
R605 commonsourceibias.n533 commonsourceibias.n532 8.11581
R606 commonsourceibias.n83 commonsourceibias.n82 7.62397
R607 commonsourceibias.n51 commonsourceibias.n29 7.62397
R608 commonsourceibias.n176 commonsourceibias.n175 7.62397
R609 commonsourceibias.n144 commonsourceibias.n122 7.62397
R610 commonsourceibias.n233 commonsourceibias.n211 7.62397
R611 commonsourceibias.n265 commonsourceibias.n264 7.62397
R612 commonsourceibias.n380 commonsourceibias.n358 7.62397
R613 commonsourceibias.n413 commonsourceibias.n412 7.62397
R614 commonsourceibias.n459 commonsourceibias.n458 7.62397
R615 commonsourceibias.n321 commonsourceibias.n299 7.62397
R616 commonsourceibias.n515 commonsourceibias.n493 7.62397
R617 commonsourceibias.n548 commonsourceibias.n547 7.62397
R618 commonsourceibias.n97 commonsourceibias.n96 7.13213
R619 commonsourceibias.n34 commonsourceibias.n33 7.13213
R620 commonsourceibias.n190 commonsourceibias.n189 7.13213
R621 commonsourceibias.n127 commonsourceibias.n126 7.13213
R622 commonsourceibias.n216 commonsourceibias.n215 7.13213
R623 commonsourceibias.n279 commonsourceibias.n278 7.13213
R624 commonsourceibias.n363 commonsourceibias.n362 7.13213
R625 commonsourceibias.n428 commonsourceibias.n427 7.13213
R626 commonsourceibias.n474 commonsourceibias.n473 7.13213
R627 commonsourceibias.n304 commonsourceibias.n303 7.13213
R628 commonsourceibias.n498 commonsourceibias.n497 7.13213
R629 commonsourceibias.n563 commonsourceibias.n562 7.13213
R630 commonsourceibias.n283 commonsourceibias.n282 5.06534
R631 commonsourceibias.n567 commonsourceibias.n566 5.06534
R632 commonsourceibias commonsourceibias.n568 4.04308
R633 commonsourceibias.n109 commonsourceibias.t55 2.82907
R634 commonsourceibias.n109 commonsourceibias.t39 2.82907
R635 commonsourceibias.n110 commonsourceibias.t43 2.82907
R636 commonsourceibias.n110 commonsourceibias.t11 2.82907
R637 commonsourceibias.n112 commonsourceibias.t1 2.82907
R638 commonsourceibias.n112 commonsourceibias.t7 2.82907
R639 commonsourceibias.n114 commonsourceibias.t37 2.82907
R640 commonsourceibias.n114 commonsourceibias.t49 2.82907
R641 commonsourceibias.n107 commonsourceibias.t5 2.82907
R642 commonsourceibias.n107 commonsourceibias.t29 2.82907
R643 commonsourceibias.n105 commonsourceibias.t47 2.82907
R644 commonsourceibias.n105 commonsourceibias.t9 2.82907
R645 commonsourceibias.n103 commonsourceibias.t27 2.82907
R646 commonsourceibias.n103 commonsourceibias.t33 2.82907
R647 commonsourceibias.n101 commonsourceibias.t35 2.82907
R648 commonsourceibias.n101 commonsourceibias.t53 2.82907
R649 commonsourceibias.n432 commonsourceibias.t59 2.82907
R650 commonsourceibias.n432 commonsourceibias.t17 2.82907
R651 commonsourceibias.n434 commonsourceibias.t57 2.82907
R652 commonsourceibias.n434 commonsourceibias.t13 2.82907
R653 commonsourceibias.n436 commonsourceibias.t21 2.82907
R654 commonsourceibias.n436 commonsourceibias.t31 2.82907
R655 commonsourceibias.n438 commonsourceibias.t3 2.82907
R656 commonsourceibias.n438 commonsourceibias.t51 2.82907
R657 commonsourceibias.n341 commonsourceibias.t45 2.82907
R658 commonsourceibias.n341 commonsourceibias.t19 2.82907
R659 commonsourceibias.n339 commonsourceibias.t63 2.82907
R660 commonsourceibias.n339 commonsourceibias.t25 2.82907
R661 commonsourceibias.n337 commonsourceibias.t23 2.82907
R662 commonsourceibias.n337 commonsourceibias.t41 2.82907
R663 commonsourceibias.n336 commonsourceibias.t15 2.82907
R664 commonsourceibias.n336 commonsourceibias.t61 2.82907
R665 commonsourceibias.n17 commonsourceibias.n15 0.738255
R666 commonsourceibias.n46 commonsourceibias.n45 0.738255
R667 commonsourceibias.n5 commonsourceibias.n3 0.738255
R668 commonsourceibias.n139 commonsourceibias.n138 0.738255
R669 commonsourceibias.n228 commonsourceibias.n227 0.738255
R670 commonsourceibias.n199 commonsourceibias.n197 0.738255
R671 commonsourceibias.n375 commonsourceibias.n374 0.738255
R672 commonsourceibias.n415 commonsourceibias.n346 0.738255
R673 commonsourceibias.n461 commonsourceibias.n287 0.738255
R674 commonsourceibias.n316 commonsourceibias.n315 0.738255
R675 commonsourceibias.n510 commonsourceibias.n509 0.738255
R676 commonsourceibias.n550 commonsourceibias.n481 0.738255
R677 commonsourceibias.n104 commonsourceibias.n102 0.573776
R678 commonsourceibias.n106 commonsourceibias.n104 0.573776
R679 commonsourceibias.n108 commonsourceibias.n106 0.573776
R680 commonsourceibias.n115 commonsourceibias.n113 0.573776
R681 commonsourceibias.n113 commonsourceibias.n111 0.573776
R682 commonsourceibias.n340 commonsourceibias.n338 0.573776
R683 commonsourceibias.n342 commonsourceibias.n340 0.573776
R684 commonsourceibias.n439 commonsourceibias.n437 0.573776
R685 commonsourceibias.n437 commonsourceibias.n435 0.573776
R686 commonsourceibias.n435 commonsourceibias.n433 0.573776
R687 commonsourceibias.n116 commonsourceibias.n108 0.287138
R688 commonsourceibias.n116 commonsourceibias.n115 0.287138
R689 commonsourceibias.n440 commonsourceibias.n342 0.287138
R690 commonsourceibias.n440 commonsourceibias.n439 0.287138
R691 commonsourceibias.n100 commonsourceibias.n12 0.285035
R692 commonsourceibias.n193 commonsourceibias.n0 0.285035
R693 commonsourceibias.n282 commonsourceibias.n194 0.285035
R694 commonsourceibias.n431 commonsourceibias.n343 0.285035
R695 commonsourceibias.n477 commonsourceibias.n284 0.285035
R696 commonsourceibias.n566 commonsourceibias.n478 0.285035
R697 commonsourceibias.n22 commonsourceibias.n20 0.246418
R698 commonsourceibias.n58 commonsourceibias.n25 0.246418
R699 commonsourceibias.n10 commonsourceibias.n8 0.246418
R700 commonsourceibias.n151 commonsourceibias.n118 0.246418
R701 commonsourceibias.n240 commonsourceibias.n207 0.246418
R702 commonsourceibias.n204 commonsourceibias.n202 0.246418
R703 commonsourceibias.n387 commonsourceibias.n354 0.246418
R704 commonsourceibias.n400 commonsourceibias.n350 0.246418
R705 commonsourceibias.n446 commonsourceibias.n291 0.246418
R706 commonsourceibias.n328 commonsourceibias.n295 0.246418
R707 commonsourceibias.n522 commonsourceibias.n489 0.246418
R708 commonsourceibias.n535 commonsourceibias.n485 0.246418
R709 commonsourceibias.n95 commonsourceibias.n12 0.189894
R710 commonsourceibias.n95 commonsourceibias.n94 0.189894
R711 commonsourceibias.n94 commonsourceibias.n93 0.189894
R712 commonsourceibias.n93 commonsourceibias.n14 0.189894
R713 commonsourceibias.n88 commonsourceibias.n14 0.189894
R714 commonsourceibias.n88 commonsourceibias.n87 0.189894
R715 commonsourceibias.n87 commonsourceibias.n86 0.189894
R716 commonsourceibias.n86 commonsourceibias.n16 0.189894
R717 commonsourceibias.n81 commonsourceibias.n16 0.189894
R718 commonsourceibias.n81 commonsourceibias.n80 0.189894
R719 commonsourceibias.n80 commonsourceibias.n79 0.189894
R720 commonsourceibias.n79 commonsourceibias.n19 0.189894
R721 commonsourceibias.n74 commonsourceibias.n19 0.189894
R722 commonsourceibias.n74 commonsourceibias.n73 0.189894
R723 commonsourceibias.n73 commonsourceibias.n72 0.189894
R724 commonsourceibias.n72 commonsourceibias.n21 0.189894
R725 commonsourceibias.n67 commonsourceibias.n21 0.189894
R726 commonsourceibias.n67 commonsourceibias.n66 0.189894
R727 commonsourceibias.n66 commonsourceibias.n65 0.189894
R728 commonsourceibias.n65 commonsourceibias.n24 0.189894
R729 commonsourceibias.n60 commonsourceibias.n24 0.189894
R730 commonsourceibias.n60 commonsourceibias.n59 0.189894
R731 commonsourceibias.n59 commonsourceibias.n26 0.189894
R732 commonsourceibias.n55 commonsourceibias.n26 0.189894
R733 commonsourceibias.n55 commonsourceibias.n54 0.189894
R734 commonsourceibias.n54 commonsourceibias.n28 0.189894
R735 commonsourceibias.n50 commonsourceibias.n28 0.189894
R736 commonsourceibias.n50 commonsourceibias.n49 0.189894
R737 commonsourceibias.n49 commonsourceibias.n30 0.189894
R738 commonsourceibias.n44 commonsourceibias.n30 0.189894
R739 commonsourceibias.n44 commonsourceibias.n43 0.189894
R740 commonsourceibias.n43 commonsourceibias.n42 0.189894
R741 commonsourceibias.n42 commonsourceibias.n32 0.189894
R742 commonsourceibias.n37 commonsourceibias.n32 0.189894
R743 commonsourceibias.n37 commonsourceibias.n36 0.189894
R744 commonsourceibias.n158 commonsourceibias.n117 0.189894
R745 commonsourceibias.n153 commonsourceibias.n117 0.189894
R746 commonsourceibias.n153 commonsourceibias.n152 0.189894
R747 commonsourceibias.n152 commonsourceibias.n119 0.189894
R748 commonsourceibias.n148 commonsourceibias.n119 0.189894
R749 commonsourceibias.n148 commonsourceibias.n147 0.189894
R750 commonsourceibias.n147 commonsourceibias.n121 0.189894
R751 commonsourceibias.n143 commonsourceibias.n121 0.189894
R752 commonsourceibias.n143 commonsourceibias.n142 0.189894
R753 commonsourceibias.n142 commonsourceibias.n123 0.189894
R754 commonsourceibias.n137 commonsourceibias.n123 0.189894
R755 commonsourceibias.n137 commonsourceibias.n136 0.189894
R756 commonsourceibias.n136 commonsourceibias.n135 0.189894
R757 commonsourceibias.n135 commonsourceibias.n125 0.189894
R758 commonsourceibias.n130 commonsourceibias.n125 0.189894
R759 commonsourceibias.n130 commonsourceibias.n129 0.189894
R760 commonsourceibias.n188 commonsourceibias.n0 0.189894
R761 commonsourceibias.n188 commonsourceibias.n187 0.189894
R762 commonsourceibias.n187 commonsourceibias.n186 0.189894
R763 commonsourceibias.n186 commonsourceibias.n2 0.189894
R764 commonsourceibias.n181 commonsourceibias.n2 0.189894
R765 commonsourceibias.n181 commonsourceibias.n180 0.189894
R766 commonsourceibias.n180 commonsourceibias.n179 0.189894
R767 commonsourceibias.n179 commonsourceibias.n4 0.189894
R768 commonsourceibias.n174 commonsourceibias.n4 0.189894
R769 commonsourceibias.n174 commonsourceibias.n173 0.189894
R770 commonsourceibias.n173 commonsourceibias.n172 0.189894
R771 commonsourceibias.n172 commonsourceibias.n7 0.189894
R772 commonsourceibias.n167 commonsourceibias.n7 0.189894
R773 commonsourceibias.n167 commonsourceibias.n166 0.189894
R774 commonsourceibias.n166 commonsourceibias.n165 0.189894
R775 commonsourceibias.n165 commonsourceibias.n9 0.189894
R776 commonsourceibias.n160 commonsourceibias.n9 0.189894
R777 commonsourceibias.n277 commonsourceibias.n194 0.189894
R778 commonsourceibias.n277 commonsourceibias.n276 0.189894
R779 commonsourceibias.n276 commonsourceibias.n275 0.189894
R780 commonsourceibias.n275 commonsourceibias.n196 0.189894
R781 commonsourceibias.n270 commonsourceibias.n196 0.189894
R782 commonsourceibias.n270 commonsourceibias.n269 0.189894
R783 commonsourceibias.n269 commonsourceibias.n268 0.189894
R784 commonsourceibias.n268 commonsourceibias.n198 0.189894
R785 commonsourceibias.n263 commonsourceibias.n198 0.189894
R786 commonsourceibias.n263 commonsourceibias.n262 0.189894
R787 commonsourceibias.n262 commonsourceibias.n261 0.189894
R788 commonsourceibias.n261 commonsourceibias.n201 0.189894
R789 commonsourceibias.n256 commonsourceibias.n201 0.189894
R790 commonsourceibias.n256 commonsourceibias.n255 0.189894
R791 commonsourceibias.n255 commonsourceibias.n254 0.189894
R792 commonsourceibias.n254 commonsourceibias.n203 0.189894
R793 commonsourceibias.n249 commonsourceibias.n203 0.189894
R794 commonsourceibias.n249 commonsourceibias.n248 0.189894
R795 commonsourceibias.n248 commonsourceibias.n247 0.189894
R796 commonsourceibias.n247 commonsourceibias.n206 0.189894
R797 commonsourceibias.n242 commonsourceibias.n206 0.189894
R798 commonsourceibias.n242 commonsourceibias.n241 0.189894
R799 commonsourceibias.n241 commonsourceibias.n208 0.189894
R800 commonsourceibias.n237 commonsourceibias.n208 0.189894
R801 commonsourceibias.n237 commonsourceibias.n236 0.189894
R802 commonsourceibias.n236 commonsourceibias.n210 0.189894
R803 commonsourceibias.n232 commonsourceibias.n210 0.189894
R804 commonsourceibias.n232 commonsourceibias.n231 0.189894
R805 commonsourceibias.n231 commonsourceibias.n212 0.189894
R806 commonsourceibias.n226 commonsourceibias.n212 0.189894
R807 commonsourceibias.n226 commonsourceibias.n225 0.189894
R808 commonsourceibias.n225 commonsourceibias.n224 0.189894
R809 commonsourceibias.n224 commonsourceibias.n214 0.189894
R810 commonsourceibias.n219 commonsourceibias.n214 0.189894
R811 commonsourceibias.n219 commonsourceibias.n218 0.189894
R812 commonsourceibias.n366 commonsourceibias.n365 0.189894
R813 commonsourceibias.n366 commonsourceibias.n361 0.189894
R814 commonsourceibias.n371 commonsourceibias.n361 0.189894
R815 commonsourceibias.n372 commonsourceibias.n371 0.189894
R816 commonsourceibias.n373 commonsourceibias.n372 0.189894
R817 commonsourceibias.n373 commonsourceibias.n359 0.189894
R818 commonsourceibias.n378 commonsourceibias.n359 0.189894
R819 commonsourceibias.n379 commonsourceibias.n378 0.189894
R820 commonsourceibias.n379 commonsourceibias.n357 0.189894
R821 commonsourceibias.n383 commonsourceibias.n357 0.189894
R822 commonsourceibias.n384 commonsourceibias.n383 0.189894
R823 commonsourceibias.n384 commonsourceibias.n355 0.189894
R824 commonsourceibias.n388 commonsourceibias.n355 0.189894
R825 commonsourceibias.n389 commonsourceibias.n388 0.189894
R826 commonsourceibias.n389 commonsourceibias.n353 0.189894
R827 commonsourceibias.n394 commonsourceibias.n353 0.189894
R828 commonsourceibias.n395 commonsourceibias.n394 0.189894
R829 commonsourceibias.n396 commonsourceibias.n395 0.189894
R830 commonsourceibias.n396 commonsourceibias.n351 0.189894
R831 commonsourceibias.n402 commonsourceibias.n351 0.189894
R832 commonsourceibias.n403 commonsourceibias.n402 0.189894
R833 commonsourceibias.n404 commonsourceibias.n403 0.189894
R834 commonsourceibias.n404 commonsourceibias.n349 0.189894
R835 commonsourceibias.n409 commonsourceibias.n349 0.189894
R836 commonsourceibias.n410 commonsourceibias.n409 0.189894
R837 commonsourceibias.n411 commonsourceibias.n410 0.189894
R838 commonsourceibias.n411 commonsourceibias.n347 0.189894
R839 commonsourceibias.n417 commonsourceibias.n347 0.189894
R840 commonsourceibias.n418 commonsourceibias.n417 0.189894
R841 commonsourceibias.n419 commonsourceibias.n418 0.189894
R842 commonsourceibias.n419 commonsourceibias.n345 0.189894
R843 commonsourceibias.n424 commonsourceibias.n345 0.189894
R844 commonsourceibias.n425 commonsourceibias.n424 0.189894
R845 commonsourceibias.n426 commonsourceibias.n425 0.189894
R846 commonsourceibias.n426 commonsourceibias.n343 0.189894
R847 commonsourceibias.n307 commonsourceibias.n306 0.189894
R848 commonsourceibias.n307 commonsourceibias.n302 0.189894
R849 commonsourceibias.n312 commonsourceibias.n302 0.189894
R850 commonsourceibias.n313 commonsourceibias.n312 0.189894
R851 commonsourceibias.n314 commonsourceibias.n313 0.189894
R852 commonsourceibias.n314 commonsourceibias.n300 0.189894
R853 commonsourceibias.n319 commonsourceibias.n300 0.189894
R854 commonsourceibias.n320 commonsourceibias.n319 0.189894
R855 commonsourceibias.n320 commonsourceibias.n298 0.189894
R856 commonsourceibias.n324 commonsourceibias.n298 0.189894
R857 commonsourceibias.n325 commonsourceibias.n324 0.189894
R858 commonsourceibias.n325 commonsourceibias.n296 0.189894
R859 commonsourceibias.n329 commonsourceibias.n296 0.189894
R860 commonsourceibias.n330 commonsourceibias.n329 0.189894
R861 commonsourceibias.n330 commonsourceibias.n294 0.189894
R862 commonsourceibias.n335 commonsourceibias.n294 0.189894
R863 commonsourceibias.n442 commonsourceibias.n292 0.189894
R864 commonsourceibias.n448 commonsourceibias.n292 0.189894
R865 commonsourceibias.n449 commonsourceibias.n448 0.189894
R866 commonsourceibias.n450 commonsourceibias.n449 0.189894
R867 commonsourceibias.n450 commonsourceibias.n290 0.189894
R868 commonsourceibias.n455 commonsourceibias.n290 0.189894
R869 commonsourceibias.n456 commonsourceibias.n455 0.189894
R870 commonsourceibias.n457 commonsourceibias.n456 0.189894
R871 commonsourceibias.n457 commonsourceibias.n288 0.189894
R872 commonsourceibias.n463 commonsourceibias.n288 0.189894
R873 commonsourceibias.n464 commonsourceibias.n463 0.189894
R874 commonsourceibias.n465 commonsourceibias.n464 0.189894
R875 commonsourceibias.n465 commonsourceibias.n286 0.189894
R876 commonsourceibias.n470 commonsourceibias.n286 0.189894
R877 commonsourceibias.n471 commonsourceibias.n470 0.189894
R878 commonsourceibias.n472 commonsourceibias.n471 0.189894
R879 commonsourceibias.n472 commonsourceibias.n284 0.189894
R880 commonsourceibias.n501 commonsourceibias.n500 0.189894
R881 commonsourceibias.n501 commonsourceibias.n496 0.189894
R882 commonsourceibias.n506 commonsourceibias.n496 0.189894
R883 commonsourceibias.n507 commonsourceibias.n506 0.189894
R884 commonsourceibias.n508 commonsourceibias.n507 0.189894
R885 commonsourceibias.n508 commonsourceibias.n494 0.189894
R886 commonsourceibias.n513 commonsourceibias.n494 0.189894
R887 commonsourceibias.n514 commonsourceibias.n513 0.189894
R888 commonsourceibias.n514 commonsourceibias.n492 0.189894
R889 commonsourceibias.n518 commonsourceibias.n492 0.189894
R890 commonsourceibias.n519 commonsourceibias.n518 0.189894
R891 commonsourceibias.n519 commonsourceibias.n490 0.189894
R892 commonsourceibias.n523 commonsourceibias.n490 0.189894
R893 commonsourceibias.n524 commonsourceibias.n523 0.189894
R894 commonsourceibias.n524 commonsourceibias.n488 0.189894
R895 commonsourceibias.n529 commonsourceibias.n488 0.189894
R896 commonsourceibias.n530 commonsourceibias.n529 0.189894
R897 commonsourceibias.n531 commonsourceibias.n530 0.189894
R898 commonsourceibias.n531 commonsourceibias.n486 0.189894
R899 commonsourceibias.n537 commonsourceibias.n486 0.189894
R900 commonsourceibias.n538 commonsourceibias.n537 0.189894
R901 commonsourceibias.n539 commonsourceibias.n538 0.189894
R902 commonsourceibias.n539 commonsourceibias.n484 0.189894
R903 commonsourceibias.n544 commonsourceibias.n484 0.189894
R904 commonsourceibias.n545 commonsourceibias.n544 0.189894
R905 commonsourceibias.n546 commonsourceibias.n545 0.189894
R906 commonsourceibias.n546 commonsourceibias.n482 0.189894
R907 commonsourceibias.n552 commonsourceibias.n482 0.189894
R908 commonsourceibias.n553 commonsourceibias.n552 0.189894
R909 commonsourceibias.n554 commonsourceibias.n553 0.189894
R910 commonsourceibias.n554 commonsourceibias.n480 0.189894
R911 commonsourceibias.n559 commonsourceibias.n480 0.189894
R912 commonsourceibias.n560 commonsourceibias.n559 0.189894
R913 commonsourceibias.n561 commonsourceibias.n560 0.189894
R914 commonsourceibias.n561 commonsourceibias.n478 0.189894
R915 commonsourceibias.n159 commonsourceibias.n158 0.170955
R916 commonsourceibias.n160 commonsourceibias.n159 0.170955
R917 commonsourceibias.n441 commonsourceibias.n335 0.170955
R918 commonsourceibias.n442 commonsourceibias.n441 0.170955
R919 CSoutput.n19 CSoutput.t188 184.661
R920 CSoutput.n78 CSoutput.n77 165.8
R921 CSoutput.n76 CSoutput.n0 165.8
R922 CSoutput.n75 CSoutput.n74 165.8
R923 CSoutput.n73 CSoutput.n72 165.8
R924 CSoutput.n71 CSoutput.n2 165.8
R925 CSoutput.n69 CSoutput.n68 165.8
R926 CSoutput.n67 CSoutput.n3 165.8
R927 CSoutput.n66 CSoutput.n65 165.8
R928 CSoutput.n63 CSoutput.n4 165.8
R929 CSoutput.n61 CSoutput.n60 165.8
R930 CSoutput.n59 CSoutput.n5 165.8
R931 CSoutput.n58 CSoutput.n57 165.8
R932 CSoutput.n55 CSoutput.n6 165.8
R933 CSoutput.n54 CSoutput.n53 165.8
R934 CSoutput.n52 CSoutput.n51 165.8
R935 CSoutput.n50 CSoutput.n8 165.8
R936 CSoutput.n48 CSoutput.n47 165.8
R937 CSoutput.n46 CSoutput.n9 165.8
R938 CSoutput.n45 CSoutput.n44 165.8
R939 CSoutput.n42 CSoutput.n10 165.8
R940 CSoutput.n41 CSoutput.n40 165.8
R941 CSoutput.n39 CSoutput.n38 165.8
R942 CSoutput.n37 CSoutput.n12 165.8
R943 CSoutput.n35 CSoutput.n34 165.8
R944 CSoutput.n33 CSoutput.n13 165.8
R945 CSoutput.n32 CSoutput.n31 165.8
R946 CSoutput.n29 CSoutput.n14 165.8
R947 CSoutput.n28 CSoutput.n27 165.8
R948 CSoutput.n26 CSoutput.n25 165.8
R949 CSoutput.n24 CSoutput.n16 165.8
R950 CSoutput.n22 CSoutput.n21 165.8
R951 CSoutput.n20 CSoutput.n17 165.8
R952 CSoutput.n77 CSoutput.t190 162.194
R953 CSoutput.n18 CSoutput.t205 120.501
R954 CSoutput.n23 CSoutput.t199 120.501
R955 CSoutput.n15 CSoutput.t196 120.501
R956 CSoutput.n30 CSoutput.t185 120.501
R957 CSoutput.n36 CSoutput.t187 120.501
R958 CSoutput.n11 CSoutput.t197 120.501
R959 CSoutput.n43 CSoutput.t195 120.501
R960 CSoutput.n49 CSoutput.t189 120.501
R961 CSoutput.n7 CSoutput.t200 120.501
R962 CSoutput.n56 CSoutput.t201 120.501
R963 CSoutput.n62 CSoutput.t192 120.501
R964 CSoutput.n64 CSoutput.t202 120.501
R965 CSoutput.n70 CSoutput.t204 120.501
R966 CSoutput.n1 CSoutput.t198 120.501
R967 CSoutput.n330 CSoutput.n328 103.469
R968 CSoutput.n310 CSoutput.n308 103.469
R969 CSoutput.n291 CSoutput.n289 103.469
R970 CSoutput.n120 CSoutput.n118 103.469
R971 CSoutput.n100 CSoutput.n98 103.469
R972 CSoutput.n81 CSoutput.n79 103.469
R973 CSoutput.n344 CSoutput.n343 103.111
R974 CSoutput.n342 CSoutput.n341 103.111
R975 CSoutput.n340 CSoutput.n339 103.111
R976 CSoutput.n338 CSoutput.n337 103.111
R977 CSoutput.n336 CSoutput.n335 103.111
R978 CSoutput.n334 CSoutput.n333 103.111
R979 CSoutput.n332 CSoutput.n331 103.111
R980 CSoutput.n330 CSoutput.n329 103.111
R981 CSoutput.n326 CSoutput.n325 103.111
R982 CSoutput.n324 CSoutput.n323 103.111
R983 CSoutput.n322 CSoutput.n321 103.111
R984 CSoutput.n320 CSoutput.n319 103.111
R985 CSoutput.n318 CSoutput.n317 103.111
R986 CSoutput.n316 CSoutput.n315 103.111
R987 CSoutput.n314 CSoutput.n313 103.111
R988 CSoutput.n312 CSoutput.n311 103.111
R989 CSoutput.n310 CSoutput.n309 103.111
R990 CSoutput.n307 CSoutput.n306 103.111
R991 CSoutput.n305 CSoutput.n304 103.111
R992 CSoutput.n303 CSoutput.n302 103.111
R993 CSoutput.n301 CSoutput.n300 103.111
R994 CSoutput.n299 CSoutput.n298 103.111
R995 CSoutput.n297 CSoutput.n296 103.111
R996 CSoutput.n295 CSoutput.n294 103.111
R997 CSoutput.n293 CSoutput.n292 103.111
R998 CSoutput.n291 CSoutput.n290 103.111
R999 CSoutput.n120 CSoutput.n119 103.111
R1000 CSoutput.n122 CSoutput.n121 103.111
R1001 CSoutput.n124 CSoutput.n123 103.111
R1002 CSoutput.n126 CSoutput.n125 103.111
R1003 CSoutput.n128 CSoutput.n127 103.111
R1004 CSoutput.n130 CSoutput.n129 103.111
R1005 CSoutput.n132 CSoutput.n131 103.111
R1006 CSoutput.n134 CSoutput.n133 103.111
R1007 CSoutput.n136 CSoutput.n135 103.111
R1008 CSoutput.n100 CSoutput.n99 103.111
R1009 CSoutput.n102 CSoutput.n101 103.111
R1010 CSoutput.n104 CSoutput.n103 103.111
R1011 CSoutput.n106 CSoutput.n105 103.111
R1012 CSoutput.n108 CSoutput.n107 103.111
R1013 CSoutput.n110 CSoutput.n109 103.111
R1014 CSoutput.n112 CSoutput.n111 103.111
R1015 CSoutput.n114 CSoutput.n113 103.111
R1016 CSoutput.n116 CSoutput.n115 103.111
R1017 CSoutput.n81 CSoutput.n80 103.111
R1018 CSoutput.n83 CSoutput.n82 103.111
R1019 CSoutput.n85 CSoutput.n84 103.111
R1020 CSoutput.n87 CSoutput.n86 103.111
R1021 CSoutput.n89 CSoutput.n88 103.111
R1022 CSoutput.n91 CSoutput.n90 103.111
R1023 CSoutput.n93 CSoutput.n92 103.111
R1024 CSoutput.n95 CSoutput.n94 103.111
R1025 CSoutput.n97 CSoutput.n96 103.111
R1026 CSoutput.n346 CSoutput.n345 103.111
R1027 CSoutput.n366 CSoutput.n364 81.5057
R1028 CSoutput.n351 CSoutput.n349 81.5057
R1029 CSoutput.n398 CSoutput.n396 81.5057
R1030 CSoutput.n383 CSoutput.n381 81.5057
R1031 CSoutput.n378 CSoutput.n377 80.9324
R1032 CSoutput.n376 CSoutput.n375 80.9324
R1033 CSoutput.n374 CSoutput.n373 80.9324
R1034 CSoutput.n372 CSoutput.n371 80.9324
R1035 CSoutput.n370 CSoutput.n369 80.9324
R1036 CSoutput.n368 CSoutput.n367 80.9324
R1037 CSoutput.n366 CSoutput.n365 80.9324
R1038 CSoutput.n363 CSoutput.n362 80.9324
R1039 CSoutput.n361 CSoutput.n360 80.9324
R1040 CSoutput.n359 CSoutput.n358 80.9324
R1041 CSoutput.n357 CSoutput.n356 80.9324
R1042 CSoutput.n355 CSoutput.n354 80.9324
R1043 CSoutput.n353 CSoutput.n352 80.9324
R1044 CSoutput.n351 CSoutput.n350 80.9324
R1045 CSoutput.n398 CSoutput.n397 80.9324
R1046 CSoutput.n400 CSoutput.n399 80.9324
R1047 CSoutput.n402 CSoutput.n401 80.9324
R1048 CSoutput.n404 CSoutput.n403 80.9324
R1049 CSoutput.n406 CSoutput.n405 80.9324
R1050 CSoutput.n408 CSoutput.n407 80.9324
R1051 CSoutput.n410 CSoutput.n409 80.9324
R1052 CSoutput.n383 CSoutput.n382 80.9324
R1053 CSoutput.n385 CSoutput.n384 80.9324
R1054 CSoutput.n387 CSoutput.n386 80.9324
R1055 CSoutput.n389 CSoutput.n388 80.9324
R1056 CSoutput.n391 CSoutput.n390 80.9324
R1057 CSoutput.n393 CSoutput.n392 80.9324
R1058 CSoutput.n395 CSoutput.n394 80.9324
R1059 CSoutput.n25 CSoutput.n24 48.1486
R1060 CSoutput.n69 CSoutput.n3 48.1486
R1061 CSoutput.n38 CSoutput.n37 48.1486
R1062 CSoutput.n42 CSoutput.n41 48.1486
R1063 CSoutput.n51 CSoutput.n50 48.1486
R1064 CSoutput.n55 CSoutput.n54 48.1486
R1065 CSoutput.n22 CSoutput.n17 46.462
R1066 CSoutput.n72 CSoutput.n71 46.462
R1067 CSoutput.n20 CSoutput.n19 44.9055
R1068 CSoutput.n29 CSoutput.n28 43.7635
R1069 CSoutput.n65 CSoutput.n63 43.7635
R1070 CSoutput.n35 CSoutput.n13 41.7396
R1071 CSoutput.n57 CSoutput.n5 41.7396
R1072 CSoutput.n44 CSoutput.n9 37.0171
R1073 CSoutput.n48 CSoutput.n9 37.0171
R1074 CSoutput.n76 CSoutput.n75 34.9932
R1075 CSoutput.n31 CSoutput.n13 32.2947
R1076 CSoutput.n61 CSoutput.n5 32.2947
R1077 CSoutput.n30 CSoutput.n29 29.6014
R1078 CSoutput.n63 CSoutput.n62 29.6014
R1079 CSoutput.n19 CSoutput.n18 28.4085
R1080 CSoutput.n18 CSoutput.n17 25.1176
R1081 CSoutput.n72 CSoutput.n1 25.1176
R1082 CSoutput.n43 CSoutput.n42 22.0922
R1083 CSoutput.n50 CSoutput.n49 22.0922
R1084 CSoutput.n77 CSoutput.n76 21.8586
R1085 CSoutput.n37 CSoutput.n36 18.9681
R1086 CSoutput.n56 CSoutput.n55 18.9681
R1087 CSoutput.n25 CSoutput.n15 17.6292
R1088 CSoutput.n64 CSoutput.n3 17.6292
R1089 CSoutput.n24 CSoutput.n23 15.844
R1090 CSoutput.n70 CSoutput.n69 15.844
R1091 CSoutput.n38 CSoutput.n11 14.5051
R1092 CSoutput.n54 CSoutput.n7 14.5051
R1093 CSoutput.n413 CSoutput.n78 11.6139
R1094 CSoutput.n41 CSoutput.n11 11.3811
R1095 CSoutput.n51 CSoutput.n7 11.3811
R1096 CSoutput.n23 CSoutput.n22 10.0422
R1097 CSoutput.n71 CSoutput.n70 10.0422
R1098 CSoutput.n327 CSoutput.n307 9.25285
R1099 CSoutput.n117 CSoutput.n97 9.25285
R1100 CSoutput.n379 CSoutput.n363 8.97993
R1101 CSoutput.n411 CSoutput.n395 8.97993
R1102 CSoutput.n380 CSoutput.n348 8.78291
R1103 CSoutput.n28 CSoutput.n15 8.25698
R1104 CSoutput.n65 CSoutput.n64 8.25698
R1105 CSoutput.n380 CSoutput.n379 7.89345
R1106 CSoutput.n412 CSoutput.n411 7.89345
R1107 CSoutput.n348 CSoutput.n347 7.12641
R1108 CSoutput.n138 CSoutput.n137 7.12641
R1109 CSoutput.n36 CSoutput.n35 6.91809
R1110 CSoutput.n57 CSoutput.n56 6.91809
R1111 CSoutput.n379 CSoutput.n378 5.25266
R1112 CSoutput.n411 CSoutput.n410 5.25266
R1113 CSoutput.n413 CSoutput.n138 5.19047
R1114 CSoutput.n347 CSoutput.n346 5.1449
R1115 CSoutput.n327 CSoutput.n326 5.1449
R1116 CSoutput.n137 CSoutput.n136 5.1449
R1117 CSoutput.n117 CSoutput.n116 5.1449
R1118 CSoutput.n229 CSoutput.n182 4.5005
R1119 CSoutput.n198 CSoutput.n182 4.5005
R1120 CSoutput.n193 CSoutput.n177 4.5005
R1121 CSoutput.n193 CSoutput.n179 4.5005
R1122 CSoutput.n193 CSoutput.n176 4.5005
R1123 CSoutput.n193 CSoutput.n180 4.5005
R1124 CSoutput.n193 CSoutput.n175 4.5005
R1125 CSoutput.n193 CSoutput.t203 4.5005
R1126 CSoutput.n193 CSoutput.n174 4.5005
R1127 CSoutput.n193 CSoutput.n181 4.5005
R1128 CSoutput.n193 CSoutput.n182 4.5005
R1129 CSoutput.n191 CSoutput.n177 4.5005
R1130 CSoutput.n191 CSoutput.n179 4.5005
R1131 CSoutput.n191 CSoutput.n176 4.5005
R1132 CSoutput.n191 CSoutput.n180 4.5005
R1133 CSoutput.n191 CSoutput.n175 4.5005
R1134 CSoutput.n191 CSoutput.t203 4.5005
R1135 CSoutput.n191 CSoutput.n174 4.5005
R1136 CSoutput.n191 CSoutput.n181 4.5005
R1137 CSoutput.n191 CSoutput.n182 4.5005
R1138 CSoutput.n190 CSoutput.n177 4.5005
R1139 CSoutput.n190 CSoutput.n179 4.5005
R1140 CSoutput.n190 CSoutput.n176 4.5005
R1141 CSoutput.n190 CSoutput.n180 4.5005
R1142 CSoutput.n190 CSoutput.n175 4.5005
R1143 CSoutput.n190 CSoutput.t203 4.5005
R1144 CSoutput.n190 CSoutput.n174 4.5005
R1145 CSoutput.n190 CSoutput.n181 4.5005
R1146 CSoutput.n190 CSoutput.n182 4.5005
R1147 CSoutput.n275 CSoutput.n177 4.5005
R1148 CSoutput.n275 CSoutput.n179 4.5005
R1149 CSoutput.n275 CSoutput.n176 4.5005
R1150 CSoutput.n275 CSoutput.n180 4.5005
R1151 CSoutput.n275 CSoutput.n175 4.5005
R1152 CSoutput.n275 CSoutput.t203 4.5005
R1153 CSoutput.n275 CSoutput.n174 4.5005
R1154 CSoutput.n275 CSoutput.n181 4.5005
R1155 CSoutput.n275 CSoutput.n182 4.5005
R1156 CSoutput.n273 CSoutput.n177 4.5005
R1157 CSoutput.n273 CSoutput.n179 4.5005
R1158 CSoutput.n273 CSoutput.n176 4.5005
R1159 CSoutput.n273 CSoutput.n180 4.5005
R1160 CSoutput.n273 CSoutput.n175 4.5005
R1161 CSoutput.n273 CSoutput.t203 4.5005
R1162 CSoutput.n273 CSoutput.n174 4.5005
R1163 CSoutput.n273 CSoutput.n181 4.5005
R1164 CSoutput.n271 CSoutput.n177 4.5005
R1165 CSoutput.n271 CSoutput.n179 4.5005
R1166 CSoutput.n271 CSoutput.n176 4.5005
R1167 CSoutput.n271 CSoutput.n180 4.5005
R1168 CSoutput.n271 CSoutput.n175 4.5005
R1169 CSoutput.n271 CSoutput.t203 4.5005
R1170 CSoutput.n271 CSoutput.n174 4.5005
R1171 CSoutput.n271 CSoutput.n181 4.5005
R1172 CSoutput.n201 CSoutput.n177 4.5005
R1173 CSoutput.n201 CSoutput.n179 4.5005
R1174 CSoutput.n201 CSoutput.n176 4.5005
R1175 CSoutput.n201 CSoutput.n180 4.5005
R1176 CSoutput.n201 CSoutput.n175 4.5005
R1177 CSoutput.n201 CSoutput.t203 4.5005
R1178 CSoutput.n201 CSoutput.n174 4.5005
R1179 CSoutput.n201 CSoutput.n181 4.5005
R1180 CSoutput.n201 CSoutput.n182 4.5005
R1181 CSoutput.n200 CSoutput.n177 4.5005
R1182 CSoutput.n200 CSoutput.n179 4.5005
R1183 CSoutput.n200 CSoutput.n176 4.5005
R1184 CSoutput.n200 CSoutput.n180 4.5005
R1185 CSoutput.n200 CSoutput.n175 4.5005
R1186 CSoutput.n200 CSoutput.t203 4.5005
R1187 CSoutput.n200 CSoutput.n174 4.5005
R1188 CSoutput.n200 CSoutput.n181 4.5005
R1189 CSoutput.n200 CSoutput.n182 4.5005
R1190 CSoutput.n204 CSoutput.n177 4.5005
R1191 CSoutput.n204 CSoutput.n179 4.5005
R1192 CSoutput.n204 CSoutput.n176 4.5005
R1193 CSoutput.n204 CSoutput.n180 4.5005
R1194 CSoutput.n204 CSoutput.n175 4.5005
R1195 CSoutput.n204 CSoutput.t203 4.5005
R1196 CSoutput.n204 CSoutput.n174 4.5005
R1197 CSoutput.n204 CSoutput.n181 4.5005
R1198 CSoutput.n204 CSoutput.n182 4.5005
R1199 CSoutput.n203 CSoutput.n177 4.5005
R1200 CSoutput.n203 CSoutput.n179 4.5005
R1201 CSoutput.n203 CSoutput.n176 4.5005
R1202 CSoutput.n203 CSoutput.n180 4.5005
R1203 CSoutput.n203 CSoutput.n175 4.5005
R1204 CSoutput.n203 CSoutput.t203 4.5005
R1205 CSoutput.n203 CSoutput.n174 4.5005
R1206 CSoutput.n203 CSoutput.n181 4.5005
R1207 CSoutput.n203 CSoutput.n182 4.5005
R1208 CSoutput.n186 CSoutput.n177 4.5005
R1209 CSoutput.n186 CSoutput.n179 4.5005
R1210 CSoutput.n186 CSoutput.n176 4.5005
R1211 CSoutput.n186 CSoutput.n180 4.5005
R1212 CSoutput.n186 CSoutput.n175 4.5005
R1213 CSoutput.n186 CSoutput.t203 4.5005
R1214 CSoutput.n186 CSoutput.n174 4.5005
R1215 CSoutput.n186 CSoutput.n181 4.5005
R1216 CSoutput.n186 CSoutput.n182 4.5005
R1217 CSoutput.n278 CSoutput.n177 4.5005
R1218 CSoutput.n278 CSoutput.n179 4.5005
R1219 CSoutput.n278 CSoutput.n176 4.5005
R1220 CSoutput.n278 CSoutput.n180 4.5005
R1221 CSoutput.n278 CSoutput.n175 4.5005
R1222 CSoutput.n278 CSoutput.t203 4.5005
R1223 CSoutput.n278 CSoutput.n174 4.5005
R1224 CSoutput.n278 CSoutput.n181 4.5005
R1225 CSoutput.n278 CSoutput.n182 4.5005
R1226 CSoutput.n265 CSoutput.n236 4.5005
R1227 CSoutput.n265 CSoutput.n242 4.5005
R1228 CSoutput.n223 CSoutput.n212 4.5005
R1229 CSoutput.n223 CSoutput.n214 4.5005
R1230 CSoutput.n223 CSoutput.n211 4.5005
R1231 CSoutput.n223 CSoutput.n215 4.5005
R1232 CSoutput.n223 CSoutput.n210 4.5005
R1233 CSoutput.n223 CSoutput.t184 4.5005
R1234 CSoutput.n223 CSoutput.n209 4.5005
R1235 CSoutput.n223 CSoutput.n216 4.5005
R1236 CSoutput.n265 CSoutput.n223 4.5005
R1237 CSoutput.n244 CSoutput.n212 4.5005
R1238 CSoutput.n244 CSoutput.n214 4.5005
R1239 CSoutput.n244 CSoutput.n211 4.5005
R1240 CSoutput.n244 CSoutput.n215 4.5005
R1241 CSoutput.n244 CSoutput.n210 4.5005
R1242 CSoutput.n244 CSoutput.t184 4.5005
R1243 CSoutput.n244 CSoutput.n209 4.5005
R1244 CSoutput.n244 CSoutput.n216 4.5005
R1245 CSoutput.n265 CSoutput.n244 4.5005
R1246 CSoutput.n222 CSoutput.n212 4.5005
R1247 CSoutput.n222 CSoutput.n214 4.5005
R1248 CSoutput.n222 CSoutput.n211 4.5005
R1249 CSoutput.n222 CSoutput.n215 4.5005
R1250 CSoutput.n222 CSoutput.n210 4.5005
R1251 CSoutput.n222 CSoutput.t184 4.5005
R1252 CSoutput.n222 CSoutput.n209 4.5005
R1253 CSoutput.n222 CSoutput.n216 4.5005
R1254 CSoutput.n265 CSoutput.n222 4.5005
R1255 CSoutput.n246 CSoutput.n212 4.5005
R1256 CSoutput.n246 CSoutput.n214 4.5005
R1257 CSoutput.n246 CSoutput.n211 4.5005
R1258 CSoutput.n246 CSoutput.n215 4.5005
R1259 CSoutput.n246 CSoutput.n210 4.5005
R1260 CSoutput.n246 CSoutput.t184 4.5005
R1261 CSoutput.n246 CSoutput.n209 4.5005
R1262 CSoutput.n246 CSoutput.n216 4.5005
R1263 CSoutput.n265 CSoutput.n246 4.5005
R1264 CSoutput.n212 CSoutput.n207 4.5005
R1265 CSoutput.n214 CSoutput.n207 4.5005
R1266 CSoutput.n211 CSoutput.n207 4.5005
R1267 CSoutput.n215 CSoutput.n207 4.5005
R1268 CSoutput.n210 CSoutput.n207 4.5005
R1269 CSoutput.t184 CSoutput.n207 4.5005
R1270 CSoutput.n209 CSoutput.n207 4.5005
R1271 CSoutput.n216 CSoutput.n207 4.5005
R1272 CSoutput.n268 CSoutput.n212 4.5005
R1273 CSoutput.n268 CSoutput.n214 4.5005
R1274 CSoutput.n268 CSoutput.n211 4.5005
R1275 CSoutput.n268 CSoutput.n215 4.5005
R1276 CSoutput.n268 CSoutput.n210 4.5005
R1277 CSoutput.n268 CSoutput.t184 4.5005
R1278 CSoutput.n268 CSoutput.n209 4.5005
R1279 CSoutput.n268 CSoutput.n216 4.5005
R1280 CSoutput.n266 CSoutput.n212 4.5005
R1281 CSoutput.n266 CSoutput.n214 4.5005
R1282 CSoutput.n266 CSoutput.n211 4.5005
R1283 CSoutput.n266 CSoutput.n215 4.5005
R1284 CSoutput.n266 CSoutput.n210 4.5005
R1285 CSoutput.n266 CSoutput.t184 4.5005
R1286 CSoutput.n266 CSoutput.n209 4.5005
R1287 CSoutput.n266 CSoutput.n216 4.5005
R1288 CSoutput.n266 CSoutput.n265 4.5005
R1289 CSoutput.n248 CSoutput.n212 4.5005
R1290 CSoutput.n248 CSoutput.n214 4.5005
R1291 CSoutput.n248 CSoutput.n211 4.5005
R1292 CSoutput.n248 CSoutput.n215 4.5005
R1293 CSoutput.n248 CSoutput.n210 4.5005
R1294 CSoutput.n248 CSoutput.t184 4.5005
R1295 CSoutput.n248 CSoutput.n209 4.5005
R1296 CSoutput.n248 CSoutput.n216 4.5005
R1297 CSoutput.n265 CSoutput.n248 4.5005
R1298 CSoutput.n220 CSoutput.n212 4.5005
R1299 CSoutput.n220 CSoutput.n214 4.5005
R1300 CSoutput.n220 CSoutput.n211 4.5005
R1301 CSoutput.n220 CSoutput.n215 4.5005
R1302 CSoutput.n220 CSoutput.n210 4.5005
R1303 CSoutput.n220 CSoutput.t184 4.5005
R1304 CSoutput.n220 CSoutput.n209 4.5005
R1305 CSoutput.n220 CSoutput.n216 4.5005
R1306 CSoutput.n265 CSoutput.n220 4.5005
R1307 CSoutput.n250 CSoutput.n212 4.5005
R1308 CSoutput.n250 CSoutput.n214 4.5005
R1309 CSoutput.n250 CSoutput.n211 4.5005
R1310 CSoutput.n250 CSoutput.n215 4.5005
R1311 CSoutput.n250 CSoutput.n210 4.5005
R1312 CSoutput.n250 CSoutput.t184 4.5005
R1313 CSoutput.n250 CSoutput.n209 4.5005
R1314 CSoutput.n250 CSoutput.n216 4.5005
R1315 CSoutput.n265 CSoutput.n250 4.5005
R1316 CSoutput.n219 CSoutput.n212 4.5005
R1317 CSoutput.n219 CSoutput.n214 4.5005
R1318 CSoutput.n219 CSoutput.n211 4.5005
R1319 CSoutput.n219 CSoutput.n215 4.5005
R1320 CSoutput.n219 CSoutput.n210 4.5005
R1321 CSoutput.n219 CSoutput.t184 4.5005
R1322 CSoutput.n219 CSoutput.n209 4.5005
R1323 CSoutput.n219 CSoutput.n216 4.5005
R1324 CSoutput.n265 CSoutput.n219 4.5005
R1325 CSoutput.n264 CSoutput.n212 4.5005
R1326 CSoutput.n264 CSoutput.n214 4.5005
R1327 CSoutput.n264 CSoutput.n211 4.5005
R1328 CSoutput.n264 CSoutput.n215 4.5005
R1329 CSoutput.n264 CSoutput.n210 4.5005
R1330 CSoutput.n264 CSoutput.t184 4.5005
R1331 CSoutput.n264 CSoutput.n209 4.5005
R1332 CSoutput.n264 CSoutput.n216 4.5005
R1333 CSoutput.n265 CSoutput.n264 4.5005
R1334 CSoutput.n263 CSoutput.n148 4.5005
R1335 CSoutput.n164 CSoutput.n148 4.5005
R1336 CSoutput.n159 CSoutput.n143 4.5005
R1337 CSoutput.n159 CSoutput.n145 4.5005
R1338 CSoutput.n159 CSoutput.n142 4.5005
R1339 CSoutput.n159 CSoutput.n146 4.5005
R1340 CSoutput.n159 CSoutput.n141 4.5005
R1341 CSoutput.n159 CSoutput.t193 4.5005
R1342 CSoutput.n159 CSoutput.n140 4.5005
R1343 CSoutput.n159 CSoutput.n147 4.5005
R1344 CSoutput.n159 CSoutput.n148 4.5005
R1345 CSoutput.n157 CSoutput.n143 4.5005
R1346 CSoutput.n157 CSoutput.n145 4.5005
R1347 CSoutput.n157 CSoutput.n142 4.5005
R1348 CSoutput.n157 CSoutput.n146 4.5005
R1349 CSoutput.n157 CSoutput.n141 4.5005
R1350 CSoutput.n157 CSoutput.t193 4.5005
R1351 CSoutput.n157 CSoutput.n140 4.5005
R1352 CSoutput.n157 CSoutput.n147 4.5005
R1353 CSoutput.n157 CSoutput.n148 4.5005
R1354 CSoutput.n156 CSoutput.n143 4.5005
R1355 CSoutput.n156 CSoutput.n145 4.5005
R1356 CSoutput.n156 CSoutput.n142 4.5005
R1357 CSoutput.n156 CSoutput.n146 4.5005
R1358 CSoutput.n156 CSoutput.n141 4.5005
R1359 CSoutput.n156 CSoutput.t193 4.5005
R1360 CSoutput.n156 CSoutput.n140 4.5005
R1361 CSoutput.n156 CSoutput.n147 4.5005
R1362 CSoutput.n156 CSoutput.n148 4.5005
R1363 CSoutput.n285 CSoutput.n143 4.5005
R1364 CSoutput.n285 CSoutput.n145 4.5005
R1365 CSoutput.n285 CSoutput.n142 4.5005
R1366 CSoutput.n285 CSoutput.n146 4.5005
R1367 CSoutput.n285 CSoutput.n141 4.5005
R1368 CSoutput.n285 CSoutput.t193 4.5005
R1369 CSoutput.n285 CSoutput.n140 4.5005
R1370 CSoutput.n285 CSoutput.n147 4.5005
R1371 CSoutput.n285 CSoutput.n148 4.5005
R1372 CSoutput.n283 CSoutput.n143 4.5005
R1373 CSoutput.n283 CSoutput.n145 4.5005
R1374 CSoutput.n283 CSoutput.n142 4.5005
R1375 CSoutput.n283 CSoutput.n146 4.5005
R1376 CSoutput.n283 CSoutput.n141 4.5005
R1377 CSoutput.n283 CSoutput.t193 4.5005
R1378 CSoutput.n283 CSoutput.n140 4.5005
R1379 CSoutput.n283 CSoutput.n147 4.5005
R1380 CSoutput.n281 CSoutput.n143 4.5005
R1381 CSoutput.n281 CSoutput.n145 4.5005
R1382 CSoutput.n281 CSoutput.n142 4.5005
R1383 CSoutput.n281 CSoutput.n146 4.5005
R1384 CSoutput.n281 CSoutput.n141 4.5005
R1385 CSoutput.n281 CSoutput.t193 4.5005
R1386 CSoutput.n281 CSoutput.n140 4.5005
R1387 CSoutput.n281 CSoutput.n147 4.5005
R1388 CSoutput.n167 CSoutput.n143 4.5005
R1389 CSoutput.n167 CSoutput.n145 4.5005
R1390 CSoutput.n167 CSoutput.n142 4.5005
R1391 CSoutput.n167 CSoutput.n146 4.5005
R1392 CSoutput.n167 CSoutput.n141 4.5005
R1393 CSoutput.n167 CSoutput.t193 4.5005
R1394 CSoutput.n167 CSoutput.n140 4.5005
R1395 CSoutput.n167 CSoutput.n147 4.5005
R1396 CSoutput.n167 CSoutput.n148 4.5005
R1397 CSoutput.n166 CSoutput.n143 4.5005
R1398 CSoutput.n166 CSoutput.n145 4.5005
R1399 CSoutput.n166 CSoutput.n142 4.5005
R1400 CSoutput.n166 CSoutput.n146 4.5005
R1401 CSoutput.n166 CSoutput.n141 4.5005
R1402 CSoutput.n166 CSoutput.t193 4.5005
R1403 CSoutput.n166 CSoutput.n140 4.5005
R1404 CSoutput.n166 CSoutput.n147 4.5005
R1405 CSoutput.n166 CSoutput.n148 4.5005
R1406 CSoutput.n170 CSoutput.n143 4.5005
R1407 CSoutput.n170 CSoutput.n145 4.5005
R1408 CSoutput.n170 CSoutput.n142 4.5005
R1409 CSoutput.n170 CSoutput.n146 4.5005
R1410 CSoutput.n170 CSoutput.n141 4.5005
R1411 CSoutput.n170 CSoutput.t193 4.5005
R1412 CSoutput.n170 CSoutput.n140 4.5005
R1413 CSoutput.n170 CSoutput.n147 4.5005
R1414 CSoutput.n170 CSoutput.n148 4.5005
R1415 CSoutput.n169 CSoutput.n143 4.5005
R1416 CSoutput.n169 CSoutput.n145 4.5005
R1417 CSoutput.n169 CSoutput.n142 4.5005
R1418 CSoutput.n169 CSoutput.n146 4.5005
R1419 CSoutput.n169 CSoutput.n141 4.5005
R1420 CSoutput.n169 CSoutput.t193 4.5005
R1421 CSoutput.n169 CSoutput.n140 4.5005
R1422 CSoutput.n169 CSoutput.n147 4.5005
R1423 CSoutput.n169 CSoutput.n148 4.5005
R1424 CSoutput.n152 CSoutput.n143 4.5005
R1425 CSoutput.n152 CSoutput.n145 4.5005
R1426 CSoutput.n152 CSoutput.n142 4.5005
R1427 CSoutput.n152 CSoutput.n146 4.5005
R1428 CSoutput.n152 CSoutput.n141 4.5005
R1429 CSoutput.n152 CSoutput.t193 4.5005
R1430 CSoutput.n152 CSoutput.n140 4.5005
R1431 CSoutput.n152 CSoutput.n147 4.5005
R1432 CSoutput.n152 CSoutput.n148 4.5005
R1433 CSoutput.n288 CSoutput.n143 4.5005
R1434 CSoutput.n288 CSoutput.n145 4.5005
R1435 CSoutput.n288 CSoutput.n142 4.5005
R1436 CSoutput.n288 CSoutput.n146 4.5005
R1437 CSoutput.n288 CSoutput.n141 4.5005
R1438 CSoutput.n288 CSoutput.t193 4.5005
R1439 CSoutput.n288 CSoutput.n140 4.5005
R1440 CSoutput.n288 CSoutput.n147 4.5005
R1441 CSoutput.n288 CSoutput.n148 4.5005
R1442 CSoutput.n347 CSoutput.n327 4.10845
R1443 CSoutput.n137 CSoutput.n117 4.10845
R1444 CSoutput.n345 CSoutput.t84 4.06363
R1445 CSoutput.n345 CSoutput.t14 4.06363
R1446 CSoutput.n343 CSoutput.t73 4.06363
R1447 CSoutput.n343 CSoutput.t96 4.06363
R1448 CSoutput.n341 CSoutput.t28 4.06363
R1449 CSoutput.n341 CSoutput.t58 4.06363
R1450 CSoutput.n339 CSoutput.t67 4.06363
R1451 CSoutput.n339 CSoutput.t60 4.06363
R1452 CSoutput.n337 CSoutput.t86 4.06363
R1453 CSoutput.n337 CSoutput.t52 4.06363
R1454 CSoutput.n335 CSoutput.t32 4.06363
R1455 CSoutput.n335 CSoutput.t43 4.06363
R1456 CSoutput.n333 CSoutput.t57 4.06363
R1457 CSoutput.n333 CSoutput.t29 4.06363
R1458 CSoutput.n331 CSoutput.t39 4.06363
R1459 CSoutput.n331 CSoutput.t65 4.06363
R1460 CSoutput.n329 CSoutput.t10 4.06363
R1461 CSoutput.n329 CSoutput.t11 4.06363
R1462 CSoutput.n328 CSoutput.t44 4.06363
R1463 CSoutput.n328 CSoutput.t94 4.06363
R1464 CSoutput.n325 CSoutput.t63 4.06363
R1465 CSoutput.n325 CSoutput.t3 4.06363
R1466 CSoutput.n323 CSoutput.t85 4.06363
R1467 CSoutput.n323 CSoutput.t21 4.06363
R1468 CSoutput.n321 CSoutput.t46 4.06363
R1469 CSoutput.n321 CSoutput.t181 4.06363
R1470 CSoutput.n319 CSoutput.t183 4.06363
R1471 CSoutput.n319 CSoutput.t179 4.06363
R1472 CSoutput.n317 CSoutput.t167 4.06363
R1473 CSoutput.n317 CSoutput.t2 4.06363
R1474 CSoutput.n315 CSoutput.t66 4.06363
R1475 CSoutput.n315 CSoutput.t16 4.06363
R1476 CSoutput.n313 CSoutput.t0 4.06363
R1477 CSoutput.n313 CSoutput.t176 4.06363
R1478 CSoutput.n311 CSoutput.t88 4.06363
R1479 CSoutput.n311 CSoutput.t42 4.06363
R1480 CSoutput.n309 CSoutput.t165 4.06363
R1481 CSoutput.n309 CSoutput.t54 4.06363
R1482 CSoutput.n308 CSoutput.t64 4.06363
R1483 CSoutput.n308 CSoutput.t53 4.06363
R1484 CSoutput.n306 CSoutput.t17 4.06363
R1485 CSoutput.n306 CSoutput.t80 4.06363
R1486 CSoutput.n304 CSoutput.t79 4.06363
R1487 CSoutput.n304 CSoutput.t8 4.06363
R1488 CSoutput.n302 CSoutput.t20 4.06363
R1489 CSoutput.n302 CSoutput.t49 4.06363
R1490 CSoutput.n300 CSoutput.t82 4.06363
R1491 CSoutput.n300 CSoutput.t61 4.06363
R1492 CSoutput.n298 CSoutput.t76 4.06363
R1493 CSoutput.n298 CSoutput.t172 4.06363
R1494 CSoutput.n296 CSoutput.t35 4.06363
R1495 CSoutput.n296 CSoutput.t173 4.06363
R1496 CSoutput.n294 CSoutput.t40 4.06363
R1497 CSoutput.n294 CSoutput.t75 4.06363
R1498 CSoutput.n292 CSoutput.t89 4.06363
R1499 CSoutput.n292 CSoutput.t51 4.06363
R1500 CSoutput.n290 CSoutput.t45 4.06363
R1501 CSoutput.n290 CSoutput.t23 4.06363
R1502 CSoutput.n289 CSoutput.t180 4.06363
R1503 CSoutput.n289 CSoutput.t33 4.06363
R1504 CSoutput.n118 CSoutput.t55 4.06363
R1505 CSoutput.n118 CSoutput.t1 4.06363
R1506 CSoutput.n119 CSoutput.t78 4.06363
R1507 CSoutput.n119 CSoutput.t38 4.06363
R1508 CSoutput.n121 CSoutput.t91 4.06363
R1509 CSoutput.n121 CSoutput.t175 4.06363
R1510 CSoutput.n123 CSoutput.t47 4.06363
R1511 CSoutput.n123 CSoutput.t30 4.06363
R1512 CSoutput.n125 CSoutput.t169 4.06363
R1513 CSoutput.n125 CSoutput.t4 4.06363
R1514 CSoutput.n127 CSoutput.t24 4.06363
R1515 CSoutput.n127 CSoutput.t48 4.06363
R1516 CSoutput.n129 CSoutput.t68 4.06363
R1517 CSoutput.n129 CSoutput.t19 4.06363
R1518 CSoutput.n131 CSoutput.t171 4.06363
R1519 CSoutput.n131 CSoutput.t12 4.06363
R1520 CSoutput.n133 CSoutput.t36 4.06363
R1521 CSoutput.n133 CSoutput.t97 4.06363
R1522 CSoutput.n135 CSoutput.t162 4.06363
R1523 CSoutput.n135 CSoutput.t177 4.06363
R1524 CSoutput.n98 CSoutput.t182 4.06363
R1525 CSoutput.n98 CSoutput.t56 4.06363
R1526 CSoutput.n99 CSoutput.t72 4.06363
R1527 CSoutput.n99 CSoutput.t178 4.06363
R1528 CSoutput.n101 CSoutput.t71 4.06363
R1529 CSoutput.n101 CSoutput.t170 4.06363
R1530 CSoutput.n103 CSoutput.t9 4.06363
R1531 CSoutput.n103 CSoutput.t74 4.06363
R1532 CSoutput.n105 CSoutput.t83 4.06363
R1533 CSoutput.n105 CSoutput.t93 4.06363
R1534 CSoutput.n107 CSoutput.t87 4.06363
R1535 CSoutput.n107 CSoutput.t62 4.06363
R1536 CSoutput.n109 CSoutput.t166 4.06363
R1537 CSoutput.n109 CSoutput.t77 4.06363
R1538 CSoutput.n111 CSoutput.t92 4.06363
R1539 CSoutput.n111 CSoutput.t26 4.06363
R1540 CSoutput.n113 CSoutput.t163 4.06363
R1541 CSoutput.n113 CSoutput.t70 4.06363
R1542 CSoutput.n115 CSoutput.t15 4.06363
R1543 CSoutput.n115 CSoutput.t31 4.06363
R1544 CSoutput.n79 CSoutput.t25 4.06363
R1545 CSoutput.n79 CSoutput.t81 4.06363
R1546 CSoutput.n80 CSoutput.t90 4.06363
R1547 CSoutput.n80 CSoutput.t50 4.06363
R1548 CSoutput.n82 CSoutput.t168 4.06363
R1549 CSoutput.n82 CSoutput.t5 4.06363
R1550 CSoutput.n84 CSoutput.t18 4.06363
R1551 CSoutput.n84 CSoutput.t164 4.06363
R1552 CSoutput.n86 CSoutput.t174 4.06363
R1553 CSoutput.n86 CSoutput.t7 4.06363
R1554 CSoutput.n88 CSoutput.t59 4.06363
R1555 CSoutput.n88 CSoutput.t13 4.06363
R1556 CSoutput.n90 CSoutput.t6 4.06363
R1557 CSoutput.n90 CSoutput.t34 4.06363
R1558 CSoutput.n92 CSoutput.t95 4.06363
R1559 CSoutput.n92 CSoutput.t27 4.06363
R1560 CSoutput.n94 CSoutput.t69 4.06363
R1561 CSoutput.n94 CSoutput.t41 4.06363
R1562 CSoutput.n96 CSoutput.t37 4.06363
R1563 CSoutput.n96 CSoutput.t22 4.06363
R1564 CSoutput.n44 CSoutput.n43 3.79402
R1565 CSoutput.n49 CSoutput.n48 3.79402
R1566 CSoutput.n413 CSoutput.n412 3.57343
R1567 CSoutput.n412 CSoutput.n380 3.08965
R1568 CSoutput.n377 CSoutput.t99 2.82907
R1569 CSoutput.n377 CSoutput.t103 2.82907
R1570 CSoutput.n375 CSoutput.t116 2.82907
R1571 CSoutput.n375 CSoutput.t146 2.82907
R1572 CSoutput.n373 CSoutput.t106 2.82907
R1573 CSoutput.n373 CSoutput.t109 2.82907
R1574 CSoutput.n371 CSoutput.t104 2.82907
R1575 CSoutput.n371 CSoutput.t123 2.82907
R1576 CSoutput.n369 CSoutput.t143 2.82907
R1577 CSoutput.n369 CSoutput.t119 2.82907
R1578 CSoutput.n367 CSoutput.t126 2.82907
R1579 CSoutput.n367 CSoutput.t133 2.82907
R1580 CSoutput.n365 CSoutput.t101 2.82907
R1581 CSoutput.n365 CSoutput.t112 2.82907
R1582 CSoutput.n364 CSoutput.t118 2.82907
R1583 CSoutput.n364 CSoutput.t148 2.82907
R1584 CSoutput.n362 CSoutput.t105 2.82907
R1585 CSoutput.n362 CSoutput.t124 2.82907
R1586 CSoutput.n360 CSoutput.t147 2.82907
R1587 CSoutput.n360 CSoutput.t160 2.82907
R1588 CSoutput.n358 CSoutput.t127 2.82907
R1589 CSoutput.n358 CSoutput.t117 2.82907
R1590 CSoutput.n356 CSoutput.t125 2.82907
R1591 CSoutput.n356 CSoutput.t132 2.82907
R1592 CSoutput.n354 CSoutput.t100 2.82907
R1593 CSoutput.n354 CSoutput.t152 2.82907
R1594 CSoutput.n352 CSoutput.t135 2.82907
R1595 CSoutput.n352 CSoutput.t141 2.82907
R1596 CSoutput.n350 CSoutput.t108 2.82907
R1597 CSoutput.n350 CSoutput.t110 2.82907
R1598 CSoutput.n349 CSoutput.t151 2.82907
R1599 CSoutput.n349 CSoutput.t129 2.82907
R1600 CSoutput.n396 CSoutput.t156 2.82907
R1601 CSoutput.n396 CSoutput.t144 2.82907
R1602 CSoutput.n397 CSoutput.t107 2.82907
R1603 CSoutput.n397 CSoutput.t142 2.82907
R1604 CSoutput.n399 CSoutput.t139 2.82907
R1605 CSoutput.n399 CSoutput.t157 2.82907
R1606 CSoutput.n401 CSoutput.t145 2.82907
R1607 CSoutput.n401 CSoutput.t153 2.82907
R1608 CSoutput.n403 CSoutput.t161 2.82907
R1609 CSoutput.n403 CSoutput.t121 2.82907
R1610 CSoutput.n405 CSoutput.t128 2.82907
R1611 CSoutput.n405 CSoutput.t111 2.82907
R1612 CSoutput.n407 CSoutput.t154 2.82907
R1613 CSoutput.n407 CSoutput.t134 2.82907
R1614 CSoutput.n409 CSoutput.t150 2.82907
R1615 CSoutput.n409 CSoutput.t149 2.82907
R1616 CSoutput.n381 CSoutput.t137 2.82907
R1617 CSoutput.n381 CSoutput.t158 2.82907
R1618 CSoutput.n382 CSoutput.t115 2.82907
R1619 CSoutput.n382 CSoutput.t98 2.82907
R1620 CSoutput.n384 CSoutput.t102 2.82907
R1621 CSoutput.n384 CSoutput.t140 2.82907
R1622 CSoutput.n386 CSoutput.t159 2.82907
R1623 CSoutput.n386 CSoutput.t113 2.82907
R1624 CSoutput.n388 CSoutput.t138 2.82907
R1625 CSoutput.n388 CSoutput.t131 2.82907
R1626 CSoutput.n390 CSoutput.t136 2.82907
R1627 CSoutput.n390 CSoutput.t120 2.82907
R1628 CSoutput.n392 CSoutput.t114 2.82907
R1629 CSoutput.n392 CSoutput.t155 2.82907
R1630 CSoutput.n394 CSoutput.t130 2.82907
R1631 CSoutput.n394 CSoutput.t122 2.82907
R1632 CSoutput.n348 CSoutput.n138 2.57547
R1633 CSoutput.n75 CSoutput.n1 2.45513
R1634 CSoutput.n229 CSoutput.n227 2.251
R1635 CSoutput.n229 CSoutput.n226 2.251
R1636 CSoutput.n229 CSoutput.n225 2.251
R1637 CSoutput.n229 CSoutput.n224 2.251
R1638 CSoutput.n198 CSoutput.n197 2.251
R1639 CSoutput.n198 CSoutput.n196 2.251
R1640 CSoutput.n198 CSoutput.n195 2.251
R1641 CSoutput.n198 CSoutput.n194 2.251
R1642 CSoutput.n271 CSoutput.n270 2.251
R1643 CSoutput.n236 CSoutput.n234 2.251
R1644 CSoutput.n236 CSoutput.n233 2.251
R1645 CSoutput.n236 CSoutput.n232 2.251
R1646 CSoutput.n254 CSoutput.n236 2.251
R1647 CSoutput.n242 CSoutput.n241 2.251
R1648 CSoutput.n242 CSoutput.n240 2.251
R1649 CSoutput.n242 CSoutput.n239 2.251
R1650 CSoutput.n242 CSoutput.n238 2.251
R1651 CSoutput.n268 CSoutput.n208 2.251
R1652 CSoutput.n263 CSoutput.n261 2.251
R1653 CSoutput.n263 CSoutput.n260 2.251
R1654 CSoutput.n263 CSoutput.n259 2.251
R1655 CSoutput.n263 CSoutput.n258 2.251
R1656 CSoutput.n164 CSoutput.n163 2.251
R1657 CSoutput.n164 CSoutput.n162 2.251
R1658 CSoutput.n164 CSoutput.n161 2.251
R1659 CSoutput.n164 CSoutput.n160 2.251
R1660 CSoutput.n281 CSoutput.n280 2.251
R1661 CSoutput.n198 CSoutput.n178 2.2505
R1662 CSoutput.n193 CSoutput.n178 2.2505
R1663 CSoutput.n191 CSoutput.n178 2.2505
R1664 CSoutput.n190 CSoutput.n178 2.2505
R1665 CSoutput.n275 CSoutput.n178 2.2505
R1666 CSoutput.n273 CSoutput.n178 2.2505
R1667 CSoutput.n271 CSoutput.n178 2.2505
R1668 CSoutput.n201 CSoutput.n178 2.2505
R1669 CSoutput.n200 CSoutput.n178 2.2505
R1670 CSoutput.n204 CSoutput.n178 2.2505
R1671 CSoutput.n203 CSoutput.n178 2.2505
R1672 CSoutput.n186 CSoutput.n178 2.2505
R1673 CSoutput.n278 CSoutput.n178 2.2505
R1674 CSoutput.n278 CSoutput.n277 2.2505
R1675 CSoutput.n242 CSoutput.n213 2.2505
R1676 CSoutput.n223 CSoutput.n213 2.2505
R1677 CSoutput.n244 CSoutput.n213 2.2505
R1678 CSoutput.n222 CSoutput.n213 2.2505
R1679 CSoutput.n246 CSoutput.n213 2.2505
R1680 CSoutput.n213 CSoutput.n207 2.2505
R1681 CSoutput.n268 CSoutput.n213 2.2505
R1682 CSoutput.n266 CSoutput.n213 2.2505
R1683 CSoutput.n248 CSoutput.n213 2.2505
R1684 CSoutput.n220 CSoutput.n213 2.2505
R1685 CSoutput.n250 CSoutput.n213 2.2505
R1686 CSoutput.n219 CSoutput.n213 2.2505
R1687 CSoutput.n264 CSoutput.n213 2.2505
R1688 CSoutput.n264 CSoutput.n217 2.2505
R1689 CSoutput.n164 CSoutput.n144 2.2505
R1690 CSoutput.n159 CSoutput.n144 2.2505
R1691 CSoutput.n157 CSoutput.n144 2.2505
R1692 CSoutput.n156 CSoutput.n144 2.2505
R1693 CSoutput.n285 CSoutput.n144 2.2505
R1694 CSoutput.n283 CSoutput.n144 2.2505
R1695 CSoutput.n281 CSoutput.n144 2.2505
R1696 CSoutput.n167 CSoutput.n144 2.2505
R1697 CSoutput.n166 CSoutput.n144 2.2505
R1698 CSoutput.n170 CSoutput.n144 2.2505
R1699 CSoutput.n169 CSoutput.n144 2.2505
R1700 CSoutput.n152 CSoutput.n144 2.2505
R1701 CSoutput.n288 CSoutput.n144 2.2505
R1702 CSoutput.n288 CSoutput.n287 2.2505
R1703 CSoutput.n206 CSoutput.n199 2.25024
R1704 CSoutput.n206 CSoutput.n192 2.25024
R1705 CSoutput.n274 CSoutput.n206 2.25024
R1706 CSoutput.n206 CSoutput.n202 2.25024
R1707 CSoutput.n206 CSoutput.n205 2.25024
R1708 CSoutput.n206 CSoutput.n173 2.25024
R1709 CSoutput.n256 CSoutput.n253 2.25024
R1710 CSoutput.n256 CSoutput.n252 2.25024
R1711 CSoutput.n256 CSoutput.n251 2.25024
R1712 CSoutput.n256 CSoutput.n218 2.25024
R1713 CSoutput.n256 CSoutput.n255 2.25024
R1714 CSoutput.n257 CSoutput.n256 2.25024
R1715 CSoutput.n172 CSoutput.n165 2.25024
R1716 CSoutput.n172 CSoutput.n158 2.25024
R1717 CSoutput.n284 CSoutput.n172 2.25024
R1718 CSoutput.n172 CSoutput.n168 2.25024
R1719 CSoutput.n172 CSoutput.n171 2.25024
R1720 CSoutput.n172 CSoutput.n139 2.25024
R1721 CSoutput.n273 CSoutput.n183 1.50111
R1722 CSoutput.n221 CSoutput.n207 1.50111
R1723 CSoutput.n283 CSoutput.n149 1.50111
R1724 CSoutput.n229 CSoutput.n228 1.501
R1725 CSoutput.n236 CSoutput.n235 1.501
R1726 CSoutput.n263 CSoutput.n262 1.501
R1727 CSoutput.n277 CSoutput.n188 1.12536
R1728 CSoutput.n277 CSoutput.n189 1.12536
R1729 CSoutput.n277 CSoutput.n276 1.12536
R1730 CSoutput.n237 CSoutput.n217 1.12536
R1731 CSoutput.n243 CSoutput.n217 1.12536
R1732 CSoutput.n245 CSoutput.n217 1.12536
R1733 CSoutput.n287 CSoutput.n154 1.12536
R1734 CSoutput.n287 CSoutput.n155 1.12536
R1735 CSoutput.n287 CSoutput.n286 1.12536
R1736 CSoutput.n277 CSoutput.n184 1.12536
R1737 CSoutput.n277 CSoutput.n185 1.12536
R1738 CSoutput.n277 CSoutput.n187 1.12536
R1739 CSoutput.n267 CSoutput.n217 1.12536
R1740 CSoutput.n247 CSoutput.n217 1.12536
R1741 CSoutput.n249 CSoutput.n217 1.12536
R1742 CSoutput.n287 CSoutput.n150 1.12536
R1743 CSoutput.n287 CSoutput.n151 1.12536
R1744 CSoutput.n287 CSoutput.n153 1.12536
R1745 CSoutput.n31 CSoutput.n30 0.669944
R1746 CSoutput.n62 CSoutput.n61 0.669944
R1747 CSoutput.n368 CSoutput.n366 0.573776
R1748 CSoutput.n370 CSoutput.n368 0.573776
R1749 CSoutput.n372 CSoutput.n370 0.573776
R1750 CSoutput.n374 CSoutput.n372 0.573776
R1751 CSoutput.n376 CSoutput.n374 0.573776
R1752 CSoutput.n378 CSoutput.n376 0.573776
R1753 CSoutput.n353 CSoutput.n351 0.573776
R1754 CSoutput.n355 CSoutput.n353 0.573776
R1755 CSoutput.n357 CSoutput.n355 0.573776
R1756 CSoutput.n359 CSoutput.n357 0.573776
R1757 CSoutput.n361 CSoutput.n359 0.573776
R1758 CSoutput.n363 CSoutput.n361 0.573776
R1759 CSoutput.n410 CSoutput.n408 0.573776
R1760 CSoutput.n408 CSoutput.n406 0.573776
R1761 CSoutput.n406 CSoutput.n404 0.573776
R1762 CSoutput.n404 CSoutput.n402 0.573776
R1763 CSoutput.n402 CSoutput.n400 0.573776
R1764 CSoutput.n400 CSoutput.n398 0.573776
R1765 CSoutput.n395 CSoutput.n393 0.573776
R1766 CSoutput.n393 CSoutput.n391 0.573776
R1767 CSoutput.n391 CSoutput.n389 0.573776
R1768 CSoutput.n389 CSoutput.n387 0.573776
R1769 CSoutput.n387 CSoutput.n385 0.573776
R1770 CSoutput.n385 CSoutput.n383 0.573776
R1771 CSoutput.n413 CSoutput.n288 0.53442
R1772 CSoutput.n332 CSoutput.n330 0.358259
R1773 CSoutput.n334 CSoutput.n332 0.358259
R1774 CSoutput.n336 CSoutput.n334 0.358259
R1775 CSoutput.n338 CSoutput.n336 0.358259
R1776 CSoutput.n340 CSoutput.n338 0.358259
R1777 CSoutput.n342 CSoutput.n340 0.358259
R1778 CSoutput.n344 CSoutput.n342 0.358259
R1779 CSoutput.n346 CSoutput.n344 0.358259
R1780 CSoutput.n312 CSoutput.n310 0.358259
R1781 CSoutput.n314 CSoutput.n312 0.358259
R1782 CSoutput.n316 CSoutput.n314 0.358259
R1783 CSoutput.n318 CSoutput.n316 0.358259
R1784 CSoutput.n320 CSoutput.n318 0.358259
R1785 CSoutput.n322 CSoutput.n320 0.358259
R1786 CSoutput.n324 CSoutput.n322 0.358259
R1787 CSoutput.n326 CSoutput.n324 0.358259
R1788 CSoutput.n293 CSoutput.n291 0.358259
R1789 CSoutput.n295 CSoutput.n293 0.358259
R1790 CSoutput.n297 CSoutput.n295 0.358259
R1791 CSoutput.n299 CSoutput.n297 0.358259
R1792 CSoutput.n301 CSoutput.n299 0.358259
R1793 CSoutput.n303 CSoutput.n301 0.358259
R1794 CSoutput.n305 CSoutput.n303 0.358259
R1795 CSoutput.n307 CSoutput.n305 0.358259
R1796 CSoutput.n136 CSoutput.n134 0.358259
R1797 CSoutput.n134 CSoutput.n132 0.358259
R1798 CSoutput.n132 CSoutput.n130 0.358259
R1799 CSoutput.n130 CSoutput.n128 0.358259
R1800 CSoutput.n128 CSoutput.n126 0.358259
R1801 CSoutput.n126 CSoutput.n124 0.358259
R1802 CSoutput.n124 CSoutput.n122 0.358259
R1803 CSoutput.n122 CSoutput.n120 0.358259
R1804 CSoutput.n116 CSoutput.n114 0.358259
R1805 CSoutput.n114 CSoutput.n112 0.358259
R1806 CSoutput.n112 CSoutput.n110 0.358259
R1807 CSoutput.n110 CSoutput.n108 0.358259
R1808 CSoutput.n108 CSoutput.n106 0.358259
R1809 CSoutput.n106 CSoutput.n104 0.358259
R1810 CSoutput.n104 CSoutput.n102 0.358259
R1811 CSoutput.n102 CSoutput.n100 0.358259
R1812 CSoutput.n97 CSoutput.n95 0.358259
R1813 CSoutput.n95 CSoutput.n93 0.358259
R1814 CSoutput.n93 CSoutput.n91 0.358259
R1815 CSoutput.n91 CSoutput.n89 0.358259
R1816 CSoutput.n89 CSoutput.n87 0.358259
R1817 CSoutput.n87 CSoutput.n85 0.358259
R1818 CSoutput.n85 CSoutput.n83 0.358259
R1819 CSoutput.n83 CSoutput.n81 0.358259
R1820 CSoutput.n21 CSoutput.n20 0.169105
R1821 CSoutput.n21 CSoutput.n16 0.169105
R1822 CSoutput.n26 CSoutput.n16 0.169105
R1823 CSoutput.n27 CSoutput.n26 0.169105
R1824 CSoutput.n27 CSoutput.n14 0.169105
R1825 CSoutput.n32 CSoutput.n14 0.169105
R1826 CSoutput.n33 CSoutput.n32 0.169105
R1827 CSoutput.n34 CSoutput.n33 0.169105
R1828 CSoutput.n34 CSoutput.n12 0.169105
R1829 CSoutput.n39 CSoutput.n12 0.169105
R1830 CSoutput.n40 CSoutput.n39 0.169105
R1831 CSoutput.n40 CSoutput.n10 0.169105
R1832 CSoutput.n45 CSoutput.n10 0.169105
R1833 CSoutput.n46 CSoutput.n45 0.169105
R1834 CSoutput.n47 CSoutput.n46 0.169105
R1835 CSoutput.n47 CSoutput.n8 0.169105
R1836 CSoutput.n52 CSoutput.n8 0.169105
R1837 CSoutput.n53 CSoutput.n52 0.169105
R1838 CSoutput.n53 CSoutput.n6 0.169105
R1839 CSoutput.n58 CSoutput.n6 0.169105
R1840 CSoutput.n59 CSoutput.n58 0.169105
R1841 CSoutput.n60 CSoutput.n59 0.169105
R1842 CSoutput.n60 CSoutput.n4 0.169105
R1843 CSoutput.n66 CSoutput.n4 0.169105
R1844 CSoutput.n67 CSoutput.n66 0.169105
R1845 CSoutput.n68 CSoutput.n67 0.169105
R1846 CSoutput.n68 CSoutput.n2 0.169105
R1847 CSoutput.n73 CSoutput.n2 0.169105
R1848 CSoutput.n74 CSoutput.n73 0.169105
R1849 CSoutput.n74 CSoutput.n0 0.169105
R1850 CSoutput.n78 CSoutput.n0 0.169105
R1851 CSoutput.n231 CSoutput.n230 0.0910737
R1852 CSoutput.n282 CSoutput.n279 0.0723685
R1853 CSoutput.n236 CSoutput.n231 0.0522944
R1854 CSoutput.n279 CSoutput.n278 0.0499135
R1855 CSoutput.n230 CSoutput.n229 0.0499135
R1856 CSoutput.n264 CSoutput.n263 0.0464294
R1857 CSoutput.n272 CSoutput.n269 0.0391444
R1858 CSoutput.n231 CSoutput.t194 0.023435
R1859 CSoutput.n279 CSoutput.t186 0.02262
R1860 CSoutput.n230 CSoutput.t191 0.02262
R1861 CSoutput CSoutput.n413 0.0052
R1862 CSoutput.n201 CSoutput.n184 0.00365111
R1863 CSoutput.n204 CSoutput.n185 0.00365111
R1864 CSoutput.n187 CSoutput.n186 0.00365111
R1865 CSoutput.n229 CSoutput.n188 0.00365111
R1866 CSoutput.n193 CSoutput.n189 0.00365111
R1867 CSoutput.n276 CSoutput.n190 0.00365111
R1868 CSoutput.n267 CSoutput.n266 0.00365111
R1869 CSoutput.n247 CSoutput.n220 0.00365111
R1870 CSoutput.n249 CSoutput.n219 0.00365111
R1871 CSoutput.n237 CSoutput.n236 0.00365111
R1872 CSoutput.n243 CSoutput.n223 0.00365111
R1873 CSoutput.n245 CSoutput.n222 0.00365111
R1874 CSoutput.n167 CSoutput.n150 0.00365111
R1875 CSoutput.n170 CSoutput.n151 0.00365111
R1876 CSoutput.n153 CSoutput.n152 0.00365111
R1877 CSoutput.n263 CSoutput.n154 0.00365111
R1878 CSoutput.n159 CSoutput.n155 0.00365111
R1879 CSoutput.n286 CSoutput.n156 0.00365111
R1880 CSoutput.n198 CSoutput.n188 0.00340054
R1881 CSoutput.n191 CSoutput.n189 0.00340054
R1882 CSoutput.n276 CSoutput.n275 0.00340054
R1883 CSoutput.n271 CSoutput.n184 0.00340054
R1884 CSoutput.n200 CSoutput.n185 0.00340054
R1885 CSoutput.n203 CSoutput.n187 0.00340054
R1886 CSoutput.n242 CSoutput.n237 0.00340054
R1887 CSoutput.n244 CSoutput.n243 0.00340054
R1888 CSoutput.n246 CSoutput.n245 0.00340054
R1889 CSoutput.n268 CSoutput.n267 0.00340054
R1890 CSoutput.n248 CSoutput.n247 0.00340054
R1891 CSoutput.n250 CSoutput.n249 0.00340054
R1892 CSoutput.n164 CSoutput.n154 0.00340054
R1893 CSoutput.n157 CSoutput.n155 0.00340054
R1894 CSoutput.n286 CSoutput.n285 0.00340054
R1895 CSoutput.n281 CSoutput.n150 0.00340054
R1896 CSoutput.n166 CSoutput.n151 0.00340054
R1897 CSoutput.n169 CSoutput.n153 0.00340054
R1898 CSoutput.n199 CSoutput.n193 0.00252698
R1899 CSoutput.n192 CSoutput.n190 0.00252698
R1900 CSoutput.n274 CSoutput.n273 0.00252698
R1901 CSoutput.n202 CSoutput.n200 0.00252698
R1902 CSoutput.n205 CSoutput.n203 0.00252698
R1903 CSoutput.n278 CSoutput.n173 0.00252698
R1904 CSoutput.n199 CSoutput.n198 0.00252698
R1905 CSoutput.n192 CSoutput.n191 0.00252698
R1906 CSoutput.n275 CSoutput.n274 0.00252698
R1907 CSoutput.n202 CSoutput.n201 0.00252698
R1908 CSoutput.n205 CSoutput.n204 0.00252698
R1909 CSoutput.n186 CSoutput.n173 0.00252698
R1910 CSoutput.n253 CSoutput.n223 0.00252698
R1911 CSoutput.n252 CSoutput.n222 0.00252698
R1912 CSoutput.n251 CSoutput.n207 0.00252698
R1913 CSoutput.n248 CSoutput.n218 0.00252698
R1914 CSoutput.n255 CSoutput.n250 0.00252698
R1915 CSoutput.n264 CSoutput.n257 0.00252698
R1916 CSoutput.n253 CSoutput.n242 0.00252698
R1917 CSoutput.n252 CSoutput.n244 0.00252698
R1918 CSoutput.n251 CSoutput.n246 0.00252698
R1919 CSoutput.n266 CSoutput.n218 0.00252698
R1920 CSoutput.n255 CSoutput.n220 0.00252698
R1921 CSoutput.n257 CSoutput.n219 0.00252698
R1922 CSoutput.n165 CSoutput.n159 0.00252698
R1923 CSoutput.n158 CSoutput.n156 0.00252698
R1924 CSoutput.n284 CSoutput.n283 0.00252698
R1925 CSoutput.n168 CSoutput.n166 0.00252698
R1926 CSoutput.n171 CSoutput.n169 0.00252698
R1927 CSoutput.n288 CSoutput.n139 0.00252698
R1928 CSoutput.n165 CSoutput.n164 0.00252698
R1929 CSoutput.n158 CSoutput.n157 0.00252698
R1930 CSoutput.n285 CSoutput.n284 0.00252698
R1931 CSoutput.n168 CSoutput.n167 0.00252698
R1932 CSoutput.n171 CSoutput.n170 0.00252698
R1933 CSoutput.n152 CSoutput.n139 0.00252698
R1934 CSoutput.n273 CSoutput.n272 0.0020275
R1935 CSoutput.n272 CSoutput.n271 0.0020275
R1936 CSoutput.n269 CSoutput.n207 0.0020275
R1937 CSoutput.n269 CSoutput.n268 0.0020275
R1938 CSoutput.n283 CSoutput.n282 0.0020275
R1939 CSoutput.n282 CSoutput.n281 0.0020275
R1940 CSoutput.n183 CSoutput.n182 0.00166668
R1941 CSoutput.n265 CSoutput.n221 0.00166668
R1942 CSoutput.n149 CSoutput.n148 0.00166668
R1943 CSoutput.n287 CSoutput.n149 0.00133328
R1944 CSoutput.n221 CSoutput.n217 0.00133328
R1945 CSoutput.n277 CSoutput.n183 0.00133328
R1946 CSoutput.n280 CSoutput.n172 0.001
R1947 CSoutput.n258 CSoutput.n172 0.001
R1948 CSoutput.n160 CSoutput.n140 0.001
R1949 CSoutput.n259 CSoutput.n140 0.001
R1950 CSoutput.n161 CSoutput.n141 0.001
R1951 CSoutput.n260 CSoutput.n141 0.001
R1952 CSoutput.n162 CSoutput.n142 0.001
R1953 CSoutput.n261 CSoutput.n142 0.001
R1954 CSoutput.n163 CSoutput.n143 0.001
R1955 CSoutput.n262 CSoutput.n143 0.001
R1956 CSoutput.n256 CSoutput.n208 0.001
R1957 CSoutput.n256 CSoutput.n254 0.001
R1958 CSoutput.n238 CSoutput.n209 0.001
R1959 CSoutput.n232 CSoutput.n209 0.001
R1960 CSoutput.n239 CSoutput.n210 0.001
R1961 CSoutput.n233 CSoutput.n210 0.001
R1962 CSoutput.n240 CSoutput.n211 0.001
R1963 CSoutput.n234 CSoutput.n211 0.001
R1964 CSoutput.n241 CSoutput.n212 0.001
R1965 CSoutput.n235 CSoutput.n212 0.001
R1966 CSoutput.n270 CSoutput.n206 0.001
R1967 CSoutput.n224 CSoutput.n206 0.001
R1968 CSoutput.n194 CSoutput.n174 0.001
R1969 CSoutput.n225 CSoutput.n174 0.001
R1970 CSoutput.n195 CSoutput.n175 0.001
R1971 CSoutput.n226 CSoutput.n175 0.001
R1972 CSoutput.n196 CSoutput.n176 0.001
R1973 CSoutput.n227 CSoutput.n176 0.001
R1974 CSoutput.n197 CSoutput.n177 0.001
R1975 CSoutput.n228 CSoutput.n177 0.001
R1976 CSoutput.n228 CSoutput.n178 0.001
R1977 CSoutput.n227 CSoutput.n179 0.001
R1978 CSoutput.n226 CSoutput.n180 0.001
R1979 CSoutput.n225 CSoutput.t203 0.001
R1980 CSoutput.n224 CSoutput.n181 0.001
R1981 CSoutput.n197 CSoutput.n179 0.001
R1982 CSoutput.n196 CSoutput.n180 0.001
R1983 CSoutput.n195 CSoutput.t203 0.001
R1984 CSoutput.n194 CSoutput.n181 0.001
R1985 CSoutput.n270 CSoutput.n182 0.001
R1986 CSoutput.n235 CSoutput.n213 0.001
R1987 CSoutput.n234 CSoutput.n214 0.001
R1988 CSoutput.n233 CSoutput.n215 0.001
R1989 CSoutput.n232 CSoutput.t184 0.001
R1990 CSoutput.n254 CSoutput.n216 0.001
R1991 CSoutput.n241 CSoutput.n214 0.001
R1992 CSoutput.n240 CSoutput.n215 0.001
R1993 CSoutput.n239 CSoutput.t184 0.001
R1994 CSoutput.n238 CSoutput.n216 0.001
R1995 CSoutput.n265 CSoutput.n208 0.001
R1996 CSoutput.n262 CSoutput.n144 0.001
R1997 CSoutput.n261 CSoutput.n145 0.001
R1998 CSoutput.n260 CSoutput.n146 0.001
R1999 CSoutput.n259 CSoutput.t193 0.001
R2000 CSoutput.n258 CSoutput.n147 0.001
R2001 CSoutput.n163 CSoutput.n145 0.001
R2002 CSoutput.n162 CSoutput.n146 0.001
R2003 CSoutput.n161 CSoutput.t193 0.001
R2004 CSoutput.n160 CSoutput.n147 0.001
R2005 CSoutput.n280 CSoutput.n148 0.001
R2006 gnd.n6609 gnd.n685 1490.86
R2007 gnd.n3920 gnd.n3919 939.716
R2008 gnd.n7178 gnd.n103 795.207
R2009 gnd.n7328 gnd.n99 795.207
R2010 gnd.n6893 gnd.n423 795.207
R2011 gnd.n5701 gnd.n386 795.207
R2012 gnd.n5934 gnd.n1267 795.207
R2013 gnd.n4564 gnd.n1270 795.207
R2014 gnd.n4172 gnd.n3922 795.207
R2015 gnd.n4213 gnd.n4097 795.207
R2016 gnd.n7326 gnd.n105 775.989
R2017 gnd.n173 gnd.n101 775.989
R2018 gnd.n6896 gnd.n6895 775.989
R2019 gnd.n6968 gnd.n390 775.989
R2020 gnd.n5932 gnd.n1272 775.989
R2021 gnd.n5863 gnd.n1269 775.989
R2022 gnd.n4061 gnd.n3921 775.989
R2023 gnd.n4215 gnd.n2456 775.989
R2024 gnd.n4555 gnd.n2199 771.183
R2025 gnd.n5707 gnd.n1474 771.183
R2026 gnd.n2281 gnd.n1367 771.183
R2027 gnd.n5709 gnd.n1470 771.183
R2028 gnd.n3827 gnd.n2458 766.379
R2029 gnd.n3830 gnd.n3829 766.379
R2030 gnd.n3069 gnd.n2972 766.379
R2031 gnd.n3065 gnd.n2970 766.379
R2032 gnd.n3918 gnd.n2480 756.769
R2033 gnd.n3821 gnd.n3820 756.769
R2034 gnd.n3162 gnd.n2879 756.769
R2035 gnd.n3160 gnd.n2882 756.769
R2036 gnd.n6190 gnd.n938 756.769
R2037 gnd.n6610 gnd.n686 756.769
R2038 gnd.n6823 gnd.n559 756.769
R2039 gnd.n6022 gnd.n1108 756.769
R2040 gnd.n6191 gnd.n6190 585
R2041 gnd.n6190 gnd.n6189 585
R2042 gnd.n942 gnd.n941 585
R2043 gnd.n6188 gnd.n942 585
R2044 gnd.n6186 gnd.n6185 585
R2045 gnd.n6187 gnd.n6186 585
R2046 gnd.n6184 gnd.n944 585
R2047 gnd.n944 gnd.n943 585
R2048 gnd.n6183 gnd.n6182 585
R2049 gnd.n6182 gnd.n6181 585
R2050 gnd.n949 gnd.n948 585
R2051 gnd.n6180 gnd.n949 585
R2052 gnd.n6178 gnd.n6177 585
R2053 gnd.n6179 gnd.n6178 585
R2054 gnd.n6176 gnd.n951 585
R2055 gnd.n951 gnd.n950 585
R2056 gnd.n6175 gnd.n6174 585
R2057 gnd.n6174 gnd.n6173 585
R2058 gnd.n957 gnd.n956 585
R2059 gnd.n6172 gnd.n957 585
R2060 gnd.n6170 gnd.n6169 585
R2061 gnd.n6171 gnd.n6170 585
R2062 gnd.n6168 gnd.n959 585
R2063 gnd.n959 gnd.n958 585
R2064 gnd.n6167 gnd.n6166 585
R2065 gnd.n6166 gnd.n6165 585
R2066 gnd.n965 gnd.n964 585
R2067 gnd.n6164 gnd.n965 585
R2068 gnd.n6162 gnd.n6161 585
R2069 gnd.n6163 gnd.n6162 585
R2070 gnd.n6160 gnd.n967 585
R2071 gnd.n967 gnd.n966 585
R2072 gnd.n6159 gnd.n6158 585
R2073 gnd.n6158 gnd.n6157 585
R2074 gnd.n973 gnd.n972 585
R2075 gnd.n6156 gnd.n973 585
R2076 gnd.n6154 gnd.n6153 585
R2077 gnd.n6155 gnd.n6154 585
R2078 gnd.n6152 gnd.n975 585
R2079 gnd.n975 gnd.n974 585
R2080 gnd.n6151 gnd.n6150 585
R2081 gnd.n6150 gnd.n6149 585
R2082 gnd.n981 gnd.n980 585
R2083 gnd.n6148 gnd.n981 585
R2084 gnd.n6146 gnd.n6145 585
R2085 gnd.n6147 gnd.n6146 585
R2086 gnd.n6144 gnd.n983 585
R2087 gnd.n983 gnd.n982 585
R2088 gnd.n6143 gnd.n6142 585
R2089 gnd.n6142 gnd.n6141 585
R2090 gnd.n989 gnd.n988 585
R2091 gnd.n6140 gnd.n989 585
R2092 gnd.n6138 gnd.n6137 585
R2093 gnd.n6139 gnd.n6138 585
R2094 gnd.n6136 gnd.n991 585
R2095 gnd.n991 gnd.n990 585
R2096 gnd.n6135 gnd.n6134 585
R2097 gnd.n6134 gnd.n6133 585
R2098 gnd.n997 gnd.n996 585
R2099 gnd.n6132 gnd.n997 585
R2100 gnd.n6130 gnd.n6129 585
R2101 gnd.n6131 gnd.n6130 585
R2102 gnd.n6128 gnd.n999 585
R2103 gnd.n999 gnd.n998 585
R2104 gnd.n6127 gnd.n6126 585
R2105 gnd.n6126 gnd.n6125 585
R2106 gnd.n1005 gnd.n1004 585
R2107 gnd.n6124 gnd.n1005 585
R2108 gnd.n6122 gnd.n6121 585
R2109 gnd.n6123 gnd.n6122 585
R2110 gnd.n6120 gnd.n1007 585
R2111 gnd.n1007 gnd.n1006 585
R2112 gnd.n6119 gnd.n6118 585
R2113 gnd.n6118 gnd.n6117 585
R2114 gnd.n1013 gnd.n1012 585
R2115 gnd.n6116 gnd.n1013 585
R2116 gnd.n6114 gnd.n6113 585
R2117 gnd.n6115 gnd.n6114 585
R2118 gnd.n6112 gnd.n1015 585
R2119 gnd.n1015 gnd.n1014 585
R2120 gnd.n6111 gnd.n6110 585
R2121 gnd.n6110 gnd.n6109 585
R2122 gnd.n1021 gnd.n1020 585
R2123 gnd.n6108 gnd.n1021 585
R2124 gnd.n6106 gnd.n6105 585
R2125 gnd.n6107 gnd.n6106 585
R2126 gnd.n6104 gnd.n1023 585
R2127 gnd.n1023 gnd.n1022 585
R2128 gnd.n6103 gnd.n6102 585
R2129 gnd.n6102 gnd.n6101 585
R2130 gnd.n1029 gnd.n1028 585
R2131 gnd.n6100 gnd.n1029 585
R2132 gnd.n6098 gnd.n6097 585
R2133 gnd.n6099 gnd.n6098 585
R2134 gnd.n6096 gnd.n1031 585
R2135 gnd.n1031 gnd.n1030 585
R2136 gnd.n6095 gnd.n6094 585
R2137 gnd.n6094 gnd.n6093 585
R2138 gnd.n1037 gnd.n1036 585
R2139 gnd.n6092 gnd.n1037 585
R2140 gnd.n6090 gnd.n6089 585
R2141 gnd.n6091 gnd.n6090 585
R2142 gnd.n6088 gnd.n1039 585
R2143 gnd.n1039 gnd.n1038 585
R2144 gnd.n6087 gnd.n6086 585
R2145 gnd.n6086 gnd.n6085 585
R2146 gnd.n1045 gnd.n1044 585
R2147 gnd.n6084 gnd.n1045 585
R2148 gnd.n6082 gnd.n6081 585
R2149 gnd.n6083 gnd.n6082 585
R2150 gnd.n6080 gnd.n1047 585
R2151 gnd.n1047 gnd.n1046 585
R2152 gnd.n6079 gnd.n6078 585
R2153 gnd.n6078 gnd.n6077 585
R2154 gnd.n1053 gnd.n1052 585
R2155 gnd.n6076 gnd.n1053 585
R2156 gnd.n6074 gnd.n6073 585
R2157 gnd.n6075 gnd.n6074 585
R2158 gnd.n6072 gnd.n1055 585
R2159 gnd.n1055 gnd.n1054 585
R2160 gnd.n6071 gnd.n6070 585
R2161 gnd.n6070 gnd.n6069 585
R2162 gnd.n1061 gnd.n1060 585
R2163 gnd.n6068 gnd.n1061 585
R2164 gnd.n6066 gnd.n6065 585
R2165 gnd.n6067 gnd.n6066 585
R2166 gnd.n6064 gnd.n1063 585
R2167 gnd.n1063 gnd.n1062 585
R2168 gnd.n6063 gnd.n6062 585
R2169 gnd.n6062 gnd.n6061 585
R2170 gnd.n1069 gnd.n1068 585
R2171 gnd.n6060 gnd.n1069 585
R2172 gnd.n6058 gnd.n6057 585
R2173 gnd.n6059 gnd.n6058 585
R2174 gnd.n6056 gnd.n1071 585
R2175 gnd.n1071 gnd.n1070 585
R2176 gnd.n6055 gnd.n6054 585
R2177 gnd.n6054 gnd.n6053 585
R2178 gnd.n1077 gnd.n1076 585
R2179 gnd.n6052 gnd.n1077 585
R2180 gnd.n6050 gnd.n6049 585
R2181 gnd.n6051 gnd.n6050 585
R2182 gnd.n6048 gnd.n1079 585
R2183 gnd.n1079 gnd.n1078 585
R2184 gnd.n6047 gnd.n6046 585
R2185 gnd.n6046 gnd.n6045 585
R2186 gnd.n1085 gnd.n1084 585
R2187 gnd.n6044 gnd.n1085 585
R2188 gnd.n6042 gnd.n6041 585
R2189 gnd.n6043 gnd.n6042 585
R2190 gnd.n6040 gnd.n1087 585
R2191 gnd.n1087 gnd.n1086 585
R2192 gnd.n6039 gnd.n6038 585
R2193 gnd.n6038 gnd.n6037 585
R2194 gnd.n1093 gnd.n1092 585
R2195 gnd.n6036 gnd.n1093 585
R2196 gnd.n6034 gnd.n6033 585
R2197 gnd.n6035 gnd.n6034 585
R2198 gnd.n6032 gnd.n1095 585
R2199 gnd.n1095 gnd.n1094 585
R2200 gnd.n6031 gnd.n6030 585
R2201 gnd.n6030 gnd.n6029 585
R2202 gnd.n1101 gnd.n1100 585
R2203 gnd.n6028 gnd.n1101 585
R2204 gnd.n6026 gnd.n6025 585
R2205 gnd.n6027 gnd.n6026 585
R2206 gnd.n6024 gnd.n1103 585
R2207 gnd.n1103 gnd.n1102 585
R2208 gnd.n939 gnd.n938 585
R2209 gnd.n938 gnd.n937 585
R2210 gnd.n6196 gnd.n6195 585
R2211 gnd.n6197 gnd.n6196 585
R2212 gnd.n936 gnd.n935 585
R2213 gnd.n6198 gnd.n936 585
R2214 gnd.n6201 gnd.n6200 585
R2215 gnd.n6200 gnd.n6199 585
R2216 gnd.n933 gnd.n932 585
R2217 gnd.n932 gnd.n931 585
R2218 gnd.n6206 gnd.n6205 585
R2219 gnd.n6207 gnd.n6206 585
R2220 gnd.n930 gnd.n929 585
R2221 gnd.n6208 gnd.n930 585
R2222 gnd.n6211 gnd.n6210 585
R2223 gnd.n6210 gnd.n6209 585
R2224 gnd.n927 gnd.n926 585
R2225 gnd.n926 gnd.n925 585
R2226 gnd.n6216 gnd.n6215 585
R2227 gnd.n6217 gnd.n6216 585
R2228 gnd.n924 gnd.n923 585
R2229 gnd.n6218 gnd.n924 585
R2230 gnd.n6221 gnd.n6220 585
R2231 gnd.n6220 gnd.n6219 585
R2232 gnd.n921 gnd.n920 585
R2233 gnd.n920 gnd.n919 585
R2234 gnd.n6226 gnd.n6225 585
R2235 gnd.n6227 gnd.n6226 585
R2236 gnd.n918 gnd.n917 585
R2237 gnd.n6228 gnd.n918 585
R2238 gnd.n6231 gnd.n6230 585
R2239 gnd.n6230 gnd.n6229 585
R2240 gnd.n915 gnd.n914 585
R2241 gnd.n914 gnd.n913 585
R2242 gnd.n6236 gnd.n6235 585
R2243 gnd.n6237 gnd.n6236 585
R2244 gnd.n912 gnd.n911 585
R2245 gnd.n6238 gnd.n912 585
R2246 gnd.n6241 gnd.n6240 585
R2247 gnd.n6240 gnd.n6239 585
R2248 gnd.n909 gnd.n908 585
R2249 gnd.n908 gnd.n907 585
R2250 gnd.n6246 gnd.n6245 585
R2251 gnd.n6247 gnd.n6246 585
R2252 gnd.n906 gnd.n905 585
R2253 gnd.n6248 gnd.n906 585
R2254 gnd.n6251 gnd.n6250 585
R2255 gnd.n6250 gnd.n6249 585
R2256 gnd.n903 gnd.n902 585
R2257 gnd.n902 gnd.n901 585
R2258 gnd.n6256 gnd.n6255 585
R2259 gnd.n6257 gnd.n6256 585
R2260 gnd.n900 gnd.n899 585
R2261 gnd.n6258 gnd.n900 585
R2262 gnd.n6261 gnd.n6260 585
R2263 gnd.n6260 gnd.n6259 585
R2264 gnd.n897 gnd.n896 585
R2265 gnd.n896 gnd.n895 585
R2266 gnd.n6266 gnd.n6265 585
R2267 gnd.n6267 gnd.n6266 585
R2268 gnd.n894 gnd.n893 585
R2269 gnd.n6268 gnd.n894 585
R2270 gnd.n6271 gnd.n6270 585
R2271 gnd.n6270 gnd.n6269 585
R2272 gnd.n891 gnd.n890 585
R2273 gnd.n890 gnd.n889 585
R2274 gnd.n6276 gnd.n6275 585
R2275 gnd.n6277 gnd.n6276 585
R2276 gnd.n888 gnd.n887 585
R2277 gnd.n6278 gnd.n888 585
R2278 gnd.n6281 gnd.n6280 585
R2279 gnd.n6280 gnd.n6279 585
R2280 gnd.n885 gnd.n884 585
R2281 gnd.n884 gnd.n883 585
R2282 gnd.n6286 gnd.n6285 585
R2283 gnd.n6287 gnd.n6286 585
R2284 gnd.n882 gnd.n881 585
R2285 gnd.n6288 gnd.n882 585
R2286 gnd.n6291 gnd.n6290 585
R2287 gnd.n6290 gnd.n6289 585
R2288 gnd.n879 gnd.n878 585
R2289 gnd.n878 gnd.n877 585
R2290 gnd.n6296 gnd.n6295 585
R2291 gnd.n6297 gnd.n6296 585
R2292 gnd.n876 gnd.n875 585
R2293 gnd.n6298 gnd.n876 585
R2294 gnd.n6301 gnd.n6300 585
R2295 gnd.n6300 gnd.n6299 585
R2296 gnd.n873 gnd.n872 585
R2297 gnd.n872 gnd.n871 585
R2298 gnd.n6306 gnd.n6305 585
R2299 gnd.n6307 gnd.n6306 585
R2300 gnd.n870 gnd.n869 585
R2301 gnd.n6308 gnd.n870 585
R2302 gnd.n6311 gnd.n6310 585
R2303 gnd.n6310 gnd.n6309 585
R2304 gnd.n867 gnd.n866 585
R2305 gnd.n866 gnd.n865 585
R2306 gnd.n6316 gnd.n6315 585
R2307 gnd.n6317 gnd.n6316 585
R2308 gnd.n864 gnd.n863 585
R2309 gnd.n6318 gnd.n864 585
R2310 gnd.n6321 gnd.n6320 585
R2311 gnd.n6320 gnd.n6319 585
R2312 gnd.n861 gnd.n860 585
R2313 gnd.n860 gnd.n859 585
R2314 gnd.n6326 gnd.n6325 585
R2315 gnd.n6327 gnd.n6326 585
R2316 gnd.n858 gnd.n857 585
R2317 gnd.n6328 gnd.n858 585
R2318 gnd.n6331 gnd.n6330 585
R2319 gnd.n6330 gnd.n6329 585
R2320 gnd.n855 gnd.n854 585
R2321 gnd.n854 gnd.n853 585
R2322 gnd.n6336 gnd.n6335 585
R2323 gnd.n6337 gnd.n6336 585
R2324 gnd.n852 gnd.n851 585
R2325 gnd.n6338 gnd.n852 585
R2326 gnd.n6341 gnd.n6340 585
R2327 gnd.n6340 gnd.n6339 585
R2328 gnd.n849 gnd.n848 585
R2329 gnd.n848 gnd.n847 585
R2330 gnd.n6346 gnd.n6345 585
R2331 gnd.n6347 gnd.n6346 585
R2332 gnd.n846 gnd.n845 585
R2333 gnd.n6348 gnd.n846 585
R2334 gnd.n6351 gnd.n6350 585
R2335 gnd.n6350 gnd.n6349 585
R2336 gnd.n843 gnd.n842 585
R2337 gnd.n842 gnd.n841 585
R2338 gnd.n6356 gnd.n6355 585
R2339 gnd.n6357 gnd.n6356 585
R2340 gnd.n840 gnd.n839 585
R2341 gnd.n6358 gnd.n840 585
R2342 gnd.n6361 gnd.n6360 585
R2343 gnd.n6360 gnd.n6359 585
R2344 gnd.n837 gnd.n836 585
R2345 gnd.n836 gnd.n835 585
R2346 gnd.n6366 gnd.n6365 585
R2347 gnd.n6367 gnd.n6366 585
R2348 gnd.n834 gnd.n833 585
R2349 gnd.n6368 gnd.n834 585
R2350 gnd.n6371 gnd.n6370 585
R2351 gnd.n6370 gnd.n6369 585
R2352 gnd.n831 gnd.n830 585
R2353 gnd.n830 gnd.n829 585
R2354 gnd.n6376 gnd.n6375 585
R2355 gnd.n6377 gnd.n6376 585
R2356 gnd.n828 gnd.n827 585
R2357 gnd.n6378 gnd.n828 585
R2358 gnd.n6381 gnd.n6380 585
R2359 gnd.n6380 gnd.n6379 585
R2360 gnd.n825 gnd.n824 585
R2361 gnd.n824 gnd.n823 585
R2362 gnd.n6386 gnd.n6385 585
R2363 gnd.n6387 gnd.n6386 585
R2364 gnd.n822 gnd.n821 585
R2365 gnd.n6388 gnd.n822 585
R2366 gnd.n6391 gnd.n6390 585
R2367 gnd.n6390 gnd.n6389 585
R2368 gnd.n819 gnd.n818 585
R2369 gnd.n818 gnd.n817 585
R2370 gnd.n6396 gnd.n6395 585
R2371 gnd.n6397 gnd.n6396 585
R2372 gnd.n816 gnd.n815 585
R2373 gnd.n6398 gnd.n816 585
R2374 gnd.n6401 gnd.n6400 585
R2375 gnd.n6400 gnd.n6399 585
R2376 gnd.n813 gnd.n812 585
R2377 gnd.n812 gnd.n811 585
R2378 gnd.n6406 gnd.n6405 585
R2379 gnd.n6407 gnd.n6406 585
R2380 gnd.n810 gnd.n809 585
R2381 gnd.n6408 gnd.n810 585
R2382 gnd.n6411 gnd.n6410 585
R2383 gnd.n6410 gnd.n6409 585
R2384 gnd.n807 gnd.n806 585
R2385 gnd.n806 gnd.n805 585
R2386 gnd.n6416 gnd.n6415 585
R2387 gnd.n6417 gnd.n6416 585
R2388 gnd.n804 gnd.n803 585
R2389 gnd.n6418 gnd.n804 585
R2390 gnd.n6421 gnd.n6420 585
R2391 gnd.n6420 gnd.n6419 585
R2392 gnd.n801 gnd.n800 585
R2393 gnd.n800 gnd.n799 585
R2394 gnd.n6426 gnd.n6425 585
R2395 gnd.n6427 gnd.n6426 585
R2396 gnd.n798 gnd.n797 585
R2397 gnd.n6428 gnd.n798 585
R2398 gnd.n6431 gnd.n6430 585
R2399 gnd.n6430 gnd.n6429 585
R2400 gnd.n795 gnd.n794 585
R2401 gnd.n794 gnd.n793 585
R2402 gnd.n6436 gnd.n6435 585
R2403 gnd.n6437 gnd.n6436 585
R2404 gnd.n792 gnd.n791 585
R2405 gnd.n6438 gnd.n792 585
R2406 gnd.n6441 gnd.n6440 585
R2407 gnd.n6440 gnd.n6439 585
R2408 gnd.n789 gnd.n788 585
R2409 gnd.n788 gnd.n787 585
R2410 gnd.n6446 gnd.n6445 585
R2411 gnd.n6447 gnd.n6446 585
R2412 gnd.n786 gnd.n785 585
R2413 gnd.n6448 gnd.n786 585
R2414 gnd.n6451 gnd.n6450 585
R2415 gnd.n6450 gnd.n6449 585
R2416 gnd.n783 gnd.n782 585
R2417 gnd.n782 gnd.n781 585
R2418 gnd.n6456 gnd.n6455 585
R2419 gnd.n6457 gnd.n6456 585
R2420 gnd.n780 gnd.n779 585
R2421 gnd.n6458 gnd.n780 585
R2422 gnd.n6461 gnd.n6460 585
R2423 gnd.n6460 gnd.n6459 585
R2424 gnd.n777 gnd.n776 585
R2425 gnd.n776 gnd.n775 585
R2426 gnd.n6466 gnd.n6465 585
R2427 gnd.n6467 gnd.n6466 585
R2428 gnd.n774 gnd.n773 585
R2429 gnd.n6468 gnd.n774 585
R2430 gnd.n6471 gnd.n6470 585
R2431 gnd.n6470 gnd.n6469 585
R2432 gnd.n771 gnd.n770 585
R2433 gnd.n770 gnd.n769 585
R2434 gnd.n6476 gnd.n6475 585
R2435 gnd.n6477 gnd.n6476 585
R2436 gnd.n768 gnd.n767 585
R2437 gnd.n6478 gnd.n768 585
R2438 gnd.n6481 gnd.n6480 585
R2439 gnd.n6480 gnd.n6479 585
R2440 gnd.n765 gnd.n764 585
R2441 gnd.n764 gnd.n763 585
R2442 gnd.n6486 gnd.n6485 585
R2443 gnd.n6487 gnd.n6486 585
R2444 gnd.n762 gnd.n761 585
R2445 gnd.n6488 gnd.n762 585
R2446 gnd.n6491 gnd.n6490 585
R2447 gnd.n6490 gnd.n6489 585
R2448 gnd.n759 gnd.n758 585
R2449 gnd.n758 gnd.n757 585
R2450 gnd.n6496 gnd.n6495 585
R2451 gnd.n6497 gnd.n6496 585
R2452 gnd.n756 gnd.n755 585
R2453 gnd.n6498 gnd.n756 585
R2454 gnd.n6501 gnd.n6500 585
R2455 gnd.n6500 gnd.n6499 585
R2456 gnd.n753 gnd.n752 585
R2457 gnd.n752 gnd.n751 585
R2458 gnd.n6506 gnd.n6505 585
R2459 gnd.n6507 gnd.n6506 585
R2460 gnd.n750 gnd.n749 585
R2461 gnd.n6508 gnd.n750 585
R2462 gnd.n6511 gnd.n6510 585
R2463 gnd.n6510 gnd.n6509 585
R2464 gnd.n747 gnd.n746 585
R2465 gnd.n746 gnd.n745 585
R2466 gnd.n6516 gnd.n6515 585
R2467 gnd.n6517 gnd.n6516 585
R2468 gnd.n744 gnd.n743 585
R2469 gnd.n6518 gnd.n744 585
R2470 gnd.n6521 gnd.n6520 585
R2471 gnd.n6520 gnd.n6519 585
R2472 gnd.n741 gnd.n740 585
R2473 gnd.n740 gnd.n739 585
R2474 gnd.n6526 gnd.n6525 585
R2475 gnd.n6527 gnd.n6526 585
R2476 gnd.n738 gnd.n737 585
R2477 gnd.n6528 gnd.n738 585
R2478 gnd.n6531 gnd.n6530 585
R2479 gnd.n6530 gnd.n6529 585
R2480 gnd.n735 gnd.n734 585
R2481 gnd.n734 gnd.n733 585
R2482 gnd.n6536 gnd.n6535 585
R2483 gnd.n6537 gnd.n6536 585
R2484 gnd.n732 gnd.n731 585
R2485 gnd.n6538 gnd.n732 585
R2486 gnd.n6541 gnd.n6540 585
R2487 gnd.n6540 gnd.n6539 585
R2488 gnd.n729 gnd.n728 585
R2489 gnd.n728 gnd.n727 585
R2490 gnd.n6546 gnd.n6545 585
R2491 gnd.n6547 gnd.n6546 585
R2492 gnd.n726 gnd.n725 585
R2493 gnd.n6548 gnd.n726 585
R2494 gnd.n6551 gnd.n6550 585
R2495 gnd.n6550 gnd.n6549 585
R2496 gnd.n723 gnd.n722 585
R2497 gnd.n722 gnd.n721 585
R2498 gnd.n6556 gnd.n6555 585
R2499 gnd.n6557 gnd.n6556 585
R2500 gnd.n720 gnd.n719 585
R2501 gnd.n6558 gnd.n720 585
R2502 gnd.n6561 gnd.n6560 585
R2503 gnd.n6560 gnd.n6559 585
R2504 gnd.n717 gnd.n716 585
R2505 gnd.n716 gnd.n715 585
R2506 gnd.n6566 gnd.n6565 585
R2507 gnd.n6567 gnd.n6566 585
R2508 gnd.n714 gnd.n713 585
R2509 gnd.n6568 gnd.n714 585
R2510 gnd.n6571 gnd.n6570 585
R2511 gnd.n6570 gnd.n6569 585
R2512 gnd.n711 gnd.n710 585
R2513 gnd.n710 gnd.n709 585
R2514 gnd.n6576 gnd.n6575 585
R2515 gnd.n6577 gnd.n6576 585
R2516 gnd.n708 gnd.n707 585
R2517 gnd.n6578 gnd.n708 585
R2518 gnd.n6581 gnd.n6580 585
R2519 gnd.n6580 gnd.n6579 585
R2520 gnd.n705 gnd.n704 585
R2521 gnd.n704 gnd.n703 585
R2522 gnd.n6586 gnd.n6585 585
R2523 gnd.n6587 gnd.n6586 585
R2524 gnd.n702 gnd.n701 585
R2525 gnd.n6588 gnd.n702 585
R2526 gnd.n6591 gnd.n6590 585
R2527 gnd.n6590 gnd.n6589 585
R2528 gnd.n699 gnd.n698 585
R2529 gnd.n698 gnd.n697 585
R2530 gnd.n6596 gnd.n6595 585
R2531 gnd.n6597 gnd.n6596 585
R2532 gnd.n696 gnd.n695 585
R2533 gnd.n6598 gnd.n696 585
R2534 gnd.n6601 gnd.n6600 585
R2535 gnd.n6600 gnd.n6599 585
R2536 gnd.n693 gnd.n692 585
R2537 gnd.n692 gnd.n691 585
R2538 gnd.n6606 gnd.n6605 585
R2539 gnd.n6607 gnd.n6606 585
R2540 gnd.n690 gnd.n689 585
R2541 gnd.n6608 gnd.n690 585
R2542 gnd.n6611 gnd.n6610 585
R2543 gnd.n6610 gnd.n6609 585
R2544 gnd.n6822 gnd.n563 585
R2545 gnd.n6822 gnd.n6821 585
R2546 gnd.n6816 gnd.n564 585
R2547 gnd.n6820 gnd.n564 585
R2548 gnd.n6818 gnd.n6817 585
R2549 gnd.n6819 gnd.n6818 585
R2550 gnd.n567 gnd.n566 585
R2551 gnd.n566 gnd.n565 585
R2552 gnd.n6811 gnd.n6810 585
R2553 gnd.n6810 gnd.n6809 585
R2554 gnd.n570 gnd.n569 585
R2555 gnd.n6808 gnd.n570 585
R2556 gnd.n6806 gnd.n6805 585
R2557 gnd.n6807 gnd.n6806 585
R2558 gnd.n573 gnd.n572 585
R2559 gnd.n572 gnd.n571 585
R2560 gnd.n6801 gnd.n6800 585
R2561 gnd.n6800 gnd.n6799 585
R2562 gnd.n576 gnd.n575 585
R2563 gnd.n6798 gnd.n576 585
R2564 gnd.n6796 gnd.n6795 585
R2565 gnd.n6797 gnd.n6796 585
R2566 gnd.n579 gnd.n578 585
R2567 gnd.n578 gnd.n577 585
R2568 gnd.n6791 gnd.n6790 585
R2569 gnd.n6790 gnd.n6789 585
R2570 gnd.n582 gnd.n581 585
R2571 gnd.n6788 gnd.n582 585
R2572 gnd.n6786 gnd.n6785 585
R2573 gnd.n6787 gnd.n6786 585
R2574 gnd.n585 gnd.n584 585
R2575 gnd.n584 gnd.n583 585
R2576 gnd.n6781 gnd.n6780 585
R2577 gnd.n6780 gnd.n6779 585
R2578 gnd.n588 gnd.n587 585
R2579 gnd.n6778 gnd.n588 585
R2580 gnd.n6776 gnd.n6775 585
R2581 gnd.n6777 gnd.n6776 585
R2582 gnd.n591 gnd.n590 585
R2583 gnd.n590 gnd.n589 585
R2584 gnd.n6771 gnd.n6770 585
R2585 gnd.n6770 gnd.n6769 585
R2586 gnd.n594 gnd.n593 585
R2587 gnd.n6768 gnd.n594 585
R2588 gnd.n6766 gnd.n6765 585
R2589 gnd.n6767 gnd.n6766 585
R2590 gnd.n597 gnd.n596 585
R2591 gnd.n596 gnd.n595 585
R2592 gnd.n6761 gnd.n6760 585
R2593 gnd.n6760 gnd.n6759 585
R2594 gnd.n600 gnd.n599 585
R2595 gnd.n6758 gnd.n600 585
R2596 gnd.n6756 gnd.n6755 585
R2597 gnd.n6757 gnd.n6756 585
R2598 gnd.n603 gnd.n602 585
R2599 gnd.n602 gnd.n601 585
R2600 gnd.n6751 gnd.n6750 585
R2601 gnd.n6750 gnd.n6749 585
R2602 gnd.n606 gnd.n605 585
R2603 gnd.n6748 gnd.n606 585
R2604 gnd.n6746 gnd.n6745 585
R2605 gnd.n6747 gnd.n6746 585
R2606 gnd.n609 gnd.n608 585
R2607 gnd.n608 gnd.n607 585
R2608 gnd.n6741 gnd.n6740 585
R2609 gnd.n6740 gnd.n6739 585
R2610 gnd.n612 gnd.n611 585
R2611 gnd.n6738 gnd.n612 585
R2612 gnd.n6736 gnd.n6735 585
R2613 gnd.n6737 gnd.n6736 585
R2614 gnd.n615 gnd.n614 585
R2615 gnd.n614 gnd.n613 585
R2616 gnd.n6731 gnd.n6730 585
R2617 gnd.n6730 gnd.n6729 585
R2618 gnd.n618 gnd.n617 585
R2619 gnd.n6728 gnd.n618 585
R2620 gnd.n6726 gnd.n6725 585
R2621 gnd.n6727 gnd.n6726 585
R2622 gnd.n621 gnd.n620 585
R2623 gnd.n620 gnd.n619 585
R2624 gnd.n6721 gnd.n6720 585
R2625 gnd.n6720 gnd.n6719 585
R2626 gnd.n624 gnd.n623 585
R2627 gnd.n6718 gnd.n624 585
R2628 gnd.n6716 gnd.n6715 585
R2629 gnd.n6717 gnd.n6716 585
R2630 gnd.n627 gnd.n626 585
R2631 gnd.n626 gnd.n625 585
R2632 gnd.n6711 gnd.n6710 585
R2633 gnd.n6710 gnd.n6709 585
R2634 gnd.n630 gnd.n629 585
R2635 gnd.n6708 gnd.n630 585
R2636 gnd.n6706 gnd.n6705 585
R2637 gnd.n6707 gnd.n6706 585
R2638 gnd.n633 gnd.n632 585
R2639 gnd.n632 gnd.n631 585
R2640 gnd.n6701 gnd.n6700 585
R2641 gnd.n6700 gnd.n6699 585
R2642 gnd.n636 gnd.n635 585
R2643 gnd.n6698 gnd.n636 585
R2644 gnd.n6696 gnd.n6695 585
R2645 gnd.n6697 gnd.n6696 585
R2646 gnd.n639 gnd.n638 585
R2647 gnd.n638 gnd.n637 585
R2648 gnd.n6691 gnd.n6690 585
R2649 gnd.n6690 gnd.n6689 585
R2650 gnd.n642 gnd.n641 585
R2651 gnd.n6688 gnd.n642 585
R2652 gnd.n6686 gnd.n6685 585
R2653 gnd.n6687 gnd.n6686 585
R2654 gnd.n645 gnd.n644 585
R2655 gnd.n644 gnd.n643 585
R2656 gnd.n6681 gnd.n6680 585
R2657 gnd.n6680 gnd.n6679 585
R2658 gnd.n648 gnd.n647 585
R2659 gnd.n6678 gnd.n648 585
R2660 gnd.n6676 gnd.n6675 585
R2661 gnd.n6677 gnd.n6676 585
R2662 gnd.n651 gnd.n650 585
R2663 gnd.n650 gnd.n649 585
R2664 gnd.n6671 gnd.n6670 585
R2665 gnd.n6670 gnd.n6669 585
R2666 gnd.n654 gnd.n653 585
R2667 gnd.n6668 gnd.n654 585
R2668 gnd.n6666 gnd.n6665 585
R2669 gnd.n6667 gnd.n6666 585
R2670 gnd.n657 gnd.n656 585
R2671 gnd.n656 gnd.n655 585
R2672 gnd.n6661 gnd.n6660 585
R2673 gnd.n6660 gnd.n6659 585
R2674 gnd.n660 gnd.n659 585
R2675 gnd.n6658 gnd.n660 585
R2676 gnd.n6656 gnd.n6655 585
R2677 gnd.n6657 gnd.n6656 585
R2678 gnd.n663 gnd.n662 585
R2679 gnd.n662 gnd.n661 585
R2680 gnd.n6651 gnd.n6650 585
R2681 gnd.n6650 gnd.n6649 585
R2682 gnd.n666 gnd.n665 585
R2683 gnd.n6648 gnd.n666 585
R2684 gnd.n6646 gnd.n6645 585
R2685 gnd.n6647 gnd.n6646 585
R2686 gnd.n669 gnd.n668 585
R2687 gnd.n668 gnd.n667 585
R2688 gnd.n6641 gnd.n6640 585
R2689 gnd.n6640 gnd.n6639 585
R2690 gnd.n672 gnd.n671 585
R2691 gnd.n6638 gnd.n672 585
R2692 gnd.n6636 gnd.n6635 585
R2693 gnd.n6637 gnd.n6636 585
R2694 gnd.n675 gnd.n674 585
R2695 gnd.n674 gnd.n673 585
R2696 gnd.n6631 gnd.n6630 585
R2697 gnd.n6630 gnd.n6629 585
R2698 gnd.n678 gnd.n677 585
R2699 gnd.n6628 gnd.n678 585
R2700 gnd.n6626 gnd.n6625 585
R2701 gnd.n6627 gnd.n6626 585
R2702 gnd.n681 gnd.n680 585
R2703 gnd.n680 gnd.n679 585
R2704 gnd.n6621 gnd.n6620 585
R2705 gnd.n6620 gnd.n6619 585
R2706 gnd.n684 gnd.n683 585
R2707 gnd.n6618 gnd.n684 585
R2708 gnd.n6616 gnd.n6615 585
R2709 gnd.n6617 gnd.n6616 585
R2710 gnd.n687 gnd.n686 585
R2711 gnd.n686 gnd.n685 585
R2712 gnd.n5935 gnd.n5934 585
R2713 gnd.n5934 gnd.n5933 585
R2714 gnd.n5936 gnd.n1262 585
R2715 gnd.n5856 gnd.n1262 585
R2716 gnd.n5938 gnd.n5937 585
R2717 gnd.n5939 gnd.n5938 585
R2718 gnd.n1246 gnd.n1245 585
R2719 gnd.n4511 gnd.n1246 585
R2720 gnd.n5947 gnd.n5946 585
R2721 gnd.n5946 gnd.n5945 585
R2722 gnd.n5948 gnd.n1240 585
R2723 gnd.n4502 gnd.n1240 585
R2724 gnd.n5950 gnd.n5949 585
R2725 gnd.n5951 gnd.n5950 585
R2726 gnd.n1225 gnd.n1224 585
R2727 gnd.n4522 gnd.n1225 585
R2728 gnd.n5959 gnd.n5958 585
R2729 gnd.n5958 gnd.n5957 585
R2730 gnd.n5960 gnd.n1219 585
R2731 gnd.n4494 gnd.n1219 585
R2732 gnd.n5962 gnd.n5961 585
R2733 gnd.n5963 gnd.n5962 585
R2734 gnd.n1204 gnd.n1203 585
R2735 gnd.n4486 gnd.n1204 585
R2736 gnd.n5971 gnd.n5970 585
R2737 gnd.n5970 gnd.n5969 585
R2738 gnd.n5972 gnd.n1198 585
R2739 gnd.n4478 gnd.n1198 585
R2740 gnd.n5974 gnd.n5973 585
R2741 gnd.n5975 gnd.n5974 585
R2742 gnd.n1183 gnd.n1182 585
R2743 gnd.n4470 gnd.n1183 585
R2744 gnd.n5983 gnd.n5982 585
R2745 gnd.n5982 gnd.n5981 585
R2746 gnd.n5984 gnd.n1177 585
R2747 gnd.n4416 gnd.n1177 585
R2748 gnd.n5986 gnd.n5985 585
R2749 gnd.n5987 gnd.n5986 585
R2750 gnd.n1163 gnd.n1162 585
R2751 gnd.n4404 gnd.n1163 585
R2752 gnd.n5995 gnd.n5994 585
R2753 gnd.n5994 gnd.n5993 585
R2754 gnd.n5996 gnd.n1157 585
R2755 gnd.n4399 gnd.n1157 585
R2756 gnd.n5998 gnd.n5997 585
R2757 gnd.n5999 gnd.n5998 585
R2758 gnd.n1158 gnd.n1156 585
R2759 gnd.n4430 gnd.n1156 585
R2760 gnd.n4384 gnd.n2350 585
R2761 gnd.n4392 gnd.n2350 585
R2762 gnd.n4386 gnd.n4385 585
R2763 gnd.n4387 gnd.n4386 585
R2764 gnd.n2354 gnd.n2353 585
R2765 gnd.n4374 gnd.n2353 585
R2766 gnd.n4351 gnd.n2368 585
R2767 gnd.n4362 gnd.n2368 585
R2768 gnd.n4352 gnd.n2375 585
R2769 gnd.n2375 gnd.n2366 585
R2770 gnd.n4354 gnd.n4353 585
R2771 gnd.n4355 gnd.n4354 585
R2772 gnd.n2376 gnd.n2374 585
R2773 gnd.n4318 gnd.n2374 585
R2774 gnd.n4346 gnd.n4345 585
R2775 gnd.n4345 gnd.n4344 585
R2776 gnd.n1133 gnd.n1132 585
R2777 gnd.n4324 gnd.n1133 585
R2778 gnd.n6010 gnd.n6009 585
R2779 gnd.n6009 gnd.n6008 585
R2780 gnd.n6011 gnd.n1127 585
R2781 gnd.n4330 gnd.n1127 585
R2782 gnd.n6013 gnd.n6012 585
R2783 gnd.n6014 gnd.n6013 585
R2784 gnd.n1128 gnd.n1126 585
R2785 gnd.n1126 gnd.n1112 585
R2786 gnd.n4265 gnd.n1113 585
R2787 gnd.n6020 gnd.n1113 585
R2788 gnd.n4267 gnd.n4266 585
R2789 gnd.n4266 gnd.n1109 585
R2790 gnd.n4268 gnd.n2404 585
R2791 gnd.n4281 gnd.n2404 585
R2792 gnd.n4269 gnd.n2413 585
R2793 gnd.n2413 gnd.n2402 585
R2794 gnd.n4271 gnd.n4270 585
R2795 gnd.n4272 gnd.n4271 585
R2796 gnd.n2414 gnd.n2412 585
R2797 gnd.n2420 gnd.n2412 585
R2798 gnd.n4256 gnd.n4255 585
R2799 gnd.n4255 gnd.n4254 585
R2800 gnd.n2417 gnd.n2416 585
R2801 gnd.n2429 gnd.n2417 585
R2802 gnd.n4245 gnd.n4244 585
R2803 gnd.n4246 gnd.n4245 585
R2804 gnd.n2431 gnd.n2430 585
R2805 gnd.n2430 gnd.n2426 585
R2806 gnd.n4240 gnd.n4239 585
R2807 gnd.n4239 gnd.n4238 585
R2808 gnd.n2434 gnd.n2433 585
R2809 gnd.n2435 gnd.n2434 585
R2810 gnd.n4229 gnd.n4228 585
R2811 gnd.n4230 gnd.n4229 585
R2812 gnd.n2447 gnd.n2446 585
R2813 gnd.n2446 gnd.n2443 585
R2814 gnd.n4224 gnd.n4223 585
R2815 gnd.n4223 gnd.n4222 585
R2816 gnd.n2450 gnd.n2449 585
R2817 gnd.n4096 gnd.n2450 585
R2818 gnd.n4213 gnd.n4212 585
R2819 gnd.n4214 gnd.n4213 585
R2820 gnd.n4209 gnd.n4097 585
R2821 gnd.n4208 gnd.n4207 585
R2822 gnd.n4205 gnd.n4099 585
R2823 gnd.n4203 gnd.n4202 585
R2824 gnd.n4201 gnd.n4100 585
R2825 gnd.n4200 gnd.n4199 585
R2826 gnd.n4197 gnd.n4105 585
R2827 gnd.n4195 gnd.n4194 585
R2828 gnd.n4193 gnd.n4106 585
R2829 gnd.n4192 gnd.n4191 585
R2830 gnd.n4189 gnd.n4111 585
R2831 gnd.n4187 gnd.n4186 585
R2832 gnd.n4185 gnd.n4112 585
R2833 gnd.n4184 gnd.n4183 585
R2834 gnd.n4181 gnd.n4117 585
R2835 gnd.n4179 gnd.n4178 585
R2836 gnd.n4177 gnd.n4118 585
R2837 gnd.n4171 gnd.n4123 585
R2838 gnd.n4173 gnd.n4172 585
R2839 gnd.n4172 gnd.n3920 585
R2840 gnd.n4565 gnd.n4564 585
R2841 gnd.n4566 gnd.n2261 585
R2842 gnd.n4567 gnd.n2257 585
R2843 gnd.n2255 gnd.n2249 585
R2844 gnd.n4574 gnd.n2248 585
R2845 gnd.n4575 gnd.n2246 585
R2846 gnd.n2245 gnd.n2238 585
R2847 gnd.n4582 gnd.n2237 585
R2848 gnd.n4583 gnd.n2236 585
R2849 gnd.n2234 gnd.n2228 585
R2850 gnd.n4590 gnd.n2227 585
R2851 gnd.n4591 gnd.n2225 585
R2852 gnd.n2224 gnd.n2217 585
R2853 gnd.n4598 gnd.n2216 585
R2854 gnd.n4599 gnd.n2215 585
R2855 gnd.n2213 gnd.n2205 585
R2856 gnd.n4606 gnd.n2204 585
R2857 gnd.n4607 gnd.n2202 585
R2858 gnd.n4608 gnd.n1267 585
R2859 gnd.n1276 gnd.n1267 585
R2860 gnd.n1345 gnd.n1270 585
R2861 gnd.n5933 gnd.n1270 585
R2862 gnd.n5855 gnd.n5854 585
R2863 gnd.n5856 gnd.n5855 585
R2864 gnd.n1344 gnd.n1260 585
R2865 gnd.n5939 gnd.n1260 585
R2866 gnd.n4514 gnd.n4512 585
R2867 gnd.n4512 gnd.n4511 585
R2868 gnd.n4515 gnd.n1249 585
R2869 gnd.n5945 gnd.n1249 585
R2870 gnd.n4516 gnd.n2305 585
R2871 gnd.n4502 gnd.n2305 585
R2872 gnd.n2302 gnd.n1238 585
R2873 gnd.n5951 gnd.n1238 585
R2874 gnd.n4521 gnd.n4520 585
R2875 gnd.n4522 gnd.n4521 585
R2876 gnd.n2301 gnd.n1228 585
R2877 gnd.n5957 gnd.n1228 585
R2878 gnd.n4493 gnd.n4492 585
R2879 gnd.n4494 gnd.n4493 585
R2880 gnd.n2311 gnd.n1217 585
R2881 gnd.n5963 gnd.n1217 585
R2882 gnd.n4488 gnd.n4487 585
R2883 gnd.n4487 gnd.n4486 585
R2884 gnd.n2313 gnd.n1207 585
R2885 gnd.n5969 gnd.n1207 585
R2886 gnd.n4477 gnd.n4476 585
R2887 gnd.n4478 gnd.n4477 585
R2888 gnd.n2318 gnd.n1196 585
R2889 gnd.n5975 gnd.n1196 585
R2890 gnd.n4472 gnd.n4471 585
R2891 gnd.n4471 gnd.n4470 585
R2892 gnd.n2320 gnd.n1186 585
R2893 gnd.n5981 gnd.n1186 585
R2894 gnd.n4418 gnd.n4417 585
R2895 gnd.n4417 gnd.n4416 585
R2896 gnd.n2342 gnd.n1175 585
R2897 gnd.n5987 gnd.n1175 585
R2898 gnd.n4422 gnd.n2341 585
R2899 gnd.n4404 gnd.n2341 585
R2900 gnd.n4423 gnd.n1166 585
R2901 gnd.n5993 gnd.n1166 585
R2902 gnd.n4424 gnd.n2340 585
R2903 gnd.n4399 gnd.n2340 585
R2904 gnd.n2337 gnd.n1154 585
R2905 gnd.n5999 gnd.n1154 585
R2906 gnd.n4429 gnd.n4428 585
R2907 gnd.n4430 gnd.n4429 585
R2908 gnd.n2336 gnd.n2335 585
R2909 gnd.n4392 gnd.n2335 585
R2910 gnd.n4307 gnd.n2352 585
R2911 gnd.n4387 gnd.n2352 585
R2912 gnd.n4311 gnd.n2361 585
R2913 gnd.n4374 gnd.n2361 585
R2914 gnd.n4312 gnd.n2367 585
R2915 gnd.n4362 gnd.n2367 585
R2916 gnd.n4314 gnd.n4313 585
R2917 gnd.n4313 gnd.n2366 585
R2918 gnd.n4315 gnd.n2372 585
R2919 gnd.n4355 gnd.n2372 585
R2920 gnd.n4317 gnd.n4316 585
R2921 gnd.n4318 gnd.n4317 585
R2922 gnd.n2395 gnd.n2380 585
R2923 gnd.n4344 gnd.n2380 585
R2924 gnd.n4326 gnd.n4325 585
R2925 gnd.n4325 gnd.n4324 585
R2926 gnd.n4327 gnd.n1135 585
R2927 gnd.n6008 gnd.n1135 585
R2928 gnd.n4329 gnd.n4328 585
R2929 gnd.n4330 gnd.n4329 585
R2930 gnd.n2391 gnd.n1124 585
R2931 gnd.n6014 gnd.n1124 585
R2932 gnd.n4144 gnd.n4143 585
R2933 gnd.n4143 gnd.n1112 585
R2934 gnd.n4145 gnd.n1111 585
R2935 gnd.n6020 gnd.n1111 585
R2936 gnd.n4147 gnd.n4146 585
R2937 gnd.n4146 gnd.n1109 585
R2938 gnd.n4148 gnd.n2403 585
R2939 gnd.n4281 gnd.n2403 585
R2940 gnd.n4150 gnd.n4149 585
R2941 gnd.n4149 gnd.n2402 585
R2942 gnd.n4151 gnd.n2411 585
R2943 gnd.n4272 gnd.n2411 585
R2944 gnd.n4153 gnd.n4152 585
R2945 gnd.n4152 gnd.n2420 585
R2946 gnd.n4154 gnd.n2419 585
R2947 gnd.n4254 gnd.n2419 585
R2948 gnd.n4156 gnd.n4155 585
R2949 gnd.n4155 gnd.n2429 585
R2950 gnd.n4157 gnd.n2428 585
R2951 gnd.n4246 gnd.n2428 585
R2952 gnd.n4159 gnd.n4158 585
R2953 gnd.n4158 gnd.n2426 585
R2954 gnd.n4160 gnd.n2437 585
R2955 gnd.n4238 gnd.n2437 585
R2956 gnd.n4162 gnd.n4161 585
R2957 gnd.n4161 gnd.n2435 585
R2958 gnd.n4163 gnd.n2445 585
R2959 gnd.n4230 gnd.n2445 585
R2960 gnd.n4165 gnd.n4164 585
R2961 gnd.n4164 gnd.n2443 585
R2962 gnd.n4166 gnd.n2452 585
R2963 gnd.n4222 gnd.n2452 585
R2964 gnd.n4167 gnd.n4125 585
R2965 gnd.n4125 gnd.n4096 585
R2966 gnd.n4168 gnd.n3922 585
R2967 gnd.n4214 gnd.n3922 585
R2968 gnd.n182 gnd.n103 585
R2969 gnd.n7327 gnd.n103 585
R2970 gnd.n7247 gnd.n7246 585
R2971 gnd.n7248 gnd.n7247 585
R2972 gnd.n181 gnd.n180 585
R2973 gnd.n189 gnd.n180 585
R2974 gnd.n7174 gnd.n7173 585
R2975 gnd.n7173 gnd.n7172 585
R2976 gnd.n185 gnd.n184 585
R2977 gnd.n186 gnd.n185 585
R2978 gnd.n7161 gnd.n7160 585
R2979 gnd.n7162 gnd.n7161 585
R2980 gnd.n199 gnd.n198 585
R2981 gnd.n198 gnd.n196 585
R2982 gnd.n7156 gnd.n7155 585
R2983 gnd.n7155 gnd.n7154 585
R2984 gnd.n202 gnd.n201 585
R2985 gnd.n203 gnd.n202 585
R2986 gnd.n7145 gnd.n7144 585
R2987 gnd.n7146 gnd.n7145 585
R2988 gnd.n213 gnd.n212 585
R2989 gnd.n219 gnd.n212 585
R2990 gnd.n7140 gnd.n7139 585
R2991 gnd.n7139 gnd.n7138 585
R2992 gnd.n216 gnd.n215 585
R2993 gnd.n227 gnd.n216 585
R2994 gnd.n7129 gnd.n7128 585
R2995 gnd.n7130 gnd.n7129 585
R2996 gnd.n229 gnd.n228 585
R2997 gnd.n228 gnd.n225 585
R2998 gnd.n7124 gnd.n7123 585
R2999 gnd.n7123 gnd.n7122 585
R3000 gnd.n232 gnd.n231 585
R3001 gnd.n243 gnd.n232 585
R3002 gnd.n7113 gnd.n7112 585
R3003 gnd.n7114 gnd.n7113 585
R3004 gnd.n245 gnd.n244 585
R3005 gnd.n545 gnd.n244 585
R3006 gnd.n7108 gnd.n7107 585
R3007 gnd.n7107 gnd.n7106 585
R3008 gnd.n248 gnd.n247 585
R3009 gnd.n549 gnd.n248 585
R3010 gnd.n7097 gnd.n7096 585
R3011 gnd.n7098 gnd.n7097 585
R3012 gnd.n262 gnd.n261 585
R3013 gnd.n6837 gnd.n261 585
R3014 gnd.n7092 gnd.n7091 585
R3015 gnd.n7091 gnd.n7090 585
R3016 gnd.n265 gnd.n264 585
R3017 gnd.n6841 gnd.n265 585
R3018 gnd.n7082 gnd.n7081 585
R3019 gnd.n7083 gnd.n7082 585
R3020 gnd.n276 gnd.n275 585
R3021 gnd.n6845 gnd.n275 585
R3022 gnd.n7076 gnd.n7075 585
R3023 gnd.n7075 gnd.n7074 585
R3024 gnd.n280 gnd.n279 585
R3025 gnd.n6851 gnd.n280 585
R3026 gnd.n7065 gnd.n7064 585
R3027 gnd.n7066 gnd.n7065 585
R3028 gnd.n293 gnd.n292 585
R3029 gnd.n5554 gnd.n292 585
R3030 gnd.n7060 gnd.n7059 585
R3031 gnd.n7059 gnd.n7058 585
R3032 gnd.n296 gnd.n295 585
R3033 gnd.n5533 gnd.n296 585
R3034 gnd.n313 gnd.n311 585
R3035 gnd.n5576 gnd.n311 585
R3036 gnd.n7047 gnd.n7046 585
R3037 gnd.n7048 gnd.n7047 585
R3038 gnd.n312 gnd.n310 585
R3039 gnd.n5582 gnd.n310 585
R3040 gnd.n7041 gnd.n7040 585
R3041 gnd.n7040 gnd.n7039 585
R3042 gnd.n316 gnd.n315 585
R3043 gnd.n5522 gnd.n316 585
R3044 gnd.n7030 gnd.n7029 585
R3045 gnd.n7031 gnd.n7030 585
R3046 gnd.n330 gnd.n329 585
R3047 gnd.n5518 gnd.n329 585
R3048 gnd.n7025 gnd.n7024 585
R3049 gnd.n7024 gnd.n7023 585
R3050 gnd.n333 gnd.n332 585
R3051 gnd.n5512 gnd.n333 585
R3052 gnd.n7014 gnd.n7013 585
R3053 gnd.n7015 gnd.n7014 585
R3054 gnd.n348 gnd.n347 585
R3055 gnd.n5598 gnd.n347 585
R3056 gnd.n7009 gnd.n7008 585
R3057 gnd.n7008 gnd.n7007 585
R3058 gnd.n351 gnd.n350 585
R3059 gnd.n5602 gnd.n351 585
R3060 gnd.n6998 gnd.n6997 585
R3061 gnd.n6999 gnd.n6998 585
R3062 gnd.n365 gnd.n364 585
R3063 gnd.n5606 gnd.n364 585
R3064 gnd.n6993 gnd.n6992 585
R3065 gnd.n6992 gnd.n6991 585
R3066 gnd.n368 gnd.n367 585
R3067 gnd.n5610 gnd.n368 585
R3068 gnd.n6982 gnd.n6981 585
R3069 gnd.n6983 gnd.n6982 585
R3070 gnd.n383 gnd.n382 585
R3071 gnd.n5616 gnd.n382 585
R3072 gnd.n6977 gnd.n6976 585
R3073 gnd.n6976 gnd.n6975 585
R3074 gnd.n386 gnd.n385 585
R3075 gnd.n6894 gnd.n386 585
R3076 gnd.n5702 gnd.n5701 585
R3077 gnd.n5700 gnd.n1478 585
R3078 gnd.n5699 gnd.n1479 585
R3079 gnd.n1488 gnd.n1480 585
R3080 gnd.n5692 gnd.n1489 585
R3081 gnd.n5691 gnd.n1490 585
R3082 gnd.n1492 gnd.n1491 585
R3083 gnd.n5684 gnd.n1498 585
R3084 gnd.n5683 gnd.n1499 585
R3085 gnd.n1506 gnd.n1500 585
R3086 gnd.n5676 gnd.n1507 585
R3087 gnd.n5675 gnd.n1508 585
R3088 gnd.n1510 gnd.n1509 585
R3089 gnd.n5668 gnd.n1516 585
R3090 gnd.n5667 gnd.n1517 585
R3091 gnd.n1524 gnd.n1518 585
R3092 gnd.n5660 gnd.n1525 585
R3093 gnd.n5659 gnd.n5656 585
R3094 gnd.n1526 gnd.n423 585
R3095 gnd.n6966 gnd.n423 585
R3096 gnd.n7216 gnd.n99 585
R3097 gnd.n7217 gnd.n7214 585
R3098 gnd.n7218 gnd.n7210 585
R3099 gnd.n7208 gnd.n7206 585
R3100 gnd.n7222 gnd.n7205 585
R3101 gnd.n7223 gnd.n7203 585
R3102 gnd.n7224 gnd.n7202 585
R3103 gnd.n7200 gnd.n7198 585
R3104 gnd.n7228 gnd.n7197 585
R3105 gnd.n7229 gnd.n7195 585
R3106 gnd.n7230 gnd.n7194 585
R3107 gnd.n7192 gnd.n7190 585
R3108 gnd.n7234 gnd.n7189 585
R3109 gnd.n7235 gnd.n7187 585
R3110 gnd.n7236 gnd.n7186 585
R3111 gnd.n7184 gnd.n7182 585
R3112 gnd.n7240 gnd.n7181 585
R3113 gnd.n7241 gnd.n7179 585
R3114 gnd.n7242 gnd.n7178 585
R3115 gnd.n7178 gnd.n102 585
R3116 gnd.n7329 gnd.n7328 585
R3117 gnd.n7328 gnd.n7327 585
R3118 gnd.n7330 gnd.n97 585
R3119 gnd.n7248 gnd.n97 585
R3120 gnd.n7331 gnd.n96 585
R3121 gnd.n189 gnd.n96 585
R3122 gnd.n188 gnd.n94 585
R3123 gnd.n7172 gnd.n188 585
R3124 gnd.n7335 gnd.n93 585
R3125 gnd.n186 gnd.n93 585
R3126 gnd.n7336 gnd.n92 585
R3127 gnd.n7162 gnd.n92 585
R3128 gnd.n7337 gnd.n91 585
R3129 gnd.n196 gnd.n91 585
R3130 gnd.n205 gnd.n89 585
R3131 gnd.n7154 gnd.n205 585
R3132 gnd.n7341 gnd.n88 585
R3133 gnd.n203 gnd.n88 585
R3134 gnd.n7342 gnd.n87 585
R3135 gnd.n7146 gnd.n87 585
R3136 gnd.n7343 gnd.n86 585
R3137 gnd.n219 gnd.n86 585
R3138 gnd.n218 gnd.n84 585
R3139 gnd.n7138 gnd.n218 585
R3140 gnd.n7347 gnd.n83 585
R3141 gnd.n227 gnd.n83 585
R3142 gnd.n7348 gnd.n82 585
R3143 gnd.n7130 gnd.n82 585
R3144 gnd.n7349 gnd.n81 585
R3145 gnd.n225 gnd.n81 585
R3146 gnd.n235 gnd.n79 585
R3147 gnd.n7122 gnd.n235 585
R3148 gnd.n7353 gnd.n78 585
R3149 gnd.n243 gnd.n78 585
R3150 gnd.n7354 gnd.n77 585
R3151 gnd.n7114 gnd.n77 585
R3152 gnd.n7355 gnd.n76 585
R3153 gnd.n545 gnd.n76 585
R3154 gnd.n251 gnd.n74 585
R3155 gnd.n7106 gnd.n251 585
R3156 gnd.n7359 gnd.n73 585
R3157 gnd.n549 gnd.n73 585
R3158 gnd.n7360 gnd.n72 585
R3159 gnd.n7098 gnd.n72 585
R3160 gnd.n7361 gnd.n71 585
R3161 gnd.n6837 gnd.n71 585
R3162 gnd.n268 gnd.n69 585
R3163 gnd.n7090 gnd.n268 585
R3164 gnd.n7365 gnd.n68 585
R3165 gnd.n6841 gnd.n68 585
R3166 gnd.n7366 gnd.n67 585
R3167 gnd.n7083 gnd.n67 585
R3168 gnd.n7367 gnd.n66 585
R3169 gnd.n6845 gnd.n66 585
R3170 gnd.n283 gnd.n65 585
R3171 gnd.n7074 gnd.n283 585
R3172 gnd.n6853 gnd.n6852 585
R3173 gnd.n6852 gnd.n6851 585
R3174 gnd.n6856 gnd.n290 585
R3175 gnd.n7066 gnd.n290 585
R3176 gnd.n6857 gnd.n494 585
R3177 gnd.n5554 gnd.n494 585
R3178 gnd.n6858 gnd.n299 585
R3179 gnd.n7058 gnd.n299 585
R3180 gnd.n5532 gnd.n492 585
R3181 gnd.n5533 gnd.n5532 585
R3182 gnd.n6862 gnd.n491 585
R3183 gnd.n5576 gnd.n491 585
R3184 gnd.n6863 gnd.n308 585
R3185 gnd.n7048 gnd.n308 585
R3186 gnd.n6864 gnd.n490 585
R3187 gnd.n5582 gnd.n490 585
R3188 gnd.n488 gnd.n319 585
R3189 gnd.n7039 gnd.n319 585
R3190 gnd.n6868 gnd.n487 585
R3191 gnd.n5522 gnd.n487 585
R3192 gnd.n6869 gnd.n327 585
R3193 gnd.n7031 gnd.n327 585
R3194 gnd.n6870 gnd.n486 585
R3195 gnd.n5518 gnd.n486 585
R3196 gnd.n484 gnd.n336 585
R3197 gnd.n7023 gnd.n336 585
R3198 gnd.n6874 gnd.n483 585
R3199 gnd.n5512 gnd.n483 585
R3200 gnd.n6875 gnd.n345 585
R3201 gnd.n7015 gnd.n345 585
R3202 gnd.n6876 gnd.n482 585
R3203 gnd.n5598 gnd.n482 585
R3204 gnd.n480 gnd.n354 585
R3205 gnd.n7007 gnd.n354 585
R3206 gnd.n6880 gnd.n479 585
R3207 gnd.n5602 gnd.n479 585
R3208 gnd.n6881 gnd.n362 585
R3209 gnd.n6999 gnd.n362 585
R3210 gnd.n6882 gnd.n478 585
R3211 gnd.n5606 gnd.n478 585
R3212 gnd.n476 gnd.n371 585
R3213 gnd.n6991 gnd.n371 585
R3214 gnd.n6886 gnd.n475 585
R3215 gnd.n5610 gnd.n475 585
R3216 gnd.n6887 gnd.n380 585
R3217 gnd.n6983 gnd.n380 585
R3218 gnd.n6888 gnd.n474 585
R3219 gnd.n5616 gnd.n474 585
R3220 gnd.n471 gnd.n389 585
R3221 gnd.n6975 gnd.n389 585
R3222 gnd.n6893 gnd.n6892 585
R3223 gnd.n6894 gnd.n6893 585
R3224 gnd.n3827 gnd.n3826 585
R3225 gnd.n3828 gnd.n3827 585
R3226 gnd.n2533 gnd.n2532 585
R3227 gnd.n2539 gnd.n2532 585
R3228 gnd.n3802 gnd.n2551 585
R3229 gnd.n2551 gnd.n2538 585
R3230 gnd.n3804 gnd.n3803 585
R3231 gnd.n3805 gnd.n3804 585
R3232 gnd.n2552 gnd.n2550 585
R3233 gnd.n2550 gnd.n2546 585
R3234 gnd.n3536 gnd.n3535 585
R3235 gnd.n3535 gnd.n3534 585
R3236 gnd.n2557 gnd.n2556 585
R3237 gnd.n3505 gnd.n2557 585
R3238 gnd.n3525 gnd.n3524 585
R3239 gnd.n3524 gnd.n3523 585
R3240 gnd.n2564 gnd.n2563 585
R3241 gnd.n3511 gnd.n2564 585
R3242 gnd.n3481 gnd.n2585 585
R3243 gnd.n2585 gnd.n2584 585
R3244 gnd.n3483 gnd.n3482 585
R3245 gnd.n3484 gnd.n3483 585
R3246 gnd.n2586 gnd.n2583 585
R3247 gnd.n2594 gnd.n2583 585
R3248 gnd.n3459 gnd.n2606 585
R3249 gnd.n2606 gnd.n2593 585
R3250 gnd.n3461 gnd.n3460 585
R3251 gnd.n3462 gnd.n3461 585
R3252 gnd.n2607 gnd.n2605 585
R3253 gnd.n2605 gnd.n2601 585
R3254 gnd.n3447 gnd.n3446 585
R3255 gnd.n3446 gnd.n3445 585
R3256 gnd.n2612 gnd.n2611 585
R3257 gnd.n2622 gnd.n2612 585
R3258 gnd.n3436 gnd.n3435 585
R3259 gnd.n3435 gnd.n3434 585
R3260 gnd.n2619 gnd.n2618 585
R3261 gnd.n3422 gnd.n2619 585
R3262 gnd.n3396 gnd.n2640 585
R3263 gnd.n2640 gnd.n2629 585
R3264 gnd.n3398 gnd.n3397 585
R3265 gnd.n3399 gnd.n3398 585
R3266 gnd.n2641 gnd.n2639 585
R3267 gnd.n2649 gnd.n2639 585
R3268 gnd.n3374 gnd.n2661 585
R3269 gnd.n2661 gnd.n2648 585
R3270 gnd.n3376 gnd.n3375 585
R3271 gnd.n3377 gnd.n3376 585
R3272 gnd.n2662 gnd.n2660 585
R3273 gnd.n2660 gnd.n2656 585
R3274 gnd.n3362 gnd.n3361 585
R3275 gnd.n3361 gnd.n3360 585
R3276 gnd.n2667 gnd.n2666 585
R3277 gnd.n2676 gnd.n2667 585
R3278 gnd.n3351 gnd.n3350 585
R3279 gnd.n3350 gnd.n3349 585
R3280 gnd.n2674 gnd.n2673 585
R3281 gnd.n3337 gnd.n2674 585
R3282 gnd.n2775 gnd.n2774 585
R3283 gnd.n2775 gnd.n2683 585
R3284 gnd.n3294 gnd.n3293 585
R3285 gnd.n3293 gnd.n3292 585
R3286 gnd.n3295 gnd.n2769 585
R3287 gnd.n2780 gnd.n2769 585
R3288 gnd.n3297 gnd.n3296 585
R3289 gnd.n3298 gnd.n3297 585
R3290 gnd.n2770 gnd.n2768 585
R3291 gnd.n2793 gnd.n2768 585
R3292 gnd.n2753 gnd.n2752 585
R3293 gnd.n2756 gnd.n2753 585
R3294 gnd.n3308 gnd.n3307 585
R3295 gnd.n3307 gnd.n3306 585
R3296 gnd.n3309 gnd.n2747 585
R3297 gnd.n3268 gnd.n2747 585
R3298 gnd.n3311 gnd.n3310 585
R3299 gnd.n3312 gnd.n3311 585
R3300 gnd.n2748 gnd.n2746 585
R3301 gnd.n2807 gnd.n2746 585
R3302 gnd.n3260 gnd.n3259 585
R3303 gnd.n3259 gnd.n3258 585
R3304 gnd.n2804 gnd.n2803 585
R3305 gnd.n3242 gnd.n2804 585
R3306 gnd.n3229 gnd.n2823 585
R3307 gnd.n2823 gnd.n2822 585
R3308 gnd.n3231 gnd.n3230 585
R3309 gnd.n3232 gnd.n3231 585
R3310 gnd.n2824 gnd.n2821 585
R3311 gnd.n2830 gnd.n2821 585
R3312 gnd.n3210 gnd.n3209 585
R3313 gnd.n3211 gnd.n3210 585
R3314 gnd.n2841 gnd.n2840 585
R3315 gnd.n2840 gnd.n2836 585
R3316 gnd.n3200 gnd.n3199 585
R3317 gnd.n3201 gnd.n3200 585
R3318 gnd.n2851 gnd.n2850 585
R3319 gnd.n2856 gnd.n2850 585
R3320 gnd.n3178 gnd.n2869 585
R3321 gnd.n2869 gnd.n2855 585
R3322 gnd.n3180 gnd.n3179 585
R3323 gnd.n3181 gnd.n3180 585
R3324 gnd.n2870 gnd.n2868 585
R3325 gnd.n2868 gnd.n2864 585
R3326 gnd.n3169 gnd.n3168 585
R3327 gnd.n3170 gnd.n3169 585
R3328 gnd.n2877 gnd.n2876 585
R3329 gnd.n2881 gnd.n2876 585
R3330 gnd.n3146 gnd.n2898 585
R3331 gnd.n2898 gnd.n2880 585
R3332 gnd.n3148 gnd.n3147 585
R3333 gnd.n3149 gnd.n3148 585
R3334 gnd.n2899 gnd.n2897 585
R3335 gnd.n2897 gnd.n2888 585
R3336 gnd.n3141 gnd.n3140 585
R3337 gnd.n3140 gnd.n3139 585
R3338 gnd.n2946 gnd.n2945 585
R3339 gnd.n2947 gnd.n2946 585
R3340 gnd.n3100 gnd.n3099 585
R3341 gnd.n3101 gnd.n3100 585
R3342 gnd.n2956 gnd.n2955 585
R3343 gnd.n2955 gnd.n2954 585
R3344 gnd.n3095 gnd.n3094 585
R3345 gnd.n3094 gnd.n3093 585
R3346 gnd.n2959 gnd.n2958 585
R3347 gnd.n2960 gnd.n2959 585
R3348 gnd.n3084 gnd.n3083 585
R3349 gnd.n3085 gnd.n3084 585
R3350 gnd.n2967 gnd.n2966 585
R3351 gnd.n3076 gnd.n2966 585
R3352 gnd.n3079 gnd.n3078 585
R3353 gnd.n3078 gnd.n3077 585
R3354 gnd.n2970 gnd.n2969 585
R3355 gnd.n2971 gnd.n2970 585
R3356 gnd.n3065 gnd.n3064 585
R3357 gnd.n3063 gnd.n2989 585
R3358 gnd.n3062 gnd.n2988 585
R3359 gnd.n3067 gnd.n2988 585
R3360 gnd.n3061 gnd.n3060 585
R3361 gnd.n3059 gnd.n3058 585
R3362 gnd.n3057 gnd.n3056 585
R3363 gnd.n3055 gnd.n3054 585
R3364 gnd.n3053 gnd.n3052 585
R3365 gnd.n3051 gnd.n3050 585
R3366 gnd.n3049 gnd.n3048 585
R3367 gnd.n3047 gnd.n3046 585
R3368 gnd.n3045 gnd.n3044 585
R3369 gnd.n3043 gnd.n3042 585
R3370 gnd.n3041 gnd.n3040 585
R3371 gnd.n3039 gnd.n3038 585
R3372 gnd.n3037 gnd.n3036 585
R3373 gnd.n3035 gnd.n3034 585
R3374 gnd.n3033 gnd.n3032 585
R3375 gnd.n3031 gnd.n3030 585
R3376 gnd.n3029 gnd.n3028 585
R3377 gnd.n3027 gnd.n3026 585
R3378 gnd.n3025 gnd.n3024 585
R3379 gnd.n3023 gnd.n3022 585
R3380 gnd.n3021 gnd.n3020 585
R3381 gnd.n3019 gnd.n3018 585
R3382 gnd.n2976 gnd.n2975 585
R3383 gnd.n3070 gnd.n3069 585
R3384 gnd.n3831 gnd.n3830 585
R3385 gnd.n3833 gnd.n3832 585
R3386 gnd.n3835 gnd.n3834 585
R3387 gnd.n3837 gnd.n3836 585
R3388 gnd.n3839 gnd.n3838 585
R3389 gnd.n3841 gnd.n3840 585
R3390 gnd.n3843 gnd.n3842 585
R3391 gnd.n3845 gnd.n3844 585
R3392 gnd.n3847 gnd.n3846 585
R3393 gnd.n3849 gnd.n3848 585
R3394 gnd.n3851 gnd.n3850 585
R3395 gnd.n3853 gnd.n3852 585
R3396 gnd.n3855 gnd.n3854 585
R3397 gnd.n3857 gnd.n3856 585
R3398 gnd.n3859 gnd.n3858 585
R3399 gnd.n3861 gnd.n3860 585
R3400 gnd.n3863 gnd.n3862 585
R3401 gnd.n3865 gnd.n3864 585
R3402 gnd.n3867 gnd.n3866 585
R3403 gnd.n3869 gnd.n3868 585
R3404 gnd.n3871 gnd.n3870 585
R3405 gnd.n3873 gnd.n3872 585
R3406 gnd.n3875 gnd.n3874 585
R3407 gnd.n3877 gnd.n3876 585
R3408 gnd.n3879 gnd.n3878 585
R3409 gnd.n3880 gnd.n2500 585
R3410 gnd.n3881 gnd.n2458 585
R3411 gnd.n3919 gnd.n2458 585
R3412 gnd.n3829 gnd.n2530 585
R3413 gnd.n3829 gnd.n3828 585
R3414 gnd.n3498 gnd.n2529 585
R3415 gnd.n2539 gnd.n2529 585
R3416 gnd.n3500 gnd.n3499 585
R3417 gnd.n3499 gnd.n2538 585
R3418 gnd.n3501 gnd.n2548 585
R3419 gnd.n3805 gnd.n2548 585
R3420 gnd.n3503 gnd.n3502 585
R3421 gnd.n3502 gnd.n2546 585
R3422 gnd.n3504 gnd.n2559 585
R3423 gnd.n3534 gnd.n2559 585
R3424 gnd.n3507 gnd.n3506 585
R3425 gnd.n3506 gnd.n3505 585
R3426 gnd.n3508 gnd.n2566 585
R3427 gnd.n3523 gnd.n2566 585
R3428 gnd.n3510 gnd.n3509 585
R3429 gnd.n3511 gnd.n3510 585
R3430 gnd.n2577 gnd.n2576 585
R3431 gnd.n2584 gnd.n2576 585
R3432 gnd.n3486 gnd.n3485 585
R3433 gnd.n3485 gnd.n3484 585
R3434 gnd.n2580 gnd.n2579 585
R3435 gnd.n2594 gnd.n2580 585
R3436 gnd.n3412 gnd.n3411 585
R3437 gnd.n3411 gnd.n2593 585
R3438 gnd.n3413 gnd.n2603 585
R3439 gnd.n3462 gnd.n2603 585
R3440 gnd.n3415 gnd.n3414 585
R3441 gnd.n3414 gnd.n2601 585
R3442 gnd.n3416 gnd.n2614 585
R3443 gnd.n3445 gnd.n2614 585
R3444 gnd.n3418 gnd.n3417 585
R3445 gnd.n3417 gnd.n2622 585
R3446 gnd.n3419 gnd.n2621 585
R3447 gnd.n3434 gnd.n2621 585
R3448 gnd.n3421 gnd.n3420 585
R3449 gnd.n3422 gnd.n3421 585
R3450 gnd.n2633 gnd.n2632 585
R3451 gnd.n2632 gnd.n2629 585
R3452 gnd.n3401 gnd.n3400 585
R3453 gnd.n3400 gnd.n3399 585
R3454 gnd.n2636 gnd.n2635 585
R3455 gnd.n2649 gnd.n2636 585
R3456 gnd.n3325 gnd.n3324 585
R3457 gnd.n3324 gnd.n2648 585
R3458 gnd.n3326 gnd.n2658 585
R3459 gnd.n3377 gnd.n2658 585
R3460 gnd.n3328 gnd.n3327 585
R3461 gnd.n3327 gnd.n2656 585
R3462 gnd.n3329 gnd.n2669 585
R3463 gnd.n3360 gnd.n2669 585
R3464 gnd.n3331 gnd.n3330 585
R3465 gnd.n3330 gnd.n2676 585
R3466 gnd.n3332 gnd.n2675 585
R3467 gnd.n3349 gnd.n2675 585
R3468 gnd.n3334 gnd.n3333 585
R3469 gnd.n3337 gnd.n3334 585
R3470 gnd.n2686 gnd.n2685 585
R3471 gnd.n2685 gnd.n2683 585
R3472 gnd.n2777 gnd.n2776 585
R3473 gnd.n3292 gnd.n2776 585
R3474 gnd.n2779 gnd.n2778 585
R3475 gnd.n2780 gnd.n2779 585
R3476 gnd.n2790 gnd.n2766 585
R3477 gnd.n3298 gnd.n2766 585
R3478 gnd.n2792 gnd.n2791 585
R3479 gnd.n2793 gnd.n2792 585
R3480 gnd.n2789 gnd.n2788 585
R3481 gnd.n2789 gnd.n2756 585
R3482 gnd.n2787 gnd.n2754 585
R3483 gnd.n3306 gnd.n2754 585
R3484 gnd.n2743 gnd.n2741 585
R3485 gnd.n3268 gnd.n2743 585
R3486 gnd.n3314 gnd.n3313 585
R3487 gnd.n3313 gnd.n3312 585
R3488 gnd.n2742 gnd.n2740 585
R3489 gnd.n2807 gnd.n2742 585
R3490 gnd.n3239 gnd.n2806 585
R3491 gnd.n3258 gnd.n2806 585
R3492 gnd.n3241 gnd.n3240 585
R3493 gnd.n3242 gnd.n3241 585
R3494 gnd.n2816 gnd.n2815 585
R3495 gnd.n2822 gnd.n2815 585
R3496 gnd.n3234 gnd.n3233 585
R3497 gnd.n3233 gnd.n3232 585
R3498 gnd.n2819 gnd.n2818 585
R3499 gnd.n2830 gnd.n2819 585
R3500 gnd.n3119 gnd.n2838 585
R3501 gnd.n3211 gnd.n2838 585
R3502 gnd.n3121 gnd.n3120 585
R3503 gnd.n3120 gnd.n2836 585
R3504 gnd.n3122 gnd.n2849 585
R3505 gnd.n3201 gnd.n2849 585
R3506 gnd.n3124 gnd.n3123 585
R3507 gnd.n3124 gnd.n2856 585
R3508 gnd.n3126 gnd.n3125 585
R3509 gnd.n3125 gnd.n2855 585
R3510 gnd.n3127 gnd.n2866 585
R3511 gnd.n3181 gnd.n2866 585
R3512 gnd.n3129 gnd.n3128 585
R3513 gnd.n3128 gnd.n2864 585
R3514 gnd.n3130 gnd.n2875 585
R3515 gnd.n3170 gnd.n2875 585
R3516 gnd.n3132 gnd.n3131 585
R3517 gnd.n3132 gnd.n2881 585
R3518 gnd.n3134 gnd.n3133 585
R3519 gnd.n3133 gnd.n2880 585
R3520 gnd.n3135 gnd.n2896 585
R3521 gnd.n3149 gnd.n2896 585
R3522 gnd.n3136 gnd.n2949 585
R3523 gnd.n2949 gnd.n2888 585
R3524 gnd.n3138 gnd.n3137 585
R3525 gnd.n3139 gnd.n3138 585
R3526 gnd.n2950 gnd.n2948 585
R3527 gnd.n2948 gnd.n2947 585
R3528 gnd.n3103 gnd.n3102 585
R3529 gnd.n3102 gnd.n3101 585
R3530 gnd.n2953 gnd.n2952 585
R3531 gnd.n2954 gnd.n2953 585
R3532 gnd.n3092 gnd.n3091 585
R3533 gnd.n3093 gnd.n3092 585
R3534 gnd.n2962 gnd.n2961 585
R3535 gnd.n2961 gnd.n2960 585
R3536 gnd.n3087 gnd.n3086 585
R3537 gnd.n3086 gnd.n3085 585
R3538 gnd.n2965 gnd.n2964 585
R3539 gnd.n3076 gnd.n2965 585
R3540 gnd.n3075 gnd.n3074 585
R3541 gnd.n3077 gnd.n3075 585
R3542 gnd.n2973 gnd.n2972 585
R3543 gnd.n2972 gnd.n2971 585
R3544 gnd.n3814 gnd.n2480 585
R3545 gnd.n2480 gnd.n2457 585
R3546 gnd.n3815 gnd.n2541 585
R3547 gnd.n2541 gnd.n2531 585
R3548 gnd.n3817 gnd.n3816 585
R3549 gnd.n3818 gnd.n3817 585
R3550 gnd.n2542 gnd.n2540 585
R3551 gnd.n2549 gnd.n2540 585
R3552 gnd.n3808 gnd.n3807 585
R3553 gnd.n3807 gnd.n3806 585
R3554 gnd.n2545 gnd.n2544 585
R3555 gnd.n3533 gnd.n2545 585
R3556 gnd.n3519 gnd.n2568 585
R3557 gnd.n2568 gnd.n2558 585
R3558 gnd.n3521 gnd.n3520 585
R3559 gnd.n3522 gnd.n3521 585
R3560 gnd.n2569 gnd.n2567 585
R3561 gnd.n2567 gnd.n2565 585
R3562 gnd.n3514 gnd.n3513 585
R3563 gnd.n3513 gnd.n3512 585
R3564 gnd.n2572 gnd.n2571 585
R3565 gnd.n2582 gnd.n2572 585
R3566 gnd.n3470 gnd.n2596 585
R3567 gnd.n2596 gnd.n2581 585
R3568 gnd.n3472 gnd.n3471 585
R3569 gnd.n3473 gnd.n3472 585
R3570 gnd.n2597 gnd.n2595 585
R3571 gnd.n2604 gnd.n2595 585
R3572 gnd.n3465 gnd.n3464 585
R3573 gnd.n3464 gnd.n3463 585
R3574 gnd.n2600 gnd.n2599 585
R3575 gnd.n3444 gnd.n2600 585
R3576 gnd.n3430 gnd.n2624 585
R3577 gnd.n2624 gnd.n2613 585
R3578 gnd.n3432 gnd.n3431 585
R3579 gnd.n3433 gnd.n3432 585
R3580 gnd.n2625 gnd.n2623 585
R3581 gnd.n2623 gnd.n2620 585
R3582 gnd.n3425 gnd.n3424 585
R3583 gnd.n3424 gnd.n3423 585
R3584 gnd.n2628 gnd.n2627 585
R3585 gnd.n2638 gnd.n2628 585
R3586 gnd.n3385 gnd.n2651 585
R3587 gnd.n2651 gnd.n2637 585
R3588 gnd.n3387 gnd.n3386 585
R3589 gnd.n3388 gnd.n3387 585
R3590 gnd.n2652 gnd.n2650 585
R3591 gnd.n2659 gnd.n2650 585
R3592 gnd.n3380 gnd.n3379 585
R3593 gnd.n3379 gnd.n3378 585
R3594 gnd.n2655 gnd.n2654 585
R3595 gnd.n3359 gnd.n2655 585
R3596 gnd.n3345 gnd.n2678 585
R3597 gnd.n2678 gnd.n2668 585
R3598 gnd.n3347 gnd.n3346 585
R3599 gnd.n3348 gnd.n3347 585
R3600 gnd.n2679 gnd.n2677 585
R3601 gnd.n3336 gnd.n2677 585
R3602 gnd.n3340 gnd.n3339 585
R3603 gnd.n3339 gnd.n3338 585
R3604 gnd.n2682 gnd.n2681 585
R3605 gnd.n3291 gnd.n2682 585
R3606 gnd.n2784 gnd.n2783 585
R3607 gnd.n2785 gnd.n2784 585
R3608 gnd.n2764 gnd.n2763 585
R3609 gnd.n2767 gnd.n2764 585
R3610 gnd.n3301 gnd.n3300 585
R3611 gnd.n3300 gnd.n3299 585
R3612 gnd.n3302 gnd.n2758 585
R3613 gnd.n2794 gnd.n2758 585
R3614 gnd.n3304 gnd.n3303 585
R3615 gnd.n3305 gnd.n3304 585
R3616 gnd.n2759 gnd.n2757 585
R3617 gnd.n3269 gnd.n2757 585
R3618 gnd.n3253 gnd.n3252 585
R3619 gnd.n3252 gnd.n2745 585
R3620 gnd.n3254 gnd.n2809 585
R3621 gnd.n2809 gnd.n2744 585
R3622 gnd.n3256 gnd.n3255 585
R3623 gnd.n3257 gnd.n3256 585
R3624 gnd.n2810 gnd.n2808 585
R3625 gnd.n2808 gnd.n2805 585
R3626 gnd.n3245 gnd.n3244 585
R3627 gnd.n3244 gnd.n3243 585
R3628 gnd.n2813 gnd.n2812 585
R3629 gnd.n2820 gnd.n2813 585
R3630 gnd.n3219 gnd.n3218 585
R3631 gnd.n3220 gnd.n3219 585
R3632 gnd.n2832 gnd.n2831 585
R3633 gnd.n2839 gnd.n2831 585
R3634 gnd.n3214 gnd.n3213 585
R3635 gnd.n3213 gnd.n3212 585
R3636 gnd.n2835 gnd.n2834 585
R3637 gnd.n3202 gnd.n2835 585
R3638 gnd.n3189 gnd.n2859 585
R3639 gnd.n2859 gnd.n2858 585
R3640 gnd.n3191 gnd.n3190 585
R3641 gnd.n3192 gnd.n3191 585
R3642 gnd.n2860 gnd.n2857 585
R3643 gnd.n2867 gnd.n2857 585
R3644 gnd.n3184 gnd.n3183 585
R3645 gnd.n3183 gnd.n3182 585
R3646 gnd.n2863 gnd.n2862 585
R3647 gnd.n3171 gnd.n2863 585
R3648 gnd.n3158 gnd.n2884 585
R3649 gnd.n2884 gnd.n2883 585
R3650 gnd.n3160 gnd.n3159 585
R3651 gnd.n3161 gnd.n3160 585
R3652 gnd.n3154 gnd.n2882 585
R3653 gnd.n3153 gnd.n3152 585
R3654 gnd.n2887 gnd.n2886 585
R3655 gnd.n3150 gnd.n2887 585
R3656 gnd.n2909 gnd.n2908 585
R3657 gnd.n2912 gnd.n2911 585
R3658 gnd.n2910 gnd.n2905 585
R3659 gnd.n2917 gnd.n2916 585
R3660 gnd.n2919 gnd.n2918 585
R3661 gnd.n2922 gnd.n2921 585
R3662 gnd.n2920 gnd.n2903 585
R3663 gnd.n2927 gnd.n2926 585
R3664 gnd.n2929 gnd.n2928 585
R3665 gnd.n2932 gnd.n2931 585
R3666 gnd.n2930 gnd.n2901 585
R3667 gnd.n2937 gnd.n2936 585
R3668 gnd.n2941 gnd.n2938 585
R3669 gnd.n2942 gnd.n2879 585
R3670 gnd.n3820 gnd.n2495 585
R3671 gnd.n3887 gnd.n3886 585
R3672 gnd.n3889 gnd.n3888 585
R3673 gnd.n3891 gnd.n3890 585
R3674 gnd.n3893 gnd.n3892 585
R3675 gnd.n3895 gnd.n3894 585
R3676 gnd.n3897 gnd.n3896 585
R3677 gnd.n3899 gnd.n3898 585
R3678 gnd.n3901 gnd.n3900 585
R3679 gnd.n3903 gnd.n3902 585
R3680 gnd.n3905 gnd.n3904 585
R3681 gnd.n3907 gnd.n3906 585
R3682 gnd.n3909 gnd.n3908 585
R3683 gnd.n3912 gnd.n3911 585
R3684 gnd.n3910 gnd.n2483 585
R3685 gnd.n3916 gnd.n2481 585
R3686 gnd.n3918 gnd.n3917 585
R3687 gnd.n3919 gnd.n3918 585
R3688 gnd.n3821 gnd.n2536 585
R3689 gnd.n3821 gnd.n2457 585
R3690 gnd.n3823 gnd.n3822 585
R3691 gnd.n3822 gnd.n2531 585
R3692 gnd.n3819 gnd.n2535 585
R3693 gnd.n3819 gnd.n3818 585
R3694 gnd.n3798 gnd.n2537 585
R3695 gnd.n2549 gnd.n2537 585
R3696 gnd.n3797 gnd.n2547 585
R3697 gnd.n3806 gnd.n2547 585
R3698 gnd.n3532 gnd.n2554 585
R3699 gnd.n3533 gnd.n3532 585
R3700 gnd.n3531 gnd.n3530 585
R3701 gnd.n3531 gnd.n2558 585
R3702 gnd.n3529 gnd.n2560 585
R3703 gnd.n3522 gnd.n2560 585
R3704 gnd.n2574 gnd.n2561 585
R3705 gnd.n2574 gnd.n2565 585
R3706 gnd.n3478 gnd.n2575 585
R3707 gnd.n3512 gnd.n2575 585
R3708 gnd.n3477 gnd.n3476 585
R3709 gnd.n3476 gnd.n2582 585
R3710 gnd.n3475 gnd.n2590 585
R3711 gnd.n3475 gnd.n2581 585
R3712 gnd.n3474 gnd.n2592 585
R3713 gnd.n3474 gnd.n3473 585
R3714 gnd.n3453 gnd.n2591 585
R3715 gnd.n2604 gnd.n2591 585
R3716 gnd.n3452 gnd.n2602 585
R3717 gnd.n3463 gnd.n2602 585
R3718 gnd.n3443 gnd.n2609 585
R3719 gnd.n3444 gnd.n3443 585
R3720 gnd.n3442 gnd.n3441 585
R3721 gnd.n3442 gnd.n2613 585
R3722 gnd.n3440 gnd.n2615 585
R3723 gnd.n3433 gnd.n2615 585
R3724 gnd.n2630 gnd.n2616 585
R3725 gnd.n2630 gnd.n2620 585
R3726 gnd.n3393 gnd.n2631 585
R3727 gnd.n3423 gnd.n2631 585
R3728 gnd.n3392 gnd.n3391 585
R3729 gnd.n3391 gnd.n2638 585
R3730 gnd.n3390 gnd.n2645 585
R3731 gnd.n3390 gnd.n2637 585
R3732 gnd.n3389 gnd.n2647 585
R3733 gnd.n3389 gnd.n3388 585
R3734 gnd.n3368 gnd.n2646 585
R3735 gnd.n2659 gnd.n2646 585
R3736 gnd.n3367 gnd.n2657 585
R3737 gnd.n3378 gnd.n2657 585
R3738 gnd.n3358 gnd.n2664 585
R3739 gnd.n3359 gnd.n3358 585
R3740 gnd.n3357 gnd.n3356 585
R3741 gnd.n3357 gnd.n2668 585
R3742 gnd.n3355 gnd.n2670 585
R3743 gnd.n3348 gnd.n2670 585
R3744 gnd.n3335 gnd.n2671 585
R3745 gnd.n3336 gnd.n3335 585
R3746 gnd.n3288 gnd.n2684 585
R3747 gnd.n3338 gnd.n2684 585
R3748 gnd.n3290 gnd.n3289 585
R3749 gnd.n3291 gnd.n3290 585
R3750 gnd.n3283 gnd.n2786 585
R3751 gnd.n2786 gnd.n2785 585
R3752 gnd.n3281 gnd.n3280 585
R3753 gnd.n3280 gnd.n2767 585
R3754 gnd.n3278 gnd.n2765 585
R3755 gnd.n3299 gnd.n2765 585
R3756 gnd.n2796 gnd.n2795 585
R3757 gnd.n2795 gnd.n2794 585
R3758 gnd.n3272 gnd.n2755 585
R3759 gnd.n3305 gnd.n2755 585
R3760 gnd.n3271 gnd.n3270 585
R3761 gnd.n3270 gnd.n3269 585
R3762 gnd.n3267 gnd.n2798 585
R3763 gnd.n3267 gnd.n2745 585
R3764 gnd.n3266 gnd.n3265 585
R3765 gnd.n3266 gnd.n2744 585
R3766 gnd.n2801 gnd.n2800 585
R3767 gnd.n3257 gnd.n2800 585
R3768 gnd.n3225 gnd.n3224 585
R3769 gnd.n3224 gnd.n2805 585
R3770 gnd.n3226 gnd.n2814 585
R3771 gnd.n3243 gnd.n2814 585
R3772 gnd.n3223 gnd.n3222 585
R3773 gnd.n3222 gnd.n2820 585
R3774 gnd.n3221 gnd.n2828 585
R3775 gnd.n3221 gnd.n3220 585
R3776 gnd.n3206 gnd.n2829 585
R3777 gnd.n2839 gnd.n2829 585
R3778 gnd.n3205 gnd.n2837 585
R3779 gnd.n3212 gnd.n2837 585
R3780 gnd.n3204 gnd.n3203 585
R3781 gnd.n3203 gnd.n3202 585
R3782 gnd.n2848 gnd.n2845 585
R3783 gnd.n2858 gnd.n2848 585
R3784 gnd.n3194 gnd.n3193 585
R3785 gnd.n3193 gnd.n3192 585
R3786 gnd.n2854 gnd.n2853 585
R3787 gnd.n2867 gnd.n2854 585
R3788 gnd.n3174 gnd.n2865 585
R3789 gnd.n3182 gnd.n2865 585
R3790 gnd.n3173 gnd.n3172 585
R3791 gnd.n3172 gnd.n3171 585
R3792 gnd.n2874 gnd.n2872 585
R3793 gnd.n2883 gnd.n2874 585
R3794 gnd.n3163 gnd.n3162 585
R3795 gnd.n3162 gnd.n3161 585
R3796 gnd.n5932 gnd.n5931 585
R3797 gnd.n5933 gnd.n5932 585
R3798 gnd.n1257 gnd.n1256 585
R3799 gnd.n5856 gnd.n1257 585
R3800 gnd.n5941 gnd.n5940 585
R3801 gnd.n5940 gnd.n5939 585
R3802 gnd.n5942 gnd.n1251 585
R3803 gnd.n4511 gnd.n1251 585
R3804 gnd.n5944 gnd.n5943 585
R3805 gnd.n5945 gnd.n5944 585
R3806 gnd.n1236 gnd.n1235 585
R3807 gnd.n4502 gnd.n1236 585
R3808 gnd.n5953 gnd.n5952 585
R3809 gnd.n5952 gnd.n5951 585
R3810 gnd.n5954 gnd.n1230 585
R3811 gnd.n4522 gnd.n1230 585
R3812 gnd.n5956 gnd.n5955 585
R3813 gnd.n5957 gnd.n5956 585
R3814 gnd.n1214 gnd.n1213 585
R3815 gnd.n4494 gnd.n1214 585
R3816 gnd.n5965 gnd.n5964 585
R3817 gnd.n5964 gnd.n5963 585
R3818 gnd.n5966 gnd.n1208 585
R3819 gnd.n4486 gnd.n1208 585
R3820 gnd.n5968 gnd.n5967 585
R3821 gnd.n5969 gnd.n5968 585
R3822 gnd.n1194 gnd.n1193 585
R3823 gnd.n4478 gnd.n1194 585
R3824 gnd.n5977 gnd.n5976 585
R3825 gnd.n5976 gnd.n5975 585
R3826 gnd.n5978 gnd.n1188 585
R3827 gnd.n4470 gnd.n1188 585
R3828 gnd.n5980 gnd.n5979 585
R3829 gnd.n5981 gnd.n5980 585
R3830 gnd.n1172 gnd.n1171 585
R3831 gnd.n4416 gnd.n1172 585
R3832 gnd.n5989 gnd.n5988 585
R3833 gnd.n5988 gnd.n5987 585
R3834 gnd.n5990 gnd.n1167 585
R3835 gnd.n4404 gnd.n1167 585
R3836 gnd.n5992 gnd.n5991 585
R3837 gnd.n5993 gnd.n5992 585
R3838 gnd.n1152 gnd.n1150 585
R3839 gnd.n4399 gnd.n1152 585
R3840 gnd.n6001 gnd.n6000 585
R3841 gnd.n6000 gnd.n5999 585
R3842 gnd.n1151 gnd.n1149 585
R3843 gnd.n4430 gnd.n1151 585
R3844 gnd.n4391 gnd.n4390 585
R3845 gnd.n4392 gnd.n4391 585
R3846 gnd.n4389 gnd.n4388 585
R3847 gnd.n4388 gnd.n4387 585
R3848 gnd.n4359 gnd.n2351 585
R3849 gnd.n4374 gnd.n2351 585
R3850 gnd.n4361 gnd.n4360 585
R3851 gnd.n4362 gnd.n4361 585
R3852 gnd.n4358 gnd.n4357 585
R3853 gnd.n4358 gnd.n2366 585
R3854 gnd.n4356 gnd.n1148 585
R3855 gnd.n4356 gnd.n4355 585
R3856 gnd.n2369 gnd.n1142 585
R3857 gnd.n4318 gnd.n2369 585
R3858 gnd.n6004 gnd.n1141 585
R3859 gnd.n4344 gnd.n1141 585
R3860 gnd.n6005 gnd.n1137 585
R3861 gnd.n4324 gnd.n1137 585
R3862 gnd.n6007 gnd.n6006 585
R3863 gnd.n6008 gnd.n6007 585
R3864 gnd.n1121 gnd.n1120 585
R3865 gnd.n4330 gnd.n1121 585
R3866 gnd.n6016 gnd.n6015 585
R3867 gnd.n6015 gnd.n6014 585
R3868 gnd.n6017 gnd.n1115 585
R3869 gnd.n1115 gnd.n1112 585
R3870 gnd.n6019 gnd.n6018 585
R3871 gnd.n6020 gnd.n6019 585
R3872 gnd.n1116 gnd.n1114 585
R3873 gnd.n1114 gnd.n1109 585
R3874 gnd.n4280 gnd.n4279 585
R3875 gnd.n4281 gnd.n4280 585
R3876 gnd.n2406 gnd.n2405 585
R3877 gnd.n2405 gnd.n2402 585
R3878 gnd.n4274 gnd.n4273 585
R3879 gnd.n4273 gnd.n4272 585
R3880 gnd.n2409 gnd.n2408 585
R3881 gnd.n2420 gnd.n2409 585
R3882 gnd.n4253 gnd.n4252 585
R3883 gnd.n4254 gnd.n4253 585
R3884 gnd.n2422 gnd.n2421 585
R3885 gnd.n2429 gnd.n2421 585
R3886 gnd.n4248 gnd.n4247 585
R3887 gnd.n4247 gnd.n4246 585
R3888 gnd.n2425 gnd.n2424 585
R3889 gnd.n2426 gnd.n2425 585
R3890 gnd.n4237 gnd.n4236 585
R3891 gnd.n4238 gnd.n4237 585
R3892 gnd.n2439 gnd.n2438 585
R3893 gnd.n2438 gnd.n2435 585
R3894 gnd.n4232 gnd.n4231 585
R3895 gnd.n4231 gnd.n4230 585
R3896 gnd.n2442 gnd.n2441 585
R3897 gnd.n2443 gnd.n2442 585
R3898 gnd.n4221 gnd.n4220 585
R3899 gnd.n4222 gnd.n4221 585
R3900 gnd.n2454 gnd.n2453 585
R3901 gnd.n4096 gnd.n2453 585
R3902 gnd.n4216 gnd.n4215 585
R3903 gnd.n4215 gnd.n4214 585
R3904 gnd.n3967 gnd.n2456 585
R3905 gnd.n3970 gnd.n3969 585
R3906 gnd.n3966 gnd.n3965 585
R3907 gnd.n3965 gnd.n3920 585
R3908 gnd.n3975 gnd.n3974 585
R3909 gnd.n3977 gnd.n3964 585
R3910 gnd.n3980 gnd.n3979 585
R3911 gnd.n3962 gnd.n3961 585
R3912 gnd.n3985 gnd.n3984 585
R3913 gnd.n3987 gnd.n3960 585
R3914 gnd.n3990 gnd.n3989 585
R3915 gnd.n3958 gnd.n3957 585
R3916 gnd.n3995 gnd.n3994 585
R3917 gnd.n3997 gnd.n3956 585
R3918 gnd.n4000 gnd.n3999 585
R3919 gnd.n3954 gnd.n3953 585
R3920 gnd.n4005 gnd.n4004 585
R3921 gnd.n4007 gnd.n3949 585
R3922 gnd.n4010 gnd.n4009 585
R3923 gnd.n3947 gnd.n3946 585
R3924 gnd.n4015 gnd.n4014 585
R3925 gnd.n4017 gnd.n3945 585
R3926 gnd.n4020 gnd.n4019 585
R3927 gnd.n3943 gnd.n3942 585
R3928 gnd.n4025 gnd.n4024 585
R3929 gnd.n4027 gnd.n3941 585
R3930 gnd.n4030 gnd.n4029 585
R3931 gnd.n3939 gnd.n3938 585
R3932 gnd.n4035 gnd.n4034 585
R3933 gnd.n4037 gnd.n3937 585
R3934 gnd.n4040 gnd.n4039 585
R3935 gnd.n3935 gnd.n3934 585
R3936 gnd.n4045 gnd.n4044 585
R3937 gnd.n4047 gnd.n3933 585
R3938 gnd.n4050 gnd.n4049 585
R3939 gnd.n3931 gnd.n3930 585
R3940 gnd.n4056 gnd.n4055 585
R3941 gnd.n4058 gnd.n3929 585
R3942 gnd.n4059 gnd.n3928 585
R3943 gnd.n4062 gnd.n4061 585
R3944 gnd.n5863 gnd.n5862 585
R3945 gnd.n5865 gnd.n1339 585
R3946 gnd.n5867 gnd.n5866 585
R3947 gnd.n5868 gnd.n1332 585
R3948 gnd.n5870 gnd.n5869 585
R3949 gnd.n5872 gnd.n1330 585
R3950 gnd.n5874 gnd.n5873 585
R3951 gnd.n5875 gnd.n1325 585
R3952 gnd.n5877 gnd.n5876 585
R3953 gnd.n5879 gnd.n1323 585
R3954 gnd.n5881 gnd.n5880 585
R3955 gnd.n5882 gnd.n1318 585
R3956 gnd.n5884 gnd.n5883 585
R3957 gnd.n5886 gnd.n1316 585
R3958 gnd.n5888 gnd.n5887 585
R3959 gnd.n5889 gnd.n1311 585
R3960 gnd.n5891 gnd.n5890 585
R3961 gnd.n5893 gnd.n1309 585
R3962 gnd.n5895 gnd.n5894 585
R3963 gnd.n5896 gnd.n1303 585
R3964 gnd.n5898 gnd.n5897 585
R3965 gnd.n5902 gnd.n1298 585
R3966 gnd.n5904 gnd.n5903 585
R3967 gnd.n5905 gnd.n1293 585
R3968 gnd.n5907 gnd.n5906 585
R3969 gnd.n5909 gnd.n1291 585
R3970 gnd.n5911 gnd.n5910 585
R3971 gnd.n5912 gnd.n1286 585
R3972 gnd.n5914 gnd.n5913 585
R3973 gnd.n5916 gnd.n1284 585
R3974 gnd.n5918 gnd.n5917 585
R3975 gnd.n5919 gnd.n1278 585
R3976 gnd.n5921 gnd.n5920 585
R3977 gnd.n5923 gnd.n1277 585
R3978 gnd.n5924 gnd.n1275 585
R3979 gnd.n5927 gnd.n5926 585
R3980 gnd.n5928 gnd.n1272 585
R3981 gnd.n1276 gnd.n1272 585
R3982 gnd.n5859 gnd.n1269 585
R3983 gnd.n5933 gnd.n1269 585
R3984 gnd.n5858 gnd.n5857 585
R3985 gnd.n5857 gnd.n5856 585
R3986 gnd.n1343 gnd.n1259 585
R3987 gnd.n5939 gnd.n1259 585
R3988 gnd.n4510 gnd.n4509 585
R3989 gnd.n4511 gnd.n4510 585
R3990 gnd.n2306 gnd.n1248 585
R3991 gnd.n5945 gnd.n1248 585
R3992 gnd.n4504 gnd.n4503 585
R3993 gnd.n4503 gnd.n4502 585
R3994 gnd.n4501 gnd.n1237 585
R3995 gnd.n5951 gnd.n1237 585
R3996 gnd.n4500 gnd.n2300 585
R3997 gnd.n4522 gnd.n2300 585
R3998 gnd.n2308 gnd.n1227 585
R3999 gnd.n5957 gnd.n1227 585
R4000 gnd.n4496 gnd.n4495 585
R4001 gnd.n4495 gnd.n4494 585
R4002 gnd.n2310 gnd.n1216 585
R4003 gnd.n5963 gnd.n1216 585
R4004 gnd.n4485 gnd.n4484 585
R4005 gnd.n4486 gnd.n4485 585
R4006 gnd.n2315 gnd.n1206 585
R4007 gnd.n5969 gnd.n1206 585
R4008 gnd.n4480 gnd.n4479 585
R4009 gnd.n4479 gnd.n4478 585
R4010 gnd.n2317 gnd.n1195 585
R4011 gnd.n5975 gnd.n1195 585
R4012 gnd.n4412 gnd.n2321 585
R4013 gnd.n4470 gnd.n2321 585
R4014 gnd.n4413 gnd.n1185 585
R4015 gnd.n5981 gnd.n1185 585
R4016 gnd.n4415 gnd.n4414 585
R4017 gnd.n4416 gnd.n4415 585
R4018 gnd.n2343 gnd.n1174 585
R4019 gnd.n5987 gnd.n1174 585
R4020 gnd.n4406 gnd.n4405 585
R4021 gnd.n4405 gnd.n4404 585
R4022 gnd.n4402 gnd.n1165 585
R4023 gnd.n5993 gnd.n1165 585
R4024 gnd.n4401 gnd.n4400 585
R4025 gnd.n4400 gnd.n4399 585
R4026 gnd.n2345 gnd.n1153 585
R4027 gnd.n5999 gnd.n1153 585
R4028 gnd.n4395 gnd.n2334 585
R4029 gnd.n4430 gnd.n2334 585
R4030 gnd.n4394 gnd.n4393 585
R4031 gnd.n4393 gnd.n4392 585
R4032 gnd.n2348 gnd.n2347 585
R4033 gnd.n4387 gnd.n2348 585
R4034 gnd.n4376 gnd.n4375 585
R4035 gnd.n4375 gnd.n4374 585
R4036 gnd.n2359 gnd.n2358 585
R4037 gnd.n4362 gnd.n2359 585
R4038 gnd.n4300 gnd.n4299 585
R4039 gnd.n4299 gnd.n2366 585
R4040 gnd.n4301 gnd.n2371 585
R4041 gnd.n4355 gnd.n2371 585
R4042 gnd.n4320 gnd.n4319 585
R4043 gnd.n4319 gnd.n4318 585
R4044 gnd.n4321 gnd.n2379 585
R4045 gnd.n4344 gnd.n2379 585
R4046 gnd.n4323 gnd.n4322 585
R4047 gnd.n4324 gnd.n4323 585
R4048 gnd.n2396 gnd.n1134 585
R4049 gnd.n6008 gnd.n1134 585
R4050 gnd.n4291 gnd.n2390 585
R4051 gnd.n4330 gnd.n2390 585
R4052 gnd.n4290 gnd.n1123 585
R4053 gnd.n6014 gnd.n1123 585
R4054 gnd.n4289 gnd.n4288 585
R4055 gnd.n4288 gnd.n1112 585
R4056 gnd.n2398 gnd.n1110 585
R4057 gnd.n6020 gnd.n1110 585
R4058 gnd.n4284 gnd.n4283 585
R4059 gnd.n4283 gnd.n1109 585
R4060 gnd.n4282 gnd.n2400 585
R4061 gnd.n4282 gnd.n4281 585
R4062 gnd.n4075 gnd.n2401 585
R4063 gnd.n2402 gnd.n2401 585
R4064 gnd.n4076 gnd.n2410 585
R4065 gnd.n4272 gnd.n2410 585
R4066 gnd.n4078 gnd.n4077 585
R4067 gnd.n4077 gnd.n2420 585
R4068 gnd.n4079 gnd.n2418 585
R4069 gnd.n4254 gnd.n2418 585
R4070 gnd.n4081 gnd.n4080 585
R4071 gnd.n4080 gnd.n2429 585
R4072 gnd.n4082 gnd.n2427 585
R4073 gnd.n4246 gnd.n2427 585
R4074 gnd.n4084 gnd.n4083 585
R4075 gnd.n4083 gnd.n2426 585
R4076 gnd.n4085 gnd.n2436 585
R4077 gnd.n4238 gnd.n2436 585
R4078 gnd.n4087 gnd.n4086 585
R4079 gnd.n4086 gnd.n2435 585
R4080 gnd.n4088 gnd.n2444 585
R4081 gnd.n4230 gnd.n2444 585
R4082 gnd.n4090 gnd.n4089 585
R4083 gnd.n4089 gnd.n2443 585
R4084 gnd.n3924 gnd.n2451 585
R4085 gnd.n4222 gnd.n2451 585
R4086 gnd.n4095 gnd.n4094 585
R4087 gnd.n4096 gnd.n4095 585
R4088 gnd.n3923 gnd.n3921 585
R4089 gnd.n4214 gnd.n3921 585
R4090 gnd.n7326 gnd.n7325 585
R4091 gnd.n7327 gnd.n7326 585
R4092 gnd.n106 gnd.n104 585
R4093 gnd.n7248 gnd.n104 585
R4094 gnd.n7169 gnd.n191 585
R4095 gnd.n191 gnd.n189 585
R4096 gnd.n7171 gnd.n7170 585
R4097 gnd.n7172 gnd.n7171 585
R4098 gnd.n192 gnd.n190 585
R4099 gnd.n190 gnd.n186 585
R4100 gnd.n7164 gnd.n7163 585
R4101 gnd.n7163 gnd.n7162 585
R4102 gnd.n195 gnd.n194 585
R4103 gnd.n196 gnd.n195 585
R4104 gnd.n7153 gnd.n7152 585
R4105 gnd.n7154 gnd.n7153 585
R4106 gnd.n207 gnd.n206 585
R4107 gnd.n206 gnd.n203 585
R4108 gnd.n7148 gnd.n7147 585
R4109 gnd.n7147 gnd.n7146 585
R4110 gnd.n210 gnd.n209 585
R4111 gnd.n219 gnd.n210 585
R4112 gnd.n7137 gnd.n7136 585
R4113 gnd.n7138 gnd.n7137 585
R4114 gnd.n221 gnd.n220 585
R4115 gnd.n227 gnd.n220 585
R4116 gnd.n7132 gnd.n7131 585
R4117 gnd.n7131 gnd.n7130 585
R4118 gnd.n224 gnd.n223 585
R4119 gnd.n225 gnd.n224 585
R4120 gnd.n7121 gnd.n7120 585
R4121 gnd.n7122 gnd.n7121 585
R4122 gnd.n237 gnd.n236 585
R4123 gnd.n243 gnd.n236 585
R4124 gnd.n7116 gnd.n7115 585
R4125 gnd.n7115 gnd.n7114 585
R4126 gnd.n240 gnd.n239 585
R4127 gnd.n545 gnd.n240 585
R4128 gnd.n7105 gnd.n7104 585
R4129 gnd.n7106 gnd.n7105 585
R4130 gnd.n254 gnd.n253 585
R4131 gnd.n549 gnd.n253 585
R4132 gnd.n7100 gnd.n7099 585
R4133 gnd.n7099 gnd.n7098 585
R4134 gnd.n257 gnd.n256 585
R4135 gnd.n6837 gnd.n257 585
R4136 gnd.n7089 gnd.n7088 585
R4137 gnd.n7090 gnd.n7089 585
R4138 gnd.n7086 gnd.n269 585
R4139 gnd.n6841 gnd.n269 585
R4140 gnd.n7085 gnd.n7084 585
R4141 gnd.n7084 gnd.n7083 585
R4142 gnd.n7071 gnd.n271 585
R4143 gnd.n6845 gnd.n271 585
R4144 gnd.n7073 gnd.n7072 585
R4145 gnd.n7074 gnd.n7073 585
R4146 gnd.n7069 gnd.n285 585
R4147 gnd.n6851 gnd.n285 585
R4148 gnd.n7068 gnd.n7067 585
R4149 gnd.n7067 gnd.n7066 585
R4150 gnd.n287 gnd.n286 585
R4151 gnd.n5554 gnd.n287 585
R4152 gnd.n7057 gnd.n7056 585
R4153 gnd.n7058 gnd.n7057 585
R4154 gnd.n7054 gnd.n300 585
R4155 gnd.n5533 gnd.n300 585
R4156 gnd.n305 gnd.n301 585
R4157 gnd.n5576 gnd.n305 585
R4158 gnd.n7050 gnd.n7049 585
R4159 gnd.n7049 gnd.n7048 585
R4160 gnd.n304 gnd.n303 585
R4161 gnd.n5582 gnd.n304 585
R4162 gnd.n7038 gnd.n7037 585
R4163 gnd.n7039 gnd.n7038 585
R4164 gnd.n321 gnd.n320 585
R4165 gnd.n5522 gnd.n320 585
R4166 gnd.n7033 gnd.n7032 585
R4167 gnd.n7032 gnd.n7031 585
R4168 gnd.n324 gnd.n323 585
R4169 gnd.n5518 gnd.n324 585
R4170 gnd.n7022 gnd.n7021 585
R4171 gnd.n7023 gnd.n7022 585
R4172 gnd.n339 gnd.n338 585
R4173 gnd.n5512 gnd.n338 585
R4174 gnd.n7017 gnd.n7016 585
R4175 gnd.n7016 gnd.n7015 585
R4176 gnd.n342 gnd.n341 585
R4177 gnd.n5598 gnd.n342 585
R4178 gnd.n7006 gnd.n7005 585
R4179 gnd.n7007 gnd.n7006 585
R4180 gnd.n356 gnd.n355 585
R4181 gnd.n5602 gnd.n355 585
R4182 gnd.n7001 gnd.n7000 585
R4183 gnd.n7000 gnd.n6999 585
R4184 gnd.n359 gnd.n358 585
R4185 gnd.n5606 gnd.n359 585
R4186 gnd.n6990 gnd.n6989 585
R4187 gnd.n6991 gnd.n6990 585
R4188 gnd.n374 gnd.n373 585
R4189 gnd.n5610 gnd.n373 585
R4190 gnd.n6985 gnd.n6984 585
R4191 gnd.n6984 gnd.n6983 585
R4192 gnd.n377 gnd.n376 585
R4193 gnd.n5616 gnd.n377 585
R4194 gnd.n6974 gnd.n6973 585
R4195 gnd.n6975 gnd.n6974 585
R4196 gnd.n391 gnd.n390 585
R4197 gnd.n6894 gnd.n390 585
R4198 gnd.n6969 gnd.n6968 585
R4199 gnd.n394 gnd.n393 585
R4200 gnd.n6965 gnd.n6964 585
R4201 gnd.n6966 gnd.n6965 585
R4202 gnd.n6963 gnd.n425 585
R4203 gnd.n6962 gnd.n6961 585
R4204 gnd.n6960 gnd.n6959 585
R4205 gnd.n6958 gnd.n6957 585
R4206 gnd.n6956 gnd.n6955 585
R4207 gnd.n6954 gnd.n6953 585
R4208 gnd.n6952 gnd.n6951 585
R4209 gnd.n6950 gnd.n6949 585
R4210 gnd.n6948 gnd.n6947 585
R4211 gnd.n6946 gnd.n6945 585
R4212 gnd.n6944 gnd.n6943 585
R4213 gnd.n6942 gnd.n6941 585
R4214 gnd.n6940 gnd.n6939 585
R4215 gnd.n6937 gnd.n6936 585
R4216 gnd.n6935 gnd.n6934 585
R4217 gnd.n6933 gnd.n6932 585
R4218 gnd.n6931 gnd.n6930 585
R4219 gnd.n6929 gnd.n6928 585
R4220 gnd.n6927 gnd.n6926 585
R4221 gnd.n6925 gnd.n6924 585
R4222 gnd.n6923 gnd.n6922 585
R4223 gnd.n6921 gnd.n6920 585
R4224 gnd.n6919 gnd.n6918 585
R4225 gnd.n6917 gnd.n6916 585
R4226 gnd.n6915 gnd.n6914 585
R4227 gnd.n6913 gnd.n6912 585
R4228 gnd.n6911 gnd.n6910 585
R4229 gnd.n6909 gnd.n6908 585
R4230 gnd.n6907 gnd.n6906 585
R4231 gnd.n6905 gnd.n6904 585
R4232 gnd.n6903 gnd.n6902 585
R4233 gnd.n6901 gnd.n463 585
R4234 gnd.n467 gnd.n464 585
R4235 gnd.n6897 gnd.n6896 585
R4236 gnd.n174 gnd.n173 585
R4237 gnd.n7255 gnd.n169 585
R4238 gnd.n7257 gnd.n7256 585
R4239 gnd.n7259 gnd.n167 585
R4240 gnd.n7261 gnd.n7260 585
R4241 gnd.n7262 gnd.n162 585
R4242 gnd.n7264 gnd.n7263 585
R4243 gnd.n7266 gnd.n160 585
R4244 gnd.n7268 gnd.n7267 585
R4245 gnd.n7269 gnd.n155 585
R4246 gnd.n7271 gnd.n7270 585
R4247 gnd.n7273 gnd.n153 585
R4248 gnd.n7275 gnd.n7274 585
R4249 gnd.n7276 gnd.n148 585
R4250 gnd.n7278 gnd.n7277 585
R4251 gnd.n7280 gnd.n146 585
R4252 gnd.n7282 gnd.n7281 585
R4253 gnd.n7283 gnd.n141 585
R4254 gnd.n7285 gnd.n7284 585
R4255 gnd.n7287 gnd.n139 585
R4256 gnd.n7289 gnd.n7288 585
R4257 gnd.n7293 gnd.n134 585
R4258 gnd.n7295 gnd.n7294 585
R4259 gnd.n7297 gnd.n132 585
R4260 gnd.n7299 gnd.n7298 585
R4261 gnd.n7300 gnd.n127 585
R4262 gnd.n7302 gnd.n7301 585
R4263 gnd.n7304 gnd.n125 585
R4264 gnd.n7306 gnd.n7305 585
R4265 gnd.n7307 gnd.n120 585
R4266 gnd.n7309 gnd.n7308 585
R4267 gnd.n7311 gnd.n118 585
R4268 gnd.n7313 gnd.n7312 585
R4269 gnd.n7314 gnd.n113 585
R4270 gnd.n7316 gnd.n7315 585
R4271 gnd.n7318 gnd.n111 585
R4272 gnd.n7320 gnd.n7319 585
R4273 gnd.n7321 gnd.n109 585
R4274 gnd.n7322 gnd.n105 585
R4275 gnd.n105 gnd.n102 585
R4276 gnd.n7251 gnd.n101 585
R4277 gnd.n7327 gnd.n101 585
R4278 gnd.n7250 gnd.n7249 585
R4279 gnd.n7249 gnd.n7248 585
R4280 gnd.n179 gnd.n178 585
R4281 gnd.n189 gnd.n179 585
R4282 gnd.n523 gnd.n187 585
R4283 gnd.n7172 gnd.n187 585
R4284 gnd.n525 gnd.n524 585
R4285 gnd.n524 gnd.n186 585
R4286 gnd.n526 gnd.n197 585
R4287 gnd.n7162 gnd.n197 585
R4288 gnd.n528 gnd.n527 585
R4289 gnd.n527 gnd.n196 585
R4290 gnd.n529 gnd.n204 585
R4291 gnd.n7154 gnd.n204 585
R4292 gnd.n531 gnd.n530 585
R4293 gnd.n530 gnd.n203 585
R4294 gnd.n532 gnd.n211 585
R4295 gnd.n7146 gnd.n211 585
R4296 gnd.n534 gnd.n533 585
R4297 gnd.n533 gnd.n219 585
R4298 gnd.n535 gnd.n217 585
R4299 gnd.n7138 gnd.n217 585
R4300 gnd.n537 gnd.n536 585
R4301 gnd.n536 gnd.n227 585
R4302 gnd.n538 gnd.n226 585
R4303 gnd.n7130 gnd.n226 585
R4304 gnd.n540 gnd.n539 585
R4305 gnd.n539 gnd.n225 585
R4306 gnd.n541 gnd.n234 585
R4307 gnd.n7122 gnd.n234 585
R4308 gnd.n543 gnd.n542 585
R4309 gnd.n542 gnd.n243 585
R4310 gnd.n544 gnd.n242 585
R4311 gnd.n7114 gnd.n242 585
R4312 gnd.n547 gnd.n546 585
R4313 gnd.n546 gnd.n545 585
R4314 gnd.n548 gnd.n250 585
R4315 gnd.n7106 gnd.n250 585
R4316 gnd.n551 gnd.n550 585
R4317 gnd.n550 gnd.n549 585
R4318 gnd.n552 gnd.n259 585
R4319 gnd.n7098 gnd.n259 585
R4320 gnd.n6839 gnd.n6838 585
R4321 gnd.n6838 gnd.n6837 585
R4322 gnd.n6840 gnd.n267 585
R4323 gnd.n7090 gnd.n267 585
R4324 gnd.n6843 gnd.n6842 585
R4325 gnd.n6842 gnd.n6841 585
R4326 gnd.n6844 gnd.n273 585
R4327 gnd.n7083 gnd.n273 585
R4328 gnd.n6847 gnd.n6846 585
R4329 gnd.n6846 gnd.n6845 585
R4330 gnd.n6848 gnd.n282 585
R4331 gnd.n7074 gnd.n282 585
R4332 gnd.n6850 gnd.n6849 585
R4333 gnd.n6851 gnd.n6850 585
R4334 gnd.n495 gnd.n289 585
R4335 gnd.n7066 gnd.n289 585
R4336 gnd.n5553 gnd.n5552 585
R4337 gnd.n5554 gnd.n5553 585
R4338 gnd.n5547 gnd.n298 585
R4339 gnd.n7058 gnd.n298 585
R4340 gnd.n5531 gnd.n5530 585
R4341 gnd.n5533 gnd.n5531 585
R4342 gnd.n5578 gnd.n5577 585
R4343 gnd.n5577 gnd.n5576 585
R4344 gnd.n5579 gnd.n307 585
R4345 gnd.n7048 gnd.n307 585
R4346 gnd.n5581 gnd.n5580 585
R4347 gnd.n5582 gnd.n5581 585
R4348 gnd.n5508 gnd.n318 585
R4349 gnd.n7039 gnd.n318 585
R4350 gnd.n5524 gnd.n5523 585
R4351 gnd.n5523 gnd.n5522 585
R4352 gnd.n5521 gnd.n326 585
R4353 gnd.n7031 gnd.n326 585
R4354 gnd.n5520 gnd.n5519 585
R4355 gnd.n5519 gnd.n5518 585
R4356 gnd.n5510 gnd.n335 585
R4357 gnd.n7023 gnd.n335 585
R4358 gnd.n5514 gnd.n5513 585
R4359 gnd.n5513 gnd.n5512 585
R4360 gnd.n5475 gnd.n344 585
R4361 gnd.n7015 gnd.n344 585
R4362 gnd.n5600 gnd.n5599 585
R4363 gnd.n5599 gnd.n5598 585
R4364 gnd.n5601 gnd.n353 585
R4365 gnd.n7007 gnd.n353 585
R4366 gnd.n5604 gnd.n5603 585
R4367 gnd.n5603 gnd.n5602 585
R4368 gnd.n5605 gnd.n361 585
R4369 gnd.n6999 gnd.n361 585
R4370 gnd.n5608 gnd.n5607 585
R4371 gnd.n5607 gnd.n5606 585
R4372 gnd.n5609 gnd.n370 585
R4373 gnd.n6991 gnd.n370 585
R4374 gnd.n5612 gnd.n5611 585
R4375 gnd.n5611 gnd.n5610 585
R4376 gnd.n5613 gnd.n379 585
R4377 gnd.n6983 gnd.n379 585
R4378 gnd.n5615 gnd.n5614 585
R4379 gnd.n5616 gnd.n5615 585
R4380 gnd.n5464 gnd.n388 585
R4381 gnd.n6975 gnd.n388 585
R4382 gnd.n6895 gnd.n469 585
R4383 gnd.n6895 gnd.n6894 585
R4384 gnd.n5325 gnd.n5324 585
R4385 gnd.n5326 gnd.n5325 585
R4386 gnd.n5236 gnd.n1650 585
R4387 gnd.n1656 gnd.n1650 585
R4388 gnd.n5235 gnd.n5234 585
R4389 gnd.n5234 gnd.n5233 585
R4390 gnd.n1653 gnd.n1652 585
R4391 gnd.n4920 gnd.n1653 585
R4392 gnd.n5198 gnd.n1663 585
R4393 gnd.n5223 gnd.n1663 585
R4394 gnd.n5199 gnd.n1677 585
R4395 gnd.n4924 gnd.n1677 585
R4396 gnd.n5201 gnd.n5200 585
R4397 gnd.n5202 gnd.n5201 585
R4398 gnd.n5197 gnd.n1676 585
R4399 gnd.n1676 gnd.n1673 585
R4400 gnd.n5196 gnd.n5195 585
R4401 gnd.n5195 gnd.n5194 585
R4402 gnd.n1679 gnd.n1678 585
R4403 gnd.n4933 gnd.n1679 585
R4404 gnd.n5183 gnd.n5182 585
R4405 gnd.n5184 gnd.n5183 585
R4406 gnd.n5181 gnd.n1689 585
R4407 gnd.n4937 gnd.n1689 585
R4408 gnd.n5180 gnd.n5179 585
R4409 gnd.n5179 gnd.n5178 585
R4410 gnd.n1691 gnd.n1690 585
R4411 gnd.n4942 gnd.n1691 585
R4412 gnd.n5165 gnd.n5164 585
R4413 gnd.n5166 gnd.n5165 585
R4414 gnd.n5163 gnd.n1703 585
R4415 gnd.n1703 gnd.n1700 585
R4416 gnd.n5162 gnd.n5161 585
R4417 gnd.n5161 gnd.n5160 585
R4418 gnd.n1705 gnd.n1704 585
R4419 gnd.n4950 gnd.n1705 585
R4420 gnd.n5135 gnd.n5134 585
R4421 gnd.n5134 gnd.n1716 585
R4422 gnd.n5136 gnd.n1725 585
R4423 gnd.n4954 gnd.n1725 585
R4424 gnd.n5138 gnd.n5137 585
R4425 gnd.n5139 gnd.n5138 585
R4426 gnd.n5133 gnd.n1724 585
R4427 gnd.n5128 gnd.n1724 585
R4428 gnd.n5132 gnd.n5131 585
R4429 gnd.n5131 gnd.n5130 585
R4430 gnd.n1727 gnd.n1726 585
R4431 gnd.n1738 gnd.n1727 585
R4432 gnd.n5105 gnd.n5104 585
R4433 gnd.n5104 gnd.n1737 585
R4434 gnd.n5106 gnd.n1747 585
R4435 gnd.n4964 gnd.n1747 585
R4436 gnd.n5108 gnd.n5107 585
R4437 gnd.n5109 gnd.n5108 585
R4438 gnd.n5103 gnd.n1746 585
R4439 gnd.n5098 gnd.n1746 585
R4440 gnd.n5102 gnd.n5101 585
R4441 gnd.n5101 gnd.n5100 585
R4442 gnd.n1749 gnd.n1748 585
R4443 gnd.n5088 gnd.n1749 585
R4444 gnd.n5075 gnd.n1770 585
R4445 gnd.n1770 gnd.n1759 585
R4446 gnd.n5077 gnd.n5076 585
R4447 gnd.n5078 gnd.n5077 585
R4448 gnd.n5074 gnd.n1769 585
R4449 gnd.n1769 gnd.n1766 585
R4450 gnd.n5073 gnd.n5072 585
R4451 gnd.n5072 gnd.n5071 585
R4452 gnd.n1772 gnd.n1771 585
R4453 gnd.n4978 gnd.n1772 585
R4454 gnd.n5060 gnd.n5059 585
R4455 gnd.n5061 gnd.n5060 585
R4456 gnd.n5058 gnd.n1784 585
R4457 gnd.n1784 gnd.n1781 585
R4458 gnd.n5057 gnd.n5056 585
R4459 gnd.n5056 gnd.n5055 585
R4460 gnd.n1786 gnd.n1785 585
R4461 gnd.n4986 gnd.n1786 585
R4462 gnd.n5042 gnd.n5041 585
R4463 gnd.n5043 gnd.n5042 585
R4464 gnd.n5040 gnd.n1799 585
R4465 gnd.n1799 gnd.n1795 585
R4466 gnd.n5039 gnd.n5038 585
R4467 gnd.n5038 gnd.n5037 585
R4468 gnd.n1801 gnd.n1800 585
R4469 gnd.n1812 gnd.n1801 585
R4470 gnd.n5012 gnd.n5011 585
R4471 gnd.n5011 gnd.n1811 585
R4472 gnd.n5013 gnd.n1821 585
R4473 gnd.n4999 gnd.n1821 585
R4474 gnd.n5015 gnd.n5014 585
R4475 gnd.n5016 gnd.n5015 585
R4476 gnd.n5010 gnd.n1820 585
R4477 gnd.n5005 gnd.n1820 585
R4478 gnd.n5009 gnd.n5008 585
R4479 gnd.n5008 gnd.n5007 585
R4480 gnd.n1823 gnd.n1822 585
R4481 gnd.n4911 gnd.n1823 585
R4482 gnd.n4897 gnd.n4896 585
R4483 gnd.n4896 gnd.n4895 585
R4484 gnd.n4898 gnd.n1836 585
R4485 gnd.n4893 gnd.n1836 585
R4486 gnd.n4900 gnd.n4899 585
R4487 gnd.n4901 gnd.n4900 585
R4488 gnd.n1837 gnd.n1835 585
R4489 gnd.n4887 gnd.n1835 585
R4490 gnd.n4852 gnd.n4851 585
R4491 gnd.n4851 gnd.n4850 585
R4492 gnd.n4853 gnd.n1851 585
R4493 gnd.n4867 gnd.n1851 585
R4494 gnd.n4854 gnd.n1863 585
R4495 gnd.n1863 gnd.n1850 585
R4496 gnd.n4856 gnd.n4855 585
R4497 gnd.n4857 gnd.n4856 585
R4498 gnd.n4848 gnd.n1862 585
R4499 gnd.n1862 gnd.n1858 585
R4500 gnd.n4847 gnd.n4846 585
R4501 gnd.n4846 gnd.n4845 585
R4502 gnd.n1865 gnd.n1864 585
R4503 gnd.n4754 gnd.n1865 585
R4504 gnd.n4834 gnd.n4833 585
R4505 gnd.n4835 gnd.n4834 585
R4506 gnd.n4832 gnd.n1876 585
R4507 gnd.n1876 gnd.n1873 585
R4508 gnd.n4831 gnd.n4830 585
R4509 gnd.n4830 gnd.n4829 585
R4510 gnd.n1878 gnd.n1877 585
R4511 gnd.n4762 gnd.n1878 585
R4512 gnd.n4816 gnd.n4815 585
R4513 gnd.n4817 gnd.n4816 585
R4514 gnd.n4814 gnd.n1891 585
R4515 gnd.n1891 gnd.n1888 585
R4516 gnd.n4813 gnd.n4812 585
R4517 gnd.n4812 gnd.n4811 585
R4518 gnd.n1893 gnd.n1892 585
R4519 gnd.n1905 gnd.n1893 585
R4520 gnd.n4786 gnd.n4785 585
R4521 gnd.n4785 gnd.n1903 585
R4522 gnd.n4787 gnd.n1915 585
R4523 gnd.n4773 gnd.n1915 585
R4524 gnd.n4789 gnd.n4788 585
R4525 gnd.n4790 gnd.n4789 585
R4526 gnd.n4784 gnd.n1914 585
R4527 gnd.n4779 gnd.n1914 585
R4528 gnd.n4783 gnd.n4782 585
R4529 gnd.n4782 gnd.n4781 585
R4530 gnd.n1917 gnd.n1916 585
R4531 gnd.n4741 gnd.n1917 585
R4532 gnd.n4727 gnd.n1935 585
R4533 gnd.n1935 gnd.n1934 585
R4534 gnd.n4729 gnd.n4728 585
R4535 gnd.n4730 gnd.n4729 585
R4536 gnd.n4726 gnd.n1931 585
R4537 gnd.n1940 gnd.n1931 585
R4538 gnd.n4725 gnd.n4724 585
R4539 gnd.n4724 gnd.n4723 585
R4540 gnd.n1937 gnd.n1936 585
R4541 gnd.n4678 gnd.n1937 585
R4542 gnd.n4693 gnd.n1949 585
R4543 gnd.n4708 gnd.n1949 585
R4544 gnd.n4694 gnd.n1958 585
R4545 gnd.n1958 gnd.n1957 585
R4546 gnd.n4696 gnd.n4695 585
R4547 gnd.n4697 gnd.n4696 585
R4548 gnd.n4692 gnd.n1955 585
R4549 gnd.n1982 gnd.n1955 585
R4550 gnd.n4691 gnd.n4690 585
R4551 gnd.n4690 gnd.n4689 585
R4552 gnd.n2024 gnd.n1980 585
R4553 gnd.n2159 gnd.n2158 585
R4554 gnd.n2157 gnd.n2023 585
R4555 gnd.n2161 gnd.n2023 585
R4556 gnd.n2156 gnd.n2155 585
R4557 gnd.n2154 gnd.n2153 585
R4558 gnd.n2152 gnd.n2151 585
R4559 gnd.n2150 gnd.n2149 585
R4560 gnd.n2148 gnd.n2147 585
R4561 gnd.n2146 gnd.n2145 585
R4562 gnd.n2144 gnd.n2143 585
R4563 gnd.n2142 gnd.n2141 585
R4564 gnd.n2140 gnd.n2139 585
R4565 gnd.n2138 gnd.n2137 585
R4566 gnd.n2136 gnd.n2135 585
R4567 gnd.n2134 gnd.n2133 585
R4568 gnd.n2132 gnd.n2131 585
R4569 gnd.n2130 gnd.n2129 585
R4570 gnd.n2128 gnd.n2127 585
R4571 gnd.n2126 gnd.n2125 585
R4572 gnd.n2124 gnd.n2123 585
R4573 gnd.n2122 gnd.n2121 585
R4574 gnd.n2120 gnd.n2119 585
R4575 gnd.n2118 gnd.n2117 585
R4576 gnd.n2116 gnd.n2115 585
R4577 gnd.n2114 gnd.n2113 585
R4578 gnd.n2112 gnd.n2111 585
R4579 gnd.n2110 gnd.n2109 585
R4580 gnd.n2108 gnd.n2107 585
R4581 gnd.n2106 gnd.n2105 585
R4582 gnd.n2104 gnd.n2103 585
R4583 gnd.n2102 gnd.n2101 585
R4584 gnd.n2100 gnd.n2099 585
R4585 gnd.n2098 gnd.n2097 585
R4586 gnd.n2096 gnd.n2094 585
R4587 gnd.n2093 gnd.n2092 585
R4588 gnd.n2091 gnd.n2090 585
R4589 gnd.n2088 gnd.n2087 585
R4590 gnd.n2086 gnd.n2085 585
R4591 gnd.n2084 gnd.n2083 585
R4592 gnd.n2082 gnd.n2081 585
R4593 gnd.n2080 gnd.n2079 585
R4594 gnd.n2078 gnd.n2077 585
R4595 gnd.n2076 gnd.n2075 585
R4596 gnd.n2074 gnd.n2073 585
R4597 gnd.n2072 gnd.n2071 585
R4598 gnd.n2070 gnd.n2069 585
R4599 gnd.n2068 gnd.n2067 585
R4600 gnd.n2066 gnd.n2065 585
R4601 gnd.n2064 gnd.n2063 585
R4602 gnd.n2062 gnd.n2061 585
R4603 gnd.n2060 gnd.n2059 585
R4604 gnd.n2058 gnd.n2057 585
R4605 gnd.n2056 gnd.n2055 585
R4606 gnd.n2054 gnd.n2053 585
R4607 gnd.n2052 gnd.n2051 585
R4608 gnd.n2050 gnd.n2049 585
R4609 gnd.n2048 gnd.n2047 585
R4610 gnd.n2046 gnd.n2045 585
R4611 gnd.n2044 gnd.n2043 585
R4612 gnd.n2042 gnd.n2041 585
R4613 gnd.n2040 gnd.n2039 585
R4614 gnd.n2038 gnd.n2037 585
R4615 gnd.n2036 gnd.n2035 585
R4616 gnd.n2034 gnd.n2033 585
R4617 gnd.n2032 gnd.n2031 585
R4618 gnd.n5329 gnd.n5328 585
R4619 gnd.n5331 gnd.n5330 585
R4620 gnd.n5333 gnd.n5332 585
R4621 gnd.n5335 gnd.n5334 585
R4622 gnd.n5337 gnd.n5336 585
R4623 gnd.n5339 gnd.n5338 585
R4624 gnd.n5341 gnd.n5340 585
R4625 gnd.n5343 gnd.n5342 585
R4626 gnd.n5345 gnd.n5344 585
R4627 gnd.n5347 gnd.n5346 585
R4628 gnd.n5349 gnd.n5348 585
R4629 gnd.n5351 gnd.n5350 585
R4630 gnd.n5353 gnd.n5352 585
R4631 gnd.n5355 gnd.n5354 585
R4632 gnd.n5357 gnd.n5356 585
R4633 gnd.n5359 gnd.n5358 585
R4634 gnd.n5361 gnd.n5360 585
R4635 gnd.n5363 gnd.n5362 585
R4636 gnd.n5365 gnd.n5364 585
R4637 gnd.n5367 gnd.n5366 585
R4638 gnd.n5369 gnd.n5368 585
R4639 gnd.n5371 gnd.n5370 585
R4640 gnd.n5373 gnd.n5372 585
R4641 gnd.n5375 gnd.n5374 585
R4642 gnd.n5377 gnd.n5376 585
R4643 gnd.n5379 gnd.n5378 585
R4644 gnd.n5381 gnd.n5380 585
R4645 gnd.n5383 gnd.n5382 585
R4646 gnd.n5385 gnd.n5384 585
R4647 gnd.n5388 gnd.n5387 585
R4648 gnd.n5390 gnd.n5389 585
R4649 gnd.n5392 gnd.n5391 585
R4650 gnd.n5394 gnd.n5393 585
R4651 gnd.n5258 gnd.n440 585
R4652 gnd.n5260 gnd.n5259 585
R4653 gnd.n5262 gnd.n5261 585
R4654 gnd.n5264 gnd.n5263 585
R4655 gnd.n5267 gnd.n5266 585
R4656 gnd.n5269 gnd.n5268 585
R4657 gnd.n5271 gnd.n5270 585
R4658 gnd.n5273 gnd.n5272 585
R4659 gnd.n5275 gnd.n5274 585
R4660 gnd.n5277 gnd.n5276 585
R4661 gnd.n5279 gnd.n5278 585
R4662 gnd.n5281 gnd.n5280 585
R4663 gnd.n5283 gnd.n5282 585
R4664 gnd.n5285 gnd.n5284 585
R4665 gnd.n5287 gnd.n5286 585
R4666 gnd.n5289 gnd.n5288 585
R4667 gnd.n5291 gnd.n5290 585
R4668 gnd.n5293 gnd.n5292 585
R4669 gnd.n5295 gnd.n5294 585
R4670 gnd.n5297 gnd.n5296 585
R4671 gnd.n5299 gnd.n5298 585
R4672 gnd.n5301 gnd.n5300 585
R4673 gnd.n5303 gnd.n5302 585
R4674 gnd.n5305 gnd.n5304 585
R4675 gnd.n5307 gnd.n5306 585
R4676 gnd.n5309 gnd.n5308 585
R4677 gnd.n5311 gnd.n5310 585
R4678 gnd.n5313 gnd.n5312 585
R4679 gnd.n5315 gnd.n5314 585
R4680 gnd.n5317 gnd.n5316 585
R4681 gnd.n5319 gnd.n5318 585
R4682 gnd.n5321 gnd.n5320 585
R4683 gnd.n5322 gnd.n1651 585
R4684 gnd.n5327 gnd.n1647 585
R4685 gnd.n5327 gnd.n5326 585
R4686 gnd.n4918 gnd.n1648 585
R4687 gnd.n1656 gnd.n1648 585
R4688 gnd.n4919 gnd.n1655 585
R4689 gnd.n5233 gnd.n1655 585
R4690 gnd.n4922 gnd.n4921 585
R4691 gnd.n4921 gnd.n4920 585
R4692 gnd.n4923 gnd.n1666 585
R4693 gnd.n5223 gnd.n1666 585
R4694 gnd.n4926 gnd.n4925 585
R4695 gnd.n4925 gnd.n4924 585
R4696 gnd.n4927 gnd.n1674 585
R4697 gnd.n5202 gnd.n1674 585
R4698 gnd.n4929 gnd.n4928 585
R4699 gnd.n4928 gnd.n1673 585
R4700 gnd.n4930 gnd.n1681 585
R4701 gnd.n5194 gnd.n1681 585
R4702 gnd.n4935 gnd.n4934 585
R4703 gnd.n4934 gnd.n4933 585
R4704 gnd.n4936 gnd.n1687 585
R4705 gnd.n5184 gnd.n1687 585
R4706 gnd.n4939 gnd.n4938 585
R4707 gnd.n4938 gnd.n4937 585
R4708 gnd.n4940 gnd.n1693 585
R4709 gnd.n5178 gnd.n1693 585
R4710 gnd.n4944 gnd.n4943 585
R4711 gnd.n4943 gnd.n4942 585
R4712 gnd.n4945 gnd.n1701 585
R4713 gnd.n5166 gnd.n1701 585
R4714 gnd.n4947 gnd.n4946 585
R4715 gnd.n4946 gnd.n1700 585
R4716 gnd.n4948 gnd.n1707 585
R4717 gnd.n5160 gnd.n1707 585
R4718 gnd.n4951 gnd.n4949 585
R4719 gnd.n4951 gnd.n4950 585
R4720 gnd.n4952 gnd.n4917 585
R4721 gnd.n4952 gnd.n1716 585
R4722 gnd.n4956 gnd.n4955 585
R4723 gnd.n4955 gnd.n4954 585
R4724 gnd.n4957 gnd.n1722 585
R4725 gnd.n5139 gnd.n1722 585
R4726 gnd.n4958 gnd.n1730 585
R4727 gnd.n5128 gnd.n1730 585
R4728 gnd.n4959 gnd.n1729 585
R4729 gnd.n5130 gnd.n1729 585
R4730 gnd.n4961 gnd.n4960 585
R4731 gnd.n4961 gnd.n1738 585
R4732 gnd.n4962 gnd.n4916 585
R4733 gnd.n4962 gnd.n1737 585
R4734 gnd.n4966 gnd.n4965 585
R4735 gnd.n4965 gnd.n4964 585
R4736 gnd.n4967 gnd.n1744 585
R4737 gnd.n5109 gnd.n1744 585
R4738 gnd.n4968 gnd.n1752 585
R4739 gnd.n5098 gnd.n1752 585
R4740 gnd.n4969 gnd.n1751 585
R4741 gnd.n5100 gnd.n1751 585
R4742 gnd.n4970 gnd.n1760 585
R4743 gnd.n5088 gnd.n1760 585
R4744 gnd.n4972 gnd.n4971 585
R4745 gnd.n4971 gnd.n1759 585
R4746 gnd.n4973 gnd.n1767 585
R4747 gnd.n5078 gnd.n1767 585
R4748 gnd.n4975 gnd.n4974 585
R4749 gnd.n4974 gnd.n1766 585
R4750 gnd.n4976 gnd.n1774 585
R4751 gnd.n5071 gnd.n1774 585
R4752 gnd.n4980 gnd.n4979 585
R4753 gnd.n4979 gnd.n4978 585
R4754 gnd.n4981 gnd.n1782 585
R4755 gnd.n5061 gnd.n1782 585
R4756 gnd.n4983 gnd.n4982 585
R4757 gnd.n4982 gnd.n1781 585
R4758 gnd.n4984 gnd.n1788 585
R4759 gnd.n5055 gnd.n1788 585
R4760 gnd.n4988 gnd.n4987 585
R4761 gnd.n4987 gnd.n4986 585
R4762 gnd.n4989 gnd.n1796 585
R4763 gnd.n5043 gnd.n1796 585
R4764 gnd.n4991 gnd.n4990 585
R4765 gnd.n4990 gnd.n1795 585
R4766 gnd.n4992 gnd.n1803 585
R4767 gnd.n5037 gnd.n1803 585
R4768 gnd.n4994 gnd.n4993 585
R4769 gnd.n4994 gnd.n1812 585
R4770 gnd.n4995 gnd.n4915 585
R4771 gnd.n4995 gnd.n1811 585
R4772 gnd.n5001 gnd.n5000 585
R4773 gnd.n5000 gnd.n4999 585
R4774 gnd.n5002 gnd.n1819 585
R4775 gnd.n5016 gnd.n1819 585
R4776 gnd.n5004 gnd.n5003 585
R4777 gnd.n5005 gnd.n5004 585
R4778 gnd.n4914 gnd.n1825 585
R4779 gnd.n5007 gnd.n1825 585
R4780 gnd.n4913 gnd.n4912 585
R4781 gnd.n4912 gnd.n4911 585
R4782 gnd.n1827 gnd.n1826 585
R4783 gnd.n4895 gnd.n1827 585
R4784 gnd.n4892 gnd.n4891 585
R4785 gnd.n4893 gnd.n4892 585
R4786 gnd.n4890 gnd.n1834 585
R4787 gnd.n4901 gnd.n1834 585
R4788 gnd.n4889 gnd.n4888 585
R4789 gnd.n4888 gnd.n4887 585
R4790 gnd.n1841 gnd.n1840 585
R4791 gnd.n4850 gnd.n1841 585
R4792 gnd.n4746 gnd.n1852 585
R4793 gnd.n4867 gnd.n1852 585
R4794 gnd.n4748 gnd.n4747 585
R4795 gnd.n4747 gnd.n1850 585
R4796 gnd.n4749 gnd.n1860 585
R4797 gnd.n4857 gnd.n1860 585
R4798 gnd.n4751 gnd.n4750 585
R4799 gnd.n4750 gnd.n1858 585
R4800 gnd.n4752 gnd.n1867 585
R4801 gnd.n4845 gnd.n1867 585
R4802 gnd.n4756 gnd.n4755 585
R4803 gnd.n4755 gnd.n4754 585
R4804 gnd.n4757 gnd.n1874 585
R4805 gnd.n4835 gnd.n1874 585
R4806 gnd.n4759 gnd.n4758 585
R4807 gnd.n4758 gnd.n1873 585
R4808 gnd.n4760 gnd.n1881 585
R4809 gnd.n4829 gnd.n1881 585
R4810 gnd.n4764 gnd.n4763 585
R4811 gnd.n4763 gnd.n4762 585
R4812 gnd.n4765 gnd.n1889 585
R4813 gnd.n4817 gnd.n1889 585
R4814 gnd.n4767 gnd.n4766 585
R4815 gnd.n4766 gnd.n1888 585
R4816 gnd.n4768 gnd.n1895 585
R4817 gnd.n4811 gnd.n1895 585
R4818 gnd.n4770 gnd.n4769 585
R4819 gnd.n4770 gnd.n1905 585
R4820 gnd.n4771 gnd.n4745 585
R4821 gnd.n4771 gnd.n1903 585
R4822 gnd.n4775 gnd.n4774 585
R4823 gnd.n4774 gnd.n4773 585
R4824 gnd.n4776 gnd.n1912 585
R4825 gnd.n4790 gnd.n1912 585
R4826 gnd.n4778 gnd.n4777 585
R4827 gnd.n4779 gnd.n4778 585
R4828 gnd.n4744 gnd.n1918 585
R4829 gnd.n4781 gnd.n1918 585
R4830 gnd.n4743 gnd.n4742 585
R4831 gnd.n4742 gnd.n4741 585
R4832 gnd.n1920 gnd.n1919 585
R4833 gnd.n1934 gnd.n1920 585
R4834 gnd.n4701 gnd.n1929 585
R4835 gnd.n4730 gnd.n1929 585
R4836 gnd.n4703 gnd.n4702 585
R4837 gnd.n4702 gnd.n1940 585
R4838 gnd.n4704 gnd.n1939 585
R4839 gnd.n4723 gnd.n1939 585
R4840 gnd.n4705 gnd.n1951 585
R4841 gnd.n4678 gnd.n1951 585
R4842 gnd.n4707 gnd.n4706 585
R4843 gnd.n4708 gnd.n4707 585
R4844 gnd.n4700 gnd.n1950 585
R4845 gnd.n1957 gnd.n1950 585
R4846 gnd.n4699 gnd.n4698 585
R4847 gnd.n4698 gnd.n4697 585
R4848 gnd.n1953 gnd.n1952 585
R4849 gnd.n1982 gnd.n1953 585
R4850 gnd.n2030 gnd.n1981 585
R4851 gnd.n4689 gnd.n1981 585
R4852 gnd.n6023 gnd.n6022 585
R4853 gnd.n6022 gnd.n6021 585
R4854 gnd.n6824 gnd.n6823 585
R4855 gnd.n6823 gnd.n233 585
R4856 gnd.n6827 gnd.n559 585
R4857 gnd.n559 gnd.n241 585
R4858 gnd.n6829 gnd.n6828 585
R4859 gnd.n6829 gnd.n252 585
R4860 gnd.n6830 gnd.n558 585
R4861 gnd.n6830 gnd.n249 585
R4862 gnd.n6832 gnd.n6831 585
R4863 gnd.n6831 gnd.n260 585
R4864 gnd.n6833 gnd.n554 585
R4865 gnd.n554 gnd.n258 585
R4866 gnd.n6835 gnd.n6834 585
R4867 gnd.n6836 gnd.n6835 585
R4868 gnd.n5557 gnd.n553 585
R4869 gnd.n553 gnd.n266 585
R4870 gnd.n5559 gnd.n5558 585
R4871 gnd.n5559 gnd.n274 585
R4872 gnd.n5561 gnd.n5560 585
R4873 gnd.n5560 gnd.n272 585
R4874 gnd.n5563 gnd.n5562 585
R4875 gnd.n5563 gnd.n284 585
R4876 gnd.n5565 gnd.n5564 585
R4877 gnd.n5565 gnd.n281 585
R4878 gnd.n5566 gnd.n5546 585
R4879 gnd.n5566 gnd.n291 585
R4880 gnd.n5568 gnd.n5567 585
R4881 gnd.n5567 gnd.n288 585
R4882 gnd.n5556 gnd.n5543 585
R4883 gnd.n5556 gnd.n5555 585
R4884 gnd.n5572 gnd.n5535 585
R4885 gnd.n5535 gnd.n297 585
R4886 gnd.n5574 gnd.n5573 585
R4887 gnd.n5575 gnd.n5574 585
R4888 gnd.n5536 gnd.n5534 585
R4889 gnd.n5534 gnd.n309 585
R4890 gnd.n5539 gnd.n5506 585
R4891 gnd.n5506 gnd.n306 585
R4892 gnd.n5584 gnd.n5507 585
R4893 gnd.n5584 gnd.n5583 585
R4894 gnd.n5585 gnd.n5505 585
R4895 gnd.n5585 gnd.n317 585
R4896 gnd.n5587 gnd.n5586 585
R4897 gnd.n5586 gnd.n328 585
R4898 gnd.n5588 gnd.n5500 585
R4899 gnd.n5500 gnd.n325 585
R4900 gnd.n5590 gnd.n5589 585
R4901 gnd.n5590 gnd.n337 585
R4902 gnd.n5591 gnd.n5499 585
R4903 gnd.n5591 gnd.n334 585
R4904 gnd.n5593 gnd.n5592 585
R4905 gnd.n5592 gnd.n346 585
R4906 gnd.n5594 gnd.n5477 585
R4907 gnd.n5477 gnd.n343 585
R4908 gnd.n5596 gnd.n5595 585
R4909 gnd.n5597 gnd.n5596 585
R4910 gnd.n5478 gnd.n5476 585
R4911 gnd.n5476 gnd.n352 585
R4912 gnd.n5493 gnd.n5492 585
R4913 gnd.n5492 gnd.n363 585
R4914 gnd.n5491 gnd.n5480 585
R4915 gnd.n5491 gnd.n360 585
R4916 gnd.n5490 gnd.n5489 585
R4917 gnd.n5490 gnd.n372 585
R4918 gnd.n5482 gnd.n5481 585
R4919 gnd.n5481 gnd.n369 585
R4920 gnd.n5485 gnd.n5484 585
R4921 gnd.n5484 gnd.n381 585
R4922 gnd.n5463 gnd.n5462 585
R4923 gnd.n5463 gnd.n378 585
R4924 gnd.n5619 gnd.n5618 585
R4925 gnd.n5618 gnd.n5617 585
R4926 gnd.n5620 gnd.n5457 585
R4927 gnd.n5457 gnd.n387 585
R4928 gnd.n5622 gnd.n5621 585
R4929 gnd.n5622 gnd.n470 585
R4930 gnd.n5623 gnd.n5456 585
R4931 gnd.n5623 gnd.n424 585
R4932 gnd.n5625 gnd.n5624 585
R4933 gnd.n5624 gnd.n395 585
R4934 gnd.n5626 gnd.n1567 585
R4935 gnd.n1567 gnd.n1565 585
R4936 gnd.n5628 gnd.n5627 585
R4937 gnd.n5629 gnd.n5628 585
R4938 gnd.n1568 gnd.n1566 585
R4939 gnd.n1566 gnd.n1544 585
R4940 gnd.n5450 gnd.n5449 585
R4941 gnd.n5449 gnd.n1472 585
R4942 gnd.n5448 gnd.n1570 585
R4943 gnd.n5448 gnd.n1471 585
R4944 gnd.n5447 gnd.n1572 585
R4945 gnd.n5447 gnd.n5446 585
R4946 gnd.n5432 gnd.n1571 585
R4947 gnd.n1573 gnd.n1571 585
R4948 gnd.n5434 gnd.n5433 585
R4949 gnd.n5435 gnd.n5434 585
R4950 gnd.n1583 gnd.n1582 585
R4951 gnd.n1582 gnd.n1579 585
R4952 gnd.n5426 gnd.n5425 585
R4953 gnd.n5425 gnd.n5424 585
R4954 gnd.n1586 gnd.n1585 585
R4955 gnd.n1594 gnd.n1586 585
R4956 gnd.n5412 gnd.n5411 585
R4957 gnd.n5413 gnd.n5412 585
R4958 gnd.n1597 gnd.n1596 585
R4959 gnd.n1596 gnd.n1592 585
R4960 gnd.n5407 gnd.n5406 585
R4961 gnd.n5406 gnd.n5405 585
R4962 gnd.n1600 gnd.n1599 585
R4963 gnd.n1601 gnd.n1600 585
R4964 gnd.n5216 gnd.n5215 585
R4965 gnd.n5216 gnd.n1627 585
R4966 gnd.n5217 gnd.n5212 585
R4967 gnd.n5217 gnd.n1607 585
R4968 gnd.n5219 gnd.n5218 585
R4969 gnd.n5218 gnd.n1657 585
R4970 gnd.n5220 gnd.n1668 585
R4971 gnd.n1668 gnd.n1654 585
R4972 gnd.n5222 gnd.n5221 585
R4973 gnd.n5223 gnd.n5222 585
R4974 gnd.n1669 gnd.n1667 585
R4975 gnd.n1675 gnd.n1667 585
R4976 gnd.n5206 gnd.n5205 585
R4977 gnd.n5205 gnd.n5204 585
R4978 gnd.n1672 gnd.n1671 585
R4979 gnd.n1680 gnd.n1672 585
R4980 gnd.n5174 gnd.n1695 585
R4981 gnd.n1695 gnd.n1688 585
R4982 gnd.n5176 gnd.n5175 585
R4983 gnd.n5177 gnd.n5176 585
R4984 gnd.n1696 gnd.n1694 585
R4985 gnd.n4941 gnd.n1694 585
R4986 gnd.n5169 gnd.n5168 585
R4987 gnd.n5168 gnd.n5167 585
R4988 gnd.n1699 gnd.n1698 585
R4989 gnd.n5159 gnd.n1699 585
R4990 gnd.n5147 gnd.n5146 585
R4991 gnd.n5148 gnd.n5147 585
R4992 gnd.n1718 gnd.n1717 585
R4993 gnd.n4953 gnd.n1717 585
R4994 gnd.n5142 gnd.n5141 585
R4995 gnd.n5141 gnd.n5140 585
R4996 gnd.n1721 gnd.n1720 585
R4997 gnd.n5129 gnd.n1721 585
R4998 gnd.n5117 gnd.n5116 585
R4999 gnd.n5118 gnd.n5117 585
R5000 gnd.n1740 gnd.n1739 585
R5001 gnd.n4963 gnd.n1739 585
R5002 gnd.n5112 gnd.n5111 585
R5003 gnd.n5111 gnd.n5110 585
R5004 gnd.n1743 gnd.n1742 585
R5005 gnd.n5099 gnd.n1743 585
R5006 gnd.n5087 gnd.n5086 585
R5007 gnd.n5088 gnd.n5087 585
R5008 gnd.n1762 gnd.n1761 585
R5009 gnd.n1768 gnd.n1761 585
R5010 gnd.n5082 gnd.n5081 585
R5011 gnd.n5081 gnd.n5080 585
R5012 gnd.n1765 gnd.n1764 585
R5013 gnd.n1773 gnd.n1765 585
R5014 gnd.n5051 gnd.n1790 585
R5015 gnd.n1790 gnd.n1783 585
R5016 gnd.n5053 gnd.n5052 585
R5017 gnd.n5054 gnd.n5053 585
R5018 gnd.n1791 gnd.n1789 585
R5019 gnd.n4985 gnd.n1789 585
R5020 gnd.n5046 gnd.n5045 585
R5021 gnd.n5045 gnd.n5044 585
R5022 gnd.n1794 gnd.n1793 585
R5023 gnd.n5036 gnd.n1794 585
R5024 gnd.n5024 gnd.n5023 585
R5025 gnd.n5025 gnd.n5024 585
R5026 gnd.n1814 gnd.n1813 585
R5027 gnd.n4998 gnd.n1813 585
R5028 gnd.n5019 gnd.n5018 585
R5029 gnd.n5018 gnd.n5017 585
R5030 gnd.n1817 gnd.n1816 585
R5031 gnd.n5006 gnd.n1817 585
R5032 gnd.n4909 gnd.n4908 585
R5033 gnd.n4910 gnd.n4909 585
R5034 gnd.n1830 gnd.n1829 585
R5035 gnd.n4894 gnd.n1829 585
R5036 gnd.n4904 gnd.n4903 585
R5037 gnd.n4903 gnd.n4902 585
R5038 gnd.n1833 gnd.n1832 585
R5039 gnd.n1842 gnd.n1833 585
R5040 gnd.n4866 gnd.n4865 585
R5041 gnd.n4867 gnd.n4866 585
R5042 gnd.n1854 gnd.n1853 585
R5043 gnd.n1861 gnd.n1853 585
R5044 gnd.n4861 gnd.n4860 585
R5045 gnd.n4860 gnd.n4859 585
R5046 gnd.n1857 gnd.n1856 585
R5047 gnd.n1866 gnd.n1857 585
R5048 gnd.n4825 gnd.n1883 585
R5049 gnd.n1883 gnd.n1875 585
R5050 gnd.n4827 gnd.n4826 585
R5051 gnd.n4828 gnd.n4827 585
R5052 gnd.n1884 gnd.n1882 585
R5053 gnd.n4761 gnd.n1882 585
R5054 gnd.n4820 gnd.n4819 585
R5055 gnd.n4819 gnd.n4818 585
R5056 gnd.n1887 gnd.n1886 585
R5057 gnd.n4810 gnd.n1887 585
R5058 gnd.n4798 gnd.n4797 585
R5059 gnd.n4799 gnd.n4798 585
R5060 gnd.n1907 gnd.n1906 585
R5061 gnd.n4772 gnd.n1906 585
R5062 gnd.n4793 gnd.n4792 585
R5063 gnd.n4792 gnd.n4791 585
R5064 gnd.n1910 gnd.n1909 585
R5065 gnd.n4780 gnd.n1910 585
R5066 gnd.n4717 gnd.n4716 585
R5067 gnd.n4716 gnd.n1921 585
R5068 gnd.n4718 gnd.n1942 585
R5069 gnd.n1942 gnd.n1930 585
R5070 gnd.n4720 gnd.n4719 585
R5071 gnd.n4721 gnd.n4720 585
R5072 gnd.n1943 gnd.n1941 585
R5073 gnd.n1941 gnd.n1938 585
R5074 gnd.n4710 gnd.n4709 585
R5075 gnd.n4709 gnd.n4708 585
R5076 gnd.n1946 gnd.n1945 585
R5077 gnd.n1956 gnd.n1946 585
R5078 gnd.n4666 gnd.n4665 585
R5079 gnd.n4665 gnd.n4664 585
R5080 gnd.n4667 gnd.n2165 585
R5081 gnd.n2165 gnd.n2164 585
R5082 gnd.n4669 gnd.n4668 585
R5083 gnd.n4670 gnd.n4669 585
R5084 gnd.n2166 gnd.n2162 585
R5085 gnd.n4654 gnd.n2162 585
R5086 gnd.n4658 gnd.n4657 585
R5087 gnd.n4657 gnd.n4656 585
R5088 gnd.n2169 gnd.n2168 585
R5089 gnd.n2170 gnd.n2169 585
R5090 gnd.n4643 gnd.n4642 585
R5091 gnd.n4644 gnd.n4643 585
R5092 gnd.n2180 gnd.n2179 585
R5093 gnd.n2179 gnd.n2176 585
R5094 gnd.n4638 gnd.n4637 585
R5095 gnd.n4637 gnd.n4636 585
R5096 gnd.n2183 gnd.n2182 585
R5097 gnd.n2184 gnd.n2183 585
R5098 gnd.n4624 gnd.n4623 585
R5099 gnd.n4625 gnd.n4624 585
R5100 gnd.n2194 gnd.n2193 585
R5101 gnd.n2193 gnd.n2190 585
R5102 gnd.n4619 gnd.n4618 585
R5103 gnd.n4618 gnd.n4617 585
R5104 gnd.n2197 gnd.n2196 585
R5105 gnd.n2198 gnd.n2197 585
R5106 gnd.n4551 gnd.n2286 585
R5107 gnd.n2286 gnd.n2284 585
R5108 gnd.n4553 gnd.n4552 585
R5109 gnd.n4554 gnd.n4553 585
R5110 gnd.n2287 gnd.n2285 585
R5111 gnd.n2285 gnd.n2264 585
R5112 gnd.n4546 gnd.n4545 585
R5113 gnd.n4545 gnd.n4544 585
R5114 gnd.n4542 gnd.n2289 585
R5115 gnd.n4543 gnd.n4542 585
R5116 gnd.n4541 gnd.n4539 585
R5117 gnd.n4541 gnd.n4540 585
R5118 gnd.n2291 gnd.n2290 585
R5119 gnd.n2290 gnd.n1271 585
R5120 gnd.n4535 gnd.n4534 585
R5121 gnd.n4534 gnd.n1268 585
R5122 gnd.n4533 gnd.n2293 585
R5123 gnd.n4533 gnd.n1261 585
R5124 gnd.n4532 gnd.n4531 585
R5125 gnd.n4532 gnd.n1258 585
R5126 gnd.n2295 gnd.n2294 585
R5127 gnd.n2294 gnd.n1250 585
R5128 gnd.n4527 gnd.n4526 585
R5129 gnd.n4526 gnd.n1247 585
R5130 gnd.n4525 gnd.n2297 585
R5131 gnd.n4525 gnd.n1239 585
R5132 gnd.n4524 gnd.n2299 585
R5133 gnd.n4524 gnd.n4523 585
R5134 gnd.n4457 gnd.n2298 585
R5135 gnd.n2298 gnd.n1229 585
R5136 gnd.n4459 gnd.n4458 585
R5137 gnd.n4458 gnd.n1226 585
R5138 gnd.n4460 gnd.n4450 585
R5139 gnd.n4450 gnd.n1218 585
R5140 gnd.n4462 gnd.n4461 585
R5141 gnd.n4462 gnd.n1215 585
R5142 gnd.n4463 gnd.n4449 585
R5143 gnd.n4463 gnd.n2314 585
R5144 gnd.n4465 gnd.n4464 585
R5145 gnd.n4464 gnd.n1205 585
R5146 gnd.n4466 gnd.n2323 585
R5147 gnd.n2323 gnd.n1197 585
R5148 gnd.n4468 gnd.n4467 585
R5149 gnd.n4469 gnd.n4468 585
R5150 gnd.n2324 gnd.n2322 585
R5151 gnd.n2322 gnd.n1187 585
R5152 gnd.n4443 gnd.n4442 585
R5153 gnd.n4442 gnd.n1184 585
R5154 gnd.n4441 gnd.n2326 585
R5155 gnd.n4441 gnd.n1176 585
R5156 gnd.n4440 gnd.n4439 585
R5157 gnd.n4440 gnd.n1173 585
R5158 gnd.n2328 gnd.n2327 585
R5159 gnd.n4403 gnd.n2327 585
R5160 gnd.n4435 gnd.n4434 585
R5161 gnd.n4434 gnd.n1164 585
R5162 gnd.n4433 gnd.n2329 585
R5163 gnd.n4433 gnd.n1155 585
R5164 gnd.n4432 gnd.n2332 585
R5165 gnd.n4432 gnd.n4431 585
R5166 gnd.n4368 gnd.n2330 585
R5167 gnd.n2333 gnd.n2330 585
R5168 gnd.n4370 gnd.n2363 585
R5169 gnd.n2363 gnd.n2349 585
R5170 gnd.n4372 gnd.n4371 585
R5171 gnd.n4373 gnd.n4372 585
R5172 gnd.n4366 gnd.n2362 585
R5173 gnd.n2362 gnd.n2360 585
R5174 gnd.n4365 gnd.n4364 585
R5175 gnd.n4364 gnd.n4363 585
R5176 gnd.n4338 gnd.n2365 585
R5177 gnd.n2373 gnd.n2365 585
R5178 gnd.n4339 gnd.n2382 585
R5179 gnd.n2382 gnd.n2370 585
R5180 gnd.n4342 gnd.n4341 585
R5181 gnd.n4343 gnd.n4342 585
R5182 gnd.n4337 gnd.n2381 585
R5183 gnd.n2381 gnd.n2378 585
R5184 gnd.n2389 gnd.n2383 585
R5185 gnd.n2389 gnd.n1136 585
R5186 gnd.n4333 gnd.n4332 585
R5187 gnd.n4332 gnd.n4331 585
R5188 gnd.n2388 gnd.n2387 585
R5189 gnd.n2388 gnd.n1125 585
R5190 gnd.n2386 gnd.n1108 585
R5191 gnd.n1122 gnd.n1108 585
R5192 gnd.n5707 gnd.n5706 585
R5193 gnd.n5708 gnd.n5707 585
R5194 gnd.n1475 gnd.n1473 585
R5195 gnd.n5445 gnd.n1473 585
R5196 gnd.n5443 gnd.n5442 585
R5197 gnd.n5444 gnd.n5443 585
R5198 gnd.n1575 gnd.n1574 585
R5199 gnd.n1581 gnd.n1574 585
R5200 gnd.n5438 gnd.n5437 585
R5201 gnd.n5437 gnd.n5436 585
R5202 gnd.n1578 gnd.n1577 585
R5203 gnd.n5423 gnd.n1578 585
R5204 gnd.n5421 gnd.n5420 585
R5205 gnd.n5422 gnd.n5421 585
R5206 gnd.n1588 gnd.n1587 585
R5207 gnd.n1595 gnd.n1587 585
R5208 gnd.n5416 gnd.n5415 585
R5209 gnd.n5415 gnd.n5414 585
R5210 gnd.n1591 gnd.n1590 585
R5211 gnd.n5404 gnd.n1591 585
R5212 gnd.n5402 gnd.n5401 585
R5213 gnd.n5403 gnd.n5402 585
R5214 gnd.n1603 gnd.n1602 585
R5215 gnd.n1626 gnd.n1602 585
R5216 gnd.n5397 gnd.n5396 585
R5217 gnd.n5396 gnd.n5395 585
R5218 gnd.n1606 gnd.n1605 585
R5219 gnd.n1649 gnd.n1606 585
R5220 gnd.n5231 gnd.n5230 585
R5221 gnd.n5232 gnd.n5231 585
R5222 gnd.n1659 gnd.n1658 585
R5223 gnd.n1665 gnd.n1658 585
R5224 gnd.n5226 gnd.n5225 585
R5225 gnd.n5225 gnd.n5224 585
R5226 gnd.n1662 gnd.n1661 585
R5227 gnd.n5203 gnd.n1662 585
R5228 gnd.n5192 gnd.n5191 585
R5229 gnd.n5193 gnd.n5192 585
R5230 gnd.n1683 gnd.n1682 585
R5231 gnd.n4932 gnd.n1682 585
R5232 gnd.n5187 gnd.n5186 585
R5233 gnd.n5186 gnd.n5185 585
R5234 gnd.n1686 gnd.n1685 585
R5235 gnd.n1692 gnd.n1686 585
R5236 gnd.n1712 gnd.n1710 585
R5237 gnd.n1710 gnd.n1702 585
R5238 gnd.n5157 gnd.n5156 585
R5239 gnd.n5158 gnd.n5157 585
R5240 gnd.n1711 gnd.n1709 585
R5241 gnd.n1709 gnd.n1706 585
R5242 gnd.n5151 gnd.n5150 585
R5243 gnd.n5150 gnd.n5149 585
R5244 gnd.n1715 gnd.n1714 585
R5245 gnd.n1723 gnd.n1715 585
R5246 gnd.n5126 gnd.n5125 585
R5247 gnd.n5127 gnd.n5126 585
R5248 gnd.n1733 gnd.n1732 585
R5249 gnd.n1732 gnd.n1728 585
R5250 gnd.n5121 gnd.n5120 585
R5251 gnd.n5120 gnd.n5119 585
R5252 gnd.n1736 gnd.n1735 585
R5253 gnd.n1745 gnd.n1736 585
R5254 gnd.n5096 gnd.n5095 585
R5255 gnd.n5097 gnd.n5096 585
R5256 gnd.n1755 gnd.n1754 585
R5257 gnd.n1754 gnd.n1750 585
R5258 gnd.n5091 gnd.n5090 585
R5259 gnd.n5090 gnd.n5089 585
R5260 gnd.n1758 gnd.n1757 585
R5261 gnd.n5079 gnd.n1758 585
R5262 gnd.n5069 gnd.n5068 585
R5263 gnd.n5070 gnd.n5069 585
R5264 gnd.n1777 gnd.n1776 585
R5265 gnd.n4977 gnd.n1776 585
R5266 gnd.n5064 gnd.n5063 585
R5267 gnd.n5063 gnd.n5062 585
R5268 gnd.n1780 gnd.n1779 585
R5269 gnd.n1787 gnd.n1780 585
R5270 gnd.n1807 gnd.n1805 585
R5271 gnd.n1805 gnd.n1798 585
R5272 gnd.n5034 gnd.n5033 585
R5273 gnd.n5035 gnd.n5034 585
R5274 gnd.n1806 gnd.n1804 585
R5275 gnd.n1804 gnd.n1802 585
R5276 gnd.n5028 gnd.n5027 585
R5277 gnd.n5027 gnd.n5026 585
R5278 gnd.n1810 gnd.n1809 585
R5279 gnd.n4997 gnd.n1810 585
R5280 gnd.n4878 gnd.n4876 585
R5281 gnd.n4876 gnd.n1818 585
R5282 gnd.n4879 gnd.n4875 585
R5283 gnd.n4875 gnd.n1824 585
R5284 gnd.n4880 gnd.n4874 585
R5285 gnd.n4874 gnd.n1828 585
R5286 gnd.n1846 gnd.n1844 585
R5287 gnd.n1844 gnd.n1839 585
R5288 gnd.n4885 gnd.n4884 585
R5289 gnd.n4886 gnd.n4885 585
R5290 gnd.n1845 gnd.n1843 585
R5291 gnd.n4849 gnd.n1843 585
R5292 gnd.n4870 gnd.n4869 585
R5293 gnd.n4869 gnd.n4868 585
R5294 gnd.n1849 gnd.n1848 585
R5295 gnd.n4858 gnd.n1849 585
R5296 gnd.n4843 gnd.n4842 585
R5297 gnd.n4844 gnd.n4843 585
R5298 gnd.n1869 gnd.n1868 585
R5299 gnd.n4753 gnd.n1868 585
R5300 gnd.n4838 gnd.n4837 585
R5301 gnd.n4837 gnd.n4836 585
R5302 gnd.n1872 gnd.n1871 585
R5303 gnd.n1880 gnd.n1872 585
R5304 gnd.n1899 gnd.n1897 585
R5305 gnd.n1897 gnd.n1890 585
R5306 gnd.n4808 gnd.n4807 585
R5307 gnd.n4809 gnd.n4808 585
R5308 gnd.n1898 gnd.n1896 585
R5309 gnd.n1896 gnd.n1894 585
R5310 gnd.n4802 gnd.n4801 585
R5311 gnd.n4801 gnd.n4800 585
R5312 gnd.n1902 gnd.n1901 585
R5313 gnd.n1913 gnd.n1902 585
R5314 gnd.n1925 gnd.n1923 585
R5315 gnd.n1923 gnd.n1911 585
R5316 gnd.n4739 gnd.n4738 585
R5317 gnd.n4740 gnd.n4739 585
R5318 gnd.n1924 gnd.n1922 585
R5319 gnd.n1933 gnd.n1922 585
R5320 gnd.n4733 gnd.n4732 585
R5321 gnd.n4732 gnd.n4731 585
R5322 gnd.n1928 gnd.n1927 585
R5323 gnd.n4722 gnd.n1928 585
R5324 gnd.n4681 gnd.n4680 585
R5325 gnd.n4680 gnd.n4679 585
R5326 gnd.n4682 gnd.n4677 585
R5327 gnd.n4677 gnd.n1948 585
R5328 gnd.n1986 gnd.n1984 585
R5329 gnd.n1984 gnd.n1954 585
R5330 gnd.n4687 gnd.n4686 585
R5331 gnd.n4688 gnd.n4687 585
R5332 gnd.n1985 gnd.n1983 585
R5333 gnd.n2163 gnd.n1983 585
R5334 gnd.n4673 gnd.n4672 585
R5335 gnd.n4672 gnd.n4671 585
R5336 gnd.n1989 gnd.n1988 585
R5337 gnd.n4655 gnd.n1989 585
R5338 gnd.n4652 gnd.n4651 585
R5339 gnd.n4653 gnd.n4652 585
R5340 gnd.n2172 gnd.n2171 585
R5341 gnd.n2178 gnd.n2171 585
R5342 gnd.n4647 gnd.n4646 585
R5343 gnd.n4646 gnd.n4645 585
R5344 gnd.n2175 gnd.n2174 585
R5345 gnd.n4635 gnd.n2175 585
R5346 gnd.n4633 gnd.n4632 585
R5347 gnd.n4634 gnd.n4633 585
R5348 gnd.n2186 gnd.n2185 585
R5349 gnd.n2192 gnd.n2185 585
R5350 gnd.n4628 gnd.n4627 585
R5351 gnd.n4627 gnd.n4626 585
R5352 gnd.n2189 gnd.n2188 585
R5353 gnd.n4616 gnd.n2189 585
R5354 gnd.n4614 gnd.n4613 585
R5355 gnd.n4615 gnd.n4614 585
R5356 gnd.n2200 gnd.n2199 585
R5357 gnd.n2283 gnd.n2199 585
R5358 gnd.n4555 gnd.n2208 585
R5359 gnd.n4603 gnd.n2209 585
R5360 gnd.n4602 gnd.n2210 585
R5361 gnd.n4557 gnd.n2210 585
R5362 gnd.n2265 gnd.n2211 585
R5363 gnd.n4595 gnd.n2219 585
R5364 gnd.n4594 gnd.n2220 585
R5365 gnd.n2267 gnd.n2221 585
R5366 gnd.n4587 gnd.n2230 585
R5367 gnd.n4586 gnd.n2231 585
R5368 gnd.n2270 gnd.n2232 585
R5369 gnd.n4579 gnd.n2240 585
R5370 gnd.n4578 gnd.n2241 585
R5371 gnd.n2272 gnd.n2242 585
R5372 gnd.n4571 gnd.n2251 585
R5373 gnd.n4570 gnd.n2252 585
R5374 gnd.n2263 gnd.n2253 585
R5375 gnd.n4560 gnd.n4559 585
R5376 gnd.n2262 gnd.n1349 585
R5377 gnd.n5849 gnd.n1350 585
R5378 gnd.n5848 gnd.n1351 585
R5379 gnd.n5847 gnd.n1352 585
R5380 gnd.n2277 gnd.n1353 585
R5381 gnd.n5843 gnd.n1355 585
R5382 gnd.n5842 gnd.n1356 585
R5383 gnd.n5841 gnd.n1357 585
R5384 gnd.n5838 gnd.n1362 585
R5385 gnd.n5837 gnd.n1363 585
R5386 gnd.n5836 gnd.n1364 585
R5387 gnd.n2281 gnd.n1365 585
R5388 gnd.n5710 gnd.n5709 585
R5389 gnd.n5709 gnd.n5708 585
R5390 gnd.n5711 gnd.n1468 585
R5391 gnd.n5445 gnd.n1468 585
R5392 gnd.n5712 gnd.n1467 585
R5393 gnd.n5444 gnd.n1467 585
R5394 gnd.n1580 gnd.n1465 585
R5395 gnd.n1581 gnd.n1580 585
R5396 gnd.n5716 gnd.n1464 585
R5397 gnd.n5436 gnd.n1464 585
R5398 gnd.n5717 gnd.n1463 585
R5399 gnd.n5423 gnd.n1463 585
R5400 gnd.n5718 gnd.n1462 585
R5401 gnd.n5422 gnd.n1462 585
R5402 gnd.n1593 gnd.n1460 585
R5403 gnd.n1595 gnd.n1593 585
R5404 gnd.n5722 gnd.n1459 585
R5405 gnd.n5414 gnd.n1459 585
R5406 gnd.n5723 gnd.n1458 585
R5407 gnd.n5404 gnd.n1458 585
R5408 gnd.n5724 gnd.n1457 585
R5409 gnd.n5403 gnd.n1457 585
R5410 gnd.n1625 gnd.n1455 585
R5411 gnd.n1626 gnd.n1625 585
R5412 gnd.n5728 gnd.n1454 585
R5413 gnd.n5395 gnd.n1454 585
R5414 gnd.n5729 gnd.n1453 585
R5415 gnd.n1649 gnd.n1453 585
R5416 gnd.n5730 gnd.n1452 585
R5417 gnd.n5232 gnd.n1452 585
R5418 gnd.n1664 gnd.n1450 585
R5419 gnd.n1665 gnd.n1664 585
R5420 gnd.n5734 gnd.n1449 585
R5421 gnd.n5224 gnd.n1449 585
R5422 gnd.n5735 gnd.n1448 585
R5423 gnd.n5203 gnd.n1448 585
R5424 gnd.n5736 gnd.n1447 585
R5425 gnd.n5193 gnd.n1447 585
R5426 gnd.n4931 gnd.n1445 585
R5427 gnd.n4932 gnd.n4931 585
R5428 gnd.n5740 gnd.n1444 585
R5429 gnd.n5185 gnd.n1444 585
R5430 gnd.n5741 gnd.n1443 585
R5431 gnd.n1692 gnd.n1443 585
R5432 gnd.n5742 gnd.n1442 585
R5433 gnd.n1702 gnd.n1442 585
R5434 gnd.n1708 gnd.n1440 585
R5435 gnd.n5158 gnd.n1708 585
R5436 gnd.n5746 gnd.n1439 585
R5437 gnd.n1706 gnd.n1439 585
R5438 gnd.n5747 gnd.n1438 585
R5439 gnd.n5149 gnd.n1438 585
R5440 gnd.n5748 gnd.n1437 585
R5441 gnd.n1723 gnd.n1437 585
R5442 gnd.n1731 gnd.n1435 585
R5443 gnd.n5127 gnd.n1731 585
R5444 gnd.n5752 gnd.n1434 585
R5445 gnd.n1728 gnd.n1434 585
R5446 gnd.n5753 gnd.n1433 585
R5447 gnd.n5119 gnd.n1433 585
R5448 gnd.n5754 gnd.n1432 585
R5449 gnd.n1745 gnd.n1432 585
R5450 gnd.n1753 gnd.n1430 585
R5451 gnd.n5097 gnd.n1753 585
R5452 gnd.n5758 gnd.n1429 585
R5453 gnd.n1750 gnd.n1429 585
R5454 gnd.n5759 gnd.n1428 585
R5455 gnd.n5089 gnd.n1428 585
R5456 gnd.n5760 gnd.n1427 585
R5457 gnd.n5079 gnd.n1427 585
R5458 gnd.n1775 gnd.n1425 585
R5459 gnd.n5070 gnd.n1775 585
R5460 gnd.n5764 gnd.n1424 585
R5461 gnd.n4977 gnd.n1424 585
R5462 gnd.n5765 gnd.n1423 585
R5463 gnd.n5062 gnd.n1423 585
R5464 gnd.n5766 gnd.n1422 585
R5465 gnd.n1787 gnd.n1422 585
R5466 gnd.n1797 gnd.n1420 585
R5467 gnd.n1798 gnd.n1797 585
R5468 gnd.n5770 gnd.n1419 585
R5469 gnd.n5035 gnd.n1419 585
R5470 gnd.n5771 gnd.n1418 585
R5471 gnd.n1802 gnd.n1418 585
R5472 gnd.n5772 gnd.n1417 585
R5473 gnd.n5026 gnd.n1417 585
R5474 gnd.n4996 gnd.n1415 585
R5475 gnd.n4997 gnd.n4996 585
R5476 gnd.n5776 gnd.n1414 585
R5477 gnd.n1818 gnd.n1414 585
R5478 gnd.n5777 gnd.n1413 585
R5479 gnd.n1824 gnd.n1413 585
R5480 gnd.n5778 gnd.n1412 585
R5481 gnd.n1828 gnd.n1412 585
R5482 gnd.n1838 gnd.n1410 585
R5483 gnd.n1839 gnd.n1838 585
R5484 gnd.n5782 gnd.n1409 585
R5485 gnd.n4886 gnd.n1409 585
R5486 gnd.n5783 gnd.n1408 585
R5487 gnd.n4849 gnd.n1408 585
R5488 gnd.n5784 gnd.n1407 585
R5489 gnd.n4868 gnd.n1407 585
R5490 gnd.n1859 gnd.n1405 585
R5491 gnd.n4858 gnd.n1859 585
R5492 gnd.n5788 gnd.n1404 585
R5493 gnd.n4844 gnd.n1404 585
R5494 gnd.n5789 gnd.n1403 585
R5495 gnd.n4753 gnd.n1403 585
R5496 gnd.n5790 gnd.n1402 585
R5497 gnd.n4836 gnd.n1402 585
R5498 gnd.n1879 gnd.n1400 585
R5499 gnd.n1880 gnd.n1879 585
R5500 gnd.n5794 gnd.n1399 585
R5501 gnd.n1890 gnd.n1399 585
R5502 gnd.n5795 gnd.n1398 585
R5503 gnd.n4809 gnd.n1398 585
R5504 gnd.n5796 gnd.n1397 585
R5505 gnd.n1894 gnd.n1397 585
R5506 gnd.n1904 gnd.n1395 585
R5507 gnd.n4800 gnd.n1904 585
R5508 gnd.n5800 gnd.n1394 585
R5509 gnd.n1913 gnd.n1394 585
R5510 gnd.n5801 gnd.n1393 585
R5511 gnd.n1911 gnd.n1393 585
R5512 gnd.n5802 gnd.n1392 585
R5513 gnd.n4740 gnd.n1392 585
R5514 gnd.n1932 gnd.n1390 585
R5515 gnd.n1933 gnd.n1932 585
R5516 gnd.n5806 gnd.n1389 585
R5517 gnd.n4731 gnd.n1389 585
R5518 gnd.n5807 gnd.n1388 585
R5519 gnd.n4722 gnd.n1388 585
R5520 gnd.n5808 gnd.n1387 585
R5521 gnd.n4679 gnd.n1387 585
R5522 gnd.n1947 gnd.n1385 585
R5523 gnd.n1948 gnd.n1947 585
R5524 gnd.n5812 gnd.n1384 585
R5525 gnd.n1954 gnd.n1384 585
R5526 gnd.n5813 gnd.n1383 585
R5527 gnd.n4688 gnd.n1383 585
R5528 gnd.n5814 gnd.n1382 585
R5529 gnd.n2163 gnd.n1382 585
R5530 gnd.n1990 gnd.n1380 585
R5531 gnd.n4671 gnd.n1990 585
R5532 gnd.n5818 gnd.n1379 585
R5533 gnd.n4655 gnd.n1379 585
R5534 gnd.n5819 gnd.n1378 585
R5535 gnd.n4653 gnd.n1378 585
R5536 gnd.n5820 gnd.n1377 585
R5537 gnd.n2178 gnd.n1377 585
R5538 gnd.n2177 gnd.n1375 585
R5539 gnd.n4645 gnd.n2177 585
R5540 gnd.n5824 gnd.n1374 585
R5541 gnd.n4635 gnd.n1374 585
R5542 gnd.n5825 gnd.n1373 585
R5543 gnd.n4634 gnd.n1373 585
R5544 gnd.n5826 gnd.n1372 585
R5545 gnd.n2192 gnd.n1372 585
R5546 gnd.n2191 gnd.n1370 585
R5547 gnd.n4626 gnd.n2191 585
R5548 gnd.n5830 gnd.n1369 585
R5549 gnd.n4616 gnd.n1369 585
R5550 gnd.n5831 gnd.n1368 585
R5551 gnd.n4615 gnd.n1368 585
R5552 gnd.n5832 gnd.n1367 585
R5553 gnd.n2283 gnd.n1367 585
R5554 gnd.n5633 gnd.n1470 585
R5555 gnd.n5630 gnd.n1470 585
R5556 gnd.n5636 gnd.n5632 585
R5557 gnd.n5637 gnd.n1543 585
R5558 gnd.n5638 gnd.n1542 585
R5559 gnd.n1563 gnd.n1537 585
R5560 gnd.n5642 gnd.n1536 585
R5561 gnd.n5643 gnd.n1535 585
R5562 gnd.n5644 gnd.n1534 585
R5563 gnd.n1560 gnd.n1532 585
R5564 gnd.n5648 gnd.n1531 585
R5565 gnd.n5649 gnd.n1530 585
R5566 gnd.n5652 gnd.n1529 585
R5567 gnd.n5653 gnd.n1528 585
R5568 gnd.n1556 gnd.n1522 585
R5569 gnd.n5663 gnd.n1521 585
R5570 gnd.n5664 gnd.n1520 585
R5571 gnd.n1554 gnd.n1514 585
R5572 gnd.n5671 gnd.n1513 585
R5573 gnd.n5672 gnd.n1512 585
R5574 gnd.n1551 gnd.n1504 585
R5575 gnd.n5679 gnd.n1503 585
R5576 gnd.n5680 gnd.n1502 585
R5577 gnd.n1549 gnd.n1496 585
R5578 gnd.n5687 gnd.n1495 585
R5579 gnd.n5688 gnd.n1494 585
R5580 gnd.n1546 gnd.n1486 585
R5581 gnd.n5695 gnd.n1485 585
R5582 gnd.n5696 gnd.n1484 585
R5583 gnd.n1483 gnd.n1474 585
R5584 gnd.n6189 gnd.n937 493.813
R5585 gnd.n5325 gnd.n1651 473.281
R5586 gnd.n5328 gnd.n5327 473.281
R5587 gnd.n2031 gnd.n1981 473.281
R5588 gnd.n4690 gnd.n1980 473.281
R5589 gnd.n2028 gnd.t110 443.966
R5590 gnd.n1645 gnd.t24 443.966
R5591 gnd.n2025 gnd.t42 443.966
R5592 gnd.n5256 gnd.t104 443.966
R5593 gnd.n1358 gnd.t90 371.625
R5594 gnd.n7211 gnd.t17 371.625
R5595 gnd.n5657 gnd.t56 371.625
R5596 gnd.n2258 gnd.t87 371.625
R5597 gnd.n443 gnd.t53 371.625
R5598 gnd.n465 gnd.t31 371.625
R5599 gnd.n175 gnd.t119 371.625
R5600 gnd.n7290 gnd.t35 371.625
R5601 gnd.n3950 gnd.t116 371.625
R5602 gnd.n3926 gnd.t107 371.625
R5603 gnd.n1337 gnd.t49 371.625
R5604 gnd.n1300 gnd.t70 371.625
R5605 gnd.n4121 gnd.t63 371.625
R5606 gnd.n1539 gnd.t73 371.625
R5607 gnd.n2939 gnd.t38 323.425
R5608 gnd.n2496 gnd.t80 323.425
R5609 gnd.n3787 gnd.n3761 289.615
R5610 gnd.n3755 gnd.n3729 289.615
R5611 gnd.n3723 gnd.n3697 289.615
R5612 gnd.n3692 gnd.n3666 289.615
R5613 gnd.n3660 gnd.n3634 289.615
R5614 gnd.n3628 gnd.n3602 289.615
R5615 gnd.n3596 gnd.n3570 289.615
R5616 gnd.n3565 gnd.n3539 289.615
R5617 gnd.n3013 gnd.t59 279.217
R5618 gnd.n2522 gnd.t100 279.217
R5619 gnd.n1965 gnd.t30 260.649
R5620 gnd.n5248 gnd.t79 260.649
R5621 gnd.n2161 gnd.n2160 256.663
R5622 gnd.n2161 gnd.n1991 256.663
R5623 gnd.n2161 gnd.n1992 256.663
R5624 gnd.n2161 gnd.n1993 256.663
R5625 gnd.n2161 gnd.n1994 256.663
R5626 gnd.n2161 gnd.n1995 256.663
R5627 gnd.n2161 gnd.n1996 256.663
R5628 gnd.n2161 gnd.n1997 256.663
R5629 gnd.n2161 gnd.n1998 256.663
R5630 gnd.n2161 gnd.n1999 256.663
R5631 gnd.n2161 gnd.n2000 256.663
R5632 gnd.n2161 gnd.n2001 256.663
R5633 gnd.n2161 gnd.n2002 256.663
R5634 gnd.n2161 gnd.n2003 256.663
R5635 gnd.n2161 gnd.n2004 256.663
R5636 gnd.n2161 gnd.n2005 256.663
R5637 gnd.n2098 gnd.n2095 256.663
R5638 gnd.n2161 gnd.n2006 256.663
R5639 gnd.n2161 gnd.n2007 256.663
R5640 gnd.n2161 gnd.n2008 256.663
R5641 gnd.n2161 gnd.n2009 256.663
R5642 gnd.n2161 gnd.n2010 256.663
R5643 gnd.n2161 gnd.n2011 256.663
R5644 gnd.n2161 gnd.n2012 256.663
R5645 gnd.n2161 gnd.n2013 256.663
R5646 gnd.n2161 gnd.n2014 256.663
R5647 gnd.n2161 gnd.n2015 256.663
R5648 gnd.n2161 gnd.n2016 256.663
R5649 gnd.n2161 gnd.n2017 256.663
R5650 gnd.n2161 gnd.n2018 256.663
R5651 gnd.n2161 gnd.n2019 256.663
R5652 gnd.n2161 gnd.n2020 256.663
R5653 gnd.n2161 gnd.n2021 256.663
R5654 gnd.n2161 gnd.n2022 256.663
R5655 gnd.n5394 gnd.n1628 256.663
R5656 gnd.n5394 gnd.n1629 256.663
R5657 gnd.n5394 gnd.n1630 256.663
R5658 gnd.n5394 gnd.n1631 256.663
R5659 gnd.n5394 gnd.n1632 256.663
R5660 gnd.n5394 gnd.n1633 256.663
R5661 gnd.n5394 gnd.n1634 256.663
R5662 gnd.n5394 gnd.n1635 256.663
R5663 gnd.n5394 gnd.n1636 256.663
R5664 gnd.n5394 gnd.n1637 256.663
R5665 gnd.n5394 gnd.n1638 256.663
R5666 gnd.n5394 gnd.n1639 256.663
R5667 gnd.n5394 gnd.n1640 256.663
R5668 gnd.n5394 gnd.n1641 256.663
R5669 gnd.n5394 gnd.n1642 256.663
R5670 gnd.n5394 gnd.n1643 256.663
R5671 gnd.n1644 gnd.n440 256.663
R5672 gnd.n5394 gnd.n1624 256.663
R5673 gnd.n5394 gnd.n1623 256.663
R5674 gnd.n5394 gnd.n1622 256.663
R5675 gnd.n5394 gnd.n1621 256.663
R5676 gnd.n5394 gnd.n1620 256.663
R5677 gnd.n5394 gnd.n1619 256.663
R5678 gnd.n5394 gnd.n1618 256.663
R5679 gnd.n5394 gnd.n1617 256.663
R5680 gnd.n5394 gnd.n1616 256.663
R5681 gnd.n5394 gnd.n1615 256.663
R5682 gnd.n5394 gnd.n1614 256.663
R5683 gnd.n5394 gnd.n1613 256.663
R5684 gnd.n5394 gnd.n1612 256.663
R5685 gnd.n5394 gnd.n1611 256.663
R5686 gnd.n5394 gnd.n1610 256.663
R5687 gnd.n5394 gnd.n1609 256.663
R5688 gnd.n5394 gnd.n1608 256.663
R5689 gnd.n4206 gnd.n3920 242.672
R5690 gnd.n4204 gnd.n3920 242.672
R5691 gnd.n4198 gnd.n3920 242.672
R5692 gnd.n4196 gnd.n3920 242.672
R5693 gnd.n4190 gnd.n3920 242.672
R5694 gnd.n4188 gnd.n3920 242.672
R5695 gnd.n4182 gnd.n3920 242.672
R5696 gnd.n4180 gnd.n3920 242.672
R5697 gnd.n4170 gnd.n3920 242.672
R5698 gnd.n4563 gnd.n1276 242.672
R5699 gnd.n2256 gnd.n1276 242.672
R5700 gnd.n2247 gnd.n1276 242.672
R5701 gnd.n2244 gnd.n1276 242.672
R5702 gnd.n2235 gnd.n1276 242.672
R5703 gnd.n2226 gnd.n1276 242.672
R5704 gnd.n2223 gnd.n1276 242.672
R5705 gnd.n2214 gnd.n1276 242.672
R5706 gnd.n2203 gnd.n1276 242.672
R5707 gnd.n6966 gnd.n414 242.672
R5708 gnd.n6966 gnd.n415 242.672
R5709 gnd.n6966 gnd.n416 242.672
R5710 gnd.n6966 gnd.n417 242.672
R5711 gnd.n6966 gnd.n418 242.672
R5712 gnd.n6966 gnd.n419 242.672
R5713 gnd.n6966 gnd.n420 242.672
R5714 gnd.n6966 gnd.n421 242.672
R5715 gnd.n6966 gnd.n422 242.672
R5716 gnd.n7213 gnd.n102 242.672
R5717 gnd.n7209 gnd.n102 242.672
R5718 gnd.n7204 gnd.n102 242.672
R5719 gnd.n7201 gnd.n102 242.672
R5720 gnd.n7196 gnd.n102 242.672
R5721 gnd.n7193 gnd.n102 242.672
R5722 gnd.n7188 gnd.n102 242.672
R5723 gnd.n7185 gnd.n102 242.672
R5724 gnd.n7180 gnd.n102 242.672
R5725 gnd.n3067 gnd.n3066 242.672
R5726 gnd.n3067 gnd.n2977 242.672
R5727 gnd.n3067 gnd.n2978 242.672
R5728 gnd.n3067 gnd.n2979 242.672
R5729 gnd.n3067 gnd.n2980 242.672
R5730 gnd.n3067 gnd.n2981 242.672
R5731 gnd.n3067 gnd.n2982 242.672
R5732 gnd.n3067 gnd.n2983 242.672
R5733 gnd.n3067 gnd.n2984 242.672
R5734 gnd.n3067 gnd.n2985 242.672
R5735 gnd.n3067 gnd.n2986 242.672
R5736 gnd.n3067 gnd.n2987 242.672
R5737 gnd.n3068 gnd.n3067 242.672
R5738 gnd.n3919 gnd.n2471 242.672
R5739 gnd.n3919 gnd.n2470 242.672
R5740 gnd.n3919 gnd.n2469 242.672
R5741 gnd.n3919 gnd.n2468 242.672
R5742 gnd.n3919 gnd.n2467 242.672
R5743 gnd.n3919 gnd.n2466 242.672
R5744 gnd.n3919 gnd.n2465 242.672
R5745 gnd.n3919 gnd.n2464 242.672
R5746 gnd.n3919 gnd.n2463 242.672
R5747 gnd.n3919 gnd.n2462 242.672
R5748 gnd.n3919 gnd.n2461 242.672
R5749 gnd.n3919 gnd.n2460 242.672
R5750 gnd.n3919 gnd.n2459 242.672
R5751 gnd.n3151 gnd.n3150 242.672
R5752 gnd.n3150 gnd.n2889 242.672
R5753 gnd.n3150 gnd.n2890 242.672
R5754 gnd.n3150 gnd.n2891 242.672
R5755 gnd.n3150 gnd.n2892 242.672
R5756 gnd.n3150 gnd.n2893 242.672
R5757 gnd.n3150 gnd.n2894 242.672
R5758 gnd.n3150 gnd.n2895 242.672
R5759 gnd.n3919 gnd.n2472 242.672
R5760 gnd.n3919 gnd.n2473 242.672
R5761 gnd.n3919 gnd.n2474 242.672
R5762 gnd.n3919 gnd.n2475 242.672
R5763 gnd.n3919 gnd.n2476 242.672
R5764 gnd.n3919 gnd.n2477 242.672
R5765 gnd.n3919 gnd.n2478 242.672
R5766 gnd.n3919 gnd.n2479 242.672
R5767 gnd.n3968 gnd.n3920 242.672
R5768 gnd.n3976 gnd.n3920 242.672
R5769 gnd.n3978 gnd.n3920 242.672
R5770 gnd.n3986 gnd.n3920 242.672
R5771 gnd.n3988 gnd.n3920 242.672
R5772 gnd.n3996 gnd.n3920 242.672
R5773 gnd.n3998 gnd.n3920 242.672
R5774 gnd.n4006 gnd.n3920 242.672
R5775 gnd.n4008 gnd.n3920 242.672
R5776 gnd.n4016 gnd.n3920 242.672
R5777 gnd.n4018 gnd.n3920 242.672
R5778 gnd.n4026 gnd.n3920 242.672
R5779 gnd.n4028 gnd.n3920 242.672
R5780 gnd.n4036 gnd.n3920 242.672
R5781 gnd.n4038 gnd.n3920 242.672
R5782 gnd.n4046 gnd.n3920 242.672
R5783 gnd.n4048 gnd.n3920 242.672
R5784 gnd.n4057 gnd.n3920 242.672
R5785 gnd.n4060 gnd.n3920 242.672
R5786 gnd.n5864 gnd.n1276 242.672
R5787 gnd.n1340 gnd.n1276 242.672
R5788 gnd.n5871 gnd.n1276 242.672
R5789 gnd.n1331 gnd.n1276 242.672
R5790 gnd.n5878 gnd.n1276 242.672
R5791 gnd.n1324 gnd.n1276 242.672
R5792 gnd.n5885 gnd.n1276 242.672
R5793 gnd.n1317 gnd.n1276 242.672
R5794 gnd.n5892 gnd.n1276 242.672
R5795 gnd.n1310 gnd.n1276 242.672
R5796 gnd.n5899 gnd.n1276 242.672
R5797 gnd.n5900 gnd.n1302 242.672
R5798 gnd.n5901 gnd.n1276 242.672
R5799 gnd.n1299 gnd.n1276 242.672
R5800 gnd.n5908 gnd.n1276 242.672
R5801 gnd.n1292 gnd.n1276 242.672
R5802 gnd.n5915 gnd.n1276 242.672
R5803 gnd.n1285 gnd.n1276 242.672
R5804 gnd.n5922 gnd.n1276 242.672
R5805 gnd.n5925 gnd.n1276 242.672
R5806 gnd.n6967 gnd.n6966 242.672
R5807 gnd.n6966 gnd.n396 242.672
R5808 gnd.n6966 gnd.n397 242.672
R5809 gnd.n6966 gnd.n398 242.672
R5810 gnd.n6966 gnd.n399 242.672
R5811 gnd.n6966 gnd.n400 242.672
R5812 gnd.n6966 gnd.n401 242.672
R5813 gnd.n6966 gnd.n402 242.672
R5814 gnd.n6938 gnd.n441 242.672
R5815 gnd.n6966 gnd.n403 242.672
R5816 gnd.n6966 gnd.n404 242.672
R5817 gnd.n6966 gnd.n405 242.672
R5818 gnd.n6966 gnd.n406 242.672
R5819 gnd.n6966 gnd.n407 242.672
R5820 gnd.n6966 gnd.n408 242.672
R5821 gnd.n6966 gnd.n409 242.672
R5822 gnd.n6966 gnd.n410 242.672
R5823 gnd.n6966 gnd.n411 242.672
R5824 gnd.n6966 gnd.n412 242.672
R5825 gnd.n6966 gnd.n413 242.672
R5826 gnd.n172 gnd.n102 242.672
R5827 gnd.n7258 gnd.n102 242.672
R5828 gnd.n168 gnd.n102 242.672
R5829 gnd.n7265 gnd.n102 242.672
R5830 gnd.n161 gnd.n102 242.672
R5831 gnd.n7272 gnd.n102 242.672
R5832 gnd.n154 gnd.n102 242.672
R5833 gnd.n7279 gnd.n102 242.672
R5834 gnd.n147 gnd.n102 242.672
R5835 gnd.n7286 gnd.n102 242.672
R5836 gnd.n140 gnd.n102 242.672
R5837 gnd.n7296 gnd.n102 242.672
R5838 gnd.n133 gnd.n102 242.672
R5839 gnd.n7303 gnd.n102 242.672
R5840 gnd.n126 gnd.n102 242.672
R5841 gnd.n7310 gnd.n102 242.672
R5842 gnd.n119 gnd.n102 242.672
R5843 gnd.n7317 gnd.n102 242.672
R5844 gnd.n112 gnd.n102 242.672
R5845 gnd.n4557 gnd.n4556 242.672
R5846 gnd.n4557 gnd.n2266 242.672
R5847 gnd.n4557 gnd.n2268 242.672
R5848 gnd.n4557 gnd.n2269 242.672
R5849 gnd.n4557 gnd.n2271 242.672
R5850 gnd.n4557 gnd.n2273 242.672
R5851 gnd.n4557 gnd.n2274 242.672
R5852 gnd.n4558 gnd.n4557 242.672
R5853 gnd.n4557 gnd.n2275 242.672
R5854 gnd.n4557 gnd.n2276 242.672
R5855 gnd.n4557 gnd.n2278 242.672
R5856 gnd.n4557 gnd.n2279 242.672
R5857 gnd.n4557 gnd.n2280 242.672
R5858 gnd.n4557 gnd.n2282 242.672
R5859 gnd.n5631 gnd.n5630 242.672
R5860 gnd.n5630 gnd.n1564 242.672
R5861 gnd.n5630 gnd.n1562 242.672
R5862 gnd.n5630 gnd.n1561 242.672
R5863 gnd.n5630 gnd.n1559 242.672
R5864 gnd.n5630 gnd.n1558 242.672
R5865 gnd.n5630 gnd.n1557 242.672
R5866 gnd.n5630 gnd.n1555 242.672
R5867 gnd.n5630 gnd.n1553 242.672
R5868 gnd.n5630 gnd.n1552 242.672
R5869 gnd.n5630 gnd.n1550 242.672
R5870 gnd.n5630 gnd.n1548 242.672
R5871 gnd.n5630 gnd.n1547 242.672
R5872 gnd.n5630 gnd.n1545 242.672
R5873 gnd.n109 gnd.n105 240.244
R5874 gnd.n7319 gnd.n7318 240.244
R5875 gnd.n7316 gnd.n113 240.244
R5876 gnd.n7312 gnd.n7311 240.244
R5877 gnd.n7309 gnd.n120 240.244
R5878 gnd.n7305 gnd.n7304 240.244
R5879 gnd.n7302 gnd.n127 240.244
R5880 gnd.n7298 gnd.n7297 240.244
R5881 gnd.n7295 gnd.n134 240.244
R5882 gnd.n7288 gnd.n7287 240.244
R5883 gnd.n7285 gnd.n141 240.244
R5884 gnd.n7281 gnd.n7280 240.244
R5885 gnd.n7278 gnd.n148 240.244
R5886 gnd.n7274 gnd.n7273 240.244
R5887 gnd.n7271 gnd.n155 240.244
R5888 gnd.n7267 gnd.n7266 240.244
R5889 gnd.n7264 gnd.n162 240.244
R5890 gnd.n7260 gnd.n7259 240.244
R5891 gnd.n7257 gnd.n169 240.244
R5892 gnd.n6895 gnd.n388 240.244
R5893 gnd.n5615 gnd.n388 240.244
R5894 gnd.n5615 gnd.n379 240.244
R5895 gnd.n5611 gnd.n379 240.244
R5896 gnd.n5611 gnd.n370 240.244
R5897 gnd.n5607 gnd.n370 240.244
R5898 gnd.n5607 gnd.n361 240.244
R5899 gnd.n5603 gnd.n361 240.244
R5900 gnd.n5603 gnd.n353 240.244
R5901 gnd.n5599 gnd.n353 240.244
R5902 gnd.n5599 gnd.n344 240.244
R5903 gnd.n5513 gnd.n344 240.244
R5904 gnd.n5513 gnd.n335 240.244
R5905 gnd.n5519 gnd.n335 240.244
R5906 gnd.n5519 gnd.n326 240.244
R5907 gnd.n5523 gnd.n326 240.244
R5908 gnd.n5523 gnd.n318 240.244
R5909 gnd.n5581 gnd.n318 240.244
R5910 gnd.n5581 gnd.n307 240.244
R5911 gnd.n5577 gnd.n307 240.244
R5912 gnd.n5577 gnd.n5531 240.244
R5913 gnd.n5531 gnd.n298 240.244
R5914 gnd.n5553 gnd.n298 240.244
R5915 gnd.n5553 gnd.n289 240.244
R5916 gnd.n6850 gnd.n289 240.244
R5917 gnd.n6850 gnd.n282 240.244
R5918 gnd.n6846 gnd.n282 240.244
R5919 gnd.n6846 gnd.n273 240.244
R5920 gnd.n6842 gnd.n273 240.244
R5921 gnd.n6842 gnd.n267 240.244
R5922 gnd.n6838 gnd.n267 240.244
R5923 gnd.n6838 gnd.n259 240.244
R5924 gnd.n550 gnd.n259 240.244
R5925 gnd.n550 gnd.n250 240.244
R5926 gnd.n546 gnd.n250 240.244
R5927 gnd.n546 gnd.n242 240.244
R5928 gnd.n542 gnd.n242 240.244
R5929 gnd.n542 gnd.n234 240.244
R5930 gnd.n539 gnd.n234 240.244
R5931 gnd.n539 gnd.n226 240.244
R5932 gnd.n536 gnd.n226 240.244
R5933 gnd.n536 gnd.n217 240.244
R5934 gnd.n533 gnd.n217 240.244
R5935 gnd.n533 gnd.n211 240.244
R5936 gnd.n530 gnd.n211 240.244
R5937 gnd.n530 gnd.n204 240.244
R5938 gnd.n527 gnd.n204 240.244
R5939 gnd.n527 gnd.n197 240.244
R5940 gnd.n524 gnd.n197 240.244
R5941 gnd.n524 gnd.n187 240.244
R5942 gnd.n187 gnd.n179 240.244
R5943 gnd.n7249 gnd.n179 240.244
R5944 gnd.n7249 gnd.n101 240.244
R5945 gnd.n6965 gnd.n394 240.244
R5946 gnd.n6965 gnd.n425 240.244
R5947 gnd.n6961 gnd.n6960 240.244
R5948 gnd.n6957 gnd.n6956 240.244
R5949 gnd.n6953 gnd.n6952 240.244
R5950 gnd.n6949 gnd.n6948 240.244
R5951 gnd.n6945 gnd.n6944 240.244
R5952 gnd.n6941 gnd.n6940 240.244
R5953 gnd.n6936 gnd.n6935 240.244
R5954 gnd.n6932 gnd.n6931 240.244
R5955 gnd.n6928 gnd.n6927 240.244
R5956 gnd.n6924 gnd.n6923 240.244
R5957 gnd.n6920 gnd.n6919 240.244
R5958 gnd.n6916 gnd.n6915 240.244
R5959 gnd.n6912 gnd.n6911 240.244
R5960 gnd.n6908 gnd.n6907 240.244
R5961 gnd.n6904 gnd.n6903 240.244
R5962 gnd.n464 gnd.n463 240.244
R5963 gnd.n6974 gnd.n390 240.244
R5964 gnd.n6974 gnd.n377 240.244
R5965 gnd.n6984 gnd.n377 240.244
R5966 gnd.n6984 gnd.n373 240.244
R5967 gnd.n6990 gnd.n373 240.244
R5968 gnd.n6990 gnd.n359 240.244
R5969 gnd.n7000 gnd.n359 240.244
R5970 gnd.n7000 gnd.n355 240.244
R5971 gnd.n7006 gnd.n355 240.244
R5972 gnd.n7006 gnd.n342 240.244
R5973 gnd.n7016 gnd.n342 240.244
R5974 gnd.n7016 gnd.n338 240.244
R5975 gnd.n7022 gnd.n338 240.244
R5976 gnd.n7022 gnd.n324 240.244
R5977 gnd.n7032 gnd.n324 240.244
R5978 gnd.n7032 gnd.n320 240.244
R5979 gnd.n7038 gnd.n320 240.244
R5980 gnd.n7038 gnd.n304 240.244
R5981 gnd.n7049 gnd.n304 240.244
R5982 gnd.n7049 gnd.n305 240.244
R5983 gnd.n305 gnd.n300 240.244
R5984 gnd.n7057 gnd.n300 240.244
R5985 gnd.n7057 gnd.n287 240.244
R5986 gnd.n7067 gnd.n287 240.244
R5987 gnd.n7067 gnd.n285 240.244
R5988 gnd.n7073 gnd.n285 240.244
R5989 gnd.n7073 gnd.n271 240.244
R5990 gnd.n7084 gnd.n271 240.244
R5991 gnd.n7084 gnd.n269 240.244
R5992 gnd.n7089 gnd.n269 240.244
R5993 gnd.n7089 gnd.n257 240.244
R5994 gnd.n7099 gnd.n257 240.244
R5995 gnd.n7099 gnd.n253 240.244
R5996 gnd.n7105 gnd.n253 240.244
R5997 gnd.n7105 gnd.n240 240.244
R5998 gnd.n7115 gnd.n240 240.244
R5999 gnd.n7115 gnd.n236 240.244
R6000 gnd.n7121 gnd.n236 240.244
R6001 gnd.n7121 gnd.n224 240.244
R6002 gnd.n7131 gnd.n224 240.244
R6003 gnd.n7131 gnd.n220 240.244
R6004 gnd.n7137 gnd.n220 240.244
R6005 gnd.n7137 gnd.n210 240.244
R6006 gnd.n7147 gnd.n210 240.244
R6007 gnd.n7147 gnd.n206 240.244
R6008 gnd.n7153 gnd.n206 240.244
R6009 gnd.n7153 gnd.n195 240.244
R6010 gnd.n7163 gnd.n195 240.244
R6011 gnd.n7163 gnd.n190 240.244
R6012 gnd.n7171 gnd.n190 240.244
R6013 gnd.n7171 gnd.n191 240.244
R6014 gnd.n191 gnd.n104 240.244
R6015 gnd.n7326 gnd.n104 240.244
R6016 gnd.n5926 gnd.n1272 240.244
R6017 gnd.n5924 gnd.n5923 240.244
R6018 gnd.n5921 gnd.n1278 240.244
R6019 gnd.n5917 gnd.n5916 240.244
R6020 gnd.n5914 gnd.n1286 240.244
R6021 gnd.n5910 gnd.n5909 240.244
R6022 gnd.n5907 gnd.n1293 240.244
R6023 gnd.n5903 gnd.n5902 240.244
R6024 gnd.n5898 gnd.n1303 240.244
R6025 gnd.n5894 gnd.n5893 240.244
R6026 gnd.n5891 gnd.n1311 240.244
R6027 gnd.n5887 gnd.n5886 240.244
R6028 gnd.n5884 gnd.n1318 240.244
R6029 gnd.n5880 gnd.n5879 240.244
R6030 gnd.n5877 gnd.n1325 240.244
R6031 gnd.n5873 gnd.n5872 240.244
R6032 gnd.n5870 gnd.n1332 240.244
R6033 gnd.n5866 gnd.n5865 240.244
R6034 gnd.n4095 gnd.n3921 240.244
R6035 gnd.n4095 gnd.n2451 240.244
R6036 gnd.n4089 gnd.n2451 240.244
R6037 gnd.n4089 gnd.n2444 240.244
R6038 gnd.n4086 gnd.n2444 240.244
R6039 gnd.n4086 gnd.n2436 240.244
R6040 gnd.n4083 gnd.n2436 240.244
R6041 gnd.n4083 gnd.n2427 240.244
R6042 gnd.n4080 gnd.n2427 240.244
R6043 gnd.n4080 gnd.n2418 240.244
R6044 gnd.n4077 gnd.n2418 240.244
R6045 gnd.n4077 gnd.n2410 240.244
R6046 gnd.n2410 gnd.n2401 240.244
R6047 gnd.n4282 gnd.n2401 240.244
R6048 gnd.n4283 gnd.n4282 240.244
R6049 gnd.n4283 gnd.n1110 240.244
R6050 gnd.n4288 gnd.n1110 240.244
R6051 gnd.n4288 gnd.n1123 240.244
R6052 gnd.n2390 gnd.n1123 240.244
R6053 gnd.n2390 gnd.n1134 240.244
R6054 gnd.n4323 gnd.n1134 240.244
R6055 gnd.n4323 gnd.n2379 240.244
R6056 gnd.n4319 gnd.n2379 240.244
R6057 gnd.n4319 gnd.n2371 240.244
R6058 gnd.n4299 gnd.n2371 240.244
R6059 gnd.n4299 gnd.n2359 240.244
R6060 gnd.n4375 gnd.n2359 240.244
R6061 gnd.n4375 gnd.n2348 240.244
R6062 gnd.n4393 gnd.n2348 240.244
R6063 gnd.n4393 gnd.n2334 240.244
R6064 gnd.n2334 gnd.n1153 240.244
R6065 gnd.n4400 gnd.n1153 240.244
R6066 gnd.n4400 gnd.n1165 240.244
R6067 gnd.n4405 gnd.n1165 240.244
R6068 gnd.n4405 gnd.n1174 240.244
R6069 gnd.n4415 gnd.n1174 240.244
R6070 gnd.n4415 gnd.n1185 240.244
R6071 gnd.n2321 gnd.n1185 240.244
R6072 gnd.n2321 gnd.n1195 240.244
R6073 gnd.n4479 gnd.n1195 240.244
R6074 gnd.n4479 gnd.n1206 240.244
R6075 gnd.n4485 gnd.n1206 240.244
R6076 gnd.n4485 gnd.n1216 240.244
R6077 gnd.n4495 gnd.n1216 240.244
R6078 gnd.n4495 gnd.n1227 240.244
R6079 gnd.n2300 gnd.n1227 240.244
R6080 gnd.n2300 gnd.n1237 240.244
R6081 gnd.n4503 gnd.n1237 240.244
R6082 gnd.n4503 gnd.n1248 240.244
R6083 gnd.n4510 gnd.n1248 240.244
R6084 gnd.n4510 gnd.n1259 240.244
R6085 gnd.n5857 gnd.n1259 240.244
R6086 gnd.n5857 gnd.n1269 240.244
R6087 gnd.n3969 gnd.n3965 240.244
R6088 gnd.n3975 gnd.n3965 240.244
R6089 gnd.n3979 gnd.n3977 240.244
R6090 gnd.n3985 gnd.n3961 240.244
R6091 gnd.n3989 gnd.n3987 240.244
R6092 gnd.n3995 gnd.n3957 240.244
R6093 gnd.n3999 gnd.n3997 240.244
R6094 gnd.n4005 gnd.n3953 240.244
R6095 gnd.n4009 gnd.n4007 240.244
R6096 gnd.n4015 gnd.n3946 240.244
R6097 gnd.n4019 gnd.n4017 240.244
R6098 gnd.n4025 gnd.n3942 240.244
R6099 gnd.n4029 gnd.n4027 240.244
R6100 gnd.n4035 gnd.n3938 240.244
R6101 gnd.n4039 gnd.n4037 240.244
R6102 gnd.n4045 gnd.n3934 240.244
R6103 gnd.n4049 gnd.n4047 240.244
R6104 gnd.n4056 gnd.n3930 240.244
R6105 gnd.n4059 gnd.n4058 240.244
R6106 gnd.n4215 gnd.n2453 240.244
R6107 gnd.n4221 gnd.n2453 240.244
R6108 gnd.n4221 gnd.n2442 240.244
R6109 gnd.n4231 gnd.n2442 240.244
R6110 gnd.n4231 gnd.n2438 240.244
R6111 gnd.n4237 gnd.n2438 240.244
R6112 gnd.n4237 gnd.n2425 240.244
R6113 gnd.n4247 gnd.n2425 240.244
R6114 gnd.n4247 gnd.n2421 240.244
R6115 gnd.n4253 gnd.n2421 240.244
R6116 gnd.n4253 gnd.n2409 240.244
R6117 gnd.n4273 gnd.n2409 240.244
R6118 gnd.n4273 gnd.n2405 240.244
R6119 gnd.n4280 gnd.n2405 240.244
R6120 gnd.n4280 gnd.n1114 240.244
R6121 gnd.n6019 gnd.n1114 240.244
R6122 gnd.n6019 gnd.n1115 240.244
R6123 gnd.n6015 gnd.n1115 240.244
R6124 gnd.n6015 gnd.n1121 240.244
R6125 gnd.n6007 gnd.n1121 240.244
R6126 gnd.n6007 gnd.n1137 240.244
R6127 gnd.n1141 gnd.n1137 240.244
R6128 gnd.n2369 gnd.n1141 240.244
R6129 gnd.n4356 gnd.n2369 240.244
R6130 gnd.n4358 gnd.n4356 240.244
R6131 gnd.n4361 gnd.n4358 240.244
R6132 gnd.n4361 gnd.n2351 240.244
R6133 gnd.n4388 gnd.n2351 240.244
R6134 gnd.n4391 gnd.n4388 240.244
R6135 gnd.n4391 gnd.n1151 240.244
R6136 gnd.n6000 gnd.n1151 240.244
R6137 gnd.n6000 gnd.n1152 240.244
R6138 gnd.n5992 gnd.n1152 240.244
R6139 gnd.n5992 gnd.n1167 240.244
R6140 gnd.n5988 gnd.n1167 240.244
R6141 gnd.n5988 gnd.n1172 240.244
R6142 gnd.n5980 gnd.n1172 240.244
R6143 gnd.n5980 gnd.n1188 240.244
R6144 gnd.n5976 gnd.n1188 240.244
R6145 gnd.n5976 gnd.n1194 240.244
R6146 gnd.n5968 gnd.n1194 240.244
R6147 gnd.n5968 gnd.n1208 240.244
R6148 gnd.n5964 gnd.n1208 240.244
R6149 gnd.n5964 gnd.n1214 240.244
R6150 gnd.n5956 gnd.n1214 240.244
R6151 gnd.n5956 gnd.n1230 240.244
R6152 gnd.n5952 gnd.n1230 240.244
R6153 gnd.n5952 gnd.n1236 240.244
R6154 gnd.n5944 gnd.n1236 240.244
R6155 gnd.n5944 gnd.n1251 240.244
R6156 gnd.n5940 gnd.n1251 240.244
R6157 gnd.n5940 gnd.n1257 240.244
R6158 gnd.n5932 gnd.n1257 240.244
R6159 gnd.n3918 gnd.n2481 240.244
R6160 gnd.n3911 gnd.n3910 240.244
R6161 gnd.n3908 gnd.n3907 240.244
R6162 gnd.n3904 gnd.n3903 240.244
R6163 gnd.n3900 gnd.n3899 240.244
R6164 gnd.n3896 gnd.n3895 240.244
R6165 gnd.n3892 gnd.n3891 240.244
R6166 gnd.n3888 gnd.n3887 240.244
R6167 gnd.n3162 gnd.n2874 240.244
R6168 gnd.n3172 gnd.n2874 240.244
R6169 gnd.n3172 gnd.n2865 240.244
R6170 gnd.n2865 gnd.n2854 240.244
R6171 gnd.n3193 gnd.n2854 240.244
R6172 gnd.n3193 gnd.n2848 240.244
R6173 gnd.n3203 gnd.n2848 240.244
R6174 gnd.n3203 gnd.n2837 240.244
R6175 gnd.n2837 gnd.n2829 240.244
R6176 gnd.n3221 gnd.n2829 240.244
R6177 gnd.n3222 gnd.n3221 240.244
R6178 gnd.n3222 gnd.n2814 240.244
R6179 gnd.n3224 gnd.n2814 240.244
R6180 gnd.n3224 gnd.n2800 240.244
R6181 gnd.n3266 gnd.n2800 240.244
R6182 gnd.n3267 gnd.n3266 240.244
R6183 gnd.n3270 gnd.n3267 240.244
R6184 gnd.n3270 gnd.n2755 240.244
R6185 gnd.n2795 gnd.n2755 240.244
R6186 gnd.n2795 gnd.n2765 240.244
R6187 gnd.n3280 gnd.n2765 240.244
R6188 gnd.n3280 gnd.n2786 240.244
R6189 gnd.n3290 gnd.n2786 240.244
R6190 gnd.n3290 gnd.n2684 240.244
R6191 gnd.n3335 gnd.n2684 240.244
R6192 gnd.n3335 gnd.n2670 240.244
R6193 gnd.n3357 gnd.n2670 240.244
R6194 gnd.n3358 gnd.n3357 240.244
R6195 gnd.n3358 gnd.n2657 240.244
R6196 gnd.n2657 gnd.n2646 240.244
R6197 gnd.n3389 gnd.n2646 240.244
R6198 gnd.n3390 gnd.n3389 240.244
R6199 gnd.n3391 gnd.n3390 240.244
R6200 gnd.n3391 gnd.n2631 240.244
R6201 gnd.n2631 gnd.n2630 240.244
R6202 gnd.n2630 gnd.n2615 240.244
R6203 gnd.n3442 gnd.n2615 240.244
R6204 gnd.n3443 gnd.n3442 240.244
R6205 gnd.n3443 gnd.n2602 240.244
R6206 gnd.n2602 gnd.n2591 240.244
R6207 gnd.n3474 gnd.n2591 240.244
R6208 gnd.n3475 gnd.n3474 240.244
R6209 gnd.n3476 gnd.n3475 240.244
R6210 gnd.n3476 gnd.n2575 240.244
R6211 gnd.n2575 gnd.n2574 240.244
R6212 gnd.n2574 gnd.n2560 240.244
R6213 gnd.n3531 gnd.n2560 240.244
R6214 gnd.n3532 gnd.n3531 240.244
R6215 gnd.n3532 gnd.n2547 240.244
R6216 gnd.n2547 gnd.n2537 240.244
R6217 gnd.n3819 gnd.n2537 240.244
R6218 gnd.n3822 gnd.n3819 240.244
R6219 gnd.n3822 gnd.n3821 240.244
R6220 gnd.n3152 gnd.n2887 240.244
R6221 gnd.n2908 gnd.n2887 240.244
R6222 gnd.n2911 gnd.n2910 240.244
R6223 gnd.n2918 gnd.n2917 240.244
R6224 gnd.n2921 gnd.n2920 240.244
R6225 gnd.n2928 gnd.n2927 240.244
R6226 gnd.n2931 gnd.n2930 240.244
R6227 gnd.n2938 gnd.n2937 240.244
R6228 gnd.n3160 gnd.n2884 240.244
R6229 gnd.n2884 gnd.n2863 240.244
R6230 gnd.n3183 gnd.n2863 240.244
R6231 gnd.n3183 gnd.n2857 240.244
R6232 gnd.n3191 gnd.n2857 240.244
R6233 gnd.n3191 gnd.n2859 240.244
R6234 gnd.n2859 gnd.n2835 240.244
R6235 gnd.n3213 gnd.n2835 240.244
R6236 gnd.n3213 gnd.n2831 240.244
R6237 gnd.n3219 gnd.n2831 240.244
R6238 gnd.n3219 gnd.n2813 240.244
R6239 gnd.n3244 gnd.n2813 240.244
R6240 gnd.n3244 gnd.n2808 240.244
R6241 gnd.n3256 gnd.n2808 240.244
R6242 gnd.n3256 gnd.n2809 240.244
R6243 gnd.n3252 gnd.n2809 240.244
R6244 gnd.n3252 gnd.n2757 240.244
R6245 gnd.n3304 gnd.n2757 240.244
R6246 gnd.n3304 gnd.n2758 240.244
R6247 gnd.n3300 gnd.n2758 240.244
R6248 gnd.n3300 gnd.n2764 240.244
R6249 gnd.n2784 gnd.n2764 240.244
R6250 gnd.n2784 gnd.n2682 240.244
R6251 gnd.n3339 gnd.n2682 240.244
R6252 gnd.n3339 gnd.n2677 240.244
R6253 gnd.n3347 gnd.n2677 240.244
R6254 gnd.n3347 gnd.n2678 240.244
R6255 gnd.n2678 gnd.n2655 240.244
R6256 gnd.n3379 gnd.n2655 240.244
R6257 gnd.n3379 gnd.n2650 240.244
R6258 gnd.n3387 gnd.n2650 240.244
R6259 gnd.n3387 gnd.n2651 240.244
R6260 gnd.n2651 gnd.n2628 240.244
R6261 gnd.n3424 gnd.n2628 240.244
R6262 gnd.n3424 gnd.n2623 240.244
R6263 gnd.n3432 gnd.n2623 240.244
R6264 gnd.n3432 gnd.n2624 240.244
R6265 gnd.n2624 gnd.n2600 240.244
R6266 gnd.n3464 gnd.n2600 240.244
R6267 gnd.n3464 gnd.n2595 240.244
R6268 gnd.n3472 gnd.n2595 240.244
R6269 gnd.n3472 gnd.n2596 240.244
R6270 gnd.n2596 gnd.n2572 240.244
R6271 gnd.n3513 gnd.n2572 240.244
R6272 gnd.n3513 gnd.n2567 240.244
R6273 gnd.n3521 gnd.n2567 240.244
R6274 gnd.n3521 gnd.n2568 240.244
R6275 gnd.n2568 gnd.n2545 240.244
R6276 gnd.n3807 gnd.n2545 240.244
R6277 gnd.n3807 gnd.n2540 240.244
R6278 gnd.n3817 gnd.n2540 240.244
R6279 gnd.n3817 gnd.n2541 240.244
R6280 gnd.n2541 gnd.n2480 240.244
R6281 gnd.n2500 gnd.n2458 240.244
R6282 gnd.n3878 gnd.n3877 240.244
R6283 gnd.n3874 gnd.n3873 240.244
R6284 gnd.n3870 gnd.n3869 240.244
R6285 gnd.n3866 gnd.n3865 240.244
R6286 gnd.n3862 gnd.n3861 240.244
R6287 gnd.n3858 gnd.n3857 240.244
R6288 gnd.n3854 gnd.n3853 240.244
R6289 gnd.n3850 gnd.n3849 240.244
R6290 gnd.n3846 gnd.n3845 240.244
R6291 gnd.n3842 gnd.n3841 240.244
R6292 gnd.n3838 gnd.n3837 240.244
R6293 gnd.n3834 gnd.n3833 240.244
R6294 gnd.n3075 gnd.n2972 240.244
R6295 gnd.n3075 gnd.n2965 240.244
R6296 gnd.n3086 gnd.n2965 240.244
R6297 gnd.n3086 gnd.n2961 240.244
R6298 gnd.n3092 gnd.n2961 240.244
R6299 gnd.n3092 gnd.n2953 240.244
R6300 gnd.n3102 gnd.n2953 240.244
R6301 gnd.n3102 gnd.n2948 240.244
R6302 gnd.n3138 gnd.n2948 240.244
R6303 gnd.n3138 gnd.n2949 240.244
R6304 gnd.n2949 gnd.n2896 240.244
R6305 gnd.n3133 gnd.n2896 240.244
R6306 gnd.n3133 gnd.n3132 240.244
R6307 gnd.n3132 gnd.n2875 240.244
R6308 gnd.n3128 gnd.n2875 240.244
R6309 gnd.n3128 gnd.n2866 240.244
R6310 gnd.n3125 gnd.n2866 240.244
R6311 gnd.n3125 gnd.n3124 240.244
R6312 gnd.n3124 gnd.n2849 240.244
R6313 gnd.n3120 gnd.n2849 240.244
R6314 gnd.n3120 gnd.n2838 240.244
R6315 gnd.n2838 gnd.n2819 240.244
R6316 gnd.n3233 gnd.n2819 240.244
R6317 gnd.n3233 gnd.n2815 240.244
R6318 gnd.n3241 gnd.n2815 240.244
R6319 gnd.n3241 gnd.n2806 240.244
R6320 gnd.n2806 gnd.n2742 240.244
R6321 gnd.n3313 gnd.n2742 240.244
R6322 gnd.n3313 gnd.n2743 240.244
R6323 gnd.n2754 gnd.n2743 240.244
R6324 gnd.n2789 gnd.n2754 240.244
R6325 gnd.n2792 gnd.n2789 240.244
R6326 gnd.n2792 gnd.n2766 240.244
R6327 gnd.n2779 gnd.n2766 240.244
R6328 gnd.n2779 gnd.n2776 240.244
R6329 gnd.n2776 gnd.n2685 240.244
R6330 gnd.n3334 gnd.n2685 240.244
R6331 gnd.n3334 gnd.n2675 240.244
R6332 gnd.n3330 gnd.n2675 240.244
R6333 gnd.n3330 gnd.n2669 240.244
R6334 gnd.n3327 gnd.n2669 240.244
R6335 gnd.n3327 gnd.n2658 240.244
R6336 gnd.n3324 gnd.n2658 240.244
R6337 gnd.n3324 gnd.n2636 240.244
R6338 gnd.n3400 gnd.n2636 240.244
R6339 gnd.n3400 gnd.n2632 240.244
R6340 gnd.n3421 gnd.n2632 240.244
R6341 gnd.n3421 gnd.n2621 240.244
R6342 gnd.n3417 gnd.n2621 240.244
R6343 gnd.n3417 gnd.n2614 240.244
R6344 gnd.n3414 gnd.n2614 240.244
R6345 gnd.n3414 gnd.n2603 240.244
R6346 gnd.n3411 gnd.n2603 240.244
R6347 gnd.n3411 gnd.n2580 240.244
R6348 gnd.n3485 gnd.n2580 240.244
R6349 gnd.n3485 gnd.n2576 240.244
R6350 gnd.n3510 gnd.n2576 240.244
R6351 gnd.n3510 gnd.n2566 240.244
R6352 gnd.n3506 gnd.n2566 240.244
R6353 gnd.n3506 gnd.n2559 240.244
R6354 gnd.n3502 gnd.n2559 240.244
R6355 gnd.n3502 gnd.n2548 240.244
R6356 gnd.n3499 gnd.n2548 240.244
R6357 gnd.n3499 gnd.n2529 240.244
R6358 gnd.n3829 gnd.n2529 240.244
R6359 gnd.n2989 gnd.n2988 240.244
R6360 gnd.n3060 gnd.n2988 240.244
R6361 gnd.n3058 gnd.n3057 240.244
R6362 gnd.n3054 gnd.n3053 240.244
R6363 gnd.n3050 gnd.n3049 240.244
R6364 gnd.n3046 gnd.n3045 240.244
R6365 gnd.n3042 gnd.n3041 240.244
R6366 gnd.n3038 gnd.n3037 240.244
R6367 gnd.n3034 gnd.n3033 240.244
R6368 gnd.n3030 gnd.n3029 240.244
R6369 gnd.n3026 gnd.n3025 240.244
R6370 gnd.n3022 gnd.n3021 240.244
R6371 gnd.n3018 gnd.n2976 240.244
R6372 gnd.n3078 gnd.n2970 240.244
R6373 gnd.n3078 gnd.n2966 240.244
R6374 gnd.n3084 gnd.n2966 240.244
R6375 gnd.n3084 gnd.n2959 240.244
R6376 gnd.n3094 gnd.n2959 240.244
R6377 gnd.n3094 gnd.n2955 240.244
R6378 gnd.n3100 gnd.n2955 240.244
R6379 gnd.n3100 gnd.n2946 240.244
R6380 gnd.n3140 gnd.n2946 240.244
R6381 gnd.n3140 gnd.n2897 240.244
R6382 gnd.n3148 gnd.n2897 240.244
R6383 gnd.n3148 gnd.n2898 240.244
R6384 gnd.n2898 gnd.n2876 240.244
R6385 gnd.n3169 gnd.n2876 240.244
R6386 gnd.n3169 gnd.n2868 240.244
R6387 gnd.n3180 gnd.n2868 240.244
R6388 gnd.n3180 gnd.n2869 240.244
R6389 gnd.n2869 gnd.n2850 240.244
R6390 gnd.n3200 gnd.n2850 240.244
R6391 gnd.n3200 gnd.n2840 240.244
R6392 gnd.n3210 gnd.n2840 240.244
R6393 gnd.n3210 gnd.n2821 240.244
R6394 gnd.n3231 gnd.n2821 240.244
R6395 gnd.n3231 gnd.n2823 240.244
R6396 gnd.n2823 gnd.n2804 240.244
R6397 gnd.n3259 gnd.n2804 240.244
R6398 gnd.n3259 gnd.n2746 240.244
R6399 gnd.n3311 gnd.n2746 240.244
R6400 gnd.n3311 gnd.n2747 240.244
R6401 gnd.n3307 gnd.n2747 240.244
R6402 gnd.n3307 gnd.n2753 240.244
R6403 gnd.n2768 gnd.n2753 240.244
R6404 gnd.n3297 gnd.n2768 240.244
R6405 gnd.n3297 gnd.n2769 240.244
R6406 gnd.n3293 gnd.n2769 240.244
R6407 gnd.n3293 gnd.n2775 240.244
R6408 gnd.n2775 gnd.n2674 240.244
R6409 gnd.n3350 gnd.n2674 240.244
R6410 gnd.n3350 gnd.n2667 240.244
R6411 gnd.n3361 gnd.n2667 240.244
R6412 gnd.n3361 gnd.n2660 240.244
R6413 gnd.n3376 gnd.n2660 240.244
R6414 gnd.n3376 gnd.n2661 240.244
R6415 gnd.n2661 gnd.n2639 240.244
R6416 gnd.n3398 gnd.n2639 240.244
R6417 gnd.n3398 gnd.n2640 240.244
R6418 gnd.n2640 gnd.n2619 240.244
R6419 gnd.n3435 gnd.n2619 240.244
R6420 gnd.n3435 gnd.n2612 240.244
R6421 gnd.n3446 gnd.n2612 240.244
R6422 gnd.n3446 gnd.n2605 240.244
R6423 gnd.n3461 gnd.n2605 240.244
R6424 gnd.n3461 gnd.n2606 240.244
R6425 gnd.n2606 gnd.n2583 240.244
R6426 gnd.n3483 gnd.n2583 240.244
R6427 gnd.n3483 gnd.n2585 240.244
R6428 gnd.n2585 gnd.n2564 240.244
R6429 gnd.n3524 gnd.n2564 240.244
R6430 gnd.n3524 gnd.n2557 240.244
R6431 gnd.n3535 gnd.n2557 240.244
R6432 gnd.n3535 gnd.n2550 240.244
R6433 gnd.n3804 gnd.n2550 240.244
R6434 gnd.n3804 gnd.n2551 240.244
R6435 gnd.n2551 gnd.n2532 240.244
R6436 gnd.n3827 gnd.n2532 240.244
R6437 gnd.n7179 gnd.n7178 240.244
R6438 gnd.n7184 gnd.n7181 240.244
R6439 gnd.n7187 gnd.n7186 240.244
R6440 gnd.n7192 gnd.n7189 240.244
R6441 gnd.n7195 gnd.n7194 240.244
R6442 gnd.n7200 gnd.n7197 240.244
R6443 gnd.n7203 gnd.n7202 240.244
R6444 gnd.n7208 gnd.n7205 240.244
R6445 gnd.n7214 gnd.n7210 240.244
R6446 gnd.n6893 gnd.n389 240.244
R6447 gnd.n474 gnd.n389 240.244
R6448 gnd.n474 gnd.n380 240.244
R6449 gnd.n475 gnd.n380 240.244
R6450 gnd.n475 gnd.n371 240.244
R6451 gnd.n478 gnd.n371 240.244
R6452 gnd.n478 gnd.n362 240.244
R6453 gnd.n479 gnd.n362 240.244
R6454 gnd.n479 gnd.n354 240.244
R6455 gnd.n482 gnd.n354 240.244
R6456 gnd.n482 gnd.n345 240.244
R6457 gnd.n483 gnd.n345 240.244
R6458 gnd.n483 gnd.n336 240.244
R6459 gnd.n486 gnd.n336 240.244
R6460 gnd.n486 gnd.n327 240.244
R6461 gnd.n487 gnd.n327 240.244
R6462 gnd.n487 gnd.n319 240.244
R6463 gnd.n490 gnd.n319 240.244
R6464 gnd.n490 gnd.n308 240.244
R6465 gnd.n491 gnd.n308 240.244
R6466 gnd.n5532 gnd.n491 240.244
R6467 gnd.n5532 gnd.n299 240.244
R6468 gnd.n494 gnd.n299 240.244
R6469 gnd.n494 gnd.n290 240.244
R6470 gnd.n6852 gnd.n290 240.244
R6471 gnd.n6852 gnd.n283 240.244
R6472 gnd.n283 gnd.n66 240.244
R6473 gnd.n67 gnd.n66 240.244
R6474 gnd.n68 gnd.n67 240.244
R6475 gnd.n268 gnd.n68 240.244
R6476 gnd.n268 gnd.n71 240.244
R6477 gnd.n72 gnd.n71 240.244
R6478 gnd.n73 gnd.n72 240.244
R6479 gnd.n251 gnd.n73 240.244
R6480 gnd.n251 gnd.n76 240.244
R6481 gnd.n77 gnd.n76 240.244
R6482 gnd.n78 gnd.n77 240.244
R6483 gnd.n235 gnd.n78 240.244
R6484 gnd.n235 gnd.n81 240.244
R6485 gnd.n82 gnd.n81 240.244
R6486 gnd.n83 gnd.n82 240.244
R6487 gnd.n218 gnd.n83 240.244
R6488 gnd.n218 gnd.n86 240.244
R6489 gnd.n87 gnd.n86 240.244
R6490 gnd.n88 gnd.n87 240.244
R6491 gnd.n205 gnd.n88 240.244
R6492 gnd.n205 gnd.n91 240.244
R6493 gnd.n92 gnd.n91 240.244
R6494 gnd.n93 gnd.n92 240.244
R6495 gnd.n188 gnd.n93 240.244
R6496 gnd.n188 gnd.n96 240.244
R6497 gnd.n97 gnd.n96 240.244
R6498 gnd.n7328 gnd.n97 240.244
R6499 gnd.n1479 gnd.n1478 240.244
R6500 gnd.n1489 gnd.n1488 240.244
R6501 gnd.n1491 gnd.n1490 240.244
R6502 gnd.n1499 gnd.n1498 240.244
R6503 gnd.n1507 gnd.n1506 240.244
R6504 gnd.n1509 gnd.n1508 240.244
R6505 gnd.n1517 gnd.n1516 240.244
R6506 gnd.n1525 gnd.n1524 240.244
R6507 gnd.n5656 gnd.n423 240.244
R6508 gnd.n6976 gnd.n386 240.244
R6509 gnd.n6976 gnd.n382 240.244
R6510 gnd.n6982 gnd.n382 240.244
R6511 gnd.n6982 gnd.n368 240.244
R6512 gnd.n6992 gnd.n368 240.244
R6513 gnd.n6992 gnd.n364 240.244
R6514 gnd.n6998 gnd.n364 240.244
R6515 gnd.n6998 gnd.n351 240.244
R6516 gnd.n7008 gnd.n351 240.244
R6517 gnd.n7008 gnd.n347 240.244
R6518 gnd.n7014 gnd.n347 240.244
R6519 gnd.n7014 gnd.n333 240.244
R6520 gnd.n7024 gnd.n333 240.244
R6521 gnd.n7024 gnd.n329 240.244
R6522 gnd.n7030 gnd.n329 240.244
R6523 gnd.n7030 gnd.n316 240.244
R6524 gnd.n7040 gnd.n316 240.244
R6525 gnd.n7040 gnd.n310 240.244
R6526 gnd.n7047 gnd.n310 240.244
R6527 gnd.n7047 gnd.n311 240.244
R6528 gnd.n311 gnd.n296 240.244
R6529 gnd.n7059 gnd.n296 240.244
R6530 gnd.n7059 gnd.n292 240.244
R6531 gnd.n7065 gnd.n292 240.244
R6532 gnd.n7065 gnd.n280 240.244
R6533 gnd.n7075 gnd.n280 240.244
R6534 gnd.n7075 gnd.n275 240.244
R6535 gnd.n7082 gnd.n275 240.244
R6536 gnd.n7082 gnd.n265 240.244
R6537 gnd.n7091 gnd.n265 240.244
R6538 gnd.n7091 gnd.n261 240.244
R6539 gnd.n7097 gnd.n261 240.244
R6540 gnd.n7097 gnd.n248 240.244
R6541 gnd.n7107 gnd.n248 240.244
R6542 gnd.n7107 gnd.n244 240.244
R6543 gnd.n7113 gnd.n244 240.244
R6544 gnd.n7113 gnd.n232 240.244
R6545 gnd.n7123 gnd.n232 240.244
R6546 gnd.n7123 gnd.n228 240.244
R6547 gnd.n7129 gnd.n228 240.244
R6548 gnd.n7129 gnd.n216 240.244
R6549 gnd.n7139 gnd.n216 240.244
R6550 gnd.n7139 gnd.n212 240.244
R6551 gnd.n7145 gnd.n212 240.244
R6552 gnd.n7145 gnd.n202 240.244
R6553 gnd.n7155 gnd.n202 240.244
R6554 gnd.n7155 gnd.n198 240.244
R6555 gnd.n7161 gnd.n198 240.244
R6556 gnd.n7161 gnd.n185 240.244
R6557 gnd.n7173 gnd.n185 240.244
R6558 gnd.n7173 gnd.n180 240.244
R6559 gnd.n7247 gnd.n180 240.244
R6560 gnd.n7247 gnd.n103 240.244
R6561 gnd.n2202 gnd.n1267 240.244
R6562 gnd.n2213 gnd.n2204 240.244
R6563 gnd.n2216 gnd.n2215 240.244
R6564 gnd.n2225 gnd.n2224 240.244
R6565 gnd.n2234 gnd.n2227 240.244
R6566 gnd.n2237 gnd.n2236 240.244
R6567 gnd.n2246 gnd.n2245 240.244
R6568 gnd.n2255 gnd.n2248 240.244
R6569 gnd.n2261 gnd.n2257 240.244
R6570 gnd.n4125 gnd.n3922 240.244
R6571 gnd.n4125 gnd.n2452 240.244
R6572 gnd.n4164 gnd.n2452 240.244
R6573 gnd.n4164 gnd.n2445 240.244
R6574 gnd.n4161 gnd.n2445 240.244
R6575 gnd.n4161 gnd.n2437 240.244
R6576 gnd.n4158 gnd.n2437 240.244
R6577 gnd.n4158 gnd.n2428 240.244
R6578 gnd.n4155 gnd.n2428 240.244
R6579 gnd.n4155 gnd.n2419 240.244
R6580 gnd.n4152 gnd.n2419 240.244
R6581 gnd.n4152 gnd.n2411 240.244
R6582 gnd.n4149 gnd.n2411 240.244
R6583 gnd.n4149 gnd.n2403 240.244
R6584 gnd.n4146 gnd.n2403 240.244
R6585 gnd.n4146 gnd.n1111 240.244
R6586 gnd.n4143 gnd.n1111 240.244
R6587 gnd.n4143 gnd.n1124 240.244
R6588 gnd.n4329 gnd.n1124 240.244
R6589 gnd.n4329 gnd.n1135 240.244
R6590 gnd.n4325 gnd.n1135 240.244
R6591 gnd.n4325 gnd.n2380 240.244
R6592 gnd.n4317 gnd.n2380 240.244
R6593 gnd.n4317 gnd.n2372 240.244
R6594 gnd.n4313 gnd.n2372 240.244
R6595 gnd.n4313 gnd.n2367 240.244
R6596 gnd.n2367 gnd.n2361 240.244
R6597 gnd.n2361 gnd.n2352 240.244
R6598 gnd.n2352 gnd.n2335 240.244
R6599 gnd.n4429 gnd.n2335 240.244
R6600 gnd.n4429 gnd.n1154 240.244
R6601 gnd.n2340 gnd.n1154 240.244
R6602 gnd.n2340 gnd.n1166 240.244
R6603 gnd.n2341 gnd.n1166 240.244
R6604 gnd.n2341 gnd.n1175 240.244
R6605 gnd.n4417 gnd.n1175 240.244
R6606 gnd.n4417 gnd.n1186 240.244
R6607 gnd.n4471 gnd.n1186 240.244
R6608 gnd.n4471 gnd.n1196 240.244
R6609 gnd.n4477 gnd.n1196 240.244
R6610 gnd.n4477 gnd.n1207 240.244
R6611 gnd.n4487 gnd.n1207 240.244
R6612 gnd.n4487 gnd.n1217 240.244
R6613 gnd.n4493 gnd.n1217 240.244
R6614 gnd.n4493 gnd.n1228 240.244
R6615 gnd.n4521 gnd.n1228 240.244
R6616 gnd.n4521 gnd.n1238 240.244
R6617 gnd.n2305 gnd.n1238 240.244
R6618 gnd.n2305 gnd.n1249 240.244
R6619 gnd.n4512 gnd.n1249 240.244
R6620 gnd.n4512 gnd.n1260 240.244
R6621 gnd.n5855 gnd.n1260 240.244
R6622 gnd.n5855 gnd.n1270 240.244
R6623 gnd.n4207 gnd.n4205 240.244
R6624 gnd.n4203 gnd.n4100 240.244
R6625 gnd.n4199 gnd.n4197 240.244
R6626 gnd.n4195 gnd.n4106 240.244
R6627 gnd.n4191 gnd.n4189 240.244
R6628 gnd.n4187 gnd.n4112 240.244
R6629 gnd.n4183 gnd.n4181 240.244
R6630 gnd.n4179 gnd.n4118 240.244
R6631 gnd.n4172 gnd.n4171 240.244
R6632 gnd.n4213 gnd.n2450 240.244
R6633 gnd.n4223 gnd.n2450 240.244
R6634 gnd.n4223 gnd.n2446 240.244
R6635 gnd.n4229 gnd.n2446 240.244
R6636 gnd.n4229 gnd.n2434 240.244
R6637 gnd.n4239 gnd.n2434 240.244
R6638 gnd.n4239 gnd.n2430 240.244
R6639 gnd.n4245 gnd.n2430 240.244
R6640 gnd.n4245 gnd.n2417 240.244
R6641 gnd.n4255 gnd.n2417 240.244
R6642 gnd.n4255 gnd.n2412 240.244
R6643 gnd.n4271 gnd.n2412 240.244
R6644 gnd.n4271 gnd.n2413 240.244
R6645 gnd.n2413 gnd.n2404 240.244
R6646 gnd.n4266 gnd.n2404 240.244
R6647 gnd.n4266 gnd.n1113 240.244
R6648 gnd.n1126 gnd.n1113 240.244
R6649 gnd.n6013 gnd.n1126 240.244
R6650 gnd.n6013 gnd.n1127 240.244
R6651 gnd.n6009 gnd.n1127 240.244
R6652 gnd.n6009 gnd.n1133 240.244
R6653 gnd.n4345 gnd.n1133 240.244
R6654 gnd.n4345 gnd.n2374 240.244
R6655 gnd.n4354 gnd.n2374 240.244
R6656 gnd.n4354 gnd.n2375 240.244
R6657 gnd.n2375 gnd.n2368 240.244
R6658 gnd.n2368 gnd.n2353 240.244
R6659 gnd.n4386 gnd.n2353 240.244
R6660 gnd.n4386 gnd.n2350 240.244
R6661 gnd.n2350 gnd.n1156 240.244
R6662 gnd.n5998 gnd.n1156 240.244
R6663 gnd.n5998 gnd.n1157 240.244
R6664 gnd.n5994 gnd.n1157 240.244
R6665 gnd.n5994 gnd.n1163 240.244
R6666 gnd.n5986 gnd.n1163 240.244
R6667 gnd.n5986 gnd.n1177 240.244
R6668 gnd.n5982 gnd.n1177 240.244
R6669 gnd.n5982 gnd.n1183 240.244
R6670 gnd.n5974 gnd.n1183 240.244
R6671 gnd.n5974 gnd.n1198 240.244
R6672 gnd.n5970 gnd.n1198 240.244
R6673 gnd.n5970 gnd.n1204 240.244
R6674 gnd.n5962 gnd.n1204 240.244
R6675 gnd.n5962 gnd.n1219 240.244
R6676 gnd.n5958 gnd.n1219 240.244
R6677 gnd.n5958 gnd.n1225 240.244
R6678 gnd.n5950 gnd.n1225 240.244
R6679 gnd.n5950 gnd.n1240 240.244
R6680 gnd.n5946 gnd.n1240 240.244
R6681 gnd.n5946 gnd.n1246 240.244
R6682 gnd.n5938 gnd.n1246 240.244
R6683 gnd.n5938 gnd.n1262 240.244
R6684 gnd.n5934 gnd.n1262 240.244
R6685 gnd.n6196 gnd.n938 240.244
R6686 gnd.n6196 gnd.n936 240.244
R6687 gnd.n6200 gnd.n936 240.244
R6688 gnd.n6200 gnd.n932 240.244
R6689 gnd.n6206 gnd.n932 240.244
R6690 gnd.n6206 gnd.n930 240.244
R6691 gnd.n6210 gnd.n930 240.244
R6692 gnd.n6210 gnd.n926 240.244
R6693 gnd.n6216 gnd.n926 240.244
R6694 gnd.n6216 gnd.n924 240.244
R6695 gnd.n6220 gnd.n924 240.244
R6696 gnd.n6220 gnd.n920 240.244
R6697 gnd.n6226 gnd.n920 240.244
R6698 gnd.n6226 gnd.n918 240.244
R6699 gnd.n6230 gnd.n918 240.244
R6700 gnd.n6230 gnd.n914 240.244
R6701 gnd.n6236 gnd.n914 240.244
R6702 gnd.n6236 gnd.n912 240.244
R6703 gnd.n6240 gnd.n912 240.244
R6704 gnd.n6240 gnd.n908 240.244
R6705 gnd.n6246 gnd.n908 240.244
R6706 gnd.n6246 gnd.n906 240.244
R6707 gnd.n6250 gnd.n906 240.244
R6708 gnd.n6250 gnd.n902 240.244
R6709 gnd.n6256 gnd.n902 240.244
R6710 gnd.n6256 gnd.n900 240.244
R6711 gnd.n6260 gnd.n900 240.244
R6712 gnd.n6260 gnd.n896 240.244
R6713 gnd.n6266 gnd.n896 240.244
R6714 gnd.n6266 gnd.n894 240.244
R6715 gnd.n6270 gnd.n894 240.244
R6716 gnd.n6270 gnd.n890 240.244
R6717 gnd.n6276 gnd.n890 240.244
R6718 gnd.n6276 gnd.n888 240.244
R6719 gnd.n6280 gnd.n888 240.244
R6720 gnd.n6280 gnd.n884 240.244
R6721 gnd.n6286 gnd.n884 240.244
R6722 gnd.n6286 gnd.n882 240.244
R6723 gnd.n6290 gnd.n882 240.244
R6724 gnd.n6290 gnd.n878 240.244
R6725 gnd.n6296 gnd.n878 240.244
R6726 gnd.n6296 gnd.n876 240.244
R6727 gnd.n6300 gnd.n876 240.244
R6728 gnd.n6300 gnd.n872 240.244
R6729 gnd.n6306 gnd.n872 240.244
R6730 gnd.n6306 gnd.n870 240.244
R6731 gnd.n6310 gnd.n870 240.244
R6732 gnd.n6310 gnd.n866 240.244
R6733 gnd.n6316 gnd.n866 240.244
R6734 gnd.n6316 gnd.n864 240.244
R6735 gnd.n6320 gnd.n864 240.244
R6736 gnd.n6320 gnd.n860 240.244
R6737 gnd.n6326 gnd.n860 240.244
R6738 gnd.n6326 gnd.n858 240.244
R6739 gnd.n6330 gnd.n858 240.244
R6740 gnd.n6330 gnd.n854 240.244
R6741 gnd.n6336 gnd.n854 240.244
R6742 gnd.n6336 gnd.n852 240.244
R6743 gnd.n6340 gnd.n852 240.244
R6744 gnd.n6340 gnd.n848 240.244
R6745 gnd.n6346 gnd.n848 240.244
R6746 gnd.n6346 gnd.n846 240.244
R6747 gnd.n6350 gnd.n846 240.244
R6748 gnd.n6350 gnd.n842 240.244
R6749 gnd.n6356 gnd.n842 240.244
R6750 gnd.n6356 gnd.n840 240.244
R6751 gnd.n6360 gnd.n840 240.244
R6752 gnd.n6360 gnd.n836 240.244
R6753 gnd.n6366 gnd.n836 240.244
R6754 gnd.n6366 gnd.n834 240.244
R6755 gnd.n6370 gnd.n834 240.244
R6756 gnd.n6370 gnd.n830 240.244
R6757 gnd.n6376 gnd.n830 240.244
R6758 gnd.n6376 gnd.n828 240.244
R6759 gnd.n6380 gnd.n828 240.244
R6760 gnd.n6380 gnd.n824 240.244
R6761 gnd.n6386 gnd.n824 240.244
R6762 gnd.n6386 gnd.n822 240.244
R6763 gnd.n6390 gnd.n822 240.244
R6764 gnd.n6390 gnd.n818 240.244
R6765 gnd.n6396 gnd.n818 240.244
R6766 gnd.n6396 gnd.n816 240.244
R6767 gnd.n6400 gnd.n816 240.244
R6768 gnd.n6400 gnd.n812 240.244
R6769 gnd.n6406 gnd.n812 240.244
R6770 gnd.n6406 gnd.n810 240.244
R6771 gnd.n6410 gnd.n810 240.244
R6772 gnd.n6410 gnd.n806 240.244
R6773 gnd.n6416 gnd.n806 240.244
R6774 gnd.n6416 gnd.n804 240.244
R6775 gnd.n6420 gnd.n804 240.244
R6776 gnd.n6420 gnd.n800 240.244
R6777 gnd.n6426 gnd.n800 240.244
R6778 gnd.n6426 gnd.n798 240.244
R6779 gnd.n6430 gnd.n798 240.244
R6780 gnd.n6430 gnd.n794 240.244
R6781 gnd.n6436 gnd.n794 240.244
R6782 gnd.n6436 gnd.n792 240.244
R6783 gnd.n6440 gnd.n792 240.244
R6784 gnd.n6440 gnd.n788 240.244
R6785 gnd.n6446 gnd.n788 240.244
R6786 gnd.n6446 gnd.n786 240.244
R6787 gnd.n6450 gnd.n786 240.244
R6788 gnd.n6450 gnd.n782 240.244
R6789 gnd.n6456 gnd.n782 240.244
R6790 gnd.n6456 gnd.n780 240.244
R6791 gnd.n6460 gnd.n780 240.244
R6792 gnd.n6460 gnd.n776 240.244
R6793 gnd.n6466 gnd.n776 240.244
R6794 gnd.n6466 gnd.n774 240.244
R6795 gnd.n6470 gnd.n774 240.244
R6796 gnd.n6470 gnd.n770 240.244
R6797 gnd.n6476 gnd.n770 240.244
R6798 gnd.n6476 gnd.n768 240.244
R6799 gnd.n6480 gnd.n768 240.244
R6800 gnd.n6480 gnd.n764 240.244
R6801 gnd.n6486 gnd.n764 240.244
R6802 gnd.n6486 gnd.n762 240.244
R6803 gnd.n6490 gnd.n762 240.244
R6804 gnd.n6490 gnd.n758 240.244
R6805 gnd.n6496 gnd.n758 240.244
R6806 gnd.n6496 gnd.n756 240.244
R6807 gnd.n6500 gnd.n756 240.244
R6808 gnd.n6500 gnd.n752 240.244
R6809 gnd.n6506 gnd.n752 240.244
R6810 gnd.n6506 gnd.n750 240.244
R6811 gnd.n6510 gnd.n750 240.244
R6812 gnd.n6510 gnd.n746 240.244
R6813 gnd.n6516 gnd.n746 240.244
R6814 gnd.n6516 gnd.n744 240.244
R6815 gnd.n6520 gnd.n744 240.244
R6816 gnd.n6520 gnd.n740 240.244
R6817 gnd.n6526 gnd.n740 240.244
R6818 gnd.n6526 gnd.n738 240.244
R6819 gnd.n6530 gnd.n738 240.244
R6820 gnd.n6530 gnd.n734 240.244
R6821 gnd.n6536 gnd.n734 240.244
R6822 gnd.n6536 gnd.n732 240.244
R6823 gnd.n6540 gnd.n732 240.244
R6824 gnd.n6540 gnd.n728 240.244
R6825 gnd.n6546 gnd.n728 240.244
R6826 gnd.n6546 gnd.n726 240.244
R6827 gnd.n6550 gnd.n726 240.244
R6828 gnd.n6550 gnd.n722 240.244
R6829 gnd.n6556 gnd.n722 240.244
R6830 gnd.n6556 gnd.n720 240.244
R6831 gnd.n6560 gnd.n720 240.244
R6832 gnd.n6560 gnd.n716 240.244
R6833 gnd.n6566 gnd.n716 240.244
R6834 gnd.n6566 gnd.n714 240.244
R6835 gnd.n6570 gnd.n714 240.244
R6836 gnd.n6570 gnd.n710 240.244
R6837 gnd.n6576 gnd.n710 240.244
R6838 gnd.n6576 gnd.n708 240.244
R6839 gnd.n6580 gnd.n708 240.244
R6840 gnd.n6580 gnd.n704 240.244
R6841 gnd.n6586 gnd.n704 240.244
R6842 gnd.n6586 gnd.n702 240.244
R6843 gnd.n6590 gnd.n702 240.244
R6844 gnd.n6590 gnd.n698 240.244
R6845 gnd.n6596 gnd.n698 240.244
R6846 gnd.n6596 gnd.n696 240.244
R6847 gnd.n6600 gnd.n696 240.244
R6848 gnd.n6600 gnd.n692 240.244
R6849 gnd.n6606 gnd.n692 240.244
R6850 gnd.n6606 gnd.n690 240.244
R6851 gnd.n6610 gnd.n690 240.244
R6852 gnd.n6616 gnd.n686 240.244
R6853 gnd.n6616 gnd.n684 240.244
R6854 gnd.n6620 gnd.n684 240.244
R6855 gnd.n6620 gnd.n680 240.244
R6856 gnd.n6626 gnd.n680 240.244
R6857 gnd.n6626 gnd.n678 240.244
R6858 gnd.n6630 gnd.n678 240.244
R6859 gnd.n6630 gnd.n674 240.244
R6860 gnd.n6636 gnd.n674 240.244
R6861 gnd.n6636 gnd.n672 240.244
R6862 gnd.n6640 gnd.n672 240.244
R6863 gnd.n6640 gnd.n668 240.244
R6864 gnd.n6646 gnd.n668 240.244
R6865 gnd.n6646 gnd.n666 240.244
R6866 gnd.n6650 gnd.n666 240.244
R6867 gnd.n6650 gnd.n662 240.244
R6868 gnd.n6656 gnd.n662 240.244
R6869 gnd.n6656 gnd.n660 240.244
R6870 gnd.n6660 gnd.n660 240.244
R6871 gnd.n6660 gnd.n656 240.244
R6872 gnd.n6666 gnd.n656 240.244
R6873 gnd.n6666 gnd.n654 240.244
R6874 gnd.n6670 gnd.n654 240.244
R6875 gnd.n6670 gnd.n650 240.244
R6876 gnd.n6676 gnd.n650 240.244
R6877 gnd.n6676 gnd.n648 240.244
R6878 gnd.n6680 gnd.n648 240.244
R6879 gnd.n6680 gnd.n644 240.244
R6880 gnd.n6686 gnd.n644 240.244
R6881 gnd.n6686 gnd.n642 240.244
R6882 gnd.n6690 gnd.n642 240.244
R6883 gnd.n6690 gnd.n638 240.244
R6884 gnd.n6696 gnd.n638 240.244
R6885 gnd.n6696 gnd.n636 240.244
R6886 gnd.n6700 gnd.n636 240.244
R6887 gnd.n6700 gnd.n632 240.244
R6888 gnd.n6706 gnd.n632 240.244
R6889 gnd.n6706 gnd.n630 240.244
R6890 gnd.n6710 gnd.n630 240.244
R6891 gnd.n6710 gnd.n626 240.244
R6892 gnd.n6716 gnd.n626 240.244
R6893 gnd.n6716 gnd.n624 240.244
R6894 gnd.n6720 gnd.n624 240.244
R6895 gnd.n6720 gnd.n620 240.244
R6896 gnd.n6726 gnd.n620 240.244
R6897 gnd.n6726 gnd.n618 240.244
R6898 gnd.n6730 gnd.n618 240.244
R6899 gnd.n6730 gnd.n614 240.244
R6900 gnd.n6736 gnd.n614 240.244
R6901 gnd.n6736 gnd.n612 240.244
R6902 gnd.n6740 gnd.n612 240.244
R6903 gnd.n6740 gnd.n608 240.244
R6904 gnd.n6746 gnd.n608 240.244
R6905 gnd.n6746 gnd.n606 240.244
R6906 gnd.n6750 gnd.n606 240.244
R6907 gnd.n6750 gnd.n602 240.244
R6908 gnd.n6756 gnd.n602 240.244
R6909 gnd.n6756 gnd.n600 240.244
R6910 gnd.n6760 gnd.n600 240.244
R6911 gnd.n6760 gnd.n596 240.244
R6912 gnd.n6766 gnd.n596 240.244
R6913 gnd.n6766 gnd.n594 240.244
R6914 gnd.n6770 gnd.n594 240.244
R6915 gnd.n6770 gnd.n590 240.244
R6916 gnd.n6776 gnd.n590 240.244
R6917 gnd.n6776 gnd.n588 240.244
R6918 gnd.n6780 gnd.n588 240.244
R6919 gnd.n6780 gnd.n584 240.244
R6920 gnd.n6786 gnd.n584 240.244
R6921 gnd.n6786 gnd.n582 240.244
R6922 gnd.n6790 gnd.n582 240.244
R6923 gnd.n6790 gnd.n578 240.244
R6924 gnd.n6796 gnd.n578 240.244
R6925 gnd.n6796 gnd.n576 240.244
R6926 gnd.n6800 gnd.n576 240.244
R6927 gnd.n6800 gnd.n572 240.244
R6928 gnd.n6806 gnd.n572 240.244
R6929 gnd.n6806 gnd.n570 240.244
R6930 gnd.n6810 gnd.n570 240.244
R6931 gnd.n6810 gnd.n566 240.244
R6932 gnd.n6818 gnd.n566 240.244
R6933 gnd.n6818 gnd.n564 240.244
R6934 gnd.n6822 gnd.n564 240.244
R6935 gnd.n6823 gnd.n6822 240.244
R6936 gnd.n2388 gnd.n1108 240.244
R6937 gnd.n4332 gnd.n2388 240.244
R6938 gnd.n4332 gnd.n2389 240.244
R6939 gnd.n2389 gnd.n2381 240.244
R6940 gnd.n4342 gnd.n2381 240.244
R6941 gnd.n4342 gnd.n2382 240.244
R6942 gnd.n2382 gnd.n2365 240.244
R6943 gnd.n4364 gnd.n2365 240.244
R6944 gnd.n4364 gnd.n2362 240.244
R6945 gnd.n4372 gnd.n2362 240.244
R6946 gnd.n4372 gnd.n2363 240.244
R6947 gnd.n2363 gnd.n2330 240.244
R6948 gnd.n4432 gnd.n2330 240.244
R6949 gnd.n4433 gnd.n4432 240.244
R6950 gnd.n4434 gnd.n4433 240.244
R6951 gnd.n4434 gnd.n2327 240.244
R6952 gnd.n4440 gnd.n2327 240.244
R6953 gnd.n4441 gnd.n4440 240.244
R6954 gnd.n4442 gnd.n4441 240.244
R6955 gnd.n4442 gnd.n2322 240.244
R6956 gnd.n4468 gnd.n2322 240.244
R6957 gnd.n4468 gnd.n2323 240.244
R6958 gnd.n4464 gnd.n2323 240.244
R6959 gnd.n4464 gnd.n4463 240.244
R6960 gnd.n4463 gnd.n4462 240.244
R6961 gnd.n4462 gnd.n4450 240.244
R6962 gnd.n4458 gnd.n4450 240.244
R6963 gnd.n4458 gnd.n2298 240.244
R6964 gnd.n4524 gnd.n2298 240.244
R6965 gnd.n4525 gnd.n4524 240.244
R6966 gnd.n4526 gnd.n4525 240.244
R6967 gnd.n4526 gnd.n2294 240.244
R6968 gnd.n4532 gnd.n2294 240.244
R6969 gnd.n4533 gnd.n4532 240.244
R6970 gnd.n4534 gnd.n4533 240.244
R6971 gnd.n4534 gnd.n2290 240.244
R6972 gnd.n4541 gnd.n2290 240.244
R6973 gnd.n4542 gnd.n4541 240.244
R6974 gnd.n4545 gnd.n4542 240.244
R6975 gnd.n4545 gnd.n2285 240.244
R6976 gnd.n4553 gnd.n2285 240.244
R6977 gnd.n4553 gnd.n2286 240.244
R6978 gnd.n2286 gnd.n2197 240.244
R6979 gnd.n4618 gnd.n2197 240.244
R6980 gnd.n4618 gnd.n2193 240.244
R6981 gnd.n4624 gnd.n2193 240.244
R6982 gnd.n4624 gnd.n2183 240.244
R6983 gnd.n4637 gnd.n2183 240.244
R6984 gnd.n4637 gnd.n2179 240.244
R6985 gnd.n4643 gnd.n2179 240.244
R6986 gnd.n4643 gnd.n2169 240.244
R6987 gnd.n4657 gnd.n2169 240.244
R6988 gnd.n4657 gnd.n2162 240.244
R6989 gnd.n4669 gnd.n2162 240.244
R6990 gnd.n4669 gnd.n2165 240.244
R6991 gnd.n4665 gnd.n2165 240.244
R6992 gnd.n4665 gnd.n1946 240.244
R6993 gnd.n4709 gnd.n1946 240.244
R6994 gnd.n4709 gnd.n1941 240.244
R6995 gnd.n4720 gnd.n1941 240.244
R6996 gnd.n4720 gnd.n1942 240.244
R6997 gnd.n4716 gnd.n1942 240.244
R6998 gnd.n4716 gnd.n1910 240.244
R6999 gnd.n4792 gnd.n1910 240.244
R7000 gnd.n4792 gnd.n1906 240.244
R7001 gnd.n4798 gnd.n1906 240.244
R7002 gnd.n4798 gnd.n1887 240.244
R7003 gnd.n4819 gnd.n1887 240.244
R7004 gnd.n4819 gnd.n1882 240.244
R7005 gnd.n4827 gnd.n1882 240.244
R7006 gnd.n4827 gnd.n1883 240.244
R7007 gnd.n1883 gnd.n1857 240.244
R7008 gnd.n4860 gnd.n1857 240.244
R7009 gnd.n4860 gnd.n1853 240.244
R7010 gnd.n4866 gnd.n1853 240.244
R7011 gnd.n4866 gnd.n1833 240.244
R7012 gnd.n4903 gnd.n1833 240.244
R7013 gnd.n4903 gnd.n1829 240.244
R7014 gnd.n4909 gnd.n1829 240.244
R7015 gnd.n4909 gnd.n1817 240.244
R7016 gnd.n5018 gnd.n1817 240.244
R7017 gnd.n5018 gnd.n1813 240.244
R7018 gnd.n5024 gnd.n1813 240.244
R7019 gnd.n5024 gnd.n1794 240.244
R7020 gnd.n5045 gnd.n1794 240.244
R7021 gnd.n5045 gnd.n1789 240.244
R7022 gnd.n5053 gnd.n1789 240.244
R7023 gnd.n5053 gnd.n1790 240.244
R7024 gnd.n1790 gnd.n1765 240.244
R7025 gnd.n5081 gnd.n1765 240.244
R7026 gnd.n5081 gnd.n1761 240.244
R7027 gnd.n5087 gnd.n1761 240.244
R7028 gnd.n5087 gnd.n1743 240.244
R7029 gnd.n5111 gnd.n1743 240.244
R7030 gnd.n5111 gnd.n1739 240.244
R7031 gnd.n5117 gnd.n1739 240.244
R7032 gnd.n5117 gnd.n1721 240.244
R7033 gnd.n5141 gnd.n1721 240.244
R7034 gnd.n5141 gnd.n1717 240.244
R7035 gnd.n5147 gnd.n1717 240.244
R7036 gnd.n5147 gnd.n1699 240.244
R7037 gnd.n5168 gnd.n1699 240.244
R7038 gnd.n5168 gnd.n1694 240.244
R7039 gnd.n5176 gnd.n1694 240.244
R7040 gnd.n5176 gnd.n1695 240.244
R7041 gnd.n1695 gnd.n1672 240.244
R7042 gnd.n5205 gnd.n1672 240.244
R7043 gnd.n5205 gnd.n1667 240.244
R7044 gnd.n5222 gnd.n1667 240.244
R7045 gnd.n5222 gnd.n1668 240.244
R7046 gnd.n5218 gnd.n1668 240.244
R7047 gnd.n5218 gnd.n5217 240.244
R7048 gnd.n5217 gnd.n5216 240.244
R7049 gnd.n5216 gnd.n1600 240.244
R7050 gnd.n5406 gnd.n1600 240.244
R7051 gnd.n5406 gnd.n1596 240.244
R7052 gnd.n5412 gnd.n1596 240.244
R7053 gnd.n5412 gnd.n1586 240.244
R7054 gnd.n5425 gnd.n1586 240.244
R7055 gnd.n5425 gnd.n1582 240.244
R7056 gnd.n5434 gnd.n1582 240.244
R7057 gnd.n5434 gnd.n1571 240.244
R7058 gnd.n5447 gnd.n1571 240.244
R7059 gnd.n5448 gnd.n5447 240.244
R7060 gnd.n5449 gnd.n5448 240.244
R7061 gnd.n5449 gnd.n1566 240.244
R7062 gnd.n5628 gnd.n1566 240.244
R7063 gnd.n5628 gnd.n1567 240.244
R7064 gnd.n5624 gnd.n1567 240.244
R7065 gnd.n5624 gnd.n5623 240.244
R7066 gnd.n5623 gnd.n5622 240.244
R7067 gnd.n5622 gnd.n5457 240.244
R7068 gnd.n5618 gnd.n5457 240.244
R7069 gnd.n5618 gnd.n5463 240.244
R7070 gnd.n5484 gnd.n5463 240.244
R7071 gnd.n5484 gnd.n5481 240.244
R7072 gnd.n5490 gnd.n5481 240.244
R7073 gnd.n5491 gnd.n5490 240.244
R7074 gnd.n5492 gnd.n5491 240.244
R7075 gnd.n5492 gnd.n5476 240.244
R7076 gnd.n5596 gnd.n5476 240.244
R7077 gnd.n5596 gnd.n5477 240.244
R7078 gnd.n5592 gnd.n5477 240.244
R7079 gnd.n5592 gnd.n5591 240.244
R7080 gnd.n5591 gnd.n5590 240.244
R7081 gnd.n5590 gnd.n5500 240.244
R7082 gnd.n5586 gnd.n5500 240.244
R7083 gnd.n5586 gnd.n5585 240.244
R7084 gnd.n5585 gnd.n5584 240.244
R7085 gnd.n5584 gnd.n5506 240.244
R7086 gnd.n5534 gnd.n5506 240.244
R7087 gnd.n5574 gnd.n5534 240.244
R7088 gnd.n5574 gnd.n5535 240.244
R7089 gnd.n5556 gnd.n5535 240.244
R7090 gnd.n5567 gnd.n5556 240.244
R7091 gnd.n5567 gnd.n5566 240.244
R7092 gnd.n5566 gnd.n5565 240.244
R7093 gnd.n5565 gnd.n5563 240.244
R7094 gnd.n5563 gnd.n5560 240.244
R7095 gnd.n5560 gnd.n5559 240.244
R7096 gnd.n5559 gnd.n553 240.244
R7097 gnd.n6835 gnd.n553 240.244
R7098 gnd.n6835 gnd.n554 240.244
R7099 gnd.n6831 gnd.n554 240.244
R7100 gnd.n6831 gnd.n6830 240.244
R7101 gnd.n6830 gnd.n6829 240.244
R7102 gnd.n6829 gnd.n559 240.244
R7103 gnd.n6190 gnd.n942 240.244
R7104 gnd.n6186 gnd.n942 240.244
R7105 gnd.n6186 gnd.n944 240.244
R7106 gnd.n6182 gnd.n944 240.244
R7107 gnd.n6182 gnd.n949 240.244
R7108 gnd.n6178 gnd.n949 240.244
R7109 gnd.n6178 gnd.n951 240.244
R7110 gnd.n6174 gnd.n951 240.244
R7111 gnd.n6174 gnd.n957 240.244
R7112 gnd.n6170 gnd.n957 240.244
R7113 gnd.n6170 gnd.n959 240.244
R7114 gnd.n6166 gnd.n959 240.244
R7115 gnd.n6166 gnd.n965 240.244
R7116 gnd.n6162 gnd.n965 240.244
R7117 gnd.n6162 gnd.n967 240.244
R7118 gnd.n6158 gnd.n967 240.244
R7119 gnd.n6158 gnd.n973 240.244
R7120 gnd.n6154 gnd.n973 240.244
R7121 gnd.n6154 gnd.n975 240.244
R7122 gnd.n6150 gnd.n975 240.244
R7123 gnd.n6150 gnd.n981 240.244
R7124 gnd.n6146 gnd.n981 240.244
R7125 gnd.n6146 gnd.n983 240.244
R7126 gnd.n6142 gnd.n983 240.244
R7127 gnd.n6142 gnd.n989 240.244
R7128 gnd.n6138 gnd.n989 240.244
R7129 gnd.n6138 gnd.n991 240.244
R7130 gnd.n6134 gnd.n991 240.244
R7131 gnd.n6134 gnd.n997 240.244
R7132 gnd.n6130 gnd.n997 240.244
R7133 gnd.n6130 gnd.n999 240.244
R7134 gnd.n6126 gnd.n999 240.244
R7135 gnd.n6126 gnd.n1005 240.244
R7136 gnd.n6122 gnd.n1005 240.244
R7137 gnd.n6122 gnd.n1007 240.244
R7138 gnd.n6118 gnd.n1007 240.244
R7139 gnd.n6118 gnd.n1013 240.244
R7140 gnd.n6114 gnd.n1013 240.244
R7141 gnd.n6114 gnd.n1015 240.244
R7142 gnd.n6110 gnd.n1015 240.244
R7143 gnd.n6110 gnd.n1021 240.244
R7144 gnd.n6106 gnd.n1021 240.244
R7145 gnd.n6106 gnd.n1023 240.244
R7146 gnd.n6102 gnd.n1023 240.244
R7147 gnd.n6102 gnd.n1029 240.244
R7148 gnd.n6098 gnd.n1029 240.244
R7149 gnd.n6098 gnd.n1031 240.244
R7150 gnd.n6094 gnd.n1031 240.244
R7151 gnd.n6094 gnd.n1037 240.244
R7152 gnd.n6090 gnd.n1037 240.244
R7153 gnd.n6090 gnd.n1039 240.244
R7154 gnd.n6086 gnd.n1039 240.244
R7155 gnd.n6086 gnd.n1045 240.244
R7156 gnd.n6082 gnd.n1045 240.244
R7157 gnd.n6082 gnd.n1047 240.244
R7158 gnd.n6078 gnd.n1047 240.244
R7159 gnd.n6078 gnd.n1053 240.244
R7160 gnd.n6074 gnd.n1053 240.244
R7161 gnd.n6074 gnd.n1055 240.244
R7162 gnd.n6070 gnd.n1055 240.244
R7163 gnd.n6070 gnd.n1061 240.244
R7164 gnd.n6066 gnd.n1061 240.244
R7165 gnd.n6066 gnd.n1063 240.244
R7166 gnd.n6062 gnd.n1063 240.244
R7167 gnd.n6062 gnd.n1069 240.244
R7168 gnd.n6058 gnd.n1069 240.244
R7169 gnd.n6058 gnd.n1071 240.244
R7170 gnd.n6054 gnd.n1071 240.244
R7171 gnd.n6054 gnd.n1077 240.244
R7172 gnd.n6050 gnd.n1077 240.244
R7173 gnd.n6050 gnd.n1079 240.244
R7174 gnd.n6046 gnd.n1079 240.244
R7175 gnd.n6046 gnd.n1085 240.244
R7176 gnd.n6042 gnd.n1085 240.244
R7177 gnd.n6042 gnd.n1087 240.244
R7178 gnd.n6038 gnd.n1087 240.244
R7179 gnd.n6038 gnd.n1093 240.244
R7180 gnd.n6034 gnd.n1093 240.244
R7181 gnd.n6034 gnd.n1095 240.244
R7182 gnd.n6030 gnd.n1095 240.244
R7183 gnd.n6030 gnd.n1101 240.244
R7184 gnd.n6026 gnd.n1101 240.244
R7185 gnd.n6026 gnd.n1103 240.244
R7186 gnd.n6022 gnd.n1103 240.244
R7187 gnd.n4614 gnd.n2199 240.244
R7188 gnd.n4614 gnd.n2189 240.244
R7189 gnd.n4627 gnd.n2189 240.244
R7190 gnd.n4627 gnd.n2185 240.244
R7191 gnd.n4633 gnd.n2185 240.244
R7192 gnd.n4633 gnd.n2175 240.244
R7193 gnd.n4646 gnd.n2175 240.244
R7194 gnd.n4646 gnd.n2171 240.244
R7195 gnd.n4652 gnd.n2171 240.244
R7196 gnd.n4652 gnd.n1989 240.244
R7197 gnd.n4672 gnd.n1989 240.244
R7198 gnd.n4672 gnd.n1983 240.244
R7199 gnd.n4687 gnd.n1983 240.244
R7200 gnd.n4687 gnd.n1984 240.244
R7201 gnd.n4677 gnd.n1984 240.244
R7202 gnd.n4680 gnd.n4677 240.244
R7203 gnd.n4680 gnd.n1928 240.244
R7204 gnd.n4732 gnd.n1928 240.244
R7205 gnd.n4732 gnd.n1922 240.244
R7206 gnd.n4739 gnd.n1922 240.244
R7207 gnd.n4739 gnd.n1923 240.244
R7208 gnd.n1923 gnd.n1902 240.244
R7209 gnd.n4801 gnd.n1902 240.244
R7210 gnd.n4801 gnd.n1896 240.244
R7211 gnd.n4808 gnd.n1896 240.244
R7212 gnd.n4808 gnd.n1897 240.244
R7213 gnd.n1897 gnd.n1872 240.244
R7214 gnd.n4837 gnd.n1872 240.244
R7215 gnd.n4837 gnd.n1868 240.244
R7216 gnd.n4843 gnd.n1868 240.244
R7217 gnd.n4843 gnd.n1849 240.244
R7218 gnd.n4869 gnd.n1849 240.244
R7219 gnd.n4869 gnd.n1843 240.244
R7220 gnd.n4885 gnd.n1843 240.244
R7221 gnd.n4885 gnd.n1844 240.244
R7222 gnd.n4874 gnd.n1844 240.244
R7223 gnd.n4875 gnd.n4874 240.244
R7224 gnd.n4876 gnd.n4875 240.244
R7225 gnd.n4876 gnd.n1810 240.244
R7226 gnd.n5027 gnd.n1810 240.244
R7227 gnd.n5027 gnd.n1804 240.244
R7228 gnd.n5034 gnd.n1804 240.244
R7229 gnd.n5034 gnd.n1805 240.244
R7230 gnd.n1805 gnd.n1780 240.244
R7231 gnd.n5063 gnd.n1780 240.244
R7232 gnd.n5063 gnd.n1776 240.244
R7233 gnd.n5069 gnd.n1776 240.244
R7234 gnd.n5069 gnd.n1758 240.244
R7235 gnd.n5090 gnd.n1758 240.244
R7236 gnd.n5090 gnd.n1754 240.244
R7237 gnd.n5096 gnd.n1754 240.244
R7238 gnd.n5096 gnd.n1736 240.244
R7239 gnd.n5120 gnd.n1736 240.244
R7240 gnd.n5120 gnd.n1732 240.244
R7241 gnd.n5126 gnd.n1732 240.244
R7242 gnd.n5126 gnd.n1715 240.244
R7243 gnd.n5150 gnd.n1715 240.244
R7244 gnd.n5150 gnd.n1709 240.244
R7245 gnd.n5157 gnd.n1709 240.244
R7246 gnd.n5157 gnd.n1710 240.244
R7247 gnd.n1710 gnd.n1686 240.244
R7248 gnd.n5186 gnd.n1686 240.244
R7249 gnd.n5186 gnd.n1682 240.244
R7250 gnd.n5192 gnd.n1682 240.244
R7251 gnd.n5192 gnd.n1662 240.244
R7252 gnd.n5225 gnd.n1662 240.244
R7253 gnd.n5225 gnd.n1658 240.244
R7254 gnd.n5231 gnd.n1658 240.244
R7255 gnd.n5231 gnd.n1606 240.244
R7256 gnd.n5396 gnd.n1606 240.244
R7257 gnd.n5396 gnd.n1602 240.244
R7258 gnd.n5402 gnd.n1602 240.244
R7259 gnd.n5402 gnd.n1591 240.244
R7260 gnd.n5415 gnd.n1591 240.244
R7261 gnd.n5415 gnd.n1587 240.244
R7262 gnd.n5421 gnd.n1587 240.244
R7263 gnd.n5421 gnd.n1578 240.244
R7264 gnd.n5437 gnd.n1578 240.244
R7265 gnd.n5437 gnd.n1574 240.244
R7266 gnd.n5443 gnd.n1574 240.244
R7267 gnd.n5443 gnd.n1473 240.244
R7268 gnd.n5707 gnd.n1473 240.244
R7269 gnd.n2210 gnd.n2209 240.244
R7270 gnd.n2265 gnd.n2210 240.244
R7271 gnd.n2220 gnd.n2219 240.244
R7272 gnd.n2267 gnd.n2230 240.244
R7273 gnd.n2270 gnd.n2231 240.244
R7274 gnd.n2241 gnd.n2240 240.244
R7275 gnd.n2272 gnd.n2251 240.244
R7276 gnd.n2263 gnd.n2252 240.244
R7277 gnd.n4559 gnd.n2262 240.244
R7278 gnd.n1351 gnd.n1350 240.244
R7279 gnd.n2277 gnd.n1352 240.244
R7280 gnd.n1356 gnd.n1355 240.244
R7281 gnd.n1362 gnd.n1357 240.244
R7282 gnd.n1364 gnd.n1363 240.244
R7283 gnd.n1368 gnd.n1367 240.244
R7284 gnd.n1369 gnd.n1368 240.244
R7285 gnd.n2191 gnd.n1369 240.244
R7286 gnd.n2191 gnd.n1372 240.244
R7287 gnd.n1373 gnd.n1372 240.244
R7288 gnd.n1374 gnd.n1373 240.244
R7289 gnd.n2177 gnd.n1374 240.244
R7290 gnd.n2177 gnd.n1377 240.244
R7291 gnd.n1378 gnd.n1377 240.244
R7292 gnd.n1379 gnd.n1378 240.244
R7293 gnd.n1990 gnd.n1379 240.244
R7294 gnd.n1990 gnd.n1382 240.244
R7295 gnd.n1383 gnd.n1382 240.244
R7296 gnd.n1384 gnd.n1383 240.244
R7297 gnd.n1947 gnd.n1384 240.244
R7298 gnd.n1947 gnd.n1387 240.244
R7299 gnd.n1388 gnd.n1387 240.244
R7300 gnd.n1389 gnd.n1388 240.244
R7301 gnd.n1932 gnd.n1389 240.244
R7302 gnd.n1932 gnd.n1392 240.244
R7303 gnd.n1393 gnd.n1392 240.244
R7304 gnd.n1394 gnd.n1393 240.244
R7305 gnd.n1904 gnd.n1394 240.244
R7306 gnd.n1904 gnd.n1397 240.244
R7307 gnd.n1398 gnd.n1397 240.244
R7308 gnd.n1399 gnd.n1398 240.244
R7309 gnd.n1879 gnd.n1399 240.244
R7310 gnd.n1879 gnd.n1402 240.244
R7311 gnd.n1403 gnd.n1402 240.244
R7312 gnd.n1404 gnd.n1403 240.244
R7313 gnd.n1859 gnd.n1404 240.244
R7314 gnd.n1859 gnd.n1407 240.244
R7315 gnd.n1408 gnd.n1407 240.244
R7316 gnd.n1409 gnd.n1408 240.244
R7317 gnd.n1838 gnd.n1409 240.244
R7318 gnd.n1838 gnd.n1412 240.244
R7319 gnd.n1413 gnd.n1412 240.244
R7320 gnd.n1414 gnd.n1413 240.244
R7321 gnd.n4996 gnd.n1414 240.244
R7322 gnd.n4996 gnd.n1417 240.244
R7323 gnd.n1418 gnd.n1417 240.244
R7324 gnd.n1419 gnd.n1418 240.244
R7325 gnd.n1797 gnd.n1419 240.244
R7326 gnd.n1797 gnd.n1422 240.244
R7327 gnd.n1423 gnd.n1422 240.244
R7328 gnd.n1424 gnd.n1423 240.244
R7329 gnd.n1775 gnd.n1424 240.244
R7330 gnd.n1775 gnd.n1427 240.244
R7331 gnd.n1428 gnd.n1427 240.244
R7332 gnd.n1429 gnd.n1428 240.244
R7333 gnd.n1753 gnd.n1429 240.244
R7334 gnd.n1753 gnd.n1432 240.244
R7335 gnd.n1433 gnd.n1432 240.244
R7336 gnd.n1434 gnd.n1433 240.244
R7337 gnd.n1731 gnd.n1434 240.244
R7338 gnd.n1731 gnd.n1437 240.244
R7339 gnd.n1438 gnd.n1437 240.244
R7340 gnd.n1439 gnd.n1438 240.244
R7341 gnd.n1708 gnd.n1439 240.244
R7342 gnd.n1708 gnd.n1442 240.244
R7343 gnd.n1443 gnd.n1442 240.244
R7344 gnd.n1444 gnd.n1443 240.244
R7345 gnd.n4931 gnd.n1444 240.244
R7346 gnd.n4931 gnd.n1447 240.244
R7347 gnd.n1448 gnd.n1447 240.244
R7348 gnd.n1449 gnd.n1448 240.244
R7349 gnd.n1664 gnd.n1449 240.244
R7350 gnd.n1664 gnd.n1452 240.244
R7351 gnd.n1453 gnd.n1452 240.244
R7352 gnd.n1454 gnd.n1453 240.244
R7353 gnd.n1625 gnd.n1454 240.244
R7354 gnd.n1625 gnd.n1457 240.244
R7355 gnd.n1458 gnd.n1457 240.244
R7356 gnd.n1459 gnd.n1458 240.244
R7357 gnd.n1593 gnd.n1459 240.244
R7358 gnd.n1593 gnd.n1462 240.244
R7359 gnd.n1463 gnd.n1462 240.244
R7360 gnd.n1464 gnd.n1463 240.244
R7361 gnd.n1580 gnd.n1464 240.244
R7362 gnd.n1580 gnd.n1467 240.244
R7363 gnd.n1468 gnd.n1467 240.244
R7364 gnd.n5709 gnd.n1468 240.244
R7365 gnd.n1485 gnd.n1484 240.244
R7366 gnd.n1546 gnd.n1494 240.244
R7367 gnd.n1549 gnd.n1495 240.244
R7368 gnd.n1503 gnd.n1502 240.244
R7369 gnd.n1551 gnd.n1512 240.244
R7370 gnd.n1554 gnd.n1513 240.244
R7371 gnd.n1521 gnd.n1520 240.244
R7372 gnd.n1556 gnd.n1528 240.244
R7373 gnd.n1530 gnd.n1529 240.244
R7374 gnd.n1560 gnd.n1531 240.244
R7375 gnd.n1535 gnd.n1534 240.244
R7376 gnd.n1563 gnd.n1536 240.244
R7377 gnd.n1543 gnd.n1542 240.244
R7378 gnd.n5632 gnd.n1470 240.244
R7379 gnd.n1965 gnd.n1964 240.132
R7380 gnd.n5248 gnd.n5247 240.132
R7381 gnd.n6197 gnd.n937 225.874
R7382 gnd.n6198 gnd.n6197 225.874
R7383 gnd.n6199 gnd.n6198 225.874
R7384 gnd.n6199 gnd.n931 225.874
R7385 gnd.n6207 gnd.n931 225.874
R7386 gnd.n6208 gnd.n6207 225.874
R7387 gnd.n6209 gnd.n6208 225.874
R7388 gnd.n6209 gnd.n925 225.874
R7389 gnd.n6217 gnd.n925 225.874
R7390 gnd.n6218 gnd.n6217 225.874
R7391 gnd.n6219 gnd.n6218 225.874
R7392 gnd.n6219 gnd.n919 225.874
R7393 gnd.n6227 gnd.n919 225.874
R7394 gnd.n6228 gnd.n6227 225.874
R7395 gnd.n6229 gnd.n6228 225.874
R7396 gnd.n6229 gnd.n913 225.874
R7397 gnd.n6237 gnd.n913 225.874
R7398 gnd.n6238 gnd.n6237 225.874
R7399 gnd.n6239 gnd.n6238 225.874
R7400 gnd.n6239 gnd.n907 225.874
R7401 gnd.n6247 gnd.n907 225.874
R7402 gnd.n6248 gnd.n6247 225.874
R7403 gnd.n6249 gnd.n6248 225.874
R7404 gnd.n6249 gnd.n901 225.874
R7405 gnd.n6257 gnd.n901 225.874
R7406 gnd.n6258 gnd.n6257 225.874
R7407 gnd.n6259 gnd.n6258 225.874
R7408 gnd.n6259 gnd.n895 225.874
R7409 gnd.n6267 gnd.n895 225.874
R7410 gnd.n6268 gnd.n6267 225.874
R7411 gnd.n6269 gnd.n6268 225.874
R7412 gnd.n6269 gnd.n889 225.874
R7413 gnd.n6277 gnd.n889 225.874
R7414 gnd.n6278 gnd.n6277 225.874
R7415 gnd.n6279 gnd.n6278 225.874
R7416 gnd.n6279 gnd.n883 225.874
R7417 gnd.n6287 gnd.n883 225.874
R7418 gnd.n6288 gnd.n6287 225.874
R7419 gnd.n6289 gnd.n6288 225.874
R7420 gnd.n6289 gnd.n877 225.874
R7421 gnd.n6297 gnd.n877 225.874
R7422 gnd.n6298 gnd.n6297 225.874
R7423 gnd.n6299 gnd.n6298 225.874
R7424 gnd.n6299 gnd.n871 225.874
R7425 gnd.n6307 gnd.n871 225.874
R7426 gnd.n6308 gnd.n6307 225.874
R7427 gnd.n6309 gnd.n6308 225.874
R7428 gnd.n6309 gnd.n865 225.874
R7429 gnd.n6317 gnd.n865 225.874
R7430 gnd.n6318 gnd.n6317 225.874
R7431 gnd.n6319 gnd.n6318 225.874
R7432 gnd.n6319 gnd.n859 225.874
R7433 gnd.n6327 gnd.n859 225.874
R7434 gnd.n6328 gnd.n6327 225.874
R7435 gnd.n6329 gnd.n6328 225.874
R7436 gnd.n6329 gnd.n853 225.874
R7437 gnd.n6337 gnd.n853 225.874
R7438 gnd.n6338 gnd.n6337 225.874
R7439 gnd.n6339 gnd.n6338 225.874
R7440 gnd.n6339 gnd.n847 225.874
R7441 gnd.n6347 gnd.n847 225.874
R7442 gnd.n6348 gnd.n6347 225.874
R7443 gnd.n6349 gnd.n6348 225.874
R7444 gnd.n6349 gnd.n841 225.874
R7445 gnd.n6357 gnd.n841 225.874
R7446 gnd.n6358 gnd.n6357 225.874
R7447 gnd.n6359 gnd.n6358 225.874
R7448 gnd.n6359 gnd.n835 225.874
R7449 gnd.n6367 gnd.n835 225.874
R7450 gnd.n6368 gnd.n6367 225.874
R7451 gnd.n6369 gnd.n6368 225.874
R7452 gnd.n6369 gnd.n829 225.874
R7453 gnd.n6377 gnd.n829 225.874
R7454 gnd.n6378 gnd.n6377 225.874
R7455 gnd.n6379 gnd.n6378 225.874
R7456 gnd.n6379 gnd.n823 225.874
R7457 gnd.n6387 gnd.n823 225.874
R7458 gnd.n6388 gnd.n6387 225.874
R7459 gnd.n6389 gnd.n6388 225.874
R7460 gnd.n6389 gnd.n817 225.874
R7461 gnd.n6397 gnd.n817 225.874
R7462 gnd.n6398 gnd.n6397 225.874
R7463 gnd.n6399 gnd.n6398 225.874
R7464 gnd.n6399 gnd.n811 225.874
R7465 gnd.n6407 gnd.n811 225.874
R7466 gnd.n6408 gnd.n6407 225.874
R7467 gnd.n6409 gnd.n6408 225.874
R7468 gnd.n6409 gnd.n805 225.874
R7469 gnd.n6417 gnd.n805 225.874
R7470 gnd.n6418 gnd.n6417 225.874
R7471 gnd.n6419 gnd.n6418 225.874
R7472 gnd.n6419 gnd.n799 225.874
R7473 gnd.n6427 gnd.n799 225.874
R7474 gnd.n6428 gnd.n6427 225.874
R7475 gnd.n6429 gnd.n6428 225.874
R7476 gnd.n6429 gnd.n793 225.874
R7477 gnd.n6437 gnd.n793 225.874
R7478 gnd.n6438 gnd.n6437 225.874
R7479 gnd.n6439 gnd.n6438 225.874
R7480 gnd.n6439 gnd.n787 225.874
R7481 gnd.n6447 gnd.n787 225.874
R7482 gnd.n6448 gnd.n6447 225.874
R7483 gnd.n6449 gnd.n6448 225.874
R7484 gnd.n6449 gnd.n781 225.874
R7485 gnd.n6457 gnd.n781 225.874
R7486 gnd.n6458 gnd.n6457 225.874
R7487 gnd.n6459 gnd.n6458 225.874
R7488 gnd.n6459 gnd.n775 225.874
R7489 gnd.n6467 gnd.n775 225.874
R7490 gnd.n6468 gnd.n6467 225.874
R7491 gnd.n6469 gnd.n6468 225.874
R7492 gnd.n6469 gnd.n769 225.874
R7493 gnd.n6477 gnd.n769 225.874
R7494 gnd.n6478 gnd.n6477 225.874
R7495 gnd.n6479 gnd.n6478 225.874
R7496 gnd.n6479 gnd.n763 225.874
R7497 gnd.n6487 gnd.n763 225.874
R7498 gnd.n6488 gnd.n6487 225.874
R7499 gnd.n6489 gnd.n6488 225.874
R7500 gnd.n6489 gnd.n757 225.874
R7501 gnd.n6497 gnd.n757 225.874
R7502 gnd.n6498 gnd.n6497 225.874
R7503 gnd.n6499 gnd.n6498 225.874
R7504 gnd.n6499 gnd.n751 225.874
R7505 gnd.n6507 gnd.n751 225.874
R7506 gnd.n6508 gnd.n6507 225.874
R7507 gnd.n6509 gnd.n6508 225.874
R7508 gnd.n6509 gnd.n745 225.874
R7509 gnd.n6517 gnd.n745 225.874
R7510 gnd.n6518 gnd.n6517 225.874
R7511 gnd.n6519 gnd.n6518 225.874
R7512 gnd.n6519 gnd.n739 225.874
R7513 gnd.n6527 gnd.n739 225.874
R7514 gnd.n6528 gnd.n6527 225.874
R7515 gnd.n6529 gnd.n6528 225.874
R7516 gnd.n6529 gnd.n733 225.874
R7517 gnd.n6537 gnd.n733 225.874
R7518 gnd.n6538 gnd.n6537 225.874
R7519 gnd.n6539 gnd.n6538 225.874
R7520 gnd.n6539 gnd.n727 225.874
R7521 gnd.n6547 gnd.n727 225.874
R7522 gnd.n6548 gnd.n6547 225.874
R7523 gnd.n6549 gnd.n6548 225.874
R7524 gnd.n6549 gnd.n721 225.874
R7525 gnd.n6557 gnd.n721 225.874
R7526 gnd.n6558 gnd.n6557 225.874
R7527 gnd.n6559 gnd.n6558 225.874
R7528 gnd.n6559 gnd.n715 225.874
R7529 gnd.n6567 gnd.n715 225.874
R7530 gnd.n6568 gnd.n6567 225.874
R7531 gnd.n6569 gnd.n6568 225.874
R7532 gnd.n6569 gnd.n709 225.874
R7533 gnd.n6577 gnd.n709 225.874
R7534 gnd.n6578 gnd.n6577 225.874
R7535 gnd.n6579 gnd.n6578 225.874
R7536 gnd.n6579 gnd.n703 225.874
R7537 gnd.n6587 gnd.n703 225.874
R7538 gnd.n6588 gnd.n6587 225.874
R7539 gnd.n6589 gnd.n6588 225.874
R7540 gnd.n6589 gnd.n697 225.874
R7541 gnd.n6597 gnd.n697 225.874
R7542 gnd.n6598 gnd.n6597 225.874
R7543 gnd.n6599 gnd.n6598 225.874
R7544 gnd.n6599 gnd.n691 225.874
R7545 gnd.n6607 gnd.n691 225.874
R7546 gnd.n6608 gnd.n6607 225.874
R7547 gnd.n6609 gnd.n6608 225.874
R7548 gnd.n3013 gnd.t62 224.174
R7549 gnd.n2522 gnd.t102 224.174
R7550 gnd.n441 gnd.n402 199.319
R7551 gnd.n441 gnd.n403 199.319
R7552 gnd.n5901 gnd.n5900 199.319
R7553 gnd.n5900 gnd.n5899 199.319
R7554 gnd.n1966 gnd.n1963 186.49
R7555 gnd.n5249 gnd.n5246 186.49
R7556 gnd.n3788 gnd.n3787 185
R7557 gnd.n3786 gnd.n3785 185
R7558 gnd.n3765 gnd.n3764 185
R7559 gnd.n3780 gnd.n3779 185
R7560 gnd.n3778 gnd.n3777 185
R7561 gnd.n3769 gnd.n3768 185
R7562 gnd.n3772 gnd.n3771 185
R7563 gnd.n3756 gnd.n3755 185
R7564 gnd.n3754 gnd.n3753 185
R7565 gnd.n3733 gnd.n3732 185
R7566 gnd.n3748 gnd.n3747 185
R7567 gnd.n3746 gnd.n3745 185
R7568 gnd.n3737 gnd.n3736 185
R7569 gnd.n3740 gnd.n3739 185
R7570 gnd.n3724 gnd.n3723 185
R7571 gnd.n3722 gnd.n3721 185
R7572 gnd.n3701 gnd.n3700 185
R7573 gnd.n3716 gnd.n3715 185
R7574 gnd.n3714 gnd.n3713 185
R7575 gnd.n3705 gnd.n3704 185
R7576 gnd.n3708 gnd.n3707 185
R7577 gnd.n3693 gnd.n3692 185
R7578 gnd.n3691 gnd.n3690 185
R7579 gnd.n3670 gnd.n3669 185
R7580 gnd.n3685 gnd.n3684 185
R7581 gnd.n3683 gnd.n3682 185
R7582 gnd.n3674 gnd.n3673 185
R7583 gnd.n3677 gnd.n3676 185
R7584 gnd.n3661 gnd.n3660 185
R7585 gnd.n3659 gnd.n3658 185
R7586 gnd.n3638 gnd.n3637 185
R7587 gnd.n3653 gnd.n3652 185
R7588 gnd.n3651 gnd.n3650 185
R7589 gnd.n3642 gnd.n3641 185
R7590 gnd.n3645 gnd.n3644 185
R7591 gnd.n3629 gnd.n3628 185
R7592 gnd.n3627 gnd.n3626 185
R7593 gnd.n3606 gnd.n3605 185
R7594 gnd.n3621 gnd.n3620 185
R7595 gnd.n3619 gnd.n3618 185
R7596 gnd.n3610 gnd.n3609 185
R7597 gnd.n3613 gnd.n3612 185
R7598 gnd.n3597 gnd.n3596 185
R7599 gnd.n3595 gnd.n3594 185
R7600 gnd.n3574 gnd.n3573 185
R7601 gnd.n3589 gnd.n3588 185
R7602 gnd.n3587 gnd.n3586 185
R7603 gnd.n3578 gnd.n3577 185
R7604 gnd.n3581 gnd.n3580 185
R7605 gnd.n3566 gnd.n3565 185
R7606 gnd.n3564 gnd.n3563 185
R7607 gnd.n3543 gnd.n3542 185
R7608 gnd.n3558 gnd.n3557 185
R7609 gnd.n3556 gnd.n3555 185
R7610 gnd.n3547 gnd.n3546 185
R7611 gnd.n3550 gnd.n3549 185
R7612 gnd.n3014 gnd.t61 178.987
R7613 gnd.n2523 gnd.t103 178.987
R7614 gnd.n1 gnd.t138 170.774
R7615 gnd.n7 gnd.t10 170.103
R7616 gnd.n6 gnd.t313 170.103
R7617 gnd.n5 gnd.t1 170.103
R7618 gnd.n4 gnd.t317 170.103
R7619 gnd.n3 gnd.t171 170.103
R7620 gnd.n2 gnd.t175 170.103
R7621 gnd.n1 gnd.t127 170.103
R7622 gnd.n5320 gnd.n5319 163.367
R7623 gnd.n5316 gnd.n5315 163.367
R7624 gnd.n5312 gnd.n5311 163.367
R7625 gnd.n5308 gnd.n5307 163.367
R7626 gnd.n5304 gnd.n5303 163.367
R7627 gnd.n5300 gnd.n5299 163.367
R7628 gnd.n5296 gnd.n5295 163.367
R7629 gnd.n5292 gnd.n5291 163.367
R7630 gnd.n5288 gnd.n5287 163.367
R7631 gnd.n5284 gnd.n5283 163.367
R7632 gnd.n5280 gnd.n5279 163.367
R7633 gnd.n5276 gnd.n5275 163.367
R7634 gnd.n5272 gnd.n5271 163.367
R7635 gnd.n5268 gnd.n5267 163.367
R7636 gnd.n5263 gnd.n5262 163.367
R7637 gnd.n5259 gnd.n5258 163.367
R7638 gnd.n5393 gnd.n5392 163.367
R7639 gnd.n5389 gnd.n5388 163.367
R7640 gnd.n5384 gnd.n5383 163.367
R7641 gnd.n5380 gnd.n5379 163.367
R7642 gnd.n5376 gnd.n5375 163.367
R7643 gnd.n5372 gnd.n5371 163.367
R7644 gnd.n5368 gnd.n5367 163.367
R7645 gnd.n5364 gnd.n5363 163.367
R7646 gnd.n5360 gnd.n5359 163.367
R7647 gnd.n5356 gnd.n5355 163.367
R7648 gnd.n5352 gnd.n5351 163.367
R7649 gnd.n5348 gnd.n5347 163.367
R7650 gnd.n5344 gnd.n5343 163.367
R7651 gnd.n5340 gnd.n5339 163.367
R7652 gnd.n5336 gnd.n5335 163.367
R7653 gnd.n5332 gnd.n5331 163.367
R7654 gnd.n1981 gnd.n1953 163.367
R7655 gnd.n4698 gnd.n1953 163.367
R7656 gnd.n4698 gnd.n1950 163.367
R7657 gnd.n4707 gnd.n1950 163.367
R7658 gnd.n4707 gnd.n1951 163.367
R7659 gnd.n1951 gnd.n1939 163.367
R7660 gnd.n4702 gnd.n1939 163.367
R7661 gnd.n4702 gnd.n1929 163.367
R7662 gnd.n1929 gnd.n1920 163.367
R7663 gnd.n4742 gnd.n1920 163.367
R7664 gnd.n4742 gnd.n1918 163.367
R7665 gnd.n4778 gnd.n1918 163.367
R7666 gnd.n4778 gnd.n1912 163.367
R7667 gnd.n4774 gnd.n1912 163.367
R7668 gnd.n4774 gnd.n4771 163.367
R7669 gnd.n4771 gnd.n4770 163.367
R7670 gnd.n4770 gnd.n1895 163.367
R7671 gnd.n4766 gnd.n1895 163.367
R7672 gnd.n4766 gnd.n1889 163.367
R7673 gnd.n4763 gnd.n1889 163.367
R7674 gnd.n4763 gnd.n1881 163.367
R7675 gnd.n4758 gnd.n1881 163.367
R7676 gnd.n4758 gnd.n1874 163.367
R7677 gnd.n4755 gnd.n1874 163.367
R7678 gnd.n4755 gnd.n1867 163.367
R7679 gnd.n4750 gnd.n1867 163.367
R7680 gnd.n4750 gnd.n1860 163.367
R7681 gnd.n4747 gnd.n1860 163.367
R7682 gnd.n4747 gnd.n1852 163.367
R7683 gnd.n1852 gnd.n1841 163.367
R7684 gnd.n4888 gnd.n1841 163.367
R7685 gnd.n4888 gnd.n1834 163.367
R7686 gnd.n4892 gnd.n1834 163.367
R7687 gnd.n4892 gnd.n1827 163.367
R7688 gnd.n4912 gnd.n1827 163.367
R7689 gnd.n4912 gnd.n1825 163.367
R7690 gnd.n5004 gnd.n1825 163.367
R7691 gnd.n5004 gnd.n1819 163.367
R7692 gnd.n5000 gnd.n1819 163.367
R7693 gnd.n5000 gnd.n4995 163.367
R7694 gnd.n4995 gnd.n4994 163.367
R7695 gnd.n4994 gnd.n1803 163.367
R7696 gnd.n4990 gnd.n1803 163.367
R7697 gnd.n4990 gnd.n1796 163.367
R7698 gnd.n4987 gnd.n1796 163.367
R7699 gnd.n4987 gnd.n1788 163.367
R7700 gnd.n4982 gnd.n1788 163.367
R7701 gnd.n4982 gnd.n1782 163.367
R7702 gnd.n4979 gnd.n1782 163.367
R7703 gnd.n4979 gnd.n1774 163.367
R7704 gnd.n4974 gnd.n1774 163.367
R7705 gnd.n4974 gnd.n1767 163.367
R7706 gnd.n4971 gnd.n1767 163.367
R7707 gnd.n4971 gnd.n1760 163.367
R7708 gnd.n1760 gnd.n1751 163.367
R7709 gnd.n1752 gnd.n1751 163.367
R7710 gnd.n1752 gnd.n1744 163.367
R7711 gnd.n4965 gnd.n1744 163.367
R7712 gnd.n4965 gnd.n4962 163.367
R7713 gnd.n4962 gnd.n4961 163.367
R7714 gnd.n4961 gnd.n1729 163.367
R7715 gnd.n1730 gnd.n1729 163.367
R7716 gnd.n1730 gnd.n1722 163.367
R7717 gnd.n4955 gnd.n1722 163.367
R7718 gnd.n4955 gnd.n4952 163.367
R7719 gnd.n4952 gnd.n4951 163.367
R7720 gnd.n4951 gnd.n1707 163.367
R7721 gnd.n4946 gnd.n1707 163.367
R7722 gnd.n4946 gnd.n1701 163.367
R7723 gnd.n4943 gnd.n1701 163.367
R7724 gnd.n4943 gnd.n1693 163.367
R7725 gnd.n4938 gnd.n1693 163.367
R7726 gnd.n4938 gnd.n1687 163.367
R7727 gnd.n4934 gnd.n1687 163.367
R7728 gnd.n4934 gnd.n1681 163.367
R7729 gnd.n4928 gnd.n1681 163.367
R7730 gnd.n4928 gnd.n1674 163.367
R7731 gnd.n4925 gnd.n1674 163.367
R7732 gnd.n4925 gnd.n1666 163.367
R7733 gnd.n4921 gnd.n1666 163.367
R7734 gnd.n4921 gnd.n1655 163.367
R7735 gnd.n1655 gnd.n1648 163.367
R7736 gnd.n5327 gnd.n1648 163.367
R7737 gnd.n2159 gnd.n2023 163.367
R7738 gnd.n2155 gnd.n2023 163.367
R7739 gnd.n2153 gnd.n2152 163.367
R7740 gnd.n2149 gnd.n2148 163.367
R7741 gnd.n2145 gnd.n2144 163.367
R7742 gnd.n2141 gnd.n2140 163.367
R7743 gnd.n2137 gnd.n2136 163.367
R7744 gnd.n2133 gnd.n2132 163.367
R7745 gnd.n2129 gnd.n2128 163.367
R7746 gnd.n2125 gnd.n2124 163.367
R7747 gnd.n2121 gnd.n2120 163.367
R7748 gnd.n2117 gnd.n2116 163.367
R7749 gnd.n2113 gnd.n2112 163.367
R7750 gnd.n2109 gnd.n2108 163.367
R7751 gnd.n2105 gnd.n2104 163.367
R7752 gnd.n2101 gnd.n2100 163.367
R7753 gnd.n2097 gnd.n2096 163.367
R7754 gnd.n2092 gnd.n2091 163.367
R7755 gnd.n2087 gnd.n2086 163.367
R7756 gnd.n2083 gnd.n2082 163.367
R7757 gnd.n2079 gnd.n2078 163.367
R7758 gnd.n2075 gnd.n2074 163.367
R7759 gnd.n2071 gnd.n2070 163.367
R7760 gnd.n2067 gnd.n2066 163.367
R7761 gnd.n2063 gnd.n2062 163.367
R7762 gnd.n2059 gnd.n2058 163.367
R7763 gnd.n2055 gnd.n2054 163.367
R7764 gnd.n2051 gnd.n2050 163.367
R7765 gnd.n2047 gnd.n2046 163.367
R7766 gnd.n2043 gnd.n2042 163.367
R7767 gnd.n2039 gnd.n2038 163.367
R7768 gnd.n2035 gnd.n2034 163.367
R7769 gnd.n4690 gnd.n1955 163.367
R7770 gnd.n4696 gnd.n1955 163.367
R7771 gnd.n4696 gnd.n1958 163.367
R7772 gnd.n1958 gnd.n1949 163.367
R7773 gnd.n1949 gnd.n1937 163.367
R7774 gnd.n4724 gnd.n1937 163.367
R7775 gnd.n4724 gnd.n1931 163.367
R7776 gnd.n4729 gnd.n1931 163.367
R7777 gnd.n4729 gnd.n1935 163.367
R7778 gnd.n1935 gnd.n1917 163.367
R7779 gnd.n4782 gnd.n1917 163.367
R7780 gnd.n4782 gnd.n1914 163.367
R7781 gnd.n4789 gnd.n1914 163.367
R7782 gnd.n4789 gnd.n1915 163.367
R7783 gnd.n4785 gnd.n1915 163.367
R7784 gnd.n4785 gnd.n1893 163.367
R7785 gnd.n4812 gnd.n1893 163.367
R7786 gnd.n4812 gnd.n1891 163.367
R7787 gnd.n4816 gnd.n1891 163.367
R7788 gnd.n4816 gnd.n1878 163.367
R7789 gnd.n4830 gnd.n1878 163.367
R7790 gnd.n4830 gnd.n1876 163.367
R7791 gnd.n4834 gnd.n1876 163.367
R7792 gnd.n4834 gnd.n1865 163.367
R7793 gnd.n4846 gnd.n1865 163.367
R7794 gnd.n4846 gnd.n1862 163.367
R7795 gnd.n4856 gnd.n1862 163.367
R7796 gnd.n4856 gnd.n1863 163.367
R7797 gnd.n1863 gnd.n1851 163.367
R7798 gnd.n4851 gnd.n1851 163.367
R7799 gnd.n4851 gnd.n1835 163.367
R7800 gnd.n4900 gnd.n1835 163.367
R7801 gnd.n4900 gnd.n1836 163.367
R7802 gnd.n4896 gnd.n1836 163.367
R7803 gnd.n4896 gnd.n1823 163.367
R7804 gnd.n5008 gnd.n1823 163.367
R7805 gnd.n5008 gnd.n1820 163.367
R7806 gnd.n5015 gnd.n1820 163.367
R7807 gnd.n5015 gnd.n1821 163.367
R7808 gnd.n5011 gnd.n1821 163.367
R7809 gnd.n5011 gnd.n1801 163.367
R7810 gnd.n5038 gnd.n1801 163.367
R7811 gnd.n5038 gnd.n1799 163.367
R7812 gnd.n5042 gnd.n1799 163.367
R7813 gnd.n5042 gnd.n1786 163.367
R7814 gnd.n5056 gnd.n1786 163.367
R7815 gnd.n5056 gnd.n1784 163.367
R7816 gnd.n5060 gnd.n1784 163.367
R7817 gnd.n5060 gnd.n1772 163.367
R7818 gnd.n5072 gnd.n1772 163.367
R7819 gnd.n5072 gnd.n1769 163.367
R7820 gnd.n5077 gnd.n1769 163.367
R7821 gnd.n5077 gnd.n1770 163.367
R7822 gnd.n1770 gnd.n1749 163.367
R7823 gnd.n5101 gnd.n1749 163.367
R7824 gnd.n5101 gnd.n1746 163.367
R7825 gnd.n5108 gnd.n1746 163.367
R7826 gnd.n5108 gnd.n1747 163.367
R7827 gnd.n5104 gnd.n1747 163.367
R7828 gnd.n5104 gnd.n1727 163.367
R7829 gnd.n5131 gnd.n1727 163.367
R7830 gnd.n5131 gnd.n1724 163.367
R7831 gnd.n5138 gnd.n1724 163.367
R7832 gnd.n5138 gnd.n1725 163.367
R7833 gnd.n5134 gnd.n1725 163.367
R7834 gnd.n5134 gnd.n1705 163.367
R7835 gnd.n5161 gnd.n1705 163.367
R7836 gnd.n5161 gnd.n1703 163.367
R7837 gnd.n5165 gnd.n1703 163.367
R7838 gnd.n5165 gnd.n1691 163.367
R7839 gnd.n5179 gnd.n1691 163.367
R7840 gnd.n5179 gnd.n1689 163.367
R7841 gnd.n5183 gnd.n1689 163.367
R7842 gnd.n5183 gnd.n1679 163.367
R7843 gnd.n5195 gnd.n1679 163.367
R7844 gnd.n5195 gnd.n1676 163.367
R7845 gnd.n5201 gnd.n1676 163.367
R7846 gnd.n5201 gnd.n1677 163.367
R7847 gnd.n1677 gnd.n1663 163.367
R7848 gnd.n1663 gnd.n1653 163.367
R7849 gnd.n5234 gnd.n1653 163.367
R7850 gnd.n5234 gnd.n1650 163.367
R7851 gnd.n5325 gnd.n1650 163.367
R7852 gnd.n5255 gnd.n5254 156.462
R7853 gnd.n3728 gnd.n3696 153.042
R7854 gnd.n3792 gnd.n3791 152.079
R7855 gnd.n3760 gnd.n3759 152.079
R7856 gnd.n3728 gnd.n3727 152.079
R7857 gnd.n1971 gnd.n1970 152
R7858 gnd.n1972 gnd.n1961 152
R7859 gnd.n1974 gnd.n1973 152
R7860 gnd.n1976 gnd.n1959 152
R7861 gnd.n1978 gnd.n1977 152
R7862 gnd.n5253 gnd.n5237 152
R7863 gnd.n5245 gnd.n5238 152
R7864 gnd.n5244 gnd.n5243 152
R7865 gnd.n5242 gnd.n5239 152
R7866 gnd.n5240 gnd.t77 150.546
R7867 gnd.t140 gnd.n3770 147.661
R7868 gnd.t173 gnd.n3738 147.661
R7869 gnd.t145 gnd.n3706 147.661
R7870 gnd.t311 gnd.n3675 147.661
R7871 gnd.t16 gnd.n3643 147.661
R7872 gnd.t147 gnd.n3611 147.661
R7873 gnd.t149 gnd.n3579 147.661
R7874 gnd.t134 gnd.n3548 147.661
R7875 gnd.n1644 gnd.n1624 143.351
R7876 gnd.n2095 gnd.n2005 143.351
R7877 gnd.n2095 gnd.n2006 143.351
R7878 gnd.n6617 gnd.n685 137.715
R7879 gnd.n6618 gnd.n6617 137.715
R7880 gnd.n6619 gnd.n6618 137.715
R7881 gnd.n6619 gnd.n679 137.715
R7882 gnd.n6627 gnd.n679 137.715
R7883 gnd.n6628 gnd.n6627 137.715
R7884 gnd.n6629 gnd.n6628 137.715
R7885 gnd.n6629 gnd.n673 137.715
R7886 gnd.n6637 gnd.n673 137.715
R7887 gnd.n6638 gnd.n6637 137.715
R7888 gnd.n6639 gnd.n6638 137.715
R7889 gnd.n6639 gnd.n667 137.715
R7890 gnd.n6647 gnd.n667 137.715
R7891 gnd.n6648 gnd.n6647 137.715
R7892 gnd.n6649 gnd.n6648 137.715
R7893 gnd.n6649 gnd.n661 137.715
R7894 gnd.n6657 gnd.n661 137.715
R7895 gnd.n6658 gnd.n6657 137.715
R7896 gnd.n6659 gnd.n6658 137.715
R7897 gnd.n6659 gnd.n655 137.715
R7898 gnd.n6667 gnd.n655 137.715
R7899 gnd.n6668 gnd.n6667 137.715
R7900 gnd.n6669 gnd.n6668 137.715
R7901 gnd.n6669 gnd.n649 137.715
R7902 gnd.n6677 gnd.n649 137.715
R7903 gnd.n6678 gnd.n6677 137.715
R7904 gnd.n6679 gnd.n6678 137.715
R7905 gnd.n6679 gnd.n643 137.715
R7906 gnd.n6687 gnd.n643 137.715
R7907 gnd.n6688 gnd.n6687 137.715
R7908 gnd.n6689 gnd.n6688 137.715
R7909 gnd.n6689 gnd.n637 137.715
R7910 gnd.n6697 gnd.n637 137.715
R7911 gnd.n6698 gnd.n6697 137.715
R7912 gnd.n6699 gnd.n6698 137.715
R7913 gnd.n6699 gnd.n631 137.715
R7914 gnd.n6707 gnd.n631 137.715
R7915 gnd.n6708 gnd.n6707 137.715
R7916 gnd.n6709 gnd.n6708 137.715
R7917 gnd.n6709 gnd.n625 137.715
R7918 gnd.n6717 gnd.n625 137.715
R7919 gnd.n6718 gnd.n6717 137.715
R7920 gnd.n6719 gnd.n6718 137.715
R7921 gnd.n6719 gnd.n619 137.715
R7922 gnd.n6727 gnd.n619 137.715
R7923 gnd.n6728 gnd.n6727 137.715
R7924 gnd.n6729 gnd.n6728 137.715
R7925 gnd.n6729 gnd.n613 137.715
R7926 gnd.n6737 gnd.n613 137.715
R7927 gnd.n6738 gnd.n6737 137.715
R7928 gnd.n6739 gnd.n6738 137.715
R7929 gnd.n6739 gnd.n607 137.715
R7930 gnd.n6747 gnd.n607 137.715
R7931 gnd.n6748 gnd.n6747 137.715
R7932 gnd.n6749 gnd.n6748 137.715
R7933 gnd.n6749 gnd.n601 137.715
R7934 gnd.n6757 gnd.n601 137.715
R7935 gnd.n6758 gnd.n6757 137.715
R7936 gnd.n6759 gnd.n6758 137.715
R7937 gnd.n6759 gnd.n595 137.715
R7938 gnd.n6767 gnd.n595 137.715
R7939 gnd.n6768 gnd.n6767 137.715
R7940 gnd.n6769 gnd.n6768 137.715
R7941 gnd.n6769 gnd.n589 137.715
R7942 gnd.n6777 gnd.n589 137.715
R7943 gnd.n6778 gnd.n6777 137.715
R7944 gnd.n6779 gnd.n6778 137.715
R7945 gnd.n6779 gnd.n583 137.715
R7946 gnd.n6787 gnd.n583 137.715
R7947 gnd.n6788 gnd.n6787 137.715
R7948 gnd.n6789 gnd.n6788 137.715
R7949 gnd.n6789 gnd.n577 137.715
R7950 gnd.n6797 gnd.n577 137.715
R7951 gnd.n6798 gnd.n6797 137.715
R7952 gnd.n6799 gnd.n6798 137.715
R7953 gnd.n6799 gnd.n571 137.715
R7954 gnd.n6807 gnd.n571 137.715
R7955 gnd.n6808 gnd.n6807 137.715
R7956 gnd.n6809 gnd.n6808 137.715
R7957 gnd.n6809 gnd.n565 137.715
R7958 gnd.n6819 gnd.n565 137.715
R7959 gnd.n6820 gnd.n6819 137.715
R7960 gnd.n6821 gnd.n6820 137.715
R7961 gnd.n1968 gnd.t21 130.484
R7962 gnd.n1977 gnd.t28 126.766
R7963 gnd.n1975 gnd.t113 126.766
R7964 gnd.n1961 gnd.t122 126.766
R7965 gnd.n1969 gnd.t84 126.766
R7966 gnd.n5241 gnd.t46 126.766
R7967 gnd.n5243 gnd.t94 126.766
R7968 gnd.n5252 gnd.t67 126.766
R7969 gnd.n5254 gnd.t97 126.766
R7970 gnd.n6938 gnd.n440 105.281
R7971 gnd.n2098 gnd.n1302 105.281
R7972 gnd.n3787 gnd.n3786 104.615
R7973 gnd.n3786 gnd.n3764 104.615
R7974 gnd.n3779 gnd.n3764 104.615
R7975 gnd.n3779 gnd.n3778 104.615
R7976 gnd.n3778 gnd.n3768 104.615
R7977 gnd.n3771 gnd.n3768 104.615
R7978 gnd.n3755 gnd.n3754 104.615
R7979 gnd.n3754 gnd.n3732 104.615
R7980 gnd.n3747 gnd.n3732 104.615
R7981 gnd.n3747 gnd.n3746 104.615
R7982 gnd.n3746 gnd.n3736 104.615
R7983 gnd.n3739 gnd.n3736 104.615
R7984 gnd.n3723 gnd.n3722 104.615
R7985 gnd.n3722 gnd.n3700 104.615
R7986 gnd.n3715 gnd.n3700 104.615
R7987 gnd.n3715 gnd.n3714 104.615
R7988 gnd.n3714 gnd.n3704 104.615
R7989 gnd.n3707 gnd.n3704 104.615
R7990 gnd.n3692 gnd.n3691 104.615
R7991 gnd.n3691 gnd.n3669 104.615
R7992 gnd.n3684 gnd.n3669 104.615
R7993 gnd.n3684 gnd.n3683 104.615
R7994 gnd.n3683 gnd.n3673 104.615
R7995 gnd.n3676 gnd.n3673 104.615
R7996 gnd.n3660 gnd.n3659 104.615
R7997 gnd.n3659 gnd.n3637 104.615
R7998 gnd.n3652 gnd.n3637 104.615
R7999 gnd.n3652 gnd.n3651 104.615
R8000 gnd.n3651 gnd.n3641 104.615
R8001 gnd.n3644 gnd.n3641 104.615
R8002 gnd.n3628 gnd.n3627 104.615
R8003 gnd.n3627 gnd.n3605 104.615
R8004 gnd.n3620 gnd.n3605 104.615
R8005 gnd.n3620 gnd.n3619 104.615
R8006 gnd.n3619 gnd.n3609 104.615
R8007 gnd.n3612 gnd.n3609 104.615
R8008 gnd.n3596 gnd.n3595 104.615
R8009 gnd.n3595 gnd.n3573 104.615
R8010 gnd.n3588 gnd.n3573 104.615
R8011 gnd.n3588 gnd.n3587 104.615
R8012 gnd.n3587 gnd.n3577 104.615
R8013 gnd.n3580 gnd.n3577 104.615
R8014 gnd.n3565 gnd.n3564 104.615
R8015 gnd.n3564 gnd.n3542 104.615
R8016 gnd.n3557 gnd.n3542 104.615
R8017 gnd.n3557 gnd.n3556 104.615
R8018 gnd.n3556 gnd.n3546 104.615
R8019 gnd.n3549 gnd.n3546 104.615
R8020 gnd.n2939 gnd.t41 100.632
R8021 gnd.n2496 gnd.t82 100.632
R8022 gnd.n7319 gnd.n112 99.6594
R8023 gnd.n7317 gnd.n7316 99.6594
R8024 gnd.n7312 gnd.n119 99.6594
R8025 gnd.n7310 gnd.n7309 99.6594
R8026 gnd.n7305 gnd.n126 99.6594
R8027 gnd.n7303 gnd.n7302 99.6594
R8028 gnd.n7298 gnd.n133 99.6594
R8029 gnd.n7296 gnd.n7295 99.6594
R8030 gnd.n7288 gnd.n140 99.6594
R8031 gnd.n7286 gnd.n7285 99.6594
R8032 gnd.n7281 gnd.n147 99.6594
R8033 gnd.n7279 gnd.n7278 99.6594
R8034 gnd.n7274 gnd.n154 99.6594
R8035 gnd.n7272 gnd.n7271 99.6594
R8036 gnd.n7267 gnd.n161 99.6594
R8037 gnd.n7265 gnd.n7264 99.6594
R8038 gnd.n7260 gnd.n168 99.6594
R8039 gnd.n7258 gnd.n7257 99.6594
R8040 gnd.n173 gnd.n172 99.6594
R8041 gnd.n6968 gnd.n6967 99.6594
R8042 gnd.n425 gnd.n396 99.6594
R8043 gnd.n6960 gnd.n397 99.6594
R8044 gnd.n6956 gnd.n398 99.6594
R8045 gnd.n6952 gnd.n399 99.6594
R8046 gnd.n6948 gnd.n400 99.6594
R8047 gnd.n6944 gnd.n401 99.6594
R8048 gnd.n6940 gnd.n402 99.6594
R8049 gnd.n6935 gnd.n404 99.6594
R8050 gnd.n6931 gnd.n405 99.6594
R8051 gnd.n6927 gnd.n406 99.6594
R8052 gnd.n6923 gnd.n407 99.6594
R8053 gnd.n6919 gnd.n408 99.6594
R8054 gnd.n6915 gnd.n409 99.6594
R8055 gnd.n6911 gnd.n410 99.6594
R8056 gnd.n6907 gnd.n411 99.6594
R8057 gnd.n6903 gnd.n412 99.6594
R8058 gnd.n464 gnd.n413 99.6594
R8059 gnd.n5925 gnd.n5924 99.6594
R8060 gnd.n5922 gnd.n5921 99.6594
R8061 gnd.n5917 gnd.n1285 99.6594
R8062 gnd.n5915 gnd.n5914 99.6594
R8063 gnd.n5910 gnd.n1292 99.6594
R8064 gnd.n5908 gnd.n5907 99.6594
R8065 gnd.n5903 gnd.n1299 99.6594
R8066 gnd.n5899 gnd.n5898 99.6594
R8067 gnd.n5894 gnd.n1310 99.6594
R8068 gnd.n5892 gnd.n5891 99.6594
R8069 gnd.n5887 gnd.n1317 99.6594
R8070 gnd.n5885 gnd.n5884 99.6594
R8071 gnd.n5880 gnd.n1324 99.6594
R8072 gnd.n5878 gnd.n5877 99.6594
R8073 gnd.n5873 gnd.n1331 99.6594
R8074 gnd.n5871 gnd.n5870 99.6594
R8075 gnd.n5866 gnd.n1340 99.6594
R8076 gnd.n5864 gnd.n5863 99.6594
R8077 gnd.n3968 gnd.n2456 99.6594
R8078 gnd.n3976 gnd.n3975 99.6594
R8079 gnd.n3979 gnd.n3978 99.6594
R8080 gnd.n3986 gnd.n3985 99.6594
R8081 gnd.n3989 gnd.n3988 99.6594
R8082 gnd.n3996 gnd.n3995 99.6594
R8083 gnd.n3999 gnd.n3998 99.6594
R8084 gnd.n4006 gnd.n4005 99.6594
R8085 gnd.n4009 gnd.n4008 99.6594
R8086 gnd.n4016 gnd.n4015 99.6594
R8087 gnd.n4019 gnd.n4018 99.6594
R8088 gnd.n4026 gnd.n4025 99.6594
R8089 gnd.n4029 gnd.n4028 99.6594
R8090 gnd.n4036 gnd.n4035 99.6594
R8091 gnd.n4039 gnd.n4038 99.6594
R8092 gnd.n4046 gnd.n4045 99.6594
R8093 gnd.n4049 gnd.n4048 99.6594
R8094 gnd.n4057 gnd.n4056 99.6594
R8095 gnd.n4060 gnd.n4059 99.6594
R8096 gnd.n3910 gnd.n2479 99.6594
R8097 gnd.n3908 gnd.n2478 99.6594
R8098 gnd.n3904 gnd.n2477 99.6594
R8099 gnd.n3900 gnd.n2476 99.6594
R8100 gnd.n3896 gnd.n2475 99.6594
R8101 gnd.n3892 gnd.n2474 99.6594
R8102 gnd.n3888 gnd.n2473 99.6594
R8103 gnd.n3820 gnd.n2472 99.6594
R8104 gnd.n3151 gnd.n2882 99.6594
R8105 gnd.n2908 gnd.n2889 99.6594
R8106 gnd.n2910 gnd.n2890 99.6594
R8107 gnd.n2918 gnd.n2891 99.6594
R8108 gnd.n2920 gnd.n2892 99.6594
R8109 gnd.n2928 gnd.n2893 99.6594
R8110 gnd.n2930 gnd.n2894 99.6594
R8111 gnd.n2938 gnd.n2895 99.6594
R8112 gnd.n3878 gnd.n2459 99.6594
R8113 gnd.n3874 gnd.n2460 99.6594
R8114 gnd.n3870 gnd.n2461 99.6594
R8115 gnd.n3866 gnd.n2462 99.6594
R8116 gnd.n3862 gnd.n2463 99.6594
R8117 gnd.n3858 gnd.n2464 99.6594
R8118 gnd.n3854 gnd.n2465 99.6594
R8119 gnd.n3850 gnd.n2466 99.6594
R8120 gnd.n3846 gnd.n2467 99.6594
R8121 gnd.n3842 gnd.n2468 99.6594
R8122 gnd.n3838 gnd.n2469 99.6594
R8123 gnd.n3834 gnd.n2470 99.6594
R8124 gnd.n3830 gnd.n2471 99.6594
R8125 gnd.n3066 gnd.n3065 99.6594
R8126 gnd.n3060 gnd.n2977 99.6594
R8127 gnd.n3057 gnd.n2978 99.6594
R8128 gnd.n3053 gnd.n2979 99.6594
R8129 gnd.n3049 gnd.n2980 99.6594
R8130 gnd.n3045 gnd.n2981 99.6594
R8131 gnd.n3041 gnd.n2982 99.6594
R8132 gnd.n3037 gnd.n2983 99.6594
R8133 gnd.n3033 gnd.n2984 99.6594
R8134 gnd.n3029 gnd.n2985 99.6594
R8135 gnd.n3025 gnd.n2986 99.6594
R8136 gnd.n3021 gnd.n2987 99.6594
R8137 gnd.n3068 gnd.n2976 99.6594
R8138 gnd.n7181 gnd.n7180 99.6594
R8139 gnd.n7186 gnd.n7185 99.6594
R8140 gnd.n7189 gnd.n7188 99.6594
R8141 gnd.n7194 gnd.n7193 99.6594
R8142 gnd.n7197 gnd.n7196 99.6594
R8143 gnd.n7202 gnd.n7201 99.6594
R8144 gnd.n7205 gnd.n7204 99.6594
R8145 gnd.n7210 gnd.n7209 99.6594
R8146 gnd.n7213 gnd.n99 99.6594
R8147 gnd.n5701 gnd.n414 99.6594
R8148 gnd.n1479 gnd.n415 99.6594
R8149 gnd.n1489 gnd.n416 99.6594
R8150 gnd.n1491 gnd.n417 99.6594
R8151 gnd.n1499 gnd.n418 99.6594
R8152 gnd.n1507 gnd.n419 99.6594
R8153 gnd.n1509 gnd.n420 99.6594
R8154 gnd.n1517 gnd.n421 99.6594
R8155 gnd.n1525 gnd.n422 99.6594
R8156 gnd.n2204 gnd.n2203 99.6594
R8157 gnd.n2215 gnd.n2214 99.6594
R8158 gnd.n2224 gnd.n2223 99.6594
R8159 gnd.n2227 gnd.n2226 99.6594
R8160 gnd.n2236 gnd.n2235 99.6594
R8161 gnd.n2245 gnd.n2244 99.6594
R8162 gnd.n2248 gnd.n2247 99.6594
R8163 gnd.n2257 gnd.n2256 99.6594
R8164 gnd.n4564 gnd.n4563 99.6594
R8165 gnd.n4206 gnd.n4097 99.6594
R8166 gnd.n4205 gnd.n4204 99.6594
R8167 gnd.n4198 gnd.n4100 99.6594
R8168 gnd.n4197 gnd.n4196 99.6594
R8169 gnd.n4190 gnd.n4106 99.6594
R8170 gnd.n4189 gnd.n4188 99.6594
R8171 gnd.n4182 gnd.n4112 99.6594
R8172 gnd.n4181 gnd.n4180 99.6594
R8173 gnd.n4170 gnd.n4118 99.6594
R8174 gnd.n4207 gnd.n4206 99.6594
R8175 gnd.n4204 gnd.n4203 99.6594
R8176 gnd.n4199 gnd.n4198 99.6594
R8177 gnd.n4196 gnd.n4195 99.6594
R8178 gnd.n4191 gnd.n4190 99.6594
R8179 gnd.n4188 gnd.n4187 99.6594
R8180 gnd.n4183 gnd.n4182 99.6594
R8181 gnd.n4180 gnd.n4179 99.6594
R8182 gnd.n4171 gnd.n4170 99.6594
R8183 gnd.n4563 gnd.n2261 99.6594
R8184 gnd.n2256 gnd.n2255 99.6594
R8185 gnd.n2247 gnd.n2246 99.6594
R8186 gnd.n2244 gnd.n2237 99.6594
R8187 gnd.n2235 gnd.n2234 99.6594
R8188 gnd.n2226 gnd.n2225 99.6594
R8189 gnd.n2223 gnd.n2216 99.6594
R8190 gnd.n2214 gnd.n2213 99.6594
R8191 gnd.n2203 gnd.n2202 99.6594
R8192 gnd.n1478 gnd.n414 99.6594
R8193 gnd.n1488 gnd.n415 99.6594
R8194 gnd.n1490 gnd.n416 99.6594
R8195 gnd.n1498 gnd.n417 99.6594
R8196 gnd.n1506 gnd.n418 99.6594
R8197 gnd.n1508 gnd.n419 99.6594
R8198 gnd.n1516 gnd.n420 99.6594
R8199 gnd.n1524 gnd.n421 99.6594
R8200 gnd.n5656 gnd.n422 99.6594
R8201 gnd.n7214 gnd.n7213 99.6594
R8202 gnd.n7209 gnd.n7208 99.6594
R8203 gnd.n7204 gnd.n7203 99.6594
R8204 gnd.n7201 gnd.n7200 99.6594
R8205 gnd.n7196 gnd.n7195 99.6594
R8206 gnd.n7193 gnd.n7192 99.6594
R8207 gnd.n7188 gnd.n7187 99.6594
R8208 gnd.n7185 gnd.n7184 99.6594
R8209 gnd.n7180 gnd.n7179 99.6594
R8210 gnd.n3066 gnd.n2989 99.6594
R8211 gnd.n3058 gnd.n2977 99.6594
R8212 gnd.n3054 gnd.n2978 99.6594
R8213 gnd.n3050 gnd.n2979 99.6594
R8214 gnd.n3046 gnd.n2980 99.6594
R8215 gnd.n3042 gnd.n2981 99.6594
R8216 gnd.n3038 gnd.n2982 99.6594
R8217 gnd.n3034 gnd.n2983 99.6594
R8218 gnd.n3030 gnd.n2984 99.6594
R8219 gnd.n3026 gnd.n2985 99.6594
R8220 gnd.n3022 gnd.n2986 99.6594
R8221 gnd.n3018 gnd.n2987 99.6594
R8222 gnd.n3069 gnd.n3068 99.6594
R8223 gnd.n3833 gnd.n2471 99.6594
R8224 gnd.n3837 gnd.n2470 99.6594
R8225 gnd.n3841 gnd.n2469 99.6594
R8226 gnd.n3845 gnd.n2468 99.6594
R8227 gnd.n3849 gnd.n2467 99.6594
R8228 gnd.n3853 gnd.n2466 99.6594
R8229 gnd.n3857 gnd.n2465 99.6594
R8230 gnd.n3861 gnd.n2464 99.6594
R8231 gnd.n3865 gnd.n2463 99.6594
R8232 gnd.n3869 gnd.n2462 99.6594
R8233 gnd.n3873 gnd.n2461 99.6594
R8234 gnd.n3877 gnd.n2460 99.6594
R8235 gnd.n2500 gnd.n2459 99.6594
R8236 gnd.n3152 gnd.n3151 99.6594
R8237 gnd.n2911 gnd.n2889 99.6594
R8238 gnd.n2917 gnd.n2890 99.6594
R8239 gnd.n2921 gnd.n2891 99.6594
R8240 gnd.n2927 gnd.n2892 99.6594
R8241 gnd.n2931 gnd.n2893 99.6594
R8242 gnd.n2937 gnd.n2894 99.6594
R8243 gnd.n2895 gnd.n2879 99.6594
R8244 gnd.n3887 gnd.n2472 99.6594
R8245 gnd.n3891 gnd.n2473 99.6594
R8246 gnd.n3895 gnd.n2474 99.6594
R8247 gnd.n3899 gnd.n2475 99.6594
R8248 gnd.n3903 gnd.n2476 99.6594
R8249 gnd.n3907 gnd.n2477 99.6594
R8250 gnd.n3911 gnd.n2478 99.6594
R8251 gnd.n2481 gnd.n2479 99.6594
R8252 gnd.n3969 gnd.n3968 99.6594
R8253 gnd.n3977 gnd.n3976 99.6594
R8254 gnd.n3978 gnd.n3961 99.6594
R8255 gnd.n3987 gnd.n3986 99.6594
R8256 gnd.n3988 gnd.n3957 99.6594
R8257 gnd.n3997 gnd.n3996 99.6594
R8258 gnd.n3998 gnd.n3953 99.6594
R8259 gnd.n4007 gnd.n4006 99.6594
R8260 gnd.n4008 gnd.n3946 99.6594
R8261 gnd.n4017 gnd.n4016 99.6594
R8262 gnd.n4018 gnd.n3942 99.6594
R8263 gnd.n4027 gnd.n4026 99.6594
R8264 gnd.n4028 gnd.n3938 99.6594
R8265 gnd.n4037 gnd.n4036 99.6594
R8266 gnd.n4038 gnd.n3934 99.6594
R8267 gnd.n4047 gnd.n4046 99.6594
R8268 gnd.n4048 gnd.n3930 99.6594
R8269 gnd.n4058 gnd.n4057 99.6594
R8270 gnd.n4061 gnd.n4060 99.6594
R8271 gnd.n5865 gnd.n5864 99.6594
R8272 gnd.n1340 gnd.n1332 99.6594
R8273 gnd.n5872 gnd.n5871 99.6594
R8274 gnd.n1331 gnd.n1325 99.6594
R8275 gnd.n5879 gnd.n5878 99.6594
R8276 gnd.n1324 gnd.n1318 99.6594
R8277 gnd.n5886 gnd.n5885 99.6594
R8278 gnd.n1317 gnd.n1311 99.6594
R8279 gnd.n5893 gnd.n5892 99.6594
R8280 gnd.n1310 gnd.n1303 99.6594
R8281 gnd.n5902 gnd.n5901 99.6594
R8282 gnd.n1299 gnd.n1293 99.6594
R8283 gnd.n5909 gnd.n5908 99.6594
R8284 gnd.n1292 gnd.n1286 99.6594
R8285 gnd.n5916 gnd.n5915 99.6594
R8286 gnd.n1285 gnd.n1278 99.6594
R8287 gnd.n5923 gnd.n5922 99.6594
R8288 gnd.n5926 gnd.n5925 99.6594
R8289 gnd.n6967 gnd.n394 99.6594
R8290 gnd.n6961 gnd.n396 99.6594
R8291 gnd.n6957 gnd.n397 99.6594
R8292 gnd.n6953 gnd.n398 99.6594
R8293 gnd.n6949 gnd.n399 99.6594
R8294 gnd.n6945 gnd.n400 99.6594
R8295 gnd.n6941 gnd.n401 99.6594
R8296 gnd.n6936 gnd.n403 99.6594
R8297 gnd.n6932 gnd.n404 99.6594
R8298 gnd.n6928 gnd.n405 99.6594
R8299 gnd.n6924 gnd.n406 99.6594
R8300 gnd.n6920 gnd.n407 99.6594
R8301 gnd.n6916 gnd.n408 99.6594
R8302 gnd.n6912 gnd.n409 99.6594
R8303 gnd.n6908 gnd.n410 99.6594
R8304 gnd.n6904 gnd.n411 99.6594
R8305 gnd.n463 gnd.n412 99.6594
R8306 gnd.n6896 gnd.n413 99.6594
R8307 gnd.n172 gnd.n169 99.6594
R8308 gnd.n7259 gnd.n7258 99.6594
R8309 gnd.n168 gnd.n162 99.6594
R8310 gnd.n7266 gnd.n7265 99.6594
R8311 gnd.n161 gnd.n155 99.6594
R8312 gnd.n7273 gnd.n7272 99.6594
R8313 gnd.n154 gnd.n148 99.6594
R8314 gnd.n7280 gnd.n7279 99.6594
R8315 gnd.n147 gnd.n141 99.6594
R8316 gnd.n7287 gnd.n7286 99.6594
R8317 gnd.n140 gnd.n134 99.6594
R8318 gnd.n7297 gnd.n7296 99.6594
R8319 gnd.n133 gnd.n127 99.6594
R8320 gnd.n7304 gnd.n7303 99.6594
R8321 gnd.n126 gnd.n120 99.6594
R8322 gnd.n7311 gnd.n7310 99.6594
R8323 gnd.n119 gnd.n113 99.6594
R8324 gnd.n7318 gnd.n7317 99.6594
R8325 gnd.n112 gnd.n109 99.6594
R8326 gnd.n4556 gnd.n4555 99.6594
R8327 gnd.n2266 gnd.n2265 99.6594
R8328 gnd.n2268 gnd.n2220 99.6594
R8329 gnd.n2269 gnd.n2230 99.6594
R8330 gnd.n2271 gnd.n2270 99.6594
R8331 gnd.n2273 gnd.n2241 99.6594
R8332 gnd.n2274 gnd.n2251 99.6594
R8333 gnd.n4558 gnd.n2263 99.6594
R8334 gnd.n2275 gnd.n2262 99.6594
R8335 gnd.n2276 gnd.n1351 99.6594
R8336 gnd.n2278 gnd.n2277 99.6594
R8337 gnd.n2279 gnd.n1356 99.6594
R8338 gnd.n2280 gnd.n1362 99.6594
R8339 gnd.n2282 gnd.n1364 99.6594
R8340 gnd.n4556 gnd.n2209 99.6594
R8341 gnd.n2266 gnd.n2219 99.6594
R8342 gnd.n2268 gnd.n2267 99.6594
R8343 gnd.n2269 gnd.n2231 99.6594
R8344 gnd.n2271 gnd.n2240 99.6594
R8345 gnd.n2273 gnd.n2272 99.6594
R8346 gnd.n2274 gnd.n2252 99.6594
R8347 gnd.n4559 gnd.n4558 99.6594
R8348 gnd.n2275 gnd.n1350 99.6594
R8349 gnd.n2276 gnd.n1352 99.6594
R8350 gnd.n2278 gnd.n1355 99.6594
R8351 gnd.n2279 gnd.n1357 99.6594
R8352 gnd.n2280 gnd.n1363 99.6594
R8353 gnd.n2282 gnd.n2281 99.6594
R8354 gnd.n1545 gnd.n1484 99.6594
R8355 gnd.n1547 gnd.n1546 99.6594
R8356 gnd.n1548 gnd.n1495 99.6594
R8357 gnd.n1550 gnd.n1502 99.6594
R8358 gnd.n1552 gnd.n1551 99.6594
R8359 gnd.n1553 gnd.n1513 99.6594
R8360 gnd.n1555 gnd.n1520 99.6594
R8361 gnd.n1557 gnd.n1556 99.6594
R8362 gnd.n1558 gnd.n1529 99.6594
R8363 gnd.n1559 gnd.n1531 99.6594
R8364 gnd.n1561 gnd.n1534 99.6594
R8365 gnd.n1562 gnd.n1536 99.6594
R8366 gnd.n1564 gnd.n1542 99.6594
R8367 gnd.n5632 gnd.n5631 99.6594
R8368 gnd.n5631 gnd.n1543 99.6594
R8369 gnd.n1564 gnd.n1563 99.6594
R8370 gnd.n1562 gnd.n1535 99.6594
R8371 gnd.n1561 gnd.n1560 99.6594
R8372 gnd.n1559 gnd.n1530 99.6594
R8373 gnd.n1558 gnd.n1528 99.6594
R8374 gnd.n1557 gnd.n1521 99.6594
R8375 gnd.n1555 gnd.n1554 99.6594
R8376 gnd.n1553 gnd.n1512 99.6594
R8377 gnd.n1552 gnd.n1503 99.6594
R8378 gnd.n1550 gnd.n1549 99.6594
R8379 gnd.n1548 gnd.n1494 99.6594
R8380 gnd.n1547 gnd.n1485 99.6594
R8381 gnd.n1545 gnd.n1474 99.6594
R8382 gnd.n1358 gnd.t93 98.63
R8383 gnd.n7211 gnd.t19 98.63
R8384 gnd.n5657 gnd.t58 98.63
R8385 gnd.n2258 gnd.t88 98.63
R8386 gnd.n443 gnd.t55 98.63
R8387 gnd.n465 gnd.t34 98.63
R8388 gnd.n175 gnd.t120 98.63
R8389 gnd.n7290 gnd.t36 98.63
R8390 gnd.n3950 gnd.t118 98.63
R8391 gnd.n3926 gnd.t109 98.63
R8392 gnd.n1337 gnd.t51 98.63
R8393 gnd.n1300 gnd.t71 98.63
R8394 gnd.n4121 gnd.t66 98.63
R8395 gnd.n1539 gnd.t75 98.63
R8396 gnd.n2028 gnd.t112 92.8196
R8397 gnd.n1645 gnd.t26 92.8196
R8398 gnd.n2025 gnd.t45 92.8118
R8399 gnd.n5256 gnd.t105 92.8118
R8400 gnd.n6821 gnd.n100 82.6296
R8401 gnd.n1968 gnd.n1967 81.8399
R8402 gnd.n2940 gnd.t40 74.8376
R8403 gnd.n2497 gnd.t83 74.8376
R8404 gnd.n2029 gnd.t111 72.8438
R8405 gnd.n1646 gnd.t27 72.8438
R8406 gnd.n1969 gnd.n1962 72.8411
R8407 gnd.n1975 gnd.n1960 72.8411
R8408 gnd.n5252 gnd.n5251 72.8411
R8409 gnd.n1359 gnd.t92 72.836
R8410 gnd.n2026 gnd.t44 72.836
R8411 gnd.n5257 gnd.t106 72.836
R8412 gnd.n7212 gnd.t20 72.836
R8413 gnd.n5658 gnd.t57 72.836
R8414 gnd.n2259 gnd.t89 72.836
R8415 gnd.n444 gnd.t54 72.836
R8416 gnd.n466 gnd.t33 72.836
R8417 gnd.n176 gnd.t121 72.836
R8418 gnd.n7291 gnd.t37 72.836
R8419 gnd.n3951 gnd.t117 72.836
R8420 gnd.n3927 gnd.t108 72.836
R8421 gnd.n1338 gnd.t52 72.836
R8422 gnd.n1301 gnd.t72 72.836
R8423 gnd.n4122 gnd.t65 72.836
R8424 gnd.n1540 gnd.t76 72.836
R8425 gnd.n5320 gnd.n1608 71.676
R8426 gnd.n5316 gnd.n1609 71.676
R8427 gnd.n5312 gnd.n1610 71.676
R8428 gnd.n5308 gnd.n1611 71.676
R8429 gnd.n5304 gnd.n1612 71.676
R8430 gnd.n5300 gnd.n1613 71.676
R8431 gnd.n5296 gnd.n1614 71.676
R8432 gnd.n5292 gnd.n1615 71.676
R8433 gnd.n5288 gnd.n1616 71.676
R8434 gnd.n5284 gnd.n1617 71.676
R8435 gnd.n5280 gnd.n1618 71.676
R8436 gnd.n5276 gnd.n1619 71.676
R8437 gnd.n5272 gnd.n1620 71.676
R8438 gnd.n5268 gnd.n1621 71.676
R8439 gnd.n5263 gnd.n1622 71.676
R8440 gnd.n5259 gnd.n1623 71.676
R8441 gnd.n5393 gnd.n1644 71.676
R8442 gnd.n5389 gnd.n1643 71.676
R8443 gnd.n5384 gnd.n1642 71.676
R8444 gnd.n5380 gnd.n1641 71.676
R8445 gnd.n5376 gnd.n1640 71.676
R8446 gnd.n5372 gnd.n1639 71.676
R8447 gnd.n5368 gnd.n1638 71.676
R8448 gnd.n5364 gnd.n1637 71.676
R8449 gnd.n5360 gnd.n1636 71.676
R8450 gnd.n5356 gnd.n1635 71.676
R8451 gnd.n5352 gnd.n1634 71.676
R8452 gnd.n5348 gnd.n1633 71.676
R8453 gnd.n5344 gnd.n1632 71.676
R8454 gnd.n5340 gnd.n1631 71.676
R8455 gnd.n5336 gnd.n1630 71.676
R8456 gnd.n5332 gnd.n1629 71.676
R8457 gnd.n5328 gnd.n1628 71.676
R8458 gnd.n2160 gnd.n1980 71.676
R8459 gnd.n2155 gnd.n1991 71.676
R8460 gnd.n2152 gnd.n1992 71.676
R8461 gnd.n2148 gnd.n1993 71.676
R8462 gnd.n2144 gnd.n1994 71.676
R8463 gnd.n2140 gnd.n1995 71.676
R8464 gnd.n2136 gnd.n1996 71.676
R8465 gnd.n2132 gnd.n1997 71.676
R8466 gnd.n2128 gnd.n1998 71.676
R8467 gnd.n2124 gnd.n1999 71.676
R8468 gnd.n2120 gnd.n2000 71.676
R8469 gnd.n2116 gnd.n2001 71.676
R8470 gnd.n2112 gnd.n2002 71.676
R8471 gnd.n2108 gnd.n2003 71.676
R8472 gnd.n2104 gnd.n2004 71.676
R8473 gnd.n2100 gnd.n2005 71.676
R8474 gnd.n2096 gnd.n2007 71.676
R8475 gnd.n2091 gnd.n2008 71.676
R8476 gnd.n2086 gnd.n2009 71.676
R8477 gnd.n2082 gnd.n2010 71.676
R8478 gnd.n2078 gnd.n2011 71.676
R8479 gnd.n2074 gnd.n2012 71.676
R8480 gnd.n2070 gnd.n2013 71.676
R8481 gnd.n2066 gnd.n2014 71.676
R8482 gnd.n2062 gnd.n2015 71.676
R8483 gnd.n2058 gnd.n2016 71.676
R8484 gnd.n2054 gnd.n2017 71.676
R8485 gnd.n2050 gnd.n2018 71.676
R8486 gnd.n2046 gnd.n2019 71.676
R8487 gnd.n2042 gnd.n2020 71.676
R8488 gnd.n2038 gnd.n2021 71.676
R8489 gnd.n2034 gnd.n2022 71.676
R8490 gnd.n2160 gnd.n2159 71.676
R8491 gnd.n2153 gnd.n1991 71.676
R8492 gnd.n2149 gnd.n1992 71.676
R8493 gnd.n2145 gnd.n1993 71.676
R8494 gnd.n2141 gnd.n1994 71.676
R8495 gnd.n2137 gnd.n1995 71.676
R8496 gnd.n2133 gnd.n1996 71.676
R8497 gnd.n2129 gnd.n1997 71.676
R8498 gnd.n2125 gnd.n1998 71.676
R8499 gnd.n2121 gnd.n1999 71.676
R8500 gnd.n2117 gnd.n2000 71.676
R8501 gnd.n2113 gnd.n2001 71.676
R8502 gnd.n2109 gnd.n2002 71.676
R8503 gnd.n2105 gnd.n2003 71.676
R8504 gnd.n2101 gnd.n2004 71.676
R8505 gnd.n2097 gnd.n2006 71.676
R8506 gnd.n2092 gnd.n2007 71.676
R8507 gnd.n2087 gnd.n2008 71.676
R8508 gnd.n2083 gnd.n2009 71.676
R8509 gnd.n2079 gnd.n2010 71.676
R8510 gnd.n2075 gnd.n2011 71.676
R8511 gnd.n2071 gnd.n2012 71.676
R8512 gnd.n2067 gnd.n2013 71.676
R8513 gnd.n2063 gnd.n2014 71.676
R8514 gnd.n2059 gnd.n2015 71.676
R8515 gnd.n2055 gnd.n2016 71.676
R8516 gnd.n2051 gnd.n2017 71.676
R8517 gnd.n2047 gnd.n2018 71.676
R8518 gnd.n2043 gnd.n2019 71.676
R8519 gnd.n2039 gnd.n2020 71.676
R8520 gnd.n2035 gnd.n2021 71.676
R8521 gnd.n2031 gnd.n2022 71.676
R8522 gnd.n5331 gnd.n1628 71.676
R8523 gnd.n5335 gnd.n1629 71.676
R8524 gnd.n5339 gnd.n1630 71.676
R8525 gnd.n5343 gnd.n1631 71.676
R8526 gnd.n5347 gnd.n1632 71.676
R8527 gnd.n5351 gnd.n1633 71.676
R8528 gnd.n5355 gnd.n1634 71.676
R8529 gnd.n5359 gnd.n1635 71.676
R8530 gnd.n5363 gnd.n1636 71.676
R8531 gnd.n5367 gnd.n1637 71.676
R8532 gnd.n5371 gnd.n1638 71.676
R8533 gnd.n5375 gnd.n1639 71.676
R8534 gnd.n5379 gnd.n1640 71.676
R8535 gnd.n5383 gnd.n1641 71.676
R8536 gnd.n5388 gnd.n1642 71.676
R8537 gnd.n5392 gnd.n1643 71.676
R8538 gnd.n5258 gnd.n1624 71.676
R8539 gnd.n5262 gnd.n1623 71.676
R8540 gnd.n5267 gnd.n1622 71.676
R8541 gnd.n5271 gnd.n1621 71.676
R8542 gnd.n5275 gnd.n1620 71.676
R8543 gnd.n5279 gnd.n1619 71.676
R8544 gnd.n5283 gnd.n1618 71.676
R8545 gnd.n5287 gnd.n1617 71.676
R8546 gnd.n5291 gnd.n1616 71.676
R8547 gnd.n5295 gnd.n1615 71.676
R8548 gnd.n5299 gnd.n1614 71.676
R8549 gnd.n5303 gnd.n1613 71.676
R8550 gnd.n5307 gnd.n1612 71.676
R8551 gnd.n5311 gnd.n1611 71.676
R8552 gnd.n5315 gnd.n1610 71.676
R8553 gnd.n5319 gnd.n1609 71.676
R8554 gnd.n1651 gnd.n1608 71.676
R8555 gnd.n8 gnd.t177 69.1507
R8556 gnd.n14 gnd.t179 68.4792
R8557 gnd.n13 gnd.t309 68.4792
R8558 gnd.n12 gnd.t12 68.4792
R8559 gnd.n11 gnd.t142 68.4792
R8560 gnd.n10 gnd.t319 68.4792
R8561 gnd.n9 gnd.t168 68.4792
R8562 gnd.n8 gnd.t315 68.4792
R8563 gnd.n3067 gnd.n2971 64.369
R8564 gnd.n2089 gnd.n2029 59.5399
R8565 gnd.n5386 gnd.n1646 59.5399
R8566 gnd.n2027 gnd.n2026 59.5399
R8567 gnd.n5265 gnd.n5257 59.5399
R8568 gnd.n1979 gnd.n1978 59.1804
R8569 gnd.n3919 gnd.n2457 57.3586
R8570 gnd.n4214 gnd.n3920 57.3586
R8571 gnd.n7327 gnd.n102 57.3586
R8572 gnd.n2722 gnd.t187 56.607
R8573 gnd.n48 gnd.t284 56.607
R8574 gnd.n2691 gnd.t246 56.407
R8575 gnd.n2706 gnd.t225 56.407
R8576 gnd.n17 gnd.t280 56.407
R8577 gnd.n32 gnd.t256 56.407
R8578 gnd.n2735 gnd.t296 55.8337
R8579 gnd.n2704 gnd.t254 55.8337
R8580 gnd.n2719 gnd.t235 55.8337
R8581 gnd.n61 gnd.t263 55.8337
R8582 gnd.n30 gnd.t286 55.8337
R8583 gnd.n45 gnd.t264 55.8337
R8584 gnd.n1966 gnd.n1965 54.358
R8585 gnd.n5249 gnd.n5248 54.358
R8586 gnd.n2722 gnd.n2721 53.0052
R8587 gnd.n2724 gnd.n2723 53.0052
R8588 gnd.n2726 gnd.n2725 53.0052
R8589 gnd.n2728 gnd.n2727 53.0052
R8590 gnd.n2730 gnd.n2729 53.0052
R8591 gnd.n2732 gnd.n2731 53.0052
R8592 gnd.n2734 gnd.n2733 53.0052
R8593 gnd.n2691 gnd.n2690 53.0052
R8594 gnd.n2693 gnd.n2692 53.0052
R8595 gnd.n2695 gnd.n2694 53.0052
R8596 gnd.n2697 gnd.n2696 53.0052
R8597 gnd.n2699 gnd.n2698 53.0052
R8598 gnd.n2701 gnd.n2700 53.0052
R8599 gnd.n2703 gnd.n2702 53.0052
R8600 gnd.n2706 gnd.n2705 53.0052
R8601 gnd.n2708 gnd.n2707 53.0052
R8602 gnd.n2710 gnd.n2709 53.0052
R8603 gnd.n2712 gnd.n2711 53.0052
R8604 gnd.n2714 gnd.n2713 53.0052
R8605 gnd.n2716 gnd.n2715 53.0052
R8606 gnd.n2718 gnd.n2717 53.0052
R8607 gnd.n60 gnd.n59 53.0052
R8608 gnd.n58 gnd.n57 53.0052
R8609 gnd.n56 gnd.n55 53.0052
R8610 gnd.n54 gnd.n53 53.0052
R8611 gnd.n52 gnd.n51 53.0052
R8612 gnd.n50 gnd.n49 53.0052
R8613 gnd.n48 gnd.n47 53.0052
R8614 gnd.n29 gnd.n28 53.0052
R8615 gnd.n27 gnd.n26 53.0052
R8616 gnd.n25 gnd.n24 53.0052
R8617 gnd.n23 gnd.n22 53.0052
R8618 gnd.n21 gnd.n20 53.0052
R8619 gnd.n19 gnd.n18 53.0052
R8620 gnd.n17 gnd.n16 53.0052
R8621 gnd.n44 gnd.n43 53.0052
R8622 gnd.n42 gnd.n41 53.0052
R8623 gnd.n40 gnd.n39 53.0052
R8624 gnd.n38 gnd.n37 53.0052
R8625 gnd.n36 gnd.n35 53.0052
R8626 gnd.n34 gnd.n33 53.0052
R8627 gnd.n32 gnd.n31 53.0052
R8628 gnd.n5240 gnd.n5239 52.4801
R8629 gnd.n3771 gnd.t140 52.3082
R8630 gnd.n3739 gnd.t173 52.3082
R8631 gnd.n3707 gnd.t145 52.3082
R8632 gnd.n3676 gnd.t311 52.3082
R8633 gnd.n3644 gnd.t16 52.3082
R8634 gnd.n3612 gnd.t147 52.3082
R8635 gnd.n3580 gnd.t149 52.3082
R8636 gnd.n3549 gnd.t134 52.3082
R8637 gnd.n3601 gnd.n3569 51.4173
R8638 gnd.n3665 gnd.n3664 50.455
R8639 gnd.n3633 gnd.n3632 50.455
R8640 gnd.n3601 gnd.n3600 50.455
R8641 gnd.n3014 gnd.n3013 45.1884
R8642 gnd.n2523 gnd.n2522 45.1884
R8643 gnd.n5323 gnd.n5255 44.3322
R8644 gnd.n1969 gnd.n1968 44.3189
R8645 gnd.n1360 gnd.n1359 42.2793
R8646 gnd.n3015 gnd.n3014 42.2793
R8647 gnd.n2524 gnd.n2523 42.2793
R8648 gnd.n2941 gnd.n2940 42.2793
R8649 gnd.n3886 gnd.n2497 42.2793
R8650 gnd.n7217 gnd.n7212 42.2793
R8651 gnd.n5659 gnd.n5658 42.2793
R8652 gnd.n4566 gnd.n2259 42.2793
R8653 gnd.n467 gnd.n466 42.2793
R8654 gnd.n7255 gnd.n176 42.2793
R8655 gnd.n7292 gnd.n7291 42.2793
R8656 gnd.n3952 gnd.n3951 42.2793
R8657 gnd.n3928 gnd.n3927 42.2793
R8658 gnd.n1339 gnd.n1338 42.2793
R8659 gnd.n4123 gnd.n4122 42.2793
R8660 gnd.n1541 gnd.n1540 42.2793
R8661 gnd.n1967 gnd.n1966 41.6274
R8662 gnd.n5250 gnd.n5249 41.6274
R8663 gnd.n1976 gnd.n1975 40.8975
R8664 gnd.n5253 gnd.n5252 40.8975
R8665 gnd.n6189 gnd.n6188 37.4091
R8666 gnd.n6188 gnd.n6187 37.4091
R8667 gnd.n6187 gnd.n943 37.4091
R8668 gnd.n6181 gnd.n943 37.4091
R8669 gnd.n6181 gnd.n6180 37.4091
R8670 gnd.n6180 gnd.n6179 37.4091
R8671 gnd.n6179 gnd.n950 37.4091
R8672 gnd.n6173 gnd.n950 37.4091
R8673 gnd.n6173 gnd.n6172 37.4091
R8674 gnd.n6172 gnd.n6171 37.4091
R8675 gnd.n6171 gnd.n958 37.4091
R8676 gnd.n6165 gnd.n958 37.4091
R8677 gnd.n6165 gnd.n6164 37.4091
R8678 gnd.n6164 gnd.n6163 37.4091
R8679 gnd.n6163 gnd.n966 37.4091
R8680 gnd.n6157 gnd.n966 37.4091
R8681 gnd.n6157 gnd.n6156 37.4091
R8682 gnd.n6156 gnd.n6155 37.4091
R8683 gnd.n6155 gnd.n974 37.4091
R8684 gnd.n6149 gnd.n974 37.4091
R8685 gnd.n6149 gnd.n6148 37.4091
R8686 gnd.n6148 gnd.n6147 37.4091
R8687 gnd.n6147 gnd.n982 37.4091
R8688 gnd.n6141 gnd.n982 37.4091
R8689 gnd.n6141 gnd.n6140 37.4091
R8690 gnd.n6140 gnd.n6139 37.4091
R8691 gnd.n6139 gnd.n990 37.4091
R8692 gnd.n6133 gnd.n990 37.4091
R8693 gnd.n6133 gnd.n6132 37.4091
R8694 gnd.n6132 gnd.n6131 37.4091
R8695 gnd.n6131 gnd.n998 37.4091
R8696 gnd.n6125 gnd.n998 37.4091
R8697 gnd.n6125 gnd.n6124 37.4091
R8698 gnd.n6124 gnd.n6123 37.4091
R8699 gnd.n6123 gnd.n1006 37.4091
R8700 gnd.n6117 gnd.n1006 37.4091
R8701 gnd.n6117 gnd.n6116 37.4091
R8702 gnd.n6116 gnd.n6115 37.4091
R8703 gnd.n6115 gnd.n1014 37.4091
R8704 gnd.n6109 gnd.n1014 37.4091
R8705 gnd.n6109 gnd.n6108 37.4091
R8706 gnd.n6108 gnd.n6107 37.4091
R8707 gnd.n6107 gnd.n1022 37.4091
R8708 gnd.n6101 gnd.n1022 37.4091
R8709 gnd.n6101 gnd.n6100 37.4091
R8710 gnd.n6100 gnd.n6099 37.4091
R8711 gnd.n6099 gnd.n1030 37.4091
R8712 gnd.n6093 gnd.n1030 37.4091
R8713 gnd.n6093 gnd.n6092 37.4091
R8714 gnd.n6092 gnd.n6091 37.4091
R8715 gnd.n6091 gnd.n1038 37.4091
R8716 gnd.n6085 gnd.n1038 37.4091
R8717 gnd.n6085 gnd.n6084 37.4091
R8718 gnd.n6084 gnd.n6083 37.4091
R8719 gnd.n6083 gnd.n1046 37.4091
R8720 gnd.n6077 gnd.n1046 37.4091
R8721 gnd.n6077 gnd.n6076 37.4091
R8722 gnd.n6076 gnd.n6075 37.4091
R8723 gnd.n6075 gnd.n1054 37.4091
R8724 gnd.n6069 gnd.n1054 37.4091
R8725 gnd.n6069 gnd.n6068 37.4091
R8726 gnd.n6068 gnd.n6067 37.4091
R8727 gnd.n6067 gnd.n1062 37.4091
R8728 gnd.n6061 gnd.n1062 37.4091
R8729 gnd.n6061 gnd.n6060 37.4091
R8730 gnd.n6060 gnd.n6059 37.4091
R8731 gnd.n6059 gnd.n1070 37.4091
R8732 gnd.n6053 gnd.n1070 37.4091
R8733 gnd.n6053 gnd.n6052 37.4091
R8734 gnd.n6052 gnd.n6051 37.4091
R8735 gnd.n6051 gnd.n1078 37.4091
R8736 gnd.n6045 gnd.n1078 37.4091
R8737 gnd.n6045 gnd.n6044 37.4091
R8738 gnd.n6044 gnd.n6043 37.4091
R8739 gnd.n6043 gnd.n1086 37.4091
R8740 gnd.n6037 gnd.n1086 37.4091
R8741 gnd.n6037 gnd.n6036 37.4091
R8742 gnd.n6036 gnd.n6035 37.4091
R8743 gnd.n6035 gnd.n1094 37.4091
R8744 gnd.n6029 gnd.n1094 37.4091
R8745 gnd.n6029 gnd.n6028 37.4091
R8746 gnd.n6028 gnd.n6027 37.4091
R8747 gnd.n6027 gnd.n1102 37.4091
R8748 gnd.n6938 gnd.n444 36.9518
R8749 gnd.n1302 gnd.n1301 36.9518
R8750 gnd.n1975 gnd.n1974 35.055
R8751 gnd.n1970 gnd.n1969 35.055
R8752 gnd.n5242 gnd.n5241 35.055
R8753 gnd.n5252 gnd.n5238 35.055
R8754 gnd.n3077 gnd.n2971 31.8661
R8755 gnd.n3077 gnd.n3076 31.8661
R8756 gnd.n3085 gnd.n2960 31.8661
R8757 gnd.n3093 gnd.n2960 31.8661
R8758 gnd.n3093 gnd.n2954 31.8661
R8759 gnd.n3101 gnd.n2954 31.8661
R8760 gnd.n3101 gnd.n2947 31.8661
R8761 gnd.n3139 gnd.n2947 31.8661
R8762 gnd.n3149 gnd.n2880 31.8661
R8763 gnd.n4214 gnd.n4096 31.8661
R8764 gnd.n4222 gnd.n2443 31.8661
R8765 gnd.n4230 gnd.n2443 31.8661
R8766 gnd.n4230 gnd.n2435 31.8661
R8767 gnd.n4238 gnd.n2435 31.8661
R8768 gnd.n4246 gnd.n2426 31.8661
R8769 gnd.n4246 gnd.n2429 31.8661
R8770 gnd.n4254 gnd.n2420 31.8661
R8771 gnd.n4272 gnd.n2402 31.8661
R8772 gnd.n4281 gnd.n2402 31.8661
R8773 gnd.n6020 gnd.n1112 31.8661
R8774 gnd.n4540 gnd.n1271 31.8661
R8775 gnd.n4544 gnd.n4543 31.8661
R8776 gnd.n4544 gnd.n2264 31.8661
R8777 gnd.n4554 gnd.n2284 31.8661
R8778 gnd.n1544 gnd.n1472 31.8661
R8779 gnd.n5629 gnd.n1565 31.8661
R8780 gnd.n1565 gnd.n395 31.8661
R8781 gnd.n470 gnd.n424 31.8661
R8782 gnd.n7114 gnd.n243 31.8661
R8783 gnd.n7130 gnd.n225 31.8661
R8784 gnd.n7130 gnd.n227 31.8661
R8785 gnd.n7138 gnd.n219 31.8661
R8786 gnd.n7146 gnd.n203 31.8661
R8787 gnd.n7154 gnd.n203 31.8661
R8788 gnd.n7162 gnd.n196 31.8661
R8789 gnd.n7162 gnd.n186 31.8661
R8790 gnd.n7172 gnd.n186 31.8661
R8791 gnd.n7172 gnd.n189 31.8661
R8792 gnd.n5329 gnd.n1647 30.7517
R8793 gnd.n2032 gnd.n2030 30.7517
R8794 gnd.n2420 gnd.t194 27.7236
R8795 gnd.n7138 gnd.t228 27.7236
R8796 gnd.n4330 gnd.n1125 26.7676
R8797 gnd.n4324 gnd.n1136 26.7676
R8798 gnd.n4344 gnd.n2378 26.7676
R8799 gnd.n4355 gnd.n2370 26.7676
R8800 gnd.n2373 gnd.n2366 26.7676
R8801 gnd.n4374 gnd.n2360 26.7676
R8802 gnd.n4392 gnd.n2349 26.7676
R8803 gnd.n4430 gnd.n2333 26.7676
R8804 gnd.n4399 gnd.n1155 26.7676
R8805 gnd.n5993 gnd.n1164 26.7676
R8806 gnd.n4404 gnd.n4403 26.7676
R8807 gnd.n5987 gnd.n1173 26.7676
R8808 gnd.n5981 gnd.n1184 26.7676
R8809 gnd.n4470 gnd.n1187 26.7676
R8810 gnd.n4478 gnd.n1197 26.7676
R8811 gnd.n5969 gnd.n1205 26.7676
R8812 gnd.n4486 gnd.n2314 26.7676
R8813 gnd.n5963 gnd.n1215 26.7676
R8814 gnd.n5957 gnd.n1226 26.7676
R8815 gnd.n4522 gnd.n1229 26.7676
R8816 gnd.n4502 gnd.n1239 26.7676
R8817 gnd.n5945 gnd.n1247 26.7676
R8818 gnd.n4511 gnd.n1250 26.7676
R8819 gnd.n5939 gnd.n1258 26.7676
R8820 gnd.n5933 gnd.n1268 26.7676
R8821 gnd.n6894 gnd.n387 26.7676
R8822 gnd.n5616 gnd.n378 26.7676
R8823 gnd.n6983 gnd.n381 26.7676
R8824 gnd.n5610 gnd.n369 26.7676
R8825 gnd.n6991 gnd.n372 26.7676
R8826 gnd.n6999 gnd.n363 26.7676
R8827 gnd.n5602 gnd.n352 26.7676
R8828 gnd.n5598 gnd.n343 26.7676
R8829 gnd.n7015 gnd.n346 26.7676
R8830 gnd.n5512 gnd.n334 26.7676
R8831 gnd.n7023 gnd.n337 26.7676
R8832 gnd.n7031 gnd.n328 26.7676
R8833 gnd.n5522 gnd.n317 26.7676
R8834 gnd.n5582 gnd.n306 26.7676
R8835 gnd.n7048 gnd.n309 26.7676
R8836 gnd.n5576 gnd.n5575 26.7676
R8837 gnd.n5533 gnd.n297 26.7676
R8838 gnd.n5554 gnd.n288 26.7676
R8839 gnd.n7066 gnd.n291 26.7676
R8840 gnd.n7074 gnd.n284 26.7676
R8841 gnd.n7083 gnd.n274 26.7676
R8842 gnd.n6841 gnd.n266 26.7676
R8843 gnd.n6837 gnd.n258 26.7676
R8844 gnd.n7098 gnd.n260 26.7676
R8845 gnd.n7106 gnd.n252 26.7676
R8846 gnd.t188 gnd.n4362 26.4489
R8847 gnd.n6845 gnd.t265 26.4489
R8848 gnd.n6014 gnd.t222 25.8116
R8849 gnd.n545 gnd.t277 25.8116
R8850 gnd.n1359 gnd.n1358 25.7944
R8851 gnd.n2940 gnd.n2939 25.7944
R8852 gnd.n2497 gnd.n2496 25.7944
R8853 gnd.n7212 gnd.n7211 25.7944
R8854 gnd.n5658 gnd.n5657 25.7944
R8855 gnd.n2259 gnd.n2258 25.7944
R8856 gnd.n444 gnd.n443 25.7944
R8857 gnd.n466 gnd.n465 25.7944
R8858 gnd.n176 gnd.n175 25.7944
R8859 gnd.n7291 gnd.n7290 25.7944
R8860 gnd.n3951 gnd.n3950 25.7944
R8861 gnd.n3927 gnd.n3926 25.7944
R8862 gnd.n1338 gnd.n1337 25.7944
R8863 gnd.n1301 gnd.n1300 25.7944
R8864 gnd.n4122 gnd.n4121 25.7944
R8865 gnd.n1540 gnd.n1539 25.7944
R8866 gnd.n4254 gnd.t251 25.1743
R8867 gnd.n6021 gnd.n6020 25.1743
R8868 gnd.n243 gnd.n233 25.1743
R8869 gnd.n219 gnd.t213 25.1743
R8870 gnd.n3161 gnd.n2881 24.8557
R8871 gnd.n3171 gnd.n2864 24.8557
R8872 gnd.n2867 gnd.n2855 24.8557
R8873 gnd.n3192 gnd.n2856 24.8557
R8874 gnd.n3202 gnd.n2836 24.8557
R8875 gnd.n3212 gnd.n3211 24.8557
R8876 gnd.n2822 gnd.n2820 24.8557
R8877 gnd.n3243 gnd.n3242 24.8557
R8878 gnd.n3258 gnd.n2805 24.8557
R8879 gnd.n3312 gnd.n2744 24.8557
R8880 gnd.n3268 gnd.n2745 24.8557
R8881 gnd.n3305 gnd.n2756 24.8557
R8882 gnd.n2794 gnd.n2793 24.8557
R8883 gnd.n3299 gnd.n3298 24.8557
R8884 gnd.n2780 gnd.n2767 24.8557
R8885 gnd.n3338 gnd.n3337 24.8557
R8886 gnd.n3348 gnd.n2676 24.8557
R8887 gnd.n3360 gnd.n2668 24.8557
R8888 gnd.n3359 gnd.n2656 24.8557
R8889 gnd.n3378 gnd.n3377 24.8557
R8890 gnd.n3388 gnd.n2649 24.8557
R8891 gnd.n3399 gnd.n2637 24.8557
R8892 gnd.n3423 gnd.n3422 24.8557
R8893 gnd.n3434 gnd.n2620 24.8557
R8894 gnd.n3433 gnd.n2622 24.8557
R8895 gnd.n3445 gnd.n2613 24.8557
R8896 gnd.n3463 gnd.n3462 24.8557
R8897 gnd.n2604 gnd.n2593 24.8557
R8898 gnd.n3484 gnd.n2581 24.8557
R8899 gnd.n3512 gnd.n3511 24.8557
R8900 gnd.n3523 gnd.n2565 24.8557
R8901 gnd.n3534 gnd.n2558 24.8557
R8902 gnd.n3533 gnd.n2546 24.8557
R8903 gnd.n3806 gnd.n3805 24.8557
R8904 gnd.n3828 gnd.n2531 24.8557
R8905 gnd.n3182 gnd.t133 23.2624
R8906 gnd.n2883 gnd.t39 22.6251
R8907 gnd.n4096 gnd.t64 22.6251
R8908 gnd.n5856 gnd.t50 22.6251
R8909 gnd.n6975 gnd.t32 22.6251
R8910 gnd.n7248 gnd.t18 22.6251
R8911 gnd.n2573 gnd.n1102 22.4457
R8912 gnd.n4331 gnd.t196 21.9878
R8913 gnd.t268 gnd.n249 21.9878
R8914 gnd.t310 gnd.n2888 21.3504
R8915 gnd.n4373 gnd.t226 21.3504
R8916 gnd.t257 gnd.n281 21.3504
R8917 gnd.t151 gnd.n2594 20.7131
R8918 gnd.t211 gnd.n1176 20.7131
R8919 gnd.n5583 gnd.t240 20.7131
R8920 gnd.n4540 gnd.n1276 20.3945
R8921 gnd.n6966 gnd.n424 20.3945
R8922 gnd.n7327 gnd.n100 20.3945
R8923 gnd.t153 gnd.n2629 20.0758
R8924 gnd.t201 gnd.n1218 20.0758
R8925 gnd.n5597 gnd.t209 20.0758
R8926 gnd.n2029 gnd.n2028 19.9763
R8927 gnd.n1646 gnd.n1645 19.9763
R8928 gnd.n2026 gnd.n2025 19.9763
R8929 gnd.n5257 gnd.n5256 19.9763
R8930 gnd.n1963 gnd.t86 19.8005
R8931 gnd.n1963 gnd.t23 19.8005
R8932 gnd.n1964 gnd.t115 19.8005
R8933 gnd.n1964 gnd.t124 19.8005
R8934 gnd.n5246 gnd.t69 19.8005
R8935 gnd.n5246 gnd.t99 19.8005
R8936 gnd.n5247 gnd.t48 19.8005
R8937 gnd.n5247 gnd.t96 19.8005
R8938 gnd.n1960 gnd.n1959 19.5087
R8939 gnd.n1973 gnd.n1960 19.5087
R8940 gnd.n1971 gnd.n1962 19.5087
R8941 gnd.n5251 gnd.n5245 19.5087
R8942 gnd.n3349 gnd.t159 19.4385
R8943 gnd.n5832 gnd.n5831 19.3944
R8944 gnd.n5831 gnd.n5830 19.3944
R8945 gnd.n5830 gnd.n1370 19.3944
R8946 gnd.n5826 gnd.n1370 19.3944
R8947 gnd.n5826 gnd.n5825 19.3944
R8948 gnd.n5825 gnd.n5824 19.3944
R8949 gnd.n5824 gnd.n1375 19.3944
R8950 gnd.n5820 gnd.n1375 19.3944
R8951 gnd.n5820 gnd.n5819 19.3944
R8952 gnd.n5819 gnd.n5818 19.3944
R8953 gnd.n5818 gnd.n1380 19.3944
R8954 gnd.n5814 gnd.n1380 19.3944
R8955 gnd.n5814 gnd.n5813 19.3944
R8956 gnd.n5813 gnd.n5812 19.3944
R8957 gnd.n5812 gnd.n1385 19.3944
R8958 gnd.n5808 gnd.n1385 19.3944
R8959 gnd.n5808 gnd.n5807 19.3944
R8960 gnd.n5807 gnd.n5806 19.3944
R8961 gnd.n5806 gnd.n1390 19.3944
R8962 gnd.n5802 gnd.n1390 19.3944
R8963 gnd.n5802 gnd.n5801 19.3944
R8964 gnd.n5801 gnd.n5800 19.3944
R8965 gnd.n5800 gnd.n1395 19.3944
R8966 gnd.n5796 gnd.n1395 19.3944
R8967 gnd.n5796 gnd.n5795 19.3944
R8968 gnd.n5795 gnd.n5794 19.3944
R8969 gnd.n5794 gnd.n1400 19.3944
R8970 gnd.n5790 gnd.n1400 19.3944
R8971 gnd.n5790 gnd.n5789 19.3944
R8972 gnd.n5789 gnd.n5788 19.3944
R8973 gnd.n5788 gnd.n1405 19.3944
R8974 gnd.n5784 gnd.n1405 19.3944
R8975 gnd.n5784 gnd.n5783 19.3944
R8976 gnd.n5783 gnd.n5782 19.3944
R8977 gnd.n5782 gnd.n1410 19.3944
R8978 gnd.n5778 gnd.n1410 19.3944
R8979 gnd.n5778 gnd.n5777 19.3944
R8980 gnd.n5777 gnd.n5776 19.3944
R8981 gnd.n5776 gnd.n1415 19.3944
R8982 gnd.n5772 gnd.n1415 19.3944
R8983 gnd.n5772 gnd.n5771 19.3944
R8984 gnd.n5771 gnd.n5770 19.3944
R8985 gnd.n5770 gnd.n1420 19.3944
R8986 gnd.n5766 gnd.n1420 19.3944
R8987 gnd.n5766 gnd.n5765 19.3944
R8988 gnd.n5765 gnd.n5764 19.3944
R8989 gnd.n5764 gnd.n1425 19.3944
R8990 gnd.n5760 gnd.n1425 19.3944
R8991 gnd.n5760 gnd.n5759 19.3944
R8992 gnd.n5759 gnd.n5758 19.3944
R8993 gnd.n5758 gnd.n1430 19.3944
R8994 gnd.n5754 gnd.n1430 19.3944
R8995 gnd.n5754 gnd.n5753 19.3944
R8996 gnd.n5753 gnd.n5752 19.3944
R8997 gnd.n5752 gnd.n1435 19.3944
R8998 gnd.n5748 gnd.n1435 19.3944
R8999 gnd.n5748 gnd.n5747 19.3944
R9000 gnd.n5747 gnd.n5746 19.3944
R9001 gnd.n5746 gnd.n1440 19.3944
R9002 gnd.n5742 gnd.n1440 19.3944
R9003 gnd.n5742 gnd.n5741 19.3944
R9004 gnd.n5741 gnd.n5740 19.3944
R9005 gnd.n5740 gnd.n1445 19.3944
R9006 gnd.n5736 gnd.n1445 19.3944
R9007 gnd.n5736 gnd.n5735 19.3944
R9008 gnd.n5735 gnd.n5734 19.3944
R9009 gnd.n5734 gnd.n1450 19.3944
R9010 gnd.n5730 gnd.n1450 19.3944
R9011 gnd.n5730 gnd.n5729 19.3944
R9012 gnd.n5729 gnd.n5728 19.3944
R9013 gnd.n5728 gnd.n1455 19.3944
R9014 gnd.n5724 gnd.n1455 19.3944
R9015 gnd.n5724 gnd.n5723 19.3944
R9016 gnd.n5723 gnd.n5722 19.3944
R9017 gnd.n5722 gnd.n1460 19.3944
R9018 gnd.n5718 gnd.n1460 19.3944
R9019 gnd.n5718 gnd.n5717 19.3944
R9020 gnd.n5717 gnd.n5716 19.3944
R9021 gnd.n5716 gnd.n1465 19.3944
R9022 gnd.n5712 gnd.n1465 19.3944
R9023 gnd.n5712 gnd.n5711 19.3944
R9024 gnd.n5711 gnd.n5710 19.3944
R9025 gnd.n5838 gnd.n5837 19.3944
R9026 gnd.n5837 gnd.n5836 19.3944
R9027 gnd.n5836 gnd.n1365 19.3944
R9028 gnd.n4603 gnd.n2208 19.3944
R9029 gnd.n4603 gnd.n4602 19.3944
R9030 gnd.n4602 gnd.n2211 19.3944
R9031 gnd.n4595 gnd.n2211 19.3944
R9032 gnd.n4595 gnd.n4594 19.3944
R9033 gnd.n4594 gnd.n2221 19.3944
R9034 gnd.n4587 gnd.n2221 19.3944
R9035 gnd.n4587 gnd.n4586 19.3944
R9036 gnd.n4586 gnd.n2232 19.3944
R9037 gnd.n4579 gnd.n2232 19.3944
R9038 gnd.n4579 gnd.n4578 19.3944
R9039 gnd.n4578 gnd.n2242 19.3944
R9040 gnd.n4571 gnd.n2242 19.3944
R9041 gnd.n4571 gnd.n4570 19.3944
R9042 gnd.n4570 gnd.n2253 19.3944
R9043 gnd.n4560 gnd.n2253 19.3944
R9044 gnd.n4560 gnd.n1349 19.3944
R9045 gnd.n5849 gnd.n1349 19.3944
R9046 gnd.n5849 gnd.n5848 19.3944
R9047 gnd.n5848 gnd.n5847 19.3944
R9048 gnd.n5847 gnd.n1353 19.3944
R9049 gnd.n5843 gnd.n1353 19.3944
R9050 gnd.n5843 gnd.n5842 19.3944
R9051 gnd.n5842 gnd.n5841 19.3944
R9052 gnd.n3064 gnd.n3063 19.3944
R9053 gnd.n3063 gnd.n3062 19.3944
R9054 gnd.n3062 gnd.n3061 19.3944
R9055 gnd.n3061 gnd.n3059 19.3944
R9056 gnd.n3059 gnd.n3056 19.3944
R9057 gnd.n3056 gnd.n3055 19.3944
R9058 gnd.n3055 gnd.n3052 19.3944
R9059 gnd.n3052 gnd.n3051 19.3944
R9060 gnd.n3051 gnd.n3048 19.3944
R9061 gnd.n3048 gnd.n3047 19.3944
R9062 gnd.n3047 gnd.n3044 19.3944
R9063 gnd.n3044 gnd.n3043 19.3944
R9064 gnd.n3043 gnd.n3040 19.3944
R9065 gnd.n3040 gnd.n3039 19.3944
R9066 gnd.n3039 gnd.n3036 19.3944
R9067 gnd.n3036 gnd.n3035 19.3944
R9068 gnd.n3035 gnd.n3032 19.3944
R9069 gnd.n3032 gnd.n3031 19.3944
R9070 gnd.n3031 gnd.n3028 19.3944
R9071 gnd.n3028 gnd.n3027 19.3944
R9072 gnd.n3027 gnd.n3024 19.3944
R9073 gnd.n3024 gnd.n3023 19.3944
R9074 gnd.n3020 gnd.n3019 19.3944
R9075 gnd.n3019 gnd.n2975 19.3944
R9076 gnd.n3070 gnd.n2975 19.3944
R9077 gnd.n3836 gnd.n3835 19.3944
R9078 gnd.n3835 gnd.n3832 19.3944
R9079 gnd.n3832 gnd.n3831 19.3944
R9080 gnd.n3881 gnd.n3880 19.3944
R9081 gnd.n3880 gnd.n3879 19.3944
R9082 gnd.n3879 gnd.n3876 19.3944
R9083 gnd.n3876 gnd.n3875 19.3944
R9084 gnd.n3875 gnd.n3872 19.3944
R9085 gnd.n3872 gnd.n3871 19.3944
R9086 gnd.n3871 gnd.n3868 19.3944
R9087 gnd.n3868 gnd.n3867 19.3944
R9088 gnd.n3867 gnd.n3864 19.3944
R9089 gnd.n3864 gnd.n3863 19.3944
R9090 gnd.n3863 gnd.n3860 19.3944
R9091 gnd.n3860 gnd.n3859 19.3944
R9092 gnd.n3859 gnd.n3856 19.3944
R9093 gnd.n3856 gnd.n3855 19.3944
R9094 gnd.n3855 gnd.n3852 19.3944
R9095 gnd.n3852 gnd.n3851 19.3944
R9096 gnd.n3851 gnd.n3848 19.3944
R9097 gnd.n3848 gnd.n3847 19.3944
R9098 gnd.n3847 gnd.n3844 19.3944
R9099 gnd.n3844 gnd.n3843 19.3944
R9100 gnd.n3843 gnd.n3840 19.3944
R9101 gnd.n3840 gnd.n3839 19.3944
R9102 gnd.n3163 gnd.n2872 19.3944
R9103 gnd.n3173 gnd.n2872 19.3944
R9104 gnd.n3174 gnd.n3173 19.3944
R9105 gnd.n3174 gnd.n2853 19.3944
R9106 gnd.n3194 gnd.n2853 19.3944
R9107 gnd.n3194 gnd.n2845 19.3944
R9108 gnd.n3204 gnd.n2845 19.3944
R9109 gnd.n3205 gnd.n3204 19.3944
R9110 gnd.n3206 gnd.n3205 19.3944
R9111 gnd.n3206 gnd.n2828 19.3944
R9112 gnd.n3223 gnd.n2828 19.3944
R9113 gnd.n3226 gnd.n3223 19.3944
R9114 gnd.n3226 gnd.n3225 19.3944
R9115 gnd.n3225 gnd.n2801 19.3944
R9116 gnd.n3265 gnd.n2801 19.3944
R9117 gnd.n3265 gnd.n2798 19.3944
R9118 gnd.n3271 gnd.n2798 19.3944
R9119 gnd.n3272 gnd.n3271 19.3944
R9120 gnd.n3272 gnd.n2796 19.3944
R9121 gnd.n3278 gnd.n2796 19.3944
R9122 gnd.n3281 gnd.n3278 19.3944
R9123 gnd.n3283 gnd.n3281 19.3944
R9124 gnd.n3289 gnd.n3283 19.3944
R9125 gnd.n3289 gnd.n3288 19.3944
R9126 gnd.n3288 gnd.n2671 19.3944
R9127 gnd.n3355 gnd.n2671 19.3944
R9128 gnd.n3356 gnd.n3355 19.3944
R9129 gnd.n3356 gnd.n2664 19.3944
R9130 gnd.n3367 gnd.n2664 19.3944
R9131 gnd.n3368 gnd.n3367 19.3944
R9132 gnd.n3368 gnd.n2647 19.3944
R9133 gnd.n2647 gnd.n2645 19.3944
R9134 gnd.n3392 gnd.n2645 19.3944
R9135 gnd.n3393 gnd.n3392 19.3944
R9136 gnd.n3393 gnd.n2616 19.3944
R9137 gnd.n3440 gnd.n2616 19.3944
R9138 gnd.n3441 gnd.n3440 19.3944
R9139 gnd.n3441 gnd.n2609 19.3944
R9140 gnd.n3452 gnd.n2609 19.3944
R9141 gnd.n3453 gnd.n3452 19.3944
R9142 gnd.n3453 gnd.n2592 19.3944
R9143 gnd.n2592 gnd.n2590 19.3944
R9144 gnd.n3477 gnd.n2590 19.3944
R9145 gnd.n3478 gnd.n3477 19.3944
R9146 gnd.n3478 gnd.n2561 19.3944
R9147 gnd.n3529 gnd.n2561 19.3944
R9148 gnd.n3530 gnd.n3529 19.3944
R9149 gnd.n3530 gnd.n2554 19.3944
R9150 gnd.n3797 gnd.n2554 19.3944
R9151 gnd.n3798 gnd.n3797 19.3944
R9152 gnd.n3798 gnd.n2535 19.3944
R9153 gnd.n3823 gnd.n2535 19.3944
R9154 gnd.n3823 gnd.n2536 19.3944
R9155 gnd.n3154 gnd.n3153 19.3944
R9156 gnd.n3153 gnd.n2886 19.3944
R9157 gnd.n2909 gnd.n2886 19.3944
R9158 gnd.n2912 gnd.n2909 19.3944
R9159 gnd.n2912 gnd.n2905 19.3944
R9160 gnd.n2916 gnd.n2905 19.3944
R9161 gnd.n2919 gnd.n2916 19.3944
R9162 gnd.n2922 gnd.n2919 19.3944
R9163 gnd.n2922 gnd.n2903 19.3944
R9164 gnd.n2926 gnd.n2903 19.3944
R9165 gnd.n2929 gnd.n2926 19.3944
R9166 gnd.n2932 gnd.n2929 19.3944
R9167 gnd.n2932 gnd.n2901 19.3944
R9168 gnd.n2936 gnd.n2901 19.3944
R9169 gnd.n3159 gnd.n3158 19.3944
R9170 gnd.n3158 gnd.n2862 19.3944
R9171 gnd.n3184 gnd.n2862 19.3944
R9172 gnd.n3184 gnd.n2860 19.3944
R9173 gnd.n3190 gnd.n2860 19.3944
R9174 gnd.n3190 gnd.n3189 19.3944
R9175 gnd.n3189 gnd.n2834 19.3944
R9176 gnd.n3214 gnd.n2834 19.3944
R9177 gnd.n3214 gnd.n2832 19.3944
R9178 gnd.n3218 gnd.n2832 19.3944
R9179 gnd.n3218 gnd.n2812 19.3944
R9180 gnd.n3245 gnd.n2812 19.3944
R9181 gnd.n3245 gnd.n2810 19.3944
R9182 gnd.n3255 gnd.n2810 19.3944
R9183 gnd.n3255 gnd.n3254 19.3944
R9184 gnd.n3254 gnd.n3253 19.3944
R9185 gnd.n3253 gnd.n2759 19.3944
R9186 gnd.n3303 gnd.n2759 19.3944
R9187 gnd.n3303 gnd.n3302 19.3944
R9188 gnd.n3302 gnd.n3301 19.3944
R9189 gnd.n3301 gnd.n2763 19.3944
R9190 gnd.n2783 gnd.n2763 19.3944
R9191 gnd.n2783 gnd.n2681 19.3944
R9192 gnd.n3340 gnd.n2681 19.3944
R9193 gnd.n3340 gnd.n2679 19.3944
R9194 gnd.n3346 gnd.n2679 19.3944
R9195 gnd.n3346 gnd.n3345 19.3944
R9196 gnd.n3345 gnd.n2654 19.3944
R9197 gnd.n3380 gnd.n2654 19.3944
R9198 gnd.n3380 gnd.n2652 19.3944
R9199 gnd.n3386 gnd.n2652 19.3944
R9200 gnd.n3386 gnd.n3385 19.3944
R9201 gnd.n3385 gnd.n2627 19.3944
R9202 gnd.n3425 gnd.n2627 19.3944
R9203 gnd.n3425 gnd.n2625 19.3944
R9204 gnd.n3431 gnd.n2625 19.3944
R9205 gnd.n3431 gnd.n3430 19.3944
R9206 gnd.n3430 gnd.n2599 19.3944
R9207 gnd.n3465 gnd.n2599 19.3944
R9208 gnd.n3465 gnd.n2597 19.3944
R9209 gnd.n3471 gnd.n2597 19.3944
R9210 gnd.n3471 gnd.n3470 19.3944
R9211 gnd.n3470 gnd.n2571 19.3944
R9212 gnd.n3514 gnd.n2571 19.3944
R9213 gnd.n3514 gnd.n2569 19.3944
R9214 gnd.n3520 gnd.n2569 19.3944
R9215 gnd.n3520 gnd.n3519 19.3944
R9216 gnd.n3519 gnd.n2544 19.3944
R9217 gnd.n3808 gnd.n2544 19.3944
R9218 gnd.n3808 gnd.n2542 19.3944
R9219 gnd.n3816 gnd.n2542 19.3944
R9220 gnd.n3816 gnd.n3815 19.3944
R9221 gnd.n3815 gnd.n3814 19.3944
R9222 gnd.n3917 gnd.n3916 19.3944
R9223 gnd.n3916 gnd.n2483 19.3944
R9224 gnd.n3912 gnd.n2483 19.3944
R9225 gnd.n3912 gnd.n3909 19.3944
R9226 gnd.n3909 gnd.n3906 19.3944
R9227 gnd.n3906 gnd.n3905 19.3944
R9228 gnd.n3905 gnd.n3902 19.3944
R9229 gnd.n3902 gnd.n3901 19.3944
R9230 gnd.n3901 gnd.n3898 19.3944
R9231 gnd.n3898 gnd.n3897 19.3944
R9232 gnd.n3897 gnd.n3894 19.3944
R9233 gnd.n3894 gnd.n3893 19.3944
R9234 gnd.n3893 gnd.n3890 19.3944
R9235 gnd.n3890 gnd.n3889 19.3944
R9236 gnd.n3074 gnd.n2973 19.3944
R9237 gnd.n3074 gnd.n2964 19.3944
R9238 gnd.n3087 gnd.n2964 19.3944
R9239 gnd.n3087 gnd.n2962 19.3944
R9240 gnd.n3091 gnd.n2962 19.3944
R9241 gnd.n3091 gnd.n2952 19.3944
R9242 gnd.n3103 gnd.n2952 19.3944
R9243 gnd.n3103 gnd.n2950 19.3944
R9244 gnd.n3137 gnd.n2950 19.3944
R9245 gnd.n3137 gnd.n3136 19.3944
R9246 gnd.n3136 gnd.n3135 19.3944
R9247 gnd.n3135 gnd.n3134 19.3944
R9248 gnd.n3134 gnd.n3131 19.3944
R9249 gnd.n3131 gnd.n3130 19.3944
R9250 gnd.n3130 gnd.n3129 19.3944
R9251 gnd.n3129 gnd.n3127 19.3944
R9252 gnd.n3127 gnd.n3126 19.3944
R9253 gnd.n3126 gnd.n3123 19.3944
R9254 gnd.n3123 gnd.n3122 19.3944
R9255 gnd.n3122 gnd.n3121 19.3944
R9256 gnd.n3121 gnd.n3119 19.3944
R9257 gnd.n3119 gnd.n2818 19.3944
R9258 gnd.n3234 gnd.n2818 19.3944
R9259 gnd.n3234 gnd.n2816 19.3944
R9260 gnd.n3240 gnd.n2816 19.3944
R9261 gnd.n3240 gnd.n3239 19.3944
R9262 gnd.n3239 gnd.n2740 19.3944
R9263 gnd.n3314 gnd.n2740 19.3944
R9264 gnd.n3314 gnd.n2741 19.3944
R9265 gnd.n2788 gnd.n2787 19.3944
R9266 gnd.n2791 gnd.n2790 19.3944
R9267 gnd.n2778 gnd.n2777 19.3944
R9268 gnd.n3333 gnd.n2686 19.3944
R9269 gnd.n3333 gnd.n3332 19.3944
R9270 gnd.n3332 gnd.n3331 19.3944
R9271 gnd.n3331 gnd.n3329 19.3944
R9272 gnd.n3329 gnd.n3328 19.3944
R9273 gnd.n3328 gnd.n3326 19.3944
R9274 gnd.n3326 gnd.n3325 19.3944
R9275 gnd.n3325 gnd.n2635 19.3944
R9276 gnd.n3401 gnd.n2635 19.3944
R9277 gnd.n3401 gnd.n2633 19.3944
R9278 gnd.n3420 gnd.n2633 19.3944
R9279 gnd.n3420 gnd.n3419 19.3944
R9280 gnd.n3419 gnd.n3418 19.3944
R9281 gnd.n3418 gnd.n3416 19.3944
R9282 gnd.n3416 gnd.n3415 19.3944
R9283 gnd.n3415 gnd.n3413 19.3944
R9284 gnd.n3413 gnd.n3412 19.3944
R9285 gnd.n3412 gnd.n2579 19.3944
R9286 gnd.n3486 gnd.n2579 19.3944
R9287 gnd.n3486 gnd.n2577 19.3944
R9288 gnd.n3509 gnd.n2577 19.3944
R9289 gnd.n3509 gnd.n3508 19.3944
R9290 gnd.n3508 gnd.n3507 19.3944
R9291 gnd.n3507 gnd.n3504 19.3944
R9292 gnd.n3504 gnd.n3503 19.3944
R9293 gnd.n3503 gnd.n3501 19.3944
R9294 gnd.n3501 gnd.n3500 19.3944
R9295 gnd.n3500 gnd.n3498 19.3944
R9296 gnd.n3498 gnd.n2530 19.3944
R9297 gnd.n3079 gnd.n2969 19.3944
R9298 gnd.n3079 gnd.n2967 19.3944
R9299 gnd.n3083 gnd.n2967 19.3944
R9300 gnd.n3083 gnd.n2958 19.3944
R9301 gnd.n3095 gnd.n2958 19.3944
R9302 gnd.n3095 gnd.n2956 19.3944
R9303 gnd.n3099 gnd.n2956 19.3944
R9304 gnd.n3099 gnd.n2945 19.3944
R9305 gnd.n3141 gnd.n2945 19.3944
R9306 gnd.n3141 gnd.n2899 19.3944
R9307 gnd.n3147 gnd.n2899 19.3944
R9308 gnd.n3147 gnd.n3146 19.3944
R9309 gnd.n3146 gnd.n2877 19.3944
R9310 gnd.n3168 gnd.n2877 19.3944
R9311 gnd.n3168 gnd.n2870 19.3944
R9312 gnd.n3179 gnd.n2870 19.3944
R9313 gnd.n3179 gnd.n3178 19.3944
R9314 gnd.n3178 gnd.n2851 19.3944
R9315 gnd.n3199 gnd.n2851 19.3944
R9316 gnd.n3199 gnd.n2841 19.3944
R9317 gnd.n3209 gnd.n2841 19.3944
R9318 gnd.n3209 gnd.n2824 19.3944
R9319 gnd.n3230 gnd.n2824 19.3944
R9320 gnd.n3230 gnd.n3229 19.3944
R9321 gnd.n3229 gnd.n2803 19.3944
R9322 gnd.n3260 gnd.n2803 19.3944
R9323 gnd.n3260 gnd.n2748 19.3944
R9324 gnd.n3310 gnd.n2748 19.3944
R9325 gnd.n3310 gnd.n3309 19.3944
R9326 gnd.n3309 gnd.n3308 19.3944
R9327 gnd.n3308 gnd.n2752 19.3944
R9328 gnd.n2770 gnd.n2752 19.3944
R9329 gnd.n3296 gnd.n2770 19.3944
R9330 gnd.n3296 gnd.n3295 19.3944
R9331 gnd.n3295 gnd.n3294 19.3944
R9332 gnd.n3294 gnd.n2774 19.3944
R9333 gnd.n2774 gnd.n2673 19.3944
R9334 gnd.n3351 gnd.n2673 19.3944
R9335 gnd.n3351 gnd.n2666 19.3944
R9336 gnd.n3362 gnd.n2666 19.3944
R9337 gnd.n3362 gnd.n2662 19.3944
R9338 gnd.n3375 gnd.n2662 19.3944
R9339 gnd.n3375 gnd.n3374 19.3944
R9340 gnd.n3374 gnd.n2641 19.3944
R9341 gnd.n3397 gnd.n2641 19.3944
R9342 gnd.n3397 gnd.n3396 19.3944
R9343 gnd.n3396 gnd.n2618 19.3944
R9344 gnd.n3436 gnd.n2618 19.3944
R9345 gnd.n3436 gnd.n2611 19.3944
R9346 gnd.n3447 gnd.n2611 19.3944
R9347 gnd.n3447 gnd.n2607 19.3944
R9348 gnd.n3460 gnd.n2607 19.3944
R9349 gnd.n3460 gnd.n3459 19.3944
R9350 gnd.n3459 gnd.n2586 19.3944
R9351 gnd.n3482 gnd.n2586 19.3944
R9352 gnd.n3482 gnd.n3481 19.3944
R9353 gnd.n3481 gnd.n2563 19.3944
R9354 gnd.n3525 gnd.n2563 19.3944
R9355 gnd.n3525 gnd.n2556 19.3944
R9356 gnd.n3536 gnd.n2556 19.3944
R9357 gnd.n3536 gnd.n2552 19.3944
R9358 gnd.n3803 gnd.n2552 19.3944
R9359 gnd.n3803 gnd.n3802 19.3944
R9360 gnd.n3802 gnd.n2533 19.3944
R9361 gnd.n3826 gnd.n2533 19.3944
R9362 gnd.n6892 gnd.n471 19.3944
R9363 gnd.n6888 gnd.n471 19.3944
R9364 gnd.n6888 gnd.n6887 19.3944
R9365 gnd.n6887 gnd.n6886 19.3944
R9366 gnd.n6886 gnd.n476 19.3944
R9367 gnd.n6882 gnd.n476 19.3944
R9368 gnd.n6882 gnd.n6881 19.3944
R9369 gnd.n6881 gnd.n6880 19.3944
R9370 gnd.n6880 gnd.n480 19.3944
R9371 gnd.n6876 gnd.n480 19.3944
R9372 gnd.n6876 gnd.n6875 19.3944
R9373 gnd.n6875 gnd.n6874 19.3944
R9374 gnd.n6874 gnd.n484 19.3944
R9375 gnd.n6870 gnd.n484 19.3944
R9376 gnd.n6870 gnd.n6869 19.3944
R9377 gnd.n6869 gnd.n6868 19.3944
R9378 gnd.n6868 gnd.n488 19.3944
R9379 gnd.n6864 gnd.n488 19.3944
R9380 gnd.n6864 gnd.n6863 19.3944
R9381 gnd.n6863 gnd.n6862 19.3944
R9382 gnd.n6862 gnd.n492 19.3944
R9383 gnd.n6858 gnd.n492 19.3944
R9384 gnd.n6858 gnd.n6857 19.3944
R9385 gnd.n6857 gnd.n6856 19.3944
R9386 gnd.n6856 gnd.n6853 19.3944
R9387 gnd.n6853 gnd.n65 19.3944
R9388 gnd.n7367 gnd.n65 19.3944
R9389 gnd.n7367 gnd.n7366 19.3944
R9390 gnd.n7366 gnd.n7365 19.3944
R9391 gnd.n7365 gnd.n69 19.3944
R9392 gnd.n7361 gnd.n69 19.3944
R9393 gnd.n7361 gnd.n7360 19.3944
R9394 gnd.n7360 gnd.n7359 19.3944
R9395 gnd.n7359 gnd.n74 19.3944
R9396 gnd.n7355 gnd.n74 19.3944
R9397 gnd.n7355 gnd.n7354 19.3944
R9398 gnd.n7354 gnd.n7353 19.3944
R9399 gnd.n7353 gnd.n79 19.3944
R9400 gnd.n7349 gnd.n79 19.3944
R9401 gnd.n7349 gnd.n7348 19.3944
R9402 gnd.n7348 gnd.n7347 19.3944
R9403 gnd.n7347 gnd.n84 19.3944
R9404 gnd.n7343 gnd.n84 19.3944
R9405 gnd.n7343 gnd.n7342 19.3944
R9406 gnd.n7342 gnd.n7341 19.3944
R9407 gnd.n7341 gnd.n89 19.3944
R9408 gnd.n7337 gnd.n89 19.3944
R9409 gnd.n7337 gnd.n7336 19.3944
R9410 gnd.n7336 gnd.n7335 19.3944
R9411 gnd.n7335 gnd.n94 19.3944
R9412 gnd.n7331 gnd.n94 19.3944
R9413 gnd.n7331 gnd.n7330 19.3944
R9414 gnd.n7330 gnd.n7329 19.3944
R9415 gnd.n7242 gnd.n7241 19.3944
R9416 gnd.n7241 gnd.n7240 19.3944
R9417 gnd.n7240 gnd.n7182 19.3944
R9418 gnd.n7236 gnd.n7182 19.3944
R9419 gnd.n7236 gnd.n7235 19.3944
R9420 gnd.n7235 gnd.n7234 19.3944
R9421 gnd.n7234 gnd.n7190 19.3944
R9422 gnd.n7230 gnd.n7190 19.3944
R9423 gnd.n7230 gnd.n7229 19.3944
R9424 gnd.n7229 gnd.n7228 19.3944
R9425 gnd.n7228 gnd.n7198 19.3944
R9426 gnd.n7224 gnd.n7198 19.3944
R9427 gnd.n7224 gnd.n7223 19.3944
R9428 gnd.n7223 gnd.n7222 19.3944
R9429 gnd.n7222 gnd.n7206 19.3944
R9430 gnd.n7218 gnd.n7206 19.3944
R9431 gnd.n5702 gnd.n5700 19.3944
R9432 gnd.n5700 gnd.n5699 19.3944
R9433 gnd.n5699 gnd.n1480 19.3944
R9434 gnd.n5692 gnd.n1480 19.3944
R9435 gnd.n5692 gnd.n5691 19.3944
R9436 gnd.n5691 gnd.n1492 19.3944
R9437 gnd.n5684 gnd.n1492 19.3944
R9438 gnd.n5684 gnd.n5683 19.3944
R9439 gnd.n5683 gnd.n1500 19.3944
R9440 gnd.n5676 gnd.n1500 19.3944
R9441 gnd.n5676 gnd.n5675 19.3944
R9442 gnd.n5675 gnd.n1510 19.3944
R9443 gnd.n5668 gnd.n1510 19.3944
R9444 gnd.n5668 gnd.n5667 19.3944
R9445 gnd.n5667 gnd.n1518 19.3944
R9446 gnd.n5660 gnd.n1518 19.3944
R9447 gnd.n6977 gnd.n385 19.3944
R9448 gnd.n6977 gnd.n383 19.3944
R9449 gnd.n6981 gnd.n383 19.3944
R9450 gnd.n6981 gnd.n367 19.3944
R9451 gnd.n6993 gnd.n367 19.3944
R9452 gnd.n6993 gnd.n365 19.3944
R9453 gnd.n6997 gnd.n365 19.3944
R9454 gnd.n6997 gnd.n350 19.3944
R9455 gnd.n7009 gnd.n350 19.3944
R9456 gnd.n7009 gnd.n348 19.3944
R9457 gnd.n7013 gnd.n348 19.3944
R9458 gnd.n7013 gnd.n332 19.3944
R9459 gnd.n7025 gnd.n332 19.3944
R9460 gnd.n7025 gnd.n330 19.3944
R9461 gnd.n7029 gnd.n330 19.3944
R9462 gnd.n7029 gnd.n315 19.3944
R9463 gnd.n7041 gnd.n315 19.3944
R9464 gnd.n7041 gnd.n312 19.3944
R9465 gnd.n7046 gnd.n312 19.3944
R9466 gnd.n7046 gnd.n313 19.3944
R9467 gnd.n313 gnd.n295 19.3944
R9468 gnd.n7060 gnd.n295 19.3944
R9469 gnd.n7060 gnd.n293 19.3944
R9470 gnd.n7064 gnd.n293 19.3944
R9471 gnd.n7064 gnd.n279 19.3944
R9472 gnd.n7076 gnd.n279 19.3944
R9473 gnd.n7076 gnd.n276 19.3944
R9474 gnd.n7081 gnd.n276 19.3944
R9475 gnd.n7081 gnd.n264 19.3944
R9476 gnd.n7092 gnd.n264 19.3944
R9477 gnd.n7092 gnd.n262 19.3944
R9478 gnd.n7096 gnd.n262 19.3944
R9479 gnd.n7096 gnd.n247 19.3944
R9480 gnd.n7108 gnd.n247 19.3944
R9481 gnd.n7108 gnd.n245 19.3944
R9482 gnd.n7112 gnd.n245 19.3944
R9483 gnd.n7112 gnd.n231 19.3944
R9484 gnd.n7124 gnd.n231 19.3944
R9485 gnd.n7124 gnd.n229 19.3944
R9486 gnd.n7128 gnd.n229 19.3944
R9487 gnd.n7128 gnd.n215 19.3944
R9488 gnd.n7140 gnd.n215 19.3944
R9489 gnd.n7140 gnd.n213 19.3944
R9490 gnd.n7144 gnd.n213 19.3944
R9491 gnd.n7144 gnd.n201 19.3944
R9492 gnd.n7156 gnd.n201 19.3944
R9493 gnd.n7156 gnd.n199 19.3944
R9494 gnd.n7160 gnd.n199 19.3944
R9495 gnd.n7160 gnd.n184 19.3944
R9496 gnd.n7174 gnd.n184 19.3944
R9497 gnd.n7174 gnd.n181 19.3944
R9498 gnd.n7246 gnd.n181 19.3944
R9499 gnd.n7246 gnd.n182 19.3944
R9500 gnd.n4608 gnd.n4607 19.3944
R9501 gnd.n4607 gnd.n4606 19.3944
R9502 gnd.n4606 gnd.n2205 19.3944
R9503 gnd.n4599 gnd.n2205 19.3944
R9504 gnd.n4599 gnd.n4598 19.3944
R9505 gnd.n4598 gnd.n2217 19.3944
R9506 gnd.n4591 gnd.n2217 19.3944
R9507 gnd.n4591 gnd.n4590 19.3944
R9508 gnd.n4590 gnd.n2228 19.3944
R9509 gnd.n4583 gnd.n2228 19.3944
R9510 gnd.n4583 gnd.n4582 19.3944
R9511 gnd.n4582 gnd.n2238 19.3944
R9512 gnd.n4575 gnd.n2238 19.3944
R9513 gnd.n4575 gnd.n4574 19.3944
R9514 gnd.n4574 gnd.n2249 19.3944
R9515 gnd.n4567 gnd.n2249 19.3944
R9516 gnd.n6615 gnd.n687 19.3944
R9517 gnd.n6615 gnd.n683 19.3944
R9518 gnd.n6621 gnd.n683 19.3944
R9519 gnd.n6621 gnd.n681 19.3944
R9520 gnd.n6625 gnd.n681 19.3944
R9521 gnd.n6625 gnd.n677 19.3944
R9522 gnd.n6631 gnd.n677 19.3944
R9523 gnd.n6631 gnd.n675 19.3944
R9524 gnd.n6635 gnd.n675 19.3944
R9525 gnd.n6635 gnd.n671 19.3944
R9526 gnd.n6641 gnd.n671 19.3944
R9527 gnd.n6641 gnd.n669 19.3944
R9528 gnd.n6645 gnd.n669 19.3944
R9529 gnd.n6645 gnd.n665 19.3944
R9530 gnd.n6651 gnd.n665 19.3944
R9531 gnd.n6651 gnd.n663 19.3944
R9532 gnd.n6655 gnd.n663 19.3944
R9533 gnd.n6655 gnd.n659 19.3944
R9534 gnd.n6661 gnd.n659 19.3944
R9535 gnd.n6661 gnd.n657 19.3944
R9536 gnd.n6665 gnd.n657 19.3944
R9537 gnd.n6665 gnd.n653 19.3944
R9538 gnd.n6671 gnd.n653 19.3944
R9539 gnd.n6671 gnd.n651 19.3944
R9540 gnd.n6675 gnd.n651 19.3944
R9541 gnd.n6675 gnd.n647 19.3944
R9542 gnd.n6681 gnd.n647 19.3944
R9543 gnd.n6681 gnd.n645 19.3944
R9544 gnd.n6685 gnd.n645 19.3944
R9545 gnd.n6685 gnd.n641 19.3944
R9546 gnd.n6691 gnd.n641 19.3944
R9547 gnd.n6691 gnd.n639 19.3944
R9548 gnd.n6695 gnd.n639 19.3944
R9549 gnd.n6695 gnd.n635 19.3944
R9550 gnd.n6701 gnd.n635 19.3944
R9551 gnd.n6701 gnd.n633 19.3944
R9552 gnd.n6705 gnd.n633 19.3944
R9553 gnd.n6705 gnd.n629 19.3944
R9554 gnd.n6711 gnd.n629 19.3944
R9555 gnd.n6711 gnd.n627 19.3944
R9556 gnd.n6715 gnd.n627 19.3944
R9557 gnd.n6715 gnd.n623 19.3944
R9558 gnd.n6721 gnd.n623 19.3944
R9559 gnd.n6721 gnd.n621 19.3944
R9560 gnd.n6725 gnd.n621 19.3944
R9561 gnd.n6725 gnd.n617 19.3944
R9562 gnd.n6731 gnd.n617 19.3944
R9563 gnd.n6731 gnd.n615 19.3944
R9564 gnd.n6735 gnd.n615 19.3944
R9565 gnd.n6735 gnd.n611 19.3944
R9566 gnd.n6741 gnd.n611 19.3944
R9567 gnd.n6741 gnd.n609 19.3944
R9568 gnd.n6745 gnd.n609 19.3944
R9569 gnd.n6745 gnd.n605 19.3944
R9570 gnd.n6751 gnd.n605 19.3944
R9571 gnd.n6751 gnd.n603 19.3944
R9572 gnd.n6755 gnd.n603 19.3944
R9573 gnd.n6755 gnd.n599 19.3944
R9574 gnd.n6761 gnd.n599 19.3944
R9575 gnd.n6761 gnd.n597 19.3944
R9576 gnd.n6765 gnd.n597 19.3944
R9577 gnd.n6765 gnd.n593 19.3944
R9578 gnd.n6771 gnd.n593 19.3944
R9579 gnd.n6771 gnd.n591 19.3944
R9580 gnd.n6775 gnd.n591 19.3944
R9581 gnd.n6775 gnd.n587 19.3944
R9582 gnd.n6781 gnd.n587 19.3944
R9583 gnd.n6781 gnd.n585 19.3944
R9584 gnd.n6785 gnd.n585 19.3944
R9585 gnd.n6785 gnd.n581 19.3944
R9586 gnd.n6791 gnd.n581 19.3944
R9587 gnd.n6791 gnd.n579 19.3944
R9588 gnd.n6795 gnd.n579 19.3944
R9589 gnd.n6795 gnd.n575 19.3944
R9590 gnd.n6801 gnd.n575 19.3944
R9591 gnd.n6801 gnd.n573 19.3944
R9592 gnd.n6805 gnd.n573 19.3944
R9593 gnd.n6805 gnd.n569 19.3944
R9594 gnd.n6811 gnd.n569 19.3944
R9595 gnd.n6811 gnd.n567 19.3944
R9596 gnd.n6817 gnd.n567 19.3944
R9597 gnd.n6817 gnd.n6816 19.3944
R9598 gnd.n6816 gnd.n563 19.3944
R9599 gnd.n6824 gnd.n563 19.3944
R9600 gnd.n6195 gnd.n939 19.3944
R9601 gnd.n6195 gnd.n935 19.3944
R9602 gnd.n6201 gnd.n935 19.3944
R9603 gnd.n6201 gnd.n933 19.3944
R9604 gnd.n6205 gnd.n933 19.3944
R9605 gnd.n6205 gnd.n929 19.3944
R9606 gnd.n6211 gnd.n929 19.3944
R9607 gnd.n6211 gnd.n927 19.3944
R9608 gnd.n6215 gnd.n927 19.3944
R9609 gnd.n6215 gnd.n923 19.3944
R9610 gnd.n6221 gnd.n923 19.3944
R9611 gnd.n6221 gnd.n921 19.3944
R9612 gnd.n6225 gnd.n921 19.3944
R9613 gnd.n6225 gnd.n917 19.3944
R9614 gnd.n6231 gnd.n917 19.3944
R9615 gnd.n6231 gnd.n915 19.3944
R9616 gnd.n6235 gnd.n915 19.3944
R9617 gnd.n6235 gnd.n911 19.3944
R9618 gnd.n6241 gnd.n911 19.3944
R9619 gnd.n6241 gnd.n909 19.3944
R9620 gnd.n6245 gnd.n909 19.3944
R9621 gnd.n6245 gnd.n905 19.3944
R9622 gnd.n6251 gnd.n905 19.3944
R9623 gnd.n6251 gnd.n903 19.3944
R9624 gnd.n6255 gnd.n903 19.3944
R9625 gnd.n6255 gnd.n899 19.3944
R9626 gnd.n6261 gnd.n899 19.3944
R9627 gnd.n6261 gnd.n897 19.3944
R9628 gnd.n6265 gnd.n897 19.3944
R9629 gnd.n6265 gnd.n893 19.3944
R9630 gnd.n6271 gnd.n893 19.3944
R9631 gnd.n6271 gnd.n891 19.3944
R9632 gnd.n6275 gnd.n891 19.3944
R9633 gnd.n6275 gnd.n887 19.3944
R9634 gnd.n6281 gnd.n887 19.3944
R9635 gnd.n6281 gnd.n885 19.3944
R9636 gnd.n6285 gnd.n885 19.3944
R9637 gnd.n6285 gnd.n881 19.3944
R9638 gnd.n6291 gnd.n881 19.3944
R9639 gnd.n6291 gnd.n879 19.3944
R9640 gnd.n6295 gnd.n879 19.3944
R9641 gnd.n6295 gnd.n875 19.3944
R9642 gnd.n6301 gnd.n875 19.3944
R9643 gnd.n6301 gnd.n873 19.3944
R9644 gnd.n6305 gnd.n873 19.3944
R9645 gnd.n6305 gnd.n869 19.3944
R9646 gnd.n6311 gnd.n869 19.3944
R9647 gnd.n6311 gnd.n867 19.3944
R9648 gnd.n6315 gnd.n867 19.3944
R9649 gnd.n6315 gnd.n863 19.3944
R9650 gnd.n6321 gnd.n863 19.3944
R9651 gnd.n6321 gnd.n861 19.3944
R9652 gnd.n6325 gnd.n861 19.3944
R9653 gnd.n6325 gnd.n857 19.3944
R9654 gnd.n6331 gnd.n857 19.3944
R9655 gnd.n6331 gnd.n855 19.3944
R9656 gnd.n6335 gnd.n855 19.3944
R9657 gnd.n6335 gnd.n851 19.3944
R9658 gnd.n6341 gnd.n851 19.3944
R9659 gnd.n6341 gnd.n849 19.3944
R9660 gnd.n6345 gnd.n849 19.3944
R9661 gnd.n6345 gnd.n845 19.3944
R9662 gnd.n6351 gnd.n845 19.3944
R9663 gnd.n6351 gnd.n843 19.3944
R9664 gnd.n6355 gnd.n843 19.3944
R9665 gnd.n6355 gnd.n839 19.3944
R9666 gnd.n6361 gnd.n839 19.3944
R9667 gnd.n6361 gnd.n837 19.3944
R9668 gnd.n6365 gnd.n837 19.3944
R9669 gnd.n6365 gnd.n833 19.3944
R9670 gnd.n6371 gnd.n833 19.3944
R9671 gnd.n6371 gnd.n831 19.3944
R9672 gnd.n6375 gnd.n831 19.3944
R9673 gnd.n6375 gnd.n827 19.3944
R9674 gnd.n6381 gnd.n827 19.3944
R9675 gnd.n6381 gnd.n825 19.3944
R9676 gnd.n6385 gnd.n825 19.3944
R9677 gnd.n6385 gnd.n821 19.3944
R9678 gnd.n6391 gnd.n821 19.3944
R9679 gnd.n6391 gnd.n819 19.3944
R9680 gnd.n6395 gnd.n819 19.3944
R9681 gnd.n6395 gnd.n815 19.3944
R9682 gnd.n6401 gnd.n815 19.3944
R9683 gnd.n6401 gnd.n813 19.3944
R9684 gnd.n6405 gnd.n813 19.3944
R9685 gnd.n6405 gnd.n809 19.3944
R9686 gnd.n6411 gnd.n809 19.3944
R9687 gnd.n6411 gnd.n807 19.3944
R9688 gnd.n6415 gnd.n807 19.3944
R9689 gnd.n6415 gnd.n803 19.3944
R9690 gnd.n6421 gnd.n803 19.3944
R9691 gnd.n6421 gnd.n801 19.3944
R9692 gnd.n6425 gnd.n801 19.3944
R9693 gnd.n6425 gnd.n797 19.3944
R9694 gnd.n6431 gnd.n797 19.3944
R9695 gnd.n6431 gnd.n795 19.3944
R9696 gnd.n6435 gnd.n795 19.3944
R9697 gnd.n6435 gnd.n791 19.3944
R9698 gnd.n6441 gnd.n791 19.3944
R9699 gnd.n6441 gnd.n789 19.3944
R9700 gnd.n6445 gnd.n789 19.3944
R9701 gnd.n6445 gnd.n785 19.3944
R9702 gnd.n6451 gnd.n785 19.3944
R9703 gnd.n6451 gnd.n783 19.3944
R9704 gnd.n6455 gnd.n783 19.3944
R9705 gnd.n6455 gnd.n779 19.3944
R9706 gnd.n6461 gnd.n779 19.3944
R9707 gnd.n6461 gnd.n777 19.3944
R9708 gnd.n6465 gnd.n777 19.3944
R9709 gnd.n6465 gnd.n773 19.3944
R9710 gnd.n6471 gnd.n773 19.3944
R9711 gnd.n6471 gnd.n771 19.3944
R9712 gnd.n6475 gnd.n771 19.3944
R9713 gnd.n6475 gnd.n767 19.3944
R9714 gnd.n6481 gnd.n767 19.3944
R9715 gnd.n6481 gnd.n765 19.3944
R9716 gnd.n6485 gnd.n765 19.3944
R9717 gnd.n6485 gnd.n761 19.3944
R9718 gnd.n6491 gnd.n761 19.3944
R9719 gnd.n6491 gnd.n759 19.3944
R9720 gnd.n6495 gnd.n759 19.3944
R9721 gnd.n6495 gnd.n755 19.3944
R9722 gnd.n6501 gnd.n755 19.3944
R9723 gnd.n6501 gnd.n753 19.3944
R9724 gnd.n6505 gnd.n753 19.3944
R9725 gnd.n6505 gnd.n749 19.3944
R9726 gnd.n6511 gnd.n749 19.3944
R9727 gnd.n6511 gnd.n747 19.3944
R9728 gnd.n6515 gnd.n747 19.3944
R9729 gnd.n6515 gnd.n743 19.3944
R9730 gnd.n6521 gnd.n743 19.3944
R9731 gnd.n6521 gnd.n741 19.3944
R9732 gnd.n6525 gnd.n741 19.3944
R9733 gnd.n6525 gnd.n737 19.3944
R9734 gnd.n6531 gnd.n737 19.3944
R9735 gnd.n6531 gnd.n735 19.3944
R9736 gnd.n6535 gnd.n735 19.3944
R9737 gnd.n6535 gnd.n731 19.3944
R9738 gnd.n6541 gnd.n731 19.3944
R9739 gnd.n6541 gnd.n729 19.3944
R9740 gnd.n6545 gnd.n729 19.3944
R9741 gnd.n6545 gnd.n725 19.3944
R9742 gnd.n6551 gnd.n725 19.3944
R9743 gnd.n6551 gnd.n723 19.3944
R9744 gnd.n6555 gnd.n723 19.3944
R9745 gnd.n6555 gnd.n719 19.3944
R9746 gnd.n6561 gnd.n719 19.3944
R9747 gnd.n6561 gnd.n717 19.3944
R9748 gnd.n6565 gnd.n717 19.3944
R9749 gnd.n6565 gnd.n713 19.3944
R9750 gnd.n6571 gnd.n713 19.3944
R9751 gnd.n6571 gnd.n711 19.3944
R9752 gnd.n6575 gnd.n711 19.3944
R9753 gnd.n6575 gnd.n707 19.3944
R9754 gnd.n6581 gnd.n707 19.3944
R9755 gnd.n6581 gnd.n705 19.3944
R9756 gnd.n6585 gnd.n705 19.3944
R9757 gnd.n6585 gnd.n701 19.3944
R9758 gnd.n6591 gnd.n701 19.3944
R9759 gnd.n6591 gnd.n699 19.3944
R9760 gnd.n6595 gnd.n699 19.3944
R9761 gnd.n6595 gnd.n695 19.3944
R9762 gnd.n6601 gnd.n695 19.3944
R9763 gnd.n6601 gnd.n693 19.3944
R9764 gnd.n6605 gnd.n693 19.3944
R9765 gnd.n6605 gnd.n689 19.3944
R9766 gnd.n6611 gnd.n689 19.3944
R9767 gnd.n6969 gnd.n393 19.3944
R9768 gnd.n6964 gnd.n393 19.3944
R9769 gnd.n6964 gnd.n6963 19.3944
R9770 gnd.n6963 gnd.n6962 19.3944
R9771 gnd.n6962 gnd.n6959 19.3944
R9772 gnd.n6959 gnd.n6958 19.3944
R9773 gnd.n6958 gnd.n6955 19.3944
R9774 gnd.n6955 gnd.n6954 19.3944
R9775 gnd.n6954 gnd.n6951 19.3944
R9776 gnd.n6951 gnd.n6950 19.3944
R9777 gnd.n6950 gnd.n6947 19.3944
R9778 gnd.n6947 gnd.n6946 19.3944
R9779 gnd.n6946 gnd.n6943 19.3944
R9780 gnd.n6943 gnd.n6942 19.3944
R9781 gnd.n6942 gnd.n6939 19.3944
R9782 gnd.n6937 gnd.n6934 19.3944
R9783 gnd.n6934 gnd.n6933 19.3944
R9784 gnd.n6933 gnd.n6930 19.3944
R9785 gnd.n6930 gnd.n6929 19.3944
R9786 gnd.n6929 gnd.n6926 19.3944
R9787 gnd.n6926 gnd.n6925 19.3944
R9788 gnd.n6925 gnd.n6922 19.3944
R9789 gnd.n6922 gnd.n6921 19.3944
R9790 gnd.n6921 gnd.n6918 19.3944
R9791 gnd.n6918 gnd.n6917 19.3944
R9792 gnd.n6917 gnd.n6914 19.3944
R9793 gnd.n6914 gnd.n6913 19.3944
R9794 gnd.n6913 gnd.n6910 19.3944
R9795 gnd.n6910 gnd.n6909 19.3944
R9796 gnd.n6909 gnd.n6906 19.3944
R9797 gnd.n6906 gnd.n6905 19.3944
R9798 gnd.n6905 gnd.n6902 19.3944
R9799 gnd.n6902 gnd.n6901 19.3944
R9800 gnd.n5464 gnd.n469 19.3944
R9801 gnd.n5614 gnd.n5464 19.3944
R9802 gnd.n5614 gnd.n5613 19.3944
R9803 gnd.n5613 gnd.n5612 19.3944
R9804 gnd.n5612 gnd.n5609 19.3944
R9805 gnd.n5609 gnd.n5608 19.3944
R9806 gnd.n5608 gnd.n5605 19.3944
R9807 gnd.n5605 gnd.n5604 19.3944
R9808 gnd.n5604 gnd.n5601 19.3944
R9809 gnd.n5601 gnd.n5600 19.3944
R9810 gnd.n5600 gnd.n5475 19.3944
R9811 gnd.n5514 gnd.n5475 19.3944
R9812 gnd.n5514 gnd.n5510 19.3944
R9813 gnd.n5520 gnd.n5510 19.3944
R9814 gnd.n5521 gnd.n5520 19.3944
R9815 gnd.n5524 gnd.n5521 19.3944
R9816 gnd.n5524 gnd.n5508 19.3944
R9817 gnd.n5580 gnd.n5508 19.3944
R9818 gnd.n5580 gnd.n5579 19.3944
R9819 gnd.n5579 gnd.n5578 19.3944
R9820 gnd.n5578 gnd.n5530 19.3944
R9821 gnd.n5547 gnd.n5530 19.3944
R9822 gnd.n5552 gnd.n5547 19.3944
R9823 gnd.n5552 gnd.n495 19.3944
R9824 gnd.n6849 gnd.n495 19.3944
R9825 gnd.n6849 gnd.n6848 19.3944
R9826 gnd.n6848 gnd.n6847 19.3944
R9827 gnd.n6847 gnd.n6844 19.3944
R9828 gnd.n6844 gnd.n6843 19.3944
R9829 gnd.n6843 gnd.n6840 19.3944
R9830 gnd.n6840 gnd.n6839 19.3944
R9831 gnd.n6839 gnd.n552 19.3944
R9832 gnd.n552 gnd.n551 19.3944
R9833 gnd.n551 gnd.n548 19.3944
R9834 gnd.n548 gnd.n547 19.3944
R9835 gnd.n547 gnd.n544 19.3944
R9836 gnd.n544 gnd.n543 19.3944
R9837 gnd.n543 gnd.n541 19.3944
R9838 gnd.n541 gnd.n540 19.3944
R9839 gnd.n540 gnd.n538 19.3944
R9840 gnd.n538 gnd.n537 19.3944
R9841 gnd.n537 gnd.n535 19.3944
R9842 gnd.n535 gnd.n534 19.3944
R9843 gnd.n534 gnd.n532 19.3944
R9844 gnd.n532 gnd.n531 19.3944
R9845 gnd.n531 gnd.n529 19.3944
R9846 gnd.n529 gnd.n528 19.3944
R9847 gnd.n528 gnd.n526 19.3944
R9848 gnd.n526 gnd.n525 19.3944
R9849 gnd.n525 gnd.n523 19.3944
R9850 gnd.n523 gnd.n178 19.3944
R9851 gnd.n7250 gnd.n178 19.3944
R9852 gnd.n7251 gnd.n7250 19.3944
R9853 gnd.n7289 gnd.n139 19.3944
R9854 gnd.n7284 gnd.n139 19.3944
R9855 gnd.n7284 gnd.n7283 19.3944
R9856 gnd.n7283 gnd.n7282 19.3944
R9857 gnd.n7282 gnd.n146 19.3944
R9858 gnd.n7277 gnd.n146 19.3944
R9859 gnd.n7277 gnd.n7276 19.3944
R9860 gnd.n7276 gnd.n7275 19.3944
R9861 gnd.n7275 gnd.n153 19.3944
R9862 gnd.n7270 gnd.n153 19.3944
R9863 gnd.n7270 gnd.n7269 19.3944
R9864 gnd.n7269 gnd.n7268 19.3944
R9865 gnd.n7268 gnd.n160 19.3944
R9866 gnd.n7263 gnd.n160 19.3944
R9867 gnd.n7263 gnd.n7262 19.3944
R9868 gnd.n7262 gnd.n7261 19.3944
R9869 gnd.n7261 gnd.n167 19.3944
R9870 gnd.n7256 gnd.n167 19.3944
R9871 gnd.n7322 gnd.n7321 19.3944
R9872 gnd.n7321 gnd.n7320 19.3944
R9873 gnd.n7320 gnd.n111 19.3944
R9874 gnd.n7315 gnd.n111 19.3944
R9875 gnd.n7315 gnd.n7314 19.3944
R9876 gnd.n7314 gnd.n7313 19.3944
R9877 gnd.n7313 gnd.n118 19.3944
R9878 gnd.n7308 gnd.n118 19.3944
R9879 gnd.n7308 gnd.n7307 19.3944
R9880 gnd.n7307 gnd.n7306 19.3944
R9881 gnd.n7306 gnd.n125 19.3944
R9882 gnd.n7301 gnd.n125 19.3944
R9883 gnd.n7301 gnd.n7300 19.3944
R9884 gnd.n7300 gnd.n7299 19.3944
R9885 gnd.n7299 gnd.n132 19.3944
R9886 gnd.n7294 gnd.n132 19.3944
R9887 gnd.n7294 gnd.n7293 19.3944
R9888 gnd.n6973 gnd.n391 19.3944
R9889 gnd.n6973 gnd.n376 19.3944
R9890 gnd.n6985 gnd.n376 19.3944
R9891 gnd.n6985 gnd.n374 19.3944
R9892 gnd.n6989 gnd.n374 19.3944
R9893 gnd.n6989 gnd.n358 19.3944
R9894 gnd.n7001 gnd.n358 19.3944
R9895 gnd.n7001 gnd.n356 19.3944
R9896 gnd.n7005 gnd.n356 19.3944
R9897 gnd.n7005 gnd.n341 19.3944
R9898 gnd.n7017 gnd.n341 19.3944
R9899 gnd.n7017 gnd.n339 19.3944
R9900 gnd.n7021 gnd.n339 19.3944
R9901 gnd.n7021 gnd.n323 19.3944
R9902 gnd.n7033 gnd.n323 19.3944
R9903 gnd.n7033 gnd.n321 19.3944
R9904 gnd.n7037 gnd.n321 19.3944
R9905 gnd.n7037 gnd.n303 19.3944
R9906 gnd.n7050 gnd.n303 19.3944
R9907 gnd.n7050 gnd.n301 19.3944
R9908 gnd.n7054 gnd.n301 19.3944
R9909 gnd.n7056 gnd.n7054 19.3944
R9910 gnd.n7068 gnd.n286 19.3944
R9911 gnd.n7069 gnd.n7068 19.3944
R9912 gnd.n7072 gnd.n7071 19.3944
R9913 gnd.n7086 gnd.n7085 19.3944
R9914 gnd.n7088 gnd.n256 19.3944
R9915 gnd.n7100 gnd.n256 19.3944
R9916 gnd.n7100 gnd.n254 19.3944
R9917 gnd.n7104 gnd.n254 19.3944
R9918 gnd.n7104 gnd.n239 19.3944
R9919 gnd.n7116 gnd.n239 19.3944
R9920 gnd.n7116 gnd.n237 19.3944
R9921 gnd.n7120 gnd.n237 19.3944
R9922 gnd.n7120 gnd.n223 19.3944
R9923 gnd.n7132 gnd.n223 19.3944
R9924 gnd.n7132 gnd.n221 19.3944
R9925 gnd.n7136 gnd.n221 19.3944
R9926 gnd.n7136 gnd.n209 19.3944
R9927 gnd.n7148 gnd.n209 19.3944
R9928 gnd.n7148 gnd.n207 19.3944
R9929 gnd.n7152 gnd.n207 19.3944
R9930 gnd.n7152 gnd.n194 19.3944
R9931 gnd.n7164 gnd.n194 19.3944
R9932 gnd.n7164 gnd.n192 19.3944
R9933 gnd.n7170 gnd.n192 19.3944
R9934 gnd.n7170 gnd.n7169 19.3944
R9935 gnd.n7169 gnd.n106 19.3944
R9936 gnd.n7325 gnd.n106 19.3944
R9937 gnd.n2387 gnd.n2386 19.3944
R9938 gnd.n4333 gnd.n2387 19.3944
R9939 gnd.n4333 gnd.n2383 19.3944
R9940 gnd.n4337 gnd.n2383 19.3944
R9941 gnd.n4341 gnd.n4337 19.3944
R9942 gnd.n4339 gnd.n4338 19.3944
R9943 gnd.n4366 gnd.n4365 19.3944
R9944 gnd.n4371 gnd.n4370 19.3944
R9945 gnd.n4368 gnd.n2332 19.3944
R9946 gnd.n4435 gnd.n2329 19.3944
R9947 gnd.n4435 gnd.n2328 19.3944
R9948 gnd.n4439 gnd.n2328 19.3944
R9949 gnd.n4439 gnd.n2326 19.3944
R9950 gnd.n4443 gnd.n2326 19.3944
R9951 gnd.n4443 gnd.n2324 19.3944
R9952 gnd.n4467 gnd.n2324 19.3944
R9953 gnd.n4467 gnd.n4466 19.3944
R9954 gnd.n4466 gnd.n4465 19.3944
R9955 gnd.n4465 gnd.n4449 19.3944
R9956 gnd.n4461 gnd.n4449 19.3944
R9957 gnd.n4461 gnd.n4460 19.3944
R9958 gnd.n4460 gnd.n4459 19.3944
R9959 gnd.n4459 gnd.n4457 19.3944
R9960 gnd.n4457 gnd.n2299 19.3944
R9961 gnd.n2299 gnd.n2297 19.3944
R9962 gnd.n4527 gnd.n2297 19.3944
R9963 gnd.n4527 gnd.n2295 19.3944
R9964 gnd.n4531 gnd.n2295 19.3944
R9965 gnd.n4531 gnd.n2293 19.3944
R9966 gnd.n4535 gnd.n2293 19.3944
R9967 gnd.n4535 gnd.n2291 19.3944
R9968 gnd.n4539 gnd.n2291 19.3944
R9969 gnd.n4539 gnd.n2289 19.3944
R9970 gnd.n4546 gnd.n2289 19.3944
R9971 gnd.n4546 gnd.n2287 19.3944
R9972 gnd.n4552 gnd.n2287 19.3944
R9973 gnd.n4552 gnd.n4551 19.3944
R9974 gnd.n4551 gnd.n2196 19.3944
R9975 gnd.n4619 gnd.n2196 19.3944
R9976 gnd.n4619 gnd.n2194 19.3944
R9977 gnd.n4623 gnd.n2194 19.3944
R9978 gnd.n4623 gnd.n2182 19.3944
R9979 gnd.n4638 gnd.n2182 19.3944
R9980 gnd.n4638 gnd.n2180 19.3944
R9981 gnd.n4642 gnd.n2180 19.3944
R9982 gnd.n4642 gnd.n2168 19.3944
R9983 gnd.n4658 gnd.n2168 19.3944
R9984 gnd.n4658 gnd.n2166 19.3944
R9985 gnd.n4668 gnd.n2166 19.3944
R9986 gnd.n4668 gnd.n4667 19.3944
R9987 gnd.n4667 gnd.n4666 19.3944
R9988 gnd.n4666 gnd.n1945 19.3944
R9989 gnd.n4710 gnd.n1945 19.3944
R9990 gnd.n4710 gnd.n1943 19.3944
R9991 gnd.n4719 gnd.n1943 19.3944
R9992 gnd.n4719 gnd.n4718 19.3944
R9993 gnd.n4718 gnd.n4717 19.3944
R9994 gnd.n4717 gnd.n1909 19.3944
R9995 gnd.n4793 gnd.n1909 19.3944
R9996 gnd.n4793 gnd.n1907 19.3944
R9997 gnd.n4797 gnd.n1907 19.3944
R9998 gnd.n4797 gnd.n1886 19.3944
R9999 gnd.n4820 gnd.n1886 19.3944
R10000 gnd.n4820 gnd.n1884 19.3944
R10001 gnd.n4826 gnd.n1884 19.3944
R10002 gnd.n4826 gnd.n4825 19.3944
R10003 gnd.n4825 gnd.n1856 19.3944
R10004 gnd.n4861 gnd.n1856 19.3944
R10005 gnd.n4861 gnd.n1854 19.3944
R10006 gnd.n4865 gnd.n1854 19.3944
R10007 gnd.n4865 gnd.n1832 19.3944
R10008 gnd.n4904 gnd.n1832 19.3944
R10009 gnd.n4904 gnd.n1830 19.3944
R10010 gnd.n4908 gnd.n1830 19.3944
R10011 gnd.n4908 gnd.n1816 19.3944
R10012 gnd.n5019 gnd.n1816 19.3944
R10013 gnd.n5019 gnd.n1814 19.3944
R10014 gnd.n5023 gnd.n1814 19.3944
R10015 gnd.n5023 gnd.n1793 19.3944
R10016 gnd.n5046 gnd.n1793 19.3944
R10017 gnd.n5046 gnd.n1791 19.3944
R10018 gnd.n5052 gnd.n1791 19.3944
R10019 gnd.n5052 gnd.n5051 19.3944
R10020 gnd.n5051 gnd.n1764 19.3944
R10021 gnd.n5082 gnd.n1764 19.3944
R10022 gnd.n5082 gnd.n1762 19.3944
R10023 gnd.n5086 gnd.n1762 19.3944
R10024 gnd.n5086 gnd.n1742 19.3944
R10025 gnd.n5112 gnd.n1742 19.3944
R10026 gnd.n5112 gnd.n1740 19.3944
R10027 gnd.n5116 gnd.n1740 19.3944
R10028 gnd.n5116 gnd.n1720 19.3944
R10029 gnd.n5142 gnd.n1720 19.3944
R10030 gnd.n5142 gnd.n1718 19.3944
R10031 gnd.n5146 gnd.n1718 19.3944
R10032 gnd.n5146 gnd.n1698 19.3944
R10033 gnd.n5169 gnd.n1698 19.3944
R10034 gnd.n5169 gnd.n1696 19.3944
R10035 gnd.n5175 gnd.n1696 19.3944
R10036 gnd.n5175 gnd.n5174 19.3944
R10037 gnd.n5174 gnd.n1671 19.3944
R10038 gnd.n5206 gnd.n1671 19.3944
R10039 gnd.n5206 gnd.n1669 19.3944
R10040 gnd.n5221 gnd.n1669 19.3944
R10041 gnd.n5221 gnd.n5220 19.3944
R10042 gnd.n5220 gnd.n5219 19.3944
R10043 gnd.n5219 gnd.n5212 19.3944
R10044 gnd.n5215 gnd.n5212 19.3944
R10045 gnd.n5215 gnd.n1599 19.3944
R10046 gnd.n5407 gnd.n1599 19.3944
R10047 gnd.n5407 gnd.n1597 19.3944
R10048 gnd.n5411 gnd.n1597 19.3944
R10049 gnd.n5411 gnd.n1585 19.3944
R10050 gnd.n5426 gnd.n1585 19.3944
R10051 gnd.n5426 gnd.n1583 19.3944
R10052 gnd.n5433 gnd.n1583 19.3944
R10053 gnd.n5433 gnd.n5432 19.3944
R10054 gnd.n5432 gnd.n1572 19.3944
R10055 gnd.n1572 gnd.n1570 19.3944
R10056 gnd.n5450 gnd.n1570 19.3944
R10057 gnd.n5450 gnd.n1568 19.3944
R10058 gnd.n5627 gnd.n1568 19.3944
R10059 gnd.n5627 gnd.n5626 19.3944
R10060 gnd.n5626 gnd.n5625 19.3944
R10061 gnd.n5625 gnd.n5456 19.3944
R10062 gnd.n5621 gnd.n5456 19.3944
R10063 gnd.n5621 gnd.n5620 19.3944
R10064 gnd.n5620 gnd.n5619 19.3944
R10065 gnd.n5619 gnd.n5462 19.3944
R10066 gnd.n5485 gnd.n5462 19.3944
R10067 gnd.n5485 gnd.n5482 19.3944
R10068 gnd.n5489 gnd.n5482 19.3944
R10069 gnd.n5489 gnd.n5480 19.3944
R10070 gnd.n5493 gnd.n5480 19.3944
R10071 gnd.n5493 gnd.n5478 19.3944
R10072 gnd.n5595 gnd.n5478 19.3944
R10073 gnd.n5595 gnd.n5594 19.3944
R10074 gnd.n5594 gnd.n5593 19.3944
R10075 gnd.n5593 gnd.n5499 19.3944
R10076 gnd.n5589 gnd.n5499 19.3944
R10077 gnd.n5589 gnd.n5588 19.3944
R10078 gnd.n5588 gnd.n5587 19.3944
R10079 gnd.n5587 gnd.n5505 19.3944
R10080 gnd.n5507 gnd.n5505 19.3944
R10081 gnd.n5539 gnd.n5507 19.3944
R10082 gnd.n5539 gnd.n5536 19.3944
R10083 gnd.n5573 gnd.n5536 19.3944
R10084 gnd.n5573 gnd.n5572 19.3944
R10085 gnd.n5568 gnd.n5543 19.3944
R10086 gnd.n5564 gnd.n5546 19.3944
R10087 gnd.n5562 gnd.n5561 19.3944
R10088 gnd.n5558 gnd.n5557 19.3944
R10089 gnd.n6834 gnd.n6833 19.3944
R10090 gnd.n6833 gnd.n6832 19.3944
R10091 gnd.n6832 gnd.n558 19.3944
R10092 gnd.n6828 gnd.n558 19.3944
R10093 gnd.n6828 gnd.n6827 19.3944
R10094 gnd.n3970 gnd.n3967 19.3944
R10095 gnd.n3970 gnd.n3966 19.3944
R10096 gnd.n3974 gnd.n3966 19.3944
R10097 gnd.n3974 gnd.n3964 19.3944
R10098 gnd.n3980 gnd.n3964 19.3944
R10099 gnd.n3980 gnd.n3962 19.3944
R10100 gnd.n3984 gnd.n3962 19.3944
R10101 gnd.n3984 gnd.n3960 19.3944
R10102 gnd.n3990 gnd.n3960 19.3944
R10103 gnd.n3990 gnd.n3958 19.3944
R10104 gnd.n3994 gnd.n3958 19.3944
R10105 gnd.n3994 gnd.n3956 19.3944
R10106 gnd.n4000 gnd.n3956 19.3944
R10107 gnd.n4000 gnd.n3954 19.3944
R10108 gnd.n4004 gnd.n3954 19.3944
R10109 gnd.n4004 gnd.n3949 19.3944
R10110 gnd.n4010 gnd.n3949 19.3944
R10111 gnd.n4014 gnd.n3947 19.3944
R10112 gnd.n4014 gnd.n3945 19.3944
R10113 gnd.n4020 gnd.n3945 19.3944
R10114 gnd.n4020 gnd.n3943 19.3944
R10115 gnd.n4024 gnd.n3943 19.3944
R10116 gnd.n4024 gnd.n3941 19.3944
R10117 gnd.n4030 gnd.n3941 19.3944
R10118 gnd.n4030 gnd.n3939 19.3944
R10119 gnd.n4034 gnd.n3939 19.3944
R10120 gnd.n4034 gnd.n3937 19.3944
R10121 gnd.n4040 gnd.n3937 19.3944
R10122 gnd.n4040 gnd.n3935 19.3944
R10123 gnd.n4044 gnd.n3935 19.3944
R10124 gnd.n4044 gnd.n3933 19.3944
R10125 gnd.n4050 gnd.n3933 19.3944
R10126 gnd.n4050 gnd.n3931 19.3944
R10127 gnd.n4055 gnd.n3931 19.3944
R10128 gnd.n4055 gnd.n3929 19.3944
R10129 gnd.n4094 gnd.n3923 19.3944
R10130 gnd.n4094 gnd.n3924 19.3944
R10131 gnd.n4090 gnd.n3924 19.3944
R10132 gnd.n4090 gnd.n4088 19.3944
R10133 gnd.n4088 gnd.n4087 19.3944
R10134 gnd.n4087 gnd.n4085 19.3944
R10135 gnd.n4085 gnd.n4084 19.3944
R10136 gnd.n4084 gnd.n4082 19.3944
R10137 gnd.n4082 gnd.n4081 19.3944
R10138 gnd.n4081 gnd.n4079 19.3944
R10139 gnd.n4079 gnd.n4078 19.3944
R10140 gnd.n4078 gnd.n4076 19.3944
R10141 gnd.n4076 gnd.n4075 19.3944
R10142 gnd.n4075 gnd.n2400 19.3944
R10143 gnd.n4284 gnd.n2400 19.3944
R10144 gnd.n4284 gnd.n2398 19.3944
R10145 gnd.n4289 gnd.n2398 19.3944
R10146 gnd.n4290 gnd.n4289 19.3944
R10147 gnd.n4291 gnd.n4290 19.3944
R10148 gnd.n4291 gnd.n2396 19.3944
R10149 gnd.n4322 gnd.n2396 19.3944
R10150 gnd.n4322 gnd.n4321 19.3944
R10151 gnd.n4321 gnd.n4320 19.3944
R10152 gnd.n4320 gnd.n4301 19.3944
R10153 gnd.n4301 gnd.n4300 19.3944
R10154 gnd.n4300 gnd.n2358 19.3944
R10155 gnd.n4376 gnd.n2358 19.3944
R10156 gnd.n4376 gnd.n2347 19.3944
R10157 gnd.n4394 gnd.n2347 19.3944
R10158 gnd.n4395 gnd.n4394 19.3944
R10159 gnd.n4395 gnd.n2345 19.3944
R10160 gnd.n4401 gnd.n2345 19.3944
R10161 gnd.n4402 gnd.n4401 19.3944
R10162 gnd.n4406 gnd.n4402 19.3944
R10163 gnd.n4406 gnd.n2343 19.3944
R10164 gnd.n4414 gnd.n2343 19.3944
R10165 gnd.n4414 gnd.n4413 19.3944
R10166 gnd.n4413 gnd.n4412 19.3944
R10167 gnd.n4412 gnd.n2317 19.3944
R10168 gnd.n4480 gnd.n2317 19.3944
R10169 gnd.n4480 gnd.n2315 19.3944
R10170 gnd.n4484 gnd.n2315 19.3944
R10171 gnd.n4484 gnd.n2310 19.3944
R10172 gnd.n4496 gnd.n2310 19.3944
R10173 gnd.n4496 gnd.n2308 19.3944
R10174 gnd.n4500 gnd.n2308 19.3944
R10175 gnd.n4501 gnd.n4500 19.3944
R10176 gnd.n4504 gnd.n4501 19.3944
R10177 gnd.n4504 gnd.n2306 19.3944
R10178 gnd.n4509 gnd.n2306 19.3944
R10179 gnd.n4509 gnd.n1343 19.3944
R10180 gnd.n5858 gnd.n1343 19.3944
R10181 gnd.n5859 gnd.n5858 19.3944
R10182 gnd.n5897 gnd.n5896 19.3944
R10183 gnd.n5896 gnd.n5895 19.3944
R10184 gnd.n5895 gnd.n1309 19.3944
R10185 gnd.n5890 gnd.n1309 19.3944
R10186 gnd.n5890 gnd.n5889 19.3944
R10187 gnd.n5889 gnd.n5888 19.3944
R10188 gnd.n5888 gnd.n1316 19.3944
R10189 gnd.n5883 gnd.n1316 19.3944
R10190 gnd.n5883 gnd.n5882 19.3944
R10191 gnd.n5882 gnd.n5881 19.3944
R10192 gnd.n5881 gnd.n1323 19.3944
R10193 gnd.n5876 gnd.n1323 19.3944
R10194 gnd.n5876 gnd.n5875 19.3944
R10195 gnd.n5875 gnd.n5874 19.3944
R10196 gnd.n5874 gnd.n1330 19.3944
R10197 gnd.n5869 gnd.n1330 19.3944
R10198 gnd.n5869 gnd.n5868 19.3944
R10199 gnd.n5868 gnd.n5867 19.3944
R10200 gnd.n5928 gnd.n5927 19.3944
R10201 gnd.n5927 gnd.n1275 19.3944
R10202 gnd.n1277 gnd.n1275 19.3944
R10203 gnd.n5920 gnd.n1277 19.3944
R10204 gnd.n5920 gnd.n5919 19.3944
R10205 gnd.n5919 gnd.n5918 19.3944
R10206 gnd.n5918 gnd.n1284 19.3944
R10207 gnd.n5913 gnd.n1284 19.3944
R10208 gnd.n5913 gnd.n5912 19.3944
R10209 gnd.n5912 gnd.n5911 19.3944
R10210 gnd.n5911 gnd.n1291 19.3944
R10211 gnd.n5906 gnd.n1291 19.3944
R10212 gnd.n5906 gnd.n5905 19.3944
R10213 gnd.n5905 gnd.n5904 19.3944
R10214 gnd.n5904 gnd.n1298 19.3944
R10215 gnd.n4212 gnd.n2449 19.3944
R10216 gnd.n4224 gnd.n2449 19.3944
R10217 gnd.n4224 gnd.n2447 19.3944
R10218 gnd.n4228 gnd.n2447 19.3944
R10219 gnd.n4228 gnd.n2433 19.3944
R10220 gnd.n4240 gnd.n2433 19.3944
R10221 gnd.n4240 gnd.n2431 19.3944
R10222 gnd.n4244 gnd.n2431 19.3944
R10223 gnd.n4244 gnd.n2416 19.3944
R10224 gnd.n4256 gnd.n2416 19.3944
R10225 gnd.n4256 gnd.n2414 19.3944
R10226 gnd.n4270 gnd.n2414 19.3944
R10227 gnd.n4270 gnd.n4269 19.3944
R10228 gnd.n4269 gnd.n4268 19.3944
R10229 gnd.n4268 gnd.n4267 19.3944
R10230 gnd.n4267 gnd.n4265 19.3944
R10231 gnd.n4265 gnd.n1128 19.3944
R10232 gnd.n6012 gnd.n1128 19.3944
R10233 gnd.n6012 gnd.n6011 19.3944
R10234 gnd.n6011 gnd.n6010 19.3944
R10235 gnd.n6010 gnd.n1132 19.3944
R10236 gnd.n4346 gnd.n1132 19.3944
R10237 gnd.n4346 gnd.n2376 19.3944
R10238 gnd.n4353 gnd.n2376 19.3944
R10239 gnd.n4353 gnd.n4352 19.3944
R10240 gnd.n4352 gnd.n4351 19.3944
R10241 gnd.n4351 gnd.n2354 19.3944
R10242 gnd.n4385 gnd.n2354 19.3944
R10243 gnd.n4385 gnd.n4384 19.3944
R10244 gnd.n4384 gnd.n1158 19.3944
R10245 gnd.n5997 gnd.n1158 19.3944
R10246 gnd.n5997 gnd.n5996 19.3944
R10247 gnd.n5996 gnd.n5995 19.3944
R10248 gnd.n5995 gnd.n1162 19.3944
R10249 gnd.n5985 gnd.n1162 19.3944
R10250 gnd.n5985 gnd.n5984 19.3944
R10251 gnd.n5984 gnd.n5983 19.3944
R10252 gnd.n5983 gnd.n1182 19.3944
R10253 gnd.n5973 gnd.n1182 19.3944
R10254 gnd.n5973 gnd.n5972 19.3944
R10255 gnd.n5972 gnd.n5971 19.3944
R10256 gnd.n5971 gnd.n1203 19.3944
R10257 gnd.n5961 gnd.n1203 19.3944
R10258 gnd.n5961 gnd.n5960 19.3944
R10259 gnd.n5960 gnd.n5959 19.3944
R10260 gnd.n5959 gnd.n1224 19.3944
R10261 gnd.n5949 gnd.n1224 19.3944
R10262 gnd.n5949 gnd.n5948 19.3944
R10263 gnd.n5948 gnd.n5947 19.3944
R10264 gnd.n5947 gnd.n1245 19.3944
R10265 gnd.n5937 gnd.n1245 19.3944
R10266 gnd.n5937 gnd.n5936 19.3944
R10267 gnd.n5936 gnd.n5935 19.3944
R10268 gnd.n4209 gnd.n4208 19.3944
R10269 gnd.n4208 gnd.n4099 19.3944
R10270 gnd.n4202 gnd.n4099 19.3944
R10271 gnd.n4202 gnd.n4201 19.3944
R10272 gnd.n4201 gnd.n4200 19.3944
R10273 gnd.n4200 gnd.n4105 19.3944
R10274 gnd.n4194 gnd.n4105 19.3944
R10275 gnd.n4194 gnd.n4193 19.3944
R10276 gnd.n4193 gnd.n4192 19.3944
R10277 gnd.n4192 gnd.n4111 19.3944
R10278 gnd.n4186 gnd.n4111 19.3944
R10279 gnd.n4186 gnd.n4185 19.3944
R10280 gnd.n4185 gnd.n4184 19.3944
R10281 gnd.n4184 gnd.n4117 19.3944
R10282 gnd.n4178 gnd.n4117 19.3944
R10283 gnd.n4178 gnd.n4177 19.3944
R10284 gnd.n4168 gnd.n4167 19.3944
R10285 gnd.n4167 gnd.n4166 19.3944
R10286 gnd.n4166 gnd.n4165 19.3944
R10287 gnd.n4165 gnd.n4163 19.3944
R10288 gnd.n4163 gnd.n4162 19.3944
R10289 gnd.n4162 gnd.n4160 19.3944
R10290 gnd.n4160 gnd.n4159 19.3944
R10291 gnd.n4159 gnd.n4157 19.3944
R10292 gnd.n4157 gnd.n4156 19.3944
R10293 gnd.n4156 gnd.n4154 19.3944
R10294 gnd.n4154 gnd.n4153 19.3944
R10295 gnd.n4153 gnd.n4151 19.3944
R10296 gnd.n4151 gnd.n4150 19.3944
R10297 gnd.n4150 gnd.n4148 19.3944
R10298 gnd.n4148 gnd.n4147 19.3944
R10299 gnd.n4147 gnd.n4145 19.3944
R10300 gnd.n4145 gnd.n4144 19.3944
R10301 gnd.n4144 gnd.n2391 19.3944
R10302 gnd.n4328 gnd.n2391 19.3944
R10303 gnd.n4328 gnd.n4327 19.3944
R10304 gnd.n4327 gnd.n4326 19.3944
R10305 gnd.n4326 gnd.n2395 19.3944
R10306 gnd.n4316 gnd.n2395 19.3944
R10307 gnd.n4316 gnd.n4315 19.3944
R10308 gnd.n4315 gnd.n4314 19.3944
R10309 gnd.n4314 gnd.n4312 19.3944
R10310 gnd.n4312 gnd.n4311 19.3944
R10311 gnd.n4311 gnd.n4307 19.3944
R10312 gnd.n4307 gnd.n2336 19.3944
R10313 gnd.n4428 gnd.n2336 19.3944
R10314 gnd.n4428 gnd.n2337 19.3944
R10315 gnd.n4424 gnd.n2337 19.3944
R10316 gnd.n4424 gnd.n4423 19.3944
R10317 gnd.n4423 gnd.n4422 19.3944
R10318 gnd.n4422 gnd.n2342 19.3944
R10319 gnd.n4418 gnd.n2342 19.3944
R10320 gnd.n4418 gnd.n2320 19.3944
R10321 gnd.n4472 gnd.n2320 19.3944
R10322 gnd.n4472 gnd.n2318 19.3944
R10323 gnd.n4476 gnd.n2318 19.3944
R10324 gnd.n4476 gnd.n2313 19.3944
R10325 gnd.n4488 gnd.n2313 19.3944
R10326 gnd.n4488 gnd.n2311 19.3944
R10327 gnd.n4492 gnd.n2311 19.3944
R10328 gnd.n4492 gnd.n2301 19.3944
R10329 gnd.n4520 gnd.n2301 19.3944
R10330 gnd.n4520 gnd.n2302 19.3944
R10331 gnd.n4516 gnd.n2302 19.3944
R10332 gnd.n4516 gnd.n4515 19.3944
R10333 gnd.n4515 gnd.n4514 19.3944
R10334 gnd.n4514 gnd.n1344 19.3944
R10335 gnd.n5854 gnd.n1344 19.3944
R10336 gnd.n5854 gnd.n1345 19.3944
R10337 gnd.n4216 gnd.n2454 19.3944
R10338 gnd.n4220 gnd.n2454 19.3944
R10339 gnd.n4220 gnd.n2441 19.3944
R10340 gnd.n4232 gnd.n2441 19.3944
R10341 gnd.n4232 gnd.n2439 19.3944
R10342 gnd.n4236 gnd.n2439 19.3944
R10343 gnd.n4236 gnd.n2424 19.3944
R10344 gnd.n4248 gnd.n2424 19.3944
R10345 gnd.n4248 gnd.n2422 19.3944
R10346 gnd.n4252 gnd.n2422 19.3944
R10347 gnd.n4252 gnd.n2408 19.3944
R10348 gnd.n4274 gnd.n2408 19.3944
R10349 gnd.n4274 gnd.n2406 19.3944
R10350 gnd.n4279 gnd.n2406 19.3944
R10351 gnd.n4279 gnd.n1116 19.3944
R10352 gnd.n6018 gnd.n1116 19.3944
R10353 gnd.n6018 gnd.n6017 19.3944
R10354 gnd.n6017 gnd.n6016 19.3944
R10355 gnd.n6016 gnd.n1120 19.3944
R10356 gnd.n6006 gnd.n1120 19.3944
R10357 gnd.n6006 gnd.n6005 19.3944
R10358 gnd.n6005 gnd.n6004 19.3944
R10359 gnd.n1148 gnd.n1142 19.3944
R10360 gnd.n4357 gnd.n1148 19.3944
R10361 gnd.n4360 gnd.n4359 19.3944
R10362 gnd.n4390 gnd.n4389 19.3944
R10363 gnd.n6001 gnd.n1149 19.3944
R10364 gnd.n6001 gnd.n1150 19.3944
R10365 gnd.n5991 gnd.n1150 19.3944
R10366 gnd.n5991 gnd.n5990 19.3944
R10367 gnd.n5990 gnd.n5989 19.3944
R10368 gnd.n5989 gnd.n1171 19.3944
R10369 gnd.n5979 gnd.n1171 19.3944
R10370 gnd.n5979 gnd.n5978 19.3944
R10371 gnd.n5978 gnd.n5977 19.3944
R10372 gnd.n5977 gnd.n1193 19.3944
R10373 gnd.n5967 gnd.n1193 19.3944
R10374 gnd.n5967 gnd.n5966 19.3944
R10375 gnd.n5966 gnd.n5965 19.3944
R10376 gnd.n5965 gnd.n1213 19.3944
R10377 gnd.n5955 gnd.n1213 19.3944
R10378 gnd.n5955 gnd.n5954 19.3944
R10379 gnd.n5954 gnd.n5953 19.3944
R10380 gnd.n5953 gnd.n1235 19.3944
R10381 gnd.n5943 gnd.n1235 19.3944
R10382 gnd.n5943 gnd.n5942 19.3944
R10383 gnd.n5942 gnd.n5941 19.3944
R10384 gnd.n5941 gnd.n1256 19.3944
R10385 gnd.n5931 gnd.n1256 19.3944
R10386 gnd.n6191 gnd.n941 19.3944
R10387 gnd.n6185 gnd.n941 19.3944
R10388 gnd.n6185 gnd.n6184 19.3944
R10389 gnd.n6184 gnd.n6183 19.3944
R10390 gnd.n6183 gnd.n948 19.3944
R10391 gnd.n6177 gnd.n948 19.3944
R10392 gnd.n6177 gnd.n6176 19.3944
R10393 gnd.n6176 gnd.n6175 19.3944
R10394 gnd.n6175 gnd.n956 19.3944
R10395 gnd.n6169 gnd.n956 19.3944
R10396 gnd.n6169 gnd.n6168 19.3944
R10397 gnd.n6168 gnd.n6167 19.3944
R10398 gnd.n6167 gnd.n964 19.3944
R10399 gnd.n6161 gnd.n964 19.3944
R10400 gnd.n6161 gnd.n6160 19.3944
R10401 gnd.n6160 gnd.n6159 19.3944
R10402 gnd.n6159 gnd.n972 19.3944
R10403 gnd.n6153 gnd.n972 19.3944
R10404 gnd.n6153 gnd.n6152 19.3944
R10405 gnd.n6152 gnd.n6151 19.3944
R10406 gnd.n6151 gnd.n980 19.3944
R10407 gnd.n6145 gnd.n980 19.3944
R10408 gnd.n6145 gnd.n6144 19.3944
R10409 gnd.n6144 gnd.n6143 19.3944
R10410 gnd.n6143 gnd.n988 19.3944
R10411 gnd.n6137 gnd.n988 19.3944
R10412 gnd.n6137 gnd.n6136 19.3944
R10413 gnd.n6136 gnd.n6135 19.3944
R10414 gnd.n6135 gnd.n996 19.3944
R10415 gnd.n6129 gnd.n996 19.3944
R10416 gnd.n6129 gnd.n6128 19.3944
R10417 gnd.n6128 gnd.n6127 19.3944
R10418 gnd.n6127 gnd.n1004 19.3944
R10419 gnd.n6121 gnd.n1004 19.3944
R10420 gnd.n6121 gnd.n6120 19.3944
R10421 gnd.n6120 gnd.n6119 19.3944
R10422 gnd.n6119 gnd.n1012 19.3944
R10423 gnd.n6113 gnd.n1012 19.3944
R10424 gnd.n6113 gnd.n6112 19.3944
R10425 gnd.n6112 gnd.n6111 19.3944
R10426 gnd.n6111 gnd.n1020 19.3944
R10427 gnd.n6105 gnd.n1020 19.3944
R10428 gnd.n6105 gnd.n6104 19.3944
R10429 gnd.n6104 gnd.n6103 19.3944
R10430 gnd.n6103 gnd.n1028 19.3944
R10431 gnd.n6097 gnd.n1028 19.3944
R10432 gnd.n6097 gnd.n6096 19.3944
R10433 gnd.n6096 gnd.n6095 19.3944
R10434 gnd.n6095 gnd.n1036 19.3944
R10435 gnd.n6089 gnd.n1036 19.3944
R10436 gnd.n6089 gnd.n6088 19.3944
R10437 gnd.n6088 gnd.n6087 19.3944
R10438 gnd.n6087 gnd.n1044 19.3944
R10439 gnd.n6081 gnd.n1044 19.3944
R10440 gnd.n6081 gnd.n6080 19.3944
R10441 gnd.n6080 gnd.n6079 19.3944
R10442 gnd.n6079 gnd.n1052 19.3944
R10443 gnd.n6073 gnd.n1052 19.3944
R10444 gnd.n6073 gnd.n6072 19.3944
R10445 gnd.n6072 gnd.n6071 19.3944
R10446 gnd.n6071 gnd.n1060 19.3944
R10447 gnd.n6065 gnd.n1060 19.3944
R10448 gnd.n6065 gnd.n6064 19.3944
R10449 gnd.n6064 gnd.n6063 19.3944
R10450 gnd.n6063 gnd.n1068 19.3944
R10451 gnd.n6057 gnd.n1068 19.3944
R10452 gnd.n6057 gnd.n6056 19.3944
R10453 gnd.n6056 gnd.n6055 19.3944
R10454 gnd.n6055 gnd.n1076 19.3944
R10455 gnd.n6049 gnd.n1076 19.3944
R10456 gnd.n6049 gnd.n6048 19.3944
R10457 gnd.n6048 gnd.n6047 19.3944
R10458 gnd.n6047 gnd.n1084 19.3944
R10459 gnd.n6041 gnd.n1084 19.3944
R10460 gnd.n6041 gnd.n6040 19.3944
R10461 gnd.n6040 gnd.n6039 19.3944
R10462 gnd.n6039 gnd.n1092 19.3944
R10463 gnd.n6033 gnd.n1092 19.3944
R10464 gnd.n6033 gnd.n6032 19.3944
R10465 gnd.n6032 gnd.n6031 19.3944
R10466 gnd.n6031 gnd.n1100 19.3944
R10467 gnd.n6025 gnd.n1100 19.3944
R10468 gnd.n6025 gnd.n6024 19.3944
R10469 gnd.n6024 gnd.n6023 19.3944
R10470 gnd.n4613 gnd.n2200 19.3944
R10471 gnd.n4613 gnd.n2188 19.3944
R10472 gnd.n4628 gnd.n2188 19.3944
R10473 gnd.n4628 gnd.n2186 19.3944
R10474 gnd.n4632 gnd.n2186 19.3944
R10475 gnd.n4632 gnd.n2174 19.3944
R10476 gnd.n4647 gnd.n2174 19.3944
R10477 gnd.n4647 gnd.n2172 19.3944
R10478 gnd.n4651 gnd.n2172 19.3944
R10479 gnd.n4651 gnd.n1988 19.3944
R10480 gnd.n4673 gnd.n1988 19.3944
R10481 gnd.n4673 gnd.n1985 19.3944
R10482 gnd.n4686 gnd.n1985 19.3944
R10483 gnd.n4686 gnd.n1986 19.3944
R10484 gnd.n4682 gnd.n1986 19.3944
R10485 gnd.n4682 gnd.n4681 19.3944
R10486 gnd.n4681 gnd.n1927 19.3944
R10487 gnd.n4733 gnd.n1927 19.3944
R10488 gnd.n4733 gnd.n1924 19.3944
R10489 gnd.n4738 gnd.n1924 19.3944
R10490 gnd.n4738 gnd.n1925 19.3944
R10491 gnd.n1925 gnd.n1901 19.3944
R10492 gnd.n4802 gnd.n1901 19.3944
R10493 gnd.n4802 gnd.n1898 19.3944
R10494 gnd.n4807 gnd.n1898 19.3944
R10495 gnd.n4807 gnd.n1899 19.3944
R10496 gnd.n1899 gnd.n1871 19.3944
R10497 gnd.n4838 gnd.n1871 19.3944
R10498 gnd.n4838 gnd.n1869 19.3944
R10499 gnd.n4842 gnd.n1869 19.3944
R10500 gnd.n4842 gnd.n1848 19.3944
R10501 gnd.n4870 gnd.n1848 19.3944
R10502 gnd.n4870 gnd.n1845 19.3944
R10503 gnd.n4884 gnd.n1845 19.3944
R10504 gnd.n4884 gnd.n1846 19.3944
R10505 gnd.n4880 gnd.n1846 19.3944
R10506 gnd.n4880 gnd.n4879 19.3944
R10507 gnd.n4879 gnd.n4878 19.3944
R10508 gnd.n4878 gnd.n1809 19.3944
R10509 gnd.n5028 gnd.n1809 19.3944
R10510 gnd.n5028 gnd.n1806 19.3944
R10511 gnd.n5033 gnd.n1806 19.3944
R10512 gnd.n5033 gnd.n1807 19.3944
R10513 gnd.n1807 gnd.n1779 19.3944
R10514 gnd.n5064 gnd.n1779 19.3944
R10515 gnd.n5064 gnd.n1777 19.3944
R10516 gnd.n5068 gnd.n1777 19.3944
R10517 gnd.n5068 gnd.n1757 19.3944
R10518 gnd.n5091 gnd.n1757 19.3944
R10519 gnd.n5091 gnd.n1755 19.3944
R10520 gnd.n5095 gnd.n1755 19.3944
R10521 gnd.n5095 gnd.n1735 19.3944
R10522 gnd.n5121 gnd.n1735 19.3944
R10523 gnd.n5121 gnd.n1733 19.3944
R10524 gnd.n5125 gnd.n1733 19.3944
R10525 gnd.n5125 gnd.n1714 19.3944
R10526 gnd.n5151 gnd.n1714 19.3944
R10527 gnd.n5151 gnd.n1711 19.3944
R10528 gnd.n5156 gnd.n1711 19.3944
R10529 gnd.n5156 gnd.n1712 19.3944
R10530 gnd.n1712 gnd.n1685 19.3944
R10531 gnd.n5187 gnd.n1685 19.3944
R10532 gnd.n5187 gnd.n1683 19.3944
R10533 gnd.n5191 gnd.n1683 19.3944
R10534 gnd.n5191 gnd.n1661 19.3944
R10535 gnd.n5226 gnd.n1661 19.3944
R10536 gnd.n5226 gnd.n1659 19.3944
R10537 gnd.n5230 gnd.n1659 19.3944
R10538 gnd.n5230 gnd.n1605 19.3944
R10539 gnd.n5397 gnd.n1605 19.3944
R10540 gnd.n5397 gnd.n1603 19.3944
R10541 gnd.n5401 gnd.n1603 19.3944
R10542 gnd.n5401 gnd.n1590 19.3944
R10543 gnd.n5416 gnd.n1590 19.3944
R10544 gnd.n5416 gnd.n1588 19.3944
R10545 gnd.n5420 gnd.n1588 19.3944
R10546 gnd.n5420 gnd.n1577 19.3944
R10547 gnd.n5438 gnd.n1577 19.3944
R10548 gnd.n5438 gnd.n1575 19.3944
R10549 gnd.n5442 gnd.n1575 19.3944
R10550 gnd.n5442 gnd.n1475 19.3944
R10551 gnd.n5706 gnd.n1475 19.3944
R10552 gnd.n5638 gnd.n5637 19.3944
R10553 gnd.n5637 gnd.n5636 19.3944
R10554 gnd.n5636 gnd.n5633 19.3944
R10555 gnd.n5696 gnd.n1483 19.3944
R10556 gnd.n5696 gnd.n5695 19.3944
R10557 gnd.n5695 gnd.n1486 19.3944
R10558 gnd.n5688 gnd.n1486 19.3944
R10559 gnd.n5688 gnd.n5687 19.3944
R10560 gnd.n5687 gnd.n1496 19.3944
R10561 gnd.n5680 gnd.n1496 19.3944
R10562 gnd.n5680 gnd.n5679 19.3944
R10563 gnd.n5679 gnd.n1504 19.3944
R10564 gnd.n5672 gnd.n1504 19.3944
R10565 gnd.n5672 gnd.n5671 19.3944
R10566 gnd.n5671 gnd.n1514 19.3944
R10567 gnd.n5664 gnd.n1514 19.3944
R10568 gnd.n5664 gnd.n5663 19.3944
R10569 gnd.n5663 gnd.n1522 19.3944
R10570 gnd.n5653 gnd.n1522 19.3944
R10571 gnd.n5653 gnd.n5652 19.3944
R10572 gnd.n5652 gnd.n5649 19.3944
R10573 gnd.n5649 gnd.n5648 19.3944
R10574 gnd.n5648 gnd.n1532 19.3944
R10575 gnd.n5644 gnd.n1532 19.3944
R10576 gnd.n5644 gnd.n5643 19.3944
R10577 gnd.n5643 gnd.n5642 19.3944
R10578 gnd.n5642 gnd.n1537 19.3944
R10579 gnd.n3306 gnd.t165 18.8012
R10580 gnd.n3291 gnd.t172 18.8012
R10581 gnd.n4691 gnd.n1979 18.5761
R10582 gnd.n5324 gnd.n5323 18.5761
R10583 gnd.n3150 gnd.n3149 18.4825
R10584 gnd.n6939 gnd.n6938 18.4247
R10585 gnd.n1302 gnd.n1298 18.4247
R10586 gnd.n7218 gnd.n7217 18.2308
R10587 gnd.n5660 gnd.n5659 18.2308
R10588 gnd.n4567 gnd.n4566 18.2308
R10589 gnd.n4177 gnd.n4123 18.2308
R10590 gnd.t150 gnd.n2830 18.1639
R10591 gnd.n2858 gnd.t163 17.5266
R10592 gnd.n4238 gnd.t234 17.5266
R10593 gnd.n5951 gnd.t186 17.5266
R10594 gnd.n5606 gnd.t255 17.5266
R10595 gnd.t262 gnd.n196 17.5266
R10596 gnd.n3257 gnd.t158 16.8893
R10597 gnd.n4281 gnd.t219 16.8893
R10598 gnd.n5975 gnd.t180 16.8893
R10599 gnd.n5518 gnd.t192 16.8893
R10600 gnd.t232 gnd.n225 16.8893
R10601 gnd.n3085 gnd.t60 16.2519
R10602 gnd.n2785 gnd.t157 16.2519
R10603 gnd.n5999 gnd.t198 16.2519
R10604 gnd.n7058 gnd.t184 16.2519
R10605 gnd.n4557 gnd.n2264 15.9333
R10606 gnd.n4557 gnd.n4554 15.9333
R10607 gnd.n2284 gnd.n2283 15.9333
R10608 gnd.n2283 gnd.n2198 15.9333
R10609 gnd.n4615 gnd.n2198 15.9333
R10610 gnd.n4617 gnd.n4615 15.9333
R10611 gnd.n4616 gnd.n2190 15.9333
R10612 gnd.n4626 gnd.n2190 15.9333
R10613 gnd.n4626 gnd.n4625 15.9333
R10614 gnd.n4625 gnd.n2192 15.9333
R10615 gnd.n2192 gnd.n2184 15.9333
R10616 gnd.n4634 gnd.n2184 15.9333
R10617 gnd.n4636 gnd.n4634 15.9333
R10618 gnd.n4636 gnd.n4635 15.9333
R10619 gnd.n4645 gnd.n2176 15.9333
R10620 gnd.n4645 gnd.n4644 15.9333
R10621 gnd.n4644 gnd.n2178 15.9333
R10622 gnd.n2178 gnd.n2170 15.9333
R10623 gnd.n4653 gnd.n2170 15.9333
R10624 gnd.n4656 gnd.n4653 15.9333
R10625 gnd.n4656 gnd.n4655 15.9333
R10626 gnd.n4655 gnd.n4654 15.9333
R10627 gnd.n4671 gnd.n4670 15.9333
R10628 gnd.n2164 gnd.n2163 15.9333
R10629 gnd.n4664 gnd.n1954 15.9333
R10630 gnd.n4708 gnd.n1948 15.9333
R10631 gnd.n4722 gnd.n4721 15.9333
R10632 gnd.n4791 gnd.n1911 15.9333
R10633 gnd.n4800 gnd.n4799 15.9333
R10634 gnd.n4868 gnd.n4867 15.9333
R10635 gnd.n4910 gnd.n1828 15.9333
R10636 gnd.n5017 gnd.n1818 15.9333
R10637 gnd.n5026 gnd.n5025 15.9333
R10638 gnd.n5036 gnd.n5035 15.9333
R10639 gnd.n4985 gnd.n1787 15.9333
R10640 gnd.n4977 gnd.n1783 15.9333
R10641 gnd.n5088 gnd.n1750 15.9333
R10642 gnd.n5159 gnd.n5158 15.9333
R10643 gnd.n4941 gnd.n1692 15.9333
R10644 gnd.n4932 gnd.n1688 15.9333
R10645 gnd.n5204 gnd.n5203 15.9333
R10646 gnd.n5223 gnd.n1665 15.9333
R10647 gnd.n5232 gnd.n1657 15.9333
R10648 gnd.n5395 gnd.n1607 15.9333
R10649 gnd.n5403 gnd.n1601 15.9333
R10650 gnd.n5405 gnd.n5403 15.9333
R10651 gnd.n5405 gnd.n5404 15.9333
R10652 gnd.n5404 gnd.n1592 15.9333
R10653 gnd.n5414 gnd.n1592 15.9333
R10654 gnd.n5414 gnd.n5413 15.9333
R10655 gnd.n5413 gnd.n1595 15.9333
R10656 gnd.n1595 gnd.n1594 15.9333
R10657 gnd.n5424 gnd.n5422 15.9333
R10658 gnd.n5424 gnd.n5423 15.9333
R10659 gnd.n5423 gnd.n1579 15.9333
R10660 gnd.n5436 gnd.n1579 15.9333
R10661 gnd.n5436 gnd.n5435 15.9333
R10662 gnd.n5435 gnd.n1581 15.9333
R10663 gnd.n1581 gnd.n1573 15.9333
R10664 gnd.n5444 gnd.n1573 15.9333
R10665 gnd.n5446 gnd.n5445 15.9333
R10666 gnd.n5445 gnd.n1471 15.9333
R10667 gnd.n5708 gnd.n1471 15.9333
R10668 gnd.n5708 gnd.n1472 15.9333
R10669 gnd.n5630 gnd.n1544 15.9333
R10670 gnd.n5630 gnd.n5629 15.9333
R10671 gnd.n3772 gnd.n3770 15.6674
R10672 gnd.n3740 gnd.n3738 15.6674
R10673 gnd.n3708 gnd.n3706 15.6674
R10674 gnd.n3677 gnd.n3675 15.6674
R10675 gnd.n3645 gnd.n3643 15.6674
R10676 gnd.n3613 gnd.n3611 15.6674
R10677 gnd.n3581 gnd.n3579 15.6674
R10678 gnd.n3550 gnd.n3548 15.6674
R10679 gnd.n3076 gnd.t60 15.6146
R10680 gnd.t101 gnd.n2538 15.6146
R10681 gnd.t81 gnd.n2539 15.6146
R10682 gnd.n4318 gnd.t206 15.6146
R10683 gnd.t91 gnd.n4616 15.6146
R10684 gnd.t74 gnd.n5444 15.6146
R10685 gnd.n7090 gnd.t203 15.6146
R10686 gnd.n4772 gnd.n1903 15.296
R10687 gnd.n4818 gnd.n1888 15.296
R10688 gnd.t136 gnd.n1880 15.296
R10689 gnd.n4998 gnd.n1811 15.296
R10690 gnd.n5044 gnd.n1795 15.296
R10691 gnd.n5127 gnd.t143 15.296
R10692 gnd.n4953 gnd.n1716 15.296
R10693 gnd.n5167 gnd.n1700 15.296
R10694 gnd.n5241 gnd.n5240 15.0827
R10695 gnd.n1967 gnd.n1962 15.0481
R10696 gnd.n5251 gnd.n5250 15.0481
R10697 gnd.n3444 gnd.t152 14.9773
R10698 gnd.t219 gnd.n1109 14.9773
R10699 gnd.n4654 gnd.t176 14.9773
R10700 gnd.t9 gnd.n1601 14.9773
R10701 gnd.n7122 gnd.t232 14.9773
R10702 gnd.n4688 gnd.n1982 14.6587
R10703 gnd.n4844 gnd.n1858 14.6587
R10704 gnd.n5109 gnd.n1745 14.6587
R10705 gnd.n5193 gnd.n1673 14.6587
R10706 gnd.t15 gnd.n2582 14.34
R10707 gnd.n3522 gnd.t161 14.34
R10708 gnd.t234 gnd.n2426 14.34
R10709 gnd.n7154 gnd.t262 14.34
R10710 gnd.n4731 gnd.t85 14.0214
R10711 gnd.n4780 gnd.n4779 14.0214
R10712 gnd.n4829 gnd.n4828 14.0214
R10713 gnd.n5006 gnd.n5005 14.0214
R10714 gnd.n5055 gnd.n5054 14.0214
R10715 gnd.n5129 gnd.n5128 14.0214
R10716 gnd.n5178 gnd.n5177 14.0214
R10717 gnd.t98 gnd.n1626 14.0214
R10718 gnd.n3232 gnd.t144 13.7027
R10719 gnd.n4902 gnd.t170 13.7027
R10720 gnd.n5080 gnd.t141 13.7027
R10721 gnd.n2942 gnd.n2941 13.5763
R10722 gnd.n3886 gnd.n2495 13.5763
R10723 gnd.n6901 gnd.n467 13.5763
R10724 gnd.n7256 gnd.n7255 13.5763
R10725 gnd.n3929 gnd.n3928 13.5763
R10726 gnd.n5867 gnd.n1339 13.5763
R10727 gnd.n3150 gnd.n2888 13.384
R10728 gnd.n4741 gnd.n4740 13.384
R10729 gnd.n4836 gnd.n4835 13.384
R10730 gnd.n4753 gnd.t128 13.384
R10731 gnd.n5119 gnd.t130 13.384
R10732 gnd.n1738 gnd.n1728 13.384
R10733 gnd.n5185 gnd.n5184 13.384
R10734 gnd.n1978 gnd.n1959 13.1884
R10735 gnd.n1973 gnd.n1972 13.1884
R10736 gnd.n1972 gnd.n1971 13.1884
R10737 gnd.n5244 gnd.n5239 13.1884
R10738 gnd.n5245 gnd.n5244 13.1884
R10739 gnd.n1974 gnd.n1961 13.146
R10740 gnd.n1970 gnd.n1961 13.146
R10741 gnd.n5243 gnd.n5242 13.146
R10742 gnd.n5243 gnd.n5238 13.146
R10743 gnd.n2163 gnd.n2161 13.0654
R10744 gnd.n5224 gnd.t308 13.0654
R10745 gnd.n5395 gnd.n5394 13.0654
R10746 gnd.n3773 gnd.n3769 12.8005
R10747 gnd.n3741 gnd.n3737 12.8005
R10748 gnd.n3709 gnd.n3705 12.8005
R10749 gnd.n3678 gnd.n3674 12.8005
R10750 gnd.n3646 gnd.n3642 12.8005
R10751 gnd.n3614 gnd.n3610 12.8005
R10752 gnd.n3582 gnd.n3578 12.8005
R10753 gnd.n3551 gnd.n3547 12.8005
R10754 gnd.n1934 gnd.n1930 12.7467
R10755 gnd.n4895 gnd.n4894 12.7467
R10756 gnd.n4978 gnd.n1773 12.7467
R10757 gnd.n4933 gnd.n1680 12.7467
R10758 gnd.n2941 gnd.n2936 12.4126
R10759 gnd.n3889 gnd.n3886 12.4126
R10760 gnd.n6897 gnd.n467 12.4126
R10761 gnd.n7255 gnd.n174 12.4126
R10762 gnd.n4062 gnd.n3928 12.4126
R10763 gnd.n5862 gnd.n1339 12.4126
R10764 gnd.n2024 gnd.n1979 12.1761
R10765 gnd.n5323 gnd.n5322 12.1761
R10766 gnd.n4790 gnd.n1913 12.1094
R10767 gnd.n4762 gnd.n1890 12.1094
R10768 gnd.n5139 gnd.n1723 12.1094
R10769 gnd.n4942 gnd.n1702 12.1094
R10770 gnd.n3777 gnd.n3776 12.0247
R10771 gnd.n3745 gnd.n3744 12.0247
R10772 gnd.n3713 gnd.n3712 12.0247
R10773 gnd.n3682 gnd.n3681 12.0247
R10774 gnd.n3650 gnd.n3649 12.0247
R10775 gnd.n3618 gnd.n3617 12.0247
R10776 gnd.n3586 gnd.n3585 12.0247
R10777 gnd.n3555 gnd.n3554 12.0247
R10778 gnd.n4543 gnd.n1276 11.4721
R10779 gnd.n4723 gnd.n1938 11.4721
R10780 gnd.t135 gnd.n4858 11.4721
R10781 gnd.n4857 gnd.n1861 11.4721
R10782 gnd.n4887 gnd.n1842 11.4721
R10783 gnd.n5078 gnd.n1768 11.4721
R10784 gnd.n5099 gnd.n5098 11.4721
R10785 gnd.n5097 gnd.t166 11.4721
R10786 gnd.n5202 gnd.n1675 11.4721
R10787 gnd.n5233 gnd.n1654 11.4721
R10788 gnd.n1656 gnd.t68 11.4721
R10789 gnd.n6966 gnd.n395 11.4721
R10790 gnd.n7248 gnd.n100 11.4721
R10791 gnd.n3780 gnd.n3767 11.249
R10792 gnd.n3748 gnd.n3735 11.249
R10793 gnd.n3716 gnd.n3703 11.249
R10794 gnd.n3685 gnd.n3672 11.249
R10795 gnd.n3653 gnd.n3640 11.249
R10796 gnd.n3621 gnd.n3608 11.249
R10797 gnd.n3589 gnd.n3576 11.249
R10798 gnd.n3558 gnd.n3545 11.249
R10799 gnd.n3220 gnd.t144 11.1535
R10800 gnd.n4343 gnd.t206 11.1535
R10801 gnd.n4635 gnd.t137 11.1535
R10802 gnd.n4754 gnd.t167 11.1535
R10803 gnd.t0 gnd.n1737 11.1535
R10804 gnd.n5422 gnd.t178 11.1535
R10805 gnd.n6836 gnd.t203 11.1535
R10806 gnd.n1905 gnd.n1894 10.8348
R10807 gnd.n4811 gnd.n1894 10.8348
R10808 gnd.n1812 gnd.n1802 10.8348
R10809 gnd.n5037 gnd.n1802 10.8348
R10810 gnd.n4950 gnd.n1706 10.8348
R10811 gnd.n5160 gnd.n1706 10.8348
R10812 gnd.n5391 gnd.n5390 10.6151
R10813 gnd.n5390 gnd.n5387 10.6151
R10814 gnd.n5385 gnd.n5382 10.6151
R10815 gnd.n5382 gnd.n5381 10.6151
R10816 gnd.n5381 gnd.n5378 10.6151
R10817 gnd.n5378 gnd.n5377 10.6151
R10818 gnd.n5377 gnd.n5374 10.6151
R10819 gnd.n5374 gnd.n5373 10.6151
R10820 gnd.n5373 gnd.n5370 10.6151
R10821 gnd.n5370 gnd.n5369 10.6151
R10822 gnd.n5369 gnd.n5366 10.6151
R10823 gnd.n5366 gnd.n5365 10.6151
R10824 gnd.n5365 gnd.n5362 10.6151
R10825 gnd.n5362 gnd.n5361 10.6151
R10826 gnd.n5361 gnd.n5358 10.6151
R10827 gnd.n5358 gnd.n5357 10.6151
R10828 gnd.n5357 gnd.n5354 10.6151
R10829 gnd.n5354 gnd.n5353 10.6151
R10830 gnd.n5353 gnd.n5350 10.6151
R10831 gnd.n5350 gnd.n5349 10.6151
R10832 gnd.n5349 gnd.n5346 10.6151
R10833 gnd.n5346 gnd.n5345 10.6151
R10834 gnd.n5345 gnd.n5342 10.6151
R10835 gnd.n5342 gnd.n5341 10.6151
R10836 gnd.n5341 gnd.n5338 10.6151
R10837 gnd.n5338 gnd.n5337 10.6151
R10838 gnd.n5337 gnd.n5334 10.6151
R10839 gnd.n5334 gnd.n5333 10.6151
R10840 gnd.n5333 gnd.n5330 10.6151
R10841 gnd.n5330 gnd.n5329 10.6151
R10842 gnd.n2030 gnd.n1952 10.6151
R10843 gnd.n4699 gnd.n1952 10.6151
R10844 gnd.n4700 gnd.n4699 10.6151
R10845 gnd.n4706 gnd.n4700 10.6151
R10846 gnd.n4706 gnd.n4705 10.6151
R10847 gnd.n4705 gnd.n4704 10.6151
R10848 gnd.n4704 gnd.n4703 10.6151
R10849 gnd.n4703 gnd.n4701 10.6151
R10850 gnd.n4701 gnd.n1919 10.6151
R10851 gnd.n4743 gnd.n1919 10.6151
R10852 gnd.n4744 gnd.n4743 10.6151
R10853 gnd.n4777 gnd.n4744 10.6151
R10854 gnd.n4777 gnd.n4776 10.6151
R10855 gnd.n4776 gnd.n4775 10.6151
R10856 gnd.n4775 gnd.n4745 10.6151
R10857 gnd.n4769 gnd.n4745 10.6151
R10858 gnd.n4769 gnd.n4768 10.6151
R10859 gnd.n4768 gnd.n4767 10.6151
R10860 gnd.n4767 gnd.n4765 10.6151
R10861 gnd.n4765 gnd.n4764 10.6151
R10862 gnd.n4764 gnd.n4760 10.6151
R10863 gnd.n4760 gnd.n4759 10.6151
R10864 gnd.n4759 gnd.n4757 10.6151
R10865 gnd.n4757 gnd.n4756 10.6151
R10866 gnd.n4756 gnd.n4752 10.6151
R10867 gnd.n4752 gnd.n4751 10.6151
R10868 gnd.n4751 gnd.n4749 10.6151
R10869 gnd.n4749 gnd.n4748 10.6151
R10870 gnd.n4748 gnd.n4746 10.6151
R10871 gnd.n4746 gnd.n1840 10.6151
R10872 gnd.n4889 gnd.n1840 10.6151
R10873 gnd.n4890 gnd.n4889 10.6151
R10874 gnd.n4891 gnd.n4890 10.6151
R10875 gnd.n4891 gnd.n1826 10.6151
R10876 gnd.n4913 gnd.n1826 10.6151
R10877 gnd.n4914 gnd.n4913 10.6151
R10878 gnd.n5003 gnd.n4914 10.6151
R10879 gnd.n5003 gnd.n5002 10.6151
R10880 gnd.n5002 gnd.n5001 10.6151
R10881 gnd.n5001 gnd.n4915 10.6151
R10882 gnd.n4993 gnd.n4915 10.6151
R10883 gnd.n4993 gnd.n4992 10.6151
R10884 gnd.n4992 gnd.n4991 10.6151
R10885 gnd.n4991 gnd.n4989 10.6151
R10886 gnd.n4989 gnd.n4988 10.6151
R10887 gnd.n4988 gnd.n4984 10.6151
R10888 gnd.n4984 gnd.n4983 10.6151
R10889 gnd.n4983 gnd.n4981 10.6151
R10890 gnd.n4981 gnd.n4980 10.6151
R10891 gnd.n4980 gnd.n4976 10.6151
R10892 gnd.n4976 gnd.n4975 10.6151
R10893 gnd.n4975 gnd.n4973 10.6151
R10894 gnd.n4973 gnd.n4972 10.6151
R10895 gnd.n4972 gnd.n4970 10.6151
R10896 gnd.n4970 gnd.n4969 10.6151
R10897 gnd.n4969 gnd.n4968 10.6151
R10898 gnd.n4968 gnd.n4967 10.6151
R10899 gnd.n4967 gnd.n4966 10.6151
R10900 gnd.n4966 gnd.n4916 10.6151
R10901 gnd.n4960 gnd.n4916 10.6151
R10902 gnd.n4960 gnd.n4959 10.6151
R10903 gnd.n4959 gnd.n4958 10.6151
R10904 gnd.n4958 gnd.n4957 10.6151
R10905 gnd.n4957 gnd.n4956 10.6151
R10906 gnd.n4956 gnd.n4917 10.6151
R10907 gnd.n4949 gnd.n4917 10.6151
R10908 gnd.n4949 gnd.n4948 10.6151
R10909 gnd.n4948 gnd.n4947 10.6151
R10910 gnd.n4947 gnd.n4945 10.6151
R10911 gnd.n4945 gnd.n4944 10.6151
R10912 gnd.n4944 gnd.n4940 10.6151
R10913 gnd.n4940 gnd.n4939 10.6151
R10914 gnd.n4939 gnd.n4936 10.6151
R10915 gnd.n4936 gnd.n4935 10.6151
R10916 gnd.n4935 gnd.n4930 10.6151
R10917 gnd.n4930 gnd.n4929 10.6151
R10918 gnd.n4929 gnd.n4927 10.6151
R10919 gnd.n4927 gnd.n4926 10.6151
R10920 gnd.n4926 gnd.n4923 10.6151
R10921 gnd.n4923 gnd.n4922 10.6151
R10922 gnd.n4922 gnd.n4919 10.6151
R10923 gnd.n4919 gnd.n4918 10.6151
R10924 gnd.n4918 gnd.n1647 10.6151
R10925 gnd.n2094 gnd.n2093 10.6151
R10926 gnd.n2093 gnd.n2090 10.6151
R10927 gnd.n2088 gnd.n2085 10.6151
R10928 gnd.n2085 gnd.n2084 10.6151
R10929 gnd.n2084 gnd.n2081 10.6151
R10930 gnd.n2081 gnd.n2080 10.6151
R10931 gnd.n2080 gnd.n2077 10.6151
R10932 gnd.n2077 gnd.n2076 10.6151
R10933 gnd.n2076 gnd.n2073 10.6151
R10934 gnd.n2073 gnd.n2072 10.6151
R10935 gnd.n2072 gnd.n2069 10.6151
R10936 gnd.n2069 gnd.n2068 10.6151
R10937 gnd.n2068 gnd.n2065 10.6151
R10938 gnd.n2065 gnd.n2064 10.6151
R10939 gnd.n2064 gnd.n2061 10.6151
R10940 gnd.n2061 gnd.n2060 10.6151
R10941 gnd.n2060 gnd.n2057 10.6151
R10942 gnd.n2057 gnd.n2056 10.6151
R10943 gnd.n2056 gnd.n2053 10.6151
R10944 gnd.n2053 gnd.n2052 10.6151
R10945 gnd.n2052 gnd.n2049 10.6151
R10946 gnd.n2049 gnd.n2048 10.6151
R10947 gnd.n2048 gnd.n2045 10.6151
R10948 gnd.n2045 gnd.n2044 10.6151
R10949 gnd.n2044 gnd.n2041 10.6151
R10950 gnd.n2041 gnd.n2040 10.6151
R10951 gnd.n2040 gnd.n2037 10.6151
R10952 gnd.n2037 gnd.n2036 10.6151
R10953 gnd.n2036 gnd.n2033 10.6151
R10954 gnd.n2033 gnd.n2032 10.6151
R10955 gnd.n2158 gnd.n2024 10.6151
R10956 gnd.n2158 gnd.n2157 10.6151
R10957 gnd.n2157 gnd.n2156 10.6151
R10958 gnd.n2156 gnd.n2154 10.6151
R10959 gnd.n2154 gnd.n2151 10.6151
R10960 gnd.n2151 gnd.n2150 10.6151
R10961 gnd.n2150 gnd.n2147 10.6151
R10962 gnd.n2147 gnd.n2146 10.6151
R10963 gnd.n2146 gnd.n2143 10.6151
R10964 gnd.n2143 gnd.n2142 10.6151
R10965 gnd.n2142 gnd.n2139 10.6151
R10966 gnd.n2139 gnd.n2138 10.6151
R10967 gnd.n2138 gnd.n2135 10.6151
R10968 gnd.n2135 gnd.n2134 10.6151
R10969 gnd.n2134 gnd.n2131 10.6151
R10970 gnd.n2131 gnd.n2130 10.6151
R10971 gnd.n2130 gnd.n2127 10.6151
R10972 gnd.n2127 gnd.n2126 10.6151
R10973 gnd.n2126 gnd.n2123 10.6151
R10974 gnd.n2123 gnd.n2122 10.6151
R10975 gnd.n2122 gnd.n2119 10.6151
R10976 gnd.n2119 gnd.n2118 10.6151
R10977 gnd.n2118 gnd.n2115 10.6151
R10978 gnd.n2115 gnd.n2114 10.6151
R10979 gnd.n2114 gnd.n2111 10.6151
R10980 gnd.n2111 gnd.n2110 10.6151
R10981 gnd.n2110 gnd.n2107 10.6151
R10982 gnd.n2107 gnd.n2106 10.6151
R10983 gnd.n2103 gnd.n2102 10.6151
R10984 gnd.n2102 gnd.n2099 10.6151
R10985 gnd.n5322 gnd.n5321 10.6151
R10986 gnd.n5321 gnd.n5318 10.6151
R10987 gnd.n5318 gnd.n5317 10.6151
R10988 gnd.n5317 gnd.n5314 10.6151
R10989 gnd.n5314 gnd.n5313 10.6151
R10990 gnd.n5313 gnd.n5310 10.6151
R10991 gnd.n5310 gnd.n5309 10.6151
R10992 gnd.n5309 gnd.n5306 10.6151
R10993 gnd.n5306 gnd.n5305 10.6151
R10994 gnd.n5305 gnd.n5302 10.6151
R10995 gnd.n5302 gnd.n5301 10.6151
R10996 gnd.n5301 gnd.n5298 10.6151
R10997 gnd.n5298 gnd.n5297 10.6151
R10998 gnd.n5297 gnd.n5294 10.6151
R10999 gnd.n5294 gnd.n5293 10.6151
R11000 gnd.n5293 gnd.n5290 10.6151
R11001 gnd.n5290 gnd.n5289 10.6151
R11002 gnd.n5289 gnd.n5286 10.6151
R11003 gnd.n5286 gnd.n5285 10.6151
R11004 gnd.n5285 gnd.n5282 10.6151
R11005 gnd.n5282 gnd.n5281 10.6151
R11006 gnd.n5281 gnd.n5278 10.6151
R11007 gnd.n5278 gnd.n5277 10.6151
R11008 gnd.n5277 gnd.n5274 10.6151
R11009 gnd.n5274 gnd.n5273 10.6151
R11010 gnd.n5273 gnd.n5270 10.6151
R11011 gnd.n5270 gnd.n5269 10.6151
R11012 gnd.n5269 gnd.n5266 10.6151
R11013 gnd.n5264 gnd.n5261 10.6151
R11014 gnd.n5261 gnd.n5260 10.6151
R11015 gnd.n4692 gnd.n4691 10.6151
R11016 gnd.n4695 gnd.n4692 10.6151
R11017 gnd.n4695 gnd.n4694 10.6151
R11018 gnd.n4694 gnd.n4693 10.6151
R11019 gnd.n4693 gnd.n1936 10.6151
R11020 gnd.n4725 gnd.n1936 10.6151
R11021 gnd.n4726 gnd.n4725 10.6151
R11022 gnd.n4728 gnd.n4726 10.6151
R11023 gnd.n4728 gnd.n4727 10.6151
R11024 gnd.n4727 gnd.n1916 10.6151
R11025 gnd.n4783 gnd.n1916 10.6151
R11026 gnd.n4784 gnd.n4783 10.6151
R11027 gnd.n4788 gnd.n4784 10.6151
R11028 gnd.n4788 gnd.n4787 10.6151
R11029 gnd.n4787 gnd.n4786 10.6151
R11030 gnd.n4786 gnd.n1892 10.6151
R11031 gnd.n4813 gnd.n1892 10.6151
R11032 gnd.n4814 gnd.n4813 10.6151
R11033 gnd.n4815 gnd.n4814 10.6151
R11034 gnd.n4815 gnd.n1877 10.6151
R11035 gnd.n4831 gnd.n1877 10.6151
R11036 gnd.n4832 gnd.n4831 10.6151
R11037 gnd.n4833 gnd.n4832 10.6151
R11038 gnd.n4833 gnd.n1864 10.6151
R11039 gnd.n4847 gnd.n1864 10.6151
R11040 gnd.n4848 gnd.n4847 10.6151
R11041 gnd.n4855 gnd.n4848 10.6151
R11042 gnd.n4855 gnd.n4854 10.6151
R11043 gnd.n4854 gnd.n4853 10.6151
R11044 gnd.n4853 gnd.n4852 10.6151
R11045 gnd.n4852 gnd.n1837 10.6151
R11046 gnd.n4899 gnd.n1837 10.6151
R11047 gnd.n4899 gnd.n4898 10.6151
R11048 gnd.n4898 gnd.n4897 10.6151
R11049 gnd.n4897 gnd.n1822 10.6151
R11050 gnd.n5009 gnd.n1822 10.6151
R11051 gnd.n5010 gnd.n5009 10.6151
R11052 gnd.n5014 gnd.n5010 10.6151
R11053 gnd.n5014 gnd.n5013 10.6151
R11054 gnd.n5013 gnd.n5012 10.6151
R11055 gnd.n5012 gnd.n1800 10.6151
R11056 gnd.n5039 gnd.n1800 10.6151
R11057 gnd.n5040 gnd.n5039 10.6151
R11058 gnd.n5041 gnd.n5040 10.6151
R11059 gnd.n5041 gnd.n1785 10.6151
R11060 gnd.n5057 gnd.n1785 10.6151
R11061 gnd.n5058 gnd.n5057 10.6151
R11062 gnd.n5059 gnd.n5058 10.6151
R11063 gnd.n5059 gnd.n1771 10.6151
R11064 gnd.n5073 gnd.n1771 10.6151
R11065 gnd.n5074 gnd.n5073 10.6151
R11066 gnd.n5076 gnd.n5074 10.6151
R11067 gnd.n5076 gnd.n5075 10.6151
R11068 gnd.n5075 gnd.n1748 10.6151
R11069 gnd.n5102 gnd.n1748 10.6151
R11070 gnd.n5103 gnd.n5102 10.6151
R11071 gnd.n5107 gnd.n5103 10.6151
R11072 gnd.n5107 gnd.n5106 10.6151
R11073 gnd.n5106 gnd.n5105 10.6151
R11074 gnd.n5105 gnd.n1726 10.6151
R11075 gnd.n5132 gnd.n1726 10.6151
R11076 gnd.n5133 gnd.n5132 10.6151
R11077 gnd.n5137 gnd.n5133 10.6151
R11078 gnd.n5137 gnd.n5136 10.6151
R11079 gnd.n5136 gnd.n5135 10.6151
R11080 gnd.n5135 gnd.n1704 10.6151
R11081 gnd.n5162 gnd.n1704 10.6151
R11082 gnd.n5163 gnd.n5162 10.6151
R11083 gnd.n5164 gnd.n5163 10.6151
R11084 gnd.n5164 gnd.n1690 10.6151
R11085 gnd.n5180 gnd.n1690 10.6151
R11086 gnd.n5181 gnd.n5180 10.6151
R11087 gnd.n5182 gnd.n5181 10.6151
R11088 gnd.n5182 gnd.n1678 10.6151
R11089 gnd.n5196 gnd.n1678 10.6151
R11090 gnd.n5197 gnd.n5196 10.6151
R11091 gnd.n5200 gnd.n5197 10.6151
R11092 gnd.n5200 gnd.n5199 10.6151
R11093 gnd.n5199 gnd.n5198 10.6151
R11094 gnd.n5198 gnd.n1652 10.6151
R11095 gnd.n5235 gnd.n1652 10.6151
R11096 gnd.n5236 gnd.n5235 10.6151
R11097 gnd.n5324 gnd.n5236 10.6151
R11098 gnd.n3139 gnd.t310 10.5161
R11099 gnd.n2584 gnd.t15 10.5161
R11100 gnd.n3505 gnd.t161 10.5161
R11101 gnd.n4431 gnd.t198 10.5161
R11102 gnd.n4810 gnd.t174 10.5161
R11103 gnd.t11 gnd.n5148 10.5161
R11104 gnd.n5555 gnd.t184 10.5161
R11105 gnd.n3781 gnd.n3765 10.4732
R11106 gnd.n3749 gnd.n3733 10.4732
R11107 gnd.n3717 gnd.n3701 10.4732
R11108 gnd.n3686 gnd.n3670 10.4732
R11109 gnd.n3654 gnd.n3638 10.4732
R11110 gnd.n3622 gnd.n3606 10.4732
R11111 gnd.n3590 gnd.n3574 10.4732
R11112 gnd.n3559 gnd.n3543 10.4732
R11113 gnd.n1957 gnd.n1956 10.1975
R11114 gnd.n4678 gnd.n1938 10.1975
R11115 gnd.n1861 gnd.n1850 10.1975
R11116 gnd.n4850 gnd.n1842 10.1975
R11117 gnd.n1768 gnd.n1759 10.1975
R11118 gnd.n5100 gnd.n5099 10.1975
R11119 gnd.t152 gnd.n2601 9.87883
R11120 gnd.n4469 gnd.t180 9.87883
R11121 gnd.t123 gnd.t126 9.87883
R11122 gnd.t192 gnd.n325 9.87883
R11123 gnd.n7370 gnd.n62 9.73455
R11124 gnd.n3785 gnd.n3784 9.69747
R11125 gnd.n3753 gnd.n3752 9.69747
R11126 gnd.n3721 gnd.n3720 9.69747
R11127 gnd.n3690 gnd.n3689 9.69747
R11128 gnd.n3658 gnd.n3657 9.69747
R11129 gnd.n3626 gnd.n3625 9.69747
R11130 gnd.n3594 gnd.n3593 9.69747
R11131 gnd.n3563 gnd.n3562 9.69747
R11132 gnd.n4773 gnd.n1913 9.56018
R11133 gnd.n4817 gnd.n1890 9.56018
R11134 gnd.n4849 gnd.t132 9.56018
R11135 gnd.n4999 gnd.n4997 9.56018
R11136 gnd.n5043 gnd.n1798 9.56018
R11137 gnd.n5089 gnd.t14 9.56018
R11138 gnd.n4954 gnd.n1723 9.56018
R11139 gnd.n5166 gnd.n1702 9.56018
R11140 gnd.n4609 gnd.n4608 9.45599
R11141 gnd.n5703 gnd.n5702 9.45599
R11142 gnd.n3791 gnd.n3790 9.45567
R11143 gnd.n3759 gnd.n3758 9.45567
R11144 gnd.n3727 gnd.n3726 9.45567
R11145 gnd.n3696 gnd.n3695 9.45567
R11146 gnd.n3664 gnd.n3663 9.45567
R11147 gnd.n3632 gnd.n3631 9.45567
R11148 gnd.n3600 gnd.n3599 9.45567
R11149 gnd.n3569 gnd.n3568 9.45567
R11150 gnd.n2737 gnd.n2736 9.39724
R11151 gnd.n3790 gnd.n3789 9.3005
R11152 gnd.n3763 gnd.n3762 9.3005
R11153 gnd.n3784 gnd.n3783 9.3005
R11154 gnd.n3782 gnd.n3781 9.3005
R11155 gnd.n3767 gnd.n3766 9.3005
R11156 gnd.n3776 gnd.n3775 9.3005
R11157 gnd.n3774 gnd.n3773 9.3005
R11158 gnd.n3758 gnd.n3757 9.3005
R11159 gnd.n3731 gnd.n3730 9.3005
R11160 gnd.n3752 gnd.n3751 9.3005
R11161 gnd.n3750 gnd.n3749 9.3005
R11162 gnd.n3735 gnd.n3734 9.3005
R11163 gnd.n3744 gnd.n3743 9.3005
R11164 gnd.n3742 gnd.n3741 9.3005
R11165 gnd.n3726 gnd.n3725 9.3005
R11166 gnd.n3699 gnd.n3698 9.3005
R11167 gnd.n3720 gnd.n3719 9.3005
R11168 gnd.n3718 gnd.n3717 9.3005
R11169 gnd.n3703 gnd.n3702 9.3005
R11170 gnd.n3712 gnd.n3711 9.3005
R11171 gnd.n3710 gnd.n3709 9.3005
R11172 gnd.n3695 gnd.n3694 9.3005
R11173 gnd.n3668 gnd.n3667 9.3005
R11174 gnd.n3689 gnd.n3688 9.3005
R11175 gnd.n3687 gnd.n3686 9.3005
R11176 gnd.n3672 gnd.n3671 9.3005
R11177 gnd.n3681 gnd.n3680 9.3005
R11178 gnd.n3679 gnd.n3678 9.3005
R11179 gnd.n3663 gnd.n3662 9.3005
R11180 gnd.n3636 gnd.n3635 9.3005
R11181 gnd.n3657 gnd.n3656 9.3005
R11182 gnd.n3655 gnd.n3654 9.3005
R11183 gnd.n3640 gnd.n3639 9.3005
R11184 gnd.n3649 gnd.n3648 9.3005
R11185 gnd.n3647 gnd.n3646 9.3005
R11186 gnd.n3631 gnd.n3630 9.3005
R11187 gnd.n3604 gnd.n3603 9.3005
R11188 gnd.n3625 gnd.n3624 9.3005
R11189 gnd.n3623 gnd.n3622 9.3005
R11190 gnd.n3608 gnd.n3607 9.3005
R11191 gnd.n3617 gnd.n3616 9.3005
R11192 gnd.n3615 gnd.n3614 9.3005
R11193 gnd.n3599 gnd.n3598 9.3005
R11194 gnd.n3572 gnd.n3571 9.3005
R11195 gnd.n3593 gnd.n3592 9.3005
R11196 gnd.n3591 gnd.n3590 9.3005
R11197 gnd.n3576 gnd.n3575 9.3005
R11198 gnd.n3585 gnd.n3584 9.3005
R11199 gnd.n3583 gnd.n3582 9.3005
R11200 gnd.n3568 gnd.n3567 9.3005
R11201 gnd.n3541 gnd.n3540 9.3005
R11202 gnd.n3562 gnd.n3561 9.3005
R11203 gnd.n3560 gnd.n3559 9.3005
R11204 gnd.n3545 gnd.n3544 9.3005
R11205 gnd.n3554 gnd.n3553 9.3005
R11206 gnd.n3552 gnd.n3551 9.3005
R11207 gnd.n3916 gnd.n3915 9.3005
R11208 gnd.n3914 gnd.n2483 9.3005
R11209 gnd.n3913 gnd.n3912 9.3005
R11210 gnd.n3909 gnd.n2484 9.3005
R11211 gnd.n3906 gnd.n2485 9.3005
R11212 gnd.n3905 gnd.n2486 9.3005
R11213 gnd.n3902 gnd.n2487 9.3005
R11214 gnd.n3901 gnd.n2488 9.3005
R11215 gnd.n3898 gnd.n2489 9.3005
R11216 gnd.n3897 gnd.n2490 9.3005
R11217 gnd.n3894 gnd.n2491 9.3005
R11218 gnd.n3893 gnd.n2492 9.3005
R11219 gnd.n3890 gnd.n2493 9.3005
R11220 gnd.n3889 gnd.n2494 9.3005
R11221 gnd.n3886 gnd.n3885 9.3005
R11222 gnd.n3884 gnd.n2495 9.3005
R11223 gnd.n3917 gnd.n2482 9.3005
R11224 gnd.n3158 gnd.n3157 9.3005
R11225 gnd.n2862 gnd.n2861 9.3005
R11226 gnd.n3185 gnd.n3184 9.3005
R11227 gnd.n3186 gnd.n2860 9.3005
R11228 gnd.n3190 gnd.n3187 9.3005
R11229 gnd.n3189 gnd.n3188 9.3005
R11230 gnd.n2834 gnd.n2833 9.3005
R11231 gnd.n3215 gnd.n3214 9.3005
R11232 gnd.n3216 gnd.n2832 9.3005
R11233 gnd.n3218 gnd.n3217 9.3005
R11234 gnd.n2812 gnd.n2811 9.3005
R11235 gnd.n3246 gnd.n3245 9.3005
R11236 gnd.n3247 gnd.n2810 9.3005
R11237 gnd.n3255 gnd.n3248 9.3005
R11238 gnd.n3254 gnd.n3249 9.3005
R11239 gnd.n3253 gnd.n3251 9.3005
R11240 gnd.n3250 gnd.n2759 9.3005
R11241 gnd.n3303 gnd.n2760 9.3005
R11242 gnd.n3302 gnd.n2761 9.3005
R11243 gnd.n3301 gnd.n2762 9.3005
R11244 gnd.n2781 gnd.n2763 9.3005
R11245 gnd.n2783 gnd.n2782 9.3005
R11246 gnd.n2681 gnd.n2680 9.3005
R11247 gnd.n3341 gnd.n3340 9.3005
R11248 gnd.n3342 gnd.n2679 9.3005
R11249 gnd.n3346 gnd.n3343 9.3005
R11250 gnd.n3345 gnd.n3344 9.3005
R11251 gnd.n2654 gnd.n2653 9.3005
R11252 gnd.n3381 gnd.n3380 9.3005
R11253 gnd.n3382 gnd.n2652 9.3005
R11254 gnd.n3386 gnd.n3383 9.3005
R11255 gnd.n3385 gnd.n3384 9.3005
R11256 gnd.n2627 gnd.n2626 9.3005
R11257 gnd.n3426 gnd.n3425 9.3005
R11258 gnd.n3427 gnd.n2625 9.3005
R11259 gnd.n3431 gnd.n3428 9.3005
R11260 gnd.n3430 gnd.n3429 9.3005
R11261 gnd.n2599 gnd.n2598 9.3005
R11262 gnd.n3466 gnd.n3465 9.3005
R11263 gnd.n3467 gnd.n2597 9.3005
R11264 gnd.n3471 gnd.n3468 9.3005
R11265 gnd.n3470 gnd.n3469 9.3005
R11266 gnd.n2571 gnd.n2570 9.3005
R11267 gnd.n3515 gnd.n3514 9.3005
R11268 gnd.n3516 gnd.n2569 9.3005
R11269 gnd.n3520 gnd.n3517 9.3005
R11270 gnd.n3519 gnd.n3518 9.3005
R11271 gnd.n2544 gnd.n2543 9.3005
R11272 gnd.n3809 gnd.n3808 9.3005
R11273 gnd.n3810 gnd.n2542 9.3005
R11274 gnd.n3816 gnd.n3811 9.3005
R11275 gnd.n3815 gnd.n3812 9.3005
R11276 gnd.n3814 gnd.n3813 9.3005
R11277 gnd.n3159 gnd.n3156 9.3005
R11278 gnd.n2941 gnd.n2900 9.3005
R11279 gnd.n2936 gnd.n2935 9.3005
R11280 gnd.n2934 gnd.n2901 9.3005
R11281 gnd.n2933 gnd.n2932 9.3005
R11282 gnd.n2929 gnd.n2902 9.3005
R11283 gnd.n2926 gnd.n2925 9.3005
R11284 gnd.n2924 gnd.n2903 9.3005
R11285 gnd.n2923 gnd.n2922 9.3005
R11286 gnd.n2919 gnd.n2904 9.3005
R11287 gnd.n2916 gnd.n2915 9.3005
R11288 gnd.n2914 gnd.n2905 9.3005
R11289 gnd.n2913 gnd.n2912 9.3005
R11290 gnd.n2909 gnd.n2907 9.3005
R11291 gnd.n2906 gnd.n2886 9.3005
R11292 gnd.n3153 gnd.n2885 9.3005
R11293 gnd.n3155 gnd.n3154 9.3005
R11294 gnd.n2943 gnd.n2942 9.3005
R11295 gnd.n3166 gnd.n2872 9.3005
R11296 gnd.n3173 gnd.n2873 9.3005
R11297 gnd.n3175 gnd.n3174 9.3005
R11298 gnd.n3176 gnd.n2853 9.3005
R11299 gnd.n3195 gnd.n3194 9.3005
R11300 gnd.n3197 gnd.n2845 9.3005
R11301 gnd.n3204 gnd.n2847 9.3005
R11302 gnd.n3205 gnd.n2842 9.3005
R11303 gnd.n3207 gnd.n3206 9.3005
R11304 gnd.n2843 gnd.n2828 9.3005
R11305 gnd.n3223 gnd.n2826 9.3005
R11306 gnd.n3227 gnd.n3226 9.3005
R11307 gnd.n3225 gnd.n2802 9.3005
R11308 gnd.n3262 gnd.n2801 9.3005
R11309 gnd.n3265 gnd.n3264 9.3005
R11310 gnd.n2798 gnd.n2797 9.3005
R11311 gnd.n3271 gnd.n2799 9.3005
R11312 gnd.n3273 gnd.n3272 9.3005
R11313 gnd.n3275 gnd.n2796 9.3005
R11314 gnd.n3278 gnd.n3277 9.3005
R11315 gnd.n3281 gnd.n3279 9.3005
R11316 gnd.n3283 gnd.n3282 9.3005
R11317 gnd.n3289 gnd.n3284 9.3005
R11318 gnd.n3288 gnd.n3287 9.3005
R11319 gnd.n2672 gnd.n2671 9.3005
R11320 gnd.n3355 gnd.n3354 9.3005
R11321 gnd.n3356 gnd.n2665 9.3005
R11322 gnd.n3364 gnd.n2664 9.3005
R11323 gnd.n3367 gnd.n3366 9.3005
R11324 gnd.n3369 gnd.n3368 9.3005
R11325 gnd.n3372 gnd.n2647 9.3005
R11326 gnd.n3370 gnd.n2645 9.3005
R11327 gnd.n3392 gnd.n2643 9.3005
R11328 gnd.n3394 gnd.n3393 9.3005
R11329 gnd.n2617 gnd.n2616 9.3005
R11330 gnd.n3440 gnd.n3439 9.3005
R11331 gnd.n3441 gnd.n2610 9.3005
R11332 gnd.n3449 gnd.n2609 9.3005
R11333 gnd.n3452 gnd.n3451 9.3005
R11334 gnd.n3454 gnd.n3453 9.3005
R11335 gnd.n3457 gnd.n2592 9.3005
R11336 gnd.n3455 gnd.n2590 9.3005
R11337 gnd.n3477 gnd.n2588 9.3005
R11338 gnd.n3479 gnd.n3478 9.3005
R11339 gnd.n2562 gnd.n2561 9.3005
R11340 gnd.n3529 gnd.n3528 9.3005
R11341 gnd.n3530 gnd.n2555 9.3005
R11342 gnd.n3538 gnd.n2554 9.3005
R11343 gnd.n3797 gnd.n3796 9.3005
R11344 gnd.n3799 gnd.n3798 9.3005
R11345 gnd.n3800 gnd.n2535 9.3005
R11346 gnd.n3824 gnd.n3823 9.3005
R11347 gnd.n2536 gnd.n2498 9.3005
R11348 gnd.n3164 gnd.n3163 9.3005
R11349 gnd.n3880 gnd.n2499 9.3005
R11350 gnd.n3879 gnd.n2501 9.3005
R11351 gnd.n3876 gnd.n2502 9.3005
R11352 gnd.n3875 gnd.n2503 9.3005
R11353 gnd.n3872 gnd.n2504 9.3005
R11354 gnd.n3871 gnd.n2505 9.3005
R11355 gnd.n3868 gnd.n2506 9.3005
R11356 gnd.n3867 gnd.n2507 9.3005
R11357 gnd.n3864 gnd.n2508 9.3005
R11358 gnd.n3863 gnd.n2509 9.3005
R11359 gnd.n3860 gnd.n2510 9.3005
R11360 gnd.n3859 gnd.n2511 9.3005
R11361 gnd.n3856 gnd.n2512 9.3005
R11362 gnd.n3855 gnd.n2513 9.3005
R11363 gnd.n3852 gnd.n2514 9.3005
R11364 gnd.n3851 gnd.n2515 9.3005
R11365 gnd.n3848 gnd.n2516 9.3005
R11366 gnd.n3847 gnd.n2517 9.3005
R11367 gnd.n3844 gnd.n2518 9.3005
R11368 gnd.n3843 gnd.n2519 9.3005
R11369 gnd.n3840 gnd.n2520 9.3005
R11370 gnd.n3839 gnd.n2521 9.3005
R11371 gnd.n3836 gnd.n2525 9.3005
R11372 gnd.n3835 gnd.n2526 9.3005
R11373 gnd.n3832 gnd.n2527 9.3005
R11374 gnd.n3831 gnd.n2528 9.3005
R11375 gnd.n3882 gnd.n3881 9.3005
R11376 gnd.n3333 gnd.n3317 9.3005
R11377 gnd.n3332 gnd.n3318 9.3005
R11378 gnd.n3331 gnd.n3319 9.3005
R11379 gnd.n3329 gnd.n3320 9.3005
R11380 gnd.n3328 gnd.n3321 9.3005
R11381 gnd.n3326 gnd.n3322 9.3005
R11382 gnd.n3325 gnd.n3323 9.3005
R11383 gnd.n2635 gnd.n2634 9.3005
R11384 gnd.n3402 gnd.n3401 9.3005
R11385 gnd.n3403 gnd.n2633 9.3005
R11386 gnd.n3420 gnd.n3404 9.3005
R11387 gnd.n3419 gnd.n3405 9.3005
R11388 gnd.n3418 gnd.n3406 9.3005
R11389 gnd.n3416 gnd.n3407 9.3005
R11390 gnd.n3415 gnd.n3408 9.3005
R11391 gnd.n3413 gnd.n3409 9.3005
R11392 gnd.n3412 gnd.n3410 9.3005
R11393 gnd.n2579 gnd.n2578 9.3005
R11394 gnd.n3487 gnd.n3486 9.3005
R11395 gnd.n3488 gnd.n2577 9.3005
R11396 gnd.n3509 gnd.n3489 9.3005
R11397 gnd.n3508 gnd.n3490 9.3005
R11398 gnd.n3507 gnd.n3491 9.3005
R11399 gnd.n3504 gnd.n3492 9.3005
R11400 gnd.n3503 gnd.n3493 9.3005
R11401 gnd.n3501 gnd.n3494 9.3005
R11402 gnd.n3500 gnd.n3495 9.3005
R11403 gnd.n3498 gnd.n3497 9.3005
R11404 gnd.n3496 gnd.n2530 9.3005
R11405 gnd.n3074 gnd.n3073 9.3005
R11406 gnd.n2964 gnd.n2963 9.3005
R11407 gnd.n3088 gnd.n3087 9.3005
R11408 gnd.n3089 gnd.n2962 9.3005
R11409 gnd.n3091 gnd.n3090 9.3005
R11410 gnd.n2952 gnd.n2951 9.3005
R11411 gnd.n3104 gnd.n3103 9.3005
R11412 gnd.n3105 gnd.n2950 9.3005
R11413 gnd.n3137 gnd.n3106 9.3005
R11414 gnd.n3136 gnd.n3107 9.3005
R11415 gnd.n3135 gnd.n3108 9.3005
R11416 gnd.n3134 gnd.n3109 9.3005
R11417 gnd.n3131 gnd.n3110 9.3005
R11418 gnd.n3130 gnd.n3111 9.3005
R11419 gnd.n3129 gnd.n3112 9.3005
R11420 gnd.n3127 gnd.n3113 9.3005
R11421 gnd.n3126 gnd.n3114 9.3005
R11422 gnd.n3123 gnd.n3115 9.3005
R11423 gnd.n3122 gnd.n3116 9.3005
R11424 gnd.n3121 gnd.n3117 9.3005
R11425 gnd.n3119 gnd.n3118 9.3005
R11426 gnd.n2818 gnd.n2817 9.3005
R11427 gnd.n3235 gnd.n3234 9.3005
R11428 gnd.n3236 gnd.n2816 9.3005
R11429 gnd.n3240 gnd.n3237 9.3005
R11430 gnd.n3239 gnd.n3238 9.3005
R11431 gnd.n2740 gnd.n2739 9.3005
R11432 gnd.n3315 gnd.n3314 9.3005
R11433 gnd.n3072 gnd.n2973 9.3005
R11434 gnd.n2975 gnd.n2974 9.3005
R11435 gnd.n3019 gnd.n3017 9.3005
R11436 gnd.n3020 gnd.n3016 9.3005
R11437 gnd.n3023 gnd.n3012 9.3005
R11438 gnd.n3024 gnd.n3011 9.3005
R11439 gnd.n3027 gnd.n3010 9.3005
R11440 gnd.n3028 gnd.n3009 9.3005
R11441 gnd.n3031 gnd.n3008 9.3005
R11442 gnd.n3032 gnd.n3007 9.3005
R11443 gnd.n3035 gnd.n3006 9.3005
R11444 gnd.n3036 gnd.n3005 9.3005
R11445 gnd.n3039 gnd.n3004 9.3005
R11446 gnd.n3040 gnd.n3003 9.3005
R11447 gnd.n3043 gnd.n3002 9.3005
R11448 gnd.n3044 gnd.n3001 9.3005
R11449 gnd.n3047 gnd.n3000 9.3005
R11450 gnd.n3048 gnd.n2999 9.3005
R11451 gnd.n3051 gnd.n2998 9.3005
R11452 gnd.n3052 gnd.n2997 9.3005
R11453 gnd.n3055 gnd.n2996 9.3005
R11454 gnd.n3056 gnd.n2995 9.3005
R11455 gnd.n3059 gnd.n2994 9.3005
R11456 gnd.n3061 gnd.n2993 9.3005
R11457 gnd.n3062 gnd.n2992 9.3005
R11458 gnd.n3063 gnd.n2991 9.3005
R11459 gnd.n3064 gnd.n2990 9.3005
R11460 gnd.n3071 gnd.n3070 9.3005
R11461 gnd.n3080 gnd.n3079 9.3005
R11462 gnd.n3081 gnd.n2967 9.3005
R11463 gnd.n3083 gnd.n3082 9.3005
R11464 gnd.n2958 gnd.n2957 9.3005
R11465 gnd.n3096 gnd.n3095 9.3005
R11466 gnd.n3097 gnd.n2956 9.3005
R11467 gnd.n3099 gnd.n3098 9.3005
R11468 gnd.n2945 gnd.n2944 9.3005
R11469 gnd.n3142 gnd.n3141 9.3005
R11470 gnd.n3143 gnd.n2899 9.3005
R11471 gnd.n3147 gnd.n3145 9.3005
R11472 gnd.n3146 gnd.n2878 9.3005
R11473 gnd.n3165 gnd.n2877 9.3005
R11474 gnd.n3168 gnd.n3167 9.3005
R11475 gnd.n2871 gnd.n2870 9.3005
R11476 gnd.n3179 gnd.n3177 9.3005
R11477 gnd.n3178 gnd.n2852 9.3005
R11478 gnd.n3196 gnd.n2851 9.3005
R11479 gnd.n3199 gnd.n3198 9.3005
R11480 gnd.n2846 gnd.n2841 9.3005
R11481 gnd.n3209 gnd.n3208 9.3005
R11482 gnd.n2844 gnd.n2824 9.3005
R11483 gnd.n3230 gnd.n2825 9.3005
R11484 gnd.n3229 gnd.n3228 9.3005
R11485 gnd.n2827 gnd.n2803 9.3005
R11486 gnd.n3261 gnd.n3260 9.3005
R11487 gnd.n3263 gnd.n2748 9.3005
R11488 gnd.n3310 gnd.n2749 9.3005
R11489 gnd.n3309 gnd.n2750 9.3005
R11490 gnd.n3308 gnd.n2751 9.3005
R11491 gnd.n3274 gnd.n2752 9.3005
R11492 gnd.n3276 gnd.n2770 9.3005
R11493 gnd.n3296 gnd.n2771 9.3005
R11494 gnd.n3295 gnd.n2772 9.3005
R11495 gnd.n3294 gnd.n2773 9.3005
R11496 gnd.n3285 gnd.n2774 9.3005
R11497 gnd.n3286 gnd.n2673 9.3005
R11498 gnd.n3352 gnd.n3351 9.3005
R11499 gnd.n3353 gnd.n2666 9.3005
R11500 gnd.n3363 gnd.n3362 9.3005
R11501 gnd.n3365 gnd.n2662 9.3005
R11502 gnd.n3375 gnd.n2663 9.3005
R11503 gnd.n3374 gnd.n3373 9.3005
R11504 gnd.n3371 gnd.n2641 9.3005
R11505 gnd.n3397 gnd.n2642 9.3005
R11506 gnd.n3396 gnd.n3395 9.3005
R11507 gnd.n2644 gnd.n2618 9.3005
R11508 gnd.n3437 gnd.n3436 9.3005
R11509 gnd.n3438 gnd.n2611 9.3005
R11510 gnd.n3448 gnd.n3447 9.3005
R11511 gnd.n3450 gnd.n2607 9.3005
R11512 gnd.n3460 gnd.n2608 9.3005
R11513 gnd.n3459 gnd.n3458 9.3005
R11514 gnd.n3456 gnd.n2586 9.3005
R11515 gnd.n3482 gnd.n2587 9.3005
R11516 gnd.n3481 gnd.n3480 9.3005
R11517 gnd.n2589 gnd.n2563 9.3005
R11518 gnd.n3526 gnd.n3525 9.3005
R11519 gnd.n3527 gnd.n2556 9.3005
R11520 gnd.n3537 gnd.n3536 9.3005
R11521 gnd.n3795 gnd.n2552 9.3005
R11522 gnd.n3803 gnd.n2553 9.3005
R11523 gnd.n3802 gnd.n3801 9.3005
R11524 gnd.n2534 gnd.n2533 9.3005
R11525 gnd.n3826 gnd.n3825 9.3005
R11526 gnd.n2969 gnd.n2968 9.3005
R11527 gnd.n6193 gnd.n939 9.3005
R11528 gnd.n6195 gnd.n6194 9.3005
R11529 gnd.n935 gnd.n934 9.3005
R11530 gnd.n6202 gnd.n6201 9.3005
R11531 gnd.n6203 gnd.n933 9.3005
R11532 gnd.n6205 gnd.n6204 9.3005
R11533 gnd.n929 gnd.n928 9.3005
R11534 gnd.n6212 gnd.n6211 9.3005
R11535 gnd.n6213 gnd.n927 9.3005
R11536 gnd.n6215 gnd.n6214 9.3005
R11537 gnd.n923 gnd.n922 9.3005
R11538 gnd.n6222 gnd.n6221 9.3005
R11539 gnd.n6223 gnd.n921 9.3005
R11540 gnd.n6225 gnd.n6224 9.3005
R11541 gnd.n917 gnd.n916 9.3005
R11542 gnd.n6232 gnd.n6231 9.3005
R11543 gnd.n6233 gnd.n915 9.3005
R11544 gnd.n6235 gnd.n6234 9.3005
R11545 gnd.n911 gnd.n910 9.3005
R11546 gnd.n6242 gnd.n6241 9.3005
R11547 gnd.n6243 gnd.n909 9.3005
R11548 gnd.n6245 gnd.n6244 9.3005
R11549 gnd.n905 gnd.n904 9.3005
R11550 gnd.n6252 gnd.n6251 9.3005
R11551 gnd.n6253 gnd.n903 9.3005
R11552 gnd.n6255 gnd.n6254 9.3005
R11553 gnd.n899 gnd.n898 9.3005
R11554 gnd.n6262 gnd.n6261 9.3005
R11555 gnd.n6263 gnd.n897 9.3005
R11556 gnd.n6265 gnd.n6264 9.3005
R11557 gnd.n893 gnd.n892 9.3005
R11558 gnd.n6272 gnd.n6271 9.3005
R11559 gnd.n6273 gnd.n891 9.3005
R11560 gnd.n6275 gnd.n6274 9.3005
R11561 gnd.n887 gnd.n886 9.3005
R11562 gnd.n6282 gnd.n6281 9.3005
R11563 gnd.n6283 gnd.n885 9.3005
R11564 gnd.n6285 gnd.n6284 9.3005
R11565 gnd.n881 gnd.n880 9.3005
R11566 gnd.n6292 gnd.n6291 9.3005
R11567 gnd.n6293 gnd.n879 9.3005
R11568 gnd.n6295 gnd.n6294 9.3005
R11569 gnd.n875 gnd.n874 9.3005
R11570 gnd.n6302 gnd.n6301 9.3005
R11571 gnd.n6303 gnd.n873 9.3005
R11572 gnd.n6305 gnd.n6304 9.3005
R11573 gnd.n869 gnd.n868 9.3005
R11574 gnd.n6312 gnd.n6311 9.3005
R11575 gnd.n6313 gnd.n867 9.3005
R11576 gnd.n6315 gnd.n6314 9.3005
R11577 gnd.n863 gnd.n862 9.3005
R11578 gnd.n6322 gnd.n6321 9.3005
R11579 gnd.n6323 gnd.n861 9.3005
R11580 gnd.n6325 gnd.n6324 9.3005
R11581 gnd.n857 gnd.n856 9.3005
R11582 gnd.n6332 gnd.n6331 9.3005
R11583 gnd.n6333 gnd.n855 9.3005
R11584 gnd.n6335 gnd.n6334 9.3005
R11585 gnd.n851 gnd.n850 9.3005
R11586 gnd.n6342 gnd.n6341 9.3005
R11587 gnd.n6343 gnd.n849 9.3005
R11588 gnd.n6345 gnd.n6344 9.3005
R11589 gnd.n845 gnd.n844 9.3005
R11590 gnd.n6352 gnd.n6351 9.3005
R11591 gnd.n6353 gnd.n843 9.3005
R11592 gnd.n6355 gnd.n6354 9.3005
R11593 gnd.n839 gnd.n838 9.3005
R11594 gnd.n6362 gnd.n6361 9.3005
R11595 gnd.n6363 gnd.n837 9.3005
R11596 gnd.n6365 gnd.n6364 9.3005
R11597 gnd.n833 gnd.n832 9.3005
R11598 gnd.n6372 gnd.n6371 9.3005
R11599 gnd.n6373 gnd.n831 9.3005
R11600 gnd.n6375 gnd.n6374 9.3005
R11601 gnd.n827 gnd.n826 9.3005
R11602 gnd.n6382 gnd.n6381 9.3005
R11603 gnd.n6383 gnd.n825 9.3005
R11604 gnd.n6385 gnd.n6384 9.3005
R11605 gnd.n821 gnd.n820 9.3005
R11606 gnd.n6392 gnd.n6391 9.3005
R11607 gnd.n6393 gnd.n819 9.3005
R11608 gnd.n6395 gnd.n6394 9.3005
R11609 gnd.n815 gnd.n814 9.3005
R11610 gnd.n6402 gnd.n6401 9.3005
R11611 gnd.n6403 gnd.n813 9.3005
R11612 gnd.n6405 gnd.n6404 9.3005
R11613 gnd.n809 gnd.n808 9.3005
R11614 gnd.n6412 gnd.n6411 9.3005
R11615 gnd.n6413 gnd.n807 9.3005
R11616 gnd.n6415 gnd.n6414 9.3005
R11617 gnd.n803 gnd.n802 9.3005
R11618 gnd.n6422 gnd.n6421 9.3005
R11619 gnd.n6423 gnd.n801 9.3005
R11620 gnd.n6425 gnd.n6424 9.3005
R11621 gnd.n797 gnd.n796 9.3005
R11622 gnd.n6432 gnd.n6431 9.3005
R11623 gnd.n6433 gnd.n795 9.3005
R11624 gnd.n6435 gnd.n6434 9.3005
R11625 gnd.n791 gnd.n790 9.3005
R11626 gnd.n6442 gnd.n6441 9.3005
R11627 gnd.n6443 gnd.n789 9.3005
R11628 gnd.n6445 gnd.n6444 9.3005
R11629 gnd.n785 gnd.n784 9.3005
R11630 gnd.n6452 gnd.n6451 9.3005
R11631 gnd.n6453 gnd.n783 9.3005
R11632 gnd.n6455 gnd.n6454 9.3005
R11633 gnd.n779 gnd.n778 9.3005
R11634 gnd.n6462 gnd.n6461 9.3005
R11635 gnd.n6463 gnd.n777 9.3005
R11636 gnd.n6465 gnd.n6464 9.3005
R11637 gnd.n773 gnd.n772 9.3005
R11638 gnd.n6472 gnd.n6471 9.3005
R11639 gnd.n6473 gnd.n771 9.3005
R11640 gnd.n6475 gnd.n6474 9.3005
R11641 gnd.n767 gnd.n766 9.3005
R11642 gnd.n6482 gnd.n6481 9.3005
R11643 gnd.n6483 gnd.n765 9.3005
R11644 gnd.n6485 gnd.n6484 9.3005
R11645 gnd.n761 gnd.n760 9.3005
R11646 gnd.n6492 gnd.n6491 9.3005
R11647 gnd.n6493 gnd.n759 9.3005
R11648 gnd.n6495 gnd.n6494 9.3005
R11649 gnd.n755 gnd.n754 9.3005
R11650 gnd.n6502 gnd.n6501 9.3005
R11651 gnd.n6503 gnd.n753 9.3005
R11652 gnd.n6505 gnd.n6504 9.3005
R11653 gnd.n749 gnd.n748 9.3005
R11654 gnd.n6512 gnd.n6511 9.3005
R11655 gnd.n6513 gnd.n747 9.3005
R11656 gnd.n6515 gnd.n6514 9.3005
R11657 gnd.n743 gnd.n742 9.3005
R11658 gnd.n6522 gnd.n6521 9.3005
R11659 gnd.n6523 gnd.n741 9.3005
R11660 gnd.n6525 gnd.n6524 9.3005
R11661 gnd.n737 gnd.n736 9.3005
R11662 gnd.n6532 gnd.n6531 9.3005
R11663 gnd.n6533 gnd.n735 9.3005
R11664 gnd.n6535 gnd.n6534 9.3005
R11665 gnd.n731 gnd.n730 9.3005
R11666 gnd.n6542 gnd.n6541 9.3005
R11667 gnd.n6543 gnd.n729 9.3005
R11668 gnd.n6545 gnd.n6544 9.3005
R11669 gnd.n725 gnd.n724 9.3005
R11670 gnd.n6552 gnd.n6551 9.3005
R11671 gnd.n6553 gnd.n723 9.3005
R11672 gnd.n6555 gnd.n6554 9.3005
R11673 gnd.n719 gnd.n718 9.3005
R11674 gnd.n6562 gnd.n6561 9.3005
R11675 gnd.n6563 gnd.n717 9.3005
R11676 gnd.n6565 gnd.n6564 9.3005
R11677 gnd.n713 gnd.n712 9.3005
R11678 gnd.n6572 gnd.n6571 9.3005
R11679 gnd.n6573 gnd.n711 9.3005
R11680 gnd.n6575 gnd.n6574 9.3005
R11681 gnd.n707 gnd.n706 9.3005
R11682 gnd.n6582 gnd.n6581 9.3005
R11683 gnd.n6583 gnd.n705 9.3005
R11684 gnd.n6585 gnd.n6584 9.3005
R11685 gnd.n701 gnd.n700 9.3005
R11686 gnd.n6592 gnd.n6591 9.3005
R11687 gnd.n6593 gnd.n699 9.3005
R11688 gnd.n6595 gnd.n6594 9.3005
R11689 gnd.n695 gnd.n694 9.3005
R11690 gnd.n6602 gnd.n6601 9.3005
R11691 gnd.n6603 gnd.n693 9.3005
R11692 gnd.n6605 gnd.n6604 9.3005
R11693 gnd.n689 gnd.n688 9.3005
R11694 gnd.n6612 gnd.n6611 9.3005
R11695 gnd.n6615 gnd.n6614 9.3005
R11696 gnd.n683 gnd.n682 9.3005
R11697 gnd.n6622 gnd.n6621 9.3005
R11698 gnd.n6623 gnd.n681 9.3005
R11699 gnd.n6625 gnd.n6624 9.3005
R11700 gnd.n677 gnd.n676 9.3005
R11701 gnd.n6632 gnd.n6631 9.3005
R11702 gnd.n6633 gnd.n675 9.3005
R11703 gnd.n6635 gnd.n6634 9.3005
R11704 gnd.n671 gnd.n670 9.3005
R11705 gnd.n6642 gnd.n6641 9.3005
R11706 gnd.n6643 gnd.n669 9.3005
R11707 gnd.n6645 gnd.n6644 9.3005
R11708 gnd.n665 gnd.n664 9.3005
R11709 gnd.n6652 gnd.n6651 9.3005
R11710 gnd.n6653 gnd.n663 9.3005
R11711 gnd.n6655 gnd.n6654 9.3005
R11712 gnd.n659 gnd.n658 9.3005
R11713 gnd.n6662 gnd.n6661 9.3005
R11714 gnd.n6663 gnd.n657 9.3005
R11715 gnd.n6665 gnd.n6664 9.3005
R11716 gnd.n653 gnd.n652 9.3005
R11717 gnd.n6672 gnd.n6671 9.3005
R11718 gnd.n6673 gnd.n651 9.3005
R11719 gnd.n6675 gnd.n6674 9.3005
R11720 gnd.n647 gnd.n646 9.3005
R11721 gnd.n6682 gnd.n6681 9.3005
R11722 gnd.n6683 gnd.n645 9.3005
R11723 gnd.n6685 gnd.n6684 9.3005
R11724 gnd.n641 gnd.n640 9.3005
R11725 gnd.n6692 gnd.n6691 9.3005
R11726 gnd.n6693 gnd.n639 9.3005
R11727 gnd.n6695 gnd.n6694 9.3005
R11728 gnd.n635 gnd.n634 9.3005
R11729 gnd.n6702 gnd.n6701 9.3005
R11730 gnd.n6703 gnd.n633 9.3005
R11731 gnd.n6705 gnd.n6704 9.3005
R11732 gnd.n629 gnd.n628 9.3005
R11733 gnd.n6712 gnd.n6711 9.3005
R11734 gnd.n6713 gnd.n627 9.3005
R11735 gnd.n6715 gnd.n6714 9.3005
R11736 gnd.n623 gnd.n622 9.3005
R11737 gnd.n6722 gnd.n6721 9.3005
R11738 gnd.n6723 gnd.n621 9.3005
R11739 gnd.n6725 gnd.n6724 9.3005
R11740 gnd.n617 gnd.n616 9.3005
R11741 gnd.n6732 gnd.n6731 9.3005
R11742 gnd.n6733 gnd.n615 9.3005
R11743 gnd.n6735 gnd.n6734 9.3005
R11744 gnd.n611 gnd.n610 9.3005
R11745 gnd.n6742 gnd.n6741 9.3005
R11746 gnd.n6743 gnd.n609 9.3005
R11747 gnd.n6745 gnd.n6744 9.3005
R11748 gnd.n605 gnd.n604 9.3005
R11749 gnd.n6752 gnd.n6751 9.3005
R11750 gnd.n6753 gnd.n603 9.3005
R11751 gnd.n6755 gnd.n6754 9.3005
R11752 gnd.n599 gnd.n598 9.3005
R11753 gnd.n6762 gnd.n6761 9.3005
R11754 gnd.n6763 gnd.n597 9.3005
R11755 gnd.n6765 gnd.n6764 9.3005
R11756 gnd.n593 gnd.n592 9.3005
R11757 gnd.n6772 gnd.n6771 9.3005
R11758 gnd.n6773 gnd.n591 9.3005
R11759 gnd.n6775 gnd.n6774 9.3005
R11760 gnd.n587 gnd.n586 9.3005
R11761 gnd.n6782 gnd.n6781 9.3005
R11762 gnd.n6783 gnd.n585 9.3005
R11763 gnd.n6785 gnd.n6784 9.3005
R11764 gnd.n581 gnd.n580 9.3005
R11765 gnd.n6792 gnd.n6791 9.3005
R11766 gnd.n6793 gnd.n579 9.3005
R11767 gnd.n6795 gnd.n6794 9.3005
R11768 gnd.n575 gnd.n574 9.3005
R11769 gnd.n6802 gnd.n6801 9.3005
R11770 gnd.n6803 gnd.n573 9.3005
R11771 gnd.n6805 gnd.n6804 9.3005
R11772 gnd.n569 gnd.n568 9.3005
R11773 gnd.n6812 gnd.n6811 9.3005
R11774 gnd.n6813 gnd.n567 9.3005
R11775 gnd.n6817 gnd.n6814 9.3005
R11776 gnd.n6816 gnd.n6815 9.3005
R11777 gnd.n563 gnd.n562 9.3005
R11778 gnd.n6825 gnd.n6824 9.3005
R11779 gnd.n6613 gnd.n687 9.3005
R11780 gnd.n7321 gnd.n108 9.3005
R11781 gnd.n7320 gnd.n110 9.3005
R11782 gnd.n114 gnd.n111 9.3005
R11783 gnd.n7315 gnd.n115 9.3005
R11784 gnd.n7314 gnd.n116 9.3005
R11785 gnd.n7313 gnd.n117 9.3005
R11786 gnd.n121 gnd.n118 9.3005
R11787 gnd.n7308 gnd.n122 9.3005
R11788 gnd.n7307 gnd.n123 9.3005
R11789 gnd.n7306 gnd.n124 9.3005
R11790 gnd.n128 gnd.n125 9.3005
R11791 gnd.n7301 gnd.n129 9.3005
R11792 gnd.n7300 gnd.n130 9.3005
R11793 gnd.n7299 gnd.n131 9.3005
R11794 gnd.n135 gnd.n132 9.3005
R11795 gnd.n7294 gnd.n136 9.3005
R11796 gnd.n7293 gnd.n137 9.3005
R11797 gnd.n7289 gnd.n138 9.3005
R11798 gnd.n142 gnd.n139 9.3005
R11799 gnd.n7284 gnd.n143 9.3005
R11800 gnd.n7283 gnd.n144 9.3005
R11801 gnd.n7282 gnd.n145 9.3005
R11802 gnd.n149 gnd.n146 9.3005
R11803 gnd.n7277 gnd.n150 9.3005
R11804 gnd.n7276 gnd.n151 9.3005
R11805 gnd.n7275 gnd.n152 9.3005
R11806 gnd.n156 gnd.n153 9.3005
R11807 gnd.n7270 gnd.n157 9.3005
R11808 gnd.n7269 gnd.n158 9.3005
R11809 gnd.n7268 gnd.n159 9.3005
R11810 gnd.n163 gnd.n160 9.3005
R11811 gnd.n7263 gnd.n164 9.3005
R11812 gnd.n7262 gnd.n165 9.3005
R11813 gnd.n7261 gnd.n166 9.3005
R11814 gnd.n170 gnd.n167 9.3005
R11815 gnd.n7256 gnd.n171 9.3005
R11816 gnd.n7255 gnd.n7254 9.3005
R11817 gnd.n7253 gnd.n174 9.3005
R11818 gnd.n7323 gnd.n7322 9.3005
R11819 gnd.n5465 gnd.n5464 9.3005
R11820 gnd.n5614 gnd.n5466 9.3005
R11821 gnd.n5613 gnd.n5467 9.3005
R11822 gnd.n5612 gnd.n5468 9.3005
R11823 gnd.n5609 gnd.n5469 9.3005
R11824 gnd.n5608 gnd.n5470 9.3005
R11825 gnd.n5605 gnd.n5471 9.3005
R11826 gnd.n5604 gnd.n5472 9.3005
R11827 gnd.n5601 gnd.n5473 9.3005
R11828 gnd.n5600 gnd.n5474 9.3005
R11829 gnd.n5511 gnd.n5475 9.3005
R11830 gnd.n5515 gnd.n5514 9.3005
R11831 gnd.n5516 gnd.n5510 9.3005
R11832 gnd.n5520 gnd.n5517 9.3005
R11833 gnd.n5521 gnd.n5509 9.3005
R11834 gnd.n5525 gnd.n5524 9.3005
R11835 gnd.n5526 gnd.n5508 9.3005
R11836 gnd.n5580 gnd.n5527 9.3005
R11837 gnd.n5579 gnd.n5528 9.3005
R11838 gnd.n5578 gnd.n5529 9.3005
R11839 gnd.n5548 gnd.n5530 9.3005
R11840 gnd.n5549 gnd.n5547 9.3005
R11841 gnd.n5552 gnd.n5551 9.3005
R11842 gnd.n5550 gnd.n495 9.3005
R11843 gnd.n6849 gnd.n496 9.3005
R11844 gnd.n6848 gnd.n497 9.3005
R11845 gnd.n6847 gnd.n498 9.3005
R11846 gnd.n6844 gnd.n499 9.3005
R11847 gnd.n6843 gnd.n500 9.3005
R11848 gnd.n6840 gnd.n501 9.3005
R11849 gnd.n6839 gnd.n502 9.3005
R11850 gnd.n552 gnd.n503 9.3005
R11851 gnd.n551 gnd.n504 9.3005
R11852 gnd.n548 gnd.n505 9.3005
R11853 gnd.n547 gnd.n506 9.3005
R11854 gnd.n544 gnd.n507 9.3005
R11855 gnd.n543 gnd.n508 9.3005
R11856 gnd.n541 gnd.n509 9.3005
R11857 gnd.n540 gnd.n510 9.3005
R11858 gnd.n538 gnd.n511 9.3005
R11859 gnd.n537 gnd.n512 9.3005
R11860 gnd.n535 gnd.n513 9.3005
R11861 gnd.n534 gnd.n514 9.3005
R11862 gnd.n532 gnd.n515 9.3005
R11863 gnd.n531 gnd.n516 9.3005
R11864 gnd.n529 gnd.n517 9.3005
R11865 gnd.n528 gnd.n518 9.3005
R11866 gnd.n526 gnd.n519 9.3005
R11867 gnd.n525 gnd.n520 9.3005
R11868 gnd.n523 gnd.n522 9.3005
R11869 gnd.n521 gnd.n178 9.3005
R11870 gnd.n7250 gnd.n177 9.3005
R11871 gnd.n7252 gnd.n7251 9.3005
R11872 gnd.n469 gnd.n468 9.3005
R11873 gnd.n6901 gnd.n6900 9.3005
R11874 gnd.n6902 gnd.n462 9.3005
R11875 gnd.n6905 gnd.n461 9.3005
R11876 gnd.n6906 gnd.n460 9.3005
R11877 gnd.n6909 gnd.n459 9.3005
R11878 gnd.n6910 gnd.n458 9.3005
R11879 gnd.n6913 gnd.n457 9.3005
R11880 gnd.n6914 gnd.n456 9.3005
R11881 gnd.n6917 gnd.n455 9.3005
R11882 gnd.n6918 gnd.n454 9.3005
R11883 gnd.n6921 gnd.n453 9.3005
R11884 gnd.n6922 gnd.n452 9.3005
R11885 gnd.n6925 gnd.n451 9.3005
R11886 gnd.n6926 gnd.n450 9.3005
R11887 gnd.n6929 gnd.n449 9.3005
R11888 gnd.n6930 gnd.n448 9.3005
R11889 gnd.n6933 gnd.n447 9.3005
R11890 gnd.n6934 gnd.n446 9.3005
R11891 gnd.n6937 gnd.n445 9.3005
R11892 gnd.n6939 gnd.n439 9.3005
R11893 gnd.n6942 gnd.n438 9.3005
R11894 gnd.n6943 gnd.n437 9.3005
R11895 gnd.n6946 gnd.n436 9.3005
R11896 gnd.n6947 gnd.n435 9.3005
R11897 gnd.n6950 gnd.n434 9.3005
R11898 gnd.n6951 gnd.n433 9.3005
R11899 gnd.n6954 gnd.n432 9.3005
R11900 gnd.n6955 gnd.n431 9.3005
R11901 gnd.n6958 gnd.n430 9.3005
R11902 gnd.n6959 gnd.n429 9.3005
R11903 gnd.n6962 gnd.n428 9.3005
R11904 gnd.n6963 gnd.n427 9.3005
R11905 gnd.n6964 gnd.n426 9.3005
R11906 gnd.n393 gnd.n392 9.3005
R11907 gnd.n6970 gnd.n6969 9.3005
R11908 gnd.n6899 gnd.n467 9.3005
R11909 gnd.n6898 gnd.n6897 9.3005
R11910 gnd.n6973 gnd.n6972 9.3005
R11911 gnd.n376 gnd.n375 9.3005
R11912 gnd.n6986 gnd.n6985 9.3005
R11913 gnd.n6987 gnd.n374 9.3005
R11914 gnd.n6989 gnd.n6988 9.3005
R11915 gnd.n358 gnd.n357 9.3005
R11916 gnd.n7002 gnd.n7001 9.3005
R11917 gnd.n7003 gnd.n356 9.3005
R11918 gnd.n7005 gnd.n7004 9.3005
R11919 gnd.n341 gnd.n340 9.3005
R11920 gnd.n7018 gnd.n7017 9.3005
R11921 gnd.n7019 gnd.n339 9.3005
R11922 gnd.n7021 gnd.n7020 9.3005
R11923 gnd.n323 gnd.n322 9.3005
R11924 gnd.n7034 gnd.n7033 9.3005
R11925 gnd.n7035 gnd.n321 9.3005
R11926 gnd.n7037 gnd.n7036 9.3005
R11927 gnd.n303 gnd.n302 9.3005
R11928 gnd.n7051 gnd.n7050 9.3005
R11929 gnd.n7052 gnd.n301 9.3005
R11930 gnd.n7054 gnd.n7053 9.3005
R11931 gnd.n7101 gnd.n7100 9.3005
R11932 gnd.n7102 gnd.n254 9.3005
R11933 gnd.n7104 gnd.n7103 9.3005
R11934 gnd.n239 gnd.n238 9.3005
R11935 gnd.n7117 gnd.n7116 9.3005
R11936 gnd.n7118 gnd.n237 9.3005
R11937 gnd.n7120 gnd.n7119 9.3005
R11938 gnd.n223 gnd.n222 9.3005
R11939 gnd.n7133 gnd.n7132 9.3005
R11940 gnd.n7134 gnd.n221 9.3005
R11941 gnd.n7136 gnd.n7135 9.3005
R11942 gnd.n209 gnd.n208 9.3005
R11943 gnd.n7149 gnd.n7148 9.3005
R11944 gnd.n7150 gnd.n207 9.3005
R11945 gnd.n7152 gnd.n7151 9.3005
R11946 gnd.n194 gnd.n193 9.3005
R11947 gnd.n7165 gnd.n7164 9.3005
R11948 gnd.n7166 gnd.n192 9.3005
R11949 gnd.n7170 gnd.n7167 9.3005
R11950 gnd.n7169 gnd.n7168 9.3005
R11951 gnd.n107 gnd.n106 9.3005
R11952 gnd.n7325 gnd.n7324 9.3005
R11953 gnd.n6971 gnd.n391 9.3005
R11954 gnd.n7068 gnd.n255 9.3005
R11955 gnd.n256 gnd.n255 9.3005
R11956 gnd.n4436 gnd.n4435 9.3005
R11957 gnd.n4437 gnd.n2328 9.3005
R11958 gnd.n4439 gnd.n4438 9.3005
R11959 gnd.n2326 gnd.n2325 9.3005
R11960 gnd.n4444 gnd.n4443 9.3005
R11961 gnd.n4445 gnd.n2324 9.3005
R11962 gnd.n4467 gnd.n4446 9.3005
R11963 gnd.n4466 gnd.n4447 9.3005
R11964 gnd.n4465 gnd.n4448 9.3005
R11965 gnd.n4451 gnd.n4449 9.3005
R11966 gnd.n4461 gnd.n4452 9.3005
R11967 gnd.n4460 gnd.n4453 9.3005
R11968 gnd.n4459 gnd.n4454 9.3005
R11969 gnd.n4457 gnd.n4456 9.3005
R11970 gnd.n4455 gnd.n2299 9.3005
R11971 gnd.n2297 gnd.n2296 9.3005
R11972 gnd.n4528 gnd.n4527 9.3005
R11973 gnd.n4529 gnd.n2295 9.3005
R11974 gnd.n4531 gnd.n4530 9.3005
R11975 gnd.n2293 gnd.n2292 9.3005
R11976 gnd.n4536 gnd.n4535 9.3005
R11977 gnd.n4537 gnd.n2291 9.3005
R11978 gnd.n4539 gnd.n4538 9.3005
R11979 gnd.n2289 gnd.n2288 9.3005
R11980 gnd.n4547 gnd.n4546 9.3005
R11981 gnd.n4548 gnd.n2287 9.3005
R11982 gnd.n4552 gnd.n4549 9.3005
R11983 gnd.n4551 gnd.n4550 9.3005
R11984 gnd.n2196 gnd.n2195 9.3005
R11985 gnd.n4620 gnd.n4619 9.3005
R11986 gnd.n4621 gnd.n2194 9.3005
R11987 gnd.n4623 gnd.n4622 9.3005
R11988 gnd.n2182 gnd.n2181 9.3005
R11989 gnd.n4639 gnd.n4638 9.3005
R11990 gnd.n4640 gnd.n2180 9.3005
R11991 gnd.n4642 gnd.n4641 9.3005
R11992 gnd.n2168 gnd.n2167 9.3005
R11993 gnd.n4659 gnd.n4658 9.3005
R11994 gnd.n4660 gnd.n2166 9.3005
R11995 gnd.n4668 gnd.n4661 9.3005
R11996 gnd.n4667 gnd.n4662 9.3005
R11997 gnd.n4666 gnd.n4663 9.3005
R11998 gnd.n1945 gnd.n1944 9.3005
R11999 gnd.n4711 gnd.n4710 9.3005
R12000 gnd.n4712 gnd.n1943 9.3005
R12001 gnd.n4719 gnd.n4713 9.3005
R12002 gnd.n4718 gnd.n4714 9.3005
R12003 gnd.n4717 gnd.n4715 9.3005
R12004 gnd.n1909 gnd.n1908 9.3005
R12005 gnd.n4794 gnd.n4793 9.3005
R12006 gnd.n4795 gnd.n1907 9.3005
R12007 gnd.n4797 gnd.n4796 9.3005
R12008 gnd.n1886 gnd.n1885 9.3005
R12009 gnd.n4821 gnd.n4820 9.3005
R12010 gnd.n4822 gnd.n1884 9.3005
R12011 gnd.n4826 gnd.n4823 9.3005
R12012 gnd.n4825 gnd.n4824 9.3005
R12013 gnd.n1856 gnd.n1855 9.3005
R12014 gnd.n4862 gnd.n4861 9.3005
R12015 gnd.n4863 gnd.n1854 9.3005
R12016 gnd.n4865 gnd.n4864 9.3005
R12017 gnd.n1832 gnd.n1831 9.3005
R12018 gnd.n4905 gnd.n4904 9.3005
R12019 gnd.n4906 gnd.n1830 9.3005
R12020 gnd.n4908 gnd.n4907 9.3005
R12021 gnd.n1816 gnd.n1815 9.3005
R12022 gnd.n5020 gnd.n5019 9.3005
R12023 gnd.n5021 gnd.n1814 9.3005
R12024 gnd.n5023 gnd.n5022 9.3005
R12025 gnd.n1793 gnd.n1792 9.3005
R12026 gnd.n5047 gnd.n5046 9.3005
R12027 gnd.n5048 gnd.n1791 9.3005
R12028 gnd.n5052 gnd.n5049 9.3005
R12029 gnd.n5051 gnd.n5050 9.3005
R12030 gnd.n1764 gnd.n1763 9.3005
R12031 gnd.n5083 gnd.n5082 9.3005
R12032 gnd.n5084 gnd.n1762 9.3005
R12033 gnd.n5086 gnd.n5085 9.3005
R12034 gnd.n1742 gnd.n1741 9.3005
R12035 gnd.n5113 gnd.n5112 9.3005
R12036 gnd.n5114 gnd.n1740 9.3005
R12037 gnd.n5116 gnd.n5115 9.3005
R12038 gnd.n1720 gnd.n1719 9.3005
R12039 gnd.n5143 gnd.n5142 9.3005
R12040 gnd.n5144 gnd.n1718 9.3005
R12041 gnd.n5146 gnd.n5145 9.3005
R12042 gnd.n1698 gnd.n1697 9.3005
R12043 gnd.n5170 gnd.n5169 9.3005
R12044 gnd.n5171 gnd.n1696 9.3005
R12045 gnd.n5175 gnd.n5172 9.3005
R12046 gnd.n5174 gnd.n5173 9.3005
R12047 gnd.n1671 gnd.n1670 9.3005
R12048 gnd.n5207 gnd.n5206 9.3005
R12049 gnd.n5208 gnd.n1669 9.3005
R12050 gnd.n5221 gnd.n5209 9.3005
R12051 gnd.n5220 gnd.n5210 9.3005
R12052 gnd.n5219 gnd.n5211 9.3005
R12053 gnd.n5213 gnd.n5212 9.3005
R12054 gnd.n5215 gnd.n5214 9.3005
R12055 gnd.n1599 gnd.n1598 9.3005
R12056 gnd.n5408 gnd.n5407 9.3005
R12057 gnd.n5409 gnd.n1597 9.3005
R12058 gnd.n5411 gnd.n5410 9.3005
R12059 gnd.n1585 gnd.n1584 9.3005
R12060 gnd.n5427 gnd.n5426 9.3005
R12061 gnd.n5428 gnd.n1583 9.3005
R12062 gnd.n5433 gnd.n5429 9.3005
R12063 gnd.n5432 gnd.n5431 9.3005
R12064 gnd.n5430 gnd.n1572 9.3005
R12065 gnd.n1570 gnd.n1569 9.3005
R12066 gnd.n5451 gnd.n5450 9.3005
R12067 gnd.n5452 gnd.n1568 9.3005
R12068 gnd.n5627 gnd.n5453 9.3005
R12069 gnd.n5626 gnd.n5454 9.3005
R12070 gnd.n5625 gnd.n5455 9.3005
R12071 gnd.n5458 gnd.n5456 9.3005
R12072 gnd.n5621 gnd.n5459 9.3005
R12073 gnd.n5620 gnd.n5460 9.3005
R12074 gnd.n5619 gnd.n5461 9.3005
R12075 gnd.n5483 gnd.n5462 9.3005
R12076 gnd.n5486 gnd.n5485 9.3005
R12077 gnd.n5487 gnd.n5482 9.3005
R12078 gnd.n5489 gnd.n5488 9.3005
R12079 gnd.n5480 gnd.n5479 9.3005
R12080 gnd.n5494 gnd.n5493 9.3005
R12081 gnd.n5495 gnd.n5478 9.3005
R12082 gnd.n5595 gnd.n5496 9.3005
R12083 gnd.n5594 gnd.n5497 9.3005
R12084 gnd.n5593 gnd.n5498 9.3005
R12085 gnd.n5501 gnd.n5499 9.3005
R12086 gnd.n5589 gnd.n5502 9.3005
R12087 gnd.n5588 gnd.n5503 9.3005
R12088 gnd.n5587 gnd.n5504 9.3005
R12089 gnd.n5537 gnd.n5505 9.3005
R12090 gnd.n5538 gnd.n5507 9.3005
R12091 gnd.n5540 gnd.n5539 9.3005
R12092 gnd.n5541 gnd.n5536 9.3005
R12093 gnd.n5573 gnd.n5542 9.3005
R12094 gnd.n6833 gnd.n556 9.3005
R12095 gnd.n6832 gnd.n557 9.3005
R12096 gnd.n560 gnd.n558 9.3005
R12097 gnd.n6828 gnd.n561 9.3005
R12098 gnd.n6827 gnd.n6826 9.3005
R12099 gnd.n1304 gnd.n1298 9.3005
R12100 gnd.n5904 gnd.n1297 9.3005
R12101 gnd.n5905 gnd.n1296 9.3005
R12102 gnd.n5906 gnd.n1295 9.3005
R12103 gnd.n1294 gnd.n1291 9.3005
R12104 gnd.n5911 gnd.n1290 9.3005
R12105 gnd.n5912 gnd.n1289 9.3005
R12106 gnd.n5913 gnd.n1288 9.3005
R12107 gnd.n1287 gnd.n1284 9.3005
R12108 gnd.n5918 gnd.n1283 9.3005
R12109 gnd.n5919 gnd.n1282 9.3005
R12110 gnd.n5920 gnd.n1281 9.3005
R12111 gnd.n1280 gnd.n1277 9.3005
R12112 gnd.n1279 gnd.n1275 9.3005
R12113 gnd.n5927 gnd.n1274 9.3005
R12114 gnd.n5929 gnd.n5928 9.3005
R12115 gnd.n5896 gnd.n1307 9.3005
R12116 gnd.n5895 gnd.n1308 9.3005
R12117 gnd.n1312 gnd.n1309 9.3005
R12118 gnd.n5890 gnd.n1313 9.3005
R12119 gnd.n5889 gnd.n1314 9.3005
R12120 gnd.n5888 gnd.n1315 9.3005
R12121 gnd.n1319 gnd.n1316 9.3005
R12122 gnd.n5883 gnd.n1320 9.3005
R12123 gnd.n5882 gnd.n1321 9.3005
R12124 gnd.n5881 gnd.n1322 9.3005
R12125 gnd.n1326 gnd.n1323 9.3005
R12126 gnd.n5876 gnd.n1327 9.3005
R12127 gnd.n5875 gnd.n1328 9.3005
R12128 gnd.n5874 gnd.n1329 9.3005
R12129 gnd.n1333 gnd.n1330 9.3005
R12130 gnd.n5869 gnd.n1334 9.3005
R12131 gnd.n5868 gnd.n1335 9.3005
R12132 gnd.n5867 gnd.n1336 9.3005
R12133 gnd.n1341 gnd.n1339 9.3005
R12134 gnd.n5862 gnd.n5861 9.3005
R12135 gnd.n5897 gnd.n1306 9.3005
R12136 gnd.n4167 gnd.n4124 9.3005
R12137 gnd.n4166 gnd.n4126 9.3005
R12138 gnd.n4165 gnd.n4127 9.3005
R12139 gnd.n4163 gnd.n4128 9.3005
R12140 gnd.n4162 gnd.n4129 9.3005
R12141 gnd.n4160 gnd.n4130 9.3005
R12142 gnd.n4159 gnd.n4131 9.3005
R12143 gnd.n4157 gnd.n4132 9.3005
R12144 gnd.n4156 gnd.n4133 9.3005
R12145 gnd.n4154 gnd.n4134 9.3005
R12146 gnd.n4153 gnd.n4135 9.3005
R12147 gnd.n4151 gnd.n4136 9.3005
R12148 gnd.n4150 gnd.n4137 9.3005
R12149 gnd.n4148 gnd.n4138 9.3005
R12150 gnd.n4147 gnd.n4139 9.3005
R12151 gnd.n4145 gnd.n4140 9.3005
R12152 gnd.n4144 gnd.n4142 9.3005
R12153 gnd.n4141 gnd.n2391 9.3005
R12154 gnd.n4328 gnd.n2392 9.3005
R12155 gnd.n4327 gnd.n2393 9.3005
R12156 gnd.n4326 gnd.n2394 9.3005
R12157 gnd.n4302 gnd.n2395 9.3005
R12158 gnd.n4316 gnd.n4303 9.3005
R12159 gnd.n4315 gnd.n4304 9.3005
R12160 gnd.n4314 gnd.n4305 9.3005
R12161 gnd.n4312 gnd.n4306 9.3005
R12162 gnd.n4169 gnd.n4168 9.3005
R12163 gnd.n4177 gnd.n4176 9.3005
R12164 gnd.n4178 gnd.n4120 9.3005
R12165 gnd.n4119 gnd.n4117 9.3005
R12166 gnd.n4184 gnd.n4116 9.3005
R12167 gnd.n4185 gnd.n4115 9.3005
R12168 gnd.n4186 gnd.n4114 9.3005
R12169 gnd.n4113 gnd.n4111 9.3005
R12170 gnd.n4192 gnd.n4110 9.3005
R12171 gnd.n4193 gnd.n4109 9.3005
R12172 gnd.n4194 gnd.n4108 9.3005
R12173 gnd.n4107 gnd.n4105 9.3005
R12174 gnd.n4200 gnd.n4104 9.3005
R12175 gnd.n4201 gnd.n4103 9.3005
R12176 gnd.n4202 gnd.n4102 9.3005
R12177 gnd.n4101 gnd.n4099 9.3005
R12178 gnd.n4208 gnd.n4098 9.3005
R12179 gnd.n4210 gnd.n4209 9.3005
R12180 gnd.n4175 gnd.n4123 9.3005
R12181 gnd.n4174 gnd.n4173 9.3005
R12182 gnd.n2449 gnd.n2448 9.3005
R12183 gnd.n4225 gnd.n4224 9.3005
R12184 gnd.n4226 gnd.n2447 9.3005
R12185 gnd.n4228 gnd.n4227 9.3005
R12186 gnd.n2433 gnd.n2432 9.3005
R12187 gnd.n4241 gnd.n4240 9.3005
R12188 gnd.n4242 gnd.n2431 9.3005
R12189 gnd.n4244 gnd.n4243 9.3005
R12190 gnd.n2416 gnd.n2415 9.3005
R12191 gnd.n4257 gnd.n4256 9.3005
R12192 gnd.n4258 gnd.n2414 9.3005
R12193 gnd.n4270 gnd.n4259 9.3005
R12194 gnd.n4269 gnd.n4260 9.3005
R12195 gnd.n4268 gnd.n4261 9.3005
R12196 gnd.n4267 gnd.n4262 9.3005
R12197 gnd.n4265 gnd.n4264 9.3005
R12198 gnd.n4263 gnd.n1128 9.3005
R12199 gnd.n6012 gnd.n1129 9.3005
R12200 gnd.n6011 gnd.n1130 9.3005
R12201 gnd.n6010 gnd.n1131 9.3005
R12202 gnd.n2377 gnd.n1132 9.3005
R12203 gnd.n4347 gnd.n4346 9.3005
R12204 gnd.n4348 gnd.n2376 9.3005
R12205 gnd.n4353 gnd.n4349 9.3005
R12206 gnd.n4352 gnd.n4350 9.3005
R12207 gnd.n4351 gnd.n2355 9.3005
R12208 gnd.n4380 gnd.n2354 9.3005
R12209 gnd.n4385 gnd.n4381 9.3005
R12210 gnd.n4384 gnd.n4383 9.3005
R12211 gnd.n4382 gnd.n1158 9.3005
R12212 gnd.n5997 gnd.n1159 9.3005
R12213 gnd.n5996 gnd.n1160 9.3005
R12214 gnd.n5995 gnd.n1161 9.3005
R12215 gnd.n1178 gnd.n1162 9.3005
R12216 gnd.n5985 gnd.n1179 9.3005
R12217 gnd.n5984 gnd.n1180 9.3005
R12218 gnd.n5983 gnd.n1181 9.3005
R12219 gnd.n1199 gnd.n1182 9.3005
R12220 gnd.n5973 gnd.n1200 9.3005
R12221 gnd.n5972 gnd.n1201 9.3005
R12222 gnd.n5971 gnd.n1202 9.3005
R12223 gnd.n1220 gnd.n1203 9.3005
R12224 gnd.n5961 gnd.n1221 9.3005
R12225 gnd.n5960 gnd.n1222 9.3005
R12226 gnd.n5959 gnd.n1223 9.3005
R12227 gnd.n1241 gnd.n1224 9.3005
R12228 gnd.n5949 gnd.n1242 9.3005
R12229 gnd.n5948 gnd.n1243 9.3005
R12230 gnd.n5947 gnd.n1244 9.3005
R12231 gnd.n1263 gnd.n1245 9.3005
R12232 gnd.n5937 gnd.n1264 9.3005
R12233 gnd.n5936 gnd.n1265 9.3005
R12234 gnd.n5935 gnd.n1266 9.3005
R12235 gnd.n4212 gnd.n4211 9.3005
R12236 gnd.n4094 gnd.n4093 9.3005
R12237 gnd.n4092 gnd.n3924 9.3005
R12238 gnd.n4091 gnd.n4090 9.3005
R12239 gnd.n4088 gnd.n4065 9.3005
R12240 gnd.n4087 gnd.n4066 9.3005
R12241 gnd.n4085 gnd.n4067 9.3005
R12242 gnd.n4084 gnd.n4068 9.3005
R12243 gnd.n4082 gnd.n4069 9.3005
R12244 gnd.n4081 gnd.n4070 9.3005
R12245 gnd.n4079 gnd.n4071 9.3005
R12246 gnd.n4078 gnd.n4072 9.3005
R12247 gnd.n4076 gnd.n4073 9.3005
R12248 gnd.n4075 gnd.n4074 9.3005
R12249 gnd.n2400 gnd.n2399 9.3005
R12250 gnd.n4285 gnd.n4284 9.3005
R12251 gnd.n4286 gnd.n2398 9.3005
R12252 gnd.n4289 gnd.n4287 9.3005
R12253 gnd.n4290 gnd.n2397 9.3005
R12254 gnd.n4292 gnd.n4291 9.3005
R12255 gnd.n4293 gnd.n2396 9.3005
R12256 gnd.n4322 gnd.n4294 9.3005
R12257 gnd.n4321 gnd.n4295 9.3005
R12258 gnd.n4320 gnd.n4296 9.3005
R12259 gnd.n4301 gnd.n4297 9.3005
R12260 gnd.n4300 gnd.n4298 9.3005
R12261 gnd.n2358 gnd.n2356 9.3005
R12262 gnd.n4377 gnd.n4376 9.3005
R12263 gnd.n2357 gnd.n2347 9.3005
R12264 gnd.n4394 gnd.n2346 9.3005
R12265 gnd.n4396 gnd.n4395 9.3005
R12266 gnd.n4397 gnd.n2345 9.3005
R12267 gnd.n4401 gnd.n4398 9.3005
R12268 gnd.n4402 gnd.n2344 9.3005
R12269 gnd.n4407 gnd.n4406 9.3005
R12270 gnd.n4408 gnd.n2343 9.3005
R12271 gnd.n4414 gnd.n4409 9.3005
R12272 gnd.n4413 gnd.n4410 9.3005
R12273 gnd.n4412 gnd.n4411 9.3005
R12274 gnd.n2317 gnd.n2316 9.3005
R12275 gnd.n4481 gnd.n4480 9.3005
R12276 gnd.n4482 gnd.n2315 9.3005
R12277 gnd.n4484 gnd.n4483 9.3005
R12278 gnd.n2310 gnd.n2309 9.3005
R12279 gnd.n4497 gnd.n4496 9.3005
R12280 gnd.n4498 gnd.n2308 9.3005
R12281 gnd.n4500 gnd.n4499 9.3005
R12282 gnd.n4501 gnd.n2307 9.3005
R12283 gnd.n4505 gnd.n4504 9.3005
R12284 gnd.n4506 gnd.n2306 9.3005
R12285 gnd.n4509 gnd.n4508 9.3005
R12286 gnd.n4507 gnd.n1343 9.3005
R12287 gnd.n5858 gnd.n1342 9.3005
R12288 gnd.n5860 gnd.n5859 9.3005
R12289 gnd.n4064 gnd.n3923 9.3005
R12290 gnd.n4053 gnd.n3929 9.3005
R12291 gnd.n4055 gnd.n4054 9.3005
R12292 gnd.n4052 gnd.n3931 9.3005
R12293 gnd.n4051 gnd.n4050 9.3005
R12294 gnd.n3933 gnd.n3932 9.3005
R12295 gnd.n4044 gnd.n4043 9.3005
R12296 gnd.n4042 gnd.n3935 9.3005
R12297 gnd.n4041 gnd.n4040 9.3005
R12298 gnd.n3937 gnd.n3936 9.3005
R12299 gnd.n4034 gnd.n4033 9.3005
R12300 gnd.n4032 gnd.n3939 9.3005
R12301 gnd.n4031 gnd.n4030 9.3005
R12302 gnd.n3941 gnd.n3940 9.3005
R12303 gnd.n4024 gnd.n4023 9.3005
R12304 gnd.n4022 gnd.n3943 9.3005
R12305 gnd.n4021 gnd.n4020 9.3005
R12306 gnd.n3945 gnd.n3944 9.3005
R12307 gnd.n4014 gnd.n4013 9.3005
R12308 gnd.n4012 gnd.n3947 9.3005
R12309 gnd.n4011 gnd.n4010 9.3005
R12310 gnd.n3949 gnd.n3948 9.3005
R12311 gnd.n4004 gnd.n4003 9.3005
R12312 gnd.n4002 gnd.n3954 9.3005
R12313 gnd.n4001 gnd.n4000 9.3005
R12314 gnd.n3956 gnd.n3955 9.3005
R12315 gnd.n3994 gnd.n3993 9.3005
R12316 gnd.n3992 gnd.n3958 9.3005
R12317 gnd.n3991 gnd.n3990 9.3005
R12318 gnd.n3960 gnd.n3959 9.3005
R12319 gnd.n3984 gnd.n3983 9.3005
R12320 gnd.n3982 gnd.n3962 9.3005
R12321 gnd.n3981 gnd.n3980 9.3005
R12322 gnd.n3964 gnd.n3963 9.3005
R12323 gnd.n3974 gnd.n3973 9.3005
R12324 gnd.n3972 gnd.n3966 9.3005
R12325 gnd.n3971 gnd.n3970 9.3005
R12326 gnd.n3967 gnd.n2455 9.3005
R12327 gnd.n3928 gnd.n3925 9.3005
R12328 gnd.n4063 gnd.n4062 9.3005
R12329 gnd.n4218 gnd.n2454 9.3005
R12330 gnd.n4220 gnd.n4219 9.3005
R12331 gnd.n2441 gnd.n2440 9.3005
R12332 gnd.n4233 gnd.n4232 9.3005
R12333 gnd.n4234 gnd.n2439 9.3005
R12334 gnd.n4236 gnd.n4235 9.3005
R12335 gnd.n2424 gnd.n2423 9.3005
R12336 gnd.n4249 gnd.n4248 9.3005
R12337 gnd.n4250 gnd.n2422 9.3005
R12338 gnd.n4252 gnd.n4251 9.3005
R12339 gnd.n2408 gnd.n2407 9.3005
R12340 gnd.n4275 gnd.n4274 9.3005
R12341 gnd.n4276 gnd.n2406 9.3005
R12342 gnd.n4279 gnd.n4278 9.3005
R12343 gnd.n4277 gnd.n1116 9.3005
R12344 gnd.n6018 gnd.n1117 9.3005
R12345 gnd.n6017 gnd.n1118 9.3005
R12346 gnd.n6016 gnd.n1119 9.3005
R12347 gnd.n1138 gnd.n1120 9.3005
R12348 gnd.n6006 gnd.n1139 9.3005
R12349 gnd.n6005 gnd.n1140 9.3005
R12350 gnd.n1150 gnd.n1143 9.3005
R12351 gnd.n5991 gnd.n1168 9.3005
R12352 gnd.n5990 gnd.n1169 9.3005
R12353 gnd.n5989 gnd.n1170 9.3005
R12354 gnd.n1189 gnd.n1171 9.3005
R12355 gnd.n5979 gnd.n1190 9.3005
R12356 gnd.n5978 gnd.n1191 9.3005
R12357 gnd.n5977 gnd.n1192 9.3005
R12358 gnd.n1209 gnd.n1193 9.3005
R12359 gnd.n5967 gnd.n1210 9.3005
R12360 gnd.n5966 gnd.n1211 9.3005
R12361 gnd.n5965 gnd.n1212 9.3005
R12362 gnd.n1231 gnd.n1213 9.3005
R12363 gnd.n5955 gnd.n1232 9.3005
R12364 gnd.n5954 gnd.n1233 9.3005
R12365 gnd.n5953 gnd.n1234 9.3005
R12366 gnd.n1252 gnd.n1235 9.3005
R12367 gnd.n5943 gnd.n1253 9.3005
R12368 gnd.n5942 gnd.n1254 9.3005
R12369 gnd.n5941 gnd.n1255 9.3005
R12370 gnd.n1273 gnd.n1256 9.3005
R12371 gnd.n5931 gnd.n5930 9.3005
R12372 gnd.n4217 gnd.n4216 9.3005
R12373 gnd.n6002 gnd.n1148 9.3005
R12374 gnd.n6002 gnd.n6001 9.3005
R12375 gnd.n2387 gnd.n2384 9.3005
R12376 gnd.n4334 gnd.n4333 9.3005
R12377 gnd.n4335 gnd.n2383 9.3005
R12378 gnd.n4337 gnd.n4336 9.3005
R12379 gnd.n2386 gnd.n2385 9.3005
R12380 gnd.n6024 gnd.n1106 9.3005
R12381 gnd.n6025 gnd.n1105 9.3005
R12382 gnd.n1104 gnd.n1100 9.3005
R12383 gnd.n6031 gnd.n1099 9.3005
R12384 gnd.n6032 gnd.n1098 9.3005
R12385 gnd.n6033 gnd.n1097 9.3005
R12386 gnd.n1096 gnd.n1092 9.3005
R12387 gnd.n6039 gnd.n1091 9.3005
R12388 gnd.n6040 gnd.n1090 9.3005
R12389 gnd.n6041 gnd.n1089 9.3005
R12390 gnd.n1088 gnd.n1084 9.3005
R12391 gnd.n6047 gnd.n1083 9.3005
R12392 gnd.n6048 gnd.n1082 9.3005
R12393 gnd.n6049 gnd.n1081 9.3005
R12394 gnd.n1080 gnd.n1076 9.3005
R12395 gnd.n6055 gnd.n1075 9.3005
R12396 gnd.n6056 gnd.n1074 9.3005
R12397 gnd.n6057 gnd.n1073 9.3005
R12398 gnd.n1072 gnd.n1068 9.3005
R12399 gnd.n6063 gnd.n1067 9.3005
R12400 gnd.n6064 gnd.n1066 9.3005
R12401 gnd.n6065 gnd.n1065 9.3005
R12402 gnd.n1064 gnd.n1060 9.3005
R12403 gnd.n6071 gnd.n1059 9.3005
R12404 gnd.n6072 gnd.n1058 9.3005
R12405 gnd.n6073 gnd.n1057 9.3005
R12406 gnd.n1056 gnd.n1052 9.3005
R12407 gnd.n6079 gnd.n1051 9.3005
R12408 gnd.n6080 gnd.n1050 9.3005
R12409 gnd.n6081 gnd.n1049 9.3005
R12410 gnd.n1048 gnd.n1044 9.3005
R12411 gnd.n6087 gnd.n1043 9.3005
R12412 gnd.n6088 gnd.n1042 9.3005
R12413 gnd.n6089 gnd.n1041 9.3005
R12414 gnd.n1040 gnd.n1036 9.3005
R12415 gnd.n6095 gnd.n1035 9.3005
R12416 gnd.n6096 gnd.n1034 9.3005
R12417 gnd.n6097 gnd.n1033 9.3005
R12418 gnd.n1032 gnd.n1028 9.3005
R12419 gnd.n6103 gnd.n1027 9.3005
R12420 gnd.n6104 gnd.n1026 9.3005
R12421 gnd.n6105 gnd.n1025 9.3005
R12422 gnd.n1024 gnd.n1020 9.3005
R12423 gnd.n6111 gnd.n1019 9.3005
R12424 gnd.n6112 gnd.n1018 9.3005
R12425 gnd.n6113 gnd.n1017 9.3005
R12426 gnd.n1016 gnd.n1012 9.3005
R12427 gnd.n6119 gnd.n1011 9.3005
R12428 gnd.n6120 gnd.n1010 9.3005
R12429 gnd.n6121 gnd.n1009 9.3005
R12430 gnd.n1008 gnd.n1004 9.3005
R12431 gnd.n6127 gnd.n1003 9.3005
R12432 gnd.n6128 gnd.n1002 9.3005
R12433 gnd.n6129 gnd.n1001 9.3005
R12434 gnd.n1000 gnd.n996 9.3005
R12435 gnd.n6135 gnd.n995 9.3005
R12436 gnd.n6136 gnd.n994 9.3005
R12437 gnd.n6137 gnd.n993 9.3005
R12438 gnd.n992 gnd.n988 9.3005
R12439 gnd.n6143 gnd.n987 9.3005
R12440 gnd.n6144 gnd.n986 9.3005
R12441 gnd.n6145 gnd.n985 9.3005
R12442 gnd.n984 gnd.n980 9.3005
R12443 gnd.n6151 gnd.n979 9.3005
R12444 gnd.n6152 gnd.n978 9.3005
R12445 gnd.n6153 gnd.n977 9.3005
R12446 gnd.n976 gnd.n972 9.3005
R12447 gnd.n6159 gnd.n971 9.3005
R12448 gnd.n6160 gnd.n970 9.3005
R12449 gnd.n6161 gnd.n969 9.3005
R12450 gnd.n968 gnd.n964 9.3005
R12451 gnd.n6167 gnd.n963 9.3005
R12452 gnd.n6168 gnd.n962 9.3005
R12453 gnd.n6169 gnd.n961 9.3005
R12454 gnd.n960 gnd.n956 9.3005
R12455 gnd.n6175 gnd.n955 9.3005
R12456 gnd.n6176 gnd.n954 9.3005
R12457 gnd.n6177 gnd.n953 9.3005
R12458 gnd.n952 gnd.n948 9.3005
R12459 gnd.n6183 gnd.n947 9.3005
R12460 gnd.n6184 gnd.n946 9.3005
R12461 gnd.n6185 gnd.n945 9.3005
R12462 gnd.n941 gnd.n940 9.3005
R12463 gnd.n6192 gnd.n6191 9.3005
R12464 gnd.n6023 gnd.n1107 9.3005
R12465 gnd.n5697 gnd.n5696 9.3005
R12466 gnd.n5695 gnd.n5694 9.3005
R12467 gnd.n1487 gnd.n1486 9.3005
R12468 gnd.n5689 gnd.n5688 9.3005
R12469 gnd.n5687 gnd.n5686 9.3005
R12470 gnd.n1497 gnd.n1496 9.3005
R12471 gnd.n5681 gnd.n5680 9.3005
R12472 gnd.n5679 gnd.n5678 9.3005
R12473 gnd.n1505 gnd.n1504 9.3005
R12474 gnd.n5673 gnd.n5672 9.3005
R12475 gnd.n5671 gnd.n5670 9.3005
R12476 gnd.n1515 gnd.n1514 9.3005
R12477 gnd.n5665 gnd.n5664 9.3005
R12478 gnd.n5663 gnd.n5662 9.3005
R12479 gnd.n1523 gnd.n1522 9.3005
R12480 gnd.n5654 gnd.n5653 9.3005
R12481 gnd.n5652 gnd.n5651 9.3005
R12482 gnd.n5650 gnd.n5649 9.3005
R12483 gnd.n1483 gnd.n1481 9.3005
R12484 gnd.n5661 gnd.n5660 9.3005
R12485 gnd.n1519 gnd.n1518 9.3005
R12486 gnd.n5667 gnd.n5666 9.3005
R12487 gnd.n5669 gnd.n5668 9.3005
R12488 gnd.n1511 gnd.n1510 9.3005
R12489 gnd.n5675 gnd.n5674 9.3005
R12490 gnd.n5677 gnd.n5676 9.3005
R12491 gnd.n1501 gnd.n1500 9.3005
R12492 gnd.n5683 gnd.n5682 9.3005
R12493 gnd.n5685 gnd.n5684 9.3005
R12494 gnd.n1493 gnd.n1492 9.3005
R12495 gnd.n5691 gnd.n5690 9.3005
R12496 gnd.n5693 gnd.n5692 9.3005
R12497 gnd.n1482 gnd.n1480 9.3005
R12498 gnd.n5699 gnd.n5698 9.3005
R12499 gnd.n5700 gnd.n1477 9.3005
R12500 gnd.n5659 gnd.n5655 9.3005
R12501 gnd.n1527 gnd.n1526 9.3005
R12502 gnd.n5648 gnd.n5647 9.3005
R12503 gnd.n5646 gnd.n1532 9.3005
R12504 gnd.n5645 gnd.n5644 9.3005
R12505 gnd.n5643 gnd.n1533 9.3005
R12506 gnd.n5642 gnd.n5641 9.3005
R12507 gnd.n5640 gnd.n1537 9.3005
R12508 gnd.n5639 gnd.n5638 9.3005
R12509 gnd.n5637 gnd.n1538 9.3005
R12510 gnd.n5636 gnd.n5635 9.3005
R12511 gnd.n5634 gnd.n5633 9.3005
R12512 gnd.n5831 gnd.n1366 9.3005
R12513 gnd.n5830 gnd.n5829 9.3005
R12514 gnd.n5828 gnd.n1370 9.3005
R12515 gnd.n5827 gnd.n5826 9.3005
R12516 gnd.n5825 gnd.n1371 9.3005
R12517 gnd.n5824 gnd.n5823 9.3005
R12518 gnd.n5822 gnd.n1375 9.3005
R12519 gnd.n5821 gnd.n5820 9.3005
R12520 gnd.n5819 gnd.n1376 9.3005
R12521 gnd.n5818 gnd.n5817 9.3005
R12522 gnd.n5816 gnd.n1380 9.3005
R12523 gnd.n5815 gnd.n5814 9.3005
R12524 gnd.n5813 gnd.n1381 9.3005
R12525 gnd.n5812 gnd.n5811 9.3005
R12526 gnd.n5810 gnd.n1385 9.3005
R12527 gnd.n5809 gnd.n5808 9.3005
R12528 gnd.n5807 gnd.n1386 9.3005
R12529 gnd.n5806 gnd.n5805 9.3005
R12530 gnd.n5804 gnd.n1390 9.3005
R12531 gnd.n5803 gnd.n5802 9.3005
R12532 gnd.n5801 gnd.n1391 9.3005
R12533 gnd.n5800 gnd.n5799 9.3005
R12534 gnd.n5798 gnd.n1395 9.3005
R12535 gnd.n5797 gnd.n5796 9.3005
R12536 gnd.n5795 gnd.n1396 9.3005
R12537 gnd.n5794 gnd.n5793 9.3005
R12538 gnd.n5792 gnd.n1400 9.3005
R12539 gnd.n5791 gnd.n5790 9.3005
R12540 gnd.n5789 gnd.n1401 9.3005
R12541 gnd.n5788 gnd.n5787 9.3005
R12542 gnd.n5786 gnd.n1405 9.3005
R12543 gnd.n5785 gnd.n5784 9.3005
R12544 gnd.n5783 gnd.n1406 9.3005
R12545 gnd.n5782 gnd.n5781 9.3005
R12546 gnd.n5780 gnd.n1410 9.3005
R12547 gnd.n5779 gnd.n5778 9.3005
R12548 gnd.n5777 gnd.n1411 9.3005
R12549 gnd.n5776 gnd.n5775 9.3005
R12550 gnd.n5774 gnd.n1415 9.3005
R12551 gnd.n5773 gnd.n5772 9.3005
R12552 gnd.n5771 gnd.n1416 9.3005
R12553 gnd.n5770 gnd.n5769 9.3005
R12554 gnd.n5768 gnd.n1420 9.3005
R12555 gnd.n5767 gnd.n5766 9.3005
R12556 gnd.n5765 gnd.n1421 9.3005
R12557 gnd.n5764 gnd.n5763 9.3005
R12558 gnd.n5762 gnd.n1425 9.3005
R12559 gnd.n5761 gnd.n5760 9.3005
R12560 gnd.n5759 gnd.n1426 9.3005
R12561 gnd.n5758 gnd.n5757 9.3005
R12562 gnd.n5756 gnd.n1430 9.3005
R12563 gnd.n5755 gnd.n5754 9.3005
R12564 gnd.n5753 gnd.n1431 9.3005
R12565 gnd.n5752 gnd.n5751 9.3005
R12566 gnd.n5750 gnd.n1435 9.3005
R12567 gnd.n5749 gnd.n5748 9.3005
R12568 gnd.n5747 gnd.n1436 9.3005
R12569 gnd.n5746 gnd.n5745 9.3005
R12570 gnd.n5744 gnd.n1440 9.3005
R12571 gnd.n5743 gnd.n5742 9.3005
R12572 gnd.n5741 gnd.n1441 9.3005
R12573 gnd.n5740 gnd.n5739 9.3005
R12574 gnd.n5738 gnd.n1445 9.3005
R12575 gnd.n5737 gnd.n5736 9.3005
R12576 gnd.n5735 gnd.n1446 9.3005
R12577 gnd.n5734 gnd.n5733 9.3005
R12578 gnd.n5732 gnd.n1450 9.3005
R12579 gnd.n5731 gnd.n5730 9.3005
R12580 gnd.n5729 gnd.n1451 9.3005
R12581 gnd.n5728 gnd.n5727 9.3005
R12582 gnd.n5726 gnd.n1455 9.3005
R12583 gnd.n5725 gnd.n5724 9.3005
R12584 gnd.n5723 gnd.n1456 9.3005
R12585 gnd.n5722 gnd.n5721 9.3005
R12586 gnd.n5720 gnd.n1460 9.3005
R12587 gnd.n5719 gnd.n5718 9.3005
R12588 gnd.n5717 gnd.n1461 9.3005
R12589 gnd.n5716 gnd.n5715 9.3005
R12590 gnd.n5714 gnd.n1465 9.3005
R12591 gnd.n5713 gnd.n5712 9.3005
R12592 gnd.n5711 gnd.n1466 9.3005
R12593 gnd.n5710 gnd.n1469 9.3005
R12594 gnd.n5833 gnd.n5832 9.3005
R12595 gnd.n5836 gnd.n5835 9.3005
R12596 gnd.n5837 gnd.n1361 9.3005
R12597 gnd.n5839 gnd.n5838 9.3005
R12598 gnd.n5841 gnd.n5840 9.3005
R12599 gnd.n5842 gnd.n1354 9.3005
R12600 gnd.n5844 gnd.n5843 9.3005
R12601 gnd.n5845 gnd.n1353 9.3005
R12602 gnd.n5847 gnd.n5846 9.3005
R12603 gnd.n5848 gnd.n1347 9.3005
R12604 gnd.n5834 gnd.n1365 9.3005
R12605 gnd.n4311 gnd.n4310 9.3005
R12606 gnd.n4309 gnd.n4307 9.3005
R12607 gnd.n2338 gnd.n2336 9.3005
R12608 gnd.n4428 gnd.n4427 9.3005
R12609 gnd.n4426 gnd.n2337 9.3005
R12610 gnd.n4425 gnd.n4424 9.3005
R12611 gnd.n4423 gnd.n2339 9.3005
R12612 gnd.n4422 gnd.n4421 9.3005
R12613 gnd.n4420 gnd.n2342 9.3005
R12614 gnd.n4419 gnd.n4418 9.3005
R12615 gnd.n2320 gnd.n2319 9.3005
R12616 gnd.n4473 gnd.n4472 9.3005
R12617 gnd.n4474 gnd.n2318 9.3005
R12618 gnd.n4476 gnd.n4475 9.3005
R12619 gnd.n2313 gnd.n2312 9.3005
R12620 gnd.n4489 gnd.n4488 9.3005
R12621 gnd.n4490 gnd.n2311 9.3005
R12622 gnd.n4492 gnd.n4491 9.3005
R12623 gnd.n2303 gnd.n2301 9.3005
R12624 gnd.n4520 gnd.n4519 9.3005
R12625 gnd.n4518 gnd.n2302 9.3005
R12626 gnd.n4517 gnd.n4516 9.3005
R12627 gnd.n4515 gnd.n2304 9.3005
R12628 gnd.n4514 gnd.n4513 9.3005
R12629 gnd.n1346 gnd.n1344 9.3005
R12630 gnd.n5854 gnd.n5853 9.3005
R12631 gnd.n5852 gnd.n1345 9.3005
R12632 gnd.n5850 gnd.n5849 9.3005
R12633 gnd.n1349 gnd.n1348 9.3005
R12634 gnd.n4561 gnd.n4560 9.3005
R12635 gnd.n2254 gnd.n2253 9.3005
R12636 gnd.n4570 gnd.n4569 9.3005
R12637 gnd.n4572 gnd.n4571 9.3005
R12638 gnd.n2243 gnd.n2242 9.3005
R12639 gnd.n4578 gnd.n4577 9.3005
R12640 gnd.n4580 gnd.n4579 9.3005
R12641 gnd.n2233 gnd.n2232 9.3005
R12642 gnd.n4586 gnd.n4585 9.3005
R12643 gnd.n4588 gnd.n4587 9.3005
R12644 gnd.n2222 gnd.n2221 9.3005
R12645 gnd.n4594 gnd.n4593 9.3005
R12646 gnd.n4596 gnd.n4595 9.3005
R12647 gnd.n2212 gnd.n2211 9.3005
R12648 gnd.n4602 gnd.n4601 9.3005
R12649 gnd.n4604 gnd.n4603 9.3005
R12650 gnd.n2208 gnd.n2206 9.3005
R12651 gnd.n4607 gnd.n2201 9.3005
R12652 gnd.n4606 gnd.n4605 9.3005
R12653 gnd.n2207 gnd.n2205 9.3005
R12654 gnd.n4600 gnd.n4599 9.3005
R12655 gnd.n4598 gnd.n4597 9.3005
R12656 gnd.n2218 gnd.n2217 9.3005
R12657 gnd.n4592 gnd.n4591 9.3005
R12658 gnd.n4590 gnd.n4589 9.3005
R12659 gnd.n2229 gnd.n2228 9.3005
R12660 gnd.n4584 gnd.n4583 9.3005
R12661 gnd.n4582 gnd.n4581 9.3005
R12662 gnd.n2239 gnd.n2238 9.3005
R12663 gnd.n4576 gnd.n4575 9.3005
R12664 gnd.n4574 gnd.n4573 9.3005
R12665 gnd.n2250 gnd.n2249 9.3005
R12666 gnd.n4568 gnd.n4567 9.3005
R12667 gnd.n4566 gnd.n2260 9.3005
R12668 gnd.n4565 gnd.n4562 9.3005
R12669 gnd.n4613 gnd.n4612 9.3005
R12670 gnd.n2188 gnd.n2187 9.3005
R12671 gnd.n4629 gnd.n4628 9.3005
R12672 gnd.n4630 gnd.n2186 9.3005
R12673 gnd.n4632 gnd.n4631 9.3005
R12674 gnd.n2174 gnd.n2173 9.3005
R12675 gnd.n4648 gnd.n4647 9.3005
R12676 gnd.n4649 gnd.n2172 9.3005
R12677 gnd.n4651 gnd.n4650 9.3005
R12678 gnd.n1988 gnd.n1987 9.3005
R12679 gnd.n4674 gnd.n4673 9.3005
R12680 gnd.n4675 gnd.n1985 9.3005
R12681 gnd.n4686 gnd.n4685 9.3005
R12682 gnd.n4684 gnd.n1986 9.3005
R12683 gnd.n4683 gnd.n4682 9.3005
R12684 gnd.n4681 gnd.n4676 9.3005
R12685 gnd.n1927 gnd.n1926 9.3005
R12686 gnd.n4734 gnd.n4733 9.3005
R12687 gnd.n4735 gnd.n1924 9.3005
R12688 gnd.n4738 gnd.n4737 9.3005
R12689 gnd.n4736 gnd.n1925 9.3005
R12690 gnd.n1901 gnd.n1900 9.3005
R12691 gnd.n4803 gnd.n4802 9.3005
R12692 gnd.n4804 gnd.n1898 9.3005
R12693 gnd.n4807 gnd.n4806 9.3005
R12694 gnd.n4805 gnd.n1899 9.3005
R12695 gnd.n1871 gnd.n1870 9.3005
R12696 gnd.n4839 gnd.n4838 9.3005
R12697 gnd.n4840 gnd.n1869 9.3005
R12698 gnd.n4842 gnd.n4841 9.3005
R12699 gnd.n1848 gnd.n1847 9.3005
R12700 gnd.n4871 gnd.n4870 9.3005
R12701 gnd.n4872 gnd.n1845 9.3005
R12702 gnd.n4884 gnd.n4883 9.3005
R12703 gnd.n4882 gnd.n1846 9.3005
R12704 gnd.n4881 gnd.n4880 9.3005
R12705 gnd.n4879 gnd.n4873 9.3005
R12706 gnd.n4878 gnd.n4877 9.3005
R12707 gnd.n1809 gnd.n1808 9.3005
R12708 gnd.n5029 gnd.n5028 9.3005
R12709 gnd.n5030 gnd.n1806 9.3005
R12710 gnd.n5033 gnd.n5032 9.3005
R12711 gnd.n5031 gnd.n1807 9.3005
R12712 gnd.n1779 gnd.n1778 9.3005
R12713 gnd.n5065 gnd.n5064 9.3005
R12714 gnd.n5066 gnd.n1777 9.3005
R12715 gnd.n5068 gnd.n5067 9.3005
R12716 gnd.n1757 gnd.n1756 9.3005
R12717 gnd.n5092 gnd.n5091 9.3005
R12718 gnd.n5093 gnd.n1755 9.3005
R12719 gnd.n5095 gnd.n5094 9.3005
R12720 gnd.n1735 gnd.n1734 9.3005
R12721 gnd.n5122 gnd.n5121 9.3005
R12722 gnd.n5123 gnd.n1733 9.3005
R12723 gnd.n5125 gnd.n5124 9.3005
R12724 gnd.n1714 gnd.n1713 9.3005
R12725 gnd.n5152 gnd.n5151 9.3005
R12726 gnd.n5153 gnd.n1711 9.3005
R12727 gnd.n5156 gnd.n5155 9.3005
R12728 gnd.n5154 gnd.n1712 9.3005
R12729 gnd.n1685 gnd.n1684 9.3005
R12730 gnd.n5188 gnd.n5187 9.3005
R12731 gnd.n5189 gnd.n1683 9.3005
R12732 gnd.n5191 gnd.n5190 9.3005
R12733 gnd.n1661 gnd.n1660 9.3005
R12734 gnd.n5227 gnd.n5226 9.3005
R12735 gnd.n5228 gnd.n1659 9.3005
R12736 gnd.n5230 gnd.n5229 9.3005
R12737 gnd.n1605 gnd.n1604 9.3005
R12738 gnd.n5398 gnd.n5397 9.3005
R12739 gnd.n5399 gnd.n1603 9.3005
R12740 gnd.n5401 gnd.n5400 9.3005
R12741 gnd.n1590 gnd.n1589 9.3005
R12742 gnd.n5417 gnd.n5416 9.3005
R12743 gnd.n5418 gnd.n1588 9.3005
R12744 gnd.n5420 gnd.n5419 9.3005
R12745 gnd.n1577 gnd.n1576 9.3005
R12746 gnd.n5439 gnd.n5438 9.3005
R12747 gnd.n5440 gnd.n1575 9.3005
R12748 gnd.n5442 gnd.n5441 9.3005
R12749 gnd.n1476 gnd.n1475 9.3005
R12750 gnd.n5706 gnd.n5705 9.3005
R12751 gnd.n4611 gnd.n2200 9.3005
R12752 gnd.n6978 gnd.n6977 9.3005
R12753 gnd.n6979 gnd.n383 9.3005
R12754 gnd.n6981 gnd.n6980 9.3005
R12755 gnd.n367 gnd.n366 9.3005
R12756 gnd.n6994 gnd.n6993 9.3005
R12757 gnd.n6995 gnd.n365 9.3005
R12758 gnd.n6997 gnd.n6996 9.3005
R12759 gnd.n350 gnd.n349 9.3005
R12760 gnd.n7010 gnd.n7009 9.3005
R12761 gnd.n7011 gnd.n348 9.3005
R12762 gnd.n7013 gnd.n7012 9.3005
R12763 gnd.n332 gnd.n331 9.3005
R12764 gnd.n7026 gnd.n7025 9.3005
R12765 gnd.n7027 gnd.n330 9.3005
R12766 gnd.n7029 gnd.n7028 9.3005
R12767 gnd.n315 gnd.n314 9.3005
R12768 gnd.n7042 gnd.n7041 9.3005
R12769 gnd.n7043 gnd.n312 9.3005
R12770 gnd.n7046 gnd.n7045 9.3005
R12771 gnd.n7044 gnd.n313 9.3005
R12772 gnd.n295 gnd.n294 9.3005
R12773 gnd.n7061 gnd.n7060 9.3005
R12774 gnd.n7062 gnd.n293 9.3005
R12775 gnd.n7064 gnd.n7063 9.3005
R12776 gnd.n279 gnd.n278 9.3005
R12777 gnd.n7077 gnd.n7076 9.3005
R12778 gnd.n7079 gnd.n276 9.3005
R12779 gnd.n7081 gnd.n7080 9.3005
R12780 gnd.n264 gnd.n263 9.3005
R12781 gnd.n7093 gnd.n7092 9.3005
R12782 gnd.n7094 gnd.n262 9.3005
R12783 gnd.n7096 gnd.n7095 9.3005
R12784 gnd.n247 gnd.n246 9.3005
R12785 gnd.n7109 gnd.n7108 9.3005
R12786 gnd.n7110 gnd.n245 9.3005
R12787 gnd.n7112 gnd.n7111 9.3005
R12788 gnd.n231 gnd.n230 9.3005
R12789 gnd.n7125 gnd.n7124 9.3005
R12790 gnd.n7126 gnd.n229 9.3005
R12791 gnd.n7128 gnd.n7127 9.3005
R12792 gnd.n215 gnd.n214 9.3005
R12793 gnd.n7141 gnd.n7140 9.3005
R12794 gnd.n7142 gnd.n213 9.3005
R12795 gnd.n7144 gnd.n7143 9.3005
R12796 gnd.n201 gnd.n200 9.3005
R12797 gnd.n7157 gnd.n7156 9.3005
R12798 gnd.n7158 gnd.n199 9.3005
R12799 gnd.n7160 gnd.n7159 9.3005
R12800 gnd.n184 gnd.n183 9.3005
R12801 gnd.n7175 gnd.n7174 9.3005
R12802 gnd.n7176 gnd.n181 9.3005
R12803 gnd.n7246 gnd.n7245 9.3005
R12804 gnd.n7244 gnd.n182 9.3005
R12805 gnd.n385 gnd.n384 9.3005
R12806 gnd.n7241 gnd.n7177 9.3005
R12807 gnd.n7240 gnd.n7239 9.3005
R12808 gnd.n7238 gnd.n7182 9.3005
R12809 gnd.n7237 gnd.n7236 9.3005
R12810 gnd.n7235 gnd.n7183 9.3005
R12811 gnd.n7234 gnd.n7233 9.3005
R12812 gnd.n7232 gnd.n7190 9.3005
R12813 gnd.n7231 gnd.n7230 9.3005
R12814 gnd.n7229 gnd.n7191 9.3005
R12815 gnd.n7228 gnd.n7227 9.3005
R12816 gnd.n7226 gnd.n7198 9.3005
R12817 gnd.n7225 gnd.n7224 9.3005
R12818 gnd.n7223 gnd.n7199 9.3005
R12819 gnd.n7222 gnd.n7221 9.3005
R12820 gnd.n7220 gnd.n7206 9.3005
R12821 gnd.n7219 gnd.n7218 9.3005
R12822 gnd.n7217 gnd.n7207 9.3005
R12823 gnd.n7216 gnd.n7215 9.3005
R12824 gnd.n7243 gnd.n7242 9.3005
R12825 gnd.n6890 gnd.n471 9.3005
R12826 gnd.n6889 gnd.n6888 9.3005
R12827 gnd.n6887 gnd.n473 9.3005
R12828 gnd.n6886 gnd.n6885 9.3005
R12829 gnd.n6884 gnd.n476 9.3005
R12830 gnd.n6883 gnd.n6882 9.3005
R12831 gnd.n6881 gnd.n477 9.3005
R12832 gnd.n6880 gnd.n6879 9.3005
R12833 gnd.n6878 gnd.n480 9.3005
R12834 gnd.n6877 gnd.n6876 9.3005
R12835 gnd.n6875 gnd.n481 9.3005
R12836 gnd.n6874 gnd.n6873 9.3005
R12837 gnd.n6872 gnd.n484 9.3005
R12838 gnd.n6871 gnd.n6870 9.3005
R12839 gnd.n6869 gnd.n485 9.3005
R12840 gnd.n6868 gnd.n6867 9.3005
R12841 gnd.n6866 gnd.n488 9.3005
R12842 gnd.n6865 gnd.n6864 9.3005
R12843 gnd.n6863 gnd.n489 9.3005
R12844 gnd.n6862 gnd.n6861 9.3005
R12845 gnd.n6860 gnd.n492 9.3005
R12846 gnd.n6859 gnd.n6858 9.3005
R12847 gnd.n6857 gnd.n493 9.3005
R12848 gnd.n6856 gnd.n6855 9.3005
R12849 gnd.n6854 gnd.n6853 9.3005
R12850 gnd.n65 gnd.n63 9.3005
R12851 gnd.n7368 gnd.n7367 9.3005
R12852 gnd.n7366 gnd.n64 9.3005
R12853 gnd.n7365 gnd.n7364 9.3005
R12854 gnd.n7363 gnd.n69 9.3005
R12855 gnd.n7362 gnd.n7361 9.3005
R12856 gnd.n7360 gnd.n70 9.3005
R12857 gnd.n7359 gnd.n7358 9.3005
R12858 gnd.n7357 gnd.n74 9.3005
R12859 gnd.n7356 gnd.n7355 9.3005
R12860 gnd.n7354 gnd.n75 9.3005
R12861 gnd.n7353 gnd.n7352 9.3005
R12862 gnd.n7351 gnd.n79 9.3005
R12863 gnd.n7350 gnd.n7349 9.3005
R12864 gnd.n7348 gnd.n80 9.3005
R12865 gnd.n7347 gnd.n7346 9.3005
R12866 gnd.n7345 gnd.n84 9.3005
R12867 gnd.n7344 gnd.n7343 9.3005
R12868 gnd.n7342 gnd.n85 9.3005
R12869 gnd.n7341 gnd.n7340 9.3005
R12870 gnd.n7339 gnd.n89 9.3005
R12871 gnd.n7338 gnd.n7337 9.3005
R12872 gnd.n7336 gnd.n90 9.3005
R12873 gnd.n7335 gnd.n7334 9.3005
R12874 gnd.n7333 gnd.n94 9.3005
R12875 gnd.n7332 gnd.n7331 9.3005
R12876 gnd.n7330 gnd.n95 9.3005
R12877 gnd.n7329 gnd.n98 9.3005
R12878 gnd.n6892 gnd.n6891 9.3005
R12879 gnd.t154 gnd.n2648 9.24152
R12880 gnd.n2549 gnd.t101 9.24152
R12881 gnd.n3818 gnd.t81 9.24152
R12882 gnd.n4222 gnd.t64 9.24152
R12883 gnd.n4523 gnd.t186 9.24152
R12884 gnd.t255 gnd.n360 9.24152
R12885 gnd.n189 gnd.t18 9.24152
R12886 gnd.t146 gnd.t154 8.92286
R12887 gnd.n4730 gnd.n1930 8.92286
R12888 gnd.t22 gnd.n1921 8.92286
R12889 gnd.n4845 gnd.n1866 8.92286
R12890 gnd.n4894 gnd.n4893 8.92286
R12891 gnd.n5071 gnd.n1773 8.92286
R12892 gnd.n4964 gnd.n4963 8.92286
R12893 gnd.n5194 gnd.n1680 8.92286
R12894 gnd.n5326 gnd.n1607 8.92286
R12895 gnd.n3788 gnd.n3763 8.92171
R12896 gnd.n3756 gnd.n3731 8.92171
R12897 gnd.n3724 gnd.n3699 8.92171
R12898 gnd.n3693 gnd.n3668 8.92171
R12899 gnd.n3661 gnd.n3636 8.92171
R12900 gnd.n3629 gnd.n3604 8.92171
R12901 gnd.n3597 gnd.n3572 8.92171
R12902 gnd.n3566 gnd.n3541 8.92171
R12903 gnd.n5255 gnd.n5237 8.72777
R12904 gnd.n3292 gnd.t157 8.60421
R12905 gnd.n2720 gnd.n2704 8.43467
R12906 gnd.n46 gnd.n30 8.43467
R12907 gnd.n4308 gnd.n0 8.41456
R12908 gnd.n7370 gnd.n7369 8.41456
R12909 gnd.n1956 gnd.t114 8.28555
R12910 gnd.n4836 gnd.n1873 8.28555
R12911 gnd.n5007 gnd.n1824 8.28555
R12912 gnd.n5062 gnd.n1781 8.28555
R12913 gnd.n5130 gnd.n1728 8.28555
R12914 gnd.t95 gnd.n1654 8.28555
R12915 gnd.n3789 gnd.n3761 8.14595
R12916 gnd.n3757 gnd.n3729 8.14595
R12917 gnd.n3725 gnd.n3697 8.14595
R12918 gnd.n3694 gnd.n3666 8.14595
R12919 gnd.n3662 gnd.n3634 8.14595
R12920 gnd.n3630 gnd.n3602 8.14595
R12921 gnd.n3598 gnd.n3570 8.14595
R12922 gnd.n3567 gnd.n3539 8.14595
R12923 gnd.n3794 gnd.n3793 7.97301
R12924 gnd.t158 gnd.n2807 7.9669
R12925 gnd.n7217 gnd.n7216 7.75808
R12926 gnd.n5659 gnd.n1526 7.75808
R12927 gnd.n4566 gnd.n4565 7.75808
R12928 gnd.n4173 gnd.n4123 7.75808
R12929 gnd.n4828 gnd.n1873 7.64824
R12930 gnd.n1839 gnd.t3 7.64824
R12931 gnd.n4911 gnd.t169 7.64824
R12932 gnd.n5007 gnd.n5006 7.64824
R12933 gnd.n5054 gnd.n1781 7.64824
R12934 gnd.t13 gnd.n5061 7.64824
R12935 gnd.n5070 gnd.t5 7.64824
R12936 gnd.n5130 gnd.n5129 7.64824
R12937 gnd.n4924 gnd.t47 7.64824
R12938 gnd.n3201 gnd.t163 7.32958
R12939 gnd.n1977 gnd.n1976 7.30353
R12940 gnd.n5254 gnd.n5253 7.30353
R12941 gnd.n3161 gnd.n2880 7.01093
R12942 gnd.n2883 gnd.n2881 7.01093
R12943 gnd.n3171 gnd.n3170 7.01093
R12944 gnd.n3182 gnd.n2864 7.01093
R12945 gnd.n3181 gnd.n2867 7.01093
R12946 gnd.n3192 gnd.n2855 7.01093
R12947 gnd.n2858 gnd.n2856 7.01093
R12948 gnd.n3202 gnd.n3201 7.01093
R12949 gnd.n3212 gnd.n2836 7.01093
R12950 gnd.n3211 gnd.n2839 7.01093
R12951 gnd.n3220 gnd.n2830 7.01093
R12952 gnd.n3232 gnd.n2820 7.01093
R12953 gnd.n3242 gnd.n2805 7.01093
R12954 gnd.n3258 gnd.n3257 7.01093
R12955 gnd.n2807 gnd.n2744 7.01093
R12956 gnd.n3312 gnd.n2745 7.01093
R12957 gnd.n3306 gnd.n3305 7.01093
R12958 gnd.n2794 gnd.n2756 7.01093
R12959 gnd.n3298 gnd.n2767 7.01093
R12960 gnd.n2785 gnd.n2780 7.01093
R12961 gnd.n3292 gnd.n3291 7.01093
R12962 gnd.n3338 gnd.n2683 7.01093
R12963 gnd.n3337 gnd.n3336 7.01093
R12964 gnd.n3349 gnd.n3348 7.01093
R12965 gnd.n2676 gnd.n2668 7.01093
R12966 gnd.n3378 gnd.n2656 7.01093
R12967 gnd.n3377 gnd.n2659 7.01093
R12968 gnd.n3388 gnd.n2648 7.01093
R12969 gnd.n2649 gnd.n2637 7.01093
R12970 gnd.n3399 gnd.n2638 7.01093
R12971 gnd.n3423 gnd.n2629 7.01093
R12972 gnd.n3422 gnd.n2620 7.01093
R12973 gnd.n3445 gnd.n3444 7.01093
R12974 gnd.n3463 gnd.n2601 7.01093
R12975 gnd.n3462 gnd.n2604 7.01093
R12976 gnd.n3473 gnd.n2593 7.01093
R12977 gnd.n2594 gnd.n2581 7.01093
R12978 gnd.n3484 gnd.n2582 7.01093
R12979 gnd.n3511 gnd.n2565 7.01093
R12980 gnd.n3523 gnd.n3522 7.01093
R12981 gnd.n3505 gnd.n2558 7.01093
R12982 gnd.n3534 gnd.n3533 7.01093
R12983 gnd.n3806 gnd.n2546 7.01093
R12984 gnd.n3805 gnd.n2549 7.01093
R12985 gnd.n3818 gnd.n2538 7.01093
R12986 gnd.n2539 gnd.n2531 7.01093
R12987 gnd.n3828 gnd.n2457 7.01093
R12988 gnd.n4689 gnd.n4688 7.01093
R12989 gnd.n4731 gnd.n4730 7.01093
R12990 gnd.n1933 gnd.t22 7.01093
R12991 gnd.n4845 gnd.n4844 7.01093
R12992 gnd.n4901 gnd.t3 7.01093
R12993 gnd.n4893 gnd.n1839 7.01093
R12994 gnd.n5071 gnd.n5070 7.01093
R12995 gnd.t5 gnd.n1766 7.01093
R12996 gnd.n4964 gnd.n1745 7.01093
R12997 gnd.n5326 gnd.n1649 7.01093
R12998 gnd.n2839 gnd.t150 6.69227
R12999 gnd.n2659 gnd.t146 6.69227
R13000 gnd.n2429 gnd.t251 6.69227
R13001 gnd.n6021 gnd.n1109 6.69227
R13002 gnd.n4494 gnd.t201 6.69227
R13003 gnd.n4740 gnd.t314 6.69227
R13004 gnd.n5185 gnd.t312 6.69227
R13005 gnd.n7007 gnd.t209 6.69227
R13006 gnd.n7122 gnd.n233 6.69227
R13007 gnd.n7146 gnd.t213 6.69227
R13008 gnd.n5387 gnd.n5386 6.5566
R13009 gnd.n2090 gnd.n2089 6.5566
R13010 gnd.n2103 gnd.n2027 6.5566
R13011 gnd.n5265 gnd.n5264 6.5566
R13012 gnd.n4689 gnd.t29 6.37362
R13013 gnd.n4818 gnd.n4817 6.37362
R13014 gnd.n4867 gnd.t132 6.37362
R13015 gnd.n4999 gnd.n4998 6.37362
R13016 gnd.n5044 gnd.n5043 6.37362
R13017 gnd.t14 gnd.n5088 6.37362
R13018 gnd.n4954 gnd.n4953 6.37362
R13019 gnd.n5838 gnd.n1360 6.20656
R13020 gnd.n7292 gnd.n7289 6.20656
R13021 gnd.n3952 gnd.n3947 6.20656
R13022 gnd.n5638 gnd.n1541 6.20656
R13023 gnd.t148 gnd.n3268 6.05496
R13024 gnd.n3269 gnd.t165 6.05496
R13025 gnd.t172 gnd.n2683 6.05496
R13026 gnd.t160 gnd.n3433 6.05496
R13027 gnd.n4416 gnd.t211 6.05496
R13028 gnd.t131 gnd.t318 6.05496
R13029 gnd.t316 gnd.t7 6.05496
R13030 gnd.n7039 gnd.t240 6.05496
R13031 gnd.n3791 gnd.n3761 5.81868
R13032 gnd.n3759 gnd.n3729 5.81868
R13033 gnd.n3727 gnd.n3697 5.81868
R13034 gnd.n3696 gnd.n3666 5.81868
R13035 gnd.n3664 gnd.n3634 5.81868
R13036 gnd.n3632 gnd.n3602 5.81868
R13037 gnd.n3600 gnd.n3570 5.81868
R13038 gnd.n3569 gnd.n3539 5.81868
R13039 gnd.n1957 gnd.n1948 5.73631
R13040 gnd.n4868 gnd.n1850 5.73631
R13041 gnd.n4850 gnd.n4849 5.73631
R13042 gnd.t169 gnd.n1824 5.73631
R13043 gnd.n5062 gnd.t13 5.73631
R13044 gnd.n5089 gnd.n1759 5.73631
R13045 gnd.n5100 gnd.n1750 5.73631
R13046 gnd.n4920 gnd.n1665 5.73631
R13047 gnd.n5391 gnd.n440 5.62001
R13048 gnd.n2098 gnd.n2094 5.62001
R13049 gnd.n2099 gnd.n2098 5.62001
R13050 gnd.n5260 gnd.n440 5.62001
R13051 gnd.n3020 gnd.n3015 5.4308
R13052 gnd.n3836 gnd.n2524 5.4308
R13053 gnd.n3336 gnd.t159 5.41765
R13054 gnd.t162 gnd.n3359 5.41765
R13055 gnd.t139 gnd.n2613 5.41765
R13056 gnd.n4387 gnd.t226 5.41765
R13057 gnd.t174 gnd.n4809 5.41765
R13058 gnd.n5149 gnd.t11 5.41765
R13059 gnd.n6851 gnd.t257 5.41765
R13060 gnd.n1122 gnd.n1112 5.09899
R13061 gnd.n6014 gnd.n1125 5.09899
R13062 gnd.n4331 gnd.n4330 5.09899
R13063 gnd.n6008 gnd.n1136 5.09899
R13064 gnd.n4324 gnd.n2378 5.09899
R13065 gnd.n4344 gnd.n4343 5.09899
R13066 gnd.n4318 gnd.n2370 5.09899
R13067 gnd.n4355 gnd.n2373 5.09899
R13068 gnd.n4363 gnd.n2366 5.09899
R13069 gnd.n4362 gnd.n2360 5.09899
R13070 gnd.n4374 gnd.n4373 5.09899
R13071 gnd.n4387 gnd.n2349 5.09899
R13072 gnd.n4392 gnd.n2333 5.09899
R13073 gnd.n4431 gnd.n4430 5.09899
R13074 gnd.n5999 gnd.n1155 5.09899
R13075 gnd.n4399 gnd.n1164 5.09899
R13076 gnd.n4404 gnd.n1173 5.09899
R13077 gnd.n5987 gnd.n1176 5.09899
R13078 gnd.n4416 gnd.n1184 5.09899
R13079 gnd.n5981 gnd.n1187 5.09899
R13080 gnd.n4470 gnd.n4469 5.09899
R13081 gnd.n5975 gnd.n1197 5.09899
R13082 gnd.n4478 gnd.n1205 5.09899
R13083 gnd.n4486 gnd.n1215 5.09899
R13084 gnd.n5963 gnd.n1218 5.09899
R13085 gnd.n4494 gnd.n1226 5.09899
R13086 gnd.n5957 gnd.n1229 5.09899
R13087 gnd.n4523 gnd.n4522 5.09899
R13088 gnd.n5951 gnd.n1239 5.09899
R13089 gnd.n4502 gnd.n1247 5.09899
R13090 gnd.n5945 gnd.n1250 5.09899
R13091 gnd.n4511 gnd.n1258 5.09899
R13092 gnd.n5939 gnd.n1261 5.09899
R13093 gnd.n5856 gnd.n1268 5.09899
R13094 gnd.n5933 gnd.n1271 5.09899
R13095 gnd.t4 gnd.n4780 5.09899
R13096 gnd.n4799 gnd.n1905 5.09899
R13097 gnd.n5025 gnd.n1812 5.09899
R13098 gnd.n5037 gnd.n5036 5.09899
R13099 gnd.n5160 gnd.n5159 5.09899
R13100 gnd.n5177 gnd.t2 5.09899
R13101 gnd.n6894 gnd.n470 5.09899
R13102 gnd.n6975 gnd.n387 5.09899
R13103 gnd.n5617 gnd.n5616 5.09899
R13104 gnd.n6983 gnd.n378 5.09899
R13105 gnd.n5610 gnd.n381 5.09899
R13106 gnd.n6991 gnd.n369 5.09899
R13107 gnd.n5606 gnd.n372 5.09899
R13108 gnd.n6999 gnd.n360 5.09899
R13109 gnd.n5602 gnd.n363 5.09899
R13110 gnd.n7007 gnd.n352 5.09899
R13111 gnd.n5598 gnd.n5597 5.09899
R13112 gnd.n7015 gnd.n343 5.09899
R13113 gnd.n7023 gnd.n334 5.09899
R13114 gnd.n5518 gnd.n337 5.09899
R13115 gnd.n7031 gnd.n325 5.09899
R13116 gnd.n5522 gnd.n328 5.09899
R13117 gnd.n7039 gnd.n317 5.09899
R13118 gnd.n5583 gnd.n5582 5.09899
R13119 gnd.n7048 gnd.n306 5.09899
R13120 gnd.n5575 gnd.n5533 5.09899
R13121 gnd.n7058 gnd.n297 5.09899
R13122 gnd.n5555 gnd.n5554 5.09899
R13123 gnd.n7066 gnd.n288 5.09899
R13124 gnd.n6851 gnd.n291 5.09899
R13125 gnd.n7074 gnd.n281 5.09899
R13126 gnd.n6845 gnd.n284 5.09899
R13127 gnd.n7083 gnd.n272 5.09899
R13128 gnd.n6841 gnd.n274 5.09899
R13129 gnd.n7090 gnd.n266 5.09899
R13130 gnd.n6837 gnd.n6836 5.09899
R13131 gnd.n7098 gnd.n258 5.09899
R13132 gnd.n549 gnd.n260 5.09899
R13133 gnd.n7106 gnd.n249 5.09899
R13134 gnd.n545 gnd.n252 5.09899
R13135 gnd.n7114 gnd.n241 5.09899
R13136 gnd.n3789 gnd.n3788 5.04292
R13137 gnd.n3757 gnd.n3756 5.04292
R13138 gnd.n3725 gnd.n3724 5.04292
R13139 gnd.n3694 gnd.n3693 5.04292
R13140 gnd.n3662 gnd.n3661 5.04292
R13141 gnd.n3630 gnd.n3629 5.04292
R13142 gnd.n3598 gnd.n3597 5.04292
R13143 gnd.n3567 gnd.n3566 5.04292
R13144 gnd.n2736 gnd.n2735 4.82753
R13145 gnd.n62 gnd.n61 4.82753
R13146 gnd.n3299 gnd.t164 4.78034
R13147 gnd.n2638 gnd.t153 4.78034
R13148 gnd.n6008 gnd.t196 4.78034
R13149 gnd.n5993 gnd.t190 4.78034
R13150 gnd.t137 gnd.n2176 4.78034
R13151 gnd.n1594 gnd.t178 4.78034
R13152 gnd.n5576 gnd.t215 4.78034
R13153 gnd.n549 gnd.t268 4.78034
R13154 gnd.n2741 gnd.n2738 4.74817
R13155 gnd.n2791 gnd.n2689 4.74817
R13156 gnd.n2778 gnd.n2688 4.74817
R13157 gnd.n2687 gnd.n2686 4.74817
R13158 gnd.n2787 gnd.n2738 4.74817
R13159 gnd.n2788 gnd.n2689 4.74817
R13160 gnd.n2790 gnd.n2688 4.74817
R13161 gnd.n2777 gnd.n2687 4.74817
R13162 gnd.n7056 gnd.n7055 4.74817
R13163 gnd.n7072 gnd.n7070 4.74817
R13164 gnd.n7085 gnd.n270 4.74817
R13165 gnd.n7088 gnd.n7087 4.74817
R13166 gnd.n7055 gnd.n286 4.74817
R13167 gnd.n7070 gnd.n7069 4.74817
R13168 gnd.n7071 gnd.n270 4.74817
R13169 gnd.n7087 gnd.n7086 4.74817
R13170 gnd.n4341 gnd.n4340 4.74817
R13171 gnd.n4365 gnd.n2364 4.74817
R13172 gnd.n4371 gnd.n4367 4.74817
R13173 gnd.n4369 gnd.n4368 4.74817
R13174 gnd.n2331 gnd.n2329 4.74817
R13175 gnd.n5571 gnd.n5543 4.74817
R13176 gnd.n5569 gnd.n5546 4.74817
R13177 gnd.n5562 gnd.n5545 4.74817
R13178 gnd.n5558 gnd.n5544 4.74817
R13179 gnd.n6834 gnd.n555 4.74817
R13180 gnd.n5572 gnd.n5571 4.74817
R13181 gnd.n5569 gnd.n5568 4.74817
R13182 gnd.n5564 gnd.n5545 4.74817
R13183 gnd.n5561 gnd.n5544 4.74817
R13184 gnd.n5557 gnd.n555 4.74817
R13185 gnd.n6004 gnd.n6003 4.74817
R13186 gnd.n4360 gnd.n1147 4.74817
R13187 gnd.n4389 gnd.n1146 4.74817
R13188 gnd.n1149 gnd.n1145 4.74817
R13189 gnd.n6003 gnd.n1142 4.74817
R13190 gnd.n4357 gnd.n1147 4.74817
R13191 gnd.n4359 gnd.n1146 4.74817
R13192 gnd.n4390 gnd.n1145 4.74817
R13193 gnd.n4340 gnd.n4339 4.74817
R13194 gnd.n4338 gnd.n2364 4.74817
R13195 gnd.n4367 gnd.n4366 4.74817
R13196 gnd.n4370 gnd.n4369 4.74817
R13197 gnd.n2332 gnd.n2331 4.74817
R13198 gnd.n2720 gnd.n2719 4.7074
R13199 gnd.n46 gnd.n45 4.7074
R13200 gnd.n2736 gnd.n2720 4.65959
R13201 gnd.n62 gnd.n46 4.65959
R13202 gnd.n6938 gnd.n442 4.6132
R13203 gnd.n1305 gnd.n1302 4.6132
R13204 gnd.n4697 gnd.n1954 4.46168
R13205 gnd.n4723 gnd.n4722 4.46168
R13206 gnd.n4859 gnd.t135 4.46168
R13207 gnd.n4858 gnd.n4857 4.46168
R13208 gnd.n4887 gnd.n4886 4.46168
R13209 gnd.n5079 gnd.n5078 4.46168
R13210 gnd.n5098 gnd.n5097 4.46168
R13211 gnd.n5110 gnd.t166 4.46168
R13212 gnd.n5194 gnd.t78 4.46168
R13213 gnd.n5203 gnd.n5202 4.46168
R13214 gnd.n5233 gnd.n5232 4.46168
R13215 gnd.n5250 gnd.n5237 4.46111
R13216 gnd.n3774 gnd.n3770 4.38594
R13217 gnd.n3742 gnd.n3738 4.38594
R13218 gnd.n3710 gnd.n3706 4.38594
R13219 gnd.n3679 gnd.n3675 4.38594
R13220 gnd.n3647 gnd.n3643 4.38594
R13221 gnd.n3615 gnd.n3611 4.38594
R13222 gnd.n3583 gnd.n3579 4.38594
R13223 gnd.n3552 gnd.n3548 4.38594
R13224 gnd.n3785 gnd.n3763 4.26717
R13225 gnd.n3753 gnd.n3731 4.26717
R13226 gnd.n3721 gnd.n3699 4.26717
R13227 gnd.n3690 gnd.n3668 4.26717
R13228 gnd.n3658 gnd.n3636 4.26717
R13229 gnd.n3626 gnd.n3604 4.26717
R13230 gnd.n3594 gnd.n3572 4.26717
R13231 gnd.n3563 gnd.n3541 4.26717
R13232 gnd.n3243 gnd.t155 4.14303
R13233 gnd.n3473 gnd.t151 4.14303
R13234 gnd.n4272 gnd.t194 4.14303
R13235 gnd.n5969 gnd.t182 4.14303
R13236 gnd.t50 gnd.n1261 4.14303
R13237 gnd.n5617 gnd.t32 4.14303
R13238 gnd.n5512 gnd.t272 4.14303
R13239 gnd.n227 gnd.t228 4.14303
R13240 gnd.n3793 gnd.n3792 4.08274
R13241 gnd.n5386 gnd.n5385 4.05904
R13242 gnd.n2089 gnd.n2088 4.05904
R13243 gnd.n2106 gnd.n2027 4.05904
R13244 gnd.n5266 gnd.n5265 4.05904
R13245 gnd.n15 gnd.n7 3.99943
R13246 gnd.n4791 gnd.n4790 3.82437
R13247 gnd.n4811 gnd.t125 3.82437
R13248 gnd.n4762 gnd.n4761 3.82437
R13249 gnd.n5017 gnd.n5016 3.82437
R13250 gnd.n4997 gnd.t131 3.82437
R13251 gnd.t7 gnd.n1798 3.82437
R13252 gnd.n4986 gnd.n4985 3.82437
R13253 gnd.n5140 gnd.n5139 3.82437
R13254 gnd.n4950 gnd.t129 3.82437
R13255 gnd.n4942 gnd.n4941 3.82437
R13256 gnd.n3793 gnd.n3665 3.70378
R13257 gnd.n3316 gnd.n2737 3.65935
R13258 gnd.n15 gnd.n14 3.60163
R13259 gnd.t156 gnd.n2573 3.50571
R13260 gnd.n3784 gnd.n3765 3.49141
R13261 gnd.n3752 gnd.n3733 3.49141
R13262 gnd.n3720 gnd.n3701 3.49141
R13263 gnd.n3689 gnd.n3670 3.49141
R13264 gnd.n3657 gnd.n3638 3.49141
R13265 gnd.n3625 gnd.n3606 3.49141
R13266 gnd.n3593 gnd.n3574 3.49141
R13267 gnd.n3562 gnd.n3543 3.49141
R13268 gnd.n3512 gnd.n2573 3.18706
R13269 gnd.n4697 gnd.t114 3.18706
R13270 gnd.n4679 gnd.t123 3.18706
R13271 gnd.n4679 gnd.t43 3.18706
R13272 gnd.n1934 gnd.n1933 3.18706
R13273 gnd.n4773 gnd.t6 3.18706
R13274 gnd.t6 gnd.n4772 3.18706
R13275 gnd.n4754 gnd.n4753 3.18706
R13276 gnd.n4895 gnd.n1828 3.18706
R13277 gnd.n4978 gnd.n4977 3.18706
R13278 gnd.n5119 gnd.n1737 3.18706
R13279 gnd.n5167 gnd.t8 3.18706
R13280 gnd.t8 gnd.n5166 3.18706
R13281 gnd.n4933 gnd.n4932 3.18706
R13282 gnd.n5224 gnd.t25 3.18706
R13283 gnd.t68 gnd.n1649 3.18706
R13284 gnd.n2822 gnd.t155 2.8684
R13285 gnd.n4670 gnd.n2161 2.8684
R13286 gnd.n4708 gnd.t126 2.8684
R13287 gnd.t308 gnd.n5223 2.8684
R13288 gnd.n5394 gnd.n1627 2.8684
R13289 gnd.n2721 gnd.t292 2.82907
R13290 gnd.n2721 gnd.t245 2.82907
R13291 gnd.n2723 gnd.t279 2.82907
R13292 gnd.n2723 gnd.t181 2.82907
R13293 gnd.n2725 gnd.t205 2.82907
R13294 gnd.n2725 gnd.t191 2.82907
R13295 gnd.n2727 gnd.t189 2.82907
R13296 gnd.n2727 gnd.t301 2.82907
R13297 gnd.n2729 gnd.t197 2.82907
R13298 gnd.n2729 gnd.t237 2.82907
R13299 gnd.n2731 gnd.t271 2.82907
R13300 gnd.n2731 gnd.t223 2.82907
R13301 gnd.n2733 gnd.t252 2.82907
R13302 gnd.n2733 gnd.t195 2.82907
R13303 gnd.n2690 gnd.t183 2.82907
R13304 gnd.n2690 gnd.t221 2.82907
R13305 gnd.n2692 gnd.t224 2.82907
R13306 gnd.n2692 gnd.t293 2.82907
R13307 gnd.n2694 gnd.t217 2.82907
R13308 gnd.n2694 gnd.t208 2.82907
R13309 gnd.n2696 gnd.t259 2.82907
R13310 gnd.n2696 gnd.t247 2.82907
R13311 gnd.n2698 gnd.t298 2.82907
R13312 gnd.n2698 gnd.t230 2.82907
R13313 gnd.n2700 gnd.t242 2.82907
R13314 gnd.n2700 gnd.t270 2.82907
R13315 gnd.n2702 gnd.t253 2.82907
R13316 gnd.n2702 gnd.t218 2.82907
R13317 gnd.n2705 gnd.t300 2.82907
R13318 gnd.n2705 gnd.t202 2.82907
R13319 gnd.n2707 gnd.t212 2.82907
R13320 gnd.n2707 gnd.t274 2.82907
R13321 gnd.n2709 gnd.t199 2.82907
R13322 gnd.n2709 gnd.t307 2.82907
R13323 gnd.n2711 gnd.t236 2.82907
R13324 gnd.n2711 gnd.t227 2.82907
R13325 gnd.n2713 gnd.t282 2.82907
R13326 gnd.n2713 gnd.t207 2.82907
R13327 gnd.n2715 gnd.t220 2.82907
R13328 gnd.n2715 gnd.t244 2.82907
R13329 gnd.n2717 gnd.t260 2.82907
R13330 gnd.n2717 gnd.t200 2.82907
R13331 gnd.n59 gnd.t290 2.82907
R13332 gnd.n59 gnd.t214 2.82907
R13333 gnd.n57 gnd.t306 2.82907
R13334 gnd.n57 gnd.t233 2.82907
R13335 gnd.n55 gnd.t204 2.82907
R13336 gnd.n55 gnd.t299 2.82907
R13337 gnd.n53 gnd.t275 2.82907
R13338 gnd.n53 gnd.t285 2.82907
R13339 gnd.n51 gnd.t288 2.82907
R13340 gnd.n51 gnd.t304 2.82907
R13341 gnd.n49 gnd.t283 2.82907
R13342 gnd.n49 gnd.t241 2.82907
R13343 gnd.n47 gnd.t210 2.82907
R13344 gnd.n47 gnd.t273 2.82907
R13345 gnd.n28 gnd.t248 2.82907
R13346 gnd.n28 gnd.t302 2.82907
R13347 gnd.n26 gnd.t295 2.82907
R13348 gnd.n26 gnd.t276 2.82907
R13349 gnd.n24 gnd.t261 2.82907
R13350 gnd.n24 gnd.t291 2.82907
R13351 gnd.n22 gnd.t281 2.82907
R13352 gnd.n22 gnd.t287 2.82907
R13353 gnd.n20 gnd.t239 2.82907
R13354 gnd.n20 gnd.t185 2.82907
R13355 gnd.n18 gnd.t193 2.82907
R13356 gnd.n18 gnd.t267 2.82907
R13357 gnd.n16 gnd.t250 2.82907
R13358 gnd.n16 gnd.t305 2.82907
R13359 gnd.n43 gnd.t229 2.82907
R13360 gnd.n43 gnd.t289 2.82907
R13361 gnd.n41 gnd.t278 2.82907
R13362 gnd.n41 gnd.t249 2.82907
R13363 gnd.n39 gnd.t238 2.82907
R13364 gnd.n39 gnd.t269 2.82907
R13365 gnd.n37 gnd.t258 2.82907
R13366 gnd.n37 gnd.t266 2.82907
R13367 gnd.n35 gnd.t216 2.82907
R13368 gnd.n35 gnd.t303 2.82907
R13369 gnd.n33 gnd.t297 2.82907
R13370 gnd.n33 gnd.t243 2.82907
R13371 gnd.n31 gnd.t231 2.82907
R13372 gnd.n31 gnd.t294 2.82907
R13373 gnd.n3781 gnd.n3780 2.71565
R13374 gnd.n3749 gnd.n3748 2.71565
R13375 gnd.n3717 gnd.n3716 2.71565
R13376 gnd.n3686 gnd.n3685 2.71565
R13377 gnd.n3654 gnd.n3653 2.71565
R13378 gnd.n3622 gnd.n3621 2.71565
R13379 gnd.n3590 gnd.n3589 2.71565
R13380 gnd.n3559 gnd.n3558 2.71565
R13381 gnd.n2164 gnd.t29 2.54975
R13382 gnd.t43 gnd.n4678 2.54975
R13383 gnd.n4741 gnd.n1921 2.54975
R13384 gnd.n4781 gnd.t4 2.54975
R13385 gnd.n4835 gnd.n1875 2.54975
R13386 gnd.t128 gnd.n1875 2.54975
R13387 gnd.n4911 gnd.n4910 2.54975
R13388 gnd.n5061 gnd.n1783 2.54975
R13389 gnd.t130 gnd.n5118 2.54975
R13390 gnd.n5118 gnd.n1738 2.54975
R13391 gnd.n4937 gnd.t2 2.54975
R13392 gnd.n5184 gnd.n1688 2.54975
R13393 gnd.t78 gnd.n5193 2.54975
R13394 gnd.t47 gnd.n1675 2.54975
R13395 gnd.n4924 gnd.t25 2.54975
R13396 gnd.n3316 gnd.n2738 2.27742
R13397 gnd.n3316 gnd.n2689 2.27742
R13398 gnd.n3316 gnd.n2688 2.27742
R13399 gnd.n3316 gnd.n2687 2.27742
R13400 gnd.n7055 gnd.n255 2.27742
R13401 gnd.n7070 gnd.n255 2.27742
R13402 gnd.n270 gnd.n255 2.27742
R13403 gnd.n7087 gnd.n255 2.27742
R13404 gnd.n5571 gnd.n5570 2.27742
R13405 gnd.n5570 gnd.n5569 2.27742
R13406 gnd.n5570 gnd.n5545 2.27742
R13407 gnd.n5570 gnd.n5544 2.27742
R13408 gnd.n5570 gnd.n555 2.27742
R13409 gnd.n6003 gnd.n6002 2.27742
R13410 gnd.n6002 gnd.n1147 2.27742
R13411 gnd.n6002 gnd.n1146 2.27742
R13412 gnd.n6002 gnd.n1145 2.27742
R13413 gnd.n4340 gnd.n1144 2.27742
R13414 gnd.n2364 gnd.n1144 2.27742
R13415 gnd.n4367 gnd.n1144 2.27742
R13416 gnd.n4369 gnd.n1144 2.27742
R13417 gnd.n2331 gnd.n1144 2.27742
R13418 gnd.n3170 gnd.t39 2.23109
R13419 gnd.n2793 gnd.t164 2.23109
R13420 gnd.n4886 gnd.t170 2.23109
R13421 gnd.n5016 gnd.t318 2.23109
R13422 gnd.n4986 gnd.t316 2.23109
R13423 gnd.t141 gnd.n5079 2.23109
R13424 gnd.n3777 gnd.n3767 1.93989
R13425 gnd.n3745 gnd.n3735 1.93989
R13426 gnd.n3713 gnd.n3703 1.93989
R13427 gnd.n3682 gnd.n3672 1.93989
R13428 gnd.n3650 gnd.n3640 1.93989
R13429 gnd.n3618 gnd.n3608 1.93989
R13430 gnd.n3586 gnd.n3576 1.93989
R13431 gnd.n3555 gnd.n3545 1.93989
R13432 gnd.n4779 gnd.n1911 1.91244
R13433 gnd.n4829 gnd.n1880 1.91244
R13434 gnd.n5005 gnd.n1818 1.91244
R13435 gnd.n5055 gnd.n1787 1.91244
R13436 gnd.n5128 gnd.n5127 1.91244
R13437 gnd.n5178 gnd.n1692 1.91244
R13438 gnd.n4920 gnd.t95 1.91244
R13439 gnd.n1627 gnd.t98 1.91244
R13440 gnd.t133 gnd.n3181 1.59378
R13441 gnd.n3360 gnd.t162 1.59378
R13442 gnd.n2622 gnd.t139 1.59378
R13443 gnd.n4781 gnd.t314 1.59378
R13444 gnd.t167 gnd.n1866 1.59378
R13445 gnd.n4963 gnd.t0 1.59378
R13446 gnd.n4937 gnd.t312 1.59378
R13447 gnd.n4664 gnd.n1982 1.27512
R13448 gnd.n4721 gnd.n1940 1.27512
R13449 gnd.t125 gnd.n4810 1.27512
R13450 gnd.n4859 gnd.n1858 1.27512
R13451 gnd.n4902 gnd.n4901 1.27512
R13452 gnd.n5080 gnd.n1766 1.27512
R13453 gnd.n5110 gnd.n5109 1.27512
R13454 gnd.n5148 gnd.t129 1.27512
R13455 gnd.n5204 gnd.n1673 1.27512
R13456 gnd.n1657 gnd.n1656 1.27512
R13457 gnd.n3023 gnd.n3015 1.16414
R13458 gnd.n3839 gnd.n2524 1.16414
R13459 gnd.n3776 gnd.n3769 1.16414
R13460 gnd.n3744 gnd.n3737 1.16414
R13461 gnd.n3712 gnd.n3705 1.16414
R13462 gnd.n3681 gnd.n3674 1.16414
R13463 gnd.n3649 gnd.n3642 1.16414
R13464 gnd.n3617 gnd.n3610 1.16414
R13465 gnd.n3585 gnd.n3578 1.16414
R13466 gnd.n3554 gnd.n3547 1.16414
R13467 gnd.n6938 gnd.n6937 0.970197
R13468 gnd.n5897 gnd.n1302 0.970197
R13469 gnd.n3760 gnd.n3728 0.962709
R13470 gnd.n3792 gnd.n3760 0.962709
R13471 gnd.n3633 gnd.n3601 0.962709
R13472 gnd.n3665 gnd.n3633 0.962709
R13473 gnd.n3269 gnd.t148 0.956468
R13474 gnd.n3434 gnd.t160 0.956468
R13475 gnd.t222 gnd.n1122 0.956468
R13476 gnd.n2314 gnd.t182 0.956468
R13477 gnd.n4671 gnd.t176 0.956468
R13478 gnd.n1626 gnd.t9 0.956468
R13479 gnd.t272 gnd.n346 0.956468
R13480 gnd.t277 gnd.n241 0.956468
R13481 gnd.n2730 gnd.n2728 0.773756
R13482 gnd.n56 gnd.n54 0.773756
R13483 gnd.n2735 gnd.n2734 0.773756
R13484 gnd.n2734 gnd.n2732 0.773756
R13485 gnd.n2732 gnd.n2730 0.773756
R13486 gnd.n2728 gnd.n2726 0.773756
R13487 gnd.n2726 gnd.n2724 0.773756
R13488 gnd.n2724 gnd.n2722 0.773756
R13489 gnd.n50 gnd.n48 0.773756
R13490 gnd.n52 gnd.n50 0.773756
R13491 gnd.n54 gnd.n52 0.773756
R13492 gnd.n58 gnd.n56 0.773756
R13493 gnd.n60 gnd.n58 0.773756
R13494 gnd.n61 gnd.n60 0.773756
R13495 gnd.n2 gnd.n1 0.672012
R13496 gnd.n3 gnd.n2 0.672012
R13497 gnd.n4 gnd.n3 0.672012
R13498 gnd.n5 gnd.n4 0.672012
R13499 gnd.n6 gnd.n5 0.672012
R13500 gnd.n7 gnd.n6 0.672012
R13501 gnd.n9 gnd.n8 0.672012
R13502 gnd.n10 gnd.n9 0.672012
R13503 gnd.n11 gnd.n10 0.672012
R13504 gnd.n12 gnd.n11 0.672012
R13505 gnd.n13 gnd.n12 0.672012
R13506 gnd.n14 gnd.n13 0.672012
R13507 gnd.n1940 gnd.t85 0.637812
R13508 gnd.n4800 gnd.n1903 0.637812
R13509 gnd.n4809 gnd.n1888 0.637812
R13510 gnd.n4761 gnd.t136 0.637812
R13511 gnd.n5026 gnd.n1811 0.637812
R13512 gnd.n5035 gnd.n1795 0.637812
R13513 gnd.n5140 gnd.t143 0.637812
R13514 gnd.n5149 gnd.n1716 0.637812
R13515 gnd.n5158 gnd.n1700 0.637812
R13516 gnd gnd.n0 0.59317
R13517 gnd.n2704 gnd.n2703 0.573776
R13518 gnd.n2703 gnd.n2701 0.573776
R13519 gnd.n2701 gnd.n2699 0.573776
R13520 gnd.n2699 gnd.n2697 0.573776
R13521 gnd.n2697 gnd.n2695 0.573776
R13522 gnd.n2695 gnd.n2693 0.573776
R13523 gnd.n2693 gnd.n2691 0.573776
R13524 gnd.n2719 gnd.n2718 0.573776
R13525 gnd.n2718 gnd.n2716 0.573776
R13526 gnd.n2716 gnd.n2714 0.573776
R13527 gnd.n2714 gnd.n2712 0.573776
R13528 gnd.n2712 gnd.n2710 0.573776
R13529 gnd.n2710 gnd.n2708 0.573776
R13530 gnd.n2708 gnd.n2706 0.573776
R13531 gnd.n19 gnd.n17 0.573776
R13532 gnd.n21 gnd.n19 0.573776
R13533 gnd.n23 gnd.n21 0.573776
R13534 gnd.n25 gnd.n23 0.573776
R13535 gnd.n27 gnd.n25 0.573776
R13536 gnd.n29 gnd.n27 0.573776
R13537 gnd.n30 gnd.n29 0.573776
R13538 gnd.n34 gnd.n32 0.573776
R13539 gnd.n36 gnd.n34 0.573776
R13540 gnd.n38 gnd.n36 0.573776
R13541 gnd.n40 gnd.n38 0.573776
R13542 gnd.n42 gnd.n40 0.573776
R13543 gnd.n44 gnd.n42 0.573776
R13544 gnd.n45 gnd.n44 0.573776
R13545 gnd.n7371 gnd.n7370 0.553533
R13546 gnd.n5570 gnd.n255 0.548625
R13547 gnd.n6002 gnd.n1144 0.548625
R13548 gnd.n4611 gnd.n4610 0.523366
R13549 gnd.n5705 gnd.n5704 0.523366
R13550 gnd.n4174 gnd.n4169 0.505073
R13551 gnd.n4211 gnd.n4210 0.505073
R13552 gnd.n7244 gnd.n7243 0.505073
R13553 gnd.n7215 gnd.n98 0.505073
R13554 gnd.n7324 gnd.n7323 0.492878
R13555 gnd.n7253 gnd.n7252 0.492878
R13556 gnd.n6898 gnd.n468 0.492878
R13557 gnd.n6971 gnd.n6970 0.492878
R13558 gnd.n5930 gnd.n5929 0.492878
R13559 gnd.n5861 gnd.n5860 0.492878
R13560 gnd.n4064 gnd.n4063 0.492878
R13561 gnd.n4217 gnd.n2455 0.492878
R13562 gnd.n5634 gnd.n1469 0.489829
R13563 gnd.n5834 gnd.n5833 0.489829
R13564 gnd.n3496 gnd.n2528 0.486781
R13565 gnd.n3072 gnd.n3071 0.48678
R13566 gnd.n3813 gnd.n2482 0.480683
R13567 gnd.n3156 gnd.n3155 0.480683
R13568 gnd.n6193 gnd.n6192 0.480683
R13569 gnd.n6613 gnd.n6612 0.480683
R13570 gnd.n6826 gnd.n6825 0.480683
R13571 gnd.n2385 gnd.n1107 0.480683
R13572 gnd.n4609 gnd.n1266 0.404992
R13573 gnd.n5703 gnd.n384 0.404992
R13574 gnd.n5841 gnd.n1360 0.388379
R13575 gnd.n3773 gnd.n3772 0.388379
R13576 gnd.n3741 gnd.n3740 0.388379
R13577 gnd.n3709 gnd.n3708 0.388379
R13578 gnd.n3678 gnd.n3677 0.388379
R13579 gnd.n3646 gnd.n3645 0.388379
R13580 gnd.n3614 gnd.n3613 0.388379
R13581 gnd.n3582 gnd.n3581 0.388379
R13582 gnd.n3551 gnd.n3550 0.388379
R13583 gnd.n7293 gnd.n7292 0.388379
R13584 gnd.n4010 gnd.n3952 0.388379
R13585 gnd.n1541 gnd.n1537 0.388379
R13586 gnd.n7371 gnd.n15 0.374463
R13587 gnd.n2584 gnd.t156 0.319156
R13588 gnd.n4363 gnd.t188 0.319156
R13589 gnd.n4403 gnd.t190 0.319156
R13590 gnd.n4617 gnd.t91 0.319156
R13591 gnd.n5446 gnd.t74 0.319156
R13592 gnd.t215 gnd.n309 0.319156
R13593 gnd.t265 gnd.n272 0.319156
R13594 gnd.n2990 gnd.n2968 0.311721
R13595 gnd gnd.n7371 0.295112
R13596 gnd.n5852 gnd.n5851 0.27489
R13597 gnd.n6891 gnd.n472 0.27489
R13598 gnd.n3884 gnd.n3883 0.268793
R13599 gnd.n3883 gnd.n3882 0.241354
R13600 gnd.n442 gnd.n439 0.229039
R13601 gnd.n445 gnd.n442 0.229039
R13602 gnd.n1305 gnd.n1304 0.229039
R13603 gnd.n1306 gnd.n1305 0.229039
R13604 gnd.n3144 gnd.n2943 0.206293
R13605 gnd.n2737 gnd.n0 0.169152
R13606 gnd.n3790 gnd.n3762 0.155672
R13607 gnd.n3783 gnd.n3762 0.155672
R13608 gnd.n3783 gnd.n3782 0.155672
R13609 gnd.n3782 gnd.n3766 0.155672
R13610 gnd.n3775 gnd.n3766 0.155672
R13611 gnd.n3775 gnd.n3774 0.155672
R13612 gnd.n3758 gnd.n3730 0.155672
R13613 gnd.n3751 gnd.n3730 0.155672
R13614 gnd.n3751 gnd.n3750 0.155672
R13615 gnd.n3750 gnd.n3734 0.155672
R13616 gnd.n3743 gnd.n3734 0.155672
R13617 gnd.n3743 gnd.n3742 0.155672
R13618 gnd.n3726 gnd.n3698 0.155672
R13619 gnd.n3719 gnd.n3698 0.155672
R13620 gnd.n3719 gnd.n3718 0.155672
R13621 gnd.n3718 gnd.n3702 0.155672
R13622 gnd.n3711 gnd.n3702 0.155672
R13623 gnd.n3711 gnd.n3710 0.155672
R13624 gnd.n3695 gnd.n3667 0.155672
R13625 gnd.n3688 gnd.n3667 0.155672
R13626 gnd.n3688 gnd.n3687 0.155672
R13627 gnd.n3687 gnd.n3671 0.155672
R13628 gnd.n3680 gnd.n3671 0.155672
R13629 gnd.n3680 gnd.n3679 0.155672
R13630 gnd.n3663 gnd.n3635 0.155672
R13631 gnd.n3656 gnd.n3635 0.155672
R13632 gnd.n3656 gnd.n3655 0.155672
R13633 gnd.n3655 gnd.n3639 0.155672
R13634 gnd.n3648 gnd.n3639 0.155672
R13635 gnd.n3648 gnd.n3647 0.155672
R13636 gnd.n3631 gnd.n3603 0.155672
R13637 gnd.n3624 gnd.n3603 0.155672
R13638 gnd.n3624 gnd.n3623 0.155672
R13639 gnd.n3623 gnd.n3607 0.155672
R13640 gnd.n3616 gnd.n3607 0.155672
R13641 gnd.n3616 gnd.n3615 0.155672
R13642 gnd.n3599 gnd.n3571 0.155672
R13643 gnd.n3592 gnd.n3571 0.155672
R13644 gnd.n3592 gnd.n3591 0.155672
R13645 gnd.n3591 gnd.n3575 0.155672
R13646 gnd.n3584 gnd.n3575 0.155672
R13647 gnd.n3584 gnd.n3583 0.155672
R13648 gnd.n3568 gnd.n3540 0.155672
R13649 gnd.n3561 gnd.n3540 0.155672
R13650 gnd.n3561 gnd.n3560 0.155672
R13651 gnd.n3560 gnd.n3544 0.155672
R13652 gnd.n3553 gnd.n3544 0.155672
R13653 gnd.n3553 gnd.n3552 0.155672
R13654 gnd.n3915 gnd.n2482 0.152939
R13655 gnd.n3915 gnd.n3914 0.152939
R13656 gnd.n3914 gnd.n3913 0.152939
R13657 gnd.n3913 gnd.n2484 0.152939
R13658 gnd.n2485 gnd.n2484 0.152939
R13659 gnd.n2486 gnd.n2485 0.152939
R13660 gnd.n2487 gnd.n2486 0.152939
R13661 gnd.n2488 gnd.n2487 0.152939
R13662 gnd.n2489 gnd.n2488 0.152939
R13663 gnd.n2490 gnd.n2489 0.152939
R13664 gnd.n2491 gnd.n2490 0.152939
R13665 gnd.n2492 gnd.n2491 0.152939
R13666 gnd.n2493 gnd.n2492 0.152939
R13667 gnd.n2494 gnd.n2493 0.152939
R13668 gnd.n3885 gnd.n2494 0.152939
R13669 gnd.n3885 gnd.n3884 0.152939
R13670 gnd.n3157 gnd.n3156 0.152939
R13671 gnd.n3157 gnd.n2861 0.152939
R13672 gnd.n3185 gnd.n2861 0.152939
R13673 gnd.n3186 gnd.n3185 0.152939
R13674 gnd.n3187 gnd.n3186 0.152939
R13675 gnd.n3188 gnd.n3187 0.152939
R13676 gnd.n3188 gnd.n2833 0.152939
R13677 gnd.n3215 gnd.n2833 0.152939
R13678 gnd.n3216 gnd.n3215 0.152939
R13679 gnd.n3217 gnd.n3216 0.152939
R13680 gnd.n3217 gnd.n2811 0.152939
R13681 gnd.n3246 gnd.n2811 0.152939
R13682 gnd.n3247 gnd.n3246 0.152939
R13683 gnd.n3248 gnd.n3247 0.152939
R13684 gnd.n3249 gnd.n3248 0.152939
R13685 gnd.n3251 gnd.n3249 0.152939
R13686 gnd.n3251 gnd.n3250 0.152939
R13687 gnd.n3250 gnd.n2760 0.152939
R13688 gnd.n2761 gnd.n2760 0.152939
R13689 gnd.n2762 gnd.n2761 0.152939
R13690 gnd.n2781 gnd.n2762 0.152939
R13691 gnd.n2782 gnd.n2781 0.152939
R13692 gnd.n2782 gnd.n2680 0.152939
R13693 gnd.n3341 gnd.n2680 0.152939
R13694 gnd.n3342 gnd.n3341 0.152939
R13695 gnd.n3343 gnd.n3342 0.152939
R13696 gnd.n3344 gnd.n3343 0.152939
R13697 gnd.n3344 gnd.n2653 0.152939
R13698 gnd.n3381 gnd.n2653 0.152939
R13699 gnd.n3382 gnd.n3381 0.152939
R13700 gnd.n3383 gnd.n3382 0.152939
R13701 gnd.n3384 gnd.n3383 0.152939
R13702 gnd.n3384 gnd.n2626 0.152939
R13703 gnd.n3426 gnd.n2626 0.152939
R13704 gnd.n3427 gnd.n3426 0.152939
R13705 gnd.n3428 gnd.n3427 0.152939
R13706 gnd.n3429 gnd.n3428 0.152939
R13707 gnd.n3429 gnd.n2598 0.152939
R13708 gnd.n3466 gnd.n2598 0.152939
R13709 gnd.n3467 gnd.n3466 0.152939
R13710 gnd.n3468 gnd.n3467 0.152939
R13711 gnd.n3469 gnd.n3468 0.152939
R13712 gnd.n3469 gnd.n2570 0.152939
R13713 gnd.n3515 gnd.n2570 0.152939
R13714 gnd.n3516 gnd.n3515 0.152939
R13715 gnd.n3517 gnd.n3516 0.152939
R13716 gnd.n3518 gnd.n3517 0.152939
R13717 gnd.n3518 gnd.n2543 0.152939
R13718 gnd.n3809 gnd.n2543 0.152939
R13719 gnd.n3810 gnd.n3809 0.152939
R13720 gnd.n3811 gnd.n3810 0.152939
R13721 gnd.n3812 gnd.n3811 0.152939
R13722 gnd.n3813 gnd.n3812 0.152939
R13723 gnd.n3155 gnd.n2885 0.152939
R13724 gnd.n2906 gnd.n2885 0.152939
R13725 gnd.n2907 gnd.n2906 0.152939
R13726 gnd.n2913 gnd.n2907 0.152939
R13727 gnd.n2914 gnd.n2913 0.152939
R13728 gnd.n2915 gnd.n2914 0.152939
R13729 gnd.n2915 gnd.n2904 0.152939
R13730 gnd.n2923 gnd.n2904 0.152939
R13731 gnd.n2924 gnd.n2923 0.152939
R13732 gnd.n2925 gnd.n2924 0.152939
R13733 gnd.n2925 gnd.n2902 0.152939
R13734 gnd.n2933 gnd.n2902 0.152939
R13735 gnd.n2934 gnd.n2933 0.152939
R13736 gnd.n2935 gnd.n2934 0.152939
R13737 gnd.n2935 gnd.n2900 0.152939
R13738 gnd.n2943 gnd.n2900 0.152939
R13739 gnd.n3882 gnd.n2499 0.152939
R13740 gnd.n2501 gnd.n2499 0.152939
R13741 gnd.n2502 gnd.n2501 0.152939
R13742 gnd.n2503 gnd.n2502 0.152939
R13743 gnd.n2504 gnd.n2503 0.152939
R13744 gnd.n2505 gnd.n2504 0.152939
R13745 gnd.n2506 gnd.n2505 0.152939
R13746 gnd.n2507 gnd.n2506 0.152939
R13747 gnd.n2508 gnd.n2507 0.152939
R13748 gnd.n2509 gnd.n2508 0.152939
R13749 gnd.n2510 gnd.n2509 0.152939
R13750 gnd.n2511 gnd.n2510 0.152939
R13751 gnd.n2512 gnd.n2511 0.152939
R13752 gnd.n2513 gnd.n2512 0.152939
R13753 gnd.n2514 gnd.n2513 0.152939
R13754 gnd.n2515 gnd.n2514 0.152939
R13755 gnd.n2516 gnd.n2515 0.152939
R13756 gnd.n2517 gnd.n2516 0.152939
R13757 gnd.n2518 gnd.n2517 0.152939
R13758 gnd.n2519 gnd.n2518 0.152939
R13759 gnd.n2520 gnd.n2519 0.152939
R13760 gnd.n2521 gnd.n2520 0.152939
R13761 gnd.n2525 gnd.n2521 0.152939
R13762 gnd.n2526 gnd.n2525 0.152939
R13763 gnd.n2527 gnd.n2526 0.152939
R13764 gnd.n2528 gnd.n2527 0.152939
R13765 gnd.n3318 gnd.n3317 0.152939
R13766 gnd.n3319 gnd.n3318 0.152939
R13767 gnd.n3320 gnd.n3319 0.152939
R13768 gnd.n3321 gnd.n3320 0.152939
R13769 gnd.n3322 gnd.n3321 0.152939
R13770 gnd.n3323 gnd.n3322 0.152939
R13771 gnd.n3323 gnd.n2634 0.152939
R13772 gnd.n3402 gnd.n2634 0.152939
R13773 gnd.n3403 gnd.n3402 0.152939
R13774 gnd.n3404 gnd.n3403 0.152939
R13775 gnd.n3405 gnd.n3404 0.152939
R13776 gnd.n3406 gnd.n3405 0.152939
R13777 gnd.n3407 gnd.n3406 0.152939
R13778 gnd.n3408 gnd.n3407 0.152939
R13779 gnd.n3409 gnd.n3408 0.152939
R13780 gnd.n3410 gnd.n3409 0.152939
R13781 gnd.n3410 gnd.n2578 0.152939
R13782 gnd.n3487 gnd.n2578 0.152939
R13783 gnd.n3488 gnd.n3487 0.152939
R13784 gnd.n3489 gnd.n3488 0.152939
R13785 gnd.n3490 gnd.n3489 0.152939
R13786 gnd.n3491 gnd.n3490 0.152939
R13787 gnd.n3492 gnd.n3491 0.152939
R13788 gnd.n3493 gnd.n3492 0.152939
R13789 gnd.n3494 gnd.n3493 0.152939
R13790 gnd.n3495 gnd.n3494 0.152939
R13791 gnd.n3497 gnd.n3495 0.152939
R13792 gnd.n3497 gnd.n3496 0.152939
R13793 gnd.n3073 gnd.n3072 0.152939
R13794 gnd.n3073 gnd.n2963 0.152939
R13795 gnd.n3088 gnd.n2963 0.152939
R13796 gnd.n3089 gnd.n3088 0.152939
R13797 gnd.n3090 gnd.n3089 0.152939
R13798 gnd.n3090 gnd.n2951 0.152939
R13799 gnd.n3104 gnd.n2951 0.152939
R13800 gnd.n3105 gnd.n3104 0.152939
R13801 gnd.n3106 gnd.n3105 0.152939
R13802 gnd.n3107 gnd.n3106 0.152939
R13803 gnd.n3108 gnd.n3107 0.152939
R13804 gnd.n3109 gnd.n3108 0.152939
R13805 gnd.n3110 gnd.n3109 0.152939
R13806 gnd.n3111 gnd.n3110 0.152939
R13807 gnd.n3112 gnd.n3111 0.152939
R13808 gnd.n3113 gnd.n3112 0.152939
R13809 gnd.n3114 gnd.n3113 0.152939
R13810 gnd.n3115 gnd.n3114 0.152939
R13811 gnd.n3116 gnd.n3115 0.152939
R13812 gnd.n3117 gnd.n3116 0.152939
R13813 gnd.n3118 gnd.n3117 0.152939
R13814 gnd.n3118 gnd.n2817 0.152939
R13815 gnd.n3235 gnd.n2817 0.152939
R13816 gnd.n3236 gnd.n3235 0.152939
R13817 gnd.n3237 gnd.n3236 0.152939
R13818 gnd.n3238 gnd.n3237 0.152939
R13819 gnd.n3238 gnd.n2739 0.152939
R13820 gnd.n3315 gnd.n2739 0.152939
R13821 gnd.n2991 gnd.n2990 0.152939
R13822 gnd.n2992 gnd.n2991 0.152939
R13823 gnd.n2993 gnd.n2992 0.152939
R13824 gnd.n2994 gnd.n2993 0.152939
R13825 gnd.n2995 gnd.n2994 0.152939
R13826 gnd.n2996 gnd.n2995 0.152939
R13827 gnd.n2997 gnd.n2996 0.152939
R13828 gnd.n2998 gnd.n2997 0.152939
R13829 gnd.n2999 gnd.n2998 0.152939
R13830 gnd.n3000 gnd.n2999 0.152939
R13831 gnd.n3001 gnd.n3000 0.152939
R13832 gnd.n3002 gnd.n3001 0.152939
R13833 gnd.n3003 gnd.n3002 0.152939
R13834 gnd.n3004 gnd.n3003 0.152939
R13835 gnd.n3005 gnd.n3004 0.152939
R13836 gnd.n3006 gnd.n3005 0.152939
R13837 gnd.n3007 gnd.n3006 0.152939
R13838 gnd.n3008 gnd.n3007 0.152939
R13839 gnd.n3009 gnd.n3008 0.152939
R13840 gnd.n3010 gnd.n3009 0.152939
R13841 gnd.n3011 gnd.n3010 0.152939
R13842 gnd.n3012 gnd.n3011 0.152939
R13843 gnd.n3016 gnd.n3012 0.152939
R13844 gnd.n3017 gnd.n3016 0.152939
R13845 gnd.n3017 gnd.n2974 0.152939
R13846 gnd.n3071 gnd.n2974 0.152939
R13847 gnd.n6194 gnd.n6193 0.152939
R13848 gnd.n6194 gnd.n934 0.152939
R13849 gnd.n6202 gnd.n934 0.152939
R13850 gnd.n6203 gnd.n6202 0.152939
R13851 gnd.n6204 gnd.n6203 0.152939
R13852 gnd.n6204 gnd.n928 0.152939
R13853 gnd.n6212 gnd.n928 0.152939
R13854 gnd.n6213 gnd.n6212 0.152939
R13855 gnd.n6214 gnd.n6213 0.152939
R13856 gnd.n6214 gnd.n922 0.152939
R13857 gnd.n6222 gnd.n922 0.152939
R13858 gnd.n6223 gnd.n6222 0.152939
R13859 gnd.n6224 gnd.n6223 0.152939
R13860 gnd.n6224 gnd.n916 0.152939
R13861 gnd.n6232 gnd.n916 0.152939
R13862 gnd.n6233 gnd.n6232 0.152939
R13863 gnd.n6234 gnd.n6233 0.152939
R13864 gnd.n6234 gnd.n910 0.152939
R13865 gnd.n6242 gnd.n910 0.152939
R13866 gnd.n6243 gnd.n6242 0.152939
R13867 gnd.n6244 gnd.n6243 0.152939
R13868 gnd.n6244 gnd.n904 0.152939
R13869 gnd.n6252 gnd.n904 0.152939
R13870 gnd.n6253 gnd.n6252 0.152939
R13871 gnd.n6254 gnd.n6253 0.152939
R13872 gnd.n6254 gnd.n898 0.152939
R13873 gnd.n6262 gnd.n898 0.152939
R13874 gnd.n6263 gnd.n6262 0.152939
R13875 gnd.n6264 gnd.n6263 0.152939
R13876 gnd.n6264 gnd.n892 0.152939
R13877 gnd.n6272 gnd.n892 0.152939
R13878 gnd.n6273 gnd.n6272 0.152939
R13879 gnd.n6274 gnd.n6273 0.152939
R13880 gnd.n6274 gnd.n886 0.152939
R13881 gnd.n6282 gnd.n886 0.152939
R13882 gnd.n6283 gnd.n6282 0.152939
R13883 gnd.n6284 gnd.n6283 0.152939
R13884 gnd.n6284 gnd.n880 0.152939
R13885 gnd.n6292 gnd.n880 0.152939
R13886 gnd.n6293 gnd.n6292 0.152939
R13887 gnd.n6294 gnd.n6293 0.152939
R13888 gnd.n6294 gnd.n874 0.152939
R13889 gnd.n6302 gnd.n874 0.152939
R13890 gnd.n6303 gnd.n6302 0.152939
R13891 gnd.n6304 gnd.n6303 0.152939
R13892 gnd.n6304 gnd.n868 0.152939
R13893 gnd.n6312 gnd.n868 0.152939
R13894 gnd.n6313 gnd.n6312 0.152939
R13895 gnd.n6314 gnd.n6313 0.152939
R13896 gnd.n6314 gnd.n862 0.152939
R13897 gnd.n6322 gnd.n862 0.152939
R13898 gnd.n6323 gnd.n6322 0.152939
R13899 gnd.n6324 gnd.n6323 0.152939
R13900 gnd.n6324 gnd.n856 0.152939
R13901 gnd.n6332 gnd.n856 0.152939
R13902 gnd.n6333 gnd.n6332 0.152939
R13903 gnd.n6334 gnd.n6333 0.152939
R13904 gnd.n6334 gnd.n850 0.152939
R13905 gnd.n6342 gnd.n850 0.152939
R13906 gnd.n6343 gnd.n6342 0.152939
R13907 gnd.n6344 gnd.n6343 0.152939
R13908 gnd.n6344 gnd.n844 0.152939
R13909 gnd.n6352 gnd.n844 0.152939
R13910 gnd.n6353 gnd.n6352 0.152939
R13911 gnd.n6354 gnd.n6353 0.152939
R13912 gnd.n6354 gnd.n838 0.152939
R13913 gnd.n6362 gnd.n838 0.152939
R13914 gnd.n6363 gnd.n6362 0.152939
R13915 gnd.n6364 gnd.n6363 0.152939
R13916 gnd.n6364 gnd.n832 0.152939
R13917 gnd.n6372 gnd.n832 0.152939
R13918 gnd.n6373 gnd.n6372 0.152939
R13919 gnd.n6374 gnd.n6373 0.152939
R13920 gnd.n6374 gnd.n826 0.152939
R13921 gnd.n6382 gnd.n826 0.152939
R13922 gnd.n6383 gnd.n6382 0.152939
R13923 gnd.n6384 gnd.n6383 0.152939
R13924 gnd.n6384 gnd.n820 0.152939
R13925 gnd.n6392 gnd.n820 0.152939
R13926 gnd.n6393 gnd.n6392 0.152939
R13927 gnd.n6394 gnd.n6393 0.152939
R13928 gnd.n6394 gnd.n814 0.152939
R13929 gnd.n6402 gnd.n814 0.152939
R13930 gnd.n6403 gnd.n6402 0.152939
R13931 gnd.n6404 gnd.n6403 0.152939
R13932 gnd.n6404 gnd.n808 0.152939
R13933 gnd.n6412 gnd.n808 0.152939
R13934 gnd.n6413 gnd.n6412 0.152939
R13935 gnd.n6414 gnd.n6413 0.152939
R13936 gnd.n6414 gnd.n802 0.152939
R13937 gnd.n6422 gnd.n802 0.152939
R13938 gnd.n6423 gnd.n6422 0.152939
R13939 gnd.n6424 gnd.n6423 0.152939
R13940 gnd.n6424 gnd.n796 0.152939
R13941 gnd.n6432 gnd.n796 0.152939
R13942 gnd.n6433 gnd.n6432 0.152939
R13943 gnd.n6434 gnd.n6433 0.152939
R13944 gnd.n6434 gnd.n790 0.152939
R13945 gnd.n6442 gnd.n790 0.152939
R13946 gnd.n6443 gnd.n6442 0.152939
R13947 gnd.n6444 gnd.n6443 0.152939
R13948 gnd.n6444 gnd.n784 0.152939
R13949 gnd.n6452 gnd.n784 0.152939
R13950 gnd.n6453 gnd.n6452 0.152939
R13951 gnd.n6454 gnd.n6453 0.152939
R13952 gnd.n6454 gnd.n778 0.152939
R13953 gnd.n6462 gnd.n778 0.152939
R13954 gnd.n6463 gnd.n6462 0.152939
R13955 gnd.n6464 gnd.n6463 0.152939
R13956 gnd.n6464 gnd.n772 0.152939
R13957 gnd.n6472 gnd.n772 0.152939
R13958 gnd.n6473 gnd.n6472 0.152939
R13959 gnd.n6474 gnd.n6473 0.152939
R13960 gnd.n6474 gnd.n766 0.152939
R13961 gnd.n6482 gnd.n766 0.152939
R13962 gnd.n6483 gnd.n6482 0.152939
R13963 gnd.n6484 gnd.n6483 0.152939
R13964 gnd.n6484 gnd.n760 0.152939
R13965 gnd.n6492 gnd.n760 0.152939
R13966 gnd.n6493 gnd.n6492 0.152939
R13967 gnd.n6494 gnd.n6493 0.152939
R13968 gnd.n6494 gnd.n754 0.152939
R13969 gnd.n6502 gnd.n754 0.152939
R13970 gnd.n6503 gnd.n6502 0.152939
R13971 gnd.n6504 gnd.n6503 0.152939
R13972 gnd.n6504 gnd.n748 0.152939
R13973 gnd.n6512 gnd.n748 0.152939
R13974 gnd.n6513 gnd.n6512 0.152939
R13975 gnd.n6514 gnd.n6513 0.152939
R13976 gnd.n6514 gnd.n742 0.152939
R13977 gnd.n6522 gnd.n742 0.152939
R13978 gnd.n6523 gnd.n6522 0.152939
R13979 gnd.n6524 gnd.n6523 0.152939
R13980 gnd.n6524 gnd.n736 0.152939
R13981 gnd.n6532 gnd.n736 0.152939
R13982 gnd.n6533 gnd.n6532 0.152939
R13983 gnd.n6534 gnd.n6533 0.152939
R13984 gnd.n6534 gnd.n730 0.152939
R13985 gnd.n6542 gnd.n730 0.152939
R13986 gnd.n6543 gnd.n6542 0.152939
R13987 gnd.n6544 gnd.n6543 0.152939
R13988 gnd.n6544 gnd.n724 0.152939
R13989 gnd.n6552 gnd.n724 0.152939
R13990 gnd.n6553 gnd.n6552 0.152939
R13991 gnd.n6554 gnd.n6553 0.152939
R13992 gnd.n6554 gnd.n718 0.152939
R13993 gnd.n6562 gnd.n718 0.152939
R13994 gnd.n6563 gnd.n6562 0.152939
R13995 gnd.n6564 gnd.n6563 0.152939
R13996 gnd.n6564 gnd.n712 0.152939
R13997 gnd.n6572 gnd.n712 0.152939
R13998 gnd.n6573 gnd.n6572 0.152939
R13999 gnd.n6574 gnd.n6573 0.152939
R14000 gnd.n6574 gnd.n706 0.152939
R14001 gnd.n6582 gnd.n706 0.152939
R14002 gnd.n6583 gnd.n6582 0.152939
R14003 gnd.n6584 gnd.n6583 0.152939
R14004 gnd.n6584 gnd.n700 0.152939
R14005 gnd.n6592 gnd.n700 0.152939
R14006 gnd.n6593 gnd.n6592 0.152939
R14007 gnd.n6594 gnd.n6593 0.152939
R14008 gnd.n6594 gnd.n694 0.152939
R14009 gnd.n6602 gnd.n694 0.152939
R14010 gnd.n6603 gnd.n6602 0.152939
R14011 gnd.n6604 gnd.n6603 0.152939
R14012 gnd.n6604 gnd.n688 0.152939
R14013 gnd.n6612 gnd.n688 0.152939
R14014 gnd.n6614 gnd.n6613 0.152939
R14015 gnd.n6614 gnd.n682 0.152939
R14016 gnd.n6622 gnd.n682 0.152939
R14017 gnd.n6623 gnd.n6622 0.152939
R14018 gnd.n6624 gnd.n6623 0.152939
R14019 gnd.n6624 gnd.n676 0.152939
R14020 gnd.n6632 gnd.n676 0.152939
R14021 gnd.n6633 gnd.n6632 0.152939
R14022 gnd.n6634 gnd.n6633 0.152939
R14023 gnd.n6634 gnd.n670 0.152939
R14024 gnd.n6642 gnd.n670 0.152939
R14025 gnd.n6643 gnd.n6642 0.152939
R14026 gnd.n6644 gnd.n6643 0.152939
R14027 gnd.n6644 gnd.n664 0.152939
R14028 gnd.n6652 gnd.n664 0.152939
R14029 gnd.n6653 gnd.n6652 0.152939
R14030 gnd.n6654 gnd.n6653 0.152939
R14031 gnd.n6654 gnd.n658 0.152939
R14032 gnd.n6662 gnd.n658 0.152939
R14033 gnd.n6663 gnd.n6662 0.152939
R14034 gnd.n6664 gnd.n6663 0.152939
R14035 gnd.n6664 gnd.n652 0.152939
R14036 gnd.n6672 gnd.n652 0.152939
R14037 gnd.n6673 gnd.n6672 0.152939
R14038 gnd.n6674 gnd.n6673 0.152939
R14039 gnd.n6674 gnd.n646 0.152939
R14040 gnd.n6682 gnd.n646 0.152939
R14041 gnd.n6683 gnd.n6682 0.152939
R14042 gnd.n6684 gnd.n6683 0.152939
R14043 gnd.n6684 gnd.n640 0.152939
R14044 gnd.n6692 gnd.n640 0.152939
R14045 gnd.n6693 gnd.n6692 0.152939
R14046 gnd.n6694 gnd.n6693 0.152939
R14047 gnd.n6694 gnd.n634 0.152939
R14048 gnd.n6702 gnd.n634 0.152939
R14049 gnd.n6703 gnd.n6702 0.152939
R14050 gnd.n6704 gnd.n6703 0.152939
R14051 gnd.n6704 gnd.n628 0.152939
R14052 gnd.n6712 gnd.n628 0.152939
R14053 gnd.n6713 gnd.n6712 0.152939
R14054 gnd.n6714 gnd.n6713 0.152939
R14055 gnd.n6714 gnd.n622 0.152939
R14056 gnd.n6722 gnd.n622 0.152939
R14057 gnd.n6723 gnd.n6722 0.152939
R14058 gnd.n6724 gnd.n6723 0.152939
R14059 gnd.n6724 gnd.n616 0.152939
R14060 gnd.n6732 gnd.n616 0.152939
R14061 gnd.n6733 gnd.n6732 0.152939
R14062 gnd.n6734 gnd.n6733 0.152939
R14063 gnd.n6734 gnd.n610 0.152939
R14064 gnd.n6742 gnd.n610 0.152939
R14065 gnd.n6743 gnd.n6742 0.152939
R14066 gnd.n6744 gnd.n6743 0.152939
R14067 gnd.n6744 gnd.n604 0.152939
R14068 gnd.n6752 gnd.n604 0.152939
R14069 gnd.n6753 gnd.n6752 0.152939
R14070 gnd.n6754 gnd.n6753 0.152939
R14071 gnd.n6754 gnd.n598 0.152939
R14072 gnd.n6762 gnd.n598 0.152939
R14073 gnd.n6763 gnd.n6762 0.152939
R14074 gnd.n6764 gnd.n6763 0.152939
R14075 gnd.n6764 gnd.n592 0.152939
R14076 gnd.n6772 gnd.n592 0.152939
R14077 gnd.n6773 gnd.n6772 0.152939
R14078 gnd.n6774 gnd.n6773 0.152939
R14079 gnd.n6774 gnd.n586 0.152939
R14080 gnd.n6782 gnd.n586 0.152939
R14081 gnd.n6783 gnd.n6782 0.152939
R14082 gnd.n6784 gnd.n6783 0.152939
R14083 gnd.n6784 gnd.n580 0.152939
R14084 gnd.n6792 gnd.n580 0.152939
R14085 gnd.n6793 gnd.n6792 0.152939
R14086 gnd.n6794 gnd.n6793 0.152939
R14087 gnd.n6794 gnd.n574 0.152939
R14088 gnd.n6802 gnd.n574 0.152939
R14089 gnd.n6803 gnd.n6802 0.152939
R14090 gnd.n6804 gnd.n6803 0.152939
R14091 gnd.n6804 gnd.n568 0.152939
R14092 gnd.n6812 gnd.n568 0.152939
R14093 gnd.n6813 gnd.n6812 0.152939
R14094 gnd.n6814 gnd.n6813 0.152939
R14095 gnd.n6815 gnd.n6814 0.152939
R14096 gnd.n6815 gnd.n562 0.152939
R14097 gnd.n6825 gnd.n562 0.152939
R14098 gnd.n557 gnd.n556 0.152939
R14099 gnd.n560 gnd.n557 0.152939
R14100 gnd.n561 gnd.n560 0.152939
R14101 gnd.n6826 gnd.n561 0.152939
R14102 gnd.n7102 gnd.n7101 0.152939
R14103 gnd.n7103 gnd.n7102 0.152939
R14104 gnd.n7103 gnd.n238 0.152939
R14105 gnd.n7117 gnd.n238 0.152939
R14106 gnd.n7118 gnd.n7117 0.152939
R14107 gnd.n7119 gnd.n7118 0.152939
R14108 gnd.n7119 gnd.n222 0.152939
R14109 gnd.n7133 gnd.n222 0.152939
R14110 gnd.n7134 gnd.n7133 0.152939
R14111 gnd.n7135 gnd.n7134 0.152939
R14112 gnd.n7135 gnd.n208 0.152939
R14113 gnd.n7149 gnd.n208 0.152939
R14114 gnd.n7150 gnd.n7149 0.152939
R14115 gnd.n7151 gnd.n7150 0.152939
R14116 gnd.n7151 gnd.n193 0.152939
R14117 gnd.n7165 gnd.n193 0.152939
R14118 gnd.n7166 gnd.n7165 0.152939
R14119 gnd.n7167 gnd.n7166 0.152939
R14120 gnd.n7168 gnd.n7167 0.152939
R14121 gnd.n7168 gnd.n107 0.152939
R14122 gnd.n7324 gnd.n107 0.152939
R14123 gnd.n7323 gnd.n108 0.152939
R14124 gnd.n110 gnd.n108 0.152939
R14125 gnd.n114 gnd.n110 0.152939
R14126 gnd.n115 gnd.n114 0.152939
R14127 gnd.n116 gnd.n115 0.152939
R14128 gnd.n117 gnd.n116 0.152939
R14129 gnd.n121 gnd.n117 0.152939
R14130 gnd.n122 gnd.n121 0.152939
R14131 gnd.n123 gnd.n122 0.152939
R14132 gnd.n124 gnd.n123 0.152939
R14133 gnd.n128 gnd.n124 0.152939
R14134 gnd.n129 gnd.n128 0.152939
R14135 gnd.n130 gnd.n129 0.152939
R14136 gnd.n131 gnd.n130 0.152939
R14137 gnd.n135 gnd.n131 0.152939
R14138 gnd.n136 gnd.n135 0.152939
R14139 gnd.n137 gnd.n136 0.152939
R14140 gnd.n138 gnd.n137 0.152939
R14141 gnd.n142 gnd.n138 0.152939
R14142 gnd.n143 gnd.n142 0.152939
R14143 gnd.n144 gnd.n143 0.152939
R14144 gnd.n145 gnd.n144 0.152939
R14145 gnd.n149 gnd.n145 0.152939
R14146 gnd.n150 gnd.n149 0.152939
R14147 gnd.n151 gnd.n150 0.152939
R14148 gnd.n152 gnd.n151 0.152939
R14149 gnd.n156 gnd.n152 0.152939
R14150 gnd.n157 gnd.n156 0.152939
R14151 gnd.n158 gnd.n157 0.152939
R14152 gnd.n159 gnd.n158 0.152939
R14153 gnd.n163 gnd.n159 0.152939
R14154 gnd.n164 gnd.n163 0.152939
R14155 gnd.n165 gnd.n164 0.152939
R14156 gnd.n166 gnd.n165 0.152939
R14157 gnd.n170 gnd.n166 0.152939
R14158 gnd.n171 gnd.n170 0.152939
R14159 gnd.n7254 gnd.n171 0.152939
R14160 gnd.n7254 gnd.n7253 0.152939
R14161 gnd.n5465 gnd.n468 0.152939
R14162 gnd.n5466 gnd.n5465 0.152939
R14163 gnd.n5467 gnd.n5466 0.152939
R14164 gnd.n5468 gnd.n5467 0.152939
R14165 gnd.n5469 gnd.n5468 0.152939
R14166 gnd.n5470 gnd.n5469 0.152939
R14167 gnd.n5471 gnd.n5470 0.152939
R14168 gnd.n5472 gnd.n5471 0.152939
R14169 gnd.n5473 gnd.n5472 0.152939
R14170 gnd.n5474 gnd.n5473 0.152939
R14171 gnd.n5511 gnd.n5474 0.152939
R14172 gnd.n5515 gnd.n5511 0.152939
R14173 gnd.n5516 gnd.n5515 0.152939
R14174 gnd.n5517 gnd.n5516 0.152939
R14175 gnd.n5517 gnd.n5509 0.152939
R14176 gnd.n5525 gnd.n5509 0.152939
R14177 gnd.n5526 gnd.n5525 0.152939
R14178 gnd.n5527 gnd.n5526 0.152939
R14179 gnd.n5528 gnd.n5527 0.152939
R14180 gnd.n5529 gnd.n5528 0.152939
R14181 gnd.n5548 gnd.n5529 0.152939
R14182 gnd.n5549 gnd.n5548 0.152939
R14183 gnd.n5551 gnd.n5549 0.152939
R14184 gnd.n5551 gnd.n5550 0.152939
R14185 gnd.n5550 gnd.n496 0.152939
R14186 gnd.n497 gnd.n496 0.152939
R14187 gnd.n499 gnd.n498 0.152939
R14188 gnd.n500 gnd.n499 0.152939
R14189 gnd.n501 gnd.n500 0.152939
R14190 gnd.n502 gnd.n501 0.152939
R14191 gnd.n503 gnd.n502 0.152939
R14192 gnd.n504 gnd.n503 0.152939
R14193 gnd.n505 gnd.n504 0.152939
R14194 gnd.n506 gnd.n505 0.152939
R14195 gnd.n507 gnd.n506 0.152939
R14196 gnd.n508 gnd.n507 0.152939
R14197 gnd.n509 gnd.n508 0.152939
R14198 gnd.n510 gnd.n509 0.152939
R14199 gnd.n511 gnd.n510 0.152939
R14200 gnd.n512 gnd.n511 0.152939
R14201 gnd.n513 gnd.n512 0.152939
R14202 gnd.n514 gnd.n513 0.152939
R14203 gnd.n515 gnd.n514 0.152939
R14204 gnd.n516 gnd.n515 0.152939
R14205 gnd.n517 gnd.n516 0.152939
R14206 gnd.n518 gnd.n517 0.152939
R14207 gnd.n519 gnd.n518 0.152939
R14208 gnd.n520 gnd.n519 0.152939
R14209 gnd.n522 gnd.n520 0.152939
R14210 gnd.n522 gnd.n521 0.152939
R14211 gnd.n521 gnd.n177 0.152939
R14212 gnd.n7252 gnd.n177 0.152939
R14213 gnd.n6970 gnd.n392 0.152939
R14214 gnd.n426 gnd.n392 0.152939
R14215 gnd.n427 gnd.n426 0.152939
R14216 gnd.n428 gnd.n427 0.152939
R14217 gnd.n429 gnd.n428 0.152939
R14218 gnd.n430 gnd.n429 0.152939
R14219 gnd.n431 gnd.n430 0.152939
R14220 gnd.n432 gnd.n431 0.152939
R14221 gnd.n433 gnd.n432 0.152939
R14222 gnd.n434 gnd.n433 0.152939
R14223 gnd.n435 gnd.n434 0.152939
R14224 gnd.n436 gnd.n435 0.152939
R14225 gnd.n437 gnd.n436 0.152939
R14226 gnd.n438 gnd.n437 0.152939
R14227 gnd.n439 gnd.n438 0.152939
R14228 gnd.n446 gnd.n445 0.152939
R14229 gnd.n447 gnd.n446 0.152939
R14230 gnd.n448 gnd.n447 0.152939
R14231 gnd.n449 gnd.n448 0.152939
R14232 gnd.n450 gnd.n449 0.152939
R14233 gnd.n451 gnd.n450 0.152939
R14234 gnd.n452 gnd.n451 0.152939
R14235 gnd.n453 gnd.n452 0.152939
R14236 gnd.n454 gnd.n453 0.152939
R14237 gnd.n455 gnd.n454 0.152939
R14238 gnd.n456 gnd.n455 0.152939
R14239 gnd.n457 gnd.n456 0.152939
R14240 gnd.n458 gnd.n457 0.152939
R14241 gnd.n459 gnd.n458 0.152939
R14242 gnd.n460 gnd.n459 0.152939
R14243 gnd.n461 gnd.n460 0.152939
R14244 gnd.n462 gnd.n461 0.152939
R14245 gnd.n6900 gnd.n462 0.152939
R14246 gnd.n6900 gnd.n6899 0.152939
R14247 gnd.n6899 gnd.n6898 0.152939
R14248 gnd.n6972 gnd.n6971 0.152939
R14249 gnd.n6972 gnd.n375 0.152939
R14250 gnd.n6986 gnd.n375 0.152939
R14251 gnd.n6987 gnd.n6986 0.152939
R14252 gnd.n6988 gnd.n6987 0.152939
R14253 gnd.n6988 gnd.n357 0.152939
R14254 gnd.n7002 gnd.n357 0.152939
R14255 gnd.n7003 gnd.n7002 0.152939
R14256 gnd.n7004 gnd.n7003 0.152939
R14257 gnd.n7004 gnd.n340 0.152939
R14258 gnd.n7018 gnd.n340 0.152939
R14259 gnd.n7019 gnd.n7018 0.152939
R14260 gnd.n7020 gnd.n7019 0.152939
R14261 gnd.n7020 gnd.n322 0.152939
R14262 gnd.n7034 gnd.n322 0.152939
R14263 gnd.n7035 gnd.n7034 0.152939
R14264 gnd.n7036 gnd.n7035 0.152939
R14265 gnd.n7036 gnd.n302 0.152939
R14266 gnd.n7051 gnd.n302 0.152939
R14267 gnd.n7052 gnd.n7051 0.152939
R14268 gnd.n7053 gnd.n7052 0.152939
R14269 gnd.n4437 gnd.n4436 0.152939
R14270 gnd.n4438 gnd.n4437 0.152939
R14271 gnd.n4438 gnd.n2325 0.152939
R14272 gnd.n4444 gnd.n2325 0.152939
R14273 gnd.n4445 gnd.n4444 0.152939
R14274 gnd.n4446 gnd.n4445 0.152939
R14275 gnd.n4447 gnd.n4446 0.152939
R14276 gnd.n4448 gnd.n4447 0.152939
R14277 gnd.n4451 gnd.n4448 0.152939
R14278 gnd.n4452 gnd.n4451 0.152939
R14279 gnd.n4453 gnd.n4452 0.152939
R14280 gnd.n4454 gnd.n4453 0.152939
R14281 gnd.n4456 gnd.n4454 0.152939
R14282 gnd.n4456 gnd.n4455 0.152939
R14283 gnd.n4455 gnd.n2296 0.152939
R14284 gnd.n4528 gnd.n2296 0.152939
R14285 gnd.n4529 gnd.n4528 0.152939
R14286 gnd.n4530 gnd.n4529 0.152939
R14287 gnd.n4530 gnd.n2292 0.152939
R14288 gnd.n4536 gnd.n2292 0.152939
R14289 gnd.n4537 gnd.n4536 0.152939
R14290 gnd.n4538 gnd.n4537 0.152939
R14291 gnd.n4538 gnd.n2288 0.152939
R14292 gnd.n4547 gnd.n2288 0.152939
R14293 gnd.n4548 gnd.n4547 0.152939
R14294 gnd.n4549 gnd.n4548 0.152939
R14295 gnd.n4550 gnd.n4549 0.152939
R14296 gnd.n4550 gnd.n2195 0.152939
R14297 gnd.n4620 gnd.n2195 0.152939
R14298 gnd.n4621 gnd.n4620 0.152939
R14299 gnd.n4622 gnd.n4621 0.152939
R14300 gnd.n4622 gnd.n2181 0.152939
R14301 gnd.n4639 gnd.n2181 0.152939
R14302 gnd.n4640 gnd.n4639 0.152939
R14303 gnd.n4641 gnd.n4640 0.152939
R14304 gnd.n4641 gnd.n2167 0.152939
R14305 gnd.n4659 gnd.n2167 0.152939
R14306 gnd.n4660 gnd.n4659 0.152939
R14307 gnd.n4661 gnd.n4660 0.152939
R14308 gnd.n4662 gnd.n4661 0.152939
R14309 gnd.n4663 gnd.n4662 0.152939
R14310 gnd.n4663 gnd.n1944 0.152939
R14311 gnd.n4711 gnd.n1944 0.152939
R14312 gnd.n4712 gnd.n4711 0.152939
R14313 gnd.n4713 gnd.n4712 0.152939
R14314 gnd.n4714 gnd.n4713 0.152939
R14315 gnd.n4715 gnd.n4714 0.152939
R14316 gnd.n4715 gnd.n1908 0.152939
R14317 gnd.n4794 gnd.n1908 0.152939
R14318 gnd.n4795 gnd.n4794 0.152939
R14319 gnd.n4796 gnd.n4795 0.152939
R14320 gnd.n4796 gnd.n1885 0.152939
R14321 gnd.n4821 gnd.n1885 0.152939
R14322 gnd.n4822 gnd.n4821 0.152939
R14323 gnd.n4823 gnd.n4822 0.152939
R14324 gnd.n4824 gnd.n4823 0.152939
R14325 gnd.n4824 gnd.n1855 0.152939
R14326 gnd.n4862 gnd.n1855 0.152939
R14327 gnd.n4863 gnd.n4862 0.152939
R14328 gnd.n4864 gnd.n4863 0.152939
R14329 gnd.n4864 gnd.n1831 0.152939
R14330 gnd.n4905 gnd.n1831 0.152939
R14331 gnd.n4906 gnd.n4905 0.152939
R14332 gnd.n4907 gnd.n4906 0.152939
R14333 gnd.n4907 gnd.n1815 0.152939
R14334 gnd.n5020 gnd.n1815 0.152939
R14335 gnd.n5021 gnd.n5020 0.152939
R14336 gnd.n5022 gnd.n5021 0.152939
R14337 gnd.n5022 gnd.n1792 0.152939
R14338 gnd.n5047 gnd.n1792 0.152939
R14339 gnd.n5048 gnd.n5047 0.152939
R14340 gnd.n5049 gnd.n5048 0.152939
R14341 gnd.n5050 gnd.n5049 0.152939
R14342 gnd.n5050 gnd.n1763 0.152939
R14343 gnd.n5083 gnd.n1763 0.152939
R14344 gnd.n5084 gnd.n5083 0.152939
R14345 gnd.n5085 gnd.n5084 0.152939
R14346 gnd.n5085 gnd.n1741 0.152939
R14347 gnd.n5113 gnd.n1741 0.152939
R14348 gnd.n5114 gnd.n5113 0.152939
R14349 gnd.n5115 gnd.n5114 0.152939
R14350 gnd.n5115 gnd.n1719 0.152939
R14351 gnd.n5143 gnd.n1719 0.152939
R14352 gnd.n5144 gnd.n5143 0.152939
R14353 gnd.n5145 gnd.n5144 0.152939
R14354 gnd.n5145 gnd.n1697 0.152939
R14355 gnd.n5170 gnd.n1697 0.152939
R14356 gnd.n5171 gnd.n5170 0.152939
R14357 gnd.n5172 gnd.n5171 0.152939
R14358 gnd.n5173 gnd.n5172 0.152939
R14359 gnd.n5173 gnd.n1670 0.152939
R14360 gnd.n5207 gnd.n1670 0.152939
R14361 gnd.n5208 gnd.n5207 0.152939
R14362 gnd.n5209 gnd.n5208 0.152939
R14363 gnd.n5210 gnd.n5209 0.152939
R14364 gnd.n5211 gnd.n5210 0.152939
R14365 gnd.n5213 gnd.n5211 0.152939
R14366 gnd.n5214 gnd.n5213 0.152939
R14367 gnd.n5214 gnd.n1598 0.152939
R14368 gnd.n5408 gnd.n1598 0.152939
R14369 gnd.n5409 gnd.n5408 0.152939
R14370 gnd.n5410 gnd.n5409 0.152939
R14371 gnd.n5410 gnd.n1584 0.152939
R14372 gnd.n5427 gnd.n1584 0.152939
R14373 gnd.n5428 gnd.n5427 0.152939
R14374 gnd.n5429 gnd.n5428 0.152939
R14375 gnd.n5431 gnd.n5429 0.152939
R14376 gnd.n5431 gnd.n5430 0.152939
R14377 gnd.n5430 gnd.n1569 0.152939
R14378 gnd.n5451 gnd.n1569 0.152939
R14379 gnd.n5452 gnd.n5451 0.152939
R14380 gnd.n5453 gnd.n5452 0.152939
R14381 gnd.n5454 gnd.n5453 0.152939
R14382 gnd.n5455 gnd.n5454 0.152939
R14383 gnd.n5458 gnd.n5455 0.152939
R14384 gnd.n5459 gnd.n5458 0.152939
R14385 gnd.n5460 gnd.n5459 0.152939
R14386 gnd.n5461 gnd.n5460 0.152939
R14387 gnd.n5483 gnd.n5461 0.152939
R14388 gnd.n5486 gnd.n5483 0.152939
R14389 gnd.n5487 gnd.n5486 0.152939
R14390 gnd.n5488 gnd.n5487 0.152939
R14391 gnd.n5488 gnd.n5479 0.152939
R14392 gnd.n5494 gnd.n5479 0.152939
R14393 gnd.n5495 gnd.n5494 0.152939
R14394 gnd.n5496 gnd.n5495 0.152939
R14395 gnd.n5497 gnd.n5496 0.152939
R14396 gnd.n5498 gnd.n5497 0.152939
R14397 gnd.n5501 gnd.n5498 0.152939
R14398 gnd.n5502 gnd.n5501 0.152939
R14399 gnd.n5503 gnd.n5502 0.152939
R14400 gnd.n5504 gnd.n5503 0.152939
R14401 gnd.n5537 gnd.n5504 0.152939
R14402 gnd.n5538 gnd.n5537 0.152939
R14403 gnd.n5540 gnd.n5538 0.152939
R14404 gnd.n5541 gnd.n5540 0.152939
R14405 gnd.n5542 gnd.n5541 0.152939
R14406 gnd.n1168 gnd.n1143 0.152939
R14407 gnd.n1169 gnd.n1168 0.152939
R14408 gnd.n1170 gnd.n1169 0.152939
R14409 gnd.n1189 gnd.n1170 0.152939
R14410 gnd.n1190 gnd.n1189 0.152939
R14411 gnd.n1191 gnd.n1190 0.152939
R14412 gnd.n1192 gnd.n1191 0.152939
R14413 gnd.n1209 gnd.n1192 0.152939
R14414 gnd.n1210 gnd.n1209 0.152939
R14415 gnd.n1211 gnd.n1210 0.152939
R14416 gnd.n1212 gnd.n1211 0.152939
R14417 gnd.n1231 gnd.n1212 0.152939
R14418 gnd.n1232 gnd.n1231 0.152939
R14419 gnd.n1233 gnd.n1232 0.152939
R14420 gnd.n1234 gnd.n1233 0.152939
R14421 gnd.n1252 gnd.n1234 0.152939
R14422 gnd.n1253 gnd.n1252 0.152939
R14423 gnd.n1254 gnd.n1253 0.152939
R14424 gnd.n1255 gnd.n1254 0.152939
R14425 gnd.n1273 gnd.n1255 0.152939
R14426 gnd.n5930 gnd.n1273 0.152939
R14427 gnd.n5929 gnd.n1274 0.152939
R14428 gnd.n1279 gnd.n1274 0.152939
R14429 gnd.n1280 gnd.n1279 0.152939
R14430 gnd.n1281 gnd.n1280 0.152939
R14431 gnd.n1282 gnd.n1281 0.152939
R14432 gnd.n1283 gnd.n1282 0.152939
R14433 gnd.n1287 gnd.n1283 0.152939
R14434 gnd.n1288 gnd.n1287 0.152939
R14435 gnd.n1289 gnd.n1288 0.152939
R14436 gnd.n1290 gnd.n1289 0.152939
R14437 gnd.n1294 gnd.n1290 0.152939
R14438 gnd.n1295 gnd.n1294 0.152939
R14439 gnd.n1296 gnd.n1295 0.152939
R14440 gnd.n1297 gnd.n1296 0.152939
R14441 gnd.n1304 gnd.n1297 0.152939
R14442 gnd.n1307 gnd.n1306 0.152939
R14443 gnd.n1308 gnd.n1307 0.152939
R14444 gnd.n1312 gnd.n1308 0.152939
R14445 gnd.n1313 gnd.n1312 0.152939
R14446 gnd.n1314 gnd.n1313 0.152939
R14447 gnd.n1315 gnd.n1314 0.152939
R14448 gnd.n1319 gnd.n1315 0.152939
R14449 gnd.n1320 gnd.n1319 0.152939
R14450 gnd.n1321 gnd.n1320 0.152939
R14451 gnd.n1322 gnd.n1321 0.152939
R14452 gnd.n1326 gnd.n1322 0.152939
R14453 gnd.n1327 gnd.n1326 0.152939
R14454 gnd.n1328 gnd.n1327 0.152939
R14455 gnd.n1329 gnd.n1328 0.152939
R14456 gnd.n1333 gnd.n1329 0.152939
R14457 gnd.n1334 gnd.n1333 0.152939
R14458 gnd.n1335 gnd.n1334 0.152939
R14459 gnd.n1336 gnd.n1335 0.152939
R14460 gnd.n1341 gnd.n1336 0.152939
R14461 gnd.n5861 gnd.n1341 0.152939
R14462 gnd.n4169 gnd.n4124 0.152939
R14463 gnd.n4126 gnd.n4124 0.152939
R14464 gnd.n4127 gnd.n4126 0.152939
R14465 gnd.n4128 gnd.n4127 0.152939
R14466 gnd.n4129 gnd.n4128 0.152939
R14467 gnd.n4130 gnd.n4129 0.152939
R14468 gnd.n4131 gnd.n4130 0.152939
R14469 gnd.n4132 gnd.n4131 0.152939
R14470 gnd.n4133 gnd.n4132 0.152939
R14471 gnd.n4134 gnd.n4133 0.152939
R14472 gnd.n4135 gnd.n4134 0.152939
R14473 gnd.n4136 gnd.n4135 0.152939
R14474 gnd.n4137 gnd.n4136 0.152939
R14475 gnd.n4138 gnd.n4137 0.152939
R14476 gnd.n4139 gnd.n4138 0.152939
R14477 gnd.n4140 gnd.n4139 0.152939
R14478 gnd.n4142 gnd.n4140 0.152939
R14479 gnd.n4142 gnd.n4141 0.152939
R14480 gnd.n4141 gnd.n2392 0.152939
R14481 gnd.n2393 gnd.n2392 0.152939
R14482 gnd.n2394 gnd.n2393 0.152939
R14483 gnd.n4302 gnd.n2394 0.152939
R14484 gnd.n4303 gnd.n4302 0.152939
R14485 gnd.n4304 gnd.n4303 0.152939
R14486 gnd.n4305 gnd.n4304 0.152939
R14487 gnd.n4306 gnd.n4305 0.152939
R14488 gnd.n4210 gnd.n4098 0.152939
R14489 gnd.n4101 gnd.n4098 0.152939
R14490 gnd.n4102 gnd.n4101 0.152939
R14491 gnd.n4103 gnd.n4102 0.152939
R14492 gnd.n4104 gnd.n4103 0.152939
R14493 gnd.n4107 gnd.n4104 0.152939
R14494 gnd.n4108 gnd.n4107 0.152939
R14495 gnd.n4109 gnd.n4108 0.152939
R14496 gnd.n4110 gnd.n4109 0.152939
R14497 gnd.n4113 gnd.n4110 0.152939
R14498 gnd.n4114 gnd.n4113 0.152939
R14499 gnd.n4115 gnd.n4114 0.152939
R14500 gnd.n4116 gnd.n4115 0.152939
R14501 gnd.n4119 gnd.n4116 0.152939
R14502 gnd.n4120 gnd.n4119 0.152939
R14503 gnd.n4176 gnd.n4120 0.152939
R14504 gnd.n4176 gnd.n4175 0.152939
R14505 gnd.n4175 gnd.n4174 0.152939
R14506 gnd.n4211 gnd.n2448 0.152939
R14507 gnd.n4225 gnd.n2448 0.152939
R14508 gnd.n4226 gnd.n4225 0.152939
R14509 gnd.n4227 gnd.n4226 0.152939
R14510 gnd.n4227 gnd.n2432 0.152939
R14511 gnd.n4241 gnd.n2432 0.152939
R14512 gnd.n4242 gnd.n4241 0.152939
R14513 gnd.n4243 gnd.n4242 0.152939
R14514 gnd.n4243 gnd.n2415 0.152939
R14515 gnd.n4257 gnd.n2415 0.152939
R14516 gnd.n4258 gnd.n4257 0.152939
R14517 gnd.n4259 gnd.n4258 0.152939
R14518 gnd.n4260 gnd.n4259 0.152939
R14519 gnd.n4261 gnd.n4260 0.152939
R14520 gnd.n4262 gnd.n4261 0.152939
R14521 gnd.n4264 gnd.n4262 0.152939
R14522 gnd.n4264 gnd.n4263 0.152939
R14523 gnd.n4263 gnd.n1129 0.152939
R14524 gnd.n1130 gnd.n1129 0.152939
R14525 gnd.n1131 gnd.n1130 0.152939
R14526 gnd.n2377 gnd.n1131 0.152939
R14527 gnd.n4347 gnd.n2377 0.152939
R14528 gnd.n4348 gnd.n4347 0.152939
R14529 gnd.n4349 gnd.n4348 0.152939
R14530 gnd.n4350 gnd.n4349 0.152939
R14531 gnd.n4350 gnd.n2355 0.152939
R14532 gnd.n4381 gnd.n4380 0.152939
R14533 gnd.n4383 gnd.n4381 0.152939
R14534 gnd.n4383 gnd.n4382 0.152939
R14535 gnd.n4382 gnd.n1159 0.152939
R14536 gnd.n1160 gnd.n1159 0.152939
R14537 gnd.n1161 gnd.n1160 0.152939
R14538 gnd.n1178 gnd.n1161 0.152939
R14539 gnd.n1179 gnd.n1178 0.152939
R14540 gnd.n1180 gnd.n1179 0.152939
R14541 gnd.n1181 gnd.n1180 0.152939
R14542 gnd.n1199 gnd.n1181 0.152939
R14543 gnd.n1200 gnd.n1199 0.152939
R14544 gnd.n1201 gnd.n1200 0.152939
R14545 gnd.n1202 gnd.n1201 0.152939
R14546 gnd.n1220 gnd.n1202 0.152939
R14547 gnd.n1221 gnd.n1220 0.152939
R14548 gnd.n1222 gnd.n1221 0.152939
R14549 gnd.n1223 gnd.n1222 0.152939
R14550 gnd.n1241 gnd.n1223 0.152939
R14551 gnd.n1242 gnd.n1241 0.152939
R14552 gnd.n1243 gnd.n1242 0.152939
R14553 gnd.n1244 gnd.n1243 0.152939
R14554 gnd.n1263 gnd.n1244 0.152939
R14555 gnd.n1264 gnd.n1263 0.152939
R14556 gnd.n1265 gnd.n1264 0.152939
R14557 gnd.n1266 gnd.n1265 0.152939
R14558 gnd.n4093 gnd.n4064 0.152939
R14559 gnd.n4093 gnd.n4092 0.152939
R14560 gnd.n4092 gnd.n4091 0.152939
R14561 gnd.n4091 gnd.n4065 0.152939
R14562 gnd.n4066 gnd.n4065 0.152939
R14563 gnd.n4067 gnd.n4066 0.152939
R14564 gnd.n4068 gnd.n4067 0.152939
R14565 gnd.n4069 gnd.n4068 0.152939
R14566 gnd.n4070 gnd.n4069 0.152939
R14567 gnd.n4071 gnd.n4070 0.152939
R14568 gnd.n4072 gnd.n4071 0.152939
R14569 gnd.n4073 gnd.n4072 0.152939
R14570 gnd.n4074 gnd.n4073 0.152939
R14571 gnd.n4074 gnd.n2399 0.152939
R14572 gnd.n4285 gnd.n2399 0.152939
R14573 gnd.n4286 gnd.n4285 0.152939
R14574 gnd.n4287 gnd.n4286 0.152939
R14575 gnd.n4287 gnd.n2397 0.152939
R14576 gnd.n4292 gnd.n2397 0.152939
R14577 gnd.n4293 gnd.n4292 0.152939
R14578 gnd.n4294 gnd.n4293 0.152939
R14579 gnd.n4295 gnd.n4294 0.152939
R14580 gnd.n4296 gnd.n4295 0.152939
R14581 gnd.n4297 gnd.n4296 0.152939
R14582 gnd.n4298 gnd.n4297 0.152939
R14583 gnd.n4298 gnd.n2356 0.152939
R14584 gnd.n4377 gnd.n2357 0.152939
R14585 gnd.n2357 gnd.n2346 0.152939
R14586 gnd.n4396 gnd.n2346 0.152939
R14587 gnd.n4397 gnd.n4396 0.152939
R14588 gnd.n4398 gnd.n4397 0.152939
R14589 gnd.n4398 gnd.n2344 0.152939
R14590 gnd.n4407 gnd.n2344 0.152939
R14591 gnd.n4408 gnd.n4407 0.152939
R14592 gnd.n4409 gnd.n4408 0.152939
R14593 gnd.n4410 gnd.n4409 0.152939
R14594 gnd.n4411 gnd.n4410 0.152939
R14595 gnd.n4411 gnd.n2316 0.152939
R14596 gnd.n4481 gnd.n2316 0.152939
R14597 gnd.n4482 gnd.n4481 0.152939
R14598 gnd.n4483 gnd.n4482 0.152939
R14599 gnd.n4483 gnd.n2309 0.152939
R14600 gnd.n4497 gnd.n2309 0.152939
R14601 gnd.n4498 gnd.n4497 0.152939
R14602 gnd.n4499 gnd.n4498 0.152939
R14603 gnd.n4499 gnd.n2307 0.152939
R14604 gnd.n4505 gnd.n2307 0.152939
R14605 gnd.n4506 gnd.n4505 0.152939
R14606 gnd.n4508 gnd.n4506 0.152939
R14607 gnd.n4508 gnd.n4507 0.152939
R14608 gnd.n4507 gnd.n1342 0.152939
R14609 gnd.n5860 gnd.n1342 0.152939
R14610 gnd.n3971 gnd.n2455 0.152939
R14611 gnd.n3972 gnd.n3971 0.152939
R14612 gnd.n3973 gnd.n3972 0.152939
R14613 gnd.n3973 gnd.n3963 0.152939
R14614 gnd.n3981 gnd.n3963 0.152939
R14615 gnd.n3982 gnd.n3981 0.152939
R14616 gnd.n3983 gnd.n3982 0.152939
R14617 gnd.n3983 gnd.n3959 0.152939
R14618 gnd.n3991 gnd.n3959 0.152939
R14619 gnd.n3992 gnd.n3991 0.152939
R14620 gnd.n3993 gnd.n3992 0.152939
R14621 gnd.n3993 gnd.n3955 0.152939
R14622 gnd.n4001 gnd.n3955 0.152939
R14623 gnd.n4002 gnd.n4001 0.152939
R14624 gnd.n4003 gnd.n4002 0.152939
R14625 gnd.n4003 gnd.n3948 0.152939
R14626 gnd.n4011 gnd.n3948 0.152939
R14627 gnd.n4012 gnd.n4011 0.152939
R14628 gnd.n4013 gnd.n4012 0.152939
R14629 gnd.n4013 gnd.n3944 0.152939
R14630 gnd.n4021 gnd.n3944 0.152939
R14631 gnd.n4022 gnd.n4021 0.152939
R14632 gnd.n4023 gnd.n4022 0.152939
R14633 gnd.n4023 gnd.n3940 0.152939
R14634 gnd.n4031 gnd.n3940 0.152939
R14635 gnd.n4032 gnd.n4031 0.152939
R14636 gnd.n4033 gnd.n4032 0.152939
R14637 gnd.n4033 gnd.n3936 0.152939
R14638 gnd.n4041 gnd.n3936 0.152939
R14639 gnd.n4042 gnd.n4041 0.152939
R14640 gnd.n4043 gnd.n4042 0.152939
R14641 gnd.n4043 gnd.n3932 0.152939
R14642 gnd.n4051 gnd.n3932 0.152939
R14643 gnd.n4052 gnd.n4051 0.152939
R14644 gnd.n4054 gnd.n4052 0.152939
R14645 gnd.n4054 gnd.n4053 0.152939
R14646 gnd.n4053 gnd.n3925 0.152939
R14647 gnd.n4063 gnd.n3925 0.152939
R14648 gnd.n4218 gnd.n4217 0.152939
R14649 gnd.n4219 gnd.n4218 0.152939
R14650 gnd.n4219 gnd.n2440 0.152939
R14651 gnd.n4233 gnd.n2440 0.152939
R14652 gnd.n4234 gnd.n4233 0.152939
R14653 gnd.n4235 gnd.n4234 0.152939
R14654 gnd.n4235 gnd.n2423 0.152939
R14655 gnd.n4249 gnd.n2423 0.152939
R14656 gnd.n4250 gnd.n4249 0.152939
R14657 gnd.n4251 gnd.n4250 0.152939
R14658 gnd.n4251 gnd.n2407 0.152939
R14659 gnd.n4275 gnd.n2407 0.152939
R14660 gnd.n4276 gnd.n4275 0.152939
R14661 gnd.n4278 gnd.n4276 0.152939
R14662 gnd.n4278 gnd.n4277 0.152939
R14663 gnd.n4277 gnd.n1117 0.152939
R14664 gnd.n1118 gnd.n1117 0.152939
R14665 gnd.n1119 gnd.n1118 0.152939
R14666 gnd.n1138 gnd.n1119 0.152939
R14667 gnd.n1139 gnd.n1138 0.152939
R14668 gnd.n1140 gnd.n1139 0.152939
R14669 gnd.n2385 gnd.n2384 0.152939
R14670 gnd.n4334 gnd.n2384 0.152939
R14671 gnd.n4335 gnd.n4334 0.152939
R14672 gnd.n4336 gnd.n4335 0.152939
R14673 gnd.n6192 gnd.n940 0.152939
R14674 gnd.n945 gnd.n940 0.152939
R14675 gnd.n946 gnd.n945 0.152939
R14676 gnd.n947 gnd.n946 0.152939
R14677 gnd.n952 gnd.n947 0.152939
R14678 gnd.n953 gnd.n952 0.152939
R14679 gnd.n954 gnd.n953 0.152939
R14680 gnd.n955 gnd.n954 0.152939
R14681 gnd.n960 gnd.n955 0.152939
R14682 gnd.n961 gnd.n960 0.152939
R14683 gnd.n962 gnd.n961 0.152939
R14684 gnd.n963 gnd.n962 0.152939
R14685 gnd.n968 gnd.n963 0.152939
R14686 gnd.n969 gnd.n968 0.152939
R14687 gnd.n970 gnd.n969 0.152939
R14688 gnd.n971 gnd.n970 0.152939
R14689 gnd.n976 gnd.n971 0.152939
R14690 gnd.n977 gnd.n976 0.152939
R14691 gnd.n978 gnd.n977 0.152939
R14692 gnd.n979 gnd.n978 0.152939
R14693 gnd.n984 gnd.n979 0.152939
R14694 gnd.n985 gnd.n984 0.152939
R14695 gnd.n986 gnd.n985 0.152939
R14696 gnd.n987 gnd.n986 0.152939
R14697 gnd.n992 gnd.n987 0.152939
R14698 gnd.n993 gnd.n992 0.152939
R14699 gnd.n994 gnd.n993 0.152939
R14700 gnd.n995 gnd.n994 0.152939
R14701 gnd.n1000 gnd.n995 0.152939
R14702 gnd.n1001 gnd.n1000 0.152939
R14703 gnd.n1002 gnd.n1001 0.152939
R14704 gnd.n1003 gnd.n1002 0.152939
R14705 gnd.n1008 gnd.n1003 0.152939
R14706 gnd.n1009 gnd.n1008 0.152939
R14707 gnd.n1010 gnd.n1009 0.152939
R14708 gnd.n1011 gnd.n1010 0.152939
R14709 gnd.n1016 gnd.n1011 0.152939
R14710 gnd.n1017 gnd.n1016 0.152939
R14711 gnd.n1018 gnd.n1017 0.152939
R14712 gnd.n1019 gnd.n1018 0.152939
R14713 gnd.n1024 gnd.n1019 0.152939
R14714 gnd.n1025 gnd.n1024 0.152939
R14715 gnd.n1026 gnd.n1025 0.152939
R14716 gnd.n1027 gnd.n1026 0.152939
R14717 gnd.n1032 gnd.n1027 0.152939
R14718 gnd.n1033 gnd.n1032 0.152939
R14719 gnd.n1034 gnd.n1033 0.152939
R14720 gnd.n1035 gnd.n1034 0.152939
R14721 gnd.n1040 gnd.n1035 0.152939
R14722 gnd.n1041 gnd.n1040 0.152939
R14723 gnd.n1042 gnd.n1041 0.152939
R14724 gnd.n1043 gnd.n1042 0.152939
R14725 gnd.n1048 gnd.n1043 0.152939
R14726 gnd.n1049 gnd.n1048 0.152939
R14727 gnd.n1050 gnd.n1049 0.152939
R14728 gnd.n1051 gnd.n1050 0.152939
R14729 gnd.n1056 gnd.n1051 0.152939
R14730 gnd.n1057 gnd.n1056 0.152939
R14731 gnd.n1058 gnd.n1057 0.152939
R14732 gnd.n1059 gnd.n1058 0.152939
R14733 gnd.n1064 gnd.n1059 0.152939
R14734 gnd.n1065 gnd.n1064 0.152939
R14735 gnd.n1066 gnd.n1065 0.152939
R14736 gnd.n1067 gnd.n1066 0.152939
R14737 gnd.n1072 gnd.n1067 0.152939
R14738 gnd.n1073 gnd.n1072 0.152939
R14739 gnd.n1074 gnd.n1073 0.152939
R14740 gnd.n1075 gnd.n1074 0.152939
R14741 gnd.n1080 gnd.n1075 0.152939
R14742 gnd.n1081 gnd.n1080 0.152939
R14743 gnd.n1082 gnd.n1081 0.152939
R14744 gnd.n1083 gnd.n1082 0.152939
R14745 gnd.n1088 gnd.n1083 0.152939
R14746 gnd.n1089 gnd.n1088 0.152939
R14747 gnd.n1090 gnd.n1089 0.152939
R14748 gnd.n1091 gnd.n1090 0.152939
R14749 gnd.n1096 gnd.n1091 0.152939
R14750 gnd.n1097 gnd.n1096 0.152939
R14751 gnd.n1098 gnd.n1097 0.152939
R14752 gnd.n1099 gnd.n1098 0.152939
R14753 gnd.n1104 gnd.n1099 0.152939
R14754 gnd.n1105 gnd.n1104 0.152939
R14755 gnd.n1106 gnd.n1105 0.152939
R14756 gnd.n1107 gnd.n1106 0.152939
R14757 gnd.n5647 gnd.n5646 0.152939
R14758 gnd.n5646 gnd.n5645 0.152939
R14759 gnd.n5645 gnd.n1533 0.152939
R14760 gnd.n5641 gnd.n1533 0.152939
R14761 gnd.n5641 gnd.n5640 0.152939
R14762 gnd.n5640 gnd.n5639 0.152939
R14763 gnd.n5639 gnd.n1538 0.152939
R14764 gnd.n5635 gnd.n1538 0.152939
R14765 gnd.n5635 gnd.n5634 0.152939
R14766 gnd.n5833 gnd.n1366 0.152939
R14767 gnd.n5829 gnd.n1366 0.152939
R14768 gnd.n5829 gnd.n5828 0.152939
R14769 gnd.n5828 gnd.n5827 0.152939
R14770 gnd.n5827 gnd.n1371 0.152939
R14771 gnd.n5823 gnd.n1371 0.152939
R14772 gnd.n5823 gnd.n5822 0.152939
R14773 gnd.n5822 gnd.n5821 0.152939
R14774 gnd.n5821 gnd.n1376 0.152939
R14775 gnd.n5817 gnd.n1376 0.152939
R14776 gnd.n5817 gnd.n5816 0.152939
R14777 gnd.n5816 gnd.n5815 0.152939
R14778 gnd.n5815 gnd.n1381 0.152939
R14779 gnd.n5811 gnd.n1381 0.152939
R14780 gnd.n5811 gnd.n5810 0.152939
R14781 gnd.n5810 gnd.n5809 0.152939
R14782 gnd.n5809 gnd.n1386 0.152939
R14783 gnd.n5805 gnd.n1386 0.152939
R14784 gnd.n5805 gnd.n5804 0.152939
R14785 gnd.n5804 gnd.n5803 0.152939
R14786 gnd.n5803 gnd.n1391 0.152939
R14787 gnd.n5799 gnd.n1391 0.152939
R14788 gnd.n5799 gnd.n5798 0.152939
R14789 gnd.n5798 gnd.n5797 0.152939
R14790 gnd.n5797 gnd.n1396 0.152939
R14791 gnd.n5793 gnd.n1396 0.152939
R14792 gnd.n5793 gnd.n5792 0.152939
R14793 gnd.n5792 gnd.n5791 0.152939
R14794 gnd.n5791 gnd.n1401 0.152939
R14795 gnd.n5787 gnd.n1401 0.152939
R14796 gnd.n5787 gnd.n5786 0.152939
R14797 gnd.n5786 gnd.n5785 0.152939
R14798 gnd.n5785 gnd.n1406 0.152939
R14799 gnd.n5781 gnd.n1406 0.152939
R14800 gnd.n5781 gnd.n5780 0.152939
R14801 gnd.n5780 gnd.n5779 0.152939
R14802 gnd.n5779 gnd.n1411 0.152939
R14803 gnd.n5775 gnd.n1411 0.152939
R14804 gnd.n5775 gnd.n5774 0.152939
R14805 gnd.n5774 gnd.n5773 0.152939
R14806 gnd.n5773 gnd.n1416 0.152939
R14807 gnd.n5769 gnd.n1416 0.152939
R14808 gnd.n5769 gnd.n5768 0.152939
R14809 gnd.n5768 gnd.n5767 0.152939
R14810 gnd.n5767 gnd.n1421 0.152939
R14811 gnd.n5763 gnd.n1421 0.152939
R14812 gnd.n5763 gnd.n5762 0.152939
R14813 gnd.n5762 gnd.n5761 0.152939
R14814 gnd.n5761 gnd.n1426 0.152939
R14815 gnd.n5757 gnd.n1426 0.152939
R14816 gnd.n5757 gnd.n5756 0.152939
R14817 gnd.n5756 gnd.n5755 0.152939
R14818 gnd.n5755 gnd.n1431 0.152939
R14819 gnd.n5751 gnd.n1431 0.152939
R14820 gnd.n5751 gnd.n5750 0.152939
R14821 gnd.n5750 gnd.n5749 0.152939
R14822 gnd.n5749 gnd.n1436 0.152939
R14823 gnd.n5745 gnd.n1436 0.152939
R14824 gnd.n5745 gnd.n5744 0.152939
R14825 gnd.n5744 gnd.n5743 0.152939
R14826 gnd.n5743 gnd.n1441 0.152939
R14827 gnd.n5739 gnd.n1441 0.152939
R14828 gnd.n5739 gnd.n5738 0.152939
R14829 gnd.n5738 gnd.n5737 0.152939
R14830 gnd.n5737 gnd.n1446 0.152939
R14831 gnd.n5733 gnd.n1446 0.152939
R14832 gnd.n5733 gnd.n5732 0.152939
R14833 gnd.n5732 gnd.n5731 0.152939
R14834 gnd.n5731 gnd.n1451 0.152939
R14835 gnd.n5727 gnd.n1451 0.152939
R14836 gnd.n5727 gnd.n5726 0.152939
R14837 gnd.n5726 gnd.n5725 0.152939
R14838 gnd.n5725 gnd.n1456 0.152939
R14839 gnd.n5721 gnd.n1456 0.152939
R14840 gnd.n5721 gnd.n5720 0.152939
R14841 gnd.n5720 gnd.n5719 0.152939
R14842 gnd.n5719 gnd.n1461 0.152939
R14843 gnd.n5715 gnd.n1461 0.152939
R14844 gnd.n5715 gnd.n5714 0.152939
R14845 gnd.n5714 gnd.n5713 0.152939
R14846 gnd.n5713 gnd.n1466 0.152939
R14847 gnd.n1469 gnd.n1466 0.152939
R14848 gnd.n5846 gnd.n1347 0.152939
R14849 gnd.n5846 gnd.n5845 0.152939
R14850 gnd.n5845 gnd.n5844 0.152939
R14851 gnd.n5844 gnd.n1354 0.152939
R14852 gnd.n5840 gnd.n1354 0.152939
R14853 gnd.n5840 gnd.n5839 0.152939
R14854 gnd.n5839 gnd.n1361 0.152939
R14855 gnd.n5835 gnd.n1361 0.152939
R14856 gnd.n5835 gnd.n5834 0.152939
R14857 gnd.n4310 gnd.n4309 0.152939
R14858 gnd.n4309 gnd.n2338 0.152939
R14859 gnd.n4427 gnd.n2338 0.152939
R14860 gnd.n4427 gnd.n4426 0.152939
R14861 gnd.n4426 gnd.n4425 0.152939
R14862 gnd.n4425 gnd.n2339 0.152939
R14863 gnd.n4421 gnd.n2339 0.152939
R14864 gnd.n4421 gnd.n4420 0.152939
R14865 gnd.n4420 gnd.n4419 0.152939
R14866 gnd.n4419 gnd.n2319 0.152939
R14867 gnd.n4473 gnd.n2319 0.152939
R14868 gnd.n4474 gnd.n4473 0.152939
R14869 gnd.n4475 gnd.n4474 0.152939
R14870 gnd.n4475 gnd.n2312 0.152939
R14871 gnd.n4489 gnd.n2312 0.152939
R14872 gnd.n4490 gnd.n4489 0.152939
R14873 gnd.n4491 gnd.n4490 0.152939
R14874 gnd.n4491 gnd.n2303 0.152939
R14875 gnd.n4519 gnd.n2303 0.152939
R14876 gnd.n4519 gnd.n4518 0.152939
R14877 gnd.n4518 gnd.n4517 0.152939
R14878 gnd.n4517 gnd.n2304 0.152939
R14879 gnd.n4513 gnd.n2304 0.152939
R14880 gnd.n4513 gnd.n1346 0.152939
R14881 gnd.n5853 gnd.n1346 0.152939
R14882 gnd.n5853 gnd.n5852 0.152939
R14883 gnd.n4612 gnd.n4611 0.152939
R14884 gnd.n4612 gnd.n2187 0.152939
R14885 gnd.n4629 gnd.n2187 0.152939
R14886 gnd.n4630 gnd.n4629 0.152939
R14887 gnd.n4631 gnd.n4630 0.152939
R14888 gnd.n4631 gnd.n2173 0.152939
R14889 gnd.n4648 gnd.n2173 0.152939
R14890 gnd.n4649 gnd.n4648 0.152939
R14891 gnd.n4650 gnd.n4649 0.152939
R14892 gnd.n4650 gnd.n1987 0.152939
R14893 gnd.n4674 gnd.n1987 0.152939
R14894 gnd.n4675 gnd.n4674 0.152939
R14895 gnd.n4685 gnd.n4675 0.152939
R14896 gnd.n4685 gnd.n4684 0.152939
R14897 gnd.n4684 gnd.n4683 0.152939
R14898 gnd.n4683 gnd.n4676 0.152939
R14899 gnd.n4676 gnd.n1926 0.152939
R14900 gnd.n4734 gnd.n1926 0.152939
R14901 gnd.n4735 gnd.n4734 0.152939
R14902 gnd.n4737 gnd.n4735 0.152939
R14903 gnd.n4737 gnd.n4736 0.152939
R14904 gnd.n4736 gnd.n1900 0.152939
R14905 gnd.n4803 gnd.n1900 0.152939
R14906 gnd.n4804 gnd.n4803 0.152939
R14907 gnd.n4806 gnd.n4804 0.152939
R14908 gnd.n4806 gnd.n4805 0.152939
R14909 gnd.n4805 gnd.n1870 0.152939
R14910 gnd.n4839 gnd.n1870 0.152939
R14911 gnd.n4840 gnd.n4839 0.152939
R14912 gnd.n4841 gnd.n4840 0.152939
R14913 gnd.n4841 gnd.n1847 0.152939
R14914 gnd.n4871 gnd.n1847 0.152939
R14915 gnd.n4872 gnd.n4871 0.152939
R14916 gnd.n4883 gnd.n4872 0.152939
R14917 gnd.n4883 gnd.n4882 0.152939
R14918 gnd.n4882 gnd.n4881 0.152939
R14919 gnd.n4881 gnd.n4873 0.152939
R14920 gnd.n4877 gnd.n4873 0.152939
R14921 gnd.n4877 gnd.n1808 0.152939
R14922 gnd.n5029 gnd.n1808 0.152939
R14923 gnd.n5030 gnd.n5029 0.152939
R14924 gnd.n5032 gnd.n5030 0.152939
R14925 gnd.n5032 gnd.n5031 0.152939
R14926 gnd.n5031 gnd.n1778 0.152939
R14927 gnd.n5065 gnd.n1778 0.152939
R14928 gnd.n5066 gnd.n5065 0.152939
R14929 gnd.n5067 gnd.n5066 0.152939
R14930 gnd.n5067 gnd.n1756 0.152939
R14931 gnd.n5092 gnd.n1756 0.152939
R14932 gnd.n5093 gnd.n5092 0.152939
R14933 gnd.n5094 gnd.n5093 0.152939
R14934 gnd.n5094 gnd.n1734 0.152939
R14935 gnd.n5122 gnd.n1734 0.152939
R14936 gnd.n5123 gnd.n5122 0.152939
R14937 gnd.n5124 gnd.n5123 0.152939
R14938 gnd.n5124 gnd.n1713 0.152939
R14939 gnd.n5152 gnd.n1713 0.152939
R14940 gnd.n5153 gnd.n5152 0.152939
R14941 gnd.n5155 gnd.n5153 0.152939
R14942 gnd.n5155 gnd.n5154 0.152939
R14943 gnd.n5154 gnd.n1684 0.152939
R14944 gnd.n5188 gnd.n1684 0.152939
R14945 gnd.n5189 gnd.n5188 0.152939
R14946 gnd.n5190 gnd.n5189 0.152939
R14947 gnd.n5190 gnd.n1660 0.152939
R14948 gnd.n5227 gnd.n1660 0.152939
R14949 gnd.n5228 gnd.n5227 0.152939
R14950 gnd.n5229 gnd.n5228 0.152939
R14951 gnd.n5229 gnd.n1604 0.152939
R14952 gnd.n5398 gnd.n1604 0.152939
R14953 gnd.n5399 gnd.n5398 0.152939
R14954 gnd.n5400 gnd.n5399 0.152939
R14955 gnd.n5400 gnd.n1589 0.152939
R14956 gnd.n5417 gnd.n1589 0.152939
R14957 gnd.n5418 gnd.n5417 0.152939
R14958 gnd.n5419 gnd.n5418 0.152939
R14959 gnd.n5419 gnd.n1576 0.152939
R14960 gnd.n5439 gnd.n1576 0.152939
R14961 gnd.n5440 gnd.n5439 0.152939
R14962 gnd.n5441 gnd.n5440 0.152939
R14963 gnd.n5441 gnd.n1476 0.152939
R14964 gnd.n5705 gnd.n1476 0.152939
R14965 gnd.n6978 gnd.n384 0.152939
R14966 gnd.n6979 gnd.n6978 0.152939
R14967 gnd.n6980 gnd.n6979 0.152939
R14968 gnd.n6980 gnd.n366 0.152939
R14969 gnd.n6994 gnd.n366 0.152939
R14970 gnd.n6995 gnd.n6994 0.152939
R14971 gnd.n6996 gnd.n6995 0.152939
R14972 gnd.n6996 gnd.n349 0.152939
R14973 gnd.n7010 gnd.n349 0.152939
R14974 gnd.n7011 gnd.n7010 0.152939
R14975 gnd.n7012 gnd.n7011 0.152939
R14976 gnd.n7012 gnd.n331 0.152939
R14977 gnd.n7026 gnd.n331 0.152939
R14978 gnd.n7027 gnd.n7026 0.152939
R14979 gnd.n7028 gnd.n7027 0.152939
R14980 gnd.n7028 gnd.n314 0.152939
R14981 gnd.n7042 gnd.n314 0.152939
R14982 gnd.n7043 gnd.n7042 0.152939
R14983 gnd.n7045 gnd.n7043 0.152939
R14984 gnd.n7045 gnd.n7044 0.152939
R14985 gnd.n7044 gnd.n294 0.152939
R14986 gnd.n7061 gnd.n294 0.152939
R14987 gnd.n7062 gnd.n7061 0.152939
R14988 gnd.n7063 gnd.n7062 0.152939
R14989 gnd.n7063 gnd.n278 0.152939
R14990 gnd.n7077 gnd.n278 0.152939
R14991 gnd.n7080 gnd.n7079 0.152939
R14992 gnd.n7080 gnd.n263 0.152939
R14993 gnd.n7093 gnd.n263 0.152939
R14994 gnd.n7094 gnd.n7093 0.152939
R14995 gnd.n7095 gnd.n7094 0.152939
R14996 gnd.n7095 gnd.n246 0.152939
R14997 gnd.n7109 gnd.n246 0.152939
R14998 gnd.n7110 gnd.n7109 0.152939
R14999 gnd.n7111 gnd.n7110 0.152939
R15000 gnd.n7111 gnd.n230 0.152939
R15001 gnd.n7125 gnd.n230 0.152939
R15002 gnd.n7126 gnd.n7125 0.152939
R15003 gnd.n7127 gnd.n7126 0.152939
R15004 gnd.n7127 gnd.n214 0.152939
R15005 gnd.n7141 gnd.n214 0.152939
R15006 gnd.n7142 gnd.n7141 0.152939
R15007 gnd.n7143 gnd.n7142 0.152939
R15008 gnd.n7143 gnd.n200 0.152939
R15009 gnd.n7157 gnd.n200 0.152939
R15010 gnd.n7158 gnd.n7157 0.152939
R15011 gnd.n7159 gnd.n7158 0.152939
R15012 gnd.n7159 gnd.n183 0.152939
R15013 gnd.n7175 gnd.n183 0.152939
R15014 gnd.n7176 gnd.n7175 0.152939
R15015 gnd.n7245 gnd.n7176 0.152939
R15016 gnd.n7245 gnd.n7244 0.152939
R15017 gnd.n7243 gnd.n7177 0.152939
R15018 gnd.n7239 gnd.n7177 0.152939
R15019 gnd.n7239 gnd.n7238 0.152939
R15020 gnd.n7238 gnd.n7237 0.152939
R15021 gnd.n7237 gnd.n7183 0.152939
R15022 gnd.n7233 gnd.n7183 0.152939
R15023 gnd.n7233 gnd.n7232 0.152939
R15024 gnd.n7232 gnd.n7231 0.152939
R15025 gnd.n7231 gnd.n7191 0.152939
R15026 gnd.n7227 gnd.n7191 0.152939
R15027 gnd.n7227 gnd.n7226 0.152939
R15028 gnd.n7226 gnd.n7225 0.152939
R15029 gnd.n7225 gnd.n7199 0.152939
R15030 gnd.n7221 gnd.n7199 0.152939
R15031 gnd.n7221 gnd.n7220 0.152939
R15032 gnd.n7220 gnd.n7219 0.152939
R15033 gnd.n7219 gnd.n7207 0.152939
R15034 gnd.n7215 gnd.n7207 0.152939
R15035 gnd.n6891 gnd.n6890 0.152939
R15036 gnd.n6890 gnd.n6889 0.152939
R15037 gnd.n6889 gnd.n473 0.152939
R15038 gnd.n6885 gnd.n473 0.152939
R15039 gnd.n6885 gnd.n6884 0.152939
R15040 gnd.n6884 gnd.n6883 0.152939
R15041 gnd.n6883 gnd.n477 0.152939
R15042 gnd.n6879 gnd.n477 0.152939
R15043 gnd.n6879 gnd.n6878 0.152939
R15044 gnd.n6878 gnd.n6877 0.152939
R15045 gnd.n6877 gnd.n481 0.152939
R15046 gnd.n6873 gnd.n481 0.152939
R15047 gnd.n6873 gnd.n6872 0.152939
R15048 gnd.n6872 gnd.n6871 0.152939
R15049 gnd.n6871 gnd.n485 0.152939
R15050 gnd.n6867 gnd.n485 0.152939
R15051 gnd.n6867 gnd.n6866 0.152939
R15052 gnd.n6866 gnd.n6865 0.152939
R15053 gnd.n6865 gnd.n489 0.152939
R15054 gnd.n6861 gnd.n489 0.152939
R15055 gnd.n6861 gnd.n6860 0.152939
R15056 gnd.n6860 gnd.n6859 0.152939
R15057 gnd.n6859 gnd.n493 0.152939
R15058 gnd.n6855 gnd.n493 0.152939
R15059 gnd.n6855 gnd.n6854 0.152939
R15060 gnd.n6854 gnd.n63 0.152939
R15061 gnd.n7368 gnd.n64 0.152939
R15062 gnd.n7364 gnd.n64 0.152939
R15063 gnd.n7364 gnd.n7363 0.152939
R15064 gnd.n7363 gnd.n7362 0.152939
R15065 gnd.n7362 gnd.n70 0.152939
R15066 gnd.n7358 gnd.n70 0.152939
R15067 gnd.n7358 gnd.n7357 0.152939
R15068 gnd.n7357 gnd.n7356 0.152939
R15069 gnd.n7356 gnd.n75 0.152939
R15070 gnd.n7352 gnd.n75 0.152939
R15071 gnd.n7352 gnd.n7351 0.152939
R15072 gnd.n7351 gnd.n7350 0.152939
R15073 gnd.n7350 gnd.n80 0.152939
R15074 gnd.n7346 gnd.n80 0.152939
R15075 gnd.n7346 gnd.n7345 0.152939
R15076 gnd.n7345 gnd.n7344 0.152939
R15077 gnd.n7344 gnd.n85 0.152939
R15078 gnd.n7340 gnd.n85 0.152939
R15079 gnd.n7340 gnd.n7339 0.152939
R15080 gnd.n7339 gnd.n7338 0.152939
R15081 gnd.n7338 gnd.n90 0.152939
R15082 gnd.n7334 gnd.n90 0.152939
R15083 gnd.n7334 gnd.n7333 0.152939
R15084 gnd.n7333 gnd.n7332 0.152939
R15085 gnd.n7332 gnd.n95 0.152939
R15086 gnd.n98 gnd.n95 0.152939
R15087 gnd.n5647 gnd.n472 0.151415
R15088 gnd.n5851 gnd.n1347 0.151415
R15089 gnd.n4436 gnd.n1144 0.10111
R15090 gnd.n5570 gnd.n5542 0.10111
R15091 gnd.n3317 gnd.n3316 0.0767195
R15092 gnd.n3316 gnd.n3315 0.0767195
R15093 gnd.n7101 gnd.n255 0.0767195
R15094 gnd.n497 gnd.n277 0.0767195
R15095 gnd.n498 gnd.n277 0.0767195
R15096 gnd.n7053 gnd.n255 0.0767195
R15097 gnd.n6002 gnd.n1143 0.0767195
R15098 gnd.n4379 gnd.n2355 0.0767195
R15099 gnd.n4380 gnd.n4379 0.0767195
R15100 gnd.n4378 gnd.n2356 0.0767195
R15101 gnd.n4378 gnd.n4377 0.0767195
R15102 gnd.n6002 gnd.n1140 0.0767195
R15103 gnd.n7078 gnd.n7077 0.0767195
R15104 gnd.n7079 gnd.n7078 0.0767195
R15105 gnd.n7369 gnd.n63 0.0767195
R15106 gnd.n7369 gnd.n7368 0.0767195
R15107 gnd.n4308 gnd.n4306 0.0695946
R15108 gnd.n4310 gnd.n4308 0.0695946
R15109 gnd.n4610 gnd.n4609 0.063
R15110 gnd.n5704 gnd.n5703 0.063
R15111 gnd.n5570 gnd.n556 0.0523293
R15112 gnd.n4336 gnd.n1144 0.0523293
R15113 gnd.n3883 gnd.n2498 0.0477147
R15114 gnd.n3080 gnd.n2968 0.0442063
R15115 gnd.n3081 gnd.n3080 0.0442063
R15116 gnd.n3082 gnd.n3081 0.0442063
R15117 gnd.n3082 gnd.n2957 0.0442063
R15118 gnd.n3096 gnd.n2957 0.0442063
R15119 gnd.n3097 gnd.n3096 0.0442063
R15120 gnd.n3098 gnd.n3097 0.0442063
R15121 gnd.n3098 gnd.n2944 0.0442063
R15122 gnd.n3142 gnd.n2944 0.0442063
R15123 gnd.n3143 gnd.n3142 0.0442063
R15124 gnd.n3145 gnd.n2878 0.0344674
R15125 gnd.n5651 gnd.n5650 0.0344674
R15126 gnd.n5850 gnd.n1348 0.0344674
R15127 gnd.n3165 gnd.n3164 0.0269946
R15128 gnd.n3167 gnd.n3166 0.0269946
R15129 gnd.n2873 gnd.n2871 0.0269946
R15130 gnd.n3177 gnd.n3175 0.0269946
R15131 gnd.n3176 gnd.n2852 0.0269946
R15132 gnd.n3196 gnd.n3195 0.0269946
R15133 gnd.n3198 gnd.n3197 0.0269946
R15134 gnd.n2847 gnd.n2846 0.0269946
R15135 gnd.n3208 gnd.n2842 0.0269946
R15136 gnd.n3207 gnd.n2844 0.0269946
R15137 gnd.n2843 gnd.n2825 0.0269946
R15138 gnd.n3228 gnd.n2826 0.0269946
R15139 gnd.n3227 gnd.n2827 0.0269946
R15140 gnd.n3261 gnd.n2802 0.0269946
R15141 gnd.n3263 gnd.n3262 0.0269946
R15142 gnd.n3264 gnd.n2749 0.0269946
R15143 gnd.n2797 gnd.n2750 0.0269946
R15144 gnd.n2799 gnd.n2751 0.0269946
R15145 gnd.n3274 gnd.n3273 0.0269946
R15146 gnd.n3276 gnd.n3275 0.0269946
R15147 gnd.n3277 gnd.n2771 0.0269946
R15148 gnd.n3279 gnd.n2772 0.0269946
R15149 gnd.n3282 gnd.n2773 0.0269946
R15150 gnd.n3285 gnd.n3284 0.0269946
R15151 gnd.n3287 gnd.n3286 0.0269946
R15152 gnd.n3352 gnd.n2672 0.0269946
R15153 gnd.n3354 gnd.n3353 0.0269946
R15154 gnd.n3363 gnd.n2665 0.0269946
R15155 gnd.n3365 gnd.n3364 0.0269946
R15156 gnd.n3366 gnd.n2663 0.0269946
R15157 gnd.n3373 gnd.n3369 0.0269946
R15158 gnd.n3372 gnd.n3371 0.0269946
R15159 gnd.n3370 gnd.n2642 0.0269946
R15160 gnd.n3395 gnd.n2643 0.0269946
R15161 gnd.n3394 gnd.n2644 0.0269946
R15162 gnd.n3437 gnd.n2617 0.0269946
R15163 gnd.n3439 gnd.n3438 0.0269946
R15164 gnd.n3448 gnd.n2610 0.0269946
R15165 gnd.n3450 gnd.n3449 0.0269946
R15166 gnd.n3451 gnd.n2608 0.0269946
R15167 gnd.n3458 gnd.n3454 0.0269946
R15168 gnd.n3457 gnd.n3456 0.0269946
R15169 gnd.n3455 gnd.n2587 0.0269946
R15170 gnd.n3480 gnd.n2588 0.0269946
R15171 gnd.n3479 gnd.n2589 0.0269946
R15172 gnd.n3526 gnd.n2562 0.0269946
R15173 gnd.n3528 gnd.n3527 0.0269946
R15174 gnd.n3537 gnd.n2555 0.0269946
R15175 gnd.n3796 gnd.n2553 0.0269946
R15176 gnd.n3801 gnd.n3799 0.0269946
R15177 gnd.n3800 gnd.n2534 0.0269946
R15178 gnd.n3825 gnd.n3824 0.0269946
R15179 gnd.n5704 gnd.n1477 0.0246168
R15180 gnd.n4610 gnd.n2201 0.0246168
R15181 gnd.n3145 gnd.n3144 0.0202011
R15182 gnd.n1481 gnd.n1477 0.0174837
R15183 gnd.n5698 gnd.n1481 0.0174837
R15184 gnd.n5698 gnd.n5697 0.0174837
R15185 gnd.n5697 gnd.n1482 0.0174837
R15186 gnd.n5694 gnd.n1482 0.0174837
R15187 gnd.n5694 gnd.n5693 0.0174837
R15188 gnd.n5693 gnd.n1487 0.0174837
R15189 gnd.n5690 gnd.n1487 0.0174837
R15190 gnd.n5690 gnd.n5689 0.0174837
R15191 gnd.n5689 gnd.n1493 0.0174837
R15192 gnd.n5686 gnd.n1493 0.0174837
R15193 gnd.n5686 gnd.n5685 0.0174837
R15194 gnd.n5685 gnd.n1497 0.0174837
R15195 gnd.n5682 gnd.n1497 0.0174837
R15196 gnd.n5682 gnd.n5681 0.0174837
R15197 gnd.n5681 gnd.n1501 0.0174837
R15198 gnd.n5678 gnd.n1501 0.0174837
R15199 gnd.n5678 gnd.n5677 0.0174837
R15200 gnd.n5677 gnd.n1505 0.0174837
R15201 gnd.n5674 gnd.n1505 0.0174837
R15202 gnd.n5674 gnd.n5673 0.0174837
R15203 gnd.n5673 gnd.n1511 0.0174837
R15204 gnd.n5670 gnd.n1511 0.0174837
R15205 gnd.n5670 gnd.n5669 0.0174837
R15206 gnd.n5669 gnd.n1515 0.0174837
R15207 gnd.n5666 gnd.n1515 0.0174837
R15208 gnd.n5666 gnd.n5665 0.0174837
R15209 gnd.n5665 gnd.n1519 0.0174837
R15210 gnd.n5662 gnd.n1519 0.0174837
R15211 gnd.n5662 gnd.n5661 0.0174837
R15212 gnd.n5661 gnd.n1523 0.0174837
R15213 gnd.n5655 gnd.n1523 0.0174837
R15214 gnd.n5655 gnd.n5654 0.0174837
R15215 gnd.n5654 gnd.n1527 0.0174837
R15216 gnd.n5651 gnd.n1527 0.0174837
R15217 gnd.n2206 gnd.n2201 0.0174837
R15218 gnd.n4605 gnd.n2206 0.0174837
R15219 gnd.n4605 gnd.n4604 0.0174837
R15220 gnd.n4604 gnd.n2207 0.0174837
R15221 gnd.n4601 gnd.n2207 0.0174837
R15222 gnd.n4601 gnd.n4600 0.0174837
R15223 gnd.n4600 gnd.n2212 0.0174837
R15224 gnd.n4597 gnd.n2212 0.0174837
R15225 gnd.n4597 gnd.n4596 0.0174837
R15226 gnd.n4596 gnd.n2218 0.0174837
R15227 gnd.n4593 gnd.n2218 0.0174837
R15228 gnd.n4593 gnd.n4592 0.0174837
R15229 gnd.n4592 gnd.n2222 0.0174837
R15230 gnd.n4589 gnd.n2222 0.0174837
R15231 gnd.n4589 gnd.n4588 0.0174837
R15232 gnd.n4588 gnd.n2229 0.0174837
R15233 gnd.n4585 gnd.n2229 0.0174837
R15234 gnd.n4585 gnd.n4584 0.0174837
R15235 gnd.n4584 gnd.n2233 0.0174837
R15236 gnd.n4581 gnd.n2233 0.0174837
R15237 gnd.n4581 gnd.n4580 0.0174837
R15238 gnd.n4580 gnd.n2239 0.0174837
R15239 gnd.n4577 gnd.n2239 0.0174837
R15240 gnd.n4577 gnd.n4576 0.0174837
R15241 gnd.n4576 gnd.n2243 0.0174837
R15242 gnd.n4573 gnd.n2243 0.0174837
R15243 gnd.n4573 gnd.n4572 0.0174837
R15244 gnd.n4572 gnd.n2250 0.0174837
R15245 gnd.n4569 gnd.n2250 0.0174837
R15246 gnd.n4569 gnd.n4568 0.0174837
R15247 gnd.n4568 gnd.n2254 0.0174837
R15248 gnd.n2260 gnd.n2254 0.0174837
R15249 gnd.n4561 gnd.n2260 0.0174837
R15250 gnd.n4562 gnd.n4561 0.0174837
R15251 gnd.n4562 gnd.n1348 0.0174837
R15252 gnd.n3144 gnd.n3143 0.0148637
R15253 gnd.n3794 gnd.n3538 0.0144266
R15254 gnd.n3795 gnd.n3794 0.0130679
R15255 gnd.n3164 gnd.n2878 0.00797283
R15256 gnd.n3166 gnd.n3165 0.00797283
R15257 gnd.n3167 gnd.n2873 0.00797283
R15258 gnd.n3175 gnd.n2871 0.00797283
R15259 gnd.n3177 gnd.n3176 0.00797283
R15260 gnd.n3195 gnd.n2852 0.00797283
R15261 gnd.n3197 gnd.n3196 0.00797283
R15262 gnd.n3198 gnd.n2847 0.00797283
R15263 gnd.n2846 gnd.n2842 0.00797283
R15264 gnd.n3208 gnd.n3207 0.00797283
R15265 gnd.n2844 gnd.n2843 0.00797283
R15266 gnd.n2826 gnd.n2825 0.00797283
R15267 gnd.n3228 gnd.n3227 0.00797283
R15268 gnd.n2827 gnd.n2802 0.00797283
R15269 gnd.n3262 gnd.n3261 0.00797283
R15270 gnd.n3264 gnd.n3263 0.00797283
R15271 gnd.n2797 gnd.n2749 0.00797283
R15272 gnd.n2799 gnd.n2750 0.00797283
R15273 gnd.n3273 gnd.n2751 0.00797283
R15274 gnd.n3275 gnd.n3274 0.00797283
R15275 gnd.n3277 gnd.n3276 0.00797283
R15276 gnd.n3279 gnd.n2771 0.00797283
R15277 gnd.n3282 gnd.n2772 0.00797283
R15278 gnd.n3284 gnd.n2773 0.00797283
R15279 gnd.n3287 gnd.n3285 0.00797283
R15280 gnd.n3286 gnd.n2672 0.00797283
R15281 gnd.n3354 gnd.n3352 0.00797283
R15282 gnd.n3353 gnd.n2665 0.00797283
R15283 gnd.n3364 gnd.n3363 0.00797283
R15284 gnd.n3366 gnd.n3365 0.00797283
R15285 gnd.n3369 gnd.n2663 0.00797283
R15286 gnd.n3373 gnd.n3372 0.00797283
R15287 gnd.n3371 gnd.n3370 0.00797283
R15288 gnd.n2643 gnd.n2642 0.00797283
R15289 gnd.n3395 gnd.n3394 0.00797283
R15290 gnd.n2644 gnd.n2617 0.00797283
R15291 gnd.n3439 gnd.n3437 0.00797283
R15292 gnd.n3438 gnd.n2610 0.00797283
R15293 gnd.n3449 gnd.n3448 0.00797283
R15294 gnd.n3451 gnd.n3450 0.00797283
R15295 gnd.n3454 gnd.n2608 0.00797283
R15296 gnd.n3458 gnd.n3457 0.00797283
R15297 gnd.n3456 gnd.n3455 0.00797283
R15298 gnd.n2588 gnd.n2587 0.00797283
R15299 gnd.n3480 gnd.n3479 0.00797283
R15300 gnd.n2589 gnd.n2562 0.00797283
R15301 gnd.n3528 gnd.n3526 0.00797283
R15302 gnd.n3527 gnd.n2555 0.00797283
R15303 gnd.n3538 gnd.n3537 0.00797283
R15304 gnd.n3796 gnd.n3795 0.00797283
R15305 gnd.n3799 gnd.n2553 0.00797283
R15306 gnd.n3801 gnd.n3800 0.00797283
R15307 gnd.n3824 gnd.n2534 0.00797283
R15308 gnd.n3825 gnd.n2498 0.00797283
R15309 gnd.n7078 gnd.n277 0.00507153
R15310 gnd.n4379 gnd.n4378 0.00507153
R15311 gnd.n5650 gnd.n472 0.000839674
R15312 gnd.n5851 gnd.n5850 0.000839674
R15313 plus.n43 plus.t18 322.512
R15314 plus.n9 plus.t13 322.512
R15315 plus.n42 plus.t17 297.12
R15316 plus.n46 plus.t22 297.12
R15317 plus.n48 plus.t21 297.12
R15318 plus.n52 plus.t23 297.12
R15319 plus.n54 plus.t8 297.12
R15320 plus.n58 plus.t7 297.12
R15321 plus.n60 plus.t12 297.12
R15322 plus.n64 plus.t10 297.12
R15323 plus.n66 plus.t24 297.12
R15324 plus.n32 plus.t14 297.12
R15325 plus.n30 plus.t15 297.12
R15326 plus.n2 plus.t9 297.12
R15327 plus.n24 plus.t5 297.12
R15328 plus.n4 plus.t6 297.12
R15329 plus.n18 plus.t19 297.12
R15330 plus.n6 plus.t20 297.12
R15331 plus.n12 plus.t16 297.12
R15332 plus.n8 plus.t11 297.12
R15333 plus.n70 plus.t0 243.97
R15334 plus.n70 plus.n69 223.454
R15335 plus.n72 plus.n71 223.454
R15336 plus.n67 plus.n66 161.3
R15337 plus.n65 plus.n34 161.3
R15338 plus.n64 plus.n63 161.3
R15339 plus.n62 plus.n35 161.3
R15340 plus.n61 plus.n60 161.3
R15341 plus.n59 plus.n36 161.3
R15342 plus.n58 plus.n57 161.3
R15343 plus.n56 plus.n37 161.3
R15344 plus.n55 plus.n54 161.3
R15345 plus.n53 plus.n38 161.3
R15346 plus.n52 plus.n51 161.3
R15347 plus.n50 plus.n39 161.3
R15348 plus.n49 plus.n48 161.3
R15349 plus.n47 plus.n40 161.3
R15350 plus.n46 plus.n45 161.3
R15351 plus.n44 plus.n41 161.3
R15352 plus.n11 plus.n10 161.3
R15353 plus.n12 plus.n7 161.3
R15354 plus.n14 plus.n13 161.3
R15355 plus.n15 plus.n6 161.3
R15356 plus.n17 plus.n16 161.3
R15357 plus.n18 plus.n5 161.3
R15358 plus.n20 plus.n19 161.3
R15359 plus.n21 plus.n4 161.3
R15360 plus.n23 plus.n22 161.3
R15361 plus.n24 plus.n3 161.3
R15362 plus.n26 plus.n25 161.3
R15363 plus.n27 plus.n2 161.3
R15364 plus.n29 plus.n28 161.3
R15365 plus.n30 plus.n1 161.3
R15366 plus.n31 plus.n0 161.3
R15367 plus.n33 plus.n32 161.3
R15368 plus.n44 plus.n43 45.0031
R15369 plus.n10 plus.n9 45.0031
R15370 plus.n66 plus.n65 41.6278
R15371 plus.n32 plus.n31 41.6278
R15372 plus.n42 plus.n41 37.246
R15373 plus.n64 plus.n35 37.246
R15374 plus.n30 plus.n29 37.246
R15375 plus.n11 plus.n8 37.246
R15376 plus.n47 plus.n46 32.8641
R15377 plus.n60 plus.n59 32.8641
R15378 plus.n25 plus.n2 32.8641
R15379 plus.n13 plus.n12 32.8641
R15380 plus.n68 plus.n67 31.6047
R15381 plus.n48 plus.n39 28.4823
R15382 plus.n58 plus.n37 28.4823
R15383 plus.n24 plus.n23 28.4823
R15384 plus.n17 plus.n6 28.4823
R15385 plus.n53 plus.n52 24.1005
R15386 plus.n54 plus.n53 24.1005
R15387 plus.n19 plus.n4 24.1005
R15388 plus.n19 plus.n18 24.1005
R15389 plus.n69 plus.t4 19.8005
R15390 plus.n69 plus.t2 19.8005
R15391 plus.n71 plus.t1 19.8005
R15392 plus.n71 plus.t3 19.8005
R15393 plus.n52 plus.n39 19.7187
R15394 plus.n54 plus.n37 19.7187
R15395 plus.n23 plus.n4 19.7187
R15396 plus.n18 plus.n17 19.7187
R15397 plus.n43 plus.n42 15.6319
R15398 plus.n9 plus.n8 15.6319
R15399 plus.n48 plus.n47 15.3369
R15400 plus.n59 plus.n58 15.3369
R15401 plus.n25 plus.n24 15.3369
R15402 plus.n13 plus.n6 15.3369
R15403 plus plus.n73 14.4446
R15404 plus.n68 plus.n33 11.866
R15405 plus.n46 plus.n41 10.955
R15406 plus.n60 plus.n35 10.955
R15407 plus.n29 plus.n2 10.955
R15408 plus.n12 plus.n11 10.955
R15409 plus.n65 plus.n64 6.57323
R15410 plus.n31 plus.n30 6.57323
R15411 plus.n73 plus.n72 5.40567
R15412 plus.n73 plus.n68 1.188
R15413 plus.n72 plus.n70 0.716017
R15414 plus.n45 plus.n44 0.189894
R15415 plus.n45 plus.n40 0.189894
R15416 plus.n49 plus.n40 0.189894
R15417 plus.n50 plus.n49 0.189894
R15418 plus.n51 plus.n50 0.189894
R15419 plus.n51 plus.n38 0.189894
R15420 plus.n55 plus.n38 0.189894
R15421 plus.n56 plus.n55 0.189894
R15422 plus.n57 plus.n56 0.189894
R15423 plus.n57 plus.n36 0.189894
R15424 plus.n61 plus.n36 0.189894
R15425 plus.n62 plus.n61 0.189894
R15426 plus.n63 plus.n62 0.189894
R15427 plus.n63 plus.n34 0.189894
R15428 plus.n67 plus.n34 0.189894
R15429 plus.n33 plus.n0 0.189894
R15430 plus.n1 plus.n0 0.189894
R15431 plus.n28 plus.n1 0.189894
R15432 plus.n28 plus.n27 0.189894
R15433 plus.n27 plus.n26 0.189894
R15434 plus.n26 plus.n3 0.189894
R15435 plus.n22 plus.n3 0.189894
R15436 plus.n22 plus.n21 0.189894
R15437 plus.n21 plus.n20 0.189894
R15438 plus.n20 plus.n5 0.189894
R15439 plus.n16 plus.n5 0.189894
R15440 plus.n16 plus.n15 0.189894
R15441 plus.n15 plus.n14 0.189894
R15442 plus.n14 plus.n7 0.189894
R15443 plus.n10 plus.n7 0.189894
R15444 a_n2903_n3924.n10 a_n2903_n3924.t31 214.944
R15445 a_n2903_n3924.n9 a_n2903_n3924.t2 214.413
R15446 a_n2903_n3924.n9 a_n2903_n3924.t46 214.321
R15447 a_n2903_n3924.n7 a_n2903_n3924.t0 214.321
R15448 a_n2903_n3924.n7 a_n2903_n3924.t47 214.321
R15449 a_n2903_n3924.n8 a_n2903_n3924.t35 214.321
R15450 a_n2903_n3924.n8 a_n2903_n3924.t37 214.321
R15451 a_n2903_n3924.n10 a_n2903_n3924.t8 214.321
R15452 a_n2903_n3924.n1 a_n2903_n3924.t14 55.8337
R15453 a_n2903_n3924.n1 a_n2903_n3924.t40 55.8337
R15454 a_n2903_n3924.n3 a_n2903_n3924.t45 55.8337
R15455 a_n2903_n3924.n0 a_n2903_n3924.t29 55.8335
R15456 a_n2903_n3924.n5 a_n2903_n3924.t5 55.8335
R15457 a_n2903_n3924.n4 a_n2903_n3924.t32 55.8335
R15458 a_n2903_n3924.n4 a_n2903_n3924.t16 55.8335
R15459 a_n2903_n3924.n6 a_n2903_n3924.t22 55.8335
R15460 a_n2903_n3924.n0 a_n2903_n3924.n24 53.0052
R15461 a_n2903_n3924.n1 a_n2903_n3924.n25 53.0052
R15462 a_n2903_n3924.n1 a_n2903_n3924.n26 53.0052
R15463 a_n2903_n3924.n1 a_n2903_n3924.n27 53.0052
R15464 a_n2903_n3924.n2 a_n2903_n3924.n11 53.0052
R15465 a_n2903_n3924.n3 a_n2903_n3924.n12 53.0052
R15466 a_n2903_n3924.n3 a_n2903_n3924.n13 53.0052
R15467 a_n2903_n3924.n5 a_n2903_n3924.n22 53.0051
R15468 a_n2903_n3924.n5 a_n2903_n3924.n21 53.0051
R15469 a_n2903_n3924.n5 a_n2903_n3924.n20 53.0051
R15470 a_n2903_n3924.n4 a_n2903_n3924.n19 53.0051
R15471 a_n2903_n3924.n4 a_n2903_n3924.n18 53.0051
R15472 a_n2903_n3924.n4 a_n2903_n3924.n17 53.0051
R15473 a_n2903_n3924.n4 a_n2903_n3924.n16 53.0051
R15474 a_n2903_n3924.n6 a_n2903_n3924.n15 53.0051
R15475 a_n2903_n3924.n28 a_n2903_n3924.n2 53.0051
R15476 a_n2903_n3924.n14 a_n2903_n3924.n3 12.1986
R15477 a_n2903_n3924.n0 a_n2903_n3924.n23 12.1986
R15478 a_n2903_n3924.n6 a_n2903_n3924.n14 5.11903
R15479 a_n2903_n3924.n23 a_n2903_n3924.n5 5.11903
R15480 a_n2903_n3924.n24 a_n2903_n3924.t18 2.82907
R15481 a_n2903_n3924.n24 a_n2903_n3924.t24 2.82907
R15482 a_n2903_n3924.n25 a_n2903_n3924.t28 2.82907
R15483 a_n2903_n3924.n25 a_n2903_n3924.t26 2.82907
R15484 a_n2903_n3924.n26 a_n2903_n3924.t17 2.82907
R15485 a_n2903_n3924.n26 a_n2903_n3924.t19 2.82907
R15486 a_n2903_n3924.n27 a_n2903_n3924.t11 2.82907
R15487 a_n2903_n3924.n27 a_n2903_n3924.t15 2.82907
R15488 a_n2903_n3924.n11 a_n2903_n3924.t36 2.82907
R15489 a_n2903_n3924.n11 a_n2903_n3924.t42 2.82907
R15490 a_n2903_n3924.n12 a_n2903_n3924.t34 2.82907
R15491 a_n2903_n3924.n12 a_n2903_n3924.t10 2.82907
R15492 a_n2903_n3924.n13 a_n2903_n3924.t7 2.82907
R15493 a_n2903_n3924.n13 a_n2903_n3924.t9 2.82907
R15494 a_n2903_n3924.n22 a_n2903_n3924.t44 2.82907
R15495 a_n2903_n3924.n22 a_n2903_n3924.t43 2.82907
R15496 a_n2903_n3924.n21 a_n2903_n3924.t38 2.82907
R15497 a_n2903_n3924.n21 a_n2903_n3924.t33 2.82907
R15498 a_n2903_n3924.n20 a_n2903_n3924.t4 2.82907
R15499 a_n2903_n3924.n20 a_n2903_n3924.t39 2.82907
R15500 a_n2903_n3924.n19 a_n2903_n3924.t3 2.82907
R15501 a_n2903_n3924.n19 a_n2903_n3924.t6 2.82907
R15502 a_n2903_n3924.n18 a_n2903_n3924.t30 2.82907
R15503 a_n2903_n3924.n18 a_n2903_n3924.t27 2.82907
R15504 a_n2903_n3924.n17 a_n2903_n3924.t21 2.82907
R15505 a_n2903_n3924.n17 a_n2903_n3924.t20 2.82907
R15506 a_n2903_n3924.n16 a_n2903_n3924.t23 2.82907
R15507 a_n2903_n3924.n16 a_n2903_n3924.t12 2.82907
R15508 a_n2903_n3924.n15 a_n2903_n3924.t13 2.82907
R15509 a_n2903_n3924.n15 a_n2903_n3924.t25 2.82907
R15510 a_n2903_n3924.t1 a_n2903_n3924.n28 2.82907
R15511 a_n2903_n3924.n28 a_n2903_n3924.t41 2.82907
R15512 a_n2903_n3924.n5 a_n2903_n3924.n4 2.45524
R15513 a_n2903_n3924.n4 a_n2903_n3924.n6 2.22033
R15514 a_n2903_n3924.n23 a_n2903_n3924.n9 1.95694
R15515 a_n2903_n3924.n14 a_n2903_n3924.n10 1.95694
R15516 a_n2903_n3924.n3 a_n2903_n3924.n2 1.77636
R15517 a_n2903_n3924.n1 a_n2903_n3924.n0 1.77636
R15518 a_n2903_n3924.n10 a_n2903_n3924.n8 1.39367
R15519 a_n2903_n3924.n8 a_n2903_n3924.n7 1.34352
R15520 a_n2903_n3924.n7 a_n2903_n3924.n9 1.25123
R15521 a_n2903_n3924.n2 a_n2903_n3924.n1 1.12334
R15522 a_n7636_8799.n217 a_n7636_8799.t60 485.149
R15523 a_n7636_8799.n279 a_n7636_8799.t72 485.149
R15524 a_n7636_8799.n342 a_n7636_8799.t109 485.149
R15525 a_n7636_8799.n27 a_n7636_8799.t131 485.149
R15526 a_n7636_8799.n89 a_n7636_8799.t146 485.149
R15527 a_n7636_8799.n152 a_n7636_8799.t108 485.149
R15528 a_n7636_8799.n260 a_n7636_8799.t82 464.166
R15529 a_n7636_8799.n259 a_n7636_8799.t81 464.166
R15530 a_n7636_8799.n201 a_n7636_8799.t54 464.166
R15531 a_n7636_8799.n253 a_n7636_8799.t130 464.166
R15532 a_n7636_8799.n252 a_n7636_8799.t85 464.166
R15533 a_n7636_8799.n204 a_n7636_8799.t61 464.166
R15534 a_n7636_8799.n246 a_n7636_8799.t136 464.166
R15535 a_n7636_8799.n245 a_n7636_8799.t102 464.166
R15536 a_n7636_8799.n207 a_n7636_8799.t100 464.166
R15537 a_n7636_8799.n239 a_n7636_8799.t35 464.166
R15538 a_n7636_8799.n238 a_n7636_8799.t106 464.166
R15539 a_n7636_8799.n210 a_n7636_8799.t105 464.166
R15540 a_n7636_8799.n232 a_n7636_8799.t37 464.166
R15541 a_n7636_8799.n231 a_n7636_8799.t36 464.166
R15542 a_n7636_8799.n213 a_n7636_8799.t122 464.166
R15543 a_n7636_8799.n225 a_n7636_8799.t56 464.166
R15544 a_n7636_8799.n224 a_n7636_8799.t40 464.166
R15545 a_n7636_8799.n216 a_n7636_8799.t126 464.166
R15546 a_n7636_8799.n218 a_n7636_8799.t84 464.166
R15547 a_n7636_8799.n322 a_n7636_8799.t92 464.166
R15548 a_n7636_8799.n321 a_n7636_8799.t91 464.166
R15549 a_n7636_8799.n263 a_n7636_8799.t69 464.166
R15550 a_n7636_8799.n315 a_n7636_8799.t145 464.166
R15551 a_n7636_8799.n314 a_n7636_8799.t98 464.166
R15552 a_n7636_8799.n266 a_n7636_8799.t71 464.166
R15553 a_n7636_8799.n308 a_n7636_8799.t151 464.166
R15554 a_n7636_8799.n307 a_n7636_8799.t115 464.166
R15555 a_n7636_8799.n269 a_n7636_8799.t114 464.166
R15556 a_n7636_8799.n301 a_n7636_8799.t45 464.166
R15557 a_n7636_8799.n300 a_n7636_8799.t118 464.166
R15558 a_n7636_8799.n272 a_n7636_8799.t117 464.166
R15559 a_n7636_8799.n294 a_n7636_8799.t49 464.166
R15560 a_n7636_8799.n293 a_n7636_8799.t48 464.166
R15561 a_n7636_8799.n275 a_n7636_8799.t139 464.166
R15562 a_n7636_8799.n287 a_n7636_8799.t70 464.166
R15563 a_n7636_8799.n286 a_n7636_8799.t52 464.166
R15564 a_n7636_8799.n278 a_n7636_8799.t140 464.166
R15565 a_n7636_8799.n280 a_n7636_8799.t99 464.166
R15566 a_n7636_8799.n385 a_n7636_8799.t150 464.166
R15567 a_n7636_8799.n384 a_n7636_8799.t47 464.166
R15568 a_n7636_8799.n326 a_n7636_8799.t97 464.166
R15569 a_n7636_8799.n378 a_n7636_8799.t34 464.166
R15570 a_n7636_8799.n377 a_n7636_8799.t121 464.166
R15571 a_n7636_8799.n329 a_n7636_8799.t58 464.166
R15572 a_n7636_8799.n371 a_n7636_8799.t104 464.166
R15573 a_n7636_8799.n370 a_n7636_8799.t39 464.166
R15574 a_n7636_8799.n332 a_n7636_8799.t64 464.166
R15575 a_n7636_8799.n364 a_n7636_8799.t144 464.166
R15576 a_n7636_8799.n363 a_n7636_8799.t113 464.166
R15577 a_n7636_8799.n335 a_n7636_8799.t138 464.166
R15578 a_n7636_8799.n357 a_n7636_8799.t95 464.166
R15579 a_n7636_8799.n356 a_n7636_8799.t116 464.166
R15580 a_n7636_8799.n338 a_n7636_8799.t51 464.166
R15581 a_n7636_8799.n350 a_n7636_8799.t135 464.166
R15582 a_n7636_8799.n349 a_n7636_8799.t76 464.166
R15583 a_n7636_8799.n341 a_n7636_8799.t127 464.166
R15584 a_n7636_8799.n343 a_n7636_8799.t63 464.166
R15585 a_n7636_8799.n28 a_n7636_8799.t133 464.166
R15586 a_n7636_8799.n30 a_n7636_8799.t83 464.166
R15587 a_n7636_8799.n34 a_n7636_8799.t112 464.166
R15588 a_n7636_8799.n35 a_n7636_8799.t129 464.166
R15589 a_n7636_8799.n23 a_n7636_8799.t79 464.166
R15590 a_n7636_8799.n41 a_n7636_8799.t80 464.166
R15591 a_n7636_8799.n42 a_n7636_8799.t110 464.166
R15592 a_n7636_8799.n46 a_n7636_8799.t67 464.166
R15593 a_n7636_8799.n48 a_n7636_8799.t68 464.166
R15594 a_n7636_8799.n19 a_n7636_8799.t107 464.166
R15595 a_n7636_8799.n53 a_n7636_8799.t32 464.166
R15596 a_n7636_8799.n17 a_n7636_8799.t65 464.166
R15597 a_n7636_8799.n58 a_n7636_8799.t88 464.166
R15598 a_n7636_8799.n60 a_n7636_8799.t132 464.166
R15599 a_n7636_8799.n64 a_n7636_8799.t44 464.166
R15600 a_n7636_8799.n65 a_n7636_8799.t62 464.166
R15601 a_n7636_8799.n13 a_n7636_8799.t128 464.166
R15602 a_n7636_8799.n71 a_n7636_8799.t41 464.166
R15603 a_n7636_8799.n72 a_n7636_8799.t42 464.166
R15604 a_n7636_8799.n90 a_n7636_8799.t149 464.166
R15605 a_n7636_8799.n92 a_n7636_8799.t93 464.166
R15606 a_n7636_8799.n96 a_n7636_8799.t125 464.166
R15607 a_n7636_8799.n97 a_n7636_8799.t143 464.166
R15608 a_n7636_8799.n85 a_n7636_8799.t89 464.166
R15609 a_n7636_8799.n103 a_n7636_8799.t90 464.166
R15610 a_n7636_8799.n104 a_n7636_8799.t123 464.166
R15611 a_n7636_8799.n108 a_n7636_8799.t77 464.166
R15612 a_n7636_8799.n110 a_n7636_8799.t78 464.166
R15613 a_n7636_8799.n81 a_n7636_8799.t119 464.166
R15614 a_n7636_8799.n115 a_n7636_8799.t43 464.166
R15615 a_n7636_8799.n79 a_n7636_8799.t74 464.166
R15616 a_n7636_8799.n120 a_n7636_8799.t101 464.166
R15617 a_n7636_8799.n122 a_n7636_8799.t147 464.166
R15618 a_n7636_8799.n126 a_n7636_8799.t59 464.166
R15619 a_n7636_8799.n127 a_n7636_8799.t73 464.166
R15620 a_n7636_8799.n75 a_n7636_8799.t141 464.166
R15621 a_n7636_8799.n133 a_n7636_8799.t53 464.166
R15622 a_n7636_8799.n134 a_n7636_8799.t55 464.166
R15623 a_n7636_8799.n153 a_n7636_8799.t86 464.166
R15624 a_n7636_8799.n155 a_n7636_8799.t124 464.166
R15625 a_n7636_8799.n159 a_n7636_8799.t75 464.166
R15626 a_n7636_8799.n160 a_n7636_8799.t134 464.166
R15627 a_n7636_8799.n148 a_n7636_8799.t50 464.166
R15628 a_n7636_8799.n166 a_n7636_8799.t33 464.166
R15629 a_n7636_8799.n167 a_n7636_8799.t94 464.166
R15630 a_n7636_8799.n171 a_n7636_8799.t137 464.166
R15631 a_n7636_8799.n173 a_n7636_8799.t111 464.166
R15632 a_n7636_8799.n144 a_n7636_8799.t142 464.166
R15633 a_n7636_8799.n178 a_n7636_8799.t87 464.166
R15634 a_n7636_8799.n142 a_n7636_8799.t38 464.166
R15635 a_n7636_8799.n183 a_n7636_8799.t103 464.166
R15636 a_n7636_8799.n185 a_n7636_8799.t57 464.166
R15637 a_n7636_8799.n189 a_n7636_8799.t120 464.166
R15638 a_n7636_8799.n190 a_n7636_8799.t66 464.166
R15639 a_n7636_8799.n138 a_n7636_8799.t96 464.166
R15640 a_n7636_8799.n196 a_n7636_8799.t46 464.166
R15641 a_n7636_8799.n197 a_n7636_8799.t148 464.166
R15642 a_n7636_8799.n220 a_n7636_8799.n219 161.3
R15643 a_n7636_8799.n221 a_n7636_8799.n216 161.3
R15644 a_n7636_8799.n223 a_n7636_8799.n222 161.3
R15645 a_n7636_8799.n224 a_n7636_8799.n215 161.3
R15646 a_n7636_8799.n225 a_n7636_8799.n214 161.3
R15647 a_n7636_8799.n227 a_n7636_8799.n226 161.3
R15648 a_n7636_8799.n228 a_n7636_8799.n213 161.3
R15649 a_n7636_8799.n230 a_n7636_8799.n229 161.3
R15650 a_n7636_8799.n231 a_n7636_8799.n212 161.3
R15651 a_n7636_8799.n232 a_n7636_8799.n211 161.3
R15652 a_n7636_8799.n234 a_n7636_8799.n233 161.3
R15653 a_n7636_8799.n235 a_n7636_8799.n210 161.3
R15654 a_n7636_8799.n237 a_n7636_8799.n236 161.3
R15655 a_n7636_8799.n238 a_n7636_8799.n209 161.3
R15656 a_n7636_8799.n239 a_n7636_8799.n208 161.3
R15657 a_n7636_8799.n241 a_n7636_8799.n240 161.3
R15658 a_n7636_8799.n242 a_n7636_8799.n207 161.3
R15659 a_n7636_8799.n244 a_n7636_8799.n243 161.3
R15660 a_n7636_8799.n245 a_n7636_8799.n206 161.3
R15661 a_n7636_8799.n246 a_n7636_8799.n205 161.3
R15662 a_n7636_8799.n248 a_n7636_8799.n247 161.3
R15663 a_n7636_8799.n249 a_n7636_8799.n204 161.3
R15664 a_n7636_8799.n251 a_n7636_8799.n250 161.3
R15665 a_n7636_8799.n252 a_n7636_8799.n203 161.3
R15666 a_n7636_8799.n253 a_n7636_8799.n202 161.3
R15667 a_n7636_8799.n255 a_n7636_8799.n254 161.3
R15668 a_n7636_8799.n256 a_n7636_8799.n201 161.3
R15669 a_n7636_8799.n258 a_n7636_8799.n257 161.3
R15670 a_n7636_8799.n259 a_n7636_8799.n200 161.3
R15671 a_n7636_8799.n261 a_n7636_8799.n260 161.3
R15672 a_n7636_8799.n282 a_n7636_8799.n281 161.3
R15673 a_n7636_8799.n283 a_n7636_8799.n278 161.3
R15674 a_n7636_8799.n285 a_n7636_8799.n284 161.3
R15675 a_n7636_8799.n286 a_n7636_8799.n277 161.3
R15676 a_n7636_8799.n287 a_n7636_8799.n276 161.3
R15677 a_n7636_8799.n289 a_n7636_8799.n288 161.3
R15678 a_n7636_8799.n290 a_n7636_8799.n275 161.3
R15679 a_n7636_8799.n292 a_n7636_8799.n291 161.3
R15680 a_n7636_8799.n293 a_n7636_8799.n274 161.3
R15681 a_n7636_8799.n294 a_n7636_8799.n273 161.3
R15682 a_n7636_8799.n296 a_n7636_8799.n295 161.3
R15683 a_n7636_8799.n297 a_n7636_8799.n272 161.3
R15684 a_n7636_8799.n299 a_n7636_8799.n298 161.3
R15685 a_n7636_8799.n300 a_n7636_8799.n271 161.3
R15686 a_n7636_8799.n301 a_n7636_8799.n270 161.3
R15687 a_n7636_8799.n303 a_n7636_8799.n302 161.3
R15688 a_n7636_8799.n304 a_n7636_8799.n269 161.3
R15689 a_n7636_8799.n306 a_n7636_8799.n305 161.3
R15690 a_n7636_8799.n307 a_n7636_8799.n268 161.3
R15691 a_n7636_8799.n308 a_n7636_8799.n267 161.3
R15692 a_n7636_8799.n310 a_n7636_8799.n309 161.3
R15693 a_n7636_8799.n311 a_n7636_8799.n266 161.3
R15694 a_n7636_8799.n313 a_n7636_8799.n312 161.3
R15695 a_n7636_8799.n314 a_n7636_8799.n265 161.3
R15696 a_n7636_8799.n315 a_n7636_8799.n264 161.3
R15697 a_n7636_8799.n317 a_n7636_8799.n316 161.3
R15698 a_n7636_8799.n318 a_n7636_8799.n263 161.3
R15699 a_n7636_8799.n320 a_n7636_8799.n319 161.3
R15700 a_n7636_8799.n321 a_n7636_8799.n262 161.3
R15701 a_n7636_8799.n323 a_n7636_8799.n322 161.3
R15702 a_n7636_8799.n345 a_n7636_8799.n344 161.3
R15703 a_n7636_8799.n346 a_n7636_8799.n341 161.3
R15704 a_n7636_8799.n348 a_n7636_8799.n347 161.3
R15705 a_n7636_8799.n349 a_n7636_8799.n340 161.3
R15706 a_n7636_8799.n350 a_n7636_8799.n339 161.3
R15707 a_n7636_8799.n352 a_n7636_8799.n351 161.3
R15708 a_n7636_8799.n353 a_n7636_8799.n338 161.3
R15709 a_n7636_8799.n355 a_n7636_8799.n354 161.3
R15710 a_n7636_8799.n356 a_n7636_8799.n337 161.3
R15711 a_n7636_8799.n357 a_n7636_8799.n336 161.3
R15712 a_n7636_8799.n359 a_n7636_8799.n358 161.3
R15713 a_n7636_8799.n360 a_n7636_8799.n335 161.3
R15714 a_n7636_8799.n362 a_n7636_8799.n361 161.3
R15715 a_n7636_8799.n363 a_n7636_8799.n334 161.3
R15716 a_n7636_8799.n364 a_n7636_8799.n333 161.3
R15717 a_n7636_8799.n366 a_n7636_8799.n365 161.3
R15718 a_n7636_8799.n367 a_n7636_8799.n332 161.3
R15719 a_n7636_8799.n369 a_n7636_8799.n368 161.3
R15720 a_n7636_8799.n370 a_n7636_8799.n331 161.3
R15721 a_n7636_8799.n371 a_n7636_8799.n330 161.3
R15722 a_n7636_8799.n373 a_n7636_8799.n372 161.3
R15723 a_n7636_8799.n374 a_n7636_8799.n329 161.3
R15724 a_n7636_8799.n376 a_n7636_8799.n375 161.3
R15725 a_n7636_8799.n377 a_n7636_8799.n328 161.3
R15726 a_n7636_8799.n378 a_n7636_8799.n327 161.3
R15727 a_n7636_8799.n380 a_n7636_8799.n379 161.3
R15728 a_n7636_8799.n381 a_n7636_8799.n326 161.3
R15729 a_n7636_8799.n383 a_n7636_8799.n382 161.3
R15730 a_n7636_8799.n384 a_n7636_8799.n325 161.3
R15731 a_n7636_8799.n386 a_n7636_8799.n385 161.3
R15732 a_n7636_8799.n73 a_n7636_8799.n72 161.3
R15733 a_n7636_8799.n71 a_n7636_8799.n12 161.3
R15734 a_n7636_8799.n70 a_n7636_8799.n69 161.3
R15735 a_n7636_8799.n68 a_n7636_8799.n13 161.3
R15736 a_n7636_8799.n67 a_n7636_8799.n66 161.3
R15737 a_n7636_8799.n65 a_n7636_8799.n14 161.3
R15738 a_n7636_8799.n64 a_n7636_8799.n63 161.3
R15739 a_n7636_8799.n62 a_n7636_8799.n15 161.3
R15740 a_n7636_8799.n61 a_n7636_8799.n60 161.3
R15741 a_n7636_8799.n59 a_n7636_8799.n16 161.3
R15742 a_n7636_8799.n58 a_n7636_8799.n57 161.3
R15743 a_n7636_8799.n56 a_n7636_8799.n17 161.3
R15744 a_n7636_8799.n55 a_n7636_8799.n54 161.3
R15745 a_n7636_8799.n53 a_n7636_8799.n18 161.3
R15746 a_n7636_8799.n52 a_n7636_8799.n51 161.3
R15747 a_n7636_8799.n50 a_n7636_8799.n19 161.3
R15748 a_n7636_8799.n49 a_n7636_8799.n48 161.3
R15749 a_n7636_8799.n47 a_n7636_8799.n20 161.3
R15750 a_n7636_8799.n46 a_n7636_8799.n45 161.3
R15751 a_n7636_8799.n44 a_n7636_8799.n21 161.3
R15752 a_n7636_8799.n43 a_n7636_8799.n42 161.3
R15753 a_n7636_8799.n41 a_n7636_8799.n22 161.3
R15754 a_n7636_8799.n40 a_n7636_8799.n39 161.3
R15755 a_n7636_8799.n38 a_n7636_8799.n23 161.3
R15756 a_n7636_8799.n37 a_n7636_8799.n36 161.3
R15757 a_n7636_8799.n35 a_n7636_8799.n24 161.3
R15758 a_n7636_8799.n34 a_n7636_8799.n33 161.3
R15759 a_n7636_8799.n32 a_n7636_8799.n25 161.3
R15760 a_n7636_8799.n31 a_n7636_8799.n30 161.3
R15761 a_n7636_8799.n29 a_n7636_8799.n26 161.3
R15762 a_n7636_8799.n135 a_n7636_8799.n134 161.3
R15763 a_n7636_8799.n133 a_n7636_8799.n74 161.3
R15764 a_n7636_8799.n132 a_n7636_8799.n131 161.3
R15765 a_n7636_8799.n130 a_n7636_8799.n75 161.3
R15766 a_n7636_8799.n129 a_n7636_8799.n128 161.3
R15767 a_n7636_8799.n127 a_n7636_8799.n76 161.3
R15768 a_n7636_8799.n126 a_n7636_8799.n125 161.3
R15769 a_n7636_8799.n124 a_n7636_8799.n77 161.3
R15770 a_n7636_8799.n123 a_n7636_8799.n122 161.3
R15771 a_n7636_8799.n121 a_n7636_8799.n78 161.3
R15772 a_n7636_8799.n120 a_n7636_8799.n119 161.3
R15773 a_n7636_8799.n118 a_n7636_8799.n79 161.3
R15774 a_n7636_8799.n117 a_n7636_8799.n116 161.3
R15775 a_n7636_8799.n115 a_n7636_8799.n80 161.3
R15776 a_n7636_8799.n114 a_n7636_8799.n113 161.3
R15777 a_n7636_8799.n112 a_n7636_8799.n81 161.3
R15778 a_n7636_8799.n111 a_n7636_8799.n110 161.3
R15779 a_n7636_8799.n109 a_n7636_8799.n82 161.3
R15780 a_n7636_8799.n108 a_n7636_8799.n107 161.3
R15781 a_n7636_8799.n106 a_n7636_8799.n83 161.3
R15782 a_n7636_8799.n105 a_n7636_8799.n104 161.3
R15783 a_n7636_8799.n103 a_n7636_8799.n84 161.3
R15784 a_n7636_8799.n102 a_n7636_8799.n101 161.3
R15785 a_n7636_8799.n100 a_n7636_8799.n85 161.3
R15786 a_n7636_8799.n99 a_n7636_8799.n98 161.3
R15787 a_n7636_8799.n97 a_n7636_8799.n86 161.3
R15788 a_n7636_8799.n96 a_n7636_8799.n95 161.3
R15789 a_n7636_8799.n94 a_n7636_8799.n87 161.3
R15790 a_n7636_8799.n93 a_n7636_8799.n92 161.3
R15791 a_n7636_8799.n91 a_n7636_8799.n88 161.3
R15792 a_n7636_8799.n198 a_n7636_8799.n197 161.3
R15793 a_n7636_8799.n196 a_n7636_8799.n137 161.3
R15794 a_n7636_8799.n195 a_n7636_8799.n194 161.3
R15795 a_n7636_8799.n193 a_n7636_8799.n138 161.3
R15796 a_n7636_8799.n192 a_n7636_8799.n191 161.3
R15797 a_n7636_8799.n190 a_n7636_8799.n139 161.3
R15798 a_n7636_8799.n189 a_n7636_8799.n188 161.3
R15799 a_n7636_8799.n187 a_n7636_8799.n140 161.3
R15800 a_n7636_8799.n186 a_n7636_8799.n185 161.3
R15801 a_n7636_8799.n184 a_n7636_8799.n141 161.3
R15802 a_n7636_8799.n183 a_n7636_8799.n182 161.3
R15803 a_n7636_8799.n181 a_n7636_8799.n142 161.3
R15804 a_n7636_8799.n180 a_n7636_8799.n179 161.3
R15805 a_n7636_8799.n178 a_n7636_8799.n143 161.3
R15806 a_n7636_8799.n177 a_n7636_8799.n176 161.3
R15807 a_n7636_8799.n175 a_n7636_8799.n144 161.3
R15808 a_n7636_8799.n174 a_n7636_8799.n173 161.3
R15809 a_n7636_8799.n172 a_n7636_8799.n145 161.3
R15810 a_n7636_8799.n171 a_n7636_8799.n170 161.3
R15811 a_n7636_8799.n169 a_n7636_8799.n146 161.3
R15812 a_n7636_8799.n168 a_n7636_8799.n167 161.3
R15813 a_n7636_8799.n166 a_n7636_8799.n147 161.3
R15814 a_n7636_8799.n165 a_n7636_8799.n164 161.3
R15815 a_n7636_8799.n163 a_n7636_8799.n148 161.3
R15816 a_n7636_8799.n162 a_n7636_8799.n161 161.3
R15817 a_n7636_8799.n160 a_n7636_8799.n149 161.3
R15818 a_n7636_8799.n159 a_n7636_8799.n158 161.3
R15819 a_n7636_8799.n157 a_n7636_8799.n150 161.3
R15820 a_n7636_8799.n156 a_n7636_8799.n155 161.3
R15821 a_n7636_8799.n154 a_n7636_8799.n151 161.3
R15822 a_n7636_8799.n8 a_n7636_8799.n6 98.9633
R15823 a_n7636_8799.n3 a_n7636_8799.n1 98.9631
R15824 a_n7636_8799.n10 a_n7636_8799.n9 98.6055
R15825 a_n7636_8799.n8 a_n7636_8799.n7 98.6055
R15826 a_n7636_8799.n3 a_n7636_8799.n2 98.6055
R15827 a_n7636_8799.n5 a_n7636_8799.n4 98.6055
R15828 a_n7636_8799.n392 a_n7636_8799.n390 81.3764
R15829 a_n7636_8799.n401 a_n7636_8799.n399 81.3764
R15830 a_n7636_8799.n404 a_n7636_8799.n0 81.3764
R15831 a_n7636_8799.n405 a_n7636_8799.n404 80.9326
R15832 a_n7636_8799.n398 a_n7636_8799.n397 80.9324
R15833 a_n7636_8799.n396 a_n7636_8799.n395 80.9324
R15834 a_n7636_8799.n394 a_n7636_8799.n393 80.9324
R15835 a_n7636_8799.n392 a_n7636_8799.n391 80.9324
R15836 a_n7636_8799.n401 a_n7636_8799.n400 80.9324
R15837 a_n7636_8799.n403 a_n7636_8799.n402 80.9324
R15838 a_n7636_8799.n220 a_n7636_8799.n217 70.4033
R15839 a_n7636_8799.n282 a_n7636_8799.n279 70.4033
R15840 a_n7636_8799.n345 a_n7636_8799.n342 70.4033
R15841 a_n7636_8799.n27 a_n7636_8799.n26 70.4033
R15842 a_n7636_8799.n89 a_n7636_8799.n88 70.4033
R15843 a_n7636_8799.n152 a_n7636_8799.n151 70.4033
R15844 a_n7636_8799.n260 a_n7636_8799.n259 48.2005
R15845 a_n7636_8799.n253 a_n7636_8799.n252 48.2005
R15846 a_n7636_8799.n246 a_n7636_8799.n245 48.2005
R15847 a_n7636_8799.n239 a_n7636_8799.n238 48.2005
R15848 a_n7636_8799.n232 a_n7636_8799.n231 48.2005
R15849 a_n7636_8799.n225 a_n7636_8799.n224 48.2005
R15850 a_n7636_8799.n322 a_n7636_8799.n321 48.2005
R15851 a_n7636_8799.n315 a_n7636_8799.n314 48.2005
R15852 a_n7636_8799.n308 a_n7636_8799.n307 48.2005
R15853 a_n7636_8799.n301 a_n7636_8799.n300 48.2005
R15854 a_n7636_8799.n294 a_n7636_8799.n293 48.2005
R15855 a_n7636_8799.n287 a_n7636_8799.n286 48.2005
R15856 a_n7636_8799.n385 a_n7636_8799.n384 48.2005
R15857 a_n7636_8799.n378 a_n7636_8799.n377 48.2005
R15858 a_n7636_8799.n371 a_n7636_8799.n370 48.2005
R15859 a_n7636_8799.n364 a_n7636_8799.n363 48.2005
R15860 a_n7636_8799.n357 a_n7636_8799.n356 48.2005
R15861 a_n7636_8799.n350 a_n7636_8799.n349 48.2005
R15862 a_n7636_8799.n35 a_n7636_8799.n34 48.2005
R15863 a_n7636_8799.n42 a_n7636_8799.n41 48.2005
R15864 a_n7636_8799.n48 a_n7636_8799.n19 48.2005
R15865 a_n7636_8799.n58 a_n7636_8799.n17 48.2005
R15866 a_n7636_8799.n65 a_n7636_8799.n64 48.2005
R15867 a_n7636_8799.n72 a_n7636_8799.n71 48.2005
R15868 a_n7636_8799.n97 a_n7636_8799.n96 48.2005
R15869 a_n7636_8799.n104 a_n7636_8799.n103 48.2005
R15870 a_n7636_8799.n110 a_n7636_8799.n81 48.2005
R15871 a_n7636_8799.n120 a_n7636_8799.n79 48.2005
R15872 a_n7636_8799.n127 a_n7636_8799.n126 48.2005
R15873 a_n7636_8799.n134 a_n7636_8799.n133 48.2005
R15874 a_n7636_8799.n160 a_n7636_8799.n159 48.2005
R15875 a_n7636_8799.n167 a_n7636_8799.n166 48.2005
R15876 a_n7636_8799.n173 a_n7636_8799.n144 48.2005
R15877 a_n7636_8799.n183 a_n7636_8799.n142 48.2005
R15878 a_n7636_8799.n190 a_n7636_8799.n189 48.2005
R15879 a_n7636_8799.n197 a_n7636_8799.n196 48.2005
R15880 a_n7636_8799.n258 a_n7636_8799.n201 40.1672
R15881 a_n7636_8799.n219 a_n7636_8799.n216 40.1672
R15882 a_n7636_8799.n320 a_n7636_8799.n263 40.1672
R15883 a_n7636_8799.n281 a_n7636_8799.n278 40.1672
R15884 a_n7636_8799.n383 a_n7636_8799.n326 40.1672
R15885 a_n7636_8799.n344 a_n7636_8799.n341 40.1672
R15886 a_n7636_8799.n30 a_n7636_8799.n29 40.1672
R15887 a_n7636_8799.n70 a_n7636_8799.n13 40.1672
R15888 a_n7636_8799.n92 a_n7636_8799.n91 40.1672
R15889 a_n7636_8799.n132 a_n7636_8799.n75 40.1672
R15890 a_n7636_8799.n155 a_n7636_8799.n154 40.1672
R15891 a_n7636_8799.n195 a_n7636_8799.n138 40.1672
R15892 a_n7636_8799.n251 a_n7636_8799.n204 38.7066
R15893 a_n7636_8799.n226 a_n7636_8799.n213 38.7066
R15894 a_n7636_8799.n313 a_n7636_8799.n266 38.7066
R15895 a_n7636_8799.n288 a_n7636_8799.n275 38.7066
R15896 a_n7636_8799.n376 a_n7636_8799.n329 38.7066
R15897 a_n7636_8799.n351 a_n7636_8799.n338 38.7066
R15898 a_n7636_8799.n36 a_n7636_8799.n23 38.7066
R15899 a_n7636_8799.n60 a_n7636_8799.n15 38.7066
R15900 a_n7636_8799.n98 a_n7636_8799.n85 38.7066
R15901 a_n7636_8799.n122 a_n7636_8799.n77 38.7066
R15902 a_n7636_8799.n161 a_n7636_8799.n148 38.7066
R15903 a_n7636_8799.n185 a_n7636_8799.n140 38.7066
R15904 a_n7636_8799.n244 a_n7636_8799.n207 37.246
R15905 a_n7636_8799.n233 a_n7636_8799.n210 37.246
R15906 a_n7636_8799.n306 a_n7636_8799.n269 37.246
R15907 a_n7636_8799.n295 a_n7636_8799.n272 37.246
R15908 a_n7636_8799.n369 a_n7636_8799.n332 37.246
R15909 a_n7636_8799.n358 a_n7636_8799.n335 37.246
R15910 a_n7636_8799.n46 a_n7636_8799.n21 37.246
R15911 a_n7636_8799.n54 a_n7636_8799.n53 37.246
R15912 a_n7636_8799.n108 a_n7636_8799.n83 37.246
R15913 a_n7636_8799.n116 a_n7636_8799.n115 37.246
R15914 a_n7636_8799.n171 a_n7636_8799.n146 37.246
R15915 a_n7636_8799.n179 a_n7636_8799.n178 37.246
R15916 a_n7636_8799.n240 a_n7636_8799.n207 35.7853
R15917 a_n7636_8799.n237 a_n7636_8799.n210 35.7853
R15918 a_n7636_8799.n302 a_n7636_8799.n269 35.7853
R15919 a_n7636_8799.n299 a_n7636_8799.n272 35.7853
R15920 a_n7636_8799.n365 a_n7636_8799.n332 35.7853
R15921 a_n7636_8799.n362 a_n7636_8799.n335 35.7853
R15922 a_n7636_8799.n47 a_n7636_8799.n46 35.7853
R15923 a_n7636_8799.n53 a_n7636_8799.n52 35.7853
R15924 a_n7636_8799.n109 a_n7636_8799.n108 35.7853
R15925 a_n7636_8799.n115 a_n7636_8799.n114 35.7853
R15926 a_n7636_8799.n172 a_n7636_8799.n171 35.7853
R15927 a_n7636_8799.n178 a_n7636_8799.n177 35.7853
R15928 a_n7636_8799.n247 a_n7636_8799.n204 34.3247
R15929 a_n7636_8799.n230 a_n7636_8799.n213 34.3247
R15930 a_n7636_8799.n309 a_n7636_8799.n266 34.3247
R15931 a_n7636_8799.n292 a_n7636_8799.n275 34.3247
R15932 a_n7636_8799.n372 a_n7636_8799.n329 34.3247
R15933 a_n7636_8799.n355 a_n7636_8799.n338 34.3247
R15934 a_n7636_8799.n40 a_n7636_8799.n23 34.3247
R15935 a_n7636_8799.n60 a_n7636_8799.n59 34.3247
R15936 a_n7636_8799.n102 a_n7636_8799.n85 34.3247
R15937 a_n7636_8799.n122 a_n7636_8799.n121 34.3247
R15938 a_n7636_8799.n165 a_n7636_8799.n148 34.3247
R15939 a_n7636_8799.n185 a_n7636_8799.n184 34.3247
R15940 a_n7636_8799.n254 a_n7636_8799.n201 32.8641
R15941 a_n7636_8799.n223 a_n7636_8799.n216 32.8641
R15942 a_n7636_8799.n316 a_n7636_8799.n263 32.8641
R15943 a_n7636_8799.n285 a_n7636_8799.n278 32.8641
R15944 a_n7636_8799.n379 a_n7636_8799.n326 32.8641
R15945 a_n7636_8799.n348 a_n7636_8799.n341 32.8641
R15946 a_n7636_8799.n30 a_n7636_8799.n25 32.8641
R15947 a_n7636_8799.n66 a_n7636_8799.n13 32.8641
R15948 a_n7636_8799.n92 a_n7636_8799.n87 32.8641
R15949 a_n7636_8799.n128 a_n7636_8799.n75 32.8641
R15950 a_n7636_8799.n155 a_n7636_8799.n150 32.8641
R15951 a_n7636_8799.n191 a_n7636_8799.n138 32.8641
R15952 a_n7636_8799.n403 a_n7636_8799.n398 32.7526
R15953 a_n7636_8799.n11 a_n7636_8799.n5 30.7135
R15954 a_n7636_8799.n218 a_n7636_8799.n217 20.9576
R15955 a_n7636_8799.n280 a_n7636_8799.n279 20.9576
R15956 a_n7636_8799.n343 a_n7636_8799.n342 20.9576
R15957 a_n7636_8799.n28 a_n7636_8799.n27 20.9576
R15958 a_n7636_8799.n90 a_n7636_8799.n89 20.9576
R15959 a_n7636_8799.n153 a_n7636_8799.n152 20.9576
R15960 a_n7636_8799.n11 a_n7636_8799.n10 17.7361
R15961 a_n7636_8799.n254 a_n7636_8799.n253 15.3369
R15962 a_n7636_8799.n224 a_n7636_8799.n223 15.3369
R15963 a_n7636_8799.n316 a_n7636_8799.n315 15.3369
R15964 a_n7636_8799.n286 a_n7636_8799.n285 15.3369
R15965 a_n7636_8799.n379 a_n7636_8799.n378 15.3369
R15966 a_n7636_8799.n349 a_n7636_8799.n348 15.3369
R15967 a_n7636_8799.n34 a_n7636_8799.n25 15.3369
R15968 a_n7636_8799.n66 a_n7636_8799.n65 15.3369
R15969 a_n7636_8799.n96 a_n7636_8799.n87 15.3369
R15970 a_n7636_8799.n128 a_n7636_8799.n127 15.3369
R15971 a_n7636_8799.n159 a_n7636_8799.n150 15.3369
R15972 a_n7636_8799.n191 a_n7636_8799.n190 15.3369
R15973 a_n7636_8799.n247 a_n7636_8799.n246 13.8763
R15974 a_n7636_8799.n231 a_n7636_8799.n230 13.8763
R15975 a_n7636_8799.n309 a_n7636_8799.n308 13.8763
R15976 a_n7636_8799.n293 a_n7636_8799.n292 13.8763
R15977 a_n7636_8799.n372 a_n7636_8799.n371 13.8763
R15978 a_n7636_8799.n356 a_n7636_8799.n355 13.8763
R15979 a_n7636_8799.n41 a_n7636_8799.n40 13.8763
R15980 a_n7636_8799.n59 a_n7636_8799.n58 13.8763
R15981 a_n7636_8799.n103 a_n7636_8799.n102 13.8763
R15982 a_n7636_8799.n121 a_n7636_8799.n120 13.8763
R15983 a_n7636_8799.n166 a_n7636_8799.n165 13.8763
R15984 a_n7636_8799.n184 a_n7636_8799.n183 13.8763
R15985 a_n7636_8799.n240 a_n7636_8799.n239 12.4157
R15986 a_n7636_8799.n238 a_n7636_8799.n237 12.4157
R15987 a_n7636_8799.n302 a_n7636_8799.n301 12.4157
R15988 a_n7636_8799.n300 a_n7636_8799.n299 12.4157
R15989 a_n7636_8799.n365 a_n7636_8799.n364 12.4157
R15990 a_n7636_8799.n363 a_n7636_8799.n362 12.4157
R15991 a_n7636_8799.n48 a_n7636_8799.n47 12.4157
R15992 a_n7636_8799.n52 a_n7636_8799.n19 12.4157
R15993 a_n7636_8799.n110 a_n7636_8799.n109 12.4157
R15994 a_n7636_8799.n114 a_n7636_8799.n81 12.4157
R15995 a_n7636_8799.n173 a_n7636_8799.n172 12.4157
R15996 a_n7636_8799.n177 a_n7636_8799.n144 12.4157
R15997 a_n7636_8799.n394 a_n7636_8799.n389 12.3339
R15998 a_n7636_8799.n389 a_n7636_8799.n11 11.4887
R15999 a_n7636_8799.n245 a_n7636_8799.n244 10.955
R16000 a_n7636_8799.n233 a_n7636_8799.n232 10.955
R16001 a_n7636_8799.n307 a_n7636_8799.n306 10.955
R16002 a_n7636_8799.n295 a_n7636_8799.n294 10.955
R16003 a_n7636_8799.n370 a_n7636_8799.n369 10.955
R16004 a_n7636_8799.n358 a_n7636_8799.n357 10.955
R16005 a_n7636_8799.n42 a_n7636_8799.n21 10.955
R16006 a_n7636_8799.n54 a_n7636_8799.n17 10.955
R16007 a_n7636_8799.n104 a_n7636_8799.n83 10.955
R16008 a_n7636_8799.n116 a_n7636_8799.n79 10.955
R16009 a_n7636_8799.n167 a_n7636_8799.n146 10.955
R16010 a_n7636_8799.n179 a_n7636_8799.n142 10.955
R16011 a_n7636_8799.n252 a_n7636_8799.n251 9.49444
R16012 a_n7636_8799.n226 a_n7636_8799.n225 9.49444
R16013 a_n7636_8799.n314 a_n7636_8799.n313 9.49444
R16014 a_n7636_8799.n288 a_n7636_8799.n287 9.49444
R16015 a_n7636_8799.n377 a_n7636_8799.n376 9.49444
R16016 a_n7636_8799.n351 a_n7636_8799.n350 9.49444
R16017 a_n7636_8799.n36 a_n7636_8799.n35 9.49444
R16018 a_n7636_8799.n64 a_n7636_8799.n15 9.49444
R16019 a_n7636_8799.n98 a_n7636_8799.n97 9.49444
R16020 a_n7636_8799.n126 a_n7636_8799.n77 9.49444
R16021 a_n7636_8799.n161 a_n7636_8799.n160 9.49444
R16022 a_n7636_8799.n189 a_n7636_8799.n140 9.49444
R16023 a_n7636_8799.n324 a_n7636_8799.n261 9.04406
R16024 a_n7636_8799.n136 a_n7636_8799.n73 9.04406
R16025 a_n7636_8799.n259 a_n7636_8799.n258 8.03383
R16026 a_n7636_8799.n219 a_n7636_8799.n218 8.03383
R16027 a_n7636_8799.n321 a_n7636_8799.n320 8.03383
R16028 a_n7636_8799.n281 a_n7636_8799.n280 8.03383
R16029 a_n7636_8799.n384 a_n7636_8799.n383 8.03383
R16030 a_n7636_8799.n344 a_n7636_8799.n343 8.03383
R16031 a_n7636_8799.n29 a_n7636_8799.n28 8.03383
R16032 a_n7636_8799.n71 a_n7636_8799.n70 8.03383
R16033 a_n7636_8799.n91 a_n7636_8799.n90 8.03383
R16034 a_n7636_8799.n133 a_n7636_8799.n132 8.03383
R16035 a_n7636_8799.n154 a_n7636_8799.n153 8.03383
R16036 a_n7636_8799.n196 a_n7636_8799.n195 8.03383
R16037 a_n7636_8799.n388 a_n7636_8799.n199 6.86985
R16038 a_n7636_8799.n388 a_n7636_8799.n387 6.51296
R16039 a_n7636_8799.n324 a_n7636_8799.n323 4.93611
R16040 a_n7636_8799.n387 a_n7636_8799.n386 4.93611
R16041 a_n7636_8799.n136 a_n7636_8799.n135 4.93611
R16042 a_n7636_8799.n199 a_n7636_8799.n198 4.93611
R16043 a_n7636_8799.n387 a_n7636_8799.n324 4.10845
R16044 a_n7636_8799.n199 a_n7636_8799.n136 4.10845
R16045 a_n7636_8799.n9 a_n7636_8799.t1 3.61217
R16046 a_n7636_8799.n9 a_n7636_8799.t27 3.61217
R16047 a_n7636_8799.n7 a_n7636_8799.t30 3.61217
R16048 a_n7636_8799.n7 a_n7636_8799.t26 3.61217
R16049 a_n7636_8799.n6 a_n7636_8799.t23 3.61217
R16050 a_n7636_8799.n6 a_n7636_8799.t25 3.61217
R16051 a_n7636_8799.n1 a_n7636_8799.t28 3.61217
R16052 a_n7636_8799.n1 a_n7636_8799.t24 3.61217
R16053 a_n7636_8799.n2 a_n7636_8799.t2 3.61217
R16054 a_n7636_8799.n2 a_n7636_8799.t29 3.61217
R16055 a_n7636_8799.n4 a_n7636_8799.t0 3.61217
R16056 a_n7636_8799.n4 a_n7636_8799.t31 3.61217
R16057 a_n7636_8799.n389 a_n7636_8799.n388 3.4105
R16058 a_n7636_8799.n399 a_n7636_8799.t16 2.82907
R16059 a_n7636_8799.n399 a_n7636_8799.t14 2.82907
R16060 a_n7636_8799.n400 a_n7636_8799.t7 2.82907
R16061 a_n7636_8799.n400 a_n7636_8799.t11 2.82907
R16062 a_n7636_8799.n402 a_n7636_8799.t21 2.82907
R16063 a_n7636_8799.n402 a_n7636_8799.t8 2.82907
R16064 a_n7636_8799.n397 a_n7636_8799.t17 2.82907
R16065 a_n7636_8799.n397 a_n7636_8799.t3 2.82907
R16066 a_n7636_8799.n395 a_n7636_8799.t20 2.82907
R16067 a_n7636_8799.n395 a_n7636_8799.t15 2.82907
R16068 a_n7636_8799.n393 a_n7636_8799.t4 2.82907
R16069 a_n7636_8799.n393 a_n7636_8799.t19 2.82907
R16070 a_n7636_8799.n391 a_n7636_8799.t5 2.82907
R16071 a_n7636_8799.n391 a_n7636_8799.t6 2.82907
R16072 a_n7636_8799.n390 a_n7636_8799.t9 2.82907
R16073 a_n7636_8799.n390 a_n7636_8799.t10 2.82907
R16074 a_n7636_8799.n0 a_n7636_8799.t13 2.82907
R16075 a_n7636_8799.n0 a_n7636_8799.t12 2.82907
R16076 a_n7636_8799.n405 a_n7636_8799.t18 2.82907
R16077 a_n7636_8799.t22 a_n7636_8799.n405 2.82907
R16078 a_n7636_8799.n394 a_n7636_8799.n392 0.444466
R16079 a_n7636_8799.n396 a_n7636_8799.n394 0.444466
R16080 a_n7636_8799.n398 a_n7636_8799.n396 0.444466
R16081 a_n7636_8799.n404 a_n7636_8799.n403 0.444466
R16082 a_n7636_8799.n403 a_n7636_8799.n401 0.444466
R16083 a_n7636_8799.n10 a_n7636_8799.n8 0.358259
R16084 a_n7636_8799.n5 a_n7636_8799.n3 0.358259
R16085 a_n7636_8799.n261 a_n7636_8799.n200 0.189894
R16086 a_n7636_8799.n257 a_n7636_8799.n200 0.189894
R16087 a_n7636_8799.n257 a_n7636_8799.n256 0.189894
R16088 a_n7636_8799.n256 a_n7636_8799.n255 0.189894
R16089 a_n7636_8799.n255 a_n7636_8799.n202 0.189894
R16090 a_n7636_8799.n203 a_n7636_8799.n202 0.189894
R16091 a_n7636_8799.n250 a_n7636_8799.n203 0.189894
R16092 a_n7636_8799.n250 a_n7636_8799.n249 0.189894
R16093 a_n7636_8799.n249 a_n7636_8799.n248 0.189894
R16094 a_n7636_8799.n248 a_n7636_8799.n205 0.189894
R16095 a_n7636_8799.n206 a_n7636_8799.n205 0.189894
R16096 a_n7636_8799.n243 a_n7636_8799.n206 0.189894
R16097 a_n7636_8799.n243 a_n7636_8799.n242 0.189894
R16098 a_n7636_8799.n242 a_n7636_8799.n241 0.189894
R16099 a_n7636_8799.n241 a_n7636_8799.n208 0.189894
R16100 a_n7636_8799.n209 a_n7636_8799.n208 0.189894
R16101 a_n7636_8799.n236 a_n7636_8799.n209 0.189894
R16102 a_n7636_8799.n236 a_n7636_8799.n235 0.189894
R16103 a_n7636_8799.n235 a_n7636_8799.n234 0.189894
R16104 a_n7636_8799.n234 a_n7636_8799.n211 0.189894
R16105 a_n7636_8799.n212 a_n7636_8799.n211 0.189894
R16106 a_n7636_8799.n229 a_n7636_8799.n212 0.189894
R16107 a_n7636_8799.n229 a_n7636_8799.n228 0.189894
R16108 a_n7636_8799.n228 a_n7636_8799.n227 0.189894
R16109 a_n7636_8799.n227 a_n7636_8799.n214 0.189894
R16110 a_n7636_8799.n215 a_n7636_8799.n214 0.189894
R16111 a_n7636_8799.n222 a_n7636_8799.n215 0.189894
R16112 a_n7636_8799.n222 a_n7636_8799.n221 0.189894
R16113 a_n7636_8799.n221 a_n7636_8799.n220 0.189894
R16114 a_n7636_8799.n323 a_n7636_8799.n262 0.189894
R16115 a_n7636_8799.n319 a_n7636_8799.n262 0.189894
R16116 a_n7636_8799.n319 a_n7636_8799.n318 0.189894
R16117 a_n7636_8799.n318 a_n7636_8799.n317 0.189894
R16118 a_n7636_8799.n317 a_n7636_8799.n264 0.189894
R16119 a_n7636_8799.n265 a_n7636_8799.n264 0.189894
R16120 a_n7636_8799.n312 a_n7636_8799.n265 0.189894
R16121 a_n7636_8799.n312 a_n7636_8799.n311 0.189894
R16122 a_n7636_8799.n311 a_n7636_8799.n310 0.189894
R16123 a_n7636_8799.n310 a_n7636_8799.n267 0.189894
R16124 a_n7636_8799.n268 a_n7636_8799.n267 0.189894
R16125 a_n7636_8799.n305 a_n7636_8799.n268 0.189894
R16126 a_n7636_8799.n305 a_n7636_8799.n304 0.189894
R16127 a_n7636_8799.n304 a_n7636_8799.n303 0.189894
R16128 a_n7636_8799.n303 a_n7636_8799.n270 0.189894
R16129 a_n7636_8799.n271 a_n7636_8799.n270 0.189894
R16130 a_n7636_8799.n298 a_n7636_8799.n271 0.189894
R16131 a_n7636_8799.n298 a_n7636_8799.n297 0.189894
R16132 a_n7636_8799.n297 a_n7636_8799.n296 0.189894
R16133 a_n7636_8799.n296 a_n7636_8799.n273 0.189894
R16134 a_n7636_8799.n274 a_n7636_8799.n273 0.189894
R16135 a_n7636_8799.n291 a_n7636_8799.n274 0.189894
R16136 a_n7636_8799.n291 a_n7636_8799.n290 0.189894
R16137 a_n7636_8799.n290 a_n7636_8799.n289 0.189894
R16138 a_n7636_8799.n289 a_n7636_8799.n276 0.189894
R16139 a_n7636_8799.n277 a_n7636_8799.n276 0.189894
R16140 a_n7636_8799.n284 a_n7636_8799.n277 0.189894
R16141 a_n7636_8799.n284 a_n7636_8799.n283 0.189894
R16142 a_n7636_8799.n283 a_n7636_8799.n282 0.189894
R16143 a_n7636_8799.n386 a_n7636_8799.n325 0.189894
R16144 a_n7636_8799.n382 a_n7636_8799.n325 0.189894
R16145 a_n7636_8799.n382 a_n7636_8799.n381 0.189894
R16146 a_n7636_8799.n381 a_n7636_8799.n380 0.189894
R16147 a_n7636_8799.n380 a_n7636_8799.n327 0.189894
R16148 a_n7636_8799.n328 a_n7636_8799.n327 0.189894
R16149 a_n7636_8799.n375 a_n7636_8799.n328 0.189894
R16150 a_n7636_8799.n375 a_n7636_8799.n374 0.189894
R16151 a_n7636_8799.n374 a_n7636_8799.n373 0.189894
R16152 a_n7636_8799.n373 a_n7636_8799.n330 0.189894
R16153 a_n7636_8799.n331 a_n7636_8799.n330 0.189894
R16154 a_n7636_8799.n368 a_n7636_8799.n331 0.189894
R16155 a_n7636_8799.n368 a_n7636_8799.n367 0.189894
R16156 a_n7636_8799.n367 a_n7636_8799.n366 0.189894
R16157 a_n7636_8799.n366 a_n7636_8799.n333 0.189894
R16158 a_n7636_8799.n334 a_n7636_8799.n333 0.189894
R16159 a_n7636_8799.n361 a_n7636_8799.n334 0.189894
R16160 a_n7636_8799.n361 a_n7636_8799.n360 0.189894
R16161 a_n7636_8799.n360 a_n7636_8799.n359 0.189894
R16162 a_n7636_8799.n359 a_n7636_8799.n336 0.189894
R16163 a_n7636_8799.n337 a_n7636_8799.n336 0.189894
R16164 a_n7636_8799.n354 a_n7636_8799.n337 0.189894
R16165 a_n7636_8799.n354 a_n7636_8799.n353 0.189894
R16166 a_n7636_8799.n353 a_n7636_8799.n352 0.189894
R16167 a_n7636_8799.n352 a_n7636_8799.n339 0.189894
R16168 a_n7636_8799.n340 a_n7636_8799.n339 0.189894
R16169 a_n7636_8799.n347 a_n7636_8799.n340 0.189894
R16170 a_n7636_8799.n347 a_n7636_8799.n346 0.189894
R16171 a_n7636_8799.n346 a_n7636_8799.n345 0.189894
R16172 a_n7636_8799.n31 a_n7636_8799.n26 0.189894
R16173 a_n7636_8799.n32 a_n7636_8799.n31 0.189894
R16174 a_n7636_8799.n33 a_n7636_8799.n32 0.189894
R16175 a_n7636_8799.n33 a_n7636_8799.n24 0.189894
R16176 a_n7636_8799.n37 a_n7636_8799.n24 0.189894
R16177 a_n7636_8799.n38 a_n7636_8799.n37 0.189894
R16178 a_n7636_8799.n39 a_n7636_8799.n38 0.189894
R16179 a_n7636_8799.n39 a_n7636_8799.n22 0.189894
R16180 a_n7636_8799.n43 a_n7636_8799.n22 0.189894
R16181 a_n7636_8799.n44 a_n7636_8799.n43 0.189894
R16182 a_n7636_8799.n45 a_n7636_8799.n44 0.189894
R16183 a_n7636_8799.n45 a_n7636_8799.n20 0.189894
R16184 a_n7636_8799.n49 a_n7636_8799.n20 0.189894
R16185 a_n7636_8799.n50 a_n7636_8799.n49 0.189894
R16186 a_n7636_8799.n51 a_n7636_8799.n50 0.189894
R16187 a_n7636_8799.n51 a_n7636_8799.n18 0.189894
R16188 a_n7636_8799.n55 a_n7636_8799.n18 0.189894
R16189 a_n7636_8799.n56 a_n7636_8799.n55 0.189894
R16190 a_n7636_8799.n57 a_n7636_8799.n56 0.189894
R16191 a_n7636_8799.n57 a_n7636_8799.n16 0.189894
R16192 a_n7636_8799.n61 a_n7636_8799.n16 0.189894
R16193 a_n7636_8799.n62 a_n7636_8799.n61 0.189894
R16194 a_n7636_8799.n63 a_n7636_8799.n62 0.189894
R16195 a_n7636_8799.n63 a_n7636_8799.n14 0.189894
R16196 a_n7636_8799.n67 a_n7636_8799.n14 0.189894
R16197 a_n7636_8799.n68 a_n7636_8799.n67 0.189894
R16198 a_n7636_8799.n69 a_n7636_8799.n68 0.189894
R16199 a_n7636_8799.n69 a_n7636_8799.n12 0.189894
R16200 a_n7636_8799.n73 a_n7636_8799.n12 0.189894
R16201 a_n7636_8799.n93 a_n7636_8799.n88 0.189894
R16202 a_n7636_8799.n94 a_n7636_8799.n93 0.189894
R16203 a_n7636_8799.n95 a_n7636_8799.n94 0.189894
R16204 a_n7636_8799.n95 a_n7636_8799.n86 0.189894
R16205 a_n7636_8799.n99 a_n7636_8799.n86 0.189894
R16206 a_n7636_8799.n100 a_n7636_8799.n99 0.189894
R16207 a_n7636_8799.n101 a_n7636_8799.n100 0.189894
R16208 a_n7636_8799.n101 a_n7636_8799.n84 0.189894
R16209 a_n7636_8799.n105 a_n7636_8799.n84 0.189894
R16210 a_n7636_8799.n106 a_n7636_8799.n105 0.189894
R16211 a_n7636_8799.n107 a_n7636_8799.n106 0.189894
R16212 a_n7636_8799.n107 a_n7636_8799.n82 0.189894
R16213 a_n7636_8799.n111 a_n7636_8799.n82 0.189894
R16214 a_n7636_8799.n112 a_n7636_8799.n111 0.189894
R16215 a_n7636_8799.n113 a_n7636_8799.n112 0.189894
R16216 a_n7636_8799.n113 a_n7636_8799.n80 0.189894
R16217 a_n7636_8799.n117 a_n7636_8799.n80 0.189894
R16218 a_n7636_8799.n118 a_n7636_8799.n117 0.189894
R16219 a_n7636_8799.n119 a_n7636_8799.n118 0.189894
R16220 a_n7636_8799.n119 a_n7636_8799.n78 0.189894
R16221 a_n7636_8799.n123 a_n7636_8799.n78 0.189894
R16222 a_n7636_8799.n124 a_n7636_8799.n123 0.189894
R16223 a_n7636_8799.n125 a_n7636_8799.n124 0.189894
R16224 a_n7636_8799.n125 a_n7636_8799.n76 0.189894
R16225 a_n7636_8799.n129 a_n7636_8799.n76 0.189894
R16226 a_n7636_8799.n130 a_n7636_8799.n129 0.189894
R16227 a_n7636_8799.n131 a_n7636_8799.n130 0.189894
R16228 a_n7636_8799.n131 a_n7636_8799.n74 0.189894
R16229 a_n7636_8799.n135 a_n7636_8799.n74 0.189894
R16230 a_n7636_8799.n156 a_n7636_8799.n151 0.189894
R16231 a_n7636_8799.n157 a_n7636_8799.n156 0.189894
R16232 a_n7636_8799.n158 a_n7636_8799.n157 0.189894
R16233 a_n7636_8799.n158 a_n7636_8799.n149 0.189894
R16234 a_n7636_8799.n162 a_n7636_8799.n149 0.189894
R16235 a_n7636_8799.n163 a_n7636_8799.n162 0.189894
R16236 a_n7636_8799.n164 a_n7636_8799.n163 0.189894
R16237 a_n7636_8799.n164 a_n7636_8799.n147 0.189894
R16238 a_n7636_8799.n168 a_n7636_8799.n147 0.189894
R16239 a_n7636_8799.n169 a_n7636_8799.n168 0.189894
R16240 a_n7636_8799.n170 a_n7636_8799.n169 0.189894
R16241 a_n7636_8799.n170 a_n7636_8799.n145 0.189894
R16242 a_n7636_8799.n174 a_n7636_8799.n145 0.189894
R16243 a_n7636_8799.n175 a_n7636_8799.n174 0.189894
R16244 a_n7636_8799.n176 a_n7636_8799.n175 0.189894
R16245 a_n7636_8799.n176 a_n7636_8799.n143 0.189894
R16246 a_n7636_8799.n180 a_n7636_8799.n143 0.189894
R16247 a_n7636_8799.n181 a_n7636_8799.n180 0.189894
R16248 a_n7636_8799.n182 a_n7636_8799.n181 0.189894
R16249 a_n7636_8799.n182 a_n7636_8799.n141 0.189894
R16250 a_n7636_8799.n186 a_n7636_8799.n141 0.189894
R16251 a_n7636_8799.n187 a_n7636_8799.n186 0.189894
R16252 a_n7636_8799.n188 a_n7636_8799.n187 0.189894
R16253 a_n7636_8799.n188 a_n7636_8799.n139 0.189894
R16254 a_n7636_8799.n192 a_n7636_8799.n139 0.189894
R16255 a_n7636_8799.n193 a_n7636_8799.n192 0.189894
R16256 a_n7636_8799.n194 a_n7636_8799.n193 0.189894
R16257 a_n7636_8799.n194 a_n7636_8799.n137 0.189894
R16258 a_n7636_8799.n198 a_n7636_8799.n137 0.189894
R16259 vdd.n327 vdd.n291 756.745
R16260 vdd.n268 vdd.n232 756.745
R16261 vdd.n225 vdd.n189 756.745
R16262 vdd.n166 vdd.n130 756.745
R16263 vdd.n124 vdd.n88 756.745
R16264 vdd.n65 vdd.n29 756.745
R16265 vdd.n1746 vdd.n1710 756.745
R16266 vdd.n1805 vdd.n1769 756.745
R16267 vdd.n1644 vdd.n1608 756.745
R16268 vdd.n1703 vdd.n1667 756.745
R16269 vdd.n1543 vdd.n1507 756.745
R16270 vdd.n1602 vdd.n1566 756.745
R16271 vdd.n2177 vdd.t260 640.208
R16272 vdd.n965 vdd.t245 640.208
R16273 vdd.n2151 vdd.t206 640.208
R16274 vdd.n957 vdd.t270 640.208
R16275 vdd.n2922 vdd.t221 640.208
R16276 vdd.n2642 vdd.t267 640.208
R16277 vdd.n832 vdd.t249 640.208
R16278 vdd.n2639 vdd.t253 640.208
R16279 vdd.n799 vdd.t257 640.208
R16280 vdd.n1027 vdd.t263 640.208
R16281 vdd.n1317 vdd.t236 592.009
R16282 vdd.n1355 vdd.t225 592.009
R16283 vdd.n1251 vdd.t239 592.009
R16284 vdd.n2333 vdd.t217 592.009
R16285 vdd.n1970 vdd.t229 592.009
R16286 vdd.n1930 vdd.t242 592.009
R16287 vdd.n426 vdd.t232 592.009
R16288 vdd.n440 vdd.t273 592.009
R16289 vdd.n452 vdd.t279 592.009
R16290 vdd.n768 vdd.t210 592.009
R16291 vdd.n3184 vdd.t214 592.009
R16292 vdd.n688 vdd.t276 592.009
R16293 vdd.n328 vdd.n327 585
R16294 vdd.n326 vdd.n293 585
R16295 vdd.n325 vdd.n324 585
R16296 vdd.n296 vdd.n294 585
R16297 vdd.n319 vdd.n318 585
R16298 vdd.n317 vdd.n316 585
R16299 vdd.n300 vdd.n299 585
R16300 vdd.n311 vdd.n310 585
R16301 vdd.n309 vdd.n308 585
R16302 vdd.n304 vdd.n303 585
R16303 vdd.n269 vdd.n268 585
R16304 vdd.n267 vdd.n234 585
R16305 vdd.n266 vdd.n265 585
R16306 vdd.n237 vdd.n235 585
R16307 vdd.n260 vdd.n259 585
R16308 vdd.n258 vdd.n257 585
R16309 vdd.n241 vdd.n240 585
R16310 vdd.n252 vdd.n251 585
R16311 vdd.n250 vdd.n249 585
R16312 vdd.n245 vdd.n244 585
R16313 vdd.n226 vdd.n225 585
R16314 vdd.n224 vdd.n191 585
R16315 vdd.n223 vdd.n222 585
R16316 vdd.n194 vdd.n192 585
R16317 vdd.n217 vdd.n216 585
R16318 vdd.n215 vdd.n214 585
R16319 vdd.n198 vdd.n197 585
R16320 vdd.n209 vdd.n208 585
R16321 vdd.n207 vdd.n206 585
R16322 vdd.n202 vdd.n201 585
R16323 vdd.n167 vdd.n166 585
R16324 vdd.n165 vdd.n132 585
R16325 vdd.n164 vdd.n163 585
R16326 vdd.n135 vdd.n133 585
R16327 vdd.n158 vdd.n157 585
R16328 vdd.n156 vdd.n155 585
R16329 vdd.n139 vdd.n138 585
R16330 vdd.n150 vdd.n149 585
R16331 vdd.n148 vdd.n147 585
R16332 vdd.n143 vdd.n142 585
R16333 vdd.n125 vdd.n124 585
R16334 vdd.n123 vdd.n90 585
R16335 vdd.n122 vdd.n121 585
R16336 vdd.n93 vdd.n91 585
R16337 vdd.n116 vdd.n115 585
R16338 vdd.n114 vdd.n113 585
R16339 vdd.n97 vdd.n96 585
R16340 vdd.n108 vdd.n107 585
R16341 vdd.n106 vdd.n105 585
R16342 vdd.n101 vdd.n100 585
R16343 vdd.n66 vdd.n65 585
R16344 vdd.n64 vdd.n31 585
R16345 vdd.n63 vdd.n62 585
R16346 vdd.n34 vdd.n32 585
R16347 vdd.n57 vdd.n56 585
R16348 vdd.n55 vdd.n54 585
R16349 vdd.n38 vdd.n37 585
R16350 vdd.n49 vdd.n48 585
R16351 vdd.n47 vdd.n46 585
R16352 vdd.n42 vdd.n41 585
R16353 vdd.n1747 vdd.n1746 585
R16354 vdd.n1745 vdd.n1712 585
R16355 vdd.n1744 vdd.n1743 585
R16356 vdd.n1715 vdd.n1713 585
R16357 vdd.n1738 vdd.n1737 585
R16358 vdd.n1736 vdd.n1735 585
R16359 vdd.n1719 vdd.n1718 585
R16360 vdd.n1730 vdd.n1729 585
R16361 vdd.n1728 vdd.n1727 585
R16362 vdd.n1723 vdd.n1722 585
R16363 vdd.n1806 vdd.n1805 585
R16364 vdd.n1804 vdd.n1771 585
R16365 vdd.n1803 vdd.n1802 585
R16366 vdd.n1774 vdd.n1772 585
R16367 vdd.n1797 vdd.n1796 585
R16368 vdd.n1795 vdd.n1794 585
R16369 vdd.n1778 vdd.n1777 585
R16370 vdd.n1789 vdd.n1788 585
R16371 vdd.n1787 vdd.n1786 585
R16372 vdd.n1782 vdd.n1781 585
R16373 vdd.n1645 vdd.n1644 585
R16374 vdd.n1643 vdd.n1610 585
R16375 vdd.n1642 vdd.n1641 585
R16376 vdd.n1613 vdd.n1611 585
R16377 vdd.n1636 vdd.n1635 585
R16378 vdd.n1634 vdd.n1633 585
R16379 vdd.n1617 vdd.n1616 585
R16380 vdd.n1628 vdd.n1627 585
R16381 vdd.n1626 vdd.n1625 585
R16382 vdd.n1621 vdd.n1620 585
R16383 vdd.n1704 vdd.n1703 585
R16384 vdd.n1702 vdd.n1669 585
R16385 vdd.n1701 vdd.n1700 585
R16386 vdd.n1672 vdd.n1670 585
R16387 vdd.n1695 vdd.n1694 585
R16388 vdd.n1693 vdd.n1692 585
R16389 vdd.n1676 vdd.n1675 585
R16390 vdd.n1687 vdd.n1686 585
R16391 vdd.n1685 vdd.n1684 585
R16392 vdd.n1680 vdd.n1679 585
R16393 vdd.n1544 vdd.n1543 585
R16394 vdd.n1542 vdd.n1509 585
R16395 vdd.n1541 vdd.n1540 585
R16396 vdd.n1512 vdd.n1510 585
R16397 vdd.n1535 vdd.n1534 585
R16398 vdd.n1533 vdd.n1532 585
R16399 vdd.n1516 vdd.n1515 585
R16400 vdd.n1527 vdd.n1526 585
R16401 vdd.n1525 vdd.n1524 585
R16402 vdd.n1520 vdd.n1519 585
R16403 vdd.n1603 vdd.n1602 585
R16404 vdd.n1601 vdd.n1568 585
R16405 vdd.n1600 vdd.n1599 585
R16406 vdd.n1571 vdd.n1569 585
R16407 vdd.n1594 vdd.n1593 585
R16408 vdd.n1592 vdd.n1591 585
R16409 vdd.n1575 vdd.n1574 585
R16410 vdd.n1586 vdd.n1585 585
R16411 vdd.n1584 vdd.n1583 585
R16412 vdd.n1579 vdd.n1578 585
R16413 vdd.n3356 vdd.n392 509.269
R16414 vdd.n3352 vdd.n393 509.269
R16415 vdd.n3224 vdd.n685 509.269
R16416 vdd.n3221 vdd.n684 509.269
R16417 vdd.n2328 vdd.n1075 509.269
R16418 vdd.n2331 vdd.n2330 509.269
R16419 vdd.n1224 vdd.n1188 509.269
R16420 vdd.n1420 vdd.n1189 509.269
R16421 vdd.n305 vdd.t141 329.043
R16422 vdd.n246 vdd.t115 329.043
R16423 vdd.n203 vdd.t128 329.043
R16424 vdd.n144 vdd.t101 329.043
R16425 vdd.n102 vdd.t80 329.043
R16426 vdd.n43 vdd.t14 329.043
R16427 vdd.n1724 vdd.t160 329.043
R16428 vdd.n1783 vdd.t47 329.043
R16429 vdd.n1622 vdd.t146 329.043
R16430 vdd.n1681 vdd.t22 329.043
R16431 vdd.n1521 vdd.t18 329.043
R16432 vdd.n1580 vdd.t81 329.043
R16433 vdd.n1317 vdd.t238 319.788
R16434 vdd.n1355 vdd.t228 319.788
R16435 vdd.n1251 vdd.t241 319.788
R16436 vdd.n2333 vdd.t219 319.788
R16437 vdd.n1970 vdd.t230 319.788
R16438 vdd.n1930 vdd.t243 319.788
R16439 vdd.n426 vdd.t234 319.788
R16440 vdd.n440 vdd.t274 319.788
R16441 vdd.n452 vdd.t280 319.788
R16442 vdd.n768 vdd.t213 319.788
R16443 vdd.n3184 vdd.t216 319.788
R16444 vdd.n688 vdd.t278 319.788
R16445 vdd.n1318 vdd.t237 303.69
R16446 vdd.n1356 vdd.t227 303.69
R16447 vdd.n1252 vdd.t240 303.69
R16448 vdd.n2334 vdd.t220 303.69
R16449 vdd.n1971 vdd.t231 303.69
R16450 vdd.n1931 vdd.t244 303.69
R16451 vdd.n427 vdd.t235 303.69
R16452 vdd.n441 vdd.t275 303.69
R16453 vdd.n453 vdd.t281 303.69
R16454 vdd.n769 vdd.t212 303.69
R16455 vdd.n3185 vdd.t215 303.69
R16456 vdd.n689 vdd.t277 303.69
R16457 vdd.n2865 vdd.n913 297.074
R16458 vdd.n3058 vdd.n809 297.074
R16459 vdd.n2995 vdd.n806 297.074
R16460 vdd.n2788 vdd.n914 297.074
R16461 vdd.n2603 vdd.n954 297.074
R16462 vdd.n2534 vdd.n2533 297.074
R16463 vdd.n2280 vdd.n1050 297.074
R16464 vdd.n2376 vdd.n1048 297.074
R16465 vdd.n2974 vdd.n807 297.074
R16466 vdd.n3061 vdd.n3060 297.074
R16467 vdd.n2637 vdd.n915 297.074
R16468 vdd.n2863 vdd.n916 297.074
R16469 vdd.n2531 vdd.n963 297.074
R16470 vdd.n961 vdd.n936 297.074
R16471 vdd.n2217 vdd.n1051 297.074
R16472 vdd.n2374 vdd.n1052 297.074
R16473 vdd.n2976 vdd.n807 185
R16474 vdd.n3059 vdd.n807 185
R16475 vdd.n2978 vdd.n2977 185
R16476 vdd.n2977 vdd.n805 185
R16477 vdd.n2979 vdd.n839 185
R16478 vdd.n2989 vdd.n839 185
R16479 vdd.n2980 vdd.n848 185
R16480 vdd.n848 vdd.n846 185
R16481 vdd.n2982 vdd.n2981 185
R16482 vdd.n2983 vdd.n2982 185
R16483 vdd.n2935 vdd.n847 185
R16484 vdd.n847 vdd.n843 185
R16485 vdd.n2934 vdd.n2933 185
R16486 vdd.n2933 vdd.n2932 185
R16487 vdd.n850 vdd.n849 185
R16488 vdd.n851 vdd.n850 185
R16489 vdd.n2925 vdd.n2924 185
R16490 vdd.n2926 vdd.n2925 185
R16491 vdd.n2921 vdd.n860 185
R16492 vdd.n860 vdd.n857 185
R16493 vdd.n2920 vdd.n2919 185
R16494 vdd.n2919 vdd.n2918 185
R16495 vdd.n862 vdd.n861 185
R16496 vdd.n870 vdd.n862 185
R16497 vdd.n2911 vdd.n2910 185
R16498 vdd.n2912 vdd.n2911 185
R16499 vdd.n2909 vdd.n871 185
R16500 vdd.n2760 vdd.n871 185
R16501 vdd.n2908 vdd.n2907 185
R16502 vdd.n2907 vdd.n2906 185
R16503 vdd.n873 vdd.n872 185
R16504 vdd.n874 vdd.n873 185
R16505 vdd.n2899 vdd.n2898 185
R16506 vdd.n2900 vdd.n2899 185
R16507 vdd.n2897 vdd.n883 185
R16508 vdd.n883 vdd.n880 185
R16509 vdd.n2896 vdd.n2895 185
R16510 vdd.n2895 vdd.n2894 185
R16511 vdd.n885 vdd.n884 185
R16512 vdd.n893 vdd.n885 185
R16513 vdd.n2887 vdd.n2886 185
R16514 vdd.n2888 vdd.n2887 185
R16515 vdd.n2885 vdd.n894 185
R16516 vdd.n900 vdd.n894 185
R16517 vdd.n2884 vdd.n2883 185
R16518 vdd.n2883 vdd.n2882 185
R16519 vdd.n896 vdd.n895 185
R16520 vdd.n897 vdd.n896 185
R16521 vdd.n2875 vdd.n2874 185
R16522 vdd.n2876 vdd.n2875 185
R16523 vdd.n2873 vdd.n906 185
R16524 vdd.n2781 vdd.n906 185
R16525 vdd.n2872 vdd.n2871 185
R16526 vdd.n2871 vdd.n2870 185
R16527 vdd.n908 vdd.n907 185
R16528 vdd.t4 vdd.n908 185
R16529 vdd.n2863 vdd.n2862 185
R16530 vdd.n2864 vdd.n2863 185
R16531 vdd.n2861 vdd.n916 185
R16532 vdd.n2860 vdd.n2859 185
R16533 vdd.n918 vdd.n917 185
R16534 vdd.n2646 vdd.n2645 185
R16535 vdd.n2648 vdd.n2647 185
R16536 vdd.n2650 vdd.n2649 185
R16537 vdd.n2652 vdd.n2651 185
R16538 vdd.n2654 vdd.n2653 185
R16539 vdd.n2656 vdd.n2655 185
R16540 vdd.n2658 vdd.n2657 185
R16541 vdd.n2660 vdd.n2659 185
R16542 vdd.n2662 vdd.n2661 185
R16543 vdd.n2664 vdd.n2663 185
R16544 vdd.n2666 vdd.n2665 185
R16545 vdd.n2668 vdd.n2667 185
R16546 vdd.n2670 vdd.n2669 185
R16547 vdd.n2672 vdd.n2671 185
R16548 vdd.n2674 vdd.n2673 185
R16549 vdd.n2676 vdd.n2675 185
R16550 vdd.n2678 vdd.n2677 185
R16551 vdd.n2680 vdd.n2679 185
R16552 vdd.n2682 vdd.n2681 185
R16553 vdd.n2684 vdd.n2683 185
R16554 vdd.n2686 vdd.n2685 185
R16555 vdd.n2688 vdd.n2687 185
R16556 vdd.n2690 vdd.n2689 185
R16557 vdd.n2692 vdd.n2691 185
R16558 vdd.n2694 vdd.n2693 185
R16559 vdd.n2696 vdd.n2695 185
R16560 vdd.n2698 vdd.n2697 185
R16561 vdd.n2700 vdd.n2699 185
R16562 vdd.n2702 vdd.n2701 185
R16563 vdd.n2704 vdd.n2703 185
R16564 vdd.n2706 vdd.n2705 185
R16565 vdd.n2707 vdd.n2637 185
R16566 vdd.n2857 vdd.n2637 185
R16567 vdd.n3062 vdd.n3061 185
R16568 vdd.n3063 vdd.n798 185
R16569 vdd.n3065 vdd.n3064 185
R16570 vdd.n3067 vdd.n796 185
R16571 vdd.n3069 vdd.n3068 185
R16572 vdd.n3070 vdd.n795 185
R16573 vdd.n3072 vdd.n3071 185
R16574 vdd.n3074 vdd.n793 185
R16575 vdd.n3076 vdd.n3075 185
R16576 vdd.n3077 vdd.n792 185
R16577 vdd.n3079 vdd.n3078 185
R16578 vdd.n3081 vdd.n790 185
R16579 vdd.n3083 vdd.n3082 185
R16580 vdd.n3084 vdd.n789 185
R16581 vdd.n3086 vdd.n3085 185
R16582 vdd.n3088 vdd.n788 185
R16583 vdd.n3089 vdd.n786 185
R16584 vdd.n3092 vdd.n3091 185
R16585 vdd.n787 vdd.n785 185
R16586 vdd.n2948 vdd.n2947 185
R16587 vdd.n2950 vdd.n2949 185
R16588 vdd.n2952 vdd.n2944 185
R16589 vdd.n2954 vdd.n2953 185
R16590 vdd.n2955 vdd.n2943 185
R16591 vdd.n2957 vdd.n2956 185
R16592 vdd.n2959 vdd.n2941 185
R16593 vdd.n2961 vdd.n2960 185
R16594 vdd.n2962 vdd.n2940 185
R16595 vdd.n2964 vdd.n2963 185
R16596 vdd.n2966 vdd.n2938 185
R16597 vdd.n2968 vdd.n2967 185
R16598 vdd.n2969 vdd.n2937 185
R16599 vdd.n2971 vdd.n2970 185
R16600 vdd.n2973 vdd.n2936 185
R16601 vdd.n2975 vdd.n2974 185
R16602 vdd.n2974 vdd.n692 185
R16603 vdd.n3060 vdd.n802 185
R16604 vdd.n3060 vdd.n3059 185
R16605 vdd.n2712 vdd.n804 185
R16606 vdd.n805 vdd.n804 185
R16607 vdd.n2713 vdd.n838 185
R16608 vdd.n2989 vdd.n838 185
R16609 vdd.n2715 vdd.n2714 185
R16610 vdd.n2714 vdd.n846 185
R16611 vdd.n2716 vdd.n845 185
R16612 vdd.n2983 vdd.n845 185
R16613 vdd.n2718 vdd.n2717 185
R16614 vdd.n2717 vdd.n843 185
R16615 vdd.n2719 vdd.n853 185
R16616 vdd.n2932 vdd.n853 185
R16617 vdd.n2721 vdd.n2720 185
R16618 vdd.n2720 vdd.n851 185
R16619 vdd.n2722 vdd.n859 185
R16620 vdd.n2926 vdd.n859 185
R16621 vdd.n2724 vdd.n2723 185
R16622 vdd.n2723 vdd.n857 185
R16623 vdd.n2725 vdd.n864 185
R16624 vdd.n2918 vdd.n864 185
R16625 vdd.n2727 vdd.n2726 185
R16626 vdd.n2726 vdd.n870 185
R16627 vdd.n2728 vdd.n869 185
R16628 vdd.n2912 vdd.n869 185
R16629 vdd.n2762 vdd.n2761 185
R16630 vdd.n2761 vdd.n2760 185
R16631 vdd.n2763 vdd.n876 185
R16632 vdd.n2906 vdd.n876 185
R16633 vdd.n2765 vdd.n2764 185
R16634 vdd.n2764 vdd.n874 185
R16635 vdd.n2766 vdd.n882 185
R16636 vdd.n2900 vdd.n882 185
R16637 vdd.n2768 vdd.n2767 185
R16638 vdd.n2767 vdd.n880 185
R16639 vdd.n2769 vdd.n887 185
R16640 vdd.n2894 vdd.n887 185
R16641 vdd.n2771 vdd.n2770 185
R16642 vdd.n2770 vdd.n893 185
R16643 vdd.n2772 vdd.n892 185
R16644 vdd.n2888 vdd.n892 185
R16645 vdd.n2774 vdd.n2773 185
R16646 vdd.n2773 vdd.n900 185
R16647 vdd.n2775 vdd.n899 185
R16648 vdd.n2882 vdd.n899 185
R16649 vdd.n2777 vdd.n2776 185
R16650 vdd.n2776 vdd.n897 185
R16651 vdd.n2778 vdd.n905 185
R16652 vdd.n2876 vdd.n905 185
R16653 vdd.n2780 vdd.n2779 185
R16654 vdd.n2781 vdd.n2780 185
R16655 vdd.n2711 vdd.n910 185
R16656 vdd.n2870 vdd.n910 185
R16657 vdd.n2710 vdd.n2709 185
R16658 vdd.n2709 vdd.t4 185
R16659 vdd.n2708 vdd.n915 185
R16660 vdd.n2864 vdd.n915 185
R16661 vdd.n2328 vdd.n2327 185
R16662 vdd.n2329 vdd.n2328 185
R16663 vdd.n1076 vdd.n1074 185
R16664 vdd.n1894 vdd.n1074 185
R16665 vdd.n1897 vdd.n1896 185
R16666 vdd.n1896 vdd.n1895 185
R16667 vdd.n1079 vdd.n1078 185
R16668 vdd.n1080 vdd.n1079 185
R16669 vdd.n1883 vdd.n1882 185
R16670 vdd.n1884 vdd.n1883 185
R16671 vdd.n1088 vdd.n1087 185
R16672 vdd.n1875 vdd.n1087 185
R16673 vdd.n1878 vdd.n1877 185
R16674 vdd.n1877 vdd.n1876 185
R16675 vdd.n1091 vdd.n1090 185
R16676 vdd.n1098 vdd.n1091 185
R16677 vdd.n1866 vdd.n1865 185
R16678 vdd.n1867 vdd.n1866 185
R16679 vdd.n1100 vdd.n1099 185
R16680 vdd.n1099 vdd.n1097 185
R16681 vdd.n1861 vdd.n1860 185
R16682 vdd.n1860 vdd.n1859 185
R16683 vdd.n1103 vdd.n1102 185
R16684 vdd.n1104 vdd.n1103 185
R16685 vdd.n1850 vdd.n1849 185
R16686 vdd.n1851 vdd.n1850 185
R16687 vdd.n1111 vdd.n1110 185
R16688 vdd.n1842 vdd.n1110 185
R16689 vdd.n1845 vdd.n1844 185
R16690 vdd.n1844 vdd.n1843 185
R16691 vdd.n1114 vdd.n1113 185
R16692 vdd.n1120 vdd.n1114 185
R16693 vdd.n1833 vdd.n1832 185
R16694 vdd.n1834 vdd.n1833 185
R16695 vdd.n1122 vdd.n1121 185
R16696 vdd.n1825 vdd.n1121 185
R16697 vdd.n1828 vdd.n1827 185
R16698 vdd.n1827 vdd.n1826 185
R16699 vdd.n1125 vdd.n1124 185
R16700 vdd.n1126 vdd.n1125 185
R16701 vdd.n1816 vdd.n1815 185
R16702 vdd.n1817 vdd.n1816 185
R16703 vdd.n1134 vdd.n1133 185
R16704 vdd.n1133 vdd.n1132 185
R16705 vdd.n1504 vdd.n1503 185
R16706 vdd.n1503 vdd.n1502 185
R16707 vdd.n1137 vdd.n1136 185
R16708 vdd.n1143 vdd.n1137 185
R16709 vdd.n1493 vdd.n1492 185
R16710 vdd.n1494 vdd.n1493 185
R16711 vdd.n1145 vdd.n1144 185
R16712 vdd.n1485 vdd.n1144 185
R16713 vdd.n1488 vdd.n1487 185
R16714 vdd.n1487 vdd.n1486 185
R16715 vdd.n1148 vdd.n1147 185
R16716 vdd.n1155 vdd.n1148 185
R16717 vdd.n1476 vdd.n1475 185
R16718 vdd.n1477 vdd.n1476 185
R16719 vdd.n1157 vdd.n1156 185
R16720 vdd.n1156 vdd.n1154 185
R16721 vdd.n1471 vdd.n1470 185
R16722 vdd.n1470 vdd.n1469 185
R16723 vdd.n1160 vdd.n1159 185
R16724 vdd.n1161 vdd.n1160 185
R16725 vdd.n1460 vdd.n1459 185
R16726 vdd.n1461 vdd.n1460 185
R16727 vdd.n1168 vdd.n1167 185
R16728 vdd.n1452 vdd.n1167 185
R16729 vdd.n1455 vdd.n1454 185
R16730 vdd.n1454 vdd.n1453 185
R16731 vdd.n1171 vdd.n1170 185
R16732 vdd.n1177 vdd.n1171 185
R16733 vdd.n1443 vdd.n1442 185
R16734 vdd.n1444 vdd.n1443 185
R16735 vdd.n1179 vdd.n1178 185
R16736 vdd.n1435 vdd.n1178 185
R16737 vdd.n1438 vdd.n1437 185
R16738 vdd.n1437 vdd.n1436 185
R16739 vdd.n1182 vdd.n1181 185
R16740 vdd.n1183 vdd.n1182 185
R16741 vdd.n1426 vdd.n1425 185
R16742 vdd.n1427 vdd.n1426 185
R16743 vdd.n1190 vdd.n1189 185
R16744 vdd.n1225 vdd.n1189 185
R16745 vdd.n1421 vdd.n1420 185
R16746 vdd.n1193 vdd.n1192 185
R16747 vdd.n1417 vdd.n1416 185
R16748 vdd.n1418 vdd.n1417 185
R16749 vdd.n1227 vdd.n1226 185
R16750 vdd.n1412 vdd.n1229 185
R16751 vdd.n1411 vdd.n1230 185
R16752 vdd.n1410 vdd.n1231 185
R16753 vdd.n1233 vdd.n1232 185
R16754 vdd.n1406 vdd.n1235 185
R16755 vdd.n1405 vdd.n1236 185
R16756 vdd.n1404 vdd.n1237 185
R16757 vdd.n1239 vdd.n1238 185
R16758 vdd.n1400 vdd.n1241 185
R16759 vdd.n1399 vdd.n1242 185
R16760 vdd.n1398 vdd.n1243 185
R16761 vdd.n1245 vdd.n1244 185
R16762 vdd.n1394 vdd.n1247 185
R16763 vdd.n1393 vdd.n1248 185
R16764 vdd.n1392 vdd.n1249 185
R16765 vdd.n1253 vdd.n1250 185
R16766 vdd.n1388 vdd.n1255 185
R16767 vdd.n1387 vdd.n1256 185
R16768 vdd.n1386 vdd.n1257 185
R16769 vdd.n1259 vdd.n1258 185
R16770 vdd.n1382 vdd.n1261 185
R16771 vdd.n1381 vdd.n1262 185
R16772 vdd.n1380 vdd.n1263 185
R16773 vdd.n1265 vdd.n1264 185
R16774 vdd.n1376 vdd.n1267 185
R16775 vdd.n1375 vdd.n1268 185
R16776 vdd.n1374 vdd.n1269 185
R16777 vdd.n1271 vdd.n1270 185
R16778 vdd.n1370 vdd.n1273 185
R16779 vdd.n1369 vdd.n1274 185
R16780 vdd.n1368 vdd.n1275 185
R16781 vdd.n1277 vdd.n1276 185
R16782 vdd.n1364 vdd.n1279 185
R16783 vdd.n1363 vdd.n1280 185
R16784 vdd.n1362 vdd.n1281 185
R16785 vdd.n1283 vdd.n1282 185
R16786 vdd.n1358 vdd.n1285 185
R16787 vdd.n1357 vdd.n1354 185
R16788 vdd.n1353 vdd.n1286 185
R16789 vdd.n1288 vdd.n1287 185
R16790 vdd.n1349 vdd.n1290 185
R16791 vdd.n1348 vdd.n1291 185
R16792 vdd.n1347 vdd.n1292 185
R16793 vdd.n1294 vdd.n1293 185
R16794 vdd.n1343 vdd.n1296 185
R16795 vdd.n1342 vdd.n1297 185
R16796 vdd.n1341 vdd.n1298 185
R16797 vdd.n1300 vdd.n1299 185
R16798 vdd.n1337 vdd.n1302 185
R16799 vdd.n1336 vdd.n1303 185
R16800 vdd.n1335 vdd.n1304 185
R16801 vdd.n1306 vdd.n1305 185
R16802 vdd.n1331 vdd.n1308 185
R16803 vdd.n1330 vdd.n1309 185
R16804 vdd.n1329 vdd.n1310 185
R16805 vdd.n1312 vdd.n1311 185
R16806 vdd.n1325 vdd.n1314 185
R16807 vdd.n1324 vdd.n1315 185
R16808 vdd.n1323 vdd.n1316 185
R16809 vdd.n1320 vdd.n1224 185
R16810 vdd.n1418 vdd.n1224 185
R16811 vdd.n2332 vdd.n2331 185
R16812 vdd.n2336 vdd.n1069 185
R16813 vdd.n1999 vdd.n1068 185
R16814 vdd.n2002 vdd.n2001 185
R16815 vdd.n2004 vdd.n2003 185
R16816 vdd.n2007 vdd.n2006 185
R16817 vdd.n2009 vdd.n2008 185
R16818 vdd.n2011 vdd.n1997 185
R16819 vdd.n2013 vdd.n2012 185
R16820 vdd.n2014 vdd.n1991 185
R16821 vdd.n2016 vdd.n2015 185
R16822 vdd.n2018 vdd.n1989 185
R16823 vdd.n2020 vdd.n2019 185
R16824 vdd.n2021 vdd.n1984 185
R16825 vdd.n2023 vdd.n2022 185
R16826 vdd.n2025 vdd.n1982 185
R16827 vdd.n2027 vdd.n2026 185
R16828 vdd.n2028 vdd.n1978 185
R16829 vdd.n2030 vdd.n2029 185
R16830 vdd.n2032 vdd.n1975 185
R16831 vdd.n2034 vdd.n2033 185
R16832 vdd.n1976 vdd.n1969 185
R16833 vdd.n2038 vdd.n1973 185
R16834 vdd.n2039 vdd.n1965 185
R16835 vdd.n2041 vdd.n2040 185
R16836 vdd.n2043 vdd.n1963 185
R16837 vdd.n2045 vdd.n2044 185
R16838 vdd.n2046 vdd.n1958 185
R16839 vdd.n2048 vdd.n2047 185
R16840 vdd.n2050 vdd.n1956 185
R16841 vdd.n2052 vdd.n2051 185
R16842 vdd.n2053 vdd.n1951 185
R16843 vdd.n2055 vdd.n2054 185
R16844 vdd.n2057 vdd.n1949 185
R16845 vdd.n2059 vdd.n2058 185
R16846 vdd.n2060 vdd.n1944 185
R16847 vdd.n2062 vdd.n2061 185
R16848 vdd.n2064 vdd.n1942 185
R16849 vdd.n2066 vdd.n2065 185
R16850 vdd.n2067 vdd.n1938 185
R16851 vdd.n2069 vdd.n2068 185
R16852 vdd.n2071 vdd.n1935 185
R16853 vdd.n2073 vdd.n2072 185
R16854 vdd.n1936 vdd.n1929 185
R16855 vdd.n2077 vdd.n1933 185
R16856 vdd.n2078 vdd.n1925 185
R16857 vdd.n2080 vdd.n2079 185
R16858 vdd.n2082 vdd.n1923 185
R16859 vdd.n2084 vdd.n2083 185
R16860 vdd.n2085 vdd.n1918 185
R16861 vdd.n2087 vdd.n2086 185
R16862 vdd.n2089 vdd.n1916 185
R16863 vdd.n2091 vdd.n2090 185
R16864 vdd.n2092 vdd.n1911 185
R16865 vdd.n2094 vdd.n2093 185
R16866 vdd.n2096 vdd.n1910 185
R16867 vdd.n2097 vdd.n1907 185
R16868 vdd.n2100 vdd.n2099 185
R16869 vdd.n1909 vdd.n1905 185
R16870 vdd.n2317 vdd.n1903 185
R16871 vdd.n2319 vdd.n2318 185
R16872 vdd.n2321 vdd.n1901 185
R16873 vdd.n2323 vdd.n2322 185
R16874 vdd.n2324 vdd.n1075 185
R16875 vdd.n2330 vdd.n1072 185
R16876 vdd.n2330 vdd.n2329 185
R16877 vdd.n1083 vdd.n1071 185
R16878 vdd.n1894 vdd.n1071 185
R16879 vdd.n1893 vdd.n1892 185
R16880 vdd.n1895 vdd.n1893 185
R16881 vdd.n1082 vdd.n1081 185
R16882 vdd.n1081 vdd.n1080 185
R16883 vdd.n1886 vdd.n1885 185
R16884 vdd.n1885 vdd.n1884 185
R16885 vdd.n1086 vdd.n1085 185
R16886 vdd.n1875 vdd.n1086 185
R16887 vdd.n1874 vdd.n1873 185
R16888 vdd.n1876 vdd.n1874 185
R16889 vdd.n1093 vdd.n1092 185
R16890 vdd.n1098 vdd.n1092 185
R16891 vdd.n1869 vdd.n1868 185
R16892 vdd.n1868 vdd.n1867 185
R16893 vdd.n1096 vdd.n1095 185
R16894 vdd.n1097 vdd.n1096 185
R16895 vdd.n1858 vdd.n1857 185
R16896 vdd.n1859 vdd.n1858 185
R16897 vdd.n1106 vdd.n1105 185
R16898 vdd.n1105 vdd.n1104 185
R16899 vdd.n1853 vdd.n1852 185
R16900 vdd.n1852 vdd.n1851 185
R16901 vdd.n1109 vdd.n1108 185
R16902 vdd.n1842 vdd.n1109 185
R16903 vdd.n1841 vdd.n1840 185
R16904 vdd.n1843 vdd.n1841 185
R16905 vdd.n1116 vdd.n1115 185
R16906 vdd.n1120 vdd.n1115 185
R16907 vdd.n1836 vdd.n1835 185
R16908 vdd.n1835 vdd.n1834 185
R16909 vdd.n1119 vdd.n1118 185
R16910 vdd.n1825 vdd.n1119 185
R16911 vdd.n1824 vdd.n1823 185
R16912 vdd.n1826 vdd.n1824 185
R16913 vdd.n1128 vdd.n1127 185
R16914 vdd.n1127 vdd.n1126 185
R16915 vdd.n1819 vdd.n1818 185
R16916 vdd.n1818 vdd.n1817 185
R16917 vdd.n1131 vdd.n1130 185
R16918 vdd.n1132 vdd.n1131 185
R16919 vdd.n1501 vdd.n1500 185
R16920 vdd.n1502 vdd.n1501 185
R16921 vdd.n1139 vdd.n1138 185
R16922 vdd.n1143 vdd.n1138 185
R16923 vdd.n1496 vdd.n1495 185
R16924 vdd.n1495 vdd.n1494 185
R16925 vdd.n1142 vdd.n1141 185
R16926 vdd.n1485 vdd.n1142 185
R16927 vdd.n1484 vdd.n1483 185
R16928 vdd.n1486 vdd.n1484 185
R16929 vdd.n1150 vdd.n1149 185
R16930 vdd.n1155 vdd.n1149 185
R16931 vdd.n1479 vdd.n1478 185
R16932 vdd.n1478 vdd.n1477 185
R16933 vdd.n1153 vdd.n1152 185
R16934 vdd.n1154 vdd.n1153 185
R16935 vdd.n1468 vdd.n1467 185
R16936 vdd.n1469 vdd.n1468 185
R16937 vdd.n1163 vdd.n1162 185
R16938 vdd.n1162 vdd.n1161 185
R16939 vdd.n1463 vdd.n1462 185
R16940 vdd.n1462 vdd.n1461 185
R16941 vdd.n1166 vdd.n1165 185
R16942 vdd.n1452 vdd.n1166 185
R16943 vdd.n1451 vdd.n1450 185
R16944 vdd.n1453 vdd.n1451 185
R16945 vdd.n1173 vdd.n1172 185
R16946 vdd.n1177 vdd.n1172 185
R16947 vdd.n1446 vdd.n1445 185
R16948 vdd.n1445 vdd.n1444 185
R16949 vdd.n1176 vdd.n1175 185
R16950 vdd.n1435 vdd.n1176 185
R16951 vdd.n1434 vdd.n1433 185
R16952 vdd.n1436 vdd.n1434 185
R16953 vdd.n1185 vdd.n1184 185
R16954 vdd.n1184 vdd.n1183 185
R16955 vdd.n1429 vdd.n1428 185
R16956 vdd.n1428 vdd.n1427 185
R16957 vdd.n1188 vdd.n1187 185
R16958 vdd.n1225 vdd.n1188 185
R16959 vdd.n956 vdd.n954 185
R16960 vdd.n2532 vdd.n954 185
R16961 vdd.n2454 vdd.n973 185
R16962 vdd.n973 vdd.t172 185
R16963 vdd.n2456 vdd.n2455 185
R16964 vdd.n2457 vdd.n2456 185
R16965 vdd.n2453 vdd.n972 185
R16966 vdd.n2156 vdd.n972 185
R16967 vdd.n2452 vdd.n2451 185
R16968 vdd.n2451 vdd.n2450 185
R16969 vdd.n975 vdd.n974 185
R16970 vdd.n976 vdd.n975 185
R16971 vdd.n2441 vdd.n2440 185
R16972 vdd.n2442 vdd.n2441 185
R16973 vdd.n2439 vdd.n986 185
R16974 vdd.n986 vdd.n983 185
R16975 vdd.n2438 vdd.n2437 185
R16976 vdd.n2437 vdd.n2436 185
R16977 vdd.n988 vdd.n987 185
R16978 vdd.n989 vdd.n988 185
R16979 vdd.n2429 vdd.n2428 185
R16980 vdd.n2430 vdd.n2429 185
R16981 vdd.n2427 vdd.n997 185
R16982 vdd.n1002 vdd.n997 185
R16983 vdd.n2426 vdd.n2425 185
R16984 vdd.n2425 vdd.n2424 185
R16985 vdd.n999 vdd.n998 185
R16986 vdd.n1008 vdd.n999 185
R16987 vdd.n2417 vdd.n2416 185
R16988 vdd.n2418 vdd.n2417 185
R16989 vdd.n2415 vdd.n1009 185
R16990 vdd.n2257 vdd.n1009 185
R16991 vdd.n2414 vdd.n2413 185
R16992 vdd.n2413 vdd.n2412 185
R16993 vdd.n1011 vdd.n1010 185
R16994 vdd.n1012 vdd.n1011 185
R16995 vdd.n2405 vdd.n2404 185
R16996 vdd.n2406 vdd.n2405 185
R16997 vdd.n2403 vdd.n1021 185
R16998 vdd.n1021 vdd.n1018 185
R16999 vdd.n2402 vdd.n2401 185
R17000 vdd.n2401 vdd.n2400 185
R17001 vdd.n1023 vdd.n1022 185
R17002 vdd.n1033 vdd.n1023 185
R17003 vdd.n2392 vdd.n2391 185
R17004 vdd.n2393 vdd.n2392 185
R17005 vdd.n2390 vdd.n1034 185
R17006 vdd.n1034 vdd.n1030 185
R17007 vdd.n2389 vdd.n2388 185
R17008 vdd.n2388 vdd.n2387 185
R17009 vdd.n1036 vdd.n1035 185
R17010 vdd.n1037 vdd.n1036 185
R17011 vdd.n2380 vdd.n2379 185
R17012 vdd.n2381 vdd.n2380 185
R17013 vdd.n2378 vdd.n1046 185
R17014 vdd.n1046 vdd.n1043 185
R17015 vdd.n2377 vdd.n2376 185
R17016 vdd.n2376 vdd.n2375 185
R17017 vdd.n1048 vdd.n1047 185
R17018 vdd.n2112 vdd.n2111 185
R17019 vdd.n2113 vdd.n2109 185
R17020 vdd.n2109 vdd.n1049 185
R17021 vdd.n2115 vdd.n2114 185
R17022 vdd.n2117 vdd.n2108 185
R17023 vdd.n2120 vdd.n2119 185
R17024 vdd.n2121 vdd.n2107 185
R17025 vdd.n2123 vdd.n2122 185
R17026 vdd.n2125 vdd.n2106 185
R17027 vdd.n2128 vdd.n2127 185
R17028 vdd.n2129 vdd.n2105 185
R17029 vdd.n2131 vdd.n2130 185
R17030 vdd.n2133 vdd.n2104 185
R17031 vdd.n2136 vdd.n2135 185
R17032 vdd.n2137 vdd.n2103 185
R17033 vdd.n2139 vdd.n2138 185
R17034 vdd.n2141 vdd.n2102 185
R17035 vdd.n2314 vdd.n2142 185
R17036 vdd.n2313 vdd.n2312 185
R17037 vdd.n2310 vdd.n2143 185
R17038 vdd.n2308 vdd.n2307 185
R17039 vdd.n2306 vdd.n2144 185
R17040 vdd.n2305 vdd.n2304 185
R17041 vdd.n2302 vdd.n2145 185
R17042 vdd.n2300 vdd.n2299 185
R17043 vdd.n2298 vdd.n2146 185
R17044 vdd.n2297 vdd.n2296 185
R17045 vdd.n2294 vdd.n2147 185
R17046 vdd.n2292 vdd.n2291 185
R17047 vdd.n2290 vdd.n2148 185
R17048 vdd.n2289 vdd.n2288 185
R17049 vdd.n2286 vdd.n2149 185
R17050 vdd.n2284 vdd.n2283 185
R17051 vdd.n2282 vdd.n2150 185
R17052 vdd.n2281 vdd.n2280 185
R17053 vdd.n2535 vdd.n2534 185
R17054 vdd.n2537 vdd.n2536 185
R17055 vdd.n2539 vdd.n2538 185
R17056 vdd.n2542 vdd.n2541 185
R17057 vdd.n2544 vdd.n2543 185
R17058 vdd.n2546 vdd.n2545 185
R17059 vdd.n2548 vdd.n2547 185
R17060 vdd.n2550 vdd.n2549 185
R17061 vdd.n2552 vdd.n2551 185
R17062 vdd.n2554 vdd.n2553 185
R17063 vdd.n2556 vdd.n2555 185
R17064 vdd.n2558 vdd.n2557 185
R17065 vdd.n2560 vdd.n2559 185
R17066 vdd.n2562 vdd.n2561 185
R17067 vdd.n2564 vdd.n2563 185
R17068 vdd.n2566 vdd.n2565 185
R17069 vdd.n2568 vdd.n2567 185
R17070 vdd.n2570 vdd.n2569 185
R17071 vdd.n2572 vdd.n2571 185
R17072 vdd.n2574 vdd.n2573 185
R17073 vdd.n2576 vdd.n2575 185
R17074 vdd.n2578 vdd.n2577 185
R17075 vdd.n2580 vdd.n2579 185
R17076 vdd.n2582 vdd.n2581 185
R17077 vdd.n2584 vdd.n2583 185
R17078 vdd.n2586 vdd.n2585 185
R17079 vdd.n2588 vdd.n2587 185
R17080 vdd.n2590 vdd.n2589 185
R17081 vdd.n2592 vdd.n2591 185
R17082 vdd.n2594 vdd.n2593 185
R17083 vdd.n2596 vdd.n2595 185
R17084 vdd.n2598 vdd.n2597 185
R17085 vdd.n2600 vdd.n2599 185
R17086 vdd.n2601 vdd.n955 185
R17087 vdd.n2603 vdd.n2602 185
R17088 vdd.n2604 vdd.n2603 185
R17089 vdd.n2533 vdd.n959 185
R17090 vdd.n2533 vdd.n2532 185
R17091 vdd.n2154 vdd.n960 185
R17092 vdd.t172 vdd.n960 185
R17093 vdd.n2155 vdd.n970 185
R17094 vdd.n2457 vdd.n970 185
R17095 vdd.n2158 vdd.n2157 185
R17096 vdd.n2157 vdd.n2156 185
R17097 vdd.n2159 vdd.n977 185
R17098 vdd.n2450 vdd.n977 185
R17099 vdd.n2161 vdd.n2160 185
R17100 vdd.n2160 vdd.n976 185
R17101 vdd.n2162 vdd.n984 185
R17102 vdd.n2442 vdd.n984 185
R17103 vdd.n2164 vdd.n2163 185
R17104 vdd.n2163 vdd.n983 185
R17105 vdd.n2165 vdd.n990 185
R17106 vdd.n2436 vdd.n990 185
R17107 vdd.n2167 vdd.n2166 185
R17108 vdd.n2166 vdd.n989 185
R17109 vdd.n2168 vdd.n995 185
R17110 vdd.n2430 vdd.n995 185
R17111 vdd.n2170 vdd.n2169 185
R17112 vdd.n2169 vdd.n1002 185
R17113 vdd.n2171 vdd.n1000 185
R17114 vdd.n2424 vdd.n1000 185
R17115 vdd.n2173 vdd.n2172 185
R17116 vdd.n2172 vdd.n1008 185
R17117 vdd.n2174 vdd.n1006 185
R17118 vdd.n2418 vdd.n1006 185
R17119 vdd.n2259 vdd.n2258 185
R17120 vdd.n2258 vdd.n2257 185
R17121 vdd.n2260 vdd.n1013 185
R17122 vdd.n2412 vdd.n1013 185
R17123 vdd.n2262 vdd.n2261 185
R17124 vdd.n2261 vdd.n1012 185
R17125 vdd.n2263 vdd.n1019 185
R17126 vdd.n2406 vdd.n1019 185
R17127 vdd.n2265 vdd.n2264 185
R17128 vdd.n2264 vdd.n1018 185
R17129 vdd.n2266 vdd.n1024 185
R17130 vdd.n2400 vdd.n1024 185
R17131 vdd.n2268 vdd.n2267 185
R17132 vdd.n2267 vdd.n1033 185
R17133 vdd.n2269 vdd.n1031 185
R17134 vdd.n2393 vdd.n1031 185
R17135 vdd.n2271 vdd.n2270 185
R17136 vdd.n2270 vdd.n1030 185
R17137 vdd.n2272 vdd.n1038 185
R17138 vdd.n2387 vdd.n1038 185
R17139 vdd.n2274 vdd.n2273 185
R17140 vdd.n2273 vdd.n1037 185
R17141 vdd.n2275 vdd.n1044 185
R17142 vdd.n2381 vdd.n1044 185
R17143 vdd.n2277 vdd.n2276 185
R17144 vdd.n2276 vdd.n1043 185
R17145 vdd.n2278 vdd.n1050 185
R17146 vdd.n2375 vdd.n1050 185
R17147 vdd.n3357 vdd.n3356 185
R17148 vdd.n3356 vdd.n3355 185
R17149 vdd.n3358 vdd.n387 185
R17150 vdd.n387 vdd.n386 185
R17151 vdd.n3360 vdd.n3359 185
R17152 vdd.n3361 vdd.n3360 185
R17153 vdd.n382 vdd.n381 185
R17154 vdd.n3362 vdd.n382 185
R17155 vdd.n3365 vdd.n3364 185
R17156 vdd.n3364 vdd.n3363 185
R17157 vdd.n3366 vdd.n376 185
R17158 vdd.n376 vdd.n375 185
R17159 vdd.n3368 vdd.n3367 185
R17160 vdd.n3369 vdd.n3368 185
R17161 vdd.n371 vdd.n370 185
R17162 vdd.n3370 vdd.n371 185
R17163 vdd.n3373 vdd.n3372 185
R17164 vdd.n3372 vdd.n3371 185
R17165 vdd.n3374 vdd.n365 185
R17166 vdd.n3331 vdd.n365 185
R17167 vdd.n3376 vdd.n3375 185
R17168 vdd.n3377 vdd.n3376 185
R17169 vdd.n360 vdd.n359 185
R17170 vdd.n3378 vdd.n360 185
R17171 vdd.n3381 vdd.n3380 185
R17172 vdd.n3380 vdd.n3379 185
R17173 vdd.n3382 vdd.n354 185
R17174 vdd.n361 vdd.n354 185
R17175 vdd.n3384 vdd.n3383 185
R17176 vdd.n3385 vdd.n3384 185
R17177 vdd.n350 vdd.n349 185
R17178 vdd.n3386 vdd.n350 185
R17179 vdd.n3389 vdd.n3388 185
R17180 vdd.n3388 vdd.n3387 185
R17181 vdd.n3390 vdd.n345 185
R17182 vdd.n345 vdd.n344 185
R17183 vdd.n3392 vdd.n3391 185
R17184 vdd.n3393 vdd.n3392 185
R17185 vdd.n339 vdd.n337 185
R17186 vdd.n3394 vdd.n339 185
R17187 vdd.n3397 vdd.n3396 185
R17188 vdd.n3396 vdd.n3395 185
R17189 vdd.n338 vdd.n336 185
R17190 vdd.n340 vdd.n338 185
R17191 vdd.n3307 vdd.n3306 185
R17192 vdd.n3308 vdd.n3307 185
R17193 vdd.n635 vdd.n634 185
R17194 vdd.n634 vdd.n633 185
R17195 vdd.n3302 vdd.n3301 185
R17196 vdd.n3301 vdd.n3300 185
R17197 vdd.n638 vdd.n637 185
R17198 vdd.n644 vdd.n638 185
R17199 vdd.n3288 vdd.n3287 185
R17200 vdd.n3289 vdd.n3288 185
R17201 vdd.n646 vdd.n645 185
R17202 vdd.n3280 vdd.n645 185
R17203 vdd.n3283 vdd.n3282 185
R17204 vdd.n3282 vdd.n3281 185
R17205 vdd.n649 vdd.n648 185
R17206 vdd.n656 vdd.n649 185
R17207 vdd.n3271 vdd.n3270 185
R17208 vdd.n3272 vdd.n3271 185
R17209 vdd.n658 vdd.n657 185
R17210 vdd.n657 vdd.n655 185
R17211 vdd.n3266 vdd.n3265 185
R17212 vdd.n3265 vdd.n3264 185
R17213 vdd.n661 vdd.n660 185
R17214 vdd.n662 vdd.n661 185
R17215 vdd.n3255 vdd.n3254 185
R17216 vdd.n3256 vdd.n3255 185
R17217 vdd.n669 vdd.n668 185
R17218 vdd.n3247 vdd.n668 185
R17219 vdd.n3250 vdd.n3249 185
R17220 vdd.n3249 vdd.n3248 185
R17221 vdd.n672 vdd.n671 185
R17222 vdd.n679 vdd.n672 185
R17223 vdd.n3238 vdd.n3237 185
R17224 vdd.n3239 vdd.n3238 185
R17225 vdd.n681 vdd.n680 185
R17226 vdd.n680 vdd.n678 185
R17227 vdd.n3233 vdd.n3232 185
R17228 vdd.n3232 vdd.n3231 185
R17229 vdd.n684 vdd.n683 185
R17230 vdd.n723 vdd.n684 185
R17231 vdd.n3221 vdd.n3220 185
R17232 vdd.n3219 vdd.n725 185
R17233 vdd.n3218 vdd.n724 185
R17234 vdd.n3223 vdd.n724 185
R17235 vdd.n729 vdd.n728 185
R17236 vdd.n733 vdd.n732 185
R17237 vdd.n3214 vdd.n734 185
R17238 vdd.n3213 vdd.n3212 185
R17239 vdd.n3211 vdd.n3210 185
R17240 vdd.n3209 vdd.n3208 185
R17241 vdd.n3207 vdd.n3206 185
R17242 vdd.n3205 vdd.n3204 185
R17243 vdd.n3203 vdd.n3202 185
R17244 vdd.n3201 vdd.n3200 185
R17245 vdd.n3199 vdd.n3198 185
R17246 vdd.n3197 vdd.n3196 185
R17247 vdd.n3195 vdd.n3194 185
R17248 vdd.n3193 vdd.n3192 185
R17249 vdd.n3191 vdd.n3190 185
R17250 vdd.n3189 vdd.n3188 185
R17251 vdd.n3187 vdd.n3186 185
R17252 vdd.n3178 vdd.n747 185
R17253 vdd.n3180 vdd.n3179 185
R17254 vdd.n3177 vdd.n3176 185
R17255 vdd.n3175 vdd.n3174 185
R17256 vdd.n3173 vdd.n3172 185
R17257 vdd.n3171 vdd.n3170 185
R17258 vdd.n3169 vdd.n3168 185
R17259 vdd.n3167 vdd.n3166 185
R17260 vdd.n3165 vdd.n3164 185
R17261 vdd.n3163 vdd.n3162 185
R17262 vdd.n3161 vdd.n3160 185
R17263 vdd.n3159 vdd.n3158 185
R17264 vdd.n3157 vdd.n3156 185
R17265 vdd.n3155 vdd.n3154 185
R17266 vdd.n3153 vdd.n3152 185
R17267 vdd.n3151 vdd.n3150 185
R17268 vdd.n3149 vdd.n3148 185
R17269 vdd.n3147 vdd.n3146 185
R17270 vdd.n3145 vdd.n3144 185
R17271 vdd.n3143 vdd.n3142 185
R17272 vdd.n3141 vdd.n3140 185
R17273 vdd.n3139 vdd.n3138 185
R17274 vdd.n3132 vdd.n767 185
R17275 vdd.n3134 vdd.n3133 185
R17276 vdd.n3131 vdd.n3130 185
R17277 vdd.n3129 vdd.n3128 185
R17278 vdd.n3127 vdd.n3126 185
R17279 vdd.n3125 vdd.n3124 185
R17280 vdd.n3123 vdd.n3122 185
R17281 vdd.n3121 vdd.n3120 185
R17282 vdd.n3119 vdd.n3118 185
R17283 vdd.n3117 vdd.n3116 185
R17284 vdd.n3115 vdd.n3114 185
R17285 vdd.n3113 vdd.n3112 185
R17286 vdd.n3111 vdd.n3110 185
R17287 vdd.n3109 vdd.n3108 185
R17288 vdd.n3107 vdd.n3106 185
R17289 vdd.n3105 vdd.n3104 185
R17290 vdd.n3103 vdd.n3102 185
R17291 vdd.n3101 vdd.n3100 185
R17292 vdd.n3099 vdd.n3098 185
R17293 vdd.n3097 vdd.n3096 185
R17294 vdd.n3095 vdd.n691 185
R17295 vdd.n3225 vdd.n3224 185
R17296 vdd.n3224 vdd.n3223 185
R17297 vdd.n3352 vdd.n3351 185
R17298 vdd.n618 vdd.n425 185
R17299 vdd.n617 vdd.n616 185
R17300 vdd.n615 vdd.n614 185
R17301 vdd.n613 vdd.n430 185
R17302 vdd.n609 vdd.n608 185
R17303 vdd.n607 vdd.n606 185
R17304 vdd.n605 vdd.n604 185
R17305 vdd.n603 vdd.n432 185
R17306 vdd.n599 vdd.n598 185
R17307 vdd.n597 vdd.n596 185
R17308 vdd.n595 vdd.n594 185
R17309 vdd.n593 vdd.n434 185
R17310 vdd.n589 vdd.n588 185
R17311 vdd.n587 vdd.n586 185
R17312 vdd.n585 vdd.n584 185
R17313 vdd.n583 vdd.n436 185
R17314 vdd.n579 vdd.n578 185
R17315 vdd.n577 vdd.n576 185
R17316 vdd.n575 vdd.n574 185
R17317 vdd.n573 vdd.n438 185
R17318 vdd.n569 vdd.n568 185
R17319 vdd.n567 vdd.n566 185
R17320 vdd.n565 vdd.n564 185
R17321 vdd.n563 vdd.n442 185
R17322 vdd.n559 vdd.n558 185
R17323 vdd.n557 vdd.n556 185
R17324 vdd.n555 vdd.n554 185
R17325 vdd.n553 vdd.n444 185
R17326 vdd.n549 vdd.n548 185
R17327 vdd.n547 vdd.n546 185
R17328 vdd.n545 vdd.n544 185
R17329 vdd.n543 vdd.n446 185
R17330 vdd.n539 vdd.n538 185
R17331 vdd.n537 vdd.n536 185
R17332 vdd.n535 vdd.n534 185
R17333 vdd.n533 vdd.n448 185
R17334 vdd.n529 vdd.n528 185
R17335 vdd.n527 vdd.n526 185
R17336 vdd.n525 vdd.n524 185
R17337 vdd.n523 vdd.n450 185
R17338 vdd.n519 vdd.n518 185
R17339 vdd.n517 vdd.n516 185
R17340 vdd.n515 vdd.n514 185
R17341 vdd.n513 vdd.n454 185
R17342 vdd.n509 vdd.n508 185
R17343 vdd.n507 vdd.n506 185
R17344 vdd.n505 vdd.n504 185
R17345 vdd.n503 vdd.n456 185
R17346 vdd.n499 vdd.n498 185
R17347 vdd.n497 vdd.n496 185
R17348 vdd.n495 vdd.n494 185
R17349 vdd.n493 vdd.n458 185
R17350 vdd.n489 vdd.n488 185
R17351 vdd.n487 vdd.n486 185
R17352 vdd.n485 vdd.n484 185
R17353 vdd.n483 vdd.n460 185
R17354 vdd.n479 vdd.n478 185
R17355 vdd.n477 vdd.n476 185
R17356 vdd.n475 vdd.n474 185
R17357 vdd.n473 vdd.n462 185
R17358 vdd.n469 vdd.n468 185
R17359 vdd.n467 vdd.n466 185
R17360 vdd.n465 vdd.n392 185
R17361 vdd.n3348 vdd.n393 185
R17362 vdd.n3355 vdd.n393 185
R17363 vdd.n3347 vdd.n3346 185
R17364 vdd.n3346 vdd.n386 185
R17365 vdd.n3345 vdd.n385 185
R17366 vdd.n3361 vdd.n385 185
R17367 vdd.n621 vdd.n384 185
R17368 vdd.n3362 vdd.n384 185
R17369 vdd.n3341 vdd.n383 185
R17370 vdd.n3363 vdd.n383 185
R17371 vdd.n3340 vdd.n3339 185
R17372 vdd.n3339 vdd.n375 185
R17373 vdd.n3338 vdd.n374 185
R17374 vdd.n3369 vdd.n374 185
R17375 vdd.n623 vdd.n373 185
R17376 vdd.n3370 vdd.n373 185
R17377 vdd.n3334 vdd.n372 185
R17378 vdd.n3371 vdd.n372 185
R17379 vdd.n3333 vdd.n3332 185
R17380 vdd.n3332 vdd.n3331 185
R17381 vdd.n3330 vdd.n364 185
R17382 vdd.n3377 vdd.n364 185
R17383 vdd.n625 vdd.n363 185
R17384 vdd.n3378 vdd.n363 185
R17385 vdd.n3326 vdd.n362 185
R17386 vdd.n3379 vdd.n362 185
R17387 vdd.n3325 vdd.n3324 185
R17388 vdd.n3324 vdd.n361 185
R17389 vdd.n3323 vdd.n353 185
R17390 vdd.n3385 vdd.n353 185
R17391 vdd.n627 vdd.n352 185
R17392 vdd.n3386 vdd.n352 185
R17393 vdd.n3319 vdd.n351 185
R17394 vdd.n3387 vdd.n351 185
R17395 vdd.n3318 vdd.n3317 185
R17396 vdd.n3317 vdd.n344 185
R17397 vdd.n3316 vdd.n343 185
R17398 vdd.n3393 vdd.n343 185
R17399 vdd.n629 vdd.n342 185
R17400 vdd.n3394 vdd.n342 185
R17401 vdd.n3312 vdd.n341 185
R17402 vdd.n3395 vdd.n341 185
R17403 vdd.n3311 vdd.n3310 185
R17404 vdd.n3310 vdd.n340 185
R17405 vdd.n3309 vdd.n631 185
R17406 vdd.n3309 vdd.n3308 185
R17407 vdd.n3297 vdd.n632 185
R17408 vdd.n633 vdd.n632 185
R17409 vdd.n3299 vdd.n3298 185
R17410 vdd.n3300 vdd.n3299 185
R17411 vdd.n640 vdd.n639 185
R17412 vdd.n644 vdd.n639 185
R17413 vdd.n3291 vdd.n3290 185
R17414 vdd.n3290 vdd.n3289 185
R17415 vdd.n643 vdd.n642 185
R17416 vdd.n3280 vdd.n643 185
R17417 vdd.n3279 vdd.n3278 185
R17418 vdd.n3281 vdd.n3279 185
R17419 vdd.n651 vdd.n650 185
R17420 vdd.n656 vdd.n650 185
R17421 vdd.n3274 vdd.n3273 185
R17422 vdd.n3273 vdd.n3272 185
R17423 vdd.n654 vdd.n653 185
R17424 vdd.n655 vdd.n654 185
R17425 vdd.n3263 vdd.n3262 185
R17426 vdd.n3264 vdd.n3263 185
R17427 vdd.n664 vdd.n663 185
R17428 vdd.n663 vdd.n662 185
R17429 vdd.n3258 vdd.n3257 185
R17430 vdd.n3257 vdd.n3256 185
R17431 vdd.n667 vdd.n666 185
R17432 vdd.n3247 vdd.n667 185
R17433 vdd.n3246 vdd.n3245 185
R17434 vdd.n3248 vdd.n3246 185
R17435 vdd.n674 vdd.n673 185
R17436 vdd.n679 vdd.n673 185
R17437 vdd.n3241 vdd.n3240 185
R17438 vdd.n3240 vdd.n3239 185
R17439 vdd.n677 vdd.n676 185
R17440 vdd.n678 vdd.n677 185
R17441 vdd.n3230 vdd.n3229 185
R17442 vdd.n3231 vdd.n3230 185
R17443 vdd.n686 vdd.n685 185
R17444 vdd.n723 vdd.n685 185
R17445 vdd.n913 vdd.n912 185
R17446 vdd.n2855 vdd.n2854 185
R17447 vdd.n2853 vdd.n2638 185
R17448 vdd.n2857 vdd.n2638 185
R17449 vdd.n2852 vdd.n2851 185
R17450 vdd.n2850 vdd.n2849 185
R17451 vdd.n2848 vdd.n2847 185
R17452 vdd.n2846 vdd.n2845 185
R17453 vdd.n2844 vdd.n2843 185
R17454 vdd.n2842 vdd.n2841 185
R17455 vdd.n2840 vdd.n2839 185
R17456 vdd.n2838 vdd.n2837 185
R17457 vdd.n2836 vdd.n2835 185
R17458 vdd.n2834 vdd.n2833 185
R17459 vdd.n2832 vdd.n2831 185
R17460 vdd.n2830 vdd.n2829 185
R17461 vdd.n2828 vdd.n2827 185
R17462 vdd.n2826 vdd.n2825 185
R17463 vdd.n2824 vdd.n2823 185
R17464 vdd.n2822 vdd.n2821 185
R17465 vdd.n2820 vdd.n2819 185
R17466 vdd.n2818 vdd.n2817 185
R17467 vdd.n2816 vdd.n2815 185
R17468 vdd.n2814 vdd.n2813 185
R17469 vdd.n2812 vdd.n2811 185
R17470 vdd.n2810 vdd.n2809 185
R17471 vdd.n2808 vdd.n2807 185
R17472 vdd.n2806 vdd.n2805 185
R17473 vdd.n2804 vdd.n2803 185
R17474 vdd.n2802 vdd.n2801 185
R17475 vdd.n2800 vdd.n2799 185
R17476 vdd.n2798 vdd.n2797 185
R17477 vdd.n2796 vdd.n2795 185
R17478 vdd.n2793 vdd.n2792 185
R17479 vdd.n2791 vdd.n2790 185
R17480 vdd.n2789 vdd.n2788 185
R17481 vdd.n2995 vdd.n2994 185
R17482 vdd.n2997 vdd.n834 185
R17483 vdd.n2999 vdd.n2998 185
R17484 vdd.n3001 vdd.n831 185
R17485 vdd.n3003 vdd.n3002 185
R17486 vdd.n3005 vdd.n829 185
R17487 vdd.n3007 vdd.n3006 185
R17488 vdd.n3008 vdd.n828 185
R17489 vdd.n3010 vdd.n3009 185
R17490 vdd.n3012 vdd.n826 185
R17491 vdd.n3014 vdd.n3013 185
R17492 vdd.n3015 vdd.n825 185
R17493 vdd.n3017 vdd.n3016 185
R17494 vdd.n3019 vdd.n823 185
R17495 vdd.n3021 vdd.n3020 185
R17496 vdd.n3022 vdd.n822 185
R17497 vdd.n3024 vdd.n3023 185
R17498 vdd.n3026 vdd.n731 185
R17499 vdd.n3028 vdd.n3027 185
R17500 vdd.n3030 vdd.n820 185
R17501 vdd.n3032 vdd.n3031 185
R17502 vdd.n3033 vdd.n819 185
R17503 vdd.n3035 vdd.n3034 185
R17504 vdd.n3037 vdd.n817 185
R17505 vdd.n3039 vdd.n3038 185
R17506 vdd.n3040 vdd.n816 185
R17507 vdd.n3042 vdd.n3041 185
R17508 vdd.n3044 vdd.n814 185
R17509 vdd.n3046 vdd.n3045 185
R17510 vdd.n3047 vdd.n813 185
R17511 vdd.n3049 vdd.n3048 185
R17512 vdd.n3051 vdd.n812 185
R17513 vdd.n3052 vdd.n811 185
R17514 vdd.n3055 vdd.n3054 185
R17515 vdd.n3056 vdd.n809 185
R17516 vdd.n809 vdd.n692 185
R17517 vdd.n2993 vdd.n806 185
R17518 vdd.n3059 vdd.n806 185
R17519 vdd.n2992 vdd.n2991 185
R17520 vdd.n2991 vdd.n805 185
R17521 vdd.n2990 vdd.n836 185
R17522 vdd.n2990 vdd.n2989 185
R17523 vdd.n2744 vdd.n837 185
R17524 vdd.n846 vdd.n837 185
R17525 vdd.n2745 vdd.n844 185
R17526 vdd.n2983 vdd.n844 185
R17527 vdd.n2747 vdd.n2746 185
R17528 vdd.n2746 vdd.n843 185
R17529 vdd.n2748 vdd.n852 185
R17530 vdd.n2932 vdd.n852 185
R17531 vdd.n2750 vdd.n2749 185
R17532 vdd.n2749 vdd.n851 185
R17533 vdd.n2751 vdd.n858 185
R17534 vdd.n2926 vdd.n858 185
R17535 vdd.n2753 vdd.n2752 185
R17536 vdd.n2752 vdd.n857 185
R17537 vdd.n2754 vdd.n863 185
R17538 vdd.n2918 vdd.n863 185
R17539 vdd.n2756 vdd.n2755 185
R17540 vdd.n2755 vdd.n870 185
R17541 vdd.n2757 vdd.n868 185
R17542 vdd.n2912 vdd.n868 185
R17543 vdd.n2759 vdd.n2758 185
R17544 vdd.n2760 vdd.n2759 185
R17545 vdd.n2743 vdd.n875 185
R17546 vdd.n2906 vdd.n875 185
R17547 vdd.n2742 vdd.n2741 185
R17548 vdd.n2741 vdd.n874 185
R17549 vdd.n2740 vdd.n881 185
R17550 vdd.n2900 vdd.n881 185
R17551 vdd.n2739 vdd.n2738 185
R17552 vdd.n2738 vdd.n880 185
R17553 vdd.n2737 vdd.n886 185
R17554 vdd.n2894 vdd.n886 185
R17555 vdd.n2736 vdd.n2735 185
R17556 vdd.n2735 vdd.n893 185
R17557 vdd.n2734 vdd.n891 185
R17558 vdd.n2888 vdd.n891 185
R17559 vdd.n2733 vdd.n2732 185
R17560 vdd.n2732 vdd.n900 185
R17561 vdd.n2731 vdd.n898 185
R17562 vdd.n2882 vdd.n898 185
R17563 vdd.n2730 vdd.n2729 185
R17564 vdd.n2729 vdd.n897 185
R17565 vdd.n2641 vdd.n904 185
R17566 vdd.n2876 vdd.n904 185
R17567 vdd.n2783 vdd.n2782 185
R17568 vdd.n2782 vdd.n2781 185
R17569 vdd.n2784 vdd.n909 185
R17570 vdd.n2870 vdd.n909 185
R17571 vdd.n2786 vdd.n2785 185
R17572 vdd.n2785 vdd.t4 185
R17573 vdd.n2787 vdd.n914 185
R17574 vdd.n2864 vdd.n914 185
R17575 vdd.n2866 vdd.n2865 185
R17576 vdd.n2865 vdd.n2864 185
R17577 vdd.n2867 vdd.n911 185
R17578 vdd.n911 vdd.t4 185
R17579 vdd.n2869 vdd.n2868 185
R17580 vdd.n2870 vdd.n2869 185
R17581 vdd.n903 vdd.n902 185
R17582 vdd.n2781 vdd.n903 185
R17583 vdd.n2878 vdd.n2877 185
R17584 vdd.n2877 vdd.n2876 185
R17585 vdd.n2879 vdd.n901 185
R17586 vdd.n901 vdd.n897 185
R17587 vdd.n2881 vdd.n2880 185
R17588 vdd.n2882 vdd.n2881 185
R17589 vdd.n890 vdd.n889 185
R17590 vdd.n900 vdd.n890 185
R17591 vdd.n2890 vdd.n2889 185
R17592 vdd.n2889 vdd.n2888 185
R17593 vdd.n2891 vdd.n888 185
R17594 vdd.n893 vdd.n888 185
R17595 vdd.n2893 vdd.n2892 185
R17596 vdd.n2894 vdd.n2893 185
R17597 vdd.n879 vdd.n878 185
R17598 vdd.n880 vdd.n879 185
R17599 vdd.n2902 vdd.n2901 185
R17600 vdd.n2901 vdd.n2900 185
R17601 vdd.n2903 vdd.n877 185
R17602 vdd.n877 vdd.n874 185
R17603 vdd.n2905 vdd.n2904 185
R17604 vdd.n2906 vdd.n2905 185
R17605 vdd.n867 vdd.n866 185
R17606 vdd.n2760 vdd.n867 185
R17607 vdd.n2914 vdd.n2913 185
R17608 vdd.n2913 vdd.n2912 185
R17609 vdd.n2915 vdd.n865 185
R17610 vdd.n870 vdd.n865 185
R17611 vdd.n2917 vdd.n2916 185
R17612 vdd.n2918 vdd.n2917 185
R17613 vdd.n856 vdd.n855 185
R17614 vdd.n857 vdd.n856 185
R17615 vdd.n2928 vdd.n2927 185
R17616 vdd.n2927 vdd.n2926 185
R17617 vdd.n2929 vdd.n854 185
R17618 vdd.n854 vdd.n851 185
R17619 vdd.n2931 vdd.n2930 185
R17620 vdd.n2932 vdd.n2931 185
R17621 vdd.n842 vdd.n841 185
R17622 vdd.n843 vdd.n842 185
R17623 vdd.n2985 vdd.n2984 185
R17624 vdd.n2984 vdd.n2983 185
R17625 vdd.n2986 vdd.n840 185
R17626 vdd.n846 vdd.n840 185
R17627 vdd.n2988 vdd.n2987 185
R17628 vdd.n2989 vdd.n2988 185
R17629 vdd.n810 vdd.n808 185
R17630 vdd.n808 vdd.n805 185
R17631 vdd.n3058 vdd.n3057 185
R17632 vdd.n3059 vdd.n3058 185
R17633 vdd.n2531 vdd.n2530 185
R17634 vdd.n2532 vdd.n2531 185
R17635 vdd.n964 vdd.n962 185
R17636 vdd.n962 vdd.t172 185
R17637 vdd.n2446 vdd.n971 185
R17638 vdd.n2457 vdd.n971 185
R17639 vdd.n2447 vdd.n980 185
R17640 vdd.n2156 vdd.n980 185
R17641 vdd.n2449 vdd.n2448 185
R17642 vdd.n2450 vdd.n2449 185
R17643 vdd.n2445 vdd.n979 185
R17644 vdd.n979 vdd.n976 185
R17645 vdd.n2444 vdd.n2443 185
R17646 vdd.n2443 vdd.n2442 185
R17647 vdd.n982 vdd.n981 185
R17648 vdd.n983 vdd.n982 185
R17649 vdd.n2435 vdd.n2434 185
R17650 vdd.n2436 vdd.n2435 185
R17651 vdd.n2433 vdd.n992 185
R17652 vdd.n992 vdd.n989 185
R17653 vdd.n2432 vdd.n2431 185
R17654 vdd.n2431 vdd.n2430 185
R17655 vdd.n994 vdd.n993 185
R17656 vdd.n1002 vdd.n994 185
R17657 vdd.n2423 vdd.n2422 185
R17658 vdd.n2424 vdd.n2423 185
R17659 vdd.n2421 vdd.n1003 185
R17660 vdd.n1008 vdd.n1003 185
R17661 vdd.n2420 vdd.n2419 185
R17662 vdd.n2419 vdd.n2418 185
R17663 vdd.n1005 vdd.n1004 185
R17664 vdd.n2257 vdd.n1005 185
R17665 vdd.n2411 vdd.n2410 185
R17666 vdd.n2412 vdd.n2411 185
R17667 vdd.n2409 vdd.n1015 185
R17668 vdd.n1015 vdd.n1012 185
R17669 vdd.n2408 vdd.n2407 185
R17670 vdd.n2407 vdd.n2406 185
R17671 vdd.n1017 vdd.n1016 185
R17672 vdd.n1018 vdd.n1017 185
R17673 vdd.n2399 vdd.n2398 185
R17674 vdd.n2400 vdd.n2399 185
R17675 vdd.n2396 vdd.n1026 185
R17676 vdd.n1033 vdd.n1026 185
R17677 vdd.n2395 vdd.n2394 185
R17678 vdd.n2394 vdd.n2393 185
R17679 vdd.n1029 vdd.n1028 185
R17680 vdd.n1030 vdd.n1029 185
R17681 vdd.n2386 vdd.n2385 185
R17682 vdd.n2387 vdd.n2386 185
R17683 vdd.n2384 vdd.n1040 185
R17684 vdd.n1040 vdd.n1037 185
R17685 vdd.n2383 vdd.n2382 185
R17686 vdd.n2382 vdd.n2381 185
R17687 vdd.n1042 vdd.n1041 185
R17688 vdd.n1043 vdd.n1042 185
R17689 vdd.n2374 vdd.n2373 185
R17690 vdd.n2375 vdd.n2374 185
R17691 vdd.n2462 vdd.n936 185
R17692 vdd.n2604 vdd.n936 185
R17693 vdd.n2464 vdd.n2463 185
R17694 vdd.n2466 vdd.n2465 185
R17695 vdd.n2468 vdd.n2467 185
R17696 vdd.n2470 vdd.n2469 185
R17697 vdd.n2472 vdd.n2471 185
R17698 vdd.n2474 vdd.n2473 185
R17699 vdd.n2476 vdd.n2475 185
R17700 vdd.n2478 vdd.n2477 185
R17701 vdd.n2480 vdd.n2479 185
R17702 vdd.n2482 vdd.n2481 185
R17703 vdd.n2484 vdd.n2483 185
R17704 vdd.n2486 vdd.n2485 185
R17705 vdd.n2488 vdd.n2487 185
R17706 vdd.n2490 vdd.n2489 185
R17707 vdd.n2492 vdd.n2491 185
R17708 vdd.n2494 vdd.n2493 185
R17709 vdd.n2496 vdd.n2495 185
R17710 vdd.n2498 vdd.n2497 185
R17711 vdd.n2500 vdd.n2499 185
R17712 vdd.n2502 vdd.n2501 185
R17713 vdd.n2504 vdd.n2503 185
R17714 vdd.n2506 vdd.n2505 185
R17715 vdd.n2508 vdd.n2507 185
R17716 vdd.n2510 vdd.n2509 185
R17717 vdd.n2512 vdd.n2511 185
R17718 vdd.n2514 vdd.n2513 185
R17719 vdd.n2516 vdd.n2515 185
R17720 vdd.n2518 vdd.n2517 185
R17721 vdd.n2520 vdd.n2519 185
R17722 vdd.n2522 vdd.n2521 185
R17723 vdd.n2524 vdd.n2523 185
R17724 vdd.n2526 vdd.n2525 185
R17725 vdd.n2528 vdd.n2527 185
R17726 vdd.n2529 vdd.n963 185
R17727 vdd.n2461 vdd.n961 185
R17728 vdd.n2532 vdd.n961 185
R17729 vdd.n2460 vdd.n2459 185
R17730 vdd.n2459 vdd.t172 185
R17731 vdd.n2458 vdd.n968 185
R17732 vdd.n2458 vdd.n2457 185
R17733 vdd.n2238 vdd.n969 185
R17734 vdd.n2156 vdd.n969 185
R17735 vdd.n2239 vdd.n978 185
R17736 vdd.n2450 vdd.n978 185
R17737 vdd.n2241 vdd.n2240 185
R17738 vdd.n2240 vdd.n976 185
R17739 vdd.n2242 vdd.n985 185
R17740 vdd.n2442 vdd.n985 185
R17741 vdd.n2244 vdd.n2243 185
R17742 vdd.n2243 vdd.n983 185
R17743 vdd.n2245 vdd.n991 185
R17744 vdd.n2436 vdd.n991 185
R17745 vdd.n2247 vdd.n2246 185
R17746 vdd.n2246 vdd.n989 185
R17747 vdd.n2248 vdd.n996 185
R17748 vdd.n2430 vdd.n996 185
R17749 vdd.n2250 vdd.n2249 185
R17750 vdd.n2249 vdd.n1002 185
R17751 vdd.n2251 vdd.n1001 185
R17752 vdd.n2424 vdd.n1001 185
R17753 vdd.n2253 vdd.n2252 185
R17754 vdd.n2252 vdd.n1008 185
R17755 vdd.n2254 vdd.n1007 185
R17756 vdd.n2418 vdd.n1007 185
R17757 vdd.n2256 vdd.n2255 185
R17758 vdd.n2257 vdd.n2256 185
R17759 vdd.n2237 vdd.n1014 185
R17760 vdd.n2412 vdd.n1014 185
R17761 vdd.n2236 vdd.n2235 185
R17762 vdd.n2235 vdd.n1012 185
R17763 vdd.n2234 vdd.n1020 185
R17764 vdd.n2406 vdd.n1020 185
R17765 vdd.n2233 vdd.n2232 185
R17766 vdd.n2232 vdd.n1018 185
R17767 vdd.n2231 vdd.n1025 185
R17768 vdd.n2400 vdd.n1025 185
R17769 vdd.n2230 vdd.n2229 185
R17770 vdd.n2229 vdd.n1033 185
R17771 vdd.n2228 vdd.n1032 185
R17772 vdd.n2393 vdd.n1032 185
R17773 vdd.n2227 vdd.n2226 185
R17774 vdd.n2226 vdd.n1030 185
R17775 vdd.n2225 vdd.n1039 185
R17776 vdd.n2387 vdd.n1039 185
R17777 vdd.n2224 vdd.n2223 185
R17778 vdd.n2223 vdd.n1037 185
R17779 vdd.n2222 vdd.n1045 185
R17780 vdd.n2381 vdd.n1045 185
R17781 vdd.n2221 vdd.n2220 185
R17782 vdd.n2220 vdd.n1043 185
R17783 vdd.n2219 vdd.n1051 185
R17784 vdd.n2375 vdd.n1051 185
R17785 vdd.n2372 vdd.n1052 185
R17786 vdd.n2371 vdd.n2370 185
R17787 vdd.n2368 vdd.n1053 185
R17788 vdd.n2366 vdd.n2365 185
R17789 vdd.n2364 vdd.n1054 185
R17790 vdd.n2363 vdd.n2362 185
R17791 vdd.n2360 vdd.n1055 185
R17792 vdd.n2358 vdd.n2357 185
R17793 vdd.n2356 vdd.n1056 185
R17794 vdd.n2355 vdd.n2354 185
R17795 vdd.n2352 vdd.n1057 185
R17796 vdd.n2350 vdd.n2349 185
R17797 vdd.n2348 vdd.n1058 185
R17798 vdd.n2347 vdd.n2346 185
R17799 vdd.n2344 vdd.n1059 185
R17800 vdd.n2342 vdd.n2341 185
R17801 vdd.n2340 vdd.n1060 185
R17802 vdd.n2339 vdd.n1062 185
R17803 vdd.n2184 vdd.n1063 185
R17804 vdd.n2187 vdd.n2186 185
R17805 vdd.n2189 vdd.n2188 185
R17806 vdd.n2191 vdd.n2183 185
R17807 vdd.n2194 vdd.n2193 185
R17808 vdd.n2195 vdd.n2182 185
R17809 vdd.n2197 vdd.n2196 185
R17810 vdd.n2199 vdd.n2181 185
R17811 vdd.n2202 vdd.n2201 185
R17812 vdd.n2203 vdd.n2180 185
R17813 vdd.n2205 vdd.n2204 185
R17814 vdd.n2207 vdd.n2179 185
R17815 vdd.n2210 vdd.n2209 185
R17816 vdd.n2211 vdd.n2176 185
R17817 vdd.n2214 vdd.n2213 185
R17818 vdd.n2216 vdd.n2175 185
R17819 vdd.n2218 vdd.n2217 185
R17820 vdd.n2217 vdd.n1049 185
R17821 vdd.n327 vdd.n326 171.744
R17822 vdd.n326 vdd.n325 171.744
R17823 vdd.n325 vdd.n294 171.744
R17824 vdd.n318 vdd.n294 171.744
R17825 vdd.n318 vdd.n317 171.744
R17826 vdd.n317 vdd.n299 171.744
R17827 vdd.n310 vdd.n299 171.744
R17828 vdd.n310 vdd.n309 171.744
R17829 vdd.n309 vdd.n303 171.744
R17830 vdd.n268 vdd.n267 171.744
R17831 vdd.n267 vdd.n266 171.744
R17832 vdd.n266 vdd.n235 171.744
R17833 vdd.n259 vdd.n235 171.744
R17834 vdd.n259 vdd.n258 171.744
R17835 vdd.n258 vdd.n240 171.744
R17836 vdd.n251 vdd.n240 171.744
R17837 vdd.n251 vdd.n250 171.744
R17838 vdd.n250 vdd.n244 171.744
R17839 vdd.n225 vdd.n224 171.744
R17840 vdd.n224 vdd.n223 171.744
R17841 vdd.n223 vdd.n192 171.744
R17842 vdd.n216 vdd.n192 171.744
R17843 vdd.n216 vdd.n215 171.744
R17844 vdd.n215 vdd.n197 171.744
R17845 vdd.n208 vdd.n197 171.744
R17846 vdd.n208 vdd.n207 171.744
R17847 vdd.n207 vdd.n201 171.744
R17848 vdd.n166 vdd.n165 171.744
R17849 vdd.n165 vdd.n164 171.744
R17850 vdd.n164 vdd.n133 171.744
R17851 vdd.n157 vdd.n133 171.744
R17852 vdd.n157 vdd.n156 171.744
R17853 vdd.n156 vdd.n138 171.744
R17854 vdd.n149 vdd.n138 171.744
R17855 vdd.n149 vdd.n148 171.744
R17856 vdd.n148 vdd.n142 171.744
R17857 vdd.n124 vdd.n123 171.744
R17858 vdd.n123 vdd.n122 171.744
R17859 vdd.n122 vdd.n91 171.744
R17860 vdd.n115 vdd.n91 171.744
R17861 vdd.n115 vdd.n114 171.744
R17862 vdd.n114 vdd.n96 171.744
R17863 vdd.n107 vdd.n96 171.744
R17864 vdd.n107 vdd.n106 171.744
R17865 vdd.n106 vdd.n100 171.744
R17866 vdd.n65 vdd.n64 171.744
R17867 vdd.n64 vdd.n63 171.744
R17868 vdd.n63 vdd.n32 171.744
R17869 vdd.n56 vdd.n32 171.744
R17870 vdd.n56 vdd.n55 171.744
R17871 vdd.n55 vdd.n37 171.744
R17872 vdd.n48 vdd.n37 171.744
R17873 vdd.n48 vdd.n47 171.744
R17874 vdd.n47 vdd.n41 171.744
R17875 vdd.n1746 vdd.n1745 171.744
R17876 vdd.n1745 vdd.n1744 171.744
R17877 vdd.n1744 vdd.n1713 171.744
R17878 vdd.n1737 vdd.n1713 171.744
R17879 vdd.n1737 vdd.n1736 171.744
R17880 vdd.n1736 vdd.n1718 171.744
R17881 vdd.n1729 vdd.n1718 171.744
R17882 vdd.n1729 vdd.n1728 171.744
R17883 vdd.n1728 vdd.n1722 171.744
R17884 vdd.n1805 vdd.n1804 171.744
R17885 vdd.n1804 vdd.n1803 171.744
R17886 vdd.n1803 vdd.n1772 171.744
R17887 vdd.n1796 vdd.n1772 171.744
R17888 vdd.n1796 vdd.n1795 171.744
R17889 vdd.n1795 vdd.n1777 171.744
R17890 vdd.n1788 vdd.n1777 171.744
R17891 vdd.n1788 vdd.n1787 171.744
R17892 vdd.n1787 vdd.n1781 171.744
R17893 vdd.n1644 vdd.n1643 171.744
R17894 vdd.n1643 vdd.n1642 171.744
R17895 vdd.n1642 vdd.n1611 171.744
R17896 vdd.n1635 vdd.n1611 171.744
R17897 vdd.n1635 vdd.n1634 171.744
R17898 vdd.n1634 vdd.n1616 171.744
R17899 vdd.n1627 vdd.n1616 171.744
R17900 vdd.n1627 vdd.n1626 171.744
R17901 vdd.n1626 vdd.n1620 171.744
R17902 vdd.n1703 vdd.n1702 171.744
R17903 vdd.n1702 vdd.n1701 171.744
R17904 vdd.n1701 vdd.n1670 171.744
R17905 vdd.n1694 vdd.n1670 171.744
R17906 vdd.n1694 vdd.n1693 171.744
R17907 vdd.n1693 vdd.n1675 171.744
R17908 vdd.n1686 vdd.n1675 171.744
R17909 vdd.n1686 vdd.n1685 171.744
R17910 vdd.n1685 vdd.n1679 171.744
R17911 vdd.n1543 vdd.n1542 171.744
R17912 vdd.n1542 vdd.n1541 171.744
R17913 vdd.n1541 vdd.n1510 171.744
R17914 vdd.n1534 vdd.n1510 171.744
R17915 vdd.n1534 vdd.n1533 171.744
R17916 vdd.n1533 vdd.n1515 171.744
R17917 vdd.n1526 vdd.n1515 171.744
R17918 vdd.n1526 vdd.n1525 171.744
R17919 vdd.n1525 vdd.n1519 171.744
R17920 vdd.n1602 vdd.n1601 171.744
R17921 vdd.n1601 vdd.n1600 171.744
R17922 vdd.n1600 vdd.n1569 171.744
R17923 vdd.n1593 vdd.n1569 171.744
R17924 vdd.n1593 vdd.n1592 171.744
R17925 vdd.n1592 vdd.n1574 171.744
R17926 vdd.n1585 vdd.n1574 171.744
R17927 vdd.n1585 vdd.n1584 171.744
R17928 vdd.n1584 vdd.n1578 171.744
R17929 vdd.n468 vdd.n467 146.341
R17930 vdd.n474 vdd.n473 146.341
R17931 vdd.n478 vdd.n477 146.341
R17932 vdd.n484 vdd.n483 146.341
R17933 vdd.n488 vdd.n487 146.341
R17934 vdd.n494 vdd.n493 146.341
R17935 vdd.n498 vdd.n497 146.341
R17936 vdd.n504 vdd.n503 146.341
R17937 vdd.n508 vdd.n507 146.341
R17938 vdd.n514 vdd.n513 146.341
R17939 vdd.n518 vdd.n517 146.341
R17940 vdd.n524 vdd.n523 146.341
R17941 vdd.n528 vdd.n527 146.341
R17942 vdd.n534 vdd.n533 146.341
R17943 vdd.n538 vdd.n537 146.341
R17944 vdd.n544 vdd.n543 146.341
R17945 vdd.n548 vdd.n547 146.341
R17946 vdd.n554 vdd.n553 146.341
R17947 vdd.n558 vdd.n557 146.341
R17948 vdd.n564 vdd.n563 146.341
R17949 vdd.n568 vdd.n567 146.341
R17950 vdd.n574 vdd.n573 146.341
R17951 vdd.n578 vdd.n577 146.341
R17952 vdd.n584 vdd.n583 146.341
R17953 vdd.n588 vdd.n587 146.341
R17954 vdd.n594 vdd.n593 146.341
R17955 vdd.n598 vdd.n597 146.341
R17956 vdd.n604 vdd.n603 146.341
R17957 vdd.n608 vdd.n607 146.341
R17958 vdd.n614 vdd.n613 146.341
R17959 vdd.n616 vdd.n425 146.341
R17960 vdd.n3230 vdd.n685 146.341
R17961 vdd.n3230 vdd.n677 146.341
R17962 vdd.n3240 vdd.n677 146.341
R17963 vdd.n3240 vdd.n673 146.341
R17964 vdd.n3246 vdd.n673 146.341
R17965 vdd.n3246 vdd.n667 146.341
R17966 vdd.n3257 vdd.n667 146.341
R17967 vdd.n3257 vdd.n663 146.341
R17968 vdd.n3263 vdd.n663 146.341
R17969 vdd.n3263 vdd.n654 146.341
R17970 vdd.n3273 vdd.n654 146.341
R17971 vdd.n3273 vdd.n650 146.341
R17972 vdd.n3279 vdd.n650 146.341
R17973 vdd.n3279 vdd.n643 146.341
R17974 vdd.n3290 vdd.n643 146.341
R17975 vdd.n3290 vdd.n639 146.341
R17976 vdd.n3299 vdd.n639 146.341
R17977 vdd.n3299 vdd.n632 146.341
R17978 vdd.n3309 vdd.n632 146.341
R17979 vdd.n3310 vdd.n3309 146.341
R17980 vdd.n3310 vdd.n341 146.341
R17981 vdd.n342 vdd.n341 146.341
R17982 vdd.n343 vdd.n342 146.341
R17983 vdd.n3317 vdd.n343 146.341
R17984 vdd.n3317 vdd.n351 146.341
R17985 vdd.n352 vdd.n351 146.341
R17986 vdd.n353 vdd.n352 146.341
R17987 vdd.n3324 vdd.n353 146.341
R17988 vdd.n3324 vdd.n362 146.341
R17989 vdd.n363 vdd.n362 146.341
R17990 vdd.n364 vdd.n363 146.341
R17991 vdd.n3332 vdd.n364 146.341
R17992 vdd.n3332 vdd.n372 146.341
R17993 vdd.n373 vdd.n372 146.341
R17994 vdd.n374 vdd.n373 146.341
R17995 vdd.n3339 vdd.n374 146.341
R17996 vdd.n3339 vdd.n383 146.341
R17997 vdd.n384 vdd.n383 146.341
R17998 vdd.n385 vdd.n384 146.341
R17999 vdd.n3346 vdd.n385 146.341
R18000 vdd.n3346 vdd.n393 146.341
R18001 vdd.n725 vdd.n724 146.341
R18002 vdd.n728 vdd.n724 146.341
R18003 vdd.n734 vdd.n733 146.341
R18004 vdd.n3212 vdd.n3211 146.341
R18005 vdd.n3208 vdd.n3207 146.341
R18006 vdd.n3204 vdd.n3203 146.341
R18007 vdd.n3200 vdd.n3199 146.341
R18008 vdd.n3196 vdd.n3195 146.341
R18009 vdd.n3192 vdd.n3191 146.341
R18010 vdd.n3188 vdd.n3187 146.341
R18011 vdd.n3179 vdd.n3178 146.341
R18012 vdd.n3176 vdd.n3175 146.341
R18013 vdd.n3172 vdd.n3171 146.341
R18014 vdd.n3168 vdd.n3167 146.341
R18015 vdd.n3164 vdd.n3163 146.341
R18016 vdd.n3160 vdd.n3159 146.341
R18017 vdd.n3156 vdd.n3155 146.341
R18018 vdd.n3152 vdd.n3151 146.341
R18019 vdd.n3148 vdd.n3147 146.341
R18020 vdd.n3144 vdd.n3143 146.341
R18021 vdd.n3140 vdd.n3139 146.341
R18022 vdd.n3133 vdd.n3132 146.341
R18023 vdd.n3130 vdd.n3129 146.341
R18024 vdd.n3126 vdd.n3125 146.341
R18025 vdd.n3122 vdd.n3121 146.341
R18026 vdd.n3118 vdd.n3117 146.341
R18027 vdd.n3114 vdd.n3113 146.341
R18028 vdd.n3110 vdd.n3109 146.341
R18029 vdd.n3106 vdd.n3105 146.341
R18030 vdd.n3102 vdd.n3101 146.341
R18031 vdd.n3098 vdd.n3097 146.341
R18032 vdd.n3224 vdd.n691 146.341
R18033 vdd.n3232 vdd.n684 146.341
R18034 vdd.n3232 vdd.n680 146.341
R18035 vdd.n3238 vdd.n680 146.341
R18036 vdd.n3238 vdd.n672 146.341
R18037 vdd.n3249 vdd.n672 146.341
R18038 vdd.n3249 vdd.n668 146.341
R18039 vdd.n3255 vdd.n668 146.341
R18040 vdd.n3255 vdd.n661 146.341
R18041 vdd.n3265 vdd.n661 146.341
R18042 vdd.n3265 vdd.n657 146.341
R18043 vdd.n3271 vdd.n657 146.341
R18044 vdd.n3271 vdd.n649 146.341
R18045 vdd.n3282 vdd.n649 146.341
R18046 vdd.n3282 vdd.n645 146.341
R18047 vdd.n3288 vdd.n645 146.341
R18048 vdd.n3288 vdd.n638 146.341
R18049 vdd.n3301 vdd.n638 146.341
R18050 vdd.n3301 vdd.n634 146.341
R18051 vdd.n3307 vdd.n634 146.341
R18052 vdd.n3307 vdd.n338 146.341
R18053 vdd.n3396 vdd.n338 146.341
R18054 vdd.n3396 vdd.n339 146.341
R18055 vdd.n3392 vdd.n339 146.341
R18056 vdd.n3392 vdd.n345 146.341
R18057 vdd.n3388 vdd.n345 146.341
R18058 vdd.n3388 vdd.n350 146.341
R18059 vdd.n3384 vdd.n350 146.341
R18060 vdd.n3384 vdd.n354 146.341
R18061 vdd.n3380 vdd.n354 146.341
R18062 vdd.n3380 vdd.n360 146.341
R18063 vdd.n3376 vdd.n360 146.341
R18064 vdd.n3376 vdd.n365 146.341
R18065 vdd.n3372 vdd.n365 146.341
R18066 vdd.n3372 vdd.n371 146.341
R18067 vdd.n3368 vdd.n371 146.341
R18068 vdd.n3368 vdd.n376 146.341
R18069 vdd.n3364 vdd.n376 146.341
R18070 vdd.n3364 vdd.n382 146.341
R18071 vdd.n3360 vdd.n382 146.341
R18072 vdd.n3360 vdd.n387 146.341
R18073 vdd.n3356 vdd.n387 146.341
R18074 vdd.n2322 vdd.n2321 146.341
R18075 vdd.n2319 vdd.n1903 146.341
R18076 vdd.n2099 vdd.n1909 146.341
R18077 vdd.n2097 vdd.n2096 146.341
R18078 vdd.n2094 vdd.n1911 146.341
R18079 vdd.n2090 vdd.n2089 146.341
R18080 vdd.n2087 vdd.n1918 146.341
R18081 vdd.n2083 vdd.n2082 146.341
R18082 vdd.n2080 vdd.n1925 146.341
R18083 vdd.n1936 vdd.n1933 146.341
R18084 vdd.n2072 vdd.n2071 146.341
R18085 vdd.n2069 vdd.n1938 146.341
R18086 vdd.n2065 vdd.n2064 146.341
R18087 vdd.n2062 vdd.n1944 146.341
R18088 vdd.n2058 vdd.n2057 146.341
R18089 vdd.n2055 vdd.n1951 146.341
R18090 vdd.n2051 vdd.n2050 146.341
R18091 vdd.n2048 vdd.n1958 146.341
R18092 vdd.n2044 vdd.n2043 146.341
R18093 vdd.n2041 vdd.n1965 146.341
R18094 vdd.n1976 vdd.n1973 146.341
R18095 vdd.n2033 vdd.n2032 146.341
R18096 vdd.n2030 vdd.n1978 146.341
R18097 vdd.n2026 vdd.n2025 146.341
R18098 vdd.n2023 vdd.n1984 146.341
R18099 vdd.n2019 vdd.n2018 146.341
R18100 vdd.n2016 vdd.n1991 146.341
R18101 vdd.n2012 vdd.n2011 146.341
R18102 vdd.n2009 vdd.n2006 146.341
R18103 vdd.n2004 vdd.n2001 146.341
R18104 vdd.n1999 vdd.n1069 146.341
R18105 vdd.n1428 vdd.n1188 146.341
R18106 vdd.n1428 vdd.n1184 146.341
R18107 vdd.n1434 vdd.n1184 146.341
R18108 vdd.n1434 vdd.n1176 146.341
R18109 vdd.n1445 vdd.n1176 146.341
R18110 vdd.n1445 vdd.n1172 146.341
R18111 vdd.n1451 vdd.n1172 146.341
R18112 vdd.n1451 vdd.n1166 146.341
R18113 vdd.n1462 vdd.n1166 146.341
R18114 vdd.n1462 vdd.n1162 146.341
R18115 vdd.n1468 vdd.n1162 146.341
R18116 vdd.n1468 vdd.n1153 146.341
R18117 vdd.n1478 vdd.n1153 146.341
R18118 vdd.n1478 vdd.n1149 146.341
R18119 vdd.n1484 vdd.n1149 146.341
R18120 vdd.n1484 vdd.n1142 146.341
R18121 vdd.n1495 vdd.n1142 146.341
R18122 vdd.n1495 vdd.n1138 146.341
R18123 vdd.n1501 vdd.n1138 146.341
R18124 vdd.n1501 vdd.n1131 146.341
R18125 vdd.n1818 vdd.n1131 146.341
R18126 vdd.n1818 vdd.n1127 146.341
R18127 vdd.n1824 vdd.n1127 146.341
R18128 vdd.n1824 vdd.n1119 146.341
R18129 vdd.n1835 vdd.n1119 146.341
R18130 vdd.n1835 vdd.n1115 146.341
R18131 vdd.n1841 vdd.n1115 146.341
R18132 vdd.n1841 vdd.n1109 146.341
R18133 vdd.n1852 vdd.n1109 146.341
R18134 vdd.n1852 vdd.n1105 146.341
R18135 vdd.n1858 vdd.n1105 146.341
R18136 vdd.n1858 vdd.n1096 146.341
R18137 vdd.n1868 vdd.n1096 146.341
R18138 vdd.n1868 vdd.n1092 146.341
R18139 vdd.n1874 vdd.n1092 146.341
R18140 vdd.n1874 vdd.n1086 146.341
R18141 vdd.n1885 vdd.n1086 146.341
R18142 vdd.n1885 vdd.n1081 146.341
R18143 vdd.n1893 vdd.n1081 146.341
R18144 vdd.n1893 vdd.n1071 146.341
R18145 vdd.n2330 vdd.n1071 146.341
R18146 vdd.n1417 vdd.n1193 146.341
R18147 vdd.n1417 vdd.n1226 146.341
R18148 vdd.n1230 vdd.n1229 146.341
R18149 vdd.n1232 vdd.n1231 146.341
R18150 vdd.n1236 vdd.n1235 146.341
R18151 vdd.n1238 vdd.n1237 146.341
R18152 vdd.n1242 vdd.n1241 146.341
R18153 vdd.n1244 vdd.n1243 146.341
R18154 vdd.n1248 vdd.n1247 146.341
R18155 vdd.n1250 vdd.n1249 146.341
R18156 vdd.n1256 vdd.n1255 146.341
R18157 vdd.n1258 vdd.n1257 146.341
R18158 vdd.n1262 vdd.n1261 146.341
R18159 vdd.n1264 vdd.n1263 146.341
R18160 vdd.n1268 vdd.n1267 146.341
R18161 vdd.n1270 vdd.n1269 146.341
R18162 vdd.n1274 vdd.n1273 146.341
R18163 vdd.n1276 vdd.n1275 146.341
R18164 vdd.n1280 vdd.n1279 146.341
R18165 vdd.n1282 vdd.n1281 146.341
R18166 vdd.n1354 vdd.n1285 146.341
R18167 vdd.n1287 vdd.n1286 146.341
R18168 vdd.n1291 vdd.n1290 146.341
R18169 vdd.n1293 vdd.n1292 146.341
R18170 vdd.n1297 vdd.n1296 146.341
R18171 vdd.n1299 vdd.n1298 146.341
R18172 vdd.n1303 vdd.n1302 146.341
R18173 vdd.n1305 vdd.n1304 146.341
R18174 vdd.n1309 vdd.n1308 146.341
R18175 vdd.n1311 vdd.n1310 146.341
R18176 vdd.n1315 vdd.n1314 146.341
R18177 vdd.n1316 vdd.n1224 146.341
R18178 vdd.n1426 vdd.n1189 146.341
R18179 vdd.n1426 vdd.n1182 146.341
R18180 vdd.n1437 vdd.n1182 146.341
R18181 vdd.n1437 vdd.n1178 146.341
R18182 vdd.n1443 vdd.n1178 146.341
R18183 vdd.n1443 vdd.n1171 146.341
R18184 vdd.n1454 vdd.n1171 146.341
R18185 vdd.n1454 vdd.n1167 146.341
R18186 vdd.n1460 vdd.n1167 146.341
R18187 vdd.n1460 vdd.n1160 146.341
R18188 vdd.n1470 vdd.n1160 146.341
R18189 vdd.n1470 vdd.n1156 146.341
R18190 vdd.n1476 vdd.n1156 146.341
R18191 vdd.n1476 vdd.n1148 146.341
R18192 vdd.n1487 vdd.n1148 146.341
R18193 vdd.n1487 vdd.n1144 146.341
R18194 vdd.n1493 vdd.n1144 146.341
R18195 vdd.n1493 vdd.n1137 146.341
R18196 vdd.n1503 vdd.n1137 146.341
R18197 vdd.n1503 vdd.n1133 146.341
R18198 vdd.n1816 vdd.n1133 146.341
R18199 vdd.n1816 vdd.n1125 146.341
R18200 vdd.n1827 vdd.n1125 146.341
R18201 vdd.n1827 vdd.n1121 146.341
R18202 vdd.n1833 vdd.n1121 146.341
R18203 vdd.n1833 vdd.n1114 146.341
R18204 vdd.n1844 vdd.n1114 146.341
R18205 vdd.n1844 vdd.n1110 146.341
R18206 vdd.n1850 vdd.n1110 146.341
R18207 vdd.n1850 vdd.n1103 146.341
R18208 vdd.n1860 vdd.n1103 146.341
R18209 vdd.n1860 vdd.n1099 146.341
R18210 vdd.n1866 vdd.n1099 146.341
R18211 vdd.n1866 vdd.n1091 146.341
R18212 vdd.n1877 vdd.n1091 146.341
R18213 vdd.n1877 vdd.n1087 146.341
R18214 vdd.n1883 vdd.n1087 146.341
R18215 vdd.n1883 vdd.n1079 146.341
R18216 vdd.n1896 vdd.n1079 146.341
R18217 vdd.n1896 vdd.n1074 146.341
R18218 vdd.n2328 vdd.n1074 146.341
R18219 vdd.n1073 vdd.n1049 141.707
R18220 vdd.n3223 vdd.n692 141.707
R18221 vdd.n2177 vdd.t262 127.284
R18222 vdd.n965 vdd.t247 127.284
R18223 vdd.n2151 vdd.t209 127.284
R18224 vdd.n957 vdd.t271 127.284
R18225 vdd.n2922 vdd.t223 127.284
R18226 vdd.n2922 vdd.t224 127.284
R18227 vdd.n2642 vdd.t269 127.284
R18228 vdd.n832 vdd.t251 127.284
R18229 vdd.n2639 vdd.t256 127.284
R18230 vdd.n799 vdd.t258 127.284
R18231 vdd.n1027 vdd.t265 127.284
R18232 vdd.n1027 vdd.t266 127.284
R18233 vdd.n22 vdd.n20 117.314
R18234 vdd.n17 vdd.n15 117.314
R18235 vdd.n27 vdd.n26 116.927
R18236 vdd.n24 vdd.n23 116.927
R18237 vdd.n22 vdd.n21 116.927
R18238 vdd.n17 vdd.n16 116.927
R18239 vdd.n19 vdd.n18 116.927
R18240 vdd.n27 vdd.n25 116.927
R18241 vdd.n2178 vdd.t261 111.188
R18242 vdd.n966 vdd.t248 111.188
R18243 vdd.n2152 vdd.t208 111.188
R18244 vdd.n958 vdd.t272 111.188
R18245 vdd.n2643 vdd.t268 111.188
R18246 vdd.n833 vdd.t252 111.188
R18247 vdd.n2640 vdd.t255 111.188
R18248 vdd.n800 vdd.t259 111.188
R18249 vdd.n2865 vdd.n911 99.5127
R18250 vdd.n2869 vdd.n911 99.5127
R18251 vdd.n2869 vdd.n903 99.5127
R18252 vdd.n2877 vdd.n903 99.5127
R18253 vdd.n2877 vdd.n901 99.5127
R18254 vdd.n2881 vdd.n901 99.5127
R18255 vdd.n2881 vdd.n890 99.5127
R18256 vdd.n2889 vdd.n890 99.5127
R18257 vdd.n2889 vdd.n888 99.5127
R18258 vdd.n2893 vdd.n888 99.5127
R18259 vdd.n2893 vdd.n879 99.5127
R18260 vdd.n2901 vdd.n879 99.5127
R18261 vdd.n2901 vdd.n877 99.5127
R18262 vdd.n2905 vdd.n877 99.5127
R18263 vdd.n2905 vdd.n867 99.5127
R18264 vdd.n2913 vdd.n867 99.5127
R18265 vdd.n2913 vdd.n865 99.5127
R18266 vdd.n2917 vdd.n865 99.5127
R18267 vdd.n2917 vdd.n856 99.5127
R18268 vdd.n2927 vdd.n856 99.5127
R18269 vdd.n2927 vdd.n854 99.5127
R18270 vdd.n2931 vdd.n854 99.5127
R18271 vdd.n2931 vdd.n842 99.5127
R18272 vdd.n2984 vdd.n842 99.5127
R18273 vdd.n2984 vdd.n840 99.5127
R18274 vdd.n2988 vdd.n840 99.5127
R18275 vdd.n2988 vdd.n808 99.5127
R18276 vdd.n3058 vdd.n808 99.5127
R18277 vdd.n3054 vdd.n809 99.5127
R18278 vdd.n3052 vdd.n3051 99.5127
R18279 vdd.n3049 vdd.n813 99.5127
R18280 vdd.n3045 vdd.n3044 99.5127
R18281 vdd.n3042 vdd.n816 99.5127
R18282 vdd.n3038 vdd.n3037 99.5127
R18283 vdd.n3035 vdd.n819 99.5127
R18284 vdd.n3031 vdd.n3030 99.5127
R18285 vdd.n3028 vdd.n3026 99.5127
R18286 vdd.n3024 vdd.n822 99.5127
R18287 vdd.n3020 vdd.n3019 99.5127
R18288 vdd.n3017 vdd.n825 99.5127
R18289 vdd.n3013 vdd.n3012 99.5127
R18290 vdd.n3010 vdd.n828 99.5127
R18291 vdd.n3006 vdd.n3005 99.5127
R18292 vdd.n3003 vdd.n831 99.5127
R18293 vdd.n2998 vdd.n2997 99.5127
R18294 vdd.n2785 vdd.n914 99.5127
R18295 vdd.n2785 vdd.n909 99.5127
R18296 vdd.n2782 vdd.n909 99.5127
R18297 vdd.n2782 vdd.n904 99.5127
R18298 vdd.n2729 vdd.n904 99.5127
R18299 vdd.n2729 vdd.n898 99.5127
R18300 vdd.n2732 vdd.n898 99.5127
R18301 vdd.n2732 vdd.n891 99.5127
R18302 vdd.n2735 vdd.n891 99.5127
R18303 vdd.n2735 vdd.n886 99.5127
R18304 vdd.n2738 vdd.n886 99.5127
R18305 vdd.n2738 vdd.n881 99.5127
R18306 vdd.n2741 vdd.n881 99.5127
R18307 vdd.n2741 vdd.n875 99.5127
R18308 vdd.n2759 vdd.n875 99.5127
R18309 vdd.n2759 vdd.n868 99.5127
R18310 vdd.n2755 vdd.n868 99.5127
R18311 vdd.n2755 vdd.n863 99.5127
R18312 vdd.n2752 vdd.n863 99.5127
R18313 vdd.n2752 vdd.n858 99.5127
R18314 vdd.n2749 vdd.n858 99.5127
R18315 vdd.n2749 vdd.n852 99.5127
R18316 vdd.n2746 vdd.n852 99.5127
R18317 vdd.n2746 vdd.n844 99.5127
R18318 vdd.n844 vdd.n837 99.5127
R18319 vdd.n2990 vdd.n837 99.5127
R18320 vdd.n2991 vdd.n2990 99.5127
R18321 vdd.n2991 vdd.n806 99.5127
R18322 vdd.n2855 vdd.n2638 99.5127
R18323 vdd.n2851 vdd.n2638 99.5127
R18324 vdd.n2849 vdd.n2848 99.5127
R18325 vdd.n2845 vdd.n2844 99.5127
R18326 vdd.n2841 vdd.n2840 99.5127
R18327 vdd.n2837 vdd.n2836 99.5127
R18328 vdd.n2833 vdd.n2832 99.5127
R18329 vdd.n2829 vdd.n2828 99.5127
R18330 vdd.n2825 vdd.n2824 99.5127
R18331 vdd.n2821 vdd.n2820 99.5127
R18332 vdd.n2817 vdd.n2816 99.5127
R18333 vdd.n2813 vdd.n2812 99.5127
R18334 vdd.n2809 vdd.n2808 99.5127
R18335 vdd.n2805 vdd.n2804 99.5127
R18336 vdd.n2801 vdd.n2800 99.5127
R18337 vdd.n2797 vdd.n2796 99.5127
R18338 vdd.n2792 vdd.n2791 99.5127
R18339 vdd.n2603 vdd.n955 99.5127
R18340 vdd.n2599 vdd.n2598 99.5127
R18341 vdd.n2595 vdd.n2594 99.5127
R18342 vdd.n2591 vdd.n2590 99.5127
R18343 vdd.n2587 vdd.n2586 99.5127
R18344 vdd.n2583 vdd.n2582 99.5127
R18345 vdd.n2579 vdd.n2578 99.5127
R18346 vdd.n2575 vdd.n2574 99.5127
R18347 vdd.n2571 vdd.n2570 99.5127
R18348 vdd.n2567 vdd.n2566 99.5127
R18349 vdd.n2563 vdd.n2562 99.5127
R18350 vdd.n2559 vdd.n2558 99.5127
R18351 vdd.n2555 vdd.n2554 99.5127
R18352 vdd.n2551 vdd.n2550 99.5127
R18353 vdd.n2547 vdd.n2546 99.5127
R18354 vdd.n2543 vdd.n2542 99.5127
R18355 vdd.n2538 vdd.n2537 99.5127
R18356 vdd.n2276 vdd.n1050 99.5127
R18357 vdd.n2276 vdd.n1044 99.5127
R18358 vdd.n2273 vdd.n1044 99.5127
R18359 vdd.n2273 vdd.n1038 99.5127
R18360 vdd.n2270 vdd.n1038 99.5127
R18361 vdd.n2270 vdd.n1031 99.5127
R18362 vdd.n2267 vdd.n1031 99.5127
R18363 vdd.n2267 vdd.n1024 99.5127
R18364 vdd.n2264 vdd.n1024 99.5127
R18365 vdd.n2264 vdd.n1019 99.5127
R18366 vdd.n2261 vdd.n1019 99.5127
R18367 vdd.n2261 vdd.n1013 99.5127
R18368 vdd.n2258 vdd.n1013 99.5127
R18369 vdd.n2258 vdd.n1006 99.5127
R18370 vdd.n2172 vdd.n1006 99.5127
R18371 vdd.n2172 vdd.n1000 99.5127
R18372 vdd.n2169 vdd.n1000 99.5127
R18373 vdd.n2169 vdd.n995 99.5127
R18374 vdd.n2166 vdd.n995 99.5127
R18375 vdd.n2166 vdd.n990 99.5127
R18376 vdd.n2163 vdd.n990 99.5127
R18377 vdd.n2163 vdd.n984 99.5127
R18378 vdd.n2160 vdd.n984 99.5127
R18379 vdd.n2160 vdd.n977 99.5127
R18380 vdd.n2157 vdd.n977 99.5127
R18381 vdd.n2157 vdd.n970 99.5127
R18382 vdd.n970 vdd.n960 99.5127
R18383 vdd.n2533 vdd.n960 99.5127
R18384 vdd.n2111 vdd.n2109 99.5127
R18385 vdd.n2115 vdd.n2109 99.5127
R18386 vdd.n2119 vdd.n2117 99.5127
R18387 vdd.n2123 vdd.n2107 99.5127
R18388 vdd.n2127 vdd.n2125 99.5127
R18389 vdd.n2131 vdd.n2105 99.5127
R18390 vdd.n2135 vdd.n2133 99.5127
R18391 vdd.n2139 vdd.n2103 99.5127
R18392 vdd.n2142 vdd.n2141 99.5127
R18393 vdd.n2312 vdd.n2310 99.5127
R18394 vdd.n2308 vdd.n2144 99.5127
R18395 vdd.n2304 vdd.n2302 99.5127
R18396 vdd.n2300 vdd.n2146 99.5127
R18397 vdd.n2296 vdd.n2294 99.5127
R18398 vdd.n2292 vdd.n2148 99.5127
R18399 vdd.n2288 vdd.n2286 99.5127
R18400 vdd.n2284 vdd.n2150 99.5127
R18401 vdd.n2376 vdd.n1046 99.5127
R18402 vdd.n2380 vdd.n1046 99.5127
R18403 vdd.n2380 vdd.n1036 99.5127
R18404 vdd.n2388 vdd.n1036 99.5127
R18405 vdd.n2388 vdd.n1034 99.5127
R18406 vdd.n2392 vdd.n1034 99.5127
R18407 vdd.n2392 vdd.n1023 99.5127
R18408 vdd.n2401 vdd.n1023 99.5127
R18409 vdd.n2401 vdd.n1021 99.5127
R18410 vdd.n2405 vdd.n1021 99.5127
R18411 vdd.n2405 vdd.n1011 99.5127
R18412 vdd.n2413 vdd.n1011 99.5127
R18413 vdd.n2413 vdd.n1009 99.5127
R18414 vdd.n2417 vdd.n1009 99.5127
R18415 vdd.n2417 vdd.n999 99.5127
R18416 vdd.n2425 vdd.n999 99.5127
R18417 vdd.n2425 vdd.n997 99.5127
R18418 vdd.n2429 vdd.n997 99.5127
R18419 vdd.n2429 vdd.n988 99.5127
R18420 vdd.n2437 vdd.n988 99.5127
R18421 vdd.n2437 vdd.n986 99.5127
R18422 vdd.n2441 vdd.n986 99.5127
R18423 vdd.n2441 vdd.n975 99.5127
R18424 vdd.n2451 vdd.n975 99.5127
R18425 vdd.n2451 vdd.n972 99.5127
R18426 vdd.n2456 vdd.n972 99.5127
R18427 vdd.n2456 vdd.n973 99.5127
R18428 vdd.n973 vdd.n954 99.5127
R18429 vdd.n2974 vdd.n2973 99.5127
R18430 vdd.n2971 vdd.n2937 99.5127
R18431 vdd.n2967 vdd.n2966 99.5127
R18432 vdd.n2964 vdd.n2940 99.5127
R18433 vdd.n2960 vdd.n2959 99.5127
R18434 vdd.n2957 vdd.n2943 99.5127
R18435 vdd.n2953 vdd.n2952 99.5127
R18436 vdd.n2950 vdd.n2947 99.5127
R18437 vdd.n3091 vdd.n787 99.5127
R18438 vdd.n3089 vdd.n3088 99.5127
R18439 vdd.n3086 vdd.n789 99.5127
R18440 vdd.n3082 vdd.n3081 99.5127
R18441 vdd.n3079 vdd.n792 99.5127
R18442 vdd.n3075 vdd.n3074 99.5127
R18443 vdd.n3072 vdd.n795 99.5127
R18444 vdd.n3068 vdd.n3067 99.5127
R18445 vdd.n3065 vdd.n798 99.5127
R18446 vdd.n2709 vdd.n915 99.5127
R18447 vdd.n2709 vdd.n910 99.5127
R18448 vdd.n2780 vdd.n910 99.5127
R18449 vdd.n2780 vdd.n905 99.5127
R18450 vdd.n2776 vdd.n905 99.5127
R18451 vdd.n2776 vdd.n899 99.5127
R18452 vdd.n2773 vdd.n899 99.5127
R18453 vdd.n2773 vdd.n892 99.5127
R18454 vdd.n2770 vdd.n892 99.5127
R18455 vdd.n2770 vdd.n887 99.5127
R18456 vdd.n2767 vdd.n887 99.5127
R18457 vdd.n2767 vdd.n882 99.5127
R18458 vdd.n2764 vdd.n882 99.5127
R18459 vdd.n2764 vdd.n876 99.5127
R18460 vdd.n2761 vdd.n876 99.5127
R18461 vdd.n2761 vdd.n869 99.5127
R18462 vdd.n2726 vdd.n869 99.5127
R18463 vdd.n2726 vdd.n864 99.5127
R18464 vdd.n2723 vdd.n864 99.5127
R18465 vdd.n2723 vdd.n859 99.5127
R18466 vdd.n2720 vdd.n859 99.5127
R18467 vdd.n2720 vdd.n853 99.5127
R18468 vdd.n2717 vdd.n853 99.5127
R18469 vdd.n2717 vdd.n845 99.5127
R18470 vdd.n2714 vdd.n845 99.5127
R18471 vdd.n2714 vdd.n838 99.5127
R18472 vdd.n838 vdd.n804 99.5127
R18473 vdd.n3060 vdd.n804 99.5127
R18474 vdd.n2859 vdd.n918 99.5127
R18475 vdd.n2647 vdd.n2646 99.5127
R18476 vdd.n2651 vdd.n2650 99.5127
R18477 vdd.n2655 vdd.n2654 99.5127
R18478 vdd.n2659 vdd.n2658 99.5127
R18479 vdd.n2663 vdd.n2662 99.5127
R18480 vdd.n2667 vdd.n2666 99.5127
R18481 vdd.n2671 vdd.n2670 99.5127
R18482 vdd.n2675 vdd.n2674 99.5127
R18483 vdd.n2679 vdd.n2678 99.5127
R18484 vdd.n2683 vdd.n2682 99.5127
R18485 vdd.n2687 vdd.n2686 99.5127
R18486 vdd.n2691 vdd.n2690 99.5127
R18487 vdd.n2695 vdd.n2694 99.5127
R18488 vdd.n2699 vdd.n2698 99.5127
R18489 vdd.n2703 vdd.n2702 99.5127
R18490 vdd.n2705 vdd.n2637 99.5127
R18491 vdd.n2863 vdd.n908 99.5127
R18492 vdd.n2871 vdd.n908 99.5127
R18493 vdd.n2871 vdd.n906 99.5127
R18494 vdd.n2875 vdd.n906 99.5127
R18495 vdd.n2875 vdd.n896 99.5127
R18496 vdd.n2883 vdd.n896 99.5127
R18497 vdd.n2883 vdd.n894 99.5127
R18498 vdd.n2887 vdd.n894 99.5127
R18499 vdd.n2887 vdd.n885 99.5127
R18500 vdd.n2895 vdd.n885 99.5127
R18501 vdd.n2895 vdd.n883 99.5127
R18502 vdd.n2899 vdd.n883 99.5127
R18503 vdd.n2899 vdd.n873 99.5127
R18504 vdd.n2907 vdd.n873 99.5127
R18505 vdd.n2907 vdd.n871 99.5127
R18506 vdd.n2911 vdd.n871 99.5127
R18507 vdd.n2911 vdd.n862 99.5127
R18508 vdd.n2919 vdd.n862 99.5127
R18509 vdd.n2919 vdd.n860 99.5127
R18510 vdd.n2925 vdd.n860 99.5127
R18511 vdd.n2925 vdd.n850 99.5127
R18512 vdd.n2933 vdd.n850 99.5127
R18513 vdd.n2933 vdd.n847 99.5127
R18514 vdd.n2982 vdd.n847 99.5127
R18515 vdd.n2982 vdd.n848 99.5127
R18516 vdd.n848 vdd.n839 99.5127
R18517 vdd.n2977 vdd.n839 99.5127
R18518 vdd.n2977 vdd.n807 99.5127
R18519 vdd.n2527 vdd.n2526 99.5127
R18520 vdd.n2523 vdd.n2522 99.5127
R18521 vdd.n2519 vdd.n2518 99.5127
R18522 vdd.n2515 vdd.n2514 99.5127
R18523 vdd.n2511 vdd.n2510 99.5127
R18524 vdd.n2507 vdd.n2506 99.5127
R18525 vdd.n2503 vdd.n2502 99.5127
R18526 vdd.n2499 vdd.n2498 99.5127
R18527 vdd.n2495 vdd.n2494 99.5127
R18528 vdd.n2491 vdd.n2490 99.5127
R18529 vdd.n2487 vdd.n2486 99.5127
R18530 vdd.n2483 vdd.n2482 99.5127
R18531 vdd.n2479 vdd.n2478 99.5127
R18532 vdd.n2475 vdd.n2474 99.5127
R18533 vdd.n2471 vdd.n2470 99.5127
R18534 vdd.n2467 vdd.n2466 99.5127
R18535 vdd.n2463 vdd.n936 99.5127
R18536 vdd.n2220 vdd.n1051 99.5127
R18537 vdd.n2220 vdd.n1045 99.5127
R18538 vdd.n2223 vdd.n1045 99.5127
R18539 vdd.n2223 vdd.n1039 99.5127
R18540 vdd.n2226 vdd.n1039 99.5127
R18541 vdd.n2226 vdd.n1032 99.5127
R18542 vdd.n2229 vdd.n1032 99.5127
R18543 vdd.n2229 vdd.n1025 99.5127
R18544 vdd.n2232 vdd.n1025 99.5127
R18545 vdd.n2232 vdd.n1020 99.5127
R18546 vdd.n2235 vdd.n1020 99.5127
R18547 vdd.n2235 vdd.n1014 99.5127
R18548 vdd.n2256 vdd.n1014 99.5127
R18549 vdd.n2256 vdd.n1007 99.5127
R18550 vdd.n2252 vdd.n1007 99.5127
R18551 vdd.n2252 vdd.n1001 99.5127
R18552 vdd.n2249 vdd.n1001 99.5127
R18553 vdd.n2249 vdd.n996 99.5127
R18554 vdd.n2246 vdd.n996 99.5127
R18555 vdd.n2246 vdd.n991 99.5127
R18556 vdd.n2243 vdd.n991 99.5127
R18557 vdd.n2243 vdd.n985 99.5127
R18558 vdd.n2240 vdd.n985 99.5127
R18559 vdd.n2240 vdd.n978 99.5127
R18560 vdd.n978 vdd.n969 99.5127
R18561 vdd.n2458 vdd.n969 99.5127
R18562 vdd.n2459 vdd.n2458 99.5127
R18563 vdd.n2459 vdd.n961 99.5127
R18564 vdd.n2370 vdd.n2368 99.5127
R18565 vdd.n2366 vdd.n1054 99.5127
R18566 vdd.n2362 vdd.n2360 99.5127
R18567 vdd.n2358 vdd.n1056 99.5127
R18568 vdd.n2354 vdd.n2352 99.5127
R18569 vdd.n2350 vdd.n1058 99.5127
R18570 vdd.n2346 vdd.n2344 99.5127
R18571 vdd.n2342 vdd.n1060 99.5127
R18572 vdd.n2184 vdd.n1062 99.5127
R18573 vdd.n2189 vdd.n2186 99.5127
R18574 vdd.n2193 vdd.n2191 99.5127
R18575 vdd.n2197 vdd.n2182 99.5127
R18576 vdd.n2201 vdd.n2199 99.5127
R18577 vdd.n2205 vdd.n2180 99.5127
R18578 vdd.n2209 vdd.n2207 99.5127
R18579 vdd.n2214 vdd.n2176 99.5127
R18580 vdd.n2217 vdd.n2216 99.5127
R18581 vdd.n2374 vdd.n1042 99.5127
R18582 vdd.n2382 vdd.n1042 99.5127
R18583 vdd.n2382 vdd.n1040 99.5127
R18584 vdd.n2386 vdd.n1040 99.5127
R18585 vdd.n2386 vdd.n1029 99.5127
R18586 vdd.n2394 vdd.n1029 99.5127
R18587 vdd.n2394 vdd.n1026 99.5127
R18588 vdd.n2399 vdd.n1026 99.5127
R18589 vdd.n2399 vdd.n1017 99.5127
R18590 vdd.n2407 vdd.n1017 99.5127
R18591 vdd.n2407 vdd.n1015 99.5127
R18592 vdd.n2411 vdd.n1015 99.5127
R18593 vdd.n2411 vdd.n1005 99.5127
R18594 vdd.n2419 vdd.n1005 99.5127
R18595 vdd.n2419 vdd.n1003 99.5127
R18596 vdd.n2423 vdd.n1003 99.5127
R18597 vdd.n2423 vdd.n994 99.5127
R18598 vdd.n2431 vdd.n994 99.5127
R18599 vdd.n2431 vdd.n992 99.5127
R18600 vdd.n2435 vdd.n992 99.5127
R18601 vdd.n2435 vdd.n982 99.5127
R18602 vdd.n2443 vdd.n982 99.5127
R18603 vdd.n2443 vdd.n979 99.5127
R18604 vdd.n2449 vdd.n979 99.5127
R18605 vdd.n2449 vdd.n980 99.5127
R18606 vdd.n980 vdd.n971 99.5127
R18607 vdd.n971 vdd.n962 99.5127
R18608 vdd.n2531 vdd.n962 99.5127
R18609 vdd.n9 vdd.n7 98.9633
R18610 vdd.n2 vdd.n0 98.9633
R18611 vdd.n9 vdd.n8 98.6055
R18612 vdd.n11 vdd.n10 98.6055
R18613 vdd.n13 vdd.n12 98.6055
R18614 vdd.n6 vdd.n5 98.6055
R18615 vdd.n4 vdd.n3 98.6055
R18616 vdd.n2 vdd.n1 98.6055
R18617 vdd.t141 vdd.n303 85.8723
R18618 vdd.t115 vdd.n244 85.8723
R18619 vdd.t128 vdd.n201 85.8723
R18620 vdd.t101 vdd.n142 85.8723
R18621 vdd.t80 vdd.n100 85.8723
R18622 vdd.t14 vdd.n41 85.8723
R18623 vdd.t160 vdd.n1722 85.8723
R18624 vdd.t47 vdd.n1781 85.8723
R18625 vdd.t146 vdd.n1620 85.8723
R18626 vdd.t22 vdd.n1679 85.8723
R18627 vdd.t18 vdd.n1519 85.8723
R18628 vdd.t81 vdd.n1578 85.8723
R18629 vdd.n2923 vdd.n2922 78.546
R18630 vdd.n2397 vdd.n1027 78.546
R18631 vdd.n290 vdd.n289 75.1835
R18632 vdd.n288 vdd.n287 75.1835
R18633 vdd.n286 vdd.n285 75.1835
R18634 vdd.n284 vdd.n283 75.1835
R18635 vdd.n282 vdd.n281 75.1835
R18636 vdd.n280 vdd.n279 75.1835
R18637 vdd.n278 vdd.n277 75.1835
R18638 vdd.n276 vdd.n275 75.1835
R18639 vdd.n274 vdd.n273 75.1835
R18640 vdd.n188 vdd.n187 75.1835
R18641 vdd.n186 vdd.n185 75.1835
R18642 vdd.n184 vdd.n183 75.1835
R18643 vdd.n182 vdd.n181 75.1835
R18644 vdd.n180 vdd.n179 75.1835
R18645 vdd.n178 vdd.n177 75.1835
R18646 vdd.n176 vdd.n175 75.1835
R18647 vdd.n174 vdd.n173 75.1835
R18648 vdd.n172 vdd.n171 75.1835
R18649 vdd.n87 vdd.n86 75.1835
R18650 vdd.n85 vdd.n84 75.1835
R18651 vdd.n83 vdd.n82 75.1835
R18652 vdd.n81 vdd.n80 75.1835
R18653 vdd.n79 vdd.n78 75.1835
R18654 vdd.n77 vdd.n76 75.1835
R18655 vdd.n75 vdd.n74 75.1835
R18656 vdd.n73 vdd.n72 75.1835
R18657 vdd.n71 vdd.n70 75.1835
R18658 vdd.n1752 vdd.n1751 75.1835
R18659 vdd.n1754 vdd.n1753 75.1835
R18660 vdd.n1756 vdd.n1755 75.1835
R18661 vdd.n1758 vdd.n1757 75.1835
R18662 vdd.n1760 vdd.n1759 75.1835
R18663 vdd.n1762 vdd.n1761 75.1835
R18664 vdd.n1764 vdd.n1763 75.1835
R18665 vdd.n1766 vdd.n1765 75.1835
R18666 vdd.n1768 vdd.n1767 75.1835
R18667 vdd.n1650 vdd.n1649 75.1835
R18668 vdd.n1652 vdd.n1651 75.1835
R18669 vdd.n1654 vdd.n1653 75.1835
R18670 vdd.n1656 vdd.n1655 75.1835
R18671 vdd.n1658 vdd.n1657 75.1835
R18672 vdd.n1660 vdd.n1659 75.1835
R18673 vdd.n1662 vdd.n1661 75.1835
R18674 vdd.n1664 vdd.n1663 75.1835
R18675 vdd.n1666 vdd.n1665 75.1835
R18676 vdd.n1549 vdd.n1548 75.1835
R18677 vdd.n1551 vdd.n1550 75.1835
R18678 vdd.n1553 vdd.n1552 75.1835
R18679 vdd.n1555 vdd.n1554 75.1835
R18680 vdd.n1557 vdd.n1556 75.1835
R18681 vdd.n1559 vdd.n1558 75.1835
R18682 vdd.n1561 vdd.n1560 75.1835
R18683 vdd.n1563 vdd.n1562 75.1835
R18684 vdd.n1565 vdd.n1564 75.1835
R18685 vdd.n2858 vdd.n2857 72.8958
R18686 vdd.n2857 vdd.n2621 72.8958
R18687 vdd.n2857 vdd.n2622 72.8958
R18688 vdd.n2857 vdd.n2623 72.8958
R18689 vdd.n2857 vdd.n2624 72.8958
R18690 vdd.n2857 vdd.n2625 72.8958
R18691 vdd.n2857 vdd.n2626 72.8958
R18692 vdd.n2857 vdd.n2627 72.8958
R18693 vdd.n2857 vdd.n2628 72.8958
R18694 vdd.n2857 vdd.n2629 72.8958
R18695 vdd.n2857 vdd.n2630 72.8958
R18696 vdd.n2857 vdd.n2631 72.8958
R18697 vdd.n2857 vdd.n2632 72.8958
R18698 vdd.n2857 vdd.n2633 72.8958
R18699 vdd.n2857 vdd.n2634 72.8958
R18700 vdd.n2857 vdd.n2635 72.8958
R18701 vdd.n2857 vdd.n2636 72.8958
R18702 vdd.n803 vdd.n692 72.8958
R18703 vdd.n3066 vdd.n692 72.8958
R18704 vdd.n797 vdd.n692 72.8958
R18705 vdd.n3073 vdd.n692 72.8958
R18706 vdd.n794 vdd.n692 72.8958
R18707 vdd.n3080 vdd.n692 72.8958
R18708 vdd.n791 vdd.n692 72.8958
R18709 vdd.n3087 vdd.n692 72.8958
R18710 vdd.n3090 vdd.n692 72.8958
R18711 vdd.n2946 vdd.n692 72.8958
R18712 vdd.n2951 vdd.n692 72.8958
R18713 vdd.n2945 vdd.n692 72.8958
R18714 vdd.n2958 vdd.n692 72.8958
R18715 vdd.n2942 vdd.n692 72.8958
R18716 vdd.n2965 vdd.n692 72.8958
R18717 vdd.n2939 vdd.n692 72.8958
R18718 vdd.n2972 vdd.n692 72.8958
R18719 vdd.n2110 vdd.n1049 72.8958
R18720 vdd.n2116 vdd.n1049 72.8958
R18721 vdd.n2118 vdd.n1049 72.8958
R18722 vdd.n2124 vdd.n1049 72.8958
R18723 vdd.n2126 vdd.n1049 72.8958
R18724 vdd.n2132 vdd.n1049 72.8958
R18725 vdd.n2134 vdd.n1049 72.8958
R18726 vdd.n2140 vdd.n1049 72.8958
R18727 vdd.n2311 vdd.n1049 72.8958
R18728 vdd.n2309 vdd.n1049 72.8958
R18729 vdd.n2303 vdd.n1049 72.8958
R18730 vdd.n2301 vdd.n1049 72.8958
R18731 vdd.n2295 vdd.n1049 72.8958
R18732 vdd.n2293 vdd.n1049 72.8958
R18733 vdd.n2287 vdd.n1049 72.8958
R18734 vdd.n2285 vdd.n1049 72.8958
R18735 vdd.n2279 vdd.n1049 72.8958
R18736 vdd.n2604 vdd.n937 72.8958
R18737 vdd.n2604 vdd.n938 72.8958
R18738 vdd.n2604 vdd.n939 72.8958
R18739 vdd.n2604 vdd.n940 72.8958
R18740 vdd.n2604 vdd.n941 72.8958
R18741 vdd.n2604 vdd.n942 72.8958
R18742 vdd.n2604 vdd.n943 72.8958
R18743 vdd.n2604 vdd.n944 72.8958
R18744 vdd.n2604 vdd.n945 72.8958
R18745 vdd.n2604 vdd.n946 72.8958
R18746 vdd.n2604 vdd.n947 72.8958
R18747 vdd.n2604 vdd.n948 72.8958
R18748 vdd.n2604 vdd.n949 72.8958
R18749 vdd.n2604 vdd.n950 72.8958
R18750 vdd.n2604 vdd.n951 72.8958
R18751 vdd.n2604 vdd.n952 72.8958
R18752 vdd.n2604 vdd.n953 72.8958
R18753 vdd.n2857 vdd.n2856 72.8958
R18754 vdd.n2857 vdd.n2605 72.8958
R18755 vdd.n2857 vdd.n2606 72.8958
R18756 vdd.n2857 vdd.n2607 72.8958
R18757 vdd.n2857 vdd.n2608 72.8958
R18758 vdd.n2857 vdd.n2609 72.8958
R18759 vdd.n2857 vdd.n2610 72.8958
R18760 vdd.n2857 vdd.n2611 72.8958
R18761 vdd.n2857 vdd.n2612 72.8958
R18762 vdd.n2857 vdd.n2613 72.8958
R18763 vdd.n2857 vdd.n2614 72.8958
R18764 vdd.n2857 vdd.n2615 72.8958
R18765 vdd.n2857 vdd.n2616 72.8958
R18766 vdd.n2857 vdd.n2617 72.8958
R18767 vdd.n2857 vdd.n2618 72.8958
R18768 vdd.n2857 vdd.n2619 72.8958
R18769 vdd.n2857 vdd.n2620 72.8958
R18770 vdd.n2996 vdd.n692 72.8958
R18771 vdd.n835 vdd.n692 72.8958
R18772 vdd.n3004 vdd.n692 72.8958
R18773 vdd.n830 vdd.n692 72.8958
R18774 vdd.n3011 vdd.n692 72.8958
R18775 vdd.n827 vdd.n692 72.8958
R18776 vdd.n3018 vdd.n692 72.8958
R18777 vdd.n824 vdd.n692 72.8958
R18778 vdd.n3025 vdd.n692 72.8958
R18779 vdd.n3029 vdd.n692 72.8958
R18780 vdd.n821 vdd.n692 72.8958
R18781 vdd.n3036 vdd.n692 72.8958
R18782 vdd.n818 vdd.n692 72.8958
R18783 vdd.n3043 vdd.n692 72.8958
R18784 vdd.n815 vdd.n692 72.8958
R18785 vdd.n3050 vdd.n692 72.8958
R18786 vdd.n3053 vdd.n692 72.8958
R18787 vdd.n2604 vdd.n935 72.8958
R18788 vdd.n2604 vdd.n934 72.8958
R18789 vdd.n2604 vdd.n933 72.8958
R18790 vdd.n2604 vdd.n932 72.8958
R18791 vdd.n2604 vdd.n931 72.8958
R18792 vdd.n2604 vdd.n930 72.8958
R18793 vdd.n2604 vdd.n929 72.8958
R18794 vdd.n2604 vdd.n928 72.8958
R18795 vdd.n2604 vdd.n927 72.8958
R18796 vdd.n2604 vdd.n926 72.8958
R18797 vdd.n2604 vdd.n925 72.8958
R18798 vdd.n2604 vdd.n924 72.8958
R18799 vdd.n2604 vdd.n923 72.8958
R18800 vdd.n2604 vdd.n922 72.8958
R18801 vdd.n2604 vdd.n921 72.8958
R18802 vdd.n2604 vdd.n920 72.8958
R18803 vdd.n2604 vdd.n919 72.8958
R18804 vdd.n2369 vdd.n1049 72.8958
R18805 vdd.n2367 vdd.n1049 72.8958
R18806 vdd.n2361 vdd.n1049 72.8958
R18807 vdd.n2359 vdd.n1049 72.8958
R18808 vdd.n2353 vdd.n1049 72.8958
R18809 vdd.n2351 vdd.n1049 72.8958
R18810 vdd.n2345 vdd.n1049 72.8958
R18811 vdd.n2343 vdd.n1049 72.8958
R18812 vdd.n1061 vdd.n1049 72.8958
R18813 vdd.n2185 vdd.n1049 72.8958
R18814 vdd.n2190 vdd.n1049 72.8958
R18815 vdd.n2192 vdd.n1049 72.8958
R18816 vdd.n2198 vdd.n1049 72.8958
R18817 vdd.n2200 vdd.n1049 72.8958
R18818 vdd.n2206 vdd.n1049 72.8958
R18819 vdd.n2208 vdd.n1049 72.8958
R18820 vdd.n2215 vdd.n1049 72.8958
R18821 vdd.n1419 vdd.n1418 66.2847
R18822 vdd.n1418 vdd.n1194 66.2847
R18823 vdd.n1418 vdd.n1195 66.2847
R18824 vdd.n1418 vdd.n1196 66.2847
R18825 vdd.n1418 vdd.n1197 66.2847
R18826 vdd.n1418 vdd.n1198 66.2847
R18827 vdd.n1418 vdd.n1199 66.2847
R18828 vdd.n1418 vdd.n1200 66.2847
R18829 vdd.n1418 vdd.n1201 66.2847
R18830 vdd.n1418 vdd.n1202 66.2847
R18831 vdd.n1418 vdd.n1203 66.2847
R18832 vdd.n1418 vdd.n1204 66.2847
R18833 vdd.n1418 vdd.n1205 66.2847
R18834 vdd.n1418 vdd.n1206 66.2847
R18835 vdd.n1418 vdd.n1207 66.2847
R18836 vdd.n1418 vdd.n1208 66.2847
R18837 vdd.n1418 vdd.n1209 66.2847
R18838 vdd.n1418 vdd.n1210 66.2847
R18839 vdd.n1418 vdd.n1211 66.2847
R18840 vdd.n1418 vdd.n1212 66.2847
R18841 vdd.n1418 vdd.n1213 66.2847
R18842 vdd.n1418 vdd.n1214 66.2847
R18843 vdd.n1418 vdd.n1215 66.2847
R18844 vdd.n1418 vdd.n1216 66.2847
R18845 vdd.n1418 vdd.n1217 66.2847
R18846 vdd.n1418 vdd.n1218 66.2847
R18847 vdd.n1418 vdd.n1219 66.2847
R18848 vdd.n1418 vdd.n1220 66.2847
R18849 vdd.n1418 vdd.n1221 66.2847
R18850 vdd.n1418 vdd.n1222 66.2847
R18851 vdd.n1418 vdd.n1223 66.2847
R18852 vdd.n1073 vdd.n1070 66.2847
R18853 vdd.n2000 vdd.n1073 66.2847
R18854 vdd.n2005 vdd.n1073 66.2847
R18855 vdd.n2010 vdd.n1073 66.2847
R18856 vdd.n1998 vdd.n1073 66.2847
R18857 vdd.n2017 vdd.n1073 66.2847
R18858 vdd.n1990 vdd.n1073 66.2847
R18859 vdd.n2024 vdd.n1073 66.2847
R18860 vdd.n1983 vdd.n1073 66.2847
R18861 vdd.n2031 vdd.n1073 66.2847
R18862 vdd.n1977 vdd.n1073 66.2847
R18863 vdd.n1972 vdd.n1073 66.2847
R18864 vdd.n2042 vdd.n1073 66.2847
R18865 vdd.n1964 vdd.n1073 66.2847
R18866 vdd.n2049 vdd.n1073 66.2847
R18867 vdd.n1957 vdd.n1073 66.2847
R18868 vdd.n2056 vdd.n1073 66.2847
R18869 vdd.n1950 vdd.n1073 66.2847
R18870 vdd.n2063 vdd.n1073 66.2847
R18871 vdd.n1943 vdd.n1073 66.2847
R18872 vdd.n2070 vdd.n1073 66.2847
R18873 vdd.n1937 vdd.n1073 66.2847
R18874 vdd.n1932 vdd.n1073 66.2847
R18875 vdd.n2081 vdd.n1073 66.2847
R18876 vdd.n1924 vdd.n1073 66.2847
R18877 vdd.n2088 vdd.n1073 66.2847
R18878 vdd.n1917 vdd.n1073 66.2847
R18879 vdd.n2095 vdd.n1073 66.2847
R18880 vdd.n2098 vdd.n1073 66.2847
R18881 vdd.n1908 vdd.n1073 66.2847
R18882 vdd.n2320 vdd.n1073 66.2847
R18883 vdd.n1902 vdd.n1073 66.2847
R18884 vdd.n3223 vdd.n3222 66.2847
R18885 vdd.n3223 vdd.n693 66.2847
R18886 vdd.n3223 vdd.n694 66.2847
R18887 vdd.n3223 vdd.n695 66.2847
R18888 vdd.n3223 vdd.n696 66.2847
R18889 vdd.n3223 vdd.n697 66.2847
R18890 vdd.n3223 vdd.n698 66.2847
R18891 vdd.n3223 vdd.n699 66.2847
R18892 vdd.n3223 vdd.n700 66.2847
R18893 vdd.n3223 vdd.n701 66.2847
R18894 vdd.n3223 vdd.n702 66.2847
R18895 vdd.n3223 vdd.n703 66.2847
R18896 vdd.n3223 vdd.n704 66.2847
R18897 vdd.n3223 vdd.n705 66.2847
R18898 vdd.n3223 vdd.n706 66.2847
R18899 vdd.n3223 vdd.n707 66.2847
R18900 vdd.n3223 vdd.n708 66.2847
R18901 vdd.n3223 vdd.n709 66.2847
R18902 vdd.n3223 vdd.n710 66.2847
R18903 vdd.n3223 vdd.n711 66.2847
R18904 vdd.n3223 vdd.n712 66.2847
R18905 vdd.n3223 vdd.n713 66.2847
R18906 vdd.n3223 vdd.n714 66.2847
R18907 vdd.n3223 vdd.n715 66.2847
R18908 vdd.n3223 vdd.n716 66.2847
R18909 vdd.n3223 vdd.n717 66.2847
R18910 vdd.n3223 vdd.n718 66.2847
R18911 vdd.n3223 vdd.n719 66.2847
R18912 vdd.n3223 vdd.n720 66.2847
R18913 vdd.n3223 vdd.n721 66.2847
R18914 vdd.n3223 vdd.n722 66.2847
R18915 vdd.n3354 vdd.n3353 66.2847
R18916 vdd.n3354 vdd.n424 66.2847
R18917 vdd.n3354 vdd.n423 66.2847
R18918 vdd.n3354 vdd.n422 66.2847
R18919 vdd.n3354 vdd.n421 66.2847
R18920 vdd.n3354 vdd.n420 66.2847
R18921 vdd.n3354 vdd.n419 66.2847
R18922 vdd.n3354 vdd.n418 66.2847
R18923 vdd.n3354 vdd.n417 66.2847
R18924 vdd.n3354 vdd.n416 66.2847
R18925 vdd.n3354 vdd.n415 66.2847
R18926 vdd.n3354 vdd.n414 66.2847
R18927 vdd.n3354 vdd.n413 66.2847
R18928 vdd.n3354 vdd.n412 66.2847
R18929 vdd.n3354 vdd.n411 66.2847
R18930 vdd.n3354 vdd.n410 66.2847
R18931 vdd.n3354 vdd.n409 66.2847
R18932 vdd.n3354 vdd.n408 66.2847
R18933 vdd.n3354 vdd.n407 66.2847
R18934 vdd.n3354 vdd.n406 66.2847
R18935 vdd.n3354 vdd.n405 66.2847
R18936 vdd.n3354 vdd.n404 66.2847
R18937 vdd.n3354 vdd.n403 66.2847
R18938 vdd.n3354 vdd.n402 66.2847
R18939 vdd.n3354 vdd.n401 66.2847
R18940 vdd.n3354 vdd.n400 66.2847
R18941 vdd.n3354 vdd.n399 66.2847
R18942 vdd.n3354 vdd.n398 66.2847
R18943 vdd.n3354 vdd.n397 66.2847
R18944 vdd.n3354 vdd.n396 66.2847
R18945 vdd.n3354 vdd.n395 66.2847
R18946 vdd.n3354 vdd.n394 66.2847
R18947 vdd.n467 vdd.n394 52.4337
R18948 vdd.n473 vdd.n395 52.4337
R18949 vdd.n477 vdd.n396 52.4337
R18950 vdd.n483 vdd.n397 52.4337
R18951 vdd.n487 vdd.n398 52.4337
R18952 vdd.n493 vdd.n399 52.4337
R18953 vdd.n497 vdd.n400 52.4337
R18954 vdd.n503 vdd.n401 52.4337
R18955 vdd.n507 vdd.n402 52.4337
R18956 vdd.n513 vdd.n403 52.4337
R18957 vdd.n517 vdd.n404 52.4337
R18958 vdd.n523 vdd.n405 52.4337
R18959 vdd.n527 vdd.n406 52.4337
R18960 vdd.n533 vdd.n407 52.4337
R18961 vdd.n537 vdd.n408 52.4337
R18962 vdd.n543 vdd.n409 52.4337
R18963 vdd.n547 vdd.n410 52.4337
R18964 vdd.n553 vdd.n411 52.4337
R18965 vdd.n557 vdd.n412 52.4337
R18966 vdd.n563 vdd.n413 52.4337
R18967 vdd.n567 vdd.n414 52.4337
R18968 vdd.n573 vdd.n415 52.4337
R18969 vdd.n577 vdd.n416 52.4337
R18970 vdd.n583 vdd.n417 52.4337
R18971 vdd.n587 vdd.n418 52.4337
R18972 vdd.n593 vdd.n419 52.4337
R18973 vdd.n597 vdd.n420 52.4337
R18974 vdd.n603 vdd.n421 52.4337
R18975 vdd.n607 vdd.n422 52.4337
R18976 vdd.n613 vdd.n423 52.4337
R18977 vdd.n616 vdd.n424 52.4337
R18978 vdd.n3353 vdd.n3352 52.4337
R18979 vdd.n3222 vdd.n3221 52.4337
R18980 vdd.n728 vdd.n693 52.4337
R18981 vdd.n734 vdd.n694 52.4337
R18982 vdd.n3211 vdd.n695 52.4337
R18983 vdd.n3207 vdd.n696 52.4337
R18984 vdd.n3203 vdd.n697 52.4337
R18985 vdd.n3199 vdd.n698 52.4337
R18986 vdd.n3195 vdd.n699 52.4337
R18987 vdd.n3191 vdd.n700 52.4337
R18988 vdd.n3187 vdd.n701 52.4337
R18989 vdd.n3179 vdd.n702 52.4337
R18990 vdd.n3175 vdd.n703 52.4337
R18991 vdd.n3171 vdd.n704 52.4337
R18992 vdd.n3167 vdd.n705 52.4337
R18993 vdd.n3163 vdd.n706 52.4337
R18994 vdd.n3159 vdd.n707 52.4337
R18995 vdd.n3155 vdd.n708 52.4337
R18996 vdd.n3151 vdd.n709 52.4337
R18997 vdd.n3147 vdd.n710 52.4337
R18998 vdd.n3143 vdd.n711 52.4337
R18999 vdd.n3139 vdd.n712 52.4337
R19000 vdd.n3133 vdd.n713 52.4337
R19001 vdd.n3129 vdd.n714 52.4337
R19002 vdd.n3125 vdd.n715 52.4337
R19003 vdd.n3121 vdd.n716 52.4337
R19004 vdd.n3117 vdd.n717 52.4337
R19005 vdd.n3113 vdd.n718 52.4337
R19006 vdd.n3109 vdd.n719 52.4337
R19007 vdd.n3105 vdd.n720 52.4337
R19008 vdd.n3101 vdd.n721 52.4337
R19009 vdd.n3097 vdd.n722 52.4337
R19010 vdd.n2322 vdd.n1902 52.4337
R19011 vdd.n2320 vdd.n2319 52.4337
R19012 vdd.n1909 vdd.n1908 52.4337
R19013 vdd.n2098 vdd.n2097 52.4337
R19014 vdd.n2095 vdd.n2094 52.4337
R19015 vdd.n2090 vdd.n1917 52.4337
R19016 vdd.n2088 vdd.n2087 52.4337
R19017 vdd.n2083 vdd.n1924 52.4337
R19018 vdd.n2081 vdd.n2080 52.4337
R19019 vdd.n1933 vdd.n1932 52.4337
R19020 vdd.n2072 vdd.n1937 52.4337
R19021 vdd.n2070 vdd.n2069 52.4337
R19022 vdd.n2065 vdd.n1943 52.4337
R19023 vdd.n2063 vdd.n2062 52.4337
R19024 vdd.n2058 vdd.n1950 52.4337
R19025 vdd.n2056 vdd.n2055 52.4337
R19026 vdd.n2051 vdd.n1957 52.4337
R19027 vdd.n2049 vdd.n2048 52.4337
R19028 vdd.n2044 vdd.n1964 52.4337
R19029 vdd.n2042 vdd.n2041 52.4337
R19030 vdd.n1973 vdd.n1972 52.4337
R19031 vdd.n2033 vdd.n1977 52.4337
R19032 vdd.n2031 vdd.n2030 52.4337
R19033 vdd.n2026 vdd.n1983 52.4337
R19034 vdd.n2024 vdd.n2023 52.4337
R19035 vdd.n2019 vdd.n1990 52.4337
R19036 vdd.n2017 vdd.n2016 52.4337
R19037 vdd.n2012 vdd.n1998 52.4337
R19038 vdd.n2010 vdd.n2009 52.4337
R19039 vdd.n2005 vdd.n2004 52.4337
R19040 vdd.n2000 vdd.n1999 52.4337
R19041 vdd.n2331 vdd.n1070 52.4337
R19042 vdd.n1420 vdd.n1419 52.4337
R19043 vdd.n1226 vdd.n1194 52.4337
R19044 vdd.n1230 vdd.n1195 52.4337
R19045 vdd.n1232 vdd.n1196 52.4337
R19046 vdd.n1236 vdd.n1197 52.4337
R19047 vdd.n1238 vdd.n1198 52.4337
R19048 vdd.n1242 vdd.n1199 52.4337
R19049 vdd.n1244 vdd.n1200 52.4337
R19050 vdd.n1248 vdd.n1201 52.4337
R19051 vdd.n1250 vdd.n1202 52.4337
R19052 vdd.n1256 vdd.n1203 52.4337
R19053 vdd.n1258 vdd.n1204 52.4337
R19054 vdd.n1262 vdd.n1205 52.4337
R19055 vdd.n1264 vdd.n1206 52.4337
R19056 vdd.n1268 vdd.n1207 52.4337
R19057 vdd.n1270 vdd.n1208 52.4337
R19058 vdd.n1274 vdd.n1209 52.4337
R19059 vdd.n1276 vdd.n1210 52.4337
R19060 vdd.n1280 vdd.n1211 52.4337
R19061 vdd.n1282 vdd.n1212 52.4337
R19062 vdd.n1354 vdd.n1213 52.4337
R19063 vdd.n1287 vdd.n1214 52.4337
R19064 vdd.n1291 vdd.n1215 52.4337
R19065 vdd.n1293 vdd.n1216 52.4337
R19066 vdd.n1297 vdd.n1217 52.4337
R19067 vdd.n1299 vdd.n1218 52.4337
R19068 vdd.n1303 vdd.n1219 52.4337
R19069 vdd.n1305 vdd.n1220 52.4337
R19070 vdd.n1309 vdd.n1221 52.4337
R19071 vdd.n1311 vdd.n1222 52.4337
R19072 vdd.n1315 vdd.n1223 52.4337
R19073 vdd.n1419 vdd.n1193 52.4337
R19074 vdd.n1229 vdd.n1194 52.4337
R19075 vdd.n1231 vdd.n1195 52.4337
R19076 vdd.n1235 vdd.n1196 52.4337
R19077 vdd.n1237 vdd.n1197 52.4337
R19078 vdd.n1241 vdd.n1198 52.4337
R19079 vdd.n1243 vdd.n1199 52.4337
R19080 vdd.n1247 vdd.n1200 52.4337
R19081 vdd.n1249 vdd.n1201 52.4337
R19082 vdd.n1255 vdd.n1202 52.4337
R19083 vdd.n1257 vdd.n1203 52.4337
R19084 vdd.n1261 vdd.n1204 52.4337
R19085 vdd.n1263 vdd.n1205 52.4337
R19086 vdd.n1267 vdd.n1206 52.4337
R19087 vdd.n1269 vdd.n1207 52.4337
R19088 vdd.n1273 vdd.n1208 52.4337
R19089 vdd.n1275 vdd.n1209 52.4337
R19090 vdd.n1279 vdd.n1210 52.4337
R19091 vdd.n1281 vdd.n1211 52.4337
R19092 vdd.n1285 vdd.n1212 52.4337
R19093 vdd.n1286 vdd.n1213 52.4337
R19094 vdd.n1290 vdd.n1214 52.4337
R19095 vdd.n1292 vdd.n1215 52.4337
R19096 vdd.n1296 vdd.n1216 52.4337
R19097 vdd.n1298 vdd.n1217 52.4337
R19098 vdd.n1302 vdd.n1218 52.4337
R19099 vdd.n1304 vdd.n1219 52.4337
R19100 vdd.n1308 vdd.n1220 52.4337
R19101 vdd.n1310 vdd.n1221 52.4337
R19102 vdd.n1314 vdd.n1222 52.4337
R19103 vdd.n1316 vdd.n1223 52.4337
R19104 vdd.n1070 vdd.n1069 52.4337
R19105 vdd.n2001 vdd.n2000 52.4337
R19106 vdd.n2006 vdd.n2005 52.4337
R19107 vdd.n2011 vdd.n2010 52.4337
R19108 vdd.n1998 vdd.n1991 52.4337
R19109 vdd.n2018 vdd.n2017 52.4337
R19110 vdd.n1990 vdd.n1984 52.4337
R19111 vdd.n2025 vdd.n2024 52.4337
R19112 vdd.n1983 vdd.n1978 52.4337
R19113 vdd.n2032 vdd.n2031 52.4337
R19114 vdd.n1977 vdd.n1976 52.4337
R19115 vdd.n1972 vdd.n1965 52.4337
R19116 vdd.n2043 vdd.n2042 52.4337
R19117 vdd.n1964 vdd.n1958 52.4337
R19118 vdd.n2050 vdd.n2049 52.4337
R19119 vdd.n1957 vdd.n1951 52.4337
R19120 vdd.n2057 vdd.n2056 52.4337
R19121 vdd.n1950 vdd.n1944 52.4337
R19122 vdd.n2064 vdd.n2063 52.4337
R19123 vdd.n1943 vdd.n1938 52.4337
R19124 vdd.n2071 vdd.n2070 52.4337
R19125 vdd.n1937 vdd.n1936 52.4337
R19126 vdd.n1932 vdd.n1925 52.4337
R19127 vdd.n2082 vdd.n2081 52.4337
R19128 vdd.n1924 vdd.n1918 52.4337
R19129 vdd.n2089 vdd.n2088 52.4337
R19130 vdd.n1917 vdd.n1911 52.4337
R19131 vdd.n2096 vdd.n2095 52.4337
R19132 vdd.n2099 vdd.n2098 52.4337
R19133 vdd.n1908 vdd.n1903 52.4337
R19134 vdd.n2321 vdd.n2320 52.4337
R19135 vdd.n1902 vdd.n1075 52.4337
R19136 vdd.n3222 vdd.n725 52.4337
R19137 vdd.n733 vdd.n693 52.4337
R19138 vdd.n3212 vdd.n694 52.4337
R19139 vdd.n3208 vdd.n695 52.4337
R19140 vdd.n3204 vdd.n696 52.4337
R19141 vdd.n3200 vdd.n697 52.4337
R19142 vdd.n3196 vdd.n698 52.4337
R19143 vdd.n3192 vdd.n699 52.4337
R19144 vdd.n3188 vdd.n700 52.4337
R19145 vdd.n3178 vdd.n701 52.4337
R19146 vdd.n3176 vdd.n702 52.4337
R19147 vdd.n3172 vdd.n703 52.4337
R19148 vdd.n3168 vdd.n704 52.4337
R19149 vdd.n3164 vdd.n705 52.4337
R19150 vdd.n3160 vdd.n706 52.4337
R19151 vdd.n3156 vdd.n707 52.4337
R19152 vdd.n3152 vdd.n708 52.4337
R19153 vdd.n3148 vdd.n709 52.4337
R19154 vdd.n3144 vdd.n710 52.4337
R19155 vdd.n3140 vdd.n711 52.4337
R19156 vdd.n3132 vdd.n712 52.4337
R19157 vdd.n3130 vdd.n713 52.4337
R19158 vdd.n3126 vdd.n714 52.4337
R19159 vdd.n3122 vdd.n715 52.4337
R19160 vdd.n3118 vdd.n716 52.4337
R19161 vdd.n3114 vdd.n717 52.4337
R19162 vdd.n3110 vdd.n718 52.4337
R19163 vdd.n3106 vdd.n719 52.4337
R19164 vdd.n3102 vdd.n720 52.4337
R19165 vdd.n3098 vdd.n721 52.4337
R19166 vdd.n722 vdd.n691 52.4337
R19167 vdd.n3353 vdd.n425 52.4337
R19168 vdd.n614 vdd.n424 52.4337
R19169 vdd.n608 vdd.n423 52.4337
R19170 vdd.n604 vdd.n422 52.4337
R19171 vdd.n598 vdd.n421 52.4337
R19172 vdd.n594 vdd.n420 52.4337
R19173 vdd.n588 vdd.n419 52.4337
R19174 vdd.n584 vdd.n418 52.4337
R19175 vdd.n578 vdd.n417 52.4337
R19176 vdd.n574 vdd.n416 52.4337
R19177 vdd.n568 vdd.n415 52.4337
R19178 vdd.n564 vdd.n414 52.4337
R19179 vdd.n558 vdd.n413 52.4337
R19180 vdd.n554 vdd.n412 52.4337
R19181 vdd.n548 vdd.n411 52.4337
R19182 vdd.n544 vdd.n410 52.4337
R19183 vdd.n538 vdd.n409 52.4337
R19184 vdd.n534 vdd.n408 52.4337
R19185 vdd.n528 vdd.n407 52.4337
R19186 vdd.n524 vdd.n406 52.4337
R19187 vdd.n518 vdd.n405 52.4337
R19188 vdd.n514 vdd.n404 52.4337
R19189 vdd.n508 vdd.n403 52.4337
R19190 vdd.n504 vdd.n402 52.4337
R19191 vdd.n498 vdd.n401 52.4337
R19192 vdd.n494 vdd.n400 52.4337
R19193 vdd.n488 vdd.n399 52.4337
R19194 vdd.n484 vdd.n398 52.4337
R19195 vdd.n478 vdd.n397 52.4337
R19196 vdd.n474 vdd.n396 52.4337
R19197 vdd.n468 vdd.n395 52.4337
R19198 vdd.n394 vdd.n392 52.4337
R19199 vdd.t292 vdd.t181 51.4683
R19200 vdd.n274 vdd.n272 42.0461
R19201 vdd.n172 vdd.n170 42.0461
R19202 vdd.n71 vdd.n69 42.0461
R19203 vdd.n1752 vdd.n1750 42.0461
R19204 vdd.n1650 vdd.n1648 42.0461
R19205 vdd.n1549 vdd.n1547 42.0461
R19206 vdd.n332 vdd.n331 41.6884
R19207 vdd.n230 vdd.n229 41.6884
R19208 vdd.n129 vdd.n128 41.6884
R19209 vdd.n1810 vdd.n1809 41.6884
R19210 vdd.n1708 vdd.n1707 41.6884
R19211 vdd.n1607 vdd.n1606 41.6884
R19212 vdd.n1319 vdd.n1318 41.1157
R19213 vdd.n1357 vdd.n1356 41.1157
R19214 vdd.n1253 vdd.n1252 41.1157
R19215 vdd.n428 vdd.n427 41.1157
R19216 vdd.n566 vdd.n441 41.1157
R19217 vdd.n454 vdd.n453 41.1157
R19218 vdd.n3053 vdd.n3052 39.2114
R19219 vdd.n3050 vdd.n3049 39.2114
R19220 vdd.n3045 vdd.n815 39.2114
R19221 vdd.n3043 vdd.n3042 39.2114
R19222 vdd.n3038 vdd.n818 39.2114
R19223 vdd.n3036 vdd.n3035 39.2114
R19224 vdd.n3031 vdd.n821 39.2114
R19225 vdd.n3029 vdd.n3028 39.2114
R19226 vdd.n3025 vdd.n3024 39.2114
R19227 vdd.n3020 vdd.n824 39.2114
R19228 vdd.n3018 vdd.n3017 39.2114
R19229 vdd.n3013 vdd.n827 39.2114
R19230 vdd.n3011 vdd.n3010 39.2114
R19231 vdd.n3006 vdd.n830 39.2114
R19232 vdd.n3004 vdd.n3003 39.2114
R19233 vdd.n2998 vdd.n835 39.2114
R19234 vdd.n2996 vdd.n2995 39.2114
R19235 vdd.n2856 vdd.n913 39.2114
R19236 vdd.n2851 vdd.n2605 39.2114
R19237 vdd.n2848 vdd.n2606 39.2114
R19238 vdd.n2844 vdd.n2607 39.2114
R19239 vdd.n2840 vdd.n2608 39.2114
R19240 vdd.n2836 vdd.n2609 39.2114
R19241 vdd.n2832 vdd.n2610 39.2114
R19242 vdd.n2828 vdd.n2611 39.2114
R19243 vdd.n2824 vdd.n2612 39.2114
R19244 vdd.n2820 vdd.n2613 39.2114
R19245 vdd.n2816 vdd.n2614 39.2114
R19246 vdd.n2812 vdd.n2615 39.2114
R19247 vdd.n2808 vdd.n2616 39.2114
R19248 vdd.n2804 vdd.n2617 39.2114
R19249 vdd.n2800 vdd.n2618 39.2114
R19250 vdd.n2796 vdd.n2619 39.2114
R19251 vdd.n2791 vdd.n2620 39.2114
R19252 vdd.n2599 vdd.n953 39.2114
R19253 vdd.n2595 vdd.n952 39.2114
R19254 vdd.n2591 vdd.n951 39.2114
R19255 vdd.n2587 vdd.n950 39.2114
R19256 vdd.n2583 vdd.n949 39.2114
R19257 vdd.n2579 vdd.n948 39.2114
R19258 vdd.n2575 vdd.n947 39.2114
R19259 vdd.n2571 vdd.n946 39.2114
R19260 vdd.n2567 vdd.n945 39.2114
R19261 vdd.n2563 vdd.n944 39.2114
R19262 vdd.n2559 vdd.n943 39.2114
R19263 vdd.n2555 vdd.n942 39.2114
R19264 vdd.n2551 vdd.n941 39.2114
R19265 vdd.n2547 vdd.n940 39.2114
R19266 vdd.n2543 vdd.n939 39.2114
R19267 vdd.n2538 vdd.n938 39.2114
R19268 vdd.n2534 vdd.n937 39.2114
R19269 vdd.n2110 vdd.n1048 39.2114
R19270 vdd.n2116 vdd.n2115 39.2114
R19271 vdd.n2119 vdd.n2118 39.2114
R19272 vdd.n2124 vdd.n2123 39.2114
R19273 vdd.n2127 vdd.n2126 39.2114
R19274 vdd.n2132 vdd.n2131 39.2114
R19275 vdd.n2135 vdd.n2134 39.2114
R19276 vdd.n2140 vdd.n2139 39.2114
R19277 vdd.n2311 vdd.n2142 39.2114
R19278 vdd.n2310 vdd.n2309 39.2114
R19279 vdd.n2303 vdd.n2144 39.2114
R19280 vdd.n2302 vdd.n2301 39.2114
R19281 vdd.n2295 vdd.n2146 39.2114
R19282 vdd.n2294 vdd.n2293 39.2114
R19283 vdd.n2287 vdd.n2148 39.2114
R19284 vdd.n2286 vdd.n2285 39.2114
R19285 vdd.n2279 vdd.n2150 39.2114
R19286 vdd.n2972 vdd.n2971 39.2114
R19287 vdd.n2967 vdd.n2939 39.2114
R19288 vdd.n2965 vdd.n2964 39.2114
R19289 vdd.n2960 vdd.n2942 39.2114
R19290 vdd.n2958 vdd.n2957 39.2114
R19291 vdd.n2953 vdd.n2945 39.2114
R19292 vdd.n2951 vdd.n2950 39.2114
R19293 vdd.n2946 vdd.n787 39.2114
R19294 vdd.n3090 vdd.n3089 39.2114
R19295 vdd.n3087 vdd.n3086 39.2114
R19296 vdd.n3082 vdd.n791 39.2114
R19297 vdd.n3080 vdd.n3079 39.2114
R19298 vdd.n3075 vdd.n794 39.2114
R19299 vdd.n3073 vdd.n3072 39.2114
R19300 vdd.n3068 vdd.n797 39.2114
R19301 vdd.n3066 vdd.n3065 39.2114
R19302 vdd.n3061 vdd.n803 39.2114
R19303 vdd.n2858 vdd.n916 39.2114
R19304 vdd.n2621 vdd.n918 39.2114
R19305 vdd.n2647 vdd.n2622 39.2114
R19306 vdd.n2651 vdd.n2623 39.2114
R19307 vdd.n2655 vdd.n2624 39.2114
R19308 vdd.n2659 vdd.n2625 39.2114
R19309 vdd.n2663 vdd.n2626 39.2114
R19310 vdd.n2667 vdd.n2627 39.2114
R19311 vdd.n2671 vdd.n2628 39.2114
R19312 vdd.n2675 vdd.n2629 39.2114
R19313 vdd.n2679 vdd.n2630 39.2114
R19314 vdd.n2683 vdd.n2631 39.2114
R19315 vdd.n2687 vdd.n2632 39.2114
R19316 vdd.n2691 vdd.n2633 39.2114
R19317 vdd.n2695 vdd.n2634 39.2114
R19318 vdd.n2699 vdd.n2635 39.2114
R19319 vdd.n2703 vdd.n2636 39.2114
R19320 vdd.n2859 vdd.n2858 39.2114
R19321 vdd.n2646 vdd.n2621 39.2114
R19322 vdd.n2650 vdd.n2622 39.2114
R19323 vdd.n2654 vdd.n2623 39.2114
R19324 vdd.n2658 vdd.n2624 39.2114
R19325 vdd.n2662 vdd.n2625 39.2114
R19326 vdd.n2666 vdd.n2626 39.2114
R19327 vdd.n2670 vdd.n2627 39.2114
R19328 vdd.n2674 vdd.n2628 39.2114
R19329 vdd.n2678 vdd.n2629 39.2114
R19330 vdd.n2682 vdd.n2630 39.2114
R19331 vdd.n2686 vdd.n2631 39.2114
R19332 vdd.n2690 vdd.n2632 39.2114
R19333 vdd.n2694 vdd.n2633 39.2114
R19334 vdd.n2698 vdd.n2634 39.2114
R19335 vdd.n2702 vdd.n2635 39.2114
R19336 vdd.n2705 vdd.n2636 39.2114
R19337 vdd.n803 vdd.n798 39.2114
R19338 vdd.n3067 vdd.n3066 39.2114
R19339 vdd.n797 vdd.n795 39.2114
R19340 vdd.n3074 vdd.n3073 39.2114
R19341 vdd.n794 vdd.n792 39.2114
R19342 vdd.n3081 vdd.n3080 39.2114
R19343 vdd.n791 vdd.n789 39.2114
R19344 vdd.n3088 vdd.n3087 39.2114
R19345 vdd.n3091 vdd.n3090 39.2114
R19346 vdd.n2947 vdd.n2946 39.2114
R19347 vdd.n2952 vdd.n2951 39.2114
R19348 vdd.n2945 vdd.n2943 39.2114
R19349 vdd.n2959 vdd.n2958 39.2114
R19350 vdd.n2942 vdd.n2940 39.2114
R19351 vdd.n2966 vdd.n2965 39.2114
R19352 vdd.n2939 vdd.n2937 39.2114
R19353 vdd.n2973 vdd.n2972 39.2114
R19354 vdd.n2111 vdd.n2110 39.2114
R19355 vdd.n2117 vdd.n2116 39.2114
R19356 vdd.n2118 vdd.n2107 39.2114
R19357 vdd.n2125 vdd.n2124 39.2114
R19358 vdd.n2126 vdd.n2105 39.2114
R19359 vdd.n2133 vdd.n2132 39.2114
R19360 vdd.n2134 vdd.n2103 39.2114
R19361 vdd.n2141 vdd.n2140 39.2114
R19362 vdd.n2312 vdd.n2311 39.2114
R19363 vdd.n2309 vdd.n2308 39.2114
R19364 vdd.n2304 vdd.n2303 39.2114
R19365 vdd.n2301 vdd.n2300 39.2114
R19366 vdd.n2296 vdd.n2295 39.2114
R19367 vdd.n2293 vdd.n2292 39.2114
R19368 vdd.n2288 vdd.n2287 39.2114
R19369 vdd.n2285 vdd.n2284 39.2114
R19370 vdd.n2280 vdd.n2279 39.2114
R19371 vdd.n2537 vdd.n937 39.2114
R19372 vdd.n2542 vdd.n938 39.2114
R19373 vdd.n2546 vdd.n939 39.2114
R19374 vdd.n2550 vdd.n940 39.2114
R19375 vdd.n2554 vdd.n941 39.2114
R19376 vdd.n2558 vdd.n942 39.2114
R19377 vdd.n2562 vdd.n943 39.2114
R19378 vdd.n2566 vdd.n944 39.2114
R19379 vdd.n2570 vdd.n945 39.2114
R19380 vdd.n2574 vdd.n946 39.2114
R19381 vdd.n2578 vdd.n947 39.2114
R19382 vdd.n2582 vdd.n948 39.2114
R19383 vdd.n2586 vdd.n949 39.2114
R19384 vdd.n2590 vdd.n950 39.2114
R19385 vdd.n2594 vdd.n951 39.2114
R19386 vdd.n2598 vdd.n952 39.2114
R19387 vdd.n955 vdd.n953 39.2114
R19388 vdd.n2856 vdd.n2855 39.2114
R19389 vdd.n2849 vdd.n2605 39.2114
R19390 vdd.n2845 vdd.n2606 39.2114
R19391 vdd.n2841 vdd.n2607 39.2114
R19392 vdd.n2837 vdd.n2608 39.2114
R19393 vdd.n2833 vdd.n2609 39.2114
R19394 vdd.n2829 vdd.n2610 39.2114
R19395 vdd.n2825 vdd.n2611 39.2114
R19396 vdd.n2821 vdd.n2612 39.2114
R19397 vdd.n2817 vdd.n2613 39.2114
R19398 vdd.n2813 vdd.n2614 39.2114
R19399 vdd.n2809 vdd.n2615 39.2114
R19400 vdd.n2805 vdd.n2616 39.2114
R19401 vdd.n2801 vdd.n2617 39.2114
R19402 vdd.n2797 vdd.n2618 39.2114
R19403 vdd.n2792 vdd.n2619 39.2114
R19404 vdd.n2788 vdd.n2620 39.2114
R19405 vdd.n2997 vdd.n2996 39.2114
R19406 vdd.n835 vdd.n831 39.2114
R19407 vdd.n3005 vdd.n3004 39.2114
R19408 vdd.n830 vdd.n828 39.2114
R19409 vdd.n3012 vdd.n3011 39.2114
R19410 vdd.n827 vdd.n825 39.2114
R19411 vdd.n3019 vdd.n3018 39.2114
R19412 vdd.n824 vdd.n822 39.2114
R19413 vdd.n3026 vdd.n3025 39.2114
R19414 vdd.n3030 vdd.n3029 39.2114
R19415 vdd.n821 vdd.n819 39.2114
R19416 vdd.n3037 vdd.n3036 39.2114
R19417 vdd.n818 vdd.n816 39.2114
R19418 vdd.n3044 vdd.n3043 39.2114
R19419 vdd.n815 vdd.n813 39.2114
R19420 vdd.n3051 vdd.n3050 39.2114
R19421 vdd.n3054 vdd.n3053 39.2114
R19422 vdd.n963 vdd.n919 39.2114
R19423 vdd.n2526 vdd.n920 39.2114
R19424 vdd.n2522 vdd.n921 39.2114
R19425 vdd.n2518 vdd.n922 39.2114
R19426 vdd.n2514 vdd.n923 39.2114
R19427 vdd.n2510 vdd.n924 39.2114
R19428 vdd.n2506 vdd.n925 39.2114
R19429 vdd.n2502 vdd.n926 39.2114
R19430 vdd.n2498 vdd.n927 39.2114
R19431 vdd.n2494 vdd.n928 39.2114
R19432 vdd.n2490 vdd.n929 39.2114
R19433 vdd.n2486 vdd.n930 39.2114
R19434 vdd.n2482 vdd.n931 39.2114
R19435 vdd.n2478 vdd.n932 39.2114
R19436 vdd.n2474 vdd.n933 39.2114
R19437 vdd.n2470 vdd.n934 39.2114
R19438 vdd.n2466 vdd.n935 39.2114
R19439 vdd.n2369 vdd.n1052 39.2114
R19440 vdd.n2368 vdd.n2367 39.2114
R19441 vdd.n2361 vdd.n1054 39.2114
R19442 vdd.n2360 vdd.n2359 39.2114
R19443 vdd.n2353 vdd.n1056 39.2114
R19444 vdd.n2352 vdd.n2351 39.2114
R19445 vdd.n2345 vdd.n1058 39.2114
R19446 vdd.n2344 vdd.n2343 39.2114
R19447 vdd.n1061 vdd.n1060 39.2114
R19448 vdd.n2185 vdd.n2184 39.2114
R19449 vdd.n2190 vdd.n2189 39.2114
R19450 vdd.n2193 vdd.n2192 39.2114
R19451 vdd.n2198 vdd.n2197 39.2114
R19452 vdd.n2201 vdd.n2200 39.2114
R19453 vdd.n2206 vdd.n2205 39.2114
R19454 vdd.n2209 vdd.n2208 39.2114
R19455 vdd.n2215 vdd.n2214 39.2114
R19456 vdd.n2463 vdd.n935 39.2114
R19457 vdd.n2467 vdd.n934 39.2114
R19458 vdd.n2471 vdd.n933 39.2114
R19459 vdd.n2475 vdd.n932 39.2114
R19460 vdd.n2479 vdd.n931 39.2114
R19461 vdd.n2483 vdd.n930 39.2114
R19462 vdd.n2487 vdd.n929 39.2114
R19463 vdd.n2491 vdd.n928 39.2114
R19464 vdd.n2495 vdd.n927 39.2114
R19465 vdd.n2499 vdd.n926 39.2114
R19466 vdd.n2503 vdd.n925 39.2114
R19467 vdd.n2507 vdd.n924 39.2114
R19468 vdd.n2511 vdd.n923 39.2114
R19469 vdd.n2515 vdd.n922 39.2114
R19470 vdd.n2519 vdd.n921 39.2114
R19471 vdd.n2523 vdd.n920 39.2114
R19472 vdd.n2527 vdd.n919 39.2114
R19473 vdd.n2370 vdd.n2369 39.2114
R19474 vdd.n2367 vdd.n2366 39.2114
R19475 vdd.n2362 vdd.n2361 39.2114
R19476 vdd.n2359 vdd.n2358 39.2114
R19477 vdd.n2354 vdd.n2353 39.2114
R19478 vdd.n2351 vdd.n2350 39.2114
R19479 vdd.n2346 vdd.n2345 39.2114
R19480 vdd.n2343 vdd.n2342 39.2114
R19481 vdd.n1062 vdd.n1061 39.2114
R19482 vdd.n2186 vdd.n2185 39.2114
R19483 vdd.n2191 vdd.n2190 39.2114
R19484 vdd.n2192 vdd.n2182 39.2114
R19485 vdd.n2199 vdd.n2198 39.2114
R19486 vdd.n2200 vdd.n2180 39.2114
R19487 vdd.n2207 vdd.n2206 39.2114
R19488 vdd.n2208 vdd.n2176 39.2114
R19489 vdd.n2216 vdd.n2215 39.2114
R19490 vdd.n2335 vdd.n2334 37.2369
R19491 vdd.n2038 vdd.n1971 37.2369
R19492 vdd.n2077 vdd.n1931 37.2369
R19493 vdd.n3138 vdd.n769 37.2369
R19494 vdd.n3186 vdd.n3185 37.2369
R19495 vdd.n690 vdd.n689 37.2369
R19496 vdd.n2377 vdd.n1047 31.6883
R19497 vdd.n2602 vdd.n956 31.6883
R19498 vdd.n2535 vdd.n959 31.6883
R19499 vdd.n2281 vdd.n2278 31.6883
R19500 vdd.n2789 vdd.n2787 31.6883
R19501 vdd.n2994 vdd.n2993 31.6883
R19502 vdd.n2866 vdd.n912 31.6883
R19503 vdd.n3057 vdd.n3056 31.6883
R19504 vdd.n2976 vdd.n2975 31.6883
R19505 vdd.n3062 vdd.n802 31.6883
R19506 vdd.n2708 vdd.n2707 31.6883
R19507 vdd.n2862 vdd.n2861 31.6883
R19508 vdd.n2373 vdd.n2372 31.6883
R19509 vdd.n2530 vdd.n2529 31.6883
R19510 vdd.n2462 vdd.n2461 31.6883
R19511 vdd.n2219 vdd.n2218 31.6883
R19512 vdd.n2212 vdd.n2178 30.449
R19513 vdd.n967 vdd.n966 30.449
R19514 vdd.n2153 vdd.n2152 30.449
R19515 vdd.n2540 vdd.n958 30.449
R19516 vdd.n2644 vdd.n2643 30.449
R19517 vdd.n3000 vdd.n833 30.449
R19518 vdd.n2794 vdd.n2640 30.449
R19519 vdd.n801 vdd.n800 30.449
R19520 vdd.n1418 vdd.n1225 22.2201
R19521 vdd.n2329 vdd.n1073 22.2201
R19522 vdd.n3223 vdd.n723 22.2201
R19523 vdd.n3355 vdd.n3354 22.2201
R19524 vdd.n1429 vdd.n1187 19.3944
R19525 vdd.n1429 vdd.n1185 19.3944
R19526 vdd.n1433 vdd.n1185 19.3944
R19527 vdd.n1433 vdd.n1175 19.3944
R19528 vdd.n1446 vdd.n1175 19.3944
R19529 vdd.n1446 vdd.n1173 19.3944
R19530 vdd.n1450 vdd.n1173 19.3944
R19531 vdd.n1450 vdd.n1165 19.3944
R19532 vdd.n1463 vdd.n1165 19.3944
R19533 vdd.n1463 vdd.n1163 19.3944
R19534 vdd.n1467 vdd.n1163 19.3944
R19535 vdd.n1467 vdd.n1152 19.3944
R19536 vdd.n1479 vdd.n1152 19.3944
R19537 vdd.n1479 vdd.n1150 19.3944
R19538 vdd.n1483 vdd.n1150 19.3944
R19539 vdd.n1483 vdd.n1141 19.3944
R19540 vdd.n1496 vdd.n1141 19.3944
R19541 vdd.n1496 vdd.n1139 19.3944
R19542 vdd.n1500 vdd.n1139 19.3944
R19543 vdd.n1500 vdd.n1130 19.3944
R19544 vdd.n1819 vdd.n1130 19.3944
R19545 vdd.n1819 vdd.n1128 19.3944
R19546 vdd.n1823 vdd.n1128 19.3944
R19547 vdd.n1823 vdd.n1118 19.3944
R19548 vdd.n1836 vdd.n1118 19.3944
R19549 vdd.n1836 vdd.n1116 19.3944
R19550 vdd.n1840 vdd.n1116 19.3944
R19551 vdd.n1840 vdd.n1108 19.3944
R19552 vdd.n1853 vdd.n1108 19.3944
R19553 vdd.n1853 vdd.n1106 19.3944
R19554 vdd.n1857 vdd.n1106 19.3944
R19555 vdd.n1857 vdd.n1095 19.3944
R19556 vdd.n1869 vdd.n1095 19.3944
R19557 vdd.n1869 vdd.n1093 19.3944
R19558 vdd.n1873 vdd.n1093 19.3944
R19559 vdd.n1873 vdd.n1085 19.3944
R19560 vdd.n1886 vdd.n1085 19.3944
R19561 vdd.n1886 vdd.n1082 19.3944
R19562 vdd.n1892 vdd.n1082 19.3944
R19563 vdd.n1892 vdd.n1083 19.3944
R19564 vdd.n1083 vdd.n1072 19.3944
R19565 vdd.n1353 vdd.n1288 19.3944
R19566 vdd.n1349 vdd.n1288 19.3944
R19567 vdd.n1349 vdd.n1348 19.3944
R19568 vdd.n1348 vdd.n1347 19.3944
R19569 vdd.n1347 vdd.n1294 19.3944
R19570 vdd.n1343 vdd.n1294 19.3944
R19571 vdd.n1343 vdd.n1342 19.3944
R19572 vdd.n1342 vdd.n1341 19.3944
R19573 vdd.n1341 vdd.n1300 19.3944
R19574 vdd.n1337 vdd.n1300 19.3944
R19575 vdd.n1337 vdd.n1336 19.3944
R19576 vdd.n1336 vdd.n1335 19.3944
R19577 vdd.n1335 vdd.n1306 19.3944
R19578 vdd.n1331 vdd.n1306 19.3944
R19579 vdd.n1331 vdd.n1330 19.3944
R19580 vdd.n1330 vdd.n1329 19.3944
R19581 vdd.n1329 vdd.n1312 19.3944
R19582 vdd.n1325 vdd.n1312 19.3944
R19583 vdd.n1325 vdd.n1324 19.3944
R19584 vdd.n1324 vdd.n1323 19.3944
R19585 vdd.n1388 vdd.n1387 19.3944
R19586 vdd.n1387 vdd.n1386 19.3944
R19587 vdd.n1386 vdd.n1259 19.3944
R19588 vdd.n1382 vdd.n1259 19.3944
R19589 vdd.n1382 vdd.n1381 19.3944
R19590 vdd.n1381 vdd.n1380 19.3944
R19591 vdd.n1380 vdd.n1265 19.3944
R19592 vdd.n1376 vdd.n1265 19.3944
R19593 vdd.n1376 vdd.n1375 19.3944
R19594 vdd.n1375 vdd.n1374 19.3944
R19595 vdd.n1374 vdd.n1271 19.3944
R19596 vdd.n1370 vdd.n1271 19.3944
R19597 vdd.n1370 vdd.n1369 19.3944
R19598 vdd.n1369 vdd.n1368 19.3944
R19599 vdd.n1368 vdd.n1277 19.3944
R19600 vdd.n1364 vdd.n1277 19.3944
R19601 vdd.n1364 vdd.n1363 19.3944
R19602 vdd.n1363 vdd.n1362 19.3944
R19603 vdd.n1362 vdd.n1283 19.3944
R19604 vdd.n1358 vdd.n1283 19.3944
R19605 vdd.n1421 vdd.n1192 19.3944
R19606 vdd.n1416 vdd.n1192 19.3944
R19607 vdd.n1416 vdd.n1227 19.3944
R19608 vdd.n1412 vdd.n1227 19.3944
R19609 vdd.n1412 vdd.n1411 19.3944
R19610 vdd.n1411 vdd.n1410 19.3944
R19611 vdd.n1410 vdd.n1233 19.3944
R19612 vdd.n1406 vdd.n1233 19.3944
R19613 vdd.n1406 vdd.n1405 19.3944
R19614 vdd.n1405 vdd.n1404 19.3944
R19615 vdd.n1404 vdd.n1239 19.3944
R19616 vdd.n1400 vdd.n1239 19.3944
R19617 vdd.n1400 vdd.n1399 19.3944
R19618 vdd.n1399 vdd.n1398 19.3944
R19619 vdd.n1398 vdd.n1245 19.3944
R19620 vdd.n1394 vdd.n1245 19.3944
R19621 vdd.n1394 vdd.n1393 19.3944
R19622 vdd.n1393 vdd.n1392 19.3944
R19623 vdd.n2034 vdd.n1969 19.3944
R19624 vdd.n2034 vdd.n1975 19.3944
R19625 vdd.n2029 vdd.n1975 19.3944
R19626 vdd.n2029 vdd.n2028 19.3944
R19627 vdd.n2028 vdd.n2027 19.3944
R19628 vdd.n2027 vdd.n1982 19.3944
R19629 vdd.n2022 vdd.n1982 19.3944
R19630 vdd.n2022 vdd.n2021 19.3944
R19631 vdd.n2021 vdd.n2020 19.3944
R19632 vdd.n2020 vdd.n1989 19.3944
R19633 vdd.n2015 vdd.n1989 19.3944
R19634 vdd.n2015 vdd.n2014 19.3944
R19635 vdd.n2014 vdd.n2013 19.3944
R19636 vdd.n2013 vdd.n1997 19.3944
R19637 vdd.n2008 vdd.n1997 19.3944
R19638 vdd.n2008 vdd.n2007 19.3944
R19639 vdd.n2003 vdd.n2002 19.3944
R19640 vdd.n2336 vdd.n1068 19.3944
R19641 vdd.n2073 vdd.n1929 19.3944
R19642 vdd.n2073 vdd.n1935 19.3944
R19643 vdd.n2068 vdd.n1935 19.3944
R19644 vdd.n2068 vdd.n2067 19.3944
R19645 vdd.n2067 vdd.n2066 19.3944
R19646 vdd.n2066 vdd.n1942 19.3944
R19647 vdd.n2061 vdd.n1942 19.3944
R19648 vdd.n2061 vdd.n2060 19.3944
R19649 vdd.n2060 vdd.n2059 19.3944
R19650 vdd.n2059 vdd.n1949 19.3944
R19651 vdd.n2054 vdd.n1949 19.3944
R19652 vdd.n2054 vdd.n2053 19.3944
R19653 vdd.n2053 vdd.n2052 19.3944
R19654 vdd.n2052 vdd.n1956 19.3944
R19655 vdd.n2047 vdd.n1956 19.3944
R19656 vdd.n2047 vdd.n2046 19.3944
R19657 vdd.n2046 vdd.n2045 19.3944
R19658 vdd.n2045 vdd.n1963 19.3944
R19659 vdd.n2040 vdd.n1963 19.3944
R19660 vdd.n2040 vdd.n2039 19.3944
R19661 vdd.n2324 vdd.n2323 19.3944
R19662 vdd.n2323 vdd.n1901 19.3944
R19663 vdd.n2318 vdd.n2317 19.3944
R19664 vdd.n2100 vdd.n1905 19.3944
R19665 vdd.n2100 vdd.n1907 19.3944
R19666 vdd.n1910 vdd.n1907 19.3944
R19667 vdd.n2093 vdd.n1910 19.3944
R19668 vdd.n2093 vdd.n2092 19.3944
R19669 vdd.n2092 vdd.n2091 19.3944
R19670 vdd.n2091 vdd.n1916 19.3944
R19671 vdd.n2086 vdd.n1916 19.3944
R19672 vdd.n2086 vdd.n2085 19.3944
R19673 vdd.n2085 vdd.n2084 19.3944
R19674 vdd.n2084 vdd.n1923 19.3944
R19675 vdd.n2079 vdd.n1923 19.3944
R19676 vdd.n2079 vdd.n2078 19.3944
R19677 vdd.n1425 vdd.n1190 19.3944
R19678 vdd.n1425 vdd.n1181 19.3944
R19679 vdd.n1438 vdd.n1181 19.3944
R19680 vdd.n1438 vdd.n1179 19.3944
R19681 vdd.n1442 vdd.n1179 19.3944
R19682 vdd.n1442 vdd.n1170 19.3944
R19683 vdd.n1455 vdd.n1170 19.3944
R19684 vdd.n1455 vdd.n1168 19.3944
R19685 vdd.n1459 vdd.n1168 19.3944
R19686 vdd.n1459 vdd.n1159 19.3944
R19687 vdd.n1471 vdd.n1159 19.3944
R19688 vdd.n1471 vdd.n1157 19.3944
R19689 vdd.n1475 vdd.n1157 19.3944
R19690 vdd.n1475 vdd.n1147 19.3944
R19691 vdd.n1488 vdd.n1147 19.3944
R19692 vdd.n1488 vdd.n1145 19.3944
R19693 vdd.n1492 vdd.n1145 19.3944
R19694 vdd.n1492 vdd.n1136 19.3944
R19695 vdd.n1504 vdd.n1136 19.3944
R19696 vdd.n1504 vdd.n1134 19.3944
R19697 vdd.n1815 vdd.n1134 19.3944
R19698 vdd.n1815 vdd.n1124 19.3944
R19699 vdd.n1828 vdd.n1124 19.3944
R19700 vdd.n1828 vdd.n1122 19.3944
R19701 vdd.n1832 vdd.n1122 19.3944
R19702 vdd.n1832 vdd.n1113 19.3944
R19703 vdd.n1845 vdd.n1113 19.3944
R19704 vdd.n1845 vdd.n1111 19.3944
R19705 vdd.n1849 vdd.n1111 19.3944
R19706 vdd.n1849 vdd.n1102 19.3944
R19707 vdd.n1861 vdd.n1102 19.3944
R19708 vdd.n1861 vdd.n1100 19.3944
R19709 vdd.n1865 vdd.n1100 19.3944
R19710 vdd.n1865 vdd.n1090 19.3944
R19711 vdd.n1878 vdd.n1090 19.3944
R19712 vdd.n1878 vdd.n1088 19.3944
R19713 vdd.n1882 vdd.n1088 19.3944
R19714 vdd.n1882 vdd.n1078 19.3944
R19715 vdd.n1897 vdd.n1078 19.3944
R19716 vdd.n1897 vdd.n1076 19.3944
R19717 vdd.n2327 vdd.n1076 19.3944
R19718 vdd.n3229 vdd.n686 19.3944
R19719 vdd.n3229 vdd.n676 19.3944
R19720 vdd.n3241 vdd.n676 19.3944
R19721 vdd.n3241 vdd.n674 19.3944
R19722 vdd.n3245 vdd.n674 19.3944
R19723 vdd.n3245 vdd.n666 19.3944
R19724 vdd.n3258 vdd.n666 19.3944
R19725 vdd.n3258 vdd.n664 19.3944
R19726 vdd.n3262 vdd.n664 19.3944
R19727 vdd.n3262 vdd.n653 19.3944
R19728 vdd.n3274 vdd.n653 19.3944
R19729 vdd.n3274 vdd.n651 19.3944
R19730 vdd.n3278 vdd.n651 19.3944
R19731 vdd.n3278 vdd.n642 19.3944
R19732 vdd.n3291 vdd.n642 19.3944
R19733 vdd.n3291 vdd.n640 19.3944
R19734 vdd.n3298 vdd.n640 19.3944
R19735 vdd.n3298 vdd.n3297 19.3944
R19736 vdd.n3297 vdd.n631 19.3944
R19737 vdd.n3311 vdd.n631 19.3944
R19738 vdd.n3312 vdd.n3311 19.3944
R19739 vdd.n3312 vdd.n629 19.3944
R19740 vdd.n3316 vdd.n629 19.3944
R19741 vdd.n3318 vdd.n3316 19.3944
R19742 vdd.n3319 vdd.n3318 19.3944
R19743 vdd.n3319 vdd.n627 19.3944
R19744 vdd.n3323 vdd.n627 19.3944
R19745 vdd.n3325 vdd.n3323 19.3944
R19746 vdd.n3326 vdd.n3325 19.3944
R19747 vdd.n3326 vdd.n625 19.3944
R19748 vdd.n3330 vdd.n625 19.3944
R19749 vdd.n3333 vdd.n3330 19.3944
R19750 vdd.n3334 vdd.n3333 19.3944
R19751 vdd.n3334 vdd.n623 19.3944
R19752 vdd.n3338 vdd.n623 19.3944
R19753 vdd.n3340 vdd.n3338 19.3944
R19754 vdd.n3341 vdd.n3340 19.3944
R19755 vdd.n3341 vdd.n621 19.3944
R19756 vdd.n3345 vdd.n621 19.3944
R19757 vdd.n3347 vdd.n3345 19.3944
R19758 vdd.n3348 vdd.n3347 19.3944
R19759 vdd.n569 vdd.n438 19.3944
R19760 vdd.n575 vdd.n438 19.3944
R19761 vdd.n576 vdd.n575 19.3944
R19762 vdd.n579 vdd.n576 19.3944
R19763 vdd.n579 vdd.n436 19.3944
R19764 vdd.n585 vdd.n436 19.3944
R19765 vdd.n586 vdd.n585 19.3944
R19766 vdd.n589 vdd.n586 19.3944
R19767 vdd.n589 vdd.n434 19.3944
R19768 vdd.n595 vdd.n434 19.3944
R19769 vdd.n596 vdd.n595 19.3944
R19770 vdd.n599 vdd.n596 19.3944
R19771 vdd.n599 vdd.n432 19.3944
R19772 vdd.n605 vdd.n432 19.3944
R19773 vdd.n606 vdd.n605 19.3944
R19774 vdd.n609 vdd.n606 19.3944
R19775 vdd.n609 vdd.n430 19.3944
R19776 vdd.n615 vdd.n430 19.3944
R19777 vdd.n617 vdd.n615 19.3944
R19778 vdd.n618 vdd.n617 19.3944
R19779 vdd.n516 vdd.n515 19.3944
R19780 vdd.n519 vdd.n516 19.3944
R19781 vdd.n519 vdd.n450 19.3944
R19782 vdd.n525 vdd.n450 19.3944
R19783 vdd.n526 vdd.n525 19.3944
R19784 vdd.n529 vdd.n526 19.3944
R19785 vdd.n529 vdd.n448 19.3944
R19786 vdd.n535 vdd.n448 19.3944
R19787 vdd.n536 vdd.n535 19.3944
R19788 vdd.n539 vdd.n536 19.3944
R19789 vdd.n539 vdd.n446 19.3944
R19790 vdd.n545 vdd.n446 19.3944
R19791 vdd.n546 vdd.n545 19.3944
R19792 vdd.n549 vdd.n546 19.3944
R19793 vdd.n549 vdd.n444 19.3944
R19794 vdd.n555 vdd.n444 19.3944
R19795 vdd.n556 vdd.n555 19.3944
R19796 vdd.n559 vdd.n556 19.3944
R19797 vdd.n559 vdd.n442 19.3944
R19798 vdd.n565 vdd.n442 19.3944
R19799 vdd.n466 vdd.n465 19.3944
R19800 vdd.n469 vdd.n466 19.3944
R19801 vdd.n469 vdd.n462 19.3944
R19802 vdd.n475 vdd.n462 19.3944
R19803 vdd.n476 vdd.n475 19.3944
R19804 vdd.n479 vdd.n476 19.3944
R19805 vdd.n479 vdd.n460 19.3944
R19806 vdd.n485 vdd.n460 19.3944
R19807 vdd.n486 vdd.n485 19.3944
R19808 vdd.n489 vdd.n486 19.3944
R19809 vdd.n489 vdd.n458 19.3944
R19810 vdd.n495 vdd.n458 19.3944
R19811 vdd.n496 vdd.n495 19.3944
R19812 vdd.n499 vdd.n496 19.3944
R19813 vdd.n499 vdd.n456 19.3944
R19814 vdd.n505 vdd.n456 19.3944
R19815 vdd.n506 vdd.n505 19.3944
R19816 vdd.n509 vdd.n506 19.3944
R19817 vdd.n3233 vdd.n683 19.3944
R19818 vdd.n3233 vdd.n681 19.3944
R19819 vdd.n3237 vdd.n681 19.3944
R19820 vdd.n3237 vdd.n671 19.3944
R19821 vdd.n3250 vdd.n671 19.3944
R19822 vdd.n3250 vdd.n669 19.3944
R19823 vdd.n3254 vdd.n669 19.3944
R19824 vdd.n3254 vdd.n660 19.3944
R19825 vdd.n3266 vdd.n660 19.3944
R19826 vdd.n3266 vdd.n658 19.3944
R19827 vdd.n3270 vdd.n658 19.3944
R19828 vdd.n3270 vdd.n648 19.3944
R19829 vdd.n3283 vdd.n648 19.3944
R19830 vdd.n3283 vdd.n646 19.3944
R19831 vdd.n3287 vdd.n646 19.3944
R19832 vdd.n3287 vdd.n637 19.3944
R19833 vdd.n3302 vdd.n637 19.3944
R19834 vdd.n3302 vdd.n635 19.3944
R19835 vdd.n3306 vdd.n635 19.3944
R19836 vdd.n3306 vdd.n336 19.3944
R19837 vdd.n3397 vdd.n336 19.3944
R19838 vdd.n3397 vdd.n337 19.3944
R19839 vdd.n3391 vdd.n337 19.3944
R19840 vdd.n3391 vdd.n3390 19.3944
R19841 vdd.n3390 vdd.n3389 19.3944
R19842 vdd.n3389 vdd.n349 19.3944
R19843 vdd.n3383 vdd.n349 19.3944
R19844 vdd.n3383 vdd.n3382 19.3944
R19845 vdd.n3382 vdd.n3381 19.3944
R19846 vdd.n3381 vdd.n359 19.3944
R19847 vdd.n3375 vdd.n359 19.3944
R19848 vdd.n3375 vdd.n3374 19.3944
R19849 vdd.n3374 vdd.n3373 19.3944
R19850 vdd.n3373 vdd.n370 19.3944
R19851 vdd.n3367 vdd.n370 19.3944
R19852 vdd.n3367 vdd.n3366 19.3944
R19853 vdd.n3366 vdd.n3365 19.3944
R19854 vdd.n3365 vdd.n381 19.3944
R19855 vdd.n3359 vdd.n381 19.3944
R19856 vdd.n3359 vdd.n3358 19.3944
R19857 vdd.n3358 vdd.n3357 19.3944
R19858 vdd.n3180 vdd.n747 19.3944
R19859 vdd.n3180 vdd.n3177 19.3944
R19860 vdd.n3177 vdd.n3174 19.3944
R19861 vdd.n3174 vdd.n3173 19.3944
R19862 vdd.n3173 vdd.n3170 19.3944
R19863 vdd.n3170 vdd.n3169 19.3944
R19864 vdd.n3169 vdd.n3166 19.3944
R19865 vdd.n3166 vdd.n3165 19.3944
R19866 vdd.n3165 vdd.n3162 19.3944
R19867 vdd.n3162 vdd.n3161 19.3944
R19868 vdd.n3161 vdd.n3158 19.3944
R19869 vdd.n3158 vdd.n3157 19.3944
R19870 vdd.n3157 vdd.n3154 19.3944
R19871 vdd.n3154 vdd.n3153 19.3944
R19872 vdd.n3153 vdd.n3150 19.3944
R19873 vdd.n3150 vdd.n3149 19.3944
R19874 vdd.n3149 vdd.n3146 19.3944
R19875 vdd.n3146 vdd.n3145 19.3944
R19876 vdd.n3145 vdd.n3142 19.3944
R19877 vdd.n3142 vdd.n3141 19.3944
R19878 vdd.n3220 vdd.n3219 19.3944
R19879 vdd.n3219 vdd.n3218 19.3944
R19880 vdd.n732 vdd.n729 19.3944
R19881 vdd.n3214 vdd.n3213 19.3944
R19882 vdd.n3213 vdd.n3210 19.3944
R19883 vdd.n3210 vdd.n3209 19.3944
R19884 vdd.n3209 vdd.n3206 19.3944
R19885 vdd.n3206 vdd.n3205 19.3944
R19886 vdd.n3205 vdd.n3202 19.3944
R19887 vdd.n3202 vdd.n3201 19.3944
R19888 vdd.n3201 vdd.n3198 19.3944
R19889 vdd.n3198 vdd.n3197 19.3944
R19890 vdd.n3197 vdd.n3194 19.3944
R19891 vdd.n3194 vdd.n3193 19.3944
R19892 vdd.n3193 vdd.n3190 19.3944
R19893 vdd.n3190 vdd.n3189 19.3944
R19894 vdd.n3134 vdd.n767 19.3944
R19895 vdd.n3134 vdd.n3131 19.3944
R19896 vdd.n3131 vdd.n3128 19.3944
R19897 vdd.n3128 vdd.n3127 19.3944
R19898 vdd.n3127 vdd.n3124 19.3944
R19899 vdd.n3124 vdd.n3123 19.3944
R19900 vdd.n3123 vdd.n3120 19.3944
R19901 vdd.n3120 vdd.n3119 19.3944
R19902 vdd.n3119 vdd.n3116 19.3944
R19903 vdd.n3116 vdd.n3115 19.3944
R19904 vdd.n3115 vdd.n3112 19.3944
R19905 vdd.n3112 vdd.n3111 19.3944
R19906 vdd.n3111 vdd.n3108 19.3944
R19907 vdd.n3108 vdd.n3107 19.3944
R19908 vdd.n3107 vdd.n3104 19.3944
R19909 vdd.n3104 vdd.n3103 19.3944
R19910 vdd.n3100 vdd.n3099 19.3944
R19911 vdd.n3096 vdd.n3095 19.3944
R19912 vdd.n1357 vdd.n1353 19.0066
R19913 vdd.n2038 vdd.n1969 19.0066
R19914 vdd.n569 vdd.n566 19.0066
R19915 vdd.n3138 vdd.n767 19.0066
R19916 vdd.n2178 vdd.n2177 16.0975
R19917 vdd.n966 vdd.n965 16.0975
R19918 vdd.n1318 vdd.n1317 16.0975
R19919 vdd.n1356 vdd.n1355 16.0975
R19920 vdd.n1252 vdd.n1251 16.0975
R19921 vdd.n2334 vdd.n2333 16.0975
R19922 vdd.n1971 vdd.n1970 16.0975
R19923 vdd.n1931 vdd.n1930 16.0975
R19924 vdd.n2152 vdd.n2151 16.0975
R19925 vdd.n958 vdd.n957 16.0975
R19926 vdd.n2643 vdd.n2642 16.0975
R19927 vdd.n427 vdd.n426 16.0975
R19928 vdd.n441 vdd.n440 16.0975
R19929 vdd.n453 vdd.n452 16.0975
R19930 vdd.n769 vdd.n768 16.0975
R19931 vdd.n3185 vdd.n3184 16.0975
R19932 vdd.n833 vdd.n832 16.0975
R19933 vdd.n2640 vdd.n2639 16.0975
R19934 vdd.n689 vdd.n688 16.0975
R19935 vdd.n800 vdd.n799 16.0975
R19936 vdd.t181 vdd.n2604 15.4182
R19937 vdd.n2857 vdd.t292 15.4182
R19938 vdd.n28 vdd.n27 14.6905
R19939 vdd.n2375 vdd.n1049 14.5112
R19940 vdd.n3059 vdd.n692 14.5112
R19941 vdd.n328 vdd.n293 13.1884
R19942 vdd.n269 vdd.n234 13.1884
R19943 vdd.n226 vdd.n191 13.1884
R19944 vdd.n167 vdd.n132 13.1884
R19945 vdd.n125 vdd.n90 13.1884
R19946 vdd.n66 vdd.n31 13.1884
R19947 vdd.n1747 vdd.n1712 13.1884
R19948 vdd.n1806 vdd.n1771 13.1884
R19949 vdd.n1645 vdd.n1610 13.1884
R19950 vdd.n1704 vdd.n1669 13.1884
R19951 vdd.n1544 vdd.n1509 13.1884
R19952 vdd.n1603 vdd.n1568 13.1884
R19953 vdd.n1388 vdd.n1253 12.9944
R19954 vdd.n1392 vdd.n1253 12.9944
R19955 vdd.n2077 vdd.n1929 12.9944
R19956 vdd.n2078 vdd.n2077 12.9944
R19957 vdd.n515 vdd.n454 12.9944
R19958 vdd.n509 vdd.n454 12.9944
R19959 vdd.n3186 vdd.n747 12.9944
R19960 vdd.n3189 vdd.n3186 12.9944
R19961 vdd.n329 vdd.n291 12.8005
R19962 vdd.n324 vdd.n295 12.8005
R19963 vdd.n270 vdd.n232 12.8005
R19964 vdd.n265 vdd.n236 12.8005
R19965 vdd.n227 vdd.n189 12.8005
R19966 vdd.n222 vdd.n193 12.8005
R19967 vdd.n168 vdd.n130 12.8005
R19968 vdd.n163 vdd.n134 12.8005
R19969 vdd.n126 vdd.n88 12.8005
R19970 vdd.n121 vdd.n92 12.8005
R19971 vdd.n67 vdd.n29 12.8005
R19972 vdd.n62 vdd.n33 12.8005
R19973 vdd.n1748 vdd.n1710 12.8005
R19974 vdd.n1743 vdd.n1714 12.8005
R19975 vdd.n1807 vdd.n1769 12.8005
R19976 vdd.n1802 vdd.n1773 12.8005
R19977 vdd.n1646 vdd.n1608 12.8005
R19978 vdd.n1641 vdd.n1612 12.8005
R19979 vdd.n1705 vdd.n1667 12.8005
R19980 vdd.n1700 vdd.n1671 12.8005
R19981 vdd.n1545 vdd.n1507 12.8005
R19982 vdd.n1540 vdd.n1511 12.8005
R19983 vdd.n1604 vdd.n1566 12.8005
R19984 vdd.n1599 vdd.n1570 12.8005
R19985 vdd.n323 vdd.n296 12.0247
R19986 vdd.n264 vdd.n237 12.0247
R19987 vdd.n221 vdd.n194 12.0247
R19988 vdd.n162 vdd.n135 12.0247
R19989 vdd.n120 vdd.n93 12.0247
R19990 vdd.n61 vdd.n34 12.0247
R19991 vdd.n1742 vdd.n1715 12.0247
R19992 vdd.n1801 vdd.n1774 12.0247
R19993 vdd.n1640 vdd.n1613 12.0247
R19994 vdd.n1699 vdd.n1672 12.0247
R19995 vdd.n1539 vdd.n1512 12.0247
R19996 vdd.n1598 vdd.n1571 12.0247
R19997 vdd.n1427 vdd.n1183 11.337
R19998 vdd.n1436 vdd.n1183 11.337
R19999 vdd.n1436 vdd.n1435 11.337
R20000 vdd.n1444 vdd.n1177 11.337
R20001 vdd.n1453 vdd.n1452 11.337
R20002 vdd.n1469 vdd.n1161 11.337
R20003 vdd.n1477 vdd.n1154 11.337
R20004 vdd.n1486 vdd.n1485 11.337
R20005 vdd.n1494 vdd.n1143 11.337
R20006 vdd.n1817 vdd.n1132 11.337
R20007 vdd.n1826 vdd.n1126 11.337
R20008 vdd.n1834 vdd.n1120 11.337
R20009 vdd.n1843 vdd.n1842 11.337
R20010 vdd.n1859 vdd.n1104 11.337
R20011 vdd.n1867 vdd.n1097 11.337
R20012 vdd.n1876 vdd.n1875 11.337
R20013 vdd.n1884 vdd.n1080 11.337
R20014 vdd.n1895 vdd.n1080 11.337
R20015 vdd.n1895 vdd.n1894 11.337
R20016 vdd.n3231 vdd.n678 11.337
R20017 vdd.n3239 vdd.n678 11.337
R20018 vdd.n3239 vdd.n679 11.337
R20019 vdd.n3248 vdd.n3247 11.337
R20020 vdd.n3264 vdd.n662 11.337
R20021 vdd.n3272 vdd.n655 11.337
R20022 vdd.n3281 vdd.n3280 11.337
R20023 vdd.n3289 vdd.n644 11.337
R20024 vdd.n3308 vdd.n633 11.337
R20025 vdd.n3395 vdd.n340 11.337
R20026 vdd.n3393 vdd.n344 11.337
R20027 vdd.n3387 vdd.n3386 11.337
R20028 vdd.n3379 vdd.n361 11.337
R20029 vdd.n3378 vdd.n3377 11.337
R20030 vdd.n3371 vdd.n3370 11.337
R20031 vdd.n3369 vdd.n375 11.337
R20032 vdd.n3363 vdd.n3362 11.337
R20033 vdd.n3362 vdd.n3361 11.337
R20034 vdd.n3361 vdd.n386 11.337
R20035 vdd.n320 vdd.n319 11.249
R20036 vdd.n261 vdd.n260 11.249
R20037 vdd.n218 vdd.n217 11.249
R20038 vdd.n159 vdd.n158 11.249
R20039 vdd.n117 vdd.n116 11.249
R20040 vdd.n58 vdd.n57 11.249
R20041 vdd.n1739 vdd.n1738 11.249
R20042 vdd.n1798 vdd.n1797 11.249
R20043 vdd.n1637 vdd.n1636 11.249
R20044 vdd.n1696 vdd.n1695 11.249
R20045 vdd.n1536 vdd.n1535 11.249
R20046 vdd.n1595 vdd.n1594 11.249
R20047 vdd.n1225 vdd.t226 11.2237
R20048 vdd.n3355 vdd.t233 11.2237
R20049 vdd.n2532 vdd.t294 11.1103
R20050 vdd.n2864 vdd.t286 11.1103
R20051 vdd.t31 vdd.n1098 10.7702
R20052 vdd.n3256 vdd.t94 10.7702
R20053 vdd.n305 vdd.n304 10.7238
R20054 vdd.n246 vdd.n245 10.7238
R20055 vdd.n203 vdd.n202 10.7238
R20056 vdd.n144 vdd.n143 10.7238
R20057 vdd.n102 vdd.n101 10.7238
R20058 vdd.n43 vdd.n42 10.7238
R20059 vdd.n1724 vdd.n1723 10.7238
R20060 vdd.n1783 vdd.n1782 10.7238
R20061 vdd.n1622 vdd.n1621 10.7238
R20062 vdd.n1681 vdd.n1680 10.7238
R20063 vdd.n1521 vdd.n1520 10.7238
R20064 vdd.n1580 vdd.n1579 10.7238
R20065 vdd.n2378 vdd.n2377 10.6151
R20066 vdd.n2379 vdd.n2378 10.6151
R20067 vdd.n2379 vdd.n1035 10.6151
R20068 vdd.n2389 vdd.n1035 10.6151
R20069 vdd.n2390 vdd.n2389 10.6151
R20070 vdd.n2391 vdd.n2390 10.6151
R20071 vdd.n2391 vdd.n1022 10.6151
R20072 vdd.n2402 vdd.n1022 10.6151
R20073 vdd.n2403 vdd.n2402 10.6151
R20074 vdd.n2404 vdd.n2403 10.6151
R20075 vdd.n2404 vdd.n1010 10.6151
R20076 vdd.n2414 vdd.n1010 10.6151
R20077 vdd.n2415 vdd.n2414 10.6151
R20078 vdd.n2416 vdd.n2415 10.6151
R20079 vdd.n2416 vdd.n998 10.6151
R20080 vdd.n2426 vdd.n998 10.6151
R20081 vdd.n2427 vdd.n2426 10.6151
R20082 vdd.n2428 vdd.n2427 10.6151
R20083 vdd.n2428 vdd.n987 10.6151
R20084 vdd.n2438 vdd.n987 10.6151
R20085 vdd.n2439 vdd.n2438 10.6151
R20086 vdd.n2440 vdd.n2439 10.6151
R20087 vdd.n2440 vdd.n974 10.6151
R20088 vdd.n2452 vdd.n974 10.6151
R20089 vdd.n2453 vdd.n2452 10.6151
R20090 vdd.n2455 vdd.n2453 10.6151
R20091 vdd.n2455 vdd.n2454 10.6151
R20092 vdd.n2454 vdd.n956 10.6151
R20093 vdd.n2602 vdd.n2601 10.6151
R20094 vdd.n2601 vdd.n2600 10.6151
R20095 vdd.n2600 vdd.n2597 10.6151
R20096 vdd.n2597 vdd.n2596 10.6151
R20097 vdd.n2596 vdd.n2593 10.6151
R20098 vdd.n2593 vdd.n2592 10.6151
R20099 vdd.n2592 vdd.n2589 10.6151
R20100 vdd.n2589 vdd.n2588 10.6151
R20101 vdd.n2588 vdd.n2585 10.6151
R20102 vdd.n2585 vdd.n2584 10.6151
R20103 vdd.n2584 vdd.n2581 10.6151
R20104 vdd.n2581 vdd.n2580 10.6151
R20105 vdd.n2580 vdd.n2577 10.6151
R20106 vdd.n2577 vdd.n2576 10.6151
R20107 vdd.n2576 vdd.n2573 10.6151
R20108 vdd.n2573 vdd.n2572 10.6151
R20109 vdd.n2572 vdd.n2569 10.6151
R20110 vdd.n2569 vdd.n2568 10.6151
R20111 vdd.n2568 vdd.n2565 10.6151
R20112 vdd.n2565 vdd.n2564 10.6151
R20113 vdd.n2564 vdd.n2561 10.6151
R20114 vdd.n2561 vdd.n2560 10.6151
R20115 vdd.n2560 vdd.n2557 10.6151
R20116 vdd.n2557 vdd.n2556 10.6151
R20117 vdd.n2556 vdd.n2553 10.6151
R20118 vdd.n2553 vdd.n2552 10.6151
R20119 vdd.n2552 vdd.n2549 10.6151
R20120 vdd.n2549 vdd.n2548 10.6151
R20121 vdd.n2548 vdd.n2545 10.6151
R20122 vdd.n2545 vdd.n2544 10.6151
R20123 vdd.n2544 vdd.n2541 10.6151
R20124 vdd.n2539 vdd.n2536 10.6151
R20125 vdd.n2536 vdd.n2535 10.6151
R20126 vdd.n2278 vdd.n2277 10.6151
R20127 vdd.n2277 vdd.n2275 10.6151
R20128 vdd.n2275 vdd.n2274 10.6151
R20129 vdd.n2274 vdd.n2272 10.6151
R20130 vdd.n2272 vdd.n2271 10.6151
R20131 vdd.n2271 vdd.n2269 10.6151
R20132 vdd.n2269 vdd.n2268 10.6151
R20133 vdd.n2268 vdd.n2266 10.6151
R20134 vdd.n2266 vdd.n2265 10.6151
R20135 vdd.n2265 vdd.n2263 10.6151
R20136 vdd.n2263 vdd.n2262 10.6151
R20137 vdd.n2262 vdd.n2260 10.6151
R20138 vdd.n2260 vdd.n2259 10.6151
R20139 vdd.n2259 vdd.n2174 10.6151
R20140 vdd.n2174 vdd.n2173 10.6151
R20141 vdd.n2173 vdd.n2171 10.6151
R20142 vdd.n2171 vdd.n2170 10.6151
R20143 vdd.n2170 vdd.n2168 10.6151
R20144 vdd.n2168 vdd.n2167 10.6151
R20145 vdd.n2167 vdd.n2165 10.6151
R20146 vdd.n2165 vdd.n2164 10.6151
R20147 vdd.n2164 vdd.n2162 10.6151
R20148 vdd.n2162 vdd.n2161 10.6151
R20149 vdd.n2161 vdd.n2159 10.6151
R20150 vdd.n2159 vdd.n2158 10.6151
R20151 vdd.n2158 vdd.n2155 10.6151
R20152 vdd.n2155 vdd.n2154 10.6151
R20153 vdd.n2154 vdd.n959 10.6151
R20154 vdd.n2112 vdd.n1047 10.6151
R20155 vdd.n2113 vdd.n2112 10.6151
R20156 vdd.n2114 vdd.n2113 10.6151
R20157 vdd.n2114 vdd.n2108 10.6151
R20158 vdd.n2120 vdd.n2108 10.6151
R20159 vdd.n2121 vdd.n2120 10.6151
R20160 vdd.n2122 vdd.n2121 10.6151
R20161 vdd.n2122 vdd.n2106 10.6151
R20162 vdd.n2128 vdd.n2106 10.6151
R20163 vdd.n2129 vdd.n2128 10.6151
R20164 vdd.n2130 vdd.n2129 10.6151
R20165 vdd.n2130 vdd.n2104 10.6151
R20166 vdd.n2136 vdd.n2104 10.6151
R20167 vdd.n2137 vdd.n2136 10.6151
R20168 vdd.n2138 vdd.n2137 10.6151
R20169 vdd.n2138 vdd.n2102 10.6151
R20170 vdd.n2314 vdd.n2102 10.6151
R20171 vdd.n2314 vdd.n2313 10.6151
R20172 vdd.n2313 vdd.n2143 10.6151
R20173 vdd.n2307 vdd.n2143 10.6151
R20174 vdd.n2307 vdd.n2306 10.6151
R20175 vdd.n2306 vdd.n2305 10.6151
R20176 vdd.n2305 vdd.n2145 10.6151
R20177 vdd.n2299 vdd.n2145 10.6151
R20178 vdd.n2299 vdd.n2298 10.6151
R20179 vdd.n2298 vdd.n2297 10.6151
R20180 vdd.n2297 vdd.n2147 10.6151
R20181 vdd.n2291 vdd.n2147 10.6151
R20182 vdd.n2291 vdd.n2290 10.6151
R20183 vdd.n2290 vdd.n2289 10.6151
R20184 vdd.n2289 vdd.n2149 10.6151
R20185 vdd.n2283 vdd.n2282 10.6151
R20186 vdd.n2282 vdd.n2281 10.6151
R20187 vdd.n2787 vdd.n2786 10.6151
R20188 vdd.n2786 vdd.n2784 10.6151
R20189 vdd.n2784 vdd.n2783 10.6151
R20190 vdd.n2783 vdd.n2641 10.6151
R20191 vdd.n2730 vdd.n2641 10.6151
R20192 vdd.n2731 vdd.n2730 10.6151
R20193 vdd.n2733 vdd.n2731 10.6151
R20194 vdd.n2734 vdd.n2733 10.6151
R20195 vdd.n2736 vdd.n2734 10.6151
R20196 vdd.n2737 vdd.n2736 10.6151
R20197 vdd.n2739 vdd.n2737 10.6151
R20198 vdd.n2740 vdd.n2739 10.6151
R20199 vdd.n2742 vdd.n2740 10.6151
R20200 vdd.n2743 vdd.n2742 10.6151
R20201 vdd.n2758 vdd.n2743 10.6151
R20202 vdd.n2758 vdd.n2757 10.6151
R20203 vdd.n2757 vdd.n2756 10.6151
R20204 vdd.n2756 vdd.n2754 10.6151
R20205 vdd.n2754 vdd.n2753 10.6151
R20206 vdd.n2753 vdd.n2751 10.6151
R20207 vdd.n2751 vdd.n2750 10.6151
R20208 vdd.n2750 vdd.n2748 10.6151
R20209 vdd.n2748 vdd.n2747 10.6151
R20210 vdd.n2747 vdd.n2745 10.6151
R20211 vdd.n2745 vdd.n2744 10.6151
R20212 vdd.n2744 vdd.n836 10.6151
R20213 vdd.n2992 vdd.n836 10.6151
R20214 vdd.n2993 vdd.n2992 10.6151
R20215 vdd.n2854 vdd.n912 10.6151
R20216 vdd.n2854 vdd.n2853 10.6151
R20217 vdd.n2853 vdd.n2852 10.6151
R20218 vdd.n2852 vdd.n2850 10.6151
R20219 vdd.n2850 vdd.n2847 10.6151
R20220 vdd.n2847 vdd.n2846 10.6151
R20221 vdd.n2846 vdd.n2843 10.6151
R20222 vdd.n2843 vdd.n2842 10.6151
R20223 vdd.n2842 vdd.n2839 10.6151
R20224 vdd.n2839 vdd.n2838 10.6151
R20225 vdd.n2838 vdd.n2835 10.6151
R20226 vdd.n2835 vdd.n2834 10.6151
R20227 vdd.n2834 vdd.n2831 10.6151
R20228 vdd.n2831 vdd.n2830 10.6151
R20229 vdd.n2830 vdd.n2827 10.6151
R20230 vdd.n2827 vdd.n2826 10.6151
R20231 vdd.n2826 vdd.n2823 10.6151
R20232 vdd.n2823 vdd.n2822 10.6151
R20233 vdd.n2822 vdd.n2819 10.6151
R20234 vdd.n2819 vdd.n2818 10.6151
R20235 vdd.n2818 vdd.n2815 10.6151
R20236 vdd.n2815 vdd.n2814 10.6151
R20237 vdd.n2814 vdd.n2811 10.6151
R20238 vdd.n2811 vdd.n2810 10.6151
R20239 vdd.n2810 vdd.n2807 10.6151
R20240 vdd.n2807 vdd.n2806 10.6151
R20241 vdd.n2806 vdd.n2803 10.6151
R20242 vdd.n2803 vdd.n2802 10.6151
R20243 vdd.n2802 vdd.n2799 10.6151
R20244 vdd.n2799 vdd.n2798 10.6151
R20245 vdd.n2798 vdd.n2795 10.6151
R20246 vdd.n2793 vdd.n2790 10.6151
R20247 vdd.n2790 vdd.n2789 10.6151
R20248 vdd.n2867 vdd.n2866 10.6151
R20249 vdd.n2868 vdd.n2867 10.6151
R20250 vdd.n2868 vdd.n902 10.6151
R20251 vdd.n2878 vdd.n902 10.6151
R20252 vdd.n2879 vdd.n2878 10.6151
R20253 vdd.n2880 vdd.n2879 10.6151
R20254 vdd.n2880 vdd.n889 10.6151
R20255 vdd.n2890 vdd.n889 10.6151
R20256 vdd.n2891 vdd.n2890 10.6151
R20257 vdd.n2892 vdd.n2891 10.6151
R20258 vdd.n2892 vdd.n878 10.6151
R20259 vdd.n2902 vdd.n878 10.6151
R20260 vdd.n2903 vdd.n2902 10.6151
R20261 vdd.n2904 vdd.n2903 10.6151
R20262 vdd.n2904 vdd.n866 10.6151
R20263 vdd.n2914 vdd.n866 10.6151
R20264 vdd.n2915 vdd.n2914 10.6151
R20265 vdd.n2916 vdd.n2915 10.6151
R20266 vdd.n2916 vdd.n855 10.6151
R20267 vdd.n2928 vdd.n855 10.6151
R20268 vdd.n2929 vdd.n2928 10.6151
R20269 vdd.n2930 vdd.n2929 10.6151
R20270 vdd.n2930 vdd.n841 10.6151
R20271 vdd.n2985 vdd.n841 10.6151
R20272 vdd.n2986 vdd.n2985 10.6151
R20273 vdd.n2987 vdd.n2986 10.6151
R20274 vdd.n2987 vdd.n810 10.6151
R20275 vdd.n3057 vdd.n810 10.6151
R20276 vdd.n3056 vdd.n3055 10.6151
R20277 vdd.n3055 vdd.n811 10.6151
R20278 vdd.n812 vdd.n811 10.6151
R20279 vdd.n3048 vdd.n812 10.6151
R20280 vdd.n3048 vdd.n3047 10.6151
R20281 vdd.n3047 vdd.n3046 10.6151
R20282 vdd.n3046 vdd.n814 10.6151
R20283 vdd.n3041 vdd.n814 10.6151
R20284 vdd.n3041 vdd.n3040 10.6151
R20285 vdd.n3040 vdd.n3039 10.6151
R20286 vdd.n3039 vdd.n817 10.6151
R20287 vdd.n3034 vdd.n817 10.6151
R20288 vdd.n3034 vdd.n3033 10.6151
R20289 vdd.n3033 vdd.n3032 10.6151
R20290 vdd.n3032 vdd.n820 10.6151
R20291 vdd.n3027 vdd.n820 10.6151
R20292 vdd.n3027 vdd.n731 10.6151
R20293 vdd.n3023 vdd.n731 10.6151
R20294 vdd.n3023 vdd.n3022 10.6151
R20295 vdd.n3022 vdd.n3021 10.6151
R20296 vdd.n3021 vdd.n823 10.6151
R20297 vdd.n3016 vdd.n823 10.6151
R20298 vdd.n3016 vdd.n3015 10.6151
R20299 vdd.n3015 vdd.n3014 10.6151
R20300 vdd.n3014 vdd.n826 10.6151
R20301 vdd.n3009 vdd.n826 10.6151
R20302 vdd.n3009 vdd.n3008 10.6151
R20303 vdd.n3008 vdd.n3007 10.6151
R20304 vdd.n3007 vdd.n829 10.6151
R20305 vdd.n3002 vdd.n829 10.6151
R20306 vdd.n3002 vdd.n3001 10.6151
R20307 vdd.n2999 vdd.n834 10.6151
R20308 vdd.n2994 vdd.n834 10.6151
R20309 vdd.n2975 vdd.n2936 10.6151
R20310 vdd.n2970 vdd.n2936 10.6151
R20311 vdd.n2970 vdd.n2969 10.6151
R20312 vdd.n2969 vdd.n2968 10.6151
R20313 vdd.n2968 vdd.n2938 10.6151
R20314 vdd.n2963 vdd.n2938 10.6151
R20315 vdd.n2963 vdd.n2962 10.6151
R20316 vdd.n2962 vdd.n2961 10.6151
R20317 vdd.n2961 vdd.n2941 10.6151
R20318 vdd.n2956 vdd.n2941 10.6151
R20319 vdd.n2956 vdd.n2955 10.6151
R20320 vdd.n2955 vdd.n2954 10.6151
R20321 vdd.n2954 vdd.n2944 10.6151
R20322 vdd.n2949 vdd.n2944 10.6151
R20323 vdd.n2949 vdd.n2948 10.6151
R20324 vdd.n2948 vdd.n785 10.6151
R20325 vdd.n3092 vdd.n785 10.6151
R20326 vdd.n3092 vdd.n786 10.6151
R20327 vdd.n788 vdd.n786 10.6151
R20328 vdd.n3085 vdd.n788 10.6151
R20329 vdd.n3085 vdd.n3084 10.6151
R20330 vdd.n3084 vdd.n3083 10.6151
R20331 vdd.n3083 vdd.n790 10.6151
R20332 vdd.n3078 vdd.n790 10.6151
R20333 vdd.n3078 vdd.n3077 10.6151
R20334 vdd.n3077 vdd.n3076 10.6151
R20335 vdd.n3076 vdd.n793 10.6151
R20336 vdd.n3071 vdd.n793 10.6151
R20337 vdd.n3071 vdd.n3070 10.6151
R20338 vdd.n3070 vdd.n3069 10.6151
R20339 vdd.n3069 vdd.n796 10.6151
R20340 vdd.n3064 vdd.n3063 10.6151
R20341 vdd.n3063 vdd.n3062 10.6151
R20342 vdd.n2710 vdd.n2708 10.6151
R20343 vdd.n2711 vdd.n2710 10.6151
R20344 vdd.n2779 vdd.n2711 10.6151
R20345 vdd.n2779 vdd.n2778 10.6151
R20346 vdd.n2778 vdd.n2777 10.6151
R20347 vdd.n2777 vdd.n2775 10.6151
R20348 vdd.n2775 vdd.n2774 10.6151
R20349 vdd.n2774 vdd.n2772 10.6151
R20350 vdd.n2772 vdd.n2771 10.6151
R20351 vdd.n2771 vdd.n2769 10.6151
R20352 vdd.n2769 vdd.n2768 10.6151
R20353 vdd.n2768 vdd.n2766 10.6151
R20354 vdd.n2766 vdd.n2765 10.6151
R20355 vdd.n2765 vdd.n2763 10.6151
R20356 vdd.n2763 vdd.n2762 10.6151
R20357 vdd.n2762 vdd.n2728 10.6151
R20358 vdd.n2728 vdd.n2727 10.6151
R20359 vdd.n2727 vdd.n2725 10.6151
R20360 vdd.n2725 vdd.n2724 10.6151
R20361 vdd.n2724 vdd.n2722 10.6151
R20362 vdd.n2722 vdd.n2721 10.6151
R20363 vdd.n2721 vdd.n2719 10.6151
R20364 vdd.n2719 vdd.n2718 10.6151
R20365 vdd.n2718 vdd.n2716 10.6151
R20366 vdd.n2716 vdd.n2715 10.6151
R20367 vdd.n2715 vdd.n2713 10.6151
R20368 vdd.n2713 vdd.n2712 10.6151
R20369 vdd.n2712 vdd.n802 10.6151
R20370 vdd.n2861 vdd.n2860 10.6151
R20371 vdd.n2860 vdd.n917 10.6151
R20372 vdd.n2645 vdd.n917 10.6151
R20373 vdd.n2648 vdd.n2645 10.6151
R20374 vdd.n2649 vdd.n2648 10.6151
R20375 vdd.n2652 vdd.n2649 10.6151
R20376 vdd.n2653 vdd.n2652 10.6151
R20377 vdd.n2656 vdd.n2653 10.6151
R20378 vdd.n2657 vdd.n2656 10.6151
R20379 vdd.n2660 vdd.n2657 10.6151
R20380 vdd.n2661 vdd.n2660 10.6151
R20381 vdd.n2664 vdd.n2661 10.6151
R20382 vdd.n2665 vdd.n2664 10.6151
R20383 vdd.n2668 vdd.n2665 10.6151
R20384 vdd.n2669 vdd.n2668 10.6151
R20385 vdd.n2672 vdd.n2669 10.6151
R20386 vdd.n2673 vdd.n2672 10.6151
R20387 vdd.n2676 vdd.n2673 10.6151
R20388 vdd.n2677 vdd.n2676 10.6151
R20389 vdd.n2680 vdd.n2677 10.6151
R20390 vdd.n2681 vdd.n2680 10.6151
R20391 vdd.n2684 vdd.n2681 10.6151
R20392 vdd.n2685 vdd.n2684 10.6151
R20393 vdd.n2688 vdd.n2685 10.6151
R20394 vdd.n2689 vdd.n2688 10.6151
R20395 vdd.n2692 vdd.n2689 10.6151
R20396 vdd.n2693 vdd.n2692 10.6151
R20397 vdd.n2696 vdd.n2693 10.6151
R20398 vdd.n2697 vdd.n2696 10.6151
R20399 vdd.n2700 vdd.n2697 10.6151
R20400 vdd.n2701 vdd.n2700 10.6151
R20401 vdd.n2706 vdd.n2704 10.6151
R20402 vdd.n2707 vdd.n2706 10.6151
R20403 vdd.n2862 vdd.n907 10.6151
R20404 vdd.n2872 vdd.n907 10.6151
R20405 vdd.n2873 vdd.n2872 10.6151
R20406 vdd.n2874 vdd.n2873 10.6151
R20407 vdd.n2874 vdd.n895 10.6151
R20408 vdd.n2884 vdd.n895 10.6151
R20409 vdd.n2885 vdd.n2884 10.6151
R20410 vdd.n2886 vdd.n2885 10.6151
R20411 vdd.n2886 vdd.n884 10.6151
R20412 vdd.n2896 vdd.n884 10.6151
R20413 vdd.n2897 vdd.n2896 10.6151
R20414 vdd.n2898 vdd.n2897 10.6151
R20415 vdd.n2898 vdd.n872 10.6151
R20416 vdd.n2908 vdd.n872 10.6151
R20417 vdd.n2909 vdd.n2908 10.6151
R20418 vdd.n2910 vdd.n2909 10.6151
R20419 vdd.n2910 vdd.n861 10.6151
R20420 vdd.n2920 vdd.n861 10.6151
R20421 vdd.n2921 vdd.n2920 10.6151
R20422 vdd.n2924 vdd.n2921 10.6151
R20423 vdd.n2934 vdd.n849 10.6151
R20424 vdd.n2935 vdd.n2934 10.6151
R20425 vdd.n2981 vdd.n2935 10.6151
R20426 vdd.n2981 vdd.n2980 10.6151
R20427 vdd.n2980 vdd.n2979 10.6151
R20428 vdd.n2979 vdd.n2978 10.6151
R20429 vdd.n2978 vdd.n2976 10.6151
R20430 vdd.n2373 vdd.n1041 10.6151
R20431 vdd.n2383 vdd.n1041 10.6151
R20432 vdd.n2384 vdd.n2383 10.6151
R20433 vdd.n2385 vdd.n2384 10.6151
R20434 vdd.n2385 vdd.n1028 10.6151
R20435 vdd.n2395 vdd.n1028 10.6151
R20436 vdd.n2396 vdd.n2395 10.6151
R20437 vdd.n2398 vdd.n1016 10.6151
R20438 vdd.n2408 vdd.n1016 10.6151
R20439 vdd.n2409 vdd.n2408 10.6151
R20440 vdd.n2410 vdd.n2409 10.6151
R20441 vdd.n2410 vdd.n1004 10.6151
R20442 vdd.n2420 vdd.n1004 10.6151
R20443 vdd.n2421 vdd.n2420 10.6151
R20444 vdd.n2422 vdd.n2421 10.6151
R20445 vdd.n2422 vdd.n993 10.6151
R20446 vdd.n2432 vdd.n993 10.6151
R20447 vdd.n2433 vdd.n2432 10.6151
R20448 vdd.n2434 vdd.n2433 10.6151
R20449 vdd.n2434 vdd.n981 10.6151
R20450 vdd.n2444 vdd.n981 10.6151
R20451 vdd.n2445 vdd.n2444 10.6151
R20452 vdd.n2448 vdd.n2445 10.6151
R20453 vdd.n2448 vdd.n2447 10.6151
R20454 vdd.n2447 vdd.n2446 10.6151
R20455 vdd.n2446 vdd.n964 10.6151
R20456 vdd.n2530 vdd.n964 10.6151
R20457 vdd.n2529 vdd.n2528 10.6151
R20458 vdd.n2528 vdd.n2525 10.6151
R20459 vdd.n2525 vdd.n2524 10.6151
R20460 vdd.n2524 vdd.n2521 10.6151
R20461 vdd.n2521 vdd.n2520 10.6151
R20462 vdd.n2520 vdd.n2517 10.6151
R20463 vdd.n2517 vdd.n2516 10.6151
R20464 vdd.n2516 vdd.n2513 10.6151
R20465 vdd.n2513 vdd.n2512 10.6151
R20466 vdd.n2512 vdd.n2509 10.6151
R20467 vdd.n2509 vdd.n2508 10.6151
R20468 vdd.n2508 vdd.n2505 10.6151
R20469 vdd.n2505 vdd.n2504 10.6151
R20470 vdd.n2504 vdd.n2501 10.6151
R20471 vdd.n2501 vdd.n2500 10.6151
R20472 vdd.n2500 vdd.n2497 10.6151
R20473 vdd.n2497 vdd.n2496 10.6151
R20474 vdd.n2496 vdd.n2493 10.6151
R20475 vdd.n2493 vdd.n2492 10.6151
R20476 vdd.n2492 vdd.n2489 10.6151
R20477 vdd.n2489 vdd.n2488 10.6151
R20478 vdd.n2488 vdd.n2485 10.6151
R20479 vdd.n2485 vdd.n2484 10.6151
R20480 vdd.n2484 vdd.n2481 10.6151
R20481 vdd.n2481 vdd.n2480 10.6151
R20482 vdd.n2480 vdd.n2477 10.6151
R20483 vdd.n2477 vdd.n2476 10.6151
R20484 vdd.n2476 vdd.n2473 10.6151
R20485 vdd.n2473 vdd.n2472 10.6151
R20486 vdd.n2472 vdd.n2469 10.6151
R20487 vdd.n2469 vdd.n2468 10.6151
R20488 vdd.n2465 vdd.n2464 10.6151
R20489 vdd.n2464 vdd.n2462 10.6151
R20490 vdd.n2221 vdd.n2219 10.6151
R20491 vdd.n2222 vdd.n2221 10.6151
R20492 vdd.n2224 vdd.n2222 10.6151
R20493 vdd.n2225 vdd.n2224 10.6151
R20494 vdd.n2227 vdd.n2225 10.6151
R20495 vdd.n2228 vdd.n2227 10.6151
R20496 vdd.n2230 vdd.n2228 10.6151
R20497 vdd.n2231 vdd.n2230 10.6151
R20498 vdd.n2233 vdd.n2231 10.6151
R20499 vdd.n2234 vdd.n2233 10.6151
R20500 vdd.n2236 vdd.n2234 10.6151
R20501 vdd.n2237 vdd.n2236 10.6151
R20502 vdd.n2255 vdd.n2237 10.6151
R20503 vdd.n2255 vdd.n2254 10.6151
R20504 vdd.n2254 vdd.n2253 10.6151
R20505 vdd.n2253 vdd.n2251 10.6151
R20506 vdd.n2251 vdd.n2250 10.6151
R20507 vdd.n2250 vdd.n2248 10.6151
R20508 vdd.n2248 vdd.n2247 10.6151
R20509 vdd.n2247 vdd.n2245 10.6151
R20510 vdd.n2245 vdd.n2244 10.6151
R20511 vdd.n2244 vdd.n2242 10.6151
R20512 vdd.n2242 vdd.n2241 10.6151
R20513 vdd.n2241 vdd.n2239 10.6151
R20514 vdd.n2239 vdd.n2238 10.6151
R20515 vdd.n2238 vdd.n968 10.6151
R20516 vdd.n2460 vdd.n968 10.6151
R20517 vdd.n2461 vdd.n2460 10.6151
R20518 vdd.n2372 vdd.n2371 10.6151
R20519 vdd.n2371 vdd.n1053 10.6151
R20520 vdd.n2365 vdd.n1053 10.6151
R20521 vdd.n2365 vdd.n2364 10.6151
R20522 vdd.n2364 vdd.n2363 10.6151
R20523 vdd.n2363 vdd.n1055 10.6151
R20524 vdd.n2357 vdd.n1055 10.6151
R20525 vdd.n2357 vdd.n2356 10.6151
R20526 vdd.n2356 vdd.n2355 10.6151
R20527 vdd.n2355 vdd.n1057 10.6151
R20528 vdd.n2349 vdd.n1057 10.6151
R20529 vdd.n2349 vdd.n2348 10.6151
R20530 vdd.n2348 vdd.n2347 10.6151
R20531 vdd.n2347 vdd.n1059 10.6151
R20532 vdd.n2341 vdd.n1059 10.6151
R20533 vdd.n2341 vdd.n2340 10.6151
R20534 vdd.n2340 vdd.n2339 10.6151
R20535 vdd.n2339 vdd.n1063 10.6151
R20536 vdd.n2187 vdd.n1063 10.6151
R20537 vdd.n2188 vdd.n2187 10.6151
R20538 vdd.n2188 vdd.n2183 10.6151
R20539 vdd.n2194 vdd.n2183 10.6151
R20540 vdd.n2195 vdd.n2194 10.6151
R20541 vdd.n2196 vdd.n2195 10.6151
R20542 vdd.n2196 vdd.n2181 10.6151
R20543 vdd.n2202 vdd.n2181 10.6151
R20544 vdd.n2203 vdd.n2202 10.6151
R20545 vdd.n2204 vdd.n2203 10.6151
R20546 vdd.n2204 vdd.n2179 10.6151
R20547 vdd.n2210 vdd.n2179 10.6151
R20548 vdd.n2211 vdd.n2210 10.6151
R20549 vdd.n2213 vdd.n2175 10.6151
R20550 vdd.n2218 vdd.n2175 10.6151
R20551 vdd.n1851 vdd.t19 10.5435
R20552 vdd.n656 vdd.t129 10.5435
R20553 vdd.n316 vdd.n298 10.4732
R20554 vdd.n257 vdd.n239 10.4732
R20555 vdd.n214 vdd.n196 10.4732
R20556 vdd.n155 vdd.n137 10.4732
R20557 vdd.n113 vdd.n95 10.4732
R20558 vdd.n54 vdd.n36 10.4732
R20559 vdd.n1735 vdd.n1717 10.4732
R20560 vdd.n1794 vdd.n1776 10.4732
R20561 vdd.n1633 vdd.n1615 10.4732
R20562 vdd.n1692 vdd.n1674 10.4732
R20563 vdd.n1532 vdd.n1514 10.4732
R20564 vdd.n1591 vdd.n1573 10.4732
R20565 vdd.t109 vdd.n1825 10.3167
R20566 vdd.n3300 vdd.t72 10.3167
R20567 vdd.n1502 vdd.t39 10.09
R20568 vdd.n3394 vdd.t37 10.09
R20569 vdd.t106 vdd.n1155 9.86327
R20570 vdd.n3385 vdd.t35 9.86327
R20571 vdd.n315 vdd.n300 9.69747
R20572 vdd.n256 vdd.n241 9.69747
R20573 vdd.n213 vdd.n198 9.69747
R20574 vdd.n154 vdd.n139 9.69747
R20575 vdd.n112 vdd.n97 9.69747
R20576 vdd.n53 vdd.n38 9.69747
R20577 vdd.n1734 vdd.n1719 9.69747
R20578 vdd.n1793 vdd.n1778 9.69747
R20579 vdd.n1632 vdd.n1617 9.69747
R20580 vdd.n1691 vdd.n1676 9.69747
R20581 vdd.n1531 vdd.n1516 9.69747
R20582 vdd.n1590 vdd.n1575 9.69747
R20583 vdd.n2315 vdd.n2314 9.67831
R20584 vdd.n3216 vdd.n731 9.67831
R20585 vdd.n3093 vdd.n3092 9.67831
R20586 vdd.n2339 vdd.n2338 9.67831
R20587 vdd.n1461 vdd.t55 9.63654
R20588 vdd.n3331 vdd.t33 9.63654
R20589 vdd.n331 vdd.n330 9.45567
R20590 vdd.n272 vdd.n271 9.45567
R20591 vdd.n229 vdd.n228 9.45567
R20592 vdd.n170 vdd.n169 9.45567
R20593 vdd.n128 vdd.n127 9.45567
R20594 vdd.n69 vdd.n68 9.45567
R20595 vdd.n1750 vdd.n1749 9.45567
R20596 vdd.n1809 vdd.n1808 9.45567
R20597 vdd.n1648 vdd.n1647 9.45567
R20598 vdd.n1707 vdd.n1706 9.45567
R20599 vdd.n1547 vdd.n1546 9.45567
R20600 vdd.n1606 vdd.n1605 9.45567
R20601 vdd.n1435 vdd.t21 9.40981
R20602 vdd.n3363 vdd.t79 9.40981
R20603 vdd.n2075 vdd.n1929 9.3005
R20604 vdd.n2074 vdd.n2073 9.3005
R20605 vdd.n1935 vdd.n1934 9.3005
R20606 vdd.n2068 vdd.n1939 9.3005
R20607 vdd.n2067 vdd.n1940 9.3005
R20608 vdd.n2066 vdd.n1941 9.3005
R20609 vdd.n1945 vdd.n1942 9.3005
R20610 vdd.n2061 vdd.n1946 9.3005
R20611 vdd.n2060 vdd.n1947 9.3005
R20612 vdd.n2059 vdd.n1948 9.3005
R20613 vdd.n1952 vdd.n1949 9.3005
R20614 vdd.n2054 vdd.n1953 9.3005
R20615 vdd.n2053 vdd.n1954 9.3005
R20616 vdd.n2052 vdd.n1955 9.3005
R20617 vdd.n1959 vdd.n1956 9.3005
R20618 vdd.n2047 vdd.n1960 9.3005
R20619 vdd.n2046 vdd.n1961 9.3005
R20620 vdd.n2045 vdd.n1962 9.3005
R20621 vdd.n1966 vdd.n1963 9.3005
R20622 vdd.n2040 vdd.n1967 9.3005
R20623 vdd.n2039 vdd.n1968 9.3005
R20624 vdd.n2038 vdd.n2037 9.3005
R20625 vdd.n2036 vdd.n1969 9.3005
R20626 vdd.n2035 vdd.n2034 9.3005
R20627 vdd.n1975 vdd.n1974 9.3005
R20628 vdd.n2029 vdd.n1979 9.3005
R20629 vdd.n2028 vdd.n1980 9.3005
R20630 vdd.n2027 vdd.n1981 9.3005
R20631 vdd.n1985 vdd.n1982 9.3005
R20632 vdd.n2022 vdd.n1986 9.3005
R20633 vdd.n2021 vdd.n1987 9.3005
R20634 vdd.n2020 vdd.n1988 9.3005
R20635 vdd.n1992 vdd.n1989 9.3005
R20636 vdd.n2015 vdd.n1993 9.3005
R20637 vdd.n2014 vdd.n1994 9.3005
R20638 vdd.n2013 vdd.n1995 9.3005
R20639 vdd.n1997 vdd.n1996 9.3005
R20640 vdd.n2008 vdd.n1064 9.3005
R20641 vdd.n2077 vdd.n2076 9.3005
R20642 vdd.n2101 vdd.n2100 9.3005
R20643 vdd.n1907 vdd.n1906 9.3005
R20644 vdd.n1912 vdd.n1910 9.3005
R20645 vdd.n2093 vdd.n1913 9.3005
R20646 vdd.n2092 vdd.n1914 9.3005
R20647 vdd.n2091 vdd.n1915 9.3005
R20648 vdd.n1919 vdd.n1916 9.3005
R20649 vdd.n2086 vdd.n1920 9.3005
R20650 vdd.n2085 vdd.n1921 9.3005
R20651 vdd.n2084 vdd.n1922 9.3005
R20652 vdd.n1926 vdd.n1923 9.3005
R20653 vdd.n2079 vdd.n1927 9.3005
R20654 vdd.n2078 vdd.n1928 9.3005
R20655 vdd.n2323 vdd.n1900 9.3005
R20656 vdd.n2325 vdd.n2324 9.3005
R20657 vdd.n1815 vdd.n1814 9.3005
R20658 vdd.n1124 vdd.n1123 9.3005
R20659 vdd.n1829 vdd.n1828 9.3005
R20660 vdd.n1830 vdd.n1122 9.3005
R20661 vdd.n1832 vdd.n1831 9.3005
R20662 vdd.n1113 vdd.n1112 9.3005
R20663 vdd.n1846 vdd.n1845 9.3005
R20664 vdd.n1847 vdd.n1111 9.3005
R20665 vdd.n1849 vdd.n1848 9.3005
R20666 vdd.n1102 vdd.n1101 9.3005
R20667 vdd.n1862 vdd.n1861 9.3005
R20668 vdd.n1863 vdd.n1100 9.3005
R20669 vdd.n1865 vdd.n1864 9.3005
R20670 vdd.n1090 vdd.n1089 9.3005
R20671 vdd.n1879 vdd.n1878 9.3005
R20672 vdd.n1880 vdd.n1088 9.3005
R20673 vdd.n1882 vdd.n1881 9.3005
R20674 vdd.n1078 vdd.n1077 9.3005
R20675 vdd.n1898 vdd.n1897 9.3005
R20676 vdd.n1899 vdd.n1076 9.3005
R20677 vdd.n2327 vdd.n2326 9.3005
R20678 vdd.n307 vdd.n306 9.3005
R20679 vdd.n302 vdd.n301 9.3005
R20680 vdd.n313 vdd.n312 9.3005
R20681 vdd.n315 vdd.n314 9.3005
R20682 vdd.n298 vdd.n297 9.3005
R20683 vdd.n321 vdd.n320 9.3005
R20684 vdd.n323 vdd.n322 9.3005
R20685 vdd.n295 vdd.n292 9.3005
R20686 vdd.n330 vdd.n329 9.3005
R20687 vdd.n248 vdd.n247 9.3005
R20688 vdd.n243 vdd.n242 9.3005
R20689 vdd.n254 vdd.n253 9.3005
R20690 vdd.n256 vdd.n255 9.3005
R20691 vdd.n239 vdd.n238 9.3005
R20692 vdd.n262 vdd.n261 9.3005
R20693 vdd.n264 vdd.n263 9.3005
R20694 vdd.n236 vdd.n233 9.3005
R20695 vdd.n271 vdd.n270 9.3005
R20696 vdd.n205 vdd.n204 9.3005
R20697 vdd.n200 vdd.n199 9.3005
R20698 vdd.n211 vdd.n210 9.3005
R20699 vdd.n213 vdd.n212 9.3005
R20700 vdd.n196 vdd.n195 9.3005
R20701 vdd.n219 vdd.n218 9.3005
R20702 vdd.n221 vdd.n220 9.3005
R20703 vdd.n193 vdd.n190 9.3005
R20704 vdd.n228 vdd.n227 9.3005
R20705 vdd.n146 vdd.n145 9.3005
R20706 vdd.n141 vdd.n140 9.3005
R20707 vdd.n152 vdd.n151 9.3005
R20708 vdd.n154 vdd.n153 9.3005
R20709 vdd.n137 vdd.n136 9.3005
R20710 vdd.n160 vdd.n159 9.3005
R20711 vdd.n162 vdd.n161 9.3005
R20712 vdd.n134 vdd.n131 9.3005
R20713 vdd.n169 vdd.n168 9.3005
R20714 vdd.n104 vdd.n103 9.3005
R20715 vdd.n99 vdd.n98 9.3005
R20716 vdd.n110 vdd.n109 9.3005
R20717 vdd.n112 vdd.n111 9.3005
R20718 vdd.n95 vdd.n94 9.3005
R20719 vdd.n118 vdd.n117 9.3005
R20720 vdd.n120 vdd.n119 9.3005
R20721 vdd.n92 vdd.n89 9.3005
R20722 vdd.n127 vdd.n126 9.3005
R20723 vdd.n45 vdd.n44 9.3005
R20724 vdd.n40 vdd.n39 9.3005
R20725 vdd.n51 vdd.n50 9.3005
R20726 vdd.n53 vdd.n52 9.3005
R20727 vdd.n36 vdd.n35 9.3005
R20728 vdd.n59 vdd.n58 9.3005
R20729 vdd.n61 vdd.n60 9.3005
R20730 vdd.n33 vdd.n30 9.3005
R20731 vdd.n68 vdd.n67 9.3005
R20732 vdd.n3138 vdd.n3137 9.3005
R20733 vdd.n3141 vdd.n766 9.3005
R20734 vdd.n3142 vdd.n765 9.3005
R20735 vdd.n3145 vdd.n764 9.3005
R20736 vdd.n3146 vdd.n763 9.3005
R20737 vdd.n3149 vdd.n762 9.3005
R20738 vdd.n3150 vdd.n761 9.3005
R20739 vdd.n3153 vdd.n760 9.3005
R20740 vdd.n3154 vdd.n759 9.3005
R20741 vdd.n3157 vdd.n758 9.3005
R20742 vdd.n3158 vdd.n757 9.3005
R20743 vdd.n3161 vdd.n756 9.3005
R20744 vdd.n3162 vdd.n755 9.3005
R20745 vdd.n3165 vdd.n754 9.3005
R20746 vdd.n3166 vdd.n753 9.3005
R20747 vdd.n3169 vdd.n752 9.3005
R20748 vdd.n3170 vdd.n751 9.3005
R20749 vdd.n3173 vdd.n750 9.3005
R20750 vdd.n3174 vdd.n749 9.3005
R20751 vdd.n3177 vdd.n748 9.3005
R20752 vdd.n3181 vdd.n3180 9.3005
R20753 vdd.n3182 vdd.n747 9.3005
R20754 vdd.n3186 vdd.n3183 9.3005
R20755 vdd.n3189 vdd.n746 9.3005
R20756 vdd.n3190 vdd.n745 9.3005
R20757 vdd.n3193 vdd.n744 9.3005
R20758 vdd.n3194 vdd.n743 9.3005
R20759 vdd.n3197 vdd.n742 9.3005
R20760 vdd.n3198 vdd.n741 9.3005
R20761 vdd.n3201 vdd.n740 9.3005
R20762 vdd.n3202 vdd.n739 9.3005
R20763 vdd.n3205 vdd.n738 9.3005
R20764 vdd.n3206 vdd.n737 9.3005
R20765 vdd.n3209 vdd.n736 9.3005
R20766 vdd.n3210 vdd.n735 9.3005
R20767 vdd.n3213 vdd.n730 9.3005
R20768 vdd.n3219 vdd.n727 9.3005
R20769 vdd.n3220 vdd.n726 9.3005
R20770 vdd.n3234 vdd.n3233 9.3005
R20771 vdd.n3235 vdd.n681 9.3005
R20772 vdd.n3237 vdd.n3236 9.3005
R20773 vdd.n671 vdd.n670 9.3005
R20774 vdd.n3251 vdd.n3250 9.3005
R20775 vdd.n3252 vdd.n669 9.3005
R20776 vdd.n3254 vdd.n3253 9.3005
R20777 vdd.n660 vdd.n659 9.3005
R20778 vdd.n3267 vdd.n3266 9.3005
R20779 vdd.n3268 vdd.n658 9.3005
R20780 vdd.n3270 vdd.n3269 9.3005
R20781 vdd.n648 vdd.n647 9.3005
R20782 vdd.n3284 vdd.n3283 9.3005
R20783 vdd.n3285 vdd.n646 9.3005
R20784 vdd.n3287 vdd.n3286 9.3005
R20785 vdd.n637 vdd.n636 9.3005
R20786 vdd.n3303 vdd.n3302 9.3005
R20787 vdd.n3304 vdd.n635 9.3005
R20788 vdd.n3306 vdd.n3305 9.3005
R20789 vdd.n336 vdd.n334 9.3005
R20790 vdd.n683 vdd.n682 9.3005
R20791 vdd.n3398 vdd.n3397 9.3005
R20792 vdd.n337 vdd.n335 9.3005
R20793 vdd.n3391 vdd.n346 9.3005
R20794 vdd.n3390 vdd.n347 9.3005
R20795 vdd.n3389 vdd.n348 9.3005
R20796 vdd.n355 vdd.n349 9.3005
R20797 vdd.n3383 vdd.n356 9.3005
R20798 vdd.n3382 vdd.n357 9.3005
R20799 vdd.n3381 vdd.n358 9.3005
R20800 vdd.n366 vdd.n359 9.3005
R20801 vdd.n3375 vdd.n367 9.3005
R20802 vdd.n3374 vdd.n368 9.3005
R20803 vdd.n3373 vdd.n369 9.3005
R20804 vdd.n377 vdd.n370 9.3005
R20805 vdd.n3367 vdd.n378 9.3005
R20806 vdd.n3366 vdd.n379 9.3005
R20807 vdd.n3365 vdd.n380 9.3005
R20808 vdd.n388 vdd.n381 9.3005
R20809 vdd.n3359 vdd.n389 9.3005
R20810 vdd.n3358 vdd.n390 9.3005
R20811 vdd.n3357 vdd.n391 9.3005
R20812 vdd.n466 vdd.n463 9.3005
R20813 vdd.n470 vdd.n469 9.3005
R20814 vdd.n471 vdd.n462 9.3005
R20815 vdd.n475 vdd.n472 9.3005
R20816 vdd.n476 vdd.n461 9.3005
R20817 vdd.n480 vdd.n479 9.3005
R20818 vdd.n481 vdd.n460 9.3005
R20819 vdd.n485 vdd.n482 9.3005
R20820 vdd.n486 vdd.n459 9.3005
R20821 vdd.n490 vdd.n489 9.3005
R20822 vdd.n491 vdd.n458 9.3005
R20823 vdd.n495 vdd.n492 9.3005
R20824 vdd.n496 vdd.n457 9.3005
R20825 vdd.n500 vdd.n499 9.3005
R20826 vdd.n501 vdd.n456 9.3005
R20827 vdd.n505 vdd.n502 9.3005
R20828 vdd.n506 vdd.n455 9.3005
R20829 vdd.n510 vdd.n509 9.3005
R20830 vdd.n511 vdd.n454 9.3005
R20831 vdd.n515 vdd.n512 9.3005
R20832 vdd.n516 vdd.n451 9.3005
R20833 vdd.n520 vdd.n519 9.3005
R20834 vdd.n521 vdd.n450 9.3005
R20835 vdd.n525 vdd.n522 9.3005
R20836 vdd.n526 vdd.n449 9.3005
R20837 vdd.n530 vdd.n529 9.3005
R20838 vdd.n531 vdd.n448 9.3005
R20839 vdd.n535 vdd.n532 9.3005
R20840 vdd.n536 vdd.n447 9.3005
R20841 vdd.n540 vdd.n539 9.3005
R20842 vdd.n541 vdd.n446 9.3005
R20843 vdd.n545 vdd.n542 9.3005
R20844 vdd.n546 vdd.n445 9.3005
R20845 vdd.n550 vdd.n549 9.3005
R20846 vdd.n551 vdd.n444 9.3005
R20847 vdd.n555 vdd.n552 9.3005
R20848 vdd.n556 vdd.n443 9.3005
R20849 vdd.n560 vdd.n559 9.3005
R20850 vdd.n561 vdd.n442 9.3005
R20851 vdd.n565 vdd.n562 9.3005
R20852 vdd.n566 vdd.n439 9.3005
R20853 vdd.n570 vdd.n569 9.3005
R20854 vdd.n571 vdd.n438 9.3005
R20855 vdd.n575 vdd.n572 9.3005
R20856 vdd.n576 vdd.n437 9.3005
R20857 vdd.n580 vdd.n579 9.3005
R20858 vdd.n581 vdd.n436 9.3005
R20859 vdd.n585 vdd.n582 9.3005
R20860 vdd.n586 vdd.n435 9.3005
R20861 vdd.n590 vdd.n589 9.3005
R20862 vdd.n591 vdd.n434 9.3005
R20863 vdd.n595 vdd.n592 9.3005
R20864 vdd.n596 vdd.n433 9.3005
R20865 vdd.n600 vdd.n599 9.3005
R20866 vdd.n601 vdd.n432 9.3005
R20867 vdd.n605 vdd.n602 9.3005
R20868 vdd.n606 vdd.n431 9.3005
R20869 vdd.n610 vdd.n609 9.3005
R20870 vdd.n611 vdd.n430 9.3005
R20871 vdd.n615 vdd.n612 9.3005
R20872 vdd.n617 vdd.n429 9.3005
R20873 vdd.n619 vdd.n618 9.3005
R20874 vdd.n3351 vdd.n3350 9.3005
R20875 vdd.n465 vdd.n464 9.3005
R20876 vdd.n3229 vdd.n3228 9.3005
R20877 vdd.n676 vdd.n675 9.3005
R20878 vdd.n3242 vdd.n3241 9.3005
R20879 vdd.n3243 vdd.n674 9.3005
R20880 vdd.n3245 vdd.n3244 9.3005
R20881 vdd.n666 vdd.n665 9.3005
R20882 vdd.n3259 vdd.n3258 9.3005
R20883 vdd.n3260 vdd.n664 9.3005
R20884 vdd.n3262 vdd.n3261 9.3005
R20885 vdd.n653 vdd.n652 9.3005
R20886 vdd.n3275 vdd.n3274 9.3005
R20887 vdd.n3276 vdd.n651 9.3005
R20888 vdd.n3278 vdd.n3277 9.3005
R20889 vdd.n642 vdd.n641 9.3005
R20890 vdd.n3292 vdd.n3291 9.3005
R20891 vdd.n3293 vdd.n640 9.3005
R20892 vdd.n3298 vdd.n3294 9.3005
R20893 vdd.n3297 vdd.n3296 9.3005
R20894 vdd.n3295 vdd.n631 9.3005
R20895 vdd.n3311 vdd.n630 9.3005
R20896 vdd.n3313 vdd.n3312 9.3005
R20897 vdd.n3314 vdd.n629 9.3005
R20898 vdd.n3316 vdd.n3315 9.3005
R20899 vdd.n3318 vdd.n628 9.3005
R20900 vdd.n3320 vdd.n3319 9.3005
R20901 vdd.n3321 vdd.n627 9.3005
R20902 vdd.n3323 vdd.n3322 9.3005
R20903 vdd.n3325 vdd.n626 9.3005
R20904 vdd.n3327 vdd.n3326 9.3005
R20905 vdd.n3328 vdd.n625 9.3005
R20906 vdd.n3330 vdd.n3329 9.3005
R20907 vdd.n3333 vdd.n624 9.3005
R20908 vdd.n3335 vdd.n3334 9.3005
R20909 vdd.n3336 vdd.n623 9.3005
R20910 vdd.n3338 vdd.n3337 9.3005
R20911 vdd.n3340 vdd.n622 9.3005
R20912 vdd.n3342 vdd.n3341 9.3005
R20913 vdd.n3343 vdd.n621 9.3005
R20914 vdd.n3345 vdd.n3344 9.3005
R20915 vdd.n3347 vdd.n620 9.3005
R20916 vdd.n3349 vdd.n3348 9.3005
R20917 vdd.n3227 vdd.n686 9.3005
R20918 vdd.n3226 vdd.n3225 9.3005
R20919 vdd.n3095 vdd.n687 9.3005
R20920 vdd.n3104 vdd.n783 9.3005
R20921 vdd.n3107 vdd.n782 9.3005
R20922 vdd.n3108 vdd.n781 9.3005
R20923 vdd.n3111 vdd.n780 9.3005
R20924 vdd.n3112 vdd.n779 9.3005
R20925 vdd.n3115 vdd.n778 9.3005
R20926 vdd.n3116 vdd.n777 9.3005
R20927 vdd.n3119 vdd.n776 9.3005
R20928 vdd.n3120 vdd.n775 9.3005
R20929 vdd.n3123 vdd.n774 9.3005
R20930 vdd.n3124 vdd.n773 9.3005
R20931 vdd.n3127 vdd.n772 9.3005
R20932 vdd.n3128 vdd.n771 9.3005
R20933 vdd.n3131 vdd.n770 9.3005
R20934 vdd.n3135 vdd.n3134 9.3005
R20935 vdd.n3136 vdd.n767 9.3005
R20936 vdd.n2337 vdd.n2336 9.3005
R20937 vdd.n2332 vdd.n1067 9.3005
R20938 vdd.n1430 vdd.n1429 9.3005
R20939 vdd.n1431 vdd.n1185 9.3005
R20940 vdd.n1433 vdd.n1432 9.3005
R20941 vdd.n1175 vdd.n1174 9.3005
R20942 vdd.n1447 vdd.n1446 9.3005
R20943 vdd.n1448 vdd.n1173 9.3005
R20944 vdd.n1450 vdd.n1449 9.3005
R20945 vdd.n1165 vdd.n1164 9.3005
R20946 vdd.n1464 vdd.n1463 9.3005
R20947 vdd.n1465 vdd.n1163 9.3005
R20948 vdd.n1467 vdd.n1466 9.3005
R20949 vdd.n1152 vdd.n1151 9.3005
R20950 vdd.n1480 vdd.n1479 9.3005
R20951 vdd.n1481 vdd.n1150 9.3005
R20952 vdd.n1483 vdd.n1482 9.3005
R20953 vdd.n1141 vdd.n1140 9.3005
R20954 vdd.n1497 vdd.n1496 9.3005
R20955 vdd.n1498 vdd.n1139 9.3005
R20956 vdd.n1500 vdd.n1499 9.3005
R20957 vdd.n1130 vdd.n1129 9.3005
R20958 vdd.n1820 vdd.n1819 9.3005
R20959 vdd.n1821 vdd.n1128 9.3005
R20960 vdd.n1823 vdd.n1822 9.3005
R20961 vdd.n1118 vdd.n1117 9.3005
R20962 vdd.n1837 vdd.n1836 9.3005
R20963 vdd.n1838 vdd.n1116 9.3005
R20964 vdd.n1840 vdd.n1839 9.3005
R20965 vdd.n1108 vdd.n1107 9.3005
R20966 vdd.n1854 vdd.n1853 9.3005
R20967 vdd.n1855 vdd.n1106 9.3005
R20968 vdd.n1857 vdd.n1856 9.3005
R20969 vdd.n1095 vdd.n1094 9.3005
R20970 vdd.n1870 vdd.n1869 9.3005
R20971 vdd.n1871 vdd.n1093 9.3005
R20972 vdd.n1873 vdd.n1872 9.3005
R20973 vdd.n1085 vdd.n1084 9.3005
R20974 vdd.n1887 vdd.n1886 9.3005
R20975 vdd.n1888 vdd.n1082 9.3005
R20976 vdd.n1892 vdd.n1891 9.3005
R20977 vdd.n1890 vdd.n1083 9.3005
R20978 vdd.n1889 vdd.n1072 9.3005
R20979 vdd.n1187 vdd.n1186 9.3005
R20980 vdd.n1323 vdd.n1322 9.3005
R20981 vdd.n1324 vdd.n1313 9.3005
R20982 vdd.n1326 vdd.n1325 9.3005
R20983 vdd.n1327 vdd.n1312 9.3005
R20984 vdd.n1329 vdd.n1328 9.3005
R20985 vdd.n1330 vdd.n1307 9.3005
R20986 vdd.n1332 vdd.n1331 9.3005
R20987 vdd.n1333 vdd.n1306 9.3005
R20988 vdd.n1335 vdd.n1334 9.3005
R20989 vdd.n1336 vdd.n1301 9.3005
R20990 vdd.n1338 vdd.n1337 9.3005
R20991 vdd.n1339 vdd.n1300 9.3005
R20992 vdd.n1341 vdd.n1340 9.3005
R20993 vdd.n1342 vdd.n1295 9.3005
R20994 vdd.n1344 vdd.n1343 9.3005
R20995 vdd.n1345 vdd.n1294 9.3005
R20996 vdd.n1347 vdd.n1346 9.3005
R20997 vdd.n1348 vdd.n1289 9.3005
R20998 vdd.n1350 vdd.n1349 9.3005
R20999 vdd.n1351 vdd.n1288 9.3005
R21000 vdd.n1353 vdd.n1352 9.3005
R21001 vdd.n1357 vdd.n1284 9.3005
R21002 vdd.n1359 vdd.n1358 9.3005
R21003 vdd.n1360 vdd.n1283 9.3005
R21004 vdd.n1362 vdd.n1361 9.3005
R21005 vdd.n1363 vdd.n1278 9.3005
R21006 vdd.n1365 vdd.n1364 9.3005
R21007 vdd.n1366 vdd.n1277 9.3005
R21008 vdd.n1368 vdd.n1367 9.3005
R21009 vdd.n1369 vdd.n1272 9.3005
R21010 vdd.n1371 vdd.n1370 9.3005
R21011 vdd.n1372 vdd.n1271 9.3005
R21012 vdd.n1374 vdd.n1373 9.3005
R21013 vdd.n1375 vdd.n1266 9.3005
R21014 vdd.n1377 vdd.n1376 9.3005
R21015 vdd.n1378 vdd.n1265 9.3005
R21016 vdd.n1380 vdd.n1379 9.3005
R21017 vdd.n1381 vdd.n1260 9.3005
R21018 vdd.n1383 vdd.n1382 9.3005
R21019 vdd.n1384 vdd.n1259 9.3005
R21020 vdd.n1386 vdd.n1385 9.3005
R21021 vdd.n1387 vdd.n1254 9.3005
R21022 vdd.n1389 vdd.n1388 9.3005
R21023 vdd.n1390 vdd.n1253 9.3005
R21024 vdd.n1392 vdd.n1391 9.3005
R21025 vdd.n1393 vdd.n1246 9.3005
R21026 vdd.n1395 vdd.n1394 9.3005
R21027 vdd.n1396 vdd.n1245 9.3005
R21028 vdd.n1398 vdd.n1397 9.3005
R21029 vdd.n1399 vdd.n1240 9.3005
R21030 vdd.n1401 vdd.n1400 9.3005
R21031 vdd.n1402 vdd.n1239 9.3005
R21032 vdd.n1404 vdd.n1403 9.3005
R21033 vdd.n1405 vdd.n1234 9.3005
R21034 vdd.n1407 vdd.n1406 9.3005
R21035 vdd.n1408 vdd.n1233 9.3005
R21036 vdd.n1410 vdd.n1409 9.3005
R21037 vdd.n1411 vdd.n1228 9.3005
R21038 vdd.n1413 vdd.n1412 9.3005
R21039 vdd.n1414 vdd.n1227 9.3005
R21040 vdd.n1416 vdd.n1415 9.3005
R21041 vdd.n1192 vdd.n1191 9.3005
R21042 vdd.n1422 vdd.n1421 9.3005
R21043 vdd.n1321 vdd.n1320 9.3005
R21044 vdd.n1425 vdd.n1424 9.3005
R21045 vdd.n1181 vdd.n1180 9.3005
R21046 vdd.n1439 vdd.n1438 9.3005
R21047 vdd.n1440 vdd.n1179 9.3005
R21048 vdd.n1442 vdd.n1441 9.3005
R21049 vdd.n1170 vdd.n1169 9.3005
R21050 vdd.n1456 vdd.n1455 9.3005
R21051 vdd.n1457 vdd.n1168 9.3005
R21052 vdd.n1459 vdd.n1458 9.3005
R21053 vdd.n1159 vdd.n1158 9.3005
R21054 vdd.n1472 vdd.n1471 9.3005
R21055 vdd.n1473 vdd.n1157 9.3005
R21056 vdd.n1475 vdd.n1474 9.3005
R21057 vdd.n1147 vdd.n1146 9.3005
R21058 vdd.n1489 vdd.n1488 9.3005
R21059 vdd.n1490 vdd.n1145 9.3005
R21060 vdd.n1492 vdd.n1491 9.3005
R21061 vdd.n1136 vdd.n1135 9.3005
R21062 vdd.n1505 vdd.n1504 9.3005
R21063 vdd.n1506 vdd.n1134 9.3005
R21064 vdd.n1423 vdd.n1190 9.3005
R21065 vdd.n1726 vdd.n1725 9.3005
R21066 vdd.n1721 vdd.n1720 9.3005
R21067 vdd.n1732 vdd.n1731 9.3005
R21068 vdd.n1734 vdd.n1733 9.3005
R21069 vdd.n1717 vdd.n1716 9.3005
R21070 vdd.n1740 vdd.n1739 9.3005
R21071 vdd.n1742 vdd.n1741 9.3005
R21072 vdd.n1714 vdd.n1711 9.3005
R21073 vdd.n1749 vdd.n1748 9.3005
R21074 vdd.n1785 vdd.n1784 9.3005
R21075 vdd.n1780 vdd.n1779 9.3005
R21076 vdd.n1791 vdd.n1790 9.3005
R21077 vdd.n1793 vdd.n1792 9.3005
R21078 vdd.n1776 vdd.n1775 9.3005
R21079 vdd.n1799 vdd.n1798 9.3005
R21080 vdd.n1801 vdd.n1800 9.3005
R21081 vdd.n1773 vdd.n1770 9.3005
R21082 vdd.n1808 vdd.n1807 9.3005
R21083 vdd.n1624 vdd.n1623 9.3005
R21084 vdd.n1619 vdd.n1618 9.3005
R21085 vdd.n1630 vdd.n1629 9.3005
R21086 vdd.n1632 vdd.n1631 9.3005
R21087 vdd.n1615 vdd.n1614 9.3005
R21088 vdd.n1638 vdd.n1637 9.3005
R21089 vdd.n1640 vdd.n1639 9.3005
R21090 vdd.n1612 vdd.n1609 9.3005
R21091 vdd.n1647 vdd.n1646 9.3005
R21092 vdd.n1683 vdd.n1682 9.3005
R21093 vdd.n1678 vdd.n1677 9.3005
R21094 vdd.n1689 vdd.n1688 9.3005
R21095 vdd.n1691 vdd.n1690 9.3005
R21096 vdd.n1674 vdd.n1673 9.3005
R21097 vdd.n1697 vdd.n1696 9.3005
R21098 vdd.n1699 vdd.n1698 9.3005
R21099 vdd.n1671 vdd.n1668 9.3005
R21100 vdd.n1706 vdd.n1705 9.3005
R21101 vdd.n1523 vdd.n1522 9.3005
R21102 vdd.n1518 vdd.n1517 9.3005
R21103 vdd.n1529 vdd.n1528 9.3005
R21104 vdd.n1531 vdd.n1530 9.3005
R21105 vdd.n1514 vdd.n1513 9.3005
R21106 vdd.n1537 vdd.n1536 9.3005
R21107 vdd.n1539 vdd.n1538 9.3005
R21108 vdd.n1511 vdd.n1508 9.3005
R21109 vdd.n1546 vdd.n1545 9.3005
R21110 vdd.n1582 vdd.n1581 9.3005
R21111 vdd.n1577 vdd.n1576 9.3005
R21112 vdd.n1588 vdd.n1587 9.3005
R21113 vdd.n1590 vdd.n1589 9.3005
R21114 vdd.n1573 vdd.n1572 9.3005
R21115 vdd.n1596 vdd.n1595 9.3005
R21116 vdd.n1598 vdd.n1597 9.3005
R21117 vdd.n1570 vdd.n1567 9.3005
R21118 vdd.n1605 vdd.n1604 9.3005
R21119 vdd.n1461 vdd.t53 9.18308
R21120 vdd.n3331 vdd.t121 9.18308
R21121 vdd.n1155 vdd.t104 8.95635
R21122 vdd.n2329 vdd.t218 8.95635
R21123 vdd.n723 vdd.t211 8.95635
R21124 vdd.t68 vdd.n3385 8.95635
R21125 vdd.n312 vdd.n311 8.92171
R21126 vdd.n253 vdd.n252 8.92171
R21127 vdd.n210 vdd.n209 8.92171
R21128 vdd.n151 vdd.n150 8.92171
R21129 vdd.n109 vdd.n108 8.92171
R21130 vdd.n50 vdd.n49 8.92171
R21131 vdd.n1731 vdd.n1730 8.92171
R21132 vdd.n1790 vdd.n1789 8.92171
R21133 vdd.n1629 vdd.n1628 8.92171
R21134 vdd.n1688 vdd.n1687 8.92171
R21135 vdd.n1528 vdd.n1527 8.92171
R21136 vdd.n1587 vdd.n1586 8.92171
R21137 vdd.n231 vdd.n129 8.81535
R21138 vdd.n1709 vdd.n1607 8.81535
R21139 vdd.n1502 vdd.t76 8.72962
R21140 vdd.t65 vdd.n3394 8.72962
R21141 vdd.n1825 vdd.t124 8.50289
R21142 vdd.n3300 vdd.t70 8.50289
R21143 vdd.n28 vdd.n14 8.42249
R21144 vdd.n1851 vdd.t62 8.27616
R21145 vdd.t60 vdd.n656 8.27616
R21146 vdd.n3400 vdd.n3399 8.16225
R21147 vdd.n1813 vdd.n1812 8.16225
R21148 vdd.n308 vdd.n302 8.14595
R21149 vdd.n249 vdd.n243 8.14595
R21150 vdd.n206 vdd.n200 8.14595
R21151 vdd.n147 vdd.n141 8.14595
R21152 vdd.n105 vdd.n99 8.14595
R21153 vdd.n46 vdd.n40 8.14595
R21154 vdd.n1727 vdd.n1721 8.14595
R21155 vdd.n1786 vdd.n1780 8.14595
R21156 vdd.n1625 vdd.n1619 8.14595
R21157 vdd.n1684 vdd.n1678 8.14595
R21158 vdd.n1524 vdd.n1518 8.14595
R21159 vdd.n1583 vdd.n1577 8.14595
R21160 vdd.n2923 vdd.n849 8.11757
R21161 vdd.n2397 vdd.n2396 8.11757
R21162 vdd.n1098 vdd.t148 8.04943
R21163 vdd.n3256 vdd.t102 8.04943
R21164 vdd.n2375 vdd.n1043 7.70933
R21165 vdd.n2381 vdd.n1043 7.70933
R21166 vdd.n2387 vdd.n1037 7.70933
R21167 vdd.n2387 vdd.n1030 7.70933
R21168 vdd.n2393 vdd.n1030 7.70933
R21169 vdd.n2393 vdd.n1033 7.70933
R21170 vdd.n2400 vdd.n1018 7.70933
R21171 vdd.n2406 vdd.n1018 7.70933
R21172 vdd.n2412 vdd.n1012 7.70933
R21173 vdd.n2418 vdd.n1008 7.70933
R21174 vdd.n2424 vdd.n1002 7.70933
R21175 vdd.n2436 vdd.n989 7.70933
R21176 vdd.n2442 vdd.n983 7.70933
R21177 vdd.n2442 vdd.n976 7.70933
R21178 vdd.n2450 vdd.n976 7.70933
R21179 vdd.n2457 vdd.t172 7.70933
R21180 vdd.n2532 vdd.t172 7.70933
R21181 vdd.n2864 vdd.t4 7.70933
R21182 vdd.n2870 vdd.t4 7.70933
R21183 vdd.n2876 vdd.n897 7.70933
R21184 vdd.n2882 vdd.n897 7.70933
R21185 vdd.n2882 vdd.n900 7.70933
R21186 vdd.n2888 vdd.n893 7.70933
R21187 vdd.n2900 vdd.n880 7.70933
R21188 vdd.n2906 vdd.n874 7.70933
R21189 vdd.n2912 vdd.n870 7.70933
R21190 vdd.n2918 vdd.n857 7.70933
R21191 vdd.n2926 vdd.n857 7.70933
R21192 vdd.n2932 vdd.n851 7.70933
R21193 vdd.n2932 vdd.n843 7.70933
R21194 vdd.n2983 vdd.n843 7.70933
R21195 vdd.n2983 vdd.n846 7.70933
R21196 vdd.n2989 vdd.n805 7.70933
R21197 vdd.n3059 vdd.n805 7.70933
R21198 vdd.n307 vdd.n304 7.3702
R21199 vdd.n248 vdd.n245 7.3702
R21200 vdd.n205 vdd.n202 7.3702
R21201 vdd.n146 vdd.n143 7.3702
R21202 vdd.n104 vdd.n101 7.3702
R21203 vdd.n45 vdd.n42 7.3702
R21204 vdd.n1726 vdd.n1723 7.3702
R21205 vdd.n1785 vdd.n1782 7.3702
R21206 vdd.n1624 vdd.n1621 7.3702
R21207 vdd.n1683 vdd.n1680 7.3702
R21208 vdd.n1523 vdd.n1520 7.3702
R21209 vdd.n1582 vdd.n1579 7.3702
R21210 vdd.n1884 vdd.t17 7.1425
R21211 vdd.n679 vdd.t13 7.1425
R21212 vdd.n1358 vdd.n1357 6.98232
R21213 vdd.n2039 vdd.n2038 6.98232
R21214 vdd.n566 vdd.n565 6.98232
R21215 vdd.n3141 vdd.n3138 6.98232
R21216 vdd.t126 vdd.n1097 6.91577
R21217 vdd.n3264 vdd.t23 6.91577
R21218 vdd.n1843 vdd.t86 6.68904
R21219 vdd.n3280 vdd.t11 6.68904
R21220 vdd.t29 vdd.n1126 6.46231
R21221 vdd.n3308 vdd.t25 6.46231
R21222 vdd.n3400 vdd.n333 6.38151
R21223 vdd.n1812 vdd.n1811 6.38151
R21224 vdd.n1494 vdd.t57 6.23558
R21225 vdd.t97 vdd.n344 6.23558
R21226 vdd.t27 vdd.n1154 6.00885
R21227 vdd.n2412 vdd.t6 6.00885
R21228 vdd.n2912 vdd.t199 6.00885
R21229 vdd.n3379 vdd.t42 6.00885
R21230 vdd.n1033 vdd.t264 5.89549
R21231 vdd.t222 vdd.n851 5.89549
R21232 vdd.n308 vdd.n307 5.81868
R21233 vdd.n249 vdd.n248 5.81868
R21234 vdd.n206 vdd.n205 5.81868
R21235 vdd.n147 vdd.n146 5.81868
R21236 vdd.n105 vdd.n104 5.81868
R21237 vdd.n46 vdd.n45 5.81868
R21238 vdd.n1727 vdd.n1726 5.81868
R21239 vdd.n1786 vdd.n1785 5.81868
R21240 vdd.n1625 vdd.n1624 5.81868
R21241 vdd.n1684 vdd.n1683 5.81868
R21242 vdd.n1524 vdd.n1523 5.81868
R21243 vdd.n1583 vdd.n1582 5.81868
R21244 vdd.n1453 vdd.t15 5.78212
R21245 vdd.t207 vdd.n1037 5.78212
R21246 vdd.n2156 vdd.t246 5.78212
R21247 vdd.n2781 vdd.t254 5.78212
R21248 vdd.n846 vdd.t250 5.78212
R21249 vdd.n3370 vdd.t91 5.78212
R21250 vdd.n2540 vdd.n2539 5.77611
R21251 vdd.n2283 vdd.n2153 5.77611
R21252 vdd.n2794 vdd.n2793 5.77611
R21253 vdd.n3000 vdd.n2999 5.77611
R21254 vdd.n3064 vdd.n801 5.77611
R21255 vdd.n2704 vdd.n2644 5.77611
R21256 vdd.n2465 vdd.n967 5.77611
R21257 vdd.n2213 vdd.n2212 5.77611
R21258 vdd.n1320 vdd.n1319 5.62474
R21259 vdd.n2335 vdd.n2332 5.62474
R21260 vdd.n3351 vdd.n428 5.62474
R21261 vdd.n3225 vdd.n690 5.62474
R21262 vdd.n1177 vdd.t15 5.55539
R21263 vdd.t91 vdd.n3369 5.55539
R21264 vdd.t179 vdd.n989 5.44203
R21265 vdd.n893 vdd.t7 5.44203
R21266 vdd.n1469 vdd.t27 5.32866
R21267 vdd.t42 vdd.n3378 5.32866
R21268 vdd.n1485 vdd.t57 5.10193
R21269 vdd.t205 vdd.n1012 5.10193
R21270 vdd.n1002 vdd.t0 5.10193
R21271 vdd.t171 vdd.n880 5.10193
R21272 vdd.n870 vdd.t1 5.10193
R21273 vdd.n3387 vdd.t97 5.10193
R21274 vdd.n311 vdd.n302 5.04292
R21275 vdd.n252 vdd.n243 5.04292
R21276 vdd.n209 vdd.n200 5.04292
R21277 vdd.n150 vdd.n141 5.04292
R21278 vdd.n108 vdd.n99 5.04292
R21279 vdd.n49 vdd.n40 5.04292
R21280 vdd.n1730 vdd.n1721 5.04292
R21281 vdd.n1789 vdd.n1780 5.04292
R21282 vdd.n1628 vdd.n1619 5.04292
R21283 vdd.n1687 vdd.n1678 5.04292
R21284 vdd.n1527 vdd.n1518 5.04292
R21285 vdd.n1586 vdd.n1577 5.04292
R21286 vdd.n1817 vdd.t29 4.8752
R21287 vdd.t3 vdd.t282 4.8752
R21288 vdd.t178 vdd.t174 4.8752
R21289 vdd.t9 vdd.t177 4.8752
R21290 vdd.t290 vdd.t204 4.8752
R21291 vdd.t25 vdd.n340 4.8752
R21292 vdd.n2541 vdd.n2540 4.83952
R21293 vdd.n2153 vdd.n2149 4.83952
R21294 vdd.n2795 vdd.n2794 4.83952
R21295 vdd.n3001 vdd.n3000 4.83952
R21296 vdd.n801 vdd.n796 4.83952
R21297 vdd.n2701 vdd.n2644 4.83952
R21298 vdd.n2468 vdd.n967 4.83952
R21299 vdd.n2212 vdd.n2211 4.83952
R21300 vdd.n2007 vdd.n1065 4.74817
R21301 vdd.n2002 vdd.n1066 4.74817
R21302 vdd.n1904 vdd.n1901 4.74817
R21303 vdd.n2316 vdd.n1905 4.74817
R21304 vdd.n2318 vdd.n1904 4.74817
R21305 vdd.n2317 vdd.n2316 4.74817
R21306 vdd.n3218 vdd.n3217 4.74817
R21307 vdd.n3215 vdd.n3214 4.74817
R21308 vdd.n3215 vdd.n732 4.74817
R21309 vdd.n3217 vdd.n729 4.74817
R21310 vdd.n3100 vdd.n784 4.74817
R21311 vdd.n3096 vdd.n3094 4.74817
R21312 vdd.n3099 vdd.n3094 4.74817
R21313 vdd.n3103 vdd.n784 4.74817
R21314 vdd.n2003 vdd.n1065 4.74817
R21315 vdd.n1068 vdd.n1066 4.74817
R21316 vdd.n333 vdd.n332 4.7074
R21317 vdd.n231 vdd.n230 4.7074
R21318 vdd.n1811 vdd.n1810 4.7074
R21319 vdd.n1709 vdd.n1708 4.7074
R21320 vdd.n1120 vdd.t86 4.64847
R21321 vdd.n3289 vdd.t11 4.64847
R21322 vdd.n2418 vdd.t202 4.53511
R21323 vdd.n2906 vdd.t284 4.53511
R21324 vdd.n1859 vdd.t126 4.42174
R21325 vdd.t23 vdd.n655 4.42174
R21326 vdd.n2450 vdd.t288 4.30838
R21327 vdd.n2876 vdd.t200 4.30838
R21328 vdd.n312 vdd.n300 4.26717
R21329 vdd.n253 vdd.n241 4.26717
R21330 vdd.n210 vdd.n198 4.26717
R21331 vdd.n151 vdd.n139 4.26717
R21332 vdd.n109 vdd.n97 4.26717
R21333 vdd.n50 vdd.n38 4.26717
R21334 vdd.n1731 vdd.n1719 4.26717
R21335 vdd.n1790 vdd.n1778 4.26717
R21336 vdd.n1629 vdd.n1617 4.26717
R21337 vdd.n1688 vdd.n1676 4.26717
R21338 vdd.n1528 vdd.n1516 4.26717
R21339 vdd.n1587 vdd.n1575 4.26717
R21340 vdd.n1875 vdd.t17 4.19501
R21341 vdd.n3248 vdd.t13 4.19501
R21342 vdd.n333 vdd.n231 4.10845
R21343 vdd.n1811 vdd.n1709 4.10845
R21344 vdd.n289 vdd.t52 4.06363
R21345 vdd.n289 vdd.t113 4.06363
R21346 vdd.n287 vdd.t145 4.06363
R21347 vdd.n287 vdd.t162 4.06363
R21348 vdd.n285 vdd.t166 4.06363
R21349 vdd.n285 vdd.t59 4.06363
R21350 vdd.n283 vdd.t84 4.06363
R21351 vdd.n283 vdd.t165 4.06363
R21352 vdd.n281 vdd.t167 4.06363
R21353 vdd.n281 vdd.t83 4.06363
R21354 vdd.n279 vdd.t88 4.06363
R21355 vdd.n279 vdd.t90 4.06363
R21356 vdd.n277 vdd.t140 4.06363
R21357 vdd.n277 vdd.t41 4.06363
R21358 vdd.n275 vdd.t48 4.06363
R21359 vdd.n275 vdd.t112 4.06363
R21360 vdd.n273 vdd.t116 4.06363
R21361 vdd.n273 vdd.t147 4.06363
R21362 vdd.n187 vdd.t34 4.06363
R21363 vdd.n187 vdd.t92 4.06363
R21364 vdd.n185 vdd.t131 4.06363
R21365 vdd.n185 vdd.t150 4.06363
R21366 vdd.n183 vdd.t154 4.06363
R21367 vdd.n183 vdd.t36 4.06363
R21368 vdd.n181 vdd.t67 4.06363
R21369 vdd.n181 vdd.t153 4.06363
R21370 vdd.n179 vdd.t157 4.06363
R21371 vdd.n179 vdd.t66 4.06363
R21372 vdd.n177 vdd.t71 4.06363
R21373 vdd.n177 vdd.t73 4.06363
R21374 vdd.n175 vdd.t130 4.06363
R21375 vdd.n175 vdd.t12 4.06363
R21376 vdd.n173 vdd.t24 4.06363
R21377 vdd.n173 vdd.t93 4.06363
R21378 vdd.n171 vdd.t103 4.06363
R21379 vdd.n171 vdd.t132 4.06363
R21380 vdd.n86 vdd.t51 4.06363
R21381 vdd.n86 vdd.t138 4.06363
R21382 vdd.n84 vdd.t43 4.06363
R21383 vdd.n84 vdd.t122 4.06363
R21384 vdd.n82 vdd.t69 4.06363
R21385 vdd.n82 vdd.t151 4.06363
R21386 vdd.n80 vdd.t38 4.06363
R21387 vdd.n80 vdd.t98 4.06363
R21388 vdd.n78 vdd.t26 4.06363
R21389 vdd.n78 vdd.t74 4.06363
R21390 vdd.n76 vdd.t163 4.06363
R21391 vdd.n76 vdd.t137 4.06363
R21392 vdd.n74 vdd.t143 4.06363
R21393 vdd.n74 vdd.t85 4.06363
R21394 vdd.n72 vdd.t168 4.06363
R21395 vdd.n72 vdd.t61 4.06363
R21396 vdd.n70 vdd.t155 4.06363
R21397 vdd.n70 vdd.t95 4.06363
R21398 vdd.n1751 vdd.t50 4.06363
R21399 vdd.n1751 vdd.t161 4.06363
R21400 vdd.n1753 vdd.t158 4.06363
R21401 vdd.n1753 vdd.t139 4.06363
R21402 vdd.n1755 vdd.t108 4.06363
R21403 vdd.n1755 vdd.t46 4.06363
R21404 vdd.n1757 vdd.t170 4.06363
R21405 vdd.n1757 vdd.t136 4.06363
R21406 vdd.n1759 vdd.t133 4.06363
R21407 vdd.n1759 vdd.t82 4.06363
R21408 vdd.n1761 vdd.t78 4.06363
R21409 vdd.n1761 vdd.t134 4.06363
R21410 vdd.n1763 vdd.t118 4.06363
R21411 vdd.n1763 vdd.t117 4.06363
R21412 vdd.n1765 vdd.t75 4.06363
R21413 vdd.n1765 vdd.t49 4.06363
R21414 vdd.n1767 vdd.t45 4.06363
R21415 vdd.n1767 vdd.t114 4.06363
R21416 vdd.n1649 vdd.t32 4.06363
R21417 vdd.n1649 vdd.t149 4.06363
R21418 vdd.n1651 vdd.t142 4.06363
R21419 vdd.n1651 vdd.t127 4.06363
R21420 vdd.n1653 vdd.t89 4.06363
R21421 vdd.n1653 vdd.t20 4.06363
R21422 vdd.n1655 vdd.t159 4.06363
R21423 vdd.n1655 vdd.t125 4.06363
R21424 vdd.n1657 vdd.t119 4.06363
R21425 vdd.n1657 vdd.t64 4.06363
R21426 vdd.n1659 vdd.t58 4.06363
R21427 vdd.n1659 vdd.t120 4.06363
R21428 vdd.n1661 vdd.t107 4.06363
R21429 vdd.n1661 vdd.t105 4.06363
R21430 vdd.n1663 vdd.t54 4.06363
R21431 vdd.n1663 vdd.t28 4.06363
R21432 vdd.n1665 vdd.t16 4.06363
R21433 vdd.n1665 vdd.t100 4.06363
R21434 vdd.n1548 vdd.t96 4.06363
R21435 vdd.n1548 vdd.t156 4.06363
R21436 vdd.n1550 vdd.t63 4.06363
R21437 vdd.n1550 vdd.t135 4.06363
R21438 vdd.n1552 vdd.t87 4.06363
R21439 vdd.n1552 vdd.t144 4.06363
R21440 vdd.n1554 vdd.t110 4.06363
R21441 vdd.n1554 vdd.t164 4.06363
R21442 vdd.n1556 vdd.t77 4.06363
R21443 vdd.n1556 vdd.t30 4.06363
R21444 vdd.n1558 vdd.t99 4.06363
R21445 vdd.n1558 vdd.t40 4.06363
R21446 vdd.n1560 vdd.t152 4.06363
R21447 vdd.n1560 vdd.t169 4.06363
R21448 vdd.n1562 vdd.t123 4.06363
R21449 vdd.n1562 vdd.t44 4.06363
R21450 vdd.n1564 vdd.t111 4.06363
R21451 vdd.n1564 vdd.t56 4.06363
R21452 vdd.n26 vdd.t193 3.9605
R21453 vdd.n26 vdd.t188 3.9605
R21454 vdd.n23 vdd.t183 3.9605
R21455 vdd.n23 vdd.t184 3.9605
R21456 vdd.n21 vdd.t186 3.9605
R21457 vdd.n21 vdd.t191 3.9605
R21458 vdd.n20 vdd.t185 3.9605
R21459 vdd.n20 vdd.t189 3.9605
R21460 vdd.n15 vdd.t198 3.9605
R21461 vdd.n15 vdd.t197 3.9605
R21462 vdd.n16 vdd.t194 3.9605
R21463 vdd.n16 vdd.t187 3.9605
R21464 vdd.n18 vdd.t190 3.9605
R21465 vdd.n18 vdd.t196 3.9605
R21466 vdd.n25 vdd.t192 3.9605
R21467 vdd.n25 vdd.t195 3.9605
R21468 vdd.n7 vdd.t291 3.61217
R21469 vdd.n7 vdd.t285 3.61217
R21470 vdd.n8 vdd.t10 3.61217
R21471 vdd.n8 vdd.t8 3.61217
R21472 vdd.n10 vdd.t5 3.61217
R21473 vdd.n10 vdd.t201 3.61217
R21474 vdd.n12 vdd.t293 3.61217
R21475 vdd.n12 vdd.t287 3.61217
R21476 vdd.n5 vdd.t295 3.61217
R21477 vdd.n5 vdd.t182 3.61217
R21478 vdd.n3 vdd.t289 3.61217
R21479 vdd.n3 vdd.t173 3.61217
R21480 vdd.n1 vdd.t180 3.61217
R21481 vdd.n1 vdd.t175 3.61217
R21482 vdd.n0 vdd.t203 3.61217
R21483 vdd.n0 vdd.t283 3.61217
R21484 vdd.n316 vdd.n315 3.49141
R21485 vdd.n257 vdd.n256 3.49141
R21486 vdd.n214 vdd.n213 3.49141
R21487 vdd.n155 vdd.n154 3.49141
R21488 vdd.n113 vdd.n112 3.49141
R21489 vdd.n54 vdd.n53 3.49141
R21490 vdd.n1735 vdd.n1734 3.49141
R21491 vdd.n1794 vdd.n1793 3.49141
R21492 vdd.n1633 vdd.n1632 3.49141
R21493 vdd.n1692 vdd.n1691 3.49141
R21494 vdd.n1532 vdd.n1531 3.49141
R21495 vdd.n1591 vdd.n1590 3.49141
R21496 vdd.n2156 vdd.t288 3.40145
R21497 vdd.n2604 vdd.t294 3.40145
R21498 vdd.n2857 vdd.t286 3.40145
R21499 vdd.n2781 vdd.t200 3.40145
R21500 vdd.n1876 vdd.t148 3.28809
R21501 vdd.n3247 vdd.t102 3.28809
R21502 vdd.n2257 vdd.t202 3.17472
R21503 vdd.n2760 vdd.t284 3.17472
R21504 vdd.t62 vdd.n1104 3.06136
R21505 vdd.n3272 vdd.t60 3.06136
R21506 vdd.n1834 vdd.t124 2.83463
R21507 vdd.n644 vdd.t70 2.83463
R21508 vdd.n319 vdd.n298 2.71565
R21509 vdd.n260 vdd.n239 2.71565
R21510 vdd.n217 vdd.n196 2.71565
R21511 vdd.n158 vdd.n137 2.71565
R21512 vdd.n116 vdd.n95 2.71565
R21513 vdd.n57 vdd.n36 2.71565
R21514 vdd.n1738 vdd.n1717 2.71565
R21515 vdd.n1797 vdd.n1776 2.71565
R21516 vdd.n1636 vdd.n1615 2.71565
R21517 vdd.n1695 vdd.n1674 2.71565
R21518 vdd.n1535 vdd.n1514 2.71565
R21519 vdd.n1594 vdd.n1573 2.71565
R21520 vdd.t76 vdd.n1132 2.6079
R21521 vdd.n2406 vdd.t205 2.6079
R21522 vdd.n2430 vdd.t0 2.6079
R21523 vdd.n2894 vdd.t171 2.6079
R21524 vdd.n2918 vdd.t1 2.6079
R21525 vdd.n3395 vdd.t65 2.6079
R21526 vdd.n2924 vdd.n2923 2.49806
R21527 vdd.n2398 vdd.n2397 2.49806
R21528 vdd.n306 vdd.n305 2.4129
R21529 vdd.n247 vdd.n246 2.4129
R21530 vdd.n204 vdd.n203 2.4129
R21531 vdd.n145 vdd.n144 2.4129
R21532 vdd.n103 vdd.n102 2.4129
R21533 vdd.n44 vdd.n43 2.4129
R21534 vdd.n1725 vdd.n1724 2.4129
R21535 vdd.n1784 vdd.n1783 2.4129
R21536 vdd.n1623 vdd.n1622 2.4129
R21537 vdd.n1682 vdd.n1681 2.4129
R21538 vdd.n1522 vdd.n1521 2.4129
R21539 vdd.n1581 vdd.n1580 2.4129
R21540 vdd.n1486 vdd.t104 2.38117
R21541 vdd.n1894 vdd.t218 2.38117
R21542 vdd.n3231 vdd.t211 2.38117
R21543 vdd.n3386 vdd.t68 2.38117
R21544 vdd.n2315 vdd.n1904 2.27742
R21545 vdd.n2316 vdd.n2315 2.27742
R21546 vdd.n3216 vdd.n3215 2.27742
R21547 vdd.n3217 vdd.n3216 2.27742
R21548 vdd.n3094 vdd.n3093 2.27742
R21549 vdd.n3093 vdd.n784 2.27742
R21550 vdd.n2338 vdd.n1065 2.27742
R21551 vdd.n2338 vdd.n1066 2.27742
R21552 vdd.n2430 vdd.t179 2.2678
R21553 vdd.n2894 vdd.t7 2.2678
R21554 vdd.t53 vdd.n1161 2.15444
R21555 vdd.n3377 vdd.t121 2.15444
R21556 vdd.t174 vdd.n983 2.04107
R21557 vdd.n900 vdd.t9 2.04107
R21558 vdd.n320 vdd.n296 1.93989
R21559 vdd.n261 vdd.n237 1.93989
R21560 vdd.n218 vdd.n194 1.93989
R21561 vdd.n159 vdd.n135 1.93989
R21562 vdd.n117 vdd.n93 1.93989
R21563 vdd.n58 vdd.n34 1.93989
R21564 vdd.n1739 vdd.n1715 1.93989
R21565 vdd.n1798 vdd.n1774 1.93989
R21566 vdd.n1637 vdd.n1613 1.93989
R21567 vdd.n1696 vdd.n1672 1.93989
R21568 vdd.n1536 vdd.n1512 1.93989
R21569 vdd.n1595 vdd.n1571 1.93989
R21570 vdd.n1444 vdd.t21 1.92771
R21571 vdd.n2381 vdd.t207 1.92771
R21572 vdd.n2457 vdd.t246 1.92771
R21573 vdd.n2870 vdd.t254 1.92771
R21574 vdd.n2989 vdd.t250 1.92771
R21575 vdd.t79 vdd.n375 1.92771
R21576 vdd.n1452 vdd.t55 1.70098
R21577 vdd.n2257 vdd.t6 1.70098
R21578 vdd.n1008 vdd.t3 1.70098
R21579 vdd.t204 vdd.n874 1.70098
R21580 vdd.n2760 vdd.t199 1.70098
R21581 vdd.n3371 vdd.t33 1.70098
R21582 vdd.n1477 vdd.t106 1.47425
R21583 vdd.n361 vdd.t35 1.47425
R21584 vdd.n1143 vdd.t39 1.24752
R21585 vdd.t37 vdd.n3393 1.24752
R21586 vdd.n331 vdd.n291 1.16414
R21587 vdd.n324 vdd.n323 1.16414
R21588 vdd.n272 vdd.n232 1.16414
R21589 vdd.n265 vdd.n264 1.16414
R21590 vdd.n229 vdd.n189 1.16414
R21591 vdd.n222 vdd.n221 1.16414
R21592 vdd.n170 vdd.n130 1.16414
R21593 vdd.n163 vdd.n162 1.16414
R21594 vdd.n128 vdd.n88 1.16414
R21595 vdd.n121 vdd.n120 1.16414
R21596 vdd.n69 vdd.n29 1.16414
R21597 vdd.n62 vdd.n61 1.16414
R21598 vdd.n1750 vdd.n1710 1.16414
R21599 vdd.n1743 vdd.n1742 1.16414
R21600 vdd.n1809 vdd.n1769 1.16414
R21601 vdd.n1802 vdd.n1801 1.16414
R21602 vdd.n1648 vdd.n1608 1.16414
R21603 vdd.n1641 vdd.n1640 1.16414
R21604 vdd.n1707 vdd.n1667 1.16414
R21605 vdd.n1700 vdd.n1699 1.16414
R21606 vdd.n1547 vdd.n1507 1.16414
R21607 vdd.n1540 vdd.n1539 1.16414
R21608 vdd.n1606 vdd.n1566 1.16414
R21609 vdd.n1599 vdd.n1598 1.16414
R21610 vdd.n2424 vdd.t282 1.13415
R21611 vdd.n2900 vdd.t290 1.13415
R21612 vdd.n1826 vdd.t109 1.02079
R21613 vdd.t264 vdd.t2 1.02079
R21614 vdd.t176 vdd.t222 1.02079
R21615 vdd.t72 vdd.n633 1.02079
R21616 vdd.n1323 vdd.n1319 0.970197
R21617 vdd.n2336 vdd.n2335 0.970197
R21618 vdd.n618 vdd.n428 0.970197
R21619 vdd.n3095 vdd.n690 0.970197
R21620 vdd.n1812 vdd.n28 0.90431
R21621 vdd vdd.n3400 0.896477
R21622 vdd.n1842 vdd.t19 0.794056
R21623 vdd.n2400 vdd.t2 0.794056
R21624 vdd.n2436 vdd.t178 0.794056
R21625 vdd.n2888 vdd.t177 0.794056
R21626 vdd.n2926 vdd.t176 0.794056
R21627 vdd.n3281 vdd.t129 0.794056
R21628 vdd.n1867 vdd.t31 0.567326
R21629 vdd.t94 vdd.n662 0.567326
R21630 vdd.n2326 vdd.n2325 0.530988
R21631 vdd.n726 vdd.n682 0.530988
R21632 vdd.n464 vdd.n391 0.530988
R21633 vdd.n3350 vdd.n3349 0.530988
R21634 vdd.n3227 vdd.n3226 0.530988
R21635 vdd.n1889 vdd.n1067 0.530988
R21636 vdd.n1321 vdd.n1186 0.530988
R21637 vdd.n1423 vdd.n1422 0.530988
R21638 vdd.n4 vdd.n2 0.459552
R21639 vdd.n11 vdd.n9 0.459552
R21640 vdd.n329 vdd.n328 0.388379
R21641 vdd.n295 vdd.n293 0.388379
R21642 vdd.n270 vdd.n269 0.388379
R21643 vdd.n236 vdd.n234 0.388379
R21644 vdd.n227 vdd.n226 0.388379
R21645 vdd.n193 vdd.n191 0.388379
R21646 vdd.n168 vdd.n167 0.388379
R21647 vdd.n134 vdd.n132 0.388379
R21648 vdd.n126 vdd.n125 0.388379
R21649 vdd.n92 vdd.n90 0.388379
R21650 vdd.n67 vdd.n66 0.388379
R21651 vdd.n33 vdd.n31 0.388379
R21652 vdd.n1748 vdd.n1747 0.388379
R21653 vdd.n1714 vdd.n1712 0.388379
R21654 vdd.n1807 vdd.n1806 0.388379
R21655 vdd.n1773 vdd.n1771 0.388379
R21656 vdd.n1646 vdd.n1645 0.388379
R21657 vdd.n1612 vdd.n1610 0.388379
R21658 vdd.n1705 vdd.n1704 0.388379
R21659 vdd.n1671 vdd.n1669 0.388379
R21660 vdd.n1545 vdd.n1544 0.388379
R21661 vdd.n1511 vdd.n1509 0.388379
R21662 vdd.n1604 vdd.n1603 0.388379
R21663 vdd.n1570 vdd.n1568 0.388379
R21664 vdd.n19 vdd.n17 0.387128
R21665 vdd.n24 vdd.n22 0.387128
R21666 vdd.n6 vdd.n4 0.358259
R21667 vdd.n13 vdd.n11 0.358259
R21668 vdd.n276 vdd.n274 0.358259
R21669 vdd.n278 vdd.n276 0.358259
R21670 vdd.n280 vdd.n278 0.358259
R21671 vdd.n282 vdd.n280 0.358259
R21672 vdd.n284 vdd.n282 0.358259
R21673 vdd.n286 vdd.n284 0.358259
R21674 vdd.n288 vdd.n286 0.358259
R21675 vdd.n290 vdd.n288 0.358259
R21676 vdd.n332 vdd.n290 0.358259
R21677 vdd.n174 vdd.n172 0.358259
R21678 vdd.n176 vdd.n174 0.358259
R21679 vdd.n178 vdd.n176 0.358259
R21680 vdd.n180 vdd.n178 0.358259
R21681 vdd.n182 vdd.n180 0.358259
R21682 vdd.n184 vdd.n182 0.358259
R21683 vdd.n186 vdd.n184 0.358259
R21684 vdd.n188 vdd.n186 0.358259
R21685 vdd.n230 vdd.n188 0.358259
R21686 vdd.n73 vdd.n71 0.358259
R21687 vdd.n75 vdd.n73 0.358259
R21688 vdd.n77 vdd.n75 0.358259
R21689 vdd.n79 vdd.n77 0.358259
R21690 vdd.n81 vdd.n79 0.358259
R21691 vdd.n83 vdd.n81 0.358259
R21692 vdd.n85 vdd.n83 0.358259
R21693 vdd.n87 vdd.n85 0.358259
R21694 vdd.n129 vdd.n87 0.358259
R21695 vdd.n1810 vdd.n1768 0.358259
R21696 vdd.n1768 vdd.n1766 0.358259
R21697 vdd.n1766 vdd.n1764 0.358259
R21698 vdd.n1764 vdd.n1762 0.358259
R21699 vdd.n1762 vdd.n1760 0.358259
R21700 vdd.n1760 vdd.n1758 0.358259
R21701 vdd.n1758 vdd.n1756 0.358259
R21702 vdd.n1756 vdd.n1754 0.358259
R21703 vdd.n1754 vdd.n1752 0.358259
R21704 vdd.n1708 vdd.n1666 0.358259
R21705 vdd.n1666 vdd.n1664 0.358259
R21706 vdd.n1664 vdd.n1662 0.358259
R21707 vdd.n1662 vdd.n1660 0.358259
R21708 vdd.n1660 vdd.n1658 0.358259
R21709 vdd.n1658 vdd.n1656 0.358259
R21710 vdd.n1656 vdd.n1654 0.358259
R21711 vdd.n1654 vdd.n1652 0.358259
R21712 vdd.n1652 vdd.n1650 0.358259
R21713 vdd.n1607 vdd.n1565 0.358259
R21714 vdd.n1565 vdd.n1563 0.358259
R21715 vdd.n1563 vdd.n1561 0.358259
R21716 vdd.n1561 vdd.n1559 0.358259
R21717 vdd.n1559 vdd.n1557 0.358259
R21718 vdd.n1557 vdd.n1555 0.358259
R21719 vdd.n1555 vdd.n1553 0.358259
R21720 vdd.n1553 vdd.n1551 0.358259
R21721 vdd.n1551 vdd.n1549 0.358259
R21722 vdd.n14 vdd.n6 0.334552
R21723 vdd.n14 vdd.n13 0.334552
R21724 vdd.n27 vdd.n19 0.21707
R21725 vdd.n27 vdd.n24 0.21707
R21726 vdd.n330 vdd.n292 0.155672
R21727 vdd.n322 vdd.n292 0.155672
R21728 vdd.n322 vdd.n321 0.155672
R21729 vdd.n321 vdd.n297 0.155672
R21730 vdd.n314 vdd.n297 0.155672
R21731 vdd.n314 vdd.n313 0.155672
R21732 vdd.n313 vdd.n301 0.155672
R21733 vdd.n306 vdd.n301 0.155672
R21734 vdd.n271 vdd.n233 0.155672
R21735 vdd.n263 vdd.n233 0.155672
R21736 vdd.n263 vdd.n262 0.155672
R21737 vdd.n262 vdd.n238 0.155672
R21738 vdd.n255 vdd.n238 0.155672
R21739 vdd.n255 vdd.n254 0.155672
R21740 vdd.n254 vdd.n242 0.155672
R21741 vdd.n247 vdd.n242 0.155672
R21742 vdd.n228 vdd.n190 0.155672
R21743 vdd.n220 vdd.n190 0.155672
R21744 vdd.n220 vdd.n219 0.155672
R21745 vdd.n219 vdd.n195 0.155672
R21746 vdd.n212 vdd.n195 0.155672
R21747 vdd.n212 vdd.n211 0.155672
R21748 vdd.n211 vdd.n199 0.155672
R21749 vdd.n204 vdd.n199 0.155672
R21750 vdd.n169 vdd.n131 0.155672
R21751 vdd.n161 vdd.n131 0.155672
R21752 vdd.n161 vdd.n160 0.155672
R21753 vdd.n160 vdd.n136 0.155672
R21754 vdd.n153 vdd.n136 0.155672
R21755 vdd.n153 vdd.n152 0.155672
R21756 vdd.n152 vdd.n140 0.155672
R21757 vdd.n145 vdd.n140 0.155672
R21758 vdd.n127 vdd.n89 0.155672
R21759 vdd.n119 vdd.n89 0.155672
R21760 vdd.n119 vdd.n118 0.155672
R21761 vdd.n118 vdd.n94 0.155672
R21762 vdd.n111 vdd.n94 0.155672
R21763 vdd.n111 vdd.n110 0.155672
R21764 vdd.n110 vdd.n98 0.155672
R21765 vdd.n103 vdd.n98 0.155672
R21766 vdd.n68 vdd.n30 0.155672
R21767 vdd.n60 vdd.n30 0.155672
R21768 vdd.n60 vdd.n59 0.155672
R21769 vdd.n59 vdd.n35 0.155672
R21770 vdd.n52 vdd.n35 0.155672
R21771 vdd.n52 vdd.n51 0.155672
R21772 vdd.n51 vdd.n39 0.155672
R21773 vdd.n44 vdd.n39 0.155672
R21774 vdd.n1749 vdd.n1711 0.155672
R21775 vdd.n1741 vdd.n1711 0.155672
R21776 vdd.n1741 vdd.n1740 0.155672
R21777 vdd.n1740 vdd.n1716 0.155672
R21778 vdd.n1733 vdd.n1716 0.155672
R21779 vdd.n1733 vdd.n1732 0.155672
R21780 vdd.n1732 vdd.n1720 0.155672
R21781 vdd.n1725 vdd.n1720 0.155672
R21782 vdd.n1808 vdd.n1770 0.155672
R21783 vdd.n1800 vdd.n1770 0.155672
R21784 vdd.n1800 vdd.n1799 0.155672
R21785 vdd.n1799 vdd.n1775 0.155672
R21786 vdd.n1792 vdd.n1775 0.155672
R21787 vdd.n1792 vdd.n1791 0.155672
R21788 vdd.n1791 vdd.n1779 0.155672
R21789 vdd.n1784 vdd.n1779 0.155672
R21790 vdd.n1647 vdd.n1609 0.155672
R21791 vdd.n1639 vdd.n1609 0.155672
R21792 vdd.n1639 vdd.n1638 0.155672
R21793 vdd.n1638 vdd.n1614 0.155672
R21794 vdd.n1631 vdd.n1614 0.155672
R21795 vdd.n1631 vdd.n1630 0.155672
R21796 vdd.n1630 vdd.n1618 0.155672
R21797 vdd.n1623 vdd.n1618 0.155672
R21798 vdd.n1706 vdd.n1668 0.155672
R21799 vdd.n1698 vdd.n1668 0.155672
R21800 vdd.n1698 vdd.n1697 0.155672
R21801 vdd.n1697 vdd.n1673 0.155672
R21802 vdd.n1690 vdd.n1673 0.155672
R21803 vdd.n1690 vdd.n1689 0.155672
R21804 vdd.n1689 vdd.n1677 0.155672
R21805 vdd.n1682 vdd.n1677 0.155672
R21806 vdd.n1546 vdd.n1508 0.155672
R21807 vdd.n1538 vdd.n1508 0.155672
R21808 vdd.n1538 vdd.n1537 0.155672
R21809 vdd.n1537 vdd.n1513 0.155672
R21810 vdd.n1530 vdd.n1513 0.155672
R21811 vdd.n1530 vdd.n1529 0.155672
R21812 vdd.n1529 vdd.n1517 0.155672
R21813 vdd.n1522 vdd.n1517 0.155672
R21814 vdd.n1605 vdd.n1567 0.155672
R21815 vdd.n1597 vdd.n1567 0.155672
R21816 vdd.n1597 vdd.n1596 0.155672
R21817 vdd.n1596 vdd.n1572 0.155672
R21818 vdd.n1589 vdd.n1572 0.155672
R21819 vdd.n1589 vdd.n1588 0.155672
R21820 vdd.n1588 vdd.n1576 0.155672
R21821 vdd.n1581 vdd.n1576 0.155672
R21822 vdd.n2101 vdd.n1906 0.152939
R21823 vdd.n1912 vdd.n1906 0.152939
R21824 vdd.n1913 vdd.n1912 0.152939
R21825 vdd.n1914 vdd.n1913 0.152939
R21826 vdd.n1915 vdd.n1914 0.152939
R21827 vdd.n1919 vdd.n1915 0.152939
R21828 vdd.n1920 vdd.n1919 0.152939
R21829 vdd.n1921 vdd.n1920 0.152939
R21830 vdd.n1922 vdd.n1921 0.152939
R21831 vdd.n1926 vdd.n1922 0.152939
R21832 vdd.n1927 vdd.n1926 0.152939
R21833 vdd.n1928 vdd.n1927 0.152939
R21834 vdd.n2076 vdd.n1928 0.152939
R21835 vdd.n2076 vdd.n2075 0.152939
R21836 vdd.n2075 vdd.n2074 0.152939
R21837 vdd.n2074 vdd.n1934 0.152939
R21838 vdd.n1939 vdd.n1934 0.152939
R21839 vdd.n1940 vdd.n1939 0.152939
R21840 vdd.n1941 vdd.n1940 0.152939
R21841 vdd.n1945 vdd.n1941 0.152939
R21842 vdd.n1946 vdd.n1945 0.152939
R21843 vdd.n1947 vdd.n1946 0.152939
R21844 vdd.n1948 vdd.n1947 0.152939
R21845 vdd.n1952 vdd.n1948 0.152939
R21846 vdd.n1953 vdd.n1952 0.152939
R21847 vdd.n1954 vdd.n1953 0.152939
R21848 vdd.n1955 vdd.n1954 0.152939
R21849 vdd.n1959 vdd.n1955 0.152939
R21850 vdd.n1960 vdd.n1959 0.152939
R21851 vdd.n1961 vdd.n1960 0.152939
R21852 vdd.n1962 vdd.n1961 0.152939
R21853 vdd.n1966 vdd.n1962 0.152939
R21854 vdd.n1967 vdd.n1966 0.152939
R21855 vdd.n1968 vdd.n1967 0.152939
R21856 vdd.n2037 vdd.n1968 0.152939
R21857 vdd.n2037 vdd.n2036 0.152939
R21858 vdd.n2036 vdd.n2035 0.152939
R21859 vdd.n2035 vdd.n1974 0.152939
R21860 vdd.n1979 vdd.n1974 0.152939
R21861 vdd.n1980 vdd.n1979 0.152939
R21862 vdd.n1981 vdd.n1980 0.152939
R21863 vdd.n1985 vdd.n1981 0.152939
R21864 vdd.n1986 vdd.n1985 0.152939
R21865 vdd.n1987 vdd.n1986 0.152939
R21866 vdd.n1988 vdd.n1987 0.152939
R21867 vdd.n1992 vdd.n1988 0.152939
R21868 vdd.n1993 vdd.n1992 0.152939
R21869 vdd.n1994 vdd.n1993 0.152939
R21870 vdd.n1995 vdd.n1994 0.152939
R21871 vdd.n1996 vdd.n1995 0.152939
R21872 vdd.n1996 vdd.n1064 0.152939
R21873 vdd.n2325 vdd.n1900 0.152939
R21874 vdd.n1814 vdd.n1123 0.152939
R21875 vdd.n1829 vdd.n1123 0.152939
R21876 vdd.n1830 vdd.n1829 0.152939
R21877 vdd.n1831 vdd.n1830 0.152939
R21878 vdd.n1831 vdd.n1112 0.152939
R21879 vdd.n1846 vdd.n1112 0.152939
R21880 vdd.n1847 vdd.n1846 0.152939
R21881 vdd.n1848 vdd.n1847 0.152939
R21882 vdd.n1848 vdd.n1101 0.152939
R21883 vdd.n1862 vdd.n1101 0.152939
R21884 vdd.n1863 vdd.n1862 0.152939
R21885 vdd.n1864 vdd.n1863 0.152939
R21886 vdd.n1864 vdd.n1089 0.152939
R21887 vdd.n1879 vdd.n1089 0.152939
R21888 vdd.n1880 vdd.n1879 0.152939
R21889 vdd.n1881 vdd.n1880 0.152939
R21890 vdd.n1881 vdd.n1077 0.152939
R21891 vdd.n1898 vdd.n1077 0.152939
R21892 vdd.n1899 vdd.n1898 0.152939
R21893 vdd.n2326 vdd.n1899 0.152939
R21894 vdd.n735 vdd.n730 0.152939
R21895 vdd.n736 vdd.n735 0.152939
R21896 vdd.n737 vdd.n736 0.152939
R21897 vdd.n738 vdd.n737 0.152939
R21898 vdd.n739 vdd.n738 0.152939
R21899 vdd.n740 vdd.n739 0.152939
R21900 vdd.n741 vdd.n740 0.152939
R21901 vdd.n742 vdd.n741 0.152939
R21902 vdd.n743 vdd.n742 0.152939
R21903 vdd.n744 vdd.n743 0.152939
R21904 vdd.n745 vdd.n744 0.152939
R21905 vdd.n746 vdd.n745 0.152939
R21906 vdd.n3183 vdd.n746 0.152939
R21907 vdd.n3183 vdd.n3182 0.152939
R21908 vdd.n3182 vdd.n3181 0.152939
R21909 vdd.n3181 vdd.n748 0.152939
R21910 vdd.n749 vdd.n748 0.152939
R21911 vdd.n750 vdd.n749 0.152939
R21912 vdd.n751 vdd.n750 0.152939
R21913 vdd.n752 vdd.n751 0.152939
R21914 vdd.n753 vdd.n752 0.152939
R21915 vdd.n754 vdd.n753 0.152939
R21916 vdd.n755 vdd.n754 0.152939
R21917 vdd.n756 vdd.n755 0.152939
R21918 vdd.n757 vdd.n756 0.152939
R21919 vdd.n758 vdd.n757 0.152939
R21920 vdd.n759 vdd.n758 0.152939
R21921 vdd.n760 vdd.n759 0.152939
R21922 vdd.n761 vdd.n760 0.152939
R21923 vdd.n762 vdd.n761 0.152939
R21924 vdd.n763 vdd.n762 0.152939
R21925 vdd.n764 vdd.n763 0.152939
R21926 vdd.n765 vdd.n764 0.152939
R21927 vdd.n766 vdd.n765 0.152939
R21928 vdd.n3137 vdd.n766 0.152939
R21929 vdd.n3137 vdd.n3136 0.152939
R21930 vdd.n3136 vdd.n3135 0.152939
R21931 vdd.n3135 vdd.n770 0.152939
R21932 vdd.n771 vdd.n770 0.152939
R21933 vdd.n772 vdd.n771 0.152939
R21934 vdd.n773 vdd.n772 0.152939
R21935 vdd.n774 vdd.n773 0.152939
R21936 vdd.n775 vdd.n774 0.152939
R21937 vdd.n776 vdd.n775 0.152939
R21938 vdd.n777 vdd.n776 0.152939
R21939 vdd.n778 vdd.n777 0.152939
R21940 vdd.n779 vdd.n778 0.152939
R21941 vdd.n780 vdd.n779 0.152939
R21942 vdd.n781 vdd.n780 0.152939
R21943 vdd.n782 vdd.n781 0.152939
R21944 vdd.n783 vdd.n782 0.152939
R21945 vdd.n727 vdd.n726 0.152939
R21946 vdd.n3234 vdd.n682 0.152939
R21947 vdd.n3235 vdd.n3234 0.152939
R21948 vdd.n3236 vdd.n3235 0.152939
R21949 vdd.n3236 vdd.n670 0.152939
R21950 vdd.n3251 vdd.n670 0.152939
R21951 vdd.n3252 vdd.n3251 0.152939
R21952 vdd.n3253 vdd.n3252 0.152939
R21953 vdd.n3253 vdd.n659 0.152939
R21954 vdd.n3267 vdd.n659 0.152939
R21955 vdd.n3268 vdd.n3267 0.152939
R21956 vdd.n3269 vdd.n3268 0.152939
R21957 vdd.n3269 vdd.n647 0.152939
R21958 vdd.n3284 vdd.n647 0.152939
R21959 vdd.n3285 vdd.n3284 0.152939
R21960 vdd.n3286 vdd.n3285 0.152939
R21961 vdd.n3286 vdd.n636 0.152939
R21962 vdd.n3303 vdd.n636 0.152939
R21963 vdd.n3304 vdd.n3303 0.152939
R21964 vdd.n3305 vdd.n3304 0.152939
R21965 vdd.n3305 vdd.n334 0.152939
R21966 vdd.n3398 vdd.n335 0.152939
R21967 vdd.n346 vdd.n335 0.152939
R21968 vdd.n347 vdd.n346 0.152939
R21969 vdd.n348 vdd.n347 0.152939
R21970 vdd.n355 vdd.n348 0.152939
R21971 vdd.n356 vdd.n355 0.152939
R21972 vdd.n357 vdd.n356 0.152939
R21973 vdd.n358 vdd.n357 0.152939
R21974 vdd.n366 vdd.n358 0.152939
R21975 vdd.n367 vdd.n366 0.152939
R21976 vdd.n368 vdd.n367 0.152939
R21977 vdd.n369 vdd.n368 0.152939
R21978 vdd.n377 vdd.n369 0.152939
R21979 vdd.n378 vdd.n377 0.152939
R21980 vdd.n379 vdd.n378 0.152939
R21981 vdd.n380 vdd.n379 0.152939
R21982 vdd.n388 vdd.n380 0.152939
R21983 vdd.n389 vdd.n388 0.152939
R21984 vdd.n390 vdd.n389 0.152939
R21985 vdd.n391 vdd.n390 0.152939
R21986 vdd.n464 vdd.n463 0.152939
R21987 vdd.n470 vdd.n463 0.152939
R21988 vdd.n471 vdd.n470 0.152939
R21989 vdd.n472 vdd.n471 0.152939
R21990 vdd.n472 vdd.n461 0.152939
R21991 vdd.n480 vdd.n461 0.152939
R21992 vdd.n481 vdd.n480 0.152939
R21993 vdd.n482 vdd.n481 0.152939
R21994 vdd.n482 vdd.n459 0.152939
R21995 vdd.n490 vdd.n459 0.152939
R21996 vdd.n491 vdd.n490 0.152939
R21997 vdd.n492 vdd.n491 0.152939
R21998 vdd.n492 vdd.n457 0.152939
R21999 vdd.n500 vdd.n457 0.152939
R22000 vdd.n501 vdd.n500 0.152939
R22001 vdd.n502 vdd.n501 0.152939
R22002 vdd.n502 vdd.n455 0.152939
R22003 vdd.n510 vdd.n455 0.152939
R22004 vdd.n511 vdd.n510 0.152939
R22005 vdd.n512 vdd.n511 0.152939
R22006 vdd.n512 vdd.n451 0.152939
R22007 vdd.n520 vdd.n451 0.152939
R22008 vdd.n521 vdd.n520 0.152939
R22009 vdd.n522 vdd.n521 0.152939
R22010 vdd.n522 vdd.n449 0.152939
R22011 vdd.n530 vdd.n449 0.152939
R22012 vdd.n531 vdd.n530 0.152939
R22013 vdd.n532 vdd.n531 0.152939
R22014 vdd.n532 vdd.n447 0.152939
R22015 vdd.n540 vdd.n447 0.152939
R22016 vdd.n541 vdd.n540 0.152939
R22017 vdd.n542 vdd.n541 0.152939
R22018 vdd.n542 vdd.n445 0.152939
R22019 vdd.n550 vdd.n445 0.152939
R22020 vdd.n551 vdd.n550 0.152939
R22021 vdd.n552 vdd.n551 0.152939
R22022 vdd.n552 vdd.n443 0.152939
R22023 vdd.n560 vdd.n443 0.152939
R22024 vdd.n561 vdd.n560 0.152939
R22025 vdd.n562 vdd.n561 0.152939
R22026 vdd.n562 vdd.n439 0.152939
R22027 vdd.n570 vdd.n439 0.152939
R22028 vdd.n571 vdd.n570 0.152939
R22029 vdd.n572 vdd.n571 0.152939
R22030 vdd.n572 vdd.n437 0.152939
R22031 vdd.n580 vdd.n437 0.152939
R22032 vdd.n581 vdd.n580 0.152939
R22033 vdd.n582 vdd.n581 0.152939
R22034 vdd.n582 vdd.n435 0.152939
R22035 vdd.n590 vdd.n435 0.152939
R22036 vdd.n591 vdd.n590 0.152939
R22037 vdd.n592 vdd.n591 0.152939
R22038 vdd.n592 vdd.n433 0.152939
R22039 vdd.n600 vdd.n433 0.152939
R22040 vdd.n601 vdd.n600 0.152939
R22041 vdd.n602 vdd.n601 0.152939
R22042 vdd.n602 vdd.n431 0.152939
R22043 vdd.n610 vdd.n431 0.152939
R22044 vdd.n611 vdd.n610 0.152939
R22045 vdd.n612 vdd.n611 0.152939
R22046 vdd.n612 vdd.n429 0.152939
R22047 vdd.n619 vdd.n429 0.152939
R22048 vdd.n3350 vdd.n619 0.152939
R22049 vdd.n3228 vdd.n3227 0.152939
R22050 vdd.n3228 vdd.n675 0.152939
R22051 vdd.n3242 vdd.n675 0.152939
R22052 vdd.n3243 vdd.n3242 0.152939
R22053 vdd.n3244 vdd.n3243 0.152939
R22054 vdd.n3244 vdd.n665 0.152939
R22055 vdd.n3259 vdd.n665 0.152939
R22056 vdd.n3260 vdd.n3259 0.152939
R22057 vdd.n3261 vdd.n3260 0.152939
R22058 vdd.n3261 vdd.n652 0.152939
R22059 vdd.n3275 vdd.n652 0.152939
R22060 vdd.n3276 vdd.n3275 0.152939
R22061 vdd.n3277 vdd.n3276 0.152939
R22062 vdd.n3277 vdd.n641 0.152939
R22063 vdd.n3292 vdd.n641 0.152939
R22064 vdd.n3293 vdd.n3292 0.152939
R22065 vdd.n3294 vdd.n3293 0.152939
R22066 vdd.n3296 vdd.n3294 0.152939
R22067 vdd.n3296 vdd.n3295 0.152939
R22068 vdd.n3295 vdd.n630 0.152939
R22069 vdd.n3313 vdd.n630 0.152939
R22070 vdd.n3314 vdd.n3313 0.152939
R22071 vdd.n3315 vdd.n3314 0.152939
R22072 vdd.n3315 vdd.n628 0.152939
R22073 vdd.n3320 vdd.n628 0.152939
R22074 vdd.n3321 vdd.n3320 0.152939
R22075 vdd.n3322 vdd.n3321 0.152939
R22076 vdd.n3322 vdd.n626 0.152939
R22077 vdd.n3327 vdd.n626 0.152939
R22078 vdd.n3328 vdd.n3327 0.152939
R22079 vdd.n3329 vdd.n3328 0.152939
R22080 vdd.n3329 vdd.n624 0.152939
R22081 vdd.n3335 vdd.n624 0.152939
R22082 vdd.n3336 vdd.n3335 0.152939
R22083 vdd.n3337 vdd.n3336 0.152939
R22084 vdd.n3337 vdd.n622 0.152939
R22085 vdd.n3342 vdd.n622 0.152939
R22086 vdd.n3343 vdd.n3342 0.152939
R22087 vdd.n3344 vdd.n3343 0.152939
R22088 vdd.n3344 vdd.n620 0.152939
R22089 vdd.n3349 vdd.n620 0.152939
R22090 vdd.n3226 vdd.n687 0.152939
R22091 vdd.n2337 vdd.n1067 0.152939
R22092 vdd.n1430 vdd.n1186 0.152939
R22093 vdd.n1431 vdd.n1430 0.152939
R22094 vdd.n1432 vdd.n1431 0.152939
R22095 vdd.n1432 vdd.n1174 0.152939
R22096 vdd.n1447 vdd.n1174 0.152939
R22097 vdd.n1448 vdd.n1447 0.152939
R22098 vdd.n1449 vdd.n1448 0.152939
R22099 vdd.n1449 vdd.n1164 0.152939
R22100 vdd.n1464 vdd.n1164 0.152939
R22101 vdd.n1465 vdd.n1464 0.152939
R22102 vdd.n1466 vdd.n1465 0.152939
R22103 vdd.n1466 vdd.n1151 0.152939
R22104 vdd.n1480 vdd.n1151 0.152939
R22105 vdd.n1481 vdd.n1480 0.152939
R22106 vdd.n1482 vdd.n1481 0.152939
R22107 vdd.n1482 vdd.n1140 0.152939
R22108 vdd.n1497 vdd.n1140 0.152939
R22109 vdd.n1498 vdd.n1497 0.152939
R22110 vdd.n1499 vdd.n1498 0.152939
R22111 vdd.n1499 vdd.n1129 0.152939
R22112 vdd.n1820 vdd.n1129 0.152939
R22113 vdd.n1821 vdd.n1820 0.152939
R22114 vdd.n1822 vdd.n1821 0.152939
R22115 vdd.n1822 vdd.n1117 0.152939
R22116 vdd.n1837 vdd.n1117 0.152939
R22117 vdd.n1838 vdd.n1837 0.152939
R22118 vdd.n1839 vdd.n1838 0.152939
R22119 vdd.n1839 vdd.n1107 0.152939
R22120 vdd.n1854 vdd.n1107 0.152939
R22121 vdd.n1855 vdd.n1854 0.152939
R22122 vdd.n1856 vdd.n1855 0.152939
R22123 vdd.n1856 vdd.n1094 0.152939
R22124 vdd.n1870 vdd.n1094 0.152939
R22125 vdd.n1871 vdd.n1870 0.152939
R22126 vdd.n1872 vdd.n1871 0.152939
R22127 vdd.n1872 vdd.n1084 0.152939
R22128 vdd.n1887 vdd.n1084 0.152939
R22129 vdd.n1888 vdd.n1887 0.152939
R22130 vdd.n1891 vdd.n1888 0.152939
R22131 vdd.n1891 vdd.n1890 0.152939
R22132 vdd.n1890 vdd.n1889 0.152939
R22133 vdd.n1422 vdd.n1191 0.152939
R22134 vdd.n1415 vdd.n1191 0.152939
R22135 vdd.n1415 vdd.n1414 0.152939
R22136 vdd.n1414 vdd.n1413 0.152939
R22137 vdd.n1413 vdd.n1228 0.152939
R22138 vdd.n1409 vdd.n1228 0.152939
R22139 vdd.n1409 vdd.n1408 0.152939
R22140 vdd.n1408 vdd.n1407 0.152939
R22141 vdd.n1407 vdd.n1234 0.152939
R22142 vdd.n1403 vdd.n1234 0.152939
R22143 vdd.n1403 vdd.n1402 0.152939
R22144 vdd.n1402 vdd.n1401 0.152939
R22145 vdd.n1401 vdd.n1240 0.152939
R22146 vdd.n1397 vdd.n1240 0.152939
R22147 vdd.n1397 vdd.n1396 0.152939
R22148 vdd.n1396 vdd.n1395 0.152939
R22149 vdd.n1395 vdd.n1246 0.152939
R22150 vdd.n1391 vdd.n1246 0.152939
R22151 vdd.n1391 vdd.n1390 0.152939
R22152 vdd.n1390 vdd.n1389 0.152939
R22153 vdd.n1389 vdd.n1254 0.152939
R22154 vdd.n1385 vdd.n1254 0.152939
R22155 vdd.n1385 vdd.n1384 0.152939
R22156 vdd.n1384 vdd.n1383 0.152939
R22157 vdd.n1383 vdd.n1260 0.152939
R22158 vdd.n1379 vdd.n1260 0.152939
R22159 vdd.n1379 vdd.n1378 0.152939
R22160 vdd.n1378 vdd.n1377 0.152939
R22161 vdd.n1377 vdd.n1266 0.152939
R22162 vdd.n1373 vdd.n1266 0.152939
R22163 vdd.n1373 vdd.n1372 0.152939
R22164 vdd.n1372 vdd.n1371 0.152939
R22165 vdd.n1371 vdd.n1272 0.152939
R22166 vdd.n1367 vdd.n1272 0.152939
R22167 vdd.n1367 vdd.n1366 0.152939
R22168 vdd.n1366 vdd.n1365 0.152939
R22169 vdd.n1365 vdd.n1278 0.152939
R22170 vdd.n1361 vdd.n1278 0.152939
R22171 vdd.n1361 vdd.n1360 0.152939
R22172 vdd.n1360 vdd.n1359 0.152939
R22173 vdd.n1359 vdd.n1284 0.152939
R22174 vdd.n1352 vdd.n1284 0.152939
R22175 vdd.n1352 vdd.n1351 0.152939
R22176 vdd.n1351 vdd.n1350 0.152939
R22177 vdd.n1350 vdd.n1289 0.152939
R22178 vdd.n1346 vdd.n1289 0.152939
R22179 vdd.n1346 vdd.n1345 0.152939
R22180 vdd.n1345 vdd.n1344 0.152939
R22181 vdd.n1344 vdd.n1295 0.152939
R22182 vdd.n1340 vdd.n1295 0.152939
R22183 vdd.n1340 vdd.n1339 0.152939
R22184 vdd.n1339 vdd.n1338 0.152939
R22185 vdd.n1338 vdd.n1301 0.152939
R22186 vdd.n1334 vdd.n1301 0.152939
R22187 vdd.n1334 vdd.n1333 0.152939
R22188 vdd.n1333 vdd.n1332 0.152939
R22189 vdd.n1332 vdd.n1307 0.152939
R22190 vdd.n1328 vdd.n1307 0.152939
R22191 vdd.n1328 vdd.n1327 0.152939
R22192 vdd.n1327 vdd.n1326 0.152939
R22193 vdd.n1326 vdd.n1313 0.152939
R22194 vdd.n1322 vdd.n1313 0.152939
R22195 vdd.n1322 vdd.n1321 0.152939
R22196 vdd.n1424 vdd.n1423 0.152939
R22197 vdd.n1424 vdd.n1180 0.152939
R22198 vdd.n1439 vdd.n1180 0.152939
R22199 vdd.n1440 vdd.n1439 0.152939
R22200 vdd.n1441 vdd.n1440 0.152939
R22201 vdd.n1441 vdd.n1169 0.152939
R22202 vdd.n1456 vdd.n1169 0.152939
R22203 vdd.n1457 vdd.n1456 0.152939
R22204 vdd.n1458 vdd.n1457 0.152939
R22205 vdd.n1458 vdd.n1158 0.152939
R22206 vdd.n1472 vdd.n1158 0.152939
R22207 vdd.n1473 vdd.n1472 0.152939
R22208 vdd.n1474 vdd.n1473 0.152939
R22209 vdd.n1474 vdd.n1146 0.152939
R22210 vdd.n1489 vdd.n1146 0.152939
R22211 vdd.n1490 vdd.n1489 0.152939
R22212 vdd.n1491 vdd.n1490 0.152939
R22213 vdd.n1491 vdd.n1135 0.152939
R22214 vdd.n1505 vdd.n1135 0.152939
R22215 vdd.n1506 vdd.n1505 0.152939
R22216 vdd.n1427 vdd.t226 0.113865
R22217 vdd.t233 vdd.n386 0.113865
R22218 vdd.n2315 vdd.n1900 0.110256
R22219 vdd.n3216 vdd.n727 0.110256
R22220 vdd.n3093 vdd.n687 0.110256
R22221 vdd.n2338 vdd.n2337 0.110256
R22222 vdd.n1814 vdd.n1813 0.0695946
R22223 vdd.n3399 vdd.n334 0.0695946
R22224 vdd.n3399 vdd.n3398 0.0695946
R22225 vdd.n1813 vdd.n1506 0.0695946
R22226 vdd.n2315 vdd.n2101 0.0431829
R22227 vdd.n2338 vdd.n1064 0.0431829
R22228 vdd.n3216 vdd.n730 0.0431829
R22229 vdd.n3093 vdd.n783 0.0431829
R22230 vdd vdd.n28 0.00833333
R22231 a_n1996_n452.n86 a_n1996_n452.t59 512.366
R22232 a_n1996_n452.n76 a_n1996_n452.t50 512.366
R22233 a_n1996_n452.n87 a_n1996_n452.t44 512.366
R22234 a_n1996_n452.n84 a_n1996_n452.t67 512.366
R22235 a_n1996_n452.n77 a_n1996_n452.t56 512.366
R22236 a_n1996_n452.n85 a_n1996_n452.t55 512.366
R22237 a_n1996_n452.n82 a_n1996_n452.t63 512.366
R22238 a_n1996_n452.n78 a_n1996_n452.t48 512.366
R22239 a_n1996_n452.n83 a_n1996_n452.t49 512.366
R22240 a_n1996_n452.n80 a_n1996_n452.t51 512.366
R22241 a_n1996_n452.n79 a_n1996_n452.t60 512.366
R22242 a_n1996_n452.n81 a_n1996_n452.t71 512.366
R22243 a_n1996_n452.n24 a_n1996_n452.t70 539.01
R22244 a_n1996_n452.n91 a_n1996_n452.t53 512.366
R22245 a_n1996_n452.n90 a_n1996_n452.t57 512.366
R22246 a_n1996_n452.n64 a_n1996_n452.t47 512.366
R22247 a_n1996_n452.n89 a_n1996_n452.t62 512.366
R22248 a_n1996_n452.n52 a_n1996_n452.t23 533.058
R22249 a_n1996_n452.n26 a_n1996_n452.t27 539.01
R22250 a_n1996_n452.n94 a_n1996_n452.t13 512.366
R22251 a_n1996_n452.n93 a_n1996_n452.t17 512.366
R22252 a_n1996_n452.n53 a_n1996_n452.t21 512.366
R22253 a_n1996_n452.n92 a_n1996_n452.t7 512.366
R22254 a_n1996_n452.n16 a_n1996_n452.t19 539.01
R22255 a_n1996_n452.n72 a_n1996_n452.t15 512.366
R22256 a_n1996_n452.n73 a_n1996_n452.t9 512.366
R22257 a_n1996_n452.n67 a_n1996_n452.t11 512.366
R22258 a_n1996_n452.n74 a_n1996_n452.t25 512.366
R22259 a_n1996_n452.n20 a_n1996_n452.t65 539.01
R22260 a_n1996_n452.n69 a_n1996_n452.t66 512.366
R22261 a_n1996_n452.n70 a_n1996_n452.t45 512.366
R22262 a_n1996_n452.n68 a_n1996_n452.t52 512.366
R22263 a_n1996_n452.n71 a_n1996_n452.t61 512.366
R22264 a_n1996_n452.n4 a_n1996_n452.n51 70.1674
R22265 a_n1996_n452.n6 a_n1996_n452.n49 70.1674
R22266 a_n1996_n452.n8 a_n1996_n452.n47 70.1674
R22267 a_n1996_n452.n11 a_n1996_n452.n45 70.1674
R22268 a_n1996_n452.n37 a_n1996_n452.n22 70.3058
R22269 a_n1996_n452.n31 a_n1996_n452.n34 70.1674
R22270 a_n1996_n452.n34 a_n1996_n452.n53 20.9683
R22271 a_n1996_n452.n33 a_n1996_n452.n32 75.0448
R22272 a_n1996_n452.n93 a_n1996_n452.n33 11.2134
R22273 a_n1996_n452.n25 a_n1996_n452.n26 44.8194
R22274 a_n1996_n452.n52 a_n1996_n452.n31 70.3058
R22275 a_n1996_n452.n23 a_n1996_n452.n36 70.1674
R22276 a_n1996_n452.n36 a_n1996_n452.n64 20.9683
R22277 a_n1996_n452.n35 a_n1996_n452.n23 75.0448
R22278 a_n1996_n452.n90 a_n1996_n452.n35 11.2134
R22279 a_n1996_n452.n21 a_n1996_n452.n24 44.8194
R22280 a_n1996_n452.n13 a_n1996_n452.n43 70.3058
R22281 a_n1996_n452.n17 a_n1996_n452.n40 70.3058
R22282 a_n1996_n452.n39 a_n1996_n452.n18 70.1674
R22283 a_n1996_n452.n39 a_n1996_n452.n68 20.9683
R22284 a_n1996_n452.n18 a_n1996_n452.n38 75.0448
R22285 a_n1996_n452.n70 a_n1996_n452.n38 11.2134
R22286 a_n1996_n452.n19 a_n1996_n452.n20 44.8194
R22287 a_n1996_n452.n42 a_n1996_n452.n14 70.1674
R22288 a_n1996_n452.n42 a_n1996_n452.n67 20.9683
R22289 a_n1996_n452.n14 a_n1996_n452.n41 75.0448
R22290 a_n1996_n452.n73 a_n1996_n452.n41 11.2134
R22291 a_n1996_n452.n15 a_n1996_n452.n16 44.8194
R22292 a_n1996_n452.n81 a_n1996_n452.n45 20.9683
R22293 a_n1996_n452.n44 a_n1996_n452.n12 75.0448
R22294 a_n1996_n452.n44 a_n1996_n452.n79 11.2134
R22295 a_n1996_n452.n12 a_n1996_n452.n80 161.3
R22296 a_n1996_n452.n83 a_n1996_n452.n47 20.9683
R22297 a_n1996_n452.n46 a_n1996_n452.n9 75.0448
R22298 a_n1996_n452.n46 a_n1996_n452.n78 11.2134
R22299 a_n1996_n452.n9 a_n1996_n452.n82 161.3
R22300 a_n1996_n452.n85 a_n1996_n452.n49 20.9683
R22301 a_n1996_n452.n48 a_n1996_n452.n7 75.0448
R22302 a_n1996_n452.n48 a_n1996_n452.n77 11.2134
R22303 a_n1996_n452.n7 a_n1996_n452.n84 161.3
R22304 a_n1996_n452.n87 a_n1996_n452.n51 20.9683
R22305 a_n1996_n452.n50 a_n1996_n452.n5 75.0448
R22306 a_n1996_n452.n50 a_n1996_n452.n76 11.2134
R22307 a_n1996_n452.n5 a_n1996_n452.n86 161.3
R22308 a_n1996_n452.n3 a_n1996_n452.n62 81.3764
R22309 a_n1996_n452.n1 a_n1996_n452.n57 81.3764
R22310 a_n1996_n452.n0 a_n1996_n452.n54 81.3764
R22311 a_n1996_n452.n3 a_n1996_n452.n63 80.9324
R22312 a_n1996_n452.n3 a_n1996_n452.n61 80.9324
R22313 a_n1996_n452.n2 a_n1996_n452.n60 80.9324
R22314 a_n1996_n452.n2 a_n1996_n452.n59 80.9324
R22315 a_n1996_n452.n1 a_n1996_n452.n58 80.9324
R22316 a_n1996_n452.n1 a_n1996_n452.n56 80.9324
R22317 a_n1996_n452.n0 a_n1996_n452.n55 80.9324
R22318 a_n1996_n452.n30 a_n1996_n452.t24 74.6477
R22319 a_n1996_n452.n27 a_n1996_n452.t20 74.6477
R22320 a_n1996_n452.n29 a_n1996_n452.t28 74.2899
R22321 a_n1996_n452.n28 a_n1996_n452.t30 74.2897
R22322 a_n1996_n452.n30 a_n1996_n452.n96 70.6783
R22323 a_n1996_n452.n28 a_n1996_n452.n66 70.6783
R22324 a_n1996_n452.n27 a_n1996_n452.n65 70.6783
R22325 a_n1996_n452.n97 a_n1996_n452.n30 70.6782
R22326 a_n1996_n452.n86 a_n1996_n452.n76 48.2005
R22327 a_n1996_n452.t64 a_n1996_n452.n51 533.335
R22328 a_n1996_n452.n84 a_n1996_n452.n77 48.2005
R22329 a_n1996_n452.t69 a_n1996_n452.n49 533.335
R22330 a_n1996_n452.n82 a_n1996_n452.n78 48.2005
R22331 a_n1996_n452.t58 a_n1996_n452.n47 533.335
R22332 a_n1996_n452.n80 a_n1996_n452.n79 48.2005
R22333 a_n1996_n452.t54 a_n1996_n452.n45 533.335
R22334 a_n1996_n452.n91 a_n1996_n452.n90 48.2005
R22335 a_n1996_n452.n89 a_n1996_n452.n36 20.9683
R22336 a_n1996_n452.n94 a_n1996_n452.n93 48.2005
R22337 a_n1996_n452.n92 a_n1996_n452.n34 20.9683
R22338 a_n1996_n452.n73 a_n1996_n452.n72 48.2005
R22339 a_n1996_n452.n74 a_n1996_n452.n42 20.9683
R22340 a_n1996_n452.n70 a_n1996_n452.n69 48.2005
R22341 a_n1996_n452.n71 a_n1996_n452.n39 20.9683
R22342 a_n1996_n452.n37 a_n1996_n452.t68 533.058
R22343 a_n1996_n452.t29 a_n1996_n452.n43 533.058
R22344 a_n1996_n452.t46 a_n1996_n452.n40 533.058
R22345 a_n1996_n452.n2 a_n1996_n452.n1 32.0139
R22346 a_n1996_n452.n87 a_n1996_n452.n50 35.3134
R22347 a_n1996_n452.n85 a_n1996_n452.n48 35.3134
R22348 a_n1996_n452.n83 a_n1996_n452.n46 35.3134
R22349 a_n1996_n452.n81 a_n1996_n452.n44 35.3134
R22350 a_n1996_n452.n35 a_n1996_n452.n64 35.3134
R22351 a_n1996_n452.n33 a_n1996_n452.n53 35.3134
R22352 a_n1996_n452.n67 a_n1996_n452.n41 35.3134
R22353 a_n1996_n452.n68 a_n1996_n452.n38 35.3134
R22354 a_n1996_n452.n31 a_n1996_n452.n3 23.891
R22355 a_n1996_n452.n19 a_n1996_n452.n10 12.046
R22356 a_n1996_n452.n22 a_n1996_n452.n88 11.8414
R22357 a_n1996_n452.n95 a_n1996_n452.n25 10.5365
R22358 a_n1996_n452.n75 a_n1996_n452.n28 9.50122
R22359 a_n1996_n452.n88 a_n1996_n452.n4 7.47588
R22360 a_n1996_n452.n12 a_n1996_n452.n10 7.47588
R22361 a_n1996_n452.n75 a_n1996_n452.n13 6.70126
R22362 a_n1996_n452.n29 a_n1996_n452.n95 5.65783
R22363 a_n1996_n452.n88 a_n1996_n452.n75 5.3452
R22364 a_n1996_n452.n31 a_n1996_n452.n21 3.95126
R22365 a_n1996_n452.n15 a_n1996_n452.n17 3.95126
R22366 a_n1996_n452.n96 a_n1996_n452.t14 3.61217
R22367 a_n1996_n452.n96 a_n1996_n452.t18 3.61217
R22368 a_n1996_n452.n66 a_n1996_n452.t12 3.61217
R22369 a_n1996_n452.n66 a_n1996_n452.t26 3.61217
R22370 a_n1996_n452.n65 a_n1996_n452.t16 3.61217
R22371 a_n1996_n452.n65 a_n1996_n452.t10 3.61217
R22372 a_n1996_n452.n97 a_n1996_n452.t22 3.61217
R22373 a_n1996_n452.t8 a_n1996_n452.n97 3.61217
R22374 a_n1996_n452.n62 a_n1996_n452.t39 2.82907
R22375 a_n1996_n452.n62 a_n1996_n452.t38 2.82907
R22376 a_n1996_n452.n63 a_n1996_n452.t40 2.82907
R22377 a_n1996_n452.n63 a_n1996_n452.t0 2.82907
R22378 a_n1996_n452.n61 a_n1996_n452.t31 2.82907
R22379 a_n1996_n452.n61 a_n1996_n452.t35 2.82907
R22380 a_n1996_n452.n60 a_n1996_n452.t6 2.82907
R22381 a_n1996_n452.n60 a_n1996_n452.t34 2.82907
R22382 a_n1996_n452.n59 a_n1996_n452.t43 2.82907
R22383 a_n1996_n452.n59 a_n1996_n452.t5 2.82907
R22384 a_n1996_n452.n57 a_n1996_n452.t41 2.82907
R22385 a_n1996_n452.n57 a_n1996_n452.t3 2.82907
R22386 a_n1996_n452.n58 a_n1996_n452.t33 2.82907
R22387 a_n1996_n452.n58 a_n1996_n452.t42 2.82907
R22388 a_n1996_n452.n56 a_n1996_n452.t37 2.82907
R22389 a_n1996_n452.n56 a_n1996_n452.t36 2.82907
R22390 a_n1996_n452.n55 a_n1996_n452.t4 2.82907
R22391 a_n1996_n452.n55 a_n1996_n452.t2 2.82907
R22392 a_n1996_n452.n54 a_n1996_n452.t32 2.82907
R22393 a_n1996_n452.n54 a_n1996_n452.t1 2.82907
R22394 a_n1996_n452.n95 a_n1996_n452.n10 1.30542
R22395 a_n1996_n452.n7 a_n1996_n452.n8 1.04595
R22396 a_n1996_n452.n24 a_n1996_n452.n91 13.657
R22397 a_n1996_n452.n89 a_n1996_n452.n37 21.4216
R22398 a_n1996_n452.n26 a_n1996_n452.n94 13.657
R22399 a_n1996_n452.n92 a_n1996_n452.n52 21.4216
R22400 a_n1996_n452.n72 a_n1996_n452.n16 13.657
R22401 a_n1996_n452.n43 a_n1996_n452.n74 21.4216
R22402 a_n1996_n452.n69 a_n1996_n452.n20 13.657
R22403 a_n1996_n452.n40 a_n1996_n452.n71 21.4216
R22404 a_n1996_n452.n3 a_n1996_n452.n2 1.3324
R22405 a_n1996_n452.n1 a_n1996_n452.n0 0.888431
R22406 a_n1996_n452.n32 a_n1996_n452.n25 0.758076
R22407 a_n1996_n452.n23 a_n1996_n452.n21 0.758076
R22408 a_n1996_n452.n23 a_n1996_n452.n22 0.758076
R22409 a_n1996_n452.n19 a_n1996_n452.n18 0.758076
R22410 a_n1996_n452.n18 a_n1996_n452.n17 0.758076
R22411 a_n1996_n452.n15 a_n1996_n452.n14 0.758076
R22412 a_n1996_n452.n14 a_n1996_n452.n13 0.758076
R22413 a_n1996_n452.n12 a_n1996_n452.n11 0.758076
R22414 a_n1996_n452.n9 a_n1996_n452.n8 0.758076
R22415 a_n1996_n452.n7 a_n1996_n452.n6 0.758076
R22416 a_n1996_n452.n5 a_n1996_n452.n4 0.758076
R22417 a_n1996_n452.n32 a_n1996_n452.n31 0.720197
R22418 a_n1996_n452.n30 a_n1996_n452.n29 0.716017
R22419 a_n1996_n452.n28 a_n1996_n452.n27 0.716017
R22420 a_n1996_n452.n9 a_n1996_n452.n11 0.67853
R22421 a_n1996_n452.n5 a_n1996_n452.n6 0.67853
R22422 a_n1808_13878.n17 a_n1808_13878.n16 98.9632
R22423 a_n1808_13878.n2 a_n1808_13878.n0 98.7517
R22424 a_n1808_13878.n16 a_n1808_13878.n15 98.6055
R22425 a_n1808_13878.n4 a_n1808_13878.n3 98.6055
R22426 a_n1808_13878.n2 a_n1808_13878.n1 98.6055
R22427 a_n1808_13878.n14 a_n1808_13878.n13 98.6054
R22428 a_n1808_13878.n6 a_n1808_13878.t13 74.6477
R22429 a_n1808_13878.n11 a_n1808_13878.t14 74.2899
R22430 a_n1808_13878.n8 a_n1808_13878.t15 74.2899
R22431 a_n1808_13878.n7 a_n1808_13878.t12 74.2899
R22432 a_n1808_13878.n10 a_n1808_13878.n9 70.6783
R22433 a_n1808_13878.n6 a_n1808_13878.n5 70.6783
R22434 a_n1808_13878.n12 a_n1808_13878.n4 13.5694
R22435 a_n1808_13878.n14 a_n1808_13878.n12 11.5762
R22436 a_n1808_13878.n12 a_n1808_13878.n11 6.2408
R22437 a_n1808_13878.n13 a_n1808_13878.t9 3.61217
R22438 a_n1808_13878.n13 a_n1808_13878.t10 3.61217
R22439 a_n1808_13878.n15 a_n1808_13878.t0 3.61217
R22440 a_n1808_13878.n15 a_n1808_13878.t5 3.61217
R22441 a_n1808_13878.n9 a_n1808_13878.t18 3.61217
R22442 a_n1808_13878.n9 a_n1808_13878.t19 3.61217
R22443 a_n1808_13878.n5 a_n1808_13878.t16 3.61217
R22444 a_n1808_13878.n5 a_n1808_13878.t17 3.61217
R22445 a_n1808_13878.n3 a_n1808_13878.t6 3.61217
R22446 a_n1808_13878.n3 a_n1808_13878.t1 3.61217
R22447 a_n1808_13878.n1 a_n1808_13878.t8 3.61217
R22448 a_n1808_13878.n1 a_n1808_13878.t3 3.61217
R22449 a_n1808_13878.n0 a_n1808_13878.t2 3.61217
R22450 a_n1808_13878.n0 a_n1808_13878.t4 3.61217
R22451 a_n1808_13878.n17 a_n1808_13878.t7 3.61217
R22452 a_n1808_13878.t11 a_n1808_13878.n17 3.61217
R22453 a_n1808_13878.n7 a_n1808_13878.n6 0.358259
R22454 a_n1808_13878.n10 a_n1808_13878.n8 0.358259
R22455 a_n1808_13878.n11 a_n1808_13878.n10 0.358259
R22456 a_n1808_13878.n16 a_n1808_13878.n14 0.358259
R22457 a_n1808_13878.n4 a_n1808_13878.n2 0.146627
R22458 a_n1808_13878.n8 a_n1808_13878.n7 0.101793
R22459 a_n1986_8322.n6 a_n1986_8322.t15 74.6477
R22460 a_n1986_8322.n1 a_n1986_8322.t1 74.6477
R22461 a_n1986_8322.n16 a_n1986_8322.t10 74.6474
R22462 a_n1986_8322.n14 a_n1986_8322.t3 74.2899
R22463 a_n1986_8322.n7 a_n1986_8322.t13 74.2899
R22464 a_n1986_8322.n8 a_n1986_8322.t16 74.2899
R22465 a_n1986_8322.n11 a_n1986_8322.t17 74.2899
R22466 a_n1986_8322.n4 a_n1986_8322.t0 74.2899
R22467 a_n1986_8322.n16 a_n1986_8322.n15 70.6783
R22468 a_n1986_8322.n6 a_n1986_8322.n5 70.6783
R22469 a_n1986_8322.n10 a_n1986_8322.n9 70.6783
R22470 a_n1986_8322.n1 a_n1986_8322.n0 70.6783
R22471 a_n1986_8322.n3 a_n1986_8322.n2 70.6783
R22472 a_n1986_8322.n18 a_n1986_8322.n17 70.6782
R22473 a_n1986_8322.n12 a_n1986_8322.n4 22.7556
R22474 a_n1986_8322.n13 a_n1986_8322.t21 9.96389
R22475 a_n1986_8322.n12 a_n1986_8322.n11 6.2408
R22476 a_n1986_8322.n14 a_n1986_8322.n13 5.83671
R22477 a_n1986_8322.n13 a_n1986_8322.n12 5.3452
R22478 a_n1986_8322.n15 a_n1986_8322.t8 3.61217
R22479 a_n1986_8322.n15 a_n1986_8322.t5 3.61217
R22480 a_n1986_8322.n5 a_n1986_8322.t19 3.61217
R22481 a_n1986_8322.n5 a_n1986_8322.t18 3.61217
R22482 a_n1986_8322.n9 a_n1986_8322.t14 3.61217
R22483 a_n1986_8322.n9 a_n1986_8322.t12 3.61217
R22484 a_n1986_8322.n0 a_n1986_8322.t9 3.61217
R22485 a_n1986_8322.n0 a_n1986_8322.t4 3.61217
R22486 a_n1986_8322.n2 a_n1986_8322.t7 3.61217
R22487 a_n1986_8322.n2 a_n1986_8322.t6 3.61217
R22488 a_n1986_8322.n18 a_n1986_8322.t2 3.61217
R22489 a_n1986_8322.t11 a_n1986_8322.n18 3.61217
R22490 a_n1986_8322.n11 a_n1986_8322.n10 0.358259
R22491 a_n1986_8322.n10 a_n1986_8322.n8 0.358259
R22492 a_n1986_8322.n7 a_n1986_8322.n6 0.358259
R22493 a_n1986_8322.n4 a_n1986_8322.n3 0.358259
R22494 a_n1986_8322.n3 a_n1986_8322.n1 0.358259
R22495 a_n1986_8322.n17 a_n1986_8322.n14 0.358259
R22496 a_n1986_8322.n17 a_n1986_8322.n16 0.358259
R22497 a_n1986_8322.n8 a_n1986_8322.n7 0.101793
R22498 a_n1986_8322.t21 a_n1986_8322.t20 0.057021
R22499 minus.n43 minus.t24 322.512
R22500 minus.n9 minus.t8 322.512
R22501 minus.n66 minus.t5 297.12
R22502 minus.n64 minus.t6 297.12
R22503 minus.n36 minus.t22 297.12
R22504 minus.n58 minus.t18 297.12
R22505 minus.n38 minus.t19 297.12
R22506 minus.n52 minus.t14 297.12
R22507 minus.n40 minus.t15 297.12
R22508 minus.n46 minus.t9 297.12
R22509 minus.n42 minus.t23 297.12
R22510 minus.n8 minus.t7 297.12
R22511 minus.n12 minus.t11 297.12
R22512 minus.n14 minus.t10 297.12
R22513 minus.n18 minus.t12 297.12
R22514 minus.n20 minus.t17 297.12
R22515 minus.n24 minus.t16 297.12
R22516 minus.n26 minus.t21 297.12
R22517 minus.n30 minus.t20 297.12
R22518 minus.n32 minus.t13 297.12
R22519 minus.n72 minus.t4 243.255
R22520 minus.n71 minus.n69 224.169
R22521 minus.n71 minus.n70 223.454
R22522 minus.n45 minus.n44 161.3
R22523 minus.n46 minus.n41 161.3
R22524 minus.n48 minus.n47 161.3
R22525 minus.n49 minus.n40 161.3
R22526 minus.n51 minus.n50 161.3
R22527 minus.n52 minus.n39 161.3
R22528 minus.n54 minus.n53 161.3
R22529 minus.n55 minus.n38 161.3
R22530 minus.n57 minus.n56 161.3
R22531 minus.n58 minus.n37 161.3
R22532 minus.n60 minus.n59 161.3
R22533 minus.n61 minus.n36 161.3
R22534 minus.n63 minus.n62 161.3
R22535 minus.n64 minus.n35 161.3
R22536 minus.n65 minus.n34 161.3
R22537 minus.n67 minus.n66 161.3
R22538 minus.n33 minus.n32 161.3
R22539 minus.n31 minus.n0 161.3
R22540 minus.n30 minus.n29 161.3
R22541 minus.n28 minus.n1 161.3
R22542 minus.n27 minus.n26 161.3
R22543 minus.n25 minus.n2 161.3
R22544 minus.n24 minus.n23 161.3
R22545 minus.n22 minus.n3 161.3
R22546 minus.n21 minus.n20 161.3
R22547 minus.n19 minus.n4 161.3
R22548 minus.n18 minus.n17 161.3
R22549 minus.n16 minus.n5 161.3
R22550 minus.n15 minus.n14 161.3
R22551 minus.n13 minus.n6 161.3
R22552 minus.n12 minus.n11 161.3
R22553 minus.n10 minus.n7 161.3
R22554 minus.n44 minus.n43 45.0031
R22555 minus.n10 minus.n9 45.0031
R22556 minus.n66 minus.n65 41.6278
R22557 minus.n32 minus.n31 41.6278
R22558 minus.n64 minus.n63 37.246
R22559 minus.n45 minus.n42 37.246
R22560 minus.n8 minus.n7 37.246
R22561 minus.n30 minus.n1 37.246
R22562 minus.n59 minus.n36 32.8641
R22563 minus.n47 minus.n46 32.8641
R22564 minus.n13 minus.n12 32.8641
R22565 minus.n26 minus.n25 32.8641
R22566 minus.n68 minus.n67 31.8206
R22567 minus.n58 minus.n57 28.4823
R22568 minus.n51 minus.n40 28.4823
R22569 minus.n14 minus.n5 28.4823
R22570 minus.n24 minus.n3 28.4823
R22571 minus.n53 minus.n38 24.1005
R22572 minus.n53 minus.n52 24.1005
R22573 minus.n19 minus.n18 24.1005
R22574 minus.n20 minus.n19 24.1005
R22575 minus.n70 minus.t3 19.8005
R22576 minus.n70 minus.t1 19.8005
R22577 minus.n69 minus.t2 19.8005
R22578 minus.n69 minus.t0 19.8005
R22579 minus.n57 minus.n38 19.7187
R22580 minus.n52 minus.n51 19.7187
R22581 minus.n18 minus.n5 19.7187
R22582 minus.n20 minus.n3 19.7187
R22583 minus.n43 minus.n42 15.6319
R22584 minus.n9 minus.n8 15.6319
R22585 minus.n59 minus.n58 15.3369
R22586 minus.n47 minus.n40 15.3369
R22587 minus.n14 minus.n13 15.3369
R22588 minus.n25 minus.n24 15.3369
R22589 minus.n68 minus.n33 12.0819
R22590 minus minus.n73 11.5399
R22591 minus.n63 minus.n36 10.955
R22592 minus.n46 minus.n45 10.955
R22593 minus.n12 minus.n7 10.955
R22594 minus.n26 minus.n1 10.955
R22595 minus.n65 minus.n64 6.57323
R22596 minus.n31 minus.n30 6.57323
R22597 minus.n73 minus.n72 4.80222
R22598 minus.n73 minus.n68 0.972091
R22599 minus.n72 minus.n71 0.716017
R22600 minus.n67 minus.n34 0.189894
R22601 minus.n35 minus.n34 0.189894
R22602 minus.n62 minus.n35 0.189894
R22603 minus.n62 minus.n61 0.189894
R22604 minus.n61 minus.n60 0.189894
R22605 minus.n60 minus.n37 0.189894
R22606 minus.n56 minus.n37 0.189894
R22607 minus.n56 minus.n55 0.189894
R22608 minus.n55 minus.n54 0.189894
R22609 minus.n54 minus.n39 0.189894
R22610 minus.n50 minus.n39 0.189894
R22611 minus.n50 minus.n49 0.189894
R22612 minus.n49 minus.n48 0.189894
R22613 minus.n48 minus.n41 0.189894
R22614 minus.n44 minus.n41 0.189894
R22615 minus.n11 minus.n10 0.189894
R22616 minus.n11 minus.n6 0.189894
R22617 minus.n15 minus.n6 0.189894
R22618 minus.n16 minus.n15 0.189894
R22619 minus.n17 minus.n16 0.189894
R22620 minus.n17 minus.n4 0.189894
R22621 minus.n21 minus.n4 0.189894
R22622 minus.n22 minus.n21 0.189894
R22623 minus.n23 minus.n22 0.189894
R22624 minus.n23 minus.n2 0.189894
R22625 minus.n27 minus.n2 0.189894
R22626 minus.n28 minus.n27 0.189894
R22627 minus.n29 minus.n28 0.189894
R22628 minus.n29 minus.n0 0.189894
R22629 minus.n33 minus.n0 0.189894
R22630 output.n41 output.n15 289.615
R22631 output.n72 output.n46 289.615
R22632 output.n104 output.n78 289.615
R22633 output.n136 output.n110 289.615
R22634 output.n77 output.n45 197.26
R22635 output.n77 output.n76 196.298
R22636 output.n109 output.n108 196.298
R22637 output.n141 output.n140 196.298
R22638 output.n42 output.n41 185
R22639 output.n40 output.n39 185
R22640 output.n19 output.n18 185
R22641 output.n34 output.n33 185
R22642 output.n32 output.n31 185
R22643 output.n23 output.n22 185
R22644 output.n26 output.n25 185
R22645 output.n73 output.n72 185
R22646 output.n71 output.n70 185
R22647 output.n50 output.n49 185
R22648 output.n65 output.n64 185
R22649 output.n63 output.n62 185
R22650 output.n54 output.n53 185
R22651 output.n57 output.n56 185
R22652 output.n105 output.n104 185
R22653 output.n103 output.n102 185
R22654 output.n82 output.n81 185
R22655 output.n97 output.n96 185
R22656 output.n95 output.n94 185
R22657 output.n86 output.n85 185
R22658 output.n89 output.n88 185
R22659 output.n137 output.n136 185
R22660 output.n135 output.n134 185
R22661 output.n114 output.n113 185
R22662 output.n129 output.n128 185
R22663 output.n127 output.n126 185
R22664 output.n118 output.n117 185
R22665 output.n121 output.n120 185
R22666 output.t0 output.n24 147.661
R22667 output.t18 output.n55 147.661
R22668 output.t1 output.n87 147.661
R22669 output.t19 output.n119 147.661
R22670 output.n41 output.n40 104.615
R22671 output.n40 output.n18 104.615
R22672 output.n33 output.n18 104.615
R22673 output.n33 output.n32 104.615
R22674 output.n32 output.n22 104.615
R22675 output.n25 output.n22 104.615
R22676 output.n72 output.n71 104.615
R22677 output.n71 output.n49 104.615
R22678 output.n64 output.n49 104.615
R22679 output.n64 output.n63 104.615
R22680 output.n63 output.n53 104.615
R22681 output.n56 output.n53 104.615
R22682 output.n104 output.n103 104.615
R22683 output.n103 output.n81 104.615
R22684 output.n96 output.n81 104.615
R22685 output.n96 output.n95 104.615
R22686 output.n95 output.n85 104.615
R22687 output.n88 output.n85 104.615
R22688 output.n136 output.n135 104.615
R22689 output.n135 output.n113 104.615
R22690 output.n128 output.n113 104.615
R22691 output.n128 output.n127 104.615
R22692 output.n127 output.n117 104.615
R22693 output.n120 output.n117 104.615
R22694 output.n1 output.t13 77.056
R22695 output.n14 output.t15 76.6694
R22696 output.n1 output.n0 72.7095
R22697 output.n3 output.n2 72.7095
R22698 output.n5 output.n4 72.7095
R22699 output.n7 output.n6 72.7095
R22700 output.n9 output.n8 72.7095
R22701 output.n11 output.n10 72.7095
R22702 output.n13 output.n12 72.7095
R22703 output.n25 output.t0 52.3082
R22704 output.n56 output.t18 52.3082
R22705 output.n88 output.t1 52.3082
R22706 output.n120 output.t19 52.3082
R22707 output.n26 output.n24 15.6674
R22708 output.n57 output.n55 15.6674
R22709 output.n89 output.n87 15.6674
R22710 output.n121 output.n119 15.6674
R22711 output.n27 output.n23 12.8005
R22712 output.n58 output.n54 12.8005
R22713 output.n90 output.n86 12.8005
R22714 output.n122 output.n118 12.8005
R22715 output.n31 output.n30 12.0247
R22716 output.n62 output.n61 12.0247
R22717 output.n94 output.n93 12.0247
R22718 output.n126 output.n125 12.0247
R22719 output.n34 output.n21 11.249
R22720 output.n65 output.n52 11.249
R22721 output.n97 output.n84 11.249
R22722 output.n129 output.n116 11.249
R22723 output.n35 output.n19 10.4732
R22724 output.n66 output.n50 10.4732
R22725 output.n98 output.n82 10.4732
R22726 output.n130 output.n114 10.4732
R22727 output.n39 output.n38 9.69747
R22728 output.n70 output.n69 9.69747
R22729 output.n102 output.n101 9.69747
R22730 output.n134 output.n133 9.69747
R22731 output.n45 output.n44 9.45567
R22732 output.n76 output.n75 9.45567
R22733 output.n108 output.n107 9.45567
R22734 output.n140 output.n139 9.45567
R22735 output.n44 output.n43 9.3005
R22736 output.n17 output.n16 9.3005
R22737 output.n38 output.n37 9.3005
R22738 output.n36 output.n35 9.3005
R22739 output.n21 output.n20 9.3005
R22740 output.n30 output.n29 9.3005
R22741 output.n28 output.n27 9.3005
R22742 output.n75 output.n74 9.3005
R22743 output.n48 output.n47 9.3005
R22744 output.n69 output.n68 9.3005
R22745 output.n67 output.n66 9.3005
R22746 output.n52 output.n51 9.3005
R22747 output.n61 output.n60 9.3005
R22748 output.n59 output.n58 9.3005
R22749 output.n107 output.n106 9.3005
R22750 output.n80 output.n79 9.3005
R22751 output.n101 output.n100 9.3005
R22752 output.n99 output.n98 9.3005
R22753 output.n84 output.n83 9.3005
R22754 output.n93 output.n92 9.3005
R22755 output.n91 output.n90 9.3005
R22756 output.n139 output.n138 9.3005
R22757 output.n112 output.n111 9.3005
R22758 output.n133 output.n132 9.3005
R22759 output.n131 output.n130 9.3005
R22760 output.n116 output.n115 9.3005
R22761 output.n125 output.n124 9.3005
R22762 output.n123 output.n122 9.3005
R22763 output.n42 output.n17 8.92171
R22764 output.n73 output.n48 8.92171
R22765 output.n105 output.n80 8.92171
R22766 output.n137 output.n112 8.92171
R22767 output output.n141 8.15037
R22768 output.n43 output.n15 8.14595
R22769 output.n74 output.n46 8.14595
R22770 output.n106 output.n78 8.14595
R22771 output.n138 output.n110 8.14595
R22772 output.n45 output.n15 5.81868
R22773 output.n76 output.n46 5.81868
R22774 output.n108 output.n78 5.81868
R22775 output.n140 output.n110 5.81868
R22776 output.n43 output.n42 5.04292
R22777 output.n74 output.n73 5.04292
R22778 output.n106 output.n105 5.04292
R22779 output.n138 output.n137 5.04292
R22780 output.n28 output.n24 4.38594
R22781 output.n59 output.n55 4.38594
R22782 output.n91 output.n87 4.38594
R22783 output.n123 output.n119 4.38594
R22784 output.n39 output.n17 4.26717
R22785 output.n70 output.n48 4.26717
R22786 output.n102 output.n80 4.26717
R22787 output.n134 output.n112 4.26717
R22788 output.n0 output.t3 3.9605
R22789 output.n0 output.t8 3.9605
R22790 output.n2 output.t12 3.9605
R22791 output.n2 output.t4 3.9605
R22792 output.n4 output.t6 3.9605
R22793 output.n4 output.t5 3.9605
R22794 output.n6 output.t11 3.9605
R22795 output.n6 output.t14 3.9605
R22796 output.n8 output.t16 3.9605
R22797 output.n8 output.t9 3.9605
R22798 output.n10 output.t10 3.9605
R22799 output.n10 output.t17 3.9605
R22800 output.n12 output.t2 3.9605
R22801 output.n12 output.t7 3.9605
R22802 output.n38 output.n19 3.49141
R22803 output.n69 output.n50 3.49141
R22804 output.n101 output.n82 3.49141
R22805 output.n133 output.n114 3.49141
R22806 output.n35 output.n34 2.71565
R22807 output.n66 output.n65 2.71565
R22808 output.n98 output.n97 2.71565
R22809 output.n130 output.n129 2.71565
R22810 output.n31 output.n21 1.93989
R22811 output.n62 output.n52 1.93989
R22812 output.n94 output.n84 1.93989
R22813 output.n126 output.n116 1.93989
R22814 output.n30 output.n23 1.16414
R22815 output.n61 output.n54 1.16414
R22816 output.n93 output.n86 1.16414
R22817 output.n125 output.n118 1.16414
R22818 output.n141 output.n109 0.962709
R22819 output.n109 output.n77 0.962709
R22820 output.n27 output.n26 0.388379
R22821 output.n58 output.n57 0.388379
R22822 output.n90 output.n89 0.388379
R22823 output.n122 output.n121 0.388379
R22824 output.n14 output.n13 0.387128
R22825 output.n13 output.n11 0.387128
R22826 output.n11 output.n9 0.387128
R22827 output.n9 output.n7 0.387128
R22828 output.n7 output.n5 0.387128
R22829 output.n5 output.n3 0.387128
R22830 output.n3 output.n1 0.387128
R22831 output.n44 output.n16 0.155672
R22832 output.n37 output.n16 0.155672
R22833 output.n37 output.n36 0.155672
R22834 output.n36 output.n20 0.155672
R22835 output.n29 output.n20 0.155672
R22836 output.n29 output.n28 0.155672
R22837 output.n75 output.n47 0.155672
R22838 output.n68 output.n47 0.155672
R22839 output.n68 output.n67 0.155672
R22840 output.n67 output.n51 0.155672
R22841 output.n60 output.n51 0.155672
R22842 output.n60 output.n59 0.155672
R22843 output.n107 output.n79 0.155672
R22844 output.n100 output.n79 0.155672
R22845 output.n100 output.n99 0.155672
R22846 output.n99 output.n83 0.155672
R22847 output.n92 output.n83 0.155672
R22848 output.n92 output.n91 0.155672
R22849 output.n139 output.n111 0.155672
R22850 output.n132 output.n111 0.155672
R22851 output.n132 output.n131 0.155672
R22852 output.n131 output.n115 0.155672
R22853 output.n124 output.n115 0.155672
R22854 output.n124 output.n123 0.155672
R22855 output output.n14 0.126227
R22856 outputibias.n27 outputibias.n1 289.615
R22857 outputibias.n58 outputibias.n32 289.615
R22858 outputibias.n90 outputibias.n64 289.615
R22859 outputibias.n122 outputibias.n96 289.615
R22860 outputibias.n28 outputibias.n27 185
R22861 outputibias.n26 outputibias.n25 185
R22862 outputibias.n5 outputibias.n4 185
R22863 outputibias.n20 outputibias.n19 185
R22864 outputibias.n18 outputibias.n17 185
R22865 outputibias.n9 outputibias.n8 185
R22866 outputibias.n12 outputibias.n11 185
R22867 outputibias.n59 outputibias.n58 185
R22868 outputibias.n57 outputibias.n56 185
R22869 outputibias.n36 outputibias.n35 185
R22870 outputibias.n51 outputibias.n50 185
R22871 outputibias.n49 outputibias.n48 185
R22872 outputibias.n40 outputibias.n39 185
R22873 outputibias.n43 outputibias.n42 185
R22874 outputibias.n91 outputibias.n90 185
R22875 outputibias.n89 outputibias.n88 185
R22876 outputibias.n68 outputibias.n67 185
R22877 outputibias.n83 outputibias.n82 185
R22878 outputibias.n81 outputibias.n80 185
R22879 outputibias.n72 outputibias.n71 185
R22880 outputibias.n75 outputibias.n74 185
R22881 outputibias.n123 outputibias.n122 185
R22882 outputibias.n121 outputibias.n120 185
R22883 outputibias.n100 outputibias.n99 185
R22884 outputibias.n115 outputibias.n114 185
R22885 outputibias.n113 outputibias.n112 185
R22886 outputibias.n104 outputibias.n103 185
R22887 outputibias.n107 outputibias.n106 185
R22888 outputibias.n0 outputibias.t8 178.945
R22889 outputibias.n133 outputibias.t9 177.018
R22890 outputibias.n132 outputibias.t10 177.018
R22891 outputibias.n0 outputibias.t11 177.018
R22892 outputibias.t7 outputibias.n10 147.661
R22893 outputibias.t5 outputibias.n41 147.661
R22894 outputibias.t1 outputibias.n73 147.661
R22895 outputibias.t3 outputibias.n105 147.661
R22896 outputibias.n128 outputibias.t6 132.363
R22897 outputibias.n128 outputibias.t4 130.436
R22898 outputibias.n129 outputibias.t0 130.436
R22899 outputibias.n130 outputibias.t2 130.436
R22900 outputibias.n27 outputibias.n26 104.615
R22901 outputibias.n26 outputibias.n4 104.615
R22902 outputibias.n19 outputibias.n4 104.615
R22903 outputibias.n19 outputibias.n18 104.615
R22904 outputibias.n18 outputibias.n8 104.615
R22905 outputibias.n11 outputibias.n8 104.615
R22906 outputibias.n58 outputibias.n57 104.615
R22907 outputibias.n57 outputibias.n35 104.615
R22908 outputibias.n50 outputibias.n35 104.615
R22909 outputibias.n50 outputibias.n49 104.615
R22910 outputibias.n49 outputibias.n39 104.615
R22911 outputibias.n42 outputibias.n39 104.615
R22912 outputibias.n90 outputibias.n89 104.615
R22913 outputibias.n89 outputibias.n67 104.615
R22914 outputibias.n82 outputibias.n67 104.615
R22915 outputibias.n82 outputibias.n81 104.615
R22916 outputibias.n81 outputibias.n71 104.615
R22917 outputibias.n74 outputibias.n71 104.615
R22918 outputibias.n122 outputibias.n121 104.615
R22919 outputibias.n121 outputibias.n99 104.615
R22920 outputibias.n114 outputibias.n99 104.615
R22921 outputibias.n114 outputibias.n113 104.615
R22922 outputibias.n113 outputibias.n103 104.615
R22923 outputibias.n106 outputibias.n103 104.615
R22924 outputibias.n63 outputibias.n31 95.6354
R22925 outputibias.n63 outputibias.n62 94.6732
R22926 outputibias.n95 outputibias.n94 94.6732
R22927 outputibias.n127 outputibias.n126 94.6732
R22928 outputibias.n11 outputibias.t7 52.3082
R22929 outputibias.n42 outputibias.t5 52.3082
R22930 outputibias.n74 outputibias.t1 52.3082
R22931 outputibias.n106 outputibias.t3 52.3082
R22932 outputibias.n12 outputibias.n10 15.6674
R22933 outputibias.n43 outputibias.n41 15.6674
R22934 outputibias.n75 outputibias.n73 15.6674
R22935 outputibias.n107 outputibias.n105 15.6674
R22936 outputibias.n13 outputibias.n9 12.8005
R22937 outputibias.n44 outputibias.n40 12.8005
R22938 outputibias.n76 outputibias.n72 12.8005
R22939 outputibias.n108 outputibias.n104 12.8005
R22940 outputibias.n17 outputibias.n16 12.0247
R22941 outputibias.n48 outputibias.n47 12.0247
R22942 outputibias.n80 outputibias.n79 12.0247
R22943 outputibias.n112 outputibias.n111 12.0247
R22944 outputibias.n20 outputibias.n7 11.249
R22945 outputibias.n51 outputibias.n38 11.249
R22946 outputibias.n83 outputibias.n70 11.249
R22947 outputibias.n115 outputibias.n102 11.249
R22948 outputibias.n21 outputibias.n5 10.4732
R22949 outputibias.n52 outputibias.n36 10.4732
R22950 outputibias.n84 outputibias.n68 10.4732
R22951 outputibias.n116 outputibias.n100 10.4732
R22952 outputibias.n25 outputibias.n24 9.69747
R22953 outputibias.n56 outputibias.n55 9.69747
R22954 outputibias.n88 outputibias.n87 9.69747
R22955 outputibias.n120 outputibias.n119 9.69747
R22956 outputibias.n31 outputibias.n30 9.45567
R22957 outputibias.n62 outputibias.n61 9.45567
R22958 outputibias.n94 outputibias.n93 9.45567
R22959 outputibias.n126 outputibias.n125 9.45567
R22960 outputibias.n30 outputibias.n29 9.3005
R22961 outputibias.n3 outputibias.n2 9.3005
R22962 outputibias.n24 outputibias.n23 9.3005
R22963 outputibias.n22 outputibias.n21 9.3005
R22964 outputibias.n7 outputibias.n6 9.3005
R22965 outputibias.n16 outputibias.n15 9.3005
R22966 outputibias.n14 outputibias.n13 9.3005
R22967 outputibias.n61 outputibias.n60 9.3005
R22968 outputibias.n34 outputibias.n33 9.3005
R22969 outputibias.n55 outputibias.n54 9.3005
R22970 outputibias.n53 outputibias.n52 9.3005
R22971 outputibias.n38 outputibias.n37 9.3005
R22972 outputibias.n47 outputibias.n46 9.3005
R22973 outputibias.n45 outputibias.n44 9.3005
R22974 outputibias.n93 outputibias.n92 9.3005
R22975 outputibias.n66 outputibias.n65 9.3005
R22976 outputibias.n87 outputibias.n86 9.3005
R22977 outputibias.n85 outputibias.n84 9.3005
R22978 outputibias.n70 outputibias.n69 9.3005
R22979 outputibias.n79 outputibias.n78 9.3005
R22980 outputibias.n77 outputibias.n76 9.3005
R22981 outputibias.n125 outputibias.n124 9.3005
R22982 outputibias.n98 outputibias.n97 9.3005
R22983 outputibias.n119 outputibias.n118 9.3005
R22984 outputibias.n117 outputibias.n116 9.3005
R22985 outputibias.n102 outputibias.n101 9.3005
R22986 outputibias.n111 outputibias.n110 9.3005
R22987 outputibias.n109 outputibias.n108 9.3005
R22988 outputibias.n28 outputibias.n3 8.92171
R22989 outputibias.n59 outputibias.n34 8.92171
R22990 outputibias.n91 outputibias.n66 8.92171
R22991 outputibias.n123 outputibias.n98 8.92171
R22992 outputibias.n29 outputibias.n1 8.14595
R22993 outputibias.n60 outputibias.n32 8.14595
R22994 outputibias.n92 outputibias.n64 8.14595
R22995 outputibias.n124 outputibias.n96 8.14595
R22996 outputibias.n31 outputibias.n1 5.81868
R22997 outputibias.n62 outputibias.n32 5.81868
R22998 outputibias.n94 outputibias.n64 5.81868
R22999 outputibias.n126 outputibias.n96 5.81868
R23000 outputibias.n131 outputibias.n130 5.20947
R23001 outputibias.n29 outputibias.n28 5.04292
R23002 outputibias.n60 outputibias.n59 5.04292
R23003 outputibias.n92 outputibias.n91 5.04292
R23004 outputibias.n124 outputibias.n123 5.04292
R23005 outputibias.n131 outputibias.n127 4.42209
R23006 outputibias.n14 outputibias.n10 4.38594
R23007 outputibias.n45 outputibias.n41 4.38594
R23008 outputibias.n77 outputibias.n73 4.38594
R23009 outputibias.n109 outputibias.n105 4.38594
R23010 outputibias.n132 outputibias.n131 4.28454
R23011 outputibias.n25 outputibias.n3 4.26717
R23012 outputibias.n56 outputibias.n34 4.26717
R23013 outputibias.n88 outputibias.n66 4.26717
R23014 outputibias.n120 outputibias.n98 4.26717
R23015 outputibias.n24 outputibias.n5 3.49141
R23016 outputibias.n55 outputibias.n36 3.49141
R23017 outputibias.n87 outputibias.n68 3.49141
R23018 outputibias.n119 outputibias.n100 3.49141
R23019 outputibias.n21 outputibias.n20 2.71565
R23020 outputibias.n52 outputibias.n51 2.71565
R23021 outputibias.n84 outputibias.n83 2.71565
R23022 outputibias.n116 outputibias.n115 2.71565
R23023 outputibias.n17 outputibias.n7 1.93989
R23024 outputibias.n48 outputibias.n38 1.93989
R23025 outputibias.n80 outputibias.n70 1.93989
R23026 outputibias.n112 outputibias.n102 1.93989
R23027 outputibias.n130 outputibias.n129 1.9266
R23028 outputibias.n129 outputibias.n128 1.9266
R23029 outputibias.n133 outputibias.n132 1.92658
R23030 outputibias.n134 outputibias.n133 1.29913
R23031 outputibias.n16 outputibias.n9 1.16414
R23032 outputibias.n47 outputibias.n40 1.16414
R23033 outputibias.n79 outputibias.n72 1.16414
R23034 outputibias.n111 outputibias.n104 1.16414
R23035 outputibias.n127 outputibias.n95 0.962709
R23036 outputibias.n95 outputibias.n63 0.962709
R23037 outputibias.n13 outputibias.n12 0.388379
R23038 outputibias.n44 outputibias.n43 0.388379
R23039 outputibias.n76 outputibias.n75 0.388379
R23040 outputibias.n108 outputibias.n107 0.388379
R23041 outputibias.n134 outputibias.n0 0.337251
R23042 outputibias outputibias.n134 0.302375
R23043 outputibias.n30 outputibias.n2 0.155672
R23044 outputibias.n23 outputibias.n2 0.155672
R23045 outputibias.n23 outputibias.n22 0.155672
R23046 outputibias.n22 outputibias.n6 0.155672
R23047 outputibias.n15 outputibias.n6 0.155672
R23048 outputibias.n15 outputibias.n14 0.155672
R23049 outputibias.n61 outputibias.n33 0.155672
R23050 outputibias.n54 outputibias.n33 0.155672
R23051 outputibias.n54 outputibias.n53 0.155672
R23052 outputibias.n53 outputibias.n37 0.155672
R23053 outputibias.n46 outputibias.n37 0.155672
R23054 outputibias.n46 outputibias.n45 0.155672
R23055 outputibias.n93 outputibias.n65 0.155672
R23056 outputibias.n86 outputibias.n65 0.155672
R23057 outputibias.n86 outputibias.n85 0.155672
R23058 outputibias.n85 outputibias.n69 0.155672
R23059 outputibias.n78 outputibias.n69 0.155672
R23060 outputibias.n78 outputibias.n77 0.155672
R23061 outputibias.n125 outputibias.n97 0.155672
R23062 outputibias.n118 outputibias.n97 0.155672
R23063 outputibias.n118 outputibias.n117 0.155672
R23064 outputibias.n117 outputibias.n101 0.155672
R23065 outputibias.n110 outputibias.n101 0.155672
R23066 outputibias.n110 outputibias.n109 0.155672
R23067 diffpairibias.n0 diffpairibias.t18 436.822
R23068 diffpairibias.n21 diffpairibias.t19 435.479
R23069 diffpairibias.n20 diffpairibias.t16 435.479
R23070 diffpairibias.n19 diffpairibias.t17 435.479
R23071 diffpairibias.n18 diffpairibias.t21 435.479
R23072 diffpairibias.n0 diffpairibias.t22 435.479
R23073 diffpairibias.n1 diffpairibias.t20 435.479
R23074 diffpairibias.n2 diffpairibias.t23 435.479
R23075 diffpairibias.n10 diffpairibias.t0 377.536
R23076 diffpairibias.n10 diffpairibias.t8 376.193
R23077 diffpairibias.n11 diffpairibias.t10 376.193
R23078 diffpairibias.n12 diffpairibias.t6 376.193
R23079 diffpairibias.n13 diffpairibias.t2 376.193
R23080 diffpairibias.n14 diffpairibias.t12 376.193
R23081 diffpairibias.n15 diffpairibias.t4 376.193
R23082 diffpairibias.n16 diffpairibias.t14 376.193
R23083 diffpairibias.n3 diffpairibias.t1 113.368
R23084 diffpairibias.n3 diffpairibias.t9 112.698
R23085 diffpairibias.n4 diffpairibias.t11 112.698
R23086 diffpairibias.n5 diffpairibias.t7 112.698
R23087 diffpairibias.n6 diffpairibias.t3 112.698
R23088 diffpairibias.n7 diffpairibias.t13 112.698
R23089 diffpairibias.n8 diffpairibias.t5 112.698
R23090 diffpairibias.n9 diffpairibias.t15 112.698
R23091 diffpairibias.n17 diffpairibias.n16 4.77242
R23092 diffpairibias.n17 diffpairibias.n9 4.30807
R23093 diffpairibias.n18 diffpairibias.n17 4.13945
R23094 diffpairibias.n16 diffpairibias.n15 1.34352
R23095 diffpairibias.n15 diffpairibias.n14 1.34352
R23096 diffpairibias.n14 diffpairibias.n13 1.34352
R23097 diffpairibias.n13 diffpairibias.n12 1.34352
R23098 diffpairibias.n12 diffpairibias.n11 1.34352
R23099 diffpairibias.n11 diffpairibias.n10 1.34352
R23100 diffpairibias.n2 diffpairibias.n1 1.34352
R23101 diffpairibias.n1 diffpairibias.n0 1.34352
R23102 diffpairibias.n19 diffpairibias.n18 1.34352
R23103 diffpairibias.n20 diffpairibias.n19 1.34352
R23104 diffpairibias.n21 diffpairibias.n20 1.34352
R23105 diffpairibias.n22 diffpairibias.n21 0.862419
R23106 diffpairibias diffpairibias.n22 0.684875
R23107 diffpairibias.n9 diffpairibias.n8 0.672012
R23108 diffpairibias.n8 diffpairibias.n7 0.672012
R23109 diffpairibias.n7 diffpairibias.n6 0.672012
R23110 diffpairibias.n6 diffpairibias.n5 0.672012
R23111 diffpairibias.n5 diffpairibias.n4 0.672012
R23112 diffpairibias.n4 diffpairibias.n3 0.672012
R23113 diffpairibias.n22 diffpairibias.n2 0.190907
C0 output outputibias 2.34152f
C1 vdd output 7.23429f
C2 CSoutput output 6.13571f
C3 CSoutput outputibias 0.032386f
C4 vdd CSoutput 0.140606p
C5 commonsourceibias output 0.006808f
C6 minus diffpairibias 3.4e-19
C7 CSoutput minus 2.76215f
C8 vdd plus 0.089709f
C9 plus diffpairibias 3.42e-19
C10 commonsourceibias outputibias 0.003832f
C11 vdd commonsourceibias 0.004218f
C12 CSoutput plus 0.858911f
C13 commonsourceibias diffpairibias 0.052851f
C14 CSoutput commonsourceibias 36.982002f
C15 minus plus 9.225019f
C16 minus commonsourceibias 0.323913f
C17 plus commonsourceibias 0.278362f
C18 diffpairibias gnd 48.96854f
C19 outputibias gnd 32.465668f
C20 output gnd 15.47879f
C21 commonsourceibias gnd 0.150128p
C22 plus gnd 33.516796f
C23 minus gnd 27.657059f
C24 CSoutput gnd 0.10126p
C25 vdd gnd 0.439524p
C26 diffpairibias.t18 gnd 0.087401f
C27 diffpairibias.t22 gnd 0.087239f
C28 diffpairibias.n0 gnd 0.102784f
C29 diffpairibias.t20 gnd 0.087239f
C30 diffpairibias.n1 gnd 0.050171f
C31 diffpairibias.t23 gnd 0.087239f
C32 diffpairibias.n2 gnd 0.039841f
C33 diffpairibias.t1 gnd 0.083757f
C34 diffpairibias.t9 gnd 0.083392f
C35 diffpairibias.n3 gnd 0.131682f
C36 diffpairibias.t11 gnd 0.083392f
C37 diffpairibias.n4 gnd 0.07027f
C38 diffpairibias.t7 gnd 0.083392f
C39 diffpairibias.n5 gnd 0.07027f
C40 diffpairibias.t3 gnd 0.083392f
C41 diffpairibias.n6 gnd 0.07027f
C42 diffpairibias.t13 gnd 0.083392f
C43 diffpairibias.n7 gnd 0.07027f
C44 diffpairibias.t5 gnd 0.083392f
C45 diffpairibias.n8 gnd 0.07027f
C46 diffpairibias.t15 gnd 0.083392f
C47 diffpairibias.n9 gnd 0.099771f
C48 diffpairibias.t0 gnd 0.08427f
C49 diffpairibias.t8 gnd 0.084123f
C50 diffpairibias.n10 gnd 0.091784f
C51 diffpairibias.t10 gnd 0.084123f
C52 diffpairibias.n11 gnd 0.050681f
C53 diffpairibias.t6 gnd 0.084123f
C54 diffpairibias.n12 gnd 0.050681f
C55 diffpairibias.t2 gnd 0.084123f
C56 diffpairibias.n13 gnd 0.050681f
C57 diffpairibias.t12 gnd 0.084123f
C58 diffpairibias.n14 gnd 0.050681f
C59 diffpairibias.t4 gnd 0.084123f
C60 diffpairibias.n15 gnd 0.050681f
C61 diffpairibias.t14 gnd 0.084123f
C62 diffpairibias.n16 gnd 0.059977f
C63 diffpairibias.n17 gnd 0.226448f
C64 diffpairibias.t21 gnd 0.087239f
C65 diffpairibias.n18 gnd 0.050181f
C66 diffpairibias.t17 gnd 0.087239f
C67 diffpairibias.n19 gnd 0.050171f
C68 diffpairibias.t16 gnd 0.087239f
C69 diffpairibias.n20 gnd 0.050171f
C70 diffpairibias.t19 gnd 0.087239f
C71 diffpairibias.n21 gnd 0.045859f
C72 diffpairibias.n22 gnd 0.046268f
C73 outputibias.t11 gnd 0.11477f
C74 outputibias.t8 gnd 0.115567f
C75 outputibias.n0 gnd 0.130108f
C76 outputibias.n1 gnd 0.001372f
C77 outputibias.n2 gnd 9.76e-19
C78 outputibias.n3 gnd 5.24e-19
C79 outputibias.n4 gnd 0.001239f
C80 outputibias.n5 gnd 5.55e-19
C81 outputibias.n6 gnd 9.76e-19
C82 outputibias.n7 gnd 5.24e-19
C83 outputibias.n8 gnd 0.001239f
C84 outputibias.n9 gnd 5.55e-19
C85 outputibias.n10 gnd 0.004176f
C86 outputibias.t7 gnd 0.00202f
C87 outputibias.n11 gnd 9.3e-19
C88 outputibias.n12 gnd 7.32e-19
C89 outputibias.n13 gnd 5.24e-19
C90 outputibias.n14 gnd 0.02322f
C91 outputibias.n15 gnd 9.76e-19
C92 outputibias.n16 gnd 5.24e-19
C93 outputibias.n17 gnd 5.55e-19
C94 outputibias.n18 gnd 0.001239f
C95 outputibias.n19 gnd 0.001239f
C96 outputibias.n20 gnd 5.55e-19
C97 outputibias.n21 gnd 5.24e-19
C98 outputibias.n22 gnd 9.76e-19
C99 outputibias.n23 gnd 9.76e-19
C100 outputibias.n24 gnd 5.24e-19
C101 outputibias.n25 gnd 5.55e-19
C102 outputibias.n26 gnd 0.001239f
C103 outputibias.n27 gnd 0.002683f
C104 outputibias.n28 gnd 5.55e-19
C105 outputibias.n29 gnd 5.24e-19
C106 outputibias.n30 gnd 0.002256f
C107 outputibias.n31 gnd 0.005781f
C108 outputibias.n32 gnd 0.001372f
C109 outputibias.n33 gnd 9.76e-19
C110 outputibias.n34 gnd 5.24e-19
C111 outputibias.n35 gnd 0.001239f
C112 outputibias.n36 gnd 5.55e-19
C113 outputibias.n37 gnd 9.76e-19
C114 outputibias.n38 gnd 5.24e-19
C115 outputibias.n39 gnd 0.001239f
C116 outputibias.n40 gnd 5.55e-19
C117 outputibias.n41 gnd 0.004176f
C118 outputibias.t5 gnd 0.00202f
C119 outputibias.n42 gnd 9.3e-19
C120 outputibias.n43 gnd 7.32e-19
C121 outputibias.n44 gnd 5.24e-19
C122 outputibias.n45 gnd 0.02322f
C123 outputibias.n46 gnd 9.76e-19
C124 outputibias.n47 gnd 5.24e-19
C125 outputibias.n48 gnd 5.55e-19
C126 outputibias.n49 gnd 0.001239f
C127 outputibias.n50 gnd 0.001239f
C128 outputibias.n51 gnd 5.55e-19
C129 outputibias.n52 gnd 5.24e-19
C130 outputibias.n53 gnd 9.76e-19
C131 outputibias.n54 gnd 9.76e-19
C132 outputibias.n55 gnd 5.24e-19
C133 outputibias.n56 gnd 5.55e-19
C134 outputibias.n57 gnd 0.001239f
C135 outputibias.n58 gnd 0.002683f
C136 outputibias.n59 gnd 5.55e-19
C137 outputibias.n60 gnd 5.24e-19
C138 outputibias.n61 gnd 0.002256f
C139 outputibias.n62 gnd 0.005197f
C140 outputibias.n63 gnd 0.121892f
C141 outputibias.n64 gnd 0.001372f
C142 outputibias.n65 gnd 9.76e-19
C143 outputibias.n66 gnd 5.24e-19
C144 outputibias.n67 gnd 0.001239f
C145 outputibias.n68 gnd 5.55e-19
C146 outputibias.n69 gnd 9.76e-19
C147 outputibias.n70 gnd 5.24e-19
C148 outputibias.n71 gnd 0.001239f
C149 outputibias.n72 gnd 5.55e-19
C150 outputibias.n73 gnd 0.004176f
C151 outputibias.t1 gnd 0.00202f
C152 outputibias.n74 gnd 9.3e-19
C153 outputibias.n75 gnd 7.32e-19
C154 outputibias.n76 gnd 5.24e-19
C155 outputibias.n77 gnd 0.02322f
C156 outputibias.n78 gnd 9.76e-19
C157 outputibias.n79 gnd 5.24e-19
C158 outputibias.n80 gnd 5.55e-19
C159 outputibias.n81 gnd 0.001239f
C160 outputibias.n82 gnd 0.001239f
C161 outputibias.n83 gnd 5.55e-19
C162 outputibias.n84 gnd 5.24e-19
C163 outputibias.n85 gnd 9.76e-19
C164 outputibias.n86 gnd 9.76e-19
C165 outputibias.n87 gnd 5.24e-19
C166 outputibias.n88 gnd 5.55e-19
C167 outputibias.n89 gnd 0.001239f
C168 outputibias.n90 gnd 0.002683f
C169 outputibias.n91 gnd 5.55e-19
C170 outputibias.n92 gnd 5.24e-19
C171 outputibias.n93 gnd 0.002256f
C172 outputibias.n94 gnd 0.005197f
C173 outputibias.n95 gnd 0.064513f
C174 outputibias.n96 gnd 0.001372f
C175 outputibias.n97 gnd 9.76e-19
C176 outputibias.n98 gnd 5.24e-19
C177 outputibias.n99 gnd 0.001239f
C178 outputibias.n100 gnd 5.55e-19
C179 outputibias.n101 gnd 9.76e-19
C180 outputibias.n102 gnd 5.24e-19
C181 outputibias.n103 gnd 0.001239f
C182 outputibias.n104 gnd 5.55e-19
C183 outputibias.n105 gnd 0.004176f
C184 outputibias.t3 gnd 0.00202f
C185 outputibias.n106 gnd 9.3e-19
C186 outputibias.n107 gnd 7.32e-19
C187 outputibias.n108 gnd 5.24e-19
C188 outputibias.n109 gnd 0.02322f
C189 outputibias.n110 gnd 9.76e-19
C190 outputibias.n111 gnd 5.24e-19
C191 outputibias.n112 gnd 5.55e-19
C192 outputibias.n113 gnd 0.001239f
C193 outputibias.n114 gnd 0.001239f
C194 outputibias.n115 gnd 5.55e-19
C195 outputibias.n116 gnd 5.24e-19
C196 outputibias.n117 gnd 9.76e-19
C197 outputibias.n118 gnd 9.76e-19
C198 outputibias.n119 gnd 5.24e-19
C199 outputibias.n120 gnd 5.55e-19
C200 outputibias.n121 gnd 0.001239f
C201 outputibias.n122 gnd 0.002683f
C202 outputibias.n123 gnd 5.55e-19
C203 outputibias.n124 gnd 5.24e-19
C204 outputibias.n125 gnd 0.002256f
C205 outputibias.n126 gnd 0.005197f
C206 outputibias.n127 gnd 0.084814f
C207 outputibias.t2 gnd 0.108319f
C208 outputibias.t0 gnd 0.108319f
C209 outputibias.t4 gnd 0.108319f
C210 outputibias.t6 gnd 0.109238f
C211 outputibias.n128 gnd 0.134674f
C212 outputibias.n129 gnd 0.07244f
C213 outputibias.n130 gnd 0.079818f
C214 outputibias.n131 gnd 0.164901f
C215 outputibias.t10 gnd 0.11477f
C216 outputibias.n132 gnd 0.067481f
C217 outputibias.t9 gnd 0.11477f
C218 outputibias.n133 gnd 0.065115f
C219 outputibias.n134 gnd 0.029159f
C220 output.t13 gnd 0.464308f
C221 output.t3 gnd 0.044422f
C222 output.t8 gnd 0.044422f
C223 output.n0 gnd 0.364624f
C224 output.n1 gnd 0.614102f
C225 output.t12 gnd 0.044422f
C226 output.t4 gnd 0.044422f
C227 output.n2 gnd 0.364624f
C228 output.n3 gnd 0.350265f
C229 output.t6 gnd 0.044422f
C230 output.t5 gnd 0.044422f
C231 output.n4 gnd 0.364624f
C232 output.n5 gnd 0.350265f
C233 output.t11 gnd 0.044422f
C234 output.t14 gnd 0.044422f
C235 output.n6 gnd 0.364624f
C236 output.n7 gnd 0.350265f
C237 output.t16 gnd 0.044422f
C238 output.t9 gnd 0.044422f
C239 output.n8 gnd 0.364624f
C240 output.n9 gnd 0.350265f
C241 output.t10 gnd 0.044422f
C242 output.t17 gnd 0.044422f
C243 output.n10 gnd 0.364624f
C244 output.n11 gnd 0.350265f
C245 output.t2 gnd 0.044422f
C246 output.t7 gnd 0.044422f
C247 output.n12 gnd 0.364624f
C248 output.n13 gnd 0.350265f
C249 output.t15 gnd 0.462979f
C250 output.n14 gnd 0.28994f
C251 output.n15 gnd 0.015803f
C252 output.n16 gnd 0.011243f
C253 output.n17 gnd 0.006041f
C254 output.n18 gnd 0.01428f
C255 output.n19 gnd 0.006397f
C256 output.n20 gnd 0.011243f
C257 output.n21 gnd 0.006041f
C258 output.n22 gnd 0.01428f
C259 output.n23 gnd 0.006397f
C260 output.n24 gnd 0.048111f
C261 output.t0 gnd 0.023274f
C262 output.n25 gnd 0.01071f
C263 output.n26 gnd 0.008435f
C264 output.n27 gnd 0.006041f
C265 output.n28 gnd 0.267512f
C266 output.n29 gnd 0.011243f
C267 output.n30 gnd 0.006041f
C268 output.n31 gnd 0.006397f
C269 output.n32 gnd 0.01428f
C270 output.n33 gnd 0.01428f
C271 output.n34 gnd 0.006397f
C272 output.n35 gnd 0.006041f
C273 output.n36 gnd 0.011243f
C274 output.n37 gnd 0.011243f
C275 output.n38 gnd 0.006041f
C276 output.n39 gnd 0.006397f
C277 output.n40 gnd 0.01428f
C278 output.n41 gnd 0.030913f
C279 output.n42 gnd 0.006397f
C280 output.n43 gnd 0.006041f
C281 output.n44 gnd 0.025987f
C282 output.n45 gnd 0.097665f
C283 output.n46 gnd 0.015803f
C284 output.n47 gnd 0.011243f
C285 output.n48 gnd 0.006041f
C286 output.n49 gnd 0.01428f
C287 output.n50 gnd 0.006397f
C288 output.n51 gnd 0.011243f
C289 output.n52 gnd 0.006041f
C290 output.n53 gnd 0.01428f
C291 output.n54 gnd 0.006397f
C292 output.n55 gnd 0.048111f
C293 output.t18 gnd 0.023274f
C294 output.n56 gnd 0.01071f
C295 output.n57 gnd 0.008435f
C296 output.n58 gnd 0.006041f
C297 output.n59 gnd 0.267512f
C298 output.n60 gnd 0.011243f
C299 output.n61 gnd 0.006041f
C300 output.n62 gnd 0.006397f
C301 output.n63 gnd 0.01428f
C302 output.n64 gnd 0.01428f
C303 output.n65 gnd 0.006397f
C304 output.n66 gnd 0.006041f
C305 output.n67 gnd 0.011243f
C306 output.n68 gnd 0.011243f
C307 output.n69 gnd 0.006041f
C308 output.n70 gnd 0.006397f
C309 output.n71 gnd 0.01428f
C310 output.n72 gnd 0.030913f
C311 output.n73 gnd 0.006397f
C312 output.n74 gnd 0.006041f
C313 output.n75 gnd 0.025987f
C314 output.n76 gnd 0.09306f
C315 output.n77 gnd 1.65264f
C316 output.n78 gnd 0.015803f
C317 output.n79 gnd 0.011243f
C318 output.n80 gnd 0.006041f
C319 output.n81 gnd 0.01428f
C320 output.n82 gnd 0.006397f
C321 output.n83 gnd 0.011243f
C322 output.n84 gnd 0.006041f
C323 output.n85 gnd 0.01428f
C324 output.n86 gnd 0.006397f
C325 output.n87 gnd 0.048111f
C326 output.t1 gnd 0.023274f
C327 output.n88 gnd 0.01071f
C328 output.n89 gnd 0.008435f
C329 output.n90 gnd 0.006041f
C330 output.n91 gnd 0.267512f
C331 output.n92 gnd 0.011243f
C332 output.n93 gnd 0.006041f
C333 output.n94 gnd 0.006397f
C334 output.n95 gnd 0.01428f
C335 output.n96 gnd 0.01428f
C336 output.n97 gnd 0.006397f
C337 output.n98 gnd 0.006041f
C338 output.n99 gnd 0.011243f
C339 output.n100 gnd 0.011243f
C340 output.n101 gnd 0.006041f
C341 output.n102 gnd 0.006397f
C342 output.n103 gnd 0.01428f
C343 output.n104 gnd 0.030913f
C344 output.n105 gnd 0.006397f
C345 output.n106 gnd 0.006041f
C346 output.n107 gnd 0.025987f
C347 output.n108 gnd 0.09306f
C348 output.n109 gnd 0.713089f
C349 output.n110 gnd 0.015803f
C350 output.n111 gnd 0.011243f
C351 output.n112 gnd 0.006041f
C352 output.n113 gnd 0.01428f
C353 output.n114 gnd 0.006397f
C354 output.n115 gnd 0.011243f
C355 output.n116 gnd 0.006041f
C356 output.n117 gnd 0.01428f
C357 output.n118 gnd 0.006397f
C358 output.n119 gnd 0.048111f
C359 output.t19 gnd 0.023274f
C360 output.n120 gnd 0.01071f
C361 output.n121 gnd 0.008435f
C362 output.n122 gnd 0.006041f
C363 output.n123 gnd 0.267512f
C364 output.n124 gnd 0.011243f
C365 output.n125 gnd 0.006041f
C366 output.n126 gnd 0.006397f
C367 output.n127 gnd 0.01428f
C368 output.n128 gnd 0.01428f
C369 output.n129 gnd 0.006397f
C370 output.n130 gnd 0.006041f
C371 output.n131 gnd 0.011243f
C372 output.n132 gnd 0.011243f
C373 output.n133 gnd 0.006041f
C374 output.n134 gnd 0.006397f
C375 output.n135 gnd 0.01428f
C376 output.n136 gnd 0.030913f
C377 output.n137 gnd 0.006397f
C378 output.n138 gnd 0.006041f
C379 output.n139 gnd 0.025987f
C380 output.n140 gnd 0.09306f
C381 output.n141 gnd 1.67353f
C382 minus.n0 gnd 0.031753f
C383 minus.n1 gnd 0.007205f
C384 minus.n2 gnd 0.031753f
C385 minus.n3 gnd 0.007205f
C386 minus.n4 gnd 0.031753f
C387 minus.n5 gnd 0.007205f
C388 minus.n6 gnd 0.031753f
C389 minus.n7 gnd 0.007205f
C390 minus.t8 gnd 0.464846f
C391 minus.t7 gnd 0.449112f
C392 minus.n8 gnd 0.204821f
C393 minus.n9 gnd 0.186055f
C394 minus.n10 gnd 0.135533f
C395 minus.n11 gnd 0.031753f
C396 minus.t11 gnd 0.449112f
C397 minus.n12 gnd 0.19951f
C398 minus.n13 gnd 0.007205f
C399 minus.t10 gnd 0.449112f
C400 minus.n14 gnd 0.19951f
C401 minus.n15 gnd 0.031753f
C402 minus.n16 gnd 0.031753f
C403 minus.n17 gnd 0.031753f
C404 minus.t12 gnd 0.449112f
C405 minus.n18 gnd 0.19951f
C406 minus.n19 gnd 0.007205f
C407 minus.t17 gnd 0.449112f
C408 minus.n20 gnd 0.19951f
C409 minus.n21 gnd 0.031753f
C410 minus.n22 gnd 0.031753f
C411 minus.n23 gnd 0.031753f
C412 minus.t16 gnd 0.449112f
C413 minus.n24 gnd 0.19951f
C414 minus.n25 gnd 0.007205f
C415 minus.t21 gnd 0.449112f
C416 minus.n26 gnd 0.19951f
C417 minus.n27 gnd 0.031753f
C418 minus.n28 gnd 0.031753f
C419 minus.n29 gnd 0.031753f
C420 minus.t20 gnd 0.449112f
C421 minus.n30 gnd 0.19951f
C422 minus.n31 gnd 0.007205f
C423 minus.t13 gnd 0.449112f
C424 minus.n32 gnd 0.199216f
C425 minus.n33 gnd 0.366878f
C426 minus.n34 gnd 0.031753f
C427 minus.t5 gnd 0.449112f
C428 minus.t6 gnd 0.449112f
C429 minus.n35 gnd 0.031753f
C430 minus.t22 gnd 0.449112f
C431 minus.n36 gnd 0.19951f
C432 minus.n37 gnd 0.031753f
C433 minus.t18 gnd 0.449112f
C434 minus.t19 gnd 0.449112f
C435 minus.n38 gnd 0.19951f
C436 minus.n39 gnd 0.031753f
C437 minus.t14 gnd 0.449112f
C438 minus.t15 gnd 0.449112f
C439 minus.n40 gnd 0.19951f
C440 minus.n41 gnd 0.031753f
C441 minus.t9 gnd 0.449112f
C442 minus.t23 gnd 0.449112f
C443 minus.n42 gnd 0.204821f
C444 minus.t24 gnd 0.464846f
C445 minus.n43 gnd 0.186055f
C446 minus.n44 gnd 0.135533f
C447 minus.n45 gnd 0.007205f
C448 minus.n46 gnd 0.19951f
C449 minus.n47 gnd 0.007205f
C450 minus.n48 gnd 0.031753f
C451 minus.n49 gnd 0.031753f
C452 minus.n50 gnd 0.031753f
C453 minus.n51 gnd 0.007205f
C454 minus.n52 gnd 0.19951f
C455 minus.n53 gnd 0.007205f
C456 minus.n54 gnd 0.031753f
C457 minus.n55 gnd 0.031753f
C458 minus.n56 gnd 0.031753f
C459 minus.n57 gnd 0.007205f
C460 minus.n58 gnd 0.19951f
C461 minus.n59 gnd 0.007205f
C462 minus.n60 gnd 0.031753f
C463 minus.n61 gnd 0.031753f
C464 minus.n62 gnd 0.031753f
C465 minus.n63 gnd 0.007205f
C466 minus.n64 gnd 0.19951f
C467 minus.n65 gnd 0.007205f
C468 minus.n66 gnd 0.199216f
C469 minus.n67 gnd 0.992181f
C470 minus.n68 gnd 1.49371f
C471 minus.t2 gnd 0.009788f
C472 minus.t0 gnd 0.009788f
C473 minus.n69 gnd 0.032187f
C474 minus.t3 gnd 0.009788f
C475 minus.t1 gnd 0.009788f
C476 minus.n70 gnd 0.031746f
C477 minus.n71 gnd 0.270934f
C478 minus.t4 gnd 0.054481f
C479 minus.n72 gnd 0.147846f
C480 minus.n73 gnd 1.99457f
C481 a_n1986_8322.t20 gnd 49.3562f
C482 a_n1986_8322.t21 gnd 75.4844f
C483 a_n1986_8322.t2 gnd 0.093529f
C484 a_n1986_8322.t1 gnd 0.875761f
C485 a_n1986_8322.t9 gnd 0.093529f
C486 a_n1986_8322.t4 gnd 0.093529f
C487 a_n1986_8322.n0 gnd 0.65882f
C488 a_n1986_8322.n1 gnd 0.736135f
C489 a_n1986_8322.t7 gnd 0.093529f
C490 a_n1986_8322.t6 gnd 0.093529f
C491 a_n1986_8322.n2 gnd 0.65882f
C492 a_n1986_8322.n3 gnd 0.374021f
C493 a_n1986_8322.t0 gnd 0.874017f
C494 a_n1986_8322.n4 gnd 1.39891f
C495 a_n1986_8322.t15 gnd 0.875761f
C496 a_n1986_8322.t19 gnd 0.093529f
C497 a_n1986_8322.t18 gnd 0.093529f
C498 a_n1986_8322.n5 gnd 0.65882f
C499 a_n1986_8322.n6 gnd 0.736135f
C500 a_n1986_8322.t13 gnd 0.874017f
C501 a_n1986_8322.n7 gnd 0.370433f
C502 a_n1986_8322.t16 gnd 0.874017f
C503 a_n1986_8322.n8 gnd 0.370433f
C504 a_n1986_8322.t14 gnd 0.093529f
C505 a_n1986_8322.t12 gnd 0.093529f
C506 a_n1986_8322.n9 gnd 0.65882f
C507 a_n1986_8322.n10 gnd 0.374021f
C508 a_n1986_8322.t17 gnd 0.874017f
C509 a_n1986_8322.n11 gnd 0.872286f
C510 a_n1986_8322.n12 gnd 1.59065f
C511 a_n1986_8322.n13 gnd 3.48702f
C512 a_n1986_8322.t3 gnd 0.874017f
C513 a_n1986_8322.n14 gnd 0.766493f
C514 a_n1986_8322.t10 gnd 0.875759f
C515 a_n1986_8322.t8 gnd 0.093529f
C516 a_n1986_8322.t5 gnd 0.093529f
C517 a_n1986_8322.n15 gnd 0.65882f
C518 a_n1986_8322.n16 gnd 0.736137f
C519 a_n1986_8322.n17 gnd 0.374019f
C520 a_n1986_8322.n18 gnd 0.658822f
C521 a_n1986_8322.t11 gnd 0.093529f
C522 a_n1808_13878.t7 gnd 0.185195f
C523 a_n1808_13878.t2 gnd 0.185195f
C524 a_n1808_13878.t4 gnd 0.185195f
C525 a_n1808_13878.n0 gnd 1.4598f
C526 a_n1808_13878.t8 gnd 0.185195f
C527 a_n1808_13878.t3 gnd 0.185195f
C528 a_n1808_13878.n1 gnd 1.45825f
C529 a_n1808_13878.n2 gnd 2.03762f
C530 a_n1808_13878.t6 gnd 0.185195f
C531 a_n1808_13878.t1 gnd 0.185195f
C532 a_n1808_13878.n3 gnd 1.45825f
C533 a_n1808_13878.n4 gnd 3.69301f
C534 a_n1808_13878.t13 gnd 1.73408f
C535 a_n1808_13878.t16 gnd 0.185195f
C536 a_n1808_13878.t17 gnd 0.185195f
C537 a_n1808_13878.n5 gnd 1.30452f
C538 a_n1808_13878.n6 gnd 1.4576f
C539 a_n1808_13878.t12 gnd 1.73062f
C540 a_n1808_13878.n7 gnd 0.733487f
C541 a_n1808_13878.t15 gnd 1.73062f
C542 a_n1808_13878.n8 gnd 0.733487f
C543 a_n1808_13878.t18 gnd 0.185195f
C544 a_n1808_13878.t19 gnd 0.185195f
C545 a_n1808_13878.n9 gnd 1.30452f
C546 a_n1808_13878.n10 gnd 0.74059f
C547 a_n1808_13878.t14 gnd 1.73062f
C548 a_n1808_13878.n11 gnd 1.7272f
C549 a_n1808_13878.n12 gnd 2.51438f
C550 a_n1808_13878.t9 gnd 0.185195f
C551 a_n1808_13878.t10 gnd 0.185195f
C552 a_n1808_13878.n13 gnd 1.45825f
C553 a_n1808_13878.n14 gnd 1.80025f
C554 a_n1808_13878.t0 gnd 0.185195f
C555 a_n1808_13878.t5 gnd 0.185195f
C556 a_n1808_13878.n15 gnd 1.45825f
C557 a_n1808_13878.n16 gnd 1.31079f
C558 a_n1808_13878.n17 gnd 1.46067f
C559 a_n1808_13878.t11 gnd 0.185195f
C560 a_n1996_n452.n0 gnd 0.822727f
C561 a_n1996_n452.n1 gnd 3.34433f
C562 a_n1996_n452.n2 gnd 3.17111f
C563 a_n1996_n452.n3 gnd 3.91594f
C564 a_n1996_n452.n4 gnd 0.527811f
C565 a_n1996_n452.n5 gnd 0.205584f
C566 a_n1996_n452.n6 gnd 0.151417f
C567 a_n1996_n452.n7 gnd 0.237979f
C568 a_n1996_n452.n8 gnd 0.183812f
C569 a_n1996_n452.n9 gnd 0.205584f
C570 a_n1996_n452.n10 gnd 1.00969f
C571 a_n1996_n452.n11 gnd 0.151417f
C572 a_n1996_n452.n12 gnd 0.581979f
C573 a_n1996_n452.n13 gnd 0.433746f
C574 a_n1996_n452.n14 gnd 0.21667f
C575 a_n1996_n452.n15 gnd 0.494132f
C576 a_n1996_n452.n16 gnd 0.283464f
C577 a_n1996_n452.n17 gnd 0.439964f
C578 a_n1996_n452.n18 gnd 0.21667f
C579 a_n1996_n452.n19 gnd 0.734001f
C580 a_n1996_n452.n20 gnd 0.283464f
C581 a_n1996_n452.n21 gnd 0.494132f
C582 a_n1996_n452.n22 gnd 0.666675f
C583 a_n1996_n452.n23 gnd 0.21667f
C584 a_n1996_n452.n24 gnd 0.283464f
C585 a_n1996_n452.n25 gnd 0.641354f
C586 a_n1996_n452.n26 gnd 0.283464f
C587 a_n1996_n452.n27 gnd 1.18284f
C588 a_n1996_n452.n28 gnd 1.92214f
C589 a_n1996_n452.n29 gnd 1.14844f
C590 a_n1996_n452.n30 gnd 1.78382f
C591 a_n1996_n452.n31 gnd 3.22512f
C592 a_n1996_n452.n32 gnd 0.108335f
C593 a_n1996_n452.n33 gnd 0.008389f
C594 a_n1996_n452.n35 gnd 0.008389f
C595 a_n1996_n452.n37 gnd 0.286629f
C596 a_n1996_n452.n38 gnd 0.008389f
C597 a_n1996_n452.n40 gnd 0.286629f
C598 a_n1996_n452.n41 gnd 0.008389f
C599 a_n1996_n452.n43 gnd 0.286629f
C600 a_n1996_n452.n44 gnd 0.008389f
C601 a_n1996_n452.n45 gnd 0.286221f
C602 a_n1996_n452.n46 gnd 0.008389f
C603 a_n1996_n452.n47 gnd 0.286221f
C604 a_n1996_n452.n48 gnd 0.008389f
C605 a_n1996_n452.n49 gnd 0.286221f
C606 a_n1996_n452.n50 gnd 0.008389f
C607 a_n1996_n452.n51 gnd 0.286221f
C608 a_n1996_n452.n52 gnd 0.286629f
C609 a_n1996_n452.t22 gnd 0.150285f
C610 a_n1996_n452.t27 gnd 0.713776f
C611 a_n1996_n452.t13 gnd 0.699053f
C612 a_n1996_n452.t17 gnd 0.699053f
C613 a_n1996_n452.t21 gnd 0.699053f
C614 a_n1996_n452.n53 gnd 0.307348f
C615 a_n1996_n452.t23 gnd 0.710611f
C616 a_n1996_n452.t32 gnd 0.116888f
C617 a_n1996_n452.t1 gnd 0.116888f
C618 a_n1996_n452.n54 gnd 1.03516f
C619 a_n1996_n452.t4 gnd 0.116888f
C620 a_n1996_n452.t2 gnd 0.116888f
C621 a_n1996_n452.n55 gnd 1.03287f
C622 a_n1996_n452.t37 gnd 0.116888f
C623 a_n1996_n452.t36 gnd 0.116888f
C624 a_n1996_n452.n56 gnd 1.03287f
C625 a_n1996_n452.t41 gnd 0.116888f
C626 a_n1996_n452.t3 gnd 0.116888f
C627 a_n1996_n452.n57 gnd 1.03516f
C628 a_n1996_n452.t33 gnd 0.116888f
C629 a_n1996_n452.t42 gnd 0.116888f
C630 a_n1996_n452.n58 gnd 1.03287f
C631 a_n1996_n452.t43 gnd 0.116888f
C632 a_n1996_n452.t5 gnd 0.116888f
C633 a_n1996_n452.n59 gnd 1.03287f
C634 a_n1996_n452.t6 gnd 0.116888f
C635 a_n1996_n452.t34 gnd 0.116888f
C636 a_n1996_n452.n60 gnd 1.03287f
C637 a_n1996_n452.t31 gnd 0.116888f
C638 a_n1996_n452.t35 gnd 0.116888f
C639 a_n1996_n452.n61 gnd 1.03287f
C640 a_n1996_n452.t39 gnd 0.116888f
C641 a_n1996_n452.t38 gnd 0.116888f
C642 a_n1996_n452.n62 gnd 1.03516f
C643 a_n1996_n452.t40 gnd 0.116888f
C644 a_n1996_n452.t0 gnd 0.116888f
C645 a_n1996_n452.n63 gnd 1.03287f
C646 a_n1996_n452.t70 gnd 0.713776f
C647 a_n1996_n452.t53 gnd 0.699053f
C648 a_n1996_n452.t57 gnd 0.699053f
C649 a_n1996_n452.t47 gnd 0.699053f
C650 a_n1996_n452.n64 gnd 0.307348f
C651 a_n1996_n452.t62 gnd 0.699053f
C652 a_n1996_n452.t68 gnd 0.710611f
C653 a_n1996_n452.t20 gnd 1.40719f
C654 a_n1996_n452.t16 gnd 0.150285f
C655 a_n1996_n452.t10 gnd 0.150285f
C656 a_n1996_n452.n65 gnd 1.05861f
C657 a_n1996_n452.t12 gnd 0.150285f
C658 a_n1996_n452.t26 gnd 0.150285f
C659 a_n1996_n452.n66 gnd 1.05861f
C660 a_n1996_n452.t30 gnd 1.40439f
C661 a_n1996_n452.t11 gnd 0.699053f
C662 a_n1996_n452.n67 gnd 0.307348f
C663 a_n1996_n452.t25 gnd 0.699053f
C664 a_n1996_n452.t15 gnd 0.699053f
C665 a_n1996_n452.t52 gnd 0.699053f
C666 a_n1996_n452.n68 gnd 0.307348f
C667 a_n1996_n452.t61 gnd 0.699053f
C668 a_n1996_n452.t66 gnd 0.699053f
C669 a_n1996_n452.t65 gnd 0.713776f
C670 a_n1996_n452.n69 gnd 0.309974f
C671 a_n1996_n452.t45 gnd 0.699053f
C672 a_n1996_n452.n70 gnd 0.303445f
C673 a_n1996_n452.n71 gnd 0.309974f
C674 a_n1996_n452.t46 gnd 0.710611f
C675 a_n1996_n452.t19 gnd 0.713776f
C676 a_n1996_n452.n72 gnd 0.309974f
C677 a_n1996_n452.t9 gnd 0.699053f
C678 a_n1996_n452.n73 gnd 0.303445f
C679 a_n1996_n452.n74 gnd 0.309974f
C680 a_n1996_n452.t29 gnd 0.710611f
C681 a_n1996_n452.n75 gnd 1.13585f
C682 a_n1996_n452.t50 gnd 0.699053f
C683 a_n1996_n452.n76 gnd 0.303445f
C684 a_n1996_n452.t56 gnd 0.699053f
C685 a_n1996_n452.n77 gnd 0.303445f
C686 a_n1996_n452.t48 gnd 0.699053f
C687 a_n1996_n452.n78 gnd 0.303445f
C688 a_n1996_n452.t60 gnd 0.699053f
C689 a_n1996_n452.n79 gnd 0.303445f
C690 a_n1996_n452.t51 gnd 0.699053f
C691 a_n1996_n452.n80 gnd 0.297934f
C692 a_n1996_n452.t71 gnd 0.699053f
C693 a_n1996_n452.n81 gnd 0.307348f
C694 a_n1996_n452.t54 gnd 0.710766f
C695 a_n1996_n452.t63 gnd 0.699053f
C696 a_n1996_n452.n82 gnd 0.297934f
C697 a_n1996_n452.t49 gnd 0.699053f
C698 a_n1996_n452.n83 gnd 0.307348f
C699 a_n1996_n452.t58 gnd 0.710766f
C700 a_n1996_n452.t67 gnd 0.699053f
C701 a_n1996_n452.n84 gnd 0.297934f
C702 a_n1996_n452.t55 gnd 0.699053f
C703 a_n1996_n452.n85 gnd 0.307348f
C704 a_n1996_n452.t69 gnd 0.710766f
C705 a_n1996_n452.t59 gnd 0.699053f
C706 a_n1996_n452.n86 gnd 0.297934f
C707 a_n1996_n452.t44 gnd 0.699053f
C708 a_n1996_n452.n87 gnd 0.307348f
C709 a_n1996_n452.t64 gnd 0.710766f
C710 a_n1996_n452.n88 gnd 1.34296f
C711 a_n1996_n452.n89 gnd 0.309974f
C712 a_n1996_n452.n90 gnd 0.303445f
C713 a_n1996_n452.n91 gnd 0.309974f
C714 a_n1996_n452.t7 gnd 0.699053f
C715 a_n1996_n452.n92 gnd 0.309974f
C716 a_n1996_n452.n93 gnd 0.303445f
C717 a_n1996_n452.n94 gnd 0.309974f
C718 a_n1996_n452.n95 gnd 0.789588f
C719 a_n1996_n452.t28 gnd 1.40439f
C720 a_n1996_n452.t14 gnd 0.150285f
C721 a_n1996_n452.t18 gnd 0.150285f
C722 a_n1996_n452.n96 gnd 1.05861f
C723 a_n1996_n452.t24 gnd 1.40719f
C724 a_n1996_n452.n97 gnd 1.05861f
C725 a_n1996_n452.t8 gnd 0.150285f
C726 vdd.t203 gnd 0.040577f
C727 vdd.t283 gnd 0.040577f
C728 vdd.n0 gnd 0.320039f
C729 vdd.t180 gnd 0.040577f
C730 vdd.t175 gnd 0.040577f
C731 vdd.n1 gnd 0.31951f
C732 vdd.n2 gnd 0.29465f
C733 vdd.t289 gnd 0.040577f
C734 vdd.t173 gnd 0.040577f
C735 vdd.n3 gnd 0.31951f
C736 vdd.n4 gnd 0.149015f
C737 vdd.t295 gnd 0.040577f
C738 vdd.t182 gnd 0.040577f
C739 vdd.n5 gnd 0.31951f
C740 vdd.n6 gnd 0.139823f
C741 vdd.t291 gnd 0.040577f
C742 vdd.t285 gnd 0.040577f
C743 vdd.n7 gnd 0.320039f
C744 vdd.t10 gnd 0.040577f
C745 vdd.t8 gnd 0.040577f
C746 vdd.n8 gnd 0.31951f
C747 vdd.n9 gnd 0.29465f
C748 vdd.t5 gnd 0.040577f
C749 vdd.t201 gnd 0.040577f
C750 vdd.n10 gnd 0.31951f
C751 vdd.n11 gnd 0.149015f
C752 vdd.t293 gnd 0.040577f
C753 vdd.t287 gnd 0.040577f
C754 vdd.n12 gnd 0.31951f
C755 vdd.n13 gnd 0.139823f
C756 vdd.n14 gnd 0.098853f
C757 vdd.t198 gnd 0.022543f
C758 vdd.t197 gnd 0.022543f
C759 vdd.n15 gnd 0.207498f
C760 vdd.t194 gnd 0.022543f
C761 vdd.t187 gnd 0.022543f
C762 vdd.n16 gnd 0.206891f
C763 vdd.n17 gnd 0.360054f
C764 vdd.t190 gnd 0.022543f
C765 vdd.t196 gnd 0.022543f
C766 vdd.n18 gnd 0.206891f
C767 vdd.n19 gnd 0.148959f
C768 vdd.t185 gnd 0.022543f
C769 vdd.t189 gnd 0.022543f
C770 vdd.n20 gnd 0.207498f
C771 vdd.t186 gnd 0.022543f
C772 vdd.t191 gnd 0.022543f
C773 vdd.n21 gnd 0.206891f
C774 vdd.n22 gnd 0.360054f
C775 vdd.t183 gnd 0.022543f
C776 vdd.t184 gnd 0.022543f
C777 vdd.n23 gnd 0.206891f
C778 vdd.n24 gnd 0.148959f
C779 vdd.t192 gnd 0.022543f
C780 vdd.t195 gnd 0.022543f
C781 vdd.n25 gnd 0.206891f
C782 vdd.t193 gnd 0.022543f
C783 vdd.t188 gnd 0.022543f
C784 vdd.n26 gnd 0.206891f
C785 vdd.n27 gnd 23.8355f
C786 vdd.n28 gnd 8.87019f
C787 vdd.n29 gnd 0.006148f
C788 vdd.n30 gnd 0.005705f
C789 vdd.n31 gnd 0.003156f
C790 vdd.n32 gnd 0.007247f
C791 vdd.n33 gnd 0.003066f
C792 vdd.n34 gnd 0.003246f
C793 vdd.n35 gnd 0.005705f
C794 vdd.n36 gnd 0.003066f
C795 vdd.n37 gnd 0.007247f
C796 vdd.n38 gnd 0.003246f
C797 vdd.n39 gnd 0.005705f
C798 vdd.n40 gnd 0.003066f
C799 vdd.n41 gnd 0.005435f
C800 vdd.n42 gnd 0.005451f
C801 vdd.t14 gnd 0.015569f
C802 vdd.n43 gnd 0.03464f
C803 vdd.n44 gnd 0.180273f
C804 vdd.n45 gnd 0.003066f
C805 vdd.n46 gnd 0.003246f
C806 vdd.n47 gnd 0.007247f
C807 vdd.n48 gnd 0.007247f
C808 vdd.n49 gnd 0.003246f
C809 vdd.n50 gnd 0.003066f
C810 vdd.n51 gnd 0.005705f
C811 vdd.n52 gnd 0.005705f
C812 vdd.n53 gnd 0.003066f
C813 vdd.n54 gnd 0.003246f
C814 vdd.n55 gnd 0.007247f
C815 vdd.n56 gnd 0.007247f
C816 vdd.n57 gnd 0.003246f
C817 vdd.n58 gnd 0.003066f
C818 vdd.n59 gnd 0.005705f
C819 vdd.n60 gnd 0.005705f
C820 vdd.n61 gnd 0.003066f
C821 vdd.n62 gnd 0.003246f
C822 vdd.n63 gnd 0.007247f
C823 vdd.n64 gnd 0.007247f
C824 vdd.n65 gnd 0.017132f
C825 vdd.n66 gnd 0.003156f
C826 vdd.n67 gnd 0.003066f
C827 vdd.n68 gnd 0.014747f
C828 vdd.n69 gnd 0.010295f
C829 vdd.t155 gnd 0.036069f
C830 vdd.t95 gnd 0.036069f
C831 vdd.n70 gnd 0.247888f
C832 vdd.n71 gnd 0.194926f
C833 vdd.t168 gnd 0.036069f
C834 vdd.t61 gnd 0.036069f
C835 vdd.n72 gnd 0.247888f
C836 vdd.n73 gnd 0.157304f
C837 vdd.t143 gnd 0.036069f
C838 vdd.t85 gnd 0.036069f
C839 vdd.n74 gnd 0.247888f
C840 vdd.n75 gnd 0.157304f
C841 vdd.t163 gnd 0.036069f
C842 vdd.t137 gnd 0.036069f
C843 vdd.n76 gnd 0.247888f
C844 vdd.n77 gnd 0.157304f
C845 vdd.t26 gnd 0.036069f
C846 vdd.t74 gnd 0.036069f
C847 vdd.n78 gnd 0.247888f
C848 vdd.n79 gnd 0.157304f
C849 vdd.t38 gnd 0.036069f
C850 vdd.t98 gnd 0.036069f
C851 vdd.n80 gnd 0.247888f
C852 vdd.n81 gnd 0.157304f
C853 vdd.t69 gnd 0.036069f
C854 vdd.t151 gnd 0.036069f
C855 vdd.n82 gnd 0.247888f
C856 vdd.n83 gnd 0.157304f
C857 vdd.t43 gnd 0.036069f
C858 vdd.t122 gnd 0.036069f
C859 vdd.n84 gnd 0.247888f
C860 vdd.n85 gnd 0.157304f
C861 vdd.t51 gnd 0.036069f
C862 vdd.t138 gnd 0.036069f
C863 vdd.n86 gnd 0.247888f
C864 vdd.n87 gnd 0.157304f
C865 vdd.n88 gnd 0.006148f
C866 vdd.n89 gnd 0.005705f
C867 vdd.n90 gnd 0.003156f
C868 vdd.n91 gnd 0.007247f
C869 vdd.n92 gnd 0.003066f
C870 vdd.n93 gnd 0.003246f
C871 vdd.n94 gnd 0.005705f
C872 vdd.n95 gnd 0.003066f
C873 vdd.n96 gnd 0.007247f
C874 vdd.n97 gnd 0.003246f
C875 vdd.n98 gnd 0.005705f
C876 vdd.n99 gnd 0.003066f
C877 vdd.n100 gnd 0.005435f
C878 vdd.n101 gnd 0.005451f
C879 vdd.t80 gnd 0.015569f
C880 vdd.n102 gnd 0.03464f
C881 vdd.n103 gnd 0.180273f
C882 vdd.n104 gnd 0.003066f
C883 vdd.n105 gnd 0.003246f
C884 vdd.n106 gnd 0.007247f
C885 vdd.n107 gnd 0.007247f
C886 vdd.n108 gnd 0.003246f
C887 vdd.n109 gnd 0.003066f
C888 vdd.n110 gnd 0.005705f
C889 vdd.n111 gnd 0.005705f
C890 vdd.n112 gnd 0.003066f
C891 vdd.n113 gnd 0.003246f
C892 vdd.n114 gnd 0.007247f
C893 vdd.n115 gnd 0.007247f
C894 vdd.n116 gnd 0.003246f
C895 vdd.n117 gnd 0.003066f
C896 vdd.n118 gnd 0.005705f
C897 vdd.n119 gnd 0.005705f
C898 vdd.n120 gnd 0.003066f
C899 vdd.n121 gnd 0.003246f
C900 vdd.n122 gnd 0.007247f
C901 vdd.n123 gnd 0.007247f
C902 vdd.n124 gnd 0.017132f
C903 vdd.n125 gnd 0.003156f
C904 vdd.n126 gnd 0.003066f
C905 vdd.n127 gnd 0.014747f
C906 vdd.n128 gnd 0.009972f
C907 vdd.n129 gnd 0.117035f
C908 vdd.n130 gnd 0.006148f
C909 vdd.n131 gnd 0.005705f
C910 vdd.n132 gnd 0.003156f
C911 vdd.n133 gnd 0.007247f
C912 vdd.n134 gnd 0.003066f
C913 vdd.n135 gnd 0.003246f
C914 vdd.n136 gnd 0.005705f
C915 vdd.n137 gnd 0.003066f
C916 vdd.n138 gnd 0.007247f
C917 vdd.n139 gnd 0.003246f
C918 vdd.n140 gnd 0.005705f
C919 vdd.n141 gnd 0.003066f
C920 vdd.n142 gnd 0.005435f
C921 vdd.n143 gnd 0.005451f
C922 vdd.t101 gnd 0.015569f
C923 vdd.n144 gnd 0.03464f
C924 vdd.n145 gnd 0.180273f
C925 vdd.n146 gnd 0.003066f
C926 vdd.n147 gnd 0.003246f
C927 vdd.n148 gnd 0.007247f
C928 vdd.n149 gnd 0.007247f
C929 vdd.n150 gnd 0.003246f
C930 vdd.n151 gnd 0.003066f
C931 vdd.n152 gnd 0.005705f
C932 vdd.n153 gnd 0.005705f
C933 vdd.n154 gnd 0.003066f
C934 vdd.n155 gnd 0.003246f
C935 vdd.n156 gnd 0.007247f
C936 vdd.n157 gnd 0.007247f
C937 vdd.n158 gnd 0.003246f
C938 vdd.n159 gnd 0.003066f
C939 vdd.n160 gnd 0.005705f
C940 vdd.n161 gnd 0.005705f
C941 vdd.n162 gnd 0.003066f
C942 vdd.n163 gnd 0.003246f
C943 vdd.n164 gnd 0.007247f
C944 vdd.n165 gnd 0.007247f
C945 vdd.n166 gnd 0.017132f
C946 vdd.n167 gnd 0.003156f
C947 vdd.n168 gnd 0.003066f
C948 vdd.n169 gnd 0.014747f
C949 vdd.n170 gnd 0.010295f
C950 vdd.t103 gnd 0.036069f
C951 vdd.t132 gnd 0.036069f
C952 vdd.n171 gnd 0.247888f
C953 vdd.n172 gnd 0.194926f
C954 vdd.t24 gnd 0.036069f
C955 vdd.t93 gnd 0.036069f
C956 vdd.n173 gnd 0.247888f
C957 vdd.n174 gnd 0.157304f
C958 vdd.t130 gnd 0.036069f
C959 vdd.t12 gnd 0.036069f
C960 vdd.n175 gnd 0.247888f
C961 vdd.n176 gnd 0.157304f
C962 vdd.t71 gnd 0.036069f
C963 vdd.t73 gnd 0.036069f
C964 vdd.n177 gnd 0.247888f
C965 vdd.n178 gnd 0.157304f
C966 vdd.t157 gnd 0.036069f
C967 vdd.t66 gnd 0.036069f
C968 vdd.n179 gnd 0.247888f
C969 vdd.n180 gnd 0.157304f
C970 vdd.t67 gnd 0.036069f
C971 vdd.t153 gnd 0.036069f
C972 vdd.n181 gnd 0.247888f
C973 vdd.n182 gnd 0.157304f
C974 vdd.t154 gnd 0.036069f
C975 vdd.t36 gnd 0.036069f
C976 vdd.n183 gnd 0.247888f
C977 vdd.n184 gnd 0.157304f
C978 vdd.t131 gnd 0.036069f
C979 vdd.t150 gnd 0.036069f
C980 vdd.n185 gnd 0.247888f
C981 vdd.n186 gnd 0.157304f
C982 vdd.t34 gnd 0.036069f
C983 vdd.t92 gnd 0.036069f
C984 vdd.n187 gnd 0.247888f
C985 vdd.n188 gnd 0.157304f
C986 vdd.n189 gnd 0.006148f
C987 vdd.n190 gnd 0.005705f
C988 vdd.n191 gnd 0.003156f
C989 vdd.n192 gnd 0.007247f
C990 vdd.n193 gnd 0.003066f
C991 vdd.n194 gnd 0.003246f
C992 vdd.n195 gnd 0.005705f
C993 vdd.n196 gnd 0.003066f
C994 vdd.n197 gnd 0.007247f
C995 vdd.n198 gnd 0.003246f
C996 vdd.n199 gnd 0.005705f
C997 vdd.n200 gnd 0.003066f
C998 vdd.n201 gnd 0.005435f
C999 vdd.n202 gnd 0.005451f
C1000 vdd.t128 gnd 0.015569f
C1001 vdd.n203 gnd 0.03464f
C1002 vdd.n204 gnd 0.180273f
C1003 vdd.n205 gnd 0.003066f
C1004 vdd.n206 gnd 0.003246f
C1005 vdd.n207 gnd 0.007247f
C1006 vdd.n208 gnd 0.007247f
C1007 vdd.n209 gnd 0.003246f
C1008 vdd.n210 gnd 0.003066f
C1009 vdd.n211 gnd 0.005705f
C1010 vdd.n212 gnd 0.005705f
C1011 vdd.n213 gnd 0.003066f
C1012 vdd.n214 gnd 0.003246f
C1013 vdd.n215 gnd 0.007247f
C1014 vdd.n216 gnd 0.007247f
C1015 vdd.n217 gnd 0.003246f
C1016 vdd.n218 gnd 0.003066f
C1017 vdd.n219 gnd 0.005705f
C1018 vdd.n220 gnd 0.005705f
C1019 vdd.n221 gnd 0.003066f
C1020 vdd.n222 gnd 0.003246f
C1021 vdd.n223 gnd 0.007247f
C1022 vdd.n224 gnd 0.007247f
C1023 vdd.n225 gnd 0.017132f
C1024 vdd.n226 gnd 0.003156f
C1025 vdd.n227 gnd 0.003066f
C1026 vdd.n228 gnd 0.014747f
C1027 vdd.n229 gnd 0.009972f
C1028 vdd.n230 gnd 0.069624f
C1029 vdd.n231 gnd 0.250874f
C1030 vdd.n232 gnd 0.006148f
C1031 vdd.n233 gnd 0.005705f
C1032 vdd.n234 gnd 0.003156f
C1033 vdd.n235 gnd 0.007247f
C1034 vdd.n236 gnd 0.003066f
C1035 vdd.n237 gnd 0.003246f
C1036 vdd.n238 gnd 0.005705f
C1037 vdd.n239 gnd 0.003066f
C1038 vdd.n240 gnd 0.007247f
C1039 vdd.n241 gnd 0.003246f
C1040 vdd.n242 gnd 0.005705f
C1041 vdd.n243 gnd 0.003066f
C1042 vdd.n244 gnd 0.005435f
C1043 vdd.n245 gnd 0.005451f
C1044 vdd.t115 gnd 0.015569f
C1045 vdd.n246 gnd 0.03464f
C1046 vdd.n247 gnd 0.180273f
C1047 vdd.n248 gnd 0.003066f
C1048 vdd.n249 gnd 0.003246f
C1049 vdd.n250 gnd 0.007247f
C1050 vdd.n251 gnd 0.007247f
C1051 vdd.n252 gnd 0.003246f
C1052 vdd.n253 gnd 0.003066f
C1053 vdd.n254 gnd 0.005705f
C1054 vdd.n255 gnd 0.005705f
C1055 vdd.n256 gnd 0.003066f
C1056 vdd.n257 gnd 0.003246f
C1057 vdd.n258 gnd 0.007247f
C1058 vdd.n259 gnd 0.007247f
C1059 vdd.n260 gnd 0.003246f
C1060 vdd.n261 gnd 0.003066f
C1061 vdd.n262 gnd 0.005705f
C1062 vdd.n263 gnd 0.005705f
C1063 vdd.n264 gnd 0.003066f
C1064 vdd.n265 gnd 0.003246f
C1065 vdd.n266 gnd 0.007247f
C1066 vdd.n267 gnd 0.007247f
C1067 vdd.n268 gnd 0.017132f
C1068 vdd.n269 gnd 0.003156f
C1069 vdd.n270 gnd 0.003066f
C1070 vdd.n271 gnd 0.014747f
C1071 vdd.n272 gnd 0.010295f
C1072 vdd.t116 gnd 0.036069f
C1073 vdd.t147 gnd 0.036069f
C1074 vdd.n273 gnd 0.247888f
C1075 vdd.n274 gnd 0.194926f
C1076 vdd.t48 gnd 0.036069f
C1077 vdd.t112 gnd 0.036069f
C1078 vdd.n275 gnd 0.247888f
C1079 vdd.n276 gnd 0.157304f
C1080 vdd.t140 gnd 0.036069f
C1081 vdd.t41 gnd 0.036069f
C1082 vdd.n277 gnd 0.247888f
C1083 vdd.n278 gnd 0.157304f
C1084 vdd.t88 gnd 0.036069f
C1085 vdd.t90 gnd 0.036069f
C1086 vdd.n279 gnd 0.247888f
C1087 vdd.n280 gnd 0.157304f
C1088 vdd.t167 gnd 0.036069f
C1089 vdd.t83 gnd 0.036069f
C1090 vdd.n281 gnd 0.247888f
C1091 vdd.n282 gnd 0.157304f
C1092 vdd.t84 gnd 0.036069f
C1093 vdd.t165 gnd 0.036069f
C1094 vdd.n283 gnd 0.247888f
C1095 vdd.n284 gnd 0.157304f
C1096 vdd.t166 gnd 0.036069f
C1097 vdd.t59 gnd 0.036069f
C1098 vdd.n285 gnd 0.247888f
C1099 vdd.n286 gnd 0.157304f
C1100 vdd.t145 gnd 0.036069f
C1101 vdd.t162 gnd 0.036069f
C1102 vdd.n287 gnd 0.247888f
C1103 vdd.n288 gnd 0.157304f
C1104 vdd.t52 gnd 0.036069f
C1105 vdd.t113 gnd 0.036069f
C1106 vdd.n289 gnd 0.247888f
C1107 vdd.n290 gnd 0.157304f
C1108 vdd.n291 gnd 0.006148f
C1109 vdd.n292 gnd 0.005705f
C1110 vdd.n293 gnd 0.003156f
C1111 vdd.n294 gnd 0.007247f
C1112 vdd.n295 gnd 0.003066f
C1113 vdd.n296 gnd 0.003246f
C1114 vdd.n297 gnd 0.005705f
C1115 vdd.n298 gnd 0.003066f
C1116 vdd.n299 gnd 0.007247f
C1117 vdd.n300 gnd 0.003246f
C1118 vdd.n301 gnd 0.005705f
C1119 vdd.n302 gnd 0.003066f
C1120 vdd.n303 gnd 0.005435f
C1121 vdd.n304 gnd 0.005451f
C1122 vdd.t141 gnd 0.015569f
C1123 vdd.n305 gnd 0.03464f
C1124 vdd.n306 gnd 0.180273f
C1125 vdd.n307 gnd 0.003066f
C1126 vdd.n308 gnd 0.003246f
C1127 vdd.n309 gnd 0.007247f
C1128 vdd.n310 gnd 0.007247f
C1129 vdd.n311 gnd 0.003246f
C1130 vdd.n312 gnd 0.003066f
C1131 vdd.n313 gnd 0.005705f
C1132 vdd.n314 gnd 0.005705f
C1133 vdd.n315 gnd 0.003066f
C1134 vdd.n316 gnd 0.003246f
C1135 vdd.n317 gnd 0.007247f
C1136 vdd.n318 gnd 0.007247f
C1137 vdd.n319 gnd 0.003246f
C1138 vdd.n320 gnd 0.003066f
C1139 vdd.n321 gnd 0.005705f
C1140 vdd.n322 gnd 0.005705f
C1141 vdd.n323 gnd 0.003066f
C1142 vdd.n324 gnd 0.003246f
C1143 vdd.n325 gnd 0.007247f
C1144 vdd.n326 gnd 0.007247f
C1145 vdd.n327 gnd 0.017132f
C1146 vdd.n328 gnd 0.003156f
C1147 vdd.n329 gnd 0.003066f
C1148 vdd.n330 gnd 0.014747f
C1149 vdd.n331 gnd 0.009972f
C1150 vdd.n332 gnd 0.069624f
C1151 vdd.n333 gnd 0.287196f
C1152 vdd.n334 gnd 0.00861f
C1153 vdd.n335 gnd 0.011203f
C1154 vdd.n336 gnd 0.009017f
C1155 vdd.n337 gnd 0.009017f
C1156 vdd.n338 gnd 0.011203f
C1157 vdd.n339 gnd 0.011203f
C1158 vdd.n340 gnd 0.818607f
C1159 vdd.n341 gnd 0.011203f
C1160 vdd.n342 gnd 0.011203f
C1161 vdd.n343 gnd 0.011203f
C1162 vdd.n344 gnd 0.887302f
C1163 vdd.n345 gnd 0.011203f
C1164 vdd.n346 gnd 0.011203f
C1165 vdd.n347 gnd 0.011203f
C1166 vdd.n348 gnd 0.011203f
C1167 vdd.n349 gnd 0.009017f
C1168 vdd.n350 gnd 0.011203f
C1169 vdd.t97 gnd 0.572453f
C1170 vdd.n351 gnd 0.011203f
C1171 vdd.n352 gnd 0.011203f
C1172 vdd.n353 gnd 0.011203f
C1173 vdd.t35 gnd 0.572453f
C1174 vdd.n354 gnd 0.011203f
C1175 vdd.n355 gnd 0.011203f
C1176 vdd.n356 gnd 0.011203f
C1177 vdd.n357 gnd 0.011203f
C1178 vdd.n358 gnd 0.011203f
C1179 vdd.n359 gnd 0.009017f
C1180 vdd.n360 gnd 0.011203f
C1181 vdd.n361 gnd 0.646871f
C1182 vdd.n362 gnd 0.011203f
C1183 vdd.n363 gnd 0.011203f
C1184 vdd.n364 gnd 0.011203f
C1185 vdd.t121 gnd 0.572453f
C1186 vdd.n365 gnd 0.011203f
C1187 vdd.n366 gnd 0.011203f
C1188 vdd.n367 gnd 0.011203f
C1189 vdd.n368 gnd 0.011203f
C1190 vdd.n369 gnd 0.011203f
C1191 vdd.n370 gnd 0.009017f
C1192 vdd.n371 gnd 0.011203f
C1193 vdd.t33 gnd 0.572453f
C1194 vdd.n372 gnd 0.011203f
C1195 vdd.n373 gnd 0.011203f
C1196 vdd.n374 gnd 0.011203f
C1197 vdd.n375 gnd 0.66977f
C1198 vdd.n376 gnd 0.011203f
C1199 vdd.n377 gnd 0.011203f
C1200 vdd.n378 gnd 0.011203f
C1201 vdd.n379 gnd 0.011203f
C1202 vdd.n380 gnd 0.011203f
C1203 vdd.n381 gnd 0.009017f
C1204 vdd.n382 gnd 0.011203f
C1205 vdd.t79 gnd 0.572453f
C1206 vdd.n383 gnd 0.011203f
C1207 vdd.n384 gnd 0.011203f
C1208 vdd.n385 gnd 0.011203f
C1209 vdd.n386 gnd 0.578177f
C1210 vdd.n387 gnd 0.011203f
C1211 vdd.n388 gnd 0.011203f
C1212 vdd.n389 gnd 0.011203f
C1213 vdd.n390 gnd 0.011203f
C1214 vdd.n391 gnd 0.027101f
C1215 vdd.n392 gnd 0.027682f
C1216 vdd.t233 gnd 0.572453f
C1217 vdd.n393 gnd 0.027101f
C1218 vdd.n425 gnd 0.011203f
C1219 vdd.t235 gnd 0.137828f
C1220 vdd.t234 gnd 0.1473f
C1221 vdd.t232 gnd 0.180001f
C1222 vdd.n426 gnd 0.230736f
C1223 vdd.n427 gnd 0.194762f
C1224 vdd.n428 gnd 0.014788f
C1225 vdd.n429 gnd 0.011203f
C1226 vdd.n430 gnd 0.009017f
C1227 vdd.n431 gnd 0.011203f
C1228 vdd.n432 gnd 0.009017f
C1229 vdd.n433 gnd 0.011203f
C1230 vdd.n434 gnd 0.009017f
C1231 vdd.n435 gnd 0.011203f
C1232 vdd.n436 gnd 0.009017f
C1233 vdd.n437 gnd 0.011203f
C1234 vdd.n438 gnd 0.009017f
C1235 vdd.n439 gnd 0.011203f
C1236 vdd.t275 gnd 0.137828f
C1237 vdd.t274 gnd 0.1473f
C1238 vdd.t273 gnd 0.180001f
C1239 vdd.n440 gnd 0.230736f
C1240 vdd.n441 gnd 0.194762f
C1241 vdd.n442 gnd 0.009017f
C1242 vdd.n443 gnd 0.011203f
C1243 vdd.n444 gnd 0.009017f
C1244 vdd.n445 gnd 0.011203f
C1245 vdd.n446 gnd 0.009017f
C1246 vdd.n447 gnd 0.011203f
C1247 vdd.n448 gnd 0.009017f
C1248 vdd.n449 gnd 0.011203f
C1249 vdd.n450 gnd 0.009017f
C1250 vdd.n451 gnd 0.011203f
C1251 vdd.t281 gnd 0.137828f
C1252 vdd.t280 gnd 0.1473f
C1253 vdd.t279 gnd 0.180001f
C1254 vdd.n452 gnd 0.230736f
C1255 vdd.n453 gnd 0.194762f
C1256 vdd.n454 gnd 0.019297f
C1257 vdd.n455 gnd 0.011203f
C1258 vdd.n456 gnd 0.009017f
C1259 vdd.n457 gnd 0.011203f
C1260 vdd.n458 gnd 0.009017f
C1261 vdd.n459 gnd 0.011203f
C1262 vdd.n460 gnd 0.009017f
C1263 vdd.n461 gnd 0.011203f
C1264 vdd.n462 gnd 0.009017f
C1265 vdd.n463 gnd 0.011203f
C1266 vdd.n464 gnd 0.027682f
C1267 vdd.n465 gnd 0.007484f
C1268 vdd.n466 gnd 0.009017f
C1269 vdd.n467 gnd 0.011203f
C1270 vdd.n468 gnd 0.011203f
C1271 vdd.n469 gnd 0.009017f
C1272 vdd.n470 gnd 0.011203f
C1273 vdd.n471 gnd 0.011203f
C1274 vdd.n472 gnd 0.011203f
C1275 vdd.n473 gnd 0.011203f
C1276 vdd.n474 gnd 0.011203f
C1277 vdd.n475 gnd 0.009017f
C1278 vdd.n476 gnd 0.009017f
C1279 vdd.n477 gnd 0.011203f
C1280 vdd.n478 gnd 0.011203f
C1281 vdd.n479 gnd 0.009017f
C1282 vdd.n480 gnd 0.011203f
C1283 vdd.n481 gnd 0.011203f
C1284 vdd.n482 gnd 0.011203f
C1285 vdd.n483 gnd 0.011203f
C1286 vdd.n484 gnd 0.011203f
C1287 vdd.n485 gnd 0.009017f
C1288 vdd.n486 gnd 0.009017f
C1289 vdd.n487 gnd 0.011203f
C1290 vdd.n488 gnd 0.011203f
C1291 vdd.n489 gnd 0.009017f
C1292 vdd.n490 gnd 0.011203f
C1293 vdd.n491 gnd 0.011203f
C1294 vdd.n492 gnd 0.011203f
C1295 vdd.n493 gnd 0.011203f
C1296 vdd.n494 gnd 0.011203f
C1297 vdd.n495 gnd 0.009017f
C1298 vdd.n496 gnd 0.009017f
C1299 vdd.n497 gnd 0.011203f
C1300 vdd.n498 gnd 0.011203f
C1301 vdd.n499 gnd 0.009017f
C1302 vdd.n500 gnd 0.011203f
C1303 vdd.n501 gnd 0.011203f
C1304 vdd.n502 gnd 0.011203f
C1305 vdd.n503 gnd 0.011203f
C1306 vdd.n504 gnd 0.011203f
C1307 vdd.n505 gnd 0.009017f
C1308 vdd.n506 gnd 0.009017f
C1309 vdd.n507 gnd 0.011203f
C1310 vdd.n508 gnd 0.011203f
C1311 vdd.n509 gnd 0.007529f
C1312 vdd.n510 gnd 0.011203f
C1313 vdd.n511 gnd 0.011203f
C1314 vdd.n512 gnd 0.011203f
C1315 vdd.n513 gnd 0.011203f
C1316 vdd.n514 gnd 0.011203f
C1317 vdd.n515 gnd 0.007529f
C1318 vdd.n516 gnd 0.009017f
C1319 vdd.n517 gnd 0.011203f
C1320 vdd.n518 gnd 0.011203f
C1321 vdd.n519 gnd 0.009017f
C1322 vdd.n520 gnd 0.011203f
C1323 vdd.n521 gnd 0.011203f
C1324 vdd.n522 gnd 0.011203f
C1325 vdd.n523 gnd 0.011203f
C1326 vdd.n524 gnd 0.011203f
C1327 vdd.n525 gnd 0.009017f
C1328 vdd.n526 gnd 0.009017f
C1329 vdd.n527 gnd 0.011203f
C1330 vdd.n528 gnd 0.011203f
C1331 vdd.n529 gnd 0.009017f
C1332 vdd.n530 gnd 0.011203f
C1333 vdd.n531 gnd 0.011203f
C1334 vdd.n532 gnd 0.011203f
C1335 vdd.n533 gnd 0.011203f
C1336 vdd.n534 gnd 0.011203f
C1337 vdd.n535 gnd 0.009017f
C1338 vdd.n536 gnd 0.009017f
C1339 vdd.n537 gnd 0.011203f
C1340 vdd.n538 gnd 0.011203f
C1341 vdd.n539 gnd 0.009017f
C1342 vdd.n540 gnd 0.011203f
C1343 vdd.n541 gnd 0.011203f
C1344 vdd.n542 gnd 0.011203f
C1345 vdd.n543 gnd 0.011203f
C1346 vdd.n544 gnd 0.011203f
C1347 vdd.n545 gnd 0.009017f
C1348 vdd.n546 gnd 0.009017f
C1349 vdd.n547 gnd 0.011203f
C1350 vdd.n548 gnd 0.011203f
C1351 vdd.n549 gnd 0.009017f
C1352 vdd.n550 gnd 0.011203f
C1353 vdd.n551 gnd 0.011203f
C1354 vdd.n552 gnd 0.011203f
C1355 vdd.n553 gnd 0.011203f
C1356 vdd.n554 gnd 0.011203f
C1357 vdd.n555 gnd 0.009017f
C1358 vdd.n556 gnd 0.009017f
C1359 vdd.n557 gnd 0.011203f
C1360 vdd.n558 gnd 0.011203f
C1361 vdd.n559 gnd 0.009017f
C1362 vdd.n560 gnd 0.011203f
C1363 vdd.n561 gnd 0.011203f
C1364 vdd.n562 gnd 0.011203f
C1365 vdd.n563 gnd 0.011203f
C1366 vdd.n564 gnd 0.011203f
C1367 vdd.n565 gnd 0.006132f
C1368 vdd.n566 gnd 0.019297f
C1369 vdd.n567 gnd 0.011203f
C1370 vdd.n568 gnd 0.011203f
C1371 vdd.n569 gnd 0.008927f
C1372 vdd.n570 gnd 0.011203f
C1373 vdd.n571 gnd 0.011203f
C1374 vdd.n572 gnd 0.011203f
C1375 vdd.n573 gnd 0.011203f
C1376 vdd.n574 gnd 0.011203f
C1377 vdd.n575 gnd 0.009017f
C1378 vdd.n576 gnd 0.009017f
C1379 vdd.n577 gnd 0.011203f
C1380 vdd.n578 gnd 0.011203f
C1381 vdd.n579 gnd 0.009017f
C1382 vdd.n580 gnd 0.011203f
C1383 vdd.n581 gnd 0.011203f
C1384 vdd.n582 gnd 0.011203f
C1385 vdd.n583 gnd 0.011203f
C1386 vdd.n584 gnd 0.011203f
C1387 vdd.n585 gnd 0.009017f
C1388 vdd.n586 gnd 0.009017f
C1389 vdd.n587 gnd 0.011203f
C1390 vdd.n588 gnd 0.011203f
C1391 vdd.n589 gnd 0.009017f
C1392 vdd.n590 gnd 0.011203f
C1393 vdd.n591 gnd 0.011203f
C1394 vdd.n592 gnd 0.011203f
C1395 vdd.n593 gnd 0.011203f
C1396 vdd.n594 gnd 0.011203f
C1397 vdd.n595 gnd 0.009017f
C1398 vdd.n596 gnd 0.009017f
C1399 vdd.n597 gnd 0.011203f
C1400 vdd.n598 gnd 0.011203f
C1401 vdd.n599 gnd 0.009017f
C1402 vdd.n600 gnd 0.011203f
C1403 vdd.n601 gnd 0.011203f
C1404 vdd.n602 gnd 0.011203f
C1405 vdd.n603 gnd 0.011203f
C1406 vdd.n604 gnd 0.011203f
C1407 vdd.n605 gnd 0.009017f
C1408 vdd.n606 gnd 0.009017f
C1409 vdd.n607 gnd 0.011203f
C1410 vdd.n608 gnd 0.011203f
C1411 vdd.n609 gnd 0.009017f
C1412 vdd.n610 gnd 0.011203f
C1413 vdd.n611 gnd 0.011203f
C1414 vdd.n612 gnd 0.011203f
C1415 vdd.n613 gnd 0.011203f
C1416 vdd.n614 gnd 0.011203f
C1417 vdd.n615 gnd 0.009017f
C1418 vdd.n616 gnd 0.011203f
C1419 vdd.n617 gnd 0.009017f
C1420 vdd.n618 gnd 0.004734f
C1421 vdd.n619 gnd 0.011203f
C1422 vdd.n620 gnd 0.011203f
C1423 vdd.n621 gnd 0.009017f
C1424 vdd.n622 gnd 0.011203f
C1425 vdd.n623 gnd 0.009017f
C1426 vdd.n624 gnd 0.011203f
C1427 vdd.n625 gnd 0.009017f
C1428 vdd.n626 gnd 0.011203f
C1429 vdd.n627 gnd 0.009017f
C1430 vdd.n628 gnd 0.011203f
C1431 vdd.n629 gnd 0.009017f
C1432 vdd.n630 gnd 0.011203f
C1433 vdd.n631 gnd 0.009017f
C1434 vdd.n632 gnd 0.011203f
C1435 vdd.n633 gnd 0.623973f
C1436 vdd.t25 gnd 0.572453f
C1437 vdd.n634 gnd 0.011203f
C1438 vdd.n635 gnd 0.009017f
C1439 vdd.n636 gnd 0.011203f
C1440 vdd.n637 gnd 0.009017f
C1441 vdd.n638 gnd 0.011203f
C1442 vdd.t70 gnd 0.572453f
C1443 vdd.n639 gnd 0.011203f
C1444 vdd.n640 gnd 0.009017f
C1445 vdd.n641 gnd 0.011203f
C1446 vdd.n642 gnd 0.009017f
C1447 vdd.n643 gnd 0.011203f
C1448 vdd.t11 gnd 0.572453f
C1449 vdd.n644 gnd 0.715566f
C1450 vdd.n645 gnd 0.011203f
C1451 vdd.n646 gnd 0.009017f
C1452 vdd.n647 gnd 0.011203f
C1453 vdd.n648 gnd 0.009017f
C1454 vdd.n649 gnd 0.011203f
C1455 vdd.t129 gnd 0.572453f
C1456 vdd.n650 gnd 0.011203f
C1457 vdd.n651 gnd 0.009017f
C1458 vdd.n652 gnd 0.011203f
C1459 vdd.n653 gnd 0.009017f
C1460 vdd.n654 gnd 0.011203f
C1461 vdd.n655 gnd 0.795709f
C1462 vdd.n656 gnd 0.950271f
C1463 vdd.t60 gnd 0.572453f
C1464 vdd.n657 gnd 0.011203f
C1465 vdd.n658 gnd 0.009017f
C1466 vdd.n659 gnd 0.011203f
C1467 vdd.n660 gnd 0.009017f
C1468 vdd.n661 gnd 0.011203f
C1469 vdd.n662 gnd 0.601075f
C1470 vdd.n663 gnd 0.011203f
C1471 vdd.n664 gnd 0.009017f
C1472 vdd.n665 gnd 0.011203f
C1473 vdd.n666 gnd 0.009017f
C1474 vdd.n667 gnd 0.011203f
C1475 vdd.t102 gnd 0.572453f
C1476 vdd.t94 gnd 0.572453f
C1477 vdd.n668 gnd 0.011203f
C1478 vdd.n669 gnd 0.009017f
C1479 vdd.n670 gnd 0.011203f
C1480 vdd.n671 gnd 0.009017f
C1481 vdd.n672 gnd 0.011203f
C1482 vdd.t13 gnd 0.572453f
C1483 vdd.n673 gnd 0.011203f
C1484 vdd.n674 gnd 0.009017f
C1485 vdd.n675 gnd 0.011203f
C1486 vdd.n676 gnd 0.009017f
C1487 vdd.n677 gnd 0.011203f
C1488 vdd.n678 gnd 1.14491f
C1489 vdd.n679 gnd 0.933098f
C1490 vdd.n680 gnd 0.011203f
C1491 vdd.n681 gnd 0.009017f
C1492 vdd.n682 gnd 0.027101f
C1493 vdd.n683 gnd 0.007484f
C1494 vdd.n684 gnd 0.027101f
C1495 vdd.t211 gnd 0.572453f
C1496 vdd.n685 gnd 0.027101f
C1497 vdd.n686 gnd 0.007484f
C1498 vdd.n687 gnd 0.009635f
C1499 vdd.t277 gnd 0.137828f
C1500 vdd.t278 gnd 0.1473f
C1501 vdd.t276 gnd 0.180001f
C1502 vdd.n688 gnd 0.230736f
C1503 vdd.n689 gnd 0.19386f
C1504 vdd.n690 gnd 0.013886f
C1505 vdd.n691 gnd 0.011203f
C1506 vdd.n692 gnd 7.8884f
C1507 vdd.n723 gnd 1.57424f
C1508 vdd.n724 gnd 0.011203f
C1509 vdd.n725 gnd 0.011203f
C1510 vdd.n726 gnd 0.027682f
C1511 vdd.n727 gnd 0.009635f
C1512 vdd.n728 gnd 0.011203f
C1513 vdd.n729 gnd 0.009017f
C1514 vdd.n730 gnd 0.00717f
C1515 vdd.n731 gnd 0.018307f
C1516 vdd.n732 gnd 0.009017f
C1517 vdd.n733 gnd 0.011203f
C1518 vdd.n734 gnd 0.011203f
C1519 vdd.n735 gnd 0.011203f
C1520 vdd.n736 gnd 0.011203f
C1521 vdd.n737 gnd 0.011203f
C1522 vdd.n738 gnd 0.011203f
C1523 vdd.n739 gnd 0.011203f
C1524 vdd.n740 gnd 0.011203f
C1525 vdd.n741 gnd 0.011203f
C1526 vdd.n742 gnd 0.011203f
C1527 vdd.n743 gnd 0.011203f
C1528 vdd.n744 gnd 0.011203f
C1529 vdd.n745 gnd 0.011203f
C1530 vdd.n746 gnd 0.011203f
C1531 vdd.n747 gnd 0.007529f
C1532 vdd.n748 gnd 0.011203f
C1533 vdd.n749 gnd 0.011203f
C1534 vdd.n750 gnd 0.011203f
C1535 vdd.n751 gnd 0.011203f
C1536 vdd.n752 gnd 0.011203f
C1537 vdd.n753 gnd 0.011203f
C1538 vdd.n754 gnd 0.011203f
C1539 vdd.n755 gnd 0.011203f
C1540 vdd.n756 gnd 0.011203f
C1541 vdd.n757 gnd 0.011203f
C1542 vdd.n758 gnd 0.011203f
C1543 vdd.n759 gnd 0.011203f
C1544 vdd.n760 gnd 0.011203f
C1545 vdd.n761 gnd 0.011203f
C1546 vdd.n762 gnd 0.011203f
C1547 vdd.n763 gnd 0.011203f
C1548 vdd.n764 gnd 0.011203f
C1549 vdd.n765 gnd 0.011203f
C1550 vdd.n766 gnd 0.011203f
C1551 vdd.n767 gnd 0.008927f
C1552 vdd.t212 gnd 0.137828f
C1553 vdd.t213 gnd 0.1473f
C1554 vdd.t210 gnd 0.180001f
C1555 vdd.n768 gnd 0.230736f
C1556 vdd.n769 gnd 0.19386f
C1557 vdd.n770 gnd 0.011203f
C1558 vdd.n771 gnd 0.011203f
C1559 vdd.n772 gnd 0.011203f
C1560 vdd.n773 gnd 0.011203f
C1561 vdd.n774 gnd 0.011203f
C1562 vdd.n775 gnd 0.011203f
C1563 vdd.n776 gnd 0.011203f
C1564 vdd.n777 gnd 0.011203f
C1565 vdd.n778 gnd 0.011203f
C1566 vdd.n779 gnd 0.011203f
C1567 vdd.n780 gnd 0.011203f
C1568 vdd.n781 gnd 0.011203f
C1569 vdd.n782 gnd 0.011203f
C1570 vdd.n783 gnd 0.00717f
C1571 vdd.n785 gnd 0.007618f
C1572 vdd.n786 gnd 0.007618f
C1573 vdd.n787 gnd 0.007618f
C1574 vdd.n788 gnd 0.007618f
C1575 vdd.n789 gnd 0.007618f
C1576 vdd.n790 gnd 0.007618f
C1577 vdd.n792 gnd 0.007618f
C1578 vdd.n793 gnd 0.007618f
C1579 vdd.n795 gnd 0.007618f
C1580 vdd.n796 gnd 0.005546f
C1581 vdd.n798 gnd 0.007618f
C1582 vdd.t259 gnd 0.307847f
C1583 vdd.t258 gnd 0.31512f
C1584 vdd.t257 gnd 0.200974f
C1585 vdd.n799 gnd 0.108616f
C1586 vdd.n800 gnd 0.06161f
C1587 vdd.n801 gnd 0.010887f
C1588 vdd.n802 gnd 0.017805f
C1589 vdd.n804 gnd 0.007618f
C1590 vdd.n805 gnd 0.778536f
C1591 vdd.n806 gnd 0.016877f
C1592 vdd.n807 gnd 0.016877f
C1593 vdd.n808 gnd 0.007618f
C1594 vdd.n809 gnd 0.018076f
C1595 vdd.n810 gnd 0.007618f
C1596 vdd.n811 gnd 0.007618f
C1597 vdd.n812 gnd 0.007618f
C1598 vdd.n813 gnd 0.007618f
C1599 vdd.n814 gnd 0.007618f
C1600 vdd.n816 gnd 0.007618f
C1601 vdd.n817 gnd 0.007618f
C1602 vdd.n819 gnd 0.007618f
C1603 vdd.n820 gnd 0.007618f
C1604 vdd.n822 gnd 0.007618f
C1605 vdd.n823 gnd 0.007618f
C1606 vdd.n825 gnd 0.007618f
C1607 vdd.n826 gnd 0.007618f
C1608 vdd.n828 gnd 0.007618f
C1609 vdd.n829 gnd 0.007618f
C1610 vdd.n831 gnd 0.007618f
C1611 vdd.t252 gnd 0.307847f
C1612 vdd.t251 gnd 0.31512f
C1613 vdd.t249 gnd 0.200974f
C1614 vdd.n832 gnd 0.108616f
C1615 vdd.n833 gnd 0.06161f
C1616 vdd.n834 gnd 0.007618f
C1617 vdd.n836 gnd 0.007618f
C1618 vdd.n837 gnd 0.007618f
C1619 vdd.t250 gnd 0.389268f
C1620 vdd.n838 gnd 0.007618f
C1621 vdd.n839 gnd 0.007618f
C1622 vdd.n840 gnd 0.007618f
C1623 vdd.n841 gnd 0.007618f
C1624 vdd.n842 gnd 0.007618f
C1625 vdd.n843 gnd 0.778536f
C1626 vdd.n844 gnd 0.007618f
C1627 vdd.n845 gnd 0.007618f
C1628 vdd.n846 gnd 0.681219f
C1629 vdd.n847 gnd 0.007618f
C1630 vdd.n848 gnd 0.007618f
C1631 vdd.n849 gnd 0.006722f
C1632 vdd.n850 gnd 0.007618f
C1633 vdd.n851 gnd 0.686943f
C1634 vdd.n852 gnd 0.007618f
C1635 vdd.n853 gnd 0.007618f
C1636 vdd.n854 gnd 0.007618f
C1637 vdd.n855 gnd 0.007618f
C1638 vdd.n856 gnd 0.007618f
C1639 vdd.n857 gnd 0.778536f
C1640 vdd.n858 gnd 0.007618f
C1641 vdd.n859 gnd 0.007618f
C1642 vdd.t222 gnd 0.349196f
C1643 vdd.t176 gnd 0.091592f
C1644 vdd.n860 gnd 0.007618f
C1645 vdd.n861 gnd 0.007618f
C1646 vdd.n862 gnd 0.007618f
C1647 vdd.t1 gnd 0.389268f
C1648 vdd.n863 gnd 0.007618f
C1649 vdd.n864 gnd 0.007618f
C1650 vdd.n865 gnd 0.007618f
C1651 vdd.n866 gnd 0.007618f
C1652 vdd.n867 gnd 0.007618f
C1653 vdd.t199 gnd 0.389268f
C1654 vdd.n868 gnd 0.007618f
C1655 vdd.n869 gnd 0.007618f
C1656 vdd.n870 gnd 0.646871f
C1657 vdd.n871 gnd 0.007618f
C1658 vdd.n872 gnd 0.007618f
C1659 vdd.n873 gnd 0.007618f
C1660 vdd.n874 gnd 0.475136f
C1661 vdd.n875 gnd 0.007618f
C1662 vdd.n876 gnd 0.007618f
C1663 vdd.t284 gnd 0.389268f
C1664 vdd.n877 gnd 0.007618f
C1665 vdd.n878 gnd 0.007618f
C1666 vdd.n879 gnd 0.007618f
C1667 vdd.n880 gnd 0.646871f
C1668 vdd.n881 gnd 0.007618f
C1669 vdd.n882 gnd 0.007618f
C1670 vdd.t204 gnd 0.332023f
C1671 vdd.t290 gnd 0.3034f
C1672 vdd.n883 gnd 0.007618f
C1673 vdd.n884 gnd 0.007618f
C1674 vdd.n885 gnd 0.007618f
C1675 vdd.t7 gnd 0.389268f
C1676 vdd.n886 gnd 0.007618f
C1677 vdd.n887 gnd 0.007618f
C1678 vdd.t171 gnd 0.389268f
C1679 vdd.n888 gnd 0.007618f
C1680 vdd.n889 gnd 0.007618f
C1681 vdd.n890 gnd 0.007618f
C1682 vdd.t177 gnd 0.286226f
C1683 vdd.n891 gnd 0.007618f
C1684 vdd.n892 gnd 0.007618f
C1685 vdd.n893 gnd 0.664045f
C1686 vdd.n894 gnd 0.007618f
C1687 vdd.n895 gnd 0.007618f
C1688 vdd.n896 gnd 0.007618f
C1689 vdd.n897 gnd 0.778536f
C1690 vdd.n898 gnd 0.007618f
C1691 vdd.n899 gnd 0.007618f
C1692 vdd.t9 gnd 0.349196f
C1693 vdd.n900 gnd 0.492309f
C1694 vdd.n901 gnd 0.007618f
C1695 vdd.n902 gnd 0.007618f
C1696 vdd.n903 gnd 0.007618f
C1697 vdd.t200 gnd 0.389268f
C1698 vdd.n904 gnd 0.007618f
C1699 vdd.n905 gnd 0.007618f
C1700 vdd.n906 gnd 0.007618f
C1701 vdd.n907 gnd 0.007618f
C1702 vdd.n908 gnd 0.007618f
C1703 vdd.t4 gnd 0.778536f
C1704 vdd.n909 gnd 0.007618f
C1705 vdd.n910 gnd 0.007618f
C1706 vdd.t254 gnd 0.389268f
C1707 vdd.n911 gnd 0.007618f
C1708 vdd.n912 gnd 0.018076f
C1709 vdd.n913 gnd 0.018076f
C1710 vdd.t286 gnd 0.732739f
C1711 vdd.n914 gnd 0.016877f
C1712 vdd.n915 gnd 0.016877f
C1713 vdd.n916 gnd 0.018076f
C1714 vdd.n917 gnd 0.007618f
C1715 vdd.n918 gnd 0.007618f
C1716 vdd.t294 gnd 0.732739f
C1717 vdd.n936 gnd 0.018076f
C1718 vdd.n954 gnd 0.016877f
C1719 vdd.n955 gnd 0.007618f
C1720 vdd.n956 gnd 0.016877f
C1721 vdd.t272 gnd 0.307847f
C1722 vdd.t271 gnd 0.31512f
C1723 vdd.t270 gnd 0.200974f
C1724 vdd.n957 gnd 0.108616f
C1725 vdd.n958 gnd 0.06161f
C1726 vdd.n959 gnd 0.017805f
C1727 vdd.n960 gnd 0.007618f
C1728 vdd.t172 gnd 0.778536f
C1729 vdd.n961 gnd 0.016877f
C1730 vdd.n962 gnd 0.007618f
C1731 vdd.n963 gnd 0.018076f
C1732 vdd.n964 gnd 0.007618f
C1733 vdd.t248 gnd 0.307847f
C1734 vdd.t247 gnd 0.31512f
C1735 vdd.t245 gnd 0.200974f
C1736 vdd.n965 gnd 0.108616f
C1737 vdd.n966 gnd 0.06161f
C1738 vdd.n967 gnd 0.010887f
C1739 vdd.n968 gnd 0.007618f
C1740 vdd.n969 gnd 0.007618f
C1741 vdd.t246 gnd 0.389268f
C1742 vdd.n970 gnd 0.007618f
C1743 vdd.n971 gnd 0.007618f
C1744 vdd.n972 gnd 0.007618f
C1745 vdd.n973 gnd 0.007618f
C1746 vdd.n974 gnd 0.007618f
C1747 vdd.n975 gnd 0.007618f
C1748 vdd.n976 gnd 0.778536f
C1749 vdd.n977 gnd 0.007618f
C1750 vdd.n978 gnd 0.007618f
C1751 vdd.t288 gnd 0.389268f
C1752 vdd.n979 gnd 0.007618f
C1753 vdd.n980 gnd 0.007618f
C1754 vdd.n981 gnd 0.007618f
C1755 vdd.n982 gnd 0.007618f
C1756 vdd.n983 gnd 0.492309f
C1757 vdd.n984 gnd 0.007618f
C1758 vdd.n985 gnd 0.007618f
C1759 vdd.n986 gnd 0.007618f
C1760 vdd.n987 gnd 0.007618f
C1761 vdd.n988 gnd 0.007618f
C1762 vdd.n989 gnd 0.664045f
C1763 vdd.n990 gnd 0.007618f
C1764 vdd.n991 gnd 0.007618f
C1765 vdd.t174 gnd 0.349196f
C1766 vdd.t178 gnd 0.286226f
C1767 vdd.n992 gnd 0.007618f
C1768 vdd.n993 gnd 0.007618f
C1769 vdd.n994 gnd 0.007618f
C1770 vdd.t0 gnd 0.389268f
C1771 vdd.n995 gnd 0.007618f
C1772 vdd.n996 gnd 0.007618f
C1773 vdd.t179 gnd 0.389268f
C1774 vdd.n997 gnd 0.007618f
C1775 vdd.n998 gnd 0.007618f
C1776 vdd.n999 gnd 0.007618f
C1777 vdd.t282 gnd 0.3034f
C1778 vdd.n1000 gnd 0.007618f
C1779 vdd.n1001 gnd 0.007618f
C1780 vdd.n1002 gnd 0.646871f
C1781 vdd.n1003 gnd 0.007618f
C1782 vdd.n1004 gnd 0.007618f
C1783 vdd.n1005 gnd 0.007618f
C1784 vdd.t202 gnd 0.389268f
C1785 vdd.n1006 gnd 0.007618f
C1786 vdd.n1007 gnd 0.007618f
C1787 vdd.t3 gnd 0.332023f
C1788 vdd.n1008 gnd 0.475136f
C1789 vdd.n1009 gnd 0.007618f
C1790 vdd.n1010 gnd 0.007618f
C1791 vdd.n1011 gnd 0.007618f
C1792 vdd.n1012 gnd 0.646871f
C1793 vdd.n1013 gnd 0.007618f
C1794 vdd.n1014 gnd 0.007618f
C1795 vdd.t6 gnd 0.389268f
C1796 vdd.n1015 gnd 0.007618f
C1797 vdd.n1016 gnd 0.007618f
C1798 vdd.n1017 gnd 0.007618f
C1799 vdd.n1018 gnd 0.778536f
C1800 vdd.n1019 gnd 0.007618f
C1801 vdd.n1020 gnd 0.007618f
C1802 vdd.t205 gnd 0.389268f
C1803 vdd.n1021 gnd 0.007618f
C1804 vdd.n1022 gnd 0.007618f
C1805 vdd.n1023 gnd 0.007618f
C1806 vdd.t2 gnd 0.091592f
C1807 vdd.n1024 gnd 0.007618f
C1808 vdd.n1025 gnd 0.007618f
C1809 vdd.n1026 gnd 0.007618f
C1810 vdd.t265 gnd 0.31512f
C1811 vdd.t263 gnd 0.200974f
C1812 vdd.t266 gnd 0.31512f
C1813 vdd.n1027 gnd 0.17711f
C1814 vdd.n1028 gnd 0.007618f
C1815 vdd.n1029 gnd 0.007618f
C1816 vdd.n1030 gnd 0.778536f
C1817 vdd.n1031 gnd 0.007618f
C1818 vdd.n1032 gnd 0.007618f
C1819 vdd.t264 gnd 0.349196f
C1820 vdd.n1033 gnd 0.686943f
C1821 vdd.n1034 gnd 0.007618f
C1822 vdd.n1035 gnd 0.007618f
C1823 vdd.n1036 gnd 0.007618f
C1824 vdd.n1037 gnd 0.681219f
C1825 vdd.n1038 gnd 0.007618f
C1826 vdd.n1039 gnd 0.007618f
C1827 vdd.n1040 gnd 0.007618f
C1828 vdd.n1041 gnd 0.007618f
C1829 vdd.n1042 gnd 0.007618f
C1830 vdd.n1043 gnd 0.778536f
C1831 vdd.n1044 gnd 0.007618f
C1832 vdd.n1045 gnd 0.007618f
C1833 vdd.t207 gnd 0.389268f
C1834 vdd.n1046 gnd 0.007618f
C1835 vdd.n1047 gnd 0.018076f
C1836 vdd.n1048 gnd 0.018076f
C1837 vdd.n1049 gnd 7.8884f
C1838 vdd.n1050 gnd 0.016877f
C1839 vdd.n1051 gnd 0.016877f
C1840 vdd.n1052 gnd 0.018076f
C1841 vdd.n1053 gnd 0.007618f
C1842 vdd.n1054 gnd 0.007618f
C1843 vdd.n1055 gnd 0.007618f
C1844 vdd.n1056 gnd 0.007618f
C1845 vdd.n1057 gnd 0.007618f
C1846 vdd.n1058 gnd 0.007618f
C1847 vdd.n1059 gnd 0.007618f
C1848 vdd.n1060 gnd 0.007618f
C1849 vdd.n1062 gnd 0.007618f
C1850 vdd.n1063 gnd 0.007618f
C1851 vdd.n1064 gnd 0.00717f
C1852 vdd.n1067 gnd 0.027682f
C1853 vdd.n1068 gnd 0.009017f
C1854 vdd.n1069 gnd 0.011203f
C1855 vdd.n1071 gnd 0.011203f
C1856 vdd.n1072 gnd 0.007484f
C1857 vdd.t218 gnd 0.572453f
C1858 vdd.n1073 gnd 8.27767f
C1859 vdd.n1074 gnd 0.011203f
C1860 vdd.n1075 gnd 0.027682f
C1861 vdd.n1076 gnd 0.009017f
C1862 vdd.n1077 gnd 0.011203f
C1863 vdd.n1078 gnd 0.009017f
C1864 vdd.n1079 gnd 0.011203f
C1865 vdd.n1080 gnd 1.14491f
C1866 vdd.n1081 gnd 0.011203f
C1867 vdd.n1082 gnd 0.009017f
C1868 vdd.n1083 gnd 0.009017f
C1869 vdd.n1084 gnd 0.011203f
C1870 vdd.n1085 gnd 0.009017f
C1871 vdd.n1086 gnd 0.011203f
C1872 vdd.t17 gnd 0.572453f
C1873 vdd.n1087 gnd 0.011203f
C1874 vdd.n1088 gnd 0.009017f
C1875 vdd.n1089 gnd 0.011203f
C1876 vdd.n1090 gnd 0.009017f
C1877 vdd.n1091 gnd 0.011203f
C1878 vdd.t148 gnd 0.572453f
C1879 vdd.n1092 gnd 0.011203f
C1880 vdd.n1093 gnd 0.009017f
C1881 vdd.n1094 gnd 0.011203f
C1882 vdd.n1095 gnd 0.009017f
C1883 vdd.n1096 gnd 0.011203f
C1884 vdd.n1097 gnd 0.921649f
C1885 vdd.n1098 gnd 0.950271f
C1886 vdd.t31 gnd 0.572453f
C1887 vdd.n1099 gnd 0.011203f
C1888 vdd.n1100 gnd 0.009017f
C1889 vdd.n1101 gnd 0.011203f
C1890 vdd.n1102 gnd 0.009017f
C1891 vdd.n1103 gnd 0.011203f
C1892 vdd.n1104 gnd 0.727015f
C1893 vdd.n1105 gnd 0.011203f
C1894 vdd.n1106 gnd 0.009017f
C1895 vdd.n1107 gnd 0.011203f
C1896 vdd.n1108 gnd 0.009017f
C1897 vdd.n1109 gnd 0.011203f
C1898 vdd.t19 gnd 0.572453f
C1899 vdd.t62 gnd 0.572453f
C1900 vdd.n1110 gnd 0.011203f
C1901 vdd.n1111 gnd 0.009017f
C1902 vdd.n1112 gnd 0.011203f
C1903 vdd.n1113 gnd 0.009017f
C1904 vdd.n1114 gnd 0.011203f
C1905 vdd.t86 gnd 0.572453f
C1906 vdd.n1115 gnd 0.011203f
C1907 vdd.n1116 gnd 0.009017f
C1908 vdd.n1117 gnd 0.011203f
C1909 vdd.n1118 gnd 0.009017f
C1910 vdd.n1119 gnd 0.011203f
C1911 vdd.t124 gnd 0.572453f
C1912 vdd.n1120 gnd 0.807158f
C1913 vdd.n1121 gnd 0.011203f
C1914 vdd.n1122 gnd 0.009017f
C1915 vdd.n1123 gnd 0.011203f
C1916 vdd.n1124 gnd 0.009017f
C1917 vdd.n1125 gnd 0.011203f
C1918 vdd.n1126 gnd 0.898751f
C1919 vdd.n1127 gnd 0.011203f
C1920 vdd.n1128 gnd 0.009017f
C1921 vdd.n1129 gnd 0.011203f
C1922 vdd.n1130 gnd 0.009017f
C1923 vdd.n1131 gnd 0.011203f
C1924 vdd.n1132 gnd 0.704117f
C1925 vdd.t29 gnd 0.572453f
C1926 vdd.n1133 gnd 0.011203f
C1927 vdd.n1134 gnd 0.009017f
C1928 vdd.n1135 gnd 0.011203f
C1929 vdd.n1136 gnd 0.009017f
C1930 vdd.n1137 gnd 0.011203f
C1931 vdd.t39 gnd 0.572453f
C1932 vdd.n1138 gnd 0.011203f
C1933 vdd.n1139 gnd 0.009017f
C1934 vdd.n1140 gnd 0.011203f
C1935 vdd.n1141 gnd 0.009017f
C1936 vdd.n1142 gnd 0.011203f
C1937 vdd.t57 gnd 0.572453f
C1938 vdd.n1143 gnd 0.635422f
C1939 vdd.n1144 gnd 0.011203f
C1940 vdd.n1145 gnd 0.009017f
C1941 vdd.n1146 gnd 0.011203f
C1942 vdd.n1147 gnd 0.009017f
C1943 vdd.n1148 gnd 0.011203f
C1944 vdd.t104 gnd 0.572453f
C1945 vdd.n1149 gnd 0.011203f
C1946 vdd.n1150 gnd 0.009017f
C1947 vdd.n1151 gnd 0.011203f
C1948 vdd.n1152 gnd 0.009017f
C1949 vdd.n1153 gnd 0.011203f
C1950 vdd.n1154 gnd 0.875853f
C1951 vdd.n1155 gnd 0.950271f
C1952 vdd.t106 gnd 0.572453f
C1953 vdd.n1156 gnd 0.011203f
C1954 vdd.n1157 gnd 0.009017f
C1955 vdd.n1158 gnd 0.011203f
C1956 vdd.n1159 gnd 0.009017f
C1957 vdd.n1160 gnd 0.011203f
C1958 vdd.n1161 gnd 0.681219f
C1959 vdd.n1162 gnd 0.011203f
C1960 vdd.n1163 gnd 0.009017f
C1961 vdd.n1164 gnd 0.011203f
C1962 vdd.n1165 gnd 0.009017f
C1963 vdd.n1166 gnd 0.011203f
C1964 vdd.t55 gnd 0.572453f
C1965 vdd.t53 gnd 0.572453f
C1966 vdd.n1167 gnd 0.011203f
C1967 vdd.n1168 gnd 0.009017f
C1968 vdd.n1169 gnd 0.011203f
C1969 vdd.n1170 gnd 0.009017f
C1970 vdd.n1171 gnd 0.011203f
C1971 vdd.t15 gnd 0.572453f
C1972 vdd.n1172 gnd 0.011203f
C1973 vdd.n1173 gnd 0.009017f
C1974 vdd.n1174 gnd 0.011203f
C1975 vdd.n1175 gnd 0.009017f
C1976 vdd.n1176 gnd 0.011203f
C1977 vdd.t21 gnd 0.572453f
C1978 vdd.n1177 gnd 0.852954f
C1979 vdd.n1178 gnd 0.011203f
C1980 vdd.n1179 gnd 0.009017f
C1981 vdd.n1180 gnd 0.011203f
C1982 vdd.n1181 gnd 0.009017f
C1983 vdd.n1182 gnd 0.011203f
C1984 vdd.n1183 gnd 1.14491f
C1985 vdd.n1184 gnd 0.011203f
C1986 vdd.n1185 gnd 0.009017f
C1987 vdd.n1186 gnd 0.027101f
C1988 vdd.n1187 gnd 0.007484f
C1989 vdd.n1188 gnd 0.027101f
C1990 vdd.t226 gnd 0.572453f
C1991 vdd.n1189 gnd 0.027101f
C1992 vdd.n1190 gnd 0.007484f
C1993 vdd.n1191 gnd 0.011203f
C1994 vdd.n1192 gnd 0.009017f
C1995 vdd.n1193 gnd 0.011203f
C1996 vdd.n1224 gnd 0.027682f
C1997 vdd.n1225 gnd 1.68874f
C1998 vdd.n1226 gnd 0.011203f
C1999 vdd.n1227 gnd 0.009017f
C2000 vdd.n1228 gnd 0.011203f
C2001 vdd.n1229 gnd 0.011203f
C2002 vdd.n1230 gnd 0.011203f
C2003 vdd.n1231 gnd 0.011203f
C2004 vdd.n1232 gnd 0.011203f
C2005 vdd.n1233 gnd 0.009017f
C2006 vdd.n1234 gnd 0.011203f
C2007 vdd.n1235 gnd 0.011203f
C2008 vdd.n1236 gnd 0.011203f
C2009 vdd.n1237 gnd 0.011203f
C2010 vdd.n1238 gnd 0.011203f
C2011 vdd.n1239 gnd 0.009017f
C2012 vdd.n1240 gnd 0.011203f
C2013 vdd.n1241 gnd 0.011203f
C2014 vdd.n1242 gnd 0.011203f
C2015 vdd.n1243 gnd 0.011203f
C2016 vdd.n1244 gnd 0.011203f
C2017 vdd.n1245 gnd 0.009017f
C2018 vdd.n1246 gnd 0.011203f
C2019 vdd.n1247 gnd 0.011203f
C2020 vdd.n1248 gnd 0.011203f
C2021 vdd.n1249 gnd 0.011203f
C2022 vdd.n1250 gnd 0.011203f
C2023 vdd.t240 gnd 0.137828f
C2024 vdd.t241 gnd 0.1473f
C2025 vdd.t239 gnd 0.180001f
C2026 vdd.n1251 gnd 0.230736f
C2027 vdd.n1252 gnd 0.194762f
C2028 vdd.n1253 gnd 0.019297f
C2029 vdd.n1254 gnd 0.011203f
C2030 vdd.n1255 gnd 0.011203f
C2031 vdd.n1256 gnd 0.011203f
C2032 vdd.n1257 gnd 0.011203f
C2033 vdd.n1258 gnd 0.011203f
C2034 vdd.n1259 gnd 0.009017f
C2035 vdd.n1260 gnd 0.011203f
C2036 vdd.n1261 gnd 0.011203f
C2037 vdd.n1262 gnd 0.011203f
C2038 vdd.n1263 gnd 0.011203f
C2039 vdd.n1264 gnd 0.011203f
C2040 vdd.n1265 gnd 0.009017f
C2041 vdd.n1266 gnd 0.011203f
C2042 vdd.n1267 gnd 0.011203f
C2043 vdd.n1268 gnd 0.011203f
C2044 vdd.n1269 gnd 0.011203f
C2045 vdd.n1270 gnd 0.011203f
C2046 vdd.n1271 gnd 0.009017f
C2047 vdd.n1272 gnd 0.011203f
C2048 vdd.n1273 gnd 0.011203f
C2049 vdd.n1274 gnd 0.011203f
C2050 vdd.n1275 gnd 0.011203f
C2051 vdd.n1276 gnd 0.011203f
C2052 vdd.n1277 gnd 0.009017f
C2053 vdd.n1278 gnd 0.011203f
C2054 vdd.n1279 gnd 0.011203f
C2055 vdd.n1280 gnd 0.011203f
C2056 vdd.n1281 gnd 0.011203f
C2057 vdd.n1282 gnd 0.011203f
C2058 vdd.n1283 gnd 0.009017f
C2059 vdd.n1284 gnd 0.011203f
C2060 vdd.n1285 gnd 0.011203f
C2061 vdd.n1286 gnd 0.011203f
C2062 vdd.n1287 gnd 0.011203f
C2063 vdd.n1288 gnd 0.009017f
C2064 vdd.n1289 gnd 0.011203f
C2065 vdd.n1290 gnd 0.011203f
C2066 vdd.n1291 gnd 0.011203f
C2067 vdd.n1292 gnd 0.011203f
C2068 vdd.n1293 gnd 0.011203f
C2069 vdd.n1294 gnd 0.009017f
C2070 vdd.n1295 gnd 0.011203f
C2071 vdd.n1296 gnd 0.011203f
C2072 vdd.n1297 gnd 0.011203f
C2073 vdd.n1298 gnd 0.011203f
C2074 vdd.n1299 gnd 0.011203f
C2075 vdd.n1300 gnd 0.009017f
C2076 vdd.n1301 gnd 0.011203f
C2077 vdd.n1302 gnd 0.011203f
C2078 vdd.n1303 gnd 0.011203f
C2079 vdd.n1304 gnd 0.011203f
C2080 vdd.n1305 gnd 0.011203f
C2081 vdd.n1306 gnd 0.009017f
C2082 vdd.n1307 gnd 0.011203f
C2083 vdd.n1308 gnd 0.011203f
C2084 vdd.n1309 gnd 0.011203f
C2085 vdd.n1310 gnd 0.011203f
C2086 vdd.n1311 gnd 0.011203f
C2087 vdd.n1312 gnd 0.009017f
C2088 vdd.n1313 gnd 0.011203f
C2089 vdd.n1314 gnd 0.011203f
C2090 vdd.n1315 gnd 0.011203f
C2091 vdd.n1316 gnd 0.011203f
C2092 vdd.t237 gnd 0.137828f
C2093 vdd.t238 gnd 0.1473f
C2094 vdd.t236 gnd 0.180001f
C2095 vdd.n1317 gnd 0.230736f
C2096 vdd.n1318 gnd 0.194762f
C2097 vdd.n1319 gnd 0.014788f
C2098 vdd.n1320 gnd 0.004283f
C2099 vdd.n1321 gnd 0.027682f
C2100 vdd.n1322 gnd 0.011203f
C2101 vdd.n1323 gnd 0.004734f
C2102 vdd.n1324 gnd 0.009017f
C2103 vdd.n1325 gnd 0.009017f
C2104 vdd.n1326 gnd 0.011203f
C2105 vdd.n1327 gnd 0.011203f
C2106 vdd.n1328 gnd 0.011203f
C2107 vdd.n1329 gnd 0.009017f
C2108 vdd.n1330 gnd 0.009017f
C2109 vdd.n1331 gnd 0.009017f
C2110 vdd.n1332 gnd 0.011203f
C2111 vdd.n1333 gnd 0.011203f
C2112 vdd.n1334 gnd 0.011203f
C2113 vdd.n1335 gnd 0.009017f
C2114 vdd.n1336 gnd 0.009017f
C2115 vdd.n1337 gnd 0.009017f
C2116 vdd.n1338 gnd 0.011203f
C2117 vdd.n1339 gnd 0.011203f
C2118 vdd.n1340 gnd 0.011203f
C2119 vdd.n1341 gnd 0.009017f
C2120 vdd.n1342 gnd 0.009017f
C2121 vdd.n1343 gnd 0.009017f
C2122 vdd.n1344 gnd 0.011203f
C2123 vdd.n1345 gnd 0.011203f
C2124 vdd.n1346 gnd 0.011203f
C2125 vdd.n1347 gnd 0.009017f
C2126 vdd.n1348 gnd 0.009017f
C2127 vdd.n1349 gnd 0.009017f
C2128 vdd.n1350 gnd 0.011203f
C2129 vdd.n1351 gnd 0.011203f
C2130 vdd.n1352 gnd 0.011203f
C2131 vdd.n1353 gnd 0.008927f
C2132 vdd.n1354 gnd 0.011203f
C2133 vdd.t227 gnd 0.137828f
C2134 vdd.t228 gnd 0.1473f
C2135 vdd.t225 gnd 0.180001f
C2136 vdd.n1355 gnd 0.230736f
C2137 vdd.n1356 gnd 0.194762f
C2138 vdd.n1357 gnd 0.019297f
C2139 vdd.n1358 gnd 0.006132f
C2140 vdd.n1359 gnd 0.011203f
C2141 vdd.n1360 gnd 0.011203f
C2142 vdd.n1361 gnd 0.011203f
C2143 vdd.n1362 gnd 0.009017f
C2144 vdd.n1363 gnd 0.009017f
C2145 vdd.n1364 gnd 0.009017f
C2146 vdd.n1365 gnd 0.011203f
C2147 vdd.n1366 gnd 0.011203f
C2148 vdd.n1367 gnd 0.011203f
C2149 vdd.n1368 gnd 0.009017f
C2150 vdd.n1369 gnd 0.009017f
C2151 vdd.n1370 gnd 0.009017f
C2152 vdd.n1371 gnd 0.011203f
C2153 vdd.n1372 gnd 0.011203f
C2154 vdd.n1373 gnd 0.011203f
C2155 vdd.n1374 gnd 0.009017f
C2156 vdd.n1375 gnd 0.009017f
C2157 vdd.n1376 gnd 0.009017f
C2158 vdd.n1377 gnd 0.011203f
C2159 vdd.n1378 gnd 0.011203f
C2160 vdd.n1379 gnd 0.011203f
C2161 vdd.n1380 gnd 0.009017f
C2162 vdd.n1381 gnd 0.009017f
C2163 vdd.n1382 gnd 0.009017f
C2164 vdd.n1383 gnd 0.011203f
C2165 vdd.n1384 gnd 0.011203f
C2166 vdd.n1385 gnd 0.011203f
C2167 vdd.n1386 gnd 0.009017f
C2168 vdd.n1387 gnd 0.009017f
C2169 vdd.n1388 gnd 0.007529f
C2170 vdd.n1389 gnd 0.011203f
C2171 vdd.n1390 gnd 0.011203f
C2172 vdd.n1391 gnd 0.011203f
C2173 vdd.n1392 gnd 0.007529f
C2174 vdd.n1393 gnd 0.009017f
C2175 vdd.n1394 gnd 0.009017f
C2176 vdd.n1395 gnd 0.011203f
C2177 vdd.n1396 gnd 0.011203f
C2178 vdd.n1397 gnd 0.011203f
C2179 vdd.n1398 gnd 0.009017f
C2180 vdd.n1399 gnd 0.009017f
C2181 vdd.n1400 gnd 0.009017f
C2182 vdd.n1401 gnd 0.011203f
C2183 vdd.n1402 gnd 0.011203f
C2184 vdd.n1403 gnd 0.011203f
C2185 vdd.n1404 gnd 0.009017f
C2186 vdd.n1405 gnd 0.009017f
C2187 vdd.n1406 gnd 0.009017f
C2188 vdd.n1407 gnd 0.011203f
C2189 vdd.n1408 gnd 0.011203f
C2190 vdd.n1409 gnd 0.011203f
C2191 vdd.n1410 gnd 0.009017f
C2192 vdd.n1411 gnd 0.009017f
C2193 vdd.n1412 gnd 0.009017f
C2194 vdd.n1413 gnd 0.011203f
C2195 vdd.n1414 gnd 0.011203f
C2196 vdd.n1415 gnd 0.011203f
C2197 vdd.n1416 gnd 0.009017f
C2198 vdd.n1417 gnd 0.011203f
C2199 vdd.n1418 gnd 2.71343f
C2200 vdd.n1420 gnd 0.027682f
C2201 vdd.n1421 gnd 0.007484f
C2202 vdd.n1422 gnd 0.027682f
C2203 vdd.n1423 gnd 0.027101f
C2204 vdd.n1424 gnd 0.011203f
C2205 vdd.n1425 gnd 0.009017f
C2206 vdd.n1426 gnd 0.011203f
C2207 vdd.n1427 gnd 0.578177f
C2208 vdd.n1428 gnd 0.011203f
C2209 vdd.n1429 gnd 0.009017f
C2210 vdd.n1430 gnd 0.011203f
C2211 vdd.n1431 gnd 0.011203f
C2212 vdd.n1432 gnd 0.011203f
C2213 vdd.n1433 gnd 0.009017f
C2214 vdd.n1434 gnd 0.011203f
C2215 vdd.n1435 gnd 1.04759f
C2216 vdd.n1436 gnd 1.14491f
C2217 vdd.n1437 gnd 0.011203f
C2218 vdd.n1438 gnd 0.009017f
C2219 vdd.n1439 gnd 0.011203f
C2220 vdd.n1440 gnd 0.011203f
C2221 vdd.n1441 gnd 0.011203f
C2222 vdd.n1442 gnd 0.009017f
C2223 vdd.n1443 gnd 0.011203f
C2224 vdd.n1444 gnd 0.66977f
C2225 vdd.n1445 gnd 0.011203f
C2226 vdd.n1446 gnd 0.009017f
C2227 vdd.n1447 gnd 0.011203f
C2228 vdd.n1448 gnd 0.011203f
C2229 vdd.n1449 gnd 0.011203f
C2230 vdd.n1450 gnd 0.009017f
C2231 vdd.n1451 gnd 0.011203f
C2232 vdd.n1452 gnd 0.658321f
C2233 vdd.n1453 gnd 0.864404f
C2234 vdd.n1454 gnd 0.011203f
C2235 vdd.n1455 gnd 0.009017f
C2236 vdd.n1456 gnd 0.011203f
C2237 vdd.n1457 gnd 0.011203f
C2238 vdd.n1458 gnd 0.011203f
C2239 vdd.n1459 gnd 0.009017f
C2240 vdd.n1460 gnd 0.011203f
C2241 vdd.n1461 gnd 0.950271f
C2242 vdd.n1462 gnd 0.011203f
C2243 vdd.n1463 gnd 0.009017f
C2244 vdd.n1464 gnd 0.011203f
C2245 vdd.n1465 gnd 0.011203f
C2246 vdd.n1466 gnd 0.011203f
C2247 vdd.n1467 gnd 0.009017f
C2248 vdd.n1468 gnd 0.011203f
C2249 vdd.t27 gnd 0.572453f
C2250 vdd.n1469 gnd 0.841505f
C2251 vdd.n1470 gnd 0.011203f
C2252 vdd.n1471 gnd 0.009017f
C2253 vdd.n1472 gnd 0.011203f
C2254 vdd.n1473 gnd 0.011203f
C2255 vdd.n1474 gnd 0.011203f
C2256 vdd.n1475 gnd 0.009017f
C2257 vdd.n1476 gnd 0.011203f
C2258 vdd.n1477 gnd 0.646871f
C2259 vdd.n1478 gnd 0.011203f
C2260 vdd.n1479 gnd 0.009017f
C2261 vdd.n1480 gnd 0.011203f
C2262 vdd.n1481 gnd 0.011203f
C2263 vdd.n1482 gnd 0.011203f
C2264 vdd.n1483 gnd 0.009017f
C2265 vdd.n1484 gnd 0.011203f
C2266 vdd.n1485 gnd 0.830056f
C2267 vdd.n1486 gnd 0.692668f
C2268 vdd.n1487 gnd 0.011203f
C2269 vdd.n1488 gnd 0.009017f
C2270 vdd.n1489 gnd 0.011203f
C2271 vdd.n1490 gnd 0.011203f
C2272 vdd.n1491 gnd 0.011203f
C2273 vdd.n1492 gnd 0.009017f
C2274 vdd.n1493 gnd 0.011203f
C2275 vdd.n1494 gnd 0.887302f
C2276 vdd.n1495 gnd 0.011203f
C2277 vdd.n1496 gnd 0.009017f
C2278 vdd.n1497 gnd 0.011203f
C2279 vdd.n1498 gnd 0.011203f
C2280 vdd.n1499 gnd 0.011203f
C2281 vdd.n1500 gnd 0.009017f
C2282 vdd.n1501 gnd 0.011203f
C2283 vdd.t76 gnd 0.572453f
C2284 vdd.n1502 gnd 0.950271f
C2285 vdd.n1503 gnd 0.011203f
C2286 vdd.n1504 gnd 0.009017f
C2287 vdd.n1505 gnd 0.011203f
C2288 vdd.n1506 gnd 0.00861f
C2289 vdd.n1507 gnd 0.006148f
C2290 vdd.n1508 gnd 0.005705f
C2291 vdd.n1509 gnd 0.003156f
C2292 vdd.n1510 gnd 0.007247f
C2293 vdd.n1511 gnd 0.003066f
C2294 vdd.n1512 gnd 0.003246f
C2295 vdd.n1513 gnd 0.005705f
C2296 vdd.n1514 gnd 0.003066f
C2297 vdd.n1515 gnd 0.007247f
C2298 vdd.n1516 gnd 0.003246f
C2299 vdd.n1517 gnd 0.005705f
C2300 vdd.n1518 gnd 0.003066f
C2301 vdd.n1519 gnd 0.005435f
C2302 vdd.n1520 gnd 0.005451f
C2303 vdd.t18 gnd 0.015569f
C2304 vdd.n1521 gnd 0.03464f
C2305 vdd.n1522 gnd 0.180273f
C2306 vdd.n1523 gnd 0.003066f
C2307 vdd.n1524 gnd 0.003246f
C2308 vdd.n1525 gnd 0.007247f
C2309 vdd.n1526 gnd 0.007247f
C2310 vdd.n1527 gnd 0.003246f
C2311 vdd.n1528 gnd 0.003066f
C2312 vdd.n1529 gnd 0.005705f
C2313 vdd.n1530 gnd 0.005705f
C2314 vdd.n1531 gnd 0.003066f
C2315 vdd.n1532 gnd 0.003246f
C2316 vdd.n1533 gnd 0.007247f
C2317 vdd.n1534 gnd 0.007247f
C2318 vdd.n1535 gnd 0.003246f
C2319 vdd.n1536 gnd 0.003066f
C2320 vdd.n1537 gnd 0.005705f
C2321 vdd.n1538 gnd 0.005705f
C2322 vdd.n1539 gnd 0.003066f
C2323 vdd.n1540 gnd 0.003246f
C2324 vdd.n1541 gnd 0.007247f
C2325 vdd.n1542 gnd 0.007247f
C2326 vdd.n1543 gnd 0.017132f
C2327 vdd.n1544 gnd 0.003156f
C2328 vdd.n1545 gnd 0.003066f
C2329 vdd.n1546 gnd 0.014747f
C2330 vdd.n1547 gnd 0.010295f
C2331 vdd.t96 gnd 0.036069f
C2332 vdd.t156 gnd 0.036069f
C2333 vdd.n1548 gnd 0.247888f
C2334 vdd.n1549 gnd 0.194926f
C2335 vdd.t63 gnd 0.036069f
C2336 vdd.t135 gnd 0.036069f
C2337 vdd.n1550 gnd 0.247888f
C2338 vdd.n1551 gnd 0.157304f
C2339 vdd.t87 gnd 0.036069f
C2340 vdd.t144 gnd 0.036069f
C2341 vdd.n1552 gnd 0.247888f
C2342 vdd.n1553 gnd 0.157304f
C2343 vdd.t110 gnd 0.036069f
C2344 vdd.t164 gnd 0.036069f
C2345 vdd.n1554 gnd 0.247888f
C2346 vdd.n1555 gnd 0.157304f
C2347 vdd.t77 gnd 0.036069f
C2348 vdd.t30 gnd 0.036069f
C2349 vdd.n1556 gnd 0.247888f
C2350 vdd.n1557 gnd 0.157304f
C2351 vdd.t99 gnd 0.036069f
C2352 vdd.t40 gnd 0.036069f
C2353 vdd.n1558 gnd 0.247888f
C2354 vdd.n1559 gnd 0.157304f
C2355 vdd.t152 gnd 0.036069f
C2356 vdd.t169 gnd 0.036069f
C2357 vdd.n1560 gnd 0.247888f
C2358 vdd.n1561 gnd 0.157304f
C2359 vdd.t123 gnd 0.036069f
C2360 vdd.t44 gnd 0.036069f
C2361 vdd.n1562 gnd 0.247888f
C2362 vdd.n1563 gnd 0.157304f
C2363 vdd.t111 gnd 0.036069f
C2364 vdd.t56 gnd 0.036069f
C2365 vdd.n1564 gnd 0.247888f
C2366 vdd.n1565 gnd 0.157304f
C2367 vdd.n1566 gnd 0.006148f
C2368 vdd.n1567 gnd 0.005705f
C2369 vdd.n1568 gnd 0.003156f
C2370 vdd.n1569 gnd 0.007247f
C2371 vdd.n1570 gnd 0.003066f
C2372 vdd.n1571 gnd 0.003246f
C2373 vdd.n1572 gnd 0.005705f
C2374 vdd.n1573 gnd 0.003066f
C2375 vdd.n1574 gnd 0.007247f
C2376 vdd.n1575 gnd 0.003246f
C2377 vdd.n1576 gnd 0.005705f
C2378 vdd.n1577 gnd 0.003066f
C2379 vdd.n1578 gnd 0.005435f
C2380 vdd.n1579 gnd 0.005451f
C2381 vdd.t81 gnd 0.015569f
C2382 vdd.n1580 gnd 0.03464f
C2383 vdd.n1581 gnd 0.180273f
C2384 vdd.n1582 gnd 0.003066f
C2385 vdd.n1583 gnd 0.003246f
C2386 vdd.n1584 gnd 0.007247f
C2387 vdd.n1585 gnd 0.007247f
C2388 vdd.n1586 gnd 0.003246f
C2389 vdd.n1587 gnd 0.003066f
C2390 vdd.n1588 gnd 0.005705f
C2391 vdd.n1589 gnd 0.005705f
C2392 vdd.n1590 gnd 0.003066f
C2393 vdd.n1591 gnd 0.003246f
C2394 vdd.n1592 gnd 0.007247f
C2395 vdd.n1593 gnd 0.007247f
C2396 vdd.n1594 gnd 0.003246f
C2397 vdd.n1595 gnd 0.003066f
C2398 vdd.n1596 gnd 0.005705f
C2399 vdd.n1597 gnd 0.005705f
C2400 vdd.n1598 gnd 0.003066f
C2401 vdd.n1599 gnd 0.003246f
C2402 vdd.n1600 gnd 0.007247f
C2403 vdd.n1601 gnd 0.007247f
C2404 vdd.n1602 gnd 0.017132f
C2405 vdd.n1603 gnd 0.003156f
C2406 vdd.n1604 gnd 0.003066f
C2407 vdd.n1605 gnd 0.014747f
C2408 vdd.n1606 gnd 0.009972f
C2409 vdd.n1607 gnd 0.117035f
C2410 vdd.n1608 gnd 0.006148f
C2411 vdd.n1609 gnd 0.005705f
C2412 vdd.n1610 gnd 0.003156f
C2413 vdd.n1611 gnd 0.007247f
C2414 vdd.n1612 gnd 0.003066f
C2415 vdd.n1613 gnd 0.003246f
C2416 vdd.n1614 gnd 0.005705f
C2417 vdd.n1615 gnd 0.003066f
C2418 vdd.n1616 gnd 0.007247f
C2419 vdd.n1617 gnd 0.003246f
C2420 vdd.n1618 gnd 0.005705f
C2421 vdd.n1619 gnd 0.003066f
C2422 vdd.n1620 gnd 0.005435f
C2423 vdd.n1621 gnd 0.005451f
C2424 vdd.t146 gnd 0.015569f
C2425 vdd.n1622 gnd 0.03464f
C2426 vdd.n1623 gnd 0.180273f
C2427 vdd.n1624 gnd 0.003066f
C2428 vdd.n1625 gnd 0.003246f
C2429 vdd.n1626 gnd 0.007247f
C2430 vdd.n1627 gnd 0.007247f
C2431 vdd.n1628 gnd 0.003246f
C2432 vdd.n1629 gnd 0.003066f
C2433 vdd.n1630 gnd 0.005705f
C2434 vdd.n1631 gnd 0.005705f
C2435 vdd.n1632 gnd 0.003066f
C2436 vdd.n1633 gnd 0.003246f
C2437 vdd.n1634 gnd 0.007247f
C2438 vdd.n1635 gnd 0.007247f
C2439 vdd.n1636 gnd 0.003246f
C2440 vdd.n1637 gnd 0.003066f
C2441 vdd.n1638 gnd 0.005705f
C2442 vdd.n1639 gnd 0.005705f
C2443 vdd.n1640 gnd 0.003066f
C2444 vdd.n1641 gnd 0.003246f
C2445 vdd.n1642 gnd 0.007247f
C2446 vdd.n1643 gnd 0.007247f
C2447 vdd.n1644 gnd 0.017132f
C2448 vdd.n1645 gnd 0.003156f
C2449 vdd.n1646 gnd 0.003066f
C2450 vdd.n1647 gnd 0.014747f
C2451 vdd.n1648 gnd 0.010295f
C2452 vdd.t32 gnd 0.036069f
C2453 vdd.t149 gnd 0.036069f
C2454 vdd.n1649 gnd 0.247888f
C2455 vdd.n1650 gnd 0.194926f
C2456 vdd.t142 gnd 0.036069f
C2457 vdd.t127 gnd 0.036069f
C2458 vdd.n1651 gnd 0.247888f
C2459 vdd.n1652 gnd 0.157304f
C2460 vdd.t89 gnd 0.036069f
C2461 vdd.t20 gnd 0.036069f
C2462 vdd.n1653 gnd 0.247888f
C2463 vdd.n1654 gnd 0.157304f
C2464 vdd.t159 gnd 0.036069f
C2465 vdd.t125 gnd 0.036069f
C2466 vdd.n1655 gnd 0.247888f
C2467 vdd.n1656 gnd 0.157304f
C2468 vdd.t119 gnd 0.036069f
C2469 vdd.t64 gnd 0.036069f
C2470 vdd.n1657 gnd 0.247888f
C2471 vdd.n1658 gnd 0.157304f
C2472 vdd.t58 gnd 0.036069f
C2473 vdd.t120 gnd 0.036069f
C2474 vdd.n1659 gnd 0.247888f
C2475 vdd.n1660 gnd 0.157304f
C2476 vdd.t107 gnd 0.036069f
C2477 vdd.t105 gnd 0.036069f
C2478 vdd.n1661 gnd 0.247888f
C2479 vdd.n1662 gnd 0.157304f
C2480 vdd.t54 gnd 0.036069f
C2481 vdd.t28 gnd 0.036069f
C2482 vdd.n1663 gnd 0.247888f
C2483 vdd.n1664 gnd 0.157304f
C2484 vdd.t16 gnd 0.036069f
C2485 vdd.t100 gnd 0.036069f
C2486 vdd.n1665 gnd 0.247888f
C2487 vdd.n1666 gnd 0.157304f
C2488 vdd.n1667 gnd 0.006148f
C2489 vdd.n1668 gnd 0.005705f
C2490 vdd.n1669 gnd 0.003156f
C2491 vdd.n1670 gnd 0.007247f
C2492 vdd.n1671 gnd 0.003066f
C2493 vdd.n1672 gnd 0.003246f
C2494 vdd.n1673 gnd 0.005705f
C2495 vdd.n1674 gnd 0.003066f
C2496 vdd.n1675 gnd 0.007247f
C2497 vdd.n1676 gnd 0.003246f
C2498 vdd.n1677 gnd 0.005705f
C2499 vdd.n1678 gnd 0.003066f
C2500 vdd.n1679 gnd 0.005435f
C2501 vdd.n1680 gnd 0.005451f
C2502 vdd.t22 gnd 0.015569f
C2503 vdd.n1681 gnd 0.03464f
C2504 vdd.n1682 gnd 0.180273f
C2505 vdd.n1683 gnd 0.003066f
C2506 vdd.n1684 gnd 0.003246f
C2507 vdd.n1685 gnd 0.007247f
C2508 vdd.n1686 gnd 0.007247f
C2509 vdd.n1687 gnd 0.003246f
C2510 vdd.n1688 gnd 0.003066f
C2511 vdd.n1689 gnd 0.005705f
C2512 vdd.n1690 gnd 0.005705f
C2513 vdd.n1691 gnd 0.003066f
C2514 vdd.n1692 gnd 0.003246f
C2515 vdd.n1693 gnd 0.007247f
C2516 vdd.n1694 gnd 0.007247f
C2517 vdd.n1695 gnd 0.003246f
C2518 vdd.n1696 gnd 0.003066f
C2519 vdd.n1697 gnd 0.005705f
C2520 vdd.n1698 gnd 0.005705f
C2521 vdd.n1699 gnd 0.003066f
C2522 vdd.n1700 gnd 0.003246f
C2523 vdd.n1701 gnd 0.007247f
C2524 vdd.n1702 gnd 0.007247f
C2525 vdd.n1703 gnd 0.017132f
C2526 vdd.n1704 gnd 0.003156f
C2527 vdd.n1705 gnd 0.003066f
C2528 vdd.n1706 gnd 0.014747f
C2529 vdd.n1707 gnd 0.009972f
C2530 vdd.n1708 gnd 0.069624f
C2531 vdd.n1709 gnd 0.250874f
C2532 vdd.n1710 gnd 0.006148f
C2533 vdd.n1711 gnd 0.005705f
C2534 vdd.n1712 gnd 0.003156f
C2535 vdd.n1713 gnd 0.007247f
C2536 vdd.n1714 gnd 0.003066f
C2537 vdd.n1715 gnd 0.003246f
C2538 vdd.n1716 gnd 0.005705f
C2539 vdd.n1717 gnd 0.003066f
C2540 vdd.n1718 gnd 0.007247f
C2541 vdd.n1719 gnd 0.003246f
C2542 vdd.n1720 gnd 0.005705f
C2543 vdd.n1721 gnd 0.003066f
C2544 vdd.n1722 gnd 0.005435f
C2545 vdd.n1723 gnd 0.005451f
C2546 vdd.t160 gnd 0.015569f
C2547 vdd.n1724 gnd 0.03464f
C2548 vdd.n1725 gnd 0.180273f
C2549 vdd.n1726 gnd 0.003066f
C2550 vdd.n1727 gnd 0.003246f
C2551 vdd.n1728 gnd 0.007247f
C2552 vdd.n1729 gnd 0.007247f
C2553 vdd.n1730 gnd 0.003246f
C2554 vdd.n1731 gnd 0.003066f
C2555 vdd.n1732 gnd 0.005705f
C2556 vdd.n1733 gnd 0.005705f
C2557 vdd.n1734 gnd 0.003066f
C2558 vdd.n1735 gnd 0.003246f
C2559 vdd.n1736 gnd 0.007247f
C2560 vdd.n1737 gnd 0.007247f
C2561 vdd.n1738 gnd 0.003246f
C2562 vdd.n1739 gnd 0.003066f
C2563 vdd.n1740 gnd 0.005705f
C2564 vdd.n1741 gnd 0.005705f
C2565 vdd.n1742 gnd 0.003066f
C2566 vdd.n1743 gnd 0.003246f
C2567 vdd.n1744 gnd 0.007247f
C2568 vdd.n1745 gnd 0.007247f
C2569 vdd.n1746 gnd 0.017132f
C2570 vdd.n1747 gnd 0.003156f
C2571 vdd.n1748 gnd 0.003066f
C2572 vdd.n1749 gnd 0.014747f
C2573 vdd.n1750 gnd 0.010295f
C2574 vdd.t50 gnd 0.036069f
C2575 vdd.t161 gnd 0.036069f
C2576 vdd.n1751 gnd 0.247888f
C2577 vdd.n1752 gnd 0.194926f
C2578 vdd.t158 gnd 0.036069f
C2579 vdd.t139 gnd 0.036069f
C2580 vdd.n1753 gnd 0.247888f
C2581 vdd.n1754 gnd 0.157304f
C2582 vdd.t108 gnd 0.036069f
C2583 vdd.t46 gnd 0.036069f
C2584 vdd.n1755 gnd 0.247888f
C2585 vdd.n1756 gnd 0.157304f
C2586 vdd.t170 gnd 0.036069f
C2587 vdd.t136 gnd 0.036069f
C2588 vdd.n1757 gnd 0.247888f
C2589 vdd.n1758 gnd 0.157304f
C2590 vdd.t133 gnd 0.036069f
C2591 vdd.t82 gnd 0.036069f
C2592 vdd.n1759 gnd 0.247888f
C2593 vdd.n1760 gnd 0.157304f
C2594 vdd.t78 gnd 0.036069f
C2595 vdd.t134 gnd 0.036069f
C2596 vdd.n1761 gnd 0.247888f
C2597 vdd.n1762 gnd 0.157304f
C2598 vdd.t118 gnd 0.036069f
C2599 vdd.t117 gnd 0.036069f
C2600 vdd.n1763 gnd 0.247888f
C2601 vdd.n1764 gnd 0.157304f
C2602 vdd.t75 gnd 0.036069f
C2603 vdd.t49 gnd 0.036069f
C2604 vdd.n1765 gnd 0.247888f
C2605 vdd.n1766 gnd 0.157304f
C2606 vdd.t45 gnd 0.036069f
C2607 vdd.t114 gnd 0.036069f
C2608 vdd.n1767 gnd 0.247888f
C2609 vdd.n1768 gnd 0.157304f
C2610 vdd.n1769 gnd 0.006148f
C2611 vdd.n1770 gnd 0.005705f
C2612 vdd.n1771 gnd 0.003156f
C2613 vdd.n1772 gnd 0.007247f
C2614 vdd.n1773 gnd 0.003066f
C2615 vdd.n1774 gnd 0.003246f
C2616 vdd.n1775 gnd 0.005705f
C2617 vdd.n1776 gnd 0.003066f
C2618 vdd.n1777 gnd 0.007247f
C2619 vdd.n1778 gnd 0.003246f
C2620 vdd.n1779 gnd 0.005705f
C2621 vdd.n1780 gnd 0.003066f
C2622 vdd.n1781 gnd 0.005435f
C2623 vdd.n1782 gnd 0.005451f
C2624 vdd.t47 gnd 0.015569f
C2625 vdd.n1783 gnd 0.03464f
C2626 vdd.n1784 gnd 0.180273f
C2627 vdd.n1785 gnd 0.003066f
C2628 vdd.n1786 gnd 0.003246f
C2629 vdd.n1787 gnd 0.007247f
C2630 vdd.n1788 gnd 0.007247f
C2631 vdd.n1789 gnd 0.003246f
C2632 vdd.n1790 gnd 0.003066f
C2633 vdd.n1791 gnd 0.005705f
C2634 vdd.n1792 gnd 0.005705f
C2635 vdd.n1793 gnd 0.003066f
C2636 vdd.n1794 gnd 0.003246f
C2637 vdd.n1795 gnd 0.007247f
C2638 vdd.n1796 gnd 0.007247f
C2639 vdd.n1797 gnd 0.003246f
C2640 vdd.n1798 gnd 0.003066f
C2641 vdd.n1799 gnd 0.005705f
C2642 vdd.n1800 gnd 0.005705f
C2643 vdd.n1801 gnd 0.003066f
C2644 vdd.n1802 gnd 0.003246f
C2645 vdd.n1803 gnd 0.007247f
C2646 vdd.n1804 gnd 0.007247f
C2647 vdd.n1805 gnd 0.017132f
C2648 vdd.n1806 gnd 0.003156f
C2649 vdd.n1807 gnd 0.003066f
C2650 vdd.n1808 gnd 0.014747f
C2651 vdd.n1809 gnd 0.009972f
C2652 vdd.n1810 gnd 0.069624f
C2653 vdd.n1811 gnd 0.287196f
C2654 vdd.n1812 gnd 2.87741f
C2655 vdd.n1813 gnd 0.660802f
C2656 vdd.n1814 gnd 0.00861f
C2657 vdd.n1815 gnd 0.009017f
C2658 vdd.n1816 gnd 0.011203f
C2659 vdd.n1817 gnd 0.818607f
C2660 vdd.n1818 gnd 0.011203f
C2661 vdd.n1819 gnd 0.009017f
C2662 vdd.n1820 gnd 0.011203f
C2663 vdd.n1821 gnd 0.011203f
C2664 vdd.n1822 gnd 0.011203f
C2665 vdd.n1823 gnd 0.009017f
C2666 vdd.n1824 gnd 0.011203f
C2667 vdd.n1825 gnd 0.950271f
C2668 vdd.t109 gnd 0.572453f
C2669 vdd.n1826 gnd 0.623973f
C2670 vdd.n1827 gnd 0.011203f
C2671 vdd.n1828 gnd 0.009017f
C2672 vdd.n1829 gnd 0.011203f
C2673 vdd.n1830 gnd 0.011203f
C2674 vdd.n1831 gnd 0.011203f
C2675 vdd.n1832 gnd 0.009017f
C2676 vdd.n1833 gnd 0.011203f
C2677 vdd.n1834 gnd 0.715566f
C2678 vdd.n1835 gnd 0.011203f
C2679 vdd.n1836 gnd 0.009017f
C2680 vdd.n1837 gnd 0.011203f
C2681 vdd.n1838 gnd 0.011203f
C2682 vdd.n1839 gnd 0.011203f
C2683 vdd.n1840 gnd 0.009017f
C2684 vdd.n1841 gnd 0.011203f
C2685 vdd.n1842 gnd 0.612524f
C2686 vdd.n1843 gnd 0.9102f
C2687 vdd.n1844 gnd 0.011203f
C2688 vdd.n1845 gnd 0.009017f
C2689 vdd.n1846 gnd 0.011203f
C2690 vdd.n1847 gnd 0.011203f
C2691 vdd.n1848 gnd 0.011203f
C2692 vdd.n1849 gnd 0.009017f
C2693 vdd.n1850 gnd 0.011203f
C2694 vdd.n1851 gnd 0.950271f
C2695 vdd.n1852 gnd 0.011203f
C2696 vdd.n1853 gnd 0.009017f
C2697 vdd.n1854 gnd 0.011203f
C2698 vdd.n1855 gnd 0.011203f
C2699 vdd.n1856 gnd 0.011203f
C2700 vdd.n1857 gnd 0.009017f
C2701 vdd.n1858 gnd 0.011203f
C2702 vdd.t126 gnd 0.572453f
C2703 vdd.n1859 gnd 0.795709f
C2704 vdd.n1860 gnd 0.011203f
C2705 vdd.n1861 gnd 0.009017f
C2706 vdd.n1862 gnd 0.011203f
C2707 vdd.n1863 gnd 0.011203f
C2708 vdd.n1864 gnd 0.011203f
C2709 vdd.n1865 gnd 0.009017f
C2710 vdd.n1866 gnd 0.011203f
C2711 vdd.n1867 gnd 0.601075f
C2712 vdd.n1868 gnd 0.011203f
C2713 vdd.n1869 gnd 0.009017f
C2714 vdd.n1870 gnd 0.011203f
C2715 vdd.n1871 gnd 0.011203f
C2716 vdd.n1872 gnd 0.011203f
C2717 vdd.n1873 gnd 0.009017f
C2718 vdd.n1874 gnd 0.011203f
C2719 vdd.n1875 gnd 0.78426f
C2720 vdd.n1876 gnd 0.738464f
C2721 vdd.n1877 gnd 0.011203f
C2722 vdd.n1878 gnd 0.009017f
C2723 vdd.n1879 gnd 0.011203f
C2724 vdd.n1880 gnd 0.011203f
C2725 vdd.n1881 gnd 0.011203f
C2726 vdd.n1882 gnd 0.009017f
C2727 vdd.n1883 gnd 0.011203f
C2728 vdd.n1884 gnd 0.933098f
C2729 vdd.n1885 gnd 0.011203f
C2730 vdd.n1886 gnd 0.009017f
C2731 vdd.n1887 gnd 0.011203f
C2732 vdd.n1888 gnd 0.011203f
C2733 vdd.n1889 gnd 0.027101f
C2734 vdd.n1890 gnd 0.011203f
C2735 vdd.n1891 gnd 0.011203f
C2736 vdd.n1892 gnd 0.009017f
C2737 vdd.n1893 gnd 0.011203f
C2738 vdd.n1894 gnd 0.692668f
C2739 vdd.n1895 gnd 1.14491f
C2740 vdd.n1896 gnd 0.011203f
C2741 vdd.n1897 gnd 0.009017f
C2742 vdd.n1898 gnd 0.011203f
C2743 vdd.n1899 gnd 0.011203f
C2744 vdd.n1900 gnd 0.009635f
C2745 vdd.n1901 gnd 0.009017f
C2746 vdd.n1903 gnd 0.011203f
C2747 vdd.n1905 gnd 0.009017f
C2748 vdd.n1906 gnd 0.011203f
C2749 vdd.n1907 gnd 0.009017f
C2750 vdd.n1909 gnd 0.011203f
C2751 vdd.n1910 gnd 0.009017f
C2752 vdd.n1911 gnd 0.011203f
C2753 vdd.n1912 gnd 0.011203f
C2754 vdd.n1913 gnd 0.011203f
C2755 vdd.n1914 gnd 0.011203f
C2756 vdd.n1915 gnd 0.011203f
C2757 vdd.n1916 gnd 0.009017f
C2758 vdd.n1918 gnd 0.011203f
C2759 vdd.n1919 gnd 0.011203f
C2760 vdd.n1920 gnd 0.011203f
C2761 vdd.n1921 gnd 0.011203f
C2762 vdd.n1922 gnd 0.011203f
C2763 vdd.n1923 gnd 0.009017f
C2764 vdd.n1925 gnd 0.011203f
C2765 vdd.n1926 gnd 0.011203f
C2766 vdd.n1927 gnd 0.011203f
C2767 vdd.n1928 gnd 0.011203f
C2768 vdd.n1929 gnd 0.007529f
C2769 vdd.t244 gnd 0.137828f
C2770 vdd.t243 gnd 0.1473f
C2771 vdd.t242 gnd 0.180001f
C2772 vdd.n1930 gnd 0.230736f
C2773 vdd.n1931 gnd 0.19386f
C2774 vdd.n1933 gnd 0.011203f
C2775 vdd.n1934 gnd 0.011203f
C2776 vdd.n1935 gnd 0.009017f
C2777 vdd.n1936 gnd 0.011203f
C2778 vdd.n1938 gnd 0.011203f
C2779 vdd.n1939 gnd 0.011203f
C2780 vdd.n1940 gnd 0.011203f
C2781 vdd.n1941 gnd 0.011203f
C2782 vdd.n1942 gnd 0.009017f
C2783 vdd.n1944 gnd 0.011203f
C2784 vdd.n1945 gnd 0.011203f
C2785 vdd.n1946 gnd 0.011203f
C2786 vdd.n1947 gnd 0.011203f
C2787 vdd.n1948 gnd 0.011203f
C2788 vdd.n1949 gnd 0.009017f
C2789 vdd.n1951 gnd 0.011203f
C2790 vdd.n1952 gnd 0.011203f
C2791 vdd.n1953 gnd 0.011203f
C2792 vdd.n1954 gnd 0.011203f
C2793 vdd.n1955 gnd 0.011203f
C2794 vdd.n1956 gnd 0.009017f
C2795 vdd.n1958 gnd 0.011203f
C2796 vdd.n1959 gnd 0.011203f
C2797 vdd.n1960 gnd 0.011203f
C2798 vdd.n1961 gnd 0.011203f
C2799 vdd.n1962 gnd 0.011203f
C2800 vdd.n1963 gnd 0.009017f
C2801 vdd.n1965 gnd 0.011203f
C2802 vdd.n1966 gnd 0.011203f
C2803 vdd.n1967 gnd 0.011203f
C2804 vdd.n1968 gnd 0.011203f
C2805 vdd.n1969 gnd 0.008927f
C2806 vdd.t231 gnd 0.137828f
C2807 vdd.t230 gnd 0.1473f
C2808 vdd.t229 gnd 0.180001f
C2809 vdd.n1970 gnd 0.230736f
C2810 vdd.n1971 gnd 0.19386f
C2811 vdd.n1973 gnd 0.011203f
C2812 vdd.n1974 gnd 0.011203f
C2813 vdd.n1975 gnd 0.009017f
C2814 vdd.n1976 gnd 0.011203f
C2815 vdd.n1978 gnd 0.011203f
C2816 vdd.n1979 gnd 0.011203f
C2817 vdd.n1980 gnd 0.011203f
C2818 vdd.n1981 gnd 0.011203f
C2819 vdd.n1982 gnd 0.009017f
C2820 vdd.n1984 gnd 0.011203f
C2821 vdd.n1985 gnd 0.011203f
C2822 vdd.n1986 gnd 0.011203f
C2823 vdd.n1987 gnd 0.011203f
C2824 vdd.n1988 gnd 0.011203f
C2825 vdd.n1989 gnd 0.009017f
C2826 vdd.n1991 gnd 0.011203f
C2827 vdd.n1992 gnd 0.011203f
C2828 vdd.n1993 gnd 0.011203f
C2829 vdd.n1994 gnd 0.011203f
C2830 vdd.n1995 gnd 0.011203f
C2831 vdd.n1996 gnd 0.011203f
C2832 vdd.n1997 gnd 0.009017f
C2833 vdd.n1999 gnd 0.011203f
C2834 vdd.n2001 gnd 0.011203f
C2835 vdd.n2002 gnd 0.009017f
C2836 vdd.n2003 gnd 0.009017f
C2837 vdd.n2004 gnd 0.011203f
C2838 vdd.n2006 gnd 0.011203f
C2839 vdd.n2007 gnd 0.009017f
C2840 vdd.n2008 gnd 0.009017f
C2841 vdd.n2009 gnd 0.011203f
C2842 vdd.n2011 gnd 0.011203f
C2843 vdd.n2012 gnd 0.011203f
C2844 vdd.n2013 gnd 0.009017f
C2845 vdd.n2014 gnd 0.009017f
C2846 vdd.n2015 gnd 0.009017f
C2847 vdd.n2016 gnd 0.011203f
C2848 vdd.n2018 gnd 0.011203f
C2849 vdd.n2019 gnd 0.011203f
C2850 vdd.n2020 gnd 0.009017f
C2851 vdd.n2021 gnd 0.009017f
C2852 vdd.n2022 gnd 0.009017f
C2853 vdd.n2023 gnd 0.011203f
C2854 vdd.n2025 gnd 0.011203f
C2855 vdd.n2026 gnd 0.011203f
C2856 vdd.n2027 gnd 0.009017f
C2857 vdd.n2028 gnd 0.009017f
C2858 vdd.n2029 gnd 0.009017f
C2859 vdd.n2030 gnd 0.011203f
C2860 vdd.n2032 gnd 0.011203f
C2861 vdd.n2033 gnd 0.011203f
C2862 vdd.n2034 gnd 0.009017f
C2863 vdd.n2035 gnd 0.011203f
C2864 vdd.n2036 gnd 0.011203f
C2865 vdd.n2037 gnd 0.011203f
C2866 vdd.n2038 gnd 0.018395f
C2867 vdd.n2039 gnd 0.006132f
C2868 vdd.n2040 gnd 0.009017f
C2869 vdd.n2041 gnd 0.011203f
C2870 vdd.n2043 gnd 0.011203f
C2871 vdd.n2044 gnd 0.011203f
C2872 vdd.n2045 gnd 0.009017f
C2873 vdd.n2046 gnd 0.009017f
C2874 vdd.n2047 gnd 0.009017f
C2875 vdd.n2048 gnd 0.011203f
C2876 vdd.n2050 gnd 0.011203f
C2877 vdd.n2051 gnd 0.011203f
C2878 vdd.n2052 gnd 0.009017f
C2879 vdd.n2053 gnd 0.009017f
C2880 vdd.n2054 gnd 0.009017f
C2881 vdd.n2055 gnd 0.011203f
C2882 vdd.n2057 gnd 0.011203f
C2883 vdd.n2058 gnd 0.011203f
C2884 vdd.n2059 gnd 0.009017f
C2885 vdd.n2060 gnd 0.009017f
C2886 vdd.n2061 gnd 0.009017f
C2887 vdd.n2062 gnd 0.011203f
C2888 vdd.n2064 gnd 0.011203f
C2889 vdd.n2065 gnd 0.011203f
C2890 vdd.n2066 gnd 0.009017f
C2891 vdd.n2067 gnd 0.009017f
C2892 vdd.n2068 gnd 0.009017f
C2893 vdd.n2069 gnd 0.011203f
C2894 vdd.n2071 gnd 0.011203f
C2895 vdd.n2072 gnd 0.011203f
C2896 vdd.n2073 gnd 0.009017f
C2897 vdd.n2074 gnd 0.011203f
C2898 vdd.n2075 gnd 0.011203f
C2899 vdd.n2076 gnd 0.011203f
C2900 vdd.n2077 gnd 0.018395f
C2901 vdd.n2078 gnd 0.007529f
C2902 vdd.n2079 gnd 0.009017f
C2903 vdd.n2080 gnd 0.011203f
C2904 vdd.n2082 gnd 0.011203f
C2905 vdd.n2083 gnd 0.011203f
C2906 vdd.n2084 gnd 0.009017f
C2907 vdd.n2085 gnd 0.009017f
C2908 vdd.n2086 gnd 0.009017f
C2909 vdd.n2087 gnd 0.011203f
C2910 vdd.n2089 gnd 0.011203f
C2911 vdd.n2090 gnd 0.011203f
C2912 vdd.n2091 gnd 0.009017f
C2913 vdd.n2092 gnd 0.009017f
C2914 vdd.n2093 gnd 0.009017f
C2915 vdd.n2094 gnd 0.011203f
C2916 vdd.n2096 gnd 0.011203f
C2917 vdd.n2097 gnd 0.011203f
C2918 vdd.n2099 gnd 0.011203f
C2919 vdd.n2100 gnd 0.009017f
C2920 vdd.n2101 gnd 0.00717f
C2921 vdd.n2102 gnd 0.007618f
C2922 vdd.n2103 gnd 0.007618f
C2923 vdd.n2104 gnd 0.007618f
C2924 vdd.n2105 gnd 0.007618f
C2925 vdd.n2106 gnd 0.007618f
C2926 vdd.n2107 gnd 0.007618f
C2927 vdd.n2108 gnd 0.007618f
C2928 vdd.n2109 gnd 0.007618f
C2929 vdd.n2111 gnd 0.007618f
C2930 vdd.n2112 gnd 0.007618f
C2931 vdd.n2113 gnd 0.007618f
C2932 vdd.n2114 gnd 0.007618f
C2933 vdd.n2115 gnd 0.007618f
C2934 vdd.n2117 gnd 0.007618f
C2935 vdd.n2119 gnd 0.007618f
C2936 vdd.n2120 gnd 0.007618f
C2937 vdd.n2121 gnd 0.007618f
C2938 vdd.n2122 gnd 0.007618f
C2939 vdd.n2123 gnd 0.007618f
C2940 vdd.n2125 gnd 0.007618f
C2941 vdd.n2127 gnd 0.007618f
C2942 vdd.n2128 gnd 0.007618f
C2943 vdd.n2129 gnd 0.007618f
C2944 vdd.n2130 gnd 0.007618f
C2945 vdd.n2131 gnd 0.007618f
C2946 vdd.n2133 gnd 0.007618f
C2947 vdd.n2135 gnd 0.007618f
C2948 vdd.n2136 gnd 0.007618f
C2949 vdd.n2137 gnd 0.007618f
C2950 vdd.n2138 gnd 0.007618f
C2951 vdd.n2139 gnd 0.007618f
C2952 vdd.n2141 gnd 0.007618f
C2953 vdd.n2142 gnd 0.007618f
C2954 vdd.n2143 gnd 0.007618f
C2955 vdd.n2144 gnd 0.007618f
C2956 vdd.n2145 gnd 0.007618f
C2957 vdd.n2146 gnd 0.007618f
C2958 vdd.n2147 gnd 0.007618f
C2959 vdd.n2148 gnd 0.007618f
C2960 vdd.n2149 gnd 0.005546f
C2961 vdd.n2150 gnd 0.007618f
C2962 vdd.t208 gnd 0.307847f
C2963 vdd.t209 gnd 0.31512f
C2964 vdd.t206 gnd 0.200974f
C2965 vdd.n2151 gnd 0.108616f
C2966 vdd.n2152 gnd 0.06161f
C2967 vdd.n2153 gnd 0.010887f
C2968 vdd.n2154 gnd 0.007618f
C2969 vdd.n2155 gnd 0.007618f
C2970 vdd.n2156 gnd 0.463687f
C2971 vdd.n2157 gnd 0.007618f
C2972 vdd.n2158 gnd 0.007618f
C2973 vdd.n2159 gnd 0.007618f
C2974 vdd.n2160 gnd 0.007618f
C2975 vdd.n2161 gnd 0.007618f
C2976 vdd.n2162 gnd 0.007618f
C2977 vdd.n2163 gnd 0.007618f
C2978 vdd.n2164 gnd 0.007618f
C2979 vdd.n2165 gnd 0.007618f
C2980 vdd.n2166 gnd 0.007618f
C2981 vdd.n2167 gnd 0.007618f
C2982 vdd.n2168 gnd 0.007618f
C2983 vdd.n2169 gnd 0.007618f
C2984 vdd.n2170 gnd 0.007618f
C2985 vdd.n2171 gnd 0.007618f
C2986 vdd.n2172 gnd 0.007618f
C2987 vdd.n2173 gnd 0.007618f
C2988 vdd.n2174 gnd 0.007618f
C2989 vdd.n2175 gnd 0.007618f
C2990 vdd.n2176 gnd 0.007618f
C2991 vdd.t261 gnd 0.307847f
C2992 vdd.t262 gnd 0.31512f
C2993 vdd.t260 gnd 0.200974f
C2994 vdd.n2177 gnd 0.108616f
C2995 vdd.n2178 gnd 0.06161f
C2996 vdd.n2179 gnd 0.007618f
C2997 vdd.n2180 gnd 0.007618f
C2998 vdd.n2181 gnd 0.007618f
C2999 vdd.n2182 gnd 0.007618f
C3000 vdd.n2183 gnd 0.007618f
C3001 vdd.n2184 gnd 0.007618f
C3002 vdd.n2186 gnd 0.007618f
C3003 vdd.n2187 gnd 0.007618f
C3004 vdd.n2188 gnd 0.007618f
C3005 vdd.n2189 gnd 0.007618f
C3006 vdd.n2191 gnd 0.007618f
C3007 vdd.n2193 gnd 0.007618f
C3008 vdd.n2194 gnd 0.007618f
C3009 vdd.n2195 gnd 0.007618f
C3010 vdd.n2196 gnd 0.007618f
C3011 vdd.n2197 gnd 0.007618f
C3012 vdd.n2199 gnd 0.007618f
C3013 vdd.n2201 gnd 0.007618f
C3014 vdd.n2202 gnd 0.007618f
C3015 vdd.n2203 gnd 0.007618f
C3016 vdd.n2204 gnd 0.007618f
C3017 vdd.n2205 gnd 0.007618f
C3018 vdd.n2207 gnd 0.007618f
C3019 vdd.n2209 gnd 0.007618f
C3020 vdd.n2210 gnd 0.007618f
C3021 vdd.n2211 gnd 0.005546f
C3022 vdd.n2212 gnd 0.010887f
C3023 vdd.n2213 gnd 0.005882f
C3024 vdd.n2214 gnd 0.007618f
C3025 vdd.n2216 gnd 0.007618f
C3026 vdd.n2217 gnd 0.018076f
C3027 vdd.n2218 gnd 0.018076f
C3028 vdd.n2219 gnd 0.016877f
C3029 vdd.n2220 gnd 0.007618f
C3030 vdd.n2221 gnd 0.007618f
C3031 vdd.n2222 gnd 0.007618f
C3032 vdd.n2223 gnd 0.007618f
C3033 vdd.n2224 gnd 0.007618f
C3034 vdd.n2225 gnd 0.007618f
C3035 vdd.n2226 gnd 0.007618f
C3036 vdd.n2227 gnd 0.007618f
C3037 vdd.n2228 gnd 0.007618f
C3038 vdd.n2229 gnd 0.007618f
C3039 vdd.n2230 gnd 0.007618f
C3040 vdd.n2231 gnd 0.007618f
C3041 vdd.n2232 gnd 0.007618f
C3042 vdd.n2233 gnd 0.007618f
C3043 vdd.n2234 gnd 0.007618f
C3044 vdd.n2235 gnd 0.007618f
C3045 vdd.n2236 gnd 0.007618f
C3046 vdd.n2237 gnd 0.007618f
C3047 vdd.n2238 gnd 0.007618f
C3048 vdd.n2239 gnd 0.007618f
C3049 vdd.n2240 gnd 0.007618f
C3050 vdd.n2241 gnd 0.007618f
C3051 vdd.n2242 gnd 0.007618f
C3052 vdd.n2243 gnd 0.007618f
C3053 vdd.n2244 gnd 0.007618f
C3054 vdd.n2245 gnd 0.007618f
C3055 vdd.n2246 gnd 0.007618f
C3056 vdd.n2247 gnd 0.007618f
C3057 vdd.n2248 gnd 0.007618f
C3058 vdd.n2249 gnd 0.007618f
C3059 vdd.n2250 gnd 0.007618f
C3060 vdd.n2251 gnd 0.007618f
C3061 vdd.n2252 gnd 0.007618f
C3062 vdd.n2253 gnd 0.007618f
C3063 vdd.n2254 gnd 0.007618f
C3064 vdd.n2255 gnd 0.007618f
C3065 vdd.n2256 gnd 0.007618f
C3066 vdd.n2257 gnd 0.246155f
C3067 vdd.n2258 gnd 0.007618f
C3068 vdd.n2259 gnd 0.007618f
C3069 vdd.n2260 gnd 0.007618f
C3070 vdd.n2261 gnd 0.007618f
C3071 vdd.n2262 gnd 0.007618f
C3072 vdd.n2263 gnd 0.007618f
C3073 vdd.n2264 gnd 0.007618f
C3074 vdd.n2265 gnd 0.007618f
C3075 vdd.n2266 gnd 0.007618f
C3076 vdd.n2267 gnd 0.007618f
C3077 vdd.n2268 gnd 0.007618f
C3078 vdd.n2269 gnd 0.007618f
C3079 vdd.n2270 gnd 0.007618f
C3080 vdd.n2271 gnd 0.007618f
C3081 vdd.n2272 gnd 0.007618f
C3082 vdd.n2273 gnd 0.007618f
C3083 vdd.n2274 gnd 0.007618f
C3084 vdd.n2275 gnd 0.007618f
C3085 vdd.n2276 gnd 0.007618f
C3086 vdd.n2277 gnd 0.007618f
C3087 vdd.n2278 gnd 0.016877f
C3088 vdd.n2280 gnd 0.018076f
C3089 vdd.n2281 gnd 0.018076f
C3090 vdd.n2282 gnd 0.007618f
C3091 vdd.n2283 gnd 0.005882f
C3092 vdd.n2284 gnd 0.007618f
C3093 vdd.n2286 gnd 0.007618f
C3094 vdd.n2288 gnd 0.007618f
C3095 vdd.n2289 gnd 0.007618f
C3096 vdd.n2290 gnd 0.007618f
C3097 vdd.n2291 gnd 0.007618f
C3098 vdd.n2292 gnd 0.007618f
C3099 vdd.n2294 gnd 0.007618f
C3100 vdd.n2296 gnd 0.007618f
C3101 vdd.n2297 gnd 0.007618f
C3102 vdd.n2298 gnd 0.007618f
C3103 vdd.n2299 gnd 0.007618f
C3104 vdd.n2300 gnd 0.007618f
C3105 vdd.n2302 gnd 0.007618f
C3106 vdd.n2304 gnd 0.007618f
C3107 vdd.n2305 gnd 0.007618f
C3108 vdd.n2306 gnd 0.007618f
C3109 vdd.n2307 gnd 0.007618f
C3110 vdd.n2308 gnd 0.007618f
C3111 vdd.n2310 gnd 0.007618f
C3112 vdd.n2312 gnd 0.007618f
C3113 vdd.n2313 gnd 0.007618f
C3114 vdd.n2314 gnd 0.022723f
C3115 vdd.n2315 gnd 0.673614f
C3116 vdd.n2317 gnd 0.009017f
C3117 vdd.n2318 gnd 0.009017f
C3118 vdd.n2319 gnd 0.011203f
C3119 vdd.n2321 gnd 0.011203f
C3120 vdd.n2322 gnd 0.011203f
C3121 vdd.n2323 gnd 0.009017f
C3122 vdd.n2324 gnd 0.007484f
C3123 vdd.n2325 gnd 0.027682f
C3124 vdd.n2326 gnd 0.027101f
C3125 vdd.n2327 gnd 0.007484f
C3126 vdd.n2328 gnd 0.027101f
C3127 vdd.n2329 gnd 1.57424f
C3128 vdd.n2330 gnd 0.027101f
C3129 vdd.n2331 gnd 0.027682f
C3130 vdd.n2332 gnd 0.004283f
C3131 vdd.t220 gnd 0.137828f
C3132 vdd.t219 gnd 0.1473f
C3133 vdd.t217 gnd 0.180001f
C3134 vdd.n2333 gnd 0.230736f
C3135 vdd.n2334 gnd 0.19386f
C3136 vdd.n2335 gnd 0.013886f
C3137 vdd.n2336 gnd 0.004734f
C3138 vdd.n2337 gnd 0.009635f
C3139 vdd.n2338 gnd 0.673614f
C3140 vdd.n2339 gnd 0.022723f
C3141 vdd.n2340 gnd 0.007618f
C3142 vdd.n2341 gnd 0.007618f
C3143 vdd.n2342 gnd 0.007618f
C3144 vdd.n2344 gnd 0.007618f
C3145 vdd.n2346 gnd 0.007618f
C3146 vdd.n2347 gnd 0.007618f
C3147 vdd.n2348 gnd 0.007618f
C3148 vdd.n2349 gnd 0.007618f
C3149 vdd.n2350 gnd 0.007618f
C3150 vdd.n2352 gnd 0.007618f
C3151 vdd.n2354 gnd 0.007618f
C3152 vdd.n2355 gnd 0.007618f
C3153 vdd.n2356 gnd 0.007618f
C3154 vdd.n2357 gnd 0.007618f
C3155 vdd.n2358 gnd 0.007618f
C3156 vdd.n2360 gnd 0.007618f
C3157 vdd.n2362 gnd 0.007618f
C3158 vdd.n2363 gnd 0.007618f
C3159 vdd.n2364 gnd 0.007618f
C3160 vdd.n2365 gnd 0.007618f
C3161 vdd.n2366 gnd 0.007618f
C3162 vdd.n2368 gnd 0.007618f
C3163 vdd.n2370 gnd 0.007618f
C3164 vdd.n2371 gnd 0.007618f
C3165 vdd.n2372 gnd 0.018076f
C3166 vdd.n2373 gnd 0.016877f
C3167 vdd.n2374 gnd 0.016877f
C3168 vdd.n2375 gnd 1.12201f
C3169 vdd.n2376 gnd 0.016877f
C3170 vdd.n2377 gnd 0.016877f
C3171 vdd.n2378 gnd 0.007618f
C3172 vdd.n2379 gnd 0.007618f
C3173 vdd.n2380 gnd 0.007618f
C3174 vdd.n2381 gnd 0.486585f
C3175 vdd.n2382 gnd 0.007618f
C3176 vdd.n2383 gnd 0.007618f
C3177 vdd.n2384 gnd 0.007618f
C3178 vdd.n2385 gnd 0.007618f
C3179 vdd.n2386 gnd 0.007618f
C3180 vdd.n2387 gnd 0.778536f
C3181 vdd.n2388 gnd 0.007618f
C3182 vdd.n2389 gnd 0.007618f
C3183 vdd.n2390 gnd 0.007618f
C3184 vdd.n2391 gnd 0.007618f
C3185 vdd.n2392 gnd 0.007618f
C3186 vdd.n2393 gnd 0.778536f
C3187 vdd.n2394 gnd 0.007618f
C3188 vdd.n2395 gnd 0.007618f
C3189 vdd.n2396 gnd 0.006722f
C3190 vdd.n2397 gnd 0.022069f
C3191 vdd.n2398 gnd 0.004705f
C3192 vdd.n2399 gnd 0.007618f
C3193 vdd.n2400 gnd 0.429339f
C3194 vdd.n2401 gnd 0.007618f
C3195 vdd.n2402 gnd 0.007618f
C3196 vdd.n2403 gnd 0.007618f
C3197 vdd.n2404 gnd 0.007618f
C3198 vdd.n2405 gnd 0.007618f
C3199 vdd.n2406 gnd 0.520932f
C3200 vdd.n2407 gnd 0.007618f
C3201 vdd.n2408 gnd 0.007618f
C3202 vdd.n2409 gnd 0.007618f
C3203 vdd.n2410 gnd 0.007618f
C3204 vdd.n2411 gnd 0.007618f
C3205 vdd.n2412 gnd 0.692668f
C3206 vdd.n2413 gnd 0.007618f
C3207 vdd.n2414 gnd 0.007618f
C3208 vdd.n2415 gnd 0.007618f
C3209 vdd.n2416 gnd 0.007618f
C3210 vdd.n2417 gnd 0.007618f
C3211 vdd.n2418 gnd 0.618249f
C3212 vdd.n2419 gnd 0.007618f
C3213 vdd.n2420 gnd 0.007618f
C3214 vdd.n2421 gnd 0.007618f
C3215 vdd.n2422 gnd 0.007618f
C3216 vdd.n2423 gnd 0.007618f
C3217 vdd.n2424 gnd 0.446513f
C3218 vdd.n2425 gnd 0.007618f
C3219 vdd.n2426 gnd 0.007618f
C3220 vdd.n2427 gnd 0.007618f
C3221 vdd.n2428 gnd 0.007618f
C3222 vdd.n2429 gnd 0.007618f
C3223 vdd.n2430 gnd 0.246155f
C3224 vdd.n2431 gnd 0.007618f
C3225 vdd.n2432 gnd 0.007618f
C3226 vdd.n2433 gnd 0.007618f
C3227 vdd.n2434 gnd 0.007618f
C3228 vdd.n2435 gnd 0.007618f
C3229 vdd.n2436 gnd 0.429339f
C3230 vdd.n2437 gnd 0.007618f
C3231 vdd.n2438 gnd 0.007618f
C3232 vdd.n2439 gnd 0.007618f
C3233 vdd.n2440 gnd 0.007618f
C3234 vdd.n2441 gnd 0.007618f
C3235 vdd.n2442 gnd 0.778536f
C3236 vdd.n2443 gnd 0.007618f
C3237 vdd.n2444 gnd 0.007618f
C3238 vdd.n2445 gnd 0.007618f
C3239 vdd.n2446 gnd 0.007618f
C3240 vdd.n2447 gnd 0.007618f
C3241 vdd.n2448 gnd 0.007618f
C3242 vdd.n2449 gnd 0.007618f
C3243 vdd.n2450 gnd 0.6068f
C3244 vdd.n2451 gnd 0.007618f
C3245 vdd.n2452 gnd 0.007618f
C3246 vdd.n2453 gnd 0.007618f
C3247 vdd.n2454 gnd 0.007618f
C3248 vdd.n2455 gnd 0.007618f
C3249 vdd.n2456 gnd 0.007618f
C3250 vdd.n2457 gnd 0.486585f
C3251 vdd.n2458 gnd 0.007618f
C3252 vdd.n2459 gnd 0.007618f
C3253 vdd.n2460 gnd 0.007618f
C3254 vdd.n2461 gnd 0.017805f
C3255 vdd.n2462 gnd 0.017149f
C3256 vdd.n2463 gnd 0.007618f
C3257 vdd.n2464 gnd 0.007618f
C3258 vdd.n2465 gnd 0.005882f
C3259 vdd.n2466 gnd 0.007618f
C3260 vdd.n2467 gnd 0.007618f
C3261 vdd.n2468 gnd 0.005546f
C3262 vdd.n2469 gnd 0.007618f
C3263 vdd.n2470 gnd 0.007618f
C3264 vdd.n2471 gnd 0.007618f
C3265 vdd.n2472 gnd 0.007618f
C3266 vdd.n2473 gnd 0.007618f
C3267 vdd.n2474 gnd 0.007618f
C3268 vdd.n2475 gnd 0.007618f
C3269 vdd.n2476 gnd 0.007618f
C3270 vdd.n2477 gnd 0.007618f
C3271 vdd.n2478 gnd 0.007618f
C3272 vdd.n2479 gnd 0.007618f
C3273 vdd.n2480 gnd 0.007618f
C3274 vdd.n2481 gnd 0.007618f
C3275 vdd.n2482 gnd 0.007618f
C3276 vdd.n2483 gnd 0.007618f
C3277 vdd.n2484 gnd 0.007618f
C3278 vdd.n2485 gnd 0.007618f
C3279 vdd.n2486 gnd 0.007618f
C3280 vdd.n2487 gnd 0.007618f
C3281 vdd.n2488 gnd 0.007618f
C3282 vdd.n2489 gnd 0.007618f
C3283 vdd.n2490 gnd 0.007618f
C3284 vdd.n2491 gnd 0.007618f
C3285 vdd.n2492 gnd 0.007618f
C3286 vdd.n2493 gnd 0.007618f
C3287 vdd.n2494 gnd 0.007618f
C3288 vdd.n2495 gnd 0.007618f
C3289 vdd.n2496 gnd 0.007618f
C3290 vdd.n2497 gnd 0.007618f
C3291 vdd.n2498 gnd 0.007618f
C3292 vdd.n2499 gnd 0.007618f
C3293 vdd.n2500 gnd 0.007618f
C3294 vdd.n2501 gnd 0.007618f
C3295 vdd.n2502 gnd 0.007618f
C3296 vdd.n2503 gnd 0.007618f
C3297 vdd.n2504 gnd 0.007618f
C3298 vdd.n2505 gnd 0.007618f
C3299 vdd.n2506 gnd 0.007618f
C3300 vdd.n2507 gnd 0.007618f
C3301 vdd.n2508 gnd 0.007618f
C3302 vdd.n2509 gnd 0.007618f
C3303 vdd.n2510 gnd 0.007618f
C3304 vdd.n2511 gnd 0.007618f
C3305 vdd.n2512 gnd 0.007618f
C3306 vdd.n2513 gnd 0.007618f
C3307 vdd.n2514 gnd 0.007618f
C3308 vdd.n2515 gnd 0.007618f
C3309 vdd.n2516 gnd 0.007618f
C3310 vdd.n2517 gnd 0.007618f
C3311 vdd.n2518 gnd 0.007618f
C3312 vdd.n2519 gnd 0.007618f
C3313 vdd.n2520 gnd 0.007618f
C3314 vdd.n2521 gnd 0.007618f
C3315 vdd.n2522 gnd 0.007618f
C3316 vdd.n2523 gnd 0.007618f
C3317 vdd.n2524 gnd 0.007618f
C3318 vdd.n2525 gnd 0.007618f
C3319 vdd.n2526 gnd 0.007618f
C3320 vdd.n2527 gnd 0.007618f
C3321 vdd.n2528 gnd 0.007618f
C3322 vdd.n2529 gnd 0.018076f
C3323 vdd.n2530 gnd 0.016877f
C3324 vdd.n2531 gnd 0.016877f
C3325 vdd.n2532 gnd 0.950271f
C3326 vdd.n2533 gnd 0.016877f
C3327 vdd.n2534 gnd 0.018076f
C3328 vdd.n2535 gnd 0.017149f
C3329 vdd.n2536 gnd 0.007618f
C3330 vdd.n2537 gnd 0.007618f
C3331 vdd.n2538 gnd 0.007618f
C3332 vdd.n2539 gnd 0.005882f
C3333 vdd.n2540 gnd 0.010887f
C3334 vdd.n2541 gnd 0.005546f
C3335 vdd.n2542 gnd 0.007618f
C3336 vdd.n2543 gnd 0.007618f
C3337 vdd.n2544 gnd 0.007618f
C3338 vdd.n2545 gnd 0.007618f
C3339 vdd.n2546 gnd 0.007618f
C3340 vdd.n2547 gnd 0.007618f
C3341 vdd.n2548 gnd 0.007618f
C3342 vdd.n2549 gnd 0.007618f
C3343 vdd.n2550 gnd 0.007618f
C3344 vdd.n2551 gnd 0.007618f
C3345 vdd.n2552 gnd 0.007618f
C3346 vdd.n2553 gnd 0.007618f
C3347 vdd.n2554 gnd 0.007618f
C3348 vdd.n2555 gnd 0.007618f
C3349 vdd.n2556 gnd 0.007618f
C3350 vdd.n2557 gnd 0.007618f
C3351 vdd.n2558 gnd 0.007618f
C3352 vdd.n2559 gnd 0.007618f
C3353 vdd.n2560 gnd 0.007618f
C3354 vdd.n2561 gnd 0.007618f
C3355 vdd.n2562 gnd 0.007618f
C3356 vdd.n2563 gnd 0.007618f
C3357 vdd.n2564 gnd 0.007618f
C3358 vdd.n2565 gnd 0.007618f
C3359 vdd.n2566 gnd 0.007618f
C3360 vdd.n2567 gnd 0.007618f
C3361 vdd.n2568 gnd 0.007618f
C3362 vdd.n2569 gnd 0.007618f
C3363 vdd.n2570 gnd 0.007618f
C3364 vdd.n2571 gnd 0.007618f
C3365 vdd.n2572 gnd 0.007618f
C3366 vdd.n2573 gnd 0.007618f
C3367 vdd.n2574 gnd 0.007618f
C3368 vdd.n2575 gnd 0.007618f
C3369 vdd.n2576 gnd 0.007618f
C3370 vdd.n2577 gnd 0.007618f
C3371 vdd.n2578 gnd 0.007618f
C3372 vdd.n2579 gnd 0.007618f
C3373 vdd.n2580 gnd 0.007618f
C3374 vdd.n2581 gnd 0.007618f
C3375 vdd.n2582 gnd 0.007618f
C3376 vdd.n2583 gnd 0.007618f
C3377 vdd.n2584 gnd 0.007618f
C3378 vdd.n2585 gnd 0.007618f
C3379 vdd.n2586 gnd 0.007618f
C3380 vdd.n2587 gnd 0.007618f
C3381 vdd.n2588 gnd 0.007618f
C3382 vdd.n2589 gnd 0.007618f
C3383 vdd.n2590 gnd 0.007618f
C3384 vdd.n2591 gnd 0.007618f
C3385 vdd.n2592 gnd 0.007618f
C3386 vdd.n2593 gnd 0.007618f
C3387 vdd.n2594 gnd 0.007618f
C3388 vdd.n2595 gnd 0.007618f
C3389 vdd.n2596 gnd 0.007618f
C3390 vdd.n2597 gnd 0.007618f
C3391 vdd.n2598 gnd 0.007618f
C3392 vdd.n2599 gnd 0.007618f
C3393 vdd.n2600 gnd 0.007618f
C3394 vdd.n2601 gnd 0.007618f
C3395 vdd.n2602 gnd 0.018076f
C3396 vdd.n2603 gnd 0.018076f
C3397 vdd.n2604 gnd 0.950271f
C3398 vdd.t181 gnd 3.37747f
C3399 vdd.t292 gnd 3.37747f
C3400 vdd.n2637 gnd 0.018076f
C3401 vdd.n2638 gnd 0.007618f
C3402 vdd.t255 gnd 0.307847f
C3403 vdd.t256 gnd 0.31512f
C3404 vdd.t253 gnd 0.200974f
C3405 vdd.n2639 gnd 0.108616f
C3406 vdd.n2640 gnd 0.06161f
C3407 vdd.n2641 gnd 0.007618f
C3408 vdd.t268 gnd 0.307847f
C3409 vdd.t269 gnd 0.31512f
C3410 vdd.t267 gnd 0.200974f
C3411 vdd.n2642 gnd 0.108616f
C3412 vdd.n2643 gnd 0.06161f
C3413 vdd.n2644 gnd 0.010887f
C3414 vdd.n2645 gnd 0.007618f
C3415 vdd.n2646 gnd 0.007618f
C3416 vdd.n2647 gnd 0.007618f
C3417 vdd.n2648 gnd 0.007618f
C3418 vdd.n2649 gnd 0.007618f
C3419 vdd.n2650 gnd 0.007618f
C3420 vdd.n2651 gnd 0.007618f
C3421 vdd.n2652 gnd 0.007618f
C3422 vdd.n2653 gnd 0.007618f
C3423 vdd.n2654 gnd 0.007618f
C3424 vdd.n2655 gnd 0.007618f
C3425 vdd.n2656 gnd 0.007618f
C3426 vdd.n2657 gnd 0.007618f
C3427 vdd.n2658 gnd 0.007618f
C3428 vdd.n2659 gnd 0.007618f
C3429 vdd.n2660 gnd 0.007618f
C3430 vdd.n2661 gnd 0.007618f
C3431 vdd.n2662 gnd 0.007618f
C3432 vdd.n2663 gnd 0.007618f
C3433 vdd.n2664 gnd 0.007618f
C3434 vdd.n2665 gnd 0.007618f
C3435 vdd.n2666 gnd 0.007618f
C3436 vdd.n2667 gnd 0.007618f
C3437 vdd.n2668 gnd 0.007618f
C3438 vdd.n2669 gnd 0.007618f
C3439 vdd.n2670 gnd 0.007618f
C3440 vdd.n2671 gnd 0.007618f
C3441 vdd.n2672 gnd 0.007618f
C3442 vdd.n2673 gnd 0.007618f
C3443 vdd.n2674 gnd 0.007618f
C3444 vdd.n2675 gnd 0.007618f
C3445 vdd.n2676 gnd 0.007618f
C3446 vdd.n2677 gnd 0.007618f
C3447 vdd.n2678 gnd 0.007618f
C3448 vdd.n2679 gnd 0.007618f
C3449 vdd.n2680 gnd 0.007618f
C3450 vdd.n2681 gnd 0.007618f
C3451 vdd.n2682 gnd 0.007618f
C3452 vdd.n2683 gnd 0.007618f
C3453 vdd.n2684 gnd 0.007618f
C3454 vdd.n2685 gnd 0.007618f
C3455 vdd.n2686 gnd 0.007618f
C3456 vdd.n2687 gnd 0.007618f
C3457 vdd.n2688 gnd 0.007618f
C3458 vdd.n2689 gnd 0.007618f
C3459 vdd.n2690 gnd 0.007618f
C3460 vdd.n2691 gnd 0.007618f
C3461 vdd.n2692 gnd 0.007618f
C3462 vdd.n2693 gnd 0.007618f
C3463 vdd.n2694 gnd 0.007618f
C3464 vdd.n2695 gnd 0.007618f
C3465 vdd.n2696 gnd 0.007618f
C3466 vdd.n2697 gnd 0.007618f
C3467 vdd.n2698 gnd 0.007618f
C3468 vdd.n2699 gnd 0.007618f
C3469 vdd.n2700 gnd 0.007618f
C3470 vdd.n2701 gnd 0.005546f
C3471 vdd.n2702 gnd 0.007618f
C3472 vdd.n2703 gnd 0.007618f
C3473 vdd.n2704 gnd 0.005882f
C3474 vdd.n2705 gnd 0.007618f
C3475 vdd.n2706 gnd 0.007618f
C3476 vdd.n2707 gnd 0.018076f
C3477 vdd.n2708 gnd 0.016877f
C3478 vdd.n2709 gnd 0.007618f
C3479 vdd.n2710 gnd 0.007618f
C3480 vdd.n2711 gnd 0.007618f
C3481 vdd.n2712 gnd 0.007618f
C3482 vdd.n2713 gnd 0.007618f
C3483 vdd.n2714 gnd 0.007618f
C3484 vdd.n2715 gnd 0.007618f
C3485 vdd.n2716 gnd 0.007618f
C3486 vdd.n2717 gnd 0.007618f
C3487 vdd.n2718 gnd 0.007618f
C3488 vdd.n2719 gnd 0.007618f
C3489 vdd.n2720 gnd 0.007618f
C3490 vdd.n2721 gnd 0.007618f
C3491 vdd.n2722 gnd 0.007618f
C3492 vdd.n2723 gnd 0.007618f
C3493 vdd.n2724 gnd 0.007618f
C3494 vdd.n2725 gnd 0.007618f
C3495 vdd.n2726 gnd 0.007618f
C3496 vdd.n2727 gnd 0.007618f
C3497 vdd.n2728 gnd 0.007618f
C3498 vdd.n2729 gnd 0.007618f
C3499 vdd.n2730 gnd 0.007618f
C3500 vdd.n2731 gnd 0.007618f
C3501 vdd.n2732 gnd 0.007618f
C3502 vdd.n2733 gnd 0.007618f
C3503 vdd.n2734 gnd 0.007618f
C3504 vdd.n2735 gnd 0.007618f
C3505 vdd.n2736 gnd 0.007618f
C3506 vdd.n2737 gnd 0.007618f
C3507 vdd.n2738 gnd 0.007618f
C3508 vdd.n2739 gnd 0.007618f
C3509 vdd.n2740 gnd 0.007618f
C3510 vdd.n2741 gnd 0.007618f
C3511 vdd.n2742 gnd 0.007618f
C3512 vdd.n2743 gnd 0.007618f
C3513 vdd.n2744 gnd 0.007618f
C3514 vdd.n2745 gnd 0.007618f
C3515 vdd.n2746 gnd 0.007618f
C3516 vdd.n2747 gnd 0.007618f
C3517 vdd.n2748 gnd 0.007618f
C3518 vdd.n2749 gnd 0.007618f
C3519 vdd.n2750 gnd 0.007618f
C3520 vdd.n2751 gnd 0.007618f
C3521 vdd.n2752 gnd 0.007618f
C3522 vdd.n2753 gnd 0.007618f
C3523 vdd.n2754 gnd 0.007618f
C3524 vdd.n2755 gnd 0.007618f
C3525 vdd.n2756 gnd 0.007618f
C3526 vdd.n2757 gnd 0.007618f
C3527 vdd.n2758 gnd 0.007618f
C3528 vdd.n2759 gnd 0.007618f
C3529 vdd.n2760 gnd 0.246155f
C3530 vdd.n2761 gnd 0.007618f
C3531 vdd.n2762 gnd 0.007618f
C3532 vdd.n2763 gnd 0.007618f
C3533 vdd.n2764 gnd 0.007618f
C3534 vdd.n2765 gnd 0.007618f
C3535 vdd.n2766 gnd 0.007618f
C3536 vdd.n2767 gnd 0.007618f
C3537 vdd.n2768 gnd 0.007618f
C3538 vdd.n2769 gnd 0.007618f
C3539 vdd.n2770 gnd 0.007618f
C3540 vdd.n2771 gnd 0.007618f
C3541 vdd.n2772 gnd 0.007618f
C3542 vdd.n2773 gnd 0.007618f
C3543 vdd.n2774 gnd 0.007618f
C3544 vdd.n2775 gnd 0.007618f
C3545 vdd.n2776 gnd 0.007618f
C3546 vdd.n2777 gnd 0.007618f
C3547 vdd.n2778 gnd 0.007618f
C3548 vdd.n2779 gnd 0.007618f
C3549 vdd.n2780 gnd 0.007618f
C3550 vdd.n2781 gnd 0.463687f
C3551 vdd.n2782 gnd 0.007618f
C3552 vdd.n2783 gnd 0.007618f
C3553 vdd.n2784 gnd 0.007618f
C3554 vdd.n2785 gnd 0.007618f
C3555 vdd.n2786 gnd 0.007618f
C3556 vdd.n2787 gnd 0.016877f
C3557 vdd.n2788 gnd 0.018076f
C3558 vdd.n2789 gnd 0.018076f
C3559 vdd.n2790 gnd 0.007618f
C3560 vdd.n2791 gnd 0.007618f
C3561 vdd.n2792 gnd 0.007618f
C3562 vdd.n2793 gnd 0.005882f
C3563 vdd.n2794 gnd 0.010887f
C3564 vdd.n2795 gnd 0.005546f
C3565 vdd.n2796 gnd 0.007618f
C3566 vdd.n2797 gnd 0.007618f
C3567 vdd.n2798 gnd 0.007618f
C3568 vdd.n2799 gnd 0.007618f
C3569 vdd.n2800 gnd 0.007618f
C3570 vdd.n2801 gnd 0.007618f
C3571 vdd.n2802 gnd 0.007618f
C3572 vdd.n2803 gnd 0.007618f
C3573 vdd.n2804 gnd 0.007618f
C3574 vdd.n2805 gnd 0.007618f
C3575 vdd.n2806 gnd 0.007618f
C3576 vdd.n2807 gnd 0.007618f
C3577 vdd.n2808 gnd 0.007618f
C3578 vdd.n2809 gnd 0.007618f
C3579 vdd.n2810 gnd 0.007618f
C3580 vdd.n2811 gnd 0.007618f
C3581 vdd.n2812 gnd 0.007618f
C3582 vdd.n2813 gnd 0.007618f
C3583 vdd.n2814 gnd 0.007618f
C3584 vdd.n2815 gnd 0.007618f
C3585 vdd.n2816 gnd 0.007618f
C3586 vdd.n2817 gnd 0.007618f
C3587 vdd.n2818 gnd 0.007618f
C3588 vdd.n2819 gnd 0.007618f
C3589 vdd.n2820 gnd 0.007618f
C3590 vdd.n2821 gnd 0.007618f
C3591 vdd.n2822 gnd 0.007618f
C3592 vdd.n2823 gnd 0.007618f
C3593 vdd.n2824 gnd 0.007618f
C3594 vdd.n2825 gnd 0.007618f
C3595 vdd.n2826 gnd 0.007618f
C3596 vdd.n2827 gnd 0.007618f
C3597 vdd.n2828 gnd 0.007618f
C3598 vdd.n2829 gnd 0.007618f
C3599 vdd.n2830 gnd 0.007618f
C3600 vdd.n2831 gnd 0.007618f
C3601 vdd.n2832 gnd 0.007618f
C3602 vdd.n2833 gnd 0.007618f
C3603 vdd.n2834 gnd 0.007618f
C3604 vdd.n2835 gnd 0.007618f
C3605 vdd.n2836 gnd 0.007618f
C3606 vdd.n2837 gnd 0.007618f
C3607 vdd.n2838 gnd 0.007618f
C3608 vdd.n2839 gnd 0.007618f
C3609 vdd.n2840 gnd 0.007618f
C3610 vdd.n2841 gnd 0.007618f
C3611 vdd.n2842 gnd 0.007618f
C3612 vdd.n2843 gnd 0.007618f
C3613 vdd.n2844 gnd 0.007618f
C3614 vdd.n2845 gnd 0.007618f
C3615 vdd.n2846 gnd 0.007618f
C3616 vdd.n2847 gnd 0.007618f
C3617 vdd.n2848 gnd 0.007618f
C3618 vdd.n2849 gnd 0.007618f
C3619 vdd.n2850 gnd 0.007618f
C3620 vdd.n2851 gnd 0.007618f
C3621 vdd.n2852 gnd 0.007618f
C3622 vdd.n2853 gnd 0.007618f
C3623 vdd.n2854 gnd 0.007618f
C3624 vdd.n2855 gnd 0.007618f
C3625 vdd.n2857 gnd 0.950271f
C3626 vdd.n2859 gnd 0.007618f
C3627 vdd.n2860 gnd 0.007618f
C3628 vdd.n2861 gnd 0.018076f
C3629 vdd.n2862 gnd 0.016877f
C3630 vdd.n2863 gnd 0.016877f
C3631 vdd.n2864 gnd 0.950271f
C3632 vdd.n2865 gnd 0.016877f
C3633 vdd.n2866 gnd 0.016877f
C3634 vdd.n2867 gnd 0.007618f
C3635 vdd.n2868 gnd 0.007618f
C3636 vdd.n2869 gnd 0.007618f
C3637 vdd.n2870 gnd 0.486585f
C3638 vdd.n2871 gnd 0.007618f
C3639 vdd.n2872 gnd 0.007618f
C3640 vdd.n2873 gnd 0.007618f
C3641 vdd.n2874 gnd 0.007618f
C3642 vdd.n2875 gnd 0.007618f
C3643 vdd.n2876 gnd 0.6068f
C3644 vdd.n2877 gnd 0.007618f
C3645 vdd.n2878 gnd 0.007618f
C3646 vdd.n2879 gnd 0.007618f
C3647 vdd.n2880 gnd 0.007618f
C3648 vdd.n2881 gnd 0.007618f
C3649 vdd.n2882 gnd 0.778536f
C3650 vdd.n2883 gnd 0.007618f
C3651 vdd.n2884 gnd 0.007618f
C3652 vdd.n2885 gnd 0.007618f
C3653 vdd.n2886 gnd 0.007618f
C3654 vdd.n2887 gnd 0.007618f
C3655 vdd.n2888 gnd 0.429339f
C3656 vdd.n2889 gnd 0.007618f
C3657 vdd.n2890 gnd 0.007618f
C3658 vdd.n2891 gnd 0.007618f
C3659 vdd.n2892 gnd 0.007618f
C3660 vdd.n2893 gnd 0.007618f
C3661 vdd.n2894 gnd 0.246155f
C3662 vdd.n2895 gnd 0.007618f
C3663 vdd.n2896 gnd 0.007618f
C3664 vdd.n2897 gnd 0.007618f
C3665 vdd.n2898 gnd 0.007618f
C3666 vdd.n2899 gnd 0.007618f
C3667 vdd.n2900 gnd 0.446513f
C3668 vdd.n2901 gnd 0.007618f
C3669 vdd.n2902 gnd 0.007618f
C3670 vdd.n2903 gnd 0.007618f
C3671 vdd.n2904 gnd 0.007618f
C3672 vdd.n2905 gnd 0.007618f
C3673 vdd.n2906 gnd 0.618249f
C3674 vdd.n2907 gnd 0.007618f
C3675 vdd.n2908 gnd 0.007618f
C3676 vdd.n2909 gnd 0.007618f
C3677 vdd.n2910 gnd 0.007618f
C3678 vdd.n2911 gnd 0.007618f
C3679 vdd.n2912 gnd 0.692668f
C3680 vdd.n2913 gnd 0.007618f
C3681 vdd.n2914 gnd 0.007618f
C3682 vdd.n2915 gnd 0.007618f
C3683 vdd.n2916 gnd 0.007618f
C3684 vdd.n2917 gnd 0.007618f
C3685 vdd.n2918 gnd 0.520932f
C3686 vdd.n2919 gnd 0.007618f
C3687 vdd.n2920 gnd 0.007618f
C3688 vdd.n2921 gnd 0.007618f
C3689 vdd.t223 gnd 0.31512f
C3690 vdd.t221 gnd 0.200974f
C3691 vdd.t224 gnd 0.31512f
C3692 vdd.n2922 gnd 0.17711f
C3693 vdd.n2923 gnd 0.022069f
C3694 vdd.n2924 gnd 0.004705f
C3695 vdd.n2925 gnd 0.007618f
C3696 vdd.n2926 gnd 0.429339f
C3697 vdd.n2927 gnd 0.007618f
C3698 vdd.n2928 gnd 0.007618f
C3699 vdd.n2929 gnd 0.007618f
C3700 vdd.n2930 gnd 0.007618f
C3701 vdd.n2931 gnd 0.007618f
C3702 vdd.n2932 gnd 0.778536f
C3703 vdd.n2933 gnd 0.007618f
C3704 vdd.n2934 gnd 0.007618f
C3705 vdd.n2935 gnd 0.007618f
C3706 vdd.n2936 gnd 0.007618f
C3707 vdd.n2937 gnd 0.007618f
C3708 vdd.n2938 gnd 0.007618f
C3709 vdd.n2940 gnd 0.007618f
C3710 vdd.n2941 gnd 0.007618f
C3711 vdd.n2943 gnd 0.007618f
C3712 vdd.n2944 gnd 0.007618f
C3713 vdd.n2947 gnd 0.007618f
C3714 vdd.n2948 gnd 0.007618f
C3715 vdd.n2949 gnd 0.007618f
C3716 vdd.n2950 gnd 0.007618f
C3717 vdd.n2952 gnd 0.007618f
C3718 vdd.n2953 gnd 0.007618f
C3719 vdd.n2954 gnd 0.007618f
C3720 vdd.n2955 gnd 0.007618f
C3721 vdd.n2956 gnd 0.007618f
C3722 vdd.n2957 gnd 0.007618f
C3723 vdd.n2959 gnd 0.007618f
C3724 vdd.n2960 gnd 0.007618f
C3725 vdd.n2961 gnd 0.007618f
C3726 vdd.n2962 gnd 0.007618f
C3727 vdd.n2963 gnd 0.007618f
C3728 vdd.n2964 gnd 0.007618f
C3729 vdd.n2966 gnd 0.007618f
C3730 vdd.n2967 gnd 0.007618f
C3731 vdd.n2968 gnd 0.007618f
C3732 vdd.n2969 gnd 0.007618f
C3733 vdd.n2970 gnd 0.007618f
C3734 vdd.n2971 gnd 0.007618f
C3735 vdd.n2973 gnd 0.007618f
C3736 vdd.n2974 gnd 0.018076f
C3737 vdd.n2975 gnd 0.018076f
C3738 vdd.n2976 gnd 0.016877f
C3739 vdd.n2977 gnd 0.007618f
C3740 vdd.n2978 gnd 0.007618f
C3741 vdd.n2979 gnd 0.007618f
C3742 vdd.n2980 gnd 0.007618f
C3743 vdd.n2981 gnd 0.007618f
C3744 vdd.n2982 gnd 0.007618f
C3745 vdd.n2983 gnd 0.778536f
C3746 vdd.n2984 gnd 0.007618f
C3747 vdd.n2985 gnd 0.007618f
C3748 vdd.n2986 gnd 0.007618f
C3749 vdd.n2987 gnd 0.007618f
C3750 vdd.n2988 gnd 0.007618f
C3751 vdd.n2989 gnd 0.486585f
C3752 vdd.n2990 gnd 0.007618f
C3753 vdd.n2991 gnd 0.007618f
C3754 vdd.n2992 gnd 0.007618f
C3755 vdd.n2993 gnd 0.017805f
C3756 vdd.n2994 gnd 0.017149f
C3757 vdd.n2995 gnd 0.018076f
C3758 vdd.n2997 gnd 0.007618f
C3759 vdd.n2998 gnd 0.007618f
C3760 vdd.n2999 gnd 0.005882f
C3761 vdd.n3000 gnd 0.010887f
C3762 vdd.n3001 gnd 0.005546f
C3763 vdd.n3002 gnd 0.007618f
C3764 vdd.n3003 gnd 0.007618f
C3765 vdd.n3005 gnd 0.007618f
C3766 vdd.n3006 gnd 0.007618f
C3767 vdd.n3007 gnd 0.007618f
C3768 vdd.n3008 gnd 0.007618f
C3769 vdd.n3009 gnd 0.007618f
C3770 vdd.n3010 gnd 0.007618f
C3771 vdd.n3012 gnd 0.007618f
C3772 vdd.n3013 gnd 0.007618f
C3773 vdd.n3014 gnd 0.007618f
C3774 vdd.n3015 gnd 0.007618f
C3775 vdd.n3016 gnd 0.007618f
C3776 vdd.n3017 gnd 0.007618f
C3777 vdd.n3019 gnd 0.007618f
C3778 vdd.n3020 gnd 0.007618f
C3779 vdd.n3021 gnd 0.007618f
C3780 vdd.n3022 gnd 0.007618f
C3781 vdd.n3023 gnd 0.007618f
C3782 vdd.n3024 gnd 0.007618f
C3783 vdd.n3026 gnd 0.007618f
C3784 vdd.n3027 gnd 0.007618f
C3785 vdd.n3028 gnd 0.007618f
C3786 vdd.n3030 gnd 0.007618f
C3787 vdd.n3031 gnd 0.007618f
C3788 vdd.n3032 gnd 0.007618f
C3789 vdd.n3033 gnd 0.007618f
C3790 vdd.n3034 gnd 0.007618f
C3791 vdd.n3035 gnd 0.007618f
C3792 vdd.n3037 gnd 0.007618f
C3793 vdd.n3038 gnd 0.007618f
C3794 vdd.n3039 gnd 0.007618f
C3795 vdd.n3040 gnd 0.007618f
C3796 vdd.n3041 gnd 0.007618f
C3797 vdd.n3042 gnd 0.007618f
C3798 vdd.n3044 gnd 0.007618f
C3799 vdd.n3045 gnd 0.007618f
C3800 vdd.n3046 gnd 0.007618f
C3801 vdd.n3047 gnd 0.007618f
C3802 vdd.n3048 gnd 0.007618f
C3803 vdd.n3049 gnd 0.007618f
C3804 vdd.n3051 gnd 0.007618f
C3805 vdd.n3052 gnd 0.007618f
C3806 vdd.n3054 gnd 0.007618f
C3807 vdd.n3055 gnd 0.007618f
C3808 vdd.n3056 gnd 0.018076f
C3809 vdd.n3057 gnd 0.016877f
C3810 vdd.n3058 gnd 0.016877f
C3811 vdd.n3059 gnd 1.12201f
C3812 vdd.n3060 gnd 0.016877f
C3813 vdd.n3061 gnd 0.018076f
C3814 vdd.n3062 gnd 0.017149f
C3815 vdd.n3063 gnd 0.007618f
C3816 vdd.n3064 gnd 0.005882f
C3817 vdd.n3065 gnd 0.007618f
C3818 vdd.n3067 gnd 0.007618f
C3819 vdd.n3068 gnd 0.007618f
C3820 vdd.n3069 gnd 0.007618f
C3821 vdd.n3070 gnd 0.007618f
C3822 vdd.n3071 gnd 0.007618f
C3823 vdd.n3072 gnd 0.007618f
C3824 vdd.n3074 gnd 0.007618f
C3825 vdd.n3075 gnd 0.007618f
C3826 vdd.n3076 gnd 0.007618f
C3827 vdd.n3077 gnd 0.007618f
C3828 vdd.n3078 gnd 0.007618f
C3829 vdd.n3079 gnd 0.007618f
C3830 vdd.n3081 gnd 0.007618f
C3831 vdd.n3082 gnd 0.007618f
C3832 vdd.n3083 gnd 0.007618f
C3833 vdd.n3084 gnd 0.007618f
C3834 vdd.n3085 gnd 0.007618f
C3835 vdd.n3086 gnd 0.007618f
C3836 vdd.n3088 gnd 0.007618f
C3837 vdd.n3089 gnd 0.007618f
C3838 vdd.n3091 gnd 0.007618f
C3839 vdd.n3092 gnd 0.018307f
C3840 vdd.n3093 gnd 0.678031f
C3841 vdd.n3095 gnd 0.004734f
C3842 vdd.n3096 gnd 0.009017f
C3843 vdd.n3097 gnd 0.011203f
C3844 vdd.n3098 gnd 0.011203f
C3845 vdd.n3099 gnd 0.009017f
C3846 vdd.n3100 gnd 0.009017f
C3847 vdd.n3101 gnd 0.011203f
C3848 vdd.n3102 gnd 0.011203f
C3849 vdd.n3103 gnd 0.009017f
C3850 vdd.n3104 gnd 0.009017f
C3851 vdd.n3105 gnd 0.011203f
C3852 vdd.n3106 gnd 0.011203f
C3853 vdd.n3107 gnd 0.009017f
C3854 vdd.n3108 gnd 0.009017f
C3855 vdd.n3109 gnd 0.011203f
C3856 vdd.n3110 gnd 0.011203f
C3857 vdd.n3111 gnd 0.009017f
C3858 vdd.n3112 gnd 0.009017f
C3859 vdd.n3113 gnd 0.011203f
C3860 vdd.n3114 gnd 0.011203f
C3861 vdd.n3115 gnd 0.009017f
C3862 vdd.n3116 gnd 0.009017f
C3863 vdd.n3117 gnd 0.011203f
C3864 vdd.n3118 gnd 0.011203f
C3865 vdd.n3119 gnd 0.009017f
C3866 vdd.n3120 gnd 0.009017f
C3867 vdd.n3121 gnd 0.011203f
C3868 vdd.n3122 gnd 0.011203f
C3869 vdd.n3123 gnd 0.009017f
C3870 vdd.n3124 gnd 0.009017f
C3871 vdd.n3125 gnd 0.011203f
C3872 vdd.n3126 gnd 0.011203f
C3873 vdd.n3127 gnd 0.009017f
C3874 vdd.n3128 gnd 0.009017f
C3875 vdd.n3129 gnd 0.011203f
C3876 vdd.n3130 gnd 0.011203f
C3877 vdd.n3131 gnd 0.009017f
C3878 vdd.n3132 gnd 0.011203f
C3879 vdd.n3133 gnd 0.011203f
C3880 vdd.n3134 gnd 0.009017f
C3881 vdd.n3135 gnd 0.011203f
C3882 vdd.n3136 gnd 0.011203f
C3883 vdd.n3137 gnd 0.011203f
C3884 vdd.n3138 gnd 0.018395f
C3885 vdd.n3139 gnd 0.011203f
C3886 vdd.n3140 gnd 0.011203f
C3887 vdd.n3141 gnd 0.006132f
C3888 vdd.n3142 gnd 0.009017f
C3889 vdd.n3143 gnd 0.011203f
C3890 vdd.n3144 gnd 0.011203f
C3891 vdd.n3145 gnd 0.009017f
C3892 vdd.n3146 gnd 0.009017f
C3893 vdd.n3147 gnd 0.011203f
C3894 vdd.n3148 gnd 0.011203f
C3895 vdd.n3149 gnd 0.009017f
C3896 vdd.n3150 gnd 0.009017f
C3897 vdd.n3151 gnd 0.011203f
C3898 vdd.n3152 gnd 0.011203f
C3899 vdd.n3153 gnd 0.009017f
C3900 vdd.n3154 gnd 0.009017f
C3901 vdd.n3155 gnd 0.011203f
C3902 vdd.n3156 gnd 0.011203f
C3903 vdd.n3157 gnd 0.009017f
C3904 vdd.n3158 gnd 0.009017f
C3905 vdd.n3159 gnd 0.011203f
C3906 vdd.n3160 gnd 0.011203f
C3907 vdd.n3161 gnd 0.009017f
C3908 vdd.n3162 gnd 0.009017f
C3909 vdd.n3163 gnd 0.011203f
C3910 vdd.n3164 gnd 0.011203f
C3911 vdd.n3165 gnd 0.009017f
C3912 vdd.n3166 gnd 0.009017f
C3913 vdd.n3167 gnd 0.011203f
C3914 vdd.n3168 gnd 0.011203f
C3915 vdd.n3169 gnd 0.009017f
C3916 vdd.n3170 gnd 0.009017f
C3917 vdd.n3171 gnd 0.011203f
C3918 vdd.n3172 gnd 0.011203f
C3919 vdd.n3173 gnd 0.009017f
C3920 vdd.n3174 gnd 0.009017f
C3921 vdd.n3175 gnd 0.011203f
C3922 vdd.n3176 gnd 0.011203f
C3923 vdd.n3177 gnd 0.009017f
C3924 vdd.n3178 gnd 0.011203f
C3925 vdd.n3179 gnd 0.011203f
C3926 vdd.n3180 gnd 0.009017f
C3927 vdd.n3181 gnd 0.011203f
C3928 vdd.n3182 gnd 0.011203f
C3929 vdd.n3183 gnd 0.011203f
C3930 vdd.t215 gnd 0.137828f
C3931 vdd.t216 gnd 0.1473f
C3932 vdd.t214 gnd 0.180001f
C3933 vdd.n3184 gnd 0.230736f
C3934 vdd.n3185 gnd 0.19386f
C3935 vdd.n3186 gnd 0.018395f
C3936 vdd.n3187 gnd 0.011203f
C3937 vdd.n3188 gnd 0.011203f
C3938 vdd.n3189 gnd 0.007529f
C3939 vdd.n3190 gnd 0.009017f
C3940 vdd.n3191 gnd 0.011203f
C3941 vdd.n3192 gnd 0.011203f
C3942 vdd.n3193 gnd 0.009017f
C3943 vdd.n3194 gnd 0.009017f
C3944 vdd.n3195 gnd 0.011203f
C3945 vdd.n3196 gnd 0.011203f
C3946 vdd.n3197 gnd 0.009017f
C3947 vdd.n3198 gnd 0.009017f
C3948 vdd.n3199 gnd 0.011203f
C3949 vdd.n3200 gnd 0.011203f
C3950 vdd.n3201 gnd 0.009017f
C3951 vdd.n3202 gnd 0.009017f
C3952 vdd.n3203 gnd 0.011203f
C3953 vdd.n3204 gnd 0.011203f
C3954 vdd.n3205 gnd 0.009017f
C3955 vdd.n3206 gnd 0.009017f
C3956 vdd.n3207 gnd 0.011203f
C3957 vdd.n3208 gnd 0.011203f
C3958 vdd.n3209 gnd 0.009017f
C3959 vdd.n3210 gnd 0.009017f
C3960 vdd.n3211 gnd 0.011203f
C3961 vdd.n3212 gnd 0.011203f
C3962 vdd.n3213 gnd 0.009017f
C3963 vdd.n3214 gnd 0.009017f
C3964 vdd.n3216 gnd 0.678031f
C3965 vdd.n3218 gnd 0.009017f
C3966 vdd.n3219 gnd 0.009017f
C3967 vdd.n3220 gnd 0.007484f
C3968 vdd.n3221 gnd 0.027682f
C3969 vdd.n3223 gnd 8.27767f
C3970 vdd.n3224 gnd 0.027682f
C3971 vdd.n3225 gnd 0.004283f
C3972 vdd.n3226 gnd 0.027682f
C3973 vdd.n3227 gnd 0.027101f
C3974 vdd.n3228 gnd 0.011203f
C3975 vdd.n3229 gnd 0.009017f
C3976 vdd.n3230 gnd 0.011203f
C3977 vdd.n3231 gnd 0.692668f
C3978 vdd.n3232 gnd 0.011203f
C3979 vdd.n3233 gnd 0.009017f
C3980 vdd.n3234 gnd 0.011203f
C3981 vdd.n3235 gnd 0.011203f
C3982 vdd.n3236 gnd 0.011203f
C3983 vdd.n3237 gnd 0.009017f
C3984 vdd.n3238 gnd 0.011203f
C3985 vdd.n3239 gnd 1.14491f
C3986 vdd.n3240 gnd 0.011203f
C3987 vdd.n3241 gnd 0.009017f
C3988 vdd.n3242 gnd 0.011203f
C3989 vdd.n3243 gnd 0.011203f
C3990 vdd.n3244 gnd 0.011203f
C3991 vdd.n3245 gnd 0.009017f
C3992 vdd.n3246 gnd 0.011203f
C3993 vdd.n3247 gnd 0.738464f
C3994 vdd.n3248 gnd 0.78426f
C3995 vdd.n3249 gnd 0.011203f
C3996 vdd.n3250 gnd 0.009017f
C3997 vdd.n3251 gnd 0.011203f
C3998 vdd.n3252 gnd 0.011203f
C3999 vdd.n3253 gnd 0.011203f
C4000 vdd.n3254 gnd 0.009017f
C4001 vdd.n3255 gnd 0.011203f
C4002 vdd.n3256 gnd 0.950271f
C4003 vdd.n3257 gnd 0.011203f
C4004 vdd.n3258 gnd 0.009017f
C4005 vdd.n3259 gnd 0.011203f
C4006 vdd.n3260 gnd 0.011203f
C4007 vdd.n3261 gnd 0.011203f
C4008 vdd.n3262 gnd 0.009017f
C4009 vdd.n3263 gnd 0.011203f
C4010 vdd.t23 gnd 0.572453f
C4011 vdd.n3264 gnd 0.921649f
C4012 vdd.n3265 gnd 0.011203f
C4013 vdd.n3266 gnd 0.009017f
C4014 vdd.n3267 gnd 0.011203f
C4015 vdd.n3268 gnd 0.011203f
C4016 vdd.n3269 gnd 0.011203f
C4017 vdd.n3270 gnd 0.009017f
C4018 vdd.n3271 gnd 0.011203f
C4019 vdd.n3272 gnd 0.727015f
C4020 vdd.n3273 gnd 0.011203f
C4021 vdd.n3274 gnd 0.009017f
C4022 vdd.n3275 gnd 0.011203f
C4023 vdd.n3276 gnd 0.011203f
C4024 vdd.n3277 gnd 0.011203f
C4025 vdd.n3278 gnd 0.009017f
C4026 vdd.n3279 gnd 0.011203f
C4027 vdd.n3280 gnd 0.9102f
C4028 vdd.n3281 gnd 0.612524f
C4029 vdd.n3282 gnd 0.011203f
C4030 vdd.n3283 gnd 0.009017f
C4031 vdd.n3284 gnd 0.011203f
C4032 vdd.n3285 gnd 0.011203f
C4033 vdd.n3286 gnd 0.011203f
C4034 vdd.n3287 gnd 0.009017f
C4035 vdd.n3288 gnd 0.011203f
C4036 vdd.n3289 gnd 0.807158f
C4037 vdd.n3290 gnd 0.011203f
C4038 vdd.n3291 gnd 0.009017f
C4039 vdd.n3292 gnd 0.011203f
C4040 vdd.n3293 gnd 0.011203f
C4041 vdd.n3294 gnd 0.011203f
C4042 vdd.n3295 gnd 0.011203f
C4043 vdd.n3296 gnd 0.011203f
C4044 vdd.n3297 gnd 0.009017f
C4045 vdd.n3298 gnd 0.009017f
C4046 vdd.n3299 gnd 0.011203f
C4047 vdd.t72 gnd 0.572453f
C4048 vdd.n3300 gnd 0.950271f
C4049 vdd.n3301 gnd 0.011203f
C4050 vdd.n3302 gnd 0.009017f
C4051 vdd.n3303 gnd 0.011203f
C4052 vdd.n3304 gnd 0.011203f
C4053 vdd.n3305 gnd 0.011203f
C4054 vdd.n3306 gnd 0.009017f
C4055 vdd.n3307 gnd 0.011203f
C4056 vdd.n3308 gnd 0.898751f
C4057 vdd.n3309 gnd 0.011203f
C4058 vdd.n3310 gnd 0.011203f
C4059 vdd.n3311 gnd 0.009017f
C4060 vdd.n3312 gnd 0.009017f
C4061 vdd.n3313 gnd 0.011203f
C4062 vdd.n3314 gnd 0.011203f
C4063 vdd.n3315 gnd 0.011203f
C4064 vdd.n3316 gnd 0.009017f
C4065 vdd.n3317 gnd 0.011203f
C4066 vdd.n3318 gnd 0.009017f
C4067 vdd.n3319 gnd 0.009017f
C4068 vdd.n3320 gnd 0.011203f
C4069 vdd.n3321 gnd 0.011203f
C4070 vdd.n3322 gnd 0.011203f
C4071 vdd.n3323 gnd 0.009017f
C4072 vdd.n3324 gnd 0.011203f
C4073 vdd.n3325 gnd 0.009017f
C4074 vdd.n3326 gnd 0.009017f
C4075 vdd.n3327 gnd 0.011203f
C4076 vdd.n3328 gnd 0.011203f
C4077 vdd.n3329 gnd 0.011203f
C4078 vdd.n3330 gnd 0.009017f
C4079 vdd.n3331 gnd 0.950271f
C4080 vdd.n3332 gnd 0.011203f
C4081 vdd.n3333 gnd 0.009017f
C4082 vdd.n3334 gnd 0.009017f
C4083 vdd.n3335 gnd 0.011203f
C4084 vdd.n3336 gnd 0.011203f
C4085 vdd.n3337 gnd 0.011203f
C4086 vdd.n3338 gnd 0.009017f
C4087 vdd.n3339 gnd 0.011203f
C4088 vdd.n3340 gnd 0.009017f
C4089 vdd.n3341 gnd 0.009017f
C4090 vdd.n3342 gnd 0.011203f
C4091 vdd.n3343 gnd 0.011203f
C4092 vdd.n3344 gnd 0.011203f
C4093 vdd.n3345 gnd 0.009017f
C4094 vdd.n3346 gnd 0.011203f
C4095 vdd.n3347 gnd 0.009017f
C4096 vdd.n3348 gnd 0.007484f
C4097 vdd.n3349 gnd 0.027101f
C4098 vdd.n3350 gnd 0.027682f
C4099 vdd.n3351 gnd 0.004283f
C4100 vdd.n3352 gnd 0.027682f
C4101 vdd.n3354 gnd 2.71343f
C4102 vdd.n3355 gnd 1.68874f
C4103 vdd.n3356 gnd 0.027101f
C4104 vdd.n3357 gnd 0.007484f
C4105 vdd.n3358 gnd 0.009017f
C4106 vdd.n3359 gnd 0.009017f
C4107 vdd.n3360 gnd 0.011203f
C4108 vdd.n3361 gnd 1.14491f
C4109 vdd.n3362 gnd 1.14491f
C4110 vdd.n3363 gnd 1.04759f
C4111 vdd.n3364 gnd 0.011203f
C4112 vdd.n3365 gnd 0.009017f
C4113 vdd.n3366 gnd 0.009017f
C4114 vdd.n3367 gnd 0.009017f
C4115 vdd.n3368 gnd 0.011203f
C4116 vdd.n3369 gnd 0.852954f
C4117 vdd.t91 gnd 0.572453f
C4118 vdd.n3370 gnd 0.864404f
C4119 vdd.n3371 gnd 0.658321f
C4120 vdd.n3372 gnd 0.011203f
C4121 vdd.n3373 gnd 0.009017f
C4122 vdd.n3374 gnd 0.009017f
C4123 vdd.n3375 gnd 0.009017f
C4124 vdd.n3376 gnd 0.011203f
C4125 vdd.n3377 gnd 0.681219f
C4126 vdd.n3378 gnd 0.841505f
C4127 vdd.t42 gnd 0.572453f
C4128 vdd.n3379 gnd 0.875853f
C4129 vdd.n3380 gnd 0.011203f
C4130 vdd.n3381 gnd 0.009017f
C4131 vdd.n3382 gnd 0.009017f
C4132 vdd.n3383 gnd 0.009017f
C4133 vdd.n3384 gnd 0.011203f
C4134 vdd.n3385 gnd 0.950271f
C4135 vdd.t68 gnd 0.572453f
C4136 vdd.n3386 gnd 0.692668f
C4137 vdd.n3387 gnd 0.830056f
C4138 vdd.n3388 gnd 0.011203f
C4139 vdd.n3389 gnd 0.009017f
C4140 vdd.n3390 gnd 0.009017f
C4141 vdd.n3391 gnd 0.009017f
C4142 vdd.n3392 gnd 0.011203f
C4143 vdd.n3393 gnd 0.635422f
C4144 vdd.t37 gnd 0.572453f
C4145 vdd.n3394 gnd 0.950271f
C4146 vdd.t65 gnd 0.572453f
C4147 vdd.n3395 gnd 0.704117f
C4148 vdd.n3396 gnd 0.011203f
C4149 vdd.n3397 gnd 0.009017f
C4150 vdd.n3398 gnd 0.00861f
C4151 vdd.n3399 gnd 0.660802f
C4152 vdd.n3400 gnd 2.8648f
C4153 a_n7636_8799.t18 gnd 0.112158f
C4154 a_n7636_8799.t13 gnd 0.112158f
C4155 a_n7636_8799.t12 gnd 0.112158f
C4156 a_n7636_8799.n0 gnd 0.993272f
C4157 a_n7636_8799.t28 gnd 0.144203f
C4158 a_n7636_8799.t24 gnd 0.144203f
C4159 a_n7636_8799.n1 gnd 1.13735f
C4160 a_n7636_8799.t2 gnd 0.144203f
C4161 a_n7636_8799.t29 gnd 0.144203f
C4162 a_n7636_8799.n2 gnd 1.13548f
C4163 a_n7636_8799.n3 gnd 1.02066f
C4164 a_n7636_8799.t0 gnd 0.144203f
C4165 a_n7636_8799.t31 gnd 0.144203f
C4166 a_n7636_8799.n4 gnd 1.13548f
C4167 a_n7636_8799.n5 gnd 2.9543f
C4168 a_n7636_8799.t23 gnd 0.144203f
C4169 a_n7636_8799.t25 gnd 0.144203f
C4170 a_n7636_8799.n6 gnd 1.13736f
C4171 a_n7636_8799.t30 gnd 0.144203f
C4172 a_n7636_8799.t26 gnd 0.144203f
C4173 a_n7636_8799.n7 gnd 1.13548f
C4174 a_n7636_8799.n8 gnd 1.02066f
C4175 a_n7636_8799.t1 gnd 0.144203f
C4176 a_n7636_8799.t27 gnd 0.144203f
C4177 a_n7636_8799.n9 gnd 1.13548f
C4178 a_n7636_8799.n10 gnd 1.81319f
C4179 a_n7636_8799.n11 gnd 5.69263f
C4180 a_n7636_8799.n12 gnd 0.051976f
C4181 a_n7636_8799.t128 gnd 0.597934f
C4182 a_n7636_8799.n13 gnd 0.267049f
C4183 a_n7636_8799.n14 gnd 0.051976f
C4184 a_n7636_8799.n15 gnd 0.011794f
C4185 a_n7636_8799.t44 gnd 0.597934f
C4186 a_n7636_8799.n16 gnd 0.051976f
C4187 a_n7636_8799.t65 gnd 0.597934f
C4188 a_n7636_8799.n17 gnd 0.264005f
C4189 a_n7636_8799.t88 gnd 0.597934f
C4190 a_n7636_8799.n18 gnd 0.051976f
C4191 a_n7636_8799.t107 gnd 0.597934f
C4192 a_n7636_8799.n19 gnd 0.264325f
C4193 a_n7636_8799.n20 gnd 0.051976f
C4194 a_n7636_8799.n21 gnd 0.011794f
C4195 a_n7636_8799.t67 gnd 0.597934f
C4196 a_n7636_8799.n22 gnd 0.051976f
C4197 a_n7636_8799.t79 gnd 0.597934f
C4198 a_n7636_8799.n23 gnd 0.267049f
C4199 a_n7636_8799.n24 gnd 0.051976f
C4200 a_n7636_8799.n25 gnd 0.011794f
C4201 a_n7636_8799.t112 gnd 0.597934f
C4202 a_n7636_8799.n26 gnd 0.164205f
C4203 a_n7636_8799.t133 gnd 0.597934f
C4204 a_n7636_8799.t131 gnd 0.609251f
C4205 a_n7636_8799.n27 gnd 0.250658f
C4206 a_n7636_8799.n28 gnd 0.263364f
C4207 a_n7636_8799.n29 gnd 0.011794f
C4208 a_n7636_8799.t83 gnd 0.597934f
C4209 a_n7636_8799.n30 gnd 0.267049f
C4210 a_n7636_8799.n31 gnd 0.051976f
C4211 a_n7636_8799.n32 gnd 0.051976f
C4212 a_n7636_8799.n33 gnd 0.051976f
C4213 a_n7636_8799.n34 gnd 0.264966f
C4214 a_n7636_8799.t129 gnd 0.597934f
C4215 a_n7636_8799.n35 gnd 0.263684f
C4216 a_n7636_8799.n36 gnd 0.011794f
C4217 a_n7636_8799.n37 gnd 0.051976f
C4218 a_n7636_8799.n38 gnd 0.051976f
C4219 a_n7636_8799.n39 gnd 0.051976f
C4220 a_n7636_8799.n40 gnd 0.011794f
C4221 a_n7636_8799.t80 gnd 0.597934f
C4222 a_n7636_8799.n41 gnd 0.264646f
C4223 a_n7636_8799.t110 gnd 0.597934f
C4224 a_n7636_8799.n42 gnd 0.264005f
C4225 a_n7636_8799.n43 gnd 0.051976f
C4226 a_n7636_8799.n44 gnd 0.051976f
C4227 a_n7636_8799.n45 gnd 0.051976f
C4228 a_n7636_8799.n46 gnd 0.267049f
C4229 a_n7636_8799.n47 gnd 0.011794f
C4230 a_n7636_8799.t68 gnd 0.597934f
C4231 a_n7636_8799.n48 gnd 0.264325f
C4232 a_n7636_8799.n49 gnd 0.051976f
C4233 a_n7636_8799.n50 gnd 0.051976f
C4234 a_n7636_8799.n51 gnd 0.051976f
C4235 a_n7636_8799.n52 gnd 0.011794f
C4236 a_n7636_8799.t32 gnd 0.597934f
C4237 a_n7636_8799.n53 gnd 0.267049f
C4238 a_n7636_8799.n54 gnd 0.011794f
C4239 a_n7636_8799.n55 gnd 0.051976f
C4240 a_n7636_8799.n56 gnd 0.051976f
C4241 a_n7636_8799.n57 gnd 0.051976f
C4242 a_n7636_8799.n58 gnd 0.264646f
C4243 a_n7636_8799.n59 gnd 0.011794f
C4244 a_n7636_8799.t132 gnd 0.597934f
C4245 a_n7636_8799.n60 gnd 0.267049f
C4246 a_n7636_8799.n61 gnd 0.051976f
C4247 a_n7636_8799.n62 gnd 0.051976f
C4248 a_n7636_8799.n63 gnd 0.051976f
C4249 a_n7636_8799.n64 gnd 0.263684f
C4250 a_n7636_8799.t62 gnd 0.597934f
C4251 a_n7636_8799.n65 gnd 0.264966f
C4252 a_n7636_8799.n66 gnd 0.011794f
C4253 a_n7636_8799.n67 gnd 0.051976f
C4254 a_n7636_8799.n68 gnd 0.051976f
C4255 a_n7636_8799.n69 gnd 0.051976f
C4256 a_n7636_8799.n70 gnd 0.011794f
C4257 a_n7636_8799.t41 gnd 0.597934f
C4258 a_n7636_8799.n71 gnd 0.263364f
C4259 a_n7636_8799.t42 gnd 0.597934f
C4260 a_n7636_8799.n72 gnd 0.261601f
C4261 a_n7636_8799.n73 gnd 0.294688f
C4262 a_n7636_8799.n74 gnd 0.051976f
C4263 a_n7636_8799.t141 gnd 0.597934f
C4264 a_n7636_8799.n75 gnd 0.267049f
C4265 a_n7636_8799.n76 gnd 0.051976f
C4266 a_n7636_8799.n77 gnd 0.011794f
C4267 a_n7636_8799.t59 gnd 0.597934f
C4268 a_n7636_8799.n78 gnd 0.051976f
C4269 a_n7636_8799.t74 gnd 0.597934f
C4270 a_n7636_8799.n79 gnd 0.264005f
C4271 a_n7636_8799.t101 gnd 0.597934f
C4272 a_n7636_8799.n80 gnd 0.051976f
C4273 a_n7636_8799.t119 gnd 0.597934f
C4274 a_n7636_8799.n81 gnd 0.264325f
C4275 a_n7636_8799.n82 gnd 0.051976f
C4276 a_n7636_8799.n83 gnd 0.011794f
C4277 a_n7636_8799.t77 gnd 0.597934f
C4278 a_n7636_8799.n84 gnd 0.051976f
C4279 a_n7636_8799.t89 gnd 0.597934f
C4280 a_n7636_8799.n85 gnd 0.267049f
C4281 a_n7636_8799.n86 gnd 0.051976f
C4282 a_n7636_8799.n87 gnd 0.011794f
C4283 a_n7636_8799.t125 gnd 0.597934f
C4284 a_n7636_8799.n88 gnd 0.164205f
C4285 a_n7636_8799.t149 gnd 0.597934f
C4286 a_n7636_8799.t146 gnd 0.609251f
C4287 a_n7636_8799.n89 gnd 0.250658f
C4288 a_n7636_8799.n90 gnd 0.263364f
C4289 a_n7636_8799.n91 gnd 0.011794f
C4290 a_n7636_8799.t93 gnd 0.597934f
C4291 a_n7636_8799.n92 gnd 0.267049f
C4292 a_n7636_8799.n93 gnd 0.051976f
C4293 a_n7636_8799.n94 gnd 0.051976f
C4294 a_n7636_8799.n95 gnd 0.051976f
C4295 a_n7636_8799.n96 gnd 0.264966f
C4296 a_n7636_8799.t143 gnd 0.597934f
C4297 a_n7636_8799.n97 gnd 0.263684f
C4298 a_n7636_8799.n98 gnd 0.011794f
C4299 a_n7636_8799.n99 gnd 0.051976f
C4300 a_n7636_8799.n100 gnd 0.051976f
C4301 a_n7636_8799.n101 gnd 0.051976f
C4302 a_n7636_8799.n102 gnd 0.011794f
C4303 a_n7636_8799.t90 gnd 0.597934f
C4304 a_n7636_8799.n103 gnd 0.264646f
C4305 a_n7636_8799.t123 gnd 0.597934f
C4306 a_n7636_8799.n104 gnd 0.264005f
C4307 a_n7636_8799.n105 gnd 0.051976f
C4308 a_n7636_8799.n106 gnd 0.051976f
C4309 a_n7636_8799.n107 gnd 0.051976f
C4310 a_n7636_8799.n108 gnd 0.267049f
C4311 a_n7636_8799.n109 gnd 0.011794f
C4312 a_n7636_8799.t78 gnd 0.597934f
C4313 a_n7636_8799.n110 gnd 0.264325f
C4314 a_n7636_8799.n111 gnd 0.051976f
C4315 a_n7636_8799.n112 gnd 0.051976f
C4316 a_n7636_8799.n113 gnd 0.051976f
C4317 a_n7636_8799.n114 gnd 0.011794f
C4318 a_n7636_8799.t43 gnd 0.597934f
C4319 a_n7636_8799.n115 gnd 0.267049f
C4320 a_n7636_8799.n116 gnd 0.011794f
C4321 a_n7636_8799.n117 gnd 0.051976f
C4322 a_n7636_8799.n118 gnd 0.051976f
C4323 a_n7636_8799.n119 gnd 0.051976f
C4324 a_n7636_8799.n120 gnd 0.264646f
C4325 a_n7636_8799.n121 gnd 0.011794f
C4326 a_n7636_8799.t147 gnd 0.597934f
C4327 a_n7636_8799.n122 gnd 0.267049f
C4328 a_n7636_8799.n123 gnd 0.051976f
C4329 a_n7636_8799.n124 gnd 0.051976f
C4330 a_n7636_8799.n125 gnd 0.051976f
C4331 a_n7636_8799.n126 gnd 0.263684f
C4332 a_n7636_8799.t73 gnd 0.597934f
C4333 a_n7636_8799.n127 gnd 0.264966f
C4334 a_n7636_8799.n128 gnd 0.011794f
C4335 a_n7636_8799.n129 gnd 0.051976f
C4336 a_n7636_8799.n130 gnd 0.051976f
C4337 a_n7636_8799.n131 gnd 0.051976f
C4338 a_n7636_8799.n132 gnd 0.011794f
C4339 a_n7636_8799.t53 gnd 0.597934f
C4340 a_n7636_8799.n133 gnd 0.263364f
C4341 a_n7636_8799.t55 gnd 0.597934f
C4342 a_n7636_8799.n134 gnd 0.261601f
C4343 a_n7636_8799.n135 gnd 0.12955f
C4344 a_n7636_8799.n136 gnd 0.898911f
C4345 a_n7636_8799.n137 gnd 0.051976f
C4346 a_n7636_8799.t96 gnd 0.597934f
C4347 a_n7636_8799.n138 gnd 0.267049f
C4348 a_n7636_8799.n139 gnd 0.051976f
C4349 a_n7636_8799.n140 gnd 0.011794f
C4350 a_n7636_8799.t120 gnd 0.597934f
C4351 a_n7636_8799.n141 gnd 0.051976f
C4352 a_n7636_8799.t38 gnd 0.597934f
C4353 a_n7636_8799.n142 gnd 0.264005f
C4354 a_n7636_8799.t103 gnd 0.597934f
C4355 a_n7636_8799.n143 gnd 0.051976f
C4356 a_n7636_8799.t142 gnd 0.597934f
C4357 a_n7636_8799.n144 gnd 0.264325f
C4358 a_n7636_8799.n145 gnd 0.051976f
C4359 a_n7636_8799.n146 gnd 0.011794f
C4360 a_n7636_8799.t137 gnd 0.597934f
C4361 a_n7636_8799.n147 gnd 0.051976f
C4362 a_n7636_8799.t50 gnd 0.597934f
C4363 a_n7636_8799.n148 gnd 0.267049f
C4364 a_n7636_8799.n149 gnd 0.051976f
C4365 a_n7636_8799.n150 gnd 0.011794f
C4366 a_n7636_8799.t75 gnd 0.597934f
C4367 a_n7636_8799.n151 gnd 0.164205f
C4368 a_n7636_8799.t86 gnd 0.597934f
C4369 a_n7636_8799.t108 gnd 0.609251f
C4370 a_n7636_8799.n152 gnd 0.250658f
C4371 a_n7636_8799.n153 gnd 0.263364f
C4372 a_n7636_8799.n154 gnd 0.011794f
C4373 a_n7636_8799.t124 gnd 0.597934f
C4374 a_n7636_8799.n155 gnd 0.267049f
C4375 a_n7636_8799.n156 gnd 0.051976f
C4376 a_n7636_8799.n157 gnd 0.051976f
C4377 a_n7636_8799.n158 gnd 0.051976f
C4378 a_n7636_8799.n159 gnd 0.264966f
C4379 a_n7636_8799.t134 gnd 0.597934f
C4380 a_n7636_8799.n160 gnd 0.263684f
C4381 a_n7636_8799.n161 gnd 0.011794f
C4382 a_n7636_8799.n162 gnd 0.051976f
C4383 a_n7636_8799.n163 gnd 0.051976f
C4384 a_n7636_8799.n164 gnd 0.051976f
C4385 a_n7636_8799.n165 gnd 0.011794f
C4386 a_n7636_8799.t33 gnd 0.597934f
C4387 a_n7636_8799.n166 gnd 0.264646f
C4388 a_n7636_8799.t94 gnd 0.597934f
C4389 a_n7636_8799.n167 gnd 0.264005f
C4390 a_n7636_8799.n168 gnd 0.051976f
C4391 a_n7636_8799.n169 gnd 0.051976f
C4392 a_n7636_8799.n170 gnd 0.051976f
C4393 a_n7636_8799.n171 gnd 0.267049f
C4394 a_n7636_8799.n172 gnd 0.011794f
C4395 a_n7636_8799.t111 gnd 0.597934f
C4396 a_n7636_8799.n173 gnd 0.264325f
C4397 a_n7636_8799.n174 gnd 0.051976f
C4398 a_n7636_8799.n175 gnd 0.051976f
C4399 a_n7636_8799.n176 gnd 0.051976f
C4400 a_n7636_8799.n177 gnd 0.011794f
C4401 a_n7636_8799.t87 gnd 0.597934f
C4402 a_n7636_8799.n178 gnd 0.267049f
C4403 a_n7636_8799.n179 gnd 0.011794f
C4404 a_n7636_8799.n180 gnd 0.051976f
C4405 a_n7636_8799.n181 gnd 0.051976f
C4406 a_n7636_8799.n182 gnd 0.051976f
C4407 a_n7636_8799.n183 gnd 0.264646f
C4408 a_n7636_8799.n184 gnd 0.011794f
C4409 a_n7636_8799.t57 gnd 0.597934f
C4410 a_n7636_8799.n185 gnd 0.267049f
C4411 a_n7636_8799.n186 gnd 0.051976f
C4412 a_n7636_8799.n187 gnd 0.051976f
C4413 a_n7636_8799.n188 gnd 0.051976f
C4414 a_n7636_8799.n189 gnd 0.263684f
C4415 a_n7636_8799.t66 gnd 0.597934f
C4416 a_n7636_8799.n190 gnd 0.264966f
C4417 a_n7636_8799.n191 gnd 0.011794f
C4418 a_n7636_8799.n192 gnd 0.051976f
C4419 a_n7636_8799.n193 gnd 0.051976f
C4420 a_n7636_8799.n194 gnd 0.051976f
C4421 a_n7636_8799.n195 gnd 0.011794f
C4422 a_n7636_8799.t46 gnd 0.597934f
C4423 a_n7636_8799.n196 gnd 0.263364f
C4424 a_n7636_8799.t148 gnd 0.597934f
C4425 a_n7636_8799.n197 gnd 0.261601f
C4426 a_n7636_8799.n198 gnd 0.12955f
C4427 a_n7636_8799.n199 gnd 1.45959f
C4428 a_n7636_8799.n200 gnd 0.051976f
C4429 a_n7636_8799.t82 gnd 0.597934f
C4430 a_n7636_8799.t81 gnd 0.597934f
C4431 a_n7636_8799.t54 gnd 0.597934f
C4432 a_n7636_8799.n201 gnd 0.267049f
C4433 a_n7636_8799.n202 gnd 0.051976f
C4434 a_n7636_8799.t130 gnd 0.597934f
C4435 a_n7636_8799.t85 gnd 0.597934f
C4436 a_n7636_8799.n203 gnd 0.051976f
C4437 a_n7636_8799.t61 gnd 0.597934f
C4438 a_n7636_8799.n204 gnd 0.267049f
C4439 a_n7636_8799.n205 gnd 0.051976f
C4440 a_n7636_8799.t136 gnd 0.597934f
C4441 a_n7636_8799.t102 gnd 0.597934f
C4442 a_n7636_8799.n206 gnd 0.051976f
C4443 a_n7636_8799.t100 gnd 0.597934f
C4444 a_n7636_8799.n207 gnd 0.267049f
C4445 a_n7636_8799.n208 gnd 0.051976f
C4446 a_n7636_8799.t35 gnd 0.597934f
C4447 a_n7636_8799.t106 gnd 0.597934f
C4448 a_n7636_8799.n209 gnd 0.051976f
C4449 a_n7636_8799.t105 gnd 0.597934f
C4450 a_n7636_8799.n210 gnd 0.267049f
C4451 a_n7636_8799.n211 gnd 0.051976f
C4452 a_n7636_8799.t37 gnd 0.597934f
C4453 a_n7636_8799.t36 gnd 0.597934f
C4454 a_n7636_8799.n212 gnd 0.051976f
C4455 a_n7636_8799.t122 gnd 0.597934f
C4456 a_n7636_8799.n213 gnd 0.267049f
C4457 a_n7636_8799.n214 gnd 0.051976f
C4458 a_n7636_8799.t56 gnd 0.597934f
C4459 a_n7636_8799.t40 gnd 0.597934f
C4460 a_n7636_8799.n215 gnd 0.051976f
C4461 a_n7636_8799.t126 gnd 0.597934f
C4462 a_n7636_8799.n216 gnd 0.267049f
C4463 a_n7636_8799.t60 gnd 0.609251f
C4464 a_n7636_8799.n217 gnd 0.250658f
C4465 a_n7636_8799.t84 gnd 0.597934f
C4466 a_n7636_8799.n218 gnd 0.263364f
C4467 a_n7636_8799.n219 gnd 0.011794f
C4468 a_n7636_8799.n220 gnd 0.164205f
C4469 a_n7636_8799.n221 gnd 0.051976f
C4470 a_n7636_8799.n222 gnd 0.051976f
C4471 a_n7636_8799.n223 gnd 0.011794f
C4472 a_n7636_8799.n224 gnd 0.264966f
C4473 a_n7636_8799.n225 gnd 0.263684f
C4474 a_n7636_8799.n226 gnd 0.011794f
C4475 a_n7636_8799.n227 gnd 0.051976f
C4476 a_n7636_8799.n228 gnd 0.051976f
C4477 a_n7636_8799.n229 gnd 0.051976f
C4478 a_n7636_8799.n230 gnd 0.011794f
C4479 a_n7636_8799.n231 gnd 0.264646f
C4480 a_n7636_8799.n232 gnd 0.264005f
C4481 a_n7636_8799.n233 gnd 0.011794f
C4482 a_n7636_8799.n234 gnd 0.051976f
C4483 a_n7636_8799.n235 gnd 0.051976f
C4484 a_n7636_8799.n236 gnd 0.051976f
C4485 a_n7636_8799.n237 gnd 0.011794f
C4486 a_n7636_8799.n238 gnd 0.264325f
C4487 a_n7636_8799.n239 gnd 0.264325f
C4488 a_n7636_8799.n240 gnd 0.011794f
C4489 a_n7636_8799.n241 gnd 0.051976f
C4490 a_n7636_8799.n242 gnd 0.051976f
C4491 a_n7636_8799.n243 gnd 0.051976f
C4492 a_n7636_8799.n244 gnd 0.011794f
C4493 a_n7636_8799.n245 gnd 0.264005f
C4494 a_n7636_8799.n246 gnd 0.264646f
C4495 a_n7636_8799.n247 gnd 0.011794f
C4496 a_n7636_8799.n248 gnd 0.051976f
C4497 a_n7636_8799.n249 gnd 0.051976f
C4498 a_n7636_8799.n250 gnd 0.051976f
C4499 a_n7636_8799.n251 gnd 0.011794f
C4500 a_n7636_8799.n252 gnd 0.263684f
C4501 a_n7636_8799.n253 gnd 0.264966f
C4502 a_n7636_8799.n254 gnd 0.011794f
C4503 a_n7636_8799.n255 gnd 0.051976f
C4504 a_n7636_8799.n256 gnd 0.051976f
C4505 a_n7636_8799.n257 gnd 0.051976f
C4506 a_n7636_8799.n258 gnd 0.011794f
C4507 a_n7636_8799.n259 gnd 0.263364f
C4508 a_n7636_8799.n260 gnd 0.261601f
C4509 a_n7636_8799.n261 gnd 0.294688f
C4510 a_n7636_8799.n262 gnd 0.051976f
C4511 a_n7636_8799.t92 gnd 0.597934f
C4512 a_n7636_8799.t91 gnd 0.597934f
C4513 a_n7636_8799.t69 gnd 0.597934f
C4514 a_n7636_8799.n263 gnd 0.267049f
C4515 a_n7636_8799.n264 gnd 0.051976f
C4516 a_n7636_8799.t145 gnd 0.597934f
C4517 a_n7636_8799.t98 gnd 0.597934f
C4518 a_n7636_8799.n265 gnd 0.051976f
C4519 a_n7636_8799.t71 gnd 0.597934f
C4520 a_n7636_8799.n266 gnd 0.267049f
C4521 a_n7636_8799.n267 gnd 0.051976f
C4522 a_n7636_8799.t151 gnd 0.597934f
C4523 a_n7636_8799.t115 gnd 0.597934f
C4524 a_n7636_8799.n268 gnd 0.051976f
C4525 a_n7636_8799.t114 gnd 0.597934f
C4526 a_n7636_8799.n269 gnd 0.267049f
C4527 a_n7636_8799.n270 gnd 0.051976f
C4528 a_n7636_8799.t45 gnd 0.597934f
C4529 a_n7636_8799.t118 gnd 0.597934f
C4530 a_n7636_8799.n271 gnd 0.051976f
C4531 a_n7636_8799.t117 gnd 0.597934f
C4532 a_n7636_8799.n272 gnd 0.267049f
C4533 a_n7636_8799.n273 gnd 0.051976f
C4534 a_n7636_8799.t49 gnd 0.597934f
C4535 a_n7636_8799.t48 gnd 0.597934f
C4536 a_n7636_8799.n274 gnd 0.051976f
C4537 a_n7636_8799.t139 gnd 0.597934f
C4538 a_n7636_8799.n275 gnd 0.267049f
C4539 a_n7636_8799.n276 gnd 0.051976f
C4540 a_n7636_8799.t70 gnd 0.597934f
C4541 a_n7636_8799.t52 gnd 0.597934f
C4542 a_n7636_8799.n277 gnd 0.051976f
C4543 a_n7636_8799.t140 gnd 0.597934f
C4544 a_n7636_8799.n278 gnd 0.267049f
C4545 a_n7636_8799.t72 gnd 0.609251f
C4546 a_n7636_8799.n279 gnd 0.250658f
C4547 a_n7636_8799.t99 gnd 0.597934f
C4548 a_n7636_8799.n280 gnd 0.263364f
C4549 a_n7636_8799.n281 gnd 0.011794f
C4550 a_n7636_8799.n282 gnd 0.164205f
C4551 a_n7636_8799.n283 gnd 0.051976f
C4552 a_n7636_8799.n284 gnd 0.051976f
C4553 a_n7636_8799.n285 gnd 0.011794f
C4554 a_n7636_8799.n286 gnd 0.264966f
C4555 a_n7636_8799.n287 gnd 0.263684f
C4556 a_n7636_8799.n288 gnd 0.011794f
C4557 a_n7636_8799.n289 gnd 0.051976f
C4558 a_n7636_8799.n290 gnd 0.051976f
C4559 a_n7636_8799.n291 gnd 0.051976f
C4560 a_n7636_8799.n292 gnd 0.011794f
C4561 a_n7636_8799.n293 gnd 0.264646f
C4562 a_n7636_8799.n294 gnd 0.264005f
C4563 a_n7636_8799.n295 gnd 0.011794f
C4564 a_n7636_8799.n296 gnd 0.051976f
C4565 a_n7636_8799.n297 gnd 0.051976f
C4566 a_n7636_8799.n298 gnd 0.051976f
C4567 a_n7636_8799.n299 gnd 0.011794f
C4568 a_n7636_8799.n300 gnd 0.264325f
C4569 a_n7636_8799.n301 gnd 0.264325f
C4570 a_n7636_8799.n302 gnd 0.011794f
C4571 a_n7636_8799.n303 gnd 0.051976f
C4572 a_n7636_8799.n304 gnd 0.051976f
C4573 a_n7636_8799.n305 gnd 0.051976f
C4574 a_n7636_8799.n306 gnd 0.011794f
C4575 a_n7636_8799.n307 gnd 0.264005f
C4576 a_n7636_8799.n308 gnd 0.264646f
C4577 a_n7636_8799.n309 gnd 0.011794f
C4578 a_n7636_8799.n310 gnd 0.051976f
C4579 a_n7636_8799.n311 gnd 0.051976f
C4580 a_n7636_8799.n312 gnd 0.051976f
C4581 a_n7636_8799.n313 gnd 0.011794f
C4582 a_n7636_8799.n314 gnd 0.263684f
C4583 a_n7636_8799.n315 gnd 0.264966f
C4584 a_n7636_8799.n316 gnd 0.011794f
C4585 a_n7636_8799.n317 gnd 0.051976f
C4586 a_n7636_8799.n318 gnd 0.051976f
C4587 a_n7636_8799.n319 gnd 0.051976f
C4588 a_n7636_8799.n320 gnd 0.011794f
C4589 a_n7636_8799.n321 gnd 0.263364f
C4590 a_n7636_8799.n322 gnd 0.261601f
C4591 a_n7636_8799.n323 gnd 0.12955f
C4592 a_n7636_8799.n324 gnd 0.898911f
C4593 a_n7636_8799.n325 gnd 0.051976f
C4594 a_n7636_8799.t150 gnd 0.597934f
C4595 a_n7636_8799.t47 gnd 0.597934f
C4596 a_n7636_8799.t97 gnd 0.597934f
C4597 a_n7636_8799.n326 gnd 0.267049f
C4598 a_n7636_8799.n327 gnd 0.051976f
C4599 a_n7636_8799.t34 gnd 0.597934f
C4600 a_n7636_8799.t121 gnd 0.597934f
C4601 a_n7636_8799.n328 gnd 0.051976f
C4602 a_n7636_8799.t58 gnd 0.597934f
C4603 a_n7636_8799.n329 gnd 0.267049f
C4604 a_n7636_8799.n330 gnd 0.051976f
C4605 a_n7636_8799.t104 gnd 0.597934f
C4606 a_n7636_8799.t39 gnd 0.597934f
C4607 a_n7636_8799.n331 gnd 0.051976f
C4608 a_n7636_8799.t64 gnd 0.597934f
C4609 a_n7636_8799.n332 gnd 0.267049f
C4610 a_n7636_8799.n333 gnd 0.051976f
C4611 a_n7636_8799.t144 gnd 0.597934f
C4612 a_n7636_8799.t113 gnd 0.597934f
C4613 a_n7636_8799.n334 gnd 0.051976f
C4614 a_n7636_8799.t138 gnd 0.597934f
C4615 a_n7636_8799.n335 gnd 0.267049f
C4616 a_n7636_8799.n336 gnd 0.051976f
C4617 a_n7636_8799.t95 gnd 0.597934f
C4618 a_n7636_8799.t116 gnd 0.597934f
C4619 a_n7636_8799.n337 gnd 0.051976f
C4620 a_n7636_8799.t51 gnd 0.597934f
C4621 a_n7636_8799.n338 gnd 0.267049f
C4622 a_n7636_8799.n339 gnd 0.051976f
C4623 a_n7636_8799.t135 gnd 0.597934f
C4624 a_n7636_8799.t76 gnd 0.597934f
C4625 a_n7636_8799.n340 gnd 0.051976f
C4626 a_n7636_8799.t127 gnd 0.597934f
C4627 a_n7636_8799.n341 gnd 0.267049f
C4628 a_n7636_8799.t109 gnd 0.609251f
C4629 a_n7636_8799.n342 gnd 0.250658f
C4630 a_n7636_8799.t63 gnd 0.597934f
C4631 a_n7636_8799.n343 gnd 0.263364f
C4632 a_n7636_8799.n344 gnd 0.011794f
C4633 a_n7636_8799.n345 gnd 0.164205f
C4634 a_n7636_8799.n346 gnd 0.051976f
C4635 a_n7636_8799.n347 gnd 0.051976f
C4636 a_n7636_8799.n348 gnd 0.011794f
C4637 a_n7636_8799.n349 gnd 0.264966f
C4638 a_n7636_8799.n350 gnd 0.263684f
C4639 a_n7636_8799.n351 gnd 0.011794f
C4640 a_n7636_8799.n352 gnd 0.051976f
C4641 a_n7636_8799.n353 gnd 0.051976f
C4642 a_n7636_8799.n354 gnd 0.051976f
C4643 a_n7636_8799.n355 gnd 0.011794f
C4644 a_n7636_8799.n356 gnd 0.264646f
C4645 a_n7636_8799.n357 gnd 0.264005f
C4646 a_n7636_8799.n358 gnd 0.011794f
C4647 a_n7636_8799.n359 gnd 0.051976f
C4648 a_n7636_8799.n360 gnd 0.051976f
C4649 a_n7636_8799.n361 gnd 0.051976f
C4650 a_n7636_8799.n362 gnd 0.011794f
C4651 a_n7636_8799.n363 gnd 0.264325f
C4652 a_n7636_8799.n364 gnd 0.264325f
C4653 a_n7636_8799.n365 gnd 0.011794f
C4654 a_n7636_8799.n366 gnd 0.051976f
C4655 a_n7636_8799.n367 gnd 0.051976f
C4656 a_n7636_8799.n368 gnd 0.051976f
C4657 a_n7636_8799.n369 gnd 0.011794f
C4658 a_n7636_8799.n370 gnd 0.264005f
C4659 a_n7636_8799.n371 gnd 0.264646f
C4660 a_n7636_8799.n372 gnd 0.011794f
C4661 a_n7636_8799.n373 gnd 0.051976f
C4662 a_n7636_8799.n374 gnd 0.051976f
C4663 a_n7636_8799.n375 gnd 0.051976f
C4664 a_n7636_8799.n376 gnd 0.011794f
C4665 a_n7636_8799.n377 gnd 0.263684f
C4666 a_n7636_8799.n378 gnd 0.264966f
C4667 a_n7636_8799.n379 gnd 0.011794f
C4668 a_n7636_8799.n380 gnd 0.051976f
C4669 a_n7636_8799.n381 gnd 0.051976f
C4670 a_n7636_8799.n382 gnd 0.051976f
C4671 a_n7636_8799.n383 gnd 0.011794f
C4672 a_n7636_8799.n384 gnd 0.263364f
C4673 a_n7636_8799.n385 gnd 0.261601f
C4674 a_n7636_8799.n386 gnd 0.12955f
C4675 a_n7636_8799.n387 gnd 1.133f
C4676 a_n7636_8799.n388 gnd 12.2459f
C4677 a_n7636_8799.n389 gnd 4.37601f
C4678 a_n7636_8799.t9 gnd 0.112158f
C4679 a_n7636_8799.t10 gnd 0.112158f
C4680 a_n7636_8799.n390 gnd 0.993273f
C4681 a_n7636_8799.t5 gnd 0.112158f
C4682 a_n7636_8799.t6 gnd 0.112158f
C4683 a_n7636_8799.n391 gnd 0.991069f
C4684 a_n7636_8799.n392 gnd 0.789432f
C4685 a_n7636_8799.t4 gnd 0.112158f
C4686 a_n7636_8799.t19 gnd 0.112158f
C4687 a_n7636_8799.n393 gnd 0.991069f
C4688 a_n7636_8799.n394 gnd 0.742248f
C4689 a_n7636_8799.t20 gnd 0.112158f
C4690 a_n7636_8799.t15 gnd 0.112158f
C4691 a_n7636_8799.n395 gnd 0.991069f
C4692 a_n7636_8799.n396 gnd 0.387651f
C4693 a_n7636_8799.t17 gnd 0.112158f
C4694 a_n7636_8799.t3 gnd 0.112158f
C4695 a_n7636_8799.n397 gnd 0.991069f
C4696 a_n7636_8799.n398 gnd 2.7113f
C4697 a_n7636_8799.t16 gnd 0.112158f
C4698 a_n7636_8799.t14 gnd 0.112158f
C4699 a_n7636_8799.n399 gnd 0.993272f
C4700 a_n7636_8799.t7 gnd 0.112158f
C4701 a_n7636_8799.t11 gnd 0.112158f
C4702 a_n7636_8799.n400 gnd 0.991068f
C4703 a_n7636_8799.n401 gnd 0.789434f
C4704 a_n7636_8799.t21 gnd 0.112158f
C4705 a_n7636_8799.t8 gnd 0.112158f
C4706 a_n7636_8799.n402 gnd 0.991068f
C4707 a_n7636_8799.n403 gnd 2.46819f
C4708 a_n7636_8799.n404 gnd 0.789436f
C4709 a_n7636_8799.n405 gnd 0.991066f
C4710 a_n7636_8799.t22 gnd 0.112158f
C4711 a_n2903_n3924.n0 gnd 1.27336f
C4712 a_n2903_n3924.n1 gnd 1.81293f
C4713 a_n2903_n3924.n2 gnd 0.724065f
C4714 a_n2903_n3924.n3 gnd 1.63539f
C4715 a_n2903_n3924.n4 gnd 2.17497f
C4716 a_n2903_n3924.n5 gnd 1.67866f
C4717 a_n2903_n3924.n6 gnd 0.954594f
C4718 a_n2903_n3924.n7 gnd 1.7731f
C4719 a_n2903_n3924.n8 gnd 1.7731f
C4720 a_n2903_n3924.n9 gnd 2.13362f
C4721 a_n2903_n3924.n10 gnd 1.60399f
C4722 a_n2903_n3924.t41 gnd 0.097476f
C4723 a_n2903_n3924.t36 gnd 0.097476f
C4724 a_n2903_n3924.t42 gnd 0.097476f
C4725 a_n2903_n3924.n11 gnd 0.796106f
C4726 a_n2903_n3924.t2 gnd 1.25909f
C4727 a_n2903_n3924.t34 gnd 0.097476f
C4728 a_n2903_n3924.t10 gnd 0.097476f
C4729 a_n2903_n3924.n12 gnd 0.796106f
C4730 a_n2903_n3924.t7 gnd 0.097476f
C4731 a_n2903_n3924.t9 gnd 0.097476f
C4732 a_n2903_n3924.n13 gnd 0.796106f
C4733 a_n2903_n3924.t45 gnd 1.01309f
C4734 a_n2903_n3924.t31 gnd 1.26033f
C4735 a_n2903_n3924.t46 gnd 1.25874f
C4736 a_n2903_n3924.t0 gnd 1.25874f
C4737 a_n2903_n3924.t47 gnd 1.25874f
C4738 a_n2903_n3924.t35 gnd 1.25874f
C4739 a_n2903_n3924.t37 gnd 1.25874f
C4740 a_n2903_n3924.t8 gnd 1.25874f
C4741 a_n2903_n3924.n14 gnd 0.914361f
C4742 a_n2903_n3924.t22 gnd 1.01309f
C4743 a_n2903_n3924.t13 gnd 0.097476f
C4744 a_n2903_n3924.t25 gnd 0.097476f
C4745 a_n2903_n3924.n15 gnd 0.796105f
C4746 a_n2903_n3924.t23 gnd 0.097476f
C4747 a_n2903_n3924.t12 gnd 0.097476f
C4748 a_n2903_n3924.n16 gnd 0.796105f
C4749 a_n2903_n3924.t21 gnd 0.097476f
C4750 a_n2903_n3924.t20 gnd 0.097476f
C4751 a_n2903_n3924.n17 gnd 0.796105f
C4752 a_n2903_n3924.t30 gnd 0.097476f
C4753 a_n2903_n3924.t27 gnd 0.097476f
C4754 a_n2903_n3924.n18 gnd 0.796105f
C4755 a_n2903_n3924.t16 gnd 1.01309f
C4756 a_n2903_n3924.t32 gnd 1.01309f
C4757 a_n2903_n3924.t3 gnd 0.097476f
C4758 a_n2903_n3924.t6 gnd 0.097476f
C4759 a_n2903_n3924.n19 gnd 0.796105f
C4760 a_n2903_n3924.t4 gnd 0.097476f
C4761 a_n2903_n3924.t39 gnd 0.097476f
C4762 a_n2903_n3924.n20 gnd 0.796105f
C4763 a_n2903_n3924.t38 gnd 0.097476f
C4764 a_n2903_n3924.t33 gnd 0.097476f
C4765 a_n2903_n3924.n21 gnd 0.796105f
C4766 a_n2903_n3924.t44 gnd 0.097476f
C4767 a_n2903_n3924.t43 gnd 0.097476f
C4768 a_n2903_n3924.n22 gnd 0.796105f
C4769 a_n2903_n3924.t5 gnd 1.01309f
C4770 a_n2903_n3924.n23 gnd 0.914361f
C4771 a_n2903_n3924.t29 gnd 1.01309f
C4772 a_n2903_n3924.t18 gnd 0.097476f
C4773 a_n2903_n3924.t24 gnd 0.097476f
C4774 a_n2903_n3924.n24 gnd 0.796106f
C4775 a_n2903_n3924.t28 gnd 0.097476f
C4776 a_n2903_n3924.t26 gnd 0.097476f
C4777 a_n2903_n3924.n25 gnd 0.796106f
C4778 a_n2903_n3924.t17 gnd 0.097476f
C4779 a_n2903_n3924.t19 gnd 0.097476f
C4780 a_n2903_n3924.n26 gnd 0.796106f
C4781 a_n2903_n3924.t11 gnd 0.097476f
C4782 a_n2903_n3924.t15 gnd 0.097476f
C4783 a_n2903_n3924.n27 gnd 0.796106f
C4784 a_n2903_n3924.t14 gnd 1.01309f
C4785 a_n2903_n3924.t40 gnd 1.01309f
C4786 a_n2903_n3924.n28 gnd 0.796107f
C4787 a_n2903_n3924.t1 gnd 0.097476f
C4788 plus.n0 gnd 0.023146f
C4789 plus.t14 gnd 0.327377f
C4790 plus.n1 gnd 0.023146f
C4791 plus.t15 gnd 0.327377f
C4792 plus.t9 gnd 0.327377f
C4793 plus.n2 gnd 0.145431f
C4794 plus.n3 gnd 0.023146f
C4795 plus.t5 gnd 0.327377f
C4796 plus.t6 gnd 0.327377f
C4797 plus.n4 gnd 0.145431f
C4798 plus.n5 gnd 0.023146f
C4799 plus.t19 gnd 0.327377f
C4800 plus.t20 gnd 0.327377f
C4801 plus.n6 gnd 0.145431f
C4802 plus.n7 gnd 0.023146f
C4803 plus.t16 gnd 0.327377f
C4804 plus.t11 gnd 0.327377f
C4805 plus.n8 gnd 0.149303f
C4806 plus.t13 gnd 0.338846f
C4807 plus.n9 gnd 0.135624f
C4808 plus.n10 gnd 0.098796f
C4809 plus.n11 gnd 0.005252f
C4810 plus.n12 gnd 0.145431f
C4811 plus.n13 gnd 0.005252f
C4812 plus.n14 gnd 0.023146f
C4813 plus.n15 gnd 0.023146f
C4814 plus.n16 gnd 0.023146f
C4815 plus.n17 gnd 0.005252f
C4816 plus.n18 gnd 0.145431f
C4817 plus.n19 gnd 0.005252f
C4818 plus.n20 gnd 0.023146f
C4819 plus.n21 gnd 0.023146f
C4820 plus.n22 gnd 0.023146f
C4821 plus.n23 gnd 0.005252f
C4822 plus.n24 gnd 0.145431f
C4823 plus.n25 gnd 0.005252f
C4824 plus.n26 gnd 0.023146f
C4825 plus.n27 gnd 0.023146f
C4826 plus.n28 gnd 0.023146f
C4827 plus.n29 gnd 0.005252f
C4828 plus.n30 gnd 0.145431f
C4829 plus.n31 gnd 0.005252f
C4830 plus.n32 gnd 0.145217f
C4831 plus.n33 gnd 0.26147f
C4832 plus.n34 gnd 0.023146f
C4833 plus.n35 gnd 0.005252f
C4834 plus.t10 gnd 0.327377f
C4835 plus.n36 gnd 0.023146f
C4836 plus.n37 gnd 0.005252f
C4837 plus.t7 gnd 0.327377f
C4838 plus.n38 gnd 0.023146f
C4839 plus.n39 gnd 0.005252f
C4840 plus.t23 gnd 0.327377f
C4841 plus.n40 gnd 0.023146f
C4842 plus.n41 gnd 0.005252f
C4843 plus.t22 gnd 0.327377f
C4844 plus.t18 gnd 0.338846f
C4845 plus.t17 gnd 0.327377f
C4846 plus.n42 gnd 0.149303f
C4847 plus.n43 gnd 0.135624f
C4848 plus.n44 gnd 0.098796f
C4849 plus.n45 gnd 0.023146f
C4850 plus.n46 gnd 0.145431f
C4851 plus.n47 gnd 0.005252f
C4852 plus.t21 gnd 0.327377f
C4853 plus.n48 gnd 0.145431f
C4854 plus.n49 gnd 0.023146f
C4855 plus.n50 gnd 0.023146f
C4856 plus.n51 gnd 0.023146f
C4857 plus.n52 gnd 0.145431f
C4858 plus.n53 gnd 0.005252f
C4859 plus.t8 gnd 0.327377f
C4860 plus.n54 gnd 0.145431f
C4861 plus.n55 gnd 0.023146f
C4862 plus.n56 gnd 0.023146f
C4863 plus.n57 gnd 0.023146f
C4864 plus.n58 gnd 0.145431f
C4865 plus.n59 gnd 0.005252f
C4866 plus.t12 gnd 0.327377f
C4867 plus.n60 gnd 0.145431f
C4868 plus.n61 gnd 0.023146f
C4869 plus.n62 gnd 0.023146f
C4870 plus.n63 gnd 0.023146f
C4871 plus.n64 gnd 0.145431f
C4872 plus.n65 gnd 0.005252f
C4873 plus.t24 gnd 0.327377f
C4874 plus.n66 gnd 0.145217f
C4875 plus.n67 gnd 0.713957f
C4876 plus.n68 gnd 1.07968f
C4877 plus.t0 gnd 0.039956f
C4878 plus.t4 gnd 0.007135f
C4879 plus.t2 gnd 0.007135f
C4880 plus.n69 gnd 0.023141f
C4881 plus.n70 gnd 0.179643f
C4882 plus.t1 gnd 0.007135f
C4883 plus.t3 gnd 0.007135f
C4884 plus.n71 gnd 0.023141f
C4885 plus.n72 gnd 0.134844f
C4886 plus.n73 gnd 2.61548f
C4887 CSoutput.n0 gnd 0.048499f
C4888 CSoutput.t198 gnd 0.320809f
C4889 CSoutput.n1 gnd 0.144861f
C4890 CSoutput.n2 gnd 0.048499f
C4891 CSoutput.t204 gnd 0.320809f
C4892 CSoutput.n3 gnd 0.038439f
C4893 CSoutput.n4 gnd 0.048499f
C4894 CSoutput.t192 gnd 0.320809f
C4895 CSoutput.n5 gnd 0.033147f
C4896 CSoutput.n6 gnd 0.048499f
C4897 CSoutput.t201 gnd 0.320809f
C4898 CSoutput.t200 gnd 0.320809f
C4899 CSoutput.n7 gnd 0.143283f
C4900 CSoutput.n8 gnd 0.048499f
C4901 CSoutput.t189 gnd 0.320809f
C4902 CSoutput.n9 gnd 0.031603f
C4903 CSoutput.n10 gnd 0.048499f
C4904 CSoutput.t195 gnd 0.320809f
C4905 CSoutput.t197 gnd 0.320809f
C4906 CSoutput.n11 gnd 0.143283f
C4907 CSoutput.n12 gnd 0.048499f
C4908 CSoutput.t187 gnd 0.320809f
C4909 CSoutput.n13 gnd 0.033147f
C4910 CSoutput.n14 gnd 0.048499f
C4911 CSoutput.t185 gnd 0.320809f
C4912 CSoutput.t196 gnd 0.320809f
C4913 CSoutput.n15 gnd 0.143283f
C4914 CSoutput.n16 gnd 0.048499f
C4915 CSoutput.t199 gnd 0.320809f
C4916 CSoutput.n17 gnd 0.035402f
C4917 CSoutput.t188 gnd 0.383375f
C4918 CSoutput.t205 gnd 0.320809f
C4919 CSoutput.n18 gnd 0.182916f
C4920 CSoutput.n19 gnd 0.177492f
C4921 CSoutput.n20 gnd 0.205912f
C4922 CSoutput.n21 gnd 0.048499f
C4923 CSoutput.n22 gnd 0.040478f
C4924 CSoutput.n23 gnd 0.143283f
C4925 CSoutput.n24 gnd 0.039019f
C4926 CSoutput.n25 gnd 0.038439f
C4927 CSoutput.n26 gnd 0.048499f
C4928 CSoutput.n27 gnd 0.048499f
C4929 CSoutput.n28 gnd 0.040166f
C4930 CSoutput.n29 gnd 0.034102f
C4931 CSoutput.n30 gnd 0.146472f
C4932 CSoutput.n31 gnd 0.034572f
C4933 CSoutput.n32 gnd 0.048499f
C4934 CSoutput.n33 gnd 0.048499f
C4935 CSoutput.n34 gnd 0.048499f
C4936 CSoutput.n35 gnd 0.039739f
C4937 CSoutput.n36 gnd 0.143283f
C4938 CSoutput.n37 gnd 0.038004f
C4939 CSoutput.n38 gnd 0.039454f
C4940 CSoutput.n39 gnd 0.048499f
C4941 CSoutput.n40 gnd 0.048499f
C4942 CSoutput.n41 gnd 0.040469f
C4943 CSoutput.n42 gnd 0.036989f
C4944 CSoutput.n43 gnd 0.143283f
C4945 CSoutput.n44 gnd 0.037927f
C4946 CSoutput.n45 gnd 0.048499f
C4947 CSoutput.n46 gnd 0.048499f
C4948 CSoutput.n47 gnd 0.048499f
C4949 CSoutput.n48 gnd 0.037927f
C4950 CSoutput.n49 gnd 0.143283f
C4951 CSoutput.n50 gnd 0.036989f
C4952 CSoutput.n51 gnd 0.040469f
C4953 CSoutput.n52 gnd 0.048499f
C4954 CSoutput.n53 gnd 0.048499f
C4955 CSoutput.n54 gnd 0.039454f
C4956 CSoutput.n55 gnd 0.038004f
C4957 CSoutput.n56 gnd 0.143283f
C4958 CSoutput.n57 gnd 0.039739f
C4959 CSoutput.n58 gnd 0.048499f
C4960 CSoutput.n59 gnd 0.048499f
C4961 CSoutput.n60 gnd 0.048499f
C4962 CSoutput.n61 gnd 0.034572f
C4963 CSoutput.n62 gnd 0.146472f
C4964 CSoutput.n63 gnd 0.034102f
C4965 CSoutput.t202 gnd 0.320809f
C4966 CSoutput.n64 gnd 0.143283f
C4967 CSoutput.n65 gnd 0.040166f
C4968 CSoutput.n66 gnd 0.048499f
C4969 CSoutput.n67 gnd 0.048499f
C4970 CSoutput.n68 gnd 0.048499f
C4971 CSoutput.n69 gnd 0.039019f
C4972 CSoutput.n70 gnd 0.143283f
C4973 CSoutput.n71 gnd 0.040478f
C4974 CSoutput.n72 gnd 0.035402f
C4975 CSoutput.n73 gnd 0.048499f
C4976 CSoutput.n74 gnd 0.048499f
C4977 CSoutput.n75 gnd 0.036715f
C4978 CSoutput.n76 gnd 0.021805f
C4979 CSoutput.t190 gnd 0.360452f
C4980 CSoutput.n77 gnd 0.179058f
C4981 CSoutput.n78 gnd 0.766173f
C4982 CSoutput.t25 gnd 0.060495f
C4983 CSoutput.t81 gnd 0.060495f
C4984 CSoutput.n79 gnd 0.468376f
C4985 CSoutput.t90 gnd 0.060495f
C4986 CSoutput.t50 gnd 0.060495f
C4987 CSoutput.n80 gnd 0.467541f
C4988 CSoutput.n81 gnd 0.474553f
C4989 CSoutput.t168 gnd 0.060495f
C4990 CSoutput.t5 gnd 0.060495f
C4991 CSoutput.n82 gnd 0.467541f
C4992 CSoutput.n83 gnd 0.23384f
C4993 CSoutput.t18 gnd 0.060495f
C4994 CSoutput.t164 gnd 0.060495f
C4995 CSoutput.n84 gnd 0.467541f
C4996 CSoutput.n85 gnd 0.23384f
C4997 CSoutput.t174 gnd 0.060495f
C4998 CSoutput.t7 gnd 0.060495f
C4999 CSoutput.n86 gnd 0.467541f
C5000 CSoutput.n87 gnd 0.23384f
C5001 CSoutput.t59 gnd 0.060495f
C5002 CSoutput.t13 gnd 0.060495f
C5003 CSoutput.n88 gnd 0.467541f
C5004 CSoutput.n89 gnd 0.23384f
C5005 CSoutput.t6 gnd 0.060495f
C5006 CSoutput.t34 gnd 0.060495f
C5007 CSoutput.n90 gnd 0.467541f
C5008 CSoutput.n91 gnd 0.23384f
C5009 CSoutput.t95 gnd 0.060495f
C5010 CSoutput.t27 gnd 0.060495f
C5011 CSoutput.n92 gnd 0.467541f
C5012 CSoutput.n93 gnd 0.23384f
C5013 CSoutput.t69 gnd 0.060495f
C5014 CSoutput.t41 gnd 0.060495f
C5015 CSoutput.n94 gnd 0.467541f
C5016 CSoutput.n95 gnd 0.23384f
C5017 CSoutput.t37 gnd 0.060495f
C5018 CSoutput.t22 gnd 0.060495f
C5019 CSoutput.n96 gnd 0.467541f
C5020 CSoutput.n97 gnd 0.428808f
C5021 CSoutput.t182 gnd 0.060495f
C5022 CSoutput.t56 gnd 0.060495f
C5023 CSoutput.n98 gnd 0.468376f
C5024 CSoutput.t72 gnd 0.060495f
C5025 CSoutput.t178 gnd 0.060495f
C5026 CSoutput.n99 gnd 0.467541f
C5027 CSoutput.n100 gnd 0.474553f
C5028 CSoutput.t71 gnd 0.060495f
C5029 CSoutput.t170 gnd 0.060495f
C5030 CSoutput.n101 gnd 0.467541f
C5031 CSoutput.n102 gnd 0.23384f
C5032 CSoutput.t9 gnd 0.060495f
C5033 CSoutput.t74 gnd 0.060495f
C5034 CSoutput.n103 gnd 0.467541f
C5035 CSoutput.n104 gnd 0.23384f
C5036 CSoutput.t83 gnd 0.060495f
C5037 CSoutput.t93 gnd 0.060495f
C5038 CSoutput.n105 gnd 0.467541f
C5039 CSoutput.n106 gnd 0.23384f
C5040 CSoutput.t87 gnd 0.060495f
C5041 CSoutput.t62 gnd 0.060495f
C5042 CSoutput.n107 gnd 0.467541f
C5043 CSoutput.n108 gnd 0.23384f
C5044 CSoutput.t166 gnd 0.060495f
C5045 CSoutput.t77 gnd 0.060495f
C5046 CSoutput.n109 gnd 0.467541f
C5047 CSoutput.n110 gnd 0.23384f
C5048 CSoutput.t92 gnd 0.060495f
C5049 CSoutput.t26 gnd 0.060495f
C5050 CSoutput.n111 gnd 0.467541f
C5051 CSoutput.n112 gnd 0.23384f
C5052 CSoutput.t163 gnd 0.060495f
C5053 CSoutput.t70 gnd 0.060495f
C5054 CSoutput.n113 gnd 0.467541f
C5055 CSoutput.n114 gnd 0.23384f
C5056 CSoutput.t15 gnd 0.060495f
C5057 CSoutput.t31 gnd 0.060495f
C5058 CSoutput.n115 gnd 0.467541f
C5059 CSoutput.n116 gnd 0.348714f
C5060 CSoutput.n117 gnd 0.439726f
C5061 CSoutput.t55 gnd 0.060495f
C5062 CSoutput.t1 gnd 0.060495f
C5063 CSoutput.n118 gnd 0.468376f
C5064 CSoutput.t78 gnd 0.060495f
C5065 CSoutput.t38 gnd 0.060495f
C5066 CSoutput.n119 gnd 0.467541f
C5067 CSoutput.n120 gnd 0.474553f
C5068 CSoutput.t91 gnd 0.060495f
C5069 CSoutput.t175 gnd 0.060495f
C5070 CSoutput.n121 gnd 0.467541f
C5071 CSoutput.n122 gnd 0.23384f
C5072 CSoutput.t47 gnd 0.060495f
C5073 CSoutput.t30 gnd 0.060495f
C5074 CSoutput.n123 gnd 0.467541f
C5075 CSoutput.n124 gnd 0.23384f
C5076 CSoutput.t169 gnd 0.060495f
C5077 CSoutput.t4 gnd 0.060495f
C5078 CSoutput.n125 gnd 0.467541f
C5079 CSoutput.n126 gnd 0.23384f
C5080 CSoutput.t24 gnd 0.060495f
C5081 CSoutput.t48 gnd 0.060495f
C5082 CSoutput.n127 gnd 0.467541f
C5083 CSoutput.n128 gnd 0.23384f
C5084 CSoutput.t68 gnd 0.060495f
C5085 CSoutput.t19 gnd 0.060495f
C5086 CSoutput.n129 gnd 0.467541f
C5087 CSoutput.n130 gnd 0.23384f
C5088 CSoutput.t171 gnd 0.060495f
C5089 CSoutput.t12 gnd 0.060495f
C5090 CSoutput.n131 gnd 0.467541f
C5091 CSoutput.n132 gnd 0.23384f
C5092 CSoutput.t36 gnd 0.060495f
C5093 CSoutput.t97 gnd 0.060495f
C5094 CSoutput.n133 gnd 0.467541f
C5095 CSoutput.n134 gnd 0.23384f
C5096 CSoutput.t162 gnd 0.060495f
C5097 CSoutput.t177 gnd 0.060495f
C5098 CSoutput.n135 gnd 0.467541f
C5099 CSoutput.n136 gnd 0.348714f
C5100 CSoutput.n137 gnd 0.491501f
C5101 CSoutput.n138 gnd 9.09265f
C5102 CSoutput.n140 gnd 0.857935f
C5103 CSoutput.n141 gnd 0.643451f
C5104 CSoutput.n142 gnd 0.857935f
C5105 CSoutput.n143 gnd 0.857935f
C5106 CSoutput.n144 gnd 2.30983f
C5107 CSoutput.n145 gnd 0.857935f
C5108 CSoutput.n146 gnd 0.857935f
C5109 CSoutput.t193 gnd 1.07242f
C5110 CSoutput.n147 gnd 0.857935f
C5111 CSoutput.n148 gnd 0.857935f
C5112 CSoutput.n152 gnd 0.857935f
C5113 CSoutput.n156 gnd 0.857935f
C5114 CSoutput.n157 gnd 0.857935f
C5115 CSoutput.n159 gnd 0.857935f
C5116 CSoutput.n164 gnd 0.857935f
C5117 CSoutput.n166 gnd 0.857935f
C5118 CSoutput.n167 gnd 0.857935f
C5119 CSoutput.n169 gnd 0.857935f
C5120 CSoutput.n170 gnd 0.857935f
C5121 CSoutput.n172 gnd 0.857935f
C5122 CSoutput.t186 gnd 14.336f
C5123 CSoutput.n174 gnd 0.857935f
C5124 CSoutput.n175 gnd 0.643451f
C5125 CSoutput.n176 gnd 0.857935f
C5126 CSoutput.n177 gnd 0.857935f
C5127 CSoutput.n178 gnd 2.30983f
C5128 CSoutput.n179 gnd 0.857935f
C5129 CSoutput.n180 gnd 0.857935f
C5130 CSoutput.t203 gnd 1.07242f
C5131 CSoutput.n181 gnd 0.857935f
C5132 CSoutput.n182 gnd 0.857935f
C5133 CSoutput.n186 gnd 0.857935f
C5134 CSoutput.n190 gnd 0.857935f
C5135 CSoutput.n191 gnd 0.857935f
C5136 CSoutput.n193 gnd 0.857935f
C5137 CSoutput.n198 gnd 0.857935f
C5138 CSoutput.n200 gnd 0.857935f
C5139 CSoutput.n201 gnd 0.857935f
C5140 CSoutput.n203 gnd 0.857935f
C5141 CSoutput.n204 gnd 0.857935f
C5142 CSoutput.n206 gnd 0.857935f
C5143 CSoutput.n207 gnd 0.643451f
C5144 CSoutput.n209 gnd 0.857935f
C5145 CSoutput.n210 gnd 0.643451f
C5146 CSoutput.n211 gnd 0.857935f
C5147 CSoutput.n212 gnd 0.857935f
C5148 CSoutput.n213 gnd 2.30983f
C5149 CSoutput.n214 gnd 0.857935f
C5150 CSoutput.n215 gnd 0.857935f
C5151 CSoutput.t184 gnd 1.07242f
C5152 CSoutput.n216 gnd 0.857935f
C5153 CSoutput.n217 gnd 2.30983f
C5154 CSoutput.n219 gnd 0.857935f
C5155 CSoutput.n220 gnd 0.857935f
C5156 CSoutput.n222 gnd 0.857935f
C5157 CSoutput.n223 gnd 0.857935f
C5158 CSoutput.t194 gnd 14.102401f
C5159 CSoutput.t191 gnd 14.336f
C5160 CSoutput.n229 gnd 2.69147f
C5161 CSoutput.n230 gnd 10.9641f
C5162 CSoutput.n231 gnd 11.4228f
C5163 CSoutput.n236 gnd 2.91559f
C5164 CSoutput.n242 gnd 0.857935f
C5165 CSoutput.n244 gnd 0.857935f
C5166 CSoutput.n246 gnd 0.857935f
C5167 CSoutput.n248 gnd 0.857935f
C5168 CSoutput.n250 gnd 0.857935f
C5169 CSoutput.n256 gnd 0.857935f
C5170 CSoutput.n263 gnd 1.57398f
C5171 CSoutput.n264 gnd 1.57398f
C5172 CSoutput.n265 gnd 0.857935f
C5173 CSoutput.n266 gnd 0.857935f
C5174 CSoutput.n268 gnd 0.643451f
C5175 CSoutput.n269 gnd 0.551058f
C5176 CSoutput.n271 gnd 0.643451f
C5177 CSoutput.n272 gnd 0.551058f
C5178 CSoutput.n273 gnd 0.643451f
C5179 CSoutput.n275 gnd 0.857935f
C5180 CSoutput.n277 gnd 2.30983f
C5181 CSoutput.n278 gnd 2.69147f
C5182 CSoutput.n279 gnd 10.0841f
C5183 CSoutput.n281 gnd 0.643451f
C5184 CSoutput.n282 gnd 1.65564f
C5185 CSoutput.n283 gnd 0.643451f
C5186 CSoutput.n285 gnd 0.857935f
C5187 CSoutput.n287 gnd 2.30983f
C5188 CSoutput.n288 gnd 5.03117f
C5189 CSoutput.t180 gnd 0.060495f
C5190 CSoutput.t33 gnd 0.060495f
C5191 CSoutput.n289 gnd 0.468376f
C5192 CSoutput.t45 gnd 0.060495f
C5193 CSoutput.t23 gnd 0.060495f
C5194 CSoutput.n290 gnd 0.467541f
C5195 CSoutput.n291 gnd 0.474553f
C5196 CSoutput.t89 gnd 0.060495f
C5197 CSoutput.t51 gnd 0.060495f
C5198 CSoutput.n292 gnd 0.467541f
C5199 CSoutput.n293 gnd 0.23384f
C5200 CSoutput.t40 gnd 0.060495f
C5201 CSoutput.t75 gnd 0.060495f
C5202 CSoutput.n294 gnd 0.467541f
C5203 CSoutput.n295 gnd 0.23384f
C5204 CSoutput.t35 gnd 0.060495f
C5205 CSoutput.t173 gnd 0.060495f
C5206 CSoutput.n296 gnd 0.467541f
C5207 CSoutput.n297 gnd 0.23384f
C5208 CSoutput.t76 gnd 0.060495f
C5209 CSoutput.t172 gnd 0.060495f
C5210 CSoutput.n298 gnd 0.467541f
C5211 CSoutput.n299 gnd 0.23384f
C5212 CSoutput.t82 gnd 0.060495f
C5213 CSoutput.t61 gnd 0.060495f
C5214 CSoutput.n300 gnd 0.467541f
C5215 CSoutput.n301 gnd 0.23384f
C5216 CSoutput.t20 gnd 0.060495f
C5217 CSoutput.t49 gnd 0.060495f
C5218 CSoutput.n302 gnd 0.467541f
C5219 CSoutput.n303 gnd 0.23384f
C5220 CSoutput.t79 gnd 0.060495f
C5221 CSoutput.t8 gnd 0.060495f
C5222 CSoutput.n304 gnd 0.467541f
C5223 CSoutput.n305 gnd 0.23384f
C5224 CSoutput.t17 gnd 0.060495f
C5225 CSoutput.t80 gnd 0.060495f
C5226 CSoutput.n306 gnd 0.467541f
C5227 CSoutput.n307 gnd 0.428808f
C5228 CSoutput.t64 gnd 0.060495f
C5229 CSoutput.t53 gnd 0.060495f
C5230 CSoutput.n308 gnd 0.468376f
C5231 CSoutput.t165 gnd 0.060495f
C5232 CSoutput.t54 gnd 0.060495f
C5233 CSoutput.n309 gnd 0.467541f
C5234 CSoutput.n310 gnd 0.474553f
C5235 CSoutput.t88 gnd 0.060495f
C5236 CSoutput.t42 gnd 0.060495f
C5237 CSoutput.n311 gnd 0.467541f
C5238 CSoutput.n312 gnd 0.23384f
C5239 CSoutput.t0 gnd 0.060495f
C5240 CSoutput.t176 gnd 0.060495f
C5241 CSoutput.n313 gnd 0.467541f
C5242 CSoutput.n314 gnd 0.23384f
C5243 CSoutput.t66 gnd 0.060495f
C5244 CSoutput.t16 gnd 0.060495f
C5245 CSoutput.n315 gnd 0.467541f
C5246 CSoutput.n316 gnd 0.23384f
C5247 CSoutput.t167 gnd 0.060495f
C5248 CSoutput.t2 gnd 0.060495f
C5249 CSoutput.n317 gnd 0.467541f
C5250 CSoutput.n318 gnd 0.23384f
C5251 CSoutput.t183 gnd 0.060495f
C5252 CSoutput.t179 gnd 0.060495f
C5253 CSoutput.n319 gnd 0.467541f
C5254 CSoutput.n320 gnd 0.23384f
C5255 CSoutput.t46 gnd 0.060495f
C5256 CSoutput.t181 gnd 0.060495f
C5257 CSoutput.n321 gnd 0.467541f
C5258 CSoutput.n322 gnd 0.23384f
C5259 CSoutput.t85 gnd 0.060495f
C5260 CSoutput.t21 gnd 0.060495f
C5261 CSoutput.n323 gnd 0.467541f
C5262 CSoutput.n324 gnd 0.23384f
C5263 CSoutput.t63 gnd 0.060495f
C5264 CSoutput.t3 gnd 0.060495f
C5265 CSoutput.n325 gnd 0.467541f
C5266 CSoutput.n326 gnd 0.348714f
C5267 CSoutput.n327 gnd 0.439726f
C5268 CSoutput.t44 gnd 0.060495f
C5269 CSoutput.t94 gnd 0.060495f
C5270 CSoutput.n328 gnd 0.468376f
C5271 CSoutput.t10 gnd 0.060495f
C5272 CSoutput.t11 gnd 0.060495f
C5273 CSoutput.n329 gnd 0.467541f
C5274 CSoutput.n330 gnd 0.474553f
C5275 CSoutput.t39 gnd 0.060495f
C5276 CSoutput.t65 gnd 0.060495f
C5277 CSoutput.n331 gnd 0.467541f
C5278 CSoutput.n332 gnd 0.23384f
C5279 CSoutput.t57 gnd 0.060495f
C5280 CSoutput.t29 gnd 0.060495f
C5281 CSoutput.n333 gnd 0.467541f
C5282 CSoutput.n334 gnd 0.23384f
C5283 CSoutput.t32 gnd 0.060495f
C5284 CSoutput.t43 gnd 0.060495f
C5285 CSoutput.n335 gnd 0.467541f
C5286 CSoutput.n336 gnd 0.23384f
C5287 CSoutput.t86 gnd 0.060495f
C5288 CSoutput.t52 gnd 0.060495f
C5289 CSoutput.n337 gnd 0.467541f
C5290 CSoutput.n338 gnd 0.23384f
C5291 CSoutput.t67 gnd 0.060495f
C5292 CSoutput.t60 gnd 0.060495f
C5293 CSoutput.n339 gnd 0.467541f
C5294 CSoutput.n340 gnd 0.23384f
C5295 CSoutput.t28 gnd 0.060495f
C5296 CSoutput.t58 gnd 0.060495f
C5297 CSoutput.n341 gnd 0.467541f
C5298 CSoutput.n342 gnd 0.23384f
C5299 CSoutput.t73 gnd 0.060495f
C5300 CSoutput.t96 gnd 0.060495f
C5301 CSoutput.n343 gnd 0.467541f
C5302 CSoutput.n344 gnd 0.23384f
C5303 CSoutput.t84 gnd 0.060495f
C5304 CSoutput.t14 gnd 0.060495f
C5305 CSoutput.n345 gnd 0.467539f
C5306 CSoutput.n346 gnd 0.348715f
C5307 CSoutput.n347 gnd 0.491501f
C5308 CSoutput.n348 gnd 12.990201f
C5309 CSoutput.t151 gnd 0.052933f
C5310 CSoutput.t129 gnd 0.052933f
C5311 CSoutput.n349 gnd 0.469304f
C5312 CSoutput.t108 gnd 0.052933f
C5313 CSoutput.t110 gnd 0.052933f
C5314 CSoutput.n350 gnd 0.467739f
C5315 CSoutput.n351 gnd 0.435845f
C5316 CSoutput.t135 gnd 0.052933f
C5317 CSoutput.t141 gnd 0.052933f
C5318 CSoutput.n352 gnd 0.467739f
C5319 CSoutput.n353 gnd 0.214851f
C5320 CSoutput.t100 gnd 0.052933f
C5321 CSoutput.t152 gnd 0.052933f
C5322 CSoutput.n354 gnd 0.467739f
C5323 CSoutput.n355 gnd 0.214851f
C5324 CSoutput.t125 gnd 0.052933f
C5325 CSoutput.t132 gnd 0.052933f
C5326 CSoutput.n356 gnd 0.467739f
C5327 CSoutput.n357 gnd 0.214851f
C5328 CSoutput.t127 gnd 0.052933f
C5329 CSoutput.t117 gnd 0.052933f
C5330 CSoutput.n358 gnd 0.467739f
C5331 CSoutput.n359 gnd 0.214851f
C5332 CSoutput.t147 gnd 0.052933f
C5333 CSoutput.t160 gnd 0.052933f
C5334 CSoutput.n360 gnd 0.467739f
C5335 CSoutput.n361 gnd 0.214851f
C5336 CSoutput.t105 gnd 0.052933f
C5337 CSoutput.t124 gnd 0.052933f
C5338 CSoutput.n362 gnd 0.467739f
C5339 CSoutput.n363 gnd 0.396229f
C5340 CSoutput.t118 gnd 0.052933f
C5341 CSoutput.t148 gnd 0.052933f
C5342 CSoutput.n364 gnd 0.469304f
C5343 CSoutput.t101 gnd 0.052933f
C5344 CSoutput.t112 gnd 0.052933f
C5345 CSoutput.n365 gnd 0.467739f
C5346 CSoutput.n366 gnd 0.435845f
C5347 CSoutput.t126 gnd 0.052933f
C5348 CSoutput.t133 gnd 0.052933f
C5349 CSoutput.n367 gnd 0.467739f
C5350 CSoutput.n368 gnd 0.214851f
C5351 CSoutput.t143 gnd 0.052933f
C5352 CSoutput.t119 gnd 0.052933f
C5353 CSoutput.n369 gnd 0.467739f
C5354 CSoutput.n370 gnd 0.214851f
C5355 CSoutput.t104 gnd 0.052933f
C5356 CSoutput.t123 gnd 0.052933f
C5357 CSoutput.n371 gnd 0.467739f
C5358 CSoutput.n372 gnd 0.214851f
C5359 CSoutput.t106 gnd 0.052933f
C5360 CSoutput.t109 gnd 0.052933f
C5361 CSoutput.n373 gnd 0.467739f
C5362 CSoutput.n374 gnd 0.214851f
C5363 CSoutput.t116 gnd 0.052933f
C5364 CSoutput.t146 gnd 0.052933f
C5365 CSoutput.n375 gnd 0.467739f
C5366 CSoutput.n376 gnd 0.214851f
C5367 CSoutput.t99 gnd 0.052933f
C5368 CSoutput.t103 gnd 0.052933f
C5369 CSoutput.n377 gnd 0.467739f
C5370 CSoutput.n378 gnd 0.32619f
C5371 CSoutput.n379 gnd 0.606086f
C5372 CSoutput.n380 gnd 13.4217f
C5373 CSoutput.t137 gnd 0.052933f
C5374 CSoutput.t158 gnd 0.052933f
C5375 CSoutput.n381 gnd 0.469304f
C5376 CSoutput.t115 gnd 0.052933f
C5377 CSoutput.t98 gnd 0.052933f
C5378 CSoutput.n382 gnd 0.467739f
C5379 CSoutput.n383 gnd 0.435845f
C5380 CSoutput.t102 gnd 0.052933f
C5381 CSoutput.t140 gnd 0.052933f
C5382 CSoutput.n384 gnd 0.467739f
C5383 CSoutput.n385 gnd 0.214851f
C5384 CSoutput.t159 gnd 0.052933f
C5385 CSoutput.t113 gnd 0.052933f
C5386 CSoutput.n386 gnd 0.467739f
C5387 CSoutput.n387 gnd 0.214851f
C5388 CSoutput.t138 gnd 0.052933f
C5389 CSoutput.t131 gnd 0.052933f
C5390 CSoutput.n388 gnd 0.467739f
C5391 CSoutput.n389 gnd 0.214851f
C5392 CSoutput.t136 gnd 0.052933f
C5393 CSoutput.t120 gnd 0.052933f
C5394 CSoutput.n390 gnd 0.467739f
C5395 CSoutput.n391 gnd 0.214851f
C5396 CSoutput.t114 gnd 0.052933f
C5397 CSoutput.t155 gnd 0.052933f
C5398 CSoutput.n392 gnd 0.467739f
C5399 CSoutput.n393 gnd 0.214851f
C5400 CSoutput.t130 gnd 0.052933f
C5401 CSoutput.t122 gnd 0.052933f
C5402 CSoutput.n394 gnd 0.467739f
C5403 CSoutput.n395 gnd 0.396229f
C5404 CSoutput.t156 gnd 0.052933f
C5405 CSoutput.t144 gnd 0.052933f
C5406 CSoutput.n396 gnd 0.469304f
C5407 CSoutput.t107 gnd 0.052933f
C5408 CSoutput.t142 gnd 0.052933f
C5409 CSoutput.n397 gnd 0.467739f
C5410 CSoutput.n398 gnd 0.435845f
C5411 CSoutput.t139 gnd 0.052933f
C5412 CSoutput.t157 gnd 0.052933f
C5413 CSoutput.n399 gnd 0.467739f
C5414 CSoutput.n400 gnd 0.214851f
C5415 CSoutput.t145 gnd 0.052933f
C5416 CSoutput.t153 gnd 0.052933f
C5417 CSoutput.n401 gnd 0.467739f
C5418 CSoutput.n402 gnd 0.214851f
C5419 CSoutput.t161 gnd 0.052933f
C5420 CSoutput.t121 gnd 0.052933f
C5421 CSoutput.n403 gnd 0.467739f
C5422 CSoutput.n404 gnd 0.214851f
C5423 CSoutput.t128 gnd 0.052933f
C5424 CSoutput.t111 gnd 0.052933f
C5425 CSoutput.n405 gnd 0.467739f
C5426 CSoutput.n406 gnd 0.214851f
C5427 CSoutput.t154 gnd 0.052933f
C5428 CSoutput.t134 gnd 0.052933f
C5429 CSoutput.n407 gnd 0.467739f
C5430 CSoutput.n408 gnd 0.214851f
C5431 CSoutput.t150 gnd 0.052933f
C5432 CSoutput.t149 gnd 0.052933f
C5433 CSoutput.n409 gnd 0.467739f
C5434 CSoutput.n410 gnd 0.32619f
C5435 CSoutput.n411 gnd 0.606086f
C5436 CSoutput.n412 gnd 7.79018f
C5437 CSoutput.n413 gnd 15.586099f
C5438 commonsourceibias.n0 gnd 0.010545f
C5439 commonsourceibias.t94 gnd 0.159685f
C5440 commonsourceibias.t109 gnd 0.147652f
C5441 commonsourceibias.n1 gnd 0.006423f
C5442 commonsourceibias.n2 gnd 0.007903f
C5443 commonsourceibias.t72 gnd 0.147652f
C5444 commonsourceibias.n3 gnd 0.008017f
C5445 commonsourceibias.n4 gnd 0.007903f
C5446 commonsourceibias.t70 gnd 0.147652f
C5447 commonsourceibias.n5 gnd 0.058913f
C5448 commonsourceibias.t102 gnd 0.147652f
C5449 commonsourceibias.n6 gnd 0.006393f
C5450 commonsourceibias.n7 gnd 0.007903f
C5451 commonsourceibias.t118 gnd 0.147652f
C5452 commonsourceibias.n8 gnd 0.00763f
C5453 commonsourceibias.n9 gnd 0.007903f
C5454 commonsourceibias.t66 gnd 0.147652f
C5455 commonsourceibias.n10 gnd 0.058913f
C5456 commonsourceibias.t93 gnd 0.147652f
C5457 commonsourceibias.n11 gnd 0.006383f
C5458 commonsourceibias.n12 gnd 0.010545f
C5459 commonsourceibias.t34 gnd 0.159685f
C5460 commonsourceibias.t52 gnd 0.147652f
C5461 commonsourceibias.n13 gnd 0.006423f
C5462 commonsourceibias.n14 gnd 0.007903f
C5463 commonsourceibias.t26 gnd 0.147652f
C5464 commonsourceibias.n15 gnd 0.008017f
C5465 commonsourceibias.n16 gnd 0.007903f
C5466 commonsourceibias.t32 gnd 0.147652f
C5467 commonsourceibias.n17 gnd 0.058913f
C5468 commonsourceibias.t46 gnd 0.147652f
C5469 commonsourceibias.n18 gnd 0.006393f
C5470 commonsourceibias.n19 gnd 0.007903f
C5471 commonsourceibias.t8 gnd 0.147652f
C5472 commonsourceibias.n20 gnd 0.00763f
C5473 commonsourceibias.n21 gnd 0.007903f
C5474 commonsourceibias.t4 gnd 0.147652f
C5475 commonsourceibias.n22 gnd 0.058913f
C5476 commonsourceibias.t28 gnd 0.147652f
C5477 commonsourceibias.n23 gnd 0.006383f
C5478 commonsourceibias.n24 gnd 0.007903f
C5479 commonsourceibias.t36 gnd 0.147652f
C5480 commonsourceibias.t48 gnd 0.147652f
C5481 commonsourceibias.n25 gnd 0.058913f
C5482 commonsourceibias.n26 gnd 0.007903f
C5483 commonsourceibias.t0 gnd 0.147652f
C5484 commonsourceibias.n27 gnd 0.058913f
C5485 commonsourceibias.n28 gnd 0.007903f
C5486 commonsourceibias.t6 gnd 0.147652f
C5487 commonsourceibias.n29 gnd 0.058913f
C5488 commonsourceibias.n30 gnd 0.007903f
C5489 commonsourceibias.t42 gnd 0.147652f
C5490 commonsourceibias.n31 gnd 0.008983f
C5491 commonsourceibias.n32 gnd 0.007903f
C5492 commonsourceibias.t10 gnd 0.147652f
C5493 commonsourceibias.n33 gnd 0.010623f
C5494 commonsourceibias.t38 gnd 0.164481f
C5495 commonsourceibias.t54 gnd 0.147652f
C5496 commonsourceibias.n34 gnd 0.065644f
C5497 commonsourceibias.n35 gnd 0.070328f
C5498 commonsourceibias.n36 gnd 0.033639f
C5499 commonsourceibias.n37 gnd 0.007903f
C5500 commonsourceibias.n38 gnd 0.006423f
C5501 commonsourceibias.n39 gnd 0.01089f
C5502 commonsourceibias.n40 gnd 0.058913f
C5503 commonsourceibias.n41 gnd 0.010937f
C5504 commonsourceibias.n42 gnd 0.007903f
C5505 commonsourceibias.n43 gnd 0.007903f
C5506 commonsourceibias.n44 gnd 0.007903f
C5507 commonsourceibias.n45 gnd 0.008017f
C5508 commonsourceibias.n46 gnd 0.058913f
C5509 commonsourceibias.n47 gnd 0.009741f
C5510 commonsourceibias.n48 gnd 0.010776f
C5511 commonsourceibias.n49 gnd 0.007903f
C5512 commonsourceibias.n50 gnd 0.007903f
C5513 commonsourceibias.n51 gnd 0.010705f
C5514 commonsourceibias.n52 gnd 0.006393f
C5515 commonsourceibias.n53 gnd 0.010838f
C5516 commonsourceibias.n54 gnd 0.007903f
C5517 commonsourceibias.n55 gnd 0.007903f
C5518 commonsourceibias.n56 gnd 0.010904f
C5519 commonsourceibias.n57 gnd 0.009403f
C5520 commonsourceibias.n58 gnd 0.00763f
C5521 commonsourceibias.n59 gnd 0.007903f
C5522 commonsourceibias.n60 gnd 0.007903f
C5523 commonsourceibias.n61 gnd 0.009667f
C5524 commonsourceibias.n62 gnd 0.01085f
C5525 commonsourceibias.n63 gnd 0.058913f
C5526 commonsourceibias.n64 gnd 0.010777f
C5527 commonsourceibias.n65 gnd 0.007903f
C5528 commonsourceibias.n66 gnd 0.007903f
C5529 commonsourceibias.n67 gnd 0.007903f
C5530 commonsourceibias.n68 gnd 0.010777f
C5531 commonsourceibias.n69 gnd 0.058913f
C5532 commonsourceibias.n70 gnd 0.01085f
C5533 commonsourceibias.n71 gnd 0.009667f
C5534 commonsourceibias.n72 gnd 0.007903f
C5535 commonsourceibias.n73 gnd 0.007903f
C5536 commonsourceibias.n74 gnd 0.007903f
C5537 commonsourceibias.n75 gnd 0.009403f
C5538 commonsourceibias.n76 gnd 0.010904f
C5539 commonsourceibias.n77 gnd 0.058913f
C5540 commonsourceibias.n78 gnd 0.010838f
C5541 commonsourceibias.n79 gnd 0.007903f
C5542 commonsourceibias.n80 gnd 0.007903f
C5543 commonsourceibias.n81 gnd 0.007903f
C5544 commonsourceibias.n82 gnd 0.010705f
C5545 commonsourceibias.n83 gnd 0.058913f
C5546 commonsourceibias.n84 gnd 0.010776f
C5547 commonsourceibias.n85 gnd 0.009741f
C5548 commonsourceibias.n86 gnd 0.007903f
C5549 commonsourceibias.n87 gnd 0.007903f
C5550 commonsourceibias.n88 gnd 0.007903f
C5551 commonsourceibias.n89 gnd 0.008983f
C5552 commonsourceibias.n90 gnd 0.010937f
C5553 commonsourceibias.n91 gnd 0.058913f
C5554 commonsourceibias.n92 gnd 0.01089f
C5555 commonsourceibias.n93 gnd 0.007903f
C5556 commonsourceibias.n94 gnd 0.007903f
C5557 commonsourceibias.n95 gnd 0.007903f
C5558 commonsourceibias.n96 gnd 0.010623f
C5559 commonsourceibias.n97 gnd 0.058913f
C5560 commonsourceibias.n98 gnd 0.010649f
C5561 commonsourceibias.n99 gnd 0.071041f
C5562 commonsourceibias.n100 gnd 0.079434f
C5563 commonsourceibias.t35 gnd 0.017054f
C5564 commonsourceibias.t53 gnd 0.017054f
C5565 commonsourceibias.n101 gnd 0.150693f
C5566 commonsourceibias.n102 gnd 0.130533f
C5567 commonsourceibias.t27 gnd 0.017054f
C5568 commonsourceibias.t33 gnd 0.017054f
C5569 commonsourceibias.n103 gnd 0.150693f
C5570 commonsourceibias.n104 gnd 0.069219f
C5571 commonsourceibias.t47 gnd 0.017054f
C5572 commonsourceibias.t9 gnd 0.017054f
C5573 commonsourceibias.n105 gnd 0.150693f
C5574 commonsourceibias.n106 gnd 0.069219f
C5575 commonsourceibias.t5 gnd 0.017054f
C5576 commonsourceibias.t29 gnd 0.017054f
C5577 commonsourceibias.n107 gnd 0.150693f
C5578 commonsourceibias.n108 gnd 0.057829f
C5579 commonsourceibias.t55 gnd 0.017054f
C5580 commonsourceibias.t39 gnd 0.017054f
C5581 commonsourceibias.n109 gnd 0.151197f
C5582 commonsourceibias.t43 gnd 0.017054f
C5583 commonsourceibias.t11 gnd 0.017054f
C5584 commonsourceibias.n110 gnd 0.150693f
C5585 commonsourceibias.n111 gnd 0.140418f
C5586 commonsourceibias.t1 gnd 0.017054f
C5587 commonsourceibias.t7 gnd 0.017054f
C5588 commonsourceibias.n112 gnd 0.150693f
C5589 commonsourceibias.n113 gnd 0.069219f
C5590 commonsourceibias.t37 gnd 0.017054f
C5591 commonsourceibias.t49 gnd 0.017054f
C5592 commonsourceibias.n114 gnd 0.150693f
C5593 commonsourceibias.n115 gnd 0.057829f
C5594 commonsourceibias.n116 gnd 0.070025f
C5595 commonsourceibias.n117 gnd 0.007903f
C5596 commonsourceibias.t88 gnd 0.147652f
C5597 commonsourceibias.t105 gnd 0.147652f
C5598 commonsourceibias.n118 gnd 0.058913f
C5599 commonsourceibias.n119 gnd 0.007903f
C5600 commonsourceibias.t86 gnd 0.147652f
C5601 commonsourceibias.n120 gnd 0.058913f
C5602 commonsourceibias.n121 gnd 0.007903f
C5603 commonsourceibias.t82 gnd 0.147652f
C5604 commonsourceibias.n122 gnd 0.058913f
C5605 commonsourceibias.n123 gnd 0.007903f
C5606 commonsourceibias.t97 gnd 0.147652f
C5607 commonsourceibias.n124 gnd 0.008983f
C5608 commonsourceibias.n125 gnd 0.007903f
C5609 commonsourceibias.t111 gnd 0.147652f
C5610 commonsourceibias.n126 gnd 0.010623f
C5611 commonsourceibias.t89 gnd 0.164481f
C5612 commonsourceibias.t75 gnd 0.147652f
C5613 commonsourceibias.n127 gnd 0.065644f
C5614 commonsourceibias.n128 gnd 0.070328f
C5615 commonsourceibias.n129 gnd 0.033639f
C5616 commonsourceibias.n130 gnd 0.007903f
C5617 commonsourceibias.n131 gnd 0.006423f
C5618 commonsourceibias.n132 gnd 0.01089f
C5619 commonsourceibias.n133 gnd 0.058913f
C5620 commonsourceibias.n134 gnd 0.010937f
C5621 commonsourceibias.n135 gnd 0.007903f
C5622 commonsourceibias.n136 gnd 0.007903f
C5623 commonsourceibias.n137 gnd 0.007903f
C5624 commonsourceibias.n138 gnd 0.008017f
C5625 commonsourceibias.n139 gnd 0.058913f
C5626 commonsourceibias.n140 gnd 0.009741f
C5627 commonsourceibias.n141 gnd 0.010776f
C5628 commonsourceibias.n142 gnd 0.007903f
C5629 commonsourceibias.n143 gnd 0.007903f
C5630 commonsourceibias.n144 gnd 0.010705f
C5631 commonsourceibias.n145 gnd 0.006393f
C5632 commonsourceibias.n146 gnd 0.010838f
C5633 commonsourceibias.n147 gnd 0.007903f
C5634 commonsourceibias.n148 gnd 0.007903f
C5635 commonsourceibias.n149 gnd 0.010904f
C5636 commonsourceibias.n150 gnd 0.009403f
C5637 commonsourceibias.n151 gnd 0.00763f
C5638 commonsourceibias.n152 gnd 0.007903f
C5639 commonsourceibias.n153 gnd 0.007903f
C5640 commonsourceibias.n154 gnd 0.009667f
C5641 commonsourceibias.n155 gnd 0.01085f
C5642 commonsourceibias.n156 gnd 0.058913f
C5643 commonsourceibias.n157 gnd 0.010777f
C5644 commonsourceibias.n158 gnd 0.007865f
C5645 commonsourceibias.n159 gnd 0.057129f
C5646 commonsourceibias.n160 gnd 0.007865f
C5647 commonsourceibias.n161 gnd 0.010777f
C5648 commonsourceibias.n162 gnd 0.058913f
C5649 commonsourceibias.n163 gnd 0.01085f
C5650 commonsourceibias.n164 gnd 0.009667f
C5651 commonsourceibias.n165 gnd 0.007903f
C5652 commonsourceibias.n166 gnd 0.007903f
C5653 commonsourceibias.n167 gnd 0.007903f
C5654 commonsourceibias.n168 gnd 0.009403f
C5655 commonsourceibias.n169 gnd 0.010904f
C5656 commonsourceibias.n170 gnd 0.058913f
C5657 commonsourceibias.n171 gnd 0.010838f
C5658 commonsourceibias.n172 gnd 0.007903f
C5659 commonsourceibias.n173 gnd 0.007903f
C5660 commonsourceibias.n174 gnd 0.007903f
C5661 commonsourceibias.n175 gnd 0.010705f
C5662 commonsourceibias.n176 gnd 0.058913f
C5663 commonsourceibias.n177 gnd 0.010776f
C5664 commonsourceibias.n178 gnd 0.009741f
C5665 commonsourceibias.n179 gnd 0.007903f
C5666 commonsourceibias.n180 gnd 0.007903f
C5667 commonsourceibias.n181 gnd 0.007903f
C5668 commonsourceibias.n182 gnd 0.008983f
C5669 commonsourceibias.n183 gnd 0.010937f
C5670 commonsourceibias.n184 gnd 0.058913f
C5671 commonsourceibias.n185 gnd 0.01089f
C5672 commonsourceibias.n186 gnd 0.007903f
C5673 commonsourceibias.n187 gnd 0.007903f
C5674 commonsourceibias.n188 gnd 0.007903f
C5675 commonsourceibias.n189 gnd 0.010623f
C5676 commonsourceibias.n190 gnd 0.058913f
C5677 commonsourceibias.n191 gnd 0.010649f
C5678 commonsourceibias.n192 gnd 0.071041f
C5679 commonsourceibias.n193 gnd 0.046914f
C5680 commonsourceibias.n194 gnd 0.010545f
C5681 commonsourceibias.t96 gnd 0.147652f
C5682 commonsourceibias.n195 gnd 0.006423f
C5683 commonsourceibias.n196 gnd 0.007903f
C5684 commonsourceibias.t65 gnd 0.147652f
C5685 commonsourceibias.n197 gnd 0.008017f
C5686 commonsourceibias.n198 gnd 0.007903f
C5687 commonsourceibias.t127 gnd 0.147652f
C5688 commonsourceibias.n199 gnd 0.058913f
C5689 commonsourceibias.t87 gnd 0.147652f
C5690 commonsourceibias.n200 gnd 0.006393f
C5691 commonsourceibias.n201 gnd 0.007903f
C5692 commonsourceibias.t104 gnd 0.147652f
C5693 commonsourceibias.n202 gnd 0.00763f
C5694 commonsourceibias.n203 gnd 0.007903f
C5695 commonsourceibias.t122 gnd 0.147652f
C5696 commonsourceibias.n204 gnd 0.058913f
C5697 commonsourceibias.t80 gnd 0.147652f
C5698 commonsourceibias.n205 gnd 0.006383f
C5699 commonsourceibias.n206 gnd 0.007903f
C5700 commonsourceibias.t76 gnd 0.147652f
C5701 commonsourceibias.t90 gnd 0.147652f
C5702 commonsourceibias.n207 gnd 0.058913f
C5703 commonsourceibias.n208 gnd 0.007903f
C5704 commonsourceibias.t74 gnd 0.147652f
C5705 commonsourceibias.n209 gnd 0.058913f
C5706 commonsourceibias.n210 gnd 0.007903f
C5707 commonsourceibias.t71 gnd 0.147652f
C5708 commonsourceibias.n211 gnd 0.058913f
C5709 commonsourceibias.n212 gnd 0.007903f
C5710 commonsourceibias.t83 gnd 0.147652f
C5711 commonsourceibias.n213 gnd 0.008983f
C5712 commonsourceibias.n214 gnd 0.007903f
C5713 commonsourceibias.t98 gnd 0.147652f
C5714 commonsourceibias.n215 gnd 0.010623f
C5715 commonsourceibias.t77 gnd 0.164481f
C5716 commonsourceibias.t67 gnd 0.147652f
C5717 commonsourceibias.n216 gnd 0.065644f
C5718 commonsourceibias.n217 gnd 0.070328f
C5719 commonsourceibias.n218 gnd 0.033639f
C5720 commonsourceibias.n219 gnd 0.007903f
C5721 commonsourceibias.n220 gnd 0.006423f
C5722 commonsourceibias.n221 gnd 0.01089f
C5723 commonsourceibias.n222 gnd 0.058913f
C5724 commonsourceibias.n223 gnd 0.010937f
C5725 commonsourceibias.n224 gnd 0.007903f
C5726 commonsourceibias.n225 gnd 0.007903f
C5727 commonsourceibias.n226 gnd 0.007903f
C5728 commonsourceibias.n227 gnd 0.008017f
C5729 commonsourceibias.n228 gnd 0.058913f
C5730 commonsourceibias.n229 gnd 0.009741f
C5731 commonsourceibias.n230 gnd 0.010776f
C5732 commonsourceibias.n231 gnd 0.007903f
C5733 commonsourceibias.n232 gnd 0.007903f
C5734 commonsourceibias.n233 gnd 0.010705f
C5735 commonsourceibias.n234 gnd 0.006393f
C5736 commonsourceibias.n235 gnd 0.010838f
C5737 commonsourceibias.n236 gnd 0.007903f
C5738 commonsourceibias.n237 gnd 0.007903f
C5739 commonsourceibias.n238 gnd 0.010904f
C5740 commonsourceibias.n239 gnd 0.009403f
C5741 commonsourceibias.n240 gnd 0.00763f
C5742 commonsourceibias.n241 gnd 0.007903f
C5743 commonsourceibias.n242 gnd 0.007903f
C5744 commonsourceibias.n243 gnd 0.009667f
C5745 commonsourceibias.n244 gnd 0.01085f
C5746 commonsourceibias.n245 gnd 0.058913f
C5747 commonsourceibias.n246 gnd 0.010777f
C5748 commonsourceibias.n247 gnd 0.007903f
C5749 commonsourceibias.n248 gnd 0.007903f
C5750 commonsourceibias.n249 gnd 0.007903f
C5751 commonsourceibias.n250 gnd 0.010777f
C5752 commonsourceibias.n251 gnd 0.058913f
C5753 commonsourceibias.n252 gnd 0.01085f
C5754 commonsourceibias.n253 gnd 0.009667f
C5755 commonsourceibias.n254 gnd 0.007903f
C5756 commonsourceibias.n255 gnd 0.007903f
C5757 commonsourceibias.n256 gnd 0.007903f
C5758 commonsourceibias.n257 gnd 0.009403f
C5759 commonsourceibias.n258 gnd 0.010904f
C5760 commonsourceibias.n259 gnd 0.058913f
C5761 commonsourceibias.n260 gnd 0.010838f
C5762 commonsourceibias.n261 gnd 0.007903f
C5763 commonsourceibias.n262 gnd 0.007903f
C5764 commonsourceibias.n263 gnd 0.007903f
C5765 commonsourceibias.n264 gnd 0.010705f
C5766 commonsourceibias.n265 gnd 0.058913f
C5767 commonsourceibias.n266 gnd 0.010776f
C5768 commonsourceibias.n267 gnd 0.009741f
C5769 commonsourceibias.n268 gnd 0.007903f
C5770 commonsourceibias.n269 gnd 0.007903f
C5771 commonsourceibias.n270 gnd 0.007903f
C5772 commonsourceibias.n271 gnd 0.008983f
C5773 commonsourceibias.n272 gnd 0.010937f
C5774 commonsourceibias.n273 gnd 0.058913f
C5775 commonsourceibias.n274 gnd 0.01089f
C5776 commonsourceibias.n275 gnd 0.007903f
C5777 commonsourceibias.n276 gnd 0.007903f
C5778 commonsourceibias.n277 gnd 0.007903f
C5779 commonsourceibias.n278 gnd 0.010623f
C5780 commonsourceibias.n279 gnd 0.058913f
C5781 commonsourceibias.n280 gnd 0.010649f
C5782 commonsourceibias.t81 gnd 0.159685f
C5783 commonsourceibias.n281 gnd 0.071041f
C5784 commonsourceibias.n282 gnd 0.02535f
C5785 commonsourceibias.n283 gnd 0.398385f
C5786 commonsourceibias.n284 gnd 0.010545f
C5787 commonsourceibias.t113 gnd 0.159685f
C5788 commonsourceibias.t123 gnd 0.147652f
C5789 commonsourceibias.n285 gnd 0.006423f
C5790 commonsourceibias.n286 gnd 0.007903f
C5791 commonsourceibias.t68 gnd 0.147652f
C5792 commonsourceibias.n287 gnd 0.008017f
C5793 commonsourceibias.n288 gnd 0.007903f
C5794 commonsourceibias.t119 gnd 0.147652f
C5795 commonsourceibias.n289 gnd 0.006393f
C5796 commonsourceibias.n290 gnd 0.007903f
C5797 commonsourceibias.t64 gnd 0.147652f
C5798 commonsourceibias.n291 gnd 0.00763f
C5799 commonsourceibias.n292 gnd 0.007903f
C5800 commonsourceibias.t112 gnd 0.147652f
C5801 commonsourceibias.n293 gnd 0.006383f
C5802 commonsourceibias.n294 gnd 0.007903f
C5803 commonsourceibias.t107 gnd 0.147652f
C5804 commonsourceibias.t121 gnd 0.147652f
C5805 commonsourceibias.n295 gnd 0.058913f
C5806 commonsourceibias.n296 gnd 0.007903f
C5807 commonsourceibias.t78 gnd 0.147652f
C5808 commonsourceibias.n297 gnd 0.058913f
C5809 commonsourceibias.n298 gnd 0.007903f
C5810 commonsourceibias.t101 gnd 0.147652f
C5811 commonsourceibias.n299 gnd 0.058913f
C5812 commonsourceibias.n300 gnd 0.007903f
C5813 commonsourceibias.t115 gnd 0.147652f
C5814 commonsourceibias.n301 gnd 0.008983f
C5815 commonsourceibias.n302 gnd 0.007903f
C5816 commonsourceibias.t125 gnd 0.147652f
C5817 commonsourceibias.n303 gnd 0.010623f
C5818 commonsourceibias.t108 gnd 0.164481f
C5819 commonsourceibias.t91 gnd 0.147652f
C5820 commonsourceibias.n304 gnd 0.065644f
C5821 commonsourceibias.n305 gnd 0.070328f
C5822 commonsourceibias.n306 gnd 0.033639f
C5823 commonsourceibias.n307 gnd 0.007903f
C5824 commonsourceibias.n308 gnd 0.006423f
C5825 commonsourceibias.n309 gnd 0.01089f
C5826 commonsourceibias.n310 gnd 0.058913f
C5827 commonsourceibias.n311 gnd 0.010937f
C5828 commonsourceibias.n312 gnd 0.007903f
C5829 commonsourceibias.n313 gnd 0.007903f
C5830 commonsourceibias.n314 gnd 0.007903f
C5831 commonsourceibias.n315 gnd 0.008017f
C5832 commonsourceibias.n316 gnd 0.058913f
C5833 commonsourceibias.n317 gnd 0.009741f
C5834 commonsourceibias.n318 gnd 0.010776f
C5835 commonsourceibias.n319 gnd 0.007903f
C5836 commonsourceibias.n320 gnd 0.007903f
C5837 commonsourceibias.n321 gnd 0.010705f
C5838 commonsourceibias.n322 gnd 0.006393f
C5839 commonsourceibias.n323 gnd 0.010838f
C5840 commonsourceibias.n324 gnd 0.007903f
C5841 commonsourceibias.n325 gnd 0.007903f
C5842 commonsourceibias.n326 gnd 0.010904f
C5843 commonsourceibias.n327 gnd 0.009403f
C5844 commonsourceibias.n328 gnd 0.00763f
C5845 commonsourceibias.n329 gnd 0.007903f
C5846 commonsourceibias.n330 gnd 0.007903f
C5847 commonsourceibias.n331 gnd 0.009667f
C5848 commonsourceibias.n332 gnd 0.01085f
C5849 commonsourceibias.n333 gnd 0.058913f
C5850 commonsourceibias.n334 gnd 0.010777f
C5851 commonsourceibias.n335 gnd 0.007865f
C5852 commonsourceibias.t15 gnd 0.017054f
C5853 commonsourceibias.t61 gnd 0.017054f
C5854 commonsourceibias.n336 gnd 0.151197f
C5855 commonsourceibias.t23 gnd 0.017054f
C5856 commonsourceibias.t41 gnd 0.017054f
C5857 commonsourceibias.n337 gnd 0.150693f
C5858 commonsourceibias.n338 gnd 0.140418f
C5859 commonsourceibias.t63 gnd 0.017054f
C5860 commonsourceibias.t25 gnd 0.017054f
C5861 commonsourceibias.n339 gnd 0.150693f
C5862 commonsourceibias.n340 gnd 0.069219f
C5863 commonsourceibias.t45 gnd 0.017054f
C5864 commonsourceibias.t19 gnd 0.017054f
C5865 commonsourceibias.n341 gnd 0.150693f
C5866 commonsourceibias.n342 gnd 0.057829f
C5867 commonsourceibias.n343 gnd 0.010545f
C5868 commonsourceibias.t58 gnd 0.147652f
C5869 commonsourceibias.n344 gnd 0.006423f
C5870 commonsourceibias.n345 gnd 0.007903f
C5871 commonsourceibias.t12 gnd 0.147652f
C5872 commonsourceibias.n346 gnd 0.008017f
C5873 commonsourceibias.n347 gnd 0.007903f
C5874 commonsourceibias.t30 gnd 0.147652f
C5875 commonsourceibias.n348 gnd 0.006393f
C5876 commonsourceibias.n349 gnd 0.007903f
C5877 commonsourceibias.t20 gnd 0.147652f
C5878 commonsourceibias.n350 gnd 0.00763f
C5879 commonsourceibias.n351 gnd 0.007903f
C5880 commonsourceibias.t2 gnd 0.147652f
C5881 commonsourceibias.n352 gnd 0.006383f
C5882 commonsourceibias.n353 gnd 0.007903f
C5883 commonsourceibias.t18 gnd 0.147652f
C5884 commonsourceibias.t44 gnd 0.147652f
C5885 commonsourceibias.n354 gnd 0.058913f
C5886 commonsourceibias.n355 gnd 0.007903f
C5887 commonsourceibias.t24 gnd 0.147652f
C5888 commonsourceibias.n356 gnd 0.058913f
C5889 commonsourceibias.n357 gnd 0.007903f
C5890 commonsourceibias.t62 gnd 0.147652f
C5891 commonsourceibias.n358 gnd 0.058913f
C5892 commonsourceibias.n359 gnd 0.007903f
C5893 commonsourceibias.t40 gnd 0.147652f
C5894 commonsourceibias.n360 gnd 0.008983f
C5895 commonsourceibias.n361 gnd 0.007903f
C5896 commonsourceibias.t22 gnd 0.147652f
C5897 commonsourceibias.n362 gnd 0.010623f
C5898 commonsourceibias.t14 gnd 0.164481f
C5899 commonsourceibias.t60 gnd 0.147652f
C5900 commonsourceibias.n363 gnd 0.065644f
C5901 commonsourceibias.n364 gnd 0.070328f
C5902 commonsourceibias.n365 gnd 0.033639f
C5903 commonsourceibias.n366 gnd 0.007903f
C5904 commonsourceibias.n367 gnd 0.006423f
C5905 commonsourceibias.n368 gnd 0.01089f
C5906 commonsourceibias.n369 gnd 0.058913f
C5907 commonsourceibias.n370 gnd 0.010937f
C5908 commonsourceibias.n371 gnd 0.007903f
C5909 commonsourceibias.n372 gnd 0.007903f
C5910 commonsourceibias.n373 gnd 0.007903f
C5911 commonsourceibias.n374 gnd 0.008017f
C5912 commonsourceibias.n375 gnd 0.058913f
C5913 commonsourceibias.n376 gnd 0.009741f
C5914 commonsourceibias.n377 gnd 0.010776f
C5915 commonsourceibias.n378 gnd 0.007903f
C5916 commonsourceibias.n379 gnd 0.007903f
C5917 commonsourceibias.n380 gnd 0.010705f
C5918 commonsourceibias.n381 gnd 0.006393f
C5919 commonsourceibias.n382 gnd 0.010838f
C5920 commonsourceibias.n383 gnd 0.007903f
C5921 commonsourceibias.n384 gnd 0.007903f
C5922 commonsourceibias.n385 gnd 0.010904f
C5923 commonsourceibias.n386 gnd 0.009403f
C5924 commonsourceibias.n387 gnd 0.00763f
C5925 commonsourceibias.n388 gnd 0.007903f
C5926 commonsourceibias.n389 gnd 0.007903f
C5927 commonsourceibias.n390 gnd 0.009667f
C5928 commonsourceibias.n391 gnd 0.01085f
C5929 commonsourceibias.n392 gnd 0.058913f
C5930 commonsourceibias.n393 gnd 0.010777f
C5931 commonsourceibias.n394 gnd 0.007903f
C5932 commonsourceibias.n395 gnd 0.007903f
C5933 commonsourceibias.n396 gnd 0.007903f
C5934 commonsourceibias.n397 gnd 0.010777f
C5935 commonsourceibias.n398 gnd 0.058913f
C5936 commonsourceibias.n399 gnd 0.01085f
C5937 commonsourceibias.t50 gnd 0.147652f
C5938 commonsourceibias.n400 gnd 0.058913f
C5939 commonsourceibias.n401 gnd 0.009667f
C5940 commonsourceibias.n402 gnd 0.007903f
C5941 commonsourceibias.n403 gnd 0.007903f
C5942 commonsourceibias.n404 gnd 0.007903f
C5943 commonsourceibias.n405 gnd 0.009403f
C5944 commonsourceibias.n406 gnd 0.010904f
C5945 commonsourceibias.n407 gnd 0.058913f
C5946 commonsourceibias.n408 gnd 0.010838f
C5947 commonsourceibias.n409 gnd 0.007903f
C5948 commonsourceibias.n410 gnd 0.007903f
C5949 commonsourceibias.n411 gnd 0.007903f
C5950 commonsourceibias.n412 gnd 0.010705f
C5951 commonsourceibias.n413 gnd 0.058913f
C5952 commonsourceibias.n414 gnd 0.010776f
C5953 commonsourceibias.t56 gnd 0.147652f
C5954 commonsourceibias.n415 gnd 0.058913f
C5955 commonsourceibias.n416 gnd 0.009741f
C5956 commonsourceibias.n417 gnd 0.007903f
C5957 commonsourceibias.n418 gnd 0.007903f
C5958 commonsourceibias.n419 gnd 0.007903f
C5959 commonsourceibias.n420 gnd 0.008983f
C5960 commonsourceibias.n421 gnd 0.010937f
C5961 commonsourceibias.n422 gnd 0.058913f
C5962 commonsourceibias.n423 gnd 0.01089f
C5963 commonsourceibias.n424 gnd 0.007903f
C5964 commonsourceibias.n425 gnd 0.007903f
C5965 commonsourceibias.n426 gnd 0.007903f
C5966 commonsourceibias.n427 gnd 0.010623f
C5967 commonsourceibias.n428 gnd 0.058913f
C5968 commonsourceibias.n429 gnd 0.010649f
C5969 commonsourceibias.t16 gnd 0.159685f
C5970 commonsourceibias.n430 gnd 0.071041f
C5971 commonsourceibias.n431 gnd 0.079434f
C5972 commonsourceibias.t59 gnd 0.017054f
C5973 commonsourceibias.t17 gnd 0.017054f
C5974 commonsourceibias.n432 gnd 0.150693f
C5975 commonsourceibias.n433 gnd 0.130533f
C5976 commonsourceibias.t57 gnd 0.017054f
C5977 commonsourceibias.t13 gnd 0.017054f
C5978 commonsourceibias.n434 gnd 0.150693f
C5979 commonsourceibias.n435 gnd 0.069219f
C5980 commonsourceibias.t21 gnd 0.017054f
C5981 commonsourceibias.t31 gnd 0.017054f
C5982 commonsourceibias.n436 gnd 0.150693f
C5983 commonsourceibias.n437 gnd 0.069219f
C5984 commonsourceibias.t3 gnd 0.017054f
C5985 commonsourceibias.t51 gnd 0.017054f
C5986 commonsourceibias.n438 gnd 0.150693f
C5987 commonsourceibias.n439 gnd 0.057829f
C5988 commonsourceibias.n440 gnd 0.070025f
C5989 commonsourceibias.n441 gnd 0.057129f
C5990 commonsourceibias.n442 gnd 0.007865f
C5991 commonsourceibias.n443 gnd 0.010777f
C5992 commonsourceibias.n444 gnd 0.058913f
C5993 commonsourceibias.n445 gnd 0.01085f
C5994 commonsourceibias.t126 gnd 0.147652f
C5995 commonsourceibias.n446 gnd 0.058913f
C5996 commonsourceibias.n447 gnd 0.009667f
C5997 commonsourceibias.n448 gnd 0.007903f
C5998 commonsourceibias.n449 gnd 0.007903f
C5999 commonsourceibias.n450 gnd 0.007903f
C6000 commonsourceibias.n451 gnd 0.009403f
C6001 commonsourceibias.n452 gnd 0.010904f
C6002 commonsourceibias.n453 gnd 0.058913f
C6003 commonsourceibias.n454 gnd 0.010838f
C6004 commonsourceibias.n455 gnd 0.007903f
C6005 commonsourceibias.n456 gnd 0.007903f
C6006 commonsourceibias.n457 gnd 0.007903f
C6007 commonsourceibias.n458 gnd 0.010705f
C6008 commonsourceibias.n459 gnd 0.058913f
C6009 commonsourceibias.n460 gnd 0.010776f
C6010 commonsourceibias.t84 gnd 0.147652f
C6011 commonsourceibias.n461 gnd 0.058913f
C6012 commonsourceibias.n462 gnd 0.009741f
C6013 commonsourceibias.n463 gnd 0.007903f
C6014 commonsourceibias.n464 gnd 0.007903f
C6015 commonsourceibias.n465 gnd 0.007903f
C6016 commonsourceibias.n466 gnd 0.008983f
C6017 commonsourceibias.n467 gnd 0.010937f
C6018 commonsourceibias.n468 gnd 0.058913f
C6019 commonsourceibias.n469 gnd 0.01089f
C6020 commonsourceibias.n470 gnd 0.007903f
C6021 commonsourceibias.n471 gnd 0.007903f
C6022 commonsourceibias.n472 gnd 0.007903f
C6023 commonsourceibias.n473 gnd 0.010623f
C6024 commonsourceibias.n474 gnd 0.058913f
C6025 commonsourceibias.n475 gnd 0.010649f
C6026 commonsourceibias.n476 gnd 0.071041f
C6027 commonsourceibias.n477 gnd 0.046914f
C6028 commonsourceibias.n478 gnd 0.010545f
C6029 commonsourceibias.t114 gnd 0.147652f
C6030 commonsourceibias.n479 gnd 0.006423f
C6031 commonsourceibias.n480 gnd 0.007903f
C6032 commonsourceibias.t124 gnd 0.147652f
C6033 commonsourceibias.n481 gnd 0.008017f
C6034 commonsourceibias.n482 gnd 0.007903f
C6035 commonsourceibias.t106 gnd 0.147652f
C6036 commonsourceibias.n483 gnd 0.006393f
C6037 commonsourceibias.n484 gnd 0.007903f
C6038 commonsourceibias.t120 gnd 0.147652f
C6039 commonsourceibias.n485 gnd 0.00763f
C6040 commonsourceibias.n486 gnd 0.007903f
C6041 commonsourceibias.t99 gnd 0.147652f
C6042 commonsourceibias.n487 gnd 0.006383f
C6043 commonsourceibias.n488 gnd 0.007903f
C6044 commonsourceibias.t92 gnd 0.147652f
C6045 commonsourceibias.t110 gnd 0.147652f
C6046 commonsourceibias.n489 gnd 0.058913f
C6047 commonsourceibias.n490 gnd 0.007903f
C6048 commonsourceibias.t69 gnd 0.147652f
C6049 commonsourceibias.n491 gnd 0.058913f
C6050 commonsourceibias.n492 gnd 0.007903f
C6051 commonsourceibias.t85 gnd 0.147652f
C6052 commonsourceibias.n493 gnd 0.058913f
C6053 commonsourceibias.n494 gnd 0.007903f
C6054 commonsourceibias.t103 gnd 0.147652f
C6055 commonsourceibias.n495 gnd 0.008983f
C6056 commonsourceibias.n496 gnd 0.007903f
C6057 commonsourceibias.t116 gnd 0.147652f
C6058 commonsourceibias.n497 gnd 0.010623f
C6059 commonsourceibias.t95 gnd 0.164481f
C6060 commonsourceibias.t79 gnd 0.147652f
C6061 commonsourceibias.n498 gnd 0.065644f
C6062 commonsourceibias.n499 gnd 0.070328f
C6063 commonsourceibias.n500 gnd 0.033639f
C6064 commonsourceibias.n501 gnd 0.007903f
C6065 commonsourceibias.n502 gnd 0.006423f
C6066 commonsourceibias.n503 gnd 0.01089f
C6067 commonsourceibias.n504 gnd 0.058913f
C6068 commonsourceibias.n505 gnd 0.010937f
C6069 commonsourceibias.n506 gnd 0.007903f
C6070 commonsourceibias.n507 gnd 0.007903f
C6071 commonsourceibias.n508 gnd 0.007903f
C6072 commonsourceibias.n509 gnd 0.008017f
C6073 commonsourceibias.n510 gnd 0.058913f
C6074 commonsourceibias.n511 gnd 0.009741f
C6075 commonsourceibias.n512 gnd 0.010776f
C6076 commonsourceibias.n513 gnd 0.007903f
C6077 commonsourceibias.n514 gnd 0.007903f
C6078 commonsourceibias.n515 gnd 0.010705f
C6079 commonsourceibias.n516 gnd 0.006393f
C6080 commonsourceibias.n517 gnd 0.010838f
C6081 commonsourceibias.n518 gnd 0.007903f
C6082 commonsourceibias.n519 gnd 0.007903f
C6083 commonsourceibias.n520 gnd 0.010904f
C6084 commonsourceibias.n521 gnd 0.009403f
C6085 commonsourceibias.n522 gnd 0.00763f
C6086 commonsourceibias.n523 gnd 0.007903f
C6087 commonsourceibias.n524 gnd 0.007903f
C6088 commonsourceibias.n525 gnd 0.009667f
C6089 commonsourceibias.n526 gnd 0.01085f
C6090 commonsourceibias.n527 gnd 0.058913f
C6091 commonsourceibias.n528 gnd 0.010777f
C6092 commonsourceibias.n529 gnd 0.007903f
C6093 commonsourceibias.n530 gnd 0.007903f
C6094 commonsourceibias.n531 gnd 0.007903f
C6095 commonsourceibias.n532 gnd 0.010777f
C6096 commonsourceibias.n533 gnd 0.058913f
C6097 commonsourceibias.n534 gnd 0.01085f
C6098 commonsourceibias.t117 gnd 0.147652f
C6099 commonsourceibias.n535 gnd 0.058913f
C6100 commonsourceibias.n536 gnd 0.009667f
C6101 commonsourceibias.n537 gnd 0.007903f
C6102 commonsourceibias.n538 gnd 0.007903f
C6103 commonsourceibias.n539 gnd 0.007903f
C6104 commonsourceibias.n540 gnd 0.009403f
C6105 commonsourceibias.n541 gnd 0.010904f
C6106 commonsourceibias.n542 gnd 0.058913f
C6107 commonsourceibias.n543 gnd 0.010838f
C6108 commonsourceibias.n544 gnd 0.007903f
C6109 commonsourceibias.n545 gnd 0.007903f
C6110 commonsourceibias.n546 gnd 0.007903f
C6111 commonsourceibias.n547 gnd 0.010705f
C6112 commonsourceibias.n548 gnd 0.058913f
C6113 commonsourceibias.n549 gnd 0.010776f
C6114 commonsourceibias.t73 gnd 0.147652f
C6115 commonsourceibias.n550 gnd 0.058913f
C6116 commonsourceibias.n551 gnd 0.009741f
C6117 commonsourceibias.n552 gnd 0.007903f
C6118 commonsourceibias.n553 gnd 0.007903f
C6119 commonsourceibias.n554 gnd 0.007903f
C6120 commonsourceibias.n555 gnd 0.008983f
C6121 commonsourceibias.n556 gnd 0.010937f
C6122 commonsourceibias.n557 gnd 0.058913f
C6123 commonsourceibias.n558 gnd 0.01089f
C6124 commonsourceibias.n559 gnd 0.007903f
C6125 commonsourceibias.n560 gnd 0.007903f
C6126 commonsourceibias.n561 gnd 0.007903f
C6127 commonsourceibias.n562 gnd 0.010623f
C6128 commonsourceibias.n563 gnd 0.058913f
C6129 commonsourceibias.n564 gnd 0.010649f
C6130 commonsourceibias.t100 gnd 0.159685f
C6131 commonsourceibias.n565 gnd 0.071041f
C6132 commonsourceibias.n566 gnd 0.02535f
C6133 commonsourceibias.n567 gnd 0.218509f
C6134 commonsourceibias.n568 gnd 4.2686f
.ends

