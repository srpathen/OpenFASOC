* NGSPICE file created from opamp.ext - technology: sky130A

.subckt opamp output vdd plus minus commonsourceibias outputibias diffpairibias gnd CSoutput
Cload output gnd 0.0p
X0 gnd.t177 gnd.t174 gnd.t176 gnd.t175 sky130_fd_pr__nfet_01v8 ad=2.34 pd=12.78 as=0 ps=0 w=6 l=2
X1 commonsourceibias.t47 commonsourceibias.t46 gnd.t271 gnd.t212 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=2.73 ps=14.78 w=7 l=1
X2 gnd.t182 commonsourceibias.t48 CSoutput.t67 gnd.t38 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X3 gnd.t173 gnd.t171 gnd.t172 gnd.t159 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=0 ps=0 w=7 l=1
X4 vdd.t160 a_n5644_8799.t36 CSoutput.t1 vdd.t107 sky130_fd_pr__pfet_01v8_lvt ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X5 a_n1986_8322.t11 a_n2848_n452.t48 vdd.t187 vdd.t186 sky130_fd_pr__pfet_01v8_lvt ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X6 a_n1808_13878.t19 a_n2848_n452.t26 a_n2848_n452.t27 vdd.t4 sky130_fd_pr__pfet_01v8_lvt ad=1.485 pd=9.33 as=3.51 ps=18.78 w=9 l=0.5
X7 a_n5644_8799.t24 plus.t5 a_n3106_n452.t40 gnd.t242 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.9
X8 output.t19 outputibias.t8 gnd.t64 gnd.t63 sky130_fd_pr__nfet_01v8 ad=2.34 pd=12.78 as=2.34 ps=12.78 w=6 l=2
X9 gnd.t263 commonsourceibias.t49 CSoutput.t66 gnd.t51 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X10 a_n3106_n452.t39 plus.t6 a_n5644_8799.t2 gnd.t19 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.9
X11 vdd.t167 CSoutput.t96 output.t15 gnd.t221 sky130_fd_pr__nfet_01v8_lvt ad=0.825 pd=5.33 as=1.95 ps=10.78 w=5 l=1
X12 a_n2848_n452.t41 a_n2848_n452.t40 a_n1808_13878.t18 vdd.t11 sky130_fd_pr__pfet_01v8_lvt ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X13 a_n1808_13878.t17 a_n2848_n452.t28 a_n2848_n452.t29 vdd.t0 sky130_fd_pr__pfet_01v8_lvt ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X14 vdd.t96 vdd.t94 vdd.t95 vdd.t69 sky130_fd_pr__pfet_01v8_lvt ad=3.51 pd=18.78 as=0 ps=0 w=9 l=0.5
X15 a_n1808_13878.t7 a_n2848_n452.t49 vdd.t189 vdd.t188 sky130_fd_pr__pfet_01v8_lvt ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X16 gnd.t194 commonsourceibias.t44 commonsourceibias.t45 gnd.t193 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X17 vdd.t165 CSoutput.t97 output.t14 gnd.t222 sky130_fd_pr__nfet_01v8_lvt ad=0.825 pd=5.33 as=0.825 ps=5.33 w=5 l=1
X18 CSoutput.t90 a_n5644_8799.t37 vdd.t159 vdd.t103 sky130_fd_pr__pfet_01v8_lvt ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X19 gnd.t291 commonsourceibias.t50 CSoutput.t65 gnd.t193 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X20 outputibias.t7 outputibias.t6 gnd.t23 gnd.t22 sky130_fd_pr__nfet_01v8 ad=2.34 pd=12.78 as=2.34 ps=12.78 w=6 l=2
X21 vdd.t93 vdd.t91 vdd.t92 vdd.t44 sky130_fd_pr__pfet_01v8_lvt ad=3.12 pd=16.78 as=0 ps=0 w=8 l=0.5
X22 a_n1986_8322.t23 a_n2848_n452.t50 a_n5644_8799.t15 vdd.t177 sky130_fd_pr__pfet_01v8_lvt ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X23 a_n2848_n452.t8 minus.t5 a_n3106_n452.t8 gnd.t37 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.9
X24 a_n5644_8799.t22 plus.t7 a_n3106_n452.t38 gnd.t235 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.9
X25 gnd.t219 commonsourceibias.t42 commonsourceibias.t43 gnd.t218 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X26 plus.t4 gnd.t168 gnd.t170 gnd.t169 sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.5
X27 a_n2848_n452.t7 minus.t6 a_n3106_n452.t7 gnd.t36 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.9
X28 CSoutput.t64 commonsourceibias.t51 gnd.t284 gnd.t44 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X29 CSoutput.t98 a_n1986_8322.t0 sky130_fd_pr__cap_mim_m3_1 l=12 w=12
X30 gnd.t41 commonsourceibias.t40 commonsourceibias.t41 gnd.t40 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X31 CSoutput.t68 a_n5644_8799.t38 vdd.t158 vdd.t116 sky130_fd_pr__pfet_01v8_lvt ad=1.32 pd=8.33 as=3.12 ps=16.78 w=8 l=0.5
X32 vdd.t157 a_n5644_8799.t39 CSoutput.t10 vdd.t134 sky130_fd_pr__pfet_01v8_lvt ad=3.12 pd=16.78 as=1.32 ps=8.33 w=8 l=0.5
X33 a_n3106_n452.t37 plus.t8 a_n5644_8799.t13 gnd.t69 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.9
X34 a_n5644_8799.t16 a_n2848_n452.t51 a_n1986_8322.t22 vdd.t4 sky130_fd_pr__pfet_01v8_lvt ad=1.485 pd=9.33 as=3.51 ps=18.78 w=9 l=0.5
X35 CSoutput.t14 a_n5644_8799.t40 vdd.t156 vdd.t97 sky130_fd_pr__pfet_01v8_lvt ad=1.32 pd=8.33 as=3.12 ps=16.78 w=8 l=0.5
X36 vdd.t155 a_n5644_8799.t41 CSoutput.t0 vdd.t150 sky130_fd_pr__pfet_01v8_lvt ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X37 a_n3106_n452.t2 minus.t7 a_n2848_n452.t2 gnd.t5 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.9
X38 CSoutput.t63 commonsourceibias.t52 gnd.t286 gnd.t232 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X39 a_n3106_n452.t11 diffpairibias.t16 gnd.t59 gnd.t58 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=2.73 ps=14.78 w=7 l=1
X40 output.t13 CSoutput.t99 vdd.t175 gnd.t187 sky130_fd_pr__nfet_01v8_lvt ad=0.825 pd=5.33 as=0.825 ps=5.33 w=5 l=1
X41 vdd.t164 CSoutput.t100 output.t12 gnd.t188 sky130_fd_pr__nfet_01v8_lvt ad=0.825 pd=5.33 as=0.825 ps=5.33 w=5 l=1
X42 CSoutput.t62 commonsourceibias.t53 gnd.t289 gnd.t34 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X43 CSoutput.t94 a_n5644_8799.t42 vdd.t154 vdd.t112 sky130_fd_pr__pfet_01v8_lvt ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X44 vdd.t90 vdd.t88 vdd.t89 vdd.t22 sky130_fd_pr__pfet_01v8_lvt ad=3.12 pd=16.78 as=0 ps=0 w=8 l=0.5
X45 CSoutput.t61 commonsourceibias.t54 gnd.t257 gnd.t212 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=2.73 ps=14.78 w=7 l=1
X46 gnd.t167 gnd.t165 gnd.t166 gnd.t117 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=0 ps=0 w=7 l=0.9
X47 a_n3106_n452.t36 plus.t9 a_n5644_8799.t14 gnd.t28 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.9
X48 a_n1808_13878.t16 a_n2848_n452.t36 a_n2848_n452.t37 vdd.t7 sky130_fd_pr__pfet_01v8_lvt ad=1.485 pd=9.33 as=3.51 ps=18.78 w=9 l=0.5
X49 vdd.t153 a_n5644_8799.t43 CSoutput.t84 vdd.t150 sky130_fd_pr__pfet_01v8_lvt ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X50 a_n3106_n452.t35 plus.t10 a_n5644_8799.t0 gnd.t0 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.9
X51 a_n3106_n452.t4 minus.t8 a_n2848_n452.t4 gnd.t11 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=1.155 ps=7.33 w=7 l=0.9
X52 diffpairibias.t15 diffpairibias.t14 gnd.t241 gnd.t240 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=2.73 ps=14.78 w=7 l=1
X53 a_n2848_n452.t35 a_n2848_n452.t34 a_n1808_13878.t15 vdd.t10 sky130_fd_pr__pfet_01v8_lvt ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X54 CSoutput.t6 a_n5644_8799.t44 vdd.t152 vdd.t128 sky130_fd_pr__pfet_01v8_lvt ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X55 gnd.t164 gnd.t162 gnd.t163 gnd.t159 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=0 ps=0 w=7 l=1
X56 vdd.t87 vdd.t85 vdd.t86 vdd.t54 sky130_fd_pr__pfet_01v8_lvt ad=3.51 pd=18.78 as=0 ps=0 w=9 l=0.5
X57 gnd.t52 commonsourceibias.t55 CSoutput.t60 gnd.t51 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X58 gnd.t249 commonsourceibias.t56 CSoutput.t59 gnd.t207 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X59 diffpairibias.t13 diffpairibias.t12 gnd.t57 gnd.t56 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=2.73 ps=14.78 w=7 l=1
X60 vdd.t84 vdd.t82 vdd.t83 vdd.t33 sky130_fd_pr__pfet_01v8_lvt ad=3.12 pd=16.78 as=0 ps=0 w=8 l=0.5
X61 gnd.t50 commonsourceibias.t57 CSoutput.t58 gnd.t40 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X62 commonsourceibias.t39 commonsourceibias.t38 gnd.t272 gnd.t44 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X63 vdd.t151 a_n5644_8799.t45 CSoutput.t76 vdd.t150 sky130_fd_pr__pfet_01v8_lvt ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X64 vdd.t171 CSoutput.t101 output.t11 gnd.t189 sky130_fd_pr__nfet_01v8_lvt ad=0.825 pd=5.33 as=0.825 ps=5.33 w=5 l=1
X65 vdd.t149 a_n5644_8799.t46 CSoutput.t75 vdd.t125 sky130_fd_pr__pfet_01v8_lvt ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X66 CSoutput.t9 a_n5644_8799.t47 vdd.t148 vdd.t97 sky130_fd_pr__pfet_01v8_lvt ad=1.32 pd=8.33 as=3.12 ps=16.78 w=8 l=0.5
X67 a_n3106_n452.t1 minus.t9 a_n2848_n452.t1 gnd.t4 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.9
X68 a_n3106_n452.t34 plus.t11 a_n5644_8799.t18 gnd.t200 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=1.155 ps=7.33 w=7 l=0.9
X69 vdd.t147 a_n5644_8799.t48 CSoutput.t72 vdd.t101 sky130_fd_pr__pfet_01v8_lvt ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X70 gnd.t179 commonsourceibias.t58 CSoutput.t57 gnd.t178 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X71 a_n5644_8799.t29 plus.t12 a_n3106_n452.t33 gnd.t266 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.9
X72 commonsourceibias.t37 commonsourceibias.t36 gnd.t214 gnd.t30 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X73 CSoutput.t79 a_n5644_8799.t49 vdd.t146 vdd.t112 sky130_fd_pr__pfet_01v8_lvt ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X74 CSoutput.t74 a_n5644_8799.t50 vdd.t145 vdd.t138 sky130_fd_pr__pfet_01v8_lvt ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X75 a_n3106_n452.t16 diffpairibias.t17 gnd.t206 gnd.t205 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=2.73 ps=14.78 w=7 l=1
X76 gnd.t211 commonsourceibias.t34 commonsourceibias.t35 gnd.t178 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X77 CSoutput.t3 a_n5644_8799.t51 vdd.t144 vdd.t138 sky130_fd_pr__pfet_01v8_lvt ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X78 a_n3106_n452.t32 plus.t13 a_n5644_8799.t1 gnd.t14 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.9
X79 vdd.t143 a_n5644_8799.t52 CSoutput.t11 vdd.t136 sky130_fd_pr__pfet_01v8_lvt ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X80 gnd.t186 commonsourceibias.t32 commonsourceibias.t33 gnd.t53 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=1.155 ps=7.33 w=7 l=1
X81 commonsourceibias.t31 commonsourceibias.t30 gnd.t35 gnd.t34 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X82 a_n2848_n452.t21 a_n2848_n452.t20 a_n1808_13878.t14 vdd.t177 sky130_fd_pr__pfet_01v8_lvt ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X83 outputibias.t5 outputibias.t4 gnd.t25 gnd.t24 sky130_fd_pr__nfet_01v8 ad=2.34 pd=12.78 as=2.34 ps=12.78 w=6 l=2
X84 a_n2848_n452.t23 a_n2848_n452.t22 a_n1808_13878.t13 vdd.t181 sky130_fd_pr__pfet_01v8_lvt ad=3.51 pd=18.78 as=1.485 ps=9.33 w=9 l=0.5
X85 vdd.t142 a_n5644_8799.t53 CSoutput.t87 vdd.t134 sky130_fd_pr__pfet_01v8_lvt ad=3.12 pd=16.78 as=1.32 ps=8.33 w=8 l=0.5
X86 a_n5644_8799.t10 a_n2848_n452.t52 a_n1986_8322.t21 vdd.t14 sky130_fd_pr__pfet_01v8_lvt ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X87 CSoutput.t56 commonsourceibias.t59 gnd.t233 gnd.t232 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X88 vdd.t141 a_n5644_8799.t54 CSoutput.t77 vdd.t136 sky130_fd_pr__pfet_01v8_lvt ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X89 a_n2848_n452.t44 minus.t10 a_n3106_n452.t52 gnd.t267 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=2.73 ps=14.78 w=7 l=0.9
X90 CSoutput.t55 commonsourceibias.t60 gnd.t290 gnd.t7 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X91 gnd.t285 commonsourceibias.t61 CSoutput.t54 gnd.t53 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=1.155 ps=7.33 w=7 l=1
X92 gnd.t161 gnd.t158 gnd.t160 gnd.t159 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=0 ps=0 w=7 l=1
X93 commonsourceibias.t29 commonsourceibias.t28 gnd.t238 gnd.t17 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X94 vdd.t81 vdd.t79 vdd.t80 vdd.t33 sky130_fd_pr__pfet_01v8_lvt ad=3.12 pd=16.78 as=0 ps=0 w=8 l=0.5
X95 CSoutput.t53 commonsourceibias.t62 gnd.t213 gnd.t212 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=2.73 ps=14.78 w=7 l=1
X96 CSoutput.t102 a_n1986_8322.t1 sky130_fd_pr__cap_mim_m3_1 l=12 w=12
X97 outputibias.t3 outputibias.t2 gnd.t288 gnd.t287 sky130_fd_pr__nfet_01v8 ad=2.34 pd=12.78 as=2.34 ps=12.78 w=6 l=2
X98 vdd.t140 a_n5644_8799.t55 CSoutput.t86 vdd.t125 sky130_fd_pr__pfet_01v8_lvt ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X99 vdd.t78 vdd.t76 vdd.t77 vdd.t62 sky130_fd_pr__pfet_01v8_lvt ad=3.51 pd=18.78 as=0 ps=0 w=9 l=0.5
X100 vdd.t75 vdd.t72 vdd.t74 vdd.t73 sky130_fd_pr__pfet_01v8_lvt ad=3.51 pd=18.78 as=0 ps=0 w=9 l=0.5
X101 a_n3106_n452.t10 diffpairibias.t18 gnd.t49 gnd.t48 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=2.73 ps=14.78 w=7 l=1
X102 vdd.t71 vdd.t68 vdd.t70 vdd.t69 sky130_fd_pr__pfet_01v8_lvt ad=3.51 pd=18.78 as=0 ps=0 w=9 l=0.5
X103 gnd.t157 gnd.t155 minus.t4 gnd.t156 sky130_fd_pr__nfet_01v8 ad=0.39 pd=2.78 as=0.165 ps=1.33 w=1 l=0.5
X104 gnd.t154 gnd.t152 gnd.t153 gnd.t99 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=0 ps=0 w=7 l=0.9
X105 commonsourceibias.t27 commonsourceibias.t26 gnd.t8 gnd.t7 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X106 vdd.t20 a_n2848_n452.t53 a_n1986_8322.t10 vdd.t19 sky130_fd_pr__pfet_01v8_lvt ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X107 vdd.t67 vdd.t65 vdd.t66 vdd.t58 sky130_fd_pr__pfet_01v8_lvt ad=3.51 pd=18.78 as=0 ps=0 w=9 l=0.5
X108 CSoutput.t95 a_n5644_8799.t56 vdd.t139 vdd.t138 sky130_fd_pr__pfet_01v8_lvt ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X109 a_n1986_8322.t9 a_n2848_n452.t54 vdd.t16 vdd.t15 sky130_fd_pr__pfet_01v8_lvt ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X110 vdd.t137 a_n5644_8799.t57 CSoutput.t73 vdd.t136 sky130_fd_pr__pfet_01v8_lvt ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X111 gnd.t244 commonsourceibias.t24 commonsourceibias.t25 gnd.t51 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X112 gnd.t208 commonsourceibias.t63 CSoutput.t52 gnd.t207 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X113 vdd.t18 a_n2848_n452.t55 a_n1808_13878.t6 vdd.t17 sky130_fd_pr__pfet_01v8_lvt ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X114 gnd.t151 gnd.t149 plus.t3 gnd.t150 sky130_fd_pr__nfet_01v8 ad=0.39 pd=2.78 as=0.165 ps=1.33 w=1 l=0.5
X115 gnd.t260 commonsourceibias.t64 CSoutput.t51 gnd.t40 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X116 a_n2848_n452.t3 minus.t11 a_n3106_n452.t3 gnd.t6 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.9
X117 a_n5644_8799.t3 plus.t14 a_n3106_n452.t31 gnd.t20 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=2.73 ps=14.78 w=7 l=0.9
X118 gnd.t181 commonsourceibias.t65 CSoutput.t50 gnd.t180 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=1.155 ps=7.33 w=7 l=1
X119 vdd.t64 vdd.t61 vdd.t63 vdd.t62 sky130_fd_pr__pfet_01v8_lvt ad=3.51 pd=18.78 as=0 ps=0 w=9 l=0.5
X120 a_n5644_8799.t9 plus.t15 a_n3106_n452.t30 gnd.t29 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.9
X121 a_n2848_n452.t42 minus.t12 a_n3106_n452.t50 gnd.t262 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.9
X122 diffpairibias.t11 diffpairibias.t10 gnd.t2 gnd.t1 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=2.73 ps=14.78 w=7 l=1
X123 vdd.t161 CSoutput.t103 output.t10 gnd.t223 sky130_fd_pr__nfet_01v8_lvt ad=0.825 pd=5.33 as=0.825 ps=5.33 w=5 l=1
X124 vdd.t60 vdd.t57 vdd.t59 vdd.t58 sky130_fd_pr__pfet_01v8_lvt ad=3.51 pd=18.78 as=0 ps=0 w=9 l=0.5
X125 vdd.t135 a_n5644_8799.t58 CSoutput.t5 vdd.t134 sky130_fd_pr__pfet_01v8_lvt ad=3.12 pd=16.78 as=1.32 ps=8.33 w=8 l=0.5
X126 gnd.t268 commonsourceibias.t66 CSoutput.t49 gnd.t246 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X127 outputibias.t1 outputibias.t0 gnd.t191 gnd.t190 sky130_fd_pr__nfet_01v8 ad=2.34 pd=12.78 as=2.34 ps=12.78 w=6 l=2
X128 a_n5644_8799.t5 a_n2848_n452.t56 a_n1986_8322.t20 vdd.t1 sky130_fd_pr__pfet_01v8_lvt ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X129 a_n1986_8322.t8 a_n2848_n452.t57 vdd.t3 vdd.t2 sky130_fd_pr__pfet_01v8_lvt ad=3.51 pd=18.78 as=1.485 ps=9.33 w=9 l=0.5
X130 vdd.t56 vdd.t53 vdd.t55 vdd.t54 sky130_fd_pr__pfet_01v8_lvt ad=3.51 pd=18.78 as=0 ps=0 w=9 l=0.5
X131 gnd.t192 commonsourceibias.t67 CSoutput.t48 gnd.t178 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X132 a_n2848_n452.t31 a_n2848_n452.t30 a_n1808_13878.t12 vdd.t193 sky130_fd_pr__pfet_01v8_lvt ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X133 a_n3106_n452.t47 minus.t13 a_n2848_n452.t17 gnd.t248 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.9
X134 CSoutput.t104 a_n1986_8322.t3 sky130_fd_pr__cap_mim_m3_1 l=12 w=12
X135 a_n5644_8799.t30 a_n2848_n452.t58 a_n1986_8322.t19 vdd.t0 sky130_fd_pr__pfet_01v8_lvt ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X136 CSoutput.t47 commonsourceibias.t68 gnd.t265 gnd.t12 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X137 CSoutput.t105 a_n1986_8322.t2 sky130_fd_pr__cap_mim_m3_1 l=12 w=12
X138 a_n1808_13878.t11 a_n2848_n452.t24 a_n2848_n452.t25 vdd.t14 sky130_fd_pr__pfet_01v8_lvt ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X139 a_n3106_n452.t29 plus.t16 a_n5644_8799.t20 gnd.t231 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.9
X140 a_n2848_n452.t12 minus.t14 a_n3106_n452.t42 gnd.t242 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.9
X141 vdd.t195 a_n2848_n452.t59 a_n1986_8322.t7 vdd.t194 sky130_fd_pr__pfet_01v8_lvt ad=1.485 pd=9.33 as=3.51 ps=18.78 w=9 l=0.5
X142 vdd.t52 vdd.t50 vdd.t51 vdd.t44 sky130_fd_pr__pfet_01v8_lvt ad=3.12 pd=16.78 as=0 ps=0 w=8 l=0.5
X143 gnd.t148 gnd.t145 gnd.t147 gnd.t146 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=0 ps=0 w=7 l=1
X144 a_n3106_n452.t41 diffpairibias.t19 gnd.t237 gnd.t236 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=2.73 ps=14.78 w=7 l=1
X145 CSoutput.t15 a_n5644_8799.t59 vdd.t133 vdd.t128 sky130_fd_pr__pfet_01v8_lvt ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X146 CSoutput.t46 commonsourceibias.t69 gnd.t42 gnd.t7 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X147 a_n5644_8799.t19 plus.t17 a_n3106_n452.t28 gnd.t228 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.9
X148 CSoutput.t45 commonsourceibias.t70 gnd.t226 gnd.t225 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X149 a_n3106_n452.t49 diffpairibias.t20 gnd.t254 gnd.t253 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=2.73 ps=14.78 w=7 l=1
X150 vdd.t132 a_n5644_8799.t60 CSoutput.t13 vdd.t99 sky130_fd_pr__pfet_01v8_lvt ad=3.12 pd=16.78 as=1.32 ps=8.33 w=8 l=0.5
X151 gnd.t54 commonsourceibias.t71 CSoutput.t44 gnd.t53 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=1.155 ps=7.33 w=7 l=1
X152 CSoutput.t43 commonsourceibias.t72 gnd.t33 gnd.t32 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X153 a_n5644_8799.t17 plus.t18 a_n3106_n452.t27 gnd.t36 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.9
X154 vdd.t131 a_n5644_8799.t61 CSoutput.t81 vdd.t114 sky130_fd_pr__pfet_01v8_lvt ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X155 minus.t3 gnd.t142 gnd.t144 gnd.t143 sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.5
X156 gnd.t141 gnd.t139 gnd.t140 gnd.t95 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=0 ps=0 w=7 l=1
X157 diffpairibias.t9 diffpairibias.t8 gnd.t256 gnd.t255 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=2.73 ps=14.78 w=7 l=1
X158 a_n2848_n452.t0 minus.t15 a_n3106_n452.t0 gnd.t3 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.9
X159 a_n3106_n452.t26 plus.t19 a_n5644_8799.t11 gnd.t5 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.9
X160 CSoutput.t92 a_n5644_8799.t62 vdd.t130 vdd.t118 sky130_fd_pr__pfet_01v8_lvt ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X161 CSoutput.t42 commonsourceibias.t73 gnd.t210 gnd.t209 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=2.73 ps=14.78 w=7 l=1
X162 gnd.t269 commonsourceibias.t74 CSoutput.t41 gnd.t218 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X163 vdd.t49 vdd.t47 vdd.t48 vdd.t29 sky130_fd_pr__pfet_01v8_lvt ad=3.12 pd=16.78 as=0 ps=0 w=8 l=0.5
X164 a_n1808_13878.t5 a_n2848_n452.t60 vdd.t197 vdd.t196 sky130_fd_pr__pfet_01v8_lvt ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X165 vdd.t199 a_n2848_n452.t61 a_n1808_13878.t4 vdd.t198 sky130_fd_pr__pfet_01v8_lvt ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X166 gnd.t220 commonsourceibias.t22 commonsourceibias.t23 gnd.t60 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X167 gnd.t264 commonsourceibias.t75 CSoutput.t40 gnd.t180 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=1.155 ps=7.33 w=7 l=1
X168 output.t9 CSoutput.t106 vdd.t168 gnd.t9 sky130_fd_pr__nfet_01v8_lvt ad=0.825 pd=5.33 as=0.825 ps=5.33 w=5 l=1
X169 vdd.t46 vdd.t43 vdd.t45 vdd.t44 sky130_fd_pr__pfet_01v8_lvt ad=3.12 pd=16.78 as=0 ps=0 w=8 l=0.5
X170 gnd.t247 commonsourceibias.t76 CSoutput.t39 gnd.t246 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X171 a_n3106_n452.t44 minus.t16 a_n2848_n452.t14 gnd.t21 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.9
X172 diffpairibias.t7 diffpairibias.t6 gnd.t230 gnd.t229 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=2.73 ps=14.78 w=7 l=1
X173 CSoutput.t91 a_n5644_8799.t63 vdd.t129 vdd.t128 sky130_fd_pr__pfet_01v8_lvt ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X174 gnd.t283 commonsourceibias.t20 commonsourceibias.t21 gnd.t246 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X175 output.t8 CSoutput.t107 vdd.t173 gnd.t10 sky130_fd_pr__nfet_01v8_lvt ad=0.825 pd=5.33 as=0.825 ps=5.33 w=5 l=1
X176 vdd.t127 a_n5644_8799.t64 CSoutput.t18 vdd.t99 sky130_fd_pr__pfet_01v8_lvt ad=3.12 pd=16.78 as=1.32 ps=8.33 w=8 l=0.5
X177 CSoutput.t38 commonsourceibias.t77 gnd.t31 gnd.t30 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X178 a_n3106_n452.t45 minus.t17 a_n2848_n452.t15 gnd.t0 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.9
X179 a_n3106_n452.t25 plus.t20 a_n5644_8799.t25 gnd.t11 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=1.155 ps=7.33 w=7 l=0.9
X180 gnd.t138 gnd.t136 gnd.t137 gnd.t95 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=0 ps=0 w=7 l=1
X181 gnd.t135 gnd.t133 gnd.t134 gnd.t74 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=0 ps=0 w=7 l=1
X182 a_n1986_8322.t18 a_n2848_n452.t62 a_n5644_8799.t8 vdd.t11 sky130_fd_pr__pfet_01v8_lvt ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X183 CSoutput.t37 commonsourceibias.t78 gnd.t65 gnd.t12 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X184 a_n3106_n452.t13 minus.t18 a_n2848_n452.t10 gnd.t19 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.9
X185 vdd.t126 a_n5644_8799.t65 CSoutput.t12 vdd.t125 sky130_fd_pr__pfet_01v8_lvt ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X186 CSoutput.t82 a_n5644_8799.t66 vdd.t124 vdd.t105 sky130_fd_pr__pfet_01v8_lvt ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X187 vdd.t123 a_n5644_8799.t67 CSoutput.t70 vdd.t114 sky130_fd_pr__pfet_01v8_lvt ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X188 vdd.t13 a_n2848_n452.t63 a_n1986_8322.t6 vdd.t12 sky130_fd_pr__pfet_01v8_lvt ad=1.485 pd=9.33 as=3.51 ps=18.78 w=9 l=0.5
X189 gnd.t227 commonsourceibias.t18 commonsourceibias.t19 gnd.t15 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X190 a_n1808_13878.t3 a_n2848_n452.t64 vdd.t192 vdd.t191 sky130_fd_pr__pfet_01v8_lvt ad=3.51 pd=18.78 as=1.485 ps=9.33 w=9 l=0.5
X191 gnd.t132 gnd.t129 gnd.t131 gnd.t130 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=0 ps=0 w=7 l=1
X192 minus.t2 gnd.t126 gnd.t128 gnd.t127 sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.5
X193 CSoutput.t36 commonsourceibias.t79 gnd.t18 gnd.t17 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X194 a_n3106_n452.t15 diffpairibias.t21 gnd.t204 gnd.t203 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=2.73 ps=14.78 w=7 l=1
X195 CSoutput.t69 a_n5644_8799.t68 vdd.t122 vdd.t118 sky130_fd_pr__pfet_01v8_lvt ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X196 a_n5644_8799.t23 plus.t21 a_n3106_n452.t24 gnd.t37 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.9
X197 a_n2848_n452.t13 minus.t19 a_n3106_n452.t43 gnd.t235 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.9
X198 CSoutput.t35 commonsourceibias.t80 gnd.t270 gnd.t225 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X199 output.t7 CSoutput.t108 vdd.t174 gnd.t67 sky130_fd_pr__nfet_01v8_lvt ad=0.825 pd=5.33 as=0.825 ps=5.33 w=5 l=1
X200 CSoutput.t7 a_n5644_8799.t69 vdd.t121 vdd.t116 sky130_fd_pr__pfet_01v8_lvt ad=1.32 pd=8.33 as=3.12 ps=16.78 w=8 l=0.5
X201 a_n3106_n452.t14 minus.t20 a_n2848_n452.t11 gnd.t200 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=1.155 ps=7.33 w=7 l=0.9
X202 CSoutput.t109 a_n1986_8322.t1 sky130_fd_pr__cap_mim_m3_1 l=12 w=12
X203 vdd.t42 vdd.t40 vdd.t41 vdd.t29 sky130_fd_pr__pfet_01v8_lvt ad=3.12 pd=16.78 as=0 ps=0 w=8 l=0.5
X204 CSoutput.t34 commonsourceibias.t81 gnd.t239 gnd.t32 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X205 gnd.t115 gnd.t112 gnd.t114 gnd.t113 sky130_fd_pr__nfet_01v8_lvt ad=1.95 pd=10.78 as=0 ps=0 w=5 l=1
X206 a_n1986_8322.t17 a_n2848_n452.t65 a_n5644_8799.t28 vdd.t193 sky130_fd_pr__pfet_01v8_lvt ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X207 vdd.t9 a_n2848_n452.t66 a_n1986_8322.t5 vdd.t8 sky130_fd_pr__pfet_01v8_lvt ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X208 vdd.t120 a_n5644_8799.t70 CSoutput.t71 vdd.t107 sky130_fd_pr__pfet_01v8_lvt ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X209 CSoutput.t80 a_n5644_8799.t71 vdd.t119 vdd.t118 sky130_fd_pr__pfet_01v8_lvt ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X210 gnd.t16 commonsourceibias.t82 CSoutput.t33 gnd.t15 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X211 output.t18 outputibias.t9 gnd.t276 gnd.t275 sky130_fd_pr__nfet_01v8 ad=2.34 pd=12.78 as=2.34 ps=12.78 w=6 l=2
X212 a_n3106_n452.t46 minus.t21 a_n2848_n452.t16 gnd.t14 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.9
X213 gnd.t125 gnd.t123 gnd.t124 gnd.t88 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=0 ps=0 w=7 l=1
X214 vdd.t169 CSoutput.t110 output.t6 gnd.t68 sky130_fd_pr__nfet_01v8_lvt ad=0.825 pd=5.33 as=0.825 ps=5.33 w=5 l=1
X215 a_n3106_n452.t12 minus.t22 a_n2848_n452.t9 gnd.t69 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.9
X216 gnd.t122 gnd.t120 gnd.t121 gnd.t88 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=0 ps=0 w=7 l=1
X217 output.t17 outputibias.t10 gnd.t279 gnd.t278 sky130_fd_pr__nfet_01v8 ad=2.34 pd=12.78 as=2.34 ps=12.78 w=6 l=2
X218 diffpairibias.t5 diffpairibias.t4 gnd.t27 gnd.t26 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=2.73 ps=14.78 w=7 l=1
X219 vdd.t39 vdd.t36 vdd.t38 vdd.t37 sky130_fd_pr__pfet_01v8_lvt ad=3.51 pd=18.78 as=0 ps=0 w=9 l=0.5
X220 vdd.t35 vdd.t32 vdd.t34 vdd.t33 sky130_fd_pr__pfet_01v8_lvt ad=3.12 pd=16.78 as=0 ps=0 w=8 l=0.5
X221 a_n1808_13878.t10 a_n2848_n452.t38 a_n2848_n452.t39 vdd.t190 sky130_fd_pr__pfet_01v8_lvt ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X222 gnd.t224 commonsourceibias.t83 CSoutput.t32 gnd.t218 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X223 CSoutput.t31 commonsourceibias.t84 gnd.t250 gnd.t209 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=2.73 ps=14.78 w=7 l=1
X224 a_n1986_8322.t16 a_n2848_n452.t67 a_n5644_8799.t7 vdd.t10 sky130_fd_pr__pfet_01v8_lvt ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X225 gnd.t119 gnd.t116 gnd.t118 gnd.t117 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=0 ps=0 w=7 l=0.9
X226 gnd.t61 commonsourceibias.t85 CSoutput.t30 gnd.t60 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X227 gnd.t258 commonsourceibias.t16 commonsourceibias.t17 gnd.t180 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=1.155 ps=7.33 w=7 l=1
X228 a_n3106_n452.t5 minus.t23 a_n2848_n452.t5 gnd.t28 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.9
X229 gnd.t111 gnd.t108 gnd.t110 gnd.t109 sky130_fd_pr__nfet_01v8 ad=2.34 pd=12.78 as=0 ps=0 w=6 l=2
X230 vdd.t176 CSoutput.t111 output.t5 gnd.t183 sky130_fd_pr__nfet_01v8_lvt ad=0.825 pd=5.33 as=0.825 ps=5.33 w=5 l=1
X231 output.t4 CSoutput.t112 vdd.t172 gnd.t184 sky130_fd_pr__nfet_01v8_lvt ad=0.825 pd=5.33 as=0.825 ps=5.33 w=5 l=1
X232 CSoutput.t4 a_n5644_8799.t72 vdd.t117 vdd.t116 sky130_fd_pr__pfet_01v8_lvt ad=1.32 pd=8.33 as=3.12 ps=16.78 w=8 l=0.5
X233 a_n1986_8322.t4 a_n2848_n452.t68 vdd.t183 vdd.t182 sky130_fd_pr__pfet_01v8_lvt ad=3.51 pd=18.78 as=1.485 ps=9.33 w=9 l=0.5
X234 gnd.t107 gnd.t105 plus.t2 gnd.t106 sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.5
X235 gnd.t104 gnd.t102 gnd.t103 gnd.t74 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=0 ps=0 w=7 l=1
X236 CSoutput.t29 commonsourceibias.t86 gnd.t55 gnd.t30 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X237 gnd.t101 gnd.t98 gnd.t100 gnd.t99 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=0 ps=0 w=7 l=0.9
X238 CSoutput.t28 commonsourceibias.t87 gnd.t274 gnd.t195 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X239 gnd.t97 gnd.t94 gnd.t96 gnd.t95 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=0 ps=0 w=7 l=1
X240 output.t3 CSoutput.t113 vdd.t162 gnd.t185 sky130_fd_pr__nfet_01v8_lvt ad=0.825 pd=5.33 as=0.825 ps=5.33 w=5 l=1
X241 vdd.t185 a_n2848_n452.t69 a_n1808_13878.t2 vdd.t184 sky130_fd_pr__pfet_01v8_lvt ad=1.485 pd=9.33 as=3.51 ps=18.78 w=9 l=0.5
X242 vdd.t31 vdd.t28 vdd.t30 vdd.t29 sky130_fd_pr__pfet_01v8_lvt ad=3.12 pd=16.78 as=0 ps=0 w=8 l=0.5
X243 a_n1986_8322.t15 a_n2848_n452.t70 a_n5644_8799.t26 vdd.t178 sky130_fd_pr__pfet_01v8_lvt ad=3.51 pd=18.78 as=1.485 ps=9.33 w=9 l=0.5
X244 a_n3106_n452.t23 plus.t22 a_n5644_8799.t35 gnd.t4 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.9
X245 output.t16 outputibias.t11 gnd.t202 gnd.t201 sky130_fd_pr__nfet_01v8 ad=2.34 pd=12.78 as=2.34 ps=12.78 w=6 l=2
X246 vdd.t27 vdd.t25 vdd.t26 vdd.t22 sky130_fd_pr__pfet_01v8_lvt ad=3.12 pd=16.78 as=0 ps=0 w=8 l=0.5
X247 a_n5644_8799.t27 a_n2848_n452.t71 a_n1986_8322.t14 vdd.t190 sky130_fd_pr__pfet_01v8_lvt ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X248 a_n1808_13878.t1 a_n2848_n452.t72 vdd.t6 vdd.t5 sky130_fd_pr__pfet_01v8_lvt ad=3.51 pd=18.78 as=1.485 ps=9.33 w=9 l=0.5
X249 vdd.t115 a_n5644_8799.t73 CSoutput.t8 vdd.t114 sky130_fd_pr__pfet_01v8_lvt ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X250 CSoutput.t85 a_n5644_8799.t74 vdd.t113 vdd.t112 sky130_fd_pr__pfet_01v8_lvt ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X251 gnd.t93 gnd.t91 minus.t1 gnd.t92 sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.39 ps=2.78 w=1 l=0.5
X252 a_n2848_n452.t6 minus.t24 a_n3106_n452.t6 gnd.t29 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.9
X253 a_n5644_8799.t31 plus.t23 a_n3106_n452.t22 gnd.t262 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.9
X254 CSoutput.t27 commonsourceibias.t88 gnd.t261 gnd.t17 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X255 a_n2848_n452.t43 minus.t25 a_n3106_n452.t51 gnd.t266 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.9
X256 commonsourceibias.t15 commonsourceibias.t14 gnd.t43 gnd.t32 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X257 gnd.t39 commonsourceibias.t89 CSoutput.t26 gnd.t38 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X258 vdd.t163 CSoutput.t114 output.t2 gnd.t198 sky130_fd_pr__nfet_01v8_lvt ad=0.825 pd=5.33 as=0.825 ps=5.33 w=5 l=1
X259 gnd.t62 commonsourceibias.t90 CSoutput.t25 gnd.t15 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X260 CSoutput.t17 a_n5644_8799.t75 vdd.t111 vdd.t105 sky130_fd_pr__pfet_01v8_lvt ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X261 a_n1808_13878.t9 a_n2848_n452.t18 a_n2848_n452.t19 vdd.t1 sky130_fd_pr__pfet_01v8_lvt ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X262 gnd.t90 gnd.t87 gnd.t89 gnd.t88 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=0 ps=0 w=7 l=1
X263 a_n3106_n452.t54 minus.t26 a_n2848_n452.t46 gnd.t231 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.9
X264 a_n3106_n452.t9 diffpairibias.t22 gnd.t47 gnd.t46 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=2.73 ps=14.78 w=7 l=1
X265 gnd.t273 commonsourceibias.t91 CSoutput.t24 gnd.t193 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X266 commonsourceibias.t13 commonsourceibias.t12 gnd.t243 gnd.t195 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X267 a_n5644_8799.t32 plus.t24 a_n3106_n452.t21 gnd.t267 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=2.73 ps=14.78 w=7 l=0.9
X268 CSoutput.t16 a_n5644_8799.t76 vdd.t110 vdd.t103 sky130_fd_pr__pfet_01v8_lvt ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X269 vdd.t109 a_n5644_8799.t77 CSoutput.t2 vdd.t101 sky130_fd_pr__pfet_01v8_lvt ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X270 diffpairibias.t3 diffpairibias.t2 gnd.t216 gnd.t215 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=2.73 ps=14.78 w=7 l=1
X271 a_n5644_8799.t6 a_n2848_n452.t73 a_n1986_8322.t13 vdd.t7 sky130_fd_pr__pfet_01v8_lvt ad=1.485 pd=9.33 as=3.51 ps=18.78 w=9 l=0.5
X272 a_n2848_n452.t33 a_n2848_n452.t32 a_n1808_13878.t8 vdd.t178 sky130_fd_pr__pfet_01v8_lvt ad=3.51 pd=18.78 as=1.485 ps=9.33 w=9 l=0.5
X273 gnd.t86 gnd.t84 plus.t1 gnd.t85 sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.39 ps=2.78 w=1 l=0.5
X274 a_n2848_n452.t47 minus.t27 a_n3106_n452.t55 gnd.t228 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.9
X275 vdd.t108 a_n5644_8799.t78 CSoutput.t78 vdd.t107 sky130_fd_pr__pfet_01v8_lvt ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X276 commonsourceibias.t11 commonsourceibias.t10 gnd.t13 gnd.t12 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X277 gnd.t66 commonsourceibias.t92 CSoutput.t23 gnd.t60 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X278 vdd.t24 vdd.t21 vdd.t23 vdd.t22 sky130_fd_pr__pfet_01v8_lvt ad=3.12 pd=16.78 as=0 ps=0 w=8 l=0.5
X279 CSoutput.t115 a_n1986_8322.t0 sky130_fd_pr__cap_mim_m3_1 l=12 w=12
X280 diffpairibias.t1 diffpairibias.t0 gnd.t281 gnd.t280 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=2.73 ps=14.78 w=7 l=1
X281 CSoutput.t22 commonsourceibias.t93 gnd.t45 gnd.t44 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X282 gnd.t83 gnd.t80 gnd.t82 gnd.t81 sky130_fd_pr__nfet_01v8_lvt ad=1.95 pd=10.78 as=0 ps=0 w=5 l=1
X283 output.t1 CSoutput.t116 vdd.t170 gnd.t199 sky130_fd_pr__nfet_01v8_lvt ad=0.825 pd=5.33 as=0.825 ps=5.33 w=5 l=1
X284 plus.t0 gnd.t77 gnd.t79 gnd.t78 sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.5
X285 gnd.t76 gnd.t73 gnd.t75 gnd.t74 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=0 ps=0 w=7 l=1
X286 CSoutput.t21 commonsourceibias.t94 gnd.t196 gnd.t195 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X287 commonsourceibias.t9 commonsourceibias.t8 gnd.t277 gnd.t232 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X288 gnd.t72 gnd.t70 minus.t0 gnd.t71 sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.5
X289 a_n5644_8799.t34 plus.t25 a_n3106_n452.t20 gnd.t3 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.9
X290 vdd.t180 a_n2848_n452.t74 a_n1808_13878.t0 vdd.t179 sky130_fd_pr__pfet_01v8_lvt ad=1.485 pd=9.33 as=3.51 ps=18.78 w=9 l=0.5
X291 CSoutput.t88 a_n5644_8799.t79 vdd.t106 vdd.t105 sky130_fd_pr__pfet_01v8_lvt ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X292 CSoutput.t20 commonsourceibias.t95 gnd.t197 gnd.t34 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X293 a_n5644_8799.t12 plus.t26 a_n3106_n452.t19 gnd.t6 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.9
X294 a_n2848_n452.t45 minus.t28 a_n3106_n452.t53 gnd.t20 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=2.73 ps=14.78 w=7 l=0.9
X295 output.t0 CSoutput.t117 vdd.t166 gnd.t282 sky130_fd_pr__nfet_01v8_lvt ad=1.95 pd=10.78 as=0.825 ps=5.33 w=5 l=1
X296 gnd.t245 commonsourceibias.t6 commonsourceibias.t7 gnd.t38 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X297 commonsourceibias.t5 commonsourceibias.t4 gnd.t259 gnd.t225 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X298 CSoutput.t19 a_n5644_8799.t80 vdd.t104 vdd.t103 sky130_fd_pr__pfet_01v8_lvt ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X299 vdd.t102 a_n5644_8799.t81 CSoutput.t83 vdd.t101 sky130_fd_pr__pfet_01v8_lvt ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X300 a_n1986_8322.t12 a_n2848_n452.t75 a_n5644_8799.t21 vdd.t181 sky130_fd_pr__pfet_01v8_lvt ad=3.51 pd=18.78 as=1.485 ps=9.33 w=9 l=0.5
X301 a_n3106_n452.t18 plus.t27 a_n5644_8799.t4 gnd.t21 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.9
X302 commonsourceibias.t3 commonsourceibias.t2 gnd.t217 gnd.t209 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=2.73 ps=14.78 w=7 l=1
X303 vdd.t100 a_n5644_8799.t82 CSoutput.t89 vdd.t99 sky130_fd_pr__pfet_01v8_lvt ad=3.12 pd=16.78 as=1.32 ps=8.33 w=8 l=0.5
X304 CSoutput.t93 a_n5644_8799.t83 vdd.t98 vdd.t97 sky130_fd_pr__pfet_01v8_lvt ad=1.32 pd=8.33 as=3.12 ps=16.78 w=8 l=0.5
X305 a_n3106_n452.t17 plus.t28 a_n5644_8799.t33 gnd.t248 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.9
X306 gnd.t234 commonsourceibias.t0 commonsourceibias.t1 gnd.t207 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X307 a_n3106_n452.t48 diffpairibias.t23 gnd.t252 gnd.t251 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=2.73 ps=14.78 w=7 l=1
R0 gnd.n5991 gnd.n635 1087.89
R1 gnd.n3878 gnd.n3570 939.716
R2 gnd.n6602 gnd.n84 838.452
R3 gnd.n6765 gnd.n80 838.452
R4 gnd.n6391 gnd.n330 838.452
R5 gnd.n6444 gnd.n332 838.452
R6 gnd.n1096 gnd.n1084 838.452
R7 gnd.n4188 gnd.n4187 838.452
R8 gnd.n3706 gnd.n3598 838.452
R9 gnd.n3880 gnd.n2115 838.452
R10 gnd.n6763 gnd.n86 819.232
R11 gnd.n154 gnd.n82 819.232
R12 gnd.n6317 gnd.n329 819.232
R13 gnd.n6446 gnd.n327 819.232
R14 gnd.n5438 gnd.n1089 819.232
R15 gnd.n4141 gnd.n1981 819.232
R16 gnd.n3800 gnd.n3799 819.232
R17 gnd.n3876 gnd.n2111 819.232
R18 gnd.n4252 gnd.n1837 771.183
R19 gnd.n5196 gnd.n337 771.183
R20 gnd.n4233 gnd.n1840 771.183
R21 gnd.n5198 gnd.n1418 771.183
R22 gnd.n3478 gnd.n2121 766.379
R23 gnd.n3481 gnd.n3480 766.379
R24 gnd.n2719 gnd.n2622 766.379
R25 gnd.n2715 gnd.n2620 766.379
R26 gnd.n3569 gnd.n2143 756.769
R27 gnd.n3472 gnd.n3471 756.769
R28 gnd.n2812 gnd.n2529 756.769
R29 gnd.n2810 gnd.n2532 756.769
R30 gnd.n5663 gnd.n827 655.866
R31 gnd.n5990 gnd.n636 655.866
R32 gnd.n6203 gnd.n6202 655.866
R33 gnd.n5495 gnd.n997 655.866
R34 gnd.n5664 gnd.n5663 585
R35 gnd.n5663 gnd.n5662 585
R36 gnd.n831 gnd.n830 585
R37 gnd.n5661 gnd.n831 585
R38 gnd.n5659 gnd.n5658 585
R39 gnd.n5660 gnd.n5659 585
R40 gnd.n5657 gnd.n833 585
R41 gnd.n833 gnd.n832 585
R42 gnd.n5656 gnd.n5655 585
R43 gnd.n5655 gnd.n5654 585
R44 gnd.n838 gnd.n837 585
R45 gnd.n5653 gnd.n838 585
R46 gnd.n5651 gnd.n5650 585
R47 gnd.n5652 gnd.n5651 585
R48 gnd.n5649 gnd.n840 585
R49 gnd.n840 gnd.n839 585
R50 gnd.n5648 gnd.n5647 585
R51 gnd.n5647 gnd.n5646 585
R52 gnd.n846 gnd.n845 585
R53 gnd.n5645 gnd.n846 585
R54 gnd.n5643 gnd.n5642 585
R55 gnd.n5644 gnd.n5643 585
R56 gnd.n5641 gnd.n848 585
R57 gnd.n848 gnd.n847 585
R58 gnd.n5640 gnd.n5639 585
R59 gnd.n5639 gnd.n5638 585
R60 gnd.n854 gnd.n853 585
R61 gnd.n5637 gnd.n854 585
R62 gnd.n5635 gnd.n5634 585
R63 gnd.n5636 gnd.n5635 585
R64 gnd.n5633 gnd.n856 585
R65 gnd.n856 gnd.n855 585
R66 gnd.n5632 gnd.n5631 585
R67 gnd.n5631 gnd.n5630 585
R68 gnd.n862 gnd.n861 585
R69 gnd.n5629 gnd.n862 585
R70 gnd.n5627 gnd.n5626 585
R71 gnd.n5628 gnd.n5627 585
R72 gnd.n5625 gnd.n864 585
R73 gnd.n864 gnd.n863 585
R74 gnd.n5624 gnd.n5623 585
R75 gnd.n5623 gnd.n5622 585
R76 gnd.n870 gnd.n869 585
R77 gnd.n5621 gnd.n870 585
R78 gnd.n5619 gnd.n5618 585
R79 gnd.n5620 gnd.n5619 585
R80 gnd.n5617 gnd.n872 585
R81 gnd.n872 gnd.n871 585
R82 gnd.n5616 gnd.n5615 585
R83 gnd.n5615 gnd.n5614 585
R84 gnd.n878 gnd.n877 585
R85 gnd.n5613 gnd.n878 585
R86 gnd.n5611 gnd.n5610 585
R87 gnd.n5612 gnd.n5611 585
R88 gnd.n5609 gnd.n880 585
R89 gnd.n880 gnd.n879 585
R90 gnd.n5608 gnd.n5607 585
R91 gnd.n5607 gnd.n5606 585
R92 gnd.n886 gnd.n885 585
R93 gnd.n5605 gnd.n886 585
R94 gnd.n5603 gnd.n5602 585
R95 gnd.n5604 gnd.n5603 585
R96 gnd.n5601 gnd.n888 585
R97 gnd.n888 gnd.n887 585
R98 gnd.n5600 gnd.n5599 585
R99 gnd.n5599 gnd.n5598 585
R100 gnd.n894 gnd.n893 585
R101 gnd.n5597 gnd.n894 585
R102 gnd.n5595 gnd.n5594 585
R103 gnd.n5596 gnd.n5595 585
R104 gnd.n5593 gnd.n896 585
R105 gnd.n896 gnd.n895 585
R106 gnd.n5592 gnd.n5591 585
R107 gnd.n5591 gnd.n5590 585
R108 gnd.n902 gnd.n901 585
R109 gnd.n5589 gnd.n902 585
R110 gnd.n5587 gnd.n5586 585
R111 gnd.n5588 gnd.n5587 585
R112 gnd.n5585 gnd.n904 585
R113 gnd.n904 gnd.n903 585
R114 gnd.n5584 gnd.n5583 585
R115 gnd.n5583 gnd.n5582 585
R116 gnd.n910 gnd.n909 585
R117 gnd.n5581 gnd.n910 585
R118 gnd.n5579 gnd.n5578 585
R119 gnd.n5580 gnd.n5579 585
R120 gnd.n5577 gnd.n912 585
R121 gnd.n912 gnd.n911 585
R122 gnd.n5576 gnd.n5575 585
R123 gnd.n5575 gnd.n5574 585
R124 gnd.n918 gnd.n917 585
R125 gnd.n5573 gnd.n918 585
R126 gnd.n5571 gnd.n5570 585
R127 gnd.n5572 gnd.n5571 585
R128 gnd.n5569 gnd.n920 585
R129 gnd.n920 gnd.n919 585
R130 gnd.n5568 gnd.n5567 585
R131 gnd.n5567 gnd.n5566 585
R132 gnd.n926 gnd.n925 585
R133 gnd.n5565 gnd.n926 585
R134 gnd.n5563 gnd.n5562 585
R135 gnd.n5564 gnd.n5563 585
R136 gnd.n5561 gnd.n928 585
R137 gnd.n928 gnd.n927 585
R138 gnd.n5560 gnd.n5559 585
R139 gnd.n5559 gnd.n5558 585
R140 gnd.n934 gnd.n933 585
R141 gnd.n5557 gnd.n934 585
R142 gnd.n5555 gnd.n5554 585
R143 gnd.n5556 gnd.n5555 585
R144 gnd.n5553 gnd.n936 585
R145 gnd.n936 gnd.n935 585
R146 gnd.n5552 gnd.n5551 585
R147 gnd.n5551 gnd.n5550 585
R148 gnd.n942 gnd.n941 585
R149 gnd.n5549 gnd.n942 585
R150 gnd.n5547 gnd.n5546 585
R151 gnd.n5548 gnd.n5547 585
R152 gnd.n5545 gnd.n944 585
R153 gnd.n944 gnd.n943 585
R154 gnd.n5544 gnd.n5543 585
R155 gnd.n5543 gnd.n5542 585
R156 gnd.n950 gnd.n949 585
R157 gnd.n5541 gnd.n950 585
R158 gnd.n5539 gnd.n5538 585
R159 gnd.n5540 gnd.n5539 585
R160 gnd.n5537 gnd.n952 585
R161 gnd.n952 gnd.n951 585
R162 gnd.n5536 gnd.n5535 585
R163 gnd.n5535 gnd.n5534 585
R164 gnd.n958 gnd.n957 585
R165 gnd.n5533 gnd.n958 585
R166 gnd.n5531 gnd.n5530 585
R167 gnd.n5532 gnd.n5531 585
R168 gnd.n5529 gnd.n960 585
R169 gnd.n960 gnd.n959 585
R170 gnd.n5528 gnd.n5527 585
R171 gnd.n5527 gnd.n5526 585
R172 gnd.n966 gnd.n965 585
R173 gnd.n5525 gnd.n966 585
R174 gnd.n5523 gnd.n5522 585
R175 gnd.n5524 gnd.n5523 585
R176 gnd.n5521 gnd.n968 585
R177 gnd.n968 gnd.n967 585
R178 gnd.n5520 gnd.n5519 585
R179 gnd.n5519 gnd.n5518 585
R180 gnd.n974 gnd.n973 585
R181 gnd.n5517 gnd.n974 585
R182 gnd.n5515 gnd.n5514 585
R183 gnd.n5516 gnd.n5515 585
R184 gnd.n5513 gnd.n976 585
R185 gnd.n976 gnd.n975 585
R186 gnd.n5512 gnd.n5511 585
R187 gnd.n5511 gnd.n5510 585
R188 gnd.n982 gnd.n981 585
R189 gnd.n5509 gnd.n982 585
R190 gnd.n5507 gnd.n5506 585
R191 gnd.n5508 gnd.n5507 585
R192 gnd.n5505 gnd.n984 585
R193 gnd.n984 gnd.n983 585
R194 gnd.n5504 gnd.n5503 585
R195 gnd.n5503 gnd.n5502 585
R196 gnd.n990 gnd.n989 585
R197 gnd.n5501 gnd.n990 585
R198 gnd.n5499 gnd.n5498 585
R199 gnd.n5500 gnd.n5499 585
R200 gnd.n5497 gnd.n992 585
R201 gnd.n992 gnd.n991 585
R202 gnd.n828 gnd.n827 585
R203 gnd.n827 gnd.n826 585
R204 gnd.n5669 gnd.n5668 585
R205 gnd.n5670 gnd.n5669 585
R206 gnd.n825 gnd.n824 585
R207 gnd.n5671 gnd.n825 585
R208 gnd.n5674 gnd.n5673 585
R209 gnd.n5673 gnd.n5672 585
R210 gnd.n822 gnd.n821 585
R211 gnd.n821 gnd.n820 585
R212 gnd.n5679 gnd.n5678 585
R213 gnd.n5680 gnd.n5679 585
R214 gnd.n819 gnd.n818 585
R215 gnd.n5681 gnd.n819 585
R216 gnd.n5684 gnd.n5683 585
R217 gnd.n5683 gnd.n5682 585
R218 gnd.n816 gnd.n815 585
R219 gnd.n815 gnd.n814 585
R220 gnd.n5689 gnd.n5688 585
R221 gnd.n5690 gnd.n5689 585
R222 gnd.n813 gnd.n812 585
R223 gnd.n5691 gnd.n813 585
R224 gnd.n5694 gnd.n5693 585
R225 gnd.n5693 gnd.n5692 585
R226 gnd.n810 gnd.n809 585
R227 gnd.n809 gnd.n808 585
R228 gnd.n5699 gnd.n5698 585
R229 gnd.n5700 gnd.n5699 585
R230 gnd.n807 gnd.n806 585
R231 gnd.n5701 gnd.n807 585
R232 gnd.n5704 gnd.n5703 585
R233 gnd.n5703 gnd.n5702 585
R234 gnd.n804 gnd.n803 585
R235 gnd.n803 gnd.n802 585
R236 gnd.n5709 gnd.n5708 585
R237 gnd.n5710 gnd.n5709 585
R238 gnd.n801 gnd.n800 585
R239 gnd.n5711 gnd.n801 585
R240 gnd.n5714 gnd.n5713 585
R241 gnd.n5713 gnd.n5712 585
R242 gnd.n798 gnd.n797 585
R243 gnd.n797 gnd.n796 585
R244 gnd.n5719 gnd.n5718 585
R245 gnd.n5720 gnd.n5719 585
R246 gnd.n795 gnd.n794 585
R247 gnd.n5721 gnd.n795 585
R248 gnd.n5724 gnd.n5723 585
R249 gnd.n5723 gnd.n5722 585
R250 gnd.n792 gnd.n791 585
R251 gnd.n791 gnd.n790 585
R252 gnd.n5729 gnd.n5728 585
R253 gnd.n5730 gnd.n5729 585
R254 gnd.n789 gnd.n788 585
R255 gnd.n5731 gnd.n789 585
R256 gnd.n5734 gnd.n5733 585
R257 gnd.n5733 gnd.n5732 585
R258 gnd.n786 gnd.n785 585
R259 gnd.n785 gnd.n784 585
R260 gnd.n5739 gnd.n5738 585
R261 gnd.n5740 gnd.n5739 585
R262 gnd.n783 gnd.n782 585
R263 gnd.n5741 gnd.n783 585
R264 gnd.n5744 gnd.n5743 585
R265 gnd.n5743 gnd.n5742 585
R266 gnd.n780 gnd.n779 585
R267 gnd.n779 gnd.n778 585
R268 gnd.n5749 gnd.n5748 585
R269 gnd.n5750 gnd.n5749 585
R270 gnd.n777 gnd.n776 585
R271 gnd.n5751 gnd.n777 585
R272 gnd.n5754 gnd.n5753 585
R273 gnd.n5753 gnd.n5752 585
R274 gnd.n774 gnd.n773 585
R275 gnd.n773 gnd.n772 585
R276 gnd.n5759 gnd.n5758 585
R277 gnd.n5760 gnd.n5759 585
R278 gnd.n771 gnd.n770 585
R279 gnd.n5761 gnd.n771 585
R280 gnd.n5764 gnd.n5763 585
R281 gnd.n5763 gnd.n5762 585
R282 gnd.n768 gnd.n767 585
R283 gnd.n767 gnd.n766 585
R284 gnd.n5769 gnd.n5768 585
R285 gnd.n5770 gnd.n5769 585
R286 gnd.n765 gnd.n764 585
R287 gnd.n5771 gnd.n765 585
R288 gnd.n5774 gnd.n5773 585
R289 gnd.n5773 gnd.n5772 585
R290 gnd.n762 gnd.n761 585
R291 gnd.n761 gnd.n760 585
R292 gnd.n5779 gnd.n5778 585
R293 gnd.n5780 gnd.n5779 585
R294 gnd.n759 gnd.n758 585
R295 gnd.n5781 gnd.n759 585
R296 gnd.n5784 gnd.n5783 585
R297 gnd.n5783 gnd.n5782 585
R298 gnd.n756 gnd.n755 585
R299 gnd.n755 gnd.n754 585
R300 gnd.n5789 gnd.n5788 585
R301 gnd.n5790 gnd.n5789 585
R302 gnd.n753 gnd.n752 585
R303 gnd.n5791 gnd.n753 585
R304 gnd.n5794 gnd.n5793 585
R305 gnd.n5793 gnd.n5792 585
R306 gnd.n750 gnd.n749 585
R307 gnd.n749 gnd.n748 585
R308 gnd.n5799 gnd.n5798 585
R309 gnd.n5800 gnd.n5799 585
R310 gnd.n747 gnd.n746 585
R311 gnd.n5801 gnd.n747 585
R312 gnd.n5804 gnd.n5803 585
R313 gnd.n5803 gnd.n5802 585
R314 gnd.n744 gnd.n743 585
R315 gnd.n743 gnd.n742 585
R316 gnd.n5809 gnd.n5808 585
R317 gnd.n5810 gnd.n5809 585
R318 gnd.n741 gnd.n740 585
R319 gnd.n5811 gnd.n741 585
R320 gnd.n5814 gnd.n5813 585
R321 gnd.n5813 gnd.n5812 585
R322 gnd.n738 gnd.n737 585
R323 gnd.n737 gnd.n736 585
R324 gnd.n5819 gnd.n5818 585
R325 gnd.n5820 gnd.n5819 585
R326 gnd.n735 gnd.n734 585
R327 gnd.n5821 gnd.n735 585
R328 gnd.n5824 gnd.n5823 585
R329 gnd.n5823 gnd.n5822 585
R330 gnd.n732 gnd.n731 585
R331 gnd.n731 gnd.n730 585
R332 gnd.n5829 gnd.n5828 585
R333 gnd.n5830 gnd.n5829 585
R334 gnd.n729 gnd.n728 585
R335 gnd.n5831 gnd.n729 585
R336 gnd.n5834 gnd.n5833 585
R337 gnd.n5833 gnd.n5832 585
R338 gnd.n726 gnd.n725 585
R339 gnd.n725 gnd.n724 585
R340 gnd.n5839 gnd.n5838 585
R341 gnd.n5840 gnd.n5839 585
R342 gnd.n723 gnd.n722 585
R343 gnd.n5841 gnd.n723 585
R344 gnd.n5844 gnd.n5843 585
R345 gnd.n5843 gnd.n5842 585
R346 gnd.n720 gnd.n719 585
R347 gnd.n719 gnd.n718 585
R348 gnd.n5849 gnd.n5848 585
R349 gnd.n5850 gnd.n5849 585
R350 gnd.n717 gnd.n716 585
R351 gnd.n5851 gnd.n717 585
R352 gnd.n5854 gnd.n5853 585
R353 gnd.n5853 gnd.n5852 585
R354 gnd.n714 gnd.n713 585
R355 gnd.n713 gnd.n712 585
R356 gnd.n5859 gnd.n5858 585
R357 gnd.n5860 gnd.n5859 585
R358 gnd.n711 gnd.n710 585
R359 gnd.n5861 gnd.n711 585
R360 gnd.n5864 gnd.n5863 585
R361 gnd.n5863 gnd.n5862 585
R362 gnd.n708 gnd.n707 585
R363 gnd.n707 gnd.n706 585
R364 gnd.n5869 gnd.n5868 585
R365 gnd.n5870 gnd.n5869 585
R366 gnd.n705 gnd.n704 585
R367 gnd.n5871 gnd.n705 585
R368 gnd.n5874 gnd.n5873 585
R369 gnd.n5873 gnd.n5872 585
R370 gnd.n702 gnd.n701 585
R371 gnd.n701 gnd.n700 585
R372 gnd.n5879 gnd.n5878 585
R373 gnd.n5880 gnd.n5879 585
R374 gnd.n699 gnd.n698 585
R375 gnd.n5881 gnd.n699 585
R376 gnd.n5884 gnd.n5883 585
R377 gnd.n5883 gnd.n5882 585
R378 gnd.n696 gnd.n695 585
R379 gnd.n695 gnd.n694 585
R380 gnd.n5889 gnd.n5888 585
R381 gnd.n5890 gnd.n5889 585
R382 gnd.n693 gnd.n692 585
R383 gnd.n5891 gnd.n693 585
R384 gnd.n5894 gnd.n5893 585
R385 gnd.n5893 gnd.n5892 585
R386 gnd.n690 gnd.n689 585
R387 gnd.n689 gnd.n688 585
R388 gnd.n5899 gnd.n5898 585
R389 gnd.n5900 gnd.n5899 585
R390 gnd.n687 gnd.n686 585
R391 gnd.n5901 gnd.n687 585
R392 gnd.n5904 gnd.n5903 585
R393 gnd.n5903 gnd.n5902 585
R394 gnd.n684 gnd.n683 585
R395 gnd.n683 gnd.n682 585
R396 gnd.n5909 gnd.n5908 585
R397 gnd.n5910 gnd.n5909 585
R398 gnd.n681 gnd.n680 585
R399 gnd.n5911 gnd.n681 585
R400 gnd.n5914 gnd.n5913 585
R401 gnd.n5913 gnd.n5912 585
R402 gnd.n678 gnd.n677 585
R403 gnd.n677 gnd.n676 585
R404 gnd.n5919 gnd.n5918 585
R405 gnd.n5920 gnd.n5919 585
R406 gnd.n675 gnd.n674 585
R407 gnd.n5921 gnd.n675 585
R408 gnd.n5924 gnd.n5923 585
R409 gnd.n5923 gnd.n5922 585
R410 gnd.n672 gnd.n671 585
R411 gnd.n671 gnd.n670 585
R412 gnd.n5929 gnd.n5928 585
R413 gnd.n5930 gnd.n5929 585
R414 gnd.n669 gnd.n668 585
R415 gnd.n5931 gnd.n669 585
R416 gnd.n5934 gnd.n5933 585
R417 gnd.n5933 gnd.n5932 585
R418 gnd.n666 gnd.n665 585
R419 gnd.n665 gnd.n664 585
R420 gnd.n5939 gnd.n5938 585
R421 gnd.n5940 gnd.n5939 585
R422 gnd.n663 gnd.n662 585
R423 gnd.n5941 gnd.n663 585
R424 gnd.n5944 gnd.n5943 585
R425 gnd.n5943 gnd.n5942 585
R426 gnd.n660 gnd.n659 585
R427 gnd.n659 gnd.n658 585
R428 gnd.n5949 gnd.n5948 585
R429 gnd.n5950 gnd.n5949 585
R430 gnd.n657 gnd.n656 585
R431 gnd.n5951 gnd.n657 585
R432 gnd.n5954 gnd.n5953 585
R433 gnd.n5953 gnd.n5952 585
R434 gnd.n654 gnd.n653 585
R435 gnd.n653 gnd.n652 585
R436 gnd.n5959 gnd.n5958 585
R437 gnd.n5960 gnd.n5959 585
R438 gnd.n651 gnd.n650 585
R439 gnd.n5961 gnd.n651 585
R440 gnd.n5964 gnd.n5963 585
R441 gnd.n5963 gnd.n5962 585
R442 gnd.n648 gnd.n647 585
R443 gnd.n647 gnd.n646 585
R444 gnd.n5969 gnd.n5968 585
R445 gnd.n5970 gnd.n5969 585
R446 gnd.n645 gnd.n644 585
R447 gnd.n5971 gnd.n645 585
R448 gnd.n5974 gnd.n5973 585
R449 gnd.n5973 gnd.n5972 585
R450 gnd.n642 gnd.n641 585
R451 gnd.n641 gnd.n640 585
R452 gnd.n5980 gnd.n5979 585
R453 gnd.n5981 gnd.n5980 585
R454 gnd.n639 gnd.n638 585
R455 gnd.n5982 gnd.n639 585
R456 gnd.n5985 gnd.n5984 585
R457 gnd.n5984 gnd.n5983 585
R458 gnd.n5986 gnd.n636 585
R459 gnd.n636 gnd.n635 585
R460 gnd.n511 gnd.n510 585
R461 gnd.n6193 gnd.n510 585
R462 gnd.n6196 gnd.n6195 585
R463 gnd.n6195 gnd.n6194 585
R464 gnd.n514 gnd.n513 585
R465 gnd.n6192 gnd.n514 585
R466 gnd.n6190 gnd.n6189 585
R467 gnd.n6191 gnd.n6190 585
R468 gnd.n517 gnd.n516 585
R469 gnd.n516 gnd.n515 585
R470 gnd.n6185 gnd.n6184 585
R471 gnd.n6184 gnd.n6183 585
R472 gnd.n520 gnd.n519 585
R473 gnd.n6182 gnd.n520 585
R474 gnd.n6180 gnd.n6179 585
R475 gnd.n6181 gnd.n6180 585
R476 gnd.n523 gnd.n522 585
R477 gnd.n522 gnd.n521 585
R478 gnd.n6175 gnd.n6174 585
R479 gnd.n6174 gnd.n6173 585
R480 gnd.n526 gnd.n525 585
R481 gnd.n6172 gnd.n526 585
R482 gnd.n6170 gnd.n6169 585
R483 gnd.n6171 gnd.n6170 585
R484 gnd.n529 gnd.n528 585
R485 gnd.n528 gnd.n527 585
R486 gnd.n6165 gnd.n6164 585
R487 gnd.n6164 gnd.n6163 585
R488 gnd.n532 gnd.n531 585
R489 gnd.n6162 gnd.n532 585
R490 gnd.n6160 gnd.n6159 585
R491 gnd.n6161 gnd.n6160 585
R492 gnd.n535 gnd.n534 585
R493 gnd.n534 gnd.n533 585
R494 gnd.n6155 gnd.n6154 585
R495 gnd.n6154 gnd.n6153 585
R496 gnd.n538 gnd.n537 585
R497 gnd.n6152 gnd.n538 585
R498 gnd.n6150 gnd.n6149 585
R499 gnd.n6151 gnd.n6150 585
R500 gnd.n541 gnd.n540 585
R501 gnd.n540 gnd.n539 585
R502 gnd.n6145 gnd.n6144 585
R503 gnd.n6144 gnd.n6143 585
R504 gnd.n544 gnd.n543 585
R505 gnd.n6142 gnd.n544 585
R506 gnd.n6140 gnd.n6139 585
R507 gnd.n6141 gnd.n6140 585
R508 gnd.n547 gnd.n546 585
R509 gnd.n546 gnd.n545 585
R510 gnd.n6135 gnd.n6134 585
R511 gnd.n6134 gnd.n6133 585
R512 gnd.n550 gnd.n549 585
R513 gnd.n6132 gnd.n550 585
R514 gnd.n6130 gnd.n6129 585
R515 gnd.n6131 gnd.n6130 585
R516 gnd.n553 gnd.n552 585
R517 gnd.n552 gnd.n551 585
R518 gnd.n6125 gnd.n6124 585
R519 gnd.n6124 gnd.n6123 585
R520 gnd.n556 gnd.n555 585
R521 gnd.n6122 gnd.n556 585
R522 gnd.n6120 gnd.n6119 585
R523 gnd.n6121 gnd.n6120 585
R524 gnd.n559 gnd.n558 585
R525 gnd.n558 gnd.n557 585
R526 gnd.n6115 gnd.n6114 585
R527 gnd.n6114 gnd.n6113 585
R528 gnd.n562 gnd.n561 585
R529 gnd.n6112 gnd.n562 585
R530 gnd.n6110 gnd.n6109 585
R531 gnd.n6111 gnd.n6110 585
R532 gnd.n565 gnd.n564 585
R533 gnd.n564 gnd.n563 585
R534 gnd.n6105 gnd.n6104 585
R535 gnd.n6104 gnd.n6103 585
R536 gnd.n568 gnd.n567 585
R537 gnd.n6102 gnd.n568 585
R538 gnd.n6100 gnd.n6099 585
R539 gnd.n6101 gnd.n6100 585
R540 gnd.n571 gnd.n570 585
R541 gnd.n570 gnd.n569 585
R542 gnd.n6095 gnd.n6094 585
R543 gnd.n6094 gnd.n6093 585
R544 gnd.n574 gnd.n573 585
R545 gnd.n6092 gnd.n574 585
R546 gnd.n6090 gnd.n6089 585
R547 gnd.n6091 gnd.n6090 585
R548 gnd.n577 gnd.n576 585
R549 gnd.n576 gnd.n575 585
R550 gnd.n6085 gnd.n6084 585
R551 gnd.n6084 gnd.n6083 585
R552 gnd.n580 gnd.n579 585
R553 gnd.n6082 gnd.n580 585
R554 gnd.n6080 gnd.n6079 585
R555 gnd.n6081 gnd.n6080 585
R556 gnd.n583 gnd.n582 585
R557 gnd.n582 gnd.n581 585
R558 gnd.n6075 gnd.n6074 585
R559 gnd.n6074 gnd.n6073 585
R560 gnd.n586 gnd.n585 585
R561 gnd.n6072 gnd.n586 585
R562 gnd.n6070 gnd.n6069 585
R563 gnd.n6071 gnd.n6070 585
R564 gnd.n589 gnd.n588 585
R565 gnd.n588 gnd.n587 585
R566 gnd.n6065 gnd.n6064 585
R567 gnd.n6064 gnd.n6063 585
R568 gnd.n592 gnd.n591 585
R569 gnd.n6062 gnd.n592 585
R570 gnd.n6060 gnd.n6059 585
R571 gnd.n6061 gnd.n6060 585
R572 gnd.n595 gnd.n594 585
R573 gnd.n594 gnd.n593 585
R574 gnd.n6055 gnd.n6054 585
R575 gnd.n6054 gnd.n6053 585
R576 gnd.n598 gnd.n597 585
R577 gnd.n6052 gnd.n598 585
R578 gnd.n6050 gnd.n6049 585
R579 gnd.n6051 gnd.n6050 585
R580 gnd.n601 gnd.n600 585
R581 gnd.n600 gnd.n599 585
R582 gnd.n6045 gnd.n6044 585
R583 gnd.n6044 gnd.n6043 585
R584 gnd.n604 gnd.n603 585
R585 gnd.n6042 gnd.n604 585
R586 gnd.n6040 gnd.n6039 585
R587 gnd.n6041 gnd.n6040 585
R588 gnd.n607 gnd.n606 585
R589 gnd.n606 gnd.n605 585
R590 gnd.n6035 gnd.n6034 585
R591 gnd.n6034 gnd.n6033 585
R592 gnd.n610 gnd.n609 585
R593 gnd.n6032 gnd.n610 585
R594 gnd.n6030 gnd.n6029 585
R595 gnd.n6031 gnd.n6030 585
R596 gnd.n613 gnd.n612 585
R597 gnd.n612 gnd.n611 585
R598 gnd.n6025 gnd.n6024 585
R599 gnd.n6024 gnd.n6023 585
R600 gnd.n616 gnd.n615 585
R601 gnd.n6022 gnd.n616 585
R602 gnd.n6020 gnd.n6019 585
R603 gnd.n6021 gnd.n6020 585
R604 gnd.n619 gnd.n618 585
R605 gnd.n618 gnd.n617 585
R606 gnd.n6015 gnd.n6014 585
R607 gnd.n6014 gnd.n6013 585
R608 gnd.n622 gnd.n621 585
R609 gnd.n6012 gnd.n622 585
R610 gnd.n6010 gnd.n6009 585
R611 gnd.n6011 gnd.n6010 585
R612 gnd.n625 gnd.n624 585
R613 gnd.n624 gnd.n623 585
R614 gnd.n6005 gnd.n6004 585
R615 gnd.n6004 gnd.n6003 585
R616 gnd.n628 gnd.n627 585
R617 gnd.n6002 gnd.n628 585
R618 gnd.n6000 gnd.n5999 585
R619 gnd.n6001 gnd.n6000 585
R620 gnd.n631 gnd.n630 585
R621 gnd.n630 gnd.n629 585
R622 gnd.n5995 gnd.n5994 585
R623 gnd.n5994 gnd.n5993 585
R624 gnd.n634 gnd.n633 585
R625 gnd.n5992 gnd.n634 585
R626 gnd.n5990 gnd.n5989 585
R627 gnd.n5991 gnd.n5990 585
R628 gnd.n1084 gnd.n1083 585
R629 gnd.n4186 gnd.n1084 585
R630 gnd.n5447 gnd.n5446 585
R631 gnd.n5446 gnd.n5445 585
R632 gnd.n5448 gnd.n1078 585
R633 gnd.n4149 gnd.n1078 585
R634 gnd.n5450 gnd.n5449 585
R635 gnd.n5451 gnd.n5450 585
R636 gnd.n1062 gnd.n1061 585
R637 gnd.n4073 gnd.n1062 585
R638 gnd.n5459 gnd.n5458 585
R639 gnd.n5458 gnd.n5457 585
R640 gnd.n5460 gnd.n1056 585
R641 gnd.n4162 gnd.n1056 585
R642 gnd.n5462 gnd.n5461 585
R643 gnd.n5463 gnd.n5462 585
R644 gnd.n1042 gnd.n1041 585
R645 gnd.n4065 gnd.n1042 585
R646 gnd.n5471 gnd.n5470 585
R647 gnd.n5470 gnd.n5469 585
R648 gnd.n5472 gnd.n1036 585
R649 gnd.n4057 gnd.n1036 585
R650 gnd.n5474 gnd.n5473 585
R651 gnd.n5475 gnd.n5474 585
R652 gnd.n1020 gnd.n1019 585
R653 gnd.n4022 gnd.n1020 585
R654 gnd.n5483 gnd.n5482 585
R655 gnd.n5482 gnd.n5481 585
R656 gnd.n5484 gnd.n1014 585
R657 gnd.n4030 gnd.n1014 585
R658 gnd.n5486 gnd.n5485 585
R659 gnd.n5487 gnd.n5486 585
R660 gnd.n1015 gnd.n1013 585
R661 gnd.n4008 gnd.n1013 585
R662 gnd.n3984 gnd.n1002 585
R663 gnd.n5493 gnd.n1002 585
R664 gnd.n3986 gnd.n3985 585
R665 gnd.n3985 gnd.n998 585
R666 gnd.n3987 gnd.n2025 585
R667 gnd.n3999 gnd.n2025 585
R668 gnd.n3988 gnd.n2034 585
R669 gnd.n2034 gnd.n2032 585
R670 gnd.n3990 gnd.n3989 585
R671 gnd.n3991 gnd.n3990 585
R672 gnd.n2035 gnd.n2033 585
R673 gnd.n2033 gnd.n2029 585
R674 gnd.n3952 gnd.n2043 585
R675 gnd.n3964 gnd.n2043 585
R676 gnd.n3953 gnd.n2051 585
R677 gnd.n2051 gnd.n2041 585
R678 gnd.n3955 gnd.n3954 585
R679 gnd.n3956 gnd.n3955 585
R680 gnd.n2052 gnd.n2050 585
R681 gnd.n2050 gnd.n2047 585
R682 gnd.n3946 gnd.n3945 585
R683 gnd.n3945 gnd.n3944 585
R684 gnd.n2055 gnd.n2054 585
R685 gnd.n2066 gnd.n2055 585
R686 gnd.n3934 gnd.n3933 585
R687 gnd.n3935 gnd.n3934 585
R688 gnd.n2068 gnd.n2067 585
R689 gnd.n2067 gnd.n2063 585
R690 gnd.n3929 gnd.n3928 585
R691 gnd.n3928 gnd.n3927 585
R692 gnd.n2071 gnd.n2070 585
R693 gnd.n2072 gnd.n2071 585
R694 gnd.n3918 gnd.n3917 585
R695 gnd.n3919 gnd.n3918 585
R696 gnd.n2084 gnd.n2083 585
R697 gnd.n2083 gnd.n2080 585
R698 gnd.n3913 gnd.n3912 585
R699 gnd.n3912 gnd.n3911 585
R700 gnd.n2087 gnd.n2086 585
R701 gnd.n2098 gnd.n2087 585
R702 gnd.n3902 gnd.n3901 585
R703 gnd.n3903 gnd.n3902 585
R704 gnd.n2100 gnd.n2099 585
R705 gnd.n2099 gnd.n2095 585
R706 gnd.n3897 gnd.n3896 585
R707 gnd.n3896 gnd.n3895 585
R708 gnd.n2103 gnd.n2102 585
R709 gnd.n2104 gnd.n2103 585
R710 gnd.n3886 gnd.n3885 585
R711 gnd.n3887 gnd.n3886 585
R712 gnd.n2116 gnd.n2115 585
R713 gnd.n2115 gnd.n2112 585
R714 gnd.n3881 gnd.n3880 585
R715 gnd.n2119 gnd.n2118 585
R716 gnd.n3611 gnd.n3610 585
R717 gnd.n3613 gnd.n3612 585
R718 gnd.n3615 gnd.n3614 585
R719 gnd.n3619 gnd.n3607 585
R720 gnd.n3621 gnd.n3620 585
R721 gnd.n3623 gnd.n3622 585
R722 gnd.n3625 gnd.n3624 585
R723 gnd.n3629 gnd.n3605 585
R724 gnd.n3631 gnd.n3630 585
R725 gnd.n3633 gnd.n3632 585
R726 gnd.n3635 gnd.n3634 585
R727 gnd.n3639 gnd.n3603 585
R728 gnd.n3641 gnd.n3640 585
R729 gnd.n3643 gnd.n3642 585
R730 gnd.n3645 gnd.n3644 585
R731 gnd.n3601 gnd.n3597 585
R732 gnd.n3706 gnd.n3705 585
R733 gnd.n3878 gnd.n3706 585
R734 gnd.n4189 gnd.n4188 585
R735 gnd.n1979 gnd.n1978 585
R736 gnd.n1977 gnd.n1974 585
R737 gnd.n1962 gnd.n1880 585
R738 gnd.n1964 gnd.n1963 585
R739 gnd.n1961 gnd.n1886 585
R740 gnd.n1885 gnd.n1884 585
R741 gnd.n1952 gnd.n1951 585
R742 gnd.n1950 gnd.n1949 585
R743 gnd.n1938 gnd.n1892 585
R744 gnd.n1940 gnd.n1939 585
R745 gnd.n1937 gnd.n1898 585
R746 gnd.n1897 gnd.n1896 585
R747 gnd.n1928 gnd.n1927 585
R748 gnd.n1926 gnd.n1925 585
R749 gnd.n1914 gnd.n1904 585
R750 gnd.n1916 gnd.n1915 585
R751 gnd.n1913 gnd.n1911 585
R752 gnd.n1910 gnd.n1096 585
R753 gnd.n5437 gnd.n1096 585
R754 gnd.n4187 gnd.n1980 585
R755 gnd.n4187 gnd.n4186 585
R756 gnd.n4151 gnd.n1087 585
R757 gnd.n5445 gnd.n1087 585
R758 gnd.n4154 gnd.n4150 585
R759 gnd.n4150 gnd.n4149 585
R760 gnd.n4155 gnd.n1076 585
R761 gnd.n5451 gnd.n1076 585
R762 gnd.n4156 gnd.n1997 585
R763 gnd.n4073 gnd.n1997 585
R764 gnd.n1994 gnd.n1065 585
R765 gnd.n5457 gnd.n1065 585
R766 gnd.n4161 gnd.n4160 585
R767 gnd.n4162 gnd.n4161 585
R768 gnd.n1993 gnd.n1055 585
R769 gnd.n5463 gnd.n1055 585
R770 gnd.n4064 gnd.n4063 585
R771 gnd.n4065 gnd.n4064 585
R772 gnd.n2003 gnd.n1044 585
R773 gnd.n5469 gnd.n1044 585
R774 gnd.n4059 gnd.n4058 585
R775 gnd.n4058 gnd.n4057 585
R776 gnd.n2005 gnd.n1034 585
R777 gnd.n5475 gnd.n1034 585
R778 gnd.n4024 gnd.n4023 585
R779 gnd.n4023 gnd.n4022 585
R780 gnd.n2014 gnd.n1023 585
R781 gnd.n5481 gnd.n1023 585
R782 gnd.n4029 gnd.n4028 585
R783 gnd.n4030 gnd.n4029 585
R784 gnd.n2013 gnd.n1012 585
R785 gnd.n5487 gnd.n1012 585
R786 gnd.n4007 gnd.n4006 585
R787 gnd.n4008 gnd.n4007 585
R788 gnd.n2020 gnd.n1000 585
R789 gnd.n5493 gnd.n1000 585
R790 gnd.n4002 gnd.n4001 585
R791 gnd.n4001 gnd.n998 585
R792 gnd.n4000 gnd.n2022 585
R793 gnd.n4000 gnd.n3999 585
R794 gnd.n3668 gnd.n2023 585
R795 gnd.n2032 gnd.n2023 585
R796 gnd.n3671 gnd.n2031 585
R797 gnd.n3991 gnd.n2031 585
R798 gnd.n3673 gnd.n3672 585
R799 gnd.n3672 gnd.n2029 585
R800 gnd.n3674 gnd.n2042 585
R801 gnd.n3964 gnd.n2042 585
R802 gnd.n3676 gnd.n3675 585
R803 gnd.n3675 gnd.n2041 585
R804 gnd.n3677 gnd.n2049 585
R805 gnd.n3956 gnd.n2049 585
R806 gnd.n3679 gnd.n3678 585
R807 gnd.n3678 gnd.n2047 585
R808 gnd.n3680 gnd.n2057 585
R809 gnd.n3944 gnd.n2057 585
R810 gnd.n3682 gnd.n3681 585
R811 gnd.n3681 gnd.n2066 585
R812 gnd.n3683 gnd.n2065 585
R813 gnd.n3935 gnd.n2065 585
R814 gnd.n3685 gnd.n3684 585
R815 gnd.n3684 gnd.n2063 585
R816 gnd.n3686 gnd.n2074 585
R817 gnd.n3927 gnd.n2074 585
R818 gnd.n3688 gnd.n3687 585
R819 gnd.n3687 gnd.n2072 585
R820 gnd.n3689 gnd.n2082 585
R821 gnd.n3919 gnd.n2082 585
R822 gnd.n3691 gnd.n3690 585
R823 gnd.n3690 gnd.n2080 585
R824 gnd.n3692 gnd.n2089 585
R825 gnd.n3911 gnd.n2089 585
R826 gnd.n3694 gnd.n3693 585
R827 gnd.n3693 gnd.n2098 585
R828 gnd.n3695 gnd.n2097 585
R829 gnd.n3903 gnd.n2097 585
R830 gnd.n3697 gnd.n3696 585
R831 gnd.n3696 gnd.n2095 585
R832 gnd.n3698 gnd.n2106 585
R833 gnd.n3895 gnd.n2106 585
R834 gnd.n3700 gnd.n3699 585
R835 gnd.n3699 gnd.n2104 585
R836 gnd.n3701 gnd.n2114 585
R837 gnd.n3887 gnd.n2114 585
R838 gnd.n3702 gnd.n3598 585
R839 gnd.n3598 gnd.n2112 585
R840 gnd.n6668 gnd.n84 585
R841 gnd.n6764 gnd.n84 585
R842 gnd.n6669 gnd.n6600 585
R843 gnd.n6600 gnd.n81 585
R844 gnd.n6670 gnd.n162 585
R845 gnd.n6684 gnd.n162 585
R846 gnd.n174 gnd.n172 585
R847 gnd.n172 gnd.n161 585
R848 gnd.n6675 gnd.n6674 585
R849 gnd.n6676 gnd.n6675 585
R850 gnd.n173 gnd.n171 585
R851 gnd.n171 gnd.n169 585
R852 gnd.n6596 gnd.n6595 585
R853 gnd.n6595 gnd.n6594 585
R854 gnd.n177 gnd.n176 585
R855 gnd.n188 gnd.n177 585
R856 gnd.n6585 gnd.n6584 585
R857 gnd.n6586 gnd.n6585 585
R858 gnd.n190 gnd.n189 585
R859 gnd.n189 gnd.n186 585
R860 gnd.n6580 gnd.n6579 585
R861 gnd.n6579 gnd.n6578 585
R862 gnd.n193 gnd.n192 585
R863 gnd.n194 gnd.n193 585
R864 gnd.n6569 gnd.n6568 585
R865 gnd.n6570 gnd.n6569 585
R866 gnd.n205 gnd.n204 585
R867 gnd.n204 gnd.n202 585
R868 gnd.n6564 gnd.n6563 585
R869 gnd.n6563 gnd.n6562 585
R870 gnd.n208 gnd.n207 585
R871 gnd.n224 gnd.n208 585
R872 gnd.n6553 gnd.n6552 585
R873 gnd.n6554 gnd.n6553 585
R874 gnd.n226 gnd.n225 585
R875 gnd.n225 gnd.n222 585
R876 gnd.n6548 gnd.n6547 585
R877 gnd.n6547 gnd.n6546 585
R878 gnd.n229 gnd.n228 585
R879 gnd.n230 gnd.n229 585
R880 gnd.n6539 gnd.n6538 585
R881 gnd.n6540 gnd.n6539 585
R882 gnd.n238 gnd.n237 585
R883 gnd.n237 gnd.n235 585
R884 gnd.n6534 gnd.n6533 585
R885 gnd.n6533 gnd.n6532 585
R886 gnd.n242 gnd.n241 585
R887 gnd.n6527 gnd.n242 585
R888 gnd.n6508 gnd.n6507 585
R889 gnd.n6507 gnd.n247 585
R890 gnd.n264 gnd.n257 585
R891 gnd.n6519 gnd.n257 585
R892 gnd.n6513 gnd.n6512 585
R893 gnd.n6514 gnd.n6513 585
R894 gnd.n263 gnd.n262 585
R895 gnd.n6287 gnd.n262 585
R896 gnd.n6504 gnd.n6503 585
R897 gnd.n6503 gnd.n6502 585
R898 gnd.n267 gnd.n266 585
R899 gnd.n6221 gnd.n267 585
R900 gnd.n6492 gnd.n6491 585
R901 gnd.n6493 gnd.n6492 585
R902 gnd.n281 gnd.n280 585
R903 gnd.n6217 gnd.n280 585
R904 gnd.n6487 gnd.n6486 585
R905 gnd.n6486 gnd.n6485 585
R906 gnd.n284 gnd.n283 585
R907 gnd.n497 gnd.n284 585
R908 gnd.n6476 gnd.n6475 585
R909 gnd.n6477 gnd.n6476 585
R910 gnd.n299 gnd.n298 585
R911 gnd.n493 gnd.n298 585
R912 gnd.n6471 gnd.n6470 585
R913 gnd.n6470 gnd.n6469 585
R914 gnd.n302 gnd.n301 585
R915 gnd.n487 gnd.n302 585
R916 gnd.n6460 gnd.n6459 585
R917 gnd.n6461 gnd.n6460 585
R918 gnd.n317 gnd.n316 585
R919 gnd.n6310 gnd.n316 585
R920 gnd.n6455 gnd.n6454 585
R921 gnd.n6454 gnd.n6453 585
R922 gnd.n320 gnd.n319 585
R923 gnd.n5150 gnd.n320 585
R924 gnd.n6444 gnd.n6443 585
R925 gnd.n6445 gnd.n6444 585
R926 gnd.n6440 gnd.n332 585
R927 gnd.n6439 gnd.n334 585
R928 gnd.n404 gnd.n335 585
R929 gnd.n6432 gnd.n341 585
R930 gnd.n6431 gnd.n342 585
R931 gnd.n406 gnd.n343 585
R932 gnd.n6424 gnd.n349 585
R933 gnd.n6423 gnd.n350 585
R934 gnd.n409 gnd.n351 585
R935 gnd.n6416 gnd.n357 585
R936 gnd.n6415 gnd.n358 585
R937 gnd.n411 gnd.n359 585
R938 gnd.n6408 gnd.n365 585
R939 gnd.n6407 gnd.n366 585
R940 gnd.n414 gnd.n367 585
R941 gnd.n6400 gnd.n373 585
R942 gnd.n6399 gnd.n374 585
R943 gnd.n383 gnd.n377 585
R944 gnd.n6392 gnd.n6391 585
R945 gnd.n6391 gnd.n6390 585
R946 gnd.n6639 gnd.n80 585
R947 gnd.n6640 gnd.n6638 585
R948 gnd.n6641 gnd.n6634 585
R949 gnd.n6632 gnd.n6630 585
R950 gnd.n6645 gnd.n6629 585
R951 gnd.n6646 gnd.n6627 585
R952 gnd.n6647 gnd.n6626 585
R953 gnd.n6624 gnd.n6622 585
R954 gnd.n6651 gnd.n6621 585
R955 gnd.n6652 gnd.n6619 585
R956 gnd.n6653 gnd.n6618 585
R957 gnd.n6616 gnd.n6614 585
R958 gnd.n6657 gnd.n6613 585
R959 gnd.n6658 gnd.n6611 585
R960 gnd.n6659 gnd.n6610 585
R961 gnd.n6608 gnd.n6606 585
R962 gnd.n6663 gnd.n6605 585
R963 gnd.n6664 gnd.n6603 585
R964 gnd.n6665 gnd.n6602 585
R965 gnd.n6602 gnd.n83 585
R966 gnd.n6766 gnd.n6765 585
R967 gnd.n6765 gnd.n6764 585
R968 gnd.n79 gnd.n77 585
R969 gnd.n81 gnd.n79 585
R970 gnd.n6770 gnd.n76 585
R971 gnd.n6684 gnd.n76 585
R972 gnd.n6771 gnd.n75 585
R973 gnd.n161 gnd.n75 585
R974 gnd.n6772 gnd.n74 585
R975 gnd.n6676 gnd.n74 585
R976 gnd.n168 gnd.n72 585
R977 gnd.n169 gnd.n168 585
R978 gnd.n6776 gnd.n71 585
R979 gnd.n6594 gnd.n71 585
R980 gnd.n6777 gnd.n70 585
R981 gnd.n188 gnd.n70 585
R982 gnd.n6778 gnd.n69 585
R983 gnd.n6586 gnd.n69 585
R984 gnd.n185 gnd.n67 585
R985 gnd.n186 gnd.n185 585
R986 gnd.n6782 gnd.n66 585
R987 gnd.n6578 gnd.n66 585
R988 gnd.n6783 gnd.n65 585
R989 gnd.n194 gnd.n65 585
R990 gnd.n6784 gnd.n64 585
R991 gnd.n6570 gnd.n64 585
R992 gnd.n201 gnd.n62 585
R993 gnd.n202 gnd.n201 585
R994 gnd.n6788 gnd.n61 585
R995 gnd.n6562 gnd.n61 585
R996 gnd.n6789 gnd.n60 585
R997 gnd.n224 gnd.n60 585
R998 gnd.n6790 gnd.n59 585
R999 gnd.n6554 gnd.n59 585
R1000 gnd.n221 gnd.n57 585
R1001 gnd.n222 gnd.n221 585
R1002 gnd.n6794 gnd.n56 585
R1003 gnd.n6546 gnd.n56 585
R1004 gnd.n6795 gnd.n55 585
R1005 gnd.n230 gnd.n55 585
R1006 gnd.n6796 gnd.n54 585
R1007 gnd.n6540 gnd.n54 585
R1008 gnd.n244 gnd.n52 585
R1009 gnd.n244 gnd.n235 585
R1010 gnd.n251 gnd.n245 585
R1011 gnd.n6532 gnd.n245 585
R1012 gnd.n6526 gnd.n6525 585
R1013 gnd.n6527 gnd.n6526 585
R1014 gnd.n250 gnd.n249 585
R1015 gnd.n249 gnd.n247 585
R1016 gnd.n6521 gnd.n6520 585
R1017 gnd.n6520 gnd.n6519 585
R1018 gnd.n254 gnd.n253 585
R1019 gnd.n6514 gnd.n254 585
R1020 gnd.n6290 gnd.n6288 585
R1021 gnd.n6288 gnd.n6287 585
R1022 gnd.n6291 gnd.n270 585
R1023 gnd.n6502 gnd.n270 585
R1024 gnd.n6292 gnd.n480 585
R1025 gnd.n6221 gnd.n480 585
R1026 gnd.n478 gnd.n278 585
R1027 gnd.n6493 gnd.n278 585
R1028 gnd.n6296 gnd.n477 585
R1029 gnd.n6217 gnd.n477 585
R1030 gnd.n6297 gnd.n287 585
R1031 gnd.n6485 gnd.n287 585
R1032 gnd.n6298 gnd.n476 585
R1033 gnd.n497 gnd.n476 585
R1034 gnd.n474 gnd.n296 585
R1035 gnd.n6477 gnd.n296 585
R1036 gnd.n6302 gnd.n473 585
R1037 gnd.n493 gnd.n473 585
R1038 gnd.n6303 gnd.n305 585
R1039 gnd.n6469 gnd.n305 585
R1040 gnd.n6304 gnd.n472 585
R1041 gnd.n487 gnd.n472 585
R1042 gnd.n469 gnd.n314 585
R1043 gnd.n6461 gnd.n314 585
R1044 gnd.n6309 gnd.n6308 585
R1045 gnd.n6310 gnd.n6309 585
R1046 gnd.n468 gnd.n322 585
R1047 gnd.n6453 gnd.n322 585
R1048 gnd.n5152 gnd.n5151 585
R1049 gnd.n5151 gnd.n5150 585
R1050 gnd.n5153 gnd.n330 585
R1051 gnd.n6445 gnd.n330 585
R1052 gnd.n3478 gnd.n3477 585
R1053 gnd.n3479 gnd.n3478 585
R1054 gnd.n2196 gnd.n2195 585
R1055 gnd.n2202 gnd.n2195 585
R1056 gnd.n3453 gnd.n2214 585
R1057 gnd.n2214 gnd.n2201 585
R1058 gnd.n3455 gnd.n3454 585
R1059 gnd.n3456 gnd.n3455 585
R1060 gnd.n2215 gnd.n2213 585
R1061 gnd.n2213 gnd.n2209 585
R1062 gnd.n3187 gnd.n3186 585
R1063 gnd.n3186 gnd.n3185 585
R1064 gnd.n2220 gnd.n2219 585
R1065 gnd.n3155 gnd.n2220 585
R1066 gnd.n3175 gnd.n3174 585
R1067 gnd.n3174 gnd.n3173 585
R1068 gnd.n2227 gnd.n2226 585
R1069 gnd.n3161 gnd.n2227 585
R1070 gnd.n3131 gnd.n2247 585
R1071 gnd.n2247 gnd.n2246 585
R1072 gnd.n3133 gnd.n3132 585
R1073 gnd.n3134 gnd.n3133 585
R1074 gnd.n2248 gnd.n2245 585
R1075 gnd.n2256 gnd.n2245 585
R1076 gnd.n3109 gnd.n2268 585
R1077 gnd.n2268 gnd.n2255 585
R1078 gnd.n3111 gnd.n3110 585
R1079 gnd.n3112 gnd.n3111 585
R1080 gnd.n2269 gnd.n2267 585
R1081 gnd.n2267 gnd.n2263 585
R1082 gnd.n3097 gnd.n3096 585
R1083 gnd.n3096 gnd.n3095 585
R1084 gnd.n2274 gnd.n2273 585
R1085 gnd.n2284 gnd.n2274 585
R1086 gnd.n3086 gnd.n3085 585
R1087 gnd.n3085 gnd.n3084 585
R1088 gnd.n2281 gnd.n2280 585
R1089 gnd.n3072 gnd.n2281 585
R1090 gnd.n3046 gnd.n2302 585
R1091 gnd.n2302 gnd.n2291 585
R1092 gnd.n3048 gnd.n3047 585
R1093 gnd.n3049 gnd.n3048 585
R1094 gnd.n2303 gnd.n2301 585
R1095 gnd.n2311 gnd.n2301 585
R1096 gnd.n3024 gnd.n2323 585
R1097 gnd.n2323 gnd.n2310 585
R1098 gnd.n3026 gnd.n3025 585
R1099 gnd.n3027 gnd.n3026 585
R1100 gnd.n2324 gnd.n2322 585
R1101 gnd.n2322 gnd.n2318 585
R1102 gnd.n3012 gnd.n3011 585
R1103 gnd.n3011 gnd.n3010 585
R1104 gnd.n2329 gnd.n2328 585
R1105 gnd.n2338 gnd.n2329 585
R1106 gnd.n3001 gnd.n3000 585
R1107 gnd.n3000 gnd.n2999 585
R1108 gnd.n2336 gnd.n2335 585
R1109 gnd.n2987 gnd.n2336 585
R1110 gnd.n2425 gnd.n2424 585
R1111 gnd.n2425 gnd.n2345 585
R1112 gnd.n2944 gnd.n2943 585
R1113 gnd.n2943 gnd.n2942 585
R1114 gnd.n2945 gnd.n2419 585
R1115 gnd.n2430 gnd.n2419 585
R1116 gnd.n2947 gnd.n2946 585
R1117 gnd.n2948 gnd.n2947 585
R1118 gnd.n2420 gnd.n2418 585
R1119 gnd.n2443 gnd.n2418 585
R1120 gnd.n2403 gnd.n2402 585
R1121 gnd.n2406 gnd.n2403 585
R1122 gnd.n2958 gnd.n2957 585
R1123 gnd.n2957 gnd.n2956 585
R1124 gnd.n2959 gnd.n2397 585
R1125 gnd.n2918 gnd.n2397 585
R1126 gnd.n2961 gnd.n2960 585
R1127 gnd.n2962 gnd.n2961 585
R1128 gnd.n2398 gnd.n2396 585
R1129 gnd.n2457 gnd.n2396 585
R1130 gnd.n2910 gnd.n2909 585
R1131 gnd.n2909 gnd.n2908 585
R1132 gnd.n2454 gnd.n2453 585
R1133 gnd.n2892 gnd.n2454 585
R1134 gnd.n2879 gnd.n2473 585
R1135 gnd.n2473 gnd.n2472 585
R1136 gnd.n2881 gnd.n2880 585
R1137 gnd.n2882 gnd.n2881 585
R1138 gnd.n2474 gnd.n2471 585
R1139 gnd.n2480 gnd.n2471 585
R1140 gnd.n2860 gnd.n2859 585
R1141 gnd.n2861 gnd.n2860 585
R1142 gnd.n2491 gnd.n2490 585
R1143 gnd.n2490 gnd.n2486 585
R1144 gnd.n2850 gnd.n2849 585
R1145 gnd.n2851 gnd.n2850 585
R1146 gnd.n2501 gnd.n2500 585
R1147 gnd.n2506 gnd.n2500 585
R1148 gnd.n2828 gnd.n2519 585
R1149 gnd.n2519 gnd.n2505 585
R1150 gnd.n2830 gnd.n2829 585
R1151 gnd.n2831 gnd.n2830 585
R1152 gnd.n2520 gnd.n2518 585
R1153 gnd.n2518 gnd.n2514 585
R1154 gnd.n2819 gnd.n2818 585
R1155 gnd.n2820 gnd.n2819 585
R1156 gnd.n2527 gnd.n2526 585
R1157 gnd.n2531 gnd.n2526 585
R1158 gnd.n2796 gnd.n2548 585
R1159 gnd.n2548 gnd.n2530 585
R1160 gnd.n2798 gnd.n2797 585
R1161 gnd.n2799 gnd.n2798 585
R1162 gnd.n2549 gnd.n2547 585
R1163 gnd.n2547 gnd.n2538 585
R1164 gnd.n2791 gnd.n2790 585
R1165 gnd.n2790 gnd.n2789 585
R1166 gnd.n2596 gnd.n2595 585
R1167 gnd.n2597 gnd.n2596 585
R1168 gnd.n2750 gnd.n2749 585
R1169 gnd.n2751 gnd.n2750 585
R1170 gnd.n2606 gnd.n2605 585
R1171 gnd.n2605 gnd.n2604 585
R1172 gnd.n2745 gnd.n2744 585
R1173 gnd.n2744 gnd.n2743 585
R1174 gnd.n2609 gnd.n2608 585
R1175 gnd.n2610 gnd.n2609 585
R1176 gnd.n2734 gnd.n2733 585
R1177 gnd.n2735 gnd.n2734 585
R1178 gnd.n2617 gnd.n2616 585
R1179 gnd.n2726 gnd.n2616 585
R1180 gnd.n2729 gnd.n2728 585
R1181 gnd.n2728 gnd.n2727 585
R1182 gnd.n2620 gnd.n2619 585
R1183 gnd.n2621 gnd.n2620 585
R1184 gnd.n2715 gnd.n2714 585
R1185 gnd.n2713 gnd.n2639 585
R1186 gnd.n2712 gnd.n2638 585
R1187 gnd.n2717 gnd.n2638 585
R1188 gnd.n2711 gnd.n2710 585
R1189 gnd.n2709 gnd.n2708 585
R1190 gnd.n2707 gnd.n2706 585
R1191 gnd.n2705 gnd.n2704 585
R1192 gnd.n2703 gnd.n2702 585
R1193 gnd.n2701 gnd.n2700 585
R1194 gnd.n2699 gnd.n2698 585
R1195 gnd.n2697 gnd.n2696 585
R1196 gnd.n2695 gnd.n2694 585
R1197 gnd.n2693 gnd.n2692 585
R1198 gnd.n2691 gnd.n2690 585
R1199 gnd.n2689 gnd.n2688 585
R1200 gnd.n2687 gnd.n2686 585
R1201 gnd.n2685 gnd.n2684 585
R1202 gnd.n2683 gnd.n2682 585
R1203 gnd.n2681 gnd.n2680 585
R1204 gnd.n2679 gnd.n2678 585
R1205 gnd.n2677 gnd.n2676 585
R1206 gnd.n2675 gnd.n2674 585
R1207 gnd.n2673 gnd.n2672 585
R1208 gnd.n2671 gnd.n2670 585
R1209 gnd.n2669 gnd.n2668 585
R1210 gnd.n2626 gnd.n2625 585
R1211 gnd.n2720 gnd.n2719 585
R1212 gnd.n3482 gnd.n3481 585
R1213 gnd.n3484 gnd.n3483 585
R1214 gnd.n3486 gnd.n3485 585
R1215 gnd.n3488 gnd.n3487 585
R1216 gnd.n3490 gnd.n3489 585
R1217 gnd.n3492 gnd.n3491 585
R1218 gnd.n3494 gnd.n3493 585
R1219 gnd.n3496 gnd.n3495 585
R1220 gnd.n3498 gnd.n3497 585
R1221 gnd.n3500 gnd.n3499 585
R1222 gnd.n3502 gnd.n3501 585
R1223 gnd.n3504 gnd.n3503 585
R1224 gnd.n3506 gnd.n3505 585
R1225 gnd.n3508 gnd.n3507 585
R1226 gnd.n3510 gnd.n3509 585
R1227 gnd.n3512 gnd.n3511 585
R1228 gnd.n3514 gnd.n3513 585
R1229 gnd.n3516 gnd.n3515 585
R1230 gnd.n3518 gnd.n3517 585
R1231 gnd.n3520 gnd.n3519 585
R1232 gnd.n3522 gnd.n3521 585
R1233 gnd.n3524 gnd.n3523 585
R1234 gnd.n3526 gnd.n3525 585
R1235 gnd.n3528 gnd.n3527 585
R1236 gnd.n3530 gnd.n3529 585
R1237 gnd.n3531 gnd.n2163 585
R1238 gnd.n3532 gnd.n2121 585
R1239 gnd.n3570 gnd.n2121 585
R1240 gnd.n3480 gnd.n2193 585
R1241 gnd.n3480 gnd.n3479 585
R1242 gnd.n3148 gnd.n2192 585
R1243 gnd.n2202 gnd.n2192 585
R1244 gnd.n3150 gnd.n3149 585
R1245 gnd.n3149 gnd.n2201 585
R1246 gnd.n3151 gnd.n2211 585
R1247 gnd.n3456 gnd.n2211 585
R1248 gnd.n3153 gnd.n3152 585
R1249 gnd.n3152 gnd.n2209 585
R1250 gnd.n3154 gnd.n2222 585
R1251 gnd.n3185 gnd.n2222 585
R1252 gnd.n3157 gnd.n3156 585
R1253 gnd.n3156 gnd.n3155 585
R1254 gnd.n3158 gnd.n2229 585
R1255 gnd.n3173 gnd.n2229 585
R1256 gnd.n3160 gnd.n3159 585
R1257 gnd.n3161 gnd.n3160 585
R1258 gnd.n2239 gnd.n2238 585
R1259 gnd.n2246 gnd.n2238 585
R1260 gnd.n3136 gnd.n3135 585
R1261 gnd.n3135 gnd.n3134 585
R1262 gnd.n2242 gnd.n2241 585
R1263 gnd.n2256 gnd.n2242 585
R1264 gnd.n3062 gnd.n3061 585
R1265 gnd.n3061 gnd.n2255 585
R1266 gnd.n3063 gnd.n2265 585
R1267 gnd.n3112 gnd.n2265 585
R1268 gnd.n3065 gnd.n3064 585
R1269 gnd.n3064 gnd.n2263 585
R1270 gnd.n3066 gnd.n2276 585
R1271 gnd.n3095 gnd.n2276 585
R1272 gnd.n3068 gnd.n3067 585
R1273 gnd.n3067 gnd.n2284 585
R1274 gnd.n3069 gnd.n2283 585
R1275 gnd.n3084 gnd.n2283 585
R1276 gnd.n3071 gnd.n3070 585
R1277 gnd.n3072 gnd.n3071 585
R1278 gnd.n2295 gnd.n2294 585
R1279 gnd.n2294 gnd.n2291 585
R1280 gnd.n3051 gnd.n3050 585
R1281 gnd.n3050 gnd.n3049 585
R1282 gnd.n2298 gnd.n2297 585
R1283 gnd.n2311 gnd.n2298 585
R1284 gnd.n2975 gnd.n2974 585
R1285 gnd.n2974 gnd.n2310 585
R1286 gnd.n2976 gnd.n2320 585
R1287 gnd.n3027 gnd.n2320 585
R1288 gnd.n2978 gnd.n2977 585
R1289 gnd.n2977 gnd.n2318 585
R1290 gnd.n2979 gnd.n2331 585
R1291 gnd.n3010 gnd.n2331 585
R1292 gnd.n2981 gnd.n2980 585
R1293 gnd.n2980 gnd.n2338 585
R1294 gnd.n2982 gnd.n2337 585
R1295 gnd.n2999 gnd.n2337 585
R1296 gnd.n2984 gnd.n2983 585
R1297 gnd.n2987 gnd.n2984 585
R1298 gnd.n2348 gnd.n2347 585
R1299 gnd.n2347 gnd.n2345 585
R1300 gnd.n2427 gnd.n2426 585
R1301 gnd.n2942 gnd.n2426 585
R1302 gnd.n2429 gnd.n2428 585
R1303 gnd.n2430 gnd.n2429 585
R1304 gnd.n2440 gnd.n2416 585
R1305 gnd.n2948 gnd.n2416 585
R1306 gnd.n2442 gnd.n2441 585
R1307 gnd.n2443 gnd.n2442 585
R1308 gnd.n2439 gnd.n2438 585
R1309 gnd.n2439 gnd.n2406 585
R1310 gnd.n2437 gnd.n2404 585
R1311 gnd.n2956 gnd.n2404 585
R1312 gnd.n2393 gnd.n2391 585
R1313 gnd.n2918 gnd.n2393 585
R1314 gnd.n2964 gnd.n2963 585
R1315 gnd.n2963 gnd.n2962 585
R1316 gnd.n2392 gnd.n2390 585
R1317 gnd.n2457 gnd.n2392 585
R1318 gnd.n2889 gnd.n2456 585
R1319 gnd.n2908 gnd.n2456 585
R1320 gnd.n2891 gnd.n2890 585
R1321 gnd.n2892 gnd.n2891 585
R1322 gnd.n2466 gnd.n2465 585
R1323 gnd.n2472 gnd.n2465 585
R1324 gnd.n2884 gnd.n2883 585
R1325 gnd.n2883 gnd.n2882 585
R1326 gnd.n2469 gnd.n2468 585
R1327 gnd.n2480 gnd.n2469 585
R1328 gnd.n2769 gnd.n2488 585
R1329 gnd.n2861 gnd.n2488 585
R1330 gnd.n2771 gnd.n2770 585
R1331 gnd.n2770 gnd.n2486 585
R1332 gnd.n2772 gnd.n2499 585
R1333 gnd.n2851 gnd.n2499 585
R1334 gnd.n2774 gnd.n2773 585
R1335 gnd.n2774 gnd.n2506 585
R1336 gnd.n2776 gnd.n2775 585
R1337 gnd.n2775 gnd.n2505 585
R1338 gnd.n2777 gnd.n2516 585
R1339 gnd.n2831 gnd.n2516 585
R1340 gnd.n2779 gnd.n2778 585
R1341 gnd.n2778 gnd.n2514 585
R1342 gnd.n2780 gnd.n2525 585
R1343 gnd.n2820 gnd.n2525 585
R1344 gnd.n2782 gnd.n2781 585
R1345 gnd.n2782 gnd.n2531 585
R1346 gnd.n2784 gnd.n2783 585
R1347 gnd.n2783 gnd.n2530 585
R1348 gnd.n2785 gnd.n2546 585
R1349 gnd.n2799 gnd.n2546 585
R1350 gnd.n2786 gnd.n2599 585
R1351 gnd.n2599 gnd.n2538 585
R1352 gnd.n2788 gnd.n2787 585
R1353 gnd.n2789 gnd.n2788 585
R1354 gnd.n2600 gnd.n2598 585
R1355 gnd.n2598 gnd.n2597 585
R1356 gnd.n2753 gnd.n2752 585
R1357 gnd.n2752 gnd.n2751 585
R1358 gnd.n2603 gnd.n2602 585
R1359 gnd.n2604 gnd.n2603 585
R1360 gnd.n2742 gnd.n2741 585
R1361 gnd.n2743 gnd.n2742 585
R1362 gnd.n2612 gnd.n2611 585
R1363 gnd.n2611 gnd.n2610 585
R1364 gnd.n2737 gnd.n2736 585
R1365 gnd.n2736 gnd.n2735 585
R1366 gnd.n2615 gnd.n2614 585
R1367 gnd.n2726 gnd.n2615 585
R1368 gnd.n2725 gnd.n2724 585
R1369 gnd.n2727 gnd.n2725 585
R1370 gnd.n2623 gnd.n2622 585
R1371 gnd.n2622 gnd.n2621 585
R1372 gnd.n3465 gnd.n2143 585
R1373 gnd.n2143 gnd.n2120 585
R1374 gnd.n3466 gnd.n2204 585
R1375 gnd.n2204 gnd.n2194 585
R1376 gnd.n3468 gnd.n3467 585
R1377 gnd.n3469 gnd.n3468 585
R1378 gnd.n2205 gnd.n2203 585
R1379 gnd.n2212 gnd.n2203 585
R1380 gnd.n3459 gnd.n3458 585
R1381 gnd.n3458 gnd.n3457 585
R1382 gnd.n2208 gnd.n2207 585
R1383 gnd.n3184 gnd.n2208 585
R1384 gnd.n3169 gnd.n2231 585
R1385 gnd.n2231 gnd.n2221 585
R1386 gnd.n3171 gnd.n3170 585
R1387 gnd.n3172 gnd.n3171 585
R1388 gnd.n2232 gnd.n2230 585
R1389 gnd.n2230 gnd.n2228 585
R1390 gnd.n3164 gnd.n3163 585
R1391 gnd.n3163 gnd.n3162 585
R1392 gnd.n2235 gnd.n2234 585
R1393 gnd.n2244 gnd.n2235 585
R1394 gnd.n3120 gnd.n2258 585
R1395 gnd.n2258 gnd.n2243 585
R1396 gnd.n3122 gnd.n3121 585
R1397 gnd.n3123 gnd.n3122 585
R1398 gnd.n2259 gnd.n2257 585
R1399 gnd.n2266 gnd.n2257 585
R1400 gnd.n3115 gnd.n3114 585
R1401 gnd.n3114 gnd.n3113 585
R1402 gnd.n2262 gnd.n2261 585
R1403 gnd.n3094 gnd.n2262 585
R1404 gnd.n3080 gnd.n2286 585
R1405 gnd.n2286 gnd.n2275 585
R1406 gnd.n3082 gnd.n3081 585
R1407 gnd.n3083 gnd.n3082 585
R1408 gnd.n2287 gnd.n2285 585
R1409 gnd.n2285 gnd.n2282 585
R1410 gnd.n3075 gnd.n3074 585
R1411 gnd.n3074 gnd.n3073 585
R1412 gnd.n2290 gnd.n2289 585
R1413 gnd.n2300 gnd.n2290 585
R1414 gnd.n3035 gnd.n2313 585
R1415 gnd.n2313 gnd.n2299 585
R1416 gnd.n3037 gnd.n3036 585
R1417 gnd.n3038 gnd.n3037 585
R1418 gnd.n2314 gnd.n2312 585
R1419 gnd.n2321 gnd.n2312 585
R1420 gnd.n3030 gnd.n3029 585
R1421 gnd.n3029 gnd.n3028 585
R1422 gnd.n2317 gnd.n2316 585
R1423 gnd.n3009 gnd.n2317 585
R1424 gnd.n2995 gnd.n2340 585
R1425 gnd.n2340 gnd.n2330 585
R1426 gnd.n2997 gnd.n2996 585
R1427 gnd.n2998 gnd.n2997 585
R1428 gnd.n2341 gnd.n2339 585
R1429 gnd.n2986 gnd.n2339 585
R1430 gnd.n2990 gnd.n2989 585
R1431 gnd.n2989 gnd.n2988 585
R1432 gnd.n2344 gnd.n2343 585
R1433 gnd.n2941 gnd.n2344 585
R1434 gnd.n2434 gnd.n2433 585
R1435 gnd.n2435 gnd.n2434 585
R1436 gnd.n2414 gnd.n2413 585
R1437 gnd.n2417 gnd.n2414 585
R1438 gnd.n2951 gnd.n2950 585
R1439 gnd.n2950 gnd.n2949 585
R1440 gnd.n2952 gnd.n2408 585
R1441 gnd.n2444 gnd.n2408 585
R1442 gnd.n2954 gnd.n2953 585
R1443 gnd.n2955 gnd.n2954 585
R1444 gnd.n2409 gnd.n2407 585
R1445 gnd.n2919 gnd.n2407 585
R1446 gnd.n2903 gnd.n2902 585
R1447 gnd.n2902 gnd.n2395 585
R1448 gnd.n2904 gnd.n2459 585
R1449 gnd.n2459 gnd.n2394 585
R1450 gnd.n2906 gnd.n2905 585
R1451 gnd.n2907 gnd.n2906 585
R1452 gnd.n2460 gnd.n2458 585
R1453 gnd.n2458 gnd.n2455 585
R1454 gnd.n2895 gnd.n2894 585
R1455 gnd.n2894 gnd.n2893 585
R1456 gnd.n2463 gnd.n2462 585
R1457 gnd.n2470 gnd.n2463 585
R1458 gnd.n2869 gnd.n2868 585
R1459 gnd.n2870 gnd.n2869 585
R1460 gnd.n2482 gnd.n2481 585
R1461 gnd.n2489 gnd.n2481 585
R1462 gnd.n2864 gnd.n2863 585
R1463 gnd.n2863 gnd.n2862 585
R1464 gnd.n2485 gnd.n2484 585
R1465 gnd.n2852 gnd.n2485 585
R1466 gnd.n2839 gnd.n2509 585
R1467 gnd.n2509 gnd.n2508 585
R1468 gnd.n2841 gnd.n2840 585
R1469 gnd.n2842 gnd.n2841 585
R1470 gnd.n2510 gnd.n2507 585
R1471 gnd.n2517 gnd.n2507 585
R1472 gnd.n2834 gnd.n2833 585
R1473 gnd.n2833 gnd.n2832 585
R1474 gnd.n2513 gnd.n2512 585
R1475 gnd.n2821 gnd.n2513 585
R1476 gnd.n2808 gnd.n2534 585
R1477 gnd.n2534 gnd.n2533 585
R1478 gnd.n2810 gnd.n2809 585
R1479 gnd.n2811 gnd.n2810 585
R1480 gnd.n2804 gnd.n2532 585
R1481 gnd.n2803 gnd.n2802 585
R1482 gnd.n2537 gnd.n2536 585
R1483 gnd.n2800 gnd.n2537 585
R1484 gnd.n2559 gnd.n2558 585
R1485 gnd.n2562 gnd.n2561 585
R1486 gnd.n2560 gnd.n2555 585
R1487 gnd.n2567 gnd.n2566 585
R1488 gnd.n2569 gnd.n2568 585
R1489 gnd.n2572 gnd.n2571 585
R1490 gnd.n2570 gnd.n2553 585
R1491 gnd.n2577 gnd.n2576 585
R1492 gnd.n2579 gnd.n2578 585
R1493 gnd.n2582 gnd.n2581 585
R1494 gnd.n2580 gnd.n2551 585
R1495 gnd.n2587 gnd.n2586 585
R1496 gnd.n2591 gnd.n2588 585
R1497 gnd.n2592 gnd.n2529 585
R1498 gnd.n3471 gnd.n2158 585
R1499 gnd.n3538 gnd.n3537 585
R1500 gnd.n3540 gnd.n3539 585
R1501 gnd.n3542 gnd.n3541 585
R1502 gnd.n3544 gnd.n3543 585
R1503 gnd.n3546 gnd.n3545 585
R1504 gnd.n3548 gnd.n3547 585
R1505 gnd.n3550 gnd.n3549 585
R1506 gnd.n3552 gnd.n3551 585
R1507 gnd.n3554 gnd.n3553 585
R1508 gnd.n3556 gnd.n3555 585
R1509 gnd.n3558 gnd.n3557 585
R1510 gnd.n3560 gnd.n3559 585
R1511 gnd.n3563 gnd.n3562 585
R1512 gnd.n3561 gnd.n2146 585
R1513 gnd.n3567 gnd.n2144 585
R1514 gnd.n3569 gnd.n3568 585
R1515 gnd.n3570 gnd.n3569 585
R1516 gnd.n3472 gnd.n2199 585
R1517 gnd.n3472 gnd.n2120 585
R1518 gnd.n3474 gnd.n3473 585
R1519 gnd.n3473 gnd.n2194 585
R1520 gnd.n3470 gnd.n2198 585
R1521 gnd.n3470 gnd.n3469 585
R1522 gnd.n3449 gnd.n2200 585
R1523 gnd.n2212 gnd.n2200 585
R1524 gnd.n3448 gnd.n2210 585
R1525 gnd.n3457 gnd.n2210 585
R1526 gnd.n3182 gnd.n2217 585
R1527 gnd.n3184 gnd.n3182 585
R1528 gnd.n3181 gnd.n3180 585
R1529 gnd.n3181 gnd.n2221 585
R1530 gnd.n3179 gnd.n2223 585
R1531 gnd.n3172 gnd.n2223 585
R1532 gnd.n2236 gnd.n2224 585
R1533 gnd.n2236 gnd.n2228 585
R1534 gnd.n3128 gnd.n2237 585
R1535 gnd.n3162 gnd.n2237 585
R1536 gnd.n3127 gnd.n3126 585
R1537 gnd.n3126 gnd.n2244 585
R1538 gnd.n3125 gnd.n2252 585
R1539 gnd.n3125 gnd.n2243 585
R1540 gnd.n3124 gnd.n2254 585
R1541 gnd.n3124 gnd.n3123 585
R1542 gnd.n3103 gnd.n2253 585
R1543 gnd.n2266 gnd.n2253 585
R1544 gnd.n3102 gnd.n2264 585
R1545 gnd.n3113 gnd.n2264 585
R1546 gnd.n3093 gnd.n2271 585
R1547 gnd.n3094 gnd.n3093 585
R1548 gnd.n3092 gnd.n3091 585
R1549 gnd.n3092 gnd.n2275 585
R1550 gnd.n3090 gnd.n2277 585
R1551 gnd.n3083 gnd.n2277 585
R1552 gnd.n2292 gnd.n2278 585
R1553 gnd.n2292 gnd.n2282 585
R1554 gnd.n3043 gnd.n2293 585
R1555 gnd.n3073 gnd.n2293 585
R1556 gnd.n3042 gnd.n3041 585
R1557 gnd.n3041 gnd.n2300 585
R1558 gnd.n3040 gnd.n2307 585
R1559 gnd.n3040 gnd.n2299 585
R1560 gnd.n3039 gnd.n2309 585
R1561 gnd.n3039 gnd.n3038 585
R1562 gnd.n3018 gnd.n2308 585
R1563 gnd.n2321 gnd.n2308 585
R1564 gnd.n3017 gnd.n2319 585
R1565 gnd.n3028 gnd.n2319 585
R1566 gnd.n3008 gnd.n2326 585
R1567 gnd.n3009 gnd.n3008 585
R1568 gnd.n3007 gnd.n3006 585
R1569 gnd.n3007 gnd.n2330 585
R1570 gnd.n3005 gnd.n2332 585
R1571 gnd.n2998 gnd.n2332 585
R1572 gnd.n2985 gnd.n2333 585
R1573 gnd.n2986 gnd.n2985 585
R1574 gnd.n2938 gnd.n2346 585
R1575 gnd.n2988 gnd.n2346 585
R1576 gnd.n2940 gnd.n2939 585
R1577 gnd.n2941 gnd.n2940 585
R1578 gnd.n2933 gnd.n2436 585
R1579 gnd.n2436 gnd.n2435 585
R1580 gnd.n2931 gnd.n2930 585
R1581 gnd.n2930 gnd.n2417 585
R1582 gnd.n2928 gnd.n2415 585
R1583 gnd.n2949 gnd.n2415 585
R1584 gnd.n2446 gnd.n2445 585
R1585 gnd.n2445 gnd.n2444 585
R1586 gnd.n2922 gnd.n2405 585
R1587 gnd.n2955 gnd.n2405 585
R1588 gnd.n2921 gnd.n2920 585
R1589 gnd.n2920 gnd.n2919 585
R1590 gnd.n2917 gnd.n2448 585
R1591 gnd.n2917 gnd.n2395 585
R1592 gnd.n2916 gnd.n2915 585
R1593 gnd.n2916 gnd.n2394 585
R1594 gnd.n2451 gnd.n2450 585
R1595 gnd.n2907 gnd.n2450 585
R1596 gnd.n2875 gnd.n2874 585
R1597 gnd.n2874 gnd.n2455 585
R1598 gnd.n2876 gnd.n2464 585
R1599 gnd.n2893 gnd.n2464 585
R1600 gnd.n2873 gnd.n2872 585
R1601 gnd.n2872 gnd.n2470 585
R1602 gnd.n2871 gnd.n2478 585
R1603 gnd.n2871 gnd.n2870 585
R1604 gnd.n2856 gnd.n2479 585
R1605 gnd.n2489 gnd.n2479 585
R1606 gnd.n2855 gnd.n2487 585
R1607 gnd.n2862 gnd.n2487 585
R1608 gnd.n2854 gnd.n2853 585
R1609 gnd.n2853 gnd.n2852 585
R1610 gnd.n2498 gnd.n2495 585
R1611 gnd.n2508 gnd.n2498 585
R1612 gnd.n2844 gnd.n2843 585
R1613 gnd.n2843 gnd.n2842 585
R1614 gnd.n2504 gnd.n2503 585
R1615 gnd.n2517 gnd.n2504 585
R1616 gnd.n2824 gnd.n2515 585
R1617 gnd.n2832 gnd.n2515 585
R1618 gnd.n2823 gnd.n2822 585
R1619 gnd.n2822 gnd.n2821 585
R1620 gnd.n2524 gnd.n2522 585
R1621 gnd.n2533 gnd.n2524 585
R1622 gnd.n2813 gnd.n2812 585
R1623 gnd.n2812 gnd.n2811 585
R1624 gnd.n5442 gnd.n1089 585
R1625 gnd.n4186 gnd.n1089 585
R1626 gnd.n5444 gnd.n5443 585
R1627 gnd.n5445 gnd.n5444 585
R1628 gnd.n1073 gnd.n1072 585
R1629 gnd.n4149 gnd.n1073 585
R1630 gnd.n5453 gnd.n5452 585
R1631 gnd.n5452 gnd.n5451 585
R1632 gnd.n5454 gnd.n1067 585
R1633 gnd.n4073 gnd.n1067 585
R1634 gnd.n5456 gnd.n5455 585
R1635 gnd.n5457 gnd.n5456 585
R1636 gnd.n1052 gnd.n1051 585
R1637 gnd.n4162 gnd.n1052 585
R1638 gnd.n5465 gnd.n5464 585
R1639 gnd.n5464 gnd.n5463 585
R1640 gnd.n5466 gnd.n1046 585
R1641 gnd.n4065 gnd.n1046 585
R1642 gnd.n5468 gnd.n5467 585
R1643 gnd.n5469 gnd.n5468 585
R1644 gnd.n1031 gnd.n1030 585
R1645 gnd.n4057 gnd.n1031 585
R1646 gnd.n5477 gnd.n5476 585
R1647 gnd.n5476 gnd.n5475 585
R1648 gnd.n5478 gnd.n1025 585
R1649 gnd.n4022 gnd.n1025 585
R1650 gnd.n5480 gnd.n5479 585
R1651 gnd.n5481 gnd.n5480 585
R1652 gnd.n1009 gnd.n1008 585
R1653 gnd.n4030 gnd.n1009 585
R1654 gnd.n5489 gnd.n5488 585
R1655 gnd.n5488 gnd.n5487 585
R1656 gnd.n5490 gnd.n1004 585
R1657 gnd.n4008 gnd.n1004 585
R1658 gnd.n5492 gnd.n5491 585
R1659 gnd.n5493 gnd.n5492 585
R1660 gnd.n3996 gnd.n1003 585
R1661 gnd.n1003 gnd.n998 585
R1662 gnd.n3998 gnd.n3997 585
R1663 gnd.n3999 gnd.n3998 585
R1664 gnd.n3994 gnd.n2026 585
R1665 gnd.n2032 gnd.n2026 585
R1666 gnd.n3993 gnd.n3992 585
R1667 gnd.n3992 gnd.n3991 585
R1668 gnd.n3961 gnd.n2028 585
R1669 gnd.n2029 gnd.n2028 585
R1670 gnd.n3963 gnd.n3962 585
R1671 gnd.n3964 gnd.n3963 585
R1672 gnd.n3959 gnd.n2044 585
R1673 gnd.n2044 gnd.n2041 585
R1674 gnd.n3958 gnd.n3957 585
R1675 gnd.n3957 gnd.n3956 585
R1676 gnd.n3941 gnd.n2046 585
R1677 gnd.n2047 gnd.n2046 585
R1678 gnd.n3943 gnd.n3942 585
R1679 gnd.n3944 gnd.n3943 585
R1680 gnd.n2059 gnd.n2058 585
R1681 gnd.n2066 gnd.n2058 585
R1682 gnd.n3937 gnd.n3936 585
R1683 gnd.n3936 gnd.n3935 585
R1684 gnd.n2062 gnd.n2061 585
R1685 gnd.n2063 gnd.n2062 585
R1686 gnd.n3926 gnd.n3925 585
R1687 gnd.n3927 gnd.n3926 585
R1688 gnd.n2076 gnd.n2075 585
R1689 gnd.n2075 gnd.n2072 585
R1690 gnd.n3921 gnd.n3920 585
R1691 gnd.n3920 gnd.n3919 585
R1692 gnd.n2079 gnd.n2078 585
R1693 gnd.n2080 gnd.n2079 585
R1694 gnd.n3910 gnd.n3909 585
R1695 gnd.n3911 gnd.n3910 585
R1696 gnd.n2091 gnd.n2090 585
R1697 gnd.n2098 gnd.n2090 585
R1698 gnd.n3905 gnd.n3904 585
R1699 gnd.n3904 gnd.n3903 585
R1700 gnd.n2094 gnd.n2093 585
R1701 gnd.n2095 gnd.n2094 585
R1702 gnd.n3894 gnd.n3893 585
R1703 gnd.n3895 gnd.n3894 585
R1704 gnd.n2108 gnd.n2107 585
R1705 gnd.n2107 gnd.n2104 585
R1706 gnd.n3889 gnd.n3888 585
R1707 gnd.n3888 gnd.n3887 585
R1708 gnd.n2111 gnd.n2110 585
R1709 gnd.n2112 gnd.n2111 585
R1710 gnd.n3876 gnd.n3875 585
R1711 gnd.n3874 gnd.n3708 585
R1712 gnd.n3873 gnd.n3707 585
R1713 gnd.n3878 gnd.n3707 585
R1714 gnd.n3872 gnd.n3871 585
R1715 gnd.n3870 gnd.n3869 585
R1716 gnd.n3868 gnd.n3867 585
R1717 gnd.n3866 gnd.n3865 585
R1718 gnd.n3864 gnd.n3863 585
R1719 gnd.n3862 gnd.n3861 585
R1720 gnd.n3860 gnd.n3859 585
R1721 gnd.n3858 gnd.n3857 585
R1722 gnd.n3856 gnd.n3855 585
R1723 gnd.n3854 gnd.n3853 585
R1724 gnd.n3852 gnd.n3851 585
R1725 gnd.n3850 gnd.n3849 585
R1726 gnd.n3848 gnd.n3847 585
R1727 gnd.n3846 gnd.n3845 585
R1728 gnd.n3844 gnd.n3843 585
R1729 gnd.n3841 gnd.n3840 585
R1730 gnd.n3839 gnd.n3838 585
R1731 gnd.n3837 gnd.n3836 585
R1732 gnd.n3835 gnd.n3834 585
R1733 gnd.n3833 gnd.n3832 585
R1734 gnd.n3831 gnd.n3830 585
R1735 gnd.n3829 gnd.n3828 585
R1736 gnd.n3827 gnd.n3826 585
R1737 gnd.n3825 gnd.n3824 585
R1738 gnd.n3823 gnd.n3822 585
R1739 gnd.n3821 gnd.n3820 585
R1740 gnd.n3819 gnd.n3818 585
R1741 gnd.n3817 gnd.n3816 585
R1742 gnd.n3815 gnd.n3814 585
R1743 gnd.n3813 gnd.n3812 585
R1744 gnd.n3811 gnd.n3810 585
R1745 gnd.n3809 gnd.n3808 585
R1746 gnd.n3807 gnd.n3806 585
R1747 gnd.n3805 gnd.n3747 585
R1748 gnd.n3751 gnd.n3748 585
R1749 gnd.n3801 gnd.n3800 585
R1750 gnd.n4142 gnd.n4141 585
R1751 gnd.n4140 gnd.n4083 585
R1752 gnd.n4139 gnd.n4138 585
R1753 gnd.n4132 gnd.n4084 585
R1754 gnd.n4134 gnd.n4133 585
R1755 gnd.n4131 gnd.n4130 585
R1756 gnd.n4129 gnd.n4128 585
R1757 gnd.n4122 gnd.n4086 585
R1758 gnd.n4124 gnd.n4123 585
R1759 gnd.n4121 gnd.n4120 585
R1760 gnd.n4119 gnd.n4118 585
R1761 gnd.n4112 gnd.n4088 585
R1762 gnd.n4114 gnd.n4113 585
R1763 gnd.n4111 gnd.n4110 585
R1764 gnd.n4109 gnd.n4108 585
R1765 gnd.n4102 gnd.n4090 585
R1766 gnd.n4104 gnd.n4103 585
R1767 gnd.n4101 gnd.n4100 585
R1768 gnd.n4099 gnd.n4098 585
R1769 gnd.n4094 gnd.n4093 585
R1770 gnd.n4092 gnd.n1140 585
R1771 gnd.n5410 gnd.n5409 585
R1772 gnd.n5412 gnd.n5411 585
R1773 gnd.n5414 gnd.n5413 585
R1774 gnd.n5416 gnd.n5415 585
R1775 gnd.n5418 gnd.n5417 585
R1776 gnd.n5420 gnd.n5419 585
R1777 gnd.n5422 gnd.n5421 585
R1778 gnd.n5424 gnd.n5423 585
R1779 gnd.n5426 gnd.n5425 585
R1780 gnd.n5428 gnd.n5427 585
R1781 gnd.n5430 gnd.n5429 585
R1782 gnd.n5432 gnd.n5431 585
R1783 gnd.n5433 gnd.n1125 585
R1784 gnd.n5435 gnd.n5434 585
R1785 gnd.n1094 gnd.n1093 585
R1786 gnd.n5439 gnd.n5438 585
R1787 gnd.n5438 gnd.n5437 585
R1788 gnd.n4145 gnd.n1981 585
R1789 gnd.n4186 gnd.n1981 585
R1790 gnd.n4146 gnd.n1086 585
R1791 gnd.n5445 gnd.n1086 585
R1792 gnd.n4148 gnd.n4147 585
R1793 gnd.n4149 gnd.n4148 585
R1794 gnd.n1998 gnd.n1075 585
R1795 gnd.n5451 gnd.n1075 585
R1796 gnd.n4075 gnd.n4074 585
R1797 gnd.n4074 gnd.n4073 585
R1798 gnd.n4072 gnd.n1064 585
R1799 gnd.n5457 gnd.n1064 585
R1800 gnd.n4071 gnd.n1992 585
R1801 gnd.n4162 gnd.n1992 585
R1802 gnd.n2000 gnd.n1054 585
R1803 gnd.n5463 gnd.n1054 585
R1804 gnd.n4067 gnd.n4066 585
R1805 gnd.n4066 gnd.n4065 585
R1806 gnd.n2002 gnd.n1043 585
R1807 gnd.n5469 gnd.n1043 585
R1808 gnd.n4018 gnd.n2006 585
R1809 gnd.n4057 gnd.n2006 585
R1810 gnd.n4019 gnd.n1033 585
R1811 gnd.n5475 gnd.n1033 585
R1812 gnd.n4021 gnd.n4020 585
R1813 gnd.n4022 gnd.n4021 585
R1814 gnd.n2016 gnd.n1022 585
R1815 gnd.n5481 gnd.n1022 585
R1816 gnd.n4012 gnd.n2012 585
R1817 gnd.n4030 gnd.n2012 585
R1818 gnd.n4011 gnd.n1011 585
R1819 gnd.n5487 gnd.n1011 585
R1820 gnd.n4010 gnd.n4009 585
R1821 gnd.n4009 gnd.n4008 585
R1822 gnd.n2018 gnd.n999 585
R1823 gnd.n5493 gnd.n999 585
R1824 gnd.n3972 gnd.n3971 585
R1825 gnd.n3971 gnd.n998 585
R1826 gnd.n3973 gnd.n2024 585
R1827 gnd.n3999 gnd.n2024 585
R1828 gnd.n3975 gnd.n3974 585
R1829 gnd.n3974 gnd.n2032 585
R1830 gnd.n3976 gnd.n2030 585
R1831 gnd.n3991 gnd.n2030 585
R1832 gnd.n3967 gnd.n3966 585
R1833 gnd.n3966 gnd.n2029 585
R1834 gnd.n3965 gnd.n2039 585
R1835 gnd.n3965 gnd.n3964 585
R1836 gnd.n3771 gnd.n2040 585
R1837 gnd.n2041 gnd.n2040 585
R1838 gnd.n3772 gnd.n2048 585
R1839 gnd.n3956 gnd.n2048 585
R1840 gnd.n3774 gnd.n3773 585
R1841 gnd.n3773 gnd.n2047 585
R1842 gnd.n3775 gnd.n2056 585
R1843 gnd.n3944 gnd.n2056 585
R1844 gnd.n3777 gnd.n3776 585
R1845 gnd.n3776 gnd.n2066 585
R1846 gnd.n3778 gnd.n2064 585
R1847 gnd.n3935 gnd.n2064 585
R1848 gnd.n3780 gnd.n3779 585
R1849 gnd.n3779 gnd.n2063 585
R1850 gnd.n3781 gnd.n2073 585
R1851 gnd.n3927 gnd.n2073 585
R1852 gnd.n3783 gnd.n3782 585
R1853 gnd.n3782 gnd.n2072 585
R1854 gnd.n3784 gnd.n2081 585
R1855 gnd.n3919 gnd.n2081 585
R1856 gnd.n3786 gnd.n3785 585
R1857 gnd.n3785 gnd.n2080 585
R1858 gnd.n3787 gnd.n2088 585
R1859 gnd.n3911 gnd.n2088 585
R1860 gnd.n3789 gnd.n3788 585
R1861 gnd.n3788 gnd.n2098 585
R1862 gnd.n3790 gnd.n2096 585
R1863 gnd.n3903 gnd.n2096 585
R1864 gnd.n3792 gnd.n3791 585
R1865 gnd.n3791 gnd.n2095 585
R1866 gnd.n3793 gnd.n2105 585
R1867 gnd.n3895 gnd.n2105 585
R1868 gnd.n3754 gnd.n3753 585
R1869 gnd.n3753 gnd.n2104 585
R1870 gnd.n3797 gnd.n2113 585
R1871 gnd.n3887 gnd.n2113 585
R1872 gnd.n3799 gnd.n3798 585
R1873 gnd.n3799 gnd.n2112 585
R1874 gnd.n6763 gnd.n6762 585
R1875 gnd.n6764 gnd.n6763 585
R1876 gnd.n87 gnd.n85 585
R1877 gnd.n85 gnd.n81 585
R1878 gnd.n6683 gnd.n6682 585
R1879 gnd.n6684 gnd.n6683 585
R1880 gnd.n164 gnd.n163 585
R1881 gnd.n163 gnd.n161 585
R1882 gnd.n6678 gnd.n6677 585
R1883 gnd.n6677 gnd.n6676 585
R1884 gnd.n167 gnd.n166 585
R1885 gnd.n169 gnd.n167 585
R1886 gnd.n6593 gnd.n6592 585
R1887 gnd.n6594 gnd.n6593 585
R1888 gnd.n181 gnd.n180 585
R1889 gnd.n188 gnd.n180 585
R1890 gnd.n6588 gnd.n6587 585
R1891 gnd.n6587 gnd.n6586 585
R1892 gnd.n184 gnd.n183 585
R1893 gnd.n186 gnd.n184 585
R1894 gnd.n6577 gnd.n6576 585
R1895 gnd.n6578 gnd.n6577 585
R1896 gnd.n197 gnd.n196 585
R1897 gnd.n196 gnd.n194 585
R1898 gnd.n6572 gnd.n6571 585
R1899 gnd.n6571 gnd.n6570 585
R1900 gnd.n200 gnd.n199 585
R1901 gnd.n202 gnd.n200 585
R1902 gnd.n6561 gnd.n6560 585
R1903 gnd.n6562 gnd.n6561 585
R1904 gnd.n211 gnd.n210 585
R1905 gnd.n224 gnd.n210 585
R1906 gnd.n6556 gnd.n6555 585
R1907 gnd.n6555 gnd.n6554 585
R1908 gnd.n220 gnd.n219 585
R1909 gnd.n222 gnd.n220 585
R1910 gnd.n6545 gnd.n6544 585
R1911 gnd.n6546 gnd.n6545 585
R1912 gnd.n6543 gnd.n6542 585
R1913 gnd.n6542 gnd.n230 585
R1914 gnd.n6541 gnd.n234 585
R1915 gnd.n6541 gnd.n6540 585
R1916 gnd.n233 gnd.n232 585
R1917 gnd.n235 gnd.n232 585
R1918 gnd.n6531 gnd.n6530 585
R1919 gnd.n6532 gnd.n6531 585
R1920 gnd.n6529 gnd.n6528 585
R1921 gnd.n6528 gnd.n6527 585
R1922 gnd.n6516 gnd.n246 585
R1923 gnd.n247 gnd.n246 585
R1924 gnd.n6518 gnd.n6517 585
R1925 gnd.n6519 gnd.n6518 585
R1926 gnd.n6515 gnd.n259 585
R1927 gnd.n6515 gnd.n6514 585
R1928 gnd.n6499 gnd.n258 585
R1929 gnd.n6287 gnd.n258 585
R1930 gnd.n6501 gnd.n6500 585
R1931 gnd.n6502 gnd.n6501 585
R1932 gnd.n273 gnd.n272 585
R1933 gnd.n6221 gnd.n272 585
R1934 gnd.n6495 gnd.n6494 585
R1935 gnd.n6494 gnd.n6493 585
R1936 gnd.n276 gnd.n275 585
R1937 gnd.n6217 gnd.n276 585
R1938 gnd.n6484 gnd.n6483 585
R1939 gnd.n6485 gnd.n6484 585
R1940 gnd.n290 gnd.n289 585
R1941 gnd.n497 gnd.n289 585
R1942 gnd.n6479 gnd.n6478 585
R1943 gnd.n6478 gnd.n6477 585
R1944 gnd.n293 gnd.n292 585
R1945 gnd.n493 gnd.n293 585
R1946 gnd.n6468 gnd.n6467 585
R1947 gnd.n6469 gnd.n6468 585
R1948 gnd.n308 gnd.n307 585
R1949 gnd.n487 gnd.n307 585
R1950 gnd.n6463 gnd.n6462 585
R1951 gnd.n6462 gnd.n6461 585
R1952 gnd.n311 gnd.n310 585
R1953 gnd.n6310 gnd.n311 585
R1954 gnd.n6452 gnd.n6451 585
R1955 gnd.n6453 gnd.n6452 585
R1956 gnd.n325 gnd.n324 585
R1957 gnd.n5150 gnd.n324 585
R1958 gnd.n6447 gnd.n6446 585
R1959 gnd.n6446 gnd.n6445 585
R1960 gnd.n419 gnd.n327 585
R1961 gnd.n6388 gnd.n6387 585
R1962 gnd.n6386 gnd.n418 585
R1963 gnd.n6390 gnd.n418 585
R1964 gnd.n6385 gnd.n6384 585
R1965 gnd.n6383 gnd.n6382 585
R1966 gnd.n6381 gnd.n6380 585
R1967 gnd.n6379 gnd.n6378 585
R1968 gnd.n6377 gnd.n6376 585
R1969 gnd.n6375 gnd.n6374 585
R1970 gnd.n6373 gnd.n6372 585
R1971 gnd.n6371 gnd.n6370 585
R1972 gnd.n6369 gnd.n6368 585
R1973 gnd.n6367 gnd.n6366 585
R1974 gnd.n6365 gnd.n6364 585
R1975 gnd.n6363 gnd.n6362 585
R1976 gnd.n6361 gnd.n6360 585
R1977 gnd.n6358 gnd.n6357 585
R1978 gnd.n6356 gnd.n6355 585
R1979 gnd.n6354 gnd.n6353 585
R1980 gnd.n6352 gnd.n6351 585
R1981 gnd.n6350 gnd.n6349 585
R1982 gnd.n6348 gnd.n6347 585
R1983 gnd.n6346 gnd.n6345 585
R1984 gnd.n6344 gnd.n6343 585
R1985 gnd.n6342 gnd.n6341 585
R1986 gnd.n6340 gnd.n6339 585
R1987 gnd.n6338 gnd.n6337 585
R1988 gnd.n6336 gnd.n6335 585
R1989 gnd.n6334 gnd.n6333 585
R1990 gnd.n6332 gnd.n6331 585
R1991 gnd.n6330 gnd.n6329 585
R1992 gnd.n6328 gnd.n6327 585
R1993 gnd.n6326 gnd.n6325 585
R1994 gnd.n6324 gnd.n6323 585
R1995 gnd.n6322 gnd.n458 585
R1996 gnd.n462 gnd.n459 585
R1997 gnd.n6318 gnd.n6317 585
R1998 gnd.n155 gnd.n154 585
R1999 gnd.n6692 gnd.n150 585
R2000 gnd.n6694 gnd.n6693 585
R2001 gnd.n6696 gnd.n148 585
R2002 gnd.n6698 gnd.n6697 585
R2003 gnd.n6699 gnd.n143 585
R2004 gnd.n6701 gnd.n6700 585
R2005 gnd.n6703 gnd.n141 585
R2006 gnd.n6705 gnd.n6704 585
R2007 gnd.n6706 gnd.n136 585
R2008 gnd.n6708 gnd.n6707 585
R2009 gnd.n6710 gnd.n134 585
R2010 gnd.n6712 gnd.n6711 585
R2011 gnd.n6713 gnd.n129 585
R2012 gnd.n6715 gnd.n6714 585
R2013 gnd.n6717 gnd.n127 585
R2014 gnd.n6719 gnd.n6718 585
R2015 gnd.n6720 gnd.n122 585
R2016 gnd.n6722 gnd.n6721 585
R2017 gnd.n6724 gnd.n120 585
R2018 gnd.n6726 gnd.n6725 585
R2019 gnd.n6730 gnd.n115 585
R2020 gnd.n6732 gnd.n6731 585
R2021 gnd.n6734 gnd.n113 585
R2022 gnd.n6736 gnd.n6735 585
R2023 gnd.n6737 gnd.n108 585
R2024 gnd.n6739 gnd.n6738 585
R2025 gnd.n6741 gnd.n106 585
R2026 gnd.n6743 gnd.n6742 585
R2027 gnd.n6744 gnd.n101 585
R2028 gnd.n6746 gnd.n6745 585
R2029 gnd.n6748 gnd.n99 585
R2030 gnd.n6750 gnd.n6749 585
R2031 gnd.n6751 gnd.n94 585
R2032 gnd.n6753 gnd.n6752 585
R2033 gnd.n6755 gnd.n92 585
R2034 gnd.n6757 gnd.n6756 585
R2035 gnd.n6758 gnd.n90 585
R2036 gnd.n6759 gnd.n86 585
R2037 gnd.n86 gnd.n83 585
R2038 gnd.n6688 gnd.n82 585
R2039 gnd.n6764 gnd.n82 585
R2040 gnd.n6687 gnd.n6686 585
R2041 gnd.n6686 gnd.n81 585
R2042 gnd.n6685 gnd.n159 585
R2043 gnd.n6685 gnd.n6684 585
R2044 gnd.n6251 gnd.n160 585
R2045 gnd.n161 gnd.n160 585
R2046 gnd.n6252 gnd.n170 585
R2047 gnd.n6676 gnd.n170 585
R2048 gnd.n6254 gnd.n6253 585
R2049 gnd.n6253 gnd.n169 585
R2050 gnd.n6255 gnd.n178 585
R2051 gnd.n6594 gnd.n178 585
R2052 gnd.n6257 gnd.n6256 585
R2053 gnd.n6256 gnd.n188 585
R2054 gnd.n6258 gnd.n187 585
R2055 gnd.n6586 gnd.n187 585
R2056 gnd.n6260 gnd.n6259 585
R2057 gnd.n6259 gnd.n186 585
R2058 gnd.n6261 gnd.n195 585
R2059 gnd.n6578 gnd.n195 585
R2060 gnd.n6263 gnd.n6262 585
R2061 gnd.n6262 gnd.n194 585
R2062 gnd.n6264 gnd.n203 585
R2063 gnd.n6570 gnd.n203 585
R2064 gnd.n6266 gnd.n6265 585
R2065 gnd.n6265 gnd.n202 585
R2066 gnd.n6267 gnd.n209 585
R2067 gnd.n6562 gnd.n209 585
R2068 gnd.n6269 gnd.n6268 585
R2069 gnd.n6268 gnd.n224 585
R2070 gnd.n6270 gnd.n223 585
R2071 gnd.n6554 gnd.n223 585
R2072 gnd.n6272 gnd.n6271 585
R2073 gnd.n6271 gnd.n222 585
R2074 gnd.n6273 gnd.n231 585
R2075 gnd.n6546 gnd.n231 585
R2076 gnd.n6275 gnd.n6274 585
R2077 gnd.n6274 gnd.n230 585
R2078 gnd.n6276 gnd.n236 585
R2079 gnd.n6540 gnd.n236 585
R2080 gnd.n6278 gnd.n6277 585
R2081 gnd.n6277 gnd.n235 585
R2082 gnd.n6279 gnd.n243 585
R2083 gnd.n6532 gnd.n243 585
R2084 gnd.n6280 gnd.n248 585
R2085 gnd.n6527 gnd.n248 585
R2086 gnd.n6282 gnd.n6281 585
R2087 gnd.n6281 gnd.n247 585
R2088 gnd.n6283 gnd.n256 585
R2089 gnd.n6519 gnd.n256 585
R2090 gnd.n6284 gnd.n261 585
R2091 gnd.n6514 gnd.n261 585
R2092 gnd.n6286 gnd.n6285 585
R2093 gnd.n6287 gnd.n6286 585
R2094 gnd.n481 gnd.n269 585
R2095 gnd.n6502 gnd.n269 585
R2096 gnd.n6223 gnd.n6222 585
R2097 gnd.n6222 gnd.n6221 585
R2098 gnd.n6220 gnd.n277 585
R2099 gnd.n6493 gnd.n277 585
R2100 gnd.n6219 gnd.n6218 585
R2101 gnd.n6218 gnd.n6217 585
R2102 gnd.n483 gnd.n286 585
R2103 gnd.n6485 gnd.n286 585
R2104 gnd.n499 gnd.n498 585
R2105 gnd.n498 gnd.n497 585
R2106 gnd.n496 gnd.n295 585
R2107 gnd.n6477 gnd.n295 585
R2108 gnd.n495 gnd.n494 585
R2109 gnd.n494 gnd.n493 585
R2110 gnd.n485 gnd.n304 585
R2111 gnd.n6469 gnd.n304 585
R2112 gnd.n489 gnd.n488 585
R2113 gnd.n488 gnd.n487 585
R2114 gnd.n467 gnd.n313 585
R2115 gnd.n6461 gnd.n313 585
R2116 gnd.n6312 gnd.n6311 585
R2117 gnd.n6311 gnd.n6310 585
R2118 gnd.n6313 gnd.n321 585
R2119 gnd.n6453 gnd.n321 585
R2120 gnd.n6314 gnd.n464 585
R2121 gnd.n5150 gnd.n464 585
R2122 gnd.n6315 gnd.n329 585
R2123 gnd.n6445 gnd.n329 585
R2124 gnd.n5062 gnd.n5061 585
R2125 gnd.n5063 gnd.n5062 585
R2126 gnd.n1439 gnd.n1437 585
R2127 gnd.n1437 gnd.n1433 585
R2128 gnd.n4935 gnd.n4934 585
R2129 gnd.n4936 gnd.n4935 585
R2130 gnd.n4933 gnd.n1514 585
R2131 gnd.n1519 gnd.n1514 585
R2132 gnd.n4932 gnd.n4931 585
R2133 gnd.n4931 gnd.n4930 585
R2134 gnd.n1516 gnd.n1515 585
R2135 gnd.n4898 gnd.n1516 585
R2136 gnd.n4919 gnd.n4918 585
R2137 gnd.n4920 gnd.n4919 585
R2138 gnd.n4917 gnd.n1528 585
R2139 gnd.n1528 gnd.n1525 585
R2140 gnd.n4916 gnd.n4915 585
R2141 gnd.n4915 gnd.n4914 585
R2142 gnd.n1530 gnd.n1529 585
R2143 gnd.n1531 gnd.n1530 585
R2144 gnd.n4885 gnd.n4884 585
R2145 gnd.n4886 gnd.n4885 585
R2146 gnd.n4883 gnd.n1541 585
R2147 gnd.n4879 gnd.n1541 585
R2148 gnd.n4882 gnd.n4881 585
R2149 gnd.n4881 gnd.n4880 585
R2150 gnd.n1543 gnd.n1542 585
R2151 gnd.n4866 gnd.n1543 585
R2152 gnd.n4855 gnd.n1560 585
R2153 gnd.n1560 gnd.n1553 585
R2154 gnd.n4857 gnd.n4856 585
R2155 gnd.n4858 gnd.n4857 585
R2156 gnd.n4854 gnd.n1559 585
R2157 gnd.n1565 gnd.n1559 585
R2158 gnd.n4853 gnd.n4852 585
R2159 gnd.n4852 gnd.n4851 585
R2160 gnd.n1562 gnd.n1561 585
R2161 gnd.n4827 gnd.n1562 585
R2162 gnd.n4839 gnd.n4838 585
R2163 gnd.n4840 gnd.n4839 585
R2164 gnd.n4837 gnd.n1575 585
R2165 gnd.n1575 gnd.n1571 585
R2166 gnd.n4836 gnd.n4835 585
R2167 gnd.n4835 gnd.n4834 585
R2168 gnd.n1577 gnd.n1576 585
R2169 gnd.n1584 gnd.n1577 585
R2170 gnd.n4821 gnd.n4820 585
R2171 gnd.n4822 gnd.n4821 585
R2172 gnd.n4819 gnd.n1585 585
R2173 gnd.n1585 gnd.n1583 585
R2174 gnd.n4818 gnd.n4817 585
R2175 gnd.n4817 gnd.n4816 585
R2176 gnd.n1587 gnd.n1586 585
R2177 gnd.n4732 gnd.n1587 585
R2178 gnd.n4803 gnd.n4802 585
R2179 gnd.n4804 gnd.n4803 585
R2180 gnd.n4801 gnd.n1601 585
R2181 gnd.n1601 gnd.n1598 585
R2182 gnd.n4800 gnd.n4799 585
R2183 gnd.n4799 gnd.n4798 585
R2184 gnd.n1603 gnd.n1602 585
R2185 gnd.n4741 gnd.n1603 585
R2186 gnd.n4743 gnd.n1625 585
R2187 gnd.n4743 gnd.n4742 585
R2188 gnd.n4745 gnd.n4744 585
R2189 gnd.n4744 gnd.n1611 585
R2190 gnd.n4746 gnd.n1623 585
R2191 gnd.n4726 gnd.n1623 585
R2192 gnd.n4748 gnd.n4747 585
R2193 gnd.n4749 gnd.n4748 585
R2194 gnd.n1624 gnd.n1622 585
R2195 gnd.n1622 gnd.n1619 585
R2196 gnd.n4718 gnd.n4717 585
R2197 gnd.n4719 gnd.n4718 585
R2198 gnd.n4716 gnd.n1631 585
R2199 gnd.n1631 gnd.n1629 585
R2200 gnd.n4715 gnd.n4714 585
R2201 gnd.n4714 gnd.n4713 585
R2202 gnd.n1633 gnd.n1632 585
R2203 gnd.n1644 gnd.n1633 585
R2204 gnd.n4702 gnd.n4701 585
R2205 gnd.n4703 gnd.n4702 585
R2206 gnd.n4700 gnd.n1645 585
R2207 gnd.n4695 gnd.n1645 585
R2208 gnd.n4699 gnd.n4698 585
R2209 gnd.n4698 gnd.n4697 585
R2210 gnd.n1647 gnd.n1646 585
R2211 gnd.n1648 gnd.n1647 585
R2212 gnd.n4682 gnd.n4681 585
R2213 gnd.n4683 gnd.n4682 585
R2214 gnd.n4680 gnd.n1655 585
R2215 gnd.n4676 gnd.n1655 585
R2216 gnd.n4679 gnd.n4678 585
R2217 gnd.n4678 gnd.n4677 585
R2218 gnd.n1657 gnd.n1656 585
R2219 gnd.n4664 gnd.n1657 585
R2220 gnd.n4653 gnd.n1675 585
R2221 gnd.n1675 gnd.n1673 585
R2222 gnd.n4655 gnd.n4654 585
R2223 gnd.n4656 gnd.n4655 585
R2224 gnd.n4652 gnd.n1674 585
R2225 gnd.n1680 gnd.n1674 585
R2226 gnd.n4651 gnd.n4650 585
R2227 gnd.n4650 gnd.n4649 585
R2228 gnd.n1677 gnd.n1676 585
R2229 gnd.n4626 gnd.n1677 585
R2230 gnd.n4638 gnd.n4637 585
R2231 gnd.n4639 gnd.n4638 585
R2232 gnd.n4636 gnd.n1690 585
R2233 gnd.n1690 gnd.n1686 585
R2234 gnd.n4635 gnd.n4634 585
R2235 gnd.n4634 gnd.n4633 585
R2236 gnd.n1692 gnd.n1691 585
R2237 gnd.n1693 gnd.n1692 585
R2238 gnd.n4620 gnd.n4619 585
R2239 gnd.n4621 gnd.n4620 585
R2240 gnd.n4618 gnd.n1702 585
R2241 gnd.n4614 gnd.n1702 585
R2242 gnd.n4617 gnd.n4616 585
R2243 gnd.n4616 gnd.n4615 585
R2244 gnd.n1704 gnd.n1703 585
R2245 gnd.n1710 gnd.n1704 585
R2246 gnd.n4607 gnd.n4606 585
R2247 gnd.n4608 gnd.n4607 585
R2248 gnd.n4605 gnd.n1713 585
R2249 gnd.n1713 gnd.n1709 585
R2250 gnd.n4604 gnd.n4603 585
R2251 gnd.n4603 gnd.n4602 585
R2252 gnd.n1715 gnd.n1714 585
R2253 gnd.n1727 gnd.n1715 585
R2254 gnd.n4580 gnd.n4579 585
R2255 gnd.n4581 gnd.n4580 585
R2256 gnd.n4578 gnd.n1728 585
R2257 gnd.n4572 gnd.n1728 585
R2258 gnd.n4577 gnd.n4576 585
R2259 gnd.n4576 gnd.n4575 585
R2260 gnd.n1730 gnd.n1729 585
R2261 gnd.n1731 gnd.n1730 585
R2262 gnd.n4560 gnd.n4559 585
R2263 gnd.n4561 gnd.n4560 585
R2264 gnd.n4558 gnd.n1737 585
R2265 gnd.n4554 gnd.n1737 585
R2266 gnd.n4557 gnd.n4556 585
R2267 gnd.n4556 gnd.n4555 585
R2268 gnd.n1739 gnd.n1738 585
R2269 gnd.n4541 gnd.n1739 585
R2270 gnd.n4530 gnd.n1756 585
R2271 gnd.n1756 gnd.n1754 585
R2272 gnd.n4532 gnd.n4531 585
R2273 gnd.n4533 gnd.n4532 585
R2274 gnd.n4529 gnd.n1755 585
R2275 gnd.n1761 gnd.n1755 585
R2276 gnd.n4528 gnd.n4527 585
R2277 gnd.n4527 gnd.n4526 585
R2278 gnd.n1758 gnd.n1757 585
R2279 gnd.n4502 gnd.n1758 585
R2280 gnd.n4514 gnd.n4513 585
R2281 gnd.n4515 gnd.n4514 585
R2282 gnd.n4512 gnd.n1770 585
R2283 gnd.n1774 gnd.n1770 585
R2284 gnd.n4511 gnd.n4510 585
R2285 gnd.n4510 gnd.n4509 585
R2286 gnd.n1772 gnd.n1771 585
R2287 gnd.n1780 gnd.n1772 585
R2288 gnd.n4496 gnd.n4495 585
R2289 gnd.n4497 gnd.n4496 585
R2290 gnd.n4494 gnd.n1782 585
R2291 gnd.n4490 gnd.n1782 585
R2292 gnd.n4493 gnd.n4492 585
R2293 gnd.n4492 gnd.n4491 585
R2294 gnd.n1784 gnd.n1783 585
R2295 gnd.n1791 gnd.n1784 585
R2296 gnd.n4483 gnd.n4482 585
R2297 gnd.n4484 gnd.n4483 585
R2298 gnd.n4481 gnd.n1793 585
R2299 gnd.n1793 gnd.n1790 585
R2300 gnd.n4480 gnd.n4479 585
R2301 gnd.n4479 gnd.n4478 585
R2302 gnd.n1795 gnd.n1794 585
R2303 gnd.n1807 gnd.n1795 585
R2304 gnd.n4456 gnd.n4455 585
R2305 gnd.n4457 gnd.n4456 585
R2306 gnd.n4454 gnd.n1808 585
R2307 gnd.n4449 gnd.n1808 585
R2308 gnd.n4453 gnd.n4452 585
R2309 gnd.n4452 gnd.n4451 585
R2310 gnd.n1810 gnd.n1809 585
R2311 gnd.n4439 gnd.n1810 585
R2312 gnd.n4295 gnd.n4294 585
R2313 gnd.n4294 gnd.n1815 585
R2314 gnd.n4297 gnd.n4296 585
R2315 gnd.n4297 gnd.n1817 585
R2316 gnd.n4312 gnd.n4293 585
R2317 gnd.n4312 gnd.n4311 585
R2318 gnd.n4314 gnd.n4313 585
R2319 gnd.n4313 gnd.n1325 585
R2320 gnd.n4315 gnd.n4292 585
R2321 gnd.n4292 gnd.n1323 585
R2322 gnd.n4317 gnd.n4316 585
R2323 gnd.n4318 gnd.n4317 585
R2324 gnd.n1307 gnd.n1306 585
R2325 gnd.n1311 gnd.n1307 585
R2326 gnd.n5316 gnd.n5315 585
R2327 gnd.n5315 gnd.n5314 585
R2328 gnd.n5317 gnd.n1304 585
R2329 gnd.n1308 gnd.n1304 585
R2330 gnd.n5319 gnd.n5318 585
R2331 gnd.n5320 gnd.n5319 585
R2332 gnd.n1305 gnd.n1303 585
R2333 gnd.n1303 gnd.n1223 585
R2334 gnd.n4269 gnd.n1221 585
R2335 gnd.n5326 gnd.n1221 585
R2336 gnd.n4271 gnd.n4270 585
R2337 gnd.n4272 gnd.n4271 585
R2338 gnd.n4268 gnd.n4267 585
R2339 gnd.n4267 gnd.n1211 585
R2340 gnd.n1206 gnd.n1205 585
R2341 gnd.n5333 gnd.n1206 585
R2342 gnd.n5336 gnd.n5335 585
R2343 gnd.n5335 gnd.n5334 585
R2344 gnd.n5337 gnd.n1184 585
R2345 gnd.n1292 gnd.n1184 585
R2346 gnd.n5402 gnd.n5401 585
R2347 gnd.n5400 gnd.n1183 585
R2348 gnd.n5399 gnd.n1182 585
R2349 gnd.n5404 gnd.n1182 585
R2350 gnd.n5398 gnd.n5397 585
R2351 gnd.n5396 gnd.n5395 585
R2352 gnd.n5394 gnd.n5393 585
R2353 gnd.n5392 gnd.n5391 585
R2354 gnd.n5390 gnd.n5389 585
R2355 gnd.n5388 gnd.n5387 585
R2356 gnd.n5386 gnd.n5385 585
R2357 gnd.n5384 gnd.n5383 585
R2358 gnd.n5382 gnd.n5381 585
R2359 gnd.n5380 gnd.n5379 585
R2360 gnd.n5378 gnd.n5377 585
R2361 gnd.n5376 gnd.n5375 585
R2362 gnd.n5374 gnd.n5373 585
R2363 gnd.n5372 gnd.n5371 585
R2364 gnd.n5370 gnd.n5369 585
R2365 gnd.n5368 gnd.n5367 585
R2366 gnd.n5366 gnd.n5365 585
R2367 gnd.n5364 gnd.n5363 585
R2368 gnd.n5362 gnd.n5361 585
R2369 gnd.n5360 gnd.n5359 585
R2370 gnd.n5358 gnd.n5357 585
R2371 gnd.n5356 gnd.n5355 585
R2372 gnd.n5354 gnd.n5353 585
R2373 gnd.n5352 gnd.n5351 585
R2374 gnd.n5350 gnd.n5349 585
R2375 gnd.n5348 gnd.n5347 585
R2376 gnd.n5346 gnd.n5345 585
R2377 gnd.n5344 gnd.n5343 585
R2378 gnd.n5342 gnd.n1146 585
R2379 gnd.n5407 gnd.n5406 585
R2380 gnd.n1148 gnd.n1145 585
R2381 gnd.n1230 gnd.n1229 585
R2382 gnd.n1232 gnd.n1231 585
R2383 gnd.n1235 gnd.n1234 585
R2384 gnd.n1237 gnd.n1236 585
R2385 gnd.n1239 gnd.n1238 585
R2386 gnd.n1241 gnd.n1240 585
R2387 gnd.n1243 gnd.n1242 585
R2388 gnd.n1245 gnd.n1244 585
R2389 gnd.n1247 gnd.n1246 585
R2390 gnd.n1249 gnd.n1248 585
R2391 gnd.n1251 gnd.n1250 585
R2392 gnd.n1253 gnd.n1252 585
R2393 gnd.n1255 gnd.n1254 585
R2394 gnd.n1257 gnd.n1256 585
R2395 gnd.n1259 gnd.n1258 585
R2396 gnd.n1261 gnd.n1260 585
R2397 gnd.n1263 gnd.n1262 585
R2398 gnd.n1265 gnd.n1264 585
R2399 gnd.n1267 gnd.n1266 585
R2400 gnd.n1269 gnd.n1268 585
R2401 gnd.n1271 gnd.n1270 585
R2402 gnd.n1273 gnd.n1272 585
R2403 gnd.n1275 gnd.n1274 585
R2404 gnd.n1277 gnd.n1276 585
R2405 gnd.n1279 gnd.n1278 585
R2406 gnd.n1281 gnd.n1280 585
R2407 gnd.n1283 gnd.n1282 585
R2408 gnd.n1285 gnd.n1284 585
R2409 gnd.n1287 gnd.n1286 585
R2410 gnd.n1289 gnd.n1288 585
R2411 gnd.n1291 gnd.n1290 585
R2412 gnd.n4943 gnd.n4942 585
R2413 gnd.n4944 gnd.n1509 585
R2414 gnd.n4946 gnd.n4945 585
R2415 gnd.n4948 gnd.n1507 585
R2416 gnd.n4950 gnd.n4949 585
R2417 gnd.n4951 gnd.n1506 585
R2418 gnd.n4953 gnd.n4952 585
R2419 gnd.n4955 gnd.n1504 585
R2420 gnd.n4957 gnd.n4956 585
R2421 gnd.n4958 gnd.n1503 585
R2422 gnd.n4960 gnd.n4959 585
R2423 gnd.n4962 gnd.n1501 585
R2424 gnd.n4964 gnd.n4963 585
R2425 gnd.n4965 gnd.n1500 585
R2426 gnd.n4967 gnd.n4966 585
R2427 gnd.n4969 gnd.n1498 585
R2428 gnd.n4971 gnd.n4970 585
R2429 gnd.n4972 gnd.n1497 585
R2430 gnd.n4974 gnd.n4973 585
R2431 gnd.n4976 gnd.n1495 585
R2432 gnd.n4978 gnd.n4977 585
R2433 gnd.n4979 gnd.n1494 585
R2434 gnd.n4981 gnd.n4980 585
R2435 gnd.n4983 gnd.n1492 585
R2436 gnd.n4985 gnd.n4984 585
R2437 gnd.n4986 gnd.n1491 585
R2438 gnd.n4988 gnd.n4987 585
R2439 gnd.n4990 gnd.n1489 585
R2440 gnd.n4992 gnd.n4991 585
R2441 gnd.n4994 gnd.n1486 585
R2442 gnd.n4996 gnd.n4995 585
R2443 gnd.n4998 gnd.n1485 585
R2444 gnd.n4999 gnd.n1461 585
R2445 gnd.n5002 gnd.n435 585
R2446 gnd.n5004 gnd.n5003 585
R2447 gnd.n5006 gnd.n1483 585
R2448 gnd.n5008 gnd.n5007 585
R2449 gnd.n5010 gnd.n1480 585
R2450 gnd.n5012 gnd.n5011 585
R2451 gnd.n5014 gnd.n1478 585
R2452 gnd.n5016 gnd.n5015 585
R2453 gnd.n5017 gnd.n1477 585
R2454 gnd.n5019 gnd.n5018 585
R2455 gnd.n5021 gnd.n1475 585
R2456 gnd.n5023 gnd.n5022 585
R2457 gnd.n5024 gnd.n1474 585
R2458 gnd.n5026 gnd.n5025 585
R2459 gnd.n5028 gnd.n1472 585
R2460 gnd.n5030 gnd.n5029 585
R2461 gnd.n5031 gnd.n1471 585
R2462 gnd.n5033 gnd.n5032 585
R2463 gnd.n5035 gnd.n1469 585
R2464 gnd.n5037 gnd.n5036 585
R2465 gnd.n5038 gnd.n1468 585
R2466 gnd.n5040 gnd.n5039 585
R2467 gnd.n5042 gnd.n1466 585
R2468 gnd.n5044 gnd.n5043 585
R2469 gnd.n5045 gnd.n1465 585
R2470 gnd.n5047 gnd.n5046 585
R2471 gnd.n5049 gnd.n1463 585
R2472 gnd.n5051 gnd.n5050 585
R2473 gnd.n5052 gnd.n1462 585
R2474 gnd.n5054 gnd.n5053 585
R2475 gnd.n5056 gnd.n1459 585
R2476 gnd.n5058 gnd.n5057 585
R2477 gnd.n5059 gnd.n1438 585
R2478 gnd.n4940 gnd.n1435 585
R2479 gnd.n5063 gnd.n1435 585
R2480 gnd.n4939 gnd.n4938 585
R2481 gnd.n4938 gnd.n1433 585
R2482 gnd.n4937 gnd.n1510 585
R2483 gnd.n4937 gnd.n4936 585
R2484 gnd.n4894 gnd.n1511 585
R2485 gnd.n1519 gnd.n1511 585
R2486 gnd.n4895 gnd.n1517 585
R2487 gnd.n4930 gnd.n1517 585
R2488 gnd.n4897 gnd.n4896 585
R2489 gnd.n4898 gnd.n4897 585
R2490 gnd.n4893 gnd.n1527 585
R2491 gnd.n4920 gnd.n1527 585
R2492 gnd.n4892 gnd.n4891 585
R2493 gnd.n4891 gnd.n1525 585
R2494 gnd.n4890 gnd.n1532 585
R2495 gnd.n4914 gnd.n1532 585
R2496 gnd.n4889 gnd.n4888 585
R2497 gnd.n4888 gnd.n1531 585
R2498 gnd.n4887 gnd.n1538 585
R2499 gnd.n4887 gnd.n4886 585
R2500 gnd.n4862 gnd.n1539 585
R2501 gnd.n4879 gnd.n1539 585
R2502 gnd.n4863 gnd.n1545 585
R2503 gnd.n4880 gnd.n1545 585
R2504 gnd.n4865 gnd.n4864 585
R2505 gnd.n4866 gnd.n4865 585
R2506 gnd.n4861 gnd.n1555 585
R2507 gnd.n1555 gnd.n1553 585
R2508 gnd.n4860 gnd.n4859 585
R2509 gnd.n4859 gnd.n4858 585
R2510 gnd.n1557 gnd.n1556 585
R2511 gnd.n1565 gnd.n1557 585
R2512 gnd.n4826 gnd.n1563 585
R2513 gnd.n4851 gnd.n1563 585
R2514 gnd.n4829 gnd.n4828 585
R2515 gnd.n4828 gnd.n4827 585
R2516 gnd.n4830 gnd.n1573 585
R2517 gnd.n4840 gnd.n1573 585
R2518 gnd.n4831 gnd.n1580 585
R2519 gnd.n1580 gnd.n1571 585
R2520 gnd.n4833 gnd.n4832 585
R2521 gnd.n4834 gnd.n4833 585
R2522 gnd.n4825 gnd.n1579 585
R2523 gnd.n1584 gnd.n1579 585
R2524 gnd.n4824 gnd.n4823 585
R2525 gnd.n4823 gnd.n4822 585
R2526 gnd.n1582 gnd.n1581 585
R2527 gnd.n1583 gnd.n1582 585
R2528 gnd.n4731 gnd.n1590 585
R2529 gnd.n4816 gnd.n1590 585
R2530 gnd.n4734 gnd.n4733 585
R2531 gnd.n4733 gnd.n4732 585
R2532 gnd.n4735 gnd.n1600 585
R2533 gnd.n4804 gnd.n1600 585
R2534 gnd.n4737 gnd.n4736 585
R2535 gnd.n4736 gnd.n1598 585
R2536 gnd.n4738 gnd.n1604 585
R2537 gnd.n4798 gnd.n1604 585
R2538 gnd.n4740 gnd.n4739 585
R2539 gnd.n4741 gnd.n4740 585
R2540 gnd.n4730 gnd.n1626 585
R2541 gnd.n4742 gnd.n1626 585
R2542 gnd.n4729 gnd.n4728 585
R2543 gnd.n4728 gnd.n1611 585
R2544 gnd.n4727 gnd.n4724 585
R2545 gnd.n4727 gnd.n4726 585
R2546 gnd.n4723 gnd.n1621 585
R2547 gnd.n4749 gnd.n1621 585
R2548 gnd.n4722 gnd.n4721 585
R2549 gnd.n4721 gnd.n1619 585
R2550 gnd.n4720 gnd.n1627 585
R2551 gnd.n4720 gnd.n4719 585
R2552 gnd.n4688 gnd.n1628 585
R2553 gnd.n1629 gnd.n1628 585
R2554 gnd.n4689 gnd.n1634 585
R2555 gnd.n4713 gnd.n1634 585
R2556 gnd.n4691 gnd.n4690 585
R2557 gnd.n4690 gnd.n1644 585
R2558 gnd.n4692 gnd.n1643 585
R2559 gnd.n4703 gnd.n1643 585
R2560 gnd.n4694 gnd.n4693 585
R2561 gnd.n4695 gnd.n4694 585
R2562 gnd.n4687 gnd.n1649 585
R2563 gnd.n4697 gnd.n1649 585
R2564 gnd.n4686 gnd.n4685 585
R2565 gnd.n4685 gnd.n1648 585
R2566 gnd.n4684 gnd.n1651 585
R2567 gnd.n4684 gnd.n4683 585
R2568 gnd.n4660 gnd.n1652 585
R2569 gnd.n4676 gnd.n1652 585
R2570 gnd.n4661 gnd.n1659 585
R2571 gnd.n4677 gnd.n1659 585
R2572 gnd.n4663 gnd.n4662 585
R2573 gnd.n4664 gnd.n4663 585
R2574 gnd.n4659 gnd.n1668 585
R2575 gnd.n1673 gnd.n1668 585
R2576 gnd.n4658 gnd.n4657 585
R2577 gnd.n4657 gnd.n4656 585
R2578 gnd.n1670 gnd.n1669 585
R2579 gnd.n1680 gnd.n1670 585
R2580 gnd.n4625 gnd.n1678 585
R2581 gnd.n4649 gnd.n1678 585
R2582 gnd.n4628 gnd.n4627 585
R2583 gnd.n4627 gnd.n4626 585
R2584 gnd.n4629 gnd.n1688 585
R2585 gnd.n4639 gnd.n1688 585
R2586 gnd.n4630 gnd.n1697 585
R2587 gnd.n1697 gnd.n1686 585
R2588 gnd.n4632 gnd.n4631 585
R2589 gnd.n4633 gnd.n4632 585
R2590 gnd.n4624 gnd.n1696 585
R2591 gnd.n1696 gnd.n1693 585
R2592 gnd.n4623 gnd.n4622 585
R2593 gnd.n4622 gnd.n4621 585
R2594 gnd.n1699 gnd.n1698 585
R2595 gnd.n4614 gnd.n1699 585
R2596 gnd.n4613 gnd.n4612 585
R2597 gnd.n4615 gnd.n4613 585
R2598 gnd.n4611 gnd.n1706 585
R2599 gnd.n1710 gnd.n1706 585
R2600 gnd.n4610 gnd.n4609 585
R2601 gnd.n4609 gnd.n4608 585
R2602 gnd.n1708 gnd.n1707 585
R2603 gnd.n1709 gnd.n1708 585
R2604 gnd.n4566 gnd.n1717 585
R2605 gnd.n4602 gnd.n1717 585
R2606 gnd.n4568 gnd.n4567 585
R2607 gnd.n4567 gnd.n1727 585
R2608 gnd.n4569 gnd.n1726 585
R2609 gnd.n4581 gnd.n1726 585
R2610 gnd.n4571 gnd.n4570 585
R2611 gnd.n4572 gnd.n4571 585
R2612 gnd.n4565 gnd.n1732 585
R2613 gnd.n4575 gnd.n1732 585
R2614 gnd.n4564 gnd.n4563 585
R2615 gnd.n4563 gnd.n1731 585
R2616 gnd.n4562 gnd.n1734 585
R2617 gnd.n4562 gnd.n4561 585
R2618 gnd.n4537 gnd.n1735 585
R2619 gnd.n4554 gnd.n1735 585
R2620 gnd.n4538 gnd.n1741 585
R2621 gnd.n4555 gnd.n1741 585
R2622 gnd.n4540 gnd.n4539 585
R2623 gnd.n4541 gnd.n4540 585
R2624 gnd.n4536 gnd.n1750 585
R2625 gnd.n1754 gnd.n1750 585
R2626 gnd.n4535 gnd.n4534 585
R2627 gnd.n4534 gnd.n4533 585
R2628 gnd.n1752 gnd.n1751 585
R2629 gnd.n1761 gnd.n1752 585
R2630 gnd.n4501 gnd.n1759 585
R2631 gnd.n4526 gnd.n1759 585
R2632 gnd.n4504 gnd.n4503 585
R2633 gnd.n4503 gnd.n4502 585
R2634 gnd.n4505 gnd.n1768 585
R2635 gnd.n4515 gnd.n1768 585
R2636 gnd.n4506 gnd.n1776 585
R2637 gnd.n1776 gnd.n1774 585
R2638 gnd.n4508 gnd.n4507 585
R2639 gnd.n4509 gnd.n4508 585
R2640 gnd.n4500 gnd.n1775 585
R2641 gnd.n1780 gnd.n1775 585
R2642 gnd.n4499 gnd.n4498 585
R2643 gnd.n4498 gnd.n4497 585
R2644 gnd.n1778 gnd.n1777 585
R2645 gnd.n4490 gnd.n1778 585
R2646 gnd.n4489 gnd.n4488 585
R2647 gnd.n4491 gnd.n4489 585
R2648 gnd.n4487 gnd.n1787 585
R2649 gnd.n1791 gnd.n1787 585
R2650 gnd.n4486 gnd.n4485 585
R2651 gnd.n4485 gnd.n4484 585
R2652 gnd.n1789 gnd.n1788 585
R2653 gnd.n1790 gnd.n1789 585
R2654 gnd.n4443 gnd.n1797 585
R2655 gnd.n4478 gnd.n1797 585
R2656 gnd.n4445 gnd.n4444 585
R2657 gnd.n4444 gnd.n1807 585
R2658 gnd.n4446 gnd.n1806 585
R2659 gnd.n4457 gnd.n1806 585
R2660 gnd.n4448 gnd.n4447 585
R2661 gnd.n4449 gnd.n4448 585
R2662 gnd.n4442 gnd.n1811 585
R2663 gnd.n4451 gnd.n1811 585
R2664 gnd.n4441 gnd.n4440 585
R2665 gnd.n4440 gnd.n4439 585
R2666 gnd.n1814 gnd.n1813 585
R2667 gnd.n1815 gnd.n1814 585
R2668 gnd.n4308 gnd.n4300 585
R2669 gnd.n4300 gnd.n1817 585
R2670 gnd.n4310 gnd.n4309 585
R2671 gnd.n4311 gnd.n4310 585
R2672 gnd.n4307 gnd.n4299 585
R2673 gnd.n4299 gnd.n1325 585
R2674 gnd.n4306 gnd.n4305 585
R2675 gnd.n4305 gnd.n1323 585
R2676 gnd.n4304 gnd.n4291 585
R2677 gnd.n4318 gnd.n4291 585
R2678 gnd.n4303 gnd.n4302 585
R2679 gnd.n4302 gnd.n1311 585
R2680 gnd.n4301 gnd.n1309 585
R2681 gnd.n5314 gnd.n1309 585
R2682 gnd.n1301 gnd.n1300 585
R2683 gnd.n1308 gnd.n1301 585
R2684 gnd.n5322 gnd.n5321 585
R2685 gnd.n5321 gnd.n5320 585
R2686 gnd.n5323 gnd.n1226 585
R2687 gnd.n1226 gnd.n1223 585
R2688 gnd.n5325 gnd.n5324 585
R2689 gnd.n5326 gnd.n5325 585
R2690 gnd.n1299 gnd.n1225 585
R2691 gnd.n4272 gnd.n1225 585
R2692 gnd.n1298 gnd.n1297 585
R2693 gnd.n1297 gnd.n1211 585
R2694 gnd.n1296 gnd.n1209 585
R2695 gnd.n5333 gnd.n1209 585
R2696 gnd.n1295 gnd.n1208 585
R2697 gnd.n5334 gnd.n1208 585
R2698 gnd.n1294 gnd.n1293 585
R2699 gnd.n1293 gnd.n1292 585
R2700 gnd.n5496 gnd.n5495 585
R2701 gnd.n5495 gnd.n5494 585
R2702 gnd.n6202 gnd.n6200 585
R2703 gnd.n6202 gnd.n6201 585
R2704 gnd.n6207 gnd.n6203 585
R2705 gnd.n6203 gnd.n255 585
R2706 gnd.n6209 gnd.n6208 585
R2707 gnd.n6209 gnd.n260 585
R2708 gnd.n6210 gnd.n509 585
R2709 gnd.n6210 gnd.n271 585
R2710 gnd.n6212 gnd.n6211 585
R2711 gnd.n6211 gnd.n268 585
R2712 gnd.n6213 gnd.n504 585
R2713 gnd.n504 gnd.n279 585
R2714 gnd.n6215 gnd.n6214 585
R2715 gnd.n6216 gnd.n6215 585
R2716 gnd.n505 gnd.n503 585
R2717 gnd.n503 gnd.n288 585
R2718 gnd.n5136 gnd.n5135 585
R2719 gnd.n5136 gnd.n285 585
R2720 gnd.n5137 gnd.n5131 585
R2721 gnd.n5137 gnd.n297 585
R2722 gnd.n5139 gnd.n5138 585
R2723 gnd.n5138 gnd.n294 585
R2724 gnd.n5140 gnd.n5126 585
R2725 gnd.n5126 gnd.n306 585
R2726 gnd.n5142 gnd.n5141 585
R2727 gnd.n5142 gnd.n303 585
R2728 gnd.n5143 gnd.n5125 585
R2729 gnd.n5143 gnd.n315 585
R2730 gnd.n5145 gnd.n5144 585
R2731 gnd.n5144 gnd.n312 585
R2732 gnd.n5146 gnd.n5107 585
R2733 gnd.n5107 gnd.n323 585
R2734 gnd.n5148 gnd.n5147 585
R2735 gnd.n5149 gnd.n5148 585
R2736 gnd.n5108 gnd.n5106 585
R2737 gnd.n5106 gnd.n331 585
R2738 gnd.n5119 gnd.n5118 585
R2739 gnd.n5118 gnd.n328 585
R2740 gnd.n5117 gnd.n5110 585
R2741 gnd.n5117 gnd.n417 585
R2742 gnd.n5116 gnd.n5115 585
R2743 gnd.n5116 gnd.n384 585
R2744 gnd.n5111 gnd.n5074 585
R2745 gnd.n5180 gnd.n5074 585
R2746 gnd.n5182 gnd.n5073 585
R2747 gnd.n5182 gnd.n5181 585
R2748 gnd.n5184 gnd.n5183 585
R2749 gnd.n5183 gnd.n1421 585
R2750 gnd.n5185 gnd.n1420 585
R2751 gnd.n5197 gnd.n1420 585
R2752 gnd.n5186 gnd.n1428 585
R2753 gnd.n1428 gnd.n1419 585
R2754 gnd.n5188 gnd.n5187 585
R2755 gnd.n5189 gnd.n5188 585
R2756 gnd.n1429 gnd.n1427 585
R2757 gnd.n1436 gnd.n1427 585
R2758 gnd.n5066 gnd.n5065 585
R2759 gnd.n5065 gnd.n5064 585
R2760 gnd.n1432 gnd.n1431 585
R2761 gnd.n1513 gnd.n1432 585
R2762 gnd.n4928 gnd.n4927 585
R2763 gnd.n4929 gnd.n4928 585
R2764 gnd.n1521 gnd.n1520 585
R2765 gnd.n4898 gnd.n1520 585
R2766 gnd.n4923 gnd.n4922 585
R2767 gnd.n4922 gnd.n4921 585
R2768 gnd.n1524 gnd.n1523 585
R2769 gnd.n4913 gnd.n1524 585
R2770 gnd.n4875 gnd.n1548 585
R2771 gnd.n1548 gnd.n1540 585
R2772 gnd.n4877 gnd.n4876 585
R2773 gnd.n4878 gnd.n4877 585
R2774 gnd.n1549 gnd.n1547 585
R2775 gnd.n1547 gnd.n1544 585
R2776 gnd.n4870 gnd.n4869 585
R2777 gnd.n4869 gnd.n4868 585
R2778 gnd.n1552 gnd.n1551 585
R2779 gnd.n1558 gnd.n1552 585
R2780 gnd.n4849 gnd.n4848 585
R2781 gnd.n4850 gnd.n4849 585
R2782 gnd.n1567 gnd.n1566 585
R2783 gnd.n1574 gnd.n1566 585
R2784 gnd.n4844 gnd.n4843 585
R2785 gnd.n4843 gnd.n4842 585
R2786 gnd.n1570 gnd.n1569 585
R2787 gnd.n1578 gnd.n1570 585
R2788 gnd.n4812 gnd.n1593 585
R2789 gnd.n1593 gnd.t0 585
R2790 gnd.n4814 gnd.n4813 585
R2791 gnd.n4815 gnd.n4814 585
R2792 gnd.n1594 gnd.n1592 585
R2793 gnd.n1592 gnd.n1589 585
R2794 gnd.n4807 gnd.n4806 585
R2795 gnd.n4806 gnd.n4805 585
R2796 gnd.n1597 gnd.n1596 585
R2797 gnd.n4797 gnd.n1597 585
R2798 gnd.n4757 gnd.n1614 585
R2799 gnd.n4741 gnd.n1614 585
R2800 gnd.n4759 gnd.n4758 585
R2801 gnd.n4760 gnd.n4759 585
R2802 gnd.n1615 gnd.n1613 585
R2803 gnd.n4725 gnd.n1613 585
R2804 gnd.n4752 gnd.n4751 585
R2805 gnd.n4751 gnd.n4750 585
R2806 gnd.n1618 gnd.n1617 585
R2807 gnd.n1630 gnd.n1618 585
R2808 gnd.n4711 gnd.n4710 585
R2809 gnd.n4712 gnd.n4711 585
R2810 gnd.n1638 gnd.n1637 585
R2811 gnd.n4362 gnd.n1637 585
R2812 gnd.n4706 gnd.n4705 585
R2813 gnd.n4705 gnd.n4704 585
R2814 gnd.n1641 gnd.n1640 585
R2815 gnd.n4696 gnd.n1641 585
R2816 gnd.n4672 gnd.n1662 585
R2817 gnd.n1662 gnd.n1654 585
R2818 gnd.n4674 gnd.n4673 585
R2819 gnd.n4675 gnd.n4674 585
R2820 gnd.n1663 gnd.n1661 585
R2821 gnd.n1661 gnd.n1658 585
R2822 gnd.n4667 gnd.n4666 585
R2823 gnd.n4666 gnd.n4665 585
R2824 gnd.n1666 gnd.n1665 585
R2825 gnd.n1672 gnd.n1666 585
R2826 gnd.n4647 gnd.n4646 585
R2827 gnd.n4648 gnd.n4647 585
R2828 gnd.n1682 gnd.n1681 585
R2829 gnd.n1689 gnd.n1681 585
R2830 gnd.n4642 gnd.n4641 585
R2831 gnd.n4641 gnd.n4640 585
R2832 gnd.n1685 gnd.n1684 585
R2833 gnd.n4633 gnd.n1685 585
R2834 gnd.n4594 gnd.n4593 585
R2835 gnd.n4594 gnd.n1701 585
R2836 gnd.n4595 gnd.n4590 585
R2837 gnd.n4595 gnd.n1700 585
R2838 gnd.n4597 gnd.n4596 585
R2839 gnd.n4596 gnd.n1705 585
R2840 gnd.n4598 gnd.n1720 585
R2841 gnd.n1720 gnd.n1712 585
R2842 gnd.n4600 gnd.n4599 585
R2843 gnd.n4601 gnd.n4600 585
R2844 gnd.n1721 gnd.n1719 585
R2845 gnd.n1719 gnd.n1716 585
R2846 gnd.n4584 gnd.n4583 585
R2847 gnd.n4583 gnd.n4582 585
R2848 gnd.n1724 gnd.n1723 585
R2849 gnd.n4574 gnd.n1724 585
R2850 gnd.n4550 gnd.n1744 585
R2851 gnd.n1744 gnd.n1736 585
R2852 gnd.n4552 gnd.n4551 585
R2853 gnd.n4553 gnd.n4552 585
R2854 gnd.n1745 gnd.n1743 585
R2855 gnd.n1743 gnd.n1740 585
R2856 gnd.n4545 gnd.n4544 585
R2857 gnd.n4544 gnd.n4543 585
R2858 gnd.n1748 gnd.n1747 585
R2859 gnd.n1753 gnd.n1748 585
R2860 gnd.n4524 gnd.n4523 585
R2861 gnd.n4525 gnd.n4524 585
R2862 gnd.n1763 gnd.n1762 585
R2863 gnd.n1769 gnd.n1762 585
R2864 gnd.n4519 gnd.n4518 585
R2865 gnd.n4518 gnd.n4517 585
R2866 gnd.n1766 gnd.n1765 585
R2867 gnd.n4509 gnd.n1766 585
R2868 gnd.n4471 gnd.n4470 585
R2869 gnd.n4471 gnd.n1781 585
R2870 gnd.n4472 gnd.n4467 585
R2871 gnd.n4472 gnd.n1779 585
R2872 gnd.n4474 gnd.n4473 585
R2873 gnd.n4473 gnd.n1786 585
R2874 gnd.n4475 gnd.n1800 585
R2875 gnd.n1800 gnd.n1792 585
R2876 gnd.n4477 gnd.n4476 585
R2877 gnd.t266 gnd.n4477 585
R2878 gnd.n1801 gnd.n1799 585
R2879 gnd.n1799 gnd.n1796 585
R2880 gnd.n4461 gnd.n4460 585
R2881 gnd.n4460 gnd.n4459 585
R2882 gnd.n1804 gnd.n1803 585
R2883 gnd.n4450 gnd.n1804 585
R2884 gnd.n4437 gnd.n4436 585
R2885 gnd.n4438 gnd.n4437 585
R2886 gnd.n4432 gnd.n4431 585
R2887 gnd.n4431 gnd.n4430 585
R2888 gnd.n1322 gnd.n1321 585
R2889 gnd.n4298 gnd.n1322 585
R2890 gnd.n5309 gnd.n5308 585
R2891 gnd.n5308 gnd.n5307 585
R2892 gnd.n5310 gnd.n1314 585
R2893 gnd.n4319 gnd.n1314 585
R2894 gnd.n5312 gnd.n5311 585
R2895 gnd.n5313 gnd.n5312 585
R2896 gnd.n1315 gnd.n1313 585
R2897 gnd.n1313 gnd.n1302 585
R2898 gnd.n1220 gnd.n1219 585
R2899 gnd.n4284 gnd.n1220 585
R2900 gnd.n5328 gnd.n5327 585
R2901 gnd.n5327 gnd.n5326 585
R2902 gnd.n5329 gnd.n1214 585
R2903 gnd.n4273 gnd.n1214 585
R2904 gnd.n5331 gnd.n5330 585
R2905 gnd.n5332 gnd.n5331 585
R2906 gnd.n1215 gnd.n1213 585
R2907 gnd.n1213 gnd.n1207 585
R2908 gnd.n4245 gnd.n4244 585
R2909 gnd.n4245 gnd.n1181 585
R2910 gnd.n4247 gnd.n4246 585
R2911 gnd.n4246 gnd.n1149 585
R2912 gnd.n4248 gnd.n1842 585
R2913 gnd.n1842 gnd.n1839 585
R2914 gnd.n4250 gnd.n4249 585
R2915 gnd.n4251 gnd.n4250 585
R2916 gnd.n1843 gnd.n1841 585
R2917 gnd.n1841 gnd.n1838 585
R2918 gnd.n4236 gnd.n4235 585
R2919 gnd.n4235 gnd.n4234 585
R2920 gnd.n1846 gnd.n1845 585
R2921 gnd.n1847 gnd.n1846 585
R2922 gnd.n4181 gnd.n4180 585
R2923 gnd.n4180 gnd.n1106 585
R2924 gnd.n4182 gnd.n1983 585
R2925 gnd.n1983 gnd.n1095 585
R2926 gnd.n4184 gnd.n4183 585
R2927 gnd.n4185 gnd.n4184 585
R2928 gnd.n1984 gnd.n1982 585
R2929 gnd.n1982 gnd.n1088 585
R2930 gnd.n4174 gnd.n4173 585
R2931 gnd.n4173 gnd.n1085 585
R2932 gnd.n4172 gnd.n1986 585
R2933 gnd.n4172 gnd.n1077 585
R2934 gnd.n4171 gnd.n4170 585
R2935 gnd.n4171 gnd.n1074 585
R2936 gnd.n1988 gnd.n1987 585
R2937 gnd.n1987 gnd.n1066 585
R2938 gnd.n4166 gnd.n4165 585
R2939 gnd.n4165 gnd.n1063 585
R2940 gnd.n4164 gnd.n1990 585
R2941 gnd.n4164 gnd.n4163 585
R2942 gnd.n4052 gnd.n1991 585
R2943 gnd.n1991 gnd.n1053 585
R2944 gnd.n4053 gnd.n2008 585
R2945 gnd.n2008 gnd.n1045 585
R2946 gnd.n4055 gnd.n4054 585
R2947 gnd.n4056 gnd.n4055 585
R2948 gnd.n2009 gnd.n2007 585
R2949 gnd.n2007 gnd.n1035 585
R2950 gnd.n4046 gnd.n4045 585
R2951 gnd.n4045 gnd.n1032 585
R2952 gnd.n4044 gnd.n2011 585
R2953 gnd.n4044 gnd.n1024 585
R2954 gnd.n4043 gnd.n4042 585
R2955 gnd.n4043 gnd.n1021 585
R2956 gnd.n4033 gnd.n4032 585
R2957 gnd.n4032 gnd.n4031 585
R2958 gnd.n4038 gnd.n4037 585
R2959 gnd.n4037 gnd.n1010 585
R2960 gnd.n4036 gnd.n997 585
R2961 gnd.n1001 gnd.n997 585
R2962 gnd.n5196 gnd.n5195 585
R2963 gnd.n5197 gnd.n5196 585
R2964 gnd.n1423 gnd.n1422 585
R2965 gnd.n1422 gnd.n1419 585
R2966 gnd.n5191 gnd.n5190 585
R2967 gnd.n5190 gnd.n5189 585
R2968 gnd.n1426 gnd.n1425 585
R2969 gnd.n1436 gnd.n1426 585
R2970 gnd.n4901 gnd.n1434 585
R2971 gnd.n5064 gnd.n1434 585
R2972 gnd.n4904 gnd.n4900 585
R2973 gnd.n4900 gnd.n1513 585
R2974 gnd.n4905 gnd.n1518 585
R2975 gnd.n4929 gnd.n1518 585
R2976 gnd.n4906 gnd.n4899 585
R2977 gnd.n4899 gnd.n4898 585
R2978 gnd.n1535 gnd.n1526 585
R2979 gnd.n4921 gnd.n1526 585
R2980 gnd.n4911 gnd.n4910 585
R2981 gnd.n4913 gnd.n4911 585
R2982 gnd.n1534 gnd.n1533 585
R2983 gnd.n1540 gnd.n1533 585
R2984 gnd.n4777 gnd.n1546 585
R2985 gnd.n4878 gnd.n1546 585
R2986 gnd.n4778 gnd.n4775 585
R2987 gnd.n4775 gnd.n1544 585
R2988 gnd.n4779 gnd.n1554 585
R2989 gnd.n4868 gnd.n1554 585
R2990 gnd.n4773 gnd.n4772 585
R2991 gnd.n4772 gnd.n1558 585
R2992 gnd.n4783 gnd.n1564 585
R2993 gnd.n4850 gnd.n1564 585
R2994 gnd.n4784 gnd.n4771 585
R2995 gnd.n4771 gnd.n1574 585
R2996 gnd.n4785 gnd.n1572 585
R2997 gnd.n4842 gnd.n1572 585
R2998 gnd.n4769 gnd.n4768 585
R2999 gnd.n4768 gnd.n1578 585
R3000 gnd.n4789 gnd.n4767 585
R3001 gnd.n4767 gnd.t0 585
R3002 gnd.n4790 gnd.n1591 585
R3003 gnd.n4815 gnd.n1591 585
R3004 gnd.n4791 gnd.n4766 585
R3005 gnd.n4766 gnd.n1589 585
R3006 gnd.n1607 gnd.n1599 585
R3007 gnd.n4805 gnd.n1599 585
R3008 gnd.n4796 gnd.n4795 585
R3009 gnd.n4797 gnd.n4796 585
R3010 gnd.n1606 gnd.n1605 585
R3011 gnd.n4741 gnd.n1605 585
R3012 gnd.n4762 gnd.n4761 585
R3013 gnd.n4761 gnd.n4760 585
R3014 gnd.n1610 gnd.n1609 585
R3015 gnd.n4725 gnd.n1610 585
R3016 gnd.n4365 gnd.n1620 585
R3017 gnd.n4750 gnd.n1620 585
R3018 gnd.n4368 gnd.n4364 585
R3019 gnd.n4364 gnd.n1630 585
R3020 gnd.n4369 gnd.n1635 585
R3021 gnd.n4712 gnd.n1635 585
R3022 gnd.n4370 gnd.n4363 585
R3023 gnd.n4363 gnd.n4362 585
R3024 gnd.n4360 gnd.n1642 585
R3025 gnd.n4704 gnd.n1642 585
R3026 gnd.n4374 gnd.n1650 585
R3027 gnd.n4696 gnd.n1650 585
R3028 gnd.n4375 gnd.n4359 585
R3029 gnd.n4359 gnd.n1654 585
R3030 gnd.n4376 gnd.n1660 585
R3031 gnd.n4675 gnd.n1660 585
R3032 gnd.n4357 gnd.n4356 585
R3033 gnd.n4356 gnd.n1658 585
R3034 gnd.n4380 gnd.n1667 585
R3035 gnd.n4665 gnd.n1667 585
R3036 gnd.n4381 gnd.n4355 585
R3037 gnd.n4355 gnd.n1672 585
R3038 gnd.n4382 gnd.n1679 585
R3039 gnd.n4648 gnd.n1679 585
R3040 gnd.n4353 gnd.n4352 585
R3041 gnd.n4352 gnd.n1689 585
R3042 gnd.n4386 gnd.n1687 585
R3043 gnd.n4640 gnd.n1687 585
R3044 gnd.n4387 gnd.n1694 585
R3045 gnd.n4633 gnd.n1694 585
R3046 gnd.n4388 gnd.n4351 585
R3047 gnd.n4351 gnd.n1701 585
R3048 gnd.n4350 gnd.n4348 585
R3049 gnd.n4350 gnd.n1700 585
R3050 gnd.n4392 gnd.n4347 585
R3051 gnd.n4347 gnd.n1705 585
R3052 gnd.n4393 gnd.n4346 585
R3053 gnd.n4346 gnd.n1712 585
R3054 gnd.n4394 gnd.n1718 585
R3055 gnd.n4601 gnd.n1718 585
R3056 gnd.n4344 gnd.n4343 585
R3057 gnd.n4343 gnd.n1716 585
R3058 gnd.n4398 gnd.n1725 585
R3059 gnd.n4582 gnd.n1725 585
R3060 gnd.n4399 gnd.n1733 585
R3061 gnd.n4574 gnd.n1733 585
R3062 gnd.n4400 gnd.n4342 585
R3063 gnd.n4342 gnd.n1736 585
R3064 gnd.n4340 gnd.n1742 585
R3065 gnd.n4553 gnd.n1742 585
R3066 gnd.n4404 gnd.n4339 585
R3067 gnd.n4339 gnd.n1740 585
R3068 gnd.n4405 gnd.n1749 585
R3069 gnd.n4543 gnd.n1749 585
R3070 gnd.n4406 gnd.n4338 585
R3071 gnd.n4338 gnd.n1753 585
R3072 gnd.n4336 gnd.n1760 585
R3073 gnd.n4525 gnd.n1760 585
R3074 gnd.n4410 gnd.n4335 585
R3075 gnd.n4335 gnd.n1769 585
R3076 gnd.n4411 gnd.n1767 585
R3077 gnd.n4517 gnd.n1767 585
R3078 gnd.n4412 gnd.n1773 585
R3079 gnd.n4509 gnd.n1773 585
R3080 gnd.n4333 gnd.n4332 585
R3081 gnd.n4332 gnd.n1781 585
R3082 gnd.n4416 gnd.n4331 585
R3083 gnd.n4331 gnd.n1779 585
R3084 gnd.n4417 gnd.n4330 585
R3085 gnd.n4330 gnd.n1786 585
R3086 gnd.n4418 gnd.n4329 585
R3087 gnd.n4329 gnd.n1792 585
R3088 gnd.n4327 gnd.n1798 585
R3089 gnd.t266 gnd.n1798 585
R3090 gnd.n4422 gnd.n4326 585
R3091 gnd.n4326 gnd.n1796 585
R3092 gnd.n4423 gnd.n1805 585
R3093 gnd.n4459 gnd.n1805 585
R3094 gnd.n4424 gnd.n1812 585
R3095 gnd.n4450 gnd.n1812 585
R3096 gnd.n1820 gnd.n1816 585
R3097 gnd.n4438 gnd.n1816 585
R3098 gnd.n4429 gnd.n4428 585
R3099 gnd.n4430 gnd.n4429 585
R3100 gnd.n1819 gnd.n1818 585
R3101 gnd.n4298 gnd.n1818 585
R3102 gnd.n4322 gnd.n1324 585
R3103 gnd.n5307 gnd.n1324 585
R3104 gnd.n4321 gnd.n4320 585
R3105 gnd.n4320 gnd.n4319 585
R3106 gnd.n4290 gnd.n1310 585
R3107 gnd.n5313 gnd.n1310 585
R3108 gnd.n1825 gnd.n1822 585
R3109 gnd.n1825 gnd.n1302 585
R3110 gnd.n4286 gnd.n4285 585
R3111 gnd.n4285 gnd.n4284 585
R3112 gnd.n1824 gnd.n1222 585
R3113 gnd.n5326 gnd.n1222 585
R3114 gnd.n4266 gnd.n4265 585
R3115 gnd.n4273 gnd.n4266 585
R3116 gnd.n1831 gnd.n1210 585
R3117 gnd.n5332 gnd.n1210 585
R3118 gnd.n4261 gnd.n4260 585
R3119 gnd.n4260 gnd.n1207 585
R3120 gnd.n4259 gnd.n1833 585
R3121 gnd.n4259 gnd.n1181 585
R3122 gnd.n4258 gnd.n4257 585
R3123 gnd.n4258 gnd.n1149 585
R3124 gnd.n1835 gnd.n1834 585
R3125 gnd.n1839 gnd.n1834 585
R3126 gnd.n4253 gnd.n4252 585
R3127 gnd.n4252 gnd.n4251 585
R3128 gnd.n1906 gnd.n1837 585
R3129 gnd.n1920 gnd.n1919 585
R3130 gnd.n1922 gnd.n1921 585
R3131 gnd.n1901 gnd.n1900 585
R3132 gnd.n1931 gnd.n1902 585
R3133 gnd.n1934 gnd.n1933 585
R3134 gnd.n1932 gnd.n1894 585
R3135 gnd.n1944 gnd.n1943 585
R3136 gnd.n1946 gnd.n1945 585
R3137 gnd.n1889 gnd.n1888 585
R3138 gnd.n1955 gnd.n1890 585
R3139 gnd.n1958 gnd.n1957 585
R3140 gnd.n1956 gnd.n1882 585
R3141 gnd.n1968 gnd.n1967 585
R3142 gnd.n1970 gnd.n1969 585
R3143 gnd.n1877 gnd.n1876 585
R3144 gnd.n4192 gnd.n1878 585
R3145 gnd.n4194 gnd.n4193 585
R3146 gnd.n4196 gnd.n4195 585
R3147 gnd.n1872 gnd.n1871 585
R3148 gnd.n4201 gnd.n1873 585
R3149 gnd.n4203 gnd.n4202 585
R3150 gnd.n4205 gnd.n4204 585
R3151 gnd.n1868 gnd.n1867 585
R3152 gnd.n4209 gnd.n1869 585
R3153 gnd.n4212 gnd.n4211 585
R3154 gnd.n4214 gnd.n4213 585
R3155 gnd.n1863 gnd.n1862 585
R3156 gnd.n4233 gnd.n4232 585
R3157 gnd.n4234 gnd.n4233 585
R3158 gnd.n5199 gnd.n5198 585
R3159 gnd.n5198 gnd.n5197 585
R3160 gnd.n1417 gnd.n1415 585
R3161 gnd.n1419 gnd.n1417 585
R3162 gnd.n5203 gnd.n1414 585
R3163 gnd.n5189 gnd.n1414 585
R3164 gnd.n5204 gnd.n1413 585
R3165 gnd.n1436 gnd.n1413 585
R3166 gnd.n5205 gnd.n1412 585
R3167 gnd.n5064 gnd.n1412 585
R3168 gnd.n1512 gnd.n1410 585
R3169 gnd.n1513 gnd.n1512 585
R3170 gnd.n5209 gnd.n1409 585
R3171 gnd.n4929 gnd.n1409 585
R3172 gnd.n5210 gnd.n1408 585
R3173 gnd.n4898 gnd.n1408 585
R3174 gnd.n5211 gnd.n1407 585
R3175 gnd.n4921 gnd.n1407 585
R3176 gnd.n4912 gnd.n1405 585
R3177 gnd.n4913 gnd.n4912 585
R3178 gnd.n5215 gnd.n1404 585
R3179 gnd.n1540 gnd.n1404 585
R3180 gnd.n5216 gnd.n1403 585
R3181 gnd.n4878 gnd.n1403 585
R3182 gnd.n5217 gnd.n1402 585
R3183 gnd.n1544 gnd.n1402 585
R3184 gnd.n4867 gnd.n1400 585
R3185 gnd.n4868 gnd.n4867 585
R3186 gnd.n5221 gnd.n1399 585
R3187 gnd.n1558 gnd.n1399 585
R3188 gnd.n5222 gnd.n1398 585
R3189 gnd.n4850 gnd.n1398 585
R3190 gnd.n5223 gnd.n1397 585
R3191 gnd.n1574 gnd.n1397 585
R3192 gnd.n4841 gnd.n1395 585
R3193 gnd.n4842 gnd.n4841 585
R3194 gnd.n5227 gnd.n1394 585
R3195 gnd.n1578 gnd.n1394 585
R3196 gnd.n5228 gnd.n1393 585
R3197 gnd.t0 gnd.n1393 585
R3198 gnd.n5229 gnd.n1392 585
R3199 gnd.n4815 gnd.n1392 585
R3200 gnd.n1588 gnd.n1390 585
R3201 gnd.n1589 gnd.n1588 585
R3202 gnd.n5233 gnd.n1389 585
R3203 gnd.n4805 gnd.n1389 585
R3204 gnd.n5234 gnd.n1388 585
R3205 gnd.n4797 gnd.n1388 585
R3206 gnd.n5235 gnd.n1387 585
R3207 gnd.n4741 gnd.n1387 585
R3208 gnd.n1612 gnd.n1385 585
R3209 gnd.n4760 gnd.n1612 585
R3210 gnd.n5239 gnd.n1384 585
R3211 gnd.n4725 gnd.n1384 585
R3212 gnd.n5240 gnd.n1383 585
R3213 gnd.n4750 gnd.n1383 585
R3214 gnd.n5241 gnd.n1382 585
R3215 gnd.n1630 gnd.n1382 585
R3216 gnd.n1636 gnd.n1380 585
R3217 gnd.n4712 gnd.n1636 585
R3218 gnd.n5245 gnd.n1379 585
R3219 gnd.n4362 gnd.n1379 585
R3220 gnd.n5246 gnd.n1378 585
R3221 gnd.n4704 gnd.n1378 585
R3222 gnd.n5247 gnd.n1377 585
R3223 gnd.n4696 gnd.n1377 585
R3224 gnd.n1653 gnd.n1375 585
R3225 gnd.n1654 gnd.n1653 585
R3226 gnd.n5251 gnd.n1374 585
R3227 gnd.n4675 gnd.n1374 585
R3228 gnd.n5252 gnd.n1373 585
R3229 gnd.n1658 gnd.n1373 585
R3230 gnd.n5253 gnd.n1372 585
R3231 gnd.n4665 gnd.n1372 585
R3232 gnd.n1671 gnd.n1370 585
R3233 gnd.n1672 gnd.n1671 585
R3234 gnd.n5257 gnd.n1369 585
R3235 gnd.n4648 gnd.n1369 585
R3236 gnd.n5258 gnd.n1368 585
R3237 gnd.n1689 gnd.n1368 585
R3238 gnd.n5259 gnd.n1367 585
R3239 gnd.n4640 gnd.n1367 585
R3240 gnd.n1695 gnd.n1365 585
R3241 gnd.n4633 gnd.n1695 585
R3242 gnd.n5263 gnd.n1364 585
R3243 gnd.n1701 gnd.n1364 585
R3244 gnd.n5264 gnd.n1363 585
R3245 gnd.n1700 gnd.n1363 585
R3246 gnd.n5265 gnd.n1362 585
R3247 gnd.n1705 gnd.n1362 585
R3248 gnd.n1711 gnd.n1360 585
R3249 gnd.n1712 gnd.n1711 585
R3250 gnd.n5269 gnd.n1359 585
R3251 gnd.n4601 gnd.n1359 585
R3252 gnd.n5270 gnd.n1358 585
R3253 gnd.n1716 gnd.n1358 585
R3254 gnd.n5271 gnd.n1357 585
R3255 gnd.n4582 gnd.n1357 585
R3256 gnd.n4573 gnd.n1355 585
R3257 gnd.n4574 gnd.n4573 585
R3258 gnd.n5275 gnd.n1354 585
R3259 gnd.n1736 gnd.n1354 585
R3260 gnd.n5276 gnd.n1353 585
R3261 gnd.n4553 gnd.n1353 585
R3262 gnd.n5277 gnd.n1352 585
R3263 gnd.n1740 gnd.n1352 585
R3264 gnd.n4542 gnd.n1350 585
R3265 gnd.n4543 gnd.n4542 585
R3266 gnd.n5281 gnd.n1349 585
R3267 gnd.n1753 gnd.n1349 585
R3268 gnd.n5282 gnd.n1348 585
R3269 gnd.n4525 gnd.n1348 585
R3270 gnd.n5283 gnd.n1347 585
R3271 gnd.n1769 gnd.n1347 585
R3272 gnd.n4516 gnd.n1345 585
R3273 gnd.n4517 gnd.n4516 585
R3274 gnd.n5287 gnd.n1344 585
R3275 gnd.n4509 gnd.n1344 585
R3276 gnd.n5288 gnd.n1343 585
R3277 gnd.n1781 gnd.n1343 585
R3278 gnd.n5289 gnd.n1342 585
R3279 gnd.n1779 gnd.n1342 585
R3280 gnd.n1785 gnd.n1340 585
R3281 gnd.n1786 gnd.n1785 585
R3282 gnd.n5293 gnd.n1339 585
R3283 gnd.n1792 gnd.n1339 585
R3284 gnd.n5294 gnd.n1338 585
R3285 gnd.t266 gnd.n1338 585
R3286 gnd.n5295 gnd.n1337 585
R3287 gnd.n1796 gnd.n1337 585
R3288 gnd.n4458 gnd.n1335 585
R3289 gnd.n4459 gnd.n4458 585
R3290 gnd.n5299 gnd.n1334 585
R3291 gnd.n4450 gnd.n1334 585
R3292 gnd.n5300 gnd.n1333 585
R3293 gnd.n4438 gnd.n1333 585
R3294 gnd.n5301 gnd.n1332 585
R3295 gnd.n4430 gnd.n1332 585
R3296 gnd.n1329 gnd.n1327 585
R3297 gnd.n4298 gnd.n1327 585
R3298 gnd.n5306 gnd.n5305 585
R3299 gnd.n5307 gnd.n5306 585
R3300 gnd.n1328 gnd.n1326 585
R3301 gnd.n4319 gnd.n1326 585
R3302 gnd.n4278 gnd.n1312 585
R3303 gnd.n5313 gnd.n1312 585
R3304 gnd.n1828 gnd.n1826 585
R3305 gnd.n1826 gnd.n1302 585
R3306 gnd.n4283 gnd.n4282 585
R3307 gnd.n4284 gnd.n4283 585
R3308 gnd.n1827 gnd.n1224 585
R3309 gnd.n5326 gnd.n1224 585
R3310 gnd.n4275 gnd.n4274 585
R3311 gnd.n4274 gnd.n4273 585
R3312 gnd.n1830 gnd.n1212 585
R3313 gnd.n5332 gnd.n1212 585
R3314 gnd.n4223 gnd.n4222 585
R3315 gnd.n4222 gnd.n1207 585
R3316 gnd.n4221 gnd.n4220 585
R3317 gnd.n4221 gnd.n1181 585
R3318 gnd.n4227 gnd.n4219 585
R3319 gnd.n4219 gnd.n1149 585
R3320 gnd.n4228 gnd.n4218 585
R3321 gnd.n4218 gnd.n1839 585
R3322 gnd.n4229 gnd.n1840 585
R3323 gnd.n4251 gnd.n1840 585
R3324 gnd.n5095 gnd.n1418 585
R3325 gnd.n5181 gnd.n1418 585
R3326 gnd.n5178 gnd.n5177 585
R3327 gnd.n5094 gnd.n5093 585
R3328 gnd.n5173 gnd.n5172 585
R3329 gnd.n5170 gnd.n5169 585
R3330 gnd.n5168 gnd.n5167 585
R3331 gnd.n5161 gnd.n5099 585
R3332 gnd.n5163 gnd.n5162 585
R3333 gnd.n5160 gnd.n5159 585
R3334 gnd.n5158 gnd.n5157 585
R3335 gnd.n5103 gnd.n5102 585
R3336 gnd.n5101 gnd.n381 585
R3337 gnd.n6395 gnd.n380 585
R3338 gnd.n6396 gnd.n379 585
R3339 gnd.n5086 gnd.n371 585
R3340 gnd.n6403 gnd.n370 585
R3341 gnd.n6404 gnd.n369 585
R3342 gnd.n5083 gnd.n363 585
R3343 gnd.n6411 gnd.n362 585
R3344 gnd.n6412 gnd.n361 585
R3345 gnd.n5081 gnd.n355 585
R3346 gnd.n6419 gnd.n354 585
R3347 gnd.n6420 gnd.n353 585
R3348 gnd.n5078 gnd.n347 585
R3349 gnd.n6427 gnd.n346 585
R3350 gnd.n6428 gnd.n345 585
R3351 gnd.n5076 gnd.n339 585
R3352 gnd.n6435 gnd.n338 585
R3353 gnd.n6436 gnd.n337 585
R3354 gnd.n5062 gnd.n1438 506.916
R3355 gnd.n4942 gnd.n1435 506.916
R3356 gnd.n1293 gnd.n1291 506.916
R3357 gnd.n5402 gnd.n1184 506.916
R3358 gnd.n1227 gnd.t165 389.64
R3359 gnd.n1487 gnd.t98 389.64
R3360 gnd.n5339 gnd.t116 389.64
R3361 gnd.n1481 gnd.t152 389.64
R3362 gnd.n5662 gnd.n826 371.755
R3363 gnd.n1865 gnd.t145 371.625
R3364 gnd.n6635 gnd.t133 371.625
R3365 gnd.n375 gnd.t123 371.625
R3366 gnd.n1975 gnd.t139 371.625
R3367 gnd.n438 gnd.t120 371.625
R3368 gnd.n460 gnd.t87 371.625
R3369 gnd.n156 gnd.t73 371.625
R3370 gnd.n6727 gnd.t102 371.625
R3371 gnd.n3727 gnd.t171 371.625
R3372 gnd.n3749 gnd.t162 371.625
R3373 gnd.n3599 gnd.t158 371.625
R3374 gnd.n4081 gnd.t94 371.625
R3375 gnd.n1141 gnd.t136 371.625
R3376 gnd.n5097 gnd.t129 371.625
R3377 gnd.n2589 gnd.t80 323.425
R3378 gnd.n2159 gnd.t112 323.425
R3379 gnd.n3438 gnd.n3412 289.615
R3380 gnd.n3406 gnd.n3380 289.615
R3381 gnd.n3374 gnd.n3348 289.615
R3382 gnd.n3343 gnd.n3317 289.615
R3383 gnd.n3311 gnd.n3285 289.615
R3384 gnd.n3279 gnd.n3253 289.615
R3385 gnd.n3247 gnd.n3221 289.615
R3386 gnd.n3216 gnd.n3190 289.615
R3387 gnd.n2663 gnd.t174 279.217
R3388 gnd.n2185 gnd.t108 279.217
R3389 gnd.n1191 gnd.t151 260.649
R3390 gnd.n1451 gnd.t157 260.649
R3391 gnd.n5404 gnd.n5403 256.663
R3392 gnd.n5404 gnd.n1150 256.663
R3393 gnd.n5404 gnd.n1151 256.663
R3394 gnd.n5404 gnd.n1152 256.663
R3395 gnd.n5404 gnd.n1153 256.663
R3396 gnd.n5404 gnd.n1154 256.663
R3397 gnd.n5404 gnd.n1155 256.663
R3398 gnd.n5404 gnd.n1156 256.663
R3399 gnd.n5404 gnd.n1157 256.663
R3400 gnd.n5404 gnd.n1158 256.663
R3401 gnd.n5404 gnd.n1159 256.663
R3402 gnd.n5404 gnd.n1160 256.663
R3403 gnd.n5404 gnd.n1161 256.663
R3404 gnd.n5404 gnd.n1162 256.663
R3405 gnd.n5404 gnd.n1163 256.663
R3406 gnd.n5404 gnd.n1164 256.663
R3407 gnd.n5407 gnd.n1147 256.663
R3408 gnd.n5405 gnd.n5404 256.663
R3409 gnd.n5404 gnd.n1165 256.663
R3410 gnd.n5404 gnd.n1166 256.663
R3411 gnd.n5404 gnd.n1167 256.663
R3412 gnd.n5404 gnd.n1168 256.663
R3413 gnd.n5404 gnd.n1169 256.663
R3414 gnd.n5404 gnd.n1170 256.663
R3415 gnd.n5404 gnd.n1171 256.663
R3416 gnd.n5404 gnd.n1172 256.663
R3417 gnd.n5404 gnd.n1173 256.663
R3418 gnd.n5404 gnd.n1174 256.663
R3419 gnd.n5404 gnd.n1175 256.663
R3420 gnd.n5404 gnd.n1176 256.663
R3421 gnd.n5404 gnd.n1177 256.663
R3422 gnd.n5404 gnd.n1178 256.663
R3423 gnd.n5404 gnd.n1179 256.663
R3424 gnd.n5404 gnd.n1180 256.663
R3425 gnd.n4941 gnd.n1461 256.663
R3426 gnd.n4947 gnd.n1461 256.663
R3427 gnd.n1508 gnd.n1461 256.663
R3428 gnd.n4954 gnd.n1461 256.663
R3429 gnd.n1505 gnd.n1461 256.663
R3430 gnd.n4961 gnd.n1461 256.663
R3431 gnd.n1502 gnd.n1461 256.663
R3432 gnd.n4968 gnd.n1461 256.663
R3433 gnd.n1499 gnd.n1461 256.663
R3434 gnd.n4975 gnd.n1461 256.663
R3435 gnd.n1496 gnd.n1461 256.663
R3436 gnd.n4982 gnd.n1461 256.663
R3437 gnd.n1493 gnd.n1461 256.663
R3438 gnd.n4989 gnd.n1461 256.663
R3439 gnd.n1490 gnd.n1461 256.663
R3440 gnd.n4997 gnd.n1461 256.663
R3441 gnd.n5000 gnd.n435 256.663
R3442 gnd.n5001 gnd.n1461 256.663
R3443 gnd.n5005 gnd.n1461 256.663
R3444 gnd.n1484 gnd.n1461 256.663
R3445 gnd.n5013 gnd.n1461 256.663
R3446 gnd.n1479 gnd.n1461 256.663
R3447 gnd.n5020 gnd.n1461 256.663
R3448 gnd.n1476 gnd.n1461 256.663
R3449 gnd.n5027 gnd.n1461 256.663
R3450 gnd.n1473 gnd.n1461 256.663
R3451 gnd.n5034 gnd.n1461 256.663
R3452 gnd.n1470 gnd.n1461 256.663
R3453 gnd.n5041 gnd.n1461 256.663
R3454 gnd.n1467 gnd.n1461 256.663
R3455 gnd.n5048 gnd.n1461 256.663
R3456 gnd.n1464 gnd.n1461 256.663
R3457 gnd.n5055 gnd.n1461 256.663
R3458 gnd.n1461 gnd.n1460 256.663
R3459 gnd.n3879 gnd.n3878 242.672
R3460 gnd.n3878 gnd.n3589 242.672
R3461 gnd.n3878 gnd.n3590 242.672
R3462 gnd.n3878 gnd.n3591 242.672
R3463 gnd.n3878 gnd.n3592 242.672
R3464 gnd.n3878 gnd.n3593 242.672
R3465 gnd.n3878 gnd.n3594 242.672
R3466 gnd.n3878 gnd.n3595 242.672
R3467 gnd.n3878 gnd.n3596 242.672
R3468 gnd.n5437 gnd.n1105 242.672
R3469 gnd.n5437 gnd.n1104 242.672
R3470 gnd.n5437 gnd.n1103 242.672
R3471 gnd.n5437 gnd.n1102 242.672
R3472 gnd.n5437 gnd.n1101 242.672
R3473 gnd.n5437 gnd.n1100 242.672
R3474 gnd.n5437 gnd.n1099 242.672
R3475 gnd.n5437 gnd.n1098 242.672
R3476 gnd.n5437 gnd.n1097 242.672
R3477 gnd.n6390 gnd.n403 242.672
R3478 gnd.n6390 gnd.n405 242.672
R3479 gnd.n6390 gnd.n407 242.672
R3480 gnd.n6390 gnd.n408 242.672
R3481 gnd.n6390 gnd.n410 242.672
R3482 gnd.n6390 gnd.n412 242.672
R3483 gnd.n6390 gnd.n413 242.672
R3484 gnd.n6390 gnd.n415 242.672
R3485 gnd.n6390 gnd.n416 242.672
R3486 gnd.n6637 gnd.n83 242.672
R3487 gnd.n6633 gnd.n83 242.672
R3488 gnd.n6628 gnd.n83 242.672
R3489 gnd.n6625 gnd.n83 242.672
R3490 gnd.n6620 gnd.n83 242.672
R3491 gnd.n6617 gnd.n83 242.672
R3492 gnd.n6612 gnd.n83 242.672
R3493 gnd.n6609 gnd.n83 242.672
R3494 gnd.n6604 gnd.n83 242.672
R3495 gnd.n2717 gnd.n2716 242.672
R3496 gnd.n2717 gnd.n2627 242.672
R3497 gnd.n2717 gnd.n2628 242.672
R3498 gnd.n2717 gnd.n2629 242.672
R3499 gnd.n2717 gnd.n2630 242.672
R3500 gnd.n2717 gnd.n2631 242.672
R3501 gnd.n2717 gnd.n2632 242.672
R3502 gnd.n2717 gnd.n2633 242.672
R3503 gnd.n2717 gnd.n2634 242.672
R3504 gnd.n2717 gnd.n2635 242.672
R3505 gnd.n2717 gnd.n2636 242.672
R3506 gnd.n2717 gnd.n2637 242.672
R3507 gnd.n2718 gnd.n2717 242.672
R3508 gnd.n3570 gnd.n2134 242.672
R3509 gnd.n3570 gnd.n2133 242.672
R3510 gnd.n3570 gnd.n2132 242.672
R3511 gnd.n3570 gnd.n2131 242.672
R3512 gnd.n3570 gnd.n2130 242.672
R3513 gnd.n3570 gnd.n2129 242.672
R3514 gnd.n3570 gnd.n2128 242.672
R3515 gnd.n3570 gnd.n2127 242.672
R3516 gnd.n3570 gnd.n2126 242.672
R3517 gnd.n3570 gnd.n2125 242.672
R3518 gnd.n3570 gnd.n2124 242.672
R3519 gnd.n3570 gnd.n2123 242.672
R3520 gnd.n3570 gnd.n2122 242.672
R3521 gnd.n2801 gnd.n2800 242.672
R3522 gnd.n2800 gnd.n2539 242.672
R3523 gnd.n2800 gnd.n2540 242.672
R3524 gnd.n2800 gnd.n2541 242.672
R3525 gnd.n2800 gnd.n2542 242.672
R3526 gnd.n2800 gnd.n2543 242.672
R3527 gnd.n2800 gnd.n2544 242.672
R3528 gnd.n2800 gnd.n2545 242.672
R3529 gnd.n3570 gnd.n2135 242.672
R3530 gnd.n3570 gnd.n2136 242.672
R3531 gnd.n3570 gnd.n2137 242.672
R3532 gnd.n3570 gnd.n2138 242.672
R3533 gnd.n3570 gnd.n2139 242.672
R3534 gnd.n3570 gnd.n2140 242.672
R3535 gnd.n3570 gnd.n2141 242.672
R3536 gnd.n3570 gnd.n2142 242.672
R3537 gnd.n3878 gnd.n3877 242.672
R3538 gnd.n3878 gnd.n3571 242.672
R3539 gnd.n3878 gnd.n3572 242.672
R3540 gnd.n3878 gnd.n3573 242.672
R3541 gnd.n3878 gnd.n3574 242.672
R3542 gnd.n3878 gnd.n3575 242.672
R3543 gnd.n3878 gnd.n3576 242.672
R3544 gnd.n3878 gnd.n3577 242.672
R3545 gnd.n3878 gnd.n3578 242.672
R3546 gnd.n3878 gnd.n3579 242.672
R3547 gnd.n3878 gnd.n3580 242.672
R3548 gnd.n3878 gnd.n3581 242.672
R3549 gnd.n3878 gnd.n3582 242.672
R3550 gnd.n3878 gnd.n3583 242.672
R3551 gnd.n3878 gnd.n3584 242.672
R3552 gnd.n3878 gnd.n3585 242.672
R3553 gnd.n3878 gnd.n3586 242.672
R3554 gnd.n3878 gnd.n3587 242.672
R3555 gnd.n3878 gnd.n3588 242.672
R3556 gnd.n5437 gnd.n1107 242.672
R3557 gnd.n5437 gnd.n1108 242.672
R3558 gnd.n5437 gnd.n1109 242.672
R3559 gnd.n5437 gnd.n1110 242.672
R3560 gnd.n5437 gnd.n1111 242.672
R3561 gnd.n5437 gnd.n1112 242.672
R3562 gnd.n5437 gnd.n1113 242.672
R3563 gnd.n5437 gnd.n1114 242.672
R3564 gnd.n5437 gnd.n1115 242.672
R3565 gnd.n5437 gnd.n1116 242.672
R3566 gnd.n5437 gnd.n1117 242.672
R3567 gnd.n5408 gnd.n1143 242.672
R3568 gnd.n5437 gnd.n1118 242.672
R3569 gnd.n5437 gnd.n1119 242.672
R3570 gnd.n5437 gnd.n1120 242.672
R3571 gnd.n5437 gnd.n1121 242.672
R3572 gnd.n5437 gnd.n1122 242.672
R3573 gnd.n5437 gnd.n1123 242.672
R3574 gnd.n5437 gnd.n1124 242.672
R3575 gnd.n5437 gnd.n5436 242.672
R3576 gnd.n6390 gnd.n6389 242.672
R3577 gnd.n6390 gnd.n385 242.672
R3578 gnd.n6390 gnd.n386 242.672
R3579 gnd.n6390 gnd.n387 242.672
R3580 gnd.n6390 gnd.n388 242.672
R3581 gnd.n6390 gnd.n389 242.672
R3582 gnd.n6390 gnd.n390 242.672
R3583 gnd.n6390 gnd.n391 242.672
R3584 gnd.n6359 gnd.n436 242.672
R3585 gnd.n6390 gnd.n392 242.672
R3586 gnd.n6390 gnd.n393 242.672
R3587 gnd.n6390 gnd.n394 242.672
R3588 gnd.n6390 gnd.n395 242.672
R3589 gnd.n6390 gnd.n396 242.672
R3590 gnd.n6390 gnd.n397 242.672
R3591 gnd.n6390 gnd.n398 242.672
R3592 gnd.n6390 gnd.n399 242.672
R3593 gnd.n6390 gnd.n400 242.672
R3594 gnd.n6390 gnd.n401 242.672
R3595 gnd.n6390 gnd.n402 242.672
R3596 gnd.n153 gnd.n83 242.672
R3597 gnd.n6695 gnd.n83 242.672
R3598 gnd.n149 gnd.n83 242.672
R3599 gnd.n6702 gnd.n83 242.672
R3600 gnd.n142 gnd.n83 242.672
R3601 gnd.n6709 gnd.n83 242.672
R3602 gnd.n135 gnd.n83 242.672
R3603 gnd.n6716 gnd.n83 242.672
R3604 gnd.n128 gnd.n83 242.672
R3605 gnd.n6723 gnd.n83 242.672
R3606 gnd.n121 gnd.n83 242.672
R3607 gnd.n6733 gnd.n83 242.672
R3608 gnd.n114 gnd.n83 242.672
R3609 gnd.n6740 gnd.n83 242.672
R3610 gnd.n107 gnd.n83 242.672
R3611 gnd.n6747 gnd.n83 242.672
R3612 gnd.n100 gnd.n83 242.672
R3613 gnd.n6754 gnd.n83 242.672
R3614 gnd.n93 gnd.n83 242.672
R3615 gnd.n4234 gnd.n1848 242.672
R3616 gnd.n4234 gnd.n1849 242.672
R3617 gnd.n4234 gnd.n1850 242.672
R3618 gnd.n4234 gnd.n1851 242.672
R3619 gnd.n4234 gnd.n1852 242.672
R3620 gnd.n4234 gnd.n1853 242.672
R3621 gnd.n4234 gnd.n1854 242.672
R3622 gnd.n4234 gnd.n1855 242.672
R3623 gnd.n4234 gnd.n1856 242.672
R3624 gnd.n4234 gnd.n1857 242.672
R3625 gnd.n4234 gnd.n1858 242.672
R3626 gnd.n4234 gnd.n1859 242.672
R3627 gnd.n4234 gnd.n1860 242.672
R3628 gnd.n4234 gnd.n1861 242.672
R3629 gnd.n5181 gnd.n5179 242.672
R3630 gnd.n5181 gnd.n5092 242.672
R3631 gnd.n5181 gnd.n5091 242.672
R3632 gnd.n5181 gnd.n5090 242.672
R3633 gnd.n5181 gnd.n5089 242.672
R3634 gnd.n5181 gnd.n5088 242.672
R3635 gnd.n5181 gnd.n5087 242.672
R3636 gnd.n5181 gnd.n5085 242.672
R3637 gnd.n5181 gnd.n5084 242.672
R3638 gnd.n5181 gnd.n5082 242.672
R3639 gnd.n5181 gnd.n5080 242.672
R3640 gnd.n5181 gnd.n5079 242.672
R3641 gnd.n5181 gnd.n5077 242.672
R3642 gnd.n5181 gnd.n5075 242.672
R3643 gnd.n90 gnd.n86 240.244
R3644 gnd.n6756 gnd.n6755 240.244
R3645 gnd.n6753 gnd.n94 240.244
R3646 gnd.n6749 gnd.n6748 240.244
R3647 gnd.n6746 gnd.n101 240.244
R3648 gnd.n6742 gnd.n6741 240.244
R3649 gnd.n6739 gnd.n108 240.244
R3650 gnd.n6735 gnd.n6734 240.244
R3651 gnd.n6732 gnd.n115 240.244
R3652 gnd.n6725 gnd.n6724 240.244
R3653 gnd.n6722 gnd.n122 240.244
R3654 gnd.n6718 gnd.n6717 240.244
R3655 gnd.n6715 gnd.n129 240.244
R3656 gnd.n6711 gnd.n6710 240.244
R3657 gnd.n6708 gnd.n136 240.244
R3658 gnd.n6704 gnd.n6703 240.244
R3659 gnd.n6701 gnd.n143 240.244
R3660 gnd.n6697 gnd.n6696 240.244
R3661 gnd.n6694 gnd.n150 240.244
R3662 gnd.n464 gnd.n329 240.244
R3663 gnd.n464 gnd.n321 240.244
R3664 gnd.n6311 gnd.n321 240.244
R3665 gnd.n6311 gnd.n313 240.244
R3666 gnd.n488 gnd.n313 240.244
R3667 gnd.n488 gnd.n304 240.244
R3668 gnd.n494 gnd.n304 240.244
R3669 gnd.n494 gnd.n295 240.244
R3670 gnd.n498 gnd.n295 240.244
R3671 gnd.n498 gnd.n286 240.244
R3672 gnd.n6218 gnd.n286 240.244
R3673 gnd.n6218 gnd.n277 240.244
R3674 gnd.n6222 gnd.n277 240.244
R3675 gnd.n6222 gnd.n269 240.244
R3676 gnd.n6286 gnd.n269 240.244
R3677 gnd.n6286 gnd.n261 240.244
R3678 gnd.n261 gnd.n256 240.244
R3679 gnd.n6281 gnd.n256 240.244
R3680 gnd.n6281 gnd.n248 240.244
R3681 gnd.n248 gnd.n243 240.244
R3682 gnd.n6277 gnd.n243 240.244
R3683 gnd.n6277 gnd.n236 240.244
R3684 gnd.n6274 gnd.n236 240.244
R3685 gnd.n6274 gnd.n231 240.244
R3686 gnd.n6271 gnd.n231 240.244
R3687 gnd.n6271 gnd.n223 240.244
R3688 gnd.n6268 gnd.n223 240.244
R3689 gnd.n6268 gnd.n209 240.244
R3690 gnd.n6265 gnd.n209 240.244
R3691 gnd.n6265 gnd.n203 240.244
R3692 gnd.n6262 gnd.n203 240.244
R3693 gnd.n6262 gnd.n195 240.244
R3694 gnd.n6259 gnd.n195 240.244
R3695 gnd.n6259 gnd.n187 240.244
R3696 gnd.n6256 gnd.n187 240.244
R3697 gnd.n6256 gnd.n178 240.244
R3698 gnd.n6253 gnd.n178 240.244
R3699 gnd.n6253 gnd.n170 240.244
R3700 gnd.n170 gnd.n160 240.244
R3701 gnd.n6685 gnd.n160 240.244
R3702 gnd.n6686 gnd.n6685 240.244
R3703 gnd.n6686 gnd.n82 240.244
R3704 gnd.n6388 gnd.n418 240.244
R3705 gnd.n6384 gnd.n418 240.244
R3706 gnd.n6382 gnd.n6381 240.244
R3707 gnd.n6378 gnd.n6377 240.244
R3708 gnd.n6374 gnd.n6373 240.244
R3709 gnd.n6370 gnd.n6369 240.244
R3710 gnd.n6366 gnd.n6365 240.244
R3711 gnd.n6362 gnd.n6361 240.244
R3712 gnd.n6357 gnd.n6356 240.244
R3713 gnd.n6353 gnd.n6352 240.244
R3714 gnd.n6349 gnd.n6348 240.244
R3715 gnd.n6345 gnd.n6344 240.244
R3716 gnd.n6341 gnd.n6340 240.244
R3717 gnd.n6337 gnd.n6336 240.244
R3718 gnd.n6333 gnd.n6332 240.244
R3719 gnd.n6329 gnd.n6328 240.244
R3720 gnd.n6325 gnd.n6324 240.244
R3721 gnd.n459 gnd.n458 240.244
R3722 gnd.n6446 gnd.n324 240.244
R3723 gnd.n6452 gnd.n324 240.244
R3724 gnd.n6452 gnd.n311 240.244
R3725 gnd.n6462 gnd.n311 240.244
R3726 gnd.n6462 gnd.n307 240.244
R3727 gnd.n6468 gnd.n307 240.244
R3728 gnd.n6468 gnd.n293 240.244
R3729 gnd.n6478 gnd.n293 240.244
R3730 gnd.n6478 gnd.n289 240.244
R3731 gnd.n6484 gnd.n289 240.244
R3732 gnd.n6484 gnd.n276 240.244
R3733 gnd.n6494 gnd.n276 240.244
R3734 gnd.n6494 gnd.n272 240.244
R3735 gnd.n6501 gnd.n272 240.244
R3736 gnd.n6501 gnd.n258 240.244
R3737 gnd.n6515 gnd.n258 240.244
R3738 gnd.n6518 gnd.n6515 240.244
R3739 gnd.n6518 gnd.n246 240.244
R3740 gnd.n6528 gnd.n246 240.244
R3741 gnd.n6531 gnd.n6528 240.244
R3742 gnd.n6531 gnd.n232 240.244
R3743 gnd.n6541 gnd.n232 240.244
R3744 gnd.n6542 gnd.n6541 240.244
R3745 gnd.n6545 gnd.n6542 240.244
R3746 gnd.n6545 gnd.n220 240.244
R3747 gnd.n6555 gnd.n220 240.244
R3748 gnd.n6555 gnd.n210 240.244
R3749 gnd.n6561 gnd.n210 240.244
R3750 gnd.n6561 gnd.n200 240.244
R3751 gnd.n6571 gnd.n200 240.244
R3752 gnd.n6571 gnd.n196 240.244
R3753 gnd.n6577 gnd.n196 240.244
R3754 gnd.n6577 gnd.n184 240.244
R3755 gnd.n6587 gnd.n184 240.244
R3756 gnd.n6587 gnd.n180 240.244
R3757 gnd.n6593 gnd.n180 240.244
R3758 gnd.n6593 gnd.n167 240.244
R3759 gnd.n6677 gnd.n167 240.244
R3760 gnd.n6677 gnd.n163 240.244
R3761 gnd.n6683 gnd.n163 240.244
R3762 gnd.n6683 gnd.n85 240.244
R3763 gnd.n6763 gnd.n85 240.244
R3764 gnd.n5438 gnd.n1094 240.244
R3765 gnd.n5435 gnd.n1125 240.244
R3766 gnd.n5431 gnd.n5430 240.244
R3767 gnd.n5427 gnd.n5426 240.244
R3768 gnd.n5423 gnd.n5422 240.244
R3769 gnd.n5419 gnd.n5418 240.244
R3770 gnd.n5415 gnd.n5414 240.244
R3771 gnd.n5411 gnd.n5410 240.244
R3772 gnd.n4093 gnd.n4092 240.244
R3773 gnd.n4100 gnd.n4099 240.244
R3774 gnd.n4103 gnd.n4102 240.244
R3775 gnd.n4110 gnd.n4109 240.244
R3776 gnd.n4113 gnd.n4112 240.244
R3777 gnd.n4120 gnd.n4119 240.244
R3778 gnd.n4123 gnd.n4122 240.244
R3779 gnd.n4130 gnd.n4129 240.244
R3780 gnd.n4133 gnd.n4132 240.244
R3781 gnd.n4138 gnd.n4083 240.244
R3782 gnd.n3799 gnd.n2113 240.244
R3783 gnd.n3753 gnd.n2113 240.244
R3784 gnd.n3753 gnd.n2105 240.244
R3785 gnd.n3791 gnd.n2105 240.244
R3786 gnd.n3791 gnd.n2096 240.244
R3787 gnd.n3788 gnd.n2096 240.244
R3788 gnd.n3788 gnd.n2088 240.244
R3789 gnd.n3785 gnd.n2088 240.244
R3790 gnd.n3785 gnd.n2081 240.244
R3791 gnd.n3782 gnd.n2081 240.244
R3792 gnd.n3782 gnd.n2073 240.244
R3793 gnd.n3779 gnd.n2073 240.244
R3794 gnd.n3779 gnd.n2064 240.244
R3795 gnd.n3776 gnd.n2064 240.244
R3796 gnd.n3776 gnd.n2056 240.244
R3797 gnd.n3773 gnd.n2056 240.244
R3798 gnd.n3773 gnd.n2048 240.244
R3799 gnd.n2048 gnd.n2040 240.244
R3800 gnd.n3965 gnd.n2040 240.244
R3801 gnd.n3966 gnd.n3965 240.244
R3802 gnd.n3966 gnd.n2030 240.244
R3803 gnd.n3974 gnd.n2030 240.244
R3804 gnd.n3974 gnd.n2024 240.244
R3805 gnd.n3971 gnd.n2024 240.244
R3806 gnd.n3971 gnd.n999 240.244
R3807 gnd.n4009 gnd.n999 240.244
R3808 gnd.n4009 gnd.n1011 240.244
R3809 gnd.n2012 gnd.n1011 240.244
R3810 gnd.n2012 gnd.n1022 240.244
R3811 gnd.n4021 gnd.n1022 240.244
R3812 gnd.n4021 gnd.n1033 240.244
R3813 gnd.n2006 gnd.n1033 240.244
R3814 gnd.n2006 gnd.n1043 240.244
R3815 gnd.n4066 gnd.n1043 240.244
R3816 gnd.n4066 gnd.n1054 240.244
R3817 gnd.n1992 gnd.n1054 240.244
R3818 gnd.n1992 gnd.n1064 240.244
R3819 gnd.n4074 gnd.n1064 240.244
R3820 gnd.n4074 gnd.n1075 240.244
R3821 gnd.n4148 gnd.n1075 240.244
R3822 gnd.n4148 gnd.n1086 240.244
R3823 gnd.n1981 gnd.n1086 240.244
R3824 gnd.n3708 gnd.n3707 240.244
R3825 gnd.n3871 gnd.n3707 240.244
R3826 gnd.n3869 gnd.n3868 240.244
R3827 gnd.n3865 gnd.n3864 240.244
R3828 gnd.n3861 gnd.n3860 240.244
R3829 gnd.n3857 gnd.n3856 240.244
R3830 gnd.n3853 gnd.n3852 240.244
R3831 gnd.n3849 gnd.n3848 240.244
R3832 gnd.n3845 gnd.n3844 240.244
R3833 gnd.n3840 gnd.n3839 240.244
R3834 gnd.n3836 gnd.n3835 240.244
R3835 gnd.n3832 gnd.n3831 240.244
R3836 gnd.n3828 gnd.n3827 240.244
R3837 gnd.n3824 gnd.n3823 240.244
R3838 gnd.n3820 gnd.n3819 240.244
R3839 gnd.n3816 gnd.n3815 240.244
R3840 gnd.n3812 gnd.n3811 240.244
R3841 gnd.n3808 gnd.n3807 240.244
R3842 gnd.n3748 gnd.n3747 240.244
R3843 gnd.n3888 gnd.n2111 240.244
R3844 gnd.n3888 gnd.n2107 240.244
R3845 gnd.n3894 gnd.n2107 240.244
R3846 gnd.n3894 gnd.n2094 240.244
R3847 gnd.n3904 gnd.n2094 240.244
R3848 gnd.n3904 gnd.n2090 240.244
R3849 gnd.n3910 gnd.n2090 240.244
R3850 gnd.n3910 gnd.n2079 240.244
R3851 gnd.n3920 gnd.n2079 240.244
R3852 gnd.n3920 gnd.n2075 240.244
R3853 gnd.n3926 gnd.n2075 240.244
R3854 gnd.n3926 gnd.n2062 240.244
R3855 gnd.n3936 gnd.n2062 240.244
R3856 gnd.n3936 gnd.n2058 240.244
R3857 gnd.n3943 gnd.n2058 240.244
R3858 gnd.n3943 gnd.n2046 240.244
R3859 gnd.n3957 gnd.n2046 240.244
R3860 gnd.n3957 gnd.n2044 240.244
R3861 gnd.n3963 gnd.n2044 240.244
R3862 gnd.n3963 gnd.n2028 240.244
R3863 gnd.n3992 gnd.n2028 240.244
R3864 gnd.n3992 gnd.n2026 240.244
R3865 gnd.n3998 gnd.n2026 240.244
R3866 gnd.n3998 gnd.n1003 240.244
R3867 gnd.n5492 gnd.n1003 240.244
R3868 gnd.n5492 gnd.n1004 240.244
R3869 gnd.n5488 gnd.n1004 240.244
R3870 gnd.n5488 gnd.n1009 240.244
R3871 gnd.n5480 gnd.n1009 240.244
R3872 gnd.n5480 gnd.n1025 240.244
R3873 gnd.n5476 gnd.n1025 240.244
R3874 gnd.n5476 gnd.n1031 240.244
R3875 gnd.n5468 gnd.n1031 240.244
R3876 gnd.n5468 gnd.n1046 240.244
R3877 gnd.n5464 gnd.n1046 240.244
R3878 gnd.n5464 gnd.n1052 240.244
R3879 gnd.n5456 gnd.n1052 240.244
R3880 gnd.n5456 gnd.n1067 240.244
R3881 gnd.n5452 gnd.n1067 240.244
R3882 gnd.n5452 gnd.n1073 240.244
R3883 gnd.n5444 gnd.n1073 240.244
R3884 gnd.n5444 gnd.n1089 240.244
R3885 gnd.n3569 gnd.n2144 240.244
R3886 gnd.n3562 gnd.n3561 240.244
R3887 gnd.n3559 gnd.n3558 240.244
R3888 gnd.n3555 gnd.n3554 240.244
R3889 gnd.n3551 gnd.n3550 240.244
R3890 gnd.n3547 gnd.n3546 240.244
R3891 gnd.n3543 gnd.n3542 240.244
R3892 gnd.n3539 gnd.n3538 240.244
R3893 gnd.n2812 gnd.n2524 240.244
R3894 gnd.n2822 gnd.n2524 240.244
R3895 gnd.n2822 gnd.n2515 240.244
R3896 gnd.n2515 gnd.n2504 240.244
R3897 gnd.n2843 gnd.n2504 240.244
R3898 gnd.n2843 gnd.n2498 240.244
R3899 gnd.n2853 gnd.n2498 240.244
R3900 gnd.n2853 gnd.n2487 240.244
R3901 gnd.n2487 gnd.n2479 240.244
R3902 gnd.n2871 gnd.n2479 240.244
R3903 gnd.n2872 gnd.n2871 240.244
R3904 gnd.n2872 gnd.n2464 240.244
R3905 gnd.n2874 gnd.n2464 240.244
R3906 gnd.n2874 gnd.n2450 240.244
R3907 gnd.n2916 gnd.n2450 240.244
R3908 gnd.n2917 gnd.n2916 240.244
R3909 gnd.n2920 gnd.n2917 240.244
R3910 gnd.n2920 gnd.n2405 240.244
R3911 gnd.n2445 gnd.n2405 240.244
R3912 gnd.n2445 gnd.n2415 240.244
R3913 gnd.n2930 gnd.n2415 240.244
R3914 gnd.n2930 gnd.n2436 240.244
R3915 gnd.n2940 gnd.n2436 240.244
R3916 gnd.n2940 gnd.n2346 240.244
R3917 gnd.n2985 gnd.n2346 240.244
R3918 gnd.n2985 gnd.n2332 240.244
R3919 gnd.n3007 gnd.n2332 240.244
R3920 gnd.n3008 gnd.n3007 240.244
R3921 gnd.n3008 gnd.n2319 240.244
R3922 gnd.n2319 gnd.n2308 240.244
R3923 gnd.n3039 gnd.n2308 240.244
R3924 gnd.n3040 gnd.n3039 240.244
R3925 gnd.n3041 gnd.n3040 240.244
R3926 gnd.n3041 gnd.n2293 240.244
R3927 gnd.n2293 gnd.n2292 240.244
R3928 gnd.n2292 gnd.n2277 240.244
R3929 gnd.n3092 gnd.n2277 240.244
R3930 gnd.n3093 gnd.n3092 240.244
R3931 gnd.n3093 gnd.n2264 240.244
R3932 gnd.n2264 gnd.n2253 240.244
R3933 gnd.n3124 gnd.n2253 240.244
R3934 gnd.n3125 gnd.n3124 240.244
R3935 gnd.n3126 gnd.n3125 240.244
R3936 gnd.n3126 gnd.n2237 240.244
R3937 gnd.n2237 gnd.n2236 240.244
R3938 gnd.n2236 gnd.n2223 240.244
R3939 gnd.n3181 gnd.n2223 240.244
R3940 gnd.n3182 gnd.n3181 240.244
R3941 gnd.n3182 gnd.n2210 240.244
R3942 gnd.n2210 gnd.n2200 240.244
R3943 gnd.n3470 gnd.n2200 240.244
R3944 gnd.n3473 gnd.n3470 240.244
R3945 gnd.n3473 gnd.n3472 240.244
R3946 gnd.n2802 gnd.n2537 240.244
R3947 gnd.n2558 gnd.n2537 240.244
R3948 gnd.n2561 gnd.n2560 240.244
R3949 gnd.n2568 gnd.n2567 240.244
R3950 gnd.n2571 gnd.n2570 240.244
R3951 gnd.n2578 gnd.n2577 240.244
R3952 gnd.n2581 gnd.n2580 240.244
R3953 gnd.n2588 gnd.n2587 240.244
R3954 gnd.n2810 gnd.n2534 240.244
R3955 gnd.n2534 gnd.n2513 240.244
R3956 gnd.n2833 gnd.n2513 240.244
R3957 gnd.n2833 gnd.n2507 240.244
R3958 gnd.n2841 gnd.n2507 240.244
R3959 gnd.n2841 gnd.n2509 240.244
R3960 gnd.n2509 gnd.n2485 240.244
R3961 gnd.n2863 gnd.n2485 240.244
R3962 gnd.n2863 gnd.n2481 240.244
R3963 gnd.n2869 gnd.n2481 240.244
R3964 gnd.n2869 gnd.n2463 240.244
R3965 gnd.n2894 gnd.n2463 240.244
R3966 gnd.n2894 gnd.n2458 240.244
R3967 gnd.n2906 gnd.n2458 240.244
R3968 gnd.n2906 gnd.n2459 240.244
R3969 gnd.n2902 gnd.n2459 240.244
R3970 gnd.n2902 gnd.n2407 240.244
R3971 gnd.n2954 gnd.n2407 240.244
R3972 gnd.n2954 gnd.n2408 240.244
R3973 gnd.n2950 gnd.n2408 240.244
R3974 gnd.n2950 gnd.n2414 240.244
R3975 gnd.n2434 gnd.n2414 240.244
R3976 gnd.n2434 gnd.n2344 240.244
R3977 gnd.n2989 gnd.n2344 240.244
R3978 gnd.n2989 gnd.n2339 240.244
R3979 gnd.n2997 gnd.n2339 240.244
R3980 gnd.n2997 gnd.n2340 240.244
R3981 gnd.n2340 gnd.n2317 240.244
R3982 gnd.n3029 gnd.n2317 240.244
R3983 gnd.n3029 gnd.n2312 240.244
R3984 gnd.n3037 gnd.n2312 240.244
R3985 gnd.n3037 gnd.n2313 240.244
R3986 gnd.n2313 gnd.n2290 240.244
R3987 gnd.n3074 gnd.n2290 240.244
R3988 gnd.n3074 gnd.n2285 240.244
R3989 gnd.n3082 gnd.n2285 240.244
R3990 gnd.n3082 gnd.n2286 240.244
R3991 gnd.n2286 gnd.n2262 240.244
R3992 gnd.n3114 gnd.n2262 240.244
R3993 gnd.n3114 gnd.n2257 240.244
R3994 gnd.n3122 gnd.n2257 240.244
R3995 gnd.n3122 gnd.n2258 240.244
R3996 gnd.n2258 gnd.n2235 240.244
R3997 gnd.n3163 gnd.n2235 240.244
R3998 gnd.n3163 gnd.n2230 240.244
R3999 gnd.n3171 gnd.n2230 240.244
R4000 gnd.n3171 gnd.n2231 240.244
R4001 gnd.n2231 gnd.n2208 240.244
R4002 gnd.n3458 gnd.n2208 240.244
R4003 gnd.n3458 gnd.n2203 240.244
R4004 gnd.n3468 gnd.n2203 240.244
R4005 gnd.n3468 gnd.n2204 240.244
R4006 gnd.n2204 gnd.n2143 240.244
R4007 gnd.n2163 gnd.n2121 240.244
R4008 gnd.n3529 gnd.n3528 240.244
R4009 gnd.n3525 gnd.n3524 240.244
R4010 gnd.n3521 gnd.n3520 240.244
R4011 gnd.n3517 gnd.n3516 240.244
R4012 gnd.n3513 gnd.n3512 240.244
R4013 gnd.n3509 gnd.n3508 240.244
R4014 gnd.n3505 gnd.n3504 240.244
R4015 gnd.n3501 gnd.n3500 240.244
R4016 gnd.n3497 gnd.n3496 240.244
R4017 gnd.n3493 gnd.n3492 240.244
R4018 gnd.n3489 gnd.n3488 240.244
R4019 gnd.n3485 gnd.n3484 240.244
R4020 gnd.n2725 gnd.n2622 240.244
R4021 gnd.n2725 gnd.n2615 240.244
R4022 gnd.n2736 gnd.n2615 240.244
R4023 gnd.n2736 gnd.n2611 240.244
R4024 gnd.n2742 gnd.n2611 240.244
R4025 gnd.n2742 gnd.n2603 240.244
R4026 gnd.n2752 gnd.n2603 240.244
R4027 gnd.n2752 gnd.n2598 240.244
R4028 gnd.n2788 gnd.n2598 240.244
R4029 gnd.n2788 gnd.n2599 240.244
R4030 gnd.n2599 gnd.n2546 240.244
R4031 gnd.n2783 gnd.n2546 240.244
R4032 gnd.n2783 gnd.n2782 240.244
R4033 gnd.n2782 gnd.n2525 240.244
R4034 gnd.n2778 gnd.n2525 240.244
R4035 gnd.n2778 gnd.n2516 240.244
R4036 gnd.n2775 gnd.n2516 240.244
R4037 gnd.n2775 gnd.n2774 240.244
R4038 gnd.n2774 gnd.n2499 240.244
R4039 gnd.n2770 gnd.n2499 240.244
R4040 gnd.n2770 gnd.n2488 240.244
R4041 gnd.n2488 gnd.n2469 240.244
R4042 gnd.n2883 gnd.n2469 240.244
R4043 gnd.n2883 gnd.n2465 240.244
R4044 gnd.n2891 gnd.n2465 240.244
R4045 gnd.n2891 gnd.n2456 240.244
R4046 gnd.n2456 gnd.n2392 240.244
R4047 gnd.n2963 gnd.n2392 240.244
R4048 gnd.n2963 gnd.n2393 240.244
R4049 gnd.n2404 gnd.n2393 240.244
R4050 gnd.n2439 gnd.n2404 240.244
R4051 gnd.n2442 gnd.n2439 240.244
R4052 gnd.n2442 gnd.n2416 240.244
R4053 gnd.n2429 gnd.n2416 240.244
R4054 gnd.n2429 gnd.n2426 240.244
R4055 gnd.n2426 gnd.n2347 240.244
R4056 gnd.n2984 gnd.n2347 240.244
R4057 gnd.n2984 gnd.n2337 240.244
R4058 gnd.n2980 gnd.n2337 240.244
R4059 gnd.n2980 gnd.n2331 240.244
R4060 gnd.n2977 gnd.n2331 240.244
R4061 gnd.n2977 gnd.n2320 240.244
R4062 gnd.n2974 gnd.n2320 240.244
R4063 gnd.n2974 gnd.n2298 240.244
R4064 gnd.n3050 gnd.n2298 240.244
R4065 gnd.n3050 gnd.n2294 240.244
R4066 gnd.n3071 gnd.n2294 240.244
R4067 gnd.n3071 gnd.n2283 240.244
R4068 gnd.n3067 gnd.n2283 240.244
R4069 gnd.n3067 gnd.n2276 240.244
R4070 gnd.n3064 gnd.n2276 240.244
R4071 gnd.n3064 gnd.n2265 240.244
R4072 gnd.n3061 gnd.n2265 240.244
R4073 gnd.n3061 gnd.n2242 240.244
R4074 gnd.n3135 gnd.n2242 240.244
R4075 gnd.n3135 gnd.n2238 240.244
R4076 gnd.n3160 gnd.n2238 240.244
R4077 gnd.n3160 gnd.n2229 240.244
R4078 gnd.n3156 gnd.n2229 240.244
R4079 gnd.n3156 gnd.n2222 240.244
R4080 gnd.n3152 gnd.n2222 240.244
R4081 gnd.n3152 gnd.n2211 240.244
R4082 gnd.n3149 gnd.n2211 240.244
R4083 gnd.n3149 gnd.n2192 240.244
R4084 gnd.n3480 gnd.n2192 240.244
R4085 gnd.n2639 gnd.n2638 240.244
R4086 gnd.n2710 gnd.n2638 240.244
R4087 gnd.n2708 gnd.n2707 240.244
R4088 gnd.n2704 gnd.n2703 240.244
R4089 gnd.n2700 gnd.n2699 240.244
R4090 gnd.n2696 gnd.n2695 240.244
R4091 gnd.n2692 gnd.n2691 240.244
R4092 gnd.n2688 gnd.n2687 240.244
R4093 gnd.n2684 gnd.n2683 240.244
R4094 gnd.n2680 gnd.n2679 240.244
R4095 gnd.n2676 gnd.n2675 240.244
R4096 gnd.n2672 gnd.n2671 240.244
R4097 gnd.n2668 gnd.n2626 240.244
R4098 gnd.n2728 gnd.n2620 240.244
R4099 gnd.n2728 gnd.n2616 240.244
R4100 gnd.n2734 gnd.n2616 240.244
R4101 gnd.n2734 gnd.n2609 240.244
R4102 gnd.n2744 gnd.n2609 240.244
R4103 gnd.n2744 gnd.n2605 240.244
R4104 gnd.n2750 gnd.n2605 240.244
R4105 gnd.n2750 gnd.n2596 240.244
R4106 gnd.n2790 gnd.n2596 240.244
R4107 gnd.n2790 gnd.n2547 240.244
R4108 gnd.n2798 gnd.n2547 240.244
R4109 gnd.n2798 gnd.n2548 240.244
R4110 gnd.n2548 gnd.n2526 240.244
R4111 gnd.n2819 gnd.n2526 240.244
R4112 gnd.n2819 gnd.n2518 240.244
R4113 gnd.n2830 gnd.n2518 240.244
R4114 gnd.n2830 gnd.n2519 240.244
R4115 gnd.n2519 gnd.n2500 240.244
R4116 gnd.n2850 gnd.n2500 240.244
R4117 gnd.n2850 gnd.n2490 240.244
R4118 gnd.n2860 gnd.n2490 240.244
R4119 gnd.n2860 gnd.n2471 240.244
R4120 gnd.n2881 gnd.n2471 240.244
R4121 gnd.n2881 gnd.n2473 240.244
R4122 gnd.n2473 gnd.n2454 240.244
R4123 gnd.n2909 gnd.n2454 240.244
R4124 gnd.n2909 gnd.n2396 240.244
R4125 gnd.n2961 gnd.n2396 240.244
R4126 gnd.n2961 gnd.n2397 240.244
R4127 gnd.n2957 gnd.n2397 240.244
R4128 gnd.n2957 gnd.n2403 240.244
R4129 gnd.n2418 gnd.n2403 240.244
R4130 gnd.n2947 gnd.n2418 240.244
R4131 gnd.n2947 gnd.n2419 240.244
R4132 gnd.n2943 gnd.n2419 240.244
R4133 gnd.n2943 gnd.n2425 240.244
R4134 gnd.n2425 gnd.n2336 240.244
R4135 gnd.n3000 gnd.n2336 240.244
R4136 gnd.n3000 gnd.n2329 240.244
R4137 gnd.n3011 gnd.n2329 240.244
R4138 gnd.n3011 gnd.n2322 240.244
R4139 gnd.n3026 gnd.n2322 240.244
R4140 gnd.n3026 gnd.n2323 240.244
R4141 gnd.n2323 gnd.n2301 240.244
R4142 gnd.n3048 gnd.n2301 240.244
R4143 gnd.n3048 gnd.n2302 240.244
R4144 gnd.n2302 gnd.n2281 240.244
R4145 gnd.n3085 gnd.n2281 240.244
R4146 gnd.n3085 gnd.n2274 240.244
R4147 gnd.n3096 gnd.n2274 240.244
R4148 gnd.n3096 gnd.n2267 240.244
R4149 gnd.n3111 gnd.n2267 240.244
R4150 gnd.n3111 gnd.n2268 240.244
R4151 gnd.n2268 gnd.n2245 240.244
R4152 gnd.n3133 gnd.n2245 240.244
R4153 gnd.n3133 gnd.n2247 240.244
R4154 gnd.n2247 gnd.n2227 240.244
R4155 gnd.n3174 gnd.n2227 240.244
R4156 gnd.n3174 gnd.n2220 240.244
R4157 gnd.n3186 gnd.n2220 240.244
R4158 gnd.n3186 gnd.n2213 240.244
R4159 gnd.n3455 gnd.n2213 240.244
R4160 gnd.n3455 gnd.n2214 240.244
R4161 gnd.n2214 gnd.n2195 240.244
R4162 gnd.n3478 gnd.n2195 240.244
R4163 gnd.n6603 gnd.n6602 240.244
R4164 gnd.n6608 gnd.n6605 240.244
R4165 gnd.n6611 gnd.n6610 240.244
R4166 gnd.n6616 gnd.n6613 240.244
R4167 gnd.n6619 gnd.n6618 240.244
R4168 gnd.n6624 gnd.n6621 240.244
R4169 gnd.n6627 gnd.n6626 240.244
R4170 gnd.n6632 gnd.n6629 240.244
R4171 gnd.n6638 gnd.n6634 240.244
R4172 gnd.n5151 gnd.n330 240.244
R4173 gnd.n5151 gnd.n322 240.244
R4174 gnd.n6309 gnd.n322 240.244
R4175 gnd.n6309 gnd.n314 240.244
R4176 gnd.n472 gnd.n314 240.244
R4177 gnd.n472 gnd.n305 240.244
R4178 gnd.n473 gnd.n305 240.244
R4179 gnd.n473 gnd.n296 240.244
R4180 gnd.n476 gnd.n296 240.244
R4181 gnd.n476 gnd.n287 240.244
R4182 gnd.n477 gnd.n287 240.244
R4183 gnd.n477 gnd.n278 240.244
R4184 gnd.n480 gnd.n278 240.244
R4185 gnd.n480 gnd.n270 240.244
R4186 gnd.n6288 gnd.n270 240.244
R4187 gnd.n6288 gnd.n254 240.244
R4188 gnd.n6520 gnd.n254 240.244
R4189 gnd.n6520 gnd.n249 240.244
R4190 gnd.n6526 gnd.n249 240.244
R4191 gnd.n6526 gnd.n245 240.244
R4192 gnd.n245 gnd.n244 240.244
R4193 gnd.n244 gnd.n54 240.244
R4194 gnd.n55 gnd.n54 240.244
R4195 gnd.n56 gnd.n55 240.244
R4196 gnd.n221 gnd.n56 240.244
R4197 gnd.n221 gnd.n59 240.244
R4198 gnd.n60 gnd.n59 240.244
R4199 gnd.n61 gnd.n60 240.244
R4200 gnd.n201 gnd.n61 240.244
R4201 gnd.n201 gnd.n64 240.244
R4202 gnd.n65 gnd.n64 240.244
R4203 gnd.n66 gnd.n65 240.244
R4204 gnd.n185 gnd.n66 240.244
R4205 gnd.n185 gnd.n69 240.244
R4206 gnd.n70 gnd.n69 240.244
R4207 gnd.n71 gnd.n70 240.244
R4208 gnd.n168 gnd.n71 240.244
R4209 gnd.n168 gnd.n74 240.244
R4210 gnd.n75 gnd.n74 240.244
R4211 gnd.n76 gnd.n75 240.244
R4212 gnd.n79 gnd.n76 240.244
R4213 gnd.n6765 gnd.n79 240.244
R4214 gnd.n404 gnd.n334 240.244
R4215 gnd.n342 gnd.n341 240.244
R4216 gnd.n406 gnd.n349 240.244
R4217 gnd.n409 gnd.n350 240.244
R4218 gnd.n358 gnd.n357 240.244
R4219 gnd.n411 gnd.n365 240.244
R4220 gnd.n414 gnd.n366 240.244
R4221 gnd.n374 gnd.n373 240.244
R4222 gnd.n6391 gnd.n383 240.244
R4223 gnd.n6444 gnd.n320 240.244
R4224 gnd.n6454 gnd.n320 240.244
R4225 gnd.n6454 gnd.n316 240.244
R4226 gnd.n6460 gnd.n316 240.244
R4227 gnd.n6460 gnd.n302 240.244
R4228 gnd.n6470 gnd.n302 240.244
R4229 gnd.n6470 gnd.n298 240.244
R4230 gnd.n6476 gnd.n298 240.244
R4231 gnd.n6476 gnd.n284 240.244
R4232 gnd.n6486 gnd.n284 240.244
R4233 gnd.n6486 gnd.n280 240.244
R4234 gnd.n6492 gnd.n280 240.244
R4235 gnd.n6492 gnd.n267 240.244
R4236 gnd.n6503 gnd.n267 240.244
R4237 gnd.n6503 gnd.n262 240.244
R4238 gnd.n6513 gnd.n262 240.244
R4239 gnd.n6513 gnd.n257 240.244
R4240 gnd.n6507 gnd.n257 240.244
R4241 gnd.n6507 gnd.n242 240.244
R4242 gnd.n6533 gnd.n242 240.244
R4243 gnd.n6533 gnd.n237 240.244
R4244 gnd.n6539 gnd.n237 240.244
R4245 gnd.n6539 gnd.n229 240.244
R4246 gnd.n6547 gnd.n229 240.244
R4247 gnd.n6547 gnd.n225 240.244
R4248 gnd.n6553 gnd.n225 240.244
R4249 gnd.n6553 gnd.n208 240.244
R4250 gnd.n6563 gnd.n208 240.244
R4251 gnd.n6563 gnd.n204 240.244
R4252 gnd.n6569 gnd.n204 240.244
R4253 gnd.n6569 gnd.n193 240.244
R4254 gnd.n6579 gnd.n193 240.244
R4255 gnd.n6579 gnd.n189 240.244
R4256 gnd.n6585 gnd.n189 240.244
R4257 gnd.n6585 gnd.n177 240.244
R4258 gnd.n6595 gnd.n177 240.244
R4259 gnd.n6595 gnd.n171 240.244
R4260 gnd.n6675 gnd.n171 240.244
R4261 gnd.n6675 gnd.n172 240.244
R4262 gnd.n172 gnd.n162 240.244
R4263 gnd.n6600 gnd.n162 240.244
R4264 gnd.n6600 gnd.n84 240.244
R4265 gnd.n1911 gnd.n1096 240.244
R4266 gnd.n1915 gnd.n1914 240.244
R4267 gnd.n1927 gnd.n1926 240.244
R4268 gnd.n1898 gnd.n1897 240.244
R4269 gnd.n1939 gnd.n1938 240.244
R4270 gnd.n1951 gnd.n1950 240.244
R4271 gnd.n1886 gnd.n1885 240.244
R4272 gnd.n1963 gnd.n1962 240.244
R4273 gnd.n1978 gnd.n1977 240.244
R4274 gnd.n3598 gnd.n2114 240.244
R4275 gnd.n3699 gnd.n2114 240.244
R4276 gnd.n3699 gnd.n2106 240.244
R4277 gnd.n3696 gnd.n2106 240.244
R4278 gnd.n3696 gnd.n2097 240.244
R4279 gnd.n3693 gnd.n2097 240.244
R4280 gnd.n3693 gnd.n2089 240.244
R4281 gnd.n3690 gnd.n2089 240.244
R4282 gnd.n3690 gnd.n2082 240.244
R4283 gnd.n3687 gnd.n2082 240.244
R4284 gnd.n3687 gnd.n2074 240.244
R4285 gnd.n3684 gnd.n2074 240.244
R4286 gnd.n3684 gnd.n2065 240.244
R4287 gnd.n3681 gnd.n2065 240.244
R4288 gnd.n3681 gnd.n2057 240.244
R4289 gnd.n3678 gnd.n2057 240.244
R4290 gnd.n3678 gnd.n2049 240.244
R4291 gnd.n3675 gnd.n2049 240.244
R4292 gnd.n3675 gnd.n2042 240.244
R4293 gnd.n3672 gnd.n2042 240.244
R4294 gnd.n3672 gnd.n2031 240.244
R4295 gnd.n2031 gnd.n2023 240.244
R4296 gnd.n4000 gnd.n2023 240.244
R4297 gnd.n4001 gnd.n4000 240.244
R4298 gnd.n4001 gnd.n1000 240.244
R4299 gnd.n4007 gnd.n1000 240.244
R4300 gnd.n4007 gnd.n1012 240.244
R4301 gnd.n4029 gnd.n1012 240.244
R4302 gnd.n4029 gnd.n1023 240.244
R4303 gnd.n4023 gnd.n1023 240.244
R4304 gnd.n4023 gnd.n1034 240.244
R4305 gnd.n4058 gnd.n1034 240.244
R4306 gnd.n4058 gnd.n1044 240.244
R4307 gnd.n4064 gnd.n1044 240.244
R4308 gnd.n4064 gnd.n1055 240.244
R4309 gnd.n4161 gnd.n1055 240.244
R4310 gnd.n4161 gnd.n1065 240.244
R4311 gnd.n1997 gnd.n1065 240.244
R4312 gnd.n1997 gnd.n1076 240.244
R4313 gnd.n4150 gnd.n1076 240.244
R4314 gnd.n4150 gnd.n1087 240.244
R4315 gnd.n4187 gnd.n1087 240.244
R4316 gnd.n3610 gnd.n2119 240.244
R4317 gnd.n3614 gnd.n3613 240.244
R4318 gnd.n3620 gnd.n3619 240.244
R4319 gnd.n3624 gnd.n3623 240.244
R4320 gnd.n3630 gnd.n3629 240.244
R4321 gnd.n3634 gnd.n3633 240.244
R4322 gnd.n3640 gnd.n3639 240.244
R4323 gnd.n3644 gnd.n3643 240.244
R4324 gnd.n3706 gnd.n3597 240.244
R4325 gnd.n3886 gnd.n2115 240.244
R4326 gnd.n3886 gnd.n2103 240.244
R4327 gnd.n3896 gnd.n2103 240.244
R4328 gnd.n3896 gnd.n2099 240.244
R4329 gnd.n3902 gnd.n2099 240.244
R4330 gnd.n3902 gnd.n2087 240.244
R4331 gnd.n3912 gnd.n2087 240.244
R4332 gnd.n3912 gnd.n2083 240.244
R4333 gnd.n3918 gnd.n2083 240.244
R4334 gnd.n3918 gnd.n2071 240.244
R4335 gnd.n3928 gnd.n2071 240.244
R4336 gnd.n3928 gnd.n2067 240.244
R4337 gnd.n3934 gnd.n2067 240.244
R4338 gnd.n3934 gnd.n2055 240.244
R4339 gnd.n3945 gnd.n2055 240.244
R4340 gnd.n3945 gnd.n2050 240.244
R4341 gnd.n3955 gnd.n2050 240.244
R4342 gnd.n3955 gnd.n2051 240.244
R4343 gnd.n2051 gnd.n2043 240.244
R4344 gnd.n2043 gnd.n2033 240.244
R4345 gnd.n3990 gnd.n2033 240.244
R4346 gnd.n3990 gnd.n2034 240.244
R4347 gnd.n2034 gnd.n2025 240.244
R4348 gnd.n3985 gnd.n2025 240.244
R4349 gnd.n3985 gnd.n1002 240.244
R4350 gnd.n1013 gnd.n1002 240.244
R4351 gnd.n5486 gnd.n1013 240.244
R4352 gnd.n5486 gnd.n1014 240.244
R4353 gnd.n5482 gnd.n1014 240.244
R4354 gnd.n5482 gnd.n1020 240.244
R4355 gnd.n5474 gnd.n1020 240.244
R4356 gnd.n5474 gnd.n1036 240.244
R4357 gnd.n5470 gnd.n1036 240.244
R4358 gnd.n5470 gnd.n1042 240.244
R4359 gnd.n5462 gnd.n1042 240.244
R4360 gnd.n5462 gnd.n1056 240.244
R4361 gnd.n5458 gnd.n1056 240.244
R4362 gnd.n5458 gnd.n1062 240.244
R4363 gnd.n5450 gnd.n1062 240.244
R4364 gnd.n5450 gnd.n1078 240.244
R4365 gnd.n5446 gnd.n1078 240.244
R4366 gnd.n5446 gnd.n1084 240.244
R4367 gnd.n5669 gnd.n827 240.244
R4368 gnd.n5669 gnd.n825 240.244
R4369 gnd.n5673 gnd.n825 240.244
R4370 gnd.n5673 gnd.n821 240.244
R4371 gnd.n5679 gnd.n821 240.244
R4372 gnd.n5679 gnd.n819 240.244
R4373 gnd.n5683 gnd.n819 240.244
R4374 gnd.n5683 gnd.n815 240.244
R4375 gnd.n5689 gnd.n815 240.244
R4376 gnd.n5689 gnd.n813 240.244
R4377 gnd.n5693 gnd.n813 240.244
R4378 gnd.n5693 gnd.n809 240.244
R4379 gnd.n5699 gnd.n809 240.244
R4380 gnd.n5699 gnd.n807 240.244
R4381 gnd.n5703 gnd.n807 240.244
R4382 gnd.n5703 gnd.n803 240.244
R4383 gnd.n5709 gnd.n803 240.244
R4384 gnd.n5709 gnd.n801 240.244
R4385 gnd.n5713 gnd.n801 240.244
R4386 gnd.n5713 gnd.n797 240.244
R4387 gnd.n5719 gnd.n797 240.244
R4388 gnd.n5719 gnd.n795 240.244
R4389 gnd.n5723 gnd.n795 240.244
R4390 gnd.n5723 gnd.n791 240.244
R4391 gnd.n5729 gnd.n791 240.244
R4392 gnd.n5729 gnd.n789 240.244
R4393 gnd.n5733 gnd.n789 240.244
R4394 gnd.n5733 gnd.n785 240.244
R4395 gnd.n5739 gnd.n785 240.244
R4396 gnd.n5739 gnd.n783 240.244
R4397 gnd.n5743 gnd.n783 240.244
R4398 gnd.n5743 gnd.n779 240.244
R4399 gnd.n5749 gnd.n779 240.244
R4400 gnd.n5749 gnd.n777 240.244
R4401 gnd.n5753 gnd.n777 240.244
R4402 gnd.n5753 gnd.n773 240.244
R4403 gnd.n5759 gnd.n773 240.244
R4404 gnd.n5759 gnd.n771 240.244
R4405 gnd.n5763 gnd.n771 240.244
R4406 gnd.n5763 gnd.n767 240.244
R4407 gnd.n5769 gnd.n767 240.244
R4408 gnd.n5769 gnd.n765 240.244
R4409 gnd.n5773 gnd.n765 240.244
R4410 gnd.n5773 gnd.n761 240.244
R4411 gnd.n5779 gnd.n761 240.244
R4412 gnd.n5779 gnd.n759 240.244
R4413 gnd.n5783 gnd.n759 240.244
R4414 gnd.n5783 gnd.n755 240.244
R4415 gnd.n5789 gnd.n755 240.244
R4416 gnd.n5789 gnd.n753 240.244
R4417 gnd.n5793 gnd.n753 240.244
R4418 gnd.n5793 gnd.n749 240.244
R4419 gnd.n5799 gnd.n749 240.244
R4420 gnd.n5799 gnd.n747 240.244
R4421 gnd.n5803 gnd.n747 240.244
R4422 gnd.n5803 gnd.n743 240.244
R4423 gnd.n5809 gnd.n743 240.244
R4424 gnd.n5809 gnd.n741 240.244
R4425 gnd.n5813 gnd.n741 240.244
R4426 gnd.n5813 gnd.n737 240.244
R4427 gnd.n5819 gnd.n737 240.244
R4428 gnd.n5819 gnd.n735 240.244
R4429 gnd.n5823 gnd.n735 240.244
R4430 gnd.n5823 gnd.n731 240.244
R4431 gnd.n5829 gnd.n731 240.244
R4432 gnd.n5829 gnd.n729 240.244
R4433 gnd.n5833 gnd.n729 240.244
R4434 gnd.n5833 gnd.n725 240.244
R4435 gnd.n5839 gnd.n725 240.244
R4436 gnd.n5839 gnd.n723 240.244
R4437 gnd.n5843 gnd.n723 240.244
R4438 gnd.n5843 gnd.n719 240.244
R4439 gnd.n5849 gnd.n719 240.244
R4440 gnd.n5849 gnd.n717 240.244
R4441 gnd.n5853 gnd.n717 240.244
R4442 gnd.n5853 gnd.n713 240.244
R4443 gnd.n5859 gnd.n713 240.244
R4444 gnd.n5859 gnd.n711 240.244
R4445 gnd.n5863 gnd.n711 240.244
R4446 gnd.n5863 gnd.n707 240.244
R4447 gnd.n5869 gnd.n707 240.244
R4448 gnd.n5869 gnd.n705 240.244
R4449 gnd.n5873 gnd.n705 240.244
R4450 gnd.n5873 gnd.n701 240.244
R4451 gnd.n5879 gnd.n701 240.244
R4452 gnd.n5879 gnd.n699 240.244
R4453 gnd.n5883 gnd.n699 240.244
R4454 gnd.n5883 gnd.n695 240.244
R4455 gnd.n5889 gnd.n695 240.244
R4456 gnd.n5889 gnd.n693 240.244
R4457 gnd.n5893 gnd.n693 240.244
R4458 gnd.n5893 gnd.n689 240.244
R4459 gnd.n5899 gnd.n689 240.244
R4460 gnd.n5899 gnd.n687 240.244
R4461 gnd.n5903 gnd.n687 240.244
R4462 gnd.n5903 gnd.n683 240.244
R4463 gnd.n5909 gnd.n683 240.244
R4464 gnd.n5909 gnd.n681 240.244
R4465 gnd.n5913 gnd.n681 240.244
R4466 gnd.n5913 gnd.n677 240.244
R4467 gnd.n5919 gnd.n677 240.244
R4468 gnd.n5919 gnd.n675 240.244
R4469 gnd.n5923 gnd.n675 240.244
R4470 gnd.n5923 gnd.n671 240.244
R4471 gnd.n5929 gnd.n671 240.244
R4472 gnd.n5929 gnd.n669 240.244
R4473 gnd.n5933 gnd.n669 240.244
R4474 gnd.n5933 gnd.n665 240.244
R4475 gnd.n5939 gnd.n665 240.244
R4476 gnd.n5939 gnd.n663 240.244
R4477 gnd.n5943 gnd.n663 240.244
R4478 gnd.n5943 gnd.n659 240.244
R4479 gnd.n5949 gnd.n659 240.244
R4480 gnd.n5949 gnd.n657 240.244
R4481 gnd.n5953 gnd.n657 240.244
R4482 gnd.n5953 gnd.n653 240.244
R4483 gnd.n5959 gnd.n653 240.244
R4484 gnd.n5959 gnd.n651 240.244
R4485 gnd.n5963 gnd.n651 240.244
R4486 gnd.n5963 gnd.n647 240.244
R4487 gnd.n5969 gnd.n647 240.244
R4488 gnd.n5969 gnd.n645 240.244
R4489 gnd.n5973 gnd.n645 240.244
R4490 gnd.n5973 gnd.n641 240.244
R4491 gnd.n5980 gnd.n641 240.244
R4492 gnd.n5980 gnd.n639 240.244
R4493 gnd.n5984 gnd.n639 240.244
R4494 gnd.n5984 gnd.n636 240.244
R4495 gnd.n5990 gnd.n634 240.244
R4496 gnd.n5994 gnd.n634 240.244
R4497 gnd.n5994 gnd.n630 240.244
R4498 gnd.n6000 gnd.n630 240.244
R4499 gnd.n6000 gnd.n628 240.244
R4500 gnd.n6004 gnd.n628 240.244
R4501 gnd.n6004 gnd.n624 240.244
R4502 gnd.n6010 gnd.n624 240.244
R4503 gnd.n6010 gnd.n622 240.244
R4504 gnd.n6014 gnd.n622 240.244
R4505 gnd.n6014 gnd.n618 240.244
R4506 gnd.n6020 gnd.n618 240.244
R4507 gnd.n6020 gnd.n616 240.244
R4508 gnd.n6024 gnd.n616 240.244
R4509 gnd.n6024 gnd.n612 240.244
R4510 gnd.n6030 gnd.n612 240.244
R4511 gnd.n6030 gnd.n610 240.244
R4512 gnd.n6034 gnd.n610 240.244
R4513 gnd.n6034 gnd.n606 240.244
R4514 gnd.n6040 gnd.n606 240.244
R4515 gnd.n6040 gnd.n604 240.244
R4516 gnd.n6044 gnd.n604 240.244
R4517 gnd.n6044 gnd.n600 240.244
R4518 gnd.n6050 gnd.n600 240.244
R4519 gnd.n6050 gnd.n598 240.244
R4520 gnd.n6054 gnd.n598 240.244
R4521 gnd.n6054 gnd.n594 240.244
R4522 gnd.n6060 gnd.n594 240.244
R4523 gnd.n6060 gnd.n592 240.244
R4524 gnd.n6064 gnd.n592 240.244
R4525 gnd.n6064 gnd.n588 240.244
R4526 gnd.n6070 gnd.n588 240.244
R4527 gnd.n6070 gnd.n586 240.244
R4528 gnd.n6074 gnd.n586 240.244
R4529 gnd.n6074 gnd.n582 240.244
R4530 gnd.n6080 gnd.n582 240.244
R4531 gnd.n6080 gnd.n580 240.244
R4532 gnd.n6084 gnd.n580 240.244
R4533 gnd.n6084 gnd.n576 240.244
R4534 gnd.n6090 gnd.n576 240.244
R4535 gnd.n6090 gnd.n574 240.244
R4536 gnd.n6094 gnd.n574 240.244
R4537 gnd.n6094 gnd.n570 240.244
R4538 gnd.n6100 gnd.n570 240.244
R4539 gnd.n6100 gnd.n568 240.244
R4540 gnd.n6104 gnd.n568 240.244
R4541 gnd.n6104 gnd.n564 240.244
R4542 gnd.n6110 gnd.n564 240.244
R4543 gnd.n6110 gnd.n562 240.244
R4544 gnd.n6114 gnd.n562 240.244
R4545 gnd.n6114 gnd.n558 240.244
R4546 gnd.n6120 gnd.n558 240.244
R4547 gnd.n6120 gnd.n556 240.244
R4548 gnd.n6124 gnd.n556 240.244
R4549 gnd.n6124 gnd.n552 240.244
R4550 gnd.n6130 gnd.n552 240.244
R4551 gnd.n6130 gnd.n550 240.244
R4552 gnd.n6134 gnd.n550 240.244
R4553 gnd.n6134 gnd.n546 240.244
R4554 gnd.n6140 gnd.n546 240.244
R4555 gnd.n6140 gnd.n544 240.244
R4556 gnd.n6144 gnd.n544 240.244
R4557 gnd.n6144 gnd.n540 240.244
R4558 gnd.n6150 gnd.n540 240.244
R4559 gnd.n6150 gnd.n538 240.244
R4560 gnd.n6154 gnd.n538 240.244
R4561 gnd.n6154 gnd.n534 240.244
R4562 gnd.n6160 gnd.n534 240.244
R4563 gnd.n6160 gnd.n532 240.244
R4564 gnd.n6164 gnd.n532 240.244
R4565 gnd.n6164 gnd.n528 240.244
R4566 gnd.n6170 gnd.n528 240.244
R4567 gnd.n6170 gnd.n526 240.244
R4568 gnd.n6174 gnd.n526 240.244
R4569 gnd.n6174 gnd.n522 240.244
R4570 gnd.n6180 gnd.n522 240.244
R4571 gnd.n6180 gnd.n520 240.244
R4572 gnd.n6184 gnd.n520 240.244
R4573 gnd.n6184 gnd.n516 240.244
R4574 gnd.n6190 gnd.n516 240.244
R4575 gnd.n6190 gnd.n514 240.244
R4576 gnd.n6195 gnd.n514 240.244
R4577 gnd.n6195 gnd.n510 240.244
R4578 gnd.n6202 gnd.n510 240.244
R4579 gnd.n4037 gnd.n997 240.244
R4580 gnd.n4037 gnd.n4032 240.244
R4581 gnd.n4043 gnd.n4032 240.244
R4582 gnd.n4044 gnd.n4043 240.244
R4583 gnd.n4045 gnd.n4044 240.244
R4584 gnd.n4045 gnd.n2007 240.244
R4585 gnd.n4055 gnd.n2007 240.244
R4586 gnd.n4055 gnd.n2008 240.244
R4587 gnd.n2008 gnd.n1991 240.244
R4588 gnd.n4164 gnd.n1991 240.244
R4589 gnd.n4165 gnd.n4164 240.244
R4590 gnd.n4165 gnd.n1987 240.244
R4591 gnd.n4171 gnd.n1987 240.244
R4592 gnd.n4172 gnd.n4171 240.244
R4593 gnd.n4173 gnd.n4172 240.244
R4594 gnd.n4173 gnd.n1982 240.244
R4595 gnd.n4184 gnd.n1982 240.244
R4596 gnd.n4184 gnd.n1983 240.244
R4597 gnd.n4180 gnd.n1983 240.244
R4598 gnd.n4180 gnd.n1846 240.244
R4599 gnd.n4235 gnd.n1846 240.244
R4600 gnd.n4235 gnd.n1841 240.244
R4601 gnd.n4250 gnd.n1841 240.244
R4602 gnd.n4250 gnd.n1842 240.244
R4603 gnd.n4246 gnd.n1842 240.244
R4604 gnd.n4246 gnd.n4245 240.244
R4605 gnd.n4245 gnd.n1213 240.244
R4606 gnd.n5331 gnd.n1213 240.244
R4607 gnd.n5331 gnd.n1214 240.244
R4608 gnd.n5327 gnd.n1214 240.244
R4609 gnd.n5327 gnd.n1220 240.244
R4610 gnd.n1313 gnd.n1220 240.244
R4611 gnd.n5312 gnd.n1313 240.244
R4612 gnd.n5312 gnd.n1314 240.244
R4613 gnd.n5308 gnd.n1314 240.244
R4614 gnd.n5308 gnd.n1322 240.244
R4615 gnd.n4431 gnd.n1322 240.244
R4616 gnd.n4437 gnd.n4431 240.244
R4617 gnd.n4437 gnd.n1804 240.244
R4618 gnd.n4460 gnd.n1804 240.244
R4619 gnd.n4460 gnd.n1799 240.244
R4620 gnd.n4477 gnd.n1799 240.244
R4621 gnd.n4477 gnd.n1800 240.244
R4622 gnd.n4473 gnd.n1800 240.244
R4623 gnd.n4473 gnd.n4472 240.244
R4624 gnd.n4472 gnd.n4471 240.244
R4625 gnd.n4471 gnd.n1766 240.244
R4626 gnd.n4518 gnd.n1766 240.244
R4627 gnd.n4518 gnd.n1762 240.244
R4628 gnd.n4524 gnd.n1762 240.244
R4629 gnd.n4524 gnd.n1748 240.244
R4630 gnd.n4544 gnd.n1748 240.244
R4631 gnd.n4544 gnd.n1743 240.244
R4632 gnd.n4552 gnd.n1743 240.244
R4633 gnd.n4552 gnd.n1744 240.244
R4634 gnd.n1744 gnd.n1724 240.244
R4635 gnd.n4583 gnd.n1724 240.244
R4636 gnd.n4583 gnd.n1719 240.244
R4637 gnd.n4600 gnd.n1719 240.244
R4638 gnd.n4600 gnd.n1720 240.244
R4639 gnd.n4596 gnd.n1720 240.244
R4640 gnd.n4596 gnd.n4595 240.244
R4641 gnd.n4595 gnd.n4594 240.244
R4642 gnd.n4594 gnd.n1685 240.244
R4643 gnd.n4641 gnd.n1685 240.244
R4644 gnd.n4641 gnd.n1681 240.244
R4645 gnd.n4647 gnd.n1681 240.244
R4646 gnd.n4647 gnd.n1666 240.244
R4647 gnd.n4666 gnd.n1666 240.244
R4648 gnd.n4666 gnd.n1661 240.244
R4649 gnd.n4674 gnd.n1661 240.244
R4650 gnd.n4674 gnd.n1662 240.244
R4651 gnd.n1662 gnd.n1641 240.244
R4652 gnd.n4705 gnd.n1641 240.244
R4653 gnd.n4705 gnd.n1637 240.244
R4654 gnd.n4711 gnd.n1637 240.244
R4655 gnd.n4711 gnd.n1618 240.244
R4656 gnd.n4751 gnd.n1618 240.244
R4657 gnd.n4751 gnd.n1613 240.244
R4658 gnd.n4759 gnd.n1613 240.244
R4659 gnd.n4759 gnd.n1614 240.244
R4660 gnd.n1614 gnd.n1597 240.244
R4661 gnd.n4806 gnd.n1597 240.244
R4662 gnd.n4806 gnd.n1592 240.244
R4663 gnd.n4814 gnd.n1592 240.244
R4664 gnd.n4814 gnd.n1593 240.244
R4665 gnd.n1593 gnd.n1570 240.244
R4666 gnd.n4843 gnd.n1570 240.244
R4667 gnd.n4843 gnd.n1566 240.244
R4668 gnd.n4849 gnd.n1566 240.244
R4669 gnd.n4849 gnd.n1552 240.244
R4670 gnd.n4869 gnd.n1552 240.244
R4671 gnd.n4869 gnd.n1547 240.244
R4672 gnd.n4877 gnd.n1547 240.244
R4673 gnd.n4877 gnd.n1548 240.244
R4674 gnd.n1548 gnd.n1524 240.244
R4675 gnd.n4922 gnd.n1524 240.244
R4676 gnd.n4922 gnd.n1520 240.244
R4677 gnd.n4928 gnd.n1520 240.244
R4678 gnd.n4928 gnd.n1432 240.244
R4679 gnd.n5065 gnd.n1432 240.244
R4680 gnd.n5065 gnd.n1427 240.244
R4681 gnd.n5188 gnd.n1427 240.244
R4682 gnd.n5188 gnd.n1428 240.244
R4683 gnd.n1428 gnd.n1420 240.244
R4684 gnd.n5183 gnd.n1420 240.244
R4685 gnd.n5183 gnd.n5182 240.244
R4686 gnd.n5182 gnd.n5074 240.244
R4687 gnd.n5116 gnd.n5074 240.244
R4688 gnd.n5117 gnd.n5116 240.244
R4689 gnd.n5118 gnd.n5117 240.244
R4690 gnd.n5118 gnd.n5106 240.244
R4691 gnd.n5148 gnd.n5106 240.244
R4692 gnd.n5148 gnd.n5107 240.244
R4693 gnd.n5144 gnd.n5107 240.244
R4694 gnd.n5144 gnd.n5143 240.244
R4695 gnd.n5143 gnd.n5142 240.244
R4696 gnd.n5142 gnd.n5126 240.244
R4697 gnd.n5138 gnd.n5126 240.244
R4698 gnd.n5138 gnd.n5137 240.244
R4699 gnd.n5137 gnd.n5136 240.244
R4700 gnd.n5136 gnd.n503 240.244
R4701 gnd.n6215 gnd.n503 240.244
R4702 gnd.n6215 gnd.n504 240.244
R4703 gnd.n6211 gnd.n504 240.244
R4704 gnd.n6211 gnd.n6210 240.244
R4705 gnd.n6210 gnd.n6209 240.244
R4706 gnd.n6209 gnd.n6203 240.244
R4707 gnd.n5663 gnd.n831 240.244
R4708 gnd.n5659 gnd.n831 240.244
R4709 gnd.n5659 gnd.n833 240.244
R4710 gnd.n5655 gnd.n833 240.244
R4711 gnd.n5655 gnd.n838 240.244
R4712 gnd.n5651 gnd.n838 240.244
R4713 gnd.n5651 gnd.n840 240.244
R4714 gnd.n5647 gnd.n840 240.244
R4715 gnd.n5647 gnd.n846 240.244
R4716 gnd.n5643 gnd.n846 240.244
R4717 gnd.n5643 gnd.n848 240.244
R4718 gnd.n5639 gnd.n848 240.244
R4719 gnd.n5639 gnd.n854 240.244
R4720 gnd.n5635 gnd.n854 240.244
R4721 gnd.n5635 gnd.n856 240.244
R4722 gnd.n5631 gnd.n856 240.244
R4723 gnd.n5631 gnd.n862 240.244
R4724 gnd.n5627 gnd.n862 240.244
R4725 gnd.n5627 gnd.n864 240.244
R4726 gnd.n5623 gnd.n864 240.244
R4727 gnd.n5623 gnd.n870 240.244
R4728 gnd.n5619 gnd.n870 240.244
R4729 gnd.n5619 gnd.n872 240.244
R4730 gnd.n5615 gnd.n872 240.244
R4731 gnd.n5615 gnd.n878 240.244
R4732 gnd.n5611 gnd.n878 240.244
R4733 gnd.n5611 gnd.n880 240.244
R4734 gnd.n5607 gnd.n880 240.244
R4735 gnd.n5607 gnd.n886 240.244
R4736 gnd.n5603 gnd.n886 240.244
R4737 gnd.n5603 gnd.n888 240.244
R4738 gnd.n5599 gnd.n888 240.244
R4739 gnd.n5599 gnd.n894 240.244
R4740 gnd.n5595 gnd.n894 240.244
R4741 gnd.n5595 gnd.n896 240.244
R4742 gnd.n5591 gnd.n896 240.244
R4743 gnd.n5591 gnd.n902 240.244
R4744 gnd.n5587 gnd.n902 240.244
R4745 gnd.n5587 gnd.n904 240.244
R4746 gnd.n5583 gnd.n904 240.244
R4747 gnd.n5583 gnd.n910 240.244
R4748 gnd.n5579 gnd.n910 240.244
R4749 gnd.n5579 gnd.n912 240.244
R4750 gnd.n5575 gnd.n912 240.244
R4751 gnd.n5575 gnd.n918 240.244
R4752 gnd.n5571 gnd.n918 240.244
R4753 gnd.n5571 gnd.n920 240.244
R4754 gnd.n5567 gnd.n920 240.244
R4755 gnd.n5567 gnd.n926 240.244
R4756 gnd.n5563 gnd.n926 240.244
R4757 gnd.n5563 gnd.n928 240.244
R4758 gnd.n5559 gnd.n928 240.244
R4759 gnd.n5559 gnd.n934 240.244
R4760 gnd.n5555 gnd.n934 240.244
R4761 gnd.n5555 gnd.n936 240.244
R4762 gnd.n5551 gnd.n936 240.244
R4763 gnd.n5551 gnd.n942 240.244
R4764 gnd.n5547 gnd.n942 240.244
R4765 gnd.n5547 gnd.n944 240.244
R4766 gnd.n5543 gnd.n944 240.244
R4767 gnd.n5543 gnd.n950 240.244
R4768 gnd.n5539 gnd.n950 240.244
R4769 gnd.n5539 gnd.n952 240.244
R4770 gnd.n5535 gnd.n952 240.244
R4771 gnd.n5535 gnd.n958 240.244
R4772 gnd.n5531 gnd.n958 240.244
R4773 gnd.n5531 gnd.n960 240.244
R4774 gnd.n5527 gnd.n960 240.244
R4775 gnd.n5527 gnd.n966 240.244
R4776 gnd.n5523 gnd.n966 240.244
R4777 gnd.n5523 gnd.n968 240.244
R4778 gnd.n5519 gnd.n968 240.244
R4779 gnd.n5519 gnd.n974 240.244
R4780 gnd.n5515 gnd.n974 240.244
R4781 gnd.n5515 gnd.n976 240.244
R4782 gnd.n5511 gnd.n976 240.244
R4783 gnd.n5511 gnd.n982 240.244
R4784 gnd.n5507 gnd.n982 240.244
R4785 gnd.n5507 gnd.n984 240.244
R4786 gnd.n5503 gnd.n984 240.244
R4787 gnd.n5503 gnd.n990 240.244
R4788 gnd.n5499 gnd.n990 240.244
R4789 gnd.n5499 gnd.n992 240.244
R4790 gnd.n5495 gnd.n992 240.244
R4791 gnd.n4252 gnd.n1834 240.244
R4792 gnd.n4258 gnd.n1834 240.244
R4793 gnd.n4259 gnd.n4258 240.244
R4794 gnd.n4260 gnd.n4259 240.244
R4795 gnd.n4260 gnd.n1210 240.244
R4796 gnd.n4266 gnd.n1210 240.244
R4797 gnd.n4266 gnd.n1222 240.244
R4798 gnd.n4285 gnd.n1222 240.244
R4799 gnd.n4285 gnd.n1825 240.244
R4800 gnd.n1825 gnd.n1310 240.244
R4801 gnd.n4320 gnd.n1310 240.244
R4802 gnd.n4320 gnd.n1324 240.244
R4803 gnd.n1818 gnd.n1324 240.244
R4804 gnd.n4429 gnd.n1818 240.244
R4805 gnd.n4429 gnd.n1816 240.244
R4806 gnd.n1816 gnd.n1812 240.244
R4807 gnd.n1812 gnd.n1805 240.244
R4808 gnd.n4326 gnd.n1805 240.244
R4809 gnd.n4326 gnd.n1798 240.244
R4810 gnd.n4329 gnd.n1798 240.244
R4811 gnd.n4330 gnd.n4329 240.244
R4812 gnd.n4331 gnd.n4330 240.244
R4813 gnd.n4332 gnd.n4331 240.244
R4814 gnd.n4332 gnd.n1773 240.244
R4815 gnd.n1773 gnd.n1767 240.244
R4816 gnd.n4335 gnd.n1767 240.244
R4817 gnd.n4335 gnd.n1760 240.244
R4818 gnd.n4338 gnd.n1760 240.244
R4819 gnd.n4338 gnd.n1749 240.244
R4820 gnd.n4339 gnd.n1749 240.244
R4821 gnd.n4339 gnd.n1742 240.244
R4822 gnd.n4342 gnd.n1742 240.244
R4823 gnd.n4342 gnd.n1733 240.244
R4824 gnd.n1733 gnd.n1725 240.244
R4825 gnd.n4343 gnd.n1725 240.244
R4826 gnd.n4343 gnd.n1718 240.244
R4827 gnd.n4346 gnd.n1718 240.244
R4828 gnd.n4347 gnd.n4346 240.244
R4829 gnd.n4350 gnd.n4347 240.244
R4830 gnd.n4351 gnd.n4350 240.244
R4831 gnd.n4351 gnd.n1694 240.244
R4832 gnd.n1694 gnd.n1687 240.244
R4833 gnd.n4352 gnd.n1687 240.244
R4834 gnd.n4352 gnd.n1679 240.244
R4835 gnd.n4355 gnd.n1679 240.244
R4836 gnd.n4355 gnd.n1667 240.244
R4837 gnd.n4356 gnd.n1667 240.244
R4838 gnd.n4356 gnd.n1660 240.244
R4839 gnd.n4359 gnd.n1660 240.244
R4840 gnd.n4359 gnd.n1650 240.244
R4841 gnd.n1650 gnd.n1642 240.244
R4842 gnd.n4363 gnd.n1642 240.244
R4843 gnd.n4363 gnd.n1635 240.244
R4844 gnd.n4364 gnd.n1635 240.244
R4845 gnd.n4364 gnd.n1620 240.244
R4846 gnd.n1620 gnd.n1610 240.244
R4847 gnd.n4761 gnd.n1610 240.244
R4848 gnd.n4761 gnd.n1605 240.244
R4849 gnd.n4796 gnd.n1605 240.244
R4850 gnd.n4796 gnd.n1599 240.244
R4851 gnd.n4766 gnd.n1599 240.244
R4852 gnd.n4766 gnd.n1591 240.244
R4853 gnd.n4767 gnd.n1591 240.244
R4854 gnd.n4768 gnd.n4767 240.244
R4855 gnd.n4768 gnd.n1572 240.244
R4856 gnd.n4771 gnd.n1572 240.244
R4857 gnd.n4771 gnd.n1564 240.244
R4858 gnd.n4772 gnd.n1564 240.244
R4859 gnd.n4772 gnd.n1554 240.244
R4860 gnd.n4775 gnd.n1554 240.244
R4861 gnd.n4775 gnd.n1546 240.244
R4862 gnd.n1546 gnd.n1533 240.244
R4863 gnd.n4911 gnd.n1533 240.244
R4864 gnd.n4911 gnd.n1526 240.244
R4865 gnd.n4899 gnd.n1526 240.244
R4866 gnd.n4899 gnd.n1518 240.244
R4867 gnd.n4900 gnd.n1518 240.244
R4868 gnd.n4900 gnd.n1434 240.244
R4869 gnd.n1434 gnd.n1426 240.244
R4870 gnd.n5190 gnd.n1426 240.244
R4871 gnd.n5190 gnd.n1422 240.244
R4872 gnd.n5196 gnd.n1422 240.244
R4873 gnd.n1921 gnd.n1920 240.244
R4874 gnd.n1902 gnd.n1901 240.244
R4875 gnd.n1933 gnd.n1932 240.244
R4876 gnd.n1945 gnd.n1944 240.244
R4877 gnd.n1890 gnd.n1889 240.244
R4878 gnd.n1957 gnd.n1956 240.244
R4879 gnd.n1969 gnd.n1968 240.244
R4880 gnd.n1878 gnd.n1877 240.244
R4881 gnd.n4195 gnd.n4194 240.244
R4882 gnd.n1873 gnd.n1872 240.244
R4883 gnd.n4204 gnd.n4203 240.244
R4884 gnd.n1869 gnd.n1868 240.244
R4885 gnd.n4213 gnd.n4212 240.244
R4886 gnd.n4233 gnd.n1862 240.244
R4887 gnd.n4218 gnd.n1840 240.244
R4888 gnd.n4219 gnd.n4218 240.244
R4889 gnd.n4221 gnd.n4219 240.244
R4890 gnd.n4222 gnd.n4221 240.244
R4891 gnd.n4222 gnd.n1212 240.244
R4892 gnd.n4274 gnd.n1212 240.244
R4893 gnd.n4274 gnd.n1224 240.244
R4894 gnd.n4283 gnd.n1224 240.244
R4895 gnd.n4283 gnd.n1826 240.244
R4896 gnd.n1826 gnd.n1312 240.244
R4897 gnd.n1326 gnd.n1312 240.244
R4898 gnd.n5306 gnd.n1326 240.244
R4899 gnd.n5306 gnd.n1327 240.244
R4900 gnd.n1332 gnd.n1327 240.244
R4901 gnd.n1333 gnd.n1332 240.244
R4902 gnd.n1334 gnd.n1333 240.244
R4903 gnd.n4458 gnd.n1334 240.244
R4904 gnd.n4458 gnd.n1337 240.244
R4905 gnd.n1338 gnd.n1337 240.244
R4906 gnd.n1339 gnd.n1338 240.244
R4907 gnd.n1785 gnd.n1339 240.244
R4908 gnd.n1785 gnd.n1342 240.244
R4909 gnd.n1343 gnd.n1342 240.244
R4910 gnd.n1344 gnd.n1343 240.244
R4911 gnd.n4516 gnd.n1344 240.244
R4912 gnd.n4516 gnd.n1347 240.244
R4913 gnd.n1348 gnd.n1347 240.244
R4914 gnd.n1349 gnd.n1348 240.244
R4915 gnd.n4542 gnd.n1349 240.244
R4916 gnd.n4542 gnd.n1352 240.244
R4917 gnd.n1353 gnd.n1352 240.244
R4918 gnd.n1354 gnd.n1353 240.244
R4919 gnd.n4573 gnd.n1354 240.244
R4920 gnd.n4573 gnd.n1357 240.244
R4921 gnd.n1358 gnd.n1357 240.244
R4922 gnd.n1359 gnd.n1358 240.244
R4923 gnd.n1711 gnd.n1359 240.244
R4924 gnd.n1711 gnd.n1362 240.244
R4925 gnd.n1363 gnd.n1362 240.244
R4926 gnd.n1364 gnd.n1363 240.244
R4927 gnd.n1695 gnd.n1364 240.244
R4928 gnd.n1695 gnd.n1367 240.244
R4929 gnd.n1368 gnd.n1367 240.244
R4930 gnd.n1369 gnd.n1368 240.244
R4931 gnd.n1671 gnd.n1369 240.244
R4932 gnd.n1671 gnd.n1372 240.244
R4933 gnd.n1373 gnd.n1372 240.244
R4934 gnd.n1374 gnd.n1373 240.244
R4935 gnd.n1653 gnd.n1374 240.244
R4936 gnd.n1653 gnd.n1377 240.244
R4937 gnd.n1378 gnd.n1377 240.244
R4938 gnd.n1379 gnd.n1378 240.244
R4939 gnd.n1636 gnd.n1379 240.244
R4940 gnd.n1636 gnd.n1382 240.244
R4941 gnd.n1383 gnd.n1382 240.244
R4942 gnd.n1384 gnd.n1383 240.244
R4943 gnd.n1612 gnd.n1384 240.244
R4944 gnd.n1612 gnd.n1387 240.244
R4945 gnd.n1388 gnd.n1387 240.244
R4946 gnd.n1389 gnd.n1388 240.244
R4947 gnd.n1588 gnd.n1389 240.244
R4948 gnd.n1588 gnd.n1392 240.244
R4949 gnd.n1393 gnd.n1392 240.244
R4950 gnd.n1394 gnd.n1393 240.244
R4951 gnd.n4841 gnd.n1394 240.244
R4952 gnd.n4841 gnd.n1397 240.244
R4953 gnd.n1398 gnd.n1397 240.244
R4954 gnd.n1399 gnd.n1398 240.244
R4955 gnd.n4867 gnd.n1399 240.244
R4956 gnd.n4867 gnd.n1402 240.244
R4957 gnd.n1403 gnd.n1402 240.244
R4958 gnd.n1404 gnd.n1403 240.244
R4959 gnd.n4912 gnd.n1404 240.244
R4960 gnd.n4912 gnd.n1407 240.244
R4961 gnd.n1408 gnd.n1407 240.244
R4962 gnd.n1409 gnd.n1408 240.244
R4963 gnd.n1512 gnd.n1409 240.244
R4964 gnd.n1512 gnd.n1412 240.244
R4965 gnd.n1413 gnd.n1412 240.244
R4966 gnd.n1414 gnd.n1413 240.244
R4967 gnd.n1417 gnd.n1414 240.244
R4968 gnd.n5198 gnd.n1417 240.244
R4969 gnd.n5076 gnd.n338 240.244
R4970 gnd.n346 gnd.n345 240.244
R4971 gnd.n5078 gnd.n353 240.244
R4972 gnd.n5081 gnd.n354 240.244
R4973 gnd.n362 gnd.n361 240.244
R4974 gnd.n5083 gnd.n369 240.244
R4975 gnd.n5086 gnd.n370 240.244
R4976 gnd.n380 gnd.n379 240.244
R4977 gnd.n5102 gnd.n5101 240.244
R4978 gnd.n5159 gnd.n5158 240.244
R4979 gnd.n5162 gnd.n5161 240.244
R4980 gnd.n5169 gnd.n5168 240.244
R4981 gnd.n5172 gnd.n5093 240.244
R4982 gnd.n5178 gnd.n1418 240.244
R4983 gnd.n1191 gnd.n1190 240.132
R4984 gnd.n1451 gnd.n1450 240.132
R4985 gnd.n5670 gnd.n826 225.874
R4986 gnd.n5671 gnd.n5670 225.874
R4987 gnd.n5672 gnd.n5671 225.874
R4988 gnd.n5672 gnd.n820 225.874
R4989 gnd.n5680 gnd.n820 225.874
R4990 gnd.n5681 gnd.n5680 225.874
R4991 gnd.n5682 gnd.n5681 225.874
R4992 gnd.n5682 gnd.n814 225.874
R4993 gnd.n5690 gnd.n814 225.874
R4994 gnd.n5691 gnd.n5690 225.874
R4995 gnd.n5692 gnd.n5691 225.874
R4996 gnd.n5692 gnd.n808 225.874
R4997 gnd.n5700 gnd.n808 225.874
R4998 gnd.n5701 gnd.n5700 225.874
R4999 gnd.n5702 gnd.n5701 225.874
R5000 gnd.n5702 gnd.n802 225.874
R5001 gnd.n5710 gnd.n802 225.874
R5002 gnd.n5711 gnd.n5710 225.874
R5003 gnd.n5712 gnd.n5711 225.874
R5004 gnd.n5712 gnd.n796 225.874
R5005 gnd.n5720 gnd.n796 225.874
R5006 gnd.n5721 gnd.n5720 225.874
R5007 gnd.n5722 gnd.n5721 225.874
R5008 gnd.n5722 gnd.n790 225.874
R5009 gnd.n5730 gnd.n790 225.874
R5010 gnd.n5731 gnd.n5730 225.874
R5011 gnd.n5732 gnd.n5731 225.874
R5012 gnd.n5732 gnd.n784 225.874
R5013 gnd.n5740 gnd.n784 225.874
R5014 gnd.n5741 gnd.n5740 225.874
R5015 gnd.n5742 gnd.n5741 225.874
R5016 gnd.n5742 gnd.n778 225.874
R5017 gnd.n5750 gnd.n778 225.874
R5018 gnd.n5751 gnd.n5750 225.874
R5019 gnd.n5752 gnd.n5751 225.874
R5020 gnd.n5752 gnd.n772 225.874
R5021 gnd.n5760 gnd.n772 225.874
R5022 gnd.n5761 gnd.n5760 225.874
R5023 gnd.n5762 gnd.n5761 225.874
R5024 gnd.n5762 gnd.n766 225.874
R5025 gnd.n5770 gnd.n766 225.874
R5026 gnd.n5771 gnd.n5770 225.874
R5027 gnd.n5772 gnd.n5771 225.874
R5028 gnd.n5772 gnd.n760 225.874
R5029 gnd.n5780 gnd.n760 225.874
R5030 gnd.n5781 gnd.n5780 225.874
R5031 gnd.n5782 gnd.n5781 225.874
R5032 gnd.n5782 gnd.n754 225.874
R5033 gnd.n5790 gnd.n754 225.874
R5034 gnd.n5791 gnd.n5790 225.874
R5035 gnd.n5792 gnd.n5791 225.874
R5036 gnd.n5792 gnd.n748 225.874
R5037 gnd.n5800 gnd.n748 225.874
R5038 gnd.n5801 gnd.n5800 225.874
R5039 gnd.n5802 gnd.n5801 225.874
R5040 gnd.n5802 gnd.n742 225.874
R5041 gnd.n5810 gnd.n742 225.874
R5042 gnd.n5811 gnd.n5810 225.874
R5043 gnd.n5812 gnd.n5811 225.874
R5044 gnd.n5812 gnd.n736 225.874
R5045 gnd.n5820 gnd.n736 225.874
R5046 gnd.n5821 gnd.n5820 225.874
R5047 gnd.n5822 gnd.n5821 225.874
R5048 gnd.n5822 gnd.n730 225.874
R5049 gnd.n5830 gnd.n730 225.874
R5050 gnd.n5831 gnd.n5830 225.874
R5051 gnd.n5832 gnd.n5831 225.874
R5052 gnd.n5832 gnd.n724 225.874
R5053 gnd.n5840 gnd.n724 225.874
R5054 gnd.n5841 gnd.n5840 225.874
R5055 gnd.n5842 gnd.n5841 225.874
R5056 gnd.n5842 gnd.n718 225.874
R5057 gnd.n5850 gnd.n718 225.874
R5058 gnd.n5851 gnd.n5850 225.874
R5059 gnd.n5852 gnd.n5851 225.874
R5060 gnd.n5852 gnd.n712 225.874
R5061 gnd.n5860 gnd.n712 225.874
R5062 gnd.n5861 gnd.n5860 225.874
R5063 gnd.n5862 gnd.n5861 225.874
R5064 gnd.n5862 gnd.n706 225.874
R5065 gnd.n5870 gnd.n706 225.874
R5066 gnd.n5871 gnd.n5870 225.874
R5067 gnd.n5872 gnd.n5871 225.874
R5068 gnd.n5872 gnd.n700 225.874
R5069 gnd.n5880 gnd.n700 225.874
R5070 gnd.n5881 gnd.n5880 225.874
R5071 gnd.n5882 gnd.n5881 225.874
R5072 gnd.n5882 gnd.n694 225.874
R5073 gnd.n5890 gnd.n694 225.874
R5074 gnd.n5891 gnd.n5890 225.874
R5075 gnd.n5892 gnd.n5891 225.874
R5076 gnd.n5892 gnd.n688 225.874
R5077 gnd.n5900 gnd.n688 225.874
R5078 gnd.n5901 gnd.n5900 225.874
R5079 gnd.n5902 gnd.n5901 225.874
R5080 gnd.n5902 gnd.n682 225.874
R5081 gnd.n5910 gnd.n682 225.874
R5082 gnd.n5911 gnd.n5910 225.874
R5083 gnd.n5912 gnd.n5911 225.874
R5084 gnd.n5912 gnd.n676 225.874
R5085 gnd.n5920 gnd.n676 225.874
R5086 gnd.n5921 gnd.n5920 225.874
R5087 gnd.n5922 gnd.n5921 225.874
R5088 gnd.n5922 gnd.n670 225.874
R5089 gnd.n5930 gnd.n670 225.874
R5090 gnd.n5931 gnd.n5930 225.874
R5091 gnd.n5932 gnd.n5931 225.874
R5092 gnd.n5932 gnd.n664 225.874
R5093 gnd.n5940 gnd.n664 225.874
R5094 gnd.n5941 gnd.n5940 225.874
R5095 gnd.n5942 gnd.n5941 225.874
R5096 gnd.n5942 gnd.n658 225.874
R5097 gnd.n5950 gnd.n658 225.874
R5098 gnd.n5951 gnd.n5950 225.874
R5099 gnd.n5952 gnd.n5951 225.874
R5100 gnd.n5952 gnd.n652 225.874
R5101 gnd.n5960 gnd.n652 225.874
R5102 gnd.n5961 gnd.n5960 225.874
R5103 gnd.n5962 gnd.n5961 225.874
R5104 gnd.n5962 gnd.n646 225.874
R5105 gnd.n5970 gnd.n646 225.874
R5106 gnd.n5971 gnd.n5970 225.874
R5107 gnd.n5972 gnd.n5971 225.874
R5108 gnd.n5972 gnd.n640 225.874
R5109 gnd.n5981 gnd.n640 225.874
R5110 gnd.n5982 gnd.n5981 225.874
R5111 gnd.n5983 gnd.n5982 225.874
R5112 gnd.n5983 gnd.n635 225.874
R5113 gnd.n2663 gnd.t177 224.174
R5114 gnd.n2185 gnd.t110 224.174
R5115 gnd.n436 gnd.n391 199.319
R5116 gnd.n436 gnd.n392 199.319
R5117 gnd.n1143 gnd.n1118 199.319
R5118 gnd.n1143 gnd.n1117 199.319
R5119 gnd.n1192 gnd.n1189 186.49
R5120 gnd.n1452 gnd.n1449 186.49
R5121 gnd.n3439 gnd.n3438 185
R5122 gnd.n3437 gnd.n3436 185
R5123 gnd.n3416 gnd.n3415 185
R5124 gnd.n3431 gnd.n3430 185
R5125 gnd.n3429 gnd.n3428 185
R5126 gnd.n3420 gnd.n3419 185
R5127 gnd.n3423 gnd.n3422 185
R5128 gnd.n3407 gnd.n3406 185
R5129 gnd.n3405 gnd.n3404 185
R5130 gnd.n3384 gnd.n3383 185
R5131 gnd.n3399 gnd.n3398 185
R5132 gnd.n3397 gnd.n3396 185
R5133 gnd.n3388 gnd.n3387 185
R5134 gnd.n3391 gnd.n3390 185
R5135 gnd.n3375 gnd.n3374 185
R5136 gnd.n3373 gnd.n3372 185
R5137 gnd.n3352 gnd.n3351 185
R5138 gnd.n3367 gnd.n3366 185
R5139 gnd.n3365 gnd.n3364 185
R5140 gnd.n3356 gnd.n3355 185
R5141 gnd.n3359 gnd.n3358 185
R5142 gnd.n3344 gnd.n3343 185
R5143 gnd.n3342 gnd.n3341 185
R5144 gnd.n3321 gnd.n3320 185
R5145 gnd.n3336 gnd.n3335 185
R5146 gnd.n3334 gnd.n3333 185
R5147 gnd.n3325 gnd.n3324 185
R5148 gnd.n3328 gnd.n3327 185
R5149 gnd.n3312 gnd.n3311 185
R5150 gnd.n3310 gnd.n3309 185
R5151 gnd.n3289 gnd.n3288 185
R5152 gnd.n3304 gnd.n3303 185
R5153 gnd.n3302 gnd.n3301 185
R5154 gnd.n3293 gnd.n3292 185
R5155 gnd.n3296 gnd.n3295 185
R5156 gnd.n3280 gnd.n3279 185
R5157 gnd.n3278 gnd.n3277 185
R5158 gnd.n3257 gnd.n3256 185
R5159 gnd.n3272 gnd.n3271 185
R5160 gnd.n3270 gnd.n3269 185
R5161 gnd.n3261 gnd.n3260 185
R5162 gnd.n3264 gnd.n3263 185
R5163 gnd.n3248 gnd.n3247 185
R5164 gnd.n3246 gnd.n3245 185
R5165 gnd.n3225 gnd.n3224 185
R5166 gnd.n3240 gnd.n3239 185
R5167 gnd.n3238 gnd.n3237 185
R5168 gnd.n3229 gnd.n3228 185
R5169 gnd.n3232 gnd.n3231 185
R5170 gnd.n3217 gnd.n3216 185
R5171 gnd.n3215 gnd.n3214 185
R5172 gnd.n3194 gnd.n3193 185
R5173 gnd.n3209 gnd.n3208 185
R5174 gnd.n3207 gnd.n3206 185
R5175 gnd.n3198 gnd.n3197 185
R5176 gnd.n3201 gnd.n3200 185
R5177 gnd.n2664 gnd.t176 178.987
R5178 gnd.n2186 gnd.t111 178.987
R5179 gnd.n1 gnd.t204 170.774
R5180 gnd.n7 gnd.t49 170.103
R5181 gnd.n6 gnd.t47 170.103
R5182 gnd.n5 gnd.t254 170.103
R5183 gnd.n4 gnd.t252 170.103
R5184 gnd.n3 gnd.t237 170.103
R5185 gnd.n2 gnd.t59 170.103
R5186 gnd.n1 gnd.t206 170.103
R5187 gnd.n5057 gnd.n5056 163.367
R5188 gnd.n5054 gnd.n1462 163.367
R5189 gnd.n5050 gnd.n5049 163.367
R5190 gnd.n5047 gnd.n1465 163.367
R5191 gnd.n5043 gnd.n5042 163.367
R5192 gnd.n5040 gnd.n1468 163.367
R5193 gnd.n5036 gnd.n5035 163.367
R5194 gnd.n5033 gnd.n1471 163.367
R5195 gnd.n5029 gnd.n5028 163.367
R5196 gnd.n5026 gnd.n1474 163.367
R5197 gnd.n5022 gnd.n5021 163.367
R5198 gnd.n5019 gnd.n1477 163.367
R5199 gnd.n5015 gnd.n5014 163.367
R5200 gnd.n5012 gnd.n1480 163.367
R5201 gnd.n5007 gnd.n5006 163.367
R5202 gnd.n5004 gnd.n5002 163.367
R5203 gnd.n4999 gnd.n4998 163.367
R5204 gnd.n4996 gnd.n1486 163.367
R5205 gnd.n4991 gnd.n4990 163.367
R5206 gnd.n4988 gnd.n1491 163.367
R5207 gnd.n4984 gnd.n4983 163.367
R5208 gnd.n4981 gnd.n1494 163.367
R5209 gnd.n4977 gnd.n4976 163.367
R5210 gnd.n4974 gnd.n1497 163.367
R5211 gnd.n4970 gnd.n4969 163.367
R5212 gnd.n4967 gnd.n1500 163.367
R5213 gnd.n4963 gnd.n4962 163.367
R5214 gnd.n4960 gnd.n1503 163.367
R5215 gnd.n4956 gnd.n4955 163.367
R5216 gnd.n4953 gnd.n1506 163.367
R5217 gnd.n4949 gnd.n4948 163.367
R5218 gnd.n4946 gnd.n1509 163.367
R5219 gnd.n1293 gnd.n1208 163.367
R5220 gnd.n1209 gnd.n1208 163.367
R5221 gnd.n1297 gnd.n1209 163.367
R5222 gnd.n1297 gnd.n1225 163.367
R5223 gnd.n5325 gnd.n1225 163.367
R5224 gnd.n5325 gnd.n1226 163.367
R5225 gnd.n5321 gnd.n1226 163.367
R5226 gnd.n5321 gnd.n1301 163.367
R5227 gnd.n1309 gnd.n1301 163.367
R5228 gnd.n4302 gnd.n1309 163.367
R5229 gnd.n4302 gnd.n4291 163.367
R5230 gnd.n4305 gnd.n4291 163.367
R5231 gnd.n4305 gnd.n4299 163.367
R5232 gnd.n4310 gnd.n4299 163.367
R5233 gnd.n4310 gnd.n4300 163.367
R5234 gnd.n4300 gnd.n1814 163.367
R5235 gnd.n4440 gnd.n1814 163.367
R5236 gnd.n4440 gnd.n1811 163.367
R5237 gnd.n4448 gnd.n1811 163.367
R5238 gnd.n4448 gnd.n1806 163.367
R5239 gnd.n4444 gnd.n1806 163.367
R5240 gnd.n4444 gnd.n1797 163.367
R5241 gnd.n1797 gnd.n1789 163.367
R5242 gnd.n4485 gnd.n1789 163.367
R5243 gnd.n4485 gnd.n1787 163.367
R5244 gnd.n4489 gnd.n1787 163.367
R5245 gnd.n4489 gnd.n1778 163.367
R5246 gnd.n4498 gnd.n1778 163.367
R5247 gnd.n4498 gnd.n1775 163.367
R5248 gnd.n4508 gnd.n1775 163.367
R5249 gnd.n4508 gnd.n1776 163.367
R5250 gnd.n1776 gnd.n1768 163.367
R5251 gnd.n4503 gnd.n1768 163.367
R5252 gnd.n4503 gnd.n1759 163.367
R5253 gnd.n1759 gnd.n1752 163.367
R5254 gnd.n4534 gnd.n1752 163.367
R5255 gnd.n4534 gnd.n1750 163.367
R5256 gnd.n4540 gnd.n1750 163.367
R5257 gnd.n4540 gnd.n1741 163.367
R5258 gnd.n1741 gnd.n1735 163.367
R5259 gnd.n4562 gnd.n1735 163.367
R5260 gnd.n4563 gnd.n4562 163.367
R5261 gnd.n4563 gnd.n1732 163.367
R5262 gnd.n4571 gnd.n1732 163.367
R5263 gnd.n4571 gnd.n1726 163.367
R5264 gnd.n4567 gnd.n1726 163.367
R5265 gnd.n4567 gnd.n1717 163.367
R5266 gnd.n1717 gnd.n1708 163.367
R5267 gnd.n4609 gnd.n1708 163.367
R5268 gnd.n4609 gnd.n1706 163.367
R5269 gnd.n4613 gnd.n1706 163.367
R5270 gnd.n4613 gnd.n1699 163.367
R5271 gnd.n4622 gnd.n1699 163.367
R5272 gnd.n4622 gnd.n1696 163.367
R5273 gnd.n4632 gnd.n1696 163.367
R5274 gnd.n4632 gnd.n1697 163.367
R5275 gnd.n1697 gnd.n1688 163.367
R5276 gnd.n4627 gnd.n1688 163.367
R5277 gnd.n4627 gnd.n1678 163.367
R5278 gnd.n1678 gnd.n1670 163.367
R5279 gnd.n4657 gnd.n1670 163.367
R5280 gnd.n4657 gnd.n1668 163.367
R5281 gnd.n4663 gnd.n1668 163.367
R5282 gnd.n4663 gnd.n1659 163.367
R5283 gnd.n1659 gnd.n1652 163.367
R5284 gnd.n4684 gnd.n1652 163.367
R5285 gnd.n4685 gnd.n4684 163.367
R5286 gnd.n4685 gnd.n1649 163.367
R5287 gnd.n4694 gnd.n1649 163.367
R5288 gnd.n4694 gnd.n1643 163.367
R5289 gnd.n4690 gnd.n1643 163.367
R5290 gnd.n4690 gnd.n1634 163.367
R5291 gnd.n1634 gnd.n1628 163.367
R5292 gnd.n4720 gnd.n1628 163.367
R5293 gnd.n4721 gnd.n4720 163.367
R5294 gnd.n4721 gnd.n1621 163.367
R5295 gnd.n4727 gnd.n1621 163.367
R5296 gnd.n4728 gnd.n4727 163.367
R5297 gnd.n4728 gnd.n1626 163.367
R5298 gnd.n4740 gnd.n1626 163.367
R5299 gnd.n4740 gnd.n1604 163.367
R5300 gnd.n4736 gnd.n1604 163.367
R5301 gnd.n4736 gnd.n1600 163.367
R5302 gnd.n4733 gnd.n1600 163.367
R5303 gnd.n4733 gnd.n1590 163.367
R5304 gnd.n1590 gnd.n1582 163.367
R5305 gnd.n4823 gnd.n1582 163.367
R5306 gnd.n4823 gnd.n1579 163.367
R5307 gnd.n4833 gnd.n1579 163.367
R5308 gnd.n4833 gnd.n1580 163.367
R5309 gnd.n1580 gnd.n1573 163.367
R5310 gnd.n4828 gnd.n1573 163.367
R5311 gnd.n4828 gnd.n1563 163.367
R5312 gnd.n1563 gnd.n1557 163.367
R5313 gnd.n4859 gnd.n1557 163.367
R5314 gnd.n4859 gnd.n1555 163.367
R5315 gnd.n4865 gnd.n1555 163.367
R5316 gnd.n4865 gnd.n1545 163.367
R5317 gnd.n1545 gnd.n1539 163.367
R5318 gnd.n4887 gnd.n1539 163.367
R5319 gnd.n4888 gnd.n4887 163.367
R5320 gnd.n4888 gnd.n1532 163.367
R5321 gnd.n4891 gnd.n1532 163.367
R5322 gnd.n4891 gnd.n1527 163.367
R5323 gnd.n4897 gnd.n1527 163.367
R5324 gnd.n4897 gnd.n1517 163.367
R5325 gnd.n1517 gnd.n1511 163.367
R5326 gnd.n4937 gnd.n1511 163.367
R5327 gnd.n4938 gnd.n4937 163.367
R5328 gnd.n4938 gnd.n1435 163.367
R5329 gnd.n1183 gnd.n1182 163.367
R5330 gnd.n5397 gnd.n1182 163.367
R5331 gnd.n5395 gnd.n5394 163.367
R5332 gnd.n5391 gnd.n5390 163.367
R5333 gnd.n5387 gnd.n5386 163.367
R5334 gnd.n5383 gnd.n5382 163.367
R5335 gnd.n5379 gnd.n5378 163.367
R5336 gnd.n5375 gnd.n5374 163.367
R5337 gnd.n5371 gnd.n5370 163.367
R5338 gnd.n5367 gnd.n5366 163.367
R5339 gnd.n5363 gnd.n5362 163.367
R5340 gnd.n5359 gnd.n5358 163.367
R5341 gnd.n5355 gnd.n5354 163.367
R5342 gnd.n5351 gnd.n5350 163.367
R5343 gnd.n5347 gnd.n5346 163.367
R5344 gnd.n5343 gnd.n5342 163.367
R5345 gnd.n5406 gnd.n1148 163.367
R5346 gnd.n1231 gnd.n1230 163.367
R5347 gnd.n1236 gnd.n1235 163.367
R5348 gnd.n1240 gnd.n1239 163.367
R5349 gnd.n1244 gnd.n1243 163.367
R5350 gnd.n1248 gnd.n1247 163.367
R5351 gnd.n1252 gnd.n1251 163.367
R5352 gnd.n1256 gnd.n1255 163.367
R5353 gnd.n1260 gnd.n1259 163.367
R5354 gnd.n1264 gnd.n1263 163.367
R5355 gnd.n1268 gnd.n1267 163.367
R5356 gnd.n1272 gnd.n1271 163.367
R5357 gnd.n1276 gnd.n1275 163.367
R5358 gnd.n1280 gnd.n1279 163.367
R5359 gnd.n1284 gnd.n1283 163.367
R5360 gnd.n1288 gnd.n1287 163.367
R5361 gnd.n5335 gnd.n1184 163.367
R5362 gnd.n5335 gnd.n1206 163.367
R5363 gnd.n4267 gnd.n1206 163.367
R5364 gnd.n4271 gnd.n4267 163.367
R5365 gnd.n4271 gnd.n1221 163.367
R5366 gnd.n1303 gnd.n1221 163.367
R5367 gnd.n5319 gnd.n1303 163.367
R5368 gnd.n5319 gnd.n1304 163.367
R5369 gnd.n5315 gnd.n1304 163.367
R5370 gnd.n5315 gnd.n1307 163.367
R5371 gnd.n4317 gnd.n1307 163.367
R5372 gnd.n4317 gnd.n4292 163.367
R5373 gnd.n4313 gnd.n4292 163.367
R5374 gnd.n4313 gnd.n4312 163.367
R5375 gnd.n4312 gnd.n4297 163.367
R5376 gnd.n4297 gnd.n4294 163.367
R5377 gnd.n4294 gnd.n1810 163.367
R5378 gnd.n4452 gnd.n1810 163.367
R5379 gnd.n4452 gnd.n1808 163.367
R5380 gnd.n4456 gnd.n1808 163.367
R5381 gnd.n4456 gnd.n1795 163.367
R5382 gnd.n4479 gnd.n1795 163.367
R5383 gnd.n4479 gnd.n1793 163.367
R5384 gnd.n4483 gnd.n1793 163.367
R5385 gnd.n4483 gnd.n1784 163.367
R5386 gnd.n4492 gnd.n1784 163.367
R5387 gnd.n4492 gnd.n1782 163.367
R5388 gnd.n4496 gnd.n1782 163.367
R5389 gnd.n4496 gnd.n1772 163.367
R5390 gnd.n4510 gnd.n1772 163.367
R5391 gnd.n4510 gnd.n1770 163.367
R5392 gnd.n4514 gnd.n1770 163.367
R5393 gnd.n4514 gnd.n1758 163.367
R5394 gnd.n4527 gnd.n1758 163.367
R5395 gnd.n4527 gnd.n1755 163.367
R5396 gnd.n4532 gnd.n1755 163.367
R5397 gnd.n4532 gnd.n1756 163.367
R5398 gnd.n1756 gnd.n1739 163.367
R5399 gnd.n4556 gnd.n1739 163.367
R5400 gnd.n4556 gnd.n1737 163.367
R5401 gnd.n4560 gnd.n1737 163.367
R5402 gnd.n4560 gnd.n1730 163.367
R5403 gnd.n4576 gnd.n1730 163.367
R5404 gnd.n4576 gnd.n1728 163.367
R5405 gnd.n4580 gnd.n1728 163.367
R5406 gnd.n4580 gnd.n1715 163.367
R5407 gnd.n4603 gnd.n1715 163.367
R5408 gnd.n4603 gnd.n1713 163.367
R5409 gnd.n4607 gnd.n1713 163.367
R5410 gnd.n4607 gnd.n1704 163.367
R5411 gnd.n4616 gnd.n1704 163.367
R5412 gnd.n4616 gnd.n1702 163.367
R5413 gnd.n4620 gnd.n1702 163.367
R5414 gnd.n4620 gnd.n1692 163.367
R5415 gnd.n4634 gnd.n1692 163.367
R5416 gnd.n4634 gnd.n1690 163.367
R5417 gnd.n4638 gnd.n1690 163.367
R5418 gnd.n4638 gnd.n1677 163.367
R5419 gnd.n4650 gnd.n1677 163.367
R5420 gnd.n4650 gnd.n1674 163.367
R5421 gnd.n4655 gnd.n1674 163.367
R5422 gnd.n4655 gnd.n1675 163.367
R5423 gnd.n1675 gnd.n1657 163.367
R5424 gnd.n4678 gnd.n1657 163.367
R5425 gnd.n4678 gnd.n1655 163.367
R5426 gnd.n4682 gnd.n1655 163.367
R5427 gnd.n4682 gnd.n1647 163.367
R5428 gnd.n4698 gnd.n1647 163.367
R5429 gnd.n4698 gnd.n1645 163.367
R5430 gnd.n4702 gnd.n1645 163.367
R5431 gnd.n4702 gnd.n1633 163.367
R5432 gnd.n4714 gnd.n1633 163.367
R5433 gnd.n4714 gnd.n1631 163.367
R5434 gnd.n4718 gnd.n1631 163.367
R5435 gnd.n4718 gnd.n1622 163.367
R5436 gnd.n4748 gnd.n1622 163.367
R5437 gnd.n4748 gnd.n1623 163.367
R5438 gnd.n4744 gnd.n1623 163.367
R5439 gnd.n4744 gnd.n4743 163.367
R5440 gnd.n4743 gnd.n1603 163.367
R5441 gnd.n4799 gnd.n1603 163.367
R5442 gnd.n4799 gnd.n1601 163.367
R5443 gnd.n4803 gnd.n1601 163.367
R5444 gnd.n4803 gnd.n1587 163.367
R5445 gnd.n4817 gnd.n1587 163.367
R5446 gnd.n4817 gnd.n1585 163.367
R5447 gnd.n4821 gnd.n1585 163.367
R5448 gnd.n4821 gnd.n1577 163.367
R5449 gnd.n4835 gnd.n1577 163.367
R5450 gnd.n4835 gnd.n1575 163.367
R5451 gnd.n4839 gnd.n1575 163.367
R5452 gnd.n4839 gnd.n1562 163.367
R5453 gnd.n4852 gnd.n1562 163.367
R5454 gnd.n4852 gnd.n1559 163.367
R5455 gnd.n4857 gnd.n1559 163.367
R5456 gnd.n4857 gnd.n1560 163.367
R5457 gnd.n1560 gnd.n1543 163.367
R5458 gnd.n4881 gnd.n1543 163.367
R5459 gnd.n4881 gnd.n1541 163.367
R5460 gnd.n4885 gnd.n1541 163.367
R5461 gnd.n4885 gnd.n1530 163.367
R5462 gnd.n4915 gnd.n1530 163.367
R5463 gnd.n4915 gnd.n1528 163.367
R5464 gnd.n4919 gnd.n1528 163.367
R5465 gnd.n4919 gnd.n1516 163.367
R5466 gnd.n4931 gnd.n1516 163.367
R5467 gnd.n4931 gnd.n1514 163.367
R5468 gnd.n4935 gnd.n1514 163.367
R5469 gnd.n4935 gnd.n1437 163.367
R5470 gnd.n5062 gnd.n1437 163.367
R5471 gnd.n1458 gnd.n1457 156.462
R5472 gnd.n3379 gnd.n3347 153.042
R5473 gnd.n3443 gnd.n3442 152.079
R5474 gnd.n3411 gnd.n3410 152.079
R5475 gnd.n3379 gnd.n3378 152.079
R5476 gnd.n1197 gnd.n1196 152
R5477 gnd.n1198 gnd.n1187 152
R5478 gnd.n1200 gnd.n1199 152
R5479 gnd.n1202 gnd.n1185 152
R5480 gnd.n1204 gnd.n1203 152
R5481 gnd.n1456 gnd.n1440 152
R5482 gnd.n1448 gnd.n1441 152
R5483 gnd.n1447 gnd.n1446 152
R5484 gnd.n1445 gnd.n1442 152
R5485 gnd.n1443 gnd.t155 150.546
R5486 gnd.t64 gnd.n3421 147.661
R5487 gnd.t276 gnd.n3389 147.661
R5488 gnd.t279 gnd.n3357 147.661
R5489 gnd.t202 gnd.n3326 147.661
R5490 gnd.t25 gnd.n3294 147.661
R5491 gnd.t23 gnd.n3262 147.661
R5492 gnd.t191 gnd.n3230 147.661
R5493 gnd.t288 gnd.n3199 147.661
R5494 gnd.n5001 gnd.n5000 143.351
R5495 gnd.n1164 gnd.n1147 143.351
R5496 gnd.n5405 gnd.n1147 143.351
R5497 gnd.n1194 gnd.t84 130.484
R5498 gnd.n1203 gnd.t149 126.766
R5499 gnd.n1201 gnd.t77 126.766
R5500 gnd.n1187 gnd.t105 126.766
R5501 gnd.n1195 gnd.t168 126.766
R5502 gnd.n1444 gnd.t142 126.766
R5503 gnd.n1446 gnd.t70 126.766
R5504 gnd.n1455 gnd.t126 126.766
R5505 gnd.n1457 gnd.t91 126.766
R5506 gnd.n5992 gnd.n5991 106.719
R5507 gnd.n5993 gnd.n5992 106.719
R5508 gnd.n5993 gnd.n629 106.719
R5509 gnd.n6001 gnd.n629 106.719
R5510 gnd.n6002 gnd.n6001 106.719
R5511 gnd.n6003 gnd.n6002 106.719
R5512 gnd.n6003 gnd.n623 106.719
R5513 gnd.n6011 gnd.n623 106.719
R5514 gnd.n6012 gnd.n6011 106.719
R5515 gnd.n6013 gnd.n6012 106.719
R5516 gnd.n6013 gnd.n617 106.719
R5517 gnd.n6021 gnd.n617 106.719
R5518 gnd.n6022 gnd.n6021 106.719
R5519 gnd.n6023 gnd.n6022 106.719
R5520 gnd.n6023 gnd.n611 106.719
R5521 gnd.n6031 gnd.n611 106.719
R5522 gnd.n6032 gnd.n6031 106.719
R5523 gnd.n6033 gnd.n6032 106.719
R5524 gnd.n6033 gnd.n605 106.719
R5525 gnd.n6041 gnd.n605 106.719
R5526 gnd.n6042 gnd.n6041 106.719
R5527 gnd.n6043 gnd.n6042 106.719
R5528 gnd.n6043 gnd.n599 106.719
R5529 gnd.n6051 gnd.n599 106.719
R5530 gnd.n6052 gnd.n6051 106.719
R5531 gnd.n6053 gnd.n6052 106.719
R5532 gnd.n6053 gnd.n593 106.719
R5533 gnd.n6061 gnd.n593 106.719
R5534 gnd.n6062 gnd.n6061 106.719
R5535 gnd.n6063 gnd.n6062 106.719
R5536 gnd.n6063 gnd.n587 106.719
R5537 gnd.n6071 gnd.n587 106.719
R5538 gnd.n6072 gnd.n6071 106.719
R5539 gnd.n6073 gnd.n6072 106.719
R5540 gnd.n6073 gnd.n581 106.719
R5541 gnd.n6081 gnd.n581 106.719
R5542 gnd.n6082 gnd.n6081 106.719
R5543 gnd.n6083 gnd.n6082 106.719
R5544 gnd.n6083 gnd.n575 106.719
R5545 gnd.n6091 gnd.n575 106.719
R5546 gnd.n6092 gnd.n6091 106.719
R5547 gnd.n6093 gnd.n6092 106.719
R5548 gnd.n6093 gnd.n569 106.719
R5549 gnd.n6101 gnd.n569 106.719
R5550 gnd.n6102 gnd.n6101 106.719
R5551 gnd.n6103 gnd.n6102 106.719
R5552 gnd.n6103 gnd.n563 106.719
R5553 gnd.n6111 gnd.n563 106.719
R5554 gnd.n6112 gnd.n6111 106.719
R5555 gnd.n6113 gnd.n6112 106.719
R5556 gnd.n6113 gnd.n557 106.719
R5557 gnd.n6121 gnd.n557 106.719
R5558 gnd.n6122 gnd.n6121 106.719
R5559 gnd.n6123 gnd.n6122 106.719
R5560 gnd.n6123 gnd.n551 106.719
R5561 gnd.n6131 gnd.n551 106.719
R5562 gnd.n6132 gnd.n6131 106.719
R5563 gnd.n6133 gnd.n6132 106.719
R5564 gnd.n6133 gnd.n545 106.719
R5565 gnd.n6141 gnd.n545 106.719
R5566 gnd.n6142 gnd.n6141 106.719
R5567 gnd.n6143 gnd.n6142 106.719
R5568 gnd.n6143 gnd.n539 106.719
R5569 gnd.n6151 gnd.n539 106.719
R5570 gnd.n6152 gnd.n6151 106.719
R5571 gnd.n6153 gnd.n6152 106.719
R5572 gnd.n6153 gnd.n533 106.719
R5573 gnd.n6161 gnd.n533 106.719
R5574 gnd.n6162 gnd.n6161 106.719
R5575 gnd.n6163 gnd.n6162 106.719
R5576 gnd.n6163 gnd.n527 106.719
R5577 gnd.n6171 gnd.n527 106.719
R5578 gnd.n6172 gnd.n6171 106.719
R5579 gnd.n6173 gnd.n6172 106.719
R5580 gnd.n6173 gnd.n521 106.719
R5581 gnd.n6181 gnd.n521 106.719
R5582 gnd.n6182 gnd.n6181 106.719
R5583 gnd.n6183 gnd.n6182 106.719
R5584 gnd.n6183 gnd.n515 106.719
R5585 gnd.n6191 gnd.n515 106.719
R5586 gnd.n6192 gnd.n6191 106.719
R5587 gnd.n6194 gnd.n6192 106.719
R5588 gnd.n6194 gnd.n6193 106.719
R5589 gnd.n3438 gnd.n3437 104.615
R5590 gnd.n3437 gnd.n3415 104.615
R5591 gnd.n3430 gnd.n3415 104.615
R5592 gnd.n3430 gnd.n3429 104.615
R5593 gnd.n3429 gnd.n3419 104.615
R5594 gnd.n3422 gnd.n3419 104.615
R5595 gnd.n3406 gnd.n3405 104.615
R5596 gnd.n3405 gnd.n3383 104.615
R5597 gnd.n3398 gnd.n3383 104.615
R5598 gnd.n3398 gnd.n3397 104.615
R5599 gnd.n3397 gnd.n3387 104.615
R5600 gnd.n3390 gnd.n3387 104.615
R5601 gnd.n3374 gnd.n3373 104.615
R5602 gnd.n3373 gnd.n3351 104.615
R5603 gnd.n3366 gnd.n3351 104.615
R5604 gnd.n3366 gnd.n3365 104.615
R5605 gnd.n3365 gnd.n3355 104.615
R5606 gnd.n3358 gnd.n3355 104.615
R5607 gnd.n3343 gnd.n3342 104.615
R5608 gnd.n3342 gnd.n3320 104.615
R5609 gnd.n3335 gnd.n3320 104.615
R5610 gnd.n3335 gnd.n3334 104.615
R5611 gnd.n3334 gnd.n3324 104.615
R5612 gnd.n3327 gnd.n3324 104.615
R5613 gnd.n3311 gnd.n3310 104.615
R5614 gnd.n3310 gnd.n3288 104.615
R5615 gnd.n3303 gnd.n3288 104.615
R5616 gnd.n3303 gnd.n3302 104.615
R5617 gnd.n3302 gnd.n3292 104.615
R5618 gnd.n3295 gnd.n3292 104.615
R5619 gnd.n3279 gnd.n3278 104.615
R5620 gnd.n3278 gnd.n3256 104.615
R5621 gnd.n3271 gnd.n3256 104.615
R5622 gnd.n3271 gnd.n3270 104.615
R5623 gnd.n3270 gnd.n3260 104.615
R5624 gnd.n3263 gnd.n3260 104.615
R5625 gnd.n3247 gnd.n3246 104.615
R5626 gnd.n3246 gnd.n3224 104.615
R5627 gnd.n3239 gnd.n3224 104.615
R5628 gnd.n3239 gnd.n3238 104.615
R5629 gnd.n3238 gnd.n3228 104.615
R5630 gnd.n3231 gnd.n3228 104.615
R5631 gnd.n3216 gnd.n3215 104.615
R5632 gnd.n3215 gnd.n3193 104.615
R5633 gnd.n3208 gnd.n3193 104.615
R5634 gnd.n3208 gnd.n3207 104.615
R5635 gnd.n3207 gnd.n3197 104.615
R5636 gnd.n3200 gnd.n3197 104.615
R5637 gnd.n2589 gnd.t83 100.632
R5638 gnd.n2159 gnd.t114 100.632
R5639 gnd.n6756 gnd.n93 99.6594
R5640 gnd.n6754 gnd.n6753 99.6594
R5641 gnd.n6749 gnd.n100 99.6594
R5642 gnd.n6747 gnd.n6746 99.6594
R5643 gnd.n6742 gnd.n107 99.6594
R5644 gnd.n6740 gnd.n6739 99.6594
R5645 gnd.n6735 gnd.n114 99.6594
R5646 gnd.n6733 gnd.n6732 99.6594
R5647 gnd.n6725 gnd.n121 99.6594
R5648 gnd.n6723 gnd.n6722 99.6594
R5649 gnd.n6718 gnd.n128 99.6594
R5650 gnd.n6716 gnd.n6715 99.6594
R5651 gnd.n6711 gnd.n135 99.6594
R5652 gnd.n6709 gnd.n6708 99.6594
R5653 gnd.n6704 gnd.n142 99.6594
R5654 gnd.n6702 gnd.n6701 99.6594
R5655 gnd.n6697 gnd.n149 99.6594
R5656 gnd.n6695 gnd.n6694 99.6594
R5657 gnd.n154 gnd.n153 99.6594
R5658 gnd.n6389 gnd.n327 99.6594
R5659 gnd.n6384 gnd.n385 99.6594
R5660 gnd.n6381 gnd.n386 99.6594
R5661 gnd.n6377 gnd.n387 99.6594
R5662 gnd.n6373 gnd.n388 99.6594
R5663 gnd.n6369 gnd.n389 99.6594
R5664 gnd.n6365 gnd.n390 99.6594
R5665 gnd.n6361 gnd.n391 99.6594
R5666 gnd.n6356 gnd.n393 99.6594
R5667 gnd.n6352 gnd.n394 99.6594
R5668 gnd.n6348 gnd.n395 99.6594
R5669 gnd.n6344 gnd.n396 99.6594
R5670 gnd.n6340 gnd.n397 99.6594
R5671 gnd.n6336 gnd.n398 99.6594
R5672 gnd.n6332 gnd.n399 99.6594
R5673 gnd.n6328 gnd.n400 99.6594
R5674 gnd.n6324 gnd.n401 99.6594
R5675 gnd.n459 gnd.n402 99.6594
R5676 gnd.n5436 gnd.n5435 99.6594
R5677 gnd.n5431 gnd.n1124 99.6594
R5678 gnd.n5427 gnd.n1123 99.6594
R5679 gnd.n5423 gnd.n1122 99.6594
R5680 gnd.n5419 gnd.n1121 99.6594
R5681 gnd.n5415 gnd.n1120 99.6594
R5682 gnd.n5411 gnd.n1119 99.6594
R5683 gnd.n4092 gnd.n1117 99.6594
R5684 gnd.n4099 gnd.n1116 99.6594
R5685 gnd.n4103 gnd.n1115 99.6594
R5686 gnd.n4109 gnd.n1114 99.6594
R5687 gnd.n4113 gnd.n1113 99.6594
R5688 gnd.n4119 gnd.n1112 99.6594
R5689 gnd.n4123 gnd.n1111 99.6594
R5690 gnd.n4129 gnd.n1110 99.6594
R5691 gnd.n4133 gnd.n1109 99.6594
R5692 gnd.n4138 gnd.n1108 99.6594
R5693 gnd.n4141 gnd.n1107 99.6594
R5694 gnd.n3877 gnd.n3876 99.6594
R5695 gnd.n3871 gnd.n3571 99.6594
R5696 gnd.n3868 gnd.n3572 99.6594
R5697 gnd.n3864 gnd.n3573 99.6594
R5698 gnd.n3860 gnd.n3574 99.6594
R5699 gnd.n3856 gnd.n3575 99.6594
R5700 gnd.n3852 gnd.n3576 99.6594
R5701 gnd.n3848 gnd.n3577 99.6594
R5702 gnd.n3844 gnd.n3578 99.6594
R5703 gnd.n3839 gnd.n3579 99.6594
R5704 gnd.n3835 gnd.n3580 99.6594
R5705 gnd.n3831 gnd.n3581 99.6594
R5706 gnd.n3827 gnd.n3582 99.6594
R5707 gnd.n3823 gnd.n3583 99.6594
R5708 gnd.n3819 gnd.n3584 99.6594
R5709 gnd.n3815 gnd.n3585 99.6594
R5710 gnd.n3811 gnd.n3586 99.6594
R5711 gnd.n3807 gnd.n3587 99.6594
R5712 gnd.n3748 gnd.n3588 99.6594
R5713 gnd.n3561 gnd.n2142 99.6594
R5714 gnd.n3559 gnd.n2141 99.6594
R5715 gnd.n3555 gnd.n2140 99.6594
R5716 gnd.n3551 gnd.n2139 99.6594
R5717 gnd.n3547 gnd.n2138 99.6594
R5718 gnd.n3543 gnd.n2137 99.6594
R5719 gnd.n3539 gnd.n2136 99.6594
R5720 gnd.n3471 gnd.n2135 99.6594
R5721 gnd.n2801 gnd.n2532 99.6594
R5722 gnd.n2558 gnd.n2539 99.6594
R5723 gnd.n2560 gnd.n2540 99.6594
R5724 gnd.n2568 gnd.n2541 99.6594
R5725 gnd.n2570 gnd.n2542 99.6594
R5726 gnd.n2578 gnd.n2543 99.6594
R5727 gnd.n2580 gnd.n2544 99.6594
R5728 gnd.n2588 gnd.n2545 99.6594
R5729 gnd.n3529 gnd.n2122 99.6594
R5730 gnd.n3525 gnd.n2123 99.6594
R5731 gnd.n3521 gnd.n2124 99.6594
R5732 gnd.n3517 gnd.n2125 99.6594
R5733 gnd.n3513 gnd.n2126 99.6594
R5734 gnd.n3509 gnd.n2127 99.6594
R5735 gnd.n3505 gnd.n2128 99.6594
R5736 gnd.n3501 gnd.n2129 99.6594
R5737 gnd.n3497 gnd.n2130 99.6594
R5738 gnd.n3493 gnd.n2131 99.6594
R5739 gnd.n3489 gnd.n2132 99.6594
R5740 gnd.n3485 gnd.n2133 99.6594
R5741 gnd.n3481 gnd.n2134 99.6594
R5742 gnd.n2716 gnd.n2715 99.6594
R5743 gnd.n2710 gnd.n2627 99.6594
R5744 gnd.n2707 gnd.n2628 99.6594
R5745 gnd.n2703 gnd.n2629 99.6594
R5746 gnd.n2699 gnd.n2630 99.6594
R5747 gnd.n2695 gnd.n2631 99.6594
R5748 gnd.n2691 gnd.n2632 99.6594
R5749 gnd.n2687 gnd.n2633 99.6594
R5750 gnd.n2683 gnd.n2634 99.6594
R5751 gnd.n2679 gnd.n2635 99.6594
R5752 gnd.n2675 gnd.n2636 99.6594
R5753 gnd.n2671 gnd.n2637 99.6594
R5754 gnd.n2718 gnd.n2626 99.6594
R5755 gnd.n6605 gnd.n6604 99.6594
R5756 gnd.n6610 gnd.n6609 99.6594
R5757 gnd.n6613 gnd.n6612 99.6594
R5758 gnd.n6618 gnd.n6617 99.6594
R5759 gnd.n6621 gnd.n6620 99.6594
R5760 gnd.n6626 gnd.n6625 99.6594
R5761 gnd.n6629 gnd.n6628 99.6594
R5762 gnd.n6634 gnd.n6633 99.6594
R5763 gnd.n6637 gnd.n80 99.6594
R5764 gnd.n403 gnd.n332 99.6594
R5765 gnd.n405 gnd.n404 99.6594
R5766 gnd.n407 gnd.n342 99.6594
R5767 gnd.n408 gnd.n349 99.6594
R5768 gnd.n410 gnd.n409 99.6594
R5769 gnd.n412 gnd.n358 99.6594
R5770 gnd.n413 gnd.n365 99.6594
R5771 gnd.n415 gnd.n414 99.6594
R5772 gnd.n416 gnd.n374 99.6594
R5773 gnd.n1915 gnd.n1097 99.6594
R5774 gnd.n1926 gnd.n1098 99.6594
R5775 gnd.n1897 gnd.n1099 99.6594
R5776 gnd.n1939 gnd.n1100 99.6594
R5777 gnd.n1950 gnd.n1101 99.6594
R5778 gnd.n1885 gnd.n1102 99.6594
R5779 gnd.n1963 gnd.n1103 99.6594
R5780 gnd.n1977 gnd.n1104 99.6594
R5781 gnd.n4188 gnd.n1105 99.6594
R5782 gnd.n3880 gnd.n3879 99.6594
R5783 gnd.n3610 gnd.n3589 99.6594
R5784 gnd.n3614 gnd.n3590 99.6594
R5785 gnd.n3620 gnd.n3591 99.6594
R5786 gnd.n3624 gnd.n3592 99.6594
R5787 gnd.n3630 gnd.n3593 99.6594
R5788 gnd.n3634 gnd.n3594 99.6594
R5789 gnd.n3640 gnd.n3595 99.6594
R5790 gnd.n3644 gnd.n3596 99.6594
R5791 gnd.n3879 gnd.n2119 99.6594
R5792 gnd.n3613 gnd.n3589 99.6594
R5793 gnd.n3619 gnd.n3590 99.6594
R5794 gnd.n3623 gnd.n3591 99.6594
R5795 gnd.n3629 gnd.n3592 99.6594
R5796 gnd.n3633 gnd.n3593 99.6594
R5797 gnd.n3639 gnd.n3594 99.6594
R5798 gnd.n3643 gnd.n3595 99.6594
R5799 gnd.n3597 gnd.n3596 99.6594
R5800 gnd.n1978 gnd.n1105 99.6594
R5801 gnd.n1962 gnd.n1104 99.6594
R5802 gnd.n1886 gnd.n1103 99.6594
R5803 gnd.n1951 gnd.n1102 99.6594
R5804 gnd.n1938 gnd.n1101 99.6594
R5805 gnd.n1898 gnd.n1100 99.6594
R5806 gnd.n1927 gnd.n1099 99.6594
R5807 gnd.n1914 gnd.n1098 99.6594
R5808 gnd.n1911 gnd.n1097 99.6594
R5809 gnd.n403 gnd.n334 99.6594
R5810 gnd.n405 gnd.n341 99.6594
R5811 gnd.n407 gnd.n406 99.6594
R5812 gnd.n408 gnd.n350 99.6594
R5813 gnd.n410 gnd.n357 99.6594
R5814 gnd.n412 gnd.n411 99.6594
R5815 gnd.n413 gnd.n366 99.6594
R5816 gnd.n415 gnd.n373 99.6594
R5817 gnd.n416 gnd.n383 99.6594
R5818 gnd.n6638 gnd.n6637 99.6594
R5819 gnd.n6633 gnd.n6632 99.6594
R5820 gnd.n6628 gnd.n6627 99.6594
R5821 gnd.n6625 gnd.n6624 99.6594
R5822 gnd.n6620 gnd.n6619 99.6594
R5823 gnd.n6617 gnd.n6616 99.6594
R5824 gnd.n6612 gnd.n6611 99.6594
R5825 gnd.n6609 gnd.n6608 99.6594
R5826 gnd.n6604 gnd.n6603 99.6594
R5827 gnd.n2716 gnd.n2639 99.6594
R5828 gnd.n2708 gnd.n2627 99.6594
R5829 gnd.n2704 gnd.n2628 99.6594
R5830 gnd.n2700 gnd.n2629 99.6594
R5831 gnd.n2696 gnd.n2630 99.6594
R5832 gnd.n2692 gnd.n2631 99.6594
R5833 gnd.n2688 gnd.n2632 99.6594
R5834 gnd.n2684 gnd.n2633 99.6594
R5835 gnd.n2680 gnd.n2634 99.6594
R5836 gnd.n2676 gnd.n2635 99.6594
R5837 gnd.n2672 gnd.n2636 99.6594
R5838 gnd.n2668 gnd.n2637 99.6594
R5839 gnd.n2719 gnd.n2718 99.6594
R5840 gnd.n3484 gnd.n2134 99.6594
R5841 gnd.n3488 gnd.n2133 99.6594
R5842 gnd.n3492 gnd.n2132 99.6594
R5843 gnd.n3496 gnd.n2131 99.6594
R5844 gnd.n3500 gnd.n2130 99.6594
R5845 gnd.n3504 gnd.n2129 99.6594
R5846 gnd.n3508 gnd.n2128 99.6594
R5847 gnd.n3512 gnd.n2127 99.6594
R5848 gnd.n3516 gnd.n2126 99.6594
R5849 gnd.n3520 gnd.n2125 99.6594
R5850 gnd.n3524 gnd.n2124 99.6594
R5851 gnd.n3528 gnd.n2123 99.6594
R5852 gnd.n2163 gnd.n2122 99.6594
R5853 gnd.n2802 gnd.n2801 99.6594
R5854 gnd.n2561 gnd.n2539 99.6594
R5855 gnd.n2567 gnd.n2540 99.6594
R5856 gnd.n2571 gnd.n2541 99.6594
R5857 gnd.n2577 gnd.n2542 99.6594
R5858 gnd.n2581 gnd.n2543 99.6594
R5859 gnd.n2587 gnd.n2544 99.6594
R5860 gnd.n2545 gnd.n2529 99.6594
R5861 gnd.n3538 gnd.n2135 99.6594
R5862 gnd.n3542 gnd.n2136 99.6594
R5863 gnd.n3546 gnd.n2137 99.6594
R5864 gnd.n3550 gnd.n2138 99.6594
R5865 gnd.n3554 gnd.n2139 99.6594
R5866 gnd.n3558 gnd.n2140 99.6594
R5867 gnd.n3562 gnd.n2141 99.6594
R5868 gnd.n2144 gnd.n2142 99.6594
R5869 gnd.n3877 gnd.n3708 99.6594
R5870 gnd.n3869 gnd.n3571 99.6594
R5871 gnd.n3865 gnd.n3572 99.6594
R5872 gnd.n3861 gnd.n3573 99.6594
R5873 gnd.n3857 gnd.n3574 99.6594
R5874 gnd.n3853 gnd.n3575 99.6594
R5875 gnd.n3849 gnd.n3576 99.6594
R5876 gnd.n3845 gnd.n3577 99.6594
R5877 gnd.n3840 gnd.n3578 99.6594
R5878 gnd.n3836 gnd.n3579 99.6594
R5879 gnd.n3832 gnd.n3580 99.6594
R5880 gnd.n3828 gnd.n3581 99.6594
R5881 gnd.n3824 gnd.n3582 99.6594
R5882 gnd.n3820 gnd.n3583 99.6594
R5883 gnd.n3816 gnd.n3584 99.6594
R5884 gnd.n3812 gnd.n3585 99.6594
R5885 gnd.n3808 gnd.n3586 99.6594
R5886 gnd.n3747 gnd.n3587 99.6594
R5887 gnd.n3800 gnd.n3588 99.6594
R5888 gnd.n4083 gnd.n1107 99.6594
R5889 gnd.n4132 gnd.n1108 99.6594
R5890 gnd.n4130 gnd.n1109 99.6594
R5891 gnd.n4122 gnd.n1110 99.6594
R5892 gnd.n4120 gnd.n1111 99.6594
R5893 gnd.n4112 gnd.n1112 99.6594
R5894 gnd.n4110 gnd.n1113 99.6594
R5895 gnd.n4102 gnd.n1114 99.6594
R5896 gnd.n4100 gnd.n1115 99.6594
R5897 gnd.n4093 gnd.n1116 99.6594
R5898 gnd.n5410 gnd.n1118 99.6594
R5899 gnd.n5414 gnd.n1119 99.6594
R5900 gnd.n5418 gnd.n1120 99.6594
R5901 gnd.n5422 gnd.n1121 99.6594
R5902 gnd.n5426 gnd.n1122 99.6594
R5903 gnd.n5430 gnd.n1123 99.6594
R5904 gnd.n1125 gnd.n1124 99.6594
R5905 gnd.n5436 gnd.n1094 99.6594
R5906 gnd.n6389 gnd.n6388 99.6594
R5907 gnd.n6382 gnd.n385 99.6594
R5908 gnd.n6378 gnd.n386 99.6594
R5909 gnd.n6374 gnd.n387 99.6594
R5910 gnd.n6370 gnd.n388 99.6594
R5911 gnd.n6366 gnd.n389 99.6594
R5912 gnd.n6362 gnd.n390 99.6594
R5913 gnd.n6357 gnd.n392 99.6594
R5914 gnd.n6353 gnd.n393 99.6594
R5915 gnd.n6349 gnd.n394 99.6594
R5916 gnd.n6345 gnd.n395 99.6594
R5917 gnd.n6341 gnd.n396 99.6594
R5918 gnd.n6337 gnd.n397 99.6594
R5919 gnd.n6333 gnd.n398 99.6594
R5920 gnd.n6329 gnd.n399 99.6594
R5921 gnd.n6325 gnd.n400 99.6594
R5922 gnd.n458 gnd.n401 99.6594
R5923 gnd.n6317 gnd.n402 99.6594
R5924 gnd.n153 gnd.n150 99.6594
R5925 gnd.n6696 gnd.n6695 99.6594
R5926 gnd.n149 gnd.n143 99.6594
R5927 gnd.n6703 gnd.n6702 99.6594
R5928 gnd.n142 gnd.n136 99.6594
R5929 gnd.n6710 gnd.n6709 99.6594
R5930 gnd.n135 gnd.n129 99.6594
R5931 gnd.n6717 gnd.n6716 99.6594
R5932 gnd.n128 gnd.n122 99.6594
R5933 gnd.n6724 gnd.n6723 99.6594
R5934 gnd.n121 gnd.n115 99.6594
R5935 gnd.n6734 gnd.n6733 99.6594
R5936 gnd.n114 gnd.n108 99.6594
R5937 gnd.n6741 gnd.n6740 99.6594
R5938 gnd.n107 gnd.n101 99.6594
R5939 gnd.n6748 gnd.n6747 99.6594
R5940 gnd.n100 gnd.n94 99.6594
R5941 gnd.n6755 gnd.n6754 99.6594
R5942 gnd.n93 gnd.n90 99.6594
R5943 gnd.n1848 gnd.n1837 99.6594
R5944 gnd.n1921 gnd.n1849 99.6594
R5945 gnd.n1902 gnd.n1850 99.6594
R5946 gnd.n1932 gnd.n1851 99.6594
R5947 gnd.n1945 gnd.n1852 99.6594
R5948 gnd.n1890 gnd.n1853 99.6594
R5949 gnd.n1956 gnd.n1854 99.6594
R5950 gnd.n1969 gnd.n1855 99.6594
R5951 gnd.n1878 gnd.n1856 99.6594
R5952 gnd.n4195 gnd.n1857 99.6594
R5953 gnd.n1873 gnd.n1858 99.6594
R5954 gnd.n4204 gnd.n1859 99.6594
R5955 gnd.n1869 gnd.n1860 99.6594
R5956 gnd.n4213 gnd.n1861 99.6594
R5957 gnd.n1920 gnd.n1848 99.6594
R5958 gnd.n1901 gnd.n1849 99.6594
R5959 gnd.n1933 gnd.n1850 99.6594
R5960 gnd.n1944 gnd.n1851 99.6594
R5961 gnd.n1889 gnd.n1852 99.6594
R5962 gnd.n1957 gnd.n1853 99.6594
R5963 gnd.n1968 gnd.n1854 99.6594
R5964 gnd.n1877 gnd.n1855 99.6594
R5965 gnd.n4194 gnd.n1856 99.6594
R5966 gnd.n1872 gnd.n1857 99.6594
R5967 gnd.n4203 gnd.n1858 99.6594
R5968 gnd.n1868 gnd.n1859 99.6594
R5969 gnd.n4212 gnd.n1860 99.6594
R5970 gnd.n1862 gnd.n1861 99.6594
R5971 gnd.n5075 gnd.n337 99.6594
R5972 gnd.n5077 gnd.n5076 99.6594
R5973 gnd.n5079 gnd.n346 99.6594
R5974 gnd.n5080 gnd.n353 99.6594
R5975 gnd.n5082 gnd.n5081 99.6594
R5976 gnd.n5084 gnd.n362 99.6594
R5977 gnd.n5085 gnd.n369 99.6594
R5978 gnd.n5087 gnd.n5086 99.6594
R5979 gnd.n5088 gnd.n380 99.6594
R5980 gnd.n5102 gnd.n5089 99.6594
R5981 gnd.n5159 gnd.n5090 99.6594
R5982 gnd.n5161 gnd.n5091 99.6594
R5983 gnd.n5169 gnd.n5092 99.6594
R5984 gnd.n5179 gnd.n5093 99.6594
R5985 gnd.n5179 gnd.n5178 99.6594
R5986 gnd.n5172 gnd.n5092 99.6594
R5987 gnd.n5168 gnd.n5091 99.6594
R5988 gnd.n5162 gnd.n5090 99.6594
R5989 gnd.n5158 gnd.n5089 99.6594
R5990 gnd.n5101 gnd.n5088 99.6594
R5991 gnd.n5087 gnd.n379 99.6594
R5992 gnd.n5085 gnd.n370 99.6594
R5993 gnd.n5084 gnd.n5083 99.6594
R5994 gnd.n5082 gnd.n361 99.6594
R5995 gnd.n5080 gnd.n354 99.6594
R5996 gnd.n5079 gnd.n5078 99.6594
R5997 gnd.n5077 gnd.n345 99.6594
R5998 gnd.n5075 gnd.n338 99.6594
R5999 gnd.n1865 gnd.t148 98.63
R6000 gnd.n6635 gnd.t134 98.63
R6001 gnd.n375 gnd.t125 98.63
R6002 gnd.n1975 gnd.t140 98.63
R6003 gnd.n438 gnd.t122 98.63
R6004 gnd.n460 gnd.t90 98.63
R6005 gnd.n156 gnd.t75 98.63
R6006 gnd.n6727 gnd.t103 98.63
R6007 gnd.n3727 gnd.t173 98.63
R6008 gnd.n3749 gnd.t164 98.63
R6009 gnd.n3599 gnd.t161 98.63
R6010 gnd.n4081 gnd.t96 98.63
R6011 gnd.n1141 gnd.t137 98.63
R6012 gnd.n5097 gnd.t131 98.63
R6013 gnd.n1227 gnd.t167 96.6984
R6014 gnd.n1487 gnd.t100 96.6984
R6015 gnd.n5339 gnd.t119 96.6906
R6016 gnd.n1481 gnd.t153 96.6906
R6017 gnd.n1194 gnd.n1193 81.8399
R6018 gnd.n2590 gnd.t82 74.8376
R6019 gnd.n2160 gnd.t115 74.8376
R6020 gnd.n1228 gnd.t166 72.8438
R6021 gnd.n1488 gnd.t101 72.8438
R6022 gnd.n1195 gnd.n1188 72.8411
R6023 gnd.n1201 gnd.n1186 72.8411
R6024 gnd.n1455 gnd.n1454 72.8411
R6025 gnd.n1866 gnd.t147 72.836
R6026 gnd.n5340 gnd.t118 72.836
R6027 gnd.n1482 gnd.t154 72.836
R6028 gnd.n6636 gnd.t135 72.836
R6029 gnd.n376 gnd.t124 72.836
R6030 gnd.n1976 gnd.t141 72.836
R6031 gnd.n439 gnd.t121 72.836
R6032 gnd.n461 gnd.t89 72.836
R6033 gnd.n157 gnd.t76 72.836
R6034 gnd.n6728 gnd.t104 72.836
R6035 gnd.n3728 gnd.t172 72.836
R6036 gnd.n3750 gnd.t163 72.836
R6037 gnd.n3600 gnd.t160 72.836
R6038 gnd.n4082 gnd.t97 72.836
R6039 gnd.n1142 gnd.t138 72.836
R6040 gnd.n5098 gnd.t132 72.836
R6041 gnd.n5057 gnd.n1460 71.676
R6042 gnd.n5055 gnd.n5054 71.676
R6043 gnd.n5050 gnd.n1464 71.676
R6044 gnd.n5048 gnd.n5047 71.676
R6045 gnd.n5043 gnd.n1467 71.676
R6046 gnd.n5041 gnd.n5040 71.676
R6047 gnd.n5036 gnd.n1470 71.676
R6048 gnd.n5034 gnd.n5033 71.676
R6049 gnd.n5029 gnd.n1473 71.676
R6050 gnd.n5027 gnd.n5026 71.676
R6051 gnd.n5022 gnd.n1476 71.676
R6052 gnd.n5020 gnd.n5019 71.676
R6053 gnd.n5015 gnd.n1479 71.676
R6054 gnd.n5013 gnd.n5012 71.676
R6055 gnd.n5007 gnd.n1484 71.676
R6056 gnd.n5005 gnd.n5004 71.676
R6057 gnd.n5000 gnd.n4999 71.676
R6058 gnd.n4997 gnd.n4996 71.676
R6059 gnd.n4991 gnd.n1490 71.676
R6060 gnd.n4989 gnd.n4988 71.676
R6061 gnd.n4984 gnd.n1493 71.676
R6062 gnd.n4982 gnd.n4981 71.676
R6063 gnd.n4977 gnd.n1496 71.676
R6064 gnd.n4975 gnd.n4974 71.676
R6065 gnd.n4970 gnd.n1499 71.676
R6066 gnd.n4968 gnd.n4967 71.676
R6067 gnd.n4963 gnd.n1502 71.676
R6068 gnd.n4961 gnd.n4960 71.676
R6069 gnd.n4956 gnd.n1505 71.676
R6070 gnd.n4954 gnd.n4953 71.676
R6071 gnd.n4949 gnd.n1508 71.676
R6072 gnd.n4947 gnd.n4946 71.676
R6073 gnd.n4942 gnd.n4941 71.676
R6074 gnd.n5403 gnd.n5402 71.676
R6075 gnd.n5397 gnd.n1150 71.676
R6076 gnd.n5394 gnd.n1151 71.676
R6077 gnd.n5390 gnd.n1152 71.676
R6078 gnd.n5386 gnd.n1153 71.676
R6079 gnd.n5382 gnd.n1154 71.676
R6080 gnd.n5378 gnd.n1155 71.676
R6081 gnd.n5374 gnd.n1156 71.676
R6082 gnd.n5370 gnd.n1157 71.676
R6083 gnd.n5366 gnd.n1158 71.676
R6084 gnd.n5362 gnd.n1159 71.676
R6085 gnd.n5358 gnd.n1160 71.676
R6086 gnd.n5354 gnd.n1161 71.676
R6087 gnd.n5350 gnd.n1162 71.676
R6088 gnd.n5346 gnd.n1163 71.676
R6089 gnd.n5342 gnd.n1164 71.676
R6090 gnd.n1165 gnd.n1148 71.676
R6091 gnd.n1231 gnd.n1166 71.676
R6092 gnd.n1236 gnd.n1167 71.676
R6093 gnd.n1240 gnd.n1168 71.676
R6094 gnd.n1244 gnd.n1169 71.676
R6095 gnd.n1248 gnd.n1170 71.676
R6096 gnd.n1252 gnd.n1171 71.676
R6097 gnd.n1256 gnd.n1172 71.676
R6098 gnd.n1260 gnd.n1173 71.676
R6099 gnd.n1264 gnd.n1174 71.676
R6100 gnd.n1268 gnd.n1175 71.676
R6101 gnd.n1272 gnd.n1176 71.676
R6102 gnd.n1276 gnd.n1177 71.676
R6103 gnd.n1280 gnd.n1178 71.676
R6104 gnd.n1284 gnd.n1179 71.676
R6105 gnd.n1288 gnd.n1180 71.676
R6106 gnd.n5403 gnd.n1183 71.676
R6107 gnd.n5395 gnd.n1150 71.676
R6108 gnd.n5391 gnd.n1151 71.676
R6109 gnd.n5387 gnd.n1152 71.676
R6110 gnd.n5383 gnd.n1153 71.676
R6111 gnd.n5379 gnd.n1154 71.676
R6112 gnd.n5375 gnd.n1155 71.676
R6113 gnd.n5371 gnd.n1156 71.676
R6114 gnd.n5367 gnd.n1157 71.676
R6115 gnd.n5363 gnd.n1158 71.676
R6116 gnd.n5359 gnd.n1159 71.676
R6117 gnd.n5355 gnd.n1160 71.676
R6118 gnd.n5351 gnd.n1161 71.676
R6119 gnd.n5347 gnd.n1162 71.676
R6120 gnd.n5343 gnd.n1163 71.676
R6121 gnd.n5406 gnd.n5405 71.676
R6122 gnd.n1230 gnd.n1165 71.676
R6123 gnd.n1235 gnd.n1166 71.676
R6124 gnd.n1239 gnd.n1167 71.676
R6125 gnd.n1243 gnd.n1168 71.676
R6126 gnd.n1247 gnd.n1169 71.676
R6127 gnd.n1251 gnd.n1170 71.676
R6128 gnd.n1255 gnd.n1171 71.676
R6129 gnd.n1259 gnd.n1172 71.676
R6130 gnd.n1263 gnd.n1173 71.676
R6131 gnd.n1267 gnd.n1174 71.676
R6132 gnd.n1271 gnd.n1175 71.676
R6133 gnd.n1275 gnd.n1176 71.676
R6134 gnd.n1279 gnd.n1177 71.676
R6135 gnd.n1283 gnd.n1178 71.676
R6136 gnd.n1287 gnd.n1179 71.676
R6137 gnd.n1291 gnd.n1180 71.676
R6138 gnd.n4941 gnd.n1509 71.676
R6139 gnd.n4948 gnd.n4947 71.676
R6140 gnd.n1508 gnd.n1506 71.676
R6141 gnd.n4955 gnd.n4954 71.676
R6142 gnd.n1505 gnd.n1503 71.676
R6143 gnd.n4962 gnd.n4961 71.676
R6144 gnd.n1502 gnd.n1500 71.676
R6145 gnd.n4969 gnd.n4968 71.676
R6146 gnd.n1499 gnd.n1497 71.676
R6147 gnd.n4976 gnd.n4975 71.676
R6148 gnd.n1496 gnd.n1494 71.676
R6149 gnd.n4983 gnd.n4982 71.676
R6150 gnd.n1493 gnd.n1491 71.676
R6151 gnd.n4990 gnd.n4989 71.676
R6152 gnd.n1490 gnd.n1486 71.676
R6153 gnd.n4998 gnd.n4997 71.676
R6154 gnd.n5002 gnd.n5001 71.676
R6155 gnd.n5006 gnd.n5005 71.676
R6156 gnd.n1484 gnd.n1480 71.676
R6157 gnd.n5014 gnd.n5013 71.676
R6158 gnd.n1479 gnd.n1477 71.676
R6159 gnd.n5021 gnd.n5020 71.676
R6160 gnd.n1476 gnd.n1474 71.676
R6161 gnd.n5028 gnd.n5027 71.676
R6162 gnd.n1473 gnd.n1471 71.676
R6163 gnd.n5035 gnd.n5034 71.676
R6164 gnd.n1470 gnd.n1468 71.676
R6165 gnd.n5042 gnd.n5041 71.676
R6166 gnd.n1467 gnd.n1465 71.676
R6167 gnd.n5049 gnd.n5048 71.676
R6168 gnd.n1464 gnd.n1462 71.676
R6169 gnd.n5056 gnd.n5055 71.676
R6170 gnd.n1460 gnd.n1438 71.676
R6171 gnd.n8 gnd.t241 69.1507
R6172 gnd.n14 gnd.t281 68.4792
R6173 gnd.n13 gnd.t256 68.4792
R6174 gnd.n12 gnd.t2 68.4792
R6175 gnd.n11 gnd.t230 68.4792
R6176 gnd.n10 gnd.t216 68.4792
R6177 gnd.n9 gnd.t57 68.4792
R6178 gnd.n8 gnd.t27 68.4792
R6179 gnd.n2717 gnd.n2621 64.369
R6180 gnd.n6193 gnd.n179 64.0315
R6181 gnd.n3878 gnd.n2112 63.0944
R6182 gnd.n6764 gnd.n83 63.0944
R6183 gnd.n1233 gnd.n1228 59.5399
R6184 gnd.n4993 gnd.n1488 59.5399
R6185 gnd.n5341 gnd.n5340 59.5399
R6186 gnd.n5009 gnd.n1482 59.5399
R6187 gnd.n5338 gnd.n1204 59.1804
R6188 gnd.n3570 gnd.n2120 57.3586
R6189 gnd.n2376 gnd.t217 56.607
R6190 gnd.n40 gnd.t186 56.607
R6191 gnd.n2353 gnd.t210 56.407
R6192 gnd.n2364 gnd.t250 56.407
R6193 gnd.n17 gnd.t285 56.407
R6194 gnd.n28 gnd.t54 56.407
R6195 gnd.n2385 gnd.t258 55.8337
R6196 gnd.n2362 gnd.t181 55.8337
R6197 gnd.n2373 gnd.t264 55.8337
R6198 gnd.n49 gnd.t271 55.8337
R6199 gnd.n26 gnd.t257 55.8337
R6200 gnd.n37 gnd.t213 55.8337
R6201 gnd.n1192 gnd.n1191 54.358
R6202 gnd.n1452 gnd.n1451 54.358
R6203 gnd.n2376 gnd.n2375 53.0052
R6204 gnd.n2378 gnd.n2377 53.0052
R6205 gnd.n2380 gnd.n2379 53.0052
R6206 gnd.n2382 gnd.n2381 53.0052
R6207 gnd.n2384 gnd.n2383 53.0052
R6208 gnd.n2353 gnd.n2352 53.0052
R6209 gnd.n2355 gnd.n2354 53.0052
R6210 gnd.n2357 gnd.n2356 53.0052
R6211 gnd.n2359 gnd.n2358 53.0052
R6212 gnd.n2361 gnd.n2360 53.0052
R6213 gnd.n2364 gnd.n2363 53.0052
R6214 gnd.n2366 gnd.n2365 53.0052
R6215 gnd.n2368 gnd.n2367 53.0052
R6216 gnd.n2370 gnd.n2369 53.0052
R6217 gnd.n2372 gnd.n2371 53.0052
R6218 gnd.n48 gnd.n47 53.0052
R6219 gnd.n46 gnd.n45 53.0052
R6220 gnd.n44 gnd.n43 53.0052
R6221 gnd.n42 gnd.n41 53.0052
R6222 gnd.n40 gnd.n39 53.0052
R6223 gnd.n25 gnd.n24 53.0052
R6224 gnd.n23 gnd.n22 53.0052
R6225 gnd.n21 gnd.n20 53.0052
R6226 gnd.n19 gnd.n18 53.0052
R6227 gnd.n17 gnd.n16 53.0052
R6228 gnd.n36 gnd.n35 53.0052
R6229 gnd.n34 gnd.n33 53.0052
R6230 gnd.n32 gnd.n31 53.0052
R6231 gnd.n30 gnd.n29 53.0052
R6232 gnd.n28 gnd.n27 53.0052
R6233 gnd.n1443 gnd.n1442 52.4801
R6234 gnd.n3422 gnd.t64 52.3082
R6235 gnd.n3390 gnd.t276 52.3082
R6236 gnd.n3358 gnd.t279 52.3082
R6237 gnd.n3327 gnd.t202 52.3082
R6238 gnd.n3295 gnd.t25 52.3082
R6239 gnd.n3263 gnd.t23 52.3082
R6240 gnd.n3231 gnd.t191 52.3082
R6241 gnd.n3200 gnd.t288 52.3082
R6242 gnd.n3252 gnd.n3220 51.4173
R6243 gnd.n3316 gnd.n3315 50.455
R6244 gnd.n3284 gnd.n3283 50.455
R6245 gnd.n3252 gnd.n3251 50.455
R6246 gnd.n6359 gnd.n435 45.6325
R6247 gnd.n5408 gnd.n5407 45.6325
R6248 gnd.n2664 gnd.n2663 45.1884
R6249 gnd.n2186 gnd.n2185 45.1884
R6250 gnd.n5060 gnd.n1458 44.3322
R6251 gnd.n1195 gnd.n1194 44.3189
R6252 gnd.n4210 gnd.n1866 42.2793
R6253 gnd.n2665 gnd.n2664 42.2793
R6254 gnd.n2187 gnd.n2186 42.2793
R6255 gnd.n2591 gnd.n2590 42.2793
R6256 gnd.n3537 gnd.n2160 42.2793
R6257 gnd.n6640 gnd.n6636 42.2793
R6258 gnd.n377 gnd.n376 42.2793
R6259 gnd.n1979 gnd.n1976 42.2793
R6260 gnd.n462 gnd.n461 42.2793
R6261 gnd.n6692 gnd.n157 42.2793
R6262 gnd.n6729 gnd.n6728 42.2793
R6263 gnd.n3842 gnd.n3728 42.2793
R6264 gnd.n3751 gnd.n3750 42.2793
R6265 gnd.n3601 gnd.n3600 42.2793
R6266 gnd.n4140 gnd.n4082 42.2793
R6267 gnd.n5171 gnd.n5098 42.2793
R6268 gnd.n1193 gnd.n1192 41.6274
R6269 gnd.n1453 gnd.n1452 41.6274
R6270 gnd.n1202 gnd.n1201 40.8975
R6271 gnd.n1456 gnd.n1455 40.8975
R6272 gnd.n6359 gnd.n439 36.9518
R6273 gnd.n5408 gnd.n1142 36.9518
R6274 gnd.n1201 gnd.n1200 35.055
R6275 gnd.n1196 gnd.n1195 35.055
R6276 gnd.n1445 gnd.n1444 35.055
R6277 gnd.n1455 gnd.n1441 35.055
R6278 gnd.n5662 gnd.n5661 34.6735
R6279 gnd.n5661 gnd.n5660 34.6735
R6280 gnd.n5660 gnd.n832 34.6735
R6281 gnd.n5654 gnd.n832 34.6735
R6282 gnd.n5654 gnd.n5653 34.6735
R6283 gnd.n5653 gnd.n5652 34.6735
R6284 gnd.n5652 gnd.n839 34.6735
R6285 gnd.n5646 gnd.n839 34.6735
R6286 gnd.n5646 gnd.n5645 34.6735
R6287 gnd.n5645 gnd.n5644 34.6735
R6288 gnd.n5644 gnd.n847 34.6735
R6289 gnd.n5638 gnd.n847 34.6735
R6290 gnd.n5638 gnd.n5637 34.6735
R6291 gnd.n5637 gnd.n5636 34.6735
R6292 gnd.n5636 gnd.n855 34.6735
R6293 gnd.n5630 gnd.n855 34.6735
R6294 gnd.n5630 gnd.n5629 34.6735
R6295 gnd.n5629 gnd.n5628 34.6735
R6296 gnd.n5628 gnd.n863 34.6735
R6297 gnd.n5622 gnd.n863 34.6735
R6298 gnd.n5622 gnd.n5621 34.6735
R6299 gnd.n5621 gnd.n5620 34.6735
R6300 gnd.n5620 gnd.n871 34.6735
R6301 gnd.n5614 gnd.n871 34.6735
R6302 gnd.n5614 gnd.n5613 34.6735
R6303 gnd.n5613 gnd.n5612 34.6735
R6304 gnd.n5612 gnd.n879 34.6735
R6305 gnd.n5606 gnd.n879 34.6735
R6306 gnd.n5606 gnd.n5605 34.6735
R6307 gnd.n5605 gnd.n5604 34.6735
R6308 gnd.n5604 gnd.n887 34.6735
R6309 gnd.n5598 gnd.n887 34.6735
R6310 gnd.n5598 gnd.n5597 34.6735
R6311 gnd.n5597 gnd.n5596 34.6735
R6312 gnd.n5596 gnd.n895 34.6735
R6313 gnd.n5590 gnd.n895 34.6735
R6314 gnd.n5590 gnd.n5589 34.6735
R6315 gnd.n5589 gnd.n5588 34.6735
R6316 gnd.n5588 gnd.n903 34.6735
R6317 gnd.n5582 gnd.n903 34.6735
R6318 gnd.n5582 gnd.n5581 34.6735
R6319 gnd.n5581 gnd.n5580 34.6735
R6320 gnd.n5580 gnd.n911 34.6735
R6321 gnd.n5574 gnd.n911 34.6735
R6322 gnd.n5574 gnd.n5573 34.6735
R6323 gnd.n5573 gnd.n5572 34.6735
R6324 gnd.n5572 gnd.n919 34.6735
R6325 gnd.n5566 gnd.n919 34.6735
R6326 gnd.n5566 gnd.n5565 34.6735
R6327 gnd.n5565 gnd.n5564 34.6735
R6328 gnd.n5564 gnd.n927 34.6735
R6329 gnd.n5558 gnd.n927 34.6735
R6330 gnd.n5558 gnd.n5557 34.6735
R6331 gnd.n5557 gnd.n5556 34.6735
R6332 gnd.n5556 gnd.n935 34.6735
R6333 gnd.n5550 gnd.n935 34.6735
R6334 gnd.n5550 gnd.n5549 34.6735
R6335 gnd.n5549 gnd.n5548 34.6735
R6336 gnd.n5548 gnd.n943 34.6735
R6337 gnd.n5542 gnd.n943 34.6735
R6338 gnd.n5542 gnd.n5541 34.6735
R6339 gnd.n5541 gnd.n5540 34.6735
R6340 gnd.n5540 gnd.n951 34.6735
R6341 gnd.n5534 gnd.n951 34.6735
R6342 gnd.n5534 gnd.n5533 34.6735
R6343 gnd.n5533 gnd.n5532 34.6735
R6344 gnd.n5532 gnd.n959 34.6735
R6345 gnd.n5526 gnd.n959 34.6735
R6346 gnd.n5526 gnd.n5525 34.6735
R6347 gnd.n5525 gnd.n5524 34.6735
R6348 gnd.n5524 gnd.n967 34.6735
R6349 gnd.n5518 gnd.n967 34.6735
R6350 gnd.n5518 gnd.n5517 34.6735
R6351 gnd.n5517 gnd.n5516 34.6735
R6352 gnd.n5516 gnd.n975 34.6735
R6353 gnd.n5510 gnd.n975 34.6735
R6354 gnd.n5510 gnd.n5509 34.6735
R6355 gnd.n5509 gnd.n5508 34.6735
R6356 gnd.n5508 gnd.n983 34.6735
R6357 gnd.n5502 gnd.n983 34.6735
R6358 gnd.n5502 gnd.n5501 34.6735
R6359 gnd.n5501 gnd.n5500 34.6735
R6360 gnd.n5500 gnd.n991 34.6735
R6361 gnd.n4943 gnd.n4940 32.9371
R6362 gnd.n1294 gnd.n1290 32.9371
R6363 gnd.n2727 gnd.n2621 31.8661
R6364 gnd.n2727 gnd.n2726 31.8661
R6365 gnd.n2735 gnd.n2610 31.8661
R6366 gnd.n2743 gnd.n2610 31.8661
R6367 gnd.n2743 gnd.n2604 31.8661
R6368 gnd.n2751 gnd.n2604 31.8661
R6369 gnd.n2751 gnd.n2597 31.8661
R6370 gnd.n2789 gnd.n2597 31.8661
R6371 gnd.n2799 gnd.n2530 31.8661
R6372 gnd.n3887 gnd.n2112 31.8661
R6373 gnd.n3895 gnd.n2104 31.8661
R6374 gnd.n3895 gnd.n2095 31.8661
R6375 gnd.n3903 gnd.n2095 31.8661
R6376 gnd.n3903 gnd.n2098 31.8661
R6377 gnd.n3911 gnd.n2080 31.8661
R6378 gnd.n3919 gnd.n2080 31.8661
R6379 gnd.n3927 gnd.n2072 31.8661
R6380 gnd.n3935 gnd.n2063 31.8661
R6381 gnd.n3935 gnd.n2066 31.8661
R6382 gnd.n3944 gnd.n2047 31.8661
R6383 gnd.n3956 gnd.n2047 31.8661
R6384 gnd.n3964 gnd.n2041 31.8661
R6385 gnd.n3991 gnd.n2029 31.8661
R6386 gnd.n3991 gnd.n2032 31.8661
R6387 gnd.n3999 gnd.n998 31.8661
R6388 gnd.n4185 gnd.n1095 31.8661
R6389 gnd.n1847 gnd.n1106 31.8661
R6390 gnd.n4234 gnd.n1847 31.8661
R6391 gnd.n4234 gnd.n1838 31.8661
R6392 gnd.n4251 gnd.n1838 31.8661
R6393 gnd.n4251 gnd.n1839 31.8661
R6394 gnd.n5197 gnd.n1419 31.8661
R6395 gnd.n5197 gnd.n1421 31.8661
R6396 gnd.n5181 gnd.n1421 31.8661
R6397 gnd.n5181 gnd.n5180 31.8661
R6398 gnd.n5180 gnd.n384 31.8661
R6399 gnd.n417 gnd.n328 31.8661
R6400 gnd.n6527 gnd.n247 31.8661
R6401 gnd.n6532 gnd.n235 31.8661
R6402 gnd.n6540 gnd.n235 31.8661
R6403 gnd.n6546 gnd.n230 31.8661
R6404 gnd.n6554 gnd.n222 31.8661
R6405 gnd.n6554 gnd.n224 31.8661
R6406 gnd.n6562 gnd.n202 31.8661
R6407 gnd.n6570 gnd.n202 31.8661
R6408 gnd.n6578 gnd.n194 31.8661
R6409 gnd.n6586 gnd.n186 31.8661
R6410 gnd.n6586 gnd.n188 31.8661
R6411 gnd.n6676 gnd.n169 31.8661
R6412 gnd.n6676 gnd.n161 31.8661
R6413 gnd.n6684 gnd.n161 31.8661
R6414 gnd.n6764 gnd.n81 31.8661
R6415 gnd.t218 gnd.n2041 31.5474
R6416 gnd.n6546 gnd.t7 31.5474
R6417 gnd.t232 gnd.n2072 30.9101
R6418 gnd.n6578 gnd.t40 30.9101
R6419 gnd.n6594 gnd.n179 28.6795
R6420 gnd.n5437 gnd.n1106 27.4049
R6421 gnd.n6390 gnd.n384 27.4049
R6422 gnd.n5493 gnd.n1001 26.7676
R6423 gnd.n4008 gnd.n1010 26.7676
R6424 gnd.n4030 gnd.n1021 26.7676
R6425 gnd.n5481 gnd.n1024 26.7676
R6426 gnd.n5475 gnd.n1035 26.7676
R6427 gnd.n4057 gnd.n4056 26.7676
R6428 gnd.n5469 gnd.n1045 26.7676
R6429 gnd.n4065 gnd.n1053 26.7676
R6430 gnd.n4162 gnd.n1063 26.7676
R6431 gnd.n5457 gnd.n1066 26.7676
R6432 gnd.n4073 gnd.n1074 26.7676
R6433 gnd.n5451 gnd.n1077 26.7676
R6434 gnd.n5445 gnd.n1088 26.7676
R6435 gnd.n4186 gnd.n4185 26.7676
R6436 gnd.n6445 gnd.n328 26.7676
R6437 gnd.n5150 gnd.n331 26.7676
R6438 gnd.n6310 gnd.n323 26.7676
R6439 gnd.n6461 gnd.n312 26.7676
R6440 gnd.n487 gnd.n315 26.7676
R6441 gnd.n6469 gnd.n303 26.7676
R6442 gnd.n6477 gnd.n294 26.7676
R6443 gnd.n497 gnd.n297 26.7676
R6444 gnd.n6485 gnd.n285 26.7676
R6445 gnd.n6217 gnd.n288 26.7676
R6446 gnd.n6221 gnd.n279 26.7676
R6447 gnd.n6502 gnd.n268 26.7676
R6448 gnd.n6514 gnd.n260 26.7676
R6449 gnd.n6519 gnd.n255 26.7676
R6450 gnd.n1866 gnd.n1865 25.7944
R6451 gnd.n2590 gnd.n2589 25.7944
R6452 gnd.n2160 gnd.n2159 25.7944
R6453 gnd.n6636 gnd.n6635 25.7944
R6454 gnd.n376 gnd.n375 25.7944
R6455 gnd.n1976 gnd.n1975 25.7944
R6456 gnd.n439 gnd.n438 25.7944
R6457 gnd.n461 gnd.n460 25.7944
R6458 gnd.n157 gnd.n156 25.7944
R6459 gnd.n6728 gnd.n6727 25.7944
R6460 gnd.n3728 gnd.n3727 25.7944
R6461 gnd.n3750 gnd.n3749 25.7944
R6462 gnd.n3600 gnd.n3599 25.7944
R6463 gnd.n4082 gnd.n4081 25.7944
R6464 gnd.n1142 gnd.n1141 25.7944
R6465 gnd.n5098 gnd.n5097 25.7944
R6466 gnd.n2811 gnd.n2531 24.8557
R6467 gnd.n2821 gnd.n2514 24.8557
R6468 gnd.n2517 gnd.n2505 24.8557
R6469 gnd.n2842 gnd.n2506 24.8557
R6470 gnd.n2852 gnd.n2486 24.8557
R6471 gnd.n2862 gnd.n2861 24.8557
R6472 gnd.n2472 gnd.n2470 24.8557
R6473 gnd.n2893 gnd.n2892 24.8557
R6474 gnd.n2908 gnd.n2455 24.8557
R6475 gnd.n2962 gnd.n2394 24.8557
R6476 gnd.n2918 gnd.n2395 24.8557
R6477 gnd.n2955 gnd.n2406 24.8557
R6478 gnd.n2444 gnd.n2443 24.8557
R6479 gnd.n2949 gnd.n2948 24.8557
R6480 gnd.n2430 gnd.n2417 24.8557
R6481 gnd.n2988 gnd.n2987 24.8557
R6482 gnd.n2998 gnd.n2338 24.8557
R6483 gnd.n3010 gnd.n2330 24.8557
R6484 gnd.n3009 gnd.n2318 24.8557
R6485 gnd.n3028 gnd.n3027 24.8557
R6486 gnd.n3038 gnd.n2311 24.8557
R6487 gnd.n3049 gnd.n2299 24.8557
R6488 gnd.n3073 gnd.n3072 24.8557
R6489 gnd.n3084 gnd.n2282 24.8557
R6490 gnd.n3083 gnd.n2284 24.8557
R6491 gnd.n3095 gnd.n2275 24.8557
R6492 gnd.n3113 gnd.n3112 24.8557
R6493 gnd.n2266 gnd.n2255 24.8557
R6494 gnd.n3134 gnd.n2243 24.8557
R6495 gnd.n3162 gnd.n3161 24.8557
R6496 gnd.n3173 gnd.n2228 24.8557
R6497 gnd.n3185 gnd.n2221 24.8557
R6498 gnd.n3457 gnd.n3456 24.8557
R6499 gnd.n3479 gnd.n2194 24.8557
R6500 gnd.n1228 gnd.n1227 23.855
R6501 gnd.n1488 gnd.n1487 23.855
R6502 gnd.n5340 gnd.n5339 23.855
R6503 gnd.n1482 gnd.n1481 23.855
R6504 gnd.n2832 gnd.t287 23.2624
R6505 gnd.n5404 gnd.n1181 23.2624
R6506 gnd.n1461 gnd.n1436 23.2624
R6507 gnd.n2533 gnd.t81 22.6251
R6508 gnd.n3927 gnd.t15 21.9878
R6509 gnd.t12 gnd.n194 21.9878
R6510 gnd.n5494 gnd.t17 21.6691
R6511 gnd.n5326 gnd.n1223 21.6691
R6512 gnd.n5314 gnd.n1308 21.6691
R6513 gnd.n4311 gnd.n1817 21.6691
R6514 gnd.n4457 gnd.n1807 21.6691
R6515 gnd.n4484 gnd.n1790 21.6691
R6516 gnd.n4509 gnd.n1774 21.6691
R6517 gnd.n4533 gnd.n1754 21.6691
R6518 gnd.n4555 gnd.n4554 21.6691
R6519 gnd.n4575 gnd.n1731 21.6691
R6520 gnd.n4581 gnd.n1727 21.6691
R6521 gnd.n4608 gnd.n1709 21.6691
R6522 gnd.n4633 gnd.n1693 21.6691
R6523 gnd.n4633 gnd.n1686 21.6691
R6524 gnd.n4656 gnd.n1673 21.6691
R6525 gnd.n4677 gnd.n4676 21.6691
R6526 gnd.n4697 gnd.n1648 21.6691
R6527 gnd.n4703 gnd.n1644 21.6691
R6528 gnd.n4719 gnd.n1629 21.6691
R6529 gnd.n4742 gnd.n4741 21.6691
R6530 gnd.n4822 gnd.n1583 21.6691
R6531 gnd.n4834 gnd.n1571 21.6691
R6532 gnd.n4858 gnd.n1553 21.6691
R6533 gnd.n4914 gnd.n1531 21.6691
R6534 gnd.n4936 gnd.n1433 21.6691
R6535 gnd.n6201 gnd.t246 21.6691
R6536 gnd.t201 gnd.n2538 21.3504
R6537 gnd.n3964 gnd.t195 21.3504
R6538 gnd.n3999 gnd.t38 21.3504
R6539 gnd.n6527 gnd.t30 21.3504
R6540 gnd.t193 gnd.n230 21.3504
R6541 gnd.n3183 gnd.n991 20.8043
R6542 gnd.n5338 gnd.n5337 20.7615
R6543 gnd.n5061 gnd.n5060 20.7615
R6544 gnd.t183 gnd.n2256 20.7131
R6545 gnd.n3944 gnd.t225 20.7131
R6546 gnd.n5487 gnd.t207 20.7131
R6547 gnd.n6287 gnd.t34 20.7131
R6548 gnd.n224 gnd.t178 20.7131
R6549 gnd.n5334 gnd.t78 20.3945
R6550 gnd.n5332 gnd.n1211 20.3945
R6551 gnd.n5320 gnd.n1302 20.3945
R6552 gnd.n4497 gnd.n1779 20.3945
R6553 gnd.n4515 gnd.n1769 20.3945
R6554 gnd.n4621 gnd.n1700 20.3945
R6555 gnd.n4639 gnd.n1689 20.3945
R6556 gnd.n4725 gnd.n1611 20.3945
R6557 gnd.n4805 gnd.n1598 20.3945
R6558 gnd.t67 gnd.n2291 20.0758
R6559 gnd.n3911 gnd.t180 20.0758
R6560 gnd.n5463 gnd.t209 20.0758
R6561 gnd.t99 gnd.t280 20.0758
R6562 gnd.n493 gnd.t53 20.0758
R6563 gnd.n188 gnd.t212 20.0758
R6564 gnd.n1189 gnd.t170 19.8005
R6565 gnd.n1189 gnd.t86 19.8005
R6566 gnd.n1190 gnd.t79 19.8005
R6567 gnd.n1190 gnd.t107 19.8005
R6568 gnd.n1449 gnd.t128 19.8005
R6569 gnd.n1449 gnd.t93 19.8005
R6570 gnd.n1450 gnd.t144 19.8005
R6571 gnd.n1450 gnd.t72 19.8005
R6572 gnd.n1186 gnd.n1185 19.5087
R6573 gnd.n1199 gnd.n1186 19.5087
R6574 gnd.n1197 gnd.n1188 19.5087
R6575 gnd.n1454 gnd.n1448 19.5087
R6576 gnd.n2999 gnd.t189 19.4385
R6577 gnd.n4229 gnd.n4228 19.3944
R6578 gnd.n4228 gnd.n4227 19.3944
R6579 gnd.n4227 gnd.n4220 19.3944
R6580 gnd.n4223 gnd.n4220 19.3944
R6581 gnd.n4223 gnd.n1830 19.3944
R6582 gnd.n4275 gnd.n1830 19.3944
R6583 gnd.n4275 gnd.n1827 19.3944
R6584 gnd.n4282 gnd.n1827 19.3944
R6585 gnd.n4282 gnd.n1828 19.3944
R6586 gnd.n4278 gnd.n1828 19.3944
R6587 gnd.n4278 gnd.n1328 19.3944
R6588 gnd.n5305 gnd.n1328 19.3944
R6589 gnd.n5305 gnd.n1329 19.3944
R6590 gnd.n5301 gnd.n1329 19.3944
R6591 gnd.n5301 gnd.n5300 19.3944
R6592 gnd.n5300 gnd.n5299 19.3944
R6593 gnd.n5299 gnd.n1335 19.3944
R6594 gnd.n5295 gnd.n1335 19.3944
R6595 gnd.n5295 gnd.n5294 19.3944
R6596 gnd.n5294 gnd.n5293 19.3944
R6597 gnd.n5293 gnd.n1340 19.3944
R6598 gnd.n5289 gnd.n1340 19.3944
R6599 gnd.n5289 gnd.n5288 19.3944
R6600 gnd.n5288 gnd.n5287 19.3944
R6601 gnd.n5287 gnd.n1345 19.3944
R6602 gnd.n5283 gnd.n1345 19.3944
R6603 gnd.n5283 gnd.n5282 19.3944
R6604 gnd.n5282 gnd.n5281 19.3944
R6605 gnd.n5281 gnd.n1350 19.3944
R6606 gnd.n5277 gnd.n1350 19.3944
R6607 gnd.n5277 gnd.n5276 19.3944
R6608 gnd.n5276 gnd.n5275 19.3944
R6609 gnd.n5275 gnd.n1355 19.3944
R6610 gnd.n5271 gnd.n1355 19.3944
R6611 gnd.n5271 gnd.n5270 19.3944
R6612 gnd.n5270 gnd.n5269 19.3944
R6613 gnd.n5269 gnd.n1360 19.3944
R6614 gnd.n5265 gnd.n1360 19.3944
R6615 gnd.n5265 gnd.n5264 19.3944
R6616 gnd.n5264 gnd.n5263 19.3944
R6617 gnd.n5263 gnd.n1365 19.3944
R6618 gnd.n5259 gnd.n1365 19.3944
R6619 gnd.n5259 gnd.n5258 19.3944
R6620 gnd.n5258 gnd.n5257 19.3944
R6621 gnd.n5257 gnd.n1370 19.3944
R6622 gnd.n5253 gnd.n1370 19.3944
R6623 gnd.n5253 gnd.n5252 19.3944
R6624 gnd.n5252 gnd.n5251 19.3944
R6625 gnd.n5251 gnd.n1375 19.3944
R6626 gnd.n5247 gnd.n1375 19.3944
R6627 gnd.n5247 gnd.n5246 19.3944
R6628 gnd.n5246 gnd.n5245 19.3944
R6629 gnd.n5245 gnd.n1380 19.3944
R6630 gnd.n5241 gnd.n1380 19.3944
R6631 gnd.n5241 gnd.n5240 19.3944
R6632 gnd.n5240 gnd.n5239 19.3944
R6633 gnd.n5239 gnd.n1385 19.3944
R6634 gnd.n5235 gnd.n1385 19.3944
R6635 gnd.n5235 gnd.n5234 19.3944
R6636 gnd.n5234 gnd.n5233 19.3944
R6637 gnd.n5233 gnd.n1390 19.3944
R6638 gnd.n5229 gnd.n1390 19.3944
R6639 gnd.n5229 gnd.n5228 19.3944
R6640 gnd.n5228 gnd.n5227 19.3944
R6641 gnd.n5227 gnd.n1395 19.3944
R6642 gnd.n5223 gnd.n1395 19.3944
R6643 gnd.n5223 gnd.n5222 19.3944
R6644 gnd.n5222 gnd.n5221 19.3944
R6645 gnd.n5221 gnd.n1400 19.3944
R6646 gnd.n5217 gnd.n1400 19.3944
R6647 gnd.n5217 gnd.n5216 19.3944
R6648 gnd.n5216 gnd.n5215 19.3944
R6649 gnd.n5215 gnd.n1405 19.3944
R6650 gnd.n5211 gnd.n1405 19.3944
R6651 gnd.n5211 gnd.n5210 19.3944
R6652 gnd.n5210 gnd.n5209 19.3944
R6653 gnd.n5209 gnd.n1410 19.3944
R6654 gnd.n5205 gnd.n1410 19.3944
R6655 gnd.n5205 gnd.n5204 19.3944
R6656 gnd.n5204 gnd.n5203 19.3944
R6657 gnd.n5203 gnd.n1415 19.3944
R6658 gnd.n5199 gnd.n1415 19.3944
R6659 gnd.n4214 gnd.n4211 19.3944
R6660 gnd.n4214 gnd.n1863 19.3944
R6661 gnd.n4232 gnd.n1863 19.3944
R6662 gnd.n1919 gnd.n1906 19.3944
R6663 gnd.n1922 gnd.n1919 19.3944
R6664 gnd.n1922 gnd.n1900 19.3944
R6665 gnd.n1931 gnd.n1900 19.3944
R6666 gnd.n1934 gnd.n1931 19.3944
R6667 gnd.n1934 gnd.n1894 19.3944
R6668 gnd.n1943 gnd.n1894 19.3944
R6669 gnd.n1946 gnd.n1943 19.3944
R6670 gnd.n1946 gnd.n1888 19.3944
R6671 gnd.n1955 gnd.n1888 19.3944
R6672 gnd.n1958 gnd.n1955 19.3944
R6673 gnd.n1958 gnd.n1882 19.3944
R6674 gnd.n1967 gnd.n1882 19.3944
R6675 gnd.n1970 gnd.n1967 19.3944
R6676 gnd.n1970 gnd.n1876 19.3944
R6677 gnd.n4192 gnd.n1876 19.3944
R6678 gnd.n4193 gnd.n4192 19.3944
R6679 gnd.n4196 gnd.n4193 19.3944
R6680 gnd.n4196 gnd.n1871 19.3944
R6681 gnd.n4201 gnd.n1871 19.3944
R6682 gnd.n4202 gnd.n4201 19.3944
R6683 gnd.n4205 gnd.n4202 19.3944
R6684 gnd.n4205 gnd.n1867 19.3944
R6685 gnd.n4209 gnd.n1867 19.3944
R6686 gnd.n2714 gnd.n2713 19.3944
R6687 gnd.n2713 gnd.n2712 19.3944
R6688 gnd.n2712 gnd.n2711 19.3944
R6689 gnd.n2711 gnd.n2709 19.3944
R6690 gnd.n2709 gnd.n2706 19.3944
R6691 gnd.n2706 gnd.n2705 19.3944
R6692 gnd.n2705 gnd.n2702 19.3944
R6693 gnd.n2702 gnd.n2701 19.3944
R6694 gnd.n2701 gnd.n2698 19.3944
R6695 gnd.n2698 gnd.n2697 19.3944
R6696 gnd.n2697 gnd.n2694 19.3944
R6697 gnd.n2694 gnd.n2693 19.3944
R6698 gnd.n2693 gnd.n2690 19.3944
R6699 gnd.n2690 gnd.n2689 19.3944
R6700 gnd.n2689 gnd.n2686 19.3944
R6701 gnd.n2686 gnd.n2685 19.3944
R6702 gnd.n2685 gnd.n2682 19.3944
R6703 gnd.n2682 gnd.n2681 19.3944
R6704 gnd.n2681 gnd.n2678 19.3944
R6705 gnd.n2678 gnd.n2677 19.3944
R6706 gnd.n2677 gnd.n2674 19.3944
R6707 gnd.n2674 gnd.n2673 19.3944
R6708 gnd.n2670 gnd.n2669 19.3944
R6709 gnd.n2669 gnd.n2625 19.3944
R6710 gnd.n2720 gnd.n2625 19.3944
R6711 gnd.n3487 gnd.n3486 19.3944
R6712 gnd.n3486 gnd.n3483 19.3944
R6713 gnd.n3483 gnd.n3482 19.3944
R6714 gnd.n3532 gnd.n3531 19.3944
R6715 gnd.n3531 gnd.n3530 19.3944
R6716 gnd.n3530 gnd.n3527 19.3944
R6717 gnd.n3527 gnd.n3526 19.3944
R6718 gnd.n3526 gnd.n3523 19.3944
R6719 gnd.n3523 gnd.n3522 19.3944
R6720 gnd.n3522 gnd.n3519 19.3944
R6721 gnd.n3519 gnd.n3518 19.3944
R6722 gnd.n3518 gnd.n3515 19.3944
R6723 gnd.n3515 gnd.n3514 19.3944
R6724 gnd.n3514 gnd.n3511 19.3944
R6725 gnd.n3511 gnd.n3510 19.3944
R6726 gnd.n3510 gnd.n3507 19.3944
R6727 gnd.n3507 gnd.n3506 19.3944
R6728 gnd.n3506 gnd.n3503 19.3944
R6729 gnd.n3503 gnd.n3502 19.3944
R6730 gnd.n3502 gnd.n3499 19.3944
R6731 gnd.n3499 gnd.n3498 19.3944
R6732 gnd.n3498 gnd.n3495 19.3944
R6733 gnd.n3495 gnd.n3494 19.3944
R6734 gnd.n3494 gnd.n3491 19.3944
R6735 gnd.n3491 gnd.n3490 19.3944
R6736 gnd.n2813 gnd.n2522 19.3944
R6737 gnd.n2823 gnd.n2522 19.3944
R6738 gnd.n2824 gnd.n2823 19.3944
R6739 gnd.n2824 gnd.n2503 19.3944
R6740 gnd.n2844 gnd.n2503 19.3944
R6741 gnd.n2844 gnd.n2495 19.3944
R6742 gnd.n2854 gnd.n2495 19.3944
R6743 gnd.n2855 gnd.n2854 19.3944
R6744 gnd.n2856 gnd.n2855 19.3944
R6745 gnd.n2856 gnd.n2478 19.3944
R6746 gnd.n2873 gnd.n2478 19.3944
R6747 gnd.n2876 gnd.n2873 19.3944
R6748 gnd.n2876 gnd.n2875 19.3944
R6749 gnd.n2875 gnd.n2451 19.3944
R6750 gnd.n2915 gnd.n2451 19.3944
R6751 gnd.n2915 gnd.n2448 19.3944
R6752 gnd.n2921 gnd.n2448 19.3944
R6753 gnd.n2922 gnd.n2921 19.3944
R6754 gnd.n2922 gnd.n2446 19.3944
R6755 gnd.n2928 gnd.n2446 19.3944
R6756 gnd.n2931 gnd.n2928 19.3944
R6757 gnd.n2933 gnd.n2931 19.3944
R6758 gnd.n2939 gnd.n2933 19.3944
R6759 gnd.n2939 gnd.n2938 19.3944
R6760 gnd.n2938 gnd.n2333 19.3944
R6761 gnd.n3005 gnd.n2333 19.3944
R6762 gnd.n3006 gnd.n3005 19.3944
R6763 gnd.n3006 gnd.n2326 19.3944
R6764 gnd.n3017 gnd.n2326 19.3944
R6765 gnd.n3018 gnd.n3017 19.3944
R6766 gnd.n3018 gnd.n2309 19.3944
R6767 gnd.n2309 gnd.n2307 19.3944
R6768 gnd.n3042 gnd.n2307 19.3944
R6769 gnd.n3043 gnd.n3042 19.3944
R6770 gnd.n3043 gnd.n2278 19.3944
R6771 gnd.n3090 gnd.n2278 19.3944
R6772 gnd.n3091 gnd.n3090 19.3944
R6773 gnd.n3091 gnd.n2271 19.3944
R6774 gnd.n3102 gnd.n2271 19.3944
R6775 gnd.n3103 gnd.n3102 19.3944
R6776 gnd.n3103 gnd.n2254 19.3944
R6777 gnd.n2254 gnd.n2252 19.3944
R6778 gnd.n3127 gnd.n2252 19.3944
R6779 gnd.n3128 gnd.n3127 19.3944
R6780 gnd.n3128 gnd.n2224 19.3944
R6781 gnd.n3179 gnd.n2224 19.3944
R6782 gnd.n3180 gnd.n3179 19.3944
R6783 gnd.n3180 gnd.n2217 19.3944
R6784 gnd.n3448 gnd.n2217 19.3944
R6785 gnd.n3449 gnd.n3448 19.3944
R6786 gnd.n3449 gnd.n2198 19.3944
R6787 gnd.n3474 gnd.n2198 19.3944
R6788 gnd.n3474 gnd.n2199 19.3944
R6789 gnd.n2804 gnd.n2803 19.3944
R6790 gnd.n2803 gnd.n2536 19.3944
R6791 gnd.n2559 gnd.n2536 19.3944
R6792 gnd.n2562 gnd.n2559 19.3944
R6793 gnd.n2562 gnd.n2555 19.3944
R6794 gnd.n2566 gnd.n2555 19.3944
R6795 gnd.n2569 gnd.n2566 19.3944
R6796 gnd.n2572 gnd.n2569 19.3944
R6797 gnd.n2572 gnd.n2553 19.3944
R6798 gnd.n2576 gnd.n2553 19.3944
R6799 gnd.n2579 gnd.n2576 19.3944
R6800 gnd.n2582 gnd.n2579 19.3944
R6801 gnd.n2582 gnd.n2551 19.3944
R6802 gnd.n2586 gnd.n2551 19.3944
R6803 gnd.n2809 gnd.n2808 19.3944
R6804 gnd.n2808 gnd.n2512 19.3944
R6805 gnd.n2834 gnd.n2512 19.3944
R6806 gnd.n2834 gnd.n2510 19.3944
R6807 gnd.n2840 gnd.n2510 19.3944
R6808 gnd.n2840 gnd.n2839 19.3944
R6809 gnd.n2839 gnd.n2484 19.3944
R6810 gnd.n2864 gnd.n2484 19.3944
R6811 gnd.n2864 gnd.n2482 19.3944
R6812 gnd.n2868 gnd.n2482 19.3944
R6813 gnd.n2868 gnd.n2462 19.3944
R6814 gnd.n2895 gnd.n2462 19.3944
R6815 gnd.n2895 gnd.n2460 19.3944
R6816 gnd.n2905 gnd.n2460 19.3944
R6817 gnd.n2905 gnd.n2904 19.3944
R6818 gnd.n2904 gnd.n2903 19.3944
R6819 gnd.n2903 gnd.n2409 19.3944
R6820 gnd.n2953 gnd.n2409 19.3944
R6821 gnd.n2953 gnd.n2952 19.3944
R6822 gnd.n2952 gnd.n2951 19.3944
R6823 gnd.n2951 gnd.n2413 19.3944
R6824 gnd.n2433 gnd.n2413 19.3944
R6825 gnd.n2433 gnd.n2343 19.3944
R6826 gnd.n2990 gnd.n2343 19.3944
R6827 gnd.n2990 gnd.n2341 19.3944
R6828 gnd.n2996 gnd.n2341 19.3944
R6829 gnd.n2996 gnd.n2995 19.3944
R6830 gnd.n2995 gnd.n2316 19.3944
R6831 gnd.n3030 gnd.n2316 19.3944
R6832 gnd.n3030 gnd.n2314 19.3944
R6833 gnd.n3036 gnd.n2314 19.3944
R6834 gnd.n3036 gnd.n3035 19.3944
R6835 gnd.n3035 gnd.n2289 19.3944
R6836 gnd.n3075 gnd.n2289 19.3944
R6837 gnd.n3075 gnd.n2287 19.3944
R6838 gnd.n3081 gnd.n2287 19.3944
R6839 gnd.n3081 gnd.n3080 19.3944
R6840 gnd.n3080 gnd.n2261 19.3944
R6841 gnd.n3115 gnd.n2261 19.3944
R6842 gnd.n3115 gnd.n2259 19.3944
R6843 gnd.n3121 gnd.n2259 19.3944
R6844 gnd.n3121 gnd.n3120 19.3944
R6845 gnd.n3120 gnd.n2234 19.3944
R6846 gnd.n3164 gnd.n2234 19.3944
R6847 gnd.n3164 gnd.n2232 19.3944
R6848 gnd.n3170 gnd.n2232 19.3944
R6849 gnd.n3170 gnd.n3169 19.3944
R6850 gnd.n3169 gnd.n2207 19.3944
R6851 gnd.n3459 gnd.n2207 19.3944
R6852 gnd.n3459 gnd.n2205 19.3944
R6853 gnd.n3467 gnd.n2205 19.3944
R6854 gnd.n3467 gnd.n3466 19.3944
R6855 gnd.n3466 gnd.n3465 19.3944
R6856 gnd.n3568 gnd.n3567 19.3944
R6857 gnd.n3567 gnd.n2146 19.3944
R6858 gnd.n3563 gnd.n2146 19.3944
R6859 gnd.n3563 gnd.n3560 19.3944
R6860 gnd.n3560 gnd.n3557 19.3944
R6861 gnd.n3557 gnd.n3556 19.3944
R6862 gnd.n3556 gnd.n3553 19.3944
R6863 gnd.n3553 gnd.n3552 19.3944
R6864 gnd.n3552 gnd.n3549 19.3944
R6865 gnd.n3549 gnd.n3548 19.3944
R6866 gnd.n3548 gnd.n3545 19.3944
R6867 gnd.n3545 gnd.n3544 19.3944
R6868 gnd.n3544 gnd.n3541 19.3944
R6869 gnd.n3541 gnd.n3540 19.3944
R6870 gnd.n2724 gnd.n2623 19.3944
R6871 gnd.n2724 gnd.n2614 19.3944
R6872 gnd.n2737 gnd.n2614 19.3944
R6873 gnd.n2737 gnd.n2612 19.3944
R6874 gnd.n2741 gnd.n2612 19.3944
R6875 gnd.n2741 gnd.n2602 19.3944
R6876 gnd.n2753 gnd.n2602 19.3944
R6877 gnd.n2753 gnd.n2600 19.3944
R6878 gnd.n2787 gnd.n2600 19.3944
R6879 gnd.n2787 gnd.n2786 19.3944
R6880 gnd.n2786 gnd.n2785 19.3944
R6881 gnd.n2785 gnd.n2784 19.3944
R6882 gnd.n2784 gnd.n2781 19.3944
R6883 gnd.n2781 gnd.n2780 19.3944
R6884 gnd.n2780 gnd.n2779 19.3944
R6885 gnd.n2779 gnd.n2777 19.3944
R6886 gnd.n2777 gnd.n2776 19.3944
R6887 gnd.n2776 gnd.n2773 19.3944
R6888 gnd.n2773 gnd.n2772 19.3944
R6889 gnd.n2772 gnd.n2771 19.3944
R6890 gnd.n2771 gnd.n2769 19.3944
R6891 gnd.n2769 gnd.n2468 19.3944
R6892 gnd.n2884 gnd.n2468 19.3944
R6893 gnd.n2884 gnd.n2466 19.3944
R6894 gnd.n2890 gnd.n2466 19.3944
R6895 gnd.n2890 gnd.n2889 19.3944
R6896 gnd.n2889 gnd.n2390 19.3944
R6897 gnd.n2964 gnd.n2390 19.3944
R6898 gnd.n2964 gnd.n2391 19.3944
R6899 gnd.n2438 gnd.n2437 19.3944
R6900 gnd.n2441 gnd.n2440 19.3944
R6901 gnd.n2428 gnd.n2427 19.3944
R6902 gnd.n2983 gnd.n2348 19.3944
R6903 gnd.n2983 gnd.n2982 19.3944
R6904 gnd.n2982 gnd.n2981 19.3944
R6905 gnd.n2981 gnd.n2979 19.3944
R6906 gnd.n2979 gnd.n2978 19.3944
R6907 gnd.n2978 gnd.n2976 19.3944
R6908 gnd.n2976 gnd.n2975 19.3944
R6909 gnd.n2975 gnd.n2297 19.3944
R6910 gnd.n3051 gnd.n2297 19.3944
R6911 gnd.n3051 gnd.n2295 19.3944
R6912 gnd.n3070 gnd.n2295 19.3944
R6913 gnd.n3070 gnd.n3069 19.3944
R6914 gnd.n3069 gnd.n3068 19.3944
R6915 gnd.n3068 gnd.n3066 19.3944
R6916 gnd.n3066 gnd.n3065 19.3944
R6917 gnd.n3065 gnd.n3063 19.3944
R6918 gnd.n3063 gnd.n3062 19.3944
R6919 gnd.n3062 gnd.n2241 19.3944
R6920 gnd.n3136 gnd.n2241 19.3944
R6921 gnd.n3136 gnd.n2239 19.3944
R6922 gnd.n3159 gnd.n2239 19.3944
R6923 gnd.n3159 gnd.n3158 19.3944
R6924 gnd.n3158 gnd.n3157 19.3944
R6925 gnd.n3157 gnd.n3154 19.3944
R6926 gnd.n3154 gnd.n3153 19.3944
R6927 gnd.n3153 gnd.n3151 19.3944
R6928 gnd.n3151 gnd.n3150 19.3944
R6929 gnd.n3150 gnd.n3148 19.3944
R6930 gnd.n3148 gnd.n2193 19.3944
R6931 gnd.n2729 gnd.n2619 19.3944
R6932 gnd.n2729 gnd.n2617 19.3944
R6933 gnd.n2733 gnd.n2617 19.3944
R6934 gnd.n2733 gnd.n2608 19.3944
R6935 gnd.n2745 gnd.n2608 19.3944
R6936 gnd.n2745 gnd.n2606 19.3944
R6937 gnd.n2749 gnd.n2606 19.3944
R6938 gnd.n2749 gnd.n2595 19.3944
R6939 gnd.n2791 gnd.n2595 19.3944
R6940 gnd.n2791 gnd.n2549 19.3944
R6941 gnd.n2797 gnd.n2549 19.3944
R6942 gnd.n2797 gnd.n2796 19.3944
R6943 gnd.n2796 gnd.n2527 19.3944
R6944 gnd.n2818 gnd.n2527 19.3944
R6945 gnd.n2818 gnd.n2520 19.3944
R6946 gnd.n2829 gnd.n2520 19.3944
R6947 gnd.n2829 gnd.n2828 19.3944
R6948 gnd.n2828 gnd.n2501 19.3944
R6949 gnd.n2849 gnd.n2501 19.3944
R6950 gnd.n2849 gnd.n2491 19.3944
R6951 gnd.n2859 gnd.n2491 19.3944
R6952 gnd.n2859 gnd.n2474 19.3944
R6953 gnd.n2880 gnd.n2474 19.3944
R6954 gnd.n2880 gnd.n2879 19.3944
R6955 gnd.n2879 gnd.n2453 19.3944
R6956 gnd.n2910 gnd.n2453 19.3944
R6957 gnd.n2910 gnd.n2398 19.3944
R6958 gnd.n2960 gnd.n2398 19.3944
R6959 gnd.n2960 gnd.n2959 19.3944
R6960 gnd.n2959 gnd.n2958 19.3944
R6961 gnd.n2958 gnd.n2402 19.3944
R6962 gnd.n2420 gnd.n2402 19.3944
R6963 gnd.n2946 gnd.n2420 19.3944
R6964 gnd.n2946 gnd.n2945 19.3944
R6965 gnd.n2945 gnd.n2944 19.3944
R6966 gnd.n2944 gnd.n2424 19.3944
R6967 gnd.n2424 gnd.n2335 19.3944
R6968 gnd.n3001 gnd.n2335 19.3944
R6969 gnd.n3001 gnd.n2328 19.3944
R6970 gnd.n3012 gnd.n2328 19.3944
R6971 gnd.n3012 gnd.n2324 19.3944
R6972 gnd.n3025 gnd.n2324 19.3944
R6973 gnd.n3025 gnd.n3024 19.3944
R6974 gnd.n3024 gnd.n2303 19.3944
R6975 gnd.n3047 gnd.n2303 19.3944
R6976 gnd.n3047 gnd.n3046 19.3944
R6977 gnd.n3046 gnd.n2280 19.3944
R6978 gnd.n3086 gnd.n2280 19.3944
R6979 gnd.n3086 gnd.n2273 19.3944
R6980 gnd.n3097 gnd.n2273 19.3944
R6981 gnd.n3097 gnd.n2269 19.3944
R6982 gnd.n3110 gnd.n2269 19.3944
R6983 gnd.n3110 gnd.n3109 19.3944
R6984 gnd.n3109 gnd.n2248 19.3944
R6985 gnd.n3132 gnd.n2248 19.3944
R6986 gnd.n3132 gnd.n3131 19.3944
R6987 gnd.n3131 gnd.n2226 19.3944
R6988 gnd.n3175 gnd.n2226 19.3944
R6989 gnd.n3175 gnd.n2219 19.3944
R6990 gnd.n3187 gnd.n2219 19.3944
R6991 gnd.n3187 gnd.n2215 19.3944
R6992 gnd.n3454 gnd.n2215 19.3944
R6993 gnd.n3454 gnd.n3453 19.3944
R6994 gnd.n3453 gnd.n2196 19.3944
R6995 gnd.n3477 gnd.n2196 19.3944
R6996 gnd.n5153 gnd.n5152 19.3944
R6997 gnd.n5152 gnd.n468 19.3944
R6998 gnd.n6308 gnd.n468 19.3944
R6999 gnd.n6308 gnd.n469 19.3944
R7000 gnd.n6304 gnd.n469 19.3944
R7001 gnd.n6304 gnd.n6303 19.3944
R7002 gnd.n6303 gnd.n6302 19.3944
R7003 gnd.n6302 gnd.n474 19.3944
R7004 gnd.n6298 gnd.n474 19.3944
R7005 gnd.n6298 gnd.n6297 19.3944
R7006 gnd.n6297 gnd.n6296 19.3944
R7007 gnd.n6296 gnd.n478 19.3944
R7008 gnd.n6292 gnd.n478 19.3944
R7009 gnd.n6292 gnd.n6291 19.3944
R7010 gnd.n6291 gnd.n6290 19.3944
R7011 gnd.n6290 gnd.n253 19.3944
R7012 gnd.n6521 gnd.n253 19.3944
R7013 gnd.n6521 gnd.n250 19.3944
R7014 gnd.n6525 gnd.n250 19.3944
R7015 gnd.n6525 gnd.n251 19.3944
R7016 gnd.n251 gnd.n52 19.3944
R7017 gnd.n6796 gnd.n52 19.3944
R7018 gnd.n6796 gnd.n6795 19.3944
R7019 gnd.n6795 gnd.n6794 19.3944
R7020 gnd.n6794 gnd.n57 19.3944
R7021 gnd.n6790 gnd.n57 19.3944
R7022 gnd.n6790 gnd.n6789 19.3944
R7023 gnd.n6789 gnd.n6788 19.3944
R7024 gnd.n6788 gnd.n62 19.3944
R7025 gnd.n6784 gnd.n62 19.3944
R7026 gnd.n6784 gnd.n6783 19.3944
R7027 gnd.n6783 gnd.n6782 19.3944
R7028 gnd.n6782 gnd.n67 19.3944
R7029 gnd.n6778 gnd.n67 19.3944
R7030 gnd.n6778 gnd.n6777 19.3944
R7031 gnd.n6777 gnd.n6776 19.3944
R7032 gnd.n6776 gnd.n72 19.3944
R7033 gnd.n6772 gnd.n72 19.3944
R7034 gnd.n6772 gnd.n6771 19.3944
R7035 gnd.n6771 gnd.n6770 19.3944
R7036 gnd.n6770 gnd.n77 19.3944
R7037 gnd.n6766 gnd.n77 19.3944
R7038 gnd.n6665 gnd.n6664 19.3944
R7039 gnd.n6664 gnd.n6663 19.3944
R7040 gnd.n6663 gnd.n6606 19.3944
R7041 gnd.n6659 gnd.n6606 19.3944
R7042 gnd.n6659 gnd.n6658 19.3944
R7043 gnd.n6658 gnd.n6657 19.3944
R7044 gnd.n6657 gnd.n6614 19.3944
R7045 gnd.n6653 gnd.n6614 19.3944
R7046 gnd.n6653 gnd.n6652 19.3944
R7047 gnd.n6652 gnd.n6651 19.3944
R7048 gnd.n6651 gnd.n6622 19.3944
R7049 gnd.n6647 gnd.n6622 19.3944
R7050 gnd.n6647 gnd.n6646 19.3944
R7051 gnd.n6646 gnd.n6645 19.3944
R7052 gnd.n6645 gnd.n6630 19.3944
R7053 gnd.n6641 gnd.n6630 19.3944
R7054 gnd.n6440 gnd.n6439 19.3944
R7055 gnd.n6439 gnd.n335 19.3944
R7056 gnd.n6432 gnd.n335 19.3944
R7057 gnd.n6432 gnd.n6431 19.3944
R7058 gnd.n6431 gnd.n343 19.3944
R7059 gnd.n6424 gnd.n343 19.3944
R7060 gnd.n6424 gnd.n6423 19.3944
R7061 gnd.n6423 gnd.n351 19.3944
R7062 gnd.n6416 gnd.n351 19.3944
R7063 gnd.n6416 gnd.n6415 19.3944
R7064 gnd.n6415 gnd.n359 19.3944
R7065 gnd.n6408 gnd.n359 19.3944
R7066 gnd.n6408 gnd.n6407 19.3944
R7067 gnd.n6407 gnd.n367 19.3944
R7068 gnd.n6400 gnd.n367 19.3944
R7069 gnd.n6400 gnd.n6399 19.3944
R7070 gnd.n6443 gnd.n319 19.3944
R7071 gnd.n6455 gnd.n319 19.3944
R7072 gnd.n6455 gnd.n317 19.3944
R7073 gnd.n6459 gnd.n317 19.3944
R7074 gnd.n6459 gnd.n301 19.3944
R7075 gnd.n6471 gnd.n301 19.3944
R7076 gnd.n6471 gnd.n299 19.3944
R7077 gnd.n6475 gnd.n299 19.3944
R7078 gnd.n6475 gnd.n283 19.3944
R7079 gnd.n6487 gnd.n283 19.3944
R7080 gnd.n6487 gnd.n281 19.3944
R7081 gnd.n6491 gnd.n281 19.3944
R7082 gnd.n6491 gnd.n266 19.3944
R7083 gnd.n6504 gnd.n266 19.3944
R7084 gnd.n6504 gnd.n263 19.3944
R7085 gnd.n6512 gnd.n263 19.3944
R7086 gnd.n6512 gnd.n264 19.3944
R7087 gnd.n6508 gnd.n264 19.3944
R7088 gnd.n6508 gnd.n241 19.3944
R7089 gnd.n6534 gnd.n241 19.3944
R7090 gnd.n6534 gnd.n238 19.3944
R7091 gnd.n6538 gnd.n238 19.3944
R7092 gnd.n6538 gnd.n228 19.3944
R7093 gnd.n6548 gnd.n228 19.3944
R7094 gnd.n6548 gnd.n226 19.3944
R7095 gnd.n6552 gnd.n226 19.3944
R7096 gnd.n6552 gnd.n207 19.3944
R7097 gnd.n6564 gnd.n207 19.3944
R7098 gnd.n6564 gnd.n205 19.3944
R7099 gnd.n6568 gnd.n205 19.3944
R7100 gnd.n6568 gnd.n192 19.3944
R7101 gnd.n6580 gnd.n192 19.3944
R7102 gnd.n6580 gnd.n190 19.3944
R7103 gnd.n6584 gnd.n190 19.3944
R7104 gnd.n6584 gnd.n176 19.3944
R7105 gnd.n6596 gnd.n176 19.3944
R7106 gnd.n6596 gnd.n173 19.3944
R7107 gnd.n6674 gnd.n173 19.3944
R7108 gnd.n6674 gnd.n174 19.3944
R7109 gnd.n6670 gnd.n174 19.3944
R7110 gnd.n6670 gnd.n6669 19.3944
R7111 gnd.n6669 gnd.n6668 19.3944
R7112 gnd.n1913 gnd.n1910 19.3944
R7113 gnd.n1916 gnd.n1913 19.3944
R7114 gnd.n1916 gnd.n1904 19.3944
R7115 gnd.n1925 gnd.n1904 19.3944
R7116 gnd.n1928 gnd.n1925 19.3944
R7117 gnd.n1928 gnd.n1896 19.3944
R7118 gnd.n1937 gnd.n1896 19.3944
R7119 gnd.n1940 gnd.n1937 19.3944
R7120 gnd.n1940 gnd.n1892 19.3944
R7121 gnd.n1949 gnd.n1892 19.3944
R7122 gnd.n1952 gnd.n1949 19.3944
R7123 gnd.n1952 gnd.n1884 19.3944
R7124 gnd.n1961 gnd.n1884 19.3944
R7125 gnd.n1964 gnd.n1961 19.3944
R7126 gnd.n1964 gnd.n1880 19.3944
R7127 gnd.n1974 gnd.n1880 19.3944
R7128 gnd.n4038 gnd.n4036 19.3944
R7129 gnd.n4038 gnd.n4033 19.3944
R7130 gnd.n4042 gnd.n4033 19.3944
R7131 gnd.n4042 gnd.n2011 19.3944
R7132 gnd.n4046 gnd.n2011 19.3944
R7133 gnd.n4046 gnd.n2009 19.3944
R7134 gnd.n4054 gnd.n2009 19.3944
R7135 gnd.n4054 gnd.n4053 19.3944
R7136 gnd.n4053 gnd.n4052 19.3944
R7137 gnd.n4052 gnd.n1990 19.3944
R7138 gnd.n4166 gnd.n1990 19.3944
R7139 gnd.n4166 gnd.n1988 19.3944
R7140 gnd.n4170 gnd.n1988 19.3944
R7141 gnd.n4170 gnd.n1986 19.3944
R7142 gnd.n4174 gnd.n1986 19.3944
R7143 gnd.n4174 gnd.n1984 19.3944
R7144 gnd.n4183 gnd.n1984 19.3944
R7145 gnd.n4183 gnd.n4182 19.3944
R7146 gnd.n4182 gnd.n4181 19.3944
R7147 gnd.n4181 gnd.n1845 19.3944
R7148 gnd.n4236 gnd.n1845 19.3944
R7149 gnd.n4236 gnd.n1843 19.3944
R7150 gnd.n4249 gnd.n1843 19.3944
R7151 gnd.n4249 gnd.n4248 19.3944
R7152 gnd.n4248 gnd.n4247 19.3944
R7153 gnd.n4247 gnd.n4244 19.3944
R7154 gnd.n4244 gnd.n1215 19.3944
R7155 gnd.n5330 gnd.n1215 19.3944
R7156 gnd.n5330 gnd.n5329 19.3944
R7157 gnd.n5329 gnd.n5328 19.3944
R7158 gnd.n5328 gnd.n1219 19.3944
R7159 gnd.n1315 gnd.n1219 19.3944
R7160 gnd.n5311 gnd.n1315 19.3944
R7161 gnd.n5311 gnd.n5310 19.3944
R7162 gnd.n5310 gnd.n5309 19.3944
R7163 gnd.n5309 gnd.n1321 19.3944
R7164 gnd.n4432 gnd.n1321 19.3944
R7165 gnd.n4436 gnd.n4432 19.3944
R7166 gnd.n4436 gnd.n1803 19.3944
R7167 gnd.n4461 gnd.n1803 19.3944
R7168 gnd.n4461 gnd.n1801 19.3944
R7169 gnd.n4476 gnd.n1801 19.3944
R7170 gnd.n4476 gnd.n4475 19.3944
R7171 gnd.n4475 gnd.n4474 19.3944
R7172 gnd.n4474 gnd.n4467 19.3944
R7173 gnd.n4470 gnd.n4467 19.3944
R7174 gnd.n4470 gnd.n1765 19.3944
R7175 gnd.n4519 gnd.n1765 19.3944
R7176 gnd.n4519 gnd.n1763 19.3944
R7177 gnd.n4523 gnd.n1763 19.3944
R7178 gnd.n4523 gnd.n1747 19.3944
R7179 gnd.n4545 gnd.n1747 19.3944
R7180 gnd.n4545 gnd.n1745 19.3944
R7181 gnd.n4551 gnd.n1745 19.3944
R7182 gnd.n4551 gnd.n4550 19.3944
R7183 gnd.n4550 gnd.n1723 19.3944
R7184 gnd.n4584 gnd.n1723 19.3944
R7185 gnd.n4584 gnd.n1721 19.3944
R7186 gnd.n4599 gnd.n1721 19.3944
R7187 gnd.n4599 gnd.n4598 19.3944
R7188 gnd.n4598 gnd.n4597 19.3944
R7189 gnd.n4597 gnd.n4590 19.3944
R7190 gnd.n4593 gnd.n4590 19.3944
R7191 gnd.n4593 gnd.n1684 19.3944
R7192 gnd.n4642 gnd.n1684 19.3944
R7193 gnd.n4642 gnd.n1682 19.3944
R7194 gnd.n4646 gnd.n1682 19.3944
R7195 gnd.n4646 gnd.n1665 19.3944
R7196 gnd.n4667 gnd.n1665 19.3944
R7197 gnd.n4667 gnd.n1663 19.3944
R7198 gnd.n4673 gnd.n1663 19.3944
R7199 gnd.n4673 gnd.n4672 19.3944
R7200 gnd.n4672 gnd.n1640 19.3944
R7201 gnd.n4706 gnd.n1640 19.3944
R7202 gnd.n4706 gnd.n1638 19.3944
R7203 gnd.n4710 gnd.n1638 19.3944
R7204 gnd.n4710 gnd.n1617 19.3944
R7205 gnd.n4752 gnd.n1617 19.3944
R7206 gnd.n4752 gnd.n1615 19.3944
R7207 gnd.n4758 gnd.n1615 19.3944
R7208 gnd.n4758 gnd.n4757 19.3944
R7209 gnd.n4757 gnd.n1596 19.3944
R7210 gnd.n4807 gnd.n1596 19.3944
R7211 gnd.n4807 gnd.n1594 19.3944
R7212 gnd.n4813 gnd.n1594 19.3944
R7213 gnd.n4813 gnd.n4812 19.3944
R7214 gnd.n4812 gnd.n1569 19.3944
R7215 gnd.n4844 gnd.n1569 19.3944
R7216 gnd.n4844 gnd.n1567 19.3944
R7217 gnd.n4848 gnd.n1567 19.3944
R7218 gnd.n4848 gnd.n1551 19.3944
R7219 gnd.n4870 gnd.n1551 19.3944
R7220 gnd.n4870 gnd.n1549 19.3944
R7221 gnd.n4876 gnd.n1549 19.3944
R7222 gnd.n4876 gnd.n4875 19.3944
R7223 gnd.n4875 gnd.n1523 19.3944
R7224 gnd.n4923 gnd.n1523 19.3944
R7225 gnd.n4923 gnd.n1521 19.3944
R7226 gnd.n4927 gnd.n1521 19.3944
R7227 gnd.n4927 gnd.n1431 19.3944
R7228 gnd.n5066 gnd.n1431 19.3944
R7229 gnd.n5066 gnd.n1429 19.3944
R7230 gnd.n5187 gnd.n1429 19.3944
R7231 gnd.n5187 gnd.n5186 19.3944
R7232 gnd.n5186 gnd.n5185 19.3944
R7233 gnd.n5185 gnd.n5184 19.3944
R7234 gnd.n5184 gnd.n5073 19.3944
R7235 gnd.n5111 gnd.n5073 19.3944
R7236 gnd.n5115 gnd.n5111 19.3944
R7237 gnd.n5115 gnd.n5110 19.3944
R7238 gnd.n5119 gnd.n5110 19.3944
R7239 gnd.n5119 gnd.n5108 19.3944
R7240 gnd.n5147 gnd.n5108 19.3944
R7241 gnd.n5147 gnd.n5146 19.3944
R7242 gnd.n5146 gnd.n5145 19.3944
R7243 gnd.n5145 gnd.n5125 19.3944
R7244 gnd.n5141 gnd.n5125 19.3944
R7245 gnd.n5141 gnd.n5140 19.3944
R7246 gnd.n5140 gnd.n5139 19.3944
R7247 gnd.n5139 gnd.n5131 19.3944
R7248 gnd.n5135 gnd.n5131 19.3944
R7249 gnd.n5135 gnd.n505 19.3944
R7250 gnd.n6214 gnd.n505 19.3944
R7251 gnd.n6214 gnd.n6213 19.3944
R7252 gnd.n6213 gnd.n6212 19.3944
R7253 gnd.n6212 gnd.n509 19.3944
R7254 gnd.n6208 gnd.n509 19.3944
R7255 gnd.n6208 gnd.n6207 19.3944
R7256 gnd.n5989 gnd.n633 19.3944
R7257 gnd.n5995 gnd.n633 19.3944
R7258 gnd.n5995 gnd.n631 19.3944
R7259 gnd.n5999 gnd.n631 19.3944
R7260 gnd.n5999 gnd.n627 19.3944
R7261 gnd.n6005 gnd.n627 19.3944
R7262 gnd.n6005 gnd.n625 19.3944
R7263 gnd.n6009 gnd.n625 19.3944
R7264 gnd.n6009 gnd.n621 19.3944
R7265 gnd.n6015 gnd.n621 19.3944
R7266 gnd.n6015 gnd.n619 19.3944
R7267 gnd.n6019 gnd.n619 19.3944
R7268 gnd.n6019 gnd.n615 19.3944
R7269 gnd.n6025 gnd.n615 19.3944
R7270 gnd.n6025 gnd.n613 19.3944
R7271 gnd.n6029 gnd.n613 19.3944
R7272 gnd.n6029 gnd.n609 19.3944
R7273 gnd.n6035 gnd.n609 19.3944
R7274 gnd.n6035 gnd.n607 19.3944
R7275 gnd.n6039 gnd.n607 19.3944
R7276 gnd.n6039 gnd.n603 19.3944
R7277 gnd.n6045 gnd.n603 19.3944
R7278 gnd.n6045 gnd.n601 19.3944
R7279 gnd.n6049 gnd.n601 19.3944
R7280 gnd.n6049 gnd.n597 19.3944
R7281 gnd.n6055 gnd.n597 19.3944
R7282 gnd.n6055 gnd.n595 19.3944
R7283 gnd.n6059 gnd.n595 19.3944
R7284 gnd.n6059 gnd.n591 19.3944
R7285 gnd.n6065 gnd.n591 19.3944
R7286 gnd.n6065 gnd.n589 19.3944
R7287 gnd.n6069 gnd.n589 19.3944
R7288 gnd.n6069 gnd.n585 19.3944
R7289 gnd.n6075 gnd.n585 19.3944
R7290 gnd.n6075 gnd.n583 19.3944
R7291 gnd.n6079 gnd.n583 19.3944
R7292 gnd.n6079 gnd.n579 19.3944
R7293 gnd.n6085 gnd.n579 19.3944
R7294 gnd.n6085 gnd.n577 19.3944
R7295 gnd.n6089 gnd.n577 19.3944
R7296 gnd.n6089 gnd.n573 19.3944
R7297 gnd.n6095 gnd.n573 19.3944
R7298 gnd.n6095 gnd.n571 19.3944
R7299 gnd.n6099 gnd.n571 19.3944
R7300 gnd.n6099 gnd.n567 19.3944
R7301 gnd.n6105 gnd.n567 19.3944
R7302 gnd.n6105 gnd.n565 19.3944
R7303 gnd.n6109 gnd.n565 19.3944
R7304 gnd.n6109 gnd.n561 19.3944
R7305 gnd.n6115 gnd.n561 19.3944
R7306 gnd.n6115 gnd.n559 19.3944
R7307 gnd.n6119 gnd.n559 19.3944
R7308 gnd.n6119 gnd.n555 19.3944
R7309 gnd.n6125 gnd.n555 19.3944
R7310 gnd.n6125 gnd.n553 19.3944
R7311 gnd.n6129 gnd.n553 19.3944
R7312 gnd.n6129 gnd.n549 19.3944
R7313 gnd.n6135 gnd.n549 19.3944
R7314 gnd.n6135 gnd.n547 19.3944
R7315 gnd.n6139 gnd.n547 19.3944
R7316 gnd.n6139 gnd.n543 19.3944
R7317 gnd.n6145 gnd.n543 19.3944
R7318 gnd.n6145 gnd.n541 19.3944
R7319 gnd.n6149 gnd.n541 19.3944
R7320 gnd.n6149 gnd.n537 19.3944
R7321 gnd.n6155 gnd.n537 19.3944
R7322 gnd.n6155 gnd.n535 19.3944
R7323 gnd.n6159 gnd.n535 19.3944
R7324 gnd.n6159 gnd.n531 19.3944
R7325 gnd.n6165 gnd.n531 19.3944
R7326 gnd.n6165 gnd.n529 19.3944
R7327 gnd.n6169 gnd.n529 19.3944
R7328 gnd.n6169 gnd.n525 19.3944
R7329 gnd.n6175 gnd.n525 19.3944
R7330 gnd.n6175 gnd.n523 19.3944
R7331 gnd.n6179 gnd.n523 19.3944
R7332 gnd.n6179 gnd.n519 19.3944
R7333 gnd.n6185 gnd.n519 19.3944
R7334 gnd.n6185 gnd.n517 19.3944
R7335 gnd.n6189 gnd.n517 19.3944
R7336 gnd.n6189 gnd.n513 19.3944
R7337 gnd.n6196 gnd.n513 19.3944
R7338 gnd.n6196 gnd.n511 19.3944
R7339 gnd.n6200 gnd.n511 19.3944
R7340 gnd.n5668 gnd.n828 19.3944
R7341 gnd.n5668 gnd.n824 19.3944
R7342 gnd.n5674 gnd.n824 19.3944
R7343 gnd.n5674 gnd.n822 19.3944
R7344 gnd.n5678 gnd.n822 19.3944
R7345 gnd.n5678 gnd.n818 19.3944
R7346 gnd.n5684 gnd.n818 19.3944
R7347 gnd.n5684 gnd.n816 19.3944
R7348 gnd.n5688 gnd.n816 19.3944
R7349 gnd.n5688 gnd.n812 19.3944
R7350 gnd.n5694 gnd.n812 19.3944
R7351 gnd.n5694 gnd.n810 19.3944
R7352 gnd.n5698 gnd.n810 19.3944
R7353 gnd.n5698 gnd.n806 19.3944
R7354 gnd.n5704 gnd.n806 19.3944
R7355 gnd.n5704 gnd.n804 19.3944
R7356 gnd.n5708 gnd.n804 19.3944
R7357 gnd.n5708 gnd.n800 19.3944
R7358 gnd.n5714 gnd.n800 19.3944
R7359 gnd.n5714 gnd.n798 19.3944
R7360 gnd.n5718 gnd.n798 19.3944
R7361 gnd.n5718 gnd.n794 19.3944
R7362 gnd.n5724 gnd.n794 19.3944
R7363 gnd.n5724 gnd.n792 19.3944
R7364 gnd.n5728 gnd.n792 19.3944
R7365 gnd.n5728 gnd.n788 19.3944
R7366 gnd.n5734 gnd.n788 19.3944
R7367 gnd.n5734 gnd.n786 19.3944
R7368 gnd.n5738 gnd.n786 19.3944
R7369 gnd.n5738 gnd.n782 19.3944
R7370 gnd.n5744 gnd.n782 19.3944
R7371 gnd.n5744 gnd.n780 19.3944
R7372 gnd.n5748 gnd.n780 19.3944
R7373 gnd.n5748 gnd.n776 19.3944
R7374 gnd.n5754 gnd.n776 19.3944
R7375 gnd.n5754 gnd.n774 19.3944
R7376 gnd.n5758 gnd.n774 19.3944
R7377 gnd.n5758 gnd.n770 19.3944
R7378 gnd.n5764 gnd.n770 19.3944
R7379 gnd.n5764 gnd.n768 19.3944
R7380 gnd.n5768 gnd.n768 19.3944
R7381 gnd.n5768 gnd.n764 19.3944
R7382 gnd.n5774 gnd.n764 19.3944
R7383 gnd.n5774 gnd.n762 19.3944
R7384 gnd.n5778 gnd.n762 19.3944
R7385 gnd.n5778 gnd.n758 19.3944
R7386 gnd.n5784 gnd.n758 19.3944
R7387 gnd.n5784 gnd.n756 19.3944
R7388 gnd.n5788 gnd.n756 19.3944
R7389 gnd.n5788 gnd.n752 19.3944
R7390 gnd.n5794 gnd.n752 19.3944
R7391 gnd.n5794 gnd.n750 19.3944
R7392 gnd.n5798 gnd.n750 19.3944
R7393 gnd.n5798 gnd.n746 19.3944
R7394 gnd.n5804 gnd.n746 19.3944
R7395 gnd.n5804 gnd.n744 19.3944
R7396 gnd.n5808 gnd.n744 19.3944
R7397 gnd.n5808 gnd.n740 19.3944
R7398 gnd.n5814 gnd.n740 19.3944
R7399 gnd.n5814 gnd.n738 19.3944
R7400 gnd.n5818 gnd.n738 19.3944
R7401 gnd.n5818 gnd.n734 19.3944
R7402 gnd.n5824 gnd.n734 19.3944
R7403 gnd.n5824 gnd.n732 19.3944
R7404 gnd.n5828 gnd.n732 19.3944
R7405 gnd.n5828 gnd.n728 19.3944
R7406 gnd.n5834 gnd.n728 19.3944
R7407 gnd.n5834 gnd.n726 19.3944
R7408 gnd.n5838 gnd.n726 19.3944
R7409 gnd.n5838 gnd.n722 19.3944
R7410 gnd.n5844 gnd.n722 19.3944
R7411 gnd.n5844 gnd.n720 19.3944
R7412 gnd.n5848 gnd.n720 19.3944
R7413 gnd.n5848 gnd.n716 19.3944
R7414 gnd.n5854 gnd.n716 19.3944
R7415 gnd.n5854 gnd.n714 19.3944
R7416 gnd.n5858 gnd.n714 19.3944
R7417 gnd.n5858 gnd.n710 19.3944
R7418 gnd.n5864 gnd.n710 19.3944
R7419 gnd.n5864 gnd.n708 19.3944
R7420 gnd.n5868 gnd.n708 19.3944
R7421 gnd.n5868 gnd.n704 19.3944
R7422 gnd.n5874 gnd.n704 19.3944
R7423 gnd.n5874 gnd.n702 19.3944
R7424 gnd.n5878 gnd.n702 19.3944
R7425 gnd.n5878 gnd.n698 19.3944
R7426 gnd.n5884 gnd.n698 19.3944
R7427 gnd.n5884 gnd.n696 19.3944
R7428 gnd.n5888 gnd.n696 19.3944
R7429 gnd.n5888 gnd.n692 19.3944
R7430 gnd.n5894 gnd.n692 19.3944
R7431 gnd.n5894 gnd.n690 19.3944
R7432 gnd.n5898 gnd.n690 19.3944
R7433 gnd.n5898 gnd.n686 19.3944
R7434 gnd.n5904 gnd.n686 19.3944
R7435 gnd.n5904 gnd.n684 19.3944
R7436 gnd.n5908 gnd.n684 19.3944
R7437 gnd.n5908 gnd.n680 19.3944
R7438 gnd.n5914 gnd.n680 19.3944
R7439 gnd.n5914 gnd.n678 19.3944
R7440 gnd.n5918 gnd.n678 19.3944
R7441 gnd.n5918 gnd.n674 19.3944
R7442 gnd.n5924 gnd.n674 19.3944
R7443 gnd.n5924 gnd.n672 19.3944
R7444 gnd.n5928 gnd.n672 19.3944
R7445 gnd.n5928 gnd.n668 19.3944
R7446 gnd.n5934 gnd.n668 19.3944
R7447 gnd.n5934 gnd.n666 19.3944
R7448 gnd.n5938 gnd.n666 19.3944
R7449 gnd.n5938 gnd.n662 19.3944
R7450 gnd.n5944 gnd.n662 19.3944
R7451 gnd.n5944 gnd.n660 19.3944
R7452 gnd.n5948 gnd.n660 19.3944
R7453 gnd.n5948 gnd.n656 19.3944
R7454 gnd.n5954 gnd.n656 19.3944
R7455 gnd.n5954 gnd.n654 19.3944
R7456 gnd.n5958 gnd.n654 19.3944
R7457 gnd.n5958 gnd.n650 19.3944
R7458 gnd.n5964 gnd.n650 19.3944
R7459 gnd.n5964 gnd.n648 19.3944
R7460 gnd.n5968 gnd.n648 19.3944
R7461 gnd.n5968 gnd.n644 19.3944
R7462 gnd.n5974 gnd.n644 19.3944
R7463 gnd.n5974 gnd.n642 19.3944
R7464 gnd.n5979 gnd.n642 19.3944
R7465 gnd.n5979 gnd.n638 19.3944
R7466 gnd.n5985 gnd.n638 19.3944
R7467 gnd.n5986 gnd.n5985 19.3944
R7468 gnd.n6387 gnd.n419 19.3944
R7469 gnd.n6387 gnd.n6386 19.3944
R7470 gnd.n6386 gnd.n6385 19.3944
R7471 gnd.n6385 gnd.n6383 19.3944
R7472 gnd.n6383 gnd.n6380 19.3944
R7473 gnd.n6380 gnd.n6379 19.3944
R7474 gnd.n6379 gnd.n6376 19.3944
R7475 gnd.n6376 gnd.n6375 19.3944
R7476 gnd.n6375 gnd.n6372 19.3944
R7477 gnd.n6372 gnd.n6371 19.3944
R7478 gnd.n6371 gnd.n6368 19.3944
R7479 gnd.n6368 gnd.n6367 19.3944
R7480 gnd.n6367 gnd.n6364 19.3944
R7481 gnd.n6364 gnd.n6363 19.3944
R7482 gnd.n6363 gnd.n6360 19.3944
R7483 gnd.n6358 gnd.n6355 19.3944
R7484 gnd.n6355 gnd.n6354 19.3944
R7485 gnd.n6354 gnd.n6351 19.3944
R7486 gnd.n6351 gnd.n6350 19.3944
R7487 gnd.n6350 gnd.n6347 19.3944
R7488 gnd.n6347 gnd.n6346 19.3944
R7489 gnd.n6346 gnd.n6343 19.3944
R7490 gnd.n6343 gnd.n6342 19.3944
R7491 gnd.n6342 gnd.n6339 19.3944
R7492 gnd.n6339 gnd.n6338 19.3944
R7493 gnd.n6338 gnd.n6335 19.3944
R7494 gnd.n6335 gnd.n6334 19.3944
R7495 gnd.n6334 gnd.n6331 19.3944
R7496 gnd.n6331 gnd.n6330 19.3944
R7497 gnd.n6330 gnd.n6327 19.3944
R7498 gnd.n6327 gnd.n6326 19.3944
R7499 gnd.n6326 gnd.n6323 19.3944
R7500 gnd.n6323 gnd.n6322 19.3944
R7501 gnd.n6315 gnd.n6314 19.3944
R7502 gnd.n6314 gnd.n6313 19.3944
R7503 gnd.n6313 gnd.n6312 19.3944
R7504 gnd.n6312 gnd.n467 19.3944
R7505 gnd.n489 gnd.n467 19.3944
R7506 gnd.n489 gnd.n485 19.3944
R7507 gnd.n495 gnd.n485 19.3944
R7508 gnd.n496 gnd.n495 19.3944
R7509 gnd.n499 gnd.n496 19.3944
R7510 gnd.n499 gnd.n483 19.3944
R7511 gnd.n6219 gnd.n483 19.3944
R7512 gnd.n6220 gnd.n6219 19.3944
R7513 gnd.n6223 gnd.n6220 19.3944
R7514 gnd.n6223 gnd.n481 19.3944
R7515 gnd.n6285 gnd.n481 19.3944
R7516 gnd.n6285 gnd.n6284 19.3944
R7517 gnd.n6284 gnd.n6283 19.3944
R7518 gnd.n6283 gnd.n6282 19.3944
R7519 gnd.n6282 gnd.n6280 19.3944
R7520 gnd.n6280 gnd.n6279 19.3944
R7521 gnd.n6279 gnd.n6278 19.3944
R7522 gnd.n6278 gnd.n6276 19.3944
R7523 gnd.n6276 gnd.n6275 19.3944
R7524 gnd.n6275 gnd.n6273 19.3944
R7525 gnd.n6273 gnd.n6272 19.3944
R7526 gnd.n6272 gnd.n6270 19.3944
R7527 gnd.n6270 gnd.n6269 19.3944
R7528 gnd.n6269 gnd.n6267 19.3944
R7529 gnd.n6267 gnd.n6266 19.3944
R7530 gnd.n6266 gnd.n6264 19.3944
R7531 gnd.n6264 gnd.n6263 19.3944
R7532 gnd.n6263 gnd.n6261 19.3944
R7533 gnd.n6261 gnd.n6260 19.3944
R7534 gnd.n6260 gnd.n6258 19.3944
R7535 gnd.n6258 gnd.n6257 19.3944
R7536 gnd.n6257 gnd.n6255 19.3944
R7537 gnd.n6255 gnd.n6254 19.3944
R7538 gnd.n6254 gnd.n6252 19.3944
R7539 gnd.n6252 gnd.n6251 19.3944
R7540 gnd.n6251 gnd.n159 19.3944
R7541 gnd.n6687 gnd.n159 19.3944
R7542 gnd.n6688 gnd.n6687 19.3944
R7543 gnd.n6726 gnd.n120 19.3944
R7544 gnd.n6721 gnd.n120 19.3944
R7545 gnd.n6721 gnd.n6720 19.3944
R7546 gnd.n6720 gnd.n6719 19.3944
R7547 gnd.n6719 gnd.n127 19.3944
R7548 gnd.n6714 gnd.n127 19.3944
R7549 gnd.n6714 gnd.n6713 19.3944
R7550 gnd.n6713 gnd.n6712 19.3944
R7551 gnd.n6712 gnd.n134 19.3944
R7552 gnd.n6707 gnd.n134 19.3944
R7553 gnd.n6707 gnd.n6706 19.3944
R7554 gnd.n6706 gnd.n6705 19.3944
R7555 gnd.n6705 gnd.n141 19.3944
R7556 gnd.n6700 gnd.n141 19.3944
R7557 gnd.n6700 gnd.n6699 19.3944
R7558 gnd.n6699 gnd.n6698 19.3944
R7559 gnd.n6698 gnd.n148 19.3944
R7560 gnd.n6693 gnd.n148 19.3944
R7561 gnd.n6759 gnd.n6758 19.3944
R7562 gnd.n6758 gnd.n6757 19.3944
R7563 gnd.n6757 gnd.n92 19.3944
R7564 gnd.n6752 gnd.n92 19.3944
R7565 gnd.n6752 gnd.n6751 19.3944
R7566 gnd.n6751 gnd.n6750 19.3944
R7567 gnd.n6750 gnd.n99 19.3944
R7568 gnd.n6745 gnd.n99 19.3944
R7569 gnd.n6745 gnd.n6744 19.3944
R7570 gnd.n6744 gnd.n6743 19.3944
R7571 gnd.n6743 gnd.n106 19.3944
R7572 gnd.n6738 gnd.n106 19.3944
R7573 gnd.n6738 gnd.n6737 19.3944
R7574 gnd.n6737 gnd.n6736 19.3944
R7575 gnd.n6736 gnd.n113 19.3944
R7576 gnd.n6731 gnd.n113 19.3944
R7577 gnd.n6731 gnd.n6730 19.3944
R7578 gnd.n6447 gnd.n325 19.3944
R7579 gnd.n6451 gnd.n325 19.3944
R7580 gnd.n6451 gnd.n310 19.3944
R7581 gnd.n6463 gnd.n310 19.3944
R7582 gnd.n6463 gnd.n308 19.3944
R7583 gnd.n6467 gnd.n308 19.3944
R7584 gnd.n6467 gnd.n292 19.3944
R7585 gnd.n6479 gnd.n292 19.3944
R7586 gnd.n6479 gnd.n290 19.3944
R7587 gnd.n6483 gnd.n290 19.3944
R7588 gnd.n6483 gnd.n275 19.3944
R7589 gnd.n6495 gnd.n275 19.3944
R7590 gnd.n6495 gnd.n273 19.3944
R7591 gnd.n6500 gnd.n273 19.3944
R7592 gnd.n6500 gnd.n6499 19.3944
R7593 gnd.n6499 gnd.n259 19.3944
R7594 gnd.n6517 gnd.n6516 19.3944
R7595 gnd.n6530 gnd.n6529 19.3944
R7596 gnd.n234 gnd.n233 19.3944
R7597 gnd.n6544 gnd.n6543 19.3944
R7598 gnd.n6556 gnd.n219 19.3944
R7599 gnd.n6556 gnd.n211 19.3944
R7600 gnd.n6560 gnd.n211 19.3944
R7601 gnd.n6560 gnd.n199 19.3944
R7602 gnd.n6572 gnd.n199 19.3944
R7603 gnd.n6572 gnd.n197 19.3944
R7604 gnd.n6576 gnd.n197 19.3944
R7605 gnd.n6576 gnd.n183 19.3944
R7606 gnd.n6588 gnd.n183 19.3944
R7607 gnd.n6588 gnd.n181 19.3944
R7608 gnd.n6592 gnd.n181 19.3944
R7609 gnd.n6592 gnd.n166 19.3944
R7610 gnd.n6678 gnd.n166 19.3944
R7611 gnd.n6678 gnd.n164 19.3944
R7612 gnd.n6682 gnd.n164 19.3944
R7613 gnd.n6682 gnd.n87 19.3944
R7614 gnd.n6762 gnd.n87 19.3944
R7615 gnd.n3875 gnd.n3874 19.3944
R7616 gnd.n3874 gnd.n3873 19.3944
R7617 gnd.n3873 gnd.n3872 19.3944
R7618 gnd.n3872 gnd.n3870 19.3944
R7619 gnd.n3870 gnd.n3867 19.3944
R7620 gnd.n3867 gnd.n3866 19.3944
R7621 gnd.n3866 gnd.n3863 19.3944
R7622 gnd.n3863 gnd.n3862 19.3944
R7623 gnd.n3862 gnd.n3859 19.3944
R7624 gnd.n3859 gnd.n3858 19.3944
R7625 gnd.n3858 gnd.n3855 19.3944
R7626 gnd.n3855 gnd.n3854 19.3944
R7627 gnd.n3854 gnd.n3851 19.3944
R7628 gnd.n3851 gnd.n3850 19.3944
R7629 gnd.n3850 gnd.n3847 19.3944
R7630 gnd.n3847 gnd.n3846 19.3944
R7631 gnd.n3846 gnd.n3843 19.3944
R7632 gnd.n3841 gnd.n3838 19.3944
R7633 gnd.n3838 gnd.n3837 19.3944
R7634 gnd.n3837 gnd.n3834 19.3944
R7635 gnd.n3834 gnd.n3833 19.3944
R7636 gnd.n3833 gnd.n3830 19.3944
R7637 gnd.n3830 gnd.n3829 19.3944
R7638 gnd.n3829 gnd.n3826 19.3944
R7639 gnd.n3826 gnd.n3825 19.3944
R7640 gnd.n3825 gnd.n3822 19.3944
R7641 gnd.n3822 gnd.n3821 19.3944
R7642 gnd.n3821 gnd.n3818 19.3944
R7643 gnd.n3818 gnd.n3817 19.3944
R7644 gnd.n3817 gnd.n3814 19.3944
R7645 gnd.n3814 gnd.n3813 19.3944
R7646 gnd.n3813 gnd.n3810 19.3944
R7647 gnd.n3810 gnd.n3809 19.3944
R7648 gnd.n3809 gnd.n3806 19.3944
R7649 gnd.n3806 gnd.n3805 19.3944
R7650 gnd.n3885 gnd.n2116 19.3944
R7651 gnd.n3885 gnd.n2102 19.3944
R7652 gnd.n3897 gnd.n2102 19.3944
R7653 gnd.n3897 gnd.n2100 19.3944
R7654 gnd.n3901 gnd.n2100 19.3944
R7655 gnd.n3901 gnd.n2086 19.3944
R7656 gnd.n3913 gnd.n2086 19.3944
R7657 gnd.n3913 gnd.n2084 19.3944
R7658 gnd.n3917 gnd.n2084 19.3944
R7659 gnd.n3917 gnd.n2070 19.3944
R7660 gnd.n3929 gnd.n2070 19.3944
R7661 gnd.n3929 gnd.n2068 19.3944
R7662 gnd.n3933 gnd.n2068 19.3944
R7663 gnd.n3933 gnd.n2054 19.3944
R7664 gnd.n3946 gnd.n2054 19.3944
R7665 gnd.n3946 gnd.n2052 19.3944
R7666 gnd.n3954 gnd.n2052 19.3944
R7667 gnd.n3954 gnd.n3953 19.3944
R7668 gnd.n3953 gnd.n3952 19.3944
R7669 gnd.n3952 gnd.n2035 19.3944
R7670 gnd.n3989 gnd.n2035 19.3944
R7671 gnd.n3989 gnd.n3988 19.3944
R7672 gnd.n3988 gnd.n3987 19.3944
R7673 gnd.n3987 gnd.n3986 19.3944
R7674 gnd.n3986 gnd.n3984 19.3944
R7675 gnd.n3984 gnd.n1015 19.3944
R7676 gnd.n5485 gnd.n1015 19.3944
R7677 gnd.n5485 gnd.n5484 19.3944
R7678 gnd.n5484 gnd.n5483 19.3944
R7679 gnd.n5483 gnd.n1019 19.3944
R7680 gnd.n5473 gnd.n1019 19.3944
R7681 gnd.n5473 gnd.n5472 19.3944
R7682 gnd.n5472 gnd.n5471 19.3944
R7683 gnd.n5471 gnd.n1041 19.3944
R7684 gnd.n5461 gnd.n1041 19.3944
R7685 gnd.n5461 gnd.n5460 19.3944
R7686 gnd.n5460 gnd.n5459 19.3944
R7687 gnd.n5459 gnd.n1061 19.3944
R7688 gnd.n5449 gnd.n1061 19.3944
R7689 gnd.n5449 gnd.n5448 19.3944
R7690 gnd.n5448 gnd.n5447 19.3944
R7691 gnd.n5447 gnd.n1083 19.3944
R7692 gnd.n3881 gnd.n2118 19.3944
R7693 gnd.n3611 gnd.n2118 19.3944
R7694 gnd.n3612 gnd.n3611 19.3944
R7695 gnd.n3615 gnd.n3612 19.3944
R7696 gnd.n3615 gnd.n3607 19.3944
R7697 gnd.n3621 gnd.n3607 19.3944
R7698 gnd.n3622 gnd.n3621 19.3944
R7699 gnd.n3625 gnd.n3622 19.3944
R7700 gnd.n3625 gnd.n3605 19.3944
R7701 gnd.n3631 gnd.n3605 19.3944
R7702 gnd.n3632 gnd.n3631 19.3944
R7703 gnd.n3635 gnd.n3632 19.3944
R7704 gnd.n3635 gnd.n3603 19.3944
R7705 gnd.n3641 gnd.n3603 19.3944
R7706 gnd.n3642 gnd.n3641 19.3944
R7707 gnd.n3645 gnd.n3642 19.3944
R7708 gnd.n3702 gnd.n3701 19.3944
R7709 gnd.n3701 gnd.n3700 19.3944
R7710 gnd.n3700 gnd.n3698 19.3944
R7711 gnd.n3698 gnd.n3697 19.3944
R7712 gnd.n3697 gnd.n3695 19.3944
R7713 gnd.n3695 gnd.n3694 19.3944
R7714 gnd.n3694 gnd.n3692 19.3944
R7715 gnd.n3692 gnd.n3691 19.3944
R7716 gnd.n3691 gnd.n3689 19.3944
R7717 gnd.n3689 gnd.n3688 19.3944
R7718 gnd.n3688 gnd.n3686 19.3944
R7719 gnd.n3686 gnd.n3685 19.3944
R7720 gnd.n3685 gnd.n3683 19.3944
R7721 gnd.n3683 gnd.n3682 19.3944
R7722 gnd.n3682 gnd.n3680 19.3944
R7723 gnd.n3680 gnd.n3679 19.3944
R7724 gnd.n3679 gnd.n3677 19.3944
R7725 gnd.n3677 gnd.n3676 19.3944
R7726 gnd.n3676 gnd.n3674 19.3944
R7727 gnd.n3674 gnd.n3673 19.3944
R7728 gnd.n3673 gnd.n3671 19.3944
R7729 gnd.n3671 gnd.n3668 19.3944
R7730 gnd.n3668 gnd.n2022 19.3944
R7731 gnd.n4002 gnd.n2022 19.3944
R7732 gnd.n4002 gnd.n2020 19.3944
R7733 gnd.n4006 gnd.n2020 19.3944
R7734 gnd.n4006 gnd.n2013 19.3944
R7735 gnd.n4028 gnd.n2013 19.3944
R7736 gnd.n4028 gnd.n2014 19.3944
R7737 gnd.n4024 gnd.n2014 19.3944
R7738 gnd.n4024 gnd.n2005 19.3944
R7739 gnd.n4059 gnd.n2005 19.3944
R7740 gnd.n4059 gnd.n2003 19.3944
R7741 gnd.n4063 gnd.n2003 19.3944
R7742 gnd.n4063 gnd.n1993 19.3944
R7743 gnd.n4160 gnd.n1993 19.3944
R7744 gnd.n4160 gnd.n1994 19.3944
R7745 gnd.n4156 gnd.n1994 19.3944
R7746 gnd.n4156 gnd.n4155 19.3944
R7747 gnd.n4155 gnd.n4154 19.3944
R7748 gnd.n4154 gnd.n4151 19.3944
R7749 gnd.n4151 gnd.n1980 19.3944
R7750 gnd.n3798 gnd.n3797 19.3944
R7751 gnd.n3797 gnd.n3754 19.3944
R7752 gnd.n3793 gnd.n3754 19.3944
R7753 gnd.n3793 gnd.n3792 19.3944
R7754 gnd.n3792 gnd.n3790 19.3944
R7755 gnd.n3790 gnd.n3789 19.3944
R7756 gnd.n3789 gnd.n3787 19.3944
R7757 gnd.n3787 gnd.n3786 19.3944
R7758 gnd.n3786 gnd.n3784 19.3944
R7759 gnd.n3784 gnd.n3783 19.3944
R7760 gnd.n3783 gnd.n3781 19.3944
R7761 gnd.n3781 gnd.n3780 19.3944
R7762 gnd.n3780 gnd.n3778 19.3944
R7763 gnd.n3778 gnd.n3777 19.3944
R7764 gnd.n3777 gnd.n3775 19.3944
R7765 gnd.n3775 gnd.n3774 19.3944
R7766 gnd.n3774 gnd.n3772 19.3944
R7767 gnd.n3772 gnd.n3771 19.3944
R7768 gnd.n3771 gnd.n2039 19.3944
R7769 gnd.n3967 gnd.n2039 19.3944
R7770 gnd.n3976 gnd.n3967 19.3944
R7771 gnd.n3976 gnd.n3975 19.3944
R7772 gnd.n3975 gnd.n3973 19.3944
R7773 gnd.n3973 gnd.n3972 19.3944
R7774 gnd.n3972 gnd.n2018 19.3944
R7775 gnd.n4010 gnd.n2018 19.3944
R7776 gnd.n4011 gnd.n4010 19.3944
R7777 gnd.n4012 gnd.n4011 19.3944
R7778 gnd.n4012 gnd.n2016 19.3944
R7779 gnd.n4020 gnd.n2016 19.3944
R7780 gnd.n4020 gnd.n4019 19.3944
R7781 gnd.n4019 gnd.n4018 19.3944
R7782 gnd.n4018 gnd.n2002 19.3944
R7783 gnd.n4067 gnd.n2002 19.3944
R7784 gnd.n4067 gnd.n2000 19.3944
R7785 gnd.n4071 gnd.n2000 19.3944
R7786 gnd.n4072 gnd.n4071 19.3944
R7787 gnd.n4075 gnd.n4072 19.3944
R7788 gnd.n4075 gnd.n1998 19.3944
R7789 gnd.n4147 gnd.n1998 19.3944
R7790 gnd.n4147 gnd.n4146 19.3944
R7791 gnd.n4146 gnd.n4145 19.3944
R7792 gnd.n4094 gnd.n1140 19.3944
R7793 gnd.n4098 gnd.n4094 19.3944
R7794 gnd.n4101 gnd.n4098 19.3944
R7795 gnd.n4104 gnd.n4101 19.3944
R7796 gnd.n4104 gnd.n4090 19.3944
R7797 gnd.n4108 gnd.n4090 19.3944
R7798 gnd.n4111 gnd.n4108 19.3944
R7799 gnd.n4114 gnd.n4111 19.3944
R7800 gnd.n4114 gnd.n4088 19.3944
R7801 gnd.n4118 gnd.n4088 19.3944
R7802 gnd.n4121 gnd.n4118 19.3944
R7803 gnd.n4124 gnd.n4121 19.3944
R7804 gnd.n4124 gnd.n4086 19.3944
R7805 gnd.n4128 gnd.n4086 19.3944
R7806 gnd.n4131 gnd.n4128 19.3944
R7807 gnd.n4134 gnd.n4131 19.3944
R7808 gnd.n4134 gnd.n4084 19.3944
R7809 gnd.n4139 gnd.n4084 19.3944
R7810 gnd.n5439 gnd.n1093 19.3944
R7811 gnd.n5434 gnd.n1093 19.3944
R7812 gnd.n5434 gnd.n5433 19.3944
R7813 gnd.n5433 gnd.n5432 19.3944
R7814 gnd.n5432 gnd.n5429 19.3944
R7815 gnd.n5429 gnd.n5428 19.3944
R7816 gnd.n5428 gnd.n5425 19.3944
R7817 gnd.n5425 gnd.n5424 19.3944
R7818 gnd.n5424 gnd.n5421 19.3944
R7819 gnd.n5421 gnd.n5420 19.3944
R7820 gnd.n5420 gnd.n5417 19.3944
R7821 gnd.n5417 gnd.n5416 19.3944
R7822 gnd.n5416 gnd.n5413 19.3944
R7823 gnd.n5413 gnd.n5412 19.3944
R7824 gnd.n5412 gnd.n5409 19.3944
R7825 gnd.n3889 gnd.n2110 19.3944
R7826 gnd.n3889 gnd.n2108 19.3944
R7827 gnd.n3893 gnd.n2108 19.3944
R7828 gnd.n3893 gnd.n2093 19.3944
R7829 gnd.n3905 gnd.n2093 19.3944
R7830 gnd.n3905 gnd.n2091 19.3944
R7831 gnd.n3909 gnd.n2091 19.3944
R7832 gnd.n3909 gnd.n2078 19.3944
R7833 gnd.n3921 gnd.n2078 19.3944
R7834 gnd.n3921 gnd.n2076 19.3944
R7835 gnd.n3925 gnd.n2076 19.3944
R7836 gnd.n3925 gnd.n2061 19.3944
R7837 gnd.n3937 gnd.n2061 19.3944
R7838 gnd.n3937 gnd.n2059 19.3944
R7839 gnd.n3942 gnd.n2059 19.3944
R7840 gnd.n3942 gnd.n3941 19.3944
R7841 gnd.n3959 gnd.n3958 19.3944
R7842 gnd.n3962 gnd.n3961 19.3944
R7843 gnd.n3994 gnd.n3993 19.3944
R7844 gnd.n3997 gnd.n3996 19.3944
R7845 gnd.n5491 gnd.n5490 19.3944
R7846 gnd.n5490 gnd.n5489 19.3944
R7847 gnd.n5489 gnd.n1008 19.3944
R7848 gnd.n5479 gnd.n1008 19.3944
R7849 gnd.n5479 gnd.n5478 19.3944
R7850 gnd.n5478 gnd.n5477 19.3944
R7851 gnd.n5477 gnd.n1030 19.3944
R7852 gnd.n5467 gnd.n1030 19.3944
R7853 gnd.n5467 gnd.n5466 19.3944
R7854 gnd.n5466 gnd.n5465 19.3944
R7855 gnd.n5465 gnd.n1051 19.3944
R7856 gnd.n5455 gnd.n1051 19.3944
R7857 gnd.n5455 gnd.n5454 19.3944
R7858 gnd.n5454 gnd.n5453 19.3944
R7859 gnd.n5453 gnd.n1072 19.3944
R7860 gnd.n5443 gnd.n1072 19.3944
R7861 gnd.n5443 gnd.n5442 19.3944
R7862 gnd.n5664 gnd.n830 19.3944
R7863 gnd.n5658 gnd.n830 19.3944
R7864 gnd.n5658 gnd.n5657 19.3944
R7865 gnd.n5657 gnd.n5656 19.3944
R7866 gnd.n5656 gnd.n837 19.3944
R7867 gnd.n5650 gnd.n837 19.3944
R7868 gnd.n5650 gnd.n5649 19.3944
R7869 gnd.n5649 gnd.n5648 19.3944
R7870 gnd.n5648 gnd.n845 19.3944
R7871 gnd.n5642 gnd.n845 19.3944
R7872 gnd.n5642 gnd.n5641 19.3944
R7873 gnd.n5641 gnd.n5640 19.3944
R7874 gnd.n5640 gnd.n853 19.3944
R7875 gnd.n5634 gnd.n853 19.3944
R7876 gnd.n5634 gnd.n5633 19.3944
R7877 gnd.n5633 gnd.n5632 19.3944
R7878 gnd.n5632 gnd.n861 19.3944
R7879 gnd.n5626 gnd.n861 19.3944
R7880 gnd.n5626 gnd.n5625 19.3944
R7881 gnd.n5625 gnd.n5624 19.3944
R7882 gnd.n5624 gnd.n869 19.3944
R7883 gnd.n5618 gnd.n869 19.3944
R7884 gnd.n5618 gnd.n5617 19.3944
R7885 gnd.n5617 gnd.n5616 19.3944
R7886 gnd.n5616 gnd.n877 19.3944
R7887 gnd.n5610 gnd.n877 19.3944
R7888 gnd.n5610 gnd.n5609 19.3944
R7889 gnd.n5609 gnd.n5608 19.3944
R7890 gnd.n5608 gnd.n885 19.3944
R7891 gnd.n5602 gnd.n885 19.3944
R7892 gnd.n5602 gnd.n5601 19.3944
R7893 gnd.n5601 gnd.n5600 19.3944
R7894 gnd.n5600 gnd.n893 19.3944
R7895 gnd.n5594 gnd.n893 19.3944
R7896 gnd.n5594 gnd.n5593 19.3944
R7897 gnd.n5593 gnd.n5592 19.3944
R7898 gnd.n5592 gnd.n901 19.3944
R7899 gnd.n5586 gnd.n901 19.3944
R7900 gnd.n5586 gnd.n5585 19.3944
R7901 gnd.n5585 gnd.n5584 19.3944
R7902 gnd.n5584 gnd.n909 19.3944
R7903 gnd.n5578 gnd.n909 19.3944
R7904 gnd.n5578 gnd.n5577 19.3944
R7905 gnd.n5577 gnd.n5576 19.3944
R7906 gnd.n5576 gnd.n917 19.3944
R7907 gnd.n5570 gnd.n917 19.3944
R7908 gnd.n5570 gnd.n5569 19.3944
R7909 gnd.n5569 gnd.n5568 19.3944
R7910 gnd.n5568 gnd.n925 19.3944
R7911 gnd.n5562 gnd.n925 19.3944
R7912 gnd.n5562 gnd.n5561 19.3944
R7913 gnd.n5561 gnd.n5560 19.3944
R7914 gnd.n5560 gnd.n933 19.3944
R7915 gnd.n5554 gnd.n933 19.3944
R7916 gnd.n5554 gnd.n5553 19.3944
R7917 gnd.n5553 gnd.n5552 19.3944
R7918 gnd.n5552 gnd.n941 19.3944
R7919 gnd.n5546 gnd.n941 19.3944
R7920 gnd.n5546 gnd.n5545 19.3944
R7921 gnd.n5545 gnd.n5544 19.3944
R7922 gnd.n5544 gnd.n949 19.3944
R7923 gnd.n5538 gnd.n949 19.3944
R7924 gnd.n5538 gnd.n5537 19.3944
R7925 gnd.n5537 gnd.n5536 19.3944
R7926 gnd.n5536 gnd.n957 19.3944
R7927 gnd.n5530 gnd.n957 19.3944
R7928 gnd.n5530 gnd.n5529 19.3944
R7929 gnd.n5529 gnd.n5528 19.3944
R7930 gnd.n5528 gnd.n965 19.3944
R7931 gnd.n5522 gnd.n965 19.3944
R7932 gnd.n5522 gnd.n5521 19.3944
R7933 gnd.n5521 gnd.n5520 19.3944
R7934 gnd.n5520 gnd.n973 19.3944
R7935 gnd.n5514 gnd.n973 19.3944
R7936 gnd.n5514 gnd.n5513 19.3944
R7937 gnd.n5513 gnd.n5512 19.3944
R7938 gnd.n5512 gnd.n981 19.3944
R7939 gnd.n5506 gnd.n981 19.3944
R7940 gnd.n5506 gnd.n5505 19.3944
R7941 gnd.n5505 gnd.n5504 19.3944
R7942 gnd.n5504 gnd.n989 19.3944
R7943 gnd.n5498 gnd.n989 19.3944
R7944 gnd.n5498 gnd.n5497 19.3944
R7945 gnd.n5497 gnd.n5496 19.3944
R7946 gnd.n4253 gnd.n1835 19.3944
R7947 gnd.n4257 gnd.n1835 19.3944
R7948 gnd.n4257 gnd.n1833 19.3944
R7949 gnd.n4261 gnd.n1833 19.3944
R7950 gnd.n4261 gnd.n1831 19.3944
R7951 gnd.n4265 gnd.n1831 19.3944
R7952 gnd.n4265 gnd.n1824 19.3944
R7953 gnd.n4286 gnd.n1824 19.3944
R7954 gnd.n4286 gnd.n1822 19.3944
R7955 gnd.n4290 gnd.n1822 19.3944
R7956 gnd.n4321 gnd.n4290 19.3944
R7957 gnd.n4322 gnd.n4321 19.3944
R7958 gnd.n4322 gnd.n1819 19.3944
R7959 gnd.n4428 gnd.n1819 19.3944
R7960 gnd.n4428 gnd.n1820 19.3944
R7961 gnd.n4424 gnd.n1820 19.3944
R7962 gnd.n4424 gnd.n4423 19.3944
R7963 gnd.n4423 gnd.n4422 19.3944
R7964 gnd.n4422 gnd.n4327 19.3944
R7965 gnd.n4418 gnd.n4327 19.3944
R7966 gnd.n4418 gnd.n4417 19.3944
R7967 gnd.n4417 gnd.n4416 19.3944
R7968 gnd.n4416 gnd.n4333 19.3944
R7969 gnd.n4412 gnd.n4333 19.3944
R7970 gnd.n4412 gnd.n4411 19.3944
R7971 gnd.n4411 gnd.n4410 19.3944
R7972 gnd.n4410 gnd.n4336 19.3944
R7973 gnd.n4406 gnd.n4336 19.3944
R7974 gnd.n4406 gnd.n4405 19.3944
R7975 gnd.n4405 gnd.n4404 19.3944
R7976 gnd.n4404 gnd.n4340 19.3944
R7977 gnd.n4400 gnd.n4340 19.3944
R7978 gnd.n4400 gnd.n4399 19.3944
R7979 gnd.n4399 gnd.n4398 19.3944
R7980 gnd.n4398 gnd.n4344 19.3944
R7981 gnd.n4394 gnd.n4344 19.3944
R7982 gnd.n4394 gnd.n4393 19.3944
R7983 gnd.n4393 gnd.n4392 19.3944
R7984 gnd.n4392 gnd.n4348 19.3944
R7985 gnd.n4388 gnd.n4348 19.3944
R7986 gnd.n4388 gnd.n4387 19.3944
R7987 gnd.n4387 gnd.n4386 19.3944
R7988 gnd.n4386 gnd.n4353 19.3944
R7989 gnd.n4382 gnd.n4353 19.3944
R7990 gnd.n4382 gnd.n4381 19.3944
R7991 gnd.n4381 gnd.n4380 19.3944
R7992 gnd.n4380 gnd.n4357 19.3944
R7993 gnd.n4376 gnd.n4357 19.3944
R7994 gnd.n4376 gnd.n4375 19.3944
R7995 gnd.n4375 gnd.n4374 19.3944
R7996 gnd.n4374 gnd.n4360 19.3944
R7997 gnd.n4370 gnd.n4360 19.3944
R7998 gnd.n4370 gnd.n4369 19.3944
R7999 gnd.n4369 gnd.n4368 19.3944
R8000 gnd.n4368 gnd.n4365 19.3944
R8001 gnd.n4365 gnd.n1609 19.3944
R8002 gnd.n4762 gnd.n1609 19.3944
R8003 gnd.n4762 gnd.n1606 19.3944
R8004 gnd.n4795 gnd.n1606 19.3944
R8005 gnd.n4795 gnd.n1607 19.3944
R8006 gnd.n4791 gnd.n1607 19.3944
R8007 gnd.n4791 gnd.n4790 19.3944
R8008 gnd.n4790 gnd.n4789 19.3944
R8009 gnd.n4789 gnd.n4769 19.3944
R8010 gnd.n4785 gnd.n4769 19.3944
R8011 gnd.n4785 gnd.n4784 19.3944
R8012 gnd.n4784 gnd.n4783 19.3944
R8013 gnd.n4783 gnd.n4773 19.3944
R8014 gnd.n4779 gnd.n4773 19.3944
R8015 gnd.n4779 gnd.n4778 19.3944
R8016 gnd.n4778 gnd.n4777 19.3944
R8017 gnd.n4777 gnd.n1534 19.3944
R8018 gnd.n4910 gnd.n1534 19.3944
R8019 gnd.n4910 gnd.n1535 19.3944
R8020 gnd.n4906 gnd.n1535 19.3944
R8021 gnd.n4906 gnd.n4905 19.3944
R8022 gnd.n4905 gnd.n4904 19.3944
R8023 gnd.n4904 gnd.n4901 19.3944
R8024 gnd.n4901 gnd.n1425 19.3944
R8025 gnd.n5191 gnd.n1425 19.3944
R8026 gnd.n5191 gnd.n1423 19.3944
R8027 gnd.n5195 gnd.n1423 19.3944
R8028 gnd.n5173 gnd.n5094 19.3944
R8029 gnd.n5177 gnd.n5094 19.3944
R8030 gnd.n5177 gnd.n5095 19.3944
R8031 gnd.n6436 gnd.n6435 19.3944
R8032 gnd.n6435 gnd.n339 19.3944
R8033 gnd.n6428 gnd.n339 19.3944
R8034 gnd.n6428 gnd.n6427 19.3944
R8035 gnd.n6427 gnd.n347 19.3944
R8036 gnd.n6420 gnd.n347 19.3944
R8037 gnd.n6420 gnd.n6419 19.3944
R8038 gnd.n6419 gnd.n355 19.3944
R8039 gnd.n6412 gnd.n355 19.3944
R8040 gnd.n6412 gnd.n6411 19.3944
R8041 gnd.n6411 gnd.n363 19.3944
R8042 gnd.n6404 gnd.n363 19.3944
R8043 gnd.n6404 gnd.n6403 19.3944
R8044 gnd.n6403 gnd.n371 19.3944
R8045 gnd.n6396 gnd.n371 19.3944
R8046 gnd.n6396 gnd.n6395 19.3944
R8047 gnd.n6395 gnd.n381 19.3944
R8048 gnd.n5103 gnd.n381 19.3944
R8049 gnd.n5157 gnd.n5103 19.3944
R8050 gnd.n5160 gnd.n5157 19.3944
R8051 gnd.n5163 gnd.n5160 19.3944
R8052 gnd.n5163 gnd.n5099 19.3944
R8053 gnd.n5167 gnd.n5099 19.3944
R8054 gnd.n5170 gnd.n5167 19.3944
R8055 gnd.n1780 gnd.t235 19.1199
R8056 gnd.n1761 gnd.n1753 19.1199
R8057 gnd.n1712 gnd.n1710 19.1199
R8058 gnd.n1680 gnd.n1672 19.1199
R8059 gnd.n1630 gnd.n1619 19.1199
R8060 gnd.n4798 gnd.t14 19.1199
R8061 gnd.n5063 gnd.n1436 19.1199
R8062 gnd.n2956 gnd.t187 18.8012
R8063 gnd.n2941 gnd.t275 18.8012
R8064 gnd.n2800 gnd.n2799 18.4825
R8065 gnd.n4920 gnd.t143 18.4825
R8066 gnd.n6360 gnd.n6359 18.4247
R8067 gnd.n5409 gnd.n5408 18.4247
R8068 gnd.n6641 gnd.n6640 18.2308
R8069 gnd.n6399 gnd.n377 18.2308
R8070 gnd.n1979 gnd.n1974 18.2308
R8071 gnd.n3645 gnd.n3601 18.2308
R8072 gnd.t222 gnd.n2480 18.1639
R8073 gnd.t240 gnd.n1311 18.1639
R8074 gnd.n4886 gnd.t48 18.1639
R8075 gnd.n4298 gnd.n1325 17.8452
R8076 gnd.n4478 gnd.n1796 17.8452
R8077 gnd.n4602 gnd.n1716 17.8452
R8078 gnd.n4664 gnd.n1658 17.8452
R8079 gnd.n1584 gnd.n1578 17.8452
R8080 gnd.n4868 gnd.n4866 17.8452
R8081 gnd.n2508 gnd.t282 17.5266
R8082 gnd.t56 gnd.n1740 17.5266
R8083 gnd.n4362 gnd.t253 17.5266
R8084 gnd.n3184 gnd.n3183 17.2079
R8085 gnd.n4318 gnd.t11 17.2079
R8086 gnd.t267 gnd.n4879 17.2079
R8087 gnd.n2907 gnd.t223 16.8893
R8088 gnd.n3887 gnd.t159 16.8893
R8089 gnd.t44 gnd.n1032 16.8893
R8090 gnd.n6216 gnd.t51 16.8893
R8091 gnd.t74 gnd.n81 16.8893
R8092 gnd.n4438 gnd.n1815 16.5706
R8093 gnd.n4450 gnd.n4449 16.5706
R8094 gnd.n4561 gnd.n1736 16.5706
R8095 gnd.n4574 gnd.n4572 16.5706
R8096 gnd.n4683 gnd.n1654 16.5706
R8097 gnd.n4696 gnd.n4695 16.5706
R8098 gnd.n4840 gnd.n1574 16.5706
R8099 gnd.n4850 gnd.n1565 16.5706
R8100 gnd.n2735 gnd.t175 16.2519
R8101 gnd.n2435 gnd.t184 16.2519
R8102 gnd.n1839 gnd.t146 16.2519
R8103 gnd.t130 gnd.n1419 16.2519
R8104 gnd.t69 gnd.n4490 15.9333
R8105 gnd.n4804 gnd.t29 15.9333
R8106 gnd.n3423 gnd.n3421 15.6674
R8107 gnd.n3391 gnd.n3389 15.6674
R8108 gnd.n3359 gnd.n3357 15.6674
R8109 gnd.n3328 gnd.n3326 15.6674
R8110 gnd.n3296 gnd.n3294 15.6674
R8111 gnd.n3264 gnd.n3262 15.6674
R8112 gnd.n3232 gnd.n3230 15.6674
R8113 gnd.n3201 gnd.n3199 15.6674
R8114 gnd.n2726 gnd.t175 15.6146
R8115 gnd.t109 gnd.n2201 15.6146
R8116 gnd.t113 gnd.n2202 15.6146
R8117 gnd.t146 gnd.n1149 15.6146
R8118 gnd.n5189 gnd.t130 15.6146
R8119 gnd.n1444 gnd.n1443 15.0827
R8120 gnd.n1193 gnd.n1188 15.0481
R8121 gnd.n1454 gnd.n1453 15.0481
R8122 gnd.n3094 gnd.t199 14.9773
R8123 gnd.t159 gnd.n2104 14.9773
R8124 gnd.n4149 gnd.t95 14.9773
R8125 gnd.n6453 gnd.t88 14.9773
R8126 gnd.n6684 gnd.t74 14.9773
R8127 gnd.n4459 gnd.t19 14.6587
R8128 gnd.n4842 gnd.t6 14.6587
R8129 gnd.t24 gnd.n2244 14.34
R8130 gnd.n3172 gnd.t221 14.34
R8131 gnd.n5307 gnd.n1325 14.0214
R8132 gnd.n4478 gnd.t266 14.0214
R8133 gnd.n4543 gnd.n4541 14.0214
R8134 gnd.n4602 gnd.n4601 14.0214
R8135 gnd.n4665 gnd.n4664 14.0214
R8136 gnd.n4713 gnd.n4712 14.0214
R8137 gnd.t0 gnd.n1584 14.0214
R8138 gnd.n4866 gnd.n1544 14.0214
R8139 gnd.t71 gnd.n1513 14.0214
R8140 gnd.n2882 gnd.t278 13.7027
R8141 gnd.n4439 gnd.t205 13.7027
R8142 gnd.n4851 gnd.t255 13.7027
R8143 gnd.n2592 gnd.n2591 13.5763
R8144 gnd.n3537 gnd.n2158 13.5763
R8145 gnd.n6322 gnd.n462 13.5763
R8146 gnd.n6693 gnd.n6692 13.5763
R8147 gnd.n3805 gnd.n3751 13.5763
R8148 gnd.n4140 gnd.n4139 13.5763
R8149 gnd.n2800 gnd.n2538 13.384
R8150 gnd.n1204 gnd.n1185 13.1884
R8151 gnd.n1199 gnd.n1198 13.1884
R8152 gnd.n1198 gnd.n1197 13.1884
R8153 gnd.n1447 gnd.n1442 13.1884
R8154 gnd.n1448 gnd.n1447 13.1884
R8155 gnd.n1200 gnd.n1187 13.146
R8156 gnd.n1196 gnd.n1187 13.146
R8157 gnd.n1446 gnd.n1445 13.146
R8158 gnd.n1446 gnd.n1441 13.146
R8159 gnd.n3424 gnd.n3420 12.8005
R8160 gnd.n3392 gnd.n3388 12.8005
R8161 gnd.n3360 gnd.n3356 12.8005
R8162 gnd.n3329 gnd.n3325 12.8005
R8163 gnd.n3297 gnd.n3293 12.8005
R8164 gnd.n3265 gnd.n3261 12.8005
R8165 gnd.n3233 gnd.n3229 12.8005
R8166 gnd.n3202 gnd.n3198 12.8005
R8167 gnd.n1292 gnd.n1207 12.7467
R8168 gnd.t106 gnd.t117 12.7467
R8169 gnd.n5313 gnd.n1311 12.7467
R8170 gnd.t262 gnd.n1815 12.7467
R8171 gnd.n1791 gnd.n1786 12.7467
R8172 gnd.n4525 gnd.n1761 12.7467
R8173 gnd.n1710 gnd.n1705 12.7467
R8174 gnd.n4615 gnd.t20 12.7467
R8175 gnd.n4649 gnd.t200 12.7467
R8176 gnd.n4648 gnd.n1680 12.7467
R8177 gnd.n4750 gnd.n1619 12.7467
R8178 gnd.n4816 gnd.n1589 12.7467
R8179 gnd.n1565 gnd.t248 12.7467
R8180 gnd.n4886 gnd.n1540 12.7467
R8181 gnd.t156 gnd.n1525 12.7467
R8182 gnd.t26 gnd.n1791 12.4281
R8183 gnd.n4816 gnd.t46 12.4281
R8184 gnd.n2591 gnd.n2586 12.4126
R8185 gnd.n3540 gnd.n3537 12.4126
R8186 gnd.n6318 gnd.n462 12.4126
R8187 gnd.n6692 gnd.n155 12.4126
R8188 gnd.n3801 gnd.n3751 12.4126
R8189 gnd.n4142 gnd.n4140 12.4126
R8190 gnd.n5401 gnd.n5338 12.1761
R8191 gnd.n5060 gnd.n5059 12.1761
R8192 gnd.n3428 gnd.n3427 12.0247
R8193 gnd.n3396 gnd.n3395 12.0247
R8194 gnd.n3364 gnd.n3363 12.0247
R8195 gnd.n3333 gnd.n3332 12.0247
R8196 gnd.n3301 gnd.n3300 12.0247
R8197 gnd.n3269 gnd.n3268 12.0247
R8198 gnd.n3237 gnd.n3236 12.0247
R8199 gnd.n3206 gnd.n3205 12.0247
R8200 gnd.n2098 gnd.t180 11.7908
R8201 gnd.t95 gnd.n1085 11.7908
R8202 gnd.n5149 gnd.t88 11.7908
R8203 gnd.n6594 gnd.t212 11.7908
R8204 gnd.n4273 gnd.n1211 11.4721
R8205 gnd.n4497 gnd.n1781 11.4721
R8206 gnd.n4517 gnd.n4515 11.4721
R8207 gnd.n4621 gnd.n1701 11.4721
R8208 gnd.n4640 gnd.n4639 11.4721
R8209 gnd.n4760 gnd.n1611 11.4721
R8210 gnd.n4797 gnd.n1598 11.4721
R8211 gnd.n4921 gnd.n1525 11.4721
R8212 gnd.n4929 gnd.n1519 11.4721
R8213 gnd.n3431 gnd.n3418 11.249
R8214 gnd.n3399 gnd.n3386 11.249
R8215 gnd.n3367 gnd.n3354 11.249
R8216 gnd.n3336 gnd.n3323 11.249
R8217 gnd.n3304 gnd.n3291 11.249
R8218 gnd.n3272 gnd.n3259 11.249
R8219 gnd.n3240 gnd.n3227 11.249
R8220 gnd.n3209 gnd.n3196 11.249
R8221 gnd.n2870 gnd.t278 11.1535
R8222 gnd.n2066 gnd.t225 11.1535
R8223 gnd.n6562 gnd.t178 11.1535
R8224 gnd.n1292 gnd.t150 10.8348
R8225 gnd.n4502 gnd.t5 10.8348
R8226 gnd.n4526 gnd.t5 10.8348
R8227 gnd.n4749 gnd.t228 10.8348
R8228 gnd.n4726 gnd.t228 10.8348
R8229 gnd.n4995 gnd.n1485 10.6151
R8230 gnd.n4995 gnd.n4994 10.6151
R8231 gnd.n4992 gnd.n1489 10.6151
R8232 gnd.n4987 gnd.n1489 10.6151
R8233 gnd.n4987 gnd.n4986 10.6151
R8234 gnd.n4986 gnd.n4985 10.6151
R8235 gnd.n4985 gnd.n1492 10.6151
R8236 gnd.n4980 gnd.n1492 10.6151
R8237 gnd.n4980 gnd.n4979 10.6151
R8238 gnd.n4979 gnd.n4978 10.6151
R8239 gnd.n4978 gnd.n1495 10.6151
R8240 gnd.n4973 gnd.n1495 10.6151
R8241 gnd.n4973 gnd.n4972 10.6151
R8242 gnd.n4972 gnd.n4971 10.6151
R8243 gnd.n4971 gnd.n1498 10.6151
R8244 gnd.n4966 gnd.n1498 10.6151
R8245 gnd.n4966 gnd.n4965 10.6151
R8246 gnd.n4965 gnd.n4964 10.6151
R8247 gnd.n4964 gnd.n1501 10.6151
R8248 gnd.n4959 gnd.n1501 10.6151
R8249 gnd.n4959 gnd.n4958 10.6151
R8250 gnd.n4958 gnd.n4957 10.6151
R8251 gnd.n4957 gnd.n1504 10.6151
R8252 gnd.n4952 gnd.n1504 10.6151
R8253 gnd.n4952 gnd.n4951 10.6151
R8254 gnd.n4951 gnd.n4950 10.6151
R8255 gnd.n4950 gnd.n1507 10.6151
R8256 gnd.n4945 gnd.n1507 10.6151
R8257 gnd.n4945 gnd.n4944 10.6151
R8258 gnd.n4944 gnd.n4943 10.6151
R8259 gnd.n1295 gnd.n1294 10.6151
R8260 gnd.n1296 gnd.n1295 10.6151
R8261 gnd.n1298 gnd.n1296 10.6151
R8262 gnd.n1299 gnd.n1298 10.6151
R8263 gnd.n5324 gnd.n1299 10.6151
R8264 gnd.n5324 gnd.n5323 10.6151
R8265 gnd.n5323 gnd.n5322 10.6151
R8266 gnd.n5322 gnd.n1300 10.6151
R8267 gnd.n4301 gnd.n1300 10.6151
R8268 gnd.n4303 gnd.n4301 10.6151
R8269 gnd.n4304 gnd.n4303 10.6151
R8270 gnd.n4306 gnd.n4304 10.6151
R8271 gnd.n4307 gnd.n4306 10.6151
R8272 gnd.n4309 gnd.n4307 10.6151
R8273 gnd.n4309 gnd.n4308 10.6151
R8274 gnd.n4308 gnd.n1813 10.6151
R8275 gnd.n4441 gnd.n1813 10.6151
R8276 gnd.n4442 gnd.n4441 10.6151
R8277 gnd.n4447 gnd.n4442 10.6151
R8278 gnd.n4447 gnd.n4446 10.6151
R8279 gnd.n4446 gnd.n4445 10.6151
R8280 gnd.n4445 gnd.n4443 10.6151
R8281 gnd.n4443 gnd.n1788 10.6151
R8282 gnd.n4486 gnd.n1788 10.6151
R8283 gnd.n4487 gnd.n4486 10.6151
R8284 gnd.n4488 gnd.n4487 10.6151
R8285 gnd.n4488 gnd.n1777 10.6151
R8286 gnd.n4499 gnd.n1777 10.6151
R8287 gnd.n4500 gnd.n4499 10.6151
R8288 gnd.n4507 gnd.n4500 10.6151
R8289 gnd.n4507 gnd.n4506 10.6151
R8290 gnd.n4506 gnd.n4505 10.6151
R8291 gnd.n4505 gnd.n4504 10.6151
R8292 gnd.n4504 gnd.n4501 10.6151
R8293 gnd.n4501 gnd.n1751 10.6151
R8294 gnd.n4535 gnd.n1751 10.6151
R8295 gnd.n4536 gnd.n4535 10.6151
R8296 gnd.n4539 gnd.n4536 10.6151
R8297 gnd.n4539 gnd.n4538 10.6151
R8298 gnd.n4538 gnd.n4537 10.6151
R8299 gnd.n4537 gnd.n1734 10.6151
R8300 gnd.n4564 gnd.n1734 10.6151
R8301 gnd.n4565 gnd.n4564 10.6151
R8302 gnd.n4570 gnd.n4565 10.6151
R8303 gnd.n4570 gnd.n4569 10.6151
R8304 gnd.n4569 gnd.n4568 10.6151
R8305 gnd.n4568 gnd.n4566 10.6151
R8306 gnd.n4566 gnd.n1707 10.6151
R8307 gnd.n4610 gnd.n1707 10.6151
R8308 gnd.n4611 gnd.n4610 10.6151
R8309 gnd.n4612 gnd.n4611 10.6151
R8310 gnd.n4612 gnd.n1698 10.6151
R8311 gnd.n4623 gnd.n1698 10.6151
R8312 gnd.n4624 gnd.n4623 10.6151
R8313 gnd.n4631 gnd.n4624 10.6151
R8314 gnd.n4631 gnd.n4630 10.6151
R8315 gnd.n4630 gnd.n4629 10.6151
R8316 gnd.n4629 gnd.n4628 10.6151
R8317 gnd.n4628 gnd.n4625 10.6151
R8318 gnd.n4625 gnd.n1669 10.6151
R8319 gnd.n4658 gnd.n1669 10.6151
R8320 gnd.n4659 gnd.n4658 10.6151
R8321 gnd.n4662 gnd.n4659 10.6151
R8322 gnd.n4662 gnd.n4661 10.6151
R8323 gnd.n4661 gnd.n4660 10.6151
R8324 gnd.n4660 gnd.n1651 10.6151
R8325 gnd.n4686 gnd.n1651 10.6151
R8326 gnd.n4687 gnd.n4686 10.6151
R8327 gnd.n4693 gnd.n4687 10.6151
R8328 gnd.n4693 gnd.n4692 10.6151
R8329 gnd.n4692 gnd.n4691 10.6151
R8330 gnd.n4691 gnd.n4689 10.6151
R8331 gnd.n4689 gnd.n4688 10.6151
R8332 gnd.n4688 gnd.n1627 10.6151
R8333 gnd.n4722 gnd.n1627 10.6151
R8334 gnd.n4723 gnd.n4722 10.6151
R8335 gnd.n4724 gnd.n4723 10.6151
R8336 gnd.n4729 gnd.n4724 10.6151
R8337 gnd.n4730 gnd.n4729 10.6151
R8338 gnd.n4739 gnd.n4730 10.6151
R8339 gnd.n4739 gnd.n4738 10.6151
R8340 gnd.n4738 gnd.n4737 10.6151
R8341 gnd.n4737 gnd.n4735 10.6151
R8342 gnd.n4735 gnd.n4734 10.6151
R8343 gnd.n4734 gnd.n4731 10.6151
R8344 gnd.n4731 gnd.n1581 10.6151
R8345 gnd.n4824 gnd.n1581 10.6151
R8346 gnd.n4825 gnd.n4824 10.6151
R8347 gnd.n4832 gnd.n4825 10.6151
R8348 gnd.n4832 gnd.n4831 10.6151
R8349 gnd.n4831 gnd.n4830 10.6151
R8350 gnd.n4830 gnd.n4829 10.6151
R8351 gnd.n4829 gnd.n4826 10.6151
R8352 gnd.n4826 gnd.n1556 10.6151
R8353 gnd.n4860 gnd.n1556 10.6151
R8354 gnd.n4861 gnd.n4860 10.6151
R8355 gnd.n4864 gnd.n4861 10.6151
R8356 gnd.n4864 gnd.n4863 10.6151
R8357 gnd.n4863 gnd.n4862 10.6151
R8358 gnd.n4862 gnd.n1538 10.6151
R8359 gnd.n4889 gnd.n1538 10.6151
R8360 gnd.n4890 gnd.n4889 10.6151
R8361 gnd.n4892 gnd.n4890 10.6151
R8362 gnd.n4893 gnd.n4892 10.6151
R8363 gnd.n4896 gnd.n4893 10.6151
R8364 gnd.n4896 gnd.n4895 10.6151
R8365 gnd.n4895 gnd.n4894 10.6151
R8366 gnd.n4894 gnd.n1510 10.6151
R8367 gnd.n4939 gnd.n1510 10.6151
R8368 gnd.n4940 gnd.n4939 10.6151
R8369 gnd.n1229 gnd.n1145 10.6151
R8370 gnd.n1232 gnd.n1229 10.6151
R8371 gnd.n1237 gnd.n1234 10.6151
R8372 gnd.n1238 gnd.n1237 10.6151
R8373 gnd.n1241 gnd.n1238 10.6151
R8374 gnd.n1242 gnd.n1241 10.6151
R8375 gnd.n1245 gnd.n1242 10.6151
R8376 gnd.n1246 gnd.n1245 10.6151
R8377 gnd.n1249 gnd.n1246 10.6151
R8378 gnd.n1250 gnd.n1249 10.6151
R8379 gnd.n1253 gnd.n1250 10.6151
R8380 gnd.n1254 gnd.n1253 10.6151
R8381 gnd.n1257 gnd.n1254 10.6151
R8382 gnd.n1258 gnd.n1257 10.6151
R8383 gnd.n1261 gnd.n1258 10.6151
R8384 gnd.n1262 gnd.n1261 10.6151
R8385 gnd.n1265 gnd.n1262 10.6151
R8386 gnd.n1266 gnd.n1265 10.6151
R8387 gnd.n1269 gnd.n1266 10.6151
R8388 gnd.n1270 gnd.n1269 10.6151
R8389 gnd.n1273 gnd.n1270 10.6151
R8390 gnd.n1274 gnd.n1273 10.6151
R8391 gnd.n1277 gnd.n1274 10.6151
R8392 gnd.n1278 gnd.n1277 10.6151
R8393 gnd.n1281 gnd.n1278 10.6151
R8394 gnd.n1282 gnd.n1281 10.6151
R8395 gnd.n1285 gnd.n1282 10.6151
R8396 gnd.n1286 gnd.n1285 10.6151
R8397 gnd.n1289 gnd.n1286 10.6151
R8398 gnd.n1290 gnd.n1289 10.6151
R8399 gnd.n5401 gnd.n5400 10.6151
R8400 gnd.n5400 gnd.n5399 10.6151
R8401 gnd.n5399 gnd.n5398 10.6151
R8402 gnd.n5398 gnd.n5396 10.6151
R8403 gnd.n5396 gnd.n5393 10.6151
R8404 gnd.n5393 gnd.n5392 10.6151
R8405 gnd.n5392 gnd.n5389 10.6151
R8406 gnd.n5389 gnd.n5388 10.6151
R8407 gnd.n5388 gnd.n5385 10.6151
R8408 gnd.n5385 gnd.n5384 10.6151
R8409 gnd.n5384 gnd.n5381 10.6151
R8410 gnd.n5381 gnd.n5380 10.6151
R8411 gnd.n5380 gnd.n5377 10.6151
R8412 gnd.n5377 gnd.n5376 10.6151
R8413 gnd.n5376 gnd.n5373 10.6151
R8414 gnd.n5373 gnd.n5372 10.6151
R8415 gnd.n5372 gnd.n5369 10.6151
R8416 gnd.n5369 gnd.n5368 10.6151
R8417 gnd.n5368 gnd.n5365 10.6151
R8418 gnd.n5365 gnd.n5364 10.6151
R8419 gnd.n5364 gnd.n5361 10.6151
R8420 gnd.n5361 gnd.n5360 10.6151
R8421 gnd.n5360 gnd.n5357 10.6151
R8422 gnd.n5357 gnd.n5356 10.6151
R8423 gnd.n5356 gnd.n5353 10.6151
R8424 gnd.n5353 gnd.n5352 10.6151
R8425 gnd.n5352 gnd.n5349 10.6151
R8426 gnd.n5349 gnd.n5348 10.6151
R8427 gnd.n5345 gnd.n5344 10.6151
R8428 gnd.n5344 gnd.n1146 10.6151
R8429 gnd.n5059 gnd.n5058 10.6151
R8430 gnd.n5058 gnd.n1459 10.6151
R8431 gnd.n5053 gnd.n1459 10.6151
R8432 gnd.n5053 gnd.n5052 10.6151
R8433 gnd.n5052 gnd.n5051 10.6151
R8434 gnd.n5051 gnd.n1463 10.6151
R8435 gnd.n5046 gnd.n1463 10.6151
R8436 gnd.n5046 gnd.n5045 10.6151
R8437 gnd.n5045 gnd.n5044 10.6151
R8438 gnd.n5044 gnd.n1466 10.6151
R8439 gnd.n5039 gnd.n1466 10.6151
R8440 gnd.n5039 gnd.n5038 10.6151
R8441 gnd.n5038 gnd.n5037 10.6151
R8442 gnd.n5037 gnd.n1469 10.6151
R8443 gnd.n5032 gnd.n1469 10.6151
R8444 gnd.n5032 gnd.n5031 10.6151
R8445 gnd.n5031 gnd.n5030 10.6151
R8446 gnd.n5030 gnd.n1472 10.6151
R8447 gnd.n5025 gnd.n1472 10.6151
R8448 gnd.n5025 gnd.n5024 10.6151
R8449 gnd.n5024 gnd.n5023 10.6151
R8450 gnd.n5023 gnd.n1475 10.6151
R8451 gnd.n5018 gnd.n1475 10.6151
R8452 gnd.n5018 gnd.n5017 10.6151
R8453 gnd.n5017 gnd.n5016 10.6151
R8454 gnd.n5016 gnd.n1478 10.6151
R8455 gnd.n5011 gnd.n1478 10.6151
R8456 gnd.n5011 gnd.n5010 10.6151
R8457 gnd.n5008 gnd.n1483 10.6151
R8458 gnd.n5003 gnd.n1483 10.6151
R8459 gnd.n5337 gnd.n5336 10.6151
R8460 gnd.n5336 gnd.n1205 10.6151
R8461 gnd.n4268 gnd.n1205 10.6151
R8462 gnd.n4270 gnd.n4268 10.6151
R8463 gnd.n4270 gnd.n4269 10.6151
R8464 gnd.n4269 gnd.n1305 10.6151
R8465 gnd.n5318 gnd.n1305 10.6151
R8466 gnd.n5318 gnd.n5317 10.6151
R8467 gnd.n5317 gnd.n5316 10.6151
R8468 gnd.n5316 gnd.n1306 10.6151
R8469 gnd.n4316 gnd.n1306 10.6151
R8470 gnd.n4316 gnd.n4315 10.6151
R8471 gnd.n4315 gnd.n4314 10.6151
R8472 gnd.n4314 gnd.n4293 10.6151
R8473 gnd.n4296 gnd.n4293 10.6151
R8474 gnd.n4296 gnd.n4295 10.6151
R8475 gnd.n4295 gnd.n1809 10.6151
R8476 gnd.n4453 gnd.n1809 10.6151
R8477 gnd.n4454 gnd.n4453 10.6151
R8478 gnd.n4455 gnd.n4454 10.6151
R8479 gnd.n4455 gnd.n1794 10.6151
R8480 gnd.n4480 gnd.n1794 10.6151
R8481 gnd.n4481 gnd.n4480 10.6151
R8482 gnd.n4482 gnd.n4481 10.6151
R8483 gnd.n4482 gnd.n1783 10.6151
R8484 gnd.n4493 gnd.n1783 10.6151
R8485 gnd.n4494 gnd.n4493 10.6151
R8486 gnd.n4495 gnd.n4494 10.6151
R8487 gnd.n4495 gnd.n1771 10.6151
R8488 gnd.n4511 gnd.n1771 10.6151
R8489 gnd.n4512 gnd.n4511 10.6151
R8490 gnd.n4513 gnd.n4512 10.6151
R8491 gnd.n4513 gnd.n1757 10.6151
R8492 gnd.n4528 gnd.n1757 10.6151
R8493 gnd.n4529 gnd.n4528 10.6151
R8494 gnd.n4531 gnd.n4529 10.6151
R8495 gnd.n4531 gnd.n4530 10.6151
R8496 gnd.n4530 gnd.n1738 10.6151
R8497 gnd.n4557 gnd.n1738 10.6151
R8498 gnd.n4558 gnd.n4557 10.6151
R8499 gnd.n4559 gnd.n4558 10.6151
R8500 gnd.n4559 gnd.n1729 10.6151
R8501 gnd.n4577 gnd.n1729 10.6151
R8502 gnd.n4578 gnd.n4577 10.6151
R8503 gnd.n4579 gnd.n4578 10.6151
R8504 gnd.n4579 gnd.n1714 10.6151
R8505 gnd.n4604 gnd.n1714 10.6151
R8506 gnd.n4605 gnd.n4604 10.6151
R8507 gnd.n4606 gnd.n4605 10.6151
R8508 gnd.n4606 gnd.n1703 10.6151
R8509 gnd.n4617 gnd.n1703 10.6151
R8510 gnd.n4618 gnd.n4617 10.6151
R8511 gnd.n4619 gnd.n4618 10.6151
R8512 gnd.n4619 gnd.n1691 10.6151
R8513 gnd.n4635 gnd.n1691 10.6151
R8514 gnd.n4636 gnd.n4635 10.6151
R8515 gnd.n4637 gnd.n4636 10.6151
R8516 gnd.n4637 gnd.n1676 10.6151
R8517 gnd.n4651 gnd.n1676 10.6151
R8518 gnd.n4652 gnd.n4651 10.6151
R8519 gnd.n4654 gnd.n4652 10.6151
R8520 gnd.n4654 gnd.n4653 10.6151
R8521 gnd.n4653 gnd.n1656 10.6151
R8522 gnd.n4679 gnd.n1656 10.6151
R8523 gnd.n4680 gnd.n4679 10.6151
R8524 gnd.n4681 gnd.n4680 10.6151
R8525 gnd.n4681 gnd.n1646 10.6151
R8526 gnd.n4699 gnd.n1646 10.6151
R8527 gnd.n4700 gnd.n4699 10.6151
R8528 gnd.n4701 gnd.n4700 10.6151
R8529 gnd.n4701 gnd.n1632 10.6151
R8530 gnd.n4715 gnd.n1632 10.6151
R8531 gnd.n4716 gnd.n4715 10.6151
R8532 gnd.n4717 gnd.n4716 10.6151
R8533 gnd.n4717 gnd.n1624 10.6151
R8534 gnd.n4747 gnd.n1624 10.6151
R8535 gnd.n4747 gnd.n4746 10.6151
R8536 gnd.n4746 gnd.n4745 10.6151
R8537 gnd.n4745 gnd.n1625 10.6151
R8538 gnd.n1625 gnd.n1602 10.6151
R8539 gnd.n4800 gnd.n1602 10.6151
R8540 gnd.n4801 gnd.n4800 10.6151
R8541 gnd.n4802 gnd.n4801 10.6151
R8542 gnd.n4802 gnd.n1586 10.6151
R8543 gnd.n4818 gnd.n1586 10.6151
R8544 gnd.n4819 gnd.n4818 10.6151
R8545 gnd.n4820 gnd.n4819 10.6151
R8546 gnd.n4820 gnd.n1576 10.6151
R8547 gnd.n4836 gnd.n1576 10.6151
R8548 gnd.n4837 gnd.n4836 10.6151
R8549 gnd.n4838 gnd.n4837 10.6151
R8550 gnd.n4838 gnd.n1561 10.6151
R8551 gnd.n4853 gnd.n1561 10.6151
R8552 gnd.n4854 gnd.n4853 10.6151
R8553 gnd.n4856 gnd.n4854 10.6151
R8554 gnd.n4856 gnd.n4855 10.6151
R8555 gnd.n4855 gnd.n1542 10.6151
R8556 gnd.n4882 gnd.n1542 10.6151
R8557 gnd.n4883 gnd.n4882 10.6151
R8558 gnd.n4884 gnd.n4883 10.6151
R8559 gnd.n4884 gnd.n1529 10.6151
R8560 gnd.n4916 gnd.n1529 10.6151
R8561 gnd.n4917 gnd.n4916 10.6151
R8562 gnd.n4918 gnd.n4917 10.6151
R8563 gnd.n4918 gnd.n1515 10.6151
R8564 gnd.n4932 gnd.n1515 10.6151
R8565 gnd.n4933 gnd.n4932 10.6151
R8566 gnd.n4934 gnd.n4933 10.6151
R8567 gnd.n4934 gnd.n1439 10.6151
R8568 gnd.n5061 gnd.n1439 10.6151
R8569 gnd.n2789 gnd.t201 10.5161
R8570 gnd.n2246 gnd.t24 10.5161
R8571 gnd.n3155 gnd.t221 10.5161
R8572 gnd.t195 gnd.n2029 10.5161
R8573 gnd.n2032 gnd.t38 10.5161
R8574 gnd.n6532 gnd.t30 10.5161
R8575 gnd.n6540 gnd.t193 10.5161
R8576 gnd.n3432 gnd.n3416 10.4732
R8577 gnd.n3400 gnd.n3384 10.4732
R8578 gnd.n3368 gnd.n3352 10.4732
R8579 gnd.n3337 gnd.n3321 10.4732
R8580 gnd.n3305 gnd.n3289 10.4732
R8581 gnd.n3273 gnd.n3257 10.4732
R8582 gnd.n3241 gnd.n3225 10.4732
R8583 gnd.n3210 gnd.n3194 10.4732
R8584 gnd.n4273 gnd.n4272 10.1975
R8585 gnd.n4284 gnd.n1223 10.1975
R8586 gnd.n1781 gnd.n1780 10.1975
R8587 gnd.n1701 gnd.n1693 10.1975
R8588 gnd.n4640 gnd.n1686 10.1975
R8589 gnd.n4798 gnd.n4797 10.1975
R8590 gnd.n4921 gnd.n4920 10.1975
R8591 gnd.n4930 gnd.n4929 10.1975
R8592 gnd.t199 gnd.n2263 9.87883
R8593 gnd.t15 gnd.n2063 9.87883
R8594 gnd.n5494 gnd.n998 9.87883
R8595 gnd.n4022 gnd.t44 9.87883
R8596 gnd.n6493 gnd.t51 9.87883
R8597 gnd.n6201 gnd.n247 9.87883
R8598 gnd.n6570 gnd.t12 9.87883
R8599 gnd.n3436 gnd.n3435 9.69747
R8600 gnd.n3404 gnd.n3403 9.69747
R8601 gnd.n3372 gnd.n3371 9.69747
R8602 gnd.n3341 gnd.n3340 9.69747
R8603 gnd.n3309 gnd.n3308 9.69747
R8604 gnd.n3277 gnd.n3276 9.69747
R8605 gnd.n3245 gnd.n3244 9.69747
R8606 gnd.n3214 gnd.n3213 9.69747
R8607 gnd.n6799 gnd.n50 9.6512
R8608 gnd.n4553 gnd.t21 9.56018
R8609 gnd.n4704 gnd.t37 9.56018
R8610 gnd.n1910 gnd.n1909 9.45599
R8611 gnd.n6441 gnd.n6440 9.45599
R8612 gnd.n3442 gnd.n3441 9.45567
R8613 gnd.n3410 gnd.n3409 9.45567
R8614 gnd.n3378 gnd.n3377 9.45567
R8615 gnd.n3347 gnd.n3346 9.45567
R8616 gnd.n3315 gnd.n3314 9.45567
R8617 gnd.n3283 gnd.n3282 9.45567
R8618 gnd.n3251 gnd.n3250 9.45567
R8619 gnd.n3220 gnd.n3219 9.45567
R8620 gnd.n2387 gnd.n2386 9.39724
R8621 gnd.n3441 gnd.n3440 9.3005
R8622 gnd.n3414 gnd.n3413 9.3005
R8623 gnd.n3435 gnd.n3434 9.3005
R8624 gnd.n3433 gnd.n3432 9.3005
R8625 gnd.n3418 gnd.n3417 9.3005
R8626 gnd.n3427 gnd.n3426 9.3005
R8627 gnd.n3425 gnd.n3424 9.3005
R8628 gnd.n3409 gnd.n3408 9.3005
R8629 gnd.n3382 gnd.n3381 9.3005
R8630 gnd.n3403 gnd.n3402 9.3005
R8631 gnd.n3401 gnd.n3400 9.3005
R8632 gnd.n3386 gnd.n3385 9.3005
R8633 gnd.n3395 gnd.n3394 9.3005
R8634 gnd.n3393 gnd.n3392 9.3005
R8635 gnd.n3377 gnd.n3376 9.3005
R8636 gnd.n3350 gnd.n3349 9.3005
R8637 gnd.n3371 gnd.n3370 9.3005
R8638 gnd.n3369 gnd.n3368 9.3005
R8639 gnd.n3354 gnd.n3353 9.3005
R8640 gnd.n3363 gnd.n3362 9.3005
R8641 gnd.n3361 gnd.n3360 9.3005
R8642 gnd.n3346 gnd.n3345 9.3005
R8643 gnd.n3319 gnd.n3318 9.3005
R8644 gnd.n3340 gnd.n3339 9.3005
R8645 gnd.n3338 gnd.n3337 9.3005
R8646 gnd.n3323 gnd.n3322 9.3005
R8647 gnd.n3332 gnd.n3331 9.3005
R8648 gnd.n3330 gnd.n3329 9.3005
R8649 gnd.n3314 gnd.n3313 9.3005
R8650 gnd.n3287 gnd.n3286 9.3005
R8651 gnd.n3308 gnd.n3307 9.3005
R8652 gnd.n3306 gnd.n3305 9.3005
R8653 gnd.n3291 gnd.n3290 9.3005
R8654 gnd.n3300 gnd.n3299 9.3005
R8655 gnd.n3298 gnd.n3297 9.3005
R8656 gnd.n3282 gnd.n3281 9.3005
R8657 gnd.n3255 gnd.n3254 9.3005
R8658 gnd.n3276 gnd.n3275 9.3005
R8659 gnd.n3274 gnd.n3273 9.3005
R8660 gnd.n3259 gnd.n3258 9.3005
R8661 gnd.n3268 gnd.n3267 9.3005
R8662 gnd.n3266 gnd.n3265 9.3005
R8663 gnd.n3250 gnd.n3249 9.3005
R8664 gnd.n3223 gnd.n3222 9.3005
R8665 gnd.n3244 gnd.n3243 9.3005
R8666 gnd.n3242 gnd.n3241 9.3005
R8667 gnd.n3227 gnd.n3226 9.3005
R8668 gnd.n3236 gnd.n3235 9.3005
R8669 gnd.n3234 gnd.n3233 9.3005
R8670 gnd.n3219 gnd.n3218 9.3005
R8671 gnd.n3192 gnd.n3191 9.3005
R8672 gnd.n3213 gnd.n3212 9.3005
R8673 gnd.n3211 gnd.n3210 9.3005
R8674 gnd.n3196 gnd.n3195 9.3005
R8675 gnd.n3205 gnd.n3204 9.3005
R8676 gnd.n3203 gnd.n3202 9.3005
R8677 gnd.n3567 gnd.n3566 9.3005
R8678 gnd.n3565 gnd.n2146 9.3005
R8679 gnd.n3564 gnd.n3563 9.3005
R8680 gnd.n3560 gnd.n2147 9.3005
R8681 gnd.n3557 gnd.n2148 9.3005
R8682 gnd.n3556 gnd.n2149 9.3005
R8683 gnd.n3553 gnd.n2150 9.3005
R8684 gnd.n3552 gnd.n2151 9.3005
R8685 gnd.n3549 gnd.n2152 9.3005
R8686 gnd.n3548 gnd.n2153 9.3005
R8687 gnd.n3545 gnd.n2154 9.3005
R8688 gnd.n3544 gnd.n2155 9.3005
R8689 gnd.n3541 gnd.n2156 9.3005
R8690 gnd.n3540 gnd.n2157 9.3005
R8691 gnd.n3537 gnd.n3536 9.3005
R8692 gnd.n3535 gnd.n2158 9.3005
R8693 gnd.n3568 gnd.n2145 9.3005
R8694 gnd.n2808 gnd.n2807 9.3005
R8695 gnd.n2512 gnd.n2511 9.3005
R8696 gnd.n2835 gnd.n2834 9.3005
R8697 gnd.n2836 gnd.n2510 9.3005
R8698 gnd.n2840 gnd.n2837 9.3005
R8699 gnd.n2839 gnd.n2838 9.3005
R8700 gnd.n2484 gnd.n2483 9.3005
R8701 gnd.n2865 gnd.n2864 9.3005
R8702 gnd.n2866 gnd.n2482 9.3005
R8703 gnd.n2868 gnd.n2867 9.3005
R8704 gnd.n2462 gnd.n2461 9.3005
R8705 gnd.n2896 gnd.n2895 9.3005
R8706 gnd.n2897 gnd.n2460 9.3005
R8707 gnd.n2905 gnd.n2898 9.3005
R8708 gnd.n2904 gnd.n2899 9.3005
R8709 gnd.n2903 gnd.n2901 9.3005
R8710 gnd.n2900 gnd.n2409 9.3005
R8711 gnd.n2953 gnd.n2410 9.3005
R8712 gnd.n2952 gnd.n2411 9.3005
R8713 gnd.n2951 gnd.n2412 9.3005
R8714 gnd.n2431 gnd.n2413 9.3005
R8715 gnd.n2433 gnd.n2432 9.3005
R8716 gnd.n2343 gnd.n2342 9.3005
R8717 gnd.n2991 gnd.n2990 9.3005
R8718 gnd.n2992 gnd.n2341 9.3005
R8719 gnd.n2996 gnd.n2993 9.3005
R8720 gnd.n2995 gnd.n2994 9.3005
R8721 gnd.n2316 gnd.n2315 9.3005
R8722 gnd.n3031 gnd.n3030 9.3005
R8723 gnd.n3032 gnd.n2314 9.3005
R8724 gnd.n3036 gnd.n3033 9.3005
R8725 gnd.n3035 gnd.n3034 9.3005
R8726 gnd.n2289 gnd.n2288 9.3005
R8727 gnd.n3076 gnd.n3075 9.3005
R8728 gnd.n3077 gnd.n2287 9.3005
R8729 gnd.n3081 gnd.n3078 9.3005
R8730 gnd.n3080 gnd.n3079 9.3005
R8731 gnd.n2261 gnd.n2260 9.3005
R8732 gnd.n3116 gnd.n3115 9.3005
R8733 gnd.n3117 gnd.n2259 9.3005
R8734 gnd.n3121 gnd.n3118 9.3005
R8735 gnd.n3120 gnd.n3119 9.3005
R8736 gnd.n2234 gnd.n2233 9.3005
R8737 gnd.n3165 gnd.n3164 9.3005
R8738 gnd.n3166 gnd.n2232 9.3005
R8739 gnd.n3170 gnd.n3167 9.3005
R8740 gnd.n3169 gnd.n3168 9.3005
R8741 gnd.n2207 gnd.n2206 9.3005
R8742 gnd.n3460 gnd.n3459 9.3005
R8743 gnd.n3461 gnd.n2205 9.3005
R8744 gnd.n3467 gnd.n3462 9.3005
R8745 gnd.n3466 gnd.n3463 9.3005
R8746 gnd.n3465 gnd.n3464 9.3005
R8747 gnd.n2809 gnd.n2806 9.3005
R8748 gnd.n2591 gnd.n2550 9.3005
R8749 gnd.n2586 gnd.n2585 9.3005
R8750 gnd.n2584 gnd.n2551 9.3005
R8751 gnd.n2583 gnd.n2582 9.3005
R8752 gnd.n2579 gnd.n2552 9.3005
R8753 gnd.n2576 gnd.n2575 9.3005
R8754 gnd.n2574 gnd.n2553 9.3005
R8755 gnd.n2573 gnd.n2572 9.3005
R8756 gnd.n2569 gnd.n2554 9.3005
R8757 gnd.n2566 gnd.n2565 9.3005
R8758 gnd.n2564 gnd.n2555 9.3005
R8759 gnd.n2563 gnd.n2562 9.3005
R8760 gnd.n2559 gnd.n2557 9.3005
R8761 gnd.n2556 gnd.n2536 9.3005
R8762 gnd.n2803 gnd.n2535 9.3005
R8763 gnd.n2805 gnd.n2804 9.3005
R8764 gnd.n2593 gnd.n2592 9.3005
R8765 gnd.n2816 gnd.n2522 9.3005
R8766 gnd.n2823 gnd.n2523 9.3005
R8767 gnd.n2825 gnd.n2824 9.3005
R8768 gnd.n2826 gnd.n2503 9.3005
R8769 gnd.n2845 gnd.n2844 9.3005
R8770 gnd.n2847 gnd.n2495 9.3005
R8771 gnd.n2854 gnd.n2497 9.3005
R8772 gnd.n2855 gnd.n2492 9.3005
R8773 gnd.n2857 gnd.n2856 9.3005
R8774 gnd.n2493 gnd.n2478 9.3005
R8775 gnd.n2873 gnd.n2476 9.3005
R8776 gnd.n2877 gnd.n2876 9.3005
R8777 gnd.n2875 gnd.n2452 9.3005
R8778 gnd.n2912 gnd.n2451 9.3005
R8779 gnd.n2915 gnd.n2914 9.3005
R8780 gnd.n2448 gnd.n2447 9.3005
R8781 gnd.n2921 gnd.n2449 9.3005
R8782 gnd.n2923 gnd.n2922 9.3005
R8783 gnd.n2925 gnd.n2446 9.3005
R8784 gnd.n2928 gnd.n2927 9.3005
R8785 gnd.n2931 gnd.n2929 9.3005
R8786 gnd.n2933 gnd.n2932 9.3005
R8787 gnd.n2939 gnd.n2934 9.3005
R8788 gnd.n2938 gnd.n2937 9.3005
R8789 gnd.n2334 gnd.n2333 9.3005
R8790 gnd.n3005 gnd.n3004 9.3005
R8791 gnd.n3006 gnd.n2327 9.3005
R8792 gnd.n3014 gnd.n2326 9.3005
R8793 gnd.n3017 gnd.n3016 9.3005
R8794 gnd.n3019 gnd.n3018 9.3005
R8795 gnd.n3022 gnd.n2309 9.3005
R8796 gnd.n3020 gnd.n2307 9.3005
R8797 gnd.n3042 gnd.n2305 9.3005
R8798 gnd.n3044 gnd.n3043 9.3005
R8799 gnd.n2279 gnd.n2278 9.3005
R8800 gnd.n3090 gnd.n3089 9.3005
R8801 gnd.n3091 gnd.n2272 9.3005
R8802 gnd.n3099 gnd.n2271 9.3005
R8803 gnd.n3102 gnd.n3101 9.3005
R8804 gnd.n3104 gnd.n3103 9.3005
R8805 gnd.n3107 gnd.n2254 9.3005
R8806 gnd.n3105 gnd.n2252 9.3005
R8807 gnd.n3127 gnd.n2250 9.3005
R8808 gnd.n3129 gnd.n3128 9.3005
R8809 gnd.n2225 gnd.n2224 9.3005
R8810 gnd.n3179 gnd.n3178 9.3005
R8811 gnd.n3180 gnd.n2218 9.3005
R8812 gnd.n3189 gnd.n2217 9.3005
R8813 gnd.n3448 gnd.n3447 9.3005
R8814 gnd.n3450 gnd.n3449 9.3005
R8815 gnd.n3451 gnd.n2198 9.3005
R8816 gnd.n3475 gnd.n3474 9.3005
R8817 gnd.n2199 gnd.n2161 9.3005
R8818 gnd.n2814 gnd.n2813 9.3005
R8819 gnd.n3531 gnd.n2162 9.3005
R8820 gnd.n3530 gnd.n2164 9.3005
R8821 gnd.n3527 gnd.n2165 9.3005
R8822 gnd.n3526 gnd.n2166 9.3005
R8823 gnd.n3523 gnd.n2167 9.3005
R8824 gnd.n3522 gnd.n2168 9.3005
R8825 gnd.n3519 gnd.n2169 9.3005
R8826 gnd.n3518 gnd.n2170 9.3005
R8827 gnd.n3515 gnd.n2171 9.3005
R8828 gnd.n3514 gnd.n2172 9.3005
R8829 gnd.n3511 gnd.n2173 9.3005
R8830 gnd.n3510 gnd.n2174 9.3005
R8831 gnd.n3507 gnd.n2175 9.3005
R8832 gnd.n3506 gnd.n2176 9.3005
R8833 gnd.n3503 gnd.n2177 9.3005
R8834 gnd.n3502 gnd.n2178 9.3005
R8835 gnd.n3499 gnd.n2179 9.3005
R8836 gnd.n3498 gnd.n2180 9.3005
R8837 gnd.n3495 gnd.n2181 9.3005
R8838 gnd.n3494 gnd.n2182 9.3005
R8839 gnd.n3491 gnd.n2183 9.3005
R8840 gnd.n3490 gnd.n2184 9.3005
R8841 gnd.n3487 gnd.n2188 9.3005
R8842 gnd.n3486 gnd.n2189 9.3005
R8843 gnd.n3483 gnd.n2190 9.3005
R8844 gnd.n3482 gnd.n2191 9.3005
R8845 gnd.n3533 gnd.n3532 9.3005
R8846 gnd.n2983 gnd.n2967 9.3005
R8847 gnd.n2982 gnd.n2968 9.3005
R8848 gnd.n2981 gnd.n2969 9.3005
R8849 gnd.n2979 gnd.n2970 9.3005
R8850 gnd.n2978 gnd.n2971 9.3005
R8851 gnd.n2976 gnd.n2972 9.3005
R8852 gnd.n2975 gnd.n2973 9.3005
R8853 gnd.n2297 gnd.n2296 9.3005
R8854 gnd.n3052 gnd.n3051 9.3005
R8855 gnd.n3053 gnd.n2295 9.3005
R8856 gnd.n3070 gnd.n3054 9.3005
R8857 gnd.n3069 gnd.n3055 9.3005
R8858 gnd.n3068 gnd.n3056 9.3005
R8859 gnd.n3066 gnd.n3057 9.3005
R8860 gnd.n3065 gnd.n3058 9.3005
R8861 gnd.n3063 gnd.n3059 9.3005
R8862 gnd.n3062 gnd.n3060 9.3005
R8863 gnd.n2241 gnd.n2240 9.3005
R8864 gnd.n3137 gnd.n3136 9.3005
R8865 gnd.n3138 gnd.n2239 9.3005
R8866 gnd.n3159 gnd.n3139 9.3005
R8867 gnd.n3158 gnd.n3140 9.3005
R8868 gnd.n3157 gnd.n3141 9.3005
R8869 gnd.n3154 gnd.n3142 9.3005
R8870 gnd.n3153 gnd.n3143 9.3005
R8871 gnd.n3151 gnd.n3144 9.3005
R8872 gnd.n3150 gnd.n3145 9.3005
R8873 gnd.n3148 gnd.n3147 9.3005
R8874 gnd.n3146 gnd.n2193 9.3005
R8875 gnd.n2724 gnd.n2723 9.3005
R8876 gnd.n2614 gnd.n2613 9.3005
R8877 gnd.n2738 gnd.n2737 9.3005
R8878 gnd.n2739 gnd.n2612 9.3005
R8879 gnd.n2741 gnd.n2740 9.3005
R8880 gnd.n2602 gnd.n2601 9.3005
R8881 gnd.n2754 gnd.n2753 9.3005
R8882 gnd.n2755 gnd.n2600 9.3005
R8883 gnd.n2787 gnd.n2756 9.3005
R8884 gnd.n2786 gnd.n2757 9.3005
R8885 gnd.n2785 gnd.n2758 9.3005
R8886 gnd.n2784 gnd.n2759 9.3005
R8887 gnd.n2781 gnd.n2760 9.3005
R8888 gnd.n2780 gnd.n2761 9.3005
R8889 gnd.n2779 gnd.n2762 9.3005
R8890 gnd.n2777 gnd.n2763 9.3005
R8891 gnd.n2776 gnd.n2764 9.3005
R8892 gnd.n2773 gnd.n2765 9.3005
R8893 gnd.n2772 gnd.n2766 9.3005
R8894 gnd.n2771 gnd.n2767 9.3005
R8895 gnd.n2769 gnd.n2768 9.3005
R8896 gnd.n2468 gnd.n2467 9.3005
R8897 gnd.n2885 gnd.n2884 9.3005
R8898 gnd.n2886 gnd.n2466 9.3005
R8899 gnd.n2890 gnd.n2887 9.3005
R8900 gnd.n2889 gnd.n2888 9.3005
R8901 gnd.n2390 gnd.n2389 9.3005
R8902 gnd.n2965 gnd.n2964 9.3005
R8903 gnd.n2722 gnd.n2623 9.3005
R8904 gnd.n2625 gnd.n2624 9.3005
R8905 gnd.n2669 gnd.n2667 9.3005
R8906 gnd.n2670 gnd.n2666 9.3005
R8907 gnd.n2673 gnd.n2662 9.3005
R8908 gnd.n2674 gnd.n2661 9.3005
R8909 gnd.n2677 gnd.n2660 9.3005
R8910 gnd.n2678 gnd.n2659 9.3005
R8911 gnd.n2681 gnd.n2658 9.3005
R8912 gnd.n2682 gnd.n2657 9.3005
R8913 gnd.n2685 gnd.n2656 9.3005
R8914 gnd.n2686 gnd.n2655 9.3005
R8915 gnd.n2689 gnd.n2654 9.3005
R8916 gnd.n2690 gnd.n2653 9.3005
R8917 gnd.n2693 gnd.n2652 9.3005
R8918 gnd.n2694 gnd.n2651 9.3005
R8919 gnd.n2697 gnd.n2650 9.3005
R8920 gnd.n2698 gnd.n2649 9.3005
R8921 gnd.n2701 gnd.n2648 9.3005
R8922 gnd.n2702 gnd.n2647 9.3005
R8923 gnd.n2705 gnd.n2646 9.3005
R8924 gnd.n2706 gnd.n2645 9.3005
R8925 gnd.n2709 gnd.n2644 9.3005
R8926 gnd.n2711 gnd.n2643 9.3005
R8927 gnd.n2712 gnd.n2642 9.3005
R8928 gnd.n2713 gnd.n2641 9.3005
R8929 gnd.n2714 gnd.n2640 9.3005
R8930 gnd.n2721 gnd.n2720 9.3005
R8931 gnd.n2730 gnd.n2729 9.3005
R8932 gnd.n2731 gnd.n2617 9.3005
R8933 gnd.n2733 gnd.n2732 9.3005
R8934 gnd.n2608 gnd.n2607 9.3005
R8935 gnd.n2746 gnd.n2745 9.3005
R8936 gnd.n2747 gnd.n2606 9.3005
R8937 gnd.n2749 gnd.n2748 9.3005
R8938 gnd.n2595 gnd.n2594 9.3005
R8939 gnd.n2792 gnd.n2791 9.3005
R8940 gnd.n2793 gnd.n2549 9.3005
R8941 gnd.n2797 gnd.n2795 9.3005
R8942 gnd.n2796 gnd.n2528 9.3005
R8943 gnd.n2815 gnd.n2527 9.3005
R8944 gnd.n2818 gnd.n2817 9.3005
R8945 gnd.n2521 gnd.n2520 9.3005
R8946 gnd.n2829 gnd.n2827 9.3005
R8947 gnd.n2828 gnd.n2502 9.3005
R8948 gnd.n2846 gnd.n2501 9.3005
R8949 gnd.n2849 gnd.n2848 9.3005
R8950 gnd.n2496 gnd.n2491 9.3005
R8951 gnd.n2859 gnd.n2858 9.3005
R8952 gnd.n2494 gnd.n2474 9.3005
R8953 gnd.n2880 gnd.n2475 9.3005
R8954 gnd.n2879 gnd.n2878 9.3005
R8955 gnd.n2477 gnd.n2453 9.3005
R8956 gnd.n2911 gnd.n2910 9.3005
R8957 gnd.n2913 gnd.n2398 9.3005
R8958 gnd.n2960 gnd.n2399 9.3005
R8959 gnd.n2959 gnd.n2400 9.3005
R8960 gnd.n2958 gnd.n2401 9.3005
R8961 gnd.n2924 gnd.n2402 9.3005
R8962 gnd.n2926 gnd.n2420 9.3005
R8963 gnd.n2946 gnd.n2421 9.3005
R8964 gnd.n2945 gnd.n2422 9.3005
R8965 gnd.n2944 gnd.n2423 9.3005
R8966 gnd.n2935 gnd.n2424 9.3005
R8967 gnd.n2936 gnd.n2335 9.3005
R8968 gnd.n3002 gnd.n3001 9.3005
R8969 gnd.n3003 gnd.n2328 9.3005
R8970 gnd.n3013 gnd.n3012 9.3005
R8971 gnd.n3015 gnd.n2324 9.3005
R8972 gnd.n3025 gnd.n2325 9.3005
R8973 gnd.n3024 gnd.n3023 9.3005
R8974 gnd.n3021 gnd.n2303 9.3005
R8975 gnd.n3047 gnd.n2304 9.3005
R8976 gnd.n3046 gnd.n3045 9.3005
R8977 gnd.n2306 gnd.n2280 9.3005
R8978 gnd.n3087 gnd.n3086 9.3005
R8979 gnd.n3088 gnd.n2273 9.3005
R8980 gnd.n3098 gnd.n3097 9.3005
R8981 gnd.n3100 gnd.n2269 9.3005
R8982 gnd.n3110 gnd.n2270 9.3005
R8983 gnd.n3109 gnd.n3108 9.3005
R8984 gnd.n3106 gnd.n2248 9.3005
R8985 gnd.n3132 gnd.n2249 9.3005
R8986 gnd.n3131 gnd.n3130 9.3005
R8987 gnd.n2251 gnd.n2226 9.3005
R8988 gnd.n3176 gnd.n3175 9.3005
R8989 gnd.n3177 gnd.n2219 9.3005
R8990 gnd.n3188 gnd.n3187 9.3005
R8991 gnd.n3446 gnd.n2215 9.3005
R8992 gnd.n3454 gnd.n2216 9.3005
R8993 gnd.n3453 gnd.n3452 9.3005
R8994 gnd.n2197 gnd.n2196 9.3005
R8995 gnd.n3477 gnd.n3476 9.3005
R8996 gnd.n2619 gnd.n2618 9.3005
R8997 gnd.n5666 gnd.n828 9.3005
R8998 gnd.n5668 gnd.n5667 9.3005
R8999 gnd.n824 gnd.n823 9.3005
R9000 gnd.n5675 gnd.n5674 9.3005
R9001 gnd.n5676 gnd.n822 9.3005
R9002 gnd.n5678 gnd.n5677 9.3005
R9003 gnd.n818 gnd.n817 9.3005
R9004 gnd.n5685 gnd.n5684 9.3005
R9005 gnd.n5686 gnd.n816 9.3005
R9006 gnd.n5688 gnd.n5687 9.3005
R9007 gnd.n812 gnd.n811 9.3005
R9008 gnd.n5695 gnd.n5694 9.3005
R9009 gnd.n5696 gnd.n810 9.3005
R9010 gnd.n5698 gnd.n5697 9.3005
R9011 gnd.n806 gnd.n805 9.3005
R9012 gnd.n5705 gnd.n5704 9.3005
R9013 gnd.n5706 gnd.n804 9.3005
R9014 gnd.n5708 gnd.n5707 9.3005
R9015 gnd.n800 gnd.n799 9.3005
R9016 gnd.n5715 gnd.n5714 9.3005
R9017 gnd.n5716 gnd.n798 9.3005
R9018 gnd.n5718 gnd.n5717 9.3005
R9019 gnd.n794 gnd.n793 9.3005
R9020 gnd.n5725 gnd.n5724 9.3005
R9021 gnd.n5726 gnd.n792 9.3005
R9022 gnd.n5728 gnd.n5727 9.3005
R9023 gnd.n788 gnd.n787 9.3005
R9024 gnd.n5735 gnd.n5734 9.3005
R9025 gnd.n5736 gnd.n786 9.3005
R9026 gnd.n5738 gnd.n5737 9.3005
R9027 gnd.n782 gnd.n781 9.3005
R9028 gnd.n5745 gnd.n5744 9.3005
R9029 gnd.n5746 gnd.n780 9.3005
R9030 gnd.n5748 gnd.n5747 9.3005
R9031 gnd.n776 gnd.n775 9.3005
R9032 gnd.n5755 gnd.n5754 9.3005
R9033 gnd.n5756 gnd.n774 9.3005
R9034 gnd.n5758 gnd.n5757 9.3005
R9035 gnd.n770 gnd.n769 9.3005
R9036 gnd.n5765 gnd.n5764 9.3005
R9037 gnd.n5766 gnd.n768 9.3005
R9038 gnd.n5768 gnd.n5767 9.3005
R9039 gnd.n764 gnd.n763 9.3005
R9040 gnd.n5775 gnd.n5774 9.3005
R9041 gnd.n5776 gnd.n762 9.3005
R9042 gnd.n5778 gnd.n5777 9.3005
R9043 gnd.n758 gnd.n757 9.3005
R9044 gnd.n5785 gnd.n5784 9.3005
R9045 gnd.n5786 gnd.n756 9.3005
R9046 gnd.n5788 gnd.n5787 9.3005
R9047 gnd.n752 gnd.n751 9.3005
R9048 gnd.n5795 gnd.n5794 9.3005
R9049 gnd.n5796 gnd.n750 9.3005
R9050 gnd.n5798 gnd.n5797 9.3005
R9051 gnd.n746 gnd.n745 9.3005
R9052 gnd.n5805 gnd.n5804 9.3005
R9053 gnd.n5806 gnd.n744 9.3005
R9054 gnd.n5808 gnd.n5807 9.3005
R9055 gnd.n740 gnd.n739 9.3005
R9056 gnd.n5815 gnd.n5814 9.3005
R9057 gnd.n5816 gnd.n738 9.3005
R9058 gnd.n5818 gnd.n5817 9.3005
R9059 gnd.n734 gnd.n733 9.3005
R9060 gnd.n5825 gnd.n5824 9.3005
R9061 gnd.n5826 gnd.n732 9.3005
R9062 gnd.n5828 gnd.n5827 9.3005
R9063 gnd.n728 gnd.n727 9.3005
R9064 gnd.n5835 gnd.n5834 9.3005
R9065 gnd.n5836 gnd.n726 9.3005
R9066 gnd.n5838 gnd.n5837 9.3005
R9067 gnd.n722 gnd.n721 9.3005
R9068 gnd.n5845 gnd.n5844 9.3005
R9069 gnd.n5846 gnd.n720 9.3005
R9070 gnd.n5848 gnd.n5847 9.3005
R9071 gnd.n716 gnd.n715 9.3005
R9072 gnd.n5855 gnd.n5854 9.3005
R9073 gnd.n5856 gnd.n714 9.3005
R9074 gnd.n5858 gnd.n5857 9.3005
R9075 gnd.n710 gnd.n709 9.3005
R9076 gnd.n5865 gnd.n5864 9.3005
R9077 gnd.n5866 gnd.n708 9.3005
R9078 gnd.n5868 gnd.n5867 9.3005
R9079 gnd.n704 gnd.n703 9.3005
R9080 gnd.n5875 gnd.n5874 9.3005
R9081 gnd.n5876 gnd.n702 9.3005
R9082 gnd.n5878 gnd.n5877 9.3005
R9083 gnd.n698 gnd.n697 9.3005
R9084 gnd.n5885 gnd.n5884 9.3005
R9085 gnd.n5886 gnd.n696 9.3005
R9086 gnd.n5888 gnd.n5887 9.3005
R9087 gnd.n692 gnd.n691 9.3005
R9088 gnd.n5895 gnd.n5894 9.3005
R9089 gnd.n5896 gnd.n690 9.3005
R9090 gnd.n5898 gnd.n5897 9.3005
R9091 gnd.n686 gnd.n685 9.3005
R9092 gnd.n5905 gnd.n5904 9.3005
R9093 gnd.n5906 gnd.n684 9.3005
R9094 gnd.n5908 gnd.n5907 9.3005
R9095 gnd.n680 gnd.n679 9.3005
R9096 gnd.n5915 gnd.n5914 9.3005
R9097 gnd.n5916 gnd.n678 9.3005
R9098 gnd.n5918 gnd.n5917 9.3005
R9099 gnd.n674 gnd.n673 9.3005
R9100 gnd.n5925 gnd.n5924 9.3005
R9101 gnd.n5926 gnd.n672 9.3005
R9102 gnd.n5928 gnd.n5927 9.3005
R9103 gnd.n668 gnd.n667 9.3005
R9104 gnd.n5935 gnd.n5934 9.3005
R9105 gnd.n5936 gnd.n666 9.3005
R9106 gnd.n5938 gnd.n5937 9.3005
R9107 gnd.n662 gnd.n661 9.3005
R9108 gnd.n5945 gnd.n5944 9.3005
R9109 gnd.n5946 gnd.n660 9.3005
R9110 gnd.n5948 gnd.n5947 9.3005
R9111 gnd.n656 gnd.n655 9.3005
R9112 gnd.n5955 gnd.n5954 9.3005
R9113 gnd.n5956 gnd.n654 9.3005
R9114 gnd.n5958 gnd.n5957 9.3005
R9115 gnd.n650 gnd.n649 9.3005
R9116 gnd.n5965 gnd.n5964 9.3005
R9117 gnd.n5966 gnd.n648 9.3005
R9118 gnd.n5968 gnd.n5967 9.3005
R9119 gnd.n644 gnd.n643 9.3005
R9120 gnd.n5975 gnd.n5974 9.3005
R9121 gnd.n5976 gnd.n642 9.3005
R9122 gnd.n5979 gnd.n5978 9.3005
R9123 gnd.n5977 gnd.n638 9.3005
R9124 gnd.n5985 gnd.n637 9.3005
R9125 gnd.n5987 gnd.n5986 9.3005
R9126 gnd.n633 gnd.n632 9.3005
R9127 gnd.n5996 gnd.n5995 9.3005
R9128 gnd.n5997 gnd.n631 9.3005
R9129 gnd.n5999 gnd.n5998 9.3005
R9130 gnd.n627 gnd.n626 9.3005
R9131 gnd.n6006 gnd.n6005 9.3005
R9132 gnd.n6007 gnd.n625 9.3005
R9133 gnd.n6009 gnd.n6008 9.3005
R9134 gnd.n621 gnd.n620 9.3005
R9135 gnd.n6016 gnd.n6015 9.3005
R9136 gnd.n6017 gnd.n619 9.3005
R9137 gnd.n6019 gnd.n6018 9.3005
R9138 gnd.n615 gnd.n614 9.3005
R9139 gnd.n6026 gnd.n6025 9.3005
R9140 gnd.n6027 gnd.n613 9.3005
R9141 gnd.n6029 gnd.n6028 9.3005
R9142 gnd.n609 gnd.n608 9.3005
R9143 gnd.n6036 gnd.n6035 9.3005
R9144 gnd.n6037 gnd.n607 9.3005
R9145 gnd.n6039 gnd.n6038 9.3005
R9146 gnd.n603 gnd.n602 9.3005
R9147 gnd.n6046 gnd.n6045 9.3005
R9148 gnd.n6047 gnd.n601 9.3005
R9149 gnd.n6049 gnd.n6048 9.3005
R9150 gnd.n597 gnd.n596 9.3005
R9151 gnd.n6056 gnd.n6055 9.3005
R9152 gnd.n6057 gnd.n595 9.3005
R9153 gnd.n6059 gnd.n6058 9.3005
R9154 gnd.n591 gnd.n590 9.3005
R9155 gnd.n6066 gnd.n6065 9.3005
R9156 gnd.n6067 gnd.n589 9.3005
R9157 gnd.n6069 gnd.n6068 9.3005
R9158 gnd.n585 gnd.n584 9.3005
R9159 gnd.n6076 gnd.n6075 9.3005
R9160 gnd.n6077 gnd.n583 9.3005
R9161 gnd.n6079 gnd.n6078 9.3005
R9162 gnd.n579 gnd.n578 9.3005
R9163 gnd.n6086 gnd.n6085 9.3005
R9164 gnd.n6087 gnd.n577 9.3005
R9165 gnd.n6089 gnd.n6088 9.3005
R9166 gnd.n573 gnd.n572 9.3005
R9167 gnd.n6096 gnd.n6095 9.3005
R9168 gnd.n6097 gnd.n571 9.3005
R9169 gnd.n6099 gnd.n6098 9.3005
R9170 gnd.n567 gnd.n566 9.3005
R9171 gnd.n6106 gnd.n6105 9.3005
R9172 gnd.n6107 gnd.n565 9.3005
R9173 gnd.n6109 gnd.n6108 9.3005
R9174 gnd.n561 gnd.n560 9.3005
R9175 gnd.n6116 gnd.n6115 9.3005
R9176 gnd.n6117 gnd.n559 9.3005
R9177 gnd.n6119 gnd.n6118 9.3005
R9178 gnd.n555 gnd.n554 9.3005
R9179 gnd.n6126 gnd.n6125 9.3005
R9180 gnd.n6127 gnd.n553 9.3005
R9181 gnd.n6129 gnd.n6128 9.3005
R9182 gnd.n549 gnd.n548 9.3005
R9183 gnd.n6136 gnd.n6135 9.3005
R9184 gnd.n6137 gnd.n547 9.3005
R9185 gnd.n6139 gnd.n6138 9.3005
R9186 gnd.n543 gnd.n542 9.3005
R9187 gnd.n6146 gnd.n6145 9.3005
R9188 gnd.n6147 gnd.n541 9.3005
R9189 gnd.n6149 gnd.n6148 9.3005
R9190 gnd.n537 gnd.n536 9.3005
R9191 gnd.n6156 gnd.n6155 9.3005
R9192 gnd.n6157 gnd.n535 9.3005
R9193 gnd.n6159 gnd.n6158 9.3005
R9194 gnd.n531 gnd.n530 9.3005
R9195 gnd.n6166 gnd.n6165 9.3005
R9196 gnd.n6167 gnd.n529 9.3005
R9197 gnd.n6169 gnd.n6168 9.3005
R9198 gnd.n525 gnd.n524 9.3005
R9199 gnd.n6176 gnd.n6175 9.3005
R9200 gnd.n6177 gnd.n523 9.3005
R9201 gnd.n6179 gnd.n6178 9.3005
R9202 gnd.n519 gnd.n518 9.3005
R9203 gnd.n6186 gnd.n6185 9.3005
R9204 gnd.n6187 gnd.n517 9.3005
R9205 gnd.n6189 gnd.n6188 9.3005
R9206 gnd.n513 gnd.n512 9.3005
R9207 gnd.n6197 gnd.n6196 9.3005
R9208 gnd.n6198 gnd.n511 9.3005
R9209 gnd.n6200 gnd.n6199 9.3005
R9210 gnd.n5989 gnd.n5988 9.3005
R9211 gnd.n6758 gnd.n89 9.3005
R9212 gnd.n6757 gnd.n91 9.3005
R9213 gnd.n95 gnd.n92 9.3005
R9214 gnd.n6752 gnd.n96 9.3005
R9215 gnd.n6751 gnd.n97 9.3005
R9216 gnd.n6750 gnd.n98 9.3005
R9217 gnd.n102 gnd.n99 9.3005
R9218 gnd.n6745 gnd.n103 9.3005
R9219 gnd.n6744 gnd.n104 9.3005
R9220 gnd.n6743 gnd.n105 9.3005
R9221 gnd.n109 gnd.n106 9.3005
R9222 gnd.n6738 gnd.n110 9.3005
R9223 gnd.n6737 gnd.n111 9.3005
R9224 gnd.n6736 gnd.n112 9.3005
R9225 gnd.n116 gnd.n113 9.3005
R9226 gnd.n6731 gnd.n117 9.3005
R9227 gnd.n6730 gnd.n118 9.3005
R9228 gnd.n6726 gnd.n119 9.3005
R9229 gnd.n123 gnd.n120 9.3005
R9230 gnd.n6721 gnd.n124 9.3005
R9231 gnd.n6720 gnd.n125 9.3005
R9232 gnd.n6719 gnd.n126 9.3005
R9233 gnd.n130 gnd.n127 9.3005
R9234 gnd.n6714 gnd.n131 9.3005
R9235 gnd.n6713 gnd.n132 9.3005
R9236 gnd.n6712 gnd.n133 9.3005
R9237 gnd.n137 gnd.n134 9.3005
R9238 gnd.n6707 gnd.n138 9.3005
R9239 gnd.n6706 gnd.n139 9.3005
R9240 gnd.n6705 gnd.n140 9.3005
R9241 gnd.n144 gnd.n141 9.3005
R9242 gnd.n6700 gnd.n145 9.3005
R9243 gnd.n6699 gnd.n146 9.3005
R9244 gnd.n6698 gnd.n147 9.3005
R9245 gnd.n151 gnd.n148 9.3005
R9246 gnd.n6693 gnd.n152 9.3005
R9247 gnd.n6692 gnd.n6691 9.3005
R9248 gnd.n6690 gnd.n155 9.3005
R9249 gnd.n6760 gnd.n6759 9.3005
R9250 gnd.n6314 gnd.n463 9.3005
R9251 gnd.n6313 gnd.n465 9.3005
R9252 gnd.n6312 gnd.n466 9.3005
R9253 gnd.n486 gnd.n467 9.3005
R9254 gnd.n490 gnd.n489 9.3005
R9255 gnd.n491 gnd.n485 9.3005
R9256 gnd.n495 gnd.n492 9.3005
R9257 gnd.n496 gnd.n484 9.3005
R9258 gnd.n500 gnd.n499 9.3005
R9259 gnd.n501 gnd.n483 9.3005
R9260 gnd.n6219 gnd.n502 9.3005
R9261 gnd.n6220 gnd.n482 9.3005
R9262 gnd.n6224 gnd.n6223 9.3005
R9263 gnd.n6225 gnd.n481 9.3005
R9264 gnd.n6285 gnd.n6226 9.3005
R9265 gnd.n6284 gnd.n6227 9.3005
R9266 gnd.n6283 gnd.n6228 9.3005
R9267 gnd.n6282 gnd.n6229 9.3005
R9268 gnd.n6280 gnd.n6230 9.3005
R9269 gnd.n6279 gnd.n6231 9.3005
R9270 gnd.n6278 gnd.n239 9.3005
R9271 gnd.n6276 gnd.n6232 9.3005
R9272 gnd.n6275 gnd.n6233 9.3005
R9273 gnd.n6273 gnd.n6234 9.3005
R9274 gnd.n6272 gnd.n6235 9.3005
R9275 gnd.n6270 gnd.n6236 9.3005
R9276 gnd.n6269 gnd.n6237 9.3005
R9277 gnd.n6267 gnd.n6238 9.3005
R9278 gnd.n6266 gnd.n6239 9.3005
R9279 gnd.n6264 gnd.n6240 9.3005
R9280 gnd.n6263 gnd.n6241 9.3005
R9281 gnd.n6261 gnd.n6242 9.3005
R9282 gnd.n6260 gnd.n6243 9.3005
R9283 gnd.n6258 gnd.n6244 9.3005
R9284 gnd.n6257 gnd.n6245 9.3005
R9285 gnd.n6255 gnd.n6246 9.3005
R9286 gnd.n6254 gnd.n6247 9.3005
R9287 gnd.n6252 gnd.n6248 9.3005
R9288 gnd.n6251 gnd.n6250 9.3005
R9289 gnd.n6249 gnd.n159 9.3005
R9290 gnd.n6687 gnd.n158 9.3005
R9291 gnd.n6689 gnd.n6688 9.3005
R9292 gnd.n6316 gnd.n6315 9.3005
R9293 gnd.n6322 gnd.n6321 9.3005
R9294 gnd.n6323 gnd.n457 9.3005
R9295 gnd.n6326 gnd.n456 9.3005
R9296 gnd.n6327 gnd.n455 9.3005
R9297 gnd.n6330 gnd.n454 9.3005
R9298 gnd.n6331 gnd.n453 9.3005
R9299 gnd.n6334 gnd.n452 9.3005
R9300 gnd.n6335 gnd.n451 9.3005
R9301 gnd.n6338 gnd.n450 9.3005
R9302 gnd.n6339 gnd.n449 9.3005
R9303 gnd.n6342 gnd.n448 9.3005
R9304 gnd.n6343 gnd.n447 9.3005
R9305 gnd.n6346 gnd.n446 9.3005
R9306 gnd.n6347 gnd.n445 9.3005
R9307 gnd.n6350 gnd.n444 9.3005
R9308 gnd.n6351 gnd.n443 9.3005
R9309 gnd.n6354 gnd.n442 9.3005
R9310 gnd.n6355 gnd.n441 9.3005
R9311 gnd.n6358 gnd.n440 9.3005
R9312 gnd.n6360 gnd.n434 9.3005
R9313 gnd.n6363 gnd.n433 9.3005
R9314 gnd.n6364 gnd.n432 9.3005
R9315 gnd.n6367 gnd.n431 9.3005
R9316 gnd.n6368 gnd.n430 9.3005
R9317 gnd.n6371 gnd.n429 9.3005
R9318 gnd.n6372 gnd.n428 9.3005
R9319 gnd.n6375 gnd.n427 9.3005
R9320 gnd.n6376 gnd.n426 9.3005
R9321 gnd.n6379 gnd.n425 9.3005
R9322 gnd.n6380 gnd.n424 9.3005
R9323 gnd.n6383 gnd.n423 9.3005
R9324 gnd.n6385 gnd.n422 9.3005
R9325 gnd.n6386 gnd.n421 9.3005
R9326 gnd.n6387 gnd.n420 9.3005
R9327 gnd.n419 gnd.n326 9.3005
R9328 gnd.n6320 gnd.n462 9.3005
R9329 gnd.n6319 gnd.n6318 9.3005
R9330 gnd.n6449 gnd.n325 9.3005
R9331 gnd.n6451 gnd.n6450 9.3005
R9332 gnd.n310 gnd.n309 9.3005
R9333 gnd.n6464 gnd.n6463 9.3005
R9334 gnd.n6465 gnd.n308 9.3005
R9335 gnd.n6467 gnd.n6466 9.3005
R9336 gnd.n292 gnd.n291 9.3005
R9337 gnd.n6480 gnd.n6479 9.3005
R9338 gnd.n6481 gnd.n290 9.3005
R9339 gnd.n6483 gnd.n6482 9.3005
R9340 gnd.n275 gnd.n274 9.3005
R9341 gnd.n6496 gnd.n6495 9.3005
R9342 gnd.n6497 gnd.n273 9.3005
R9343 gnd.n6500 gnd.n6498 9.3005
R9344 gnd.n6499 gnd.n212 9.3005
R9345 gnd.n6558 gnd.n211 9.3005
R9346 gnd.n6560 gnd.n6559 9.3005
R9347 gnd.n199 gnd.n198 9.3005
R9348 gnd.n6573 gnd.n6572 9.3005
R9349 gnd.n6574 gnd.n197 9.3005
R9350 gnd.n6576 gnd.n6575 9.3005
R9351 gnd.n183 gnd.n182 9.3005
R9352 gnd.n6589 gnd.n6588 9.3005
R9353 gnd.n6590 gnd.n181 9.3005
R9354 gnd.n6592 gnd.n6591 9.3005
R9355 gnd.n166 gnd.n165 9.3005
R9356 gnd.n6679 gnd.n6678 9.3005
R9357 gnd.n6680 gnd.n164 9.3005
R9358 gnd.n6682 gnd.n6681 9.3005
R9359 gnd.n88 gnd.n87 9.3005
R9360 gnd.n6762 gnd.n6761 9.3005
R9361 gnd.n6448 gnd.n6447 9.3005
R9362 gnd.n6557 gnd.n6556 9.3005
R9363 gnd.n6207 gnd.n6206 9.3005
R9364 gnd.n4039 gnd.n4038 9.3005
R9365 gnd.n4040 gnd.n4033 9.3005
R9366 gnd.n4042 gnd.n4041 9.3005
R9367 gnd.n2011 gnd.n2010 9.3005
R9368 gnd.n4047 gnd.n4046 9.3005
R9369 gnd.n4048 gnd.n2009 9.3005
R9370 gnd.n4054 gnd.n4049 9.3005
R9371 gnd.n4053 gnd.n4050 9.3005
R9372 gnd.n4052 gnd.n4051 9.3005
R9373 gnd.n1990 gnd.n1989 9.3005
R9374 gnd.n4167 gnd.n4166 9.3005
R9375 gnd.n4168 gnd.n1988 9.3005
R9376 gnd.n4170 gnd.n4169 9.3005
R9377 gnd.n1986 gnd.n1985 9.3005
R9378 gnd.n4175 gnd.n4174 9.3005
R9379 gnd.n4176 gnd.n1984 9.3005
R9380 gnd.n4183 gnd.n4177 9.3005
R9381 gnd.n4182 gnd.n4178 9.3005
R9382 gnd.n4181 gnd.n4179 9.3005
R9383 gnd.n1845 gnd.n1844 9.3005
R9384 gnd.n4237 gnd.n4236 9.3005
R9385 gnd.n4238 gnd.n1843 9.3005
R9386 gnd.n4249 gnd.n4239 9.3005
R9387 gnd.n4248 gnd.n4240 9.3005
R9388 gnd.n4247 gnd.n4241 9.3005
R9389 gnd.n4244 gnd.n4243 9.3005
R9390 gnd.n4242 gnd.n1215 9.3005
R9391 gnd.n5330 gnd.n1216 9.3005
R9392 gnd.n5329 gnd.n1217 9.3005
R9393 gnd.n5328 gnd.n1218 9.3005
R9394 gnd.n1316 gnd.n1219 9.3005
R9395 gnd.n1317 gnd.n1315 9.3005
R9396 gnd.n5311 gnd.n1318 9.3005
R9397 gnd.n5310 gnd.n1319 9.3005
R9398 gnd.n5309 gnd.n1320 9.3005
R9399 gnd.n4433 gnd.n1321 9.3005
R9400 gnd.n4434 gnd.n4432 9.3005
R9401 gnd.n4436 gnd.n4435 9.3005
R9402 gnd.n1803 gnd.n1802 9.3005
R9403 gnd.n4462 gnd.n4461 9.3005
R9404 gnd.n4463 gnd.n1801 9.3005
R9405 gnd.n4476 gnd.n4464 9.3005
R9406 gnd.n4475 gnd.n4465 9.3005
R9407 gnd.n4474 gnd.n4466 9.3005
R9408 gnd.n4468 gnd.n4467 9.3005
R9409 gnd.n4470 gnd.n4469 9.3005
R9410 gnd.n1765 gnd.n1764 9.3005
R9411 gnd.n4520 gnd.n4519 9.3005
R9412 gnd.n4521 gnd.n1763 9.3005
R9413 gnd.n4523 gnd.n4522 9.3005
R9414 gnd.n1747 gnd.n1746 9.3005
R9415 gnd.n4546 gnd.n4545 9.3005
R9416 gnd.n4547 gnd.n1745 9.3005
R9417 gnd.n4551 gnd.n4548 9.3005
R9418 gnd.n4550 gnd.n4549 9.3005
R9419 gnd.n1723 gnd.n1722 9.3005
R9420 gnd.n4585 gnd.n4584 9.3005
R9421 gnd.n4586 gnd.n1721 9.3005
R9422 gnd.n4599 gnd.n4587 9.3005
R9423 gnd.n4598 gnd.n4588 9.3005
R9424 gnd.n4597 gnd.n4589 9.3005
R9425 gnd.n4591 gnd.n4590 9.3005
R9426 gnd.n4593 gnd.n4592 9.3005
R9427 gnd.n1684 gnd.n1683 9.3005
R9428 gnd.n4643 gnd.n4642 9.3005
R9429 gnd.n4644 gnd.n1682 9.3005
R9430 gnd.n4646 gnd.n4645 9.3005
R9431 gnd.n1665 gnd.n1664 9.3005
R9432 gnd.n4668 gnd.n4667 9.3005
R9433 gnd.n4669 gnd.n1663 9.3005
R9434 gnd.n4673 gnd.n4670 9.3005
R9435 gnd.n4672 gnd.n4671 9.3005
R9436 gnd.n1640 gnd.n1639 9.3005
R9437 gnd.n4707 gnd.n4706 9.3005
R9438 gnd.n4708 gnd.n1638 9.3005
R9439 gnd.n4710 gnd.n4709 9.3005
R9440 gnd.n1617 gnd.n1616 9.3005
R9441 gnd.n4753 gnd.n4752 9.3005
R9442 gnd.n4754 gnd.n1615 9.3005
R9443 gnd.n4758 gnd.n4755 9.3005
R9444 gnd.n4757 gnd.n4756 9.3005
R9445 gnd.n1596 gnd.n1595 9.3005
R9446 gnd.n4808 gnd.n4807 9.3005
R9447 gnd.n4809 gnd.n1594 9.3005
R9448 gnd.n4813 gnd.n4810 9.3005
R9449 gnd.n4812 gnd.n4811 9.3005
R9450 gnd.n1569 gnd.n1568 9.3005
R9451 gnd.n4845 gnd.n4844 9.3005
R9452 gnd.n4846 gnd.n1567 9.3005
R9453 gnd.n4848 gnd.n4847 9.3005
R9454 gnd.n1551 gnd.n1550 9.3005
R9455 gnd.n4871 gnd.n4870 9.3005
R9456 gnd.n4872 gnd.n1549 9.3005
R9457 gnd.n4876 gnd.n4873 9.3005
R9458 gnd.n4875 gnd.n4874 9.3005
R9459 gnd.n1523 gnd.n1522 9.3005
R9460 gnd.n4924 gnd.n4923 9.3005
R9461 gnd.n4925 gnd.n1521 9.3005
R9462 gnd.n4927 gnd.n4926 9.3005
R9463 gnd.n1431 gnd.n1430 9.3005
R9464 gnd.n5067 gnd.n5066 9.3005
R9465 gnd.n5068 gnd.n1429 9.3005
R9466 gnd.n5187 gnd.n5069 9.3005
R9467 gnd.n5186 gnd.n5070 9.3005
R9468 gnd.n5185 gnd.n5071 9.3005
R9469 gnd.n5184 gnd.n5072 9.3005
R9470 gnd.n5112 gnd.n5073 9.3005
R9471 gnd.n5113 gnd.n5111 9.3005
R9472 gnd.n5115 gnd.n5114 9.3005
R9473 gnd.n5110 gnd.n5109 9.3005
R9474 gnd.n5120 gnd.n5119 9.3005
R9475 gnd.n5121 gnd.n5108 9.3005
R9476 gnd.n5147 gnd.n5122 9.3005
R9477 gnd.n5146 gnd.n5123 9.3005
R9478 gnd.n5145 gnd.n5124 9.3005
R9479 gnd.n5127 gnd.n5125 9.3005
R9480 gnd.n5141 gnd.n5128 9.3005
R9481 gnd.n5140 gnd.n5129 9.3005
R9482 gnd.n5139 gnd.n5130 9.3005
R9483 gnd.n5132 gnd.n5131 9.3005
R9484 gnd.n5135 gnd.n5134 9.3005
R9485 gnd.n5133 gnd.n505 9.3005
R9486 gnd.n6214 gnd.n506 9.3005
R9487 gnd.n6213 gnd.n507 9.3005
R9488 gnd.n6212 gnd.n508 9.3005
R9489 gnd.n6204 gnd.n509 9.3005
R9490 gnd.n6208 gnd.n6205 9.3005
R9491 gnd.n3671 gnd.n3670 9.3005
R9492 gnd.n3701 gnd.n3648 9.3005
R9493 gnd.n3700 gnd.n3649 9.3005
R9494 gnd.n3698 gnd.n3650 9.3005
R9495 gnd.n3697 gnd.n3651 9.3005
R9496 gnd.n3695 gnd.n3652 9.3005
R9497 gnd.n3694 gnd.n3653 9.3005
R9498 gnd.n3692 gnd.n3654 9.3005
R9499 gnd.n3691 gnd.n3655 9.3005
R9500 gnd.n3689 gnd.n3656 9.3005
R9501 gnd.n3688 gnd.n3657 9.3005
R9502 gnd.n3686 gnd.n3658 9.3005
R9503 gnd.n3685 gnd.n3659 9.3005
R9504 gnd.n3683 gnd.n3660 9.3005
R9505 gnd.n3682 gnd.n3661 9.3005
R9506 gnd.n3680 gnd.n3662 9.3005
R9507 gnd.n3679 gnd.n3663 9.3005
R9508 gnd.n3677 gnd.n3664 9.3005
R9509 gnd.n3676 gnd.n3665 9.3005
R9510 gnd.n3674 gnd.n3666 9.3005
R9511 gnd.n3673 gnd.n3667 9.3005
R9512 gnd.n3703 gnd.n3702 9.3005
R9513 gnd.n3646 gnd.n3645 9.3005
R9514 gnd.n3642 gnd.n3602 9.3005
R9515 gnd.n3641 gnd.n3638 9.3005
R9516 gnd.n3637 gnd.n3603 9.3005
R9517 gnd.n3636 gnd.n3635 9.3005
R9518 gnd.n3632 gnd.n3604 9.3005
R9519 gnd.n3631 gnd.n3628 9.3005
R9520 gnd.n3627 gnd.n3605 9.3005
R9521 gnd.n3626 gnd.n3625 9.3005
R9522 gnd.n3622 gnd.n3606 9.3005
R9523 gnd.n3621 gnd.n3618 9.3005
R9524 gnd.n3617 gnd.n3607 9.3005
R9525 gnd.n3616 gnd.n3615 9.3005
R9526 gnd.n3612 gnd.n3608 9.3005
R9527 gnd.n3611 gnd.n3609 9.3005
R9528 gnd.n2118 gnd.n2117 9.3005
R9529 gnd.n3882 gnd.n3881 9.3005
R9530 gnd.n3647 gnd.n3601 9.3005
R9531 gnd.n3705 gnd.n3704 9.3005
R9532 gnd.n3885 gnd.n3884 9.3005
R9533 gnd.n2102 gnd.n2101 9.3005
R9534 gnd.n3898 gnd.n3897 9.3005
R9535 gnd.n3899 gnd.n2100 9.3005
R9536 gnd.n3901 gnd.n3900 9.3005
R9537 gnd.n2086 gnd.n2085 9.3005
R9538 gnd.n3914 gnd.n3913 9.3005
R9539 gnd.n3915 gnd.n2084 9.3005
R9540 gnd.n3917 gnd.n3916 9.3005
R9541 gnd.n2070 gnd.n2069 9.3005
R9542 gnd.n3930 gnd.n3929 9.3005
R9543 gnd.n3931 gnd.n2068 9.3005
R9544 gnd.n3933 gnd.n3932 9.3005
R9545 gnd.n2054 gnd.n2053 9.3005
R9546 gnd.n3947 gnd.n3946 9.3005
R9547 gnd.n3948 gnd.n2052 9.3005
R9548 gnd.n3954 gnd.n3949 9.3005
R9549 gnd.n3953 gnd.n3950 9.3005
R9550 gnd.n3952 gnd.n3951 9.3005
R9551 gnd.n2036 gnd.n2035 9.3005
R9552 gnd.n3989 gnd.n3978 9.3005
R9553 gnd.n3988 gnd.n3979 9.3005
R9554 gnd.n3987 gnd.n3980 9.3005
R9555 gnd.n3986 gnd.n3981 9.3005
R9556 gnd.n3984 gnd.n3983 9.3005
R9557 gnd.n3982 gnd.n1015 9.3005
R9558 gnd.n5485 gnd.n1016 9.3005
R9559 gnd.n5484 gnd.n1017 9.3005
R9560 gnd.n5483 gnd.n1018 9.3005
R9561 gnd.n1037 gnd.n1019 9.3005
R9562 gnd.n5473 gnd.n1038 9.3005
R9563 gnd.n5472 gnd.n1039 9.3005
R9564 gnd.n5471 gnd.n1040 9.3005
R9565 gnd.n1057 gnd.n1041 9.3005
R9566 gnd.n5461 gnd.n1058 9.3005
R9567 gnd.n5460 gnd.n1059 9.3005
R9568 gnd.n5459 gnd.n1060 9.3005
R9569 gnd.n1079 gnd.n1061 9.3005
R9570 gnd.n5449 gnd.n1080 9.3005
R9571 gnd.n5448 gnd.n1081 9.3005
R9572 gnd.n5447 gnd.n1082 9.3005
R9573 gnd.n1908 gnd.n1083 9.3005
R9574 gnd.n3883 gnd.n2116 9.3005
R9575 gnd.n5409 gnd.n1139 9.3005
R9576 gnd.n5412 gnd.n1138 9.3005
R9577 gnd.n5413 gnd.n1137 9.3005
R9578 gnd.n5416 gnd.n1136 9.3005
R9579 gnd.n5417 gnd.n1135 9.3005
R9580 gnd.n5420 gnd.n1134 9.3005
R9581 gnd.n5421 gnd.n1133 9.3005
R9582 gnd.n5424 gnd.n1132 9.3005
R9583 gnd.n5425 gnd.n1131 9.3005
R9584 gnd.n5428 gnd.n1130 9.3005
R9585 gnd.n5429 gnd.n1129 9.3005
R9586 gnd.n5432 gnd.n1128 9.3005
R9587 gnd.n5433 gnd.n1127 9.3005
R9588 gnd.n5434 gnd.n1126 9.3005
R9589 gnd.n1093 gnd.n1092 9.3005
R9590 gnd.n5440 gnd.n5439 9.3005
R9591 gnd.n4096 gnd.n4094 9.3005
R9592 gnd.n4098 gnd.n4097 9.3005
R9593 gnd.n4101 gnd.n4091 9.3005
R9594 gnd.n4105 gnd.n4104 9.3005
R9595 gnd.n4106 gnd.n4090 9.3005
R9596 gnd.n4108 gnd.n4107 9.3005
R9597 gnd.n4111 gnd.n4089 9.3005
R9598 gnd.n4115 gnd.n4114 9.3005
R9599 gnd.n4116 gnd.n4088 9.3005
R9600 gnd.n4118 gnd.n4117 9.3005
R9601 gnd.n4121 gnd.n4087 9.3005
R9602 gnd.n4125 gnd.n4124 9.3005
R9603 gnd.n4126 gnd.n4086 9.3005
R9604 gnd.n4128 gnd.n4127 9.3005
R9605 gnd.n4131 gnd.n4085 9.3005
R9606 gnd.n4135 gnd.n4134 9.3005
R9607 gnd.n4136 gnd.n4084 9.3005
R9608 gnd.n4139 gnd.n4137 9.3005
R9609 gnd.n4140 gnd.n4080 9.3005
R9610 gnd.n4143 gnd.n4142 9.3005
R9611 gnd.n4095 gnd.n1140 9.3005
R9612 gnd.n3797 gnd.n3796 9.3005
R9613 gnd.n3795 gnd.n3754 9.3005
R9614 gnd.n3794 gnd.n3793 9.3005
R9615 gnd.n3792 gnd.n3755 9.3005
R9616 gnd.n3790 gnd.n3756 9.3005
R9617 gnd.n3789 gnd.n3757 9.3005
R9618 gnd.n3787 gnd.n3758 9.3005
R9619 gnd.n3786 gnd.n3759 9.3005
R9620 gnd.n3784 gnd.n3760 9.3005
R9621 gnd.n3783 gnd.n3761 9.3005
R9622 gnd.n3781 gnd.n3762 9.3005
R9623 gnd.n3780 gnd.n3763 9.3005
R9624 gnd.n3778 gnd.n3764 9.3005
R9625 gnd.n3777 gnd.n3765 9.3005
R9626 gnd.n3775 gnd.n3766 9.3005
R9627 gnd.n3774 gnd.n3767 9.3005
R9628 gnd.n3772 gnd.n3768 9.3005
R9629 gnd.n3771 gnd.n3770 9.3005
R9630 gnd.n3769 gnd.n2039 9.3005
R9631 gnd.n3967 gnd.n2037 9.3005
R9632 gnd.n3977 gnd.n3976 9.3005
R9633 gnd.n3975 gnd.n2038 9.3005
R9634 gnd.n3973 gnd.n3968 9.3005
R9635 gnd.n3972 gnd.n3970 9.3005
R9636 gnd.n3969 gnd.n2018 9.3005
R9637 gnd.n4010 gnd.n2019 9.3005
R9638 gnd.n4011 gnd.n2017 9.3005
R9639 gnd.n4013 gnd.n4012 9.3005
R9640 gnd.n4014 gnd.n2016 9.3005
R9641 gnd.n4020 gnd.n4015 9.3005
R9642 gnd.n4019 gnd.n4016 9.3005
R9643 gnd.n4018 gnd.n4017 9.3005
R9644 gnd.n2002 gnd.n2001 9.3005
R9645 gnd.n4068 gnd.n4067 9.3005
R9646 gnd.n4069 gnd.n2000 9.3005
R9647 gnd.n4071 gnd.n4070 9.3005
R9648 gnd.n4072 gnd.n1999 9.3005
R9649 gnd.n4076 gnd.n4075 9.3005
R9650 gnd.n4077 gnd.n1998 9.3005
R9651 gnd.n4147 gnd.n4078 9.3005
R9652 gnd.n4146 gnd.n4079 9.3005
R9653 gnd.n4145 gnd.n4144 9.3005
R9654 gnd.n3798 gnd.n3752 9.3005
R9655 gnd.n3805 gnd.n3804 9.3005
R9656 gnd.n3806 gnd.n3746 9.3005
R9657 gnd.n3809 gnd.n3745 9.3005
R9658 gnd.n3810 gnd.n3744 9.3005
R9659 gnd.n3813 gnd.n3743 9.3005
R9660 gnd.n3814 gnd.n3742 9.3005
R9661 gnd.n3817 gnd.n3741 9.3005
R9662 gnd.n3818 gnd.n3740 9.3005
R9663 gnd.n3821 gnd.n3739 9.3005
R9664 gnd.n3822 gnd.n3738 9.3005
R9665 gnd.n3825 gnd.n3737 9.3005
R9666 gnd.n3826 gnd.n3736 9.3005
R9667 gnd.n3829 gnd.n3735 9.3005
R9668 gnd.n3830 gnd.n3734 9.3005
R9669 gnd.n3833 gnd.n3733 9.3005
R9670 gnd.n3834 gnd.n3732 9.3005
R9671 gnd.n3837 gnd.n3731 9.3005
R9672 gnd.n3838 gnd.n3730 9.3005
R9673 gnd.n3841 gnd.n3729 9.3005
R9674 gnd.n3843 gnd.n3726 9.3005
R9675 gnd.n3846 gnd.n3725 9.3005
R9676 gnd.n3847 gnd.n3724 9.3005
R9677 gnd.n3850 gnd.n3723 9.3005
R9678 gnd.n3851 gnd.n3722 9.3005
R9679 gnd.n3854 gnd.n3721 9.3005
R9680 gnd.n3855 gnd.n3720 9.3005
R9681 gnd.n3858 gnd.n3719 9.3005
R9682 gnd.n3859 gnd.n3718 9.3005
R9683 gnd.n3862 gnd.n3717 9.3005
R9684 gnd.n3863 gnd.n3716 9.3005
R9685 gnd.n3866 gnd.n3715 9.3005
R9686 gnd.n3867 gnd.n3714 9.3005
R9687 gnd.n3870 gnd.n3713 9.3005
R9688 gnd.n3872 gnd.n3712 9.3005
R9689 gnd.n3873 gnd.n3711 9.3005
R9690 gnd.n3874 gnd.n3710 9.3005
R9691 gnd.n3875 gnd.n3709 9.3005
R9692 gnd.n3803 gnd.n3751 9.3005
R9693 gnd.n3802 gnd.n3801 9.3005
R9694 gnd.n3890 gnd.n3889 9.3005
R9695 gnd.n3891 gnd.n2108 9.3005
R9696 gnd.n3893 gnd.n3892 9.3005
R9697 gnd.n2093 gnd.n2092 9.3005
R9698 gnd.n3906 gnd.n3905 9.3005
R9699 gnd.n3907 gnd.n2091 9.3005
R9700 gnd.n3909 gnd.n3908 9.3005
R9701 gnd.n2078 gnd.n2077 9.3005
R9702 gnd.n3922 gnd.n3921 9.3005
R9703 gnd.n3923 gnd.n2076 9.3005
R9704 gnd.n3925 gnd.n3924 9.3005
R9705 gnd.n2061 gnd.n2060 9.3005
R9706 gnd.n3938 gnd.n3937 9.3005
R9707 gnd.n3939 gnd.n2059 9.3005
R9708 gnd.n3942 gnd.n3940 9.3005
R9709 gnd.n5489 gnd.n1007 9.3005
R9710 gnd.n1026 gnd.n1008 9.3005
R9711 gnd.n5479 gnd.n1027 9.3005
R9712 gnd.n5478 gnd.n1028 9.3005
R9713 gnd.n5477 gnd.n1029 9.3005
R9714 gnd.n1047 gnd.n1030 9.3005
R9715 gnd.n5467 gnd.n1048 9.3005
R9716 gnd.n5466 gnd.n1049 9.3005
R9717 gnd.n5465 gnd.n1050 9.3005
R9718 gnd.n1068 gnd.n1051 9.3005
R9719 gnd.n5455 gnd.n1069 9.3005
R9720 gnd.n5454 gnd.n1070 9.3005
R9721 gnd.n5453 gnd.n1071 9.3005
R9722 gnd.n1090 gnd.n1072 9.3005
R9723 gnd.n5443 gnd.n1091 9.3005
R9724 gnd.n5442 gnd.n5441 9.3005
R9725 gnd.n2110 gnd.n2109 9.3005
R9726 gnd.n5490 gnd.n1006 9.3005
R9727 gnd.n4036 gnd.n4035 9.3005
R9728 gnd.n5497 gnd.n995 9.3005
R9729 gnd.n5498 gnd.n994 9.3005
R9730 gnd.n993 gnd.n989 9.3005
R9731 gnd.n5504 gnd.n988 9.3005
R9732 gnd.n5505 gnd.n987 9.3005
R9733 gnd.n5506 gnd.n986 9.3005
R9734 gnd.n985 gnd.n981 9.3005
R9735 gnd.n5512 gnd.n980 9.3005
R9736 gnd.n5513 gnd.n979 9.3005
R9737 gnd.n5514 gnd.n978 9.3005
R9738 gnd.n977 gnd.n973 9.3005
R9739 gnd.n5520 gnd.n972 9.3005
R9740 gnd.n5521 gnd.n971 9.3005
R9741 gnd.n5522 gnd.n970 9.3005
R9742 gnd.n969 gnd.n965 9.3005
R9743 gnd.n5528 gnd.n964 9.3005
R9744 gnd.n5529 gnd.n963 9.3005
R9745 gnd.n5530 gnd.n962 9.3005
R9746 gnd.n961 gnd.n957 9.3005
R9747 gnd.n5536 gnd.n956 9.3005
R9748 gnd.n5537 gnd.n955 9.3005
R9749 gnd.n5538 gnd.n954 9.3005
R9750 gnd.n953 gnd.n949 9.3005
R9751 gnd.n5544 gnd.n948 9.3005
R9752 gnd.n5545 gnd.n947 9.3005
R9753 gnd.n5546 gnd.n946 9.3005
R9754 gnd.n945 gnd.n941 9.3005
R9755 gnd.n5552 gnd.n940 9.3005
R9756 gnd.n5553 gnd.n939 9.3005
R9757 gnd.n5554 gnd.n938 9.3005
R9758 gnd.n937 gnd.n933 9.3005
R9759 gnd.n5560 gnd.n932 9.3005
R9760 gnd.n5561 gnd.n931 9.3005
R9761 gnd.n5562 gnd.n930 9.3005
R9762 gnd.n929 gnd.n925 9.3005
R9763 gnd.n5568 gnd.n924 9.3005
R9764 gnd.n5569 gnd.n923 9.3005
R9765 gnd.n5570 gnd.n922 9.3005
R9766 gnd.n921 gnd.n917 9.3005
R9767 gnd.n5576 gnd.n916 9.3005
R9768 gnd.n5577 gnd.n915 9.3005
R9769 gnd.n5578 gnd.n914 9.3005
R9770 gnd.n913 gnd.n909 9.3005
R9771 gnd.n5584 gnd.n908 9.3005
R9772 gnd.n5585 gnd.n907 9.3005
R9773 gnd.n5586 gnd.n906 9.3005
R9774 gnd.n905 gnd.n901 9.3005
R9775 gnd.n5592 gnd.n900 9.3005
R9776 gnd.n5593 gnd.n899 9.3005
R9777 gnd.n5594 gnd.n898 9.3005
R9778 gnd.n897 gnd.n893 9.3005
R9779 gnd.n5600 gnd.n892 9.3005
R9780 gnd.n5601 gnd.n891 9.3005
R9781 gnd.n5602 gnd.n890 9.3005
R9782 gnd.n889 gnd.n885 9.3005
R9783 gnd.n5608 gnd.n884 9.3005
R9784 gnd.n5609 gnd.n883 9.3005
R9785 gnd.n5610 gnd.n882 9.3005
R9786 gnd.n881 gnd.n877 9.3005
R9787 gnd.n5616 gnd.n876 9.3005
R9788 gnd.n5617 gnd.n875 9.3005
R9789 gnd.n5618 gnd.n874 9.3005
R9790 gnd.n873 gnd.n869 9.3005
R9791 gnd.n5624 gnd.n868 9.3005
R9792 gnd.n5625 gnd.n867 9.3005
R9793 gnd.n5626 gnd.n866 9.3005
R9794 gnd.n865 gnd.n861 9.3005
R9795 gnd.n5632 gnd.n860 9.3005
R9796 gnd.n5633 gnd.n859 9.3005
R9797 gnd.n5634 gnd.n858 9.3005
R9798 gnd.n857 gnd.n853 9.3005
R9799 gnd.n5640 gnd.n852 9.3005
R9800 gnd.n5641 gnd.n851 9.3005
R9801 gnd.n5642 gnd.n850 9.3005
R9802 gnd.n849 gnd.n845 9.3005
R9803 gnd.n5648 gnd.n844 9.3005
R9804 gnd.n5649 gnd.n843 9.3005
R9805 gnd.n5650 gnd.n842 9.3005
R9806 gnd.n841 gnd.n837 9.3005
R9807 gnd.n5656 gnd.n836 9.3005
R9808 gnd.n5657 gnd.n835 9.3005
R9809 gnd.n5658 gnd.n834 9.3005
R9810 gnd.n830 gnd.n829 9.3005
R9811 gnd.n5665 gnd.n5664 9.3005
R9812 gnd.n5496 gnd.n996 9.3005
R9813 gnd.n6435 gnd.n6434 9.3005
R9814 gnd.n340 gnd.n339 9.3005
R9815 gnd.n6429 gnd.n6428 9.3005
R9816 gnd.n6427 gnd.n6426 9.3005
R9817 gnd.n348 gnd.n347 9.3005
R9818 gnd.n6421 gnd.n6420 9.3005
R9819 gnd.n6419 gnd.n6418 9.3005
R9820 gnd.n356 gnd.n355 9.3005
R9821 gnd.n6413 gnd.n6412 9.3005
R9822 gnd.n6411 gnd.n6410 9.3005
R9823 gnd.n364 gnd.n363 9.3005
R9824 gnd.n6405 gnd.n6404 9.3005
R9825 gnd.n6403 gnd.n6402 9.3005
R9826 gnd.n372 gnd.n371 9.3005
R9827 gnd.n6397 gnd.n6396 9.3005
R9828 gnd.n6395 gnd.n6394 9.3005
R9829 gnd.n382 gnd.n381 9.3005
R9830 gnd.n5104 gnd.n5103 9.3005
R9831 gnd.n6437 gnd.n6436 9.3005
R9832 gnd.n6399 gnd.n6398 9.3005
R9833 gnd.n6401 gnd.n6400 9.3005
R9834 gnd.n368 gnd.n367 9.3005
R9835 gnd.n6407 gnd.n6406 9.3005
R9836 gnd.n6409 gnd.n6408 9.3005
R9837 gnd.n360 gnd.n359 9.3005
R9838 gnd.n6415 gnd.n6414 9.3005
R9839 gnd.n6417 gnd.n6416 9.3005
R9840 gnd.n352 gnd.n351 9.3005
R9841 gnd.n6423 gnd.n6422 9.3005
R9842 gnd.n6425 gnd.n6424 9.3005
R9843 gnd.n344 gnd.n343 9.3005
R9844 gnd.n6431 gnd.n6430 9.3005
R9845 gnd.n6433 gnd.n6432 9.3005
R9846 gnd.n336 gnd.n335 9.3005
R9847 gnd.n6439 gnd.n6438 9.3005
R9848 gnd.n378 gnd.n377 9.3005
R9849 gnd.n6393 gnd.n6392 9.3005
R9850 gnd.n5157 gnd.n5156 9.3005
R9851 gnd.n5160 gnd.n5100 9.3005
R9852 gnd.n5164 gnd.n5163 9.3005
R9853 gnd.n5165 gnd.n5099 9.3005
R9854 gnd.n5167 gnd.n5166 9.3005
R9855 gnd.n5170 gnd.n5096 9.3005
R9856 gnd.n5174 gnd.n5173 9.3005
R9857 gnd.n5175 gnd.n5094 9.3005
R9858 gnd.n5177 gnd.n5176 9.3005
R9859 gnd.n5095 gnd.n1416 9.3005
R9860 gnd.n4228 gnd.n4217 9.3005
R9861 gnd.n4227 gnd.n4226 9.3005
R9862 gnd.n4225 gnd.n4220 9.3005
R9863 gnd.n4224 gnd.n4223 9.3005
R9864 gnd.n1830 gnd.n1829 9.3005
R9865 gnd.n4276 gnd.n4275 9.3005
R9866 gnd.n4277 gnd.n1827 9.3005
R9867 gnd.n4282 gnd.n4281 9.3005
R9868 gnd.n4280 gnd.n1828 9.3005
R9869 gnd.n4279 gnd.n4278 9.3005
R9870 gnd.n1330 gnd.n1328 9.3005
R9871 gnd.n5305 gnd.n5304 9.3005
R9872 gnd.n5303 gnd.n1329 9.3005
R9873 gnd.n5302 gnd.n5301 9.3005
R9874 gnd.n5300 gnd.n1331 9.3005
R9875 gnd.n5299 gnd.n5298 9.3005
R9876 gnd.n5297 gnd.n1335 9.3005
R9877 gnd.n5296 gnd.n5295 9.3005
R9878 gnd.n5294 gnd.n1336 9.3005
R9879 gnd.n5293 gnd.n5292 9.3005
R9880 gnd.n5291 gnd.n1340 9.3005
R9881 gnd.n5290 gnd.n5289 9.3005
R9882 gnd.n5288 gnd.n1341 9.3005
R9883 gnd.n5287 gnd.n5286 9.3005
R9884 gnd.n5285 gnd.n1345 9.3005
R9885 gnd.n5284 gnd.n5283 9.3005
R9886 gnd.n5282 gnd.n1346 9.3005
R9887 gnd.n5281 gnd.n5280 9.3005
R9888 gnd.n5279 gnd.n1350 9.3005
R9889 gnd.n5278 gnd.n5277 9.3005
R9890 gnd.n5276 gnd.n1351 9.3005
R9891 gnd.n5275 gnd.n5274 9.3005
R9892 gnd.n5273 gnd.n1355 9.3005
R9893 gnd.n5272 gnd.n5271 9.3005
R9894 gnd.n5270 gnd.n1356 9.3005
R9895 gnd.n5269 gnd.n5268 9.3005
R9896 gnd.n5267 gnd.n1360 9.3005
R9897 gnd.n5266 gnd.n5265 9.3005
R9898 gnd.n5264 gnd.n1361 9.3005
R9899 gnd.n5263 gnd.n5262 9.3005
R9900 gnd.n5261 gnd.n1365 9.3005
R9901 gnd.n5260 gnd.n5259 9.3005
R9902 gnd.n5258 gnd.n1366 9.3005
R9903 gnd.n5257 gnd.n5256 9.3005
R9904 gnd.n5255 gnd.n1370 9.3005
R9905 gnd.n5254 gnd.n5253 9.3005
R9906 gnd.n5252 gnd.n1371 9.3005
R9907 gnd.n5251 gnd.n5250 9.3005
R9908 gnd.n5249 gnd.n1375 9.3005
R9909 gnd.n5248 gnd.n5247 9.3005
R9910 gnd.n5246 gnd.n1376 9.3005
R9911 gnd.n5245 gnd.n5244 9.3005
R9912 gnd.n5243 gnd.n1380 9.3005
R9913 gnd.n5242 gnd.n5241 9.3005
R9914 gnd.n5240 gnd.n1381 9.3005
R9915 gnd.n5239 gnd.n5238 9.3005
R9916 gnd.n5237 gnd.n1385 9.3005
R9917 gnd.n5236 gnd.n5235 9.3005
R9918 gnd.n5234 gnd.n1386 9.3005
R9919 gnd.n5233 gnd.n5232 9.3005
R9920 gnd.n5231 gnd.n1390 9.3005
R9921 gnd.n5230 gnd.n5229 9.3005
R9922 gnd.n5228 gnd.n1391 9.3005
R9923 gnd.n5227 gnd.n5226 9.3005
R9924 gnd.n5225 gnd.n1395 9.3005
R9925 gnd.n5224 gnd.n5223 9.3005
R9926 gnd.n5222 gnd.n1396 9.3005
R9927 gnd.n5221 gnd.n5220 9.3005
R9928 gnd.n5219 gnd.n1400 9.3005
R9929 gnd.n5218 gnd.n5217 9.3005
R9930 gnd.n5216 gnd.n1401 9.3005
R9931 gnd.n5215 gnd.n5214 9.3005
R9932 gnd.n5213 gnd.n1405 9.3005
R9933 gnd.n5212 gnd.n5211 9.3005
R9934 gnd.n5210 gnd.n1406 9.3005
R9935 gnd.n5209 gnd.n5208 9.3005
R9936 gnd.n5207 gnd.n1410 9.3005
R9937 gnd.n5206 gnd.n5205 9.3005
R9938 gnd.n5204 gnd.n1411 9.3005
R9939 gnd.n5203 gnd.n5202 9.3005
R9940 gnd.n5201 gnd.n1415 9.3005
R9941 gnd.n5200 gnd.n5199 9.3005
R9942 gnd.n4230 gnd.n4229 9.3005
R9943 gnd.n4216 gnd.n1863 9.3005
R9944 gnd.n4215 gnd.n4214 9.3005
R9945 gnd.n4211 gnd.n1864 9.3005
R9946 gnd.n4209 gnd.n4208 9.3005
R9947 gnd.n4207 gnd.n1867 9.3005
R9948 gnd.n4206 gnd.n4205 9.3005
R9949 gnd.n4202 gnd.n1870 9.3005
R9950 gnd.n4201 gnd.n4200 9.3005
R9951 gnd.n4199 gnd.n1871 9.3005
R9952 gnd.n4232 gnd.n4231 9.3005
R9953 gnd.n3669 gnd.n3668 9.3005
R9954 gnd.n2022 gnd.n2021 9.3005
R9955 gnd.n4003 gnd.n4002 9.3005
R9956 gnd.n4004 gnd.n2020 9.3005
R9957 gnd.n4006 gnd.n4005 9.3005
R9958 gnd.n2015 gnd.n2013 9.3005
R9959 gnd.n4028 gnd.n4027 9.3005
R9960 gnd.n4026 gnd.n2014 9.3005
R9961 gnd.n4025 gnd.n4024 9.3005
R9962 gnd.n2005 gnd.n2004 9.3005
R9963 gnd.n4060 gnd.n4059 9.3005
R9964 gnd.n4061 gnd.n2003 9.3005
R9965 gnd.n4063 gnd.n4062 9.3005
R9966 gnd.n1995 gnd.n1993 9.3005
R9967 gnd.n4160 gnd.n4159 9.3005
R9968 gnd.n4158 gnd.n1994 9.3005
R9969 gnd.n4157 gnd.n4156 9.3005
R9970 gnd.n4155 gnd.n1996 9.3005
R9971 gnd.n4154 gnd.n4153 9.3005
R9972 gnd.n4152 gnd.n4151 9.3005
R9973 gnd.n1980 gnd.n1874 9.3005
R9974 gnd.n4197 gnd.n4196 9.3005
R9975 gnd.n4193 gnd.n1875 9.3005
R9976 gnd.n4192 gnd.n4191 9.3005
R9977 gnd.n1972 gnd.n1876 9.3005
R9978 gnd.n1971 gnd.n1970 9.3005
R9979 gnd.n1967 gnd.n1966 9.3005
R9980 gnd.n1883 gnd.n1882 9.3005
R9981 gnd.n1959 gnd.n1958 9.3005
R9982 gnd.n1955 gnd.n1954 9.3005
R9983 gnd.n1891 gnd.n1888 9.3005
R9984 gnd.n1947 gnd.n1946 9.3005
R9985 gnd.n1943 gnd.n1942 9.3005
R9986 gnd.n1895 gnd.n1894 9.3005
R9987 gnd.n1935 gnd.n1934 9.3005
R9988 gnd.n1931 gnd.n1930 9.3005
R9989 gnd.n1903 gnd.n1900 9.3005
R9990 gnd.n1923 gnd.n1922 9.3005
R9991 gnd.n1919 gnd.n1918 9.3005
R9992 gnd.n1907 gnd.n1906 9.3005
R9993 gnd.n1913 gnd.n1912 9.3005
R9994 gnd.n1917 gnd.n1916 9.3005
R9995 gnd.n1905 gnd.n1904 9.3005
R9996 gnd.n1925 gnd.n1924 9.3005
R9997 gnd.n1929 gnd.n1928 9.3005
R9998 gnd.n1899 gnd.n1896 9.3005
R9999 gnd.n1937 gnd.n1936 9.3005
R10000 gnd.n1941 gnd.n1940 9.3005
R10001 gnd.n1893 gnd.n1892 9.3005
R10002 gnd.n1949 gnd.n1948 9.3005
R10003 gnd.n1953 gnd.n1952 9.3005
R10004 gnd.n1887 gnd.n1884 9.3005
R10005 gnd.n1961 gnd.n1960 9.3005
R10006 gnd.n1965 gnd.n1964 9.3005
R10007 gnd.n1881 gnd.n1880 9.3005
R10008 gnd.n1974 gnd.n1973 9.3005
R10009 gnd.n1979 gnd.n1879 9.3005
R10010 gnd.n4190 gnd.n4189 9.3005
R10011 gnd.n4255 gnd.n1835 9.3005
R10012 gnd.n4257 gnd.n4256 9.3005
R10013 gnd.n1833 gnd.n1832 9.3005
R10014 gnd.n4262 gnd.n4261 9.3005
R10015 gnd.n4263 gnd.n1831 9.3005
R10016 gnd.n4265 gnd.n4264 9.3005
R10017 gnd.n1824 gnd.n1823 9.3005
R10018 gnd.n4287 gnd.n4286 9.3005
R10019 gnd.n4288 gnd.n1822 9.3005
R10020 gnd.n4290 gnd.n4289 9.3005
R10021 gnd.n4321 gnd.n1821 9.3005
R10022 gnd.n4323 gnd.n4322 9.3005
R10023 gnd.n4324 gnd.n1819 9.3005
R10024 gnd.n4428 gnd.n4427 9.3005
R10025 gnd.n4426 gnd.n1820 9.3005
R10026 gnd.n4425 gnd.n4424 9.3005
R10027 gnd.n4423 gnd.n4325 9.3005
R10028 gnd.n4422 gnd.n4421 9.3005
R10029 gnd.n4420 gnd.n4327 9.3005
R10030 gnd.n4419 gnd.n4418 9.3005
R10031 gnd.n4417 gnd.n4328 9.3005
R10032 gnd.n4416 gnd.n4415 9.3005
R10033 gnd.n4414 gnd.n4333 9.3005
R10034 gnd.n4413 gnd.n4412 9.3005
R10035 gnd.n4411 gnd.n4334 9.3005
R10036 gnd.n4410 gnd.n4409 9.3005
R10037 gnd.n4408 gnd.n4336 9.3005
R10038 gnd.n4407 gnd.n4406 9.3005
R10039 gnd.n4405 gnd.n4337 9.3005
R10040 gnd.n4404 gnd.n4403 9.3005
R10041 gnd.n4402 gnd.n4340 9.3005
R10042 gnd.n4401 gnd.n4400 9.3005
R10043 gnd.n4399 gnd.n4341 9.3005
R10044 gnd.n4398 gnd.n4397 9.3005
R10045 gnd.n4396 gnd.n4344 9.3005
R10046 gnd.n4395 gnd.n4394 9.3005
R10047 gnd.n4393 gnd.n4345 9.3005
R10048 gnd.n4392 gnd.n4391 9.3005
R10049 gnd.n4390 gnd.n4348 9.3005
R10050 gnd.n4389 gnd.n4388 9.3005
R10051 gnd.n4387 gnd.n4349 9.3005
R10052 gnd.n4386 gnd.n4385 9.3005
R10053 gnd.n4384 gnd.n4353 9.3005
R10054 gnd.n4383 gnd.n4382 9.3005
R10055 gnd.n4381 gnd.n4354 9.3005
R10056 gnd.n4380 gnd.n4379 9.3005
R10057 gnd.n4378 gnd.n4357 9.3005
R10058 gnd.n4377 gnd.n4376 9.3005
R10059 gnd.n4375 gnd.n4358 9.3005
R10060 gnd.n4374 gnd.n4373 9.3005
R10061 gnd.n4372 gnd.n4360 9.3005
R10062 gnd.n4371 gnd.n4370 9.3005
R10063 gnd.n4369 gnd.n4361 9.3005
R10064 gnd.n4368 gnd.n4367 9.3005
R10065 gnd.n4366 gnd.n4365 9.3005
R10066 gnd.n1609 gnd.n1608 9.3005
R10067 gnd.n4763 gnd.n4762 9.3005
R10068 gnd.n4764 gnd.n1606 9.3005
R10069 gnd.n4795 gnd.n4794 9.3005
R10070 gnd.n4793 gnd.n1607 9.3005
R10071 gnd.n4792 gnd.n4791 9.3005
R10072 gnd.n4790 gnd.n4765 9.3005
R10073 gnd.n4789 gnd.n4788 9.3005
R10074 gnd.n4787 gnd.n4769 9.3005
R10075 gnd.n4786 gnd.n4785 9.3005
R10076 gnd.n4784 gnd.n4770 9.3005
R10077 gnd.n4783 gnd.n4782 9.3005
R10078 gnd.n4781 gnd.n4773 9.3005
R10079 gnd.n4780 gnd.n4779 9.3005
R10080 gnd.n4778 gnd.n4774 9.3005
R10081 gnd.n4777 gnd.n4776 9.3005
R10082 gnd.n1536 gnd.n1534 9.3005
R10083 gnd.n4910 gnd.n4909 9.3005
R10084 gnd.n4908 gnd.n1535 9.3005
R10085 gnd.n4907 gnd.n4906 9.3005
R10086 gnd.n4905 gnd.n1537 9.3005
R10087 gnd.n4904 gnd.n4903 9.3005
R10088 gnd.n4902 gnd.n4901 9.3005
R10089 gnd.n1425 gnd.n1424 9.3005
R10090 gnd.n5192 gnd.n5191 9.3005
R10091 gnd.n5193 gnd.n1423 9.3005
R10092 gnd.n5195 gnd.n5194 9.3005
R10093 gnd.n4254 gnd.n4253 9.3005
R10094 gnd.n319 gnd.n318 9.3005
R10095 gnd.n6456 gnd.n6455 9.3005
R10096 gnd.n6457 gnd.n317 9.3005
R10097 gnd.n6459 gnd.n6458 9.3005
R10098 gnd.n301 gnd.n300 9.3005
R10099 gnd.n6472 gnd.n6471 9.3005
R10100 gnd.n6473 gnd.n299 9.3005
R10101 gnd.n6475 gnd.n6474 9.3005
R10102 gnd.n283 gnd.n282 9.3005
R10103 gnd.n6488 gnd.n6487 9.3005
R10104 gnd.n6489 gnd.n281 9.3005
R10105 gnd.n6491 gnd.n6490 9.3005
R10106 gnd.n266 gnd.n265 9.3005
R10107 gnd.n6505 gnd.n6504 9.3005
R10108 gnd.n6506 gnd.n263 9.3005
R10109 gnd.n6512 gnd.n6511 9.3005
R10110 gnd.n6510 gnd.n264 9.3005
R10111 gnd.n6509 gnd.n6508 9.3005
R10112 gnd.n241 gnd.n240 9.3005
R10113 gnd.n6535 gnd.n6534 9.3005
R10114 gnd.n6536 gnd.n238 9.3005
R10115 gnd.n6538 gnd.n6537 9.3005
R10116 gnd.n228 gnd.n227 9.3005
R10117 gnd.n6549 gnd.n6548 9.3005
R10118 gnd.n6550 gnd.n226 9.3005
R10119 gnd.n6552 gnd.n6551 9.3005
R10120 gnd.n207 gnd.n206 9.3005
R10121 gnd.n6565 gnd.n6564 9.3005
R10122 gnd.n6566 gnd.n205 9.3005
R10123 gnd.n6568 gnd.n6567 9.3005
R10124 gnd.n192 gnd.n191 9.3005
R10125 gnd.n6581 gnd.n6580 9.3005
R10126 gnd.n6582 gnd.n190 9.3005
R10127 gnd.n6584 gnd.n6583 9.3005
R10128 gnd.n176 gnd.n175 9.3005
R10129 gnd.n6597 gnd.n6596 9.3005
R10130 gnd.n6598 gnd.n173 9.3005
R10131 gnd.n6674 gnd.n6673 9.3005
R10132 gnd.n6672 gnd.n174 9.3005
R10133 gnd.n6671 gnd.n6670 9.3005
R10134 gnd.n6669 gnd.n6599 9.3005
R10135 gnd.n6668 gnd.n6667 9.3005
R10136 gnd.n6443 gnd.n6442 9.3005
R10137 gnd.n6664 gnd.n6601 9.3005
R10138 gnd.n6663 gnd.n6662 9.3005
R10139 gnd.n6661 gnd.n6606 9.3005
R10140 gnd.n6660 gnd.n6659 9.3005
R10141 gnd.n6658 gnd.n6607 9.3005
R10142 gnd.n6657 gnd.n6656 9.3005
R10143 gnd.n6655 gnd.n6614 9.3005
R10144 gnd.n6654 gnd.n6653 9.3005
R10145 gnd.n6652 gnd.n6615 9.3005
R10146 gnd.n6651 gnd.n6650 9.3005
R10147 gnd.n6649 gnd.n6622 9.3005
R10148 gnd.n6648 gnd.n6647 9.3005
R10149 gnd.n6646 gnd.n6623 9.3005
R10150 gnd.n6645 gnd.n6644 9.3005
R10151 gnd.n6643 gnd.n6630 9.3005
R10152 gnd.n6642 gnd.n6641 9.3005
R10153 gnd.n6640 gnd.n6631 9.3005
R10154 gnd.n6639 gnd.n78 9.3005
R10155 gnd.n6666 gnd.n6665 9.3005
R10156 gnd.n5152 gnd.n5105 9.3005
R10157 gnd.n470 gnd.n468 9.3005
R10158 gnd.n6308 gnd.n6307 9.3005
R10159 gnd.n6306 gnd.n469 9.3005
R10160 gnd.n6305 gnd.n6304 9.3005
R10161 gnd.n6303 gnd.n471 9.3005
R10162 gnd.n6302 gnd.n6301 9.3005
R10163 gnd.n6300 gnd.n474 9.3005
R10164 gnd.n6299 gnd.n6298 9.3005
R10165 gnd.n6297 gnd.n475 9.3005
R10166 gnd.n6296 gnd.n6295 9.3005
R10167 gnd.n6294 gnd.n478 9.3005
R10168 gnd.n6293 gnd.n6292 9.3005
R10169 gnd.n6291 gnd.n479 9.3005
R10170 gnd.n6290 gnd.n6289 9.3005
R10171 gnd.n253 gnd.n252 9.3005
R10172 gnd.n6522 gnd.n6521 9.3005
R10173 gnd.n6523 gnd.n250 9.3005
R10174 gnd.n6525 gnd.n6524 9.3005
R10175 gnd.n251 gnd.n51 9.3005
R10176 gnd.n6798 gnd.n52 9.3005
R10177 gnd.n6797 gnd.n6796 9.3005
R10178 gnd.n6795 gnd.n53 9.3005
R10179 gnd.n6794 gnd.n6793 9.3005
R10180 gnd.n6792 gnd.n57 9.3005
R10181 gnd.n6791 gnd.n6790 9.3005
R10182 gnd.n6789 gnd.n58 9.3005
R10183 gnd.n6788 gnd.n6787 9.3005
R10184 gnd.n6786 gnd.n62 9.3005
R10185 gnd.n6785 gnd.n6784 9.3005
R10186 gnd.n6783 gnd.n63 9.3005
R10187 gnd.n6782 gnd.n6781 9.3005
R10188 gnd.n6780 gnd.n67 9.3005
R10189 gnd.n6779 gnd.n6778 9.3005
R10190 gnd.n6777 gnd.n68 9.3005
R10191 gnd.n6776 gnd.n6775 9.3005
R10192 gnd.n6774 gnd.n72 9.3005
R10193 gnd.n6773 gnd.n6772 9.3005
R10194 gnd.n6771 gnd.n73 9.3005
R10195 gnd.n6770 gnd.n6769 9.3005
R10196 gnd.n6768 gnd.n77 9.3005
R10197 gnd.n6767 gnd.n6766 9.3005
R10198 gnd.n5154 gnd.n5153 9.3005
R10199 gnd.t198 gnd.n2310 9.24152
R10200 gnd.n2212 gnd.t109 9.24152
R10201 gnd.n3469 gnd.t113 9.24152
R10202 gnd.t22 gnd.t198 8.92286
R10203 gnd.n5334 gnd.n1207 8.92286
R10204 gnd.n4491 gnd.n1786 8.92286
R10205 gnd.n4526 gnd.n4525 8.92286
R10206 gnd.n4615 gnd.n1705 8.92286
R10207 gnd.n4649 gnd.n4648 8.92286
R10208 gnd.n4750 gnd.n4749 8.92286
R10209 gnd.n4732 gnd.n1589 8.92286
R10210 gnd.n1540 gnd.n1531 8.92286
R10211 gnd.n5064 gnd.n1433 8.92286
R10212 gnd.n3439 gnd.n3414 8.92171
R10213 gnd.n3407 gnd.n3382 8.92171
R10214 gnd.n3375 gnd.n3350 8.92171
R10215 gnd.n3344 gnd.n3319 8.92171
R10216 gnd.n3312 gnd.n3287 8.92171
R10217 gnd.n3280 gnd.n3255 8.92171
R10218 gnd.n3248 gnd.n3223 8.92171
R10219 gnd.n3217 gnd.n3192 8.92171
R10220 gnd.n1458 gnd.n1440 8.72777
R10221 gnd.n2942 gnd.t184 8.60421
R10222 gnd.n5404 gnd.n1149 8.60421
R10223 gnd.t215 gnd.n4614 8.60421
R10224 gnd.n4626 gnd.t251 8.60421
R10225 gnd.n2374 gnd.n2362 8.43467
R10226 gnd.n38 gnd.n26 8.43467
R10227 gnd.n3670 gnd.n0 8.41456
R10228 gnd.n6799 gnd.n6798 8.41456
R10229 gnd.t150 gnd.n1181 8.28555
R10230 gnd.n3440 gnd.n3412 8.14595
R10231 gnd.n3408 gnd.n3380 8.14595
R10232 gnd.n3376 gnd.n3348 8.14595
R10233 gnd.n3345 gnd.n3317 8.14595
R10234 gnd.n3313 gnd.n3285 8.14595
R10235 gnd.n3281 gnd.n3253 8.14595
R10236 gnd.n3249 gnd.n3221 8.14595
R10237 gnd.n3218 gnd.n3190 8.14595
R10238 gnd.n3445 gnd.n3444 7.97301
R10239 gnd.t223 gnd.n2457 7.9669
R10240 gnd.n4451 gnd.t205 7.9669
R10241 gnd.n4827 gnd.t255 7.9669
R10242 gnd.n6640 gnd.n6639 7.75808
R10243 gnd.n6392 gnd.n377 7.75808
R10244 gnd.n4189 gnd.n1979 7.75808
R10245 gnd.n3705 gnd.n3601 7.75808
R10246 gnd.n3183 gnd.n2209 7.64824
R10247 gnd.n4284 gnd.t169 7.64824
R10248 gnd.n5307 gnd.n1323 7.64824
R10249 gnd.t266 gnd.n1790 7.64824
R10250 gnd.n4572 gnd.t3 7.64824
R10251 gnd.n4582 gnd.t3 7.64824
R10252 gnd.n4675 gnd.t4 7.64824
R10253 gnd.n4683 gnd.t4 7.64824
R10254 gnd.n4822 gnd.t0 7.64824
R10255 gnd.n4880 gnd.n1544 7.64824
R10256 gnd.n4913 gnd.t156 7.64824
R10257 gnd.n2851 gnd.t282 7.32958
R10258 gnd.t203 gnd.t106 7.32958
R10259 gnd.n1203 gnd.n1202 7.30353
R10260 gnd.n1457 gnd.n1456 7.30353
R10261 gnd.n2811 gnd.n2530 7.01093
R10262 gnd.n2533 gnd.n2531 7.01093
R10263 gnd.n2821 gnd.n2820 7.01093
R10264 gnd.n2832 gnd.n2514 7.01093
R10265 gnd.n2831 gnd.n2517 7.01093
R10266 gnd.n2842 gnd.n2505 7.01093
R10267 gnd.n2508 gnd.n2506 7.01093
R10268 gnd.n2852 gnd.n2851 7.01093
R10269 gnd.n2862 gnd.n2486 7.01093
R10270 gnd.n2861 gnd.n2489 7.01093
R10271 gnd.n2870 gnd.n2480 7.01093
R10272 gnd.n2882 gnd.n2470 7.01093
R10273 gnd.n2892 gnd.n2455 7.01093
R10274 gnd.n2908 gnd.n2907 7.01093
R10275 gnd.n2457 gnd.n2394 7.01093
R10276 gnd.n2962 gnd.n2395 7.01093
R10277 gnd.n2956 gnd.n2955 7.01093
R10278 gnd.n2444 gnd.n2406 7.01093
R10279 gnd.n2948 gnd.n2417 7.01093
R10280 gnd.n2435 gnd.n2430 7.01093
R10281 gnd.n2942 gnd.n2941 7.01093
R10282 gnd.n2988 gnd.n2345 7.01093
R10283 gnd.n2987 gnd.n2986 7.01093
R10284 gnd.n2999 gnd.n2998 7.01093
R10285 gnd.n2338 gnd.n2330 7.01093
R10286 gnd.n3028 gnd.n2318 7.01093
R10287 gnd.n3027 gnd.n2321 7.01093
R10288 gnd.n3038 gnd.n2310 7.01093
R10289 gnd.n2311 gnd.n2299 7.01093
R10290 gnd.n3049 gnd.n2300 7.01093
R10291 gnd.n3073 gnd.n2291 7.01093
R10292 gnd.n3072 gnd.n2282 7.01093
R10293 gnd.n3095 gnd.n3094 7.01093
R10294 gnd.n3113 gnd.n2263 7.01093
R10295 gnd.n3112 gnd.n2266 7.01093
R10296 gnd.n3123 gnd.n2255 7.01093
R10297 gnd.n2256 gnd.n2243 7.01093
R10298 gnd.n3134 gnd.n2244 7.01093
R10299 gnd.n3161 gnd.n2228 7.01093
R10300 gnd.n3173 gnd.n3172 7.01093
R10301 gnd.n3155 gnd.n2221 7.01093
R10302 gnd.n3185 gnd.n3184 7.01093
R10303 gnd.n3457 gnd.n2209 7.01093
R10304 gnd.n3456 gnd.n2212 7.01093
R10305 gnd.n3469 gnd.n2201 7.01093
R10306 gnd.n2202 gnd.n2194 7.01093
R10307 gnd.n3479 gnd.n2120 7.01093
R10308 gnd.n4601 gnd.t28 7.01093
R10309 gnd.n4665 gnd.t242 7.01093
R10310 gnd.n5064 gnd.t127 7.01093
R10311 gnd.n2489 gnd.t222 6.69227
R10312 gnd.n2321 gnd.t22 6.69227
R10313 gnd.n3162 gnd.t9 6.69227
R10314 gnd.n4163 gnd.t209 6.69227
R10315 gnd.n1792 gnd.t26 6.69227
R10316 gnd.t46 gnd.n4815 6.69227
R10317 gnd.t53 gnd.n306 6.69227
R10318 gnd.n4994 gnd.n4993 6.5566
R10319 gnd.n1233 gnd.n1232 6.5566
R10320 gnd.n5345 gnd.n5341 6.5566
R10321 gnd.n5009 gnd.n5008 6.5566
R10322 gnd.n4430 gnd.n1817 6.37362
R10323 gnd.n4459 gnd.n4457 6.37362
R10324 gnd.n4554 gnd.n4553 6.37362
R10325 gnd.n4704 gnd.n4703 6.37362
R10326 gnd.n4842 gnd.n1571 6.37362
R10327 gnd.n4858 gnd.n1558 6.37362
R10328 gnd.n1519 gnd.t71 6.37362
R10329 gnd.n4211 gnd.n4210 6.20656
R10330 gnd.n6729 gnd.n6726 6.20656
R10331 gnd.n3842 gnd.n3841 6.20656
R10332 gnd.n5173 gnd.n5171 6.20656
R10333 gnd.t190 gnd.n2918 6.05496
R10334 gnd.n2919 gnd.t187 6.05496
R10335 gnd.t275 gnd.n2345 6.05496
R10336 gnd.t188 gnd.n3083 6.05496
R10337 gnd.n4031 gnd.t207 6.05496
R10338 gnd.t34 gnd.n271 6.05496
R10339 gnd.n3442 gnd.n3412 5.81868
R10340 gnd.n3410 gnd.n3380 5.81868
R10341 gnd.n3378 gnd.n3348 5.81868
R10342 gnd.n3347 gnd.n3317 5.81868
R10343 gnd.n3315 gnd.n3285 5.81868
R10344 gnd.n3283 gnd.n3253 5.81868
R10345 gnd.n3251 gnd.n3221 5.81868
R10346 gnd.n3220 gnd.n3190 5.81868
R10347 gnd.n5314 gnd.t85 5.73631
R10348 gnd.n4491 gnd.t69 5.73631
R10349 gnd.n4561 gnd.t21 5.73631
R10350 gnd.n4695 gnd.t37 5.73631
R10351 gnd.n4732 gnd.t29 5.73631
R10352 gnd.t127 gnd.n5063 5.73631
R10353 gnd.n1485 gnd.n435 5.62001
R10354 gnd.n5407 gnd.n1145 5.62001
R10355 gnd.n5407 gnd.n1146 5.62001
R10356 gnd.n5003 gnd.n435 5.62001
R10357 gnd.n2670 gnd.n2665 5.4308
R10358 gnd.n3487 gnd.n2187 5.4308
R10359 gnd.n2986 gnd.t189 5.41765
R10360 gnd.t185 gnd.n3009 5.41765
R10361 gnd.t63 gnd.n2275 5.41765
R10362 gnd.n4517 gnd.t58 5.41765
R10363 gnd.n4760 gnd.t1 5.41765
R10364 gnd.n4008 gnd.n1001 5.09899
R10365 gnd.n5487 gnd.n1010 5.09899
R10366 gnd.n4031 gnd.n4030 5.09899
R10367 gnd.n5481 gnd.n1021 5.09899
R10368 gnd.n4022 gnd.n1024 5.09899
R10369 gnd.n5475 gnd.n1032 5.09899
R10370 gnd.n4057 gnd.n1035 5.09899
R10371 gnd.n4065 gnd.n1045 5.09899
R10372 gnd.n5463 gnd.n1053 5.09899
R10373 gnd.n4163 gnd.n4162 5.09899
R10374 gnd.n5457 gnd.n1063 5.09899
R10375 gnd.n4073 gnd.n1066 5.09899
R10376 gnd.n5451 gnd.n1074 5.09899
R10377 gnd.n4149 gnd.n1077 5.09899
R10378 gnd.n5445 gnd.n1085 5.09899
R10379 gnd.n4186 gnd.n1088 5.09899
R10380 gnd.n4439 gnd.n4438 5.09899
R10381 gnd.n4451 gnd.n4450 5.09899
R10382 gnd.n4543 gnd.t36 5.09899
R10383 gnd.n1736 gnd.n1731 5.09899
R10384 gnd.n4575 gnd.n4574 5.09899
R10385 gnd.n1654 gnd.n1648 5.09899
R10386 gnd.n4697 gnd.n4696 5.09899
R10387 gnd.n4712 gnd.t231 5.09899
R10388 gnd.n4827 gnd.n1574 5.09899
R10389 gnd.n4851 gnd.n4850 5.09899
R10390 gnd.n6445 gnd.n331 5.09899
R10391 gnd.n5150 gnd.n5149 5.09899
R10392 gnd.n6453 gnd.n323 5.09899
R10393 gnd.n6310 gnd.n312 5.09899
R10394 gnd.n6461 gnd.n315 5.09899
R10395 gnd.n487 gnd.n303 5.09899
R10396 gnd.n6469 gnd.n306 5.09899
R10397 gnd.n493 gnd.n294 5.09899
R10398 gnd.n6477 gnd.n297 5.09899
R10399 gnd.n6485 gnd.n288 5.09899
R10400 gnd.n6217 gnd.n6216 5.09899
R10401 gnd.n6493 gnd.n279 5.09899
R10402 gnd.n6221 gnd.n268 5.09899
R10403 gnd.n6502 gnd.n271 5.09899
R10404 gnd.n6287 gnd.n260 5.09899
R10405 gnd.n6514 gnd.n255 5.09899
R10406 gnd.n3440 gnd.n3439 5.04292
R10407 gnd.n3408 gnd.n3407 5.04292
R10408 gnd.n3376 gnd.n3375 5.04292
R10409 gnd.n3345 gnd.n3344 5.04292
R10410 gnd.n3313 gnd.n3312 5.04292
R10411 gnd.n3281 gnd.n3280 5.04292
R10412 gnd.n3249 gnd.n3248 5.04292
R10413 gnd.n3218 gnd.n3217 5.04292
R10414 gnd.n2386 gnd.n2385 4.82753
R10415 gnd.n50 gnd.n49 4.82753
R10416 gnd.n2949 gnd.t68 4.78034
R10417 gnd.n2300 gnd.t67 4.78034
R10418 gnd.n1774 gnd.t58 4.78034
R10419 gnd.n4742 gnd.t1 4.78034
R10420 gnd.n1461 gnd.t92 4.78034
R10421 gnd.n2391 gnd.n2388 4.74817
R10422 gnd.n2441 gnd.n2351 4.74817
R10423 gnd.n2428 gnd.n2350 4.74817
R10424 gnd.n2349 gnd.n2348 4.74817
R10425 gnd.n2437 gnd.n2388 4.74817
R10426 gnd.n2438 gnd.n2351 4.74817
R10427 gnd.n2440 gnd.n2350 4.74817
R10428 gnd.n2427 gnd.n2349 4.74817
R10429 gnd.n6517 gnd.n218 4.74817
R10430 gnd.n6529 gnd.n217 4.74817
R10431 gnd.n233 gnd.n216 4.74817
R10432 gnd.n6543 gnd.n215 4.74817
R10433 gnd.n219 gnd.n214 4.74817
R10434 gnd.n259 gnd.n218 4.74817
R10435 gnd.n6516 gnd.n217 4.74817
R10436 gnd.n6530 gnd.n216 4.74817
R10437 gnd.n234 gnd.n215 4.74817
R10438 gnd.n6544 gnd.n214 4.74817
R10439 gnd.n3958 gnd.n2045 4.74817
R10440 gnd.n3962 gnd.n3960 4.74817
R10441 gnd.n3993 gnd.n2027 4.74817
R10442 gnd.n3997 gnd.n3995 4.74817
R10443 gnd.n5491 gnd.n1005 4.74817
R10444 gnd.n3941 gnd.n2045 4.74817
R10445 gnd.n3960 gnd.n3959 4.74817
R10446 gnd.n3961 gnd.n2027 4.74817
R10447 gnd.n3995 gnd.n3994 4.74817
R10448 gnd.n3996 gnd.n1005 4.74817
R10449 gnd.n2374 gnd.n2373 4.7074
R10450 gnd.n38 gnd.n37 4.7074
R10451 gnd.n2386 gnd.n2374 4.65959
R10452 gnd.n50 gnd.n38 4.65959
R10453 gnd.n6359 gnd.n437 4.6132
R10454 gnd.n5408 gnd.n1144 4.6132
R10455 gnd.n5437 gnd.n1095 4.46168
R10456 gnd.t11 gnd.n1323 4.46168
R10457 gnd.n4880 gnd.t267 4.46168
R10458 gnd.n6390 gnd.n417 4.46168
R10459 gnd.n1453 gnd.n1440 4.46111
R10460 gnd.n3425 gnd.n3421 4.38594
R10461 gnd.n3393 gnd.n3389 4.38594
R10462 gnd.n3361 gnd.n3357 4.38594
R10463 gnd.n3330 gnd.n3326 4.38594
R10464 gnd.n3298 gnd.n3294 4.38594
R10465 gnd.n3266 gnd.n3262 4.38594
R10466 gnd.n3234 gnd.n3230 4.38594
R10467 gnd.n3203 gnd.n3199 4.38594
R10468 gnd.n3436 gnd.n3414 4.26717
R10469 gnd.n3404 gnd.n3382 4.26717
R10470 gnd.n3372 gnd.n3350 4.26717
R10471 gnd.n3341 gnd.n3319 4.26717
R10472 gnd.n3309 gnd.n3287 4.26717
R10473 gnd.n3277 gnd.n3255 4.26717
R10474 gnd.n3245 gnd.n3223 4.26717
R10475 gnd.n3214 gnd.n3192 4.26717
R10476 gnd.n2893 gnd.t10 4.14303
R10477 gnd.n3123 gnd.t183 4.14303
R10478 gnd.n4056 gnd.t60 4.14303
R10479 gnd.t236 gnd.n4581 4.14303
R10480 gnd.n4676 gnd.t229 4.14303
R10481 gnd.t32 gnd.n285 4.14303
R10482 gnd.n3444 gnd.n3443 4.08274
R10483 gnd.n4993 gnd.n4992 4.05904
R10484 gnd.n1234 gnd.n1233 4.05904
R10485 gnd.n5348 gnd.n5341 4.05904
R10486 gnd.n5010 gnd.n5009 4.05904
R10487 gnd.n15 gnd.n7 3.99943
R10488 gnd.n5320 gnd.t169 3.82437
R10489 gnd.n4311 gnd.n4298 3.82437
R10490 gnd.n1807 gnd.n1796 3.82437
R10491 gnd.n4555 gnd.n1740 3.82437
R10492 gnd.n1727 gnd.n1716 3.82437
R10493 gnd.n4677 gnd.n1658 3.82437
R10494 gnd.n4362 gnd.n1644 3.82437
R10495 gnd.n4834 gnd.n1578 3.82437
R10496 gnd.n4868 gnd.n1553 3.82437
R10497 gnd.n5189 gnd.t92 3.82437
R10498 gnd.n3444 gnd.n3316 3.70378
R10499 gnd.n2966 gnd.n2387 3.65935
R10500 gnd.n15 gnd.n14 3.60163
R10501 gnd.n3435 gnd.n3416 3.49141
R10502 gnd.n3403 gnd.n3384 3.49141
R10503 gnd.n3371 gnd.n3352 3.49141
R10504 gnd.n3340 gnd.n3321 3.49141
R10505 gnd.n3308 gnd.n3289 3.49141
R10506 gnd.n3276 gnd.n3257 3.49141
R10507 gnd.n3244 gnd.n3225 3.49141
R10508 gnd.n3213 gnd.n3194 3.49141
R10509 gnd.t85 gnd.n5313 3.18706
R10510 gnd.n4898 gnd.t143 3.18706
R10511 gnd.n179 gnd.n169 3.18706
R10512 gnd.n2472 gnd.t10 2.8684
R10513 gnd.n2375 gnd.t272 2.82907
R10514 gnd.n2375 gnd.t220 2.82907
R10515 gnd.n2377 gnd.t238 2.82907
R10516 gnd.n2377 gnd.t234 2.82907
R10517 gnd.n2379 gnd.t243 2.82907
R10518 gnd.n2379 gnd.t245 2.82907
R10519 gnd.n2381 gnd.t259 2.82907
R10520 gnd.n2381 gnd.t219 2.82907
R10521 gnd.n2383 gnd.t277 2.82907
R10522 gnd.n2383 gnd.t227 2.82907
R10523 gnd.n2352 gnd.t45 2.82907
R10524 gnd.n2352 gnd.t61 2.82907
R10525 gnd.n2354 gnd.t18 2.82907
R10526 gnd.n2354 gnd.t249 2.82907
R10527 gnd.n2356 gnd.t274 2.82907
R10528 gnd.n2356 gnd.t39 2.82907
R10529 gnd.n2358 gnd.t226 2.82907
R10530 gnd.n2358 gnd.t269 2.82907
R10531 gnd.n2360 gnd.t286 2.82907
R10532 gnd.n2360 gnd.t16 2.82907
R10533 gnd.n2363 gnd.t284 2.82907
R10534 gnd.n2363 gnd.t66 2.82907
R10535 gnd.n2365 gnd.t261 2.82907
R10536 gnd.n2365 gnd.t208 2.82907
R10537 gnd.n2367 gnd.t196 2.82907
R10538 gnd.n2367 gnd.t182 2.82907
R10539 gnd.n2369 gnd.t270 2.82907
R10540 gnd.n2369 gnd.t224 2.82907
R10541 gnd.n2371 gnd.t233 2.82907
R10542 gnd.n2371 gnd.t62 2.82907
R10543 gnd.n47 gnd.t13 2.82907
R10544 gnd.n47 gnd.t41 2.82907
R10545 gnd.n45 gnd.t8 2.82907
R10546 gnd.n45 gnd.t211 2.82907
R10547 gnd.n43 gnd.t214 2.82907
R10548 gnd.n43 gnd.t194 2.82907
R10549 gnd.n41 gnd.t35 2.82907
R10550 gnd.n41 gnd.t283 2.82907
R10551 gnd.n39 gnd.t43 2.82907
R10552 gnd.n39 gnd.t244 2.82907
R10553 gnd.n24 gnd.t265 2.82907
R10554 gnd.n24 gnd.t50 2.82907
R10555 gnd.n22 gnd.t290 2.82907
R10556 gnd.n22 gnd.t179 2.82907
R10557 gnd.n20 gnd.t31 2.82907
R10558 gnd.n20 gnd.t273 2.82907
R10559 gnd.n18 gnd.t197 2.82907
R10560 gnd.n18 gnd.t268 2.82907
R10561 gnd.n16 gnd.t33 2.82907
R10562 gnd.n16 gnd.t263 2.82907
R10563 gnd.n35 gnd.t65 2.82907
R10564 gnd.n35 gnd.t260 2.82907
R10565 gnd.n33 gnd.t42 2.82907
R10566 gnd.n33 gnd.t192 2.82907
R10567 gnd.n31 gnd.t55 2.82907
R10568 gnd.n31 gnd.t291 2.82907
R10569 gnd.n29 gnd.t289 2.82907
R10570 gnd.n29 gnd.t247 2.82907
R10571 gnd.n27 gnd.t239 2.82907
R10572 gnd.n27 gnd.t52 2.82907
R10573 gnd.n3432 gnd.n3431 2.71565
R10574 gnd.n3400 gnd.n3399 2.71565
R10575 gnd.n3368 gnd.n3367 2.71565
R10576 gnd.n3337 gnd.n3336 2.71565
R10577 gnd.n3305 gnd.n3304 2.71565
R10578 gnd.n3273 gnd.n3272 2.71565
R10579 gnd.n3241 gnd.n3240 2.71565
R10580 gnd.n3210 gnd.n3209 2.71565
R10581 gnd.n4319 gnd.n4318 2.54975
R10582 gnd.n4430 gnd.t262 2.54975
R10583 gnd.n4484 gnd.n1792 2.54975
R10584 gnd.n4509 gnd.t235 2.54975
R10585 gnd.n4533 gnd.n1753 2.54975
R10586 gnd.n1754 gnd.t36 2.54975
R10587 gnd.n4608 gnd.n1712 2.54975
R10588 gnd.n4656 gnd.n1672 2.54975
R10589 gnd.t231 gnd.n1629 2.54975
R10590 gnd.n4719 gnd.n1630 2.54975
R10591 gnd.n4741 gnd.t14 2.54975
R10592 gnd.n4815 gnd.n1583 2.54975
R10593 gnd.t248 gnd.n1558 2.54975
R10594 gnd.n4879 gnd.n4878 2.54975
R10595 gnd.n2966 gnd.n2388 2.27742
R10596 gnd.n2966 gnd.n2351 2.27742
R10597 gnd.n2966 gnd.n2350 2.27742
R10598 gnd.n2966 gnd.n2349 2.27742
R10599 gnd.n6557 gnd.n218 2.27742
R10600 gnd.n6557 gnd.n217 2.27742
R10601 gnd.n6557 gnd.n216 2.27742
R10602 gnd.n6557 gnd.n215 2.27742
R10603 gnd.n6557 gnd.n214 2.27742
R10604 gnd.n2045 gnd.n1006 2.27742
R10605 gnd.n3960 gnd.n1006 2.27742
R10606 gnd.n2027 gnd.n1006 2.27742
R10607 gnd.n3995 gnd.n1006 2.27742
R10608 gnd.n1006 gnd.n1005 2.27742
R10609 gnd.n2820 gnd.t81 2.23109
R10610 gnd.n2443 gnd.t68 2.23109
R10611 gnd.n4582 gnd.t236 2.23109
R10612 gnd.t229 gnd.n4675 2.23109
R10613 gnd.n3428 gnd.n3418 1.93989
R10614 gnd.n3396 gnd.n3386 1.93989
R10615 gnd.n3364 gnd.n3354 1.93989
R10616 gnd.n3333 gnd.n3323 1.93989
R10617 gnd.n3301 gnd.n3291 1.93989
R10618 gnd.n3269 gnd.n3259 1.93989
R10619 gnd.n3237 gnd.n3227 1.93989
R10620 gnd.n3206 gnd.n3196 1.93989
R10621 gnd.t287 gnd.n2831 1.59378
R10622 gnd.n3010 gnd.t185 1.59378
R10623 gnd.n2284 gnd.t63 1.59378
R10624 gnd.t78 gnd.n5333 1.27512
R10625 gnd.n5333 gnd.n5332 1.27512
R10626 gnd.n1308 gnd.n1302 1.27512
R10627 gnd.n4490 gnd.n1779 1.27512
R10628 gnd.n4502 gnd.n1769 1.27512
R10629 gnd.n4614 gnd.n1700 1.27512
R10630 gnd.n4626 gnd.n1689 1.27512
R10631 gnd.n4726 gnd.n4725 1.27512
R10632 gnd.n4805 gnd.n4804 1.27512
R10633 gnd.n4914 gnd.n4913 1.27512
R10634 gnd.n4936 gnd.n1513 1.27512
R10635 gnd.n2673 gnd.n2665 1.16414
R10636 gnd.n3490 gnd.n2187 1.16414
R10637 gnd.n3427 gnd.n3420 1.16414
R10638 gnd.n3395 gnd.n3388 1.16414
R10639 gnd.n3363 gnd.n3356 1.16414
R10640 gnd.n3332 gnd.n3325 1.16414
R10641 gnd.n3300 gnd.n3293 1.16414
R10642 gnd.n3268 gnd.n3261 1.16414
R10643 gnd.n3236 gnd.n3229 1.16414
R10644 gnd.n3205 gnd.n3198 1.16414
R10645 gnd.n6359 gnd.n6358 0.970197
R10646 gnd.n5408 gnd.n1140 0.970197
R10647 gnd.n3411 gnd.n3379 0.962709
R10648 gnd.n3443 gnd.n3411 0.962709
R10649 gnd.n3284 gnd.n3252 0.962709
R10650 gnd.n3316 gnd.n3284 0.962709
R10651 gnd.n2919 gnd.t190 0.956468
R10652 gnd.n3084 gnd.t188 0.956468
R10653 gnd.n3919 gnd.t232 0.956468
R10654 gnd.n5469 gnd.t60 0.956468
R10655 gnd.n4272 gnd.t203 0.956468
R10656 gnd.n4319 gnd.t240 0.956468
R10657 gnd.n4878 gnd.t48 0.956468
R10658 gnd.n4930 gnd.t280 0.956468
R10659 gnd.n497 gnd.t32 0.956468
R10660 gnd.t40 gnd.n186 0.956468
R10661 gnd.n2382 gnd.n2380 0.773756
R10662 gnd.n46 gnd.n44 0.773756
R10663 gnd.n2385 gnd.n2384 0.773756
R10664 gnd.n2384 gnd.n2382 0.773756
R10665 gnd.n2380 gnd.n2378 0.773756
R10666 gnd.n2378 gnd.n2376 0.773756
R10667 gnd.n42 gnd.n40 0.773756
R10668 gnd.n44 gnd.n42 0.773756
R10669 gnd.n48 gnd.n46 0.773756
R10670 gnd.n49 gnd.n48 0.773756
R10671 gnd.n2 gnd.n1 0.672012
R10672 gnd.n3 gnd.n2 0.672012
R10673 gnd.n4 gnd.n3 0.672012
R10674 gnd.n5 gnd.n4 0.672012
R10675 gnd.n6 gnd.n5 0.672012
R10676 gnd.n7 gnd.n6 0.672012
R10677 gnd.n9 gnd.n8 0.672012
R10678 gnd.n10 gnd.n9 0.672012
R10679 gnd.n11 gnd.n10 0.672012
R10680 gnd.n12 gnd.n11 0.672012
R10681 gnd.n13 gnd.n12 0.672012
R10682 gnd.n14 gnd.n13 0.672012
R10683 gnd.n5326 gnd.t117 0.637812
R10684 gnd.n4449 gnd.t19 0.637812
R10685 gnd.t28 gnd.n1709 0.637812
R10686 gnd.n1673 gnd.t242 0.637812
R10687 gnd.t6 gnd.n4840 0.637812
R10688 gnd.n4898 gnd.t99 0.637812
R10689 gnd.n2362 gnd.n2361 0.573776
R10690 gnd.n2361 gnd.n2359 0.573776
R10691 gnd.n2359 gnd.n2357 0.573776
R10692 gnd.n2357 gnd.n2355 0.573776
R10693 gnd.n2355 gnd.n2353 0.573776
R10694 gnd.n2373 gnd.n2372 0.573776
R10695 gnd.n2372 gnd.n2370 0.573776
R10696 gnd.n2370 gnd.n2368 0.573776
R10697 gnd.n2368 gnd.n2366 0.573776
R10698 gnd.n2366 gnd.n2364 0.573776
R10699 gnd.n19 gnd.n17 0.573776
R10700 gnd.n21 gnd.n19 0.573776
R10701 gnd.n23 gnd.n21 0.573776
R10702 gnd.n25 gnd.n23 0.573776
R10703 gnd.n26 gnd.n25 0.573776
R10704 gnd.n30 gnd.n28 0.573776
R10705 gnd.n32 gnd.n30 0.573776
R10706 gnd.n34 gnd.n32 0.573776
R10707 gnd.n36 gnd.n34 0.573776
R10708 gnd.n37 gnd.n36 0.573776
R10709 gnd gnd.n0 0.551497
R10710 gnd.n6557 gnd.n213 0.5435
R10711 gnd.n4034 gnd.n1006 0.5435
R10712 gnd.n3704 gnd.n3703 0.532512
R10713 gnd.n3883 gnd.n3882 0.532512
R10714 gnd.n6667 gnd.n6666 0.532512
R10715 gnd.n6767 gnd.n78 0.532512
R10716 gnd.n4254 gnd.n1836 0.523366
R10717 gnd.n5194 gnd.n333 0.523366
R10718 gnd.n6761 gnd.n6760 0.520317
R10719 gnd.n6690 gnd.n6689 0.520317
R10720 gnd.n6319 gnd.n6316 0.520317
R10721 gnd.n6448 gnd.n326 0.520317
R10722 gnd.n5441 gnd.n5440 0.520317
R10723 gnd.n4144 gnd.n4143 0.520317
R10724 gnd.n3802 gnd.n3752 0.520317
R10725 gnd.n3709 gnd.n2109 0.520317
R10726 gnd.n5200 gnd.n1416 0.489829
R10727 gnd.n4231 gnd.n4230 0.489829
R10728 gnd.n3146 gnd.n2191 0.486781
R10729 gnd.n2722 gnd.n2721 0.48678
R10730 gnd.n3464 gnd.n2145 0.480683
R10731 gnd.n2806 gnd.n2805 0.480683
R10732 gnd.n6800 gnd.n6799 0.470187
R10733 gnd.n1909 gnd.n1908 0.432431
R10734 gnd.n6442 gnd.n6441 0.432431
R10735 gnd.n5666 gnd.n5665 0.416659
R10736 gnd.n5988 gnd.n5987 0.416659
R10737 gnd.n4210 gnd.n4209 0.388379
R10738 gnd.n3424 gnd.n3423 0.388379
R10739 gnd.n3392 gnd.n3391 0.388379
R10740 gnd.n3360 gnd.n3359 0.388379
R10741 gnd.n3329 gnd.n3328 0.388379
R10742 gnd.n3297 gnd.n3296 0.388379
R10743 gnd.n3265 gnd.n3264 0.388379
R10744 gnd.n3233 gnd.n3232 0.388379
R10745 gnd.n3202 gnd.n3201 0.388379
R10746 gnd.n6730 gnd.n6729 0.388379
R10747 gnd.n3843 gnd.n3842 0.388379
R10748 gnd.n5171 gnd.n5170 0.388379
R10749 gnd.n6800 gnd.n15 0.374463
R10750 gnd.n2246 gnd.t9 0.319156
R10751 gnd.n3956 gnd.t218 0.319156
R10752 gnd.t17 gnd.n5493 0.319156
R10753 gnd.n4541 gnd.t56 0.319156
R10754 gnd.t20 gnd.t215 0.319156
R10755 gnd.t251 gnd.t200 0.319156
R10756 gnd.n4713 gnd.t253 0.319156
R10757 gnd.n6519 gnd.t246 0.319156
R10758 gnd.t7 gnd.n222 0.319156
R10759 gnd.n2640 gnd.n2618 0.311721
R10760 gnd.n4198 gnd.n1874 0.302329
R10761 gnd.n5155 gnd.n5154 0.302329
R10762 gnd gnd.n6800 0.295112
R10763 gnd.n6199 gnd.n213 0.280988
R10764 gnd.n4034 gnd.n996 0.280988
R10765 gnd.n3535 gnd.n3534 0.268793
R10766 gnd.n3534 gnd.n3533 0.241354
R10767 gnd.n437 gnd.n434 0.229039
R10768 gnd.n440 gnd.n437 0.229039
R10769 gnd.n1144 gnd.n1139 0.229039
R10770 gnd.n4095 gnd.n1144 0.229039
R10771 gnd.n2794 gnd.n2593 0.206293
R10772 gnd.n3441 gnd.n3413 0.155672
R10773 gnd.n3434 gnd.n3413 0.155672
R10774 gnd.n3434 gnd.n3433 0.155672
R10775 gnd.n3433 gnd.n3417 0.155672
R10776 gnd.n3426 gnd.n3417 0.155672
R10777 gnd.n3426 gnd.n3425 0.155672
R10778 gnd.n3409 gnd.n3381 0.155672
R10779 gnd.n3402 gnd.n3381 0.155672
R10780 gnd.n3402 gnd.n3401 0.155672
R10781 gnd.n3401 gnd.n3385 0.155672
R10782 gnd.n3394 gnd.n3385 0.155672
R10783 gnd.n3394 gnd.n3393 0.155672
R10784 gnd.n3377 gnd.n3349 0.155672
R10785 gnd.n3370 gnd.n3349 0.155672
R10786 gnd.n3370 gnd.n3369 0.155672
R10787 gnd.n3369 gnd.n3353 0.155672
R10788 gnd.n3362 gnd.n3353 0.155672
R10789 gnd.n3362 gnd.n3361 0.155672
R10790 gnd.n3346 gnd.n3318 0.155672
R10791 gnd.n3339 gnd.n3318 0.155672
R10792 gnd.n3339 gnd.n3338 0.155672
R10793 gnd.n3338 gnd.n3322 0.155672
R10794 gnd.n3331 gnd.n3322 0.155672
R10795 gnd.n3331 gnd.n3330 0.155672
R10796 gnd.n3314 gnd.n3286 0.155672
R10797 gnd.n3307 gnd.n3286 0.155672
R10798 gnd.n3307 gnd.n3306 0.155672
R10799 gnd.n3306 gnd.n3290 0.155672
R10800 gnd.n3299 gnd.n3290 0.155672
R10801 gnd.n3299 gnd.n3298 0.155672
R10802 gnd.n3282 gnd.n3254 0.155672
R10803 gnd.n3275 gnd.n3254 0.155672
R10804 gnd.n3275 gnd.n3274 0.155672
R10805 gnd.n3274 gnd.n3258 0.155672
R10806 gnd.n3267 gnd.n3258 0.155672
R10807 gnd.n3267 gnd.n3266 0.155672
R10808 gnd.n3250 gnd.n3222 0.155672
R10809 gnd.n3243 gnd.n3222 0.155672
R10810 gnd.n3243 gnd.n3242 0.155672
R10811 gnd.n3242 gnd.n3226 0.155672
R10812 gnd.n3235 gnd.n3226 0.155672
R10813 gnd.n3235 gnd.n3234 0.155672
R10814 gnd.n3219 gnd.n3191 0.155672
R10815 gnd.n3212 gnd.n3191 0.155672
R10816 gnd.n3212 gnd.n3211 0.155672
R10817 gnd.n3211 gnd.n3195 0.155672
R10818 gnd.n3204 gnd.n3195 0.155672
R10819 gnd.n3204 gnd.n3203 0.155672
R10820 gnd.n3566 gnd.n2145 0.152939
R10821 gnd.n3566 gnd.n3565 0.152939
R10822 gnd.n3565 gnd.n3564 0.152939
R10823 gnd.n3564 gnd.n2147 0.152939
R10824 gnd.n2148 gnd.n2147 0.152939
R10825 gnd.n2149 gnd.n2148 0.152939
R10826 gnd.n2150 gnd.n2149 0.152939
R10827 gnd.n2151 gnd.n2150 0.152939
R10828 gnd.n2152 gnd.n2151 0.152939
R10829 gnd.n2153 gnd.n2152 0.152939
R10830 gnd.n2154 gnd.n2153 0.152939
R10831 gnd.n2155 gnd.n2154 0.152939
R10832 gnd.n2156 gnd.n2155 0.152939
R10833 gnd.n2157 gnd.n2156 0.152939
R10834 gnd.n3536 gnd.n2157 0.152939
R10835 gnd.n3536 gnd.n3535 0.152939
R10836 gnd.n2807 gnd.n2806 0.152939
R10837 gnd.n2807 gnd.n2511 0.152939
R10838 gnd.n2835 gnd.n2511 0.152939
R10839 gnd.n2836 gnd.n2835 0.152939
R10840 gnd.n2837 gnd.n2836 0.152939
R10841 gnd.n2838 gnd.n2837 0.152939
R10842 gnd.n2838 gnd.n2483 0.152939
R10843 gnd.n2865 gnd.n2483 0.152939
R10844 gnd.n2866 gnd.n2865 0.152939
R10845 gnd.n2867 gnd.n2866 0.152939
R10846 gnd.n2867 gnd.n2461 0.152939
R10847 gnd.n2896 gnd.n2461 0.152939
R10848 gnd.n2897 gnd.n2896 0.152939
R10849 gnd.n2898 gnd.n2897 0.152939
R10850 gnd.n2899 gnd.n2898 0.152939
R10851 gnd.n2901 gnd.n2899 0.152939
R10852 gnd.n2901 gnd.n2900 0.152939
R10853 gnd.n2900 gnd.n2410 0.152939
R10854 gnd.n2411 gnd.n2410 0.152939
R10855 gnd.n2412 gnd.n2411 0.152939
R10856 gnd.n2431 gnd.n2412 0.152939
R10857 gnd.n2432 gnd.n2431 0.152939
R10858 gnd.n2432 gnd.n2342 0.152939
R10859 gnd.n2991 gnd.n2342 0.152939
R10860 gnd.n2992 gnd.n2991 0.152939
R10861 gnd.n2993 gnd.n2992 0.152939
R10862 gnd.n2994 gnd.n2993 0.152939
R10863 gnd.n2994 gnd.n2315 0.152939
R10864 gnd.n3031 gnd.n2315 0.152939
R10865 gnd.n3032 gnd.n3031 0.152939
R10866 gnd.n3033 gnd.n3032 0.152939
R10867 gnd.n3034 gnd.n3033 0.152939
R10868 gnd.n3034 gnd.n2288 0.152939
R10869 gnd.n3076 gnd.n2288 0.152939
R10870 gnd.n3077 gnd.n3076 0.152939
R10871 gnd.n3078 gnd.n3077 0.152939
R10872 gnd.n3079 gnd.n3078 0.152939
R10873 gnd.n3079 gnd.n2260 0.152939
R10874 gnd.n3116 gnd.n2260 0.152939
R10875 gnd.n3117 gnd.n3116 0.152939
R10876 gnd.n3118 gnd.n3117 0.152939
R10877 gnd.n3119 gnd.n3118 0.152939
R10878 gnd.n3119 gnd.n2233 0.152939
R10879 gnd.n3165 gnd.n2233 0.152939
R10880 gnd.n3166 gnd.n3165 0.152939
R10881 gnd.n3167 gnd.n3166 0.152939
R10882 gnd.n3168 gnd.n3167 0.152939
R10883 gnd.n3168 gnd.n2206 0.152939
R10884 gnd.n3460 gnd.n2206 0.152939
R10885 gnd.n3461 gnd.n3460 0.152939
R10886 gnd.n3462 gnd.n3461 0.152939
R10887 gnd.n3463 gnd.n3462 0.152939
R10888 gnd.n3464 gnd.n3463 0.152939
R10889 gnd.n2805 gnd.n2535 0.152939
R10890 gnd.n2556 gnd.n2535 0.152939
R10891 gnd.n2557 gnd.n2556 0.152939
R10892 gnd.n2563 gnd.n2557 0.152939
R10893 gnd.n2564 gnd.n2563 0.152939
R10894 gnd.n2565 gnd.n2564 0.152939
R10895 gnd.n2565 gnd.n2554 0.152939
R10896 gnd.n2573 gnd.n2554 0.152939
R10897 gnd.n2574 gnd.n2573 0.152939
R10898 gnd.n2575 gnd.n2574 0.152939
R10899 gnd.n2575 gnd.n2552 0.152939
R10900 gnd.n2583 gnd.n2552 0.152939
R10901 gnd.n2584 gnd.n2583 0.152939
R10902 gnd.n2585 gnd.n2584 0.152939
R10903 gnd.n2585 gnd.n2550 0.152939
R10904 gnd.n2593 gnd.n2550 0.152939
R10905 gnd.n3533 gnd.n2162 0.152939
R10906 gnd.n2164 gnd.n2162 0.152939
R10907 gnd.n2165 gnd.n2164 0.152939
R10908 gnd.n2166 gnd.n2165 0.152939
R10909 gnd.n2167 gnd.n2166 0.152939
R10910 gnd.n2168 gnd.n2167 0.152939
R10911 gnd.n2169 gnd.n2168 0.152939
R10912 gnd.n2170 gnd.n2169 0.152939
R10913 gnd.n2171 gnd.n2170 0.152939
R10914 gnd.n2172 gnd.n2171 0.152939
R10915 gnd.n2173 gnd.n2172 0.152939
R10916 gnd.n2174 gnd.n2173 0.152939
R10917 gnd.n2175 gnd.n2174 0.152939
R10918 gnd.n2176 gnd.n2175 0.152939
R10919 gnd.n2177 gnd.n2176 0.152939
R10920 gnd.n2178 gnd.n2177 0.152939
R10921 gnd.n2179 gnd.n2178 0.152939
R10922 gnd.n2180 gnd.n2179 0.152939
R10923 gnd.n2181 gnd.n2180 0.152939
R10924 gnd.n2182 gnd.n2181 0.152939
R10925 gnd.n2183 gnd.n2182 0.152939
R10926 gnd.n2184 gnd.n2183 0.152939
R10927 gnd.n2188 gnd.n2184 0.152939
R10928 gnd.n2189 gnd.n2188 0.152939
R10929 gnd.n2190 gnd.n2189 0.152939
R10930 gnd.n2191 gnd.n2190 0.152939
R10931 gnd.n2968 gnd.n2967 0.152939
R10932 gnd.n2969 gnd.n2968 0.152939
R10933 gnd.n2970 gnd.n2969 0.152939
R10934 gnd.n2971 gnd.n2970 0.152939
R10935 gnd.n2972 gnd.n2971 0.152939
R10936 gnd.n2973 gnd.n2972 0.152939
R10937 gnd.n2973 gnd.n2296 0.152939
R10938 gnd.n3052 gnd.n2296 0.152939
R10939 gnd.n3053 gnd.n3052 0.152939
R10940 gnd.n3054 gnd.n3053 0.152939
R10941 gnd.n3055 gnd.n3054 0.152939
R10942 gnd.n3056 gnd.n3055 0.152939
R10943 gnd.n3057 gnd.n3056 0.152939
R10944 gnd.n3058 gnd.n3057 0.152939
R10945 gnd.n3059 gnd.n3058 0.152939
R10946 gnd.n3060 gnd.n3059 0.152939
R10947 gnd.n3060 gnd.n2240 0.152939
R10948 gnd.n3137 gnd.n2240 0.152939
R10949 gnd.n3138 gnd.n3137 0.152939
R10950 gnd.n3139 gnd.n3138 0.152939
R10951 gnd.n3140 gnd.n3139 0.152939
R10952 gnd.n3141 gnd.n3140 0.152939
R10953 gnd.n3142 gnd.n3141 0.152939
R10954 gnd.n3143 gnd.n3142 0.152939
R10955 gnd.n3144 gnd.n3143 0.152939
R10956 gnd.n3145 gnd.n3144 0.152939
R10957 gnd.n3147 gnd.n3145 0.152939
R10958 gnd.n3147 gnd.n3146 0.152939
R10959 gnd.n2723 gnd.n2722 0.152939
R10960 gnd.n2723 gnd.n2613 0.152939
R10961 gnd.n2738 gnd.n2613 0.152939
R10962 gnd.n2739 gnd.n2738 0.152939
R10963 gnd.n2740 gnd.n2739 0.152939
R10964 gnd.n2740 gnd.n2601 0.152939
R10965 gnd.n2754 gnd.n2601 0.152939
R10966 gnd.n2755 gnd.n2754 0.152939
R10967 gnd.n2756 gnd.n2755 0.152939
R10968 gnd.n2757 gnd.n2756 0.152939
R10969 gnd.n2758 gnd.n2757 0.152939
R10970 gnd.n2759 gnd.n2758 0.152939
R10971 gnd.n2760 gnd.n2759 0.152939
R10972 gnd.n2761 gnd.n2760 0.152939
R10973 gnd.n2762 gnd.n2761 0.152939
R10974 gnd.n2763 gnd.n2762 0.152939
R10975 gnd.n2764 gnd.n2763 0.152939
R10976 gnd.n2765 gnd.n2764 0.152939
R10977 gnd.n2766 gnd.n2765 0.152939
R10978 gnd.n2767 gnd.n2766 0.152939
R10979 gnd.n2768 gnd.n2767 0.152939
R10980 gnd.n2768 gnd.n2467 0.152939
R10981 gnd.n2885 gnd.n2467 0.152939
R10982 gnd.n2886 gnd.n2885 0.152939
R10983 gnd.n2887 gnd.n2886 0.152939
R10984 gnd.n2888 gnd.n2887 0.152939
R10985 gnd.n2888 gnd.n2389 0.152939
R10986 gnd.n2965 gnd.n2389 0.152939
R10987 gnd.n2641 gnd.n2640 0.152939
R10988 gnd.n2642 gnd.n2641 0.152939
R10989 gnd.n2643 gnd.n2642 0.152939
R10990 gnd.n2644 gnd.n2643 0.152939
R10991 gnd.n2645 gnd.n2644 0.152939
R10992 gnd.n2646 gnd.n2645 0.152939
R10993 gnd.n2647 gnd.n2646 0.152939
R10994 gnd.n2648 gnd.n2647 0.152939
R10995 gnd.n2649 gnd.n2648 0.152939
R10996 gnd.n2650 gnd.n2649 0.152939
R10997 gnd.n2651 gnd.n2650 0.152939
R10998 gnd.n2652 gnd.n2651 0.152939
R10999 gnd.n2653 gnd.n2652 0.152939
R11000 gnd.n2654 gnd.n2653 0.152939
R11001 gnd.n2655 gnd.n2654 0.152939
R11002 gnd.n2656 gnd.n2655 0.152939
R11003 gnd.n2657 gnd.n2656 0.152939
R11004 gnd.n2658 gnd.n2657 0.152939
R11005 gnd.n2659 gnd.n2658 0.152939
R11006 gnd.n2660 gnd.n2659 0.152939
R11007 gnd.n2661 gnd.n2660 0.152939
R11008 gnd.n2662 gnd.n2661 0.152939
R11009 gnd.n2666 gnd.n2662 0.152939
R11010 gnd.n2667 gnd.n2666 0.152939
R11011 gnd.n2667 gnd.n2624 0.152939
R11012 gnd.n2721 gnd.n2624 0.152939
R11013 gnd.n5667 gnd.n5666 0.152939
R11014 gnd.n5667 gnd.n823 0.152939
R11015 gnd.n5675 gnd.n823 0.152939
R11016 gnd.n5676 gnd.n5675 0.152939
R11017 gnd.n5677 gnd.n5676 0.152939
R11018 gnd.n5677 gnd.n817 0.152939
R11019 gnd.n5685 gnd.n817 0.152939
R11020 gnd.n5686 gnd.n5685 0.152939
R11021 gnd.n5687 gnd.n5686 0.152939
R11022 gnd.n5687 gnd.n811 0.152939
R11023 gnd.n5695 gnd.n811 0.152939
R11024 gnd.n5696 gnd.n5695 0.152939
R11025 gnd.n5697 gnd.n5696 0.152939
R11026 gnd.n5697 gnd.n805 0.152939
R11027 gnd.n5705 gnd.n805 0.152939
R11028 gnd.n5706 gnd.n5705 0.152939
R11029 gnd.n5707 gnd.n5706 0.152939
R11030 gnd.n5707 gnd.n799 0.152939
R11031 gnd.n5715 gnd.n799 0.152939
R11032 gnd.n5716 gnd.n5715 0.152939
R11033 gnd.n5717 gnd.n5716 0.152939
R11034 gnd.n5717 gnd.n793 0.152939
R11035 gnd.n5725 gnd.n793 0.152939
R11036 gnd.n5726 gnd.n5725 0.152939
R11037 gnd.n5727 gnd.n5726 0.152939
R11038 gnd.n5727 gnd.n787 0.152939
R11039 gnd.n5735 gnd.n787 0.152939
R11040 gnd.n5736 gnd.n5735 0.152939
R11041 gnd.n5737 gnd.n5736 0.152939
R11042 gnd.n5737 gnd.n781 0.152939
R11043 gnd.n5745 gnd.n781 0.152939
R11044 gnd.n5746 gnd.n5745 0.152939
R11045 gnd.n5747 gnd.n5746 0.152939
R11046 gnd.n5747 gnd.n775 0.152939
R11047 gnd.n5755 gnd.n775 0.152939
R11048 gnd.n5756 gnd.n5755 0.152939
R11049 gnd.n5757 gnd.n5756 0.152939
R11050 gnd.n5757 gnd.n769 0.152939
R11051 gnd.n5765 gnd.n769 0.152939
R11052 gnd.n5766 gnd.n5765 0.152939
R11053 gnd.n5767 gnd.n5766 0.152939
R11054 gnd.n5767 gnd.n763 0.152939
R11055 gnd.n5775 gnd.n763 0.152939
R11056 gnd.n5776 gnd.n5775 0.152939
R11057 gnd.n5777 gnd.n5776 0.152939
R11058 gnd.n5777 gnd.n757 0.152939
R11059 gnd.n5785 gnd.n757 0.152939
R11060 gnd.n5786 gnd.n5785 0.152939
R11061 gnd.n5787 gnd.n5786 0.152939
R11062 gnd.n5787 gnd.n751 0.152939
R11063 gnd.n5795 gnd.n751 0.152939
R11064 gnd.n5796 gnd.n5795 0.152939
R11065 gnd.n5797 gnd.n5796 0.152939
R11066 gnd.n5797 gnd.n745 0.152939
R11067 gnd.n5805 gnd.n745 0.152939
R11068 gnd.n5806 gnd.n5805 0.152939
R11069 gnd.n5807 gnd.n5806 0.152939
R11070 gnd.n5807 gnd.n739 0.152939
R11071 gnd.n5815 gnd.n739 0.152939
R11072 gnd.n5816 gnd.n5815 0.152939
R11073 gnd.n5817 gnd.n5816 0.152939
R11074 gnd.n5817 gnd.n733 0.152939
R11075 gnd.n5825 gnd.n733 0.152939
R11076 gnd.n5826 gnd.n5825 0.152939
R11077 gnd.n5827 gnd.n5826 0.152939
R11078 gnd.n5827 gnd.n727 0.152939
R11079 gnd.n5835 gnd.n727 0.152939
R11080 gnd.n5836 gnd.n5835 0.152939
R11081 gnd.n5837 gnd.n5836 0.152939
R11082 gnd.n5837 gnd.n721 0.152939
R11083 gnd.n5845 gnd.n721 0.152939
R11084 gnd.n5846 gnd.n5845 0.152939
R11085 gnd.n5847 gnd.n5846 0.152939
R11086 gnd.n5847 gnd.n715 0.152939
R11087 gnd.n5855 gnd.n715 0.152939
R11088 gnd.n5856 gnd.n5855 0.152939
R11089 gnd.n5857 gnd.n5856 0.152939
R11090 gnd.n5857 gnd.n709 0.152939
R11091 gnd.n5865 gnd.n709 0.152939
R11092 gnd.n5866 gnd.n5865 0.152939
R11093 gnd.n5867 gnd.n5866 0.152939
R11094 gnd.n5867 gnd.n703 0.152939
R11095 gnd.n5875 gnd.n703 0.152939
R11096 gnd.n5876 gnd.n5875 0.152939
R11097 gnd.n5877 gnd.n5876 0.152939
R11098 gnd.n5877 gnd.n697 0.152939
R11099 gnd.n5885 gnd.n697 0.152939
R11100 gnd.n5886 gnd.n5885 0.152939
R11101 gnd.n5887 gnd.n5886 0.152939
R11102 gnd.n5887 gnd.n691 0.152939
R11103 gnd.n5895 gnd.n691 0.152939
R11104 gnd.n5896 gnd.n5895 0.152939
R11105 gnd.n5897 gnd.n5896 0.152939
R11106 gnd.n5897 gnd.n685 0.152939
R11107 gnd.n5905 gnd.n685 0.152939
R11108 gnd.n5906 gnd.n5905 0.152939
R11109 gnd.n5907 gnd.n5906 0.152939
R11110 gnd.n5907 gnd.n679 0.152939
R11111 gnd.n5915 gnd.n679 0.152939
R11112 gnd.n5916 gnd.n5915 0.152939
R11113 gnd.n5917 gnd.n5916 0.152939
R11114 gnd.n5917 gnd.n673 0.152939
R11115 gnd.n5925 gnd.n673 0.152939
R11116 gnd.n5926 gnd.n5925 0.152939
R11117 gnd.n5927 gnd.n5926 0.152939
R11118 gnd.n5927 gnd.n667 0.152939
R11119 gnd.n5935 gnd.n667 0.152939
R11120 gnd.n5936 gnd.n5935 0.152939
R11121 gnd.n5937 gnd.n5936 0.152939
R11122 gnd.n5937 gnd.n661 0.152939
R11123 gnd.n5945 gnd.n661 0.152939
R11124 gnd.n5946 gnd.n5945 0.152939
R11125 gnd.n5947 gnd.n5946 0.152939
R11126 gnd.n5947 gnd.n655 0.152939
R11127 gnd.n5955 gnd.n655 0.152939
R11128 gnd.n5956 gnd.n5955 0.152939
R11129 gnd.n5957 gnd.n5956 0.152939
R11130 gnd.n5957 gnd.n649 0.152939
R11131 gnd.n5965 gnd.n649 0.152939
R11132 gnd.n5966 gnd.n5965 0.152939
R11133 gnd.n5967 gnd.n5966 0.152939
R11134 gnd.n5967 gnd.n643 0.152939
R11135 gnd.n5975 gnd.n643 0.152939
R11136 gnd.n5976 gnd.n5975 0.152939
R11137 gnd.n5978 gnd.n5976 0.152939
R11138 gnd.n5978 gnd.n5977 0.152939
R11139 gnd.n5977 gnd.n637 0.152939
R11140 gnd.n5987 gnd.n637 0.152939
R11141 gnd.n5988 gnd.n632 0.152939
R11142 gnd.n5996 gnd.n632 0.152939
R11143 gnd.n5997 gnd.n5996 0.152939
R11144 gnd.n5998 gnd.n5997 0.152939
R11145 gnd.n5998 gnd.n626 0.152939
R11146 gnd.n6006 gnd.n626 0.152939
R11147 gnd.n6007 gnd.n6006 0.152939
R11148 gnd.n6008 gnd.n6007 0.152939
R11149 gnd.n6008 gnd.n620 0.152939
R11150 gnd.n6016 gnd.n620 0.152939
R11151 gnd.n6017 gnd.n6016 0.152939
R11152 gnd.n6018 gnd.n6017 0.152939
R11153 gnd.n6018 gnd.n614 0.152939
R11154 gnd.n6026 gnd.n614 0.152939
R11155 gnd.n6027 gnd.n6026 0.152939
R11156 gnd.n6028 gnd.n6027 0.152939
R11157 gnd.n6028 gnd.n608 0.152939
R11158 gnd.n6036 gnd.n608 0.152939
R11159 gnd.n6037 gnd.n6036 0.152939
R11160 gnd.n6038 gnd.n6037 0.152939
R11161 gnd.n6038 gnd.n602 0.152939
R11162 gnd.n6046 gnd.n602 0.152939
R11163 gnd.n6047 gnd.n6046 0.152939
R11164 gnd.n6048 gnd.n6047 0.152939
R11165 gnd.n6048 gnd.n596 0.152939
R11166 gnd.n6056 gnd.n596 0.152939
R11167 gnd.n6057 gnd.n6056 0.152939
R11168 gnd.n6058 gnd.n6057 0.152939
R11169 gnd.n6058 gnd.n590 0.152939
R11170 gnd.n6066 gnd.n590 0.152939
R11171 gnd.n6067 gnd.n6066 0.152939
R11172 gnd.n6068 gnd.n6067 0.152939
R11173 gnd.n6068 gnd.n584 0.152939
R11174 gnd.n6076 gnd.n584 0.152939
R11175 gnd.n6077 gnd.n6076 0.152939
R11176 gnd.n6078 gnd.n6077 0.152939
R11177 gnd.n6078 gnd.n578 0.152939
R11178 gnd.n6086 gnd.n578 0.152939
R11179 gnd.n6087 gnd.n6086 0.152939
R11180 gnd.n6088 gnd.n6087 0.152939
R11181 gnd.n6088 gnd.n572 0.152939
R11182 gnd.n6096 gnd.n572 0.152939
R11183 gnd.n6097 gnd.n6096 0.152939
R11184 gnd.n6098 gnd.n6097 0.152939
R11185 gnd.n6098 gnd.n566 0.152939
R11186 gnd.n6106 gnd.n566 0.152939
R11187 gnd.n6107 gnd.n6106 0.152939
R11188 gnd.n6108 gnd.n6107 0.152939
R11189 gnd.n6108 gnd.n560 0.152939
R11190 gnd.n6116 gnd.n560 0.152939
R11191 gnd.n6117 gnd.n6116 0.152939
R11192 gnd.n6118 gnd.n6117 0.152939
R11193 gnd.n6118 gnd.n554 0.152939
R11194 gnd.n6126 gnd.n554 0.152939
R11195 gnd.n6127 gnd.n6126 0.152939
R11196 gnd.n6128 gnd.n6127 0.152939
R11197 gnd.n6128 gnd.n548 0.152939
R11198 gnd.n6136 gnd.n548 0.152939
R11199 gnd.n6137 gnd.n6136 0.152939
R11200 gnd.n6138 gnd.n6137 0.152939
R11201 gnd.n6138 gnd.n542 0.152939
R11202 gnd.n6146 gnd.n542 0.152939
R11203 gnd.n6147 gnd.n6146 0.152939
R11204 gnd.n6148 gnd.n6147 0.152939
R11205 gnd.n6148 gnd.n536 0.152939
R11206 gnd.n6156 gnd.n536 0.152939
R11207 gnd.n6157 gnd.n6156 0.152939
R11208 gnd.n6158 gnd.n6157 0.152939
R11209 gnd.n6158 gnd.n530 0.152939
R11210 gnd.n6166 gnd.n530 0.152939
R11211 gnd.n6167 gnd.n6166 0.152939
R11212 gnd.n6168 gnd.n6167 0.152939
R11213 gnd.n6168 gnd.n524 0.152939
R11214 gnd.n6176 gnd.n524 0.152939
R11215 gnd.n6177 gnd.n6176 0.152939
R11216 gnd.n6178 gnd.n6177 0.152939
R11217 gnd.n6178 gnd.n518 0.152939
R11218 gnd.n6186 gnd.n518 0.152939
R11219 gnd.n6187 gnd.n6186 0.152939
R11220 gnd.n6188 gnd.n6187 0.152939
R11221 gnd.n6188 gnd.n512 0.152939
R11222 gnd.n6197 gnd.n512 0.152939
R11223 gnd.n6198 gnd.n6197 0.152939
R11224 gnd.n6199 gnd.n6198 0.152939
R11225 gnd.n6558 gnd.n6557 0.152939
R11226 gnd.n6559 gnd.n6558 0.152939
R11227 gnd.n6559 gnd.n198 0.152939
R11228 gnd.n6573 gnd.n198 0.152939
R11229 gnd.n6574 gnd.n6573 0.152939
R11230 gnd.n6575 gnd.n6574 0.152939
R11231 gnd.n6575 gnd.n182 0.152939
R11232 gnd.n6589 gnd.n182 0.152939
R11233 gnd.n6590 gnd.n6589 0.152939
R11234 gnd.n6591 gnd.n6590 0.152939
R11235 gnd.n6591 gnd.n165 0.152939
R11236 gnd.n6679 gnd.n165 0.152939
R11237 gnd.n6680 gnd.n6679 0.152939
R11238 gnd.n6681 gnd.n6680 0.152939
R11239 gnd.n6681 gnd.n88 0.152939
R11240 gnd.n6761 gnd.n88 0.152939
R11241 gnd.n6760 gnd.n89 0.152939
R11242 gnd.n91 gnd.n89 0.152939
R11243 gnd.n95 gnd.n91 0.152939
R11244 gnd.n96 gnd.n95 0.152939
R11245 gnd.n97 gnd.n96 0.152939
R11246 gnd.n98 gnd.n97 0.152939
R11247 gnd.n102 gnd.n98 0.152939
R11248 gnd.n103 gnd.n102 0.152939
R11249 gnd.n104 gnd.n103 0.152939
R11250 gnd.n105 gnd.n104 0.152939
R11251 gnd.n109 gnd.n105 0.152939
R11252 gnd.n110 gnd.n109 0.152939
R11253 gnd.n111 gnd.n110 0.152939
R11254 gnd.n112 gnd.n111 0.152939
R11255 gnd.n116 gnd.n112 0.152939
R11256 gnd.n117 gnd.n116 0.152939
R11257 gnd.n118 gnd.n117 0.152939
R11258 gnd.n119 gnd.n118 0.152939
R11259 gnd.n123 gnd.n119 0.152939
R11260 gnd.n124 gnd.n123 0.152939
R11261 gnd.n125 gnd.n124 0.152939
R11262 gnd.n126 gnd.n125 0.152939
R11263 gnd.n130 gnd.n126 0.152939
R11264 gnd.n131 gnd.n130 0.152939
R11265 gnd.n132 gnd.n131 0.152939
R11266 gnd.n133 gnd.n132 0.152939
R11267 gnd.n137 gnd.n133 0.152939
R11268 gnd.n138 gnd.n137 0.152939
R11269 gnd.n139 gnd.n138 0.152939
R11270 gnd.n140 gnd.n139 0.152939
R11271 gnd.n144 gnd.n140 0.152939
R11272 gnd.n145 gnd.n144 0.152939
R11273 gnd.n146 gnd.n145 0.152939
R11274 gnd.n147 gnd.n146 0.152939
R11275 gnd.n151 gnd.n147 0.152939
R11276 gnd.n152 gnd.n151 0.152939
R11277 gnd.n6691 gnd.n152 0.152939
R11278 gnd.n6691 gnd.n6690 0.152939
R11279 gnd.n6316 gnd.n463 0.152939
R11280 gnd.n465 gnd.n463 0.152939
R11281 gnd.n466 gnd.n465 0.152939
R11282 gnd.n486 gnd.n466 0.152939
R11283 gnd.n490 gnd.n486 0.152939
R11284 gnd.n491 gnd.n490 0.152939
R11285 gnd.n492 gnd.n491 0.152939
R11286 gnd.n492 gnd.n484 0.152939
R11287 gnd.n500 gnd.n484 0.152939
R11288 gnd.n501 gnd.n500 0.152939
R11289 gnd.n502 gnd.n501 0.152939
R11290 gnd.n502 gnd.n482 0.152939
R11291 gnd.n6224 gnd.n482 0.152939
R11292 gnd.n6225 gnd.n6224 0.152939
R11293 gnd.n6226 gnd.n6225 0.152939
R11294 gnd.n6227 gnd.n6226 0.152939
R11295 gnd.n6228 gnd.n6227 0.152939
R11296 gnd.n6229 gnd.n6228 0.152939
R11297 gnd.n6230 gnd.n6229 0.152939
R11298 gnd.n6231 gnd.n6230 0.152939
R11299 gnd.n6231 gnd.n239 0.152939
R11300 gnd.n6232 gnd.n239 0.152939
R11301 gnd.n6233 gnd.n6232 0.152939
R11302 gnd.n6234 gnd.n6233 0.152939
R11303 gnd.n6235 gnd.n6234 0.152939
R11304 gnd.n6236 gnd.n6235 0.152939
R11305 gnd.n6237 gnd.n6236 0.152939
R11306 gnd.n6238 gnd.n6237 0.152939
R11307 gnd.n6239 gnd.n6238 0.152939
R11308 gnd.n6240 gnd.n6239 0.152939
R11309 gnd.n6241 gnd.n6240 0.152939
R11310 gnd.n6242 gnd.n6241 0.152939
R11311 gnd.n6243 gnd.n6242 0.152939
R11312 gnd.n6244 gnd.n6243 0.152939
R11313 gnd.n6245 gnd.n6244 0.152939
R11314 gnd.n6246 gnd.n6245 0.152939
R11315 gnd.n6247 gnd.n6246 0.152939
R11316 gnd.n6248 gnd.n6247 0.152939
R11317 gnd.n6250 gnd.n6248 0.152939
R11318 gnd.n6250 gnd.n6249 0.152939
R11319 gnd.n6249 gnd.n158 0.152939
R11320 gnd.n6689 gnd.n158 0.152939
R11321 gnd.n420 gnd.n326 0.152939
R11322 gnd.n421 gnd.n420 0.152939
R11323 gnd.n422 gnd.n421 0.152939
R11324 gnd.n423 gnd.n422 0.152939
R11325 gnd.n424 gnd.n423 0.152939
R11326 gnd.n425 gnd.n424 0.152939
R11327 gnd.n426 gnd.n425 0.152939
R11328 gnd.n427 gnd.n426 0.152939
R11329 gnd.n428 gnd.n427 0.152939
R11330 gnd.n429 gnd.n428 0.152939
R11331 gnd.n430 gnd.n429 0.152939
R11332 gnd.n431 gnd.n430 0.152939
R11333 gnd.n432 gnd.n431 0.152939
R11334 gnd.n433 gnd.n432 0.152939
R11335 gnd.n434 gnd.n433 0.152939
R11336 gnd.n441 gnd.n440 0.152939
R11337 gnd.n442 gnd.n441 0.152939
R11338 gnd.n443 gnd.n442 0.152939
R11339 gnd.n444 gnd.n443 0.152939
R11340 gnd.n445 gnd.n444 0.152939
R11341 gnd.n446 gnd.n445 0.152939
R11342 gnd.n447 gnd.n446 0.152939
R11343 gnd.n448 gnd.n447 0.152939
R11344 gnd.n449 gnd.n448 0.152939
R11345 gnd.n450 gnd.n449 0.152939
R11346 gnd.n451 gnd.n450 0.152939
R11347 gnd.n452 gnd.n451 0.152939
R11348 gnd.n453 gnd.n452 0.152939
R11349 gnd.n454 gnd.n453 0.152939
R11350 gnd.n455 gnd.n454 0.152939
R11351 gnd.n456 gnd.n455 0.152939
R11352 gnd.n457 gnd.n456 0.152939
R11353 gnd.n6321 gnd.n457 0.152939
R11354 gnd.n6321 gnd.n6320 0.152939
R11355 gnd.n6320 gnd.n6319 0.152939
R11356 gnd.n6449 gnd.n6448 0.152939
R11357 gnd.n6450 gnd.n6449 0.152939
R11358 gnd.n6450 gnd.n309 0.152939
R11359 gnd.n6464 gnd.n309 0.152939
R11360 gnd.n6465 gnd.n6464 0.152939
R11361 gnd.n6466 gnd.n6465 0.152939
R11362 gnd.n6466 gnd.n291 0.152939
R11363 gnd.n6480 gnd.n291 0.152939
R11364 gnd.n6481 gnd.n6480 0.152939
R11365 gnd.n6482 gnd.n6481 0.152939
R11366 gnd.n6482 gnd.n274 0.152939
R11367 gnd.n6496 gnd.n274 0.152939
R11368 gnd.n6497 gnd.n6496 0.152939
R11369 gnd.n6498 gnd.n6497 0.152939
R11370 gnd.n6498 gnd.n212 0.152939
R11371 gnd.n6557 gnd.n212 0.152939
R11372 gnd.n6206 gnd.n6205 0.152939
R11373 gnd.n4039 gnd.n4035 0.152939
R11374 gnd.n4040 gnd.n4039 0.152939
R11375 gnd.n4041 gnd.n4040 0.152939
R11376 gnd.n4041 gnd.n2010 0.152939
R11377 gnd.n4047 gnd.n2010 0.152939
R11378 gnd.n4048 gnd.n4047 0.152939
R11379 gnd.n4049 gnd.n4048 0.152939
R11380 gnd.n4050 gnd.n4049 0.152939
R11381 gnd.n4051 gnd.n4050 0.152939
R11382 gnd.n4051 gnd.n1989 0.152939
R11383 gnd.n4167 gnd.n1989 0.152939
R11384 gnd.n4168 gnd.n4167 0.152939
R11385 gnd.n4169 gnd.n4168 0.152939
R11386 gnd.n4169 gnd.n1985 0.152939
R11387 gnd.n4175 gnd.n1985 0.152939
R11388 gnd.n4176 gnd.n4175 0.152939
R11389 gnd.n4177 gnd.n4176 0.152939
R11390 gnd.n4178 gnd.n4177 0.152939
R11391 gnd.n4179 gnd.n4178 0.152939
R11392 gnd.n4179 gnd.n1844 0.152939
R11393 gnd.n4237 gnd.n1844 0.152939
R11394 gnd.n4238 gnd.n4237 0.152939
R11395 gnd.n4239 gnd.n4238 0.152939
R11396 gnd.n4240 gnd.n4239 0.152939
R11397 gnd.n4241 gnd.n4240 0.152939
R11398 gnd.n4243 gnd.n4241 0.152939
R11399 gnd.n4243 gnd.n4242 0.152939
R11400 gnd.n4242 gnd.n1216 0.152939
R11401 gnd.n1217 gnd.n1216 0.152939
R11402 gnd.n1218 gnd.n1217 0.152939
R11403 gnd.n1316 gnd.n1218 0.152939
R11404 gnd.n1317 gnd.n1316 0.152939
R11405 gnd.n1318 gnd.n1317 0.152939
R11406 gnd.n1319 gnd.n1318 0.152939
R11407 gnd.n1320 gnd.n1319 0.152939
R11408 gnd.n4433 gnd.n1320 0.152939
R11409 gnd.n4434 gnd.n4433 0.152939
R11410 gnd.n4435 gnd.n4434 0.152939
R11411 gnd.n4435 gnd.n1802 0.152939
R11412 gnd.n4462 gnd.n1802 0.152939
R11413 gnd.n4463 gnd.n4462 0.152939
R11414 gnd.n4464 gnd.n4463 0.152939
R11415 gnd.n4465 gnd.n4464 0.152939
R11416 gnd.n4466 gnd.n4465 0.152939
R11417 gnd.n4468 gnd.n4466 0.152939
R11418 gnd.n4469 gnd.n4468 0.152939
R11419 gnd.n4469 gnd.n1764 0.152939
R11420 gnd.n4520 gnd.n1764 0.152939
R11421 gnd.n4521 gnd.n4520 0.152939
R11422 gnd.n4522 gnd.n4521 0.152939
R11423 gnd.n4522 gnd.n1746 0.152939
R11424 gnd.n4546 gnd.n1746 0.152939
R11425 gnd.n4547 gnd.n4546 0.152939
R11426 gnd.n4548 gnd.n4547 0.152939
R11427 gnd.n4549 gnd.n4548 0.152939
R11428 gnd.n4549 gnd.n1722 0.152939
R11429 gnd.n4585 gnd.n1722 0.152939
R11430 gnd.n4586 gnd.n4585 0.152939
R11431 gnd.n4587 gnd.n4586 0.152939
R11432 gnd.n4588 gnd.n4587 0.152939
R11433 gnd.n4589 gnd.n4588 0.152939
R11434 gnd.n4591 gnd.n4589 0.152939
R11435 gnd.n4592 gnd.n4591 0.152939
R11436 gnd.n4592 gnd.n1683 0.152939
R11437 gnd.n4643 gnd.n1683 0.152939
R11438 gnd.n4644 gnd.n4643 0.152939
R11439 gnd.n4645 gnd.n4644 0.152939
R11440 gnd.n4645 gnd.n1664 0.152939
R11441 gnd.n4668 gnd.n1664 0.152939
R11442 gnd.n4669 gnd.n4668 0.152939
R11443 gnd.n4670 gnd.n4669 0.152939
R11444 gnd.n4671 gnd.n4670 0.152939
R11445 gnd.n4671 gnd.n1639 0.152939
R11446 gnd.n4707 gnd.n1639 0.152939
R11447 gnd.n4708 gnd.n4707 0.152939
R11448 gnd.n4709 gnd.n4708 0.152939
R11449 gnd.n4709 gnd.n1616 0.152939
R11450 gnd.n4753 gnd.n1616 0.152939
R11451 gnd.n4754 gnd.n4753 0.152939
R11452 gnd.n4755 gnd.n4754 0.152939
R11453 gnd.n4756 gnd.n4755 0.152939
R11454 gnd.n4756 gnd.n1595 0.152939
R11455 gnd.n4808 gnd.n1595 0.152939
R11456 gnd.n4809 gnd.n4808 0.152939
R11457 gnd.n4810 gnd.n4809 0.152939
R11458 gnd.n4811 gnd.n4810 0.152939
R11459 gnd.n4811 gnd.n1568 0.152939
R11460 gnd.n4845 gnd.n1568 0.152939
R11461 gnd.n4846 gnd.n4845 0.152939
R11462 gnd.n4847 gnd.n4846 0.152939
R11463 gnd.n4847 gnd.n1550 0.152939
R11464 gnd.n4871 gnd.n1550 0.152939
R11465 gnd.n4872 gnd.n4871 0.152939
R11466 gnd.n4873 gnd.n4872 0.152939
R11467 gnd.n4874 gnd.n4873 0.152939
R11468 gnd.n4874 gnd.n1522 0.152939
R11469 gnd.n4924 gnd.n1522 0.152939
R11470 gnd.n4925 gnd.n4924 0.152939
R11471 gnd.n4926 gnd.n4925 0.152939
R11472 gnd.n4926 gnd.n1430 0.152939
R11473 gnd.n5067 gnd.n1430 0.152939
R11474 gnd.n5068 gnd.n5067 0.152939
R11475 gnd.n5069 gnd.n5068 0.152939
R11476 gnd.n5070 gnd.n5069 0.152939
R11477 gnd.n5071 gnd.n5070 0.152939
R11478 gnd.n5072 gnd.n5071 0.152939
R11479 gnd.n5112 gnd.n5072 0.152939
R11480 gnd.n5113 gnd.n5112 0.152939
R11481 gnd.n5114 gnd.n5113 0.152939
R11482 gnd.n5114 gnd.n5109 0.152939
R11483 gnd.n5120 gnd.n5109 0.152939
R11484 gnd.n5121 gnd.n5120 0.152939
R11485 gnd.n5122 gnd.n5121 0.152939
R11486 gnd.n5123 gnd.n5122 0.152939
R11487 gnd.n5124 gnd.n5123 0.152939
R11488 gnd.n5127 gnd.n5124 0.152939
R11489 gnd.n5128 gnd.n5127 0.152939
R11490 gnd.n5129 gnd.n5128 0.152939
R11491 gnd.n5130 gnd.n5129 0.152939
R11492 gnd.n5132 gnd.n5130 0.152939
R11493 gnd.n5134 gnd.n5132 0.152939
R11494 gnd.n5134 gnd.n5133 0.152939
R11495 gnd.n5133 gnd.n506 0.152939
R11496 gnd.n507 gnd.n506 0.152939
R11497 gnd.n508 gnd.n507 0.152939
R11498 gnd.n6204 gnd.n508 0.152939
R11499 gnd.n6205 gnd.n6204 0.152939
R11500 gnd.n3703 gnd.n3648 0.152939
R11501 gnd.n3649 gnd.n3648 0.152939
R11502 gnd.n3650 gnd.n3649 0.152939
R11503 gnd.n3651 gnd.n3650 0.152939
R11504 gnd.n3652 gnd.n3651 0.152939
R11505 gnd.n3653 gnd.n3652 0.152939
R11506 gnd.n3654 gnd.n3653 0.152939
R11507 gnd.n3655 gnd.n3654 0.152939
R11508 gnd.n3656 gnd.n3655 0.152939
R11509 gnd.n3657 gnd.n3656 0.152939
R11510 gnd.n3658 gnd.n3657 0.152939
R11511 gnd.n3659 gnd.n3658 0.152939
R11512 gnd.n3660 gnd.n3659 0.152939
R11513 gnd.n3661 gnd.n3660 0.152939
R11514 gnd.n3662 gnd.n3661 0.152939
R11515 gnd.n3663 gnd.n3662 0.152939
R11516 gnd.n3664 gnd.n3663 0.152939
R11517 gnd.n3665 gnd.n3664 0.152939
R11518 gnd.n3666 gnd.n3665 0.152939
R11519 gnd.n3667 gnd.n3666 0.152939
R11520 gnd.n3882 gnd.n2117 0.152939
R11521 gnd.n3609 gnd.n2117 0.152939
R11522 gnd.n3609 gnd.n3608 0.152939
R11523 gnd.n3616 gnd.n3608 0.152939
R11524 gnd.n3617 gnd.n3616 0.152939
R11525 gnd.n3618 gnd.n3617 0.152939
R11526 gnd.n3618 gnd.n3606 0.152939
R11527 gnd.n3626 gnd.n3606 0.152939
R11528 gnd.n3627 gnd.n3626 0.152939
R11529 gnd.n3628 gnd.n3627 0.152939
R11530 gnd.n3628 gnd.n3604 0.152939
R11531 gnd.n3636 gnd.n3604 0.152939
R11532 gnd.n3637 gnd.n3636 0.152939
R11533 gnd.n3638 gnd.n3637 0.152939
R11534 gnd.n3638 gnd.n3602 0.152939
R11535 gnd.n3646 gnd.n3602 0.152939
R11536 gnd.n3647 gnd.n3646 0.152939
R11537 gnd.n3704 gnd.n3647 0.152939
R11538 gnd.n3884 gnd.n3883 0.152939
R11539 gnd.n3884 gnd.n2101 0.152939
R11540 gnd.n3898 gnd.n2101 0.152939
R11541 gnd.n3899 gnd.n3898 0.152939
R11542 gnd.n3900 gnd.n3899 0.152939
R11543 gnd.n3900 gnd.n2085 0.152939
R11544 gnd.n3914 gnd.n2085 0.152939
R11545 gnd.n3915 gnd.n3914 0.152939
R11546 gnd.n3916 gnd.n3915 0.152939
R11547 gnd.n3916 gnd.n2069 0.152939
R11548 gnd.n3930 gnd.n2069 0.152939
R11549 gnd.n3931 gnd.n3930 0.152939
R11550 gnd.n3932 gnd.n3931 0.152939
R11551 gnd.n3932 gnd.n2053 0.152939
R11552 gnd.n3947 gnd.n2053 0.152939
R11553 gnd.n3948 gnd.n3947 0.152939
R11554 gnd.n3949 gnd.n3948 0.152939
R11555 gnd.n3950 gnd.n3949 0.152939
R11556 gnd.n3951 gnd.n3950 0.152939
R11557 gnd.n3951 gnd.n2036 0.152939
R11558 gnd.n3978 gnd.n2036 0.152939
R11559 gnd.n3979 gnd.n3978 0.152939
R11560 gnd.n3980 gnd.n3979 0.152939
R11561 gnd.n3981 gnd.n3980 0.152939
R11562 gnd.n3983 gnd.n3981 0.152939
R11563 gnd.n3983 gnd.n3982 0.152939
R11564 gnd.n3982 gnd.n1016 0.152939
R11565 gnd.n1017 gnd.n1016 0.152939
R11566 gnd.n1018 gnd.n1017 0.152939
R11567 gnd.n1037 gnd.n1018 0.152939
R11568 gnd.n1038 gnd.n1037 0.152939
R11569 gnd.n1039 gnd.n1038 0.152939
R11570 gnd.n1040 gnd.n1039 0.152939
R11571 gnd.n1057 gnd.n1040 0.152939
R11572 gnd.n1058 gnd.n1057 0.152939
R11573 gnd.n1059 gnd.n1058 0.152939
R11574 gnd.n1060 gnd.n1059 0.152939
R11575 gnd.n1079 gnd.n1060 0.152939
R11576 gnd.n1080 gnd.n1079 0.152939
R11577 gnd.n1081 gnd.n1080 0.152939
R11578 gnd.n1082 gnd.n1081 0.152939
R11579 gnd.n1908 gnd.n1082 0.152939
R11580 gnd.n1007 gnd.n1006 0.152939
R11581 gnd.n1026 gnd.n1007 0.152939
R11582 gnd.n1027 gnd.n1026 0.152939
R11583 gnd.n1028 gnd.n1027 0.152939
R11584 gnd.n1029 gnd.n1028 0.152939
R11585 gnd.n1047 gnd.n1029 0.152939
R11586 gnd.n1048 gnd.n1047 0.152939
R11587 gnd.n1049 gnd.n1048 0.152939
R11588 gnd.n1050 gnd.n1049 0.152939
R11589 gnd.n1068 gnd.n1050 0.152939
R11590 gnd.n1069 gnd.n1068 0.152939
R11591 gnd.n1070 gnd.n1069 0.152939
R11592 gnd.n1071 gnd.n1070 0.152939
R11593 gnd.n1090 gnd.n1071 0.152939
R11594 gnd.n1091 gnd.n1090 0.152939
R11595 gnd.n5441 gnd.n1091 0.152939
R11596 gnd.n5440 gnd.n1092 0.152939
R11597 gnd.n1126 gnd.n1092 0.152939
R11598 gnd.n1127 gnd.n1126 0.152939
R11599 gnd.n1128 gnd.n1127 0.152939
R11600 gnd.n1129 gnd.n1128 0.152939
R11601 gnd.n1130 gnd.n1129 0.152939
R11602 gnd.n1131 gnd.n1130 0.152939
R11603 gnd.n1132 gnd.n1131 0.152939
R11604 gnd.n1133 gnd.n1132 0.152939
R11605 gnd.n1134 gnd.n1133 0.152939
R11606 gnd.n1135 gnd.n1134 0.152939
R11607 gnd.n1136 gnd.n1135 0.152939
R11608 gnd.n1137 gnd.n1136 0.152939
R11609 gnd.n1138 gnd.n1137 0.152939
R11610 gnd.n1139 gnd.n1138 0.152939
R11611 gnd.n4096 gnd.n4095 0.152939
R11612 gnd.n4097 gnd.n4096 0.152939
R11613 gnd.n4097 gnd.n4091 0.152939
R11614 gnd.n4105 gnd.n4091 0.152939
R11615 gnd.n4106 gnd.n4105 0.152939
R11616 gnd.n4107 gnd.n4106 0.152939
R11617 gnd.n4107 gnd.n4089 0.152939
R11618 gnd.n4115 gnd.n4089 0.152939
R11619 gnd.n4116 gnd.n4115 0.152939
R11620 gnd.n4117 gnd.n4116 0.152939
R11621 gnd.n4117 gnd.n4087 0.152939
R11622 gnd.n4125 gnd.n4087 0.152939
R11623 gnd.n4126 gnd.n4125 0.152939
R11624 gnd.n4127 gnd.n4126 0.152939
R11625 gnd.n4127 gnd.n4085 0.152939
R11626 gnd.n4135 gnd.n4085 0.152939
R11627 gnd.n4136 gnd.n4135 0.152939
R11628 gnd.n4137 gnd.n4136 0.152939
R11629 gnd.n4137 gnd.n4080 0.152939
R11630 gnd.n4143 gnd.n4080 0.152939
R11631 gnd.n3796 gnd.n3752 0.152939
R11632 gnd.n3796 gnd.n3795 0.152939
R11633 gnd.n3795 gnd.n3794 0.152939
R11634 gnd.n3794 gnd.n3755 0.152939
R11635 gnd.n3756 gnd.n3755 0.152939
R11636 gnd.n3757 gnd.n3756 0.152939
R11637 gnd.n3758 gnd.n3757 0.152939
R11638 gnd.n3759 gnd.n3758 0.152939
R11639 gnd.n3760 gnd.n3759 0.152939
R11640 gnd.n3761 gnd.n3760 0.152939
R11641 gnd.n3762 gnd.n3761 0.152939
R11642 gnd.n3763 gnd.n3762 0.152939
R11643 gnd.n3764 gnd.n3763 0.152939
R11644 gnd.n3765 gnd.n3764 0.152939
R11645 gnd.n3766 gnd.n3765 0.152939
R11646 gnd.n3767 gnd.n3766 0.152939
R11647 gnd.n3768 gnd.n3767 0.152939
R11648 gnd.n3770 gnd.n3768 0.152939
R11649 gnd.n3770 gnd.n3769 0.152939
R11650 gnd.n3769 gnd.n2037 0.152939
R11651 gnd.n3977 gnd.n2037 0.152939
R11652 gnd.n3977 gnd.n2038 0.152939
R11653 gnd.n3968 gnd.n2038 0.152939
R11654 gnd.n3970 gnd.n3968 0.152939
R11655 gnd.n3970 gnd.n3969 0.152939
R11656 gnd.n3969 gnd.n2019 0.152939
R11657 gnd.n2019 gnd.n2017 0.152939
R11658 gnd.n4013 gnd.n2017 0.152939
R11659 gnd.n4014 gnd.n4013 0.152939
R11660 gnd.n4015 gnd.n4014 0.152939
R11661 gnd.n4016 gnd.n4015 0.152939
R11662 gnd.n4017 gnd.n4016 0.152939
R11663 gnd.n4017 gnd.n2001 0.152939
R11664 gnd.n4068 gnd.n2001 0.152939
R11665 gnd.n4069 gnd.n4068 0.152939
R11666 gnd.n4070 gnd.n4069 0.152939
R11667 gnd.n4070 gnd.n1999 0.152939
R11668 gnd.n4076 gnd.n1999 0.152939
R11669 gnd.n4077 gnd.n4076 0.152939
R11670 gnd.n4078 gnd.n4077 0.152939
R11671 gnd.n4079 gnd.n4078 0.152939
R11672 gnd.n4144 gnd.n4079 0.152939
R11673 gnd.n3710 gnd.n3709 0.152939
R11674 gnd.n3711 gnd.n3710 0.152939
R11675 gnd.n3712 gnd.n3711 0.152939
R11676 gnd.n3713 gnd.n3712 0.152939
R11677 gnd.n3714 gnd.n3713 0.152939
R11678 gnd.n3715 gnd.n3714 0.152939
R11679 gnd.n3716 gnd.n3715 0.152939
R11680 gnd.n3717 gnd.n3716 0.152939
R11681 gnd.n3718 gnd.n3717 0.152939
R11682 gnd.n3719 gnd.n3718 0.152939
R11683 gnd.n3720 gnd.n3719 0.152939
R11684 gnd.n3721 gnd.n3720 0.152939
R11685 gnd.n3722 gnd.n3721 0.152939
R11686 gnd.n3723 gnd.n3722 0.152939
R11687 gnd.n3724 gnd.n3723 0.152939
R11688 gnd.n3725 gnd.n3724 0.152939
R11689 gnd.n3726 gnd.n3725 0.152939
R11690 gnd.n3729 gnd.n3726 0.152939
R11691 gnd.n3730 gnd.n3729 0.152939
R11692 gnd.n3731 gnd.n3730 0.152939
R11693 gnd.n3732 gnd.n3731 0.152939
R11694 gnd.n3733 gnd.n3732 0.152939
R11695 gnd.n3734 gnd.n3733 0.152939
R11696 gnd.n3735 gnd.n3734 0.152939
R11697 gnd.n3736 gnd.n3735 0.152939
R11698 gnd.n3737 gnd.n3736 0.152939
R11699 gnd.n3738 gnd.n3737 0.152939
R11700 gnd.n3739 gnd.n3738 0.152939
R11701 gnd.n3740 gnd.n3739 0.152939
R11702 gnd.n3741 gnd.n3740 0.152939
R11703 gnd.n3742 gnd.n3741 0.152939
R11704 gnd.n3743 gnd.n3742 0.152939
R11705 gnd.n3744 gnd.n3743 0.152939
R11706 gnd.n3745 gnd.n3744 0.152939
R11707 gnd.n3746 gnd.n3745 0.152939
R11708 gnd.n3804 gnd.n3746 0.152939
R11709 gnd.n3804 gnd.n3803 0.152939
R11710 gnd.n3803 gnd.n3802 0.152939
R11711 gnd.n3890 gnd.n2109 0.152939
R11712 gnd.n3891 gnd.n3890 0.152939
R11713 gnd.n3892 gnd.n3891 0.152939
R11714 gnd.n3892 gnd.n2092 0.152939
R11715 gnd.n3906 gnd.n2092 0.152939
R11716 gnd.n3907 gnd.n3906 0.152939
R11717 gnd.n3908 gnd.n3907 0.152939
R11718 gnd.n3908 gnd.n2077 0.152939
R11719 gnd.n3922 gnd.n2077 0.152939
R11720 gnd.n3923 gnd.n3922 0.152939
R11721 gnd.n3924 gnd.n3923 0.152939
R11722 gnd.n3924 gnd.n2060 0.152939
R11723 gnd.n3938 gnd.n2060 0.152939
R11724 gnd.n3939 gnd.n3938 0.152939
R11725 gnd.n3940 gnd.n3939 0.152939
R11726 gnd.n3940 gnd.n1006 0.152939
R11727 gnd.n5665 gnd.n829 0.152939
R11728 gnd.n834 gnd.n829 0.152939
R11729 gnd.n835 gnd.n834 0.152939
R11730 gnd.n836 gnd.n835 0.152939
R11731 gnd.n841 gnd.n836 0.152939
R11732 gnd.n842 gnd.n841 0.152939
R11733 gnd.n843 gnd.n842 0.152939
R11734 gnd.n844 gnd.n843 0.152939
R11735 gnd.n849 gnd.n844 0.152939
R11736 gnd.n850 gnd.n849 0.152939
R11737 gnd.n851 gnd.n850 0.152939
R11738 gnd.n852 gnd.n851 0.152939
R11739 gnd.n857 gnd.n852 0.152939
R11740 gnd.n858 gnd.n857 0.152939
R11741 gnd.n859 gnd.n858 0.152939
R11742 gnd.n860 gnd.n859 0.152939
R11743 gnd.n865 gnd.n860 0.152939
R11744 gnd.n866 gnd.n865 0.152939
R11745 gnd.n867 gnd.n866 0.152939
R11746 gnd.n868 gnd.n867 0.152939
R11747 gnd.n873 gnd.n868 0.152939
R11748 gnd.n874 gnd.n873 0.152939
R11749 gnd.n875 gnd.n874 0.152939
R11750 gnd.n876 gnd.n875 0.152939
R11751 gnd.n881 gnd.n876 0.152939
R11752 gnd.n882 gnd.n881 0.152939
R11753 gnd.n883 gnd.n882 0.152939
R11754 gnd.n884 gnd.n883 0.152939
R11755 gnd.n889 gnd.n884 0.152939
R11756 gnd.n890 gnd.n889 0.152939
R11757 gnd.n891 gnd.n890 0.152939
R11758 gnd.n892 gnd.n891 0.152939
R11759 gnd.n897 gnd.n892 0.152939
R11760 gnd.n898 gnd.n897 0.152939
R11761 gnd.n899 gnd.n898 0.152939
R11762 gnd.n900 gnd.n899 0.152939
R11763 gnd.n905 gnd.n900 0.152939
R11764 gnd.n906 gnd.n905 0.152939
R11765 gnd.n907 gnd.n906 0.152939
R11766 gnd.n908 gnd.n907 0.152939
R11767 gnd.n913 gnd.n908 0.152939
R11768 gnd.n914 gnd.n913 0.152939
R11769 gnd.n915 gnd.n914 0.152939
R11770 gnd.n916 gnd.n915 0.152939
R11771 gnd.n921 gnd.n916 0.152939
R11772 gnd.n922 gnd.n921 0.152939
R11773 gnd.n923 gnd.n922 0.152939
R11774 gnd.n924 gnd.n923 0.152939
R11775 gnd.n929 gnd.n924 0.152939
R11776 gnd.n930 gnd.n929 0.152939
R11777 gnd.n931 gnd.n930 0.152939
R11778 gnd.n932 gnd.n931 0.152939
R11779 gnd.n937 gnd.n932 0.152939
R11780 gnd.n938 gnd.n937 0.152939
R11781 gnd.n939 gnd.n938 0.152939
R11782 gnd.n940 gnd.n939 0.152939
R11783 gnd.n945 gnd.n940 0.152939
R11784 gnd.n946 gnd.n945 0.152939
R11785 gnd.n947 gnd.n946 0.152939
R11786 gnd.n948 gnd.n947 0.152939
R11787 gnd.n953 gnd.n948 0.152939
R11788 gnd.n954 gnd.n953 0.152939
R11789 gnd.n955 gnd.n954 0.152939
R11790 gnd.n956 gnd.n955 0.152939
R11791 gnd.n961 gnd.n956 0.152939
R11792 gnd.n962 gnd.n961 0.152939
R11793 gnd.n963 gnd.n962 0.152939
R11794 gnd.n964 gnd.n963 0.152939
R11795 gnd.n969 gnd.n964 0.152939
R11796 gnd.n970 gnd.n969 0.152939
R11797 gnd.n971 gnd.n970 0.152939
R11798 gnd.n972 gnd.n971 0.152939
R11799 gnd.n977 gnd.n972 0.152939
R11800 gnd.n978 gnd.n977 0.152939
R11801 gnd.n979 gnd.n978 0.152939
R11802 gnd.n980 gnd.n979 0.152939
R11803 gnd.n985 gnd.n980 0.152939
R11804 gnd.n986 gnd.n985 0.152939
R11805 gnd.n987 gnd.n986 0.152939
R11806 gnd.n988 gnd.n987 0.152939
R11807 gnd.n993 gnd.n988 0.152939
R11808 gnd.n994 gnd.n993 0.152939
R11809 gnd.n995 gnd.n994 0.152939
R11810 gnd.n996 gnd.n995 0.152939
R11811 gnd.n5156 gnd.n5100 0.152939
R11812 gnd.n5164 gnd.n5100 0.152939
R11813 gnd.n5165 gnd.n5164 0.152939
R11814 gnd.n5166 gnd.n5165 0.152939
R11815 gnd.n5166 gnd.n5096 0.152939
R11816 gnd.n5174 gnd.n5096 0.152939
R11817 gnd.n5175 gnd.n5174 0.152939
R11818 gnd.n5176 gnd.n5175 0.152939
R11819 gnd.n5176 gnd.n1416 0.152939
R11820 gnd.n4230 gnd.n4217 0.152939
R11821 gnd.n4226 gnd.n4217 0.152939
R11822 gnd.n4226 gnd.n4225 0.152939
R11823 gnd.n4225 gnd.n4224 0.152939
R11824 gnd.n4224 gnd.n1829 0.152939
R11825 gnd.n4276 gnd.n1829 0.152939
R11826 gnd.n4277 gnd.n4276 0.152939
R11827 gnd.n4281 gnd.n4277 0.152939
R11828 gnd.n4281 gnd.n4280 0.152939
R11829 gnd.n4280 gnd.n4279 0.152939
R11830 gnd.n4279 gnd.n1330 0.152939
R11831 gnd.n5304 gnd.n1330 0.152939
R11832 gnd.n5304 gnd.n5303 0.152939
R11833 gnd.n5303 gnd.n5302 0.152939
R11834 gnd.n5302 gnd.n1331 0.152939
R11835 gnd.n5298 gnd.n1331 0.152939
R11836 gnd.n5298 gnd.n5297 0.152939
R11837 gnd.n5297 gnd.n5296 0.152939
R11838 gnd.n5296 gnd.n1336 0.152939
R11839 gnd.n5292 gnd.n1336 0.152939
R11840 gnd.n5292 gnd.n5291 0.152939
R11841 gnd.n5291 gnd.n5290 0.152939
R11842 gnd.n5290 gnd.n1341 0.152939
R11843 gnd.n5286 gnd.n1341 0.152939
R11844 gnd.n5286 gnd.n5285 0.152939
R11845 gnd.n5285 gnd.n5284 0.152939
R11846 gnd.n5284 gnd.n1346 0.152939
R11847 gnd.n5280 gnd.n1346 0.152939
R11848 gnd.n5280 gnd.n5279 0.152939
R11849 gnd.n5279 gnd.n5278 0.152939
R11850 gnd.n5278 gnd.n1351 0.152939
R11851 gnd.n5274 gnd.n1351 0.152939
R11852 gnd.n5274 gnd.n5273 0.152939
R11853 gnd.n5273 gnd.n5272 0.152939
R11854 gnd.n5272 gnd.n1356 0.152939
R11855 gnd.n5268 gnd.n1356 0.152939
R11856 gnd.n5268 gnd.n5267 0.152939
R11857 gnd.n5267 gnd.n5266 0.152939
R11858 gnd.n5266 gnd.n1361 0.152939
R11859 gnd.n5262 gnd.n1361 0.152939
R11860 gnd.n5262 gnd.n5261 0.152939
R11861 gnd.n5261 gnd.n5260 0.152939
R11862 gnd.n5260 gnd.n1366 0.152939
R11863 gnd.n5256 gnd.n1366 0.152939
R11864 gnd.n5256 gnd.n5255 0.152939
R11865 gnd.n5255 gnd.n5254 0.152939
R11866 gnd.n5254 gnd.n1371 0.152939
R11867 gnd.n5250 gnd.n1371 0.152939
R11868 gnd.n5250 gnd.n5249 0.152939
R11869 gnd.n5249 gnd.n5248 0.152939
R11870 gnd.n5248 gnd.n1376 0.152939
R11871 gnd.n5244 gnd.n1376 0.152939
R11872 gnd.n5244 gnd.n5243 0.152939
R11873 gnd.n5243 gnd.n5242 0.152939
R11874 gnd.n5242 gnd.n1381 0.152939
R11875 gnd.n5238 gnd.n1381 0.152939
R11876 gnd.n5238 gnd.n5237 0.152939
R11877 gnd.n5237 gnd.n5236 0.152939
R11878 gnd.n5236 gnd.n1386 0.152939
R11879 gnd.n5232 gnd.n1386 0.152939
R11880 gnd.n5232 gnd.n5231 0.152939
R11881 gnd.n5231 gnd.n5230 0.152939
R11882 gnd.n5230 gnd.n1391 0.152939
R11883 gnd.n5226 gnd.n1391 0.152939
R11884 gnd.n5226 gnd.n5225 0.152939
R11885 gnd.n5225 gnd.n5224 0.152939
R11886 gnd.n5224 gnd.n1396 0.152939
R11887 gnd.n5220 gnd.n1396 0.152939
R11888 gnd.n5220 gnd.n5219 0.152939
R11889 gnd.n5219 gnd.n5218 0.152939
R11890 gnd.n5218 gnd.n1401 0.152939
R11891 gnd.n5214 gnd.n1401 0.152939
R11892 gnd.n5214 gnd.n5213 0.152939
R11893 gnd.n5213 gnd.n5212 0.152939
R11894 gnd.n5212 gnd.n1406 0.152939
R11895 gnd.n5208 gnd.n1406 0.152939
R11896 gnd.n5208 gnd.n5207 0.152939
R11897 gnd.n5207 gnd.n5206 0.152939
R11898 gnd.n5206 gnd.n1411 0.152939
R11899 gnd.n5202 gnd.n1411 0.152939
R11900 gnd.n5202 gnd.n5201 0.152939
R11901 gnd.n5201 gnd.n5200 0.152939
R11902 gnd.n4200 gnd.n4199 0.152939
R11903 gnd.n4200 gnd.n1870 0.152939
R11904 gnd.n4206 gnd.n1870 0.152939
R11905 gnd.n4207 gnd.n4206 0.152939
R11906 gnd.n4208 gnd.n4207 0.152939
R11907 gnd.n4208 gnd.n1864 0.152939
R11908 gnd.n4215 gnd.n1864 0.152939
R11909 gnd.n4216 gnd.n4215 0.152939
R11910 gnd.n4231 gnd.n4216 0.152939
R11911 gnd.n3669 gnd.n2021 0.152939
R11912 gnd.n4003 gnd.n2021 0.152939
R11913 gnd.n4004 gnd.n4003 0.152939
R11914 gnd.n4005 gnd.n4004 0.152939
R11915 gnd.n4005 gnd.n2015 0.152939
R11916 gnd.n4027 gnd.n2015 0.152939
R11917 gnd.n4027 gnd.n4026 0.152939
R11918 gnd.n4026 gnd.n4025 0.152939
R11919 gnd.n4025 gnd.n2004 0.152939
R11920 gnd.n4060 gnd.n2004 0.152939
R11921 gnd.n4061 gnd.n4060 0.152939
R11922 gnd.n4062 gnd.n4061 0.152939
R11923 gnd.n4062 gnd.n1995 0.152939
R11924 gnd.n4159 gnd.n1995 0.152939
R11925 gnd.n4159 gnd.n4158 0.152939
R11926 gnd.n4158 gnd.n4157 0.152939
R11927 gnd.n4157 gnd.n1996 0.152939
R11928 gnd.n4153 gnd.n1996 0.152939
R11929 gnd.n4153 gnd.n4152 0.152939
R11930 gnd.n4152 gnd.n1874 0.152939
R11931 gnd.n4255 gnd.n4254 0.152939
R11932 gnd.n4256 gnd.n4255 0.152939
R11933 gnd.n4256 gnd.n1832 0.152939
R11934 gnd.n4262 gnd.n1832 0.152939
R11935 gnd.n4263 gnd.n4262 0.152939
R11936 gnd.n4264 gnd.n4263 0.152939
R11937 gnd.n4264 gnd.n1823 0.152939
R11938 gnd.n4287 gnd.n1823 0.152939
R11939 gnd.n4288 gnd.n4287 0.152939
R11940 gnd.n4289 gnd.n4288 0.152939
R11941 gnd.n4289 gnd.n1821 0.152939
R11942 gnd.n4323 gnd.n1821 0.152939
R11943 gnd.n4324 gnd.n4323 0.152939
R11944 gnd.n4427 gnd.n4324 0.152939
R11945 gnd.n4427 gnd.n4426 0.152939
R11946 gnd.n4426 gnd.n4425 0.152939
R11947 gnd.n4425 gnd.n4325 0.152939
R11948 gnd.n4421 gnd.n4325 0.152939
R11949 gnd.n4421 gnd.n4420 0.152939
R11950 gnd.n4420 gnd.n4419 0.152939
R11951 gnd.n4419 gnd.n4328 0.152939
R11952 gnd.n4415 gnd.n4328 0.152939
R11953 gnd.n4415 gnd.n4414 0.152939
R11954 gnd.n4414 gnd.n4413 0.152939
R11955 gnd.n4413 gnd.n4334 0.152939
R11956 gnd.n4409 gnd.n4334 0.152939
R11957 gnd.n4409 gnd.n4408 0.152939
R11958 gnd.n4408 gnd.n4407 0.152939
R11959 gnd.n4407 gnd.n4337 0.152939
R11960 gnd.n4403 gnd.n4337 0.152939
R11961 gnd.n4403 gnd.n4402 0.152939
R11962 gnd.n4402 gnd.n4401 0.152939
R11963 gnd.n4401 gnd.n4341 0.152939
R11964 gnd.n4397 gnd.n4341 0.152939
R11965 gnd.n4397 gnd.n4396 0.152939
R11966 gnd.n4396 gnd.n4395 0.152939
R11967 gnd.n4395 gnd.n4345 0.152939
R11968 gnd.n4391 gnd.n4345 0.152939
R11969 gnd.n4391 gnd.n4390 0.152939
R11970 gnd.n4390 gnd.n4389 0.152939
R11971 gnd.n4389 gnd.n4349 0.152939
R11972 gnd.n4385 gnd.n4349 0.152939
R11973 gnd.n4385 gnd.n4384 0.152939
R11974 gnd.n4384 gnd.n4383 0.152939
R11975 gnd.n4383 gnd.n4354 0.152939
R11976 gnd.n4379 gnd.n4354 0.152939
R11977 gnd.n4379 gnd.n4378 0.152939
R11978 gnd.n4378 gnd.n4377 0.152939
R11979 gnd.n4377 gnd.n4358 0.152939
R11980 gnd.n4373 gnd.n4358 0.152939
R11981 gnd.n4373 gnd.n4372 0.152939
R11982 gnd.n4372 gnd.n4371 0.152939
R11983 gnd.n4371 gnd.n4361 0.152939
R11984 gnd.n4367 gnd.n4361 0.152939
R11985 gnd.n4367 gnd.n4366 0.152939
R11986 gnd.n4366 gnd.n1608 0.152939
R11987 gnd.n4763 gnd.n1608 0.152939
R11988 gnd.n4764 gnd.n4763 0.152939
R11989 gnd.n4794 gnd.n4764 0.152939
R11990 gnd.n4794 gnd.n4793 0.152939
R11991 gnd.n4793 gnd.n4792 0.152939
R11992 gnd.n4792 gnd.n4765 0.152939
R11993 gnd.n4788 gnd.n4765 0.152939
R11994 gnd.n4788 gnd.n4787 0.152939
R11995 gnd.n4787 gnd.n4786 0.152939
R11996 gnd.n4786 gnd.n4770 0.152939
R11997 gnd.n4782 gnd.n4770 0.152939
R11998 gnd.n4782 gnd.n4781 0.152939
R11999 gnd.n4781 gnd.n4780 0.152939
R12000 gnd.n4780 gnd.n4774 0.152939
R12001 gnd.n4776 gnd.n4774 0.152939
R12002 gnd.n4776 gnd.n1536 0.152939
R12003 gnd.n4909 gnd.n1536 0.152939
R12004 gnd.n4909 gnd.n4908 0.152939
R12005 gnd.n4908 gnd.n4907 0.152939
R12006 gnd.n4907 gnd.n1537 0.152939
R12007 gnd.n4903 gnd.n1537 0.152939
R12008 gnd.n4903 gnd.n4902 0.152939
R12009 gnd.n4902 gnd.n1424 0.152939
R12010 gnd.n5192 gnd.n1424 0.152939
R12011 gnd.n5193 gnd.n5192 0.152939
R12012 gnd.n5194 gnd.n5193 0.152939
R12013 gnd.n6442 gnd.n318 0.152939
R12014 gnd.n6456 gnd.n318 0.152939
R12015 gnd.n6457 gnd.n6456 0.152939
R12016 gnd.n6458 gnd.n6457 0.152939
R12017 gnd.n6458 gnd.n300 0.152939
R12018 gnd.n6472 gnd.n300 0.152939
R12019 gnd.n6473 gnd.n6472 0.152939
R12020 gnd.n6474 gnd.n6473 0.152939
R12021 gnd.n6474 gnd.n282 0.152939
R12022 gnd.n6488 gnd.n282 0.152939
R12023 gnd.n6489 gnd.n6488 0.152939
R12024 gnd.n6490 gnd.n6489 0.152939
R12025 gnd.n6490 gnd.n265 0.152939
R12026 gnd.n6505 gnd.n265 0.152939
R12027 gnd.n6506 gnd.n6505 0.152939
R12028 gnd.n6511 gnd.n6506 0.152939
R12029 gnd.n6511 gnd.n6510 0.152939
R12030 gnd.n6510 gnd.n6509 0.152939
R12031 gnd.n6509 gnd.n240 0.152939
R12032 gnd.n6535 gnd.n240 0.152939
R12033 gnd.n6536 gnd.n6535 0.152939
R12034 gnd.n6537 gnd.n6536 0.152939
R12035 gnd.n6537 gnd.n227 0.152939
R12036 gnd.n6549 gnd.n227 0.152939
R12037 gnd.n6550 gnd.n6549 0.152939
R12038 gnd.n6551 gnd.n6550 0.152939
R12039 gnd.n6551 gnd.n206 0.152939
R12040 gnd.n6565 gnd.n206 0.152939
R12041 gnd.n6566 gnd.n6565 0.152939
R12042 gnd.n6567 gnd.n6566 0.152939
R12043 gnd.n6567 gnd.n191 0.152939
R12044 gnd.n6581 gnd.n191 0.152939
R12045 gnd.n6582 gnd.n6581 0.152939
R12046 gnd.n6583 gnd.n6582 0.152939
R12047 gnd.n6583 gnd.n175 0.152939
R12048 gnd.n6597 gnd.n175 0.152939
R12049 gnd.n6598 gnd.n6597 0.152939
R12050 gnd.n6673 gnd.n6598 0.152939
R12051 gnd.n6673 gnd.n6672 0.152939
R12052 gnd.n6672 gnd.n6671 0.152939
R12053 gnd.n6671 gnd.n6599 0.152939
R12054 gnd.n6667 gnd.n6599 0.152939
R12055 gnd.n6666 gnd.n6601 0.152939
R12056 gnd.n6662 gnd.n6601 0.152939
R12057 gnd.n6662 gnd.n6661 0.152939
R12058 gnd.n6661 gnd.n6660 0.152939
R12059 gnd.n6660 gnd.n6607 0.152939
R12060 gnd.n6656 gnd.n6607 0.152939
R12061 gnd.n6656 gnd.n6655 0.152939
R12062 gnd.n6655 gnd.n6654 0.152939
R12063 gnd.n6654 gnd.n6615 0.152939
R12064 gnd.n6650 gnd.n6615 0.152939
R12065 gnd.n6650 gnd.n6649 0.152939
R12066 gnd.n6649 gnd.n6648 0.152939
R12067 gnd.n6648 gnd.n6623 0.152939
R12068 gnd.n6644 gnd.n6623 0.152939
R12069 gnd.n6644 gnd.n6643 0.152939
R12070 gnd.n6643 gnd.n6642 0.152939
R12071 gnd.n6642 gnd.n6631 0.152939
R12072 gnd.n6631 gnd.n78 0.152939
R12073 gnd.n5154 gnd.n5105 0.152939
R12074 gnd.n5105 gnd.n470 0.152939
R12075 gnd.n6307 gnd.n470 0.152939
R12076 gnd.n6307 gnd.n6306 0.152939
R12077 gnd.n6306 gnd.n6305 0.152939
R12078 gnd.n6305 gnd.n471 0.152939
R12079 gnd.n6301 gnd.n471 0.152939
R12080 gnd.n6301 gnd.n6300 0.152939
R12081 gnd.n6300 gnd.n6299 0.152939
R12082 gnd.n6299 gnd.n475 0.152939
R12083 gnd.n6295 gnd.n475 0.152939
R12084 gnd.n6295 gnd.n6294 0.152939
R12085 gnd.n6294 gnd.n6293 0.152939
R12086 gnd.n6293 gnd.n479 0.152939
R12087 gnd.n6289 gnd.n479 0.152939
R12088 gnd.n6289 gnd.n252 0.152939
R12089 gnd.n6522 gnd.n252 0.152939
R12090 gnd.n6523 gnd.n6522 0.152939
R12091 gnd.n6524 gnd.n6523 0.152939
R12092 gnd.n6524 gnd.n51 0.152939
R12093 gnd.n6798 gnd.n51 0.152939
R12094 gnd.n6798 gnd.n6797 0.152939
R12095 gnd.n6797 gnd.n53 0.152939
R12096 gnd.n6793 gnd.n53 0.152939
R12097 gnd.n6793 gnd.n6792 0.152939
R12098 gnd.n6792 gnd.n6791 0.152939
R12099 gnd.n6791 gnd.n58 0.152939
R12100 gnd.n6787 gnd.n58 0.152939
R12101 gnd.n6787 gnd.n6786 0.152939
R12102 gnd.n6786 gnd.n6785 0.152939
R12103 gnd.n6785 gnd.n63 0.152939
R12104 gnd.n6781 gnd.n63 0.152939
R12105 gnd.n6781 gnd.n6780 0.152939
R12106 gnd.n6780 gnd.n6779 0.152939
R12107 gnd.n6779 gnd.n68 0.152939
R12108 gnd.n6775 gnd.n68 0.152939
R12109 gnd.n6775 gnd.n6774 0.152939
R12110 gnd.n6774 gnd.n6773 0.152939
R12111 gnd.n6773 gnd.n73 0.152939
R12112 gnd.n6769 gnd.n73 0.152939
R12113 gnd.n6769 gnd.n6768 0.152939
R12114 gnd.n6768 gnd.n6767 0.152939
R12115 gnd.n5156 gnd.n5155 0.151415
R12116 gnd.n4199 gnd.n4198 0.151415
R12117 gnd.n3670 gnd.n3667 0.145814
R12118 gnd.n3670 gnd.n3669 0.145814
R12119 gnd.n6206 gnd.n213 0.136171
R12120 gnd.n4035 gnd.n4034 0.136171
R12121 gnd.n2387 gnd.n0 0.127478
R12122 gnd.n2967 gnd.n2966 0.0767195
R12123 gnd.n2966 gnd.n2965 0.0767195
R12124 gnd.n1909 gnd.n1836 0.063
R12125 gnd.n6441 gnd.n333 0.063
R12126 gnd.n3534 gnd.n2161 0.0477147
R12127 gnd.n2730 gnd.n2618 0.0442063
R12128 gnd.n2731 gnd.n2730 0.0442063
R12129 gnd.n2732 gnd.n2731 0.0442063
R12130 gnd.n2732 gnd.n2607 0.0442063
R12131 gnd.n2746 gnd.n2607 0.0442063
R12132 gnd.n2747 gnd.n2746 0.0442063
R12133 gnd.n2748 gnd.n2747 0.0442063
R12134 gnd.n2748 gnd.n2594 0.0442063
R12135 gnd.n2792 gnd.n2594 0.0442063
R12136 gnd.n2793 gnd.n2792 0.0442063
R12137 gnd.n2795 gnd.n2528 0.0344674
R12138 gnd.n5104 gnd.n382 0.0344674
R12139 gnd.n4197 gnd.n1875 0.0344674
R12140 gnd.n2815 gnd.n2814 0.0269946
R12141 gnd.n2817 gnd.n2816 0.0269946
R12142 gnd.n2523 gnd.n2521 0.0269946
R12143 gnd.n2827 gnd.n2825 0.0269946
R12144 gnd.n2826 gnd.n2502 0.0269946
R12145 gnd.n2846 gnd.n2845 0.0269946
R12146 gnd.n2848 gnd.n2847 0.0269946
R12147 gnd.n2497 gnd.n2496 0.0269946
R12148 gnd.n2858 gnd.n2492 0.0269946
R12149 gnd.n2857 gnd.n2494 0.0269946
R12150 gnd.n2493 gnd.n2475 0.0269946
R12151 gnd.n2878 gnd.n2476 0.0269946
R12152 gnd.n2877 gnd.n2477 0.0269946
R12153 gnd.n2911 gnd.n2452 0.0269946
R12154 gnd.n2913 gnd.n2912 0.0269946
R12155 gnd.n2914 gnd.n2399 0.0269946
R12156 gnd.n2447 gnd.n2400 0.0269946
R12157 gnd.n2449 gnd.n2401 0.0269946
R12158 gnd.n2924 gnd.n2923 0.0269946
R12159 gnd.n2926 gnd.n2925 0.0269946
R12160 gnd.n2927 gnd.n2421 0.0269946
R12161 gnd.n2929 gnd.n2422 0.0269946
R12162 gnd.n2932 gnd.n2423 0.0269946
R12163 gnd.n2935 gnd.n2934 0.0269946
R12164 gnd.n2937 gnd.n2936 0.0269946
R12165 gnd.n3002 gnd.n2334 0.0269946
R12166 gnd.n3004 gnd.n3003 0.0269946
R12167 gnd.n3013 gnd.n2327 0.0269946
R12168 gnd.n3015 gnd.n3014 0.0269946
R12169 gnd.n3016 gnd.n2325 0.0269946
R12170 gnd.n3023 gnd.n3019 0.0269946
R12171 gnd.n3022 gnd.n3021 0.0269946
R12172 gnd.n3020 gnd.n2304 0.0269946
R12173 gnd.n3045 gnd.n2305 0.0269946
R12174 gnd.n3044 gnd.n2306 0.0269946
R12175 gnd.n3087 gnd.n2279 0.0269946
R12176 gnd.n3089 gnd.n3088 0.0269946
R12177 gnd.n3098 gnd.n2272 0.0269946
R12178 gnd.n3100 gnd.n3099 0.0269946
R12179 gnd.n3101 gnd.n2270 0.0269946
R12180 gnd.n3108 gnd.n3104 0.0269946
R12181 gnd.n3107 gnd.n3106 0.0269946
R12182 gnd.n3105 gnd.n2249 0.0269946
R12183 gnd.n3130 gnd.n2250 0.0269946
R12184 gnd.n3129 gnd.n2251 0.0269946
R12185 gnd.n3176 gnd.n2225 0.0269946
R12186 gnd.n3178 gnd.n3177 0.0269946
R12187 gnd.n3188 gnd.n2218 0.0269946
R12188 gnd.n3447 gnd.n2216 0.0269946
R12189 gnd.n3452 gnd.n3450 0.0269946
R12190 gnd.n3451 gnd.n2197 0.0269946
R12191 gnd.n3476 gnd.n3475 0.0269946
R12192 gnd.n6438 gnd.n333 0.0246168
R12193 gnd.n1912 gnd.n1836 0.0246168
R12194 gnd.n2795 gnd.n2794 0.0202011
R12195 gnd.n6438 gnd.n6437 0.0174837
R12196 gnd.n6437 gnd.n336 0.0174837
R12197 gnd.n6434 gnd.n336 0.0174837
R12198 gnd.n6434 gnd.n6433 0.0174837
R12199 gnd.n6433 gnd.n340 0.0174837
R12200 gnd.n6430 gnd.n340 0.0174837
R12201 gnd.n6430 gnd.n6429 0.0174837
R12202 gnd.n6429 gnd.n344 0.0174837
R12203 gnd.n6426 gnd.n344 0.0174837
R12204 gnd.n6426 gnd.n6425 0.0174837
R12205 gnd.n6425 gnd.n348 0.0174837
R12206 gnd.n6422 gnd.n348 0.0174837
R12207 gnd.n6422 gnd.n6421 0.0174837
R12208 gnd.n6421 gnd.n352 0.0174837
R12209 gnd.n6418 gnd.n352 0.0174837
R12210 gnd.n6418 gnd.n6417 0.0174837
R12211 gnd.n6417 gnd.n356 0.0174837
R12212 gnd.n6414 gnd.n356 0.0174837
R12213 gnd.n6414 gnd.n6413 0.0174837
R12214 gnd.n6413 gnd.n360 0.0174837
R12215 gnd.n6410 gnd.n360 0.0174837
R12216 gnd.n6410 gnd.n6409 0.0174837
R12217 gnd.n6409 gnd.n364 0.0174837
R12218 gnd.n6406 gnd.n364 0.0174837
R12219 gnd.n6406 gnd.n6405 0.0174837
R12220 gnd.n6405 gnd.n368 0.0174837
R12221 gnd.n6402 gnd.n368 0.0174837
R12222 gnd.n6402 gnd.n6401 0.0174837
R12223 gnd.n6401 gnd.n372 0.0174837
R12224 gnd.n6398 gnd.n372 0.0174837
R12225 gnd.n6398 gnd.n6397 0.0174837
R12226 gnd.n6397 gnd.n378 0.0174837
R12227 gnd.n6394 gnd.n378 0.0174837
R12228 gnd.n6394 gnd.n6393 0.0174837
R12229 gnd.n6393 gnd.n382 0.0174837
R12230 gnd.n1912 gnd.n1907 0.0174837
R12231 gnd.n1917 gnd.n1907 0.0174837
R12232 gnd.n1918 gnd.n1917 0.0174837
R12233 gnd.n1918 gnd.n1905 0.0174837
R12234 gnd.n1923 gnd.n1905 0.0174837
R12235 gnd.n1924 gnd.n1923 0.0174837
R12236 gnd.n1924 gnd.n1903 0.0174837
R12237 gnd.n1929 gnd.n1903 0.0174837
R12238 gnd.n1930 gnd.n1929 0.0174837
R12239 gnd.n1930 gnd.n1899 0.0174837
R12240 gnd.n1935 gnd.n1899 0.0174837
R12241 gnd.n1936 gnd.n1935 0.0174837
R12242 gnd.n1936 gnd.n1895 0.0174837
R12243 gnd.n1941 gnd.n1895 0.0174837
R12244 gnd.n1942 gnd.n1941 0.0174837
R12245 gnd.n1942 gnd.n1893 0.0174837
R12246 gnd.n1947 gnd.n1893 0.0174837
R12247 gnd.n1948 gnd.n1947 0.0174837
R12248 gnd.n1948 gnd.n1891 0.0174837
R12249 gnd.n1953 gnd.n1891 0.0174837
R12250 gnd.n1954 gnd.n1953 0.0174837
R12251 gnd.n1954 gnd.n1887 0.0174837
R12252 gnd.n1959 gnd.n1887 0.0174837
R12253 gnd.n1960 gnd.n1959 0.0174837
R12254 gnd.n1960 gnd.n1883 0.0174837
R12255 gnd.n1965 gnd.n1883 0.0174837
R12256 gnd.n1966 gnd.n1965 0.0174837
R12257 gnd.n1966 gnd.n1881 0.0174837
R12258 gnd.n1971 gnd.n1881 0.0174837
R12259 gnd.n1973 gnd.n1971 0.0174837
R12260 gnd.n1973 gnd.n1972 0.0174837
R12261 gnd.n1972 gnd.n1879 0.0174837
R12262 gnd.n4191 gnd.n1879 0.0174837
R12263 gnd.n4191 gnd.n4190 0.0174837
R12264 gnd.n4190 gnd.n1875 0.0174837
R12265 gnd.n2794 gnd.n2793 0.0148637
R12266 gnd.n3445 gnd.n3189 0.0144266
R12267 gnd.n3446 gnd.n3445 0.0130679
R12268 gnd.n2814 gnd.n2528 0.00797283
R12269 gnd.n2816 gnd.n2815 0.00797283
R12270 gnd.n2817 gnd.n2523 0.00797283
R12271 gnd.n2825 gnd.n2521 0.00797283
R12272 gnd.n2827 gnd.n2826 0.00797283
R12273 gnd.n2845 gnd.n2502 0.00797283
R12274 gnd.n2847 gnd.n2846 0.00797283
R12275 gnd.n2848 gnd.n2497 0.00797283
R12276 gnd.n2496 gnd.n2492 0.00797283
R12277 gnd.n2858 gnd.n2857 0.00797283
R12278 gnd.n2494 gnd.n2493 0.00797283
R12279 gnd.n2476 gnd.n2475 0.00797283
R12280 gnd.n2878 gnd.n2877 0.00797283
R12281 gnd.n2477 gnd.n2452 0.00797283
R12282 gnd.n2912 gnd.n2911 0.00797283
R12283 gnd.n2914 gnd.n2913 0.00797283
R12284 gnd.n2447 gnd.n2399 0.00797283
R12285 gnd.n2449 gnd.n2400 0.00797283
R12286 gnd.n2923 gnd.n2401 0.00797283
R12287 gnd.n2925 gnd.n2924 0.00797283
R12288 gnd.n2927 gnd.n2926 0.00797283
R12289 gnd.n2929 gnd.n2421 0.00797283
R12290 gnd.n2932 gnd.n2422 0.00797283
R12291 gnd.n2934 gnd.n2423 0.00797283
R12292 gnd.n2937 gnd.n2935 0.00797283
R12293 gnd.n2936 gnd.n2334 0.00797283
R12294 gnd.n3004 gnd.n3002 0.00797283
R12295 gnd.n3003 gnd.n2327 0.00797283
R12296 gnd.n3014 gnd.n3013 0.00797283
R12297 gnd.n3016 gnd.n3015 0.00797283
R12298 gnd.n3019 gnd.n2325 0.00797283
R12299 gnd.n3023 gnd.n3022 0.00797283
R12300 gnd.n3021 gnd.n3020 0.00797283
R12301 gnd.n2305 gnd.n2304 0.00797283
R12302 gnd.n3045 gnd.n3044 0.00797283
R12303 gnd.n2306 gnd.n2279 0.00797283
R12304 gnd.n3089 gnd.n3087 0.00797283
R12305 gnd.n3088 gnd.n2272 0.00797283
R12306 gnd.n3099 gnd.n3098 0.00797283
R12307 gnd.n3101 gnd.n3100 0.00797283
R12308 gnd.n3104 gnd.n2270 0.00797283
R12309 gnd.n3108 gnd.n3107 0.00797283
R12310 gnd.n3106 gnd.n3105 0.00797283
R12311 gnd.n2250 gnd.n2249 0.00797283
R12312 gnd.n3130 gnd.n3129 0.00797283
R12313 gnd.n2251 gnd.n2225 0.00797283
R12314 gnd.n3178 gnd.n3176 0.00797283
R12315 gnd.n3177 gnd.n2218 0.00797283
R12316 gnd.n3189 gnd.n3188 0.00797283
R12317 gnd.n3447 gnd.n3446 0.00797283
R12318 gnd.n3450 gnd.n2216 0.00797283
R12319 gnd.n3452 gnd.n3451 0.00797283
R12320 gnd.n3475 gnd.n2197 0.00797283
R12321 gnd.n3476 gnd.n2161 0.00797283
R12322 gnd.n6536 gnd.n239 0.00614909
R12323 gnd.n3978 gnd.n3977 0.00614909
R12324 gnd.n5155 gnd.n5104 0.000839674
R12325 gnd.n4198 gnd.n4197 0.000839674
R12326 commonsourceibias.n25 commonsourceibias.t46 230.006
R12327 commonsourceibias.n91 commonsourceibias.t62 230.006
R12328 commonsourceibias.n154 commonsourceibias.t54 230.006
R12329 commonsourceibias.n258 commonsourceibias.t16 230.006
R12330 commonsourceibias.n217 commonsourceibias.t75 230.006
R12331 commonsourceibias.n355 commonsourceibias.t65 230.006
R12332 commonsourceibias.n70 commonsourceibias.t32 207.983
R12333 commonsourceibias.n136 commonsourceibias.t71 207.983
R12334 commonsourceibias.n199 commonsourceibias.t61 207.983
R12335 commonsourceibias.n304 commonsourceibias.t2 207.983
R12336 commonsourceibias.n338 commonsourceibias.t84 207.983
R12337 commonsourceibias.n401 commonsourceibias.t73 207.983
R12338 commonsourceibias.n10 commonsourceibias.t14 168.701
R12339 commonsourceibias.n63 commonsourceibias.t24 168.701
R12340 commonsourceibias.n57 commonsourceibias.t30 168.701
R12341 commonsourceibias.n16 commonsourceibias.t20 168.701
R12342 commonsourceibias.n49 commonsourceibias.t36 168.701
R12343 commonsourceibias.n43 commonsourceibias.t44 168.701
R12344 commonsourceibias.n19 commonsourceibias.t26 168.701
R12345 commonsourceibias.n21 commonsourceibias.t34 168.701
R12346 commonsourceibias.n23 commonsourceibias.t10 168.701
R12347 commonsourceibias.n26 commonsourceibias.t40 168.701
R12348 commonsourceibias.n1 commonsourceibias.t81 168.701
R12349 commonsourceibias.n129 commonsourceibias.t55 168.701
R12350 commonsourceibias.n123 commonsourceibias.t53 168.701
R12351 commonsourceibias.n7 commonsourceibias.t76 168.701
R12352 commonsourceibias.n115 commonsourceibias.t86 168.701
R12353 commonsourceibias.n109 commonsourceibias.t50 168.701
R12354 commonsourceibias.n85 commonsourceibias.t69 168.701
R12355 commonsourceibias.n87 commonsourceibias.t67 168.701
R12356 commonsourceibias.n89 commonsourceibias.t78 168.701
R12357 commonsourceibias.n92 commonsourceibias.t64 168.701
R12358 commonsourceibias.n155 commonsourceibias.t57 168.701
R12359 commonsourceibias.n152 commonsourceibias.t68 168.701
R12360 commonsourceibias.n150 commonsourceibias.t58 168.701
R12361 commonsourceibias.n148 commonsourceibias.t60 168.701
R12362 commonsourceibias.n172 commonsourceibias.t91 168.701
R12363 commonsourceibias.n178 commonsourceibias.t77 168.701
R12364 commonsourceibias.n145 commonsourceibias.t66 168.701
R12365 commonsourceibias.n186 commonsourceibias.t95 168.701
R12366 commonsourceibias.n192 commonsourceibias.t49 168.701
R12367 commonsourceibias.n139 commonsourceibias.t72 168.701
R12368 commonsourceibias.n259 commonsourceibias.t8 168.701
R12369 commonsourceibias.n256 commonsourceibias.t18 168.701
R12370 commonsourceibias.n254 commonsourceibias.t4 168.701
R12371 commonsourceibias.n252 commonsourceibias.t42 168.701
R12372 commonsourceibias.n276 commonsourceibias.t12 168.701
R12373 commonsourceibias.n282 commonsourceibias.t6 168.701
R12374 commonsourceibias.n284 commonsourceibias.t28 168.701
R12375 commonsourceibias.n291 commonsourceibias.t0 168.701
R12376 commonsourceibias.n297 commonsourceibias.t38 168.701
R12377 commonsourceibias.n244 commonsourceibias.t22 168.701
R12378 commonsourceibias.n203 commonsourceibias.t92 168.701
R12379 commonsourceibias.n331 commonsourceibias.t51 168.701
R12380 commonsourceibias.n325 commonsourceibias.t63 168.701
R12381 commonsourceibias.n318 commonsourceibias.t88 168.701
R12382 commonsourceibias.n316 commonsourceibias.t48 168.701
R12383 commonsourceibias.n218 commonsourceibias.t59 168.701
R12384 commonsourceibias.n215 commonsourceibias.t90 168.701
R12385 commonsourceibias.n213 commonsourceibias.t80 168.701
R12386 commonsourceibias.n211 commonsourceibias.t83 168.701
R12387 commonsourceibias.n235 commonsourceibias.t94 168.701
R12388 commonsourceibias.n356 commonsourceibias.t52 168.701
R12389 commonsourceibias.n353 commonsourceibias.t82 168.701
R12390 commonsourceibias.n351 commonsourceibias.t70 168.701
R12391 commonsourceibias.n349 commonsourceibias.t74 168.701
R12392 commonsourceibias.n373 commonsourceibias.t87 168.701
R12393 commonsourceibias.n379 commonsourceibias.t89 168.701
R12394 commonsourceibias.n381 commonsourceibias.t79 168.701
R12395 commonsourceibias.n388 commonsourceibias.t56 168.701
R12396 commonsourceibias.n394 commonsourceibias.t93 168.701
R12397 commonsourceibias.n341 commonsourceibias.t85 168.701
R12398 commonsourceibias.n27 commonsourceibias.n24 161.3
R12399 commonsourceibias.n29 commonsourceibias.n28 161.3
R12400 commonsourceibias.n31 commonsourceibias.n30 161.3
R12401 commonsourceibias.n32 commonsourceibias.n22 161.3
R12402 commonsourceibias.n34 commonsourceibias.n33 161.3
R12403 commonsourceibias.n36 commonsourceibias.n35 161.3
R12404 commonsourceibias.n37 commonsourceibias.n20 161.3
R12405 commonsourceibias.n39 commonsourceibias.n38 161.3
R12406 commonsourceibias.n41 commonsourceibias.n40 161.3
R12407 commonsourceibias.n42 commonsourceibias.n18 161.3
R12408 commonsourceibias.n45 commonsourceibias.n44 161.3
R12409 commonsourceibias.n46 commonsourceibias.n17 161.3
R12410 commonsourceibias.n48 commonsourceibias.n47 161.3
R12411 commonsourceibias.n50 commonsourceibias.n15 161.3
R12412 commonsourceibias.n52 commonsourceibias.n51 161.3
R12413 commonsourceibias.n53 commonsourceibias.n14 161.3
R12414 commonsourceibias.n55 commonsourceibias.n54 161.3
R12415 commonsourceibias.n56 commonsourceibias.n13 161.3
R12416 commonsourceibias.n59 commonsourceibias.n58 161.3
R12417 commonsourceibias.n60 commonsourceibias.n12 161.3
R12418 commonsourceibias.n62 commonsourceibias.n61 161.3
R12419 commonsourceibias.n64 commonsourceibias.n11 161.3
R12420 commonsourceibias.n66 commonsourceibias.n65 161.3
R12421 commonsourceibias.n68 commonsourceibias.n67 161.3
R12422 commonsourceibias.n69 commonsourceibias.n9 161.3
R12423 commonsourceibias.n93 commonsourceibias.n90 161.3
R12424 commonsourceibias.n95 commonsourceibias.n94 161.3
R12425 commonsourceibias.n97 commonsourceibias.n96 161.3
R12426 commonsourceibias.n98 commonsourceibias.n88 161.3
R12427 commonsourceibias.n100 commonsourceibias.n99 161.3
R12428 commonsourceibias.n102 commonsourceibias.n101 161.3
R12429 commonsourceibias.n103 commonsourceibias.n86 161.3
R12430 commonsourceibias.n105 commonsourceibias.n104 161.3
R12431 commonsourceibias.n107 commonsourceibias.n106 161.3
R12432 commonsourceibias.n108 commonsourceibias.n84 161.3
R12433 commonsourceibias.n111 commonsourceibias.n110 161.3
R12434 commonsourceibias.n112 commonsourceibias.n8 161.3
R12435 commonsourceibias.n114 commonsourceibias.n113 161.3
R12436 commonsourceibias.n116 commonsourceibias.n6 161.3
R12437 commonsourceibias.n118 commonsourceibias.n117 161.3
R12438 commonsourceibias.n119 commonsourceibias.n5 161.3
R12439 commonsourceibias.n121 commonsourceibias.n120 161.3
R12440 commonsourceibias.n122 commonsourceibias.n4 161.3
R12441 commonsourceibias.n125 commonsourceibias.n124 161.3
R12442 commonsourceibias.n126 commonsourceibias.n3 161.3
R12443 commonsourceibias.n128 commonsourceibias.n127 161.3
R12444 commonsourceibias.n130 commonsourceibias.n2 161.3
R12445 commonsourceibias.n132 commonsourceibias.n131 161.3
R12446 commonsourceibias.n134 commonsourceibias.n133 161.3
R12447 commonsourceibias.n135 commonsourceibias.n0 161.3
R12448 commonsourceibias.n198 commonsourceibias.n138 161.3
R12449 commonsourceibias.n197 commonsourceibias.n196 161.3
R12450 commonsourceibias.n195 commonsourceibias.n194 161.3
R12451 commonsourceibias.n193 commonsourceibias.n140 161.3
R12452 commonsourceibias.n191 commonsourceibias.n190 161.3
R12453 commonsourceibias.n189 commonsourceibias.n141 161.3
R12454 commonsourceibias.n188 commonsourceibias.n187 161.3
R12455 commonsourceibias.n185 commonsourceibias.n142 161.3
R12456 commonsourceibias.n184 commonsourceibias.n183 161.3
R12457 commonsourceibias.n182 commonsourceibias.n143 161.3
R12458 commonsourceibias.n181 commonsourceibias.n180 161.3
R12459 commonsourceibias.n179 commonsourceibias.n144 161.3
R12460 commonsourceibias.n177 commonsourceibias.n176 161.3
R12461 commonsourceibias.n175 commonsourceibias.n146 161.3
R12462 commonsourceibias.n174 commonsourceibias.n173 161.3
R12463 commonsourceibias.n171 commonsourceibias.n147 161.3
R12464 commonsourceibias.n170 commonsourceibias.n169 161.3
R12465 commonsourceibias.n168 commonsourceibias.n167 161.3
R12466 commonsourceibias.n166 commonsourceibias.n149 161.3
R12467 commonsourceibias.n165 commonsourceibias.n164 161.3
R12468 commonsourceibias.n163 commonsourceibias.n162 161.3
R12469 commonsourceibias.n161 commonsourceibias.n151 161.3
R12470 commonsourceibias.n160 commonsourceibias.n159 161.3
R12471 commonsourceibias.n158 commonsourceibias.n157 161.3
R12472 commonsourceibias.n156 commonsourceibias.n153 161.3
R12473 commonsourceibias.n303 commonsourceibias.n243 161.3
R12474 commonsourceibias.n302 commonsourceibias.n301 161.3
R12475 commonsourceibias.n300 commonsourceibias.n299 161.3
R12476 commonsourceibias.n298 commonsourceibias.n245 161.3
R12477 commonsourceibias.n296 commonsourceibias.n295 161.3
R12478 commonsourceibias.n294 commonsourceibias.n246 161.3
R12479 commonsourceibias.n293 commonsourceibias.n292 161.3
R12480 commonsourceibias.n290 commonsourceibias.n247 161.3
R12481 commonsourceibias.n289 commonsourceibias.n288 161.3
R12482 commonsourceibias.n287 commonsourceibias.n248 161.3
R12483 commonsourceibias.n286 commonsourceibias.n285 161.3
R12484 commonsourceibias.n283 commonsourceibias.n249 161.3
R12485 commonsourceibias.n281 commonsourceibias.n280 161.3
R12486 commonsourceibias.n279 commonsourceibias.n250 161.3
R12487 commonsourceibias.n278 commonsourceibias.n277 161.3
R12488 commonsourceibias.n275 commonsourceibias.n251 161.3
R12489 commonsourceibias.n274 commonsourceibias.n273 161.3
R12490 commonsourceibias.n272 commonsourceibias.n271 161.3
R12491 commonsourceibias.n270 commonsourceibias.n253 161.3
R12492 commonsourceibias.n269 commonsourceibias.n268 161.3
R12493 commonsourceibias.n267 commonsourceibias.n266 161.3
R12494 commonsourceibias.n265 commonsourceibias.n255 161.3
R12495 commonsourceibias.n264 commonsourceibias.n263 161.3
R12496 commonsourceibias.n262 commonsourceibias.n261 161.3
R12497 commonsourceibias.n260 commonsourceibias.n257 161.3
R12498 commonsourceibias.n237 commonsourceibias.n236 161.3
R12499 commonsourceibias.n234 commonsourceibias.n210 161.3
R12500 commonsourceibias.n233 commonsourceibias.n232 161.3
R12501 commonsourceibias.n231 commonsourceibias.n230 161.3
R12502 commonsourceibias.n229 commonsourceibias.n212 161.3
R12503 commonsourceibias.n228 commonsourceibias.n227 161.3
R12504 commonsourceibias.n226 commonsourceibias.n225 161.3
R12505 commonsourceibias.n224 commonsourceibias.n214 161.3
R12506 commonsourceibias.n223 commonsourceibias.n222 161.3
R12507 commonsourceibias.n221 commonsourceibias.n220 161.3
R12508 commonsourceibias.n219 commonsourceibias.n216 161.3
R12509 commonsourceibias.n313 commonsourceibias.n209 161.3
R12510 commonsourceibias.n337 commonsourceibias.n202 161.3
R12511 commonsourceibias.n336 commonsourceibias.n335 161.3
R12512 commonsourceibias.n334 commonsourceibias.n333 161.3
R12513 commonsourceibias.n332 commonsourceibias.n204 161.3
R12514 commonsourceibias.n330 commonsourceibias.n329 161.3
R12515 commonsourceibias.n328 commonsourceibias.n205 161.3
R12516 commonsourceibias.n327 commonsourceibias.n326 161.3
R12517 commonsourceibias.n324 commonsourceibias.n206 161.3
R12518 commonsourceibias.n323 commonsourceibias.n322 161.3
R12519 commonsourceibias.n321 commonsourceibias.n207 161.3
R12520 commonsourceibias.n320 commonsourceibias.n319 161.3
R12521 commonsourceibias.n317 commonsourceibias.n208 161.3
R12522 commonsourceibias.n315 commonsourceibias.n314 161.3
R12523 commonsourceibias.n400 commonsourceibias.n340 161.3
R12524 commonsourceibias.n399 commonsourceibias.n398 161.3
R12525 commonsourceibias.n397 commonsourceibias.n396 161.3
R12526 commonsourceibias.n395 commonsourceibias.n342 161.3
R12527 commonsourceibias.n393 commonsourceibias.n392 161.3
R12528 commonsourceibias.n391 commonsourceibias.n343 161.3
R12529 commonsourceibias.n390 commonsourceibias.n389 161.3
R12530 commonsourceibias.n387 commonsourceibias.n344 161.3
R12531 commonsourceibias.n386 commonsourceibias.n385 161.3
R12532 commonsourceibias.n384 commonsourceibias.n345 161.3
R12533 commonsourceibias.n383 commonsourceibias.n382 161.3
R12534 commonsourceibias.n380 commonsourceibias.n346 161.3
R12535 commonsourceibias.n378 commonsourceibias.n377 161.3
R12536 commonsourceibias.n376 commonsourceibias.n347 161.3
R12537 commonsourceibias.n375 commonsourceibias.n374 161.3
R12538 commonsourceibias.n372 commonsourceibias.n348 161.3
R12539 commonsourceibias.n371 commonsourceibias.n370 161.3
R12540 commonsourceibias.n369 commonsourceibias.n368 161.3
R12541 commonsourceibias.n367 commonsourceibias.n350 161.3
R12542 commonsourceibias.n366 commonsourceibias.n365 161.3
R12543 commonsourceibias.n364 commonsourceibias.n363 161.3
R12544 commonsourceibias.n362 commonsourceibias.n352 161.3
R12545 commonsourceibias.n361 commonsourceibias.n360 161.3
R12546 commonsourceibias.n359 commonsourceibias.n358 161.3
R12547 commonsourceibias.n357 commonsourceibias.n354 161.3
R12548 commonsourceibias.n80 commonsourceibias.n78 81.5057
R12549 commonsourceibias.n240 commonsourceibias.n238 81.5057
R12550 commonsourceibias.n80 commonsourceibias.n79 80.9324
R12551 commonsourceibias.n82 commonsourceibias.n81 80.9324
R12552 commonsourceibias.n77 commonsourceibias.n76 80.9324
R12553 commonsourceibias.n75 commonsourceibias.n74 80.9324
R12554 commonsourceibias.n73 commonsourceibias.n72 80.9324
R12555 commonsourceibias.n307 commonsourceibias.n306 80.9324
R12556 commonsourceibias.n309 commonsourceibias.n308 80.9324
R12557 commonsourceibias.n311 commonsourceibias.n310 80.9324
R12558 commonsourceibias.n242 commonsourceibias.n241 80.9324
R12559 commonsourceibias.n240 commonsourceibias.n239 80.9324
R12560 commonsourceibias.n71 commonsourceibias.n70 80.6037
R12561 commonsourceibias.n137 commonsourceibias.n136 80.6037
R12562 commonsourceibias.n200 commonsourceibias.n199 80.6037
R12563 commonsourceibias.n305 commonsourceibias.n304 80.6037
R12564 commonsourceibias.n339 commonsourceibias.n338 80.6037
R12565 commonsourceibias.n402 commonsourceibias.n401 80.6037
R12566 commonsourceibias.n65 commonsourceibias.n64 56.5617
R12567 commonsourceibias.n51 commonsourceibias.n50 56.5617
R12568 commonsourceibias.n42 commonsourceibias.n41 56.5617
R12569 commonsourceibias.n28 commonsourceibias.n27 56.5617
R12570 commonsourceibias.n131 commonsourceibias.n130 56.5617
R12571 commonsourceibias.n117 commonsourceibias.n116 56.5617
R12572 commonsourceibias.n108 commonsourceibias.n107 56.5617
R12573 commonsourceibias.n94 commonsourceibias.n93 56.5617
R12574 commonsourceibias.n157 commonsourceibias.n156 56.5617
R12575 commonsourceibias.n171 commonsourceibias.n170 56.5617
R12576 commonsourceibias.n180 commonsourceibias.n179 56.5617
R12577 commonsourceibias.n194 commonsourceibias.n193 56.5617
R12578 commonsourceibias.n261 commonsourceibias.n260 56.5617
R12579 commonsourceibias.n275 commonsourceibias.n274 56.5617
R12580 commonsourceibias.n285 commonsourceibias.n283 56.5617
R12581 commonsourceibias.n299 commonsourceibias.n298 56.5617
R12582 commonsourceibias.n333 commonsourceibias.n332 56.5617
R12583 commonsourceibias.n319 commonsourceibias.n317 56.5617
R12584 commonsourceibias.n220 commonsourceibias.n219 56.5617
R12585 commonsourceibias.n234 commonsourceibias.n233 56.5617
R12586 commonsourceibias.n358 commonsourceibias.n357 56.5617
R12587 commonsourceibias.n372 commonsourceibias.n371 56.5617
R12588 commonsourceibias.n382 commonsourceibias.n380 56.5617
R12589 commonsourceibias.n396 commonsourceibias.n395 56.5617
R12590 commonsourceibias.n56 commonsourceibias.n55 56.0773
R12591 commonsourceibias.n37 commonsourceibias.n36 56.0773
R12592 commonsourceibias.n122 commonsourceibias.n121 56.0773
R12593 commonsourceibias.n103 commonsourceibias.n102 56.0773
R12594 commonsourceibias.n166 commonsourceibias.n165 56.0773
R12595 commonsourceibias.n185 commonsourceibias.n184 56.0773
R12596 commonsourceibias.n270 commonsourceibias.n269 56.0773
R12597 commonsourceibias.n290 commonsourceibias.n289 56.0773
R12598 commonsourceibias.n324 commonsourceibias.n323 56.0773
R12599 commonsourceibias.n229 commonsourceibias.n228 56.0773
R12600 commonsourceibias.n367 commonsourceibias.n366 56.0773
R12601 commonsourceibias.n387 commonsourceibias.n386 56.0773
R12602 commonsourceibias.n70 commonsourceibias.n69 46.0096
R12603 commonsourceibias.n136 commonsourceibias.n135 46.0096
R12604 commonsourceibias.n199 commonsourceibias.n198 46.0096
R12605 commonsourceibias.n304 commonsourceibias.n303 46.0096
R12606 commonsourceibias.n338 commonsourceibias.n337 46.0096
R12607 commonsourceibias.n401 commonsourceibias.n400 46.0096
R12608 commonsourceibias.n58 commonsourceibias.n12 41.5458
R12609 commonsourceibias.n33 commonsourceibias.n32 41.5458
R12610 commonsourceibias.n124 commonsourceibias.n3 41.5458
R12611 commonsourceibias.n99 commonsourceibias.n98 41.5458
R12612 commonsourceibias.n162 commonsourceibias.n161 41.5458
R12613 commonsourceibias.n187 commonsourceibias.n141 41.5458
R12614 commonsourceibias.n266 commonsourceibias.n265 41.5458
R12615 commonsourceibias.n292 commonsourceibias.n246 41.5458
R12616 commonsourceibias.n326 commonsourceibias.n205 41.5458
R12617 commonsourceibias.n225 commonsourceibias.n224 41.5458
R12618 commonsourceibias.n363 commonsourceibias.n362 41.5458
R12619 commonsourceibias.n389 commonsourceibias.n343 41.5458
R12620 commonsourceibias.n48 commonsourceibias.n17 40.577
R12621 commonsourceibias.n44 commonsourceibias.n17 40.577
R12622 commonsourceibias.n114 commonsourceibias.n8 40.577
R12623 commonsourceibias.n110 commonsourceibias.n8 40.577
R12624 commonsourceibias.n173 commonsourceibias.n146 40.577
R12625 commonsourceibias.n177 commonsourceibias.n146 40.577
R12626 commonsourceibias.n277 commonsourceibias.n250 40.577
R12627 commonsourceibias.n281 commonsourceibias.n250 40.577
R12628 commonsourceibias.n315 commonsourceibias.n209 40.577
R12629 commonsourceibias.n236 commonsourceibias.n209 40.577
R12630 commonsourceibias.n374 commonsourceibias.n347 40.577
R12631 commonsourceibias.n378 commonsourceibias.n347 40.577
R12632 commonsourceibias.n62 commonsourceibias.n12 39.6083
R12633 commonsourceibias.n32 commonsourceibias.n31 39.6083
R12634 commonsourceibias.n128 commonsourceibias.n3 39.6083
R12635 commonsourceibias.n98 commonsourceibias.n97 39.6083
R12636 commonsourceibias.n161 commonsourceibias.n160 39.6083
R12637 commonsourceibias.n191 commonsourceibias.n141 39.6083
R12638 commonsourceibias.n265 commonsourceibias.n264 39.6083
R12639 commonsourceibias.n296 commonsourceibias.n246 39.6083
R12640 commonsourceibias.n330 commonsourceibias.n205 39.6083
R12641 commonsourceibias.n224 commonsourceibias.n223 39.6083
R12642 commonsourceibias.n362 commonsourceibias.n361 39.6083
R12643 commonsourceibias.n393 commonsourceibias.n343 39.6083
R12644 commonsourceibias.n26 commonsourceibias.n25 33.0515
R12645 commonsourceibias.n92 commonsourceibias.n91 33.0515
R12646 commonsourceibias.n155 commonsourceibias.n154 33.0515
R12647 commonsourceibias.n259 commonsourceibias.n258 33.0515
R12648 commonsourceibias.n218 commonsourceibias.n217 33.0515
R12649 commonsourceibias.n356 commonsourceibias.n355 33.0515
R12650 commonsourceibias.n25 commonsourceibias.n24 28.5514
R12651 commonsourceibias.n91 commonsourceibias.n90 28.5514
R12652 commonsourceibias.n154 commonsourceibias.n153 28.5514
R12653 commonsourceibias.n258 commonsourceibias.n257 28.5514
R12654 commonsourceibias.n217 commonsourceibias.n216 28.5514
R12655 commonsourceibias.n355 commonsourceibias.n354 28.5514
R12656 commonsourceibias.n69 commonsourceibias.n68 26.0455
R12657 commonsourceibias.n135 commonsourceibias.n134 26.0455
R12658 commonsourceibias.n198 commonsourceibias.n197 26.0455
R12659 commonsourceibias.n303 commonsourceibias.n302 26.0455
R12660 commonsourceibias.n337 commonsourceibias.n336 26.0455
R12661 commonsourceibias.n400 commonsourceibias.n399 26.0455
R12662 commonsourceibias.n55 commonsourceibias.n14 25.0767
R12663 commonsourceibias.n38 commonsourceibias.n37 25.0767
R12664 commonsourceibias.n121 commonsourceibias.n5 25.0767
R12665 commonsourceibias.n104 commonsourceibias.n103 25.0767
R12666 commonsourceibias.n167 commonsourceibias.n166 25.0767
R12667 commonsourceibias.n184 commonsourceibias.n143 25.0767
R12668 commonsourceibias.n271 commonsourceibias.n270 25.0767
R12669 commonsourceibias.n289 commonsourceibias.n248 25.0767
R12670 commonsourceibias.n323 commonsourceibias.n207 25.0767
R12671 commonsourceibias.n230 commonsourceibias.n229 25.0767
R12672 commonsourceibias.n368 commonsourceibias.n367 25.0767
R12673 commonsourceibias.n386 commonsourceibias.n345 25.0767
R12674 commonsourceibias.n51 commonsourceibias.n16 24.3464
R12675 commonsourceibias.n41 commonsourceibias.n19 24.3464
R12676 commonsourceibias.n117 commonsourceibias.n7 24.3464
R12677 commonsourceibias.n107 commonsourceibias.n85 24.3464
R12678 commonsourceibias.n170 commonsourceibias.n148 24.3464
R12679 commonsourceibias.n180 commonsourceibias.n145 24.3464
R12680 commonsourceibias.n274 commonsourceibias.n252 24.3464
R12681 commonsourceibias.n285 commonsourceibias.n284 24.3464
R12682 commonsourceibias.n319 commonsourceibias.n318 24.3464
R12683 commonsourceibias.n233 commonsourceibias.n211 24.3464
R12684 commonsourceibias.n371 commonsourceibias.n349 24.3464
R12685 commonsourceibias.n382 commonsourceibias.n381 24.3464
R12686 commonsourceibias.n65 commonsourceibias.n10 23.8546
R12687 commonsourceibias.n27 commonsourceibias.n26 23.8546
R12688 commonsourceibias.n131 commonsourceibias.n1 23.8546
R12689 commonsourceibias.n93 commonsourceibias.n92 23.8546
R12690 commonsourceibias.n156 commonsourceibias.n155 23.8546
R12691 commonsourceibias.n194 commonsourceibias.n139 23.8546
R12692 commonsourceibias.n260 commonsourceibias.n259 23.8546
R12693 commonsourceibias.n299 commonsourceibias.n244 23.8546
R12694 commonsourceibias.n333 commonsourceibias.n203 23.8546
R12695 commonsourceibias.n219 commonsourceibias.n218 23.8546
R12696 commonsourceibias.n357 commonsourceibias.n356 23.8546
R12697 commonsourceibias.n396 commonsourceibias.n341 23.8546
R12698 commonsourceibias.n64 commonsourceibias.n63 16.9689
R12699 commonsourceibias.n28 commonsourceibias.n23 16.9689
R12700 commonsourceibias.n130 commonsourceibias.n129 16.9689
R12701 commonsourceibias.n94 commonsourceibias.n89 16.9689
R12702 commonsourceibias.n157 commonsourceibias.n152 16.9689
R12703 commonsourceibias.n193 commonsourceibias.n192 16.9689
R12704 commonsourceibias.n261 commonsourceibias.n256 16.9689
R12705 commonsourceibias.n298 commonsourceibias.n297 16.9689
R12706 commonsourceibias.n332 commonsourceibias.n331 16.9689
R12707 commonsourceibias.n220 commonsourceibias.n215 16.9689
R12708 commonsourceibias.n358 commonsourceibias.n353 16.9689
R12709 commonsourceibias.n395 commonsourceibias.n394 16.9689
R12710 commonsourceibias.n50 commonsourceibias.n49 16.477
R12711 commonsourceibias.n43 commonsourceibias.n42 16.477
R12712 commonsourceibias.n116 commonsourceibias.n115 16.477
R12713 commonsourceibias.n109 commonsourceibias.n108 16.477
R12714 commonsourceibias.n172 commonsourceibias.n171 16.477
R12715 commonsourceibias.n179 commonsourceibias.n178 16.477
R12716 commonsourceibias.n276 commonsourceibias.n275 16.477
R12717 commonsourceibias.n283 commonsourceibias.n282 16.477
R12718 commonsourceibias.n317 commonsourceibias.n316 16.477
R12719 commonsourceibias.n235 commonsourceibias.n234 16.477
R12720 commonsourceibias.n373 commonsourceibias.n372 16.477
R12721 commonsourceibias.n380 commonsourceibias.n379 16.477
R12722 commonsourceibias.n57 commonsourceibias.n56 15.9852
R12723 commonsourceibias.n36 commonsourceibias.n21 15.9852
R12724 commonsourceibias.n123 commonsourceibias.n122 15.9852
R12725 commonsourceibias.n102 commonsourceibias.n87 15.9852
R12726 commonsourceibias.n165 commonsourceibias.n150 15.9852
R12727 commonsourceibias.n186 commonsourceibias.n185 15.9852
R12728 commonsourceibias.n269 commonsourceibias.n254 15.9852
R12729 commonsourceibias.n291 commonsourceibias.n290 15.9852
R12730 commonsourceibias.n325 commonsourceibias.n324 15.9852
R12731 commonsourceibias.n228 commonsourceibias.n213 15.9852
R12732 commonsourceibias.n366 commonsourceibias.n351 15.9852
R12733 commonsourceibias.n388 commonsourceibias.n387 15.9852
R12734 commonsourceibias.n73 commonsourceibias.n71 13.2057
R12735 commonsourceibias.n307 commonsourceibias.n305 13.2057
R12736 commonsourceibias.n404 commonsourceibias.n201 11.9876
R12737 commonsourceibias.n404 commonsourceibias.n403 10.3347
R12738 commonsourceibias.n112 commonsourceibias.n83 9.50363
R12739 commonsourceibias.n313 commonsourceibias.n312 9.50363
R12740 commonsourceibias.n201 commonsourceibias.n137 8.732
R12741 commonsourceibias.n403 commonsourceibias.n339 8.732
R12742 commonsourceibias.n58 commonsourceibias.n57 8.60764
R12743 commonsourceibias.n33 commonsourceibias.n21 8.60764
R12744 commonsourceibias.n124 commonsourceibias.n123 8.60764
R12745 commonsourceibias.n99 commonsourceibias.n87 8.60764
R12746 commonsourceibias.n162 commonsourceibias.n150 8.60764
R12747 commonsourceibias.n187 commonsourceibias.n186 8.60764
R12748 commonsourceibias.n266 commonsourceibias.n254 8.60764
R12749 commonsourceibias.n292 commonsourceibias.n291 8.60764
R12750 commonsourceibias.n326 commonsourceibias.n325 8.60764
R12751 commonsourceibias.n225 commonsourceibias.n213 8.60764
R12752 commonsourceibias.n363 commonsourceibias.n351 8.60764
R12753 commonsourceibias.n389 commonsourceibias.n388 8.60764
R12754 commonsourceibias.n49 commonsourceibias.n48 8.11581
R12755 commonsourceibias.n44 commonsourceibias.n43 8.11581
R12756 commonsourceibias.n115 commonsourceibias.n114 8.11581
R12757 commonsourceibias.n110 commonsourceibias.n109 8.11581
R12758 commonsourceibias.n173 commonsourceibias.n172 8.11581
R12759 commonsourceibias.n178 commonsourceibias.n177 8.11581
R12760 commonsourceibias.n277 commonsourceibias.n276 8.11581
R12761 commonsourceibias.n282 commonsourceibias.n281 8.11581
R12762 commonsourceibias.n316 commonsourceibias.n315 8.11581
R12763 commonsourceibias.n236 commonsourceibias.n235 8.11581
R12764 commonsourceibias.n374 commonsourceibias.n373 8.11581
R12765 commonsourceibias.n379 commonsourceibias.n378 8.11581
R12766 commonsourceibias.n63 commonsourceibias.n62 7.62397
R12767 commonsourceibias.n31 commonsourceibias.n23 7.62397
R12768 commonsourceibias.n129 commonsourceibias.n128 7.62397
R12769 commonsourceibias.n97 commonsourceibias.n89 7.62397
R12770 commonsourceibias.n160 commonsourceibias.n152 7.62397
R12771 commonsourceibias.n192 commonsourceibias.n191 7.62397
R12772 commonsourceibias.n264 commonsourceibias.n256 7.62397
R12773 commonsourceibias.n297 commonsourceibias.n296 7.62397
R12774 commonsourceibias.n331 commonsourceibias.n330 7.62397
R12775 commonsourceibias.n223 commonsourceibias.n215 7.62397
R12776 commonsourceibias.n361 commonsourceibias.n353 7.62397
R12777 commonsourceibias.n394 commonsourceibias.n393 7.62397
R12778 commonsourceibias.n201 commonsourceibias.n200 5.00473
R12779 commonsourceibias.n403 commonsourceibias.n402 5.00473
R12780 commonsourceibias commonsourceibias.n404 3.87639
R12781 commonsourceibias.n78 commonsourceibias.t41 2.82907
R12782 commonsourceibias.n78 commonsourceibias.t47 2.82907
R12783 commonsourceibias.n79 commonsourceibias.t35 2.82907
R12784 commonsourceibias.n79 commonsourceibias.t11 2.82907
R12785 commonsourceibias.n81 commonsourceibias.t45 2.82907
R12786 commonsourceibias.n81 commonsourceibias.t27 2.82907
R12787 commonsourceibias.n76 commonsourceibias.t21 2.82907
R12788 commonsourceibias.n76 commonsourceibias.t37 2.82907
R12789 commonsourceibias.n74 commonsourceibias.t25 2.82907
R12790 commonsourceibias.n74 commonsourceibias.t31 2.82907
R12791 commonsourceibias.n72 commonsourceibias.t33 2.82907
R12792 commonsourceibias.n72 commonsourceibias.t15 2.82907
R12793 commonsourceibias.n306 commonsourceibias.t23 2.82907
R12794 commonsourceibias.n306 commonsourceibias.t3 2.82907
R12795 commonsourceibias.n308 commonsourceibias.t1 2.82907
R12796 commonsourceibias.n308 commonsourceibias.t39 2.82907
R12797 commonsourceibias.n310 commonsourceibias.t7 2.82907
R12798 commonsourceibias.n310 commonsourceibias.t29 2.82907
R12799 commonsourceibias.n241 commonsourceibias.t43 2.82907
R12800 commonsourceibias.n241 commonsourceibias.t13 2.82907
R12801 commonsourceibias.n239 commonsourceibias.t19 2.82907
R12802 commonsourceibias.n239 commonsourceibias.t5 2.82907
R12803 commonsourceibias.n238 commonsourceibias.t17 2.82907
R12804 commonsourceibias.n238 commonsourceibias.t9 2.82907
R12805 commonsourceibias.n68 commonsourceibias.n10 0.738255
R12806 commonsourceibias.n134 commonsourceibias.n1 0.738255
R12807 commonsourceibias.n197 commonsourceibias.n139 0.738255
R12808 commonsourceibias.n302 commonsourceibias.n244 0.738255
R12809 commonsourceibias.n336 commonsourceibias.n203 0.738255
R12810 commonsourceibias.n399 commonsourceibias.n341 0.738255
R12811 commonsourceibias.n75 commonsourceibias.n73 0.573776
R12812 commonsourceibias.n77 commonsourceibias.n75 0.573776
R12813 commonsourceibias.n82 commonsourceibias.n80 0.573776
R12814 commonsourceibias.n242 commonsourceibias.n240 0.573776
R12815 commonsourceibias.n311 commonsourceibias.n309 0.573776
R12816 commonsourceibias.n309 commonsourceibias.n307 0.573776
R12817 commonsourceibias.n83 commonsourceibias.n77 0.287138
R12818 commonsourceibias.n83 commonsourceibias.n82 0.287138
R12819 commonsourceibias.n312 commonsourceibias.n242 0.287138
R12820 commonsourceibias.n312 commonsourceibias.n311 0.287138
R12821 commonsourceibias.n71 commonsourceibias.n9 0.285035
R12822 commonsourceibias.n137 commonsourceibias.n0 0.285035
R12823 commonsourceibias.n200 commonsourceibias.n138 0.285035
R12824 commonsourceibias.n305 commonsourceibias.n243 0.285035
R12825 commonsourceibias.n339 commonsourceibias.n202 0.285035
R12826 commonsourceibias.n402 commonsourceibias.n340 0.285035
R12827 commonsourceibias.n16 commonsourceibias.n14 0.246418
R12828 commonsourceibias.n38 commonsourceibias.n19 0.246418
R12829 commonsourceibias.n7 commonsourceibias.n5 0.246418
R12830 commonsourceibias.n104 commonsourceibias.n85 0.246418
R12831 commonsourceibias.n167 commonsourceibias.n148 0.246418
R12832 commonsourceibias.n145 commonsourceibias.n143 0.246418
R12833 commonsourceibias.n271 commonsourceibias.n252 0.246418
R12834 commonsourceibias.n284 commonsourceibias.n248 0.246418
R12835 commonsourceibias.n318 commonsourceibias.n207 0.246418
R12836 commonsourceibias.n230 commonsourceibias.n211 0.246418
R12837 commonsourceibias.n368 commonsourceibias.n349 0.246418
R12838 commonsourceibias.n381 commonsourceibias.n345 0.246418
R12839 commonsourceibias.n67 commonsourceibias.n9 0.189894
R12840 commonsourceibias.n67 commonsourceibias.n66 0.189894
R12841 commonsourceibias.n66 commonsourceibias.n11 0.189894
R12842 commonsourceibias.n61 commonsourceibias.n11 0.189894
R12843 commonsourceibias.n61 commonsourceibias.n60 0.189894
R12844 commonsourceibias.n60 commonsourceibias.n59 0.189894
R12845 commonsourceibias.n59 commonsourceibias.n13 0.189894
R12846 commonsourceibias.n54 commonsourceibias.n13 0.189894
R12847 commonsourceibias.n54 commonsourceibias.n53 0.189894
R12848 commonsourceibias.n53 commonsourceibias.n52 0.189894
R12849 commonsourceibias.n52 commonsourceibias.n15 0.189894
R12850 commonsourceibias.n47 commonsourceibias.n15 0.189894
R12851 commonsourceibias.n47 commonsourceibias.n46 0.189894
R12852 commonsourceibias.n46 commonsourceibias.n45 0.189894
R12853 commonsourceibias.n45 commonsourceibias.n18 0.189894
R12854 commonsourceibias.n40 commonsourceibias.n18 0.189894
R12855 commonsourceibias.n40 commonsourceibias.n39 0.189894
R12856 commonsourceibias.n39 commonsourceibias.n20 0.189894
R12857 commonsourceibias.n35 commonsourceibias.n20 0.189894
R12858 commonsourceibias.n35 commonsourceibias.n34 0.189894
R12859 commonsourceibias.n34 commonsourceibias.n22 0.189894
R12860 commonsourceibias.n30 commonsourceibias.n22 0.189894
R12861 commonsourceibias.n30 commonsourceibias.n29 0.189894
R12862 commonsourceibias.n29 commonsourceibias.n24 0.189894
R12863 commonsourceibias.n111 commonsourceibias.n84 0.189894
R12864 commonsourceibias.n106 commonsourceibias.n84 0.189894
R12865 commonsourceibias.n106 commonsourceibias.n105 0.189894
R12866 commonsourceibias.n105 commonsourceibias.n86 0.189894
R12867 commonsourceibias.n101 commonsourceibias.n86 0.189894
R12868 commonsourceibias.n101 commonsourceibias.n100 0.189894
R12869 commonsourceibias.n100 commonsourceibias.n88 0.189894
R12870 commonsourceibias.n96 commonsourceibias.n88 0.189894
R12871 commonsourceibias.n96 commonsourceibias.n95 0.189894
R12872 commonsourceibias.n95 commonsourceibias.n90 0.189894
R12873 commonsourceibias.n133 commonsourceibias.n0 0.189894
R12874 commonsourceibias.n133 commonsourceibias.n132 0.189894
R12875 commonsourceibias.n132 commonsourceibias.n2 0.189894
R12876 commonsourceibias.n127 commonsourceibias.n2 0.189894
R12877 commonsourceibias.n127 commonsourceibias.n126 0.189894
R12878 commonsourceibias.n126 commonsourceibias.n125 0.189894
R12879 commonsourceibias.n125 commonsourceibias.n4 0.189894
R12880 commonsourceibias.n120 commonsourceibias.n4 0.189894
R12881 commonsourceibias.n120 commonsourceibias.n119 0.189894
R12882 commonsourceibias.n119 commonsourceibias.n118 0.189894
R12883 commonsourceibias.n118 commonsourceibias.n6 0.189894
R12884 commonsourceibias.n113 commonsourceibias.n6 0.189894
R12885 commonsourceibias.n196 commonsourceibias.n138 0.189894
R12886 commonsourceibias.n196 commonsourceibias.n195 0.189894
R12887 commonsourceibias.n195 commonsourceibias.n140 0.189894
R12888 commonsourceibias.n190 commonsourceibias.n140 0.189894
R12889 commonsourceibias.n190 commonsourceibias.n189 0.189894
R12890 commonsourceibias.n189 commonsourceibias.n188 0.189894
R12891 commonsourceibias.n188 commonsourceibias.n142 0.189894
R12892 commonsourceibias.n183 commonsourceibias.n142 0.189894
R12893 commonsourceibias.n183 commonsourceibias.n182 0.189894
R12894 commonsourceibias.n182 commonsourceibias.n181 0.189894
R12895 commonsourceibias.n181 commonsourceibias.n144 0.189894
R12896 commonsourceibias.n176 commonsourceibias.n144 0.189894
R12897 commonsourceibias.n176 commonsourceibias.n175 0.189894
R12898 commonsourceibias.n175 commonsourceibias.n174 0.189894
R12899 commonsourceibias.n174 commonsourceibias.n147 0.189894
R12900 commonsourceibias.n169 commonsourceibias.n147 0.189894
R12901 commonsourceibias.n169 commonsourceibias.n168 0.189894
R12902 commonsourceibias.n168 commonsourceibias.n149 0.189894
R12903 commonsourceibias.n164 commonsourceibias.n149 0.189894
R12904 commonsourceibias.n164 commonsourceibias.n163 0.189894
R12905 commonsourceibias.n163 commonsourceibias.n151 0.189894
R12906 commonsourceibias.n159 commonsourceibias.n151 0.189894
R12907 commonsourceibias.n159 commonsourceibias.n158 0.189894
R12908 commonsourceibias.n158 commonsourceibias.n153 0.189894
R12909 commonsourceibias.n262 commonsourceibias.n257 0.189894
R12910 commonsourceibias.n263 commonsourceibias.n262 0.189894
R12911 commonsourceibias.n263 commonsourceibias.n255 0.189894
R12912 commonsourceibias.n267 commonsourceibias.n255 0.189894
R12913 commonsourceibias.n268 commonsourceibias.n267 0.189894
R12914 commonsourceibias.n268 commonsourceibias.n253 0.189894
R12915 commonsourceibias.n272 commonsourceibias.n253 0.189894
R12916 commonsourceibias.n273 commonsourceibias.n272 0.189894
R12917 commonsourceibias.n273 commonsourceibias.n251 0.189894
R12918 commonsourceibias.n278 commonsourceibias.n251 0.189894
R12919 commonsourceibias.n279 commonsourceibias.n278 0.189894
R12920 commonsourceibias.n280 commonsourceibias.n279 0.189894
R12921 commonsourceibias.n280 commonsourceibias.n249 0.189894
R12922 commonsourceibias.n286 commonsourceibias.n249 0.189894
R12923 commonsourceibias.n287 commonsourceibias.n286 0.189894
R12924 commonsourceibias.n288 commonsourceibias.n287 0.189894
R12925 commonsourceibias.n288 commonsourceibias.n247 0.189894
R12926 commonsourceibias.n293 commonsourceibias.n247 0.189894
R12927 commonsourceibias.n294 commonsourceibias.n293 0.189894
R12928 commonsourceibias.n295 commonsourceibias.n294 0.189894
R12929 commonsourceibias.n295 commonsourceibias.n245 0.189894
R12930 commonsourceibias.n300 commonsourceibias.n245 0.189894
R12931 commonsourceibias.n301 commonsourceibias.n300 0.189894
R12932 commonsourceibias.n301 commonsourceibias.n243 0.189894
R12933 commonsourceibias.n221 commonsourceibias.n216 0.189894
R12934 commonsourceibias.n222 commonsourceibias.n221 0.189894
R12935 commonsourceibias.n222 commonsourceibias.n214 0.189894
R12936 commonsourceibias.n226 commonsourceibias.n214 0.189894
R12937 commonsourceibias.n227 commonsourceibias.n226 0.189894
R12938 commonsourceibias.n227 commonsourceibias.n212 0.189894
R12939 commonsourceibias.n231 commonsourceibias.n212 0.189894
R12940 commonsourceibias.n232 commonsourceibias.n231 0.189894
R12941 commonsourceibias.n232 commonsourceibias.n210 0.189894
R12942 commonsourceibias.n237 commonsourceibias.n210 0.189894
R12943 commonsourceibias.n314 commonsourceibias.n208 0.189894
R12944 commonsourceibias.n320 commonsourceibias.n208 0.189894
R12945 commonsourceibias.n321 commonsourceibias.n320 0.189894
R12946 commonsourceibias.n322 commonsourceibias.n321 0.189894
R12947 commonsourceibias.n322 commonsourceibias.n206 0.189894
R12948 commonsourceibias.n327 commonsourceibias.n206 0.189894
R12949 commonsourceibias.n328 commonsourceibias.n327 0.189894
R12950 commonsourceibias.n329 commonsourceibias.n328 0.189894
R12951 commonsourceibias.n329 commonsourceibias.n204 0.189894
R12952 commonsourceibias.n334 commonsourceibias.n204 0.189894
R12953 commonsourceibias.n335 commonsourceibias.n334 0.189894
R12954 commonsourceibias.n335 commonsourceibias.n202 0.189894
R12955 commonsourceibias.n359 commonsourceibias.n354 0.189894
R12956 commonsourceibias.n360 commonsourceibias.n359 0.189894
R12957 commonsourceibias.n360 commonsourceibias.n352 0.189894
R12958 commonsourceibias.n364 commonsourceibias.n352 0.189894
R12959 commonsourceibias.n365 commonsourceibias.n364 0.189894
R12960 commonsourceibias.n365 commonsourceibias.n350 0.189894
R12961 commonsourceibias.n369 commonsourceibias.n350 0.189894
R12962 commonsourceibias.n370 commonsourceibias.n369 0.189894
R12963 commonsourceibias.n370 commonsourceibias.n348 0.189894
R12964 commonsourceibias.n375 commonsourceibias.n348 0.189894
R12965 commonsourceibias.n376 commonsourceibias.n375 0.189894
R12966 commonsourceibias.n377 commonsourceibias.n376 0.189894
R12967 commonsourceibias.n377 commonsourceibias.n346 0.189894
R12968 commonsourceibias.n383 commonsourceibias.n346 0.189894
R12969 commonsourceibias.n384 commonsourceibias.n383 0.189894
R12970 commonsourceibias.n385 commonsourceibias.n384 0.189894
R12971 commonsourceibias.n385 commonsourceibias.n344 0.189894
R12972 commonsourceibias.n390 commonsourceibias.n344 0.189894
R12973 commonsourceibias.n391 commonsourceibias.n390 0.189894
R12974 commonsourceibias.n392 commonsourceibias.n391 0.189894
R12975 commonsourceibias.n392 commonsourceibias.n342 0.189894
R12976 commonsourceibias.n397 commonsourceibias.n342 0.189894
R12977 commonsourceibias.n398 commonsourceibias.n397 0.189894
R12978 commonsourceibias.n398 commonsourceibias.n340 0.189894
R12979 commonsourceibias.n112 commonsourceibias.n111 0.170955
R12980 commonsourceibias.n113 commonsourceibias.n112 0.170955
R12981 commonsourceibias.n313 commonsourceibias.n237 0.170955
R12982 commonsourceibias.n314 commonsourceibias.n313 0.170955
R12983 CSoutput.n19 CSoutput.t117 184.661
R12984 CSoutput.n78 CSoutput.n77 165.8
R12985 CSoutput.n76 CSoutput.n0 165.8
R12986 CSoutput.n75 CSoutput.n74 165.8
R12987 CSoutput.n73 CSoutput.n72 165.8
R12988 CSoutput.n71 CSoutput.n2 165.8
R12989 CSoutput.n69 CSoutput.n68 165.8
R12990 CSoutput.n67 CSoutput.n3 165.8
R12991 CSoutput.n66 CSoutput.n65 165.8
R12992 CSoutput.n63 CSoutput.n4 165.8
R12993 CSoutput.n61 CSoutput.n60 165.8
R12994 CSoutput.n59 CSoutput.n5 165.8
R12995 CSoutput.n58 CSoutput.n57 165.8
R12996 CSoutput.n55 CSoutput.n6 165.8
R12997 CSoutput.n54 CSoutput.n53 165.8
R12998 CSoutput.n52 CSoutput.n51 165.8
R12999 CSoutput.n50 CSoutput.n8 165.8
R13000 CSoutput.n48 CSoutput.n47 165.8
R13001 CSoutput.n46 CSoutput.n9 165.8
R13002 CSoutput.n45 CSoutput.n44 165.8
R13003 CSoutput.n42 CSoutput.n10 165.8
R13004 CSoutput.n41 CSoutput.n40 165.8
R13005 CSoutput.n39 CSoutput.n38 165.8
R13006 CSoutput.n37 CSoutput.n12 165.8
R13007 CSoutput.n35 CSoutput.n34 165.8
R13008 CSoutput.n33 CSoutput.n13 165.8
R13009 CSoutput.n32 CSoutput.n31 165.8
R13010 CSoutput.n29 CSoutput.n14 165.8
R13011 CSoutput.n28 CSoutput.n27 165.8
R13012 CSoutput.n26 CSoutput.n25 165.8
R13013 CSoutput.n24 CSoutput.n16 165.8
R13014 CSoutput.n22 CSoutput.n21 165.8
R13015 CSoutput.n20 CSoutput.n17 165.8
R13016 CSoutput.n77 CSoutput.t96 162.194
R13017 CSoutput.n18 CSoutput.t97 120.501
R13018 CSoutput.n23 CSoutput.t107 120.501
R13019 CSoutput.n15 CSoutput.t103 120.501
R13020 CSoutput.n30 CSoutput.t99 120.501
R13021 CSoutput.n36 CSoutput.t110 120.501
R13022 CSoutput.n11 CSoutput.t112 120.501
R13023 CSoutput.n43 CSoutput.t101 120.501
R13024 CSoutput.n49 CSoutput.t113 120.501
R13025 CSoutput.n7 CSoutput.t114 120.501
R13026 CSoutput.n56 CSoutput.t108 120.501
R13027 CSoutput.n62 CSoutput.t100 120.501
R13028 CSoutput.n64 CSoutput.t116 120.501
R13029 CSoutput.n70 CSoutput.t111 120.501
R13030 CSoutput.n1 CSoutput.t106 120.501
R13031 CSoutput.n270 CSoutput.n268 103.469
R13032 CSoutput.n262 CSoutput.n260 103.469
R13033 CSoutput.n255 CSoutput.n253 103.469
R13034 CSoutput.n96 CSoutput.n94 103.469
R13035 CSoutput.n88 CSoutput.n86 103.469
R13036 CSoutput.n81 CSoutput.n79 103.469
R13037 CSoutput.n272 CSoutput.n271 103.111
R13038 CSoutput.n270 CSoutput.n269 103.111
R13039 CSoutput.n266 CSoutput.n265 103.111
R13040 CSoutput.n264 CSoutput.n263 103.111
R13041 CSoutput.n262 CSoutput.n261 103.111
R13042 CSoutput.n259 CSoutput.n258 103.111
R13043 CSoutput.n257 CSoutput.n256 103.111
R13044 CSoutput.n255 CSoutput.n254 103.111
R13045 CSoutput.n96 CSoutput.n95 103.111
R13046 CSoutput.n98 CSoutput.n97 103.111
R13047 CSoutput.n100 CSoutput.n99 103.111
R13048 CSoutput.n88 CSoutput.n87 103.111
R13049 CSoutput.n90 CSoutput.n89 103.111
R13050 CSoutput.n92 CSoutput.n91 103.111
R13051 CSoutput.n81 CSoutput.n80 103.111
R13052 CSoutput.n83 CSoutput.n82 103.111
R13053 CSoutput.n85 CSoutput.n84 103.111
R13054 CSoutput.n274 CSoutput.n273 103.111
R13055 CSoutput.n290 CSoutput.n288 81.5057
R13056 CSoutput.n279 CSoutput.n277 81.5057
R13057 CSoutput.n314 CSoutput.n312 81.5057
R13058 CSoutput.n303 CSoutput.n301 81.5057
R13059 CSoutput.n298 CSoutput.n297 80.9324
R13060 CSoutput.n296 CSoutput.n295 80.9324
R13061 CSoutput.n294 CSoutput.n293 80.9324
R13062 CSoutput.n292 CSoutput.n291 80.9324
R13063 CSoutput.n290 CSoutput.n289 80.9324
R13064 CSoutput.n287 CSoutput.n286 80.9324
R13065 CSoutput.n285 CSoutput.n284 80.9324
R13066 CSoutput.n283 CSoutput.n282 80.9324
R13067 CSoutput.n281 CSoutput.n280 80.9324
R13068 CSoutput.n279 CSoutput.n278 80.9324
R13069 CSoutput.n314 CSoutput.n313 80.9324
R13070 CSoutput.n316 CSoutput.n315 80.9324
R13071 CSoutput.n318 CSoutput.n317 80.9324
R13072 CSoutput.n320 CSoutput.n319 80.9324
R13073 CSoutput.n322 CSoutput.n321 80.9324
R13074 CSoutput.n303 CSoutput.n302 80.9324
R13075 CSoutput.n305 CSoutput.n304 80.9324
R13076 CSoutput.n307 CSoutput.n306 80.9324
R13077 CSoutput.n309 CSoutput.n308 80.9324
R13078 CSoutput.n311 CSoutput.n310 80.9324
R13079 CSoutput.n25 CSoutput.n24 48.1486
R13080 CSoutput.n69 CSoutput.n3 48.1486
R13081 CSoutput.n38 CSoutput.n37 48.1486
R13082 CSoutput.n42 CSoutput.n41 48.1486
R13083 CSoutput.n51 CSoutput.n50 48.1486
R13084 CSoutput.n55 CSoutput.n54 48.1486
R13085 CSoutput.n22 CSoutput.n17 46.462
R13086 CSoutput.n72 CSoutput.n71 46.462
R13087 CSoutput.n20 CSoutput.n19 44.9055
R13088 CSoutput.n29 CSoutput.n28 43.7635
R13089 CSoutput.n65 CSoutput.n63 43.7635
R13090 CSoutput.n35 CSoutput.n13 41.7396
R13091 CSoutput.n57 CSoutput.n5 41.7396
R13092 CSoutput.n44 CSoutput.n9 37.0171
R13093 CSoutput.n48 CSoutput.n9 37.0171
R13094 CSoutput.n76 CSoutput.n75 34.9932
R13095 CSoutput.n31 CSoutput.n13 32.2947
R13096 CSoutput.n61 CSoutput.n5 32.2947
R13097 CSoutput.n30 CSoutput.n29 29.6014
R13098 CSoutput.n63 CSoutput.n62 29.6014
R13099 CSoutput.n19 CSoutput.n18 28.4085
R13100 CSoutput.n18 CSoutput.n17 25.1176
R13101 CSoutput.n72 CSoutput.n1 25.1176
R13102 CSoutput.n43 CSoutput.n42 22.0922
R13103 CSoutput.n50 CSoutput.n49 22.0922
R13104 CSoutput.n77 CSoutput.n76 21.8586
R13105 CSoutput.n37 CSoutput.n36 18.9681
R13106 CSoutput.n56 CSoutput.n55 18.9681
R13107 CSoutput.n25 CSoutput.n15 17.6292
R13108 CSoutput.n64 CSoutput.n3 17.6292
R13109 CSoutput.n24 CSoutput.n23 15.844
R13110 CSoutput.n70 CSoutput.n69 15.844
R13111 CSoutput.n38 CSoutput.n11 14.5051
R13112 CSoutput.n54 CSoutput.n7 14.5051
R13113 CSoutput.n325 CSoutput.n78 11.6139
R13114 CSoutput.n41 CSoutput.n11 11.3811
R13115 CSoutput.n51 CSoutput.n7 11.3811
R13116 CSoutput.n23 CSoutput.n22 10.0422
R13117 CSoutput.n71 CSoutput.n70 10.0422
R13118 CSoutput.n267 CSoutput.n259 9.25285
R13119 CSoutput.n93 CSoutput.n85 9.25285
R13120 CSoutput.n299 CSoutput.n287 8.97993
R13121 CSoutput.n323 CSoutput.n311 8.97993
R13122 CSoutput.n300 CSoutput.n276 8.92829
R13123 CSoutput.n28 CSoutput.n15 8.25698
R13124 CSoutput.n65 CSoutput.n64 8.25698
R13125 CSoutput.n300 CSoutput.n299 7.89345
R13126 CSoutput.n324 CSoutput.n323 7.89345
R13127 CSoutput.n276 CSoutput.n275 7.12641
R13128 CSoutput.n102 CSoutput.n101 7.12641
R13129 CSoutput.n36 CSoutput.n35 6.91809
R13130 CSoutput.n57 CSoutput.n56 6.91809
R13131 CSoutput.n325 CSoutput.n102 5.33585
R13132 CSoutput.n299 CSoutput.n298 5.25266
R13133 CSoutput.n323 CSoutput.n322 5.25266
R13134 CSoutput.n275 CSoutput.n274 5.1449
R13135 CSoutput.n267 CSoutput.n266 5.1449
R13136 CSoutput.n101 CSoutput.n100 5.1449
R13137 CSoutput.n93 CSoutput.n92 5.1449
R13138 CSoutput.n193 CSoutput.n146 4.5005
R13139 CSoutput.n162 CSoutput.n146 4.5005
R13140 CSoutput.n157 CSoutput.n141 4.5005
R13141 CSoutput.n157 CSoutput.n143 4.5005
R13142 CSoutput.n157 CSoutput.n140 4.5005
R13143 CSoutput.n157 CSoutput.n144 4.5005
R13144 CSoutput.n157 CSoutput.n139 4.5005
R13145 CSoutput.n157 CSoutput.t102 4.5005
R13146 CSoutput.n157 CSoutput.n138 4.5005
R13147 CSoutput.n157 CSoutput.n145 4.5005
R13148 CSoutput.n157 CSoutput.n146 4.5005
R13149 CSoutput.n155 CSoutput.n141 4.5005
R13150 CSoutput.n155 CSoutput.n143 4.5005
R13151 CSoutput.n155 CSoutput.n140 4.5005
R13152 CSoutput.n155 CSoutput.n144 4.5005
R13153 CSoutput.n155 CSoutput.n139 4.5005
R13154 CSoutput.n155 CSoutput.t102 4.5005
R13155 CSoutput.n155 CSoutput.n138 4.5005
R13156 CSoutput.n155 CSoutput.n145 4.5005
R13157 CSoutput.n155 CSoutput.n146 4.5005
R13158 CSoutput.n154 CSoutput.n141 4.5005
R13159 CSoutput.n154 CSoutput.n143 4.5005
R13160 CSoutput.n154 CSoutput.n140 4.5005
R13161 CSoutput.n154 CSoutput.n144 4.5005
R13162 CSoutput.n154 CSoutput.n139 4.5005
R13163 CSoutput.n154 CSoutput.t102 4.5005
R13164 CSoutput.n154 CSoutput.n138 4.5005
R13165 CSoutput.n154 CSoutput.n145 4.5005
R13166 CSoutput.n154 CSoutput.n146 4.5005
R13167 CSoutput.n239 CSoutput.n141 4.5005
R13168 CSoutput.n239 CSoutput.n143 4.5005
R13169 CSoutput.n239 CSoutput.n140 4.5005
R13170 CSoutput.n239 CSoutput.n144 4.5005
R13171 CSoutput.n239 CSoutput.n139 4.5005
R13172 CSoutput.n239 CSoutput.t102 4.5005
R13173 CSoutput.n239 CSoutput.n138 4.5005
R13174 CSoutput.n239 CSoutput.n145 4.5005
R13175 CSoutput.n239 CSoutput.n146 4.5005
R13176 CSoutput.n237 CSoutput.n141 4.5005
R13177 CSoutput.n237 CSoutput.n143 4.5005
R13178 CSoutput.n237 CSoutput.n140 4.5005
R13179 CSoutput.n237 CSoutput.n144 4.5005
R13180 CSoutput.n237 CSoutput.n139 4.5005
R13181 CSoutput.n237 CSoutput.t102 4.5005
R13182 CSoutput.n237 CSoutput.n138 4.5005
R13183 CSoutput.n237 CSoutput.n145 4.5005
R13184 CSoutput.n235 CSoutput.n141 4.5005
R13185 CSoutput.n235 CSoutput.n143 4.5005
R13186 CSoutput.n235 CSoutput.n140 4.5005
R13187 CSoutput.n235 CSoutput.n144 4.5005
R13188 CSoutput.n235 CSoutput.n139 4.5005
R13189 CSoutput.n235 CSoutput.t102 4.5005
R13190 CSoutput.n235 CSoutput.n138 4.5005
R13191 CSoutput.n235 CSoutput.n145 4.5005
R13192 CSoutput.n165 CSoutput.n141 4.5005
R13193 CSoutput.n165 CSoutput.n143 4.5005
R13194 CSoutput.n165 CSoutput.n140 4.5005
R13195 CSoutput.n165 CSoutput.n144 4.5005
R13196 CSoutput.n165 CSoutput.n139 4.5005
R13197 CSoutput.n165 CSoutput.t102 4.5005
R13198 CSoutput.n165 CSoutput.n138 4.5005
R13199 CSoutput.n165 CSoutput.n145 4.5005
R13200 CSoutput.n165 CSoutput.n146 4.5005
R13201 CSoutput.n164 CSoutput.n141 4.5005
R13202 CSoutput.n164 CSoutput.n143 4.5005
R13203 CSoutput.n164 CSoutput.n140 4.5005
R13204 CSoutput.n164 CSoutput.n144 4.5005
R13205 CSoutput.n164 CSoutput.n139 4.5005
R13206 CSoutput.n164 CSoutput.t102 4.5005
R13207 CSoutput.n164 CSoutput.n138 4.5005
R13208 CSoutput.n164 CSoutput.n145 4.5005
R13209 CSoutput.n164 CSoutput.n146 4.5005
R13210 CSoutput.n168 CSoutput.n141 4.5005
R13211 CSoutput.n168 CSoutput.n143 4.5005
R13212 CSoutput.n168 CSoutput.n140 4.5005
R13213 CSoutput.n168 CSoutput.n144 4.5005
R13214 CSoutput.n168 CSoutput.n139 4.5005
R13215 CSoutput.n168 CSoutput.t102 4.5005
R13216 CSoutput.n168 CSoutput.n138 4.5005
R13217 CSoutput.n168 CSoutput.n145 4.5005
R13218 CSoutput.n168 CSoutput.n146 4.5005
R13219 CSoutput.n167 CSoutput.n141 4.5005
R13220 CSoutput.n167 CSoutput.n143 4.5005
R13221 CSoutput.n167 CSoutput.n140 4.5005
R13222 CSoutput.n167 CSoutput.n144 4.5005
R13223 CSoutput.n167 CSoutput.n139 4.5005
R13224 CSoutput.n167 CSoutput.t102 4.5005
R13225 CSoutput.n167 CSoutput.n138 4.5005
R13226 CSoutput.n167 CSoutput.n145 4.5005
R13227 CSoutput.n167 CSoutput.n146 4.5005
R13228 CSoutput.n150 CSoutput.n141 4.5005
R13229 CSoutput.n150 CSoutput.n143 4.5005
R13230 CSoutput.n150 CSoutput.n140 4.5005
R13231 CSoutput.n150 CSoutput.n144 4.5005
R13232 CSoutput.n150 CSoutput.n139 4.5005
R13233 CSoutput.n150 CSoutput.t102 4.5005
R13234 CSoutput.n150 CSoutput.n138 4.5005
R13235 CSoutput.n150 CSoutput.n145 4.5005
R13236 CSoutput.n150 CSoutput.n146 4.5005
R13237 CSoutput.n242 CSoutput.n141 4.5005
R13238 CSoutput.n242 CSoutput.n143 4.5005
R13239 CSoutput.n242 CSoutput.n140 4.5005
R13240 CSoutput.n242 CSoutput.n144 4.5005
R13241 CSoutput.n242 CSoutput.n139 4.5005
R13242 CSoutput.n242 CSoutput.t102 4.5005
R13243 CSoutput.n242 CSoutput.n138 4.5005
R13244 CSoutput.n242 CSoutput.n145 4.5005
R13245 CSoutput.n242 CSoutput.n146 4.5005
R13246 CSoutput.n229 CSoutput.n200 4.5005
R13247 CSoutput.n229 CSoutput.n206 4.5005
R13248 CSoutput.n187 CSoutput.n176 4.5005
R13249 CSoutput.n187 CSoutput.n178 4.5005
R13250 CSoutput.n187 CSoutput.n175 4.5005
R13251 CSoutput.n187 CSoutput.n179 4.5005
R13252 CSoutput.n187 CSoutput.n174 4.5005
R13253 CSoutput.n187 CSoutput.t98 4.5005
R13254 CSoutput.n187 CSoutput.n173 4.5005
R13255 CSoutput.n187 CSoutput.n180 4.5005
R13256 CSoutput.n229 CSoutput.n187 4.5005
R13257 CSoutput.n208 CSoutput.n176 4.5005
R13258 CSoutput.n208 CSoutput.n178 4.5005
R13259 CSoutput.n208 CSoutput.n175 4.5005
R13260 CSoutput.n208 CSoutput.n179 4.5005
R13261 CSoutput.n208 CSoutput.n174 4.5005
R13262 CSoutput.n208 CSoutput.t98 4.5005
R13263 CSoutput.n208 CSoutput.n173 4.5005
R13264 CSoutput.n208 CSoutput.n180 4.5005
R13265 CSoutput.n229 CSoutput.n208 4.5005
R13266 CSoutput.n186 CSoutput.n176 4.5005
R13267 CSoutput.n186 CSoutput.n178 4.5005
R13268 CSoutput.n186 CSoutput.n175 4.5005
R13269 CSoutput.n186 CSoutput.n179 4.5005
R13270 CSoutput.n186 CSoutput.n174 4.5005
R13271 CSoutput.n186 CSoutput.t98 4.5005
R13272 CSoutput.n186 CSoutput.n173 4.5005
R13273 CSoutput.n186 CSoutput.n180 4.5005
R13274 CSoutput.n229 CSoutput.n186 4.5005
R13275 CSoutput.n210 CSoutput.n176 4.5005
R13276 CSoutput.n210 CSoutput.n178 4.5005
R13277 CSoutput.n210 CSoutput.n175 4.5005
R13278 CSoutput.n210 CSoutput.n179 4.5005
R13279 CSoutput.n210 CSoutput.n174 4.5005
R13280 CSoutput.n210 CSoutput.t98 4.5005
R13281 CSoutput.n210 CSoutput.n173 4.5005
R13282 CSoutput.n210 CSoutput.n180 4.5005
R13283 CSoutput.n229 CSoutput.n210 4.5005
R13284 CSoutput.n176 CSoutput.n171 4.5005
R13285 CSoutput.n178 CSoutput.n171 4.5005
R13286 CSoutput.n175 CSoutput.n171 4.5005
R13287 CSoutput.n179 CSoutput.n171 4.5005
R13288 CSoutput.n174 CSoutput.n171 4.5005
R13289 CSoutput.t98 CSoutput.n171 4.5005
R13290 CSoutput.n173 CSoutput.n171 4.5005
R13291 CSoutput.n180 CSoutput.n171 4.5005
R13292 CSoutput.n232 CSoutput.n176 4.5005
R13293 CSoutput.n232 CSoutput.n178 4.5005
R13294 CSoutput.n232 CSoutput.n175 4.5005
R13295 CSoutput.n232 CSoutput.n179 4.5005
R13296 CSoutput.n232 CSoutput.n174 4.5005
R13297 CSoutput.n232 CSoutput.t98 4.5005
R13298 CSoutput.n232 CSoutput.n173 4.5005
R13299 CSoutput.n232 CSoutput.n180 4.5005
R13300 CSoutput.n230 CSoutput.n176 4.5005
R13301 CSoutput.n230 CSoutput.n178 4.5005
R13302 CSoutput.n230 CSoutput.n175 4.5005
R13303 CSoutput.n230 CSoutput.n179 4.5005
R13304 CSoutput.n230 CSoutput.n174 4.5005
R13305 CSoutput.n230 CSoutput.t98 4.5005
R13306 CSoutput.n230 CSoutput.n173 4.5005
R13307 CSoutput.n230 CSoutput.n180 4.5005
R13308 CSoutput.n230 CSoutput.n229 4.5005
R13309 CSoutput.n212 CSoutput.n176 4.5005
R13310 CSoutput.n212 CSoutput.n178 4.5005
R13311 CSoutput.n212 CSoutput.n175 4.5005
R13312 CSoutput.n212 CSoutput.n179 4.5005
R13313 CSoutput.n212 CSoutput.n174 4.5005
R13314 CSoutput.n212 CSoutput.t98 4.5005
R13315 CSoutput.n212 CSoutput.n173 4.5005
R13316 CSoutput.n212 CSoutput.n180 4.5005
R13317 CSoutput.n229 CSoutput.n212 4.5005
R13318 CSoutput.n184 CSoutput.n176 4.5005
R13319 CSoutput.n184 CSoutput.n178 4.5005
R13320 CSoutput.n184 CSoutput.n175 4.5005
R13321 CSoutput.n184 CSoutput.n179 4.5005
R13322 CSoutput.n184 CSoutput.n174 4.5005
R13323 CSoutput.n184 CSoutput.t98 4.5005
R13324 CSoutput.n184 CSoutput.n173 4.5005
R13325 CSoutput.n184 CSoutput.n180 4.5005
R13326 CSoutput.n229 CSoutput.n184 4.5005
R13327 CSoutput.n214 CSoutput.n176 4.5005
R13328 CSoutput.n214 CSoutput.n178 4.5005
R13329 CSoutput.n214 CSoutput.n175 4.5005
R13330 CSoutput.n214 CSoutput.n179 4.5005
R13331 CSoutput.n214 CSoutput.n174 4.5005
R13332 CSoutput.n214 CSoutput.t98 4.5005
R13333 CSoutput.n214 CSoutput.n173 4.5005
R13334 CSoutput.n214 CSoutput.n180 4.5005
R13335 CSoutput.n229 CSoutput.n214 4.5005
R13336 CSoutput.n183 CSoutput.n176 4.5005
R13337 CSoutput.n183 CSoutput.n178 4.5005
R13338 CSoutput.n183 CSoutput.n175 4.5005
R13339 CSoutput.n183 CSoutput.n179 4.5005
R13340 CSoutput.n183 CSoutput.n174 4.5005
R13341 CSoutput.n183 CSoutput.t98 4.5005
R13342 CSoutput.n183 CSoutput.n173 4.5005
R13343 CSoutput.n183 CSoutput.n180 4.5005
R13344 CSoutput.n229 CSoutput.n183 4.5005
R13345 CSoutput.n228 CSoutput.n176 4.5005
R13346 CSoutput.n228 CSoutput.n178 4.5005
R13347 CSoutput.n228 CSoutput.n175 4.5005
R13348 CSoutput.n228 CSoutput.n179 4.5005
R13349 CSoutput.n228 CSoutput.n174 4.5005
R13350 CSoutput.n228 CSoutput.t98 4.5005
R13351 CSoutput.n228 CSoutput.n173 4.5005
R13352 CSoutput.n228 CSoutput.n180 4.5005
R13353 CSoutput.n229 CSoutput.n228 4.5005
R13354 CSoutput.n227 CSoutput.n112 4.5005
R13355 CSoutput.n128 CSoutput.n112 4.5005
R13356 CSoutput.n123 CSoutput.n107 4.5005
R13357 CSoutput.n123 CSoutput.n109 4.5005
R13358 CSoutput.n123 CSoutput.n106 4.5005
R13359 CSoutput.n123 CSoutput.n110 4.5005
R13360 CSoutput.n123 CSoutput.n105 4.5005
R13361 CSoutput.n123 CSoutput.t115 4.5005
R13362 CSoutput.n123 CSoutput.n104 4.5005
R13363 CSoutput.n123 CSoutput.n111 4.5005
R13364 CSoutput.n123 CSoutput.n112 4.5005
R13365 CSoutput.n121 CSoutput.n107 4.5005
R13366 CSoutput.n121 CSoutput.n109 4.5005
R13367 CSoutput.n121 CSoutput.n106 4.5005
R13368 CSoutput.n121 CSoutput.n110 4.5005
R13369 CSoutput.n121 CSoutput.n105 4.5005
R13370 CSoutput.n121 CSoutput.t115 4.5005
R13371 CSoutput.n121 CSoutput.n104 4.5005
R13372 CSoutput.n121 CSoutput.n111 4.5005
R13373 CSoutput.n121 CSoutput.n112 4.5005
R13374 CSoutput.n120 CSoutput.n107 4.5005
R13375 CSoutput.n120 CSoutput.n109 4.5005
R13376 CSoutput.n120 CSoutput.n106 4.5005
R13377 CSoutput.n120 CSoutput.n110 4.5005
R13378 CSoutput.n120 CSoutput.n105 4.5005
R13379 CSoutput.n120 CSoutput.t115 4.5005
R13380 CSoutput.n120 CSoutput.n104 4.5005
R13381 CSoutput.n120 CSoutput.n111 4.5005
R13382 CSoutput.n120 CSoutput.n112 4.5005
R13383 CSoutput.n249 CSoutput.n107 4.5005
R13384 CSoutput.n249 CSoutput.n109 4.5005
R13385 CSoutput.n249 CSoutput.n106 4.5005
R13386 CSoutput.n249 CSoutput.n110 4.5005
R13387 CSoutput.n249 CSoutput.n105 4.5005
R13388 CSoutput.n249 CSoutput.t115 4.5005
R13389 CSoutput.n249 CSoutput.n104 4.5005
R13390 CSoutput.n249 CSoutput.n111 4.5005
R13391 CSoutput.n249 CSoutput.n112 4.5005
R13392 CSoutput.n247 CSoutput.n107 4.5005
R13393 CSoutput.n247 CSoutput.n109 4.5005
R13394 CSoutput.n247 CSoutput.n106 4.5005
R13395 CSoutput.n247 CSoutput.n110 4.5005
R13396 CSoutput.n247 CSoutput.n105 4.5005
R13397 CSoutput.n247 CSoutput.t115 4.5005
R13398 CSoutput.n247 CSoutput.n104 4.5005
R13399 CSoutput.n247 CSoutput.n111 4.5005
R13400 CSoutput.n245 CSoutput.n107 4.5005
R13401 CSoutput.n245 CSoutput.n109 4.5005
R13402 CSoutput.n245 CSoutput.n106 4.5005
R13403 CSoutput.n245 CSoutput.n110 4.5005
R13404 CSoutput.n245 CSoutput.n105 4.5005
R13405 CSoutput.n245 CSoutput.t115 4.5005
R13406 CSoutput.n245 CSoutput.n104 4.5005
R13407 CSoutput.n245 CSoutput.n111 4.5005
R13408 CSoutput.n131 CSoutput.n107 4.5005
R13409 CSoutput.n131 CSoutput.n109 4.5005
R13410 CSoutput.n131 CSoutput.n106 4.5005
R13411 CSoutput.n131 CSoutput.n110 4.5005
R13412 CSoutput.n131 CSoutput.n105 4.5005
R13413 CSoutput.n131 CSoutput.t115 4.5005
R13414 CSoutput.n131 CSoutput.n104 4.5005
R13415 CSoutput.n131 CSoutput.n111 4.5005
R13416 CSoutput.n131 CSoutput.n112 4.5005
R13417 CSoutput.n130 CSoutput.n107 4.5005
R13418 CSoutput.n130 CSoutput.n109 4.5005
R13419 CSoutput.n130 CSoutput.n106 4.5005
R13420 CSoutput.n130 CSoutput.n110 4.5005
R13421 CSoutput.n130 CSoutput.n105 4.5005
R13422 CSoutput.n130 CSoutput.t115 4.5005
R13423 CSoutput.n130 CSoutput.n104 4.5005
R13424 CSoutput.n130 CSoutput.n111 4.5005
R13425 CSoutput.n130 CSoutput.n112 4.5005
R13426 CSoutput.n134 CSoutput.n107 4.5005
R13427 CSoutput.n134 CSoutput.n109 4.5005
R13428 CSoutput.n134 CSoutput.n106 4.5005
R13429 CSoutput.n134 CSoutput.n110 4.5005
R13430 CSoutput.n134 CSoutput.n105 4.5005
R13431 CSoutput.n134 CSoutput.t115 4.5005
R13432 CSoutput.n134 CSoutput.n104 4.5005
R13433 CSoutput.n134 CSoutput.n111 4.5005
R13434 CSoutput.n134 CSoutput.n112 4.5005
R13435 CSoutput.n133 CSoutput.n107 4.5005
R13436 CSoutput.n133 CSoutput.n109 4.5005
R13437 CSoutput.n133 CSoutput.n106 4.5005
R13438 CSoutput.n133 CSoutput.n110 4.5005
R13439 CSoutput.n133 CSoutput.n105 4.5005
R13440 CSoutput.n133 CSoutput.t115 4.5005
R13441 CSoutput.n133 CSoutput.n104 4.5005
R13442 CSoutput.n133 CSoutput.n111 4.5005
R13443 CSoutput.n133 CSoutput.n112 4.5005
R13444 CSoutput.n116 CSoutput.n107 4.5005
R13445 CSoutput.n116 CSoutput.n109 4.5005
R13446 CSoutput.n116 CSoutput.n106 4.5005
R13447 CSoutput.n116 CSoutput.n110 4.5005
R13448 CSoutput.n116 CSoutput.n105 4.5005
R13449 CSoutput.n116 CSoutput.t115 4.5005
R13450 CSoutput.n116 CSoutput.n104 4.5005
R13451 CSoutput.n116 CSoutput.n111 4.5005
R13452 CSoutput.n116 CSoutput.n112 4.5005
R13453 CSoutput.n252 CSoutput.n107 4.5005
R13454 CSoutput.n252 CSoutput.n109 4.5005
R13455 CSoutput.n252 CSoutput.n106 4.5005
R13456 CSoutput.n252 CSoutput.n110 4.5005
R13457 CSoutput.n252 CSoutput.n105 4.5005
R13458 CSoutput.n252 CSoutput.t115 4.5005
R13459 CSoutput.n252 CSoutput.n104 4.5005
R13460 CSoutput.n252 CSoutput.n111 4.5005
R13461 CSoutput.n252 CSoutput.n112 4.5005
R13462 CSoutput.n275 CSoutput.n267 4.10845
R13463 CSoutput.n101 CSoutput.n93 4.10845
R13464 CSoutput.n273 CSoutput.t78 4.06363
R13465 CSoutput.n273 CSoutput.t7 4.06363
R13466 CSoutput.n271 CSoutput.t81 4.06363
R13467 CSoutput.n271 CSoutput.t3 4.06363
R13468 CSoutput.n269 CSoutput.t75 4.06363
R13469 CSoutput.n269 CSoutput.t16 4.06363
R13470 CSoutput.n268 CSoutput.t13 4.06363
R13471 CSoutput.n268 CSoutput.t15 4.06363
R13472 CSoutput.n265 CSoutput.t1 4.06363
R13473 CSoutput.n265 CSoutput.t4 4.06363
R13474 CSoutput.n263 CSoutput.t70 4.06363
R13475 CSoutput.n263 CSoutput.t95 4.06363
R13476 CSoutput.n261 CSoutput.t86 4.06363
R13477 CSoutput.n261 CSoutput.t19 4.06363
R13478 CSoutput.n260 CSoutput.t18 4.06363
R13479 CSoutput.n260 CSoutput.t91 4.06363
R13480 CSoutput.n258 CSoutput.t71 4.06363
R13481 CSoutput.n258 CSoutput.t68 4.06363
R13482 CSoutput.n256 CSoutput.t8 4.06363
R13483 CSoutput.n256 CSoutput.t74 4.06363
R13484 CSoutput.n254 CSoutput.t12 4.06363
R13485 CSoutput.n254 CSoutput.t90 4.06363
R13486 CSoutput.n253 CSoutput.t89 4.06363
R13487 CSoutput.n253 CSoutput.t6 4.06363
R13488 CSoutput.n94 CSoutput.t0 4.06363
R13489 CSoutput.n94 CSoutput.t14 4.06363
R13490 CSoutput.n95 CSoutput.t11 4.06363
R13491 CSoutput.n95 CSoutput.t17 4.06363
R13492 CSoutput.n97 CSoutput.t2 4.06363
R13493 CSoutput.n97 CSoutput.t94 4.06363
R13494 CSoutput.n99 CSoutput.t87 4.06363
R13495 CSoutput.n99 CSoutput.t92 4.06363
R13496 CSoutput.n86 CSoutput.t76 4.06363
R13497 CSoutput.n86 CSoutput.t9 4.06363
R13498 CSoutput.n87 CSoutput.t73 4.06363
R13499 CSoutput.n87 CSoutput.t88 4.06363
R13500 CSoutput.n89 CSoutput.t83 4.06363
R13501 CSoutput.n89 CSoutput.t79 4.06363
R13502 CSoutput.n91 CSoutput.t5 4.06363
R13503 CSoutput.n91 CSoutput.t69 4.06363
R13504 CSoutput.n79 CSoutput.t84 4.06363
R13505 CSoutput.n79 CSoutput.t93 4.06363
R13506 CSoutput.n80 CSoutput.t77 4.06363
R13507 CSoutput.n80 CSoutput.t82 4.06363
R13508 CSoutput.n82 CSoutput.t72 4.06363
R13509 CSoutput.n82 CSoutput.t85 4.06363
R13510 CSoutput.n84 CSoutput.t10 4.06363
R13511 CSoutput.n84 CSoutput.t80 4.06363
R13512 CSoutput.n44 CSoutput.n43 3.79402
R13513 CSoutput.n49 CSoutput.n48 3.79402
R13514 CSoutput.n325 CSoutput.n324 3.57343
R13515 CSoutput.n297 CSoutput.t58 2.82907
R13516 CSoutput.n297 CSoutput.t61 2.82907
R13517 CSoutput.n295 CSoutput.t57 2.82907
R13518 CSoutput.n295 CSoutput.t47 2.82907
R13519 CSoutput.n293 CSoutput.t24 2.82907
R13520 CSoutput.n293 CSoutput.t55 2.82907
R13521 CSoutput.n291 CSoutput.t49 2.82907
R13522 CSoutput.n291 CSoutput.t38 2.82907
R13523 CSoutput.n289 CSoutput.t66 2.82907
R13524 CSoutput.n289 CSoutput.t20 2.82907
R13525 CSoutput.n288 CSoutput.t54 2.82907
R13526 CSoutput.n288 CSoutput.t43 2.82907
R13527 CSoutput.n286 CSoutput.t51 2.82907
R13528 CSoutput.n286 CSoutput.t53 2.82907
R13529 CSoutput.n284 CSoutput.t48 2.82907
R13530 CSoutput.n284 CSoutput.t37 2.82907
R13531 CSoutput.n282 CSoutput.t65 2.82907
R13532 CSoutput.n282 CSoutput.t46 2.82907
R13533 CSoutput.n280 CSoutput.t39 2.82907
R13534 CSoutput.n280 CSoutput.t29 2.82907
R13535 CSoutput.n278 CSoutput.t60 2.82907
R13536 CSoutput.n278 CSoutput.t62 2.82907
R13537 CSoutput.n277 CSoutput.t44 2.82907
R13538 CSoutput.n277 CSoutput.t34 2.82907
R13539 CSoutput.n312 CSoutput.t30 2.82907
R13540 CSoutput.n312 CSoutput.t42 2.82907
R13541 CSoutput.n313 CSoutput.t59 2.82907
R13542 CSoutput.n313 CSoutput.t22 2.82907
R13543 CSoutput.n315 CSoutput.t26 2.82907
R13544 CSoutput.n315 CSoutput.t36 2.82907
R13545 CSoutput.n317 CSoutput.t41 2.82907
R13546 CSoutput.n317 CSoutput.t28 2.82907
R13547 CSoutput.n319 CSoutput.t33 2.82907
R13548 CSoutput.n319 CSoutput.t45 2.82907
R13549 CSoutput.n321 CSoutput.t50 2.82907
R13550 CSoutput.n321 CSoutput.t63 2.82907
R13551 CSoutput.n301 CSoutput.t23 2.82907
R13552 CSoutput.n301 CSoutput.t31 2.82907
R13553 CSoutput.n302 CSoutput.t52 2.82907
R13554 CSoutput.n302 CSoutput.t64 2.82907
R13555 CSoutput.n304 CSoutput.t67 2.82907
R13556 CSoutput.n304 CSoutput.t27 2.82907
R13557 CSoutput.n306 CSoutput.t32 2.82907
R13558 CSoutput.n306 CSoutput.t21 2.82907
R13559 CSoutput.n308 CSoutput.t25 2.82907
R13560 CSoutput.n308 CSoutput.t35 2.82907
R13561 CSoutput.n310 CSoutput.t40 2.82907
R13562 CSoutput.n310 CSoutput.t56 2.82907
R13563 CSoutput.n324 CSoutput.n300 2.75627
R13564 CSoutput.n75 CSoutput.n1 2.45513
R13565 CSoutput.n193 CSoutput.n191 2.251
R13566 CSoutput.n193 CSoutput.n190 2.251
R13567 CSoutput.n193 CSoutput.n189 2.251
R13568 CSoutput.n193 CSoutput.n188 2.251
R13569 CSoutput.n162 CSoutput.n161 2.251
R13570 CSoutput.n162 CSoutput.n160 2.251
R13571 CSoutput.n162 CSoutput.n159 2.251
R13572 CSoutput.n162 CSoutput.n158 2.251
R13573 CSoutput.n235 CSoutput.n234 2.251
R13574 CSoutput.n200 CSoutput.n198 2.251
R13575 CSoutput.n200 CSoutput.n197 2.251
R13576 CSoutput.n200 CSoutput.n196 2.251
R13577 CSoutput.n218 CSoutput.n200 2.251
R13578 CSoutput.n206 CSoutput.n205 2.251
R13579 CSoutput.n206 CSoutput.n204 2.251
R13580 CSoutput.n206 CSoutput.n203 2.251
R13581 CSoutput.n206 CSoutput.n202 2.251
R13582 CSoutput.n232 CSoutput.n172 2.251
R13583 CSoutput.n227 CSoutput.n225 2.251
R13584 CSoutput.n227 CSoutput.n224 2.251
R13585 CSoutput.n227 CSoutput.n223 2.251
R13586 CSoutput.n227 CSoutput.n222 2.251
R13587 CSoutput.n128 CSoutput.n127 2.251
R13588 CSoutput.n128 CSoutput.n126 2.251
R13589 CSoutput.n128 CSoutput.n125 2.251
R13590 CSoutput.n128 CSoutput.n124 2.251
R13591 CSoutput.n245 CSoutput.n244 2.251
R13592 CSoutput.n162 CSoutput.n142 2.2505
R13593 CSoutput.n157 CSoutput.n142 2.2505
R13594 CSoutput.n155 CSoutput.n142 2.2505
R13595 CSoutput.n154 CSoutput.n142 2.2505
R13596 CSoutput.n239 CSoutput.n142 2.2505
R13597 CSoutput.n237 CSoutput.n142 2.2505
R13598 CSoutput.n235 CSoutput.n142 2.2505
R13599 CSoutput.n165 CSoutput.n142 2.2505
R13600 CSoutput.n164 CSoutput.n142 2.2505
R13601 CSoutput.n168 CSoutput.n142 2.2505
R13602 CSoutput.n167 CSoutput.n142 2.2505
R13603 CSoutput.n150 CSoutput.n142 2.2505
R13604 CSoutput.n242 CSoutput.n142 2.2505
R13605 CSoutput.n242 CSoutput.n241 2.2505
R13606 CSoutput.n206 CSoutput.n177 2.2505
R13607 CSoutput.n187 CSoutput.n177 2.2505
R13608 CSoutput.n208 CSoutput.n177 2.2505
R13609 CSoutput.n186 CSoutput.n177 2.2505
R13610 CSoutput.n210 CSoutput.n177 2.2505
R13611 CSoutput.n177 CSoutput.n171 2.2505
R13612 CSoutput.n232 CSoutput.n177 2.2505
R13613 CSoutput.n230 CSoutput.n177 2.2505
R13614 CSoutput.n212 CSoutput.n177 2.2505
R13615 CSoutput.n184 CSoutput.n177 2.2505
R13616 CSoutput.n214 CSoutput.n177 2.2505
R13617 CSoutput.n183 CSoutput.n177 2.2505
R13618 CSoutput.n228 CSoutput.n177 2.2505
R13619 CSoutput.n228 CSoutput.n181 2.2505
R13620 CSoutput.n128 CSoutput.n108 2.2505
R13621 CSoutput.n123 CSoutput.n108 2.2505
R13622 CSoutput.n121 CSoutput.n108 2.2505
R13623 CSoutput.n120 CSoutput.n108 2.2505
R13624 CSoutput.n249 CSoutput.n108 2.2505
R13625 CSoutput.n247 CSoutput.n108 2.2505
R13626 CSoutput.n245 CSoutput.n108 2.2505
R13627 CSoutput.n131 CSoutput.n108 2.2505
R13628 CSoutput.n130 CSoutput.n108 2.2505
R13629 CSoutput.n134 CSoutput.n108 2.2505
R13630 CSoutput.n133 CSoutput.n108 2.2505
R13631 CSoutput.n116 CSoutput.n108 2.2505
R13632 CSoutput.n252 CSoutput.n108 2.2505
R13633 CSoutput.n252 CSoutput.n251 2.2505
R13634 CSoutput.n170 CSoutput.n163 2.25024
R13635 CSoutput.n170 CSoutput.n156 2.25024
R13636 CSoutput.n238 CSoutput.n170 2.25024
R13637 CSoutput.n170 CSoutput.n166 2.25024
R13638 CSoutput.n170 CSoutput.n169 2.25024
R13639 CSoutput.n170 CSoutput.n137 2.25024
R13640 CSoutput.n220 CSoutput.n217 2.25024
R13641 CSoutput.n220 CSoutput.n216 2.25024
R13642 CSoutput.n220 CSoutput.n215 2.25024
R13643 CSoutput.n220 CSoutput.n182 2.25024
R13644 CSoutput.n220 CSoutput.n219 2.25024
R13645 CSoutput.n221 CSoutput.n220 2.25024
R13646 CSoutput.n136 CSoutput.n129 2.25024
R13647 CSoutput.n136 CSoutput.n122 2.25024
R13648 CSoutput.n248 CSoutput.n136 2.25024
R13649 CSoutput.n136 CSoutput.n132 2.25024
R13650 CSoutput.n136 CSoutput.n135 2.25024
R13651 CSoutput.n136 CSoutput.n103 2.25024
R13652 CSoutput.n276 CSoutput.n102 1.95131
R13653 CSoutput.n237 CSoutput.n147 1.50111
R13654 CSoutput.n185 CSoutput.n171 1.50111
R13655 CSoutput.n247 CSoutput.n113 1.50111
R13656 CSoutput.n193 CSoutput.n192 1.501
R13657 CSoutput.n200 CSoutput.n199 1.501
R13658 CSoutput.n227 CSoutput.n226 1.501
R13659 CSoutput.n241 CSoutput.n152 1.12536
R13660 CSoutput.n241 CSoutput.n153 1.12536
R13661 CSoutput.n241 CSoutput.n240 1.12536
R13662 CSoutput.n201 CSoutput.n181 1.12536
R13663 CSoutput.n207 CSoutput.n181 1.12536
R13664 CSoutput.n209 CSoutput.n181 1.12536
R13665 CSoutput.n251 CSoutput.n118 1.12536
R13666 CSoutput.n251 CSoutput.n119 1.12536
R13667 CSoutput.n251 CSoutput.n250 1.12536
R13668 CSoutput.n241 CSoutput.n148 1.12536
R13669 CSoutput.n241 CSoutput.n149 1.12536
R13670 CSoutput.n241 CSoutput.n151 1.12536
R13671 CSoutput.n231 CSoutput.n181 1.12536
R13672 CSoutput.n211 CSoutput.n181 1.12536
R13673 CSoutput.n213 CSoutput.n181 1.12536
R13674 CSoutput.n251 CSoutput.n114 1.12536
R13675 CSoutput.n251 CSoutput.n115 1.12536
R13676 CSoutput.n251 CSoutput.n117 1.12536
R13677 CSoutput.n31 CSoutput.n30 0.669944
R13678 CSoutput.n62 CSoutput.n61 0.669944
R13679 CSoutput.n292 CSoutput.n290 0.573776
R13680 CSoutput.n294 CSoutput.n292 0.573776
R13681 CSoutput.n296 CSoutput.n294 0.573776
R13682 CSoutput.n298 CSoutput.n296 0.573776
R13683 CSoutput.n281 CSoutput.n279 0.573776
R13684 CSoutput.n283 CSoutput.n281 0.573776
R13685 CSoutput.n285 CSoutput.n283 0.573776
R13686 CSoutput.n287 CSoutput.n285 0.573776
R13687 CSoutput.n322 CSoutput.n320 0.573776
R13688 CSoutput.n320 CSoutput.n318 0.573776
R13689 CSoutput.n318 CSoutput.n316 0.573776
R13690 CSoutput.n316 CSoutput.n314 0.573776
R13691 CSoutput.n311 CSoutput.n309 0.573776
R13692 CSoutput.n309 CSoutput.n307 0.573776
R13693 CSoutput.n307 CSoutput.n305 0.573776
R13694 CSoutput.n305 CSoutput.n303 0.573776
R13695 CSoutput.n325 CSoutput.n252 0.53442
R13696 CSoutput.n272 CSoutput.n270 0.358259
R13697 CSoutput.n274 CSoutput.n272 0.358259
R13698 CSoutput.n264 CSoutput.n262 0.358259
R13699 CSoutput.n266 CSoutput.n264 0.358259
R13700 CSoutput.n257 CSoutput.n255 0.358259
R13701 CSoutput.n259 CSoutput.n257 0.358259
R13702 CSoutput.n100 CSoutput.n98 0.358259
R13703 CSoutput.n98 CSoutput.n96 0.358259
R13704 CSoutput.n92 CSoutput.n90 0.358259
R13705 CSoutput.n90 CSoutput.n88 0.358259
R13706 CSoutput.n85 CSoutput.n83 0.358259
R13707 CSoutput.n83 CSoutput.n81 0.358259
R13708 CSoutput.n21 CSoutput.n20 0.169105
R13709 CSoutput.n21 CSoutput.n16 0.169105
R13710 CSoutput.n26 CSoutput.n16 0.169105
R13711 CSoutput.n27 CSoutput.n26 0.169105
R13712 CSoutput.n27 CSoutput.n14 0.169105
R13713 CSoutput.n32 CSoutput.n14 0.169105
R13714 CSoutput.n33 CSoutput.n32 0.169105
R13715 CSoutput.n34 CSoutput.n33 0.169105
R13716 CSoutput.n34 CSoutput.n12 0.169105
R13717 CSoutput.n39 CSoutput.n12 0.169105
R13718 CSoutput.n40 CSoutput.n39 0.169105
R13719 CSoutput.n40 CSoutput.n10 0.169105
R13720 CSoutput.n45 CSoutput.n10 0.169105
R13721 CSoutput.n46 CSoutput.n45 0.169105
R13722 CSoutput.n47 CSoutput.n46 0.169105
R13723 CSoutput.n47 CSoutput.n8 0.169105
R13724 CSoutput.n52 CSoutput.n8 0.169105
R13725 CSoutput.n53 CSoutput.n52 0.169105
R13726 CSoutput.n53 CSoutput.n6 0.169105
R13727 CSoutput.n58 CSoutput.n6 0.169105
R13728 CSoutput.n59 CSoutput.n58 0.169105
R13729 CSoutput.n60 CSoutput.n59 0.169105
R13730 CSoutput.n60 CSoutput.n4 0.169105
R13731 CSoutput.n66 CSoutput.n4 0.169105
R13732 CSoutput.n67 CSoutput.n66 0.169105
R13733 CSoutput.n68 CSoutput.n67 0.169105
R13734 CSoutput.n68 CSoutput.n2 0.169105
R13735 CSoutput.n73 CSoutput.n2 0.169105
R13736 CSoutput.n74 CSoutput.n73 0.169105
R13737 CSoutput.n74 CSoutput.n0 0.169105
R13738 CSoutput.n78 CSoutput.n0 0.169105
R13739 CSoutput.n195 CSoutput.n194 0.0910737
R13740 CSoutput.n246 CSoutput.n243 0.0723685
R13741 CSoutput.n200 CSoutput.n195 0.0522944
R13742 CSoutput.n243 CSoutput.n242 0.0499135
R13743 CSoutput.n194 CSoutput.n193 0.0499135
R13744 CSoutput.n228 CSoutput.n227 0.0464294
R13745 CSoutput.n236 CSoutput.n233 0.0391444
R13746 CSoutput.n195 CSoutput.t105 0.023435
R13747 CSoutput.n243 CSoutput.t104 0.02262
R13748 CSoutput.n194 CSoutput.t109 0.02262
R13749 CSoutput CSoutput.n325 0.0052
R13750 CSoutput.n165 CSoutput.n148 0.00365111
R13751 CSoutput.n168 CSoutput.n149 0.00365111
R13752 CSoutput.n151 CSoutput.n150 0.00365111
R13753 CSoutput.n193 CSoutput.n152 0.00365111
R13754 CSoutput.n157 CSoutput.n153 0.00365111
R13755 CSoutput.n240 CSoutput.n154 0.00365111
R13756 CSoutput.n231 CSoutput.n230 0.00365111
R13757 CSoutput.n211 CSoutput.n184 0.00365111
R13758 CSoutput.n213 CSoutput.n183 0.00365111
R13759 CSoutput.n201 CSoutput.n200 0.00365111
R13760 CSoutput.n207 CSoutput.n187 0.00365111
R13761 CSoutput.n209 CSoutput.n186 0.00365111
R13762 CSoutput.n131 CSoutput.n114 0.00365111
R13763 CSoutput.n134 CSoutput.n115 0.00365111
R13764 CSoutput.n117 CSoutput.n116 0.00365111
R13765 CSoutput.n227 CSoutput.n118 0.00365111
R13766 CSoutput.n123 CSoutput.n119 0.00365111
R13767 CSoutput.n250 CSoutput.n120 0.00365111
R13768 CSoutput.n162 CSoutput.n152 0.00340054
R13769 CSoutput.n155 CSoutput.n153 0.00340054
R13770 CSoutput.n240 CSoutput.n239 0.00340054
R13771 CSoutput.n235 CSoutput.n148 0.00340054
R13772 CSoutput.n164 CSoutput.n149 0.00340054
R13773 CSoutput.n167 CSoutput.n151 0.00340054
R13774 CSoutput.n206 CSoutput.n201 0.00340054
R13775 CSoutput.n208 CSoutput.n207 0.00340054
R13776 CSoutput.n210 CSoutput.n209 0.00340054
R13777 CSoutput.n232 CSoutput.n231 0.00340054
R13778 CSoutput.n212 CSoutput.n211 0.00340054
R13779 CSoutput.n214 CSoutput.n213 0.00340054
R13780 CSoutput.n128 CSoutput.n118 0.00340054
R13781 CSoutput.n121 CSoutput.n119 0.00340054
R13782 CSoutput.n250 CSoutput.n249 0.00340054
R13783 CSoutput.n245 CSoutput.n114 0.00340054
R13784 CSoutput.n130 CSoutput.n115 0.00340054
R13785 CSoutput.n133 CSoutput.n117 0.00340054
R13786 CSoutput.n163 CSoutput.n157 0.00252698
R13787 CSoutput.n156 CSoutput.n154 0.00252698
R13788 CSoutput.n238 CSoutput.n237 0.00252698
R13789 CSoutput.n166 CSoutput.n164 0.00252698
R13790 CSoutput.n169 CSoutput.n167 0.00252698
R13791 CSoutput.n242 CSoutput.n137 0.00252698
R13792 CSoutput.n163 CSoutput.n162 0.00252698
R13793 CSoutput.n156 CSoutput.n155 0.00252698
R13794 CSoutput.n239 CSoutput.n238 0.00252698
R13795 CSoutput.n166 CSoutput.n165 0.00252698
R13796 CSoutput.n169 CSoutput.n168 0.00252698
R13797 CSoutput.n150 CSoutput.n137 0.00252698
R13798 CSoutput.n217 CSoutput.n187 0.00252698
R13799 CSoutput.n216 CSoutput.n186 0.00252698
R13800 CSoutput.n215 CSoutput.n171 0.00252698
R13801 CSoutput.n212 CSoutput.n182 0.00252698
R13802 CSoutput.n219 CSoutput.n214 0.00252698
R13803 CSoutput.n228 CSoutput.n221 0.00252698
R13804 CSoutput.n217 CSoutput.n206 0.00252698
R13805 CSoutput.n216 CSoutput.n208 0.00252698
R13806 CSoutput.n215 CSoutput.n210 0.00252698
R13807 CSoutput.n230 CSoutput.n182 0.00252698
R13808 CSoutput.n219 CSoutput.n184 0.00252698
R13809 CSoutput.n221 CSoutput.n183 0.00252698
R13810 CSoutput.n129 CSoutput.n123 0.00252698
R13811 CSoutput.n122 CSoutput.n120 0.00252698
R13812 CSoutput.n248 CSoutput.n247 0.00252698
R13813 CSoutput.n132 CSoutput.n130 0.00252698
R13814 CSoutput.n135 CSoutput.n133 0.00252698
R13815 CSoutput.n252 CSoutput.n103 0.00252698
R13816 CSoutput.n129 CSoutput.n128 0.00252698
R13817 CSoutput.n122 CSoutput.n121 0.00252698
R13818 CSoutput.n249 CSoutput.n248 0.00252698
R13819 CSoutput.n132 CSoutput.n131 0.00252698
R13820 CSoutput.n135 CSoutput.n134 0.00252698
R13821 CSoutput.n116 CSoutput.n103 0.00252698
R13822 CSoutput.n237 CSoutput.n236 0.0020275
R13823 CSoutput.n236 CSoutput.n235 0.0020275
R13824 CSoutput.n233 CSoutput.n171 0.0020275
R13825 CSoutput.n233 CSoutput.n232 0.0020275
R13826 CSoutput.n247 CSoutput.n246 0.0020275
R13827 CSoutput.n246 CSoutput.n245 0.0020275
R13828 CSoutput.n147 CSoutput.n146 0.00166668
R13829 CSoutput.n229 CSoutput.n185 0.00166668
R13830 CSoutput.n113 CSoutput.n112 0.00166668
R13831 CSoutput.n251 CSoutput.n113 0.00133328
R13832 CSoutput.n185 CSoutput.n181 0.00133328
R13833 CSoutput.n241 CSoutput.n147 0.00133328
R13834 CSoutput.n244 CSoutput.n136 0.001
R13835 CSoutput.n222 CSoutput.n136 0.001
R13836 CSoutput.n124 CSoutput.n104 0.001
R13837 CSoutput.n223 CSoutput.n104 0.001
R13838 CSoutput.n125 CSoutput.n105 0.001
R13839 CSoutput.n224 CSoutput.n105 0.001
R13840 CSoutput.n126 CSoutput.n106 0.001
R13841 CSoutput.n225 CSoutput.n106 0.001
R13842 CSoutput.n127 CSoutput.n107 0.001
R13843 CSoutput.n226 CSoutput.n107 0.001
R13844 CSoutput.n220 CSoutput.n172 0.001
R13845 CSoutput.n220 CSoutput.n218 0.001
R13846 CSoutput.n202 CSoutput.n173 0.001
R13847 CSoutput.n196 CSoutput.n173 0.001
R13848 CSoutput.n203 CSoutput.n174 0.001
R13849 CSoutput.n197 CSoutput.n174 0.001
R13850 CSoutput.n204 CSoutput.n175 0.001
R13851 CSoutput.n198 CSoutput.n175 0.001
R13852 CSoutput.n205 CSoutput.n176 0.001
R13853 CSoutput.n199 CSoutput.n176 0.001
R13854 CSoutput.n234 CSoutput.n170 0.001
R13855 CSoutput.n188 CSoutput.n170 0.001
R13856 CSoutput.n158 CSoutput.n138 0.001
R13857 CSoutput.n189 CSoutput.n138 0.001
R13858 CSoutput.n159 CSoutput.n139 0.001
R13859 CSoutput.n190 CSoutput.n139 0.001
R13860 CSoutput.n160 CSoutput.n140 0.001
R13861 CSoutput.n191 CSoutput.n140 0.001
R13862 CSoutput.n161 CSoutput.n141 0.001
R13863 CSoutput.n192 CSoutput.n141 0.001
R13864 CSoutput.n192 CSoutput.n142 0.001
R13865 CSoutput.n191 CSoutput.n143 0.001
R13866 CSoutput.n190 CSoutput.n144 0.001
R13867 CSoutput.n189 CSoutput.t102 0.001
R13868 CSoutput.n188 CSoutput.n145 0.001
R13869 CSoutput.n161 CSoutput.n143 0.001
R13870 CSoutput.n160 CSoutput.n144 0.001
R13871 CSoutput.n159 CSoutput.t102 0.001
R13872 CSoutput.n158 CSoutput.n145 0.001
R13873 CSoutput.n234 CSoutput.n146 0.001
R13874 CSoutput.n199 CSoutput.n177 0.001
R13875 CSoutput.n198 CSoutput.n178 0.001
R13876 CSoutput.n197 CSoutput.n179 0.001
R13877 CSoutput.n196 CSoutput.t98 0.001
R13878 CSoutput.n218 CSoutput.n180 0.001
R13879 CSoutput.n205 CSoutput.n178 0.001
R13880 CSoutput.n204 CSoutput.n179 0.001
R13881 CSoutput.n203 CSoutput.t98 0.001
R13882 CSoutput.n202 CSoutput.n180 0.001
R13883 CSoutput.n229 CSoutput.n172 0.001
R13884 CSoutput.n226 CSoutput.n108 0.001
R13885 CSoutput.n225 CSoutput.n109 0.001
R13886 CSoutput.n224 CSoutput.n110 0.001
R13887 CSoutput.n223 CSoutput.t115 0.001
R13888 CSoutput.n222 CSoutput.n111 0.001
R13889 CSoutput.n127 CSoutput.n109 0.001
R13890 CSoutput.n126 CSoutput.n110 0.001
R13891 CSoutput.n125 CSoutput.t115 0.001
R13892 CSoutput.n124 CSoutput.n111 0.001
R13893 CSoutput.n244 CSoutput.n112 0.001
R13894 a_n5644_8799.n99 a_n5644_8799.t69 485.149
R13895 a_n5644_8799.n106 a_n5644_8799.t72 485.149
R13896 a_n5644_8799.n114 a_n5644_8799.t38 485.149
R13897 a_n5644_8799.n75 a_n5644_8799.t53 485.149
R13898 a_n5644_8799.n82 a_n5644_8799.t58 485.149
R13899 a_n5644_8799.n90 a_n5644_8799.t39 485.149
R13900 a_n5644_8799.n24 a_n5644_8799.t60 485.135
R13901 a_n5644_8799.n103 a_n5644_8799.t59 464.166
R13902 a_n5644_8799.n97 a_n5644_8799.t46 464.166
R13903 a_n5644_8799.n102 a_n5644_8799.t76 464.166
R13904 a_n5644_8799.n101 a_n5644_8799.t61 464.166
R13905 a_n5644_8799.n98 a_n5644_8799.t51 464.166
R13906 a_n5644_8799.n100 a_n5644_8799.t78 464.166
R13907 a_n5644_8799.n29 a_n5644_8799.t64 485.135
R13908 a_n5644_8799.n110 a_n5644_8799.t63 464.166
R13909 a_n5644_8799.n104 a_n5644_8799.t55 464.166
R13910 a_n5644_8799.n109 a_n5644_8799.t80 464.166
R13911 a_n5644_8799.n108 a_n5644_8799.t67 464.166
R13912 a_n5644_8799.n105 a_n5644_8799.t56 464.166
R13913 a_n5644_8799.n107 a_n5644_8799.t36 464.166
R13914 a_n5644_8799.n34 a_n5644_8799.t82 485.135
R13915 a_n5644_8799.n118 a_n5644_8799.t44 464.166
R13916 a_n5644_8799.n112 a_n5644_8799.t65 464.166
R13917 a_n5644_8799.n117 a_n5644_8799.t37 464.166
R13918 a_n5644_8799.n116 a_n5644_8799.t73 464.166
R13919 a_n5644_8799.n113 a_n5644_8799.t50 464.166
R13920 a_n5644_8799.n115 a_n5644_8799.t70 464.166
R13921 a_n5644_8799.n76 a_n5644_8799.t62 464.166
R13922 a_n5644_8799.n77 a_n5644_8799.t77 464.166
R13923 a_n5644_8799.n78 a_n5644_8799.t42 464.166
R13924 a_n5644_8799.n79 a_n5644_8799.t52 464.166
R13925 a_n5644_8799.n74 a_n5644_8799.t75 464.166
R13926 a_n5644_8799.n80 a_n5644_8799.t41 464.166
R13927 a_n5644_8799.n83 a_n5644_8799.t68 464.166
R13928 a_n5644_8799.n84 a_n5644_8799.t81 464.166
R13929 a_n5644_8799.n85 a_n5644_8799.t49 464.166
R13930 a_n5644_8799.n86 a_n5644_8799.t57 464.166
R13931 a_n5644_8799.n81 a_n5644_8799.t79 464.166
R13932 a_n5644_8799.n87 a_n5644_8799.t45 464.166
R13933 a_n5644_8799.n91 a_n5644_8799.t71 464.166
R13934 a_n5644_8799.n92 a_n5644_8799.t48 464.166
R13935 a_n5644_8799.n93 a_n5644_8799.t74 464.166
R13936 a_n5644_8799.n94 a_n5644_8799.t54 464.166
R13937 a_n5644_8799.n89 a_n5644_8799.t66 464.166
R13938 a_n5644_8799.n95 a_n5644_8799.t43 464.166
R13939 a_n5644_8799.n16 a_n5644_8799.n28 72.3034
R13940 a_n5644_8799.n28 a_n5644_8799.n98 16.6962
R13941 a_n5644_8799.n27 a_n5644_8799.n16 77.6622
R13942 a_n5644_8799.n101 a_n5644_8799.n27 5.97853
R13943 a_n5644_8799.n26 a_n5644_8799.n15 77.6622
R13944 a_n5644_8799.n15 a_n5644_8799.n25 72.3034
R13945 a_n5644_8799.n103 a_n5644_8799.n24 20.9683
R13946 a_n5644_8799.n17 a_n5644_8799.n24 70.1674
R13947 a_n5644_8799.n13 a_n5644_8799.n33 72.3034
R13948 a_n5644_8799.n33 a_n5644_8799.n105 16.6962
R13949 a_n5644_8799.n32 a_n5644_8799.n13 77.6622
R13950 a_n5644_8799.n108 a_n5644_8799.n32 5.97853
R13951 a_n5644_8799.n31 a_n5644_8799.n12 77.6622
R13952 a_n5644_8799.n12 a_n5644_8799.n30 72.3034
R13953 a_n5644_8799.n110 a_n5644_8799.n29 20.9683
R13954 a_n5644_8799.n14 a_n5644_8799.n29 70.1674
R13955 a_n5644_8799.n10 a_n5644_8799.n38 72.3034
R13956 a_n5644_8799.n38 a_n5644_8799.n113 16.6962
R13957 a_n5644_8799.n37 a_n5644_8799.n10 77.6622
R13958 a_n5644_8799.n116 a_n5644_8799.n37 5.97853
R13959 a_n5644_8799.n36 a_n5644_8799.n9 77.6622
R13960 a_n5644_8799.n9 a_n5644_8799.n35 72.3034
R13961 a_n5644_8799.n118 a_n5644_8799.n34 20.9683
R13962 a_n5644_8799.n11 a_n5644_8799.n34 70.1674
R13963 a_n5644_8799.n7 a_n5644_8799.n43 70.1674
R13964 a_n5644_8799.n80 a_n5644_8799.n43 20.9683
R13965 a_n5644_8799.n42 a_n5644_8799.n7 72.3034
R13966 a_n5644_8799.n42 a_n5644_8799.n74 16.6962
R13967 a_n5644_8799.n6 a_n5644_8799.n41 77.6622
R13968 a_n5644_8799.n79 a_n5644_8799.n41 5.97853
R13969 a_n5644_8799.n40 a_n5644_8799.n6 77.6622
R13970 a_n5644_8799.n39 a_n5644_8799.n77 16.6962
R13971 a_n5644_8799.n39 a_n5644_8799.n8 72.3034
R13972 a_n5644_8799.n4 a_n5644_8799.n48 70.1674
R13973 a_n5644_8799.n87 a_n5644_8799.n48 20.9683
R13974 a_n5644_8799.n47 a_n5644_8799.n4 72.3034
R13975 a_n5644_8799.n47 a_n5644_8799.n81 16.6962
R13976 a_n5644_8799.n3 a_n5644_8799.n46 77.6622
R13977 a_n5644_8799.n86 a_n5644_8799.n46 5.97853
R13978 a_n5644_8799.n45 a_n5644_8799.n3 77.6622
R13979 a_n5644_8799.n44 a_n5644_8799.n84 16.6962
R13980 a_n5644_8799.n44 a_n5644_8799.n5 72.3034
R13981 a_n5644_8799.n1 a_n5644_8799.n53 70.1674
R13982 a_n5644_8799.n95 a_n5644_8799.n53 20.9683
R13983 a_n5644_8799.n52 a_n5644_8799.n1 72.3034
R13984 a_n5644_8799.n52 a_n5644_8799.n89 16.6962
R13985 a_n5644_8799.n0 a_n5644_8799.n51 77.6622
R13986 a_n5644_8799.n94 a_n5644_8799.n51 5.97853
R13987 a_n5644_8799.n50 a_n5644_8799.n0 77.6622
R13988 a_n5644_8799.n49 a_n5644_8799.n92 16.6962
R13989 a_n5644_8799.n49 a_n5644_8799.n2 72.3034
R13990 a_n5644_8799.n18 a_n5644_8799.n54 98.9633
R13991 a_n5644_8799.n19 a_n5644_8799.n124 98.9631
R13992 a_n5644_8799.n19 a_n5644_8799.n123 98.6055
R13993 a_n5644_8799.n18 a_n5644_8799.n56 98.6055
R13994 a_n5644_8799.n18 a_n5644_8799.n55 98.6055
R13995 a_n5644_8799.n125 a_n5644_8799.n19 98.6054
R13996 a_n5644_8799.n59 a_n5644_8799.n57 81.4626
R13997 a_n5644_8799.n67 a_n5644_8799.n65 81.4626
R13998 a_n5644_8799.n63 a_n5644_8799.n61 81.4626
R13999 a_n5644_8799.n70 a_n5644_8799.n69 80.9324
R14000 a_n5644_8799.n72 a_n5644_8799.n71 80.9324
R14001 a_n5644_8799.n23 a_n5644_8799.n73 80.9324
R14002 a_n5644_8799.n22 a_n5644_8799.n60 80.9324
R14003 a_n5644_8799.n59 a_n5644_8799.n58 80.9324
R14004 a_n5644_8799.n67 a_n5644_8799.n66 80.9324
R14005 a_n5644_8799.n21 a_n5644_8799.n68 80.9324
R14006 a_n5644_8799.n20 a_n5644_8799.n64 80.9324
R14007 a_n5644_8799.n63 a_n5644_8799.n62 80.9324
R14008 a_n5644_8799.n16 a_n5644_8799.n99 70.4033
R14009 a_n5644_8799.n13 a_n5644_8799.n106 70.4033
R14010 a_n5644_8799.n10 a_n5644_8799.n114 70.4033
R14011 a_n5644_8799.n75 a_n5644_8799.n8 70.4033
R14012 a_n5644_8799.n82 a_n5644_8799.n5 70.4033
R14013 a_n5644_8799.n90 a_n5644_8799.n2 70.4033
R14014 a_n5644_8799.n102 a_n5644_8799.n101 48.2005
R14015 a_n5644_8799.n109 a_n5644_8799.n108 48.2005
R14016 a_n5644_8799.n117 a_n5644_8799.n116 48.2005
R14017 a_n5644_8799.n79 a_n5644_8799.n78 48.2005
R14018 a_n5644_8799.t40 a_n5644_8799.n43 485.135
R14019 a_n5644_8799.n86 a_n5644_8799.n85 48.2005
R14020 a_n5644_8799.t47 a_n5644_8799.n48 485.135
R14021 a_n5644_8799.n94 a_n5644_8799.n93 48.2005
R14022 a_n5644_8799.t83 a_n5644_8799.n53 485.135
R14023 a_n5644_8799.n25 a_n5644_8799.n97 16.6962
R14024 a_n5644_8799.n100 a_n5644_8799.n28 27.6507
R14025 a_n5644_8799.n30 a_n5644_8799.n104 16.6962
R14026 a_n5644_8799.n107 a_n5644_8799.n33 27.6507
R14027 a_n5644_8799.n35 a_n5644_8799.n112 16.6962
R14028 a_n5644_8799.n115 a_n5644_8799.n38 27.6507
R14029 a_n5644_8799.n80 a_n5644_8799.n42 27.6507
R14030 a_n5644_8799.n87 a_n5644_8799.n47 27.6507
R14031 a_n5644_8799.n95 a_n5644_8799.n52 27.6507
R14032 a_n5644_8799.n26 a_n5644_8799.n97 41.7634
R14033 a_n5644_8799.n31 a_n5644_8799.n104 41.7634
R14034 a_n5644_8799.n36 a_n5644_8799.n112 41.7634
R14035 a_n5644_8799.n77 a_n5644_8799.n40 41.7634
R14036 a_n5644_8799.n84 a_n5644_8799.n45 41.7634
R14037 a_n5644_8799.n92 a_n5644_8799.n50 41.7634
R14038 a_n5644_8799.n70 a_n5644_8799.n21 34.3237
R14039 a_n5644_8799.n100 a_n5644_8799.n99 20.9576
R14040 a_n5644_8799.n107 a_n5644_8799.n106 20.9576
R14041 a_n5644_8799.n115 a_n5644_8799.n114 20.9576
R14042 a_n5644_8799.n76 a_n5644_8799.n75 20.9576
R14043 a_n5644_8799.n83 a_n5644_8799.n82 20.9576
R14044 a_n5644_8799.n91 a_n5644_8799.n90 20.9576
R14045 a_n5644_8799.n26 a_n5644_8799.n102 5.97853
R14046 a_n5644_8799.n27 a_n5644_8799.n98 41.7634
R14047 a_n5644_8799.n31 a_n5644_8799.n109 5.97853
R14048 a_n5644_8799.n32 a_n5644_8799.n105 41.7634
R14049 a_n5644_8799.n36 a_n5644_8799.n117 5.97853
R14050 a_n5644_8799.n37 a_n5644_8799.n113 41.7634
R14051 a_n5644_8799.n78 a_n5644_8799.n40 5.97853
R14052 a_n5644_8799.n74 a_n5644_8799.n41 41.7634
R14053 a_n5644_8799.n85 a_n5644_8799.n45 5.97853
R14054 a_n5644_8799.n81 a_n5644_8799.n46 41.7634
R14055 a_n5644_8799.n93 a_n5644_8799.n50 5.97853
R14056 a_n5644_8799.n89 a_n5644_8799.n51 41.7634
R14057 a_n5644_8799.n19 a_n5644_8799.n122 31.5519
R14058 a_n5644_8799.n121 a_n5644_8799.n23 12.3339
R14059 a_n5644_8799.n122 a_n5644_8799.n121 11.4887
R14060 a_n5644_8799.n103 a_n5644_8799.n25 27.6507
R14061 a_n5644_8799.n110 a_n5644_8799.n30 27.6507
R14062 a_n5644_8799.n118 a_n5644_8799.n35 27.6507
R14063 a_n5644_8799.n39 a_n5644_8799.n76 27.6507
R14064 a_n5644_8799.n44 a_n5644_8799.n83 27.6507
R14065 a_n5644_8799.n49 a_n5644_8799.n91 27.6507
R14066 a_n5644_8799.n122 a_n5644_8799.n18 17.6132
R14067 a_n5644_8799.n111 a_n5644_8799.n17 9.05164
R14068 a_n5644_8799.n88 a_n5644_8799.n7 9.05164
R14069 a_n5644_8799.n120 a_n5644_8799.n96 6.93972
R14070 a_n5644_8799.n120 a_n5644_8799.n119 6.44309
R14071 a_n5644_8799.n111 a_n5644_8799.n14 4.94368
R14072 a_n5644_8799.n119 a_n5644_8799.n11 4.94368
R14073 a_n5644_8799.n88 a_n5644_8799.n4 4.94368
R14074 a_n5644_8799.n96 a_n5644_8799.n1 4.94368
R14075 a_n5644_8799.n119 a_n5644_8799.n111 4.10845
R14076 a_n5644_8799.n96 a_n5644_8799.n88 4.10845
R14077 a_n5644_8799.n124 a_n5644_8799.t28 3.61217
R14078 a_n5644_8799.n124 a_n5644_8799.t16 3.61217
R14079 a_n5644_8799.n123 a_n5644_8799.t26 3.61217
R14080 a_n5644_8799.n123 a_n5644_8799.t27 3.61217
R14081 a_n5644_8799.n56 a_n5644_8799.t7 3.61217
R14082 a_n5644_8799.n56 a_n5644_8799.t6 3.61217
R14083 a_n5644_8799.n55 a_n5644_8799.t8 3.61217
R14084 a_n5644_8799.n55 a_n5644_8799.t10 3.61217
R14085 a_n5644_8799.n54 a_n5644_8799.t21 3.61217
R14086 a_n5644_8799.n54 a_n5644_8799.t30 3.61217
R14087 a_n5644_8799.n125 a_n5644_8799.t15 3.61217
R14088 a_n5644_8799.t5 a_n5644_8799.n125 3.61217
R14089 a_n5644_8799.n121 a_n5644_8799.n120 3.4105
R14090 a_n5644_8799.n69 a_n5644_8799.t33 2.82907
R14091 a_n5644_8799.n69 a_n5644_8799.t32 2.82907
R14092 a_n5644_8799.n71 a_n5644_8799.t0 2.82907
R14093 a_n5644_8799.n71 a_n5644_8799.t12 2.82907
R14094 a_n5644_8799.n73 a_n5644_8799.t1 2.82907
R14095 a_n5644_8799.n73 a_n5644_8799.t9 2.82907
R14096 a_n5644_8799.n60 a_n5644_8799.t20 2.82907
R14097 a_n5644_8799.n60 a_n5644_8799.t19 2.82907
R14098 a_n5644_8799.n58 a_n5644_8799.t35 2.82907
R14099 a_n5644_8799.n58 a_n5644_8799.t23 2.82907
R14100 a_n5644_8799.n57 a_n5644_8799.t18 2.82907
R14101 a_n5644_8799.n57 a_n5644_8799.t24 2.82907
R14102 a_n5644_8799.n65 a_n5644_8799.t14 2.82907
R14103 a_n5644_8799.n65 a_n5644_8799.t3 2.82907
R14104 a_n5644_8799.n66 a_n5644_8799.t4 2.82907
R14105 a_n5644_8799.n66 a_n5644_8799.t34 2.82907
R14106 a_n5644_8799.n68 a_n5644_8799.t11 2.82907
R14107 a_n5644_8799.n68 a_n5644_8799.t17 2.82907
R14108 a_n5644_8799.n64 a_n5644_8799.t13 2.82907
R14109 a_n5644_8799.n64 a_n5644_8799.t22 2.82907
R14110 a_n5644_8799.n62 a_n5644_8799.t2 2.82907
R14111 a_n5644_8799.n62 a_n5644_8799.t29 2.82907
R14112 a_n5644_8799.n61 a_n5644_8799.t25 2.82907
R14113 a_n5644_8799.n61 a_n5644_8799.t31 2.82907
R14114 a_n5644_8799.n16 a_n5644_8799.n15 1.13686
R14115 a_n5644_8799.n13 a_n5644_8799.n12 1.13686
R14116 a_n5644_8799.n10 a_n5644_8799.n9 1.13686
R14117 a_n5644_8799.n7 a_n5644_8799.n6 1.13686
R14118 a_n5644_8799.n4 a_n5644_8799.n3 1.13686
R14119 a_n5644_8799.n1 a_n5644_8799.n0 1.13686
R14120 a_n5644_8799.n0 a_n5644_8799.n2 0.568682
R14121 a_n5644_8799.n3 a_n5644_8799.n5 0.568682
R14122 a_n5644_8799.n6 a_n5644_8799.n8 0.568682
R14123 a_n5644_8799.n9 a_n5644_8799.n11 0.568682
R14124 a_n5644_8799.n12 a_n5644_8799.n14 0.568682
R14125 a_n5644_8799.n15 a_n5644_8799.n17 0.568682
R14126 a_n5644_8799.n20 a_n5644_8799.n63 0.530672
R14127 a_n5644_8799.n21 a_n5644_8799.n67 0.530672
R14128 a_n5644_8799.n22 a_n5644_8799.n59 0.530672
R14129 a_n5644_8799.n23 a_n5644_8799.n72 0.530672
R14130 a_n5644_8799.n72 a_n5644_8799.n70 0.530672
R14131 a_n5644_8799.n23 a_n5644_8799.n22 0.530672
R14132 a_n5644_8799.n21 a_n5644_8799.n20 0.530672
R14133 vdd.n291 vdd.n255 756.745
R14134 vdd.n244 vdd.n208 756.745
R14135 vdd.n201 vdd.n165 756.745
R14136 vdd.n154 vdd.n118 756.745
R14137 vdd.n112 vdd.n76 756.745
R14138 vdd.n65 vdd.n29 756.745
R14139 vdd.n1106 vdd.n1070 756.745
R14140 vdd.n1153 vdd.n1117 756.745
R14141 vdd.n1016 vdd.n980 756.745
R14142 vdd.n1063 vdd.n1027 756.745
R14143 vdd.n927 vdd.n891 756.745
R14144 vdd.n974 vdd.n938 756.745
R14145 vdd.n1791 vdd.t68 640.208
R14146 vdd.n755 vdd.t53 640.208
R14147 vdd.n1765 vdd.t94 640.208
R14148 vdd.n747 vdd.t85 640.208
R14149 vdd.n2536 vdd.t36 640.208
R14150 vdd.n2256 vdd.t76 640.208
R14151 vdd.n622 vdd.t57 640.208
R14152 vdd.n2253 vdd.t61 640.208
R14153 vdd.n589 vdd.t65 640.208
R14154 vdd.n817 vdd.t72 640.208
R14155 vdd.n1320 vdd.t32 592.009
R14156 vdd.n1358 vdd.t79 592.009
R14157 vdd.n1254 vdd.t82 592.009
R14158 vdd.n1947 vdd.t28 592.009
R14159 vdd.n1584 vdd.t40 592.009
R14160 vdd.n1544 vdd.t47 592.009
R14161 vdd.n2908 vdd.t91 592.009
R14162 vdd.n405 vdd.t43 592.009
R14163 vdd.n365 vdd.t50 592.009
R14164 vdd.n557 vdd.t21 592.009
R14165 vdd.n2804 vdd.t25 592.009
R14166 vdd.n2711 vdd.t88 592.009
R14167 vdd.n292 vdd.n291 585
R14168 vdd.n290 vdd.n257 585
R14169 vdd.n289 vdd.n288 585
R14170 vdd.n260 vdd.n258 585
R14171 vdd.n283 vdd.n282 585
R14172 vdd.n281 vdd.n280 585
R14173 vdd.n264 vdd.n263 585
R14174 vdd.n275 vdd.n274 585
R14175 vdd.n273 vdd.n272 585
R14176 vdd.n268 vdd.n267 585
R14177 vdd.n245 vdd.n244 585
R14178 vdd.n243 vdd.n210 585
R14179 vdd.n242 vdd.n241 585
R14180 vdd.n213 vdd.n211 585
R14181 vdd.n236 vdd.n235 585
R14182 vdd.n234 vdd.n233 585
R14183 vdd.n217 vdd.n216 585
R14184 vdd.n228 vdd.n227 585
R14185 vdd.n226 vdd.n225 585
R14186 vdd.n221 vdd.n220 585
R14187 vdd.n202 vdd.n201 585
R14188 vdd.n200 vdd.n167 585
R14189 vdd.n199 vdd.n198 585
R14190 vdd.n170 vdd.n168 585
R14191 vdd.n193 vdd.n192 585
R14192 vdd.n191 vdd.n190 585
R14193 vdd.n174 vdd.n173 585
R14194 vdd.n185 vdd.n184 585
R14195 vdd.n183 vdd.n182 585
R14196 vdd.n178 vdd.n177 585
R14197 vdd.n155 vdd.n154 585
R14198 vdd.n153 vdd.n120 585
R14199 vdd.n152 vdd.n151 585
R14200 vdd.n123 vdd.n121 585
R14201 vdd.n146 vdd.n145 585
R14202 vdd.n144 vdd.n143 585
R14203 vdd.n127 vdd.n126 585
R14204 vdd.n138 vdd.n137 585
R14205 vdd.n136 vdd.n135 585
R14206 vdd.n131 vdd.n130 585
R14207 vdd.n113 vdd.n112 585
R14208 vdd.n111 vdd.n78 585
R14209 vdd.n110 vdd.n109 585
R14210 vdd.n81 vdd.n79 585
R14211 vdd.n104 vdd.n103 585
R14212 vdd.n102 vdd.n101 585
R14213 vdd.n85 vdd.n84 585
R14214 vdd.n96 vdd.n95 585
R14215 vdd.n94 vdd.n93 585
R14216 vdd.n89 vdd.n88 585
R14217 vdd.n66 vdd.n65 585
R14218 vdd.n64 vdd.n31 585
R14219 vdd.n63 vdd.n62 585
R14220 vdd.n34 vdd.n32 585
R14221 vdd.n57 vdd.n56 585
R14222 vdd.n55 vdd.n54 585
R14223 vdd.n38 vdd.n37 585
R14224 vdd.n49 vdd.n48 585
R14225 vdd.n47 vdd.n46 585
R14226 vdd.n42 vdd.n41 585
R14227 vdd.n1107 vdd.n1106 585
R14228 vdd.n1105 vdd.n1072 585
R14229 vdd.n1104 vdd.n1103 585
R14230 vdd.n1075 vdd.n1073 585
R14231 vdd.n1098 vdd.n1097 585
R14232 vdd.n1096 vdd.n1095 585
R14233 vdd.n1079 vdd.n1078 585
R14234 vdd.n1090 vdd.n1089 585
R14235 vdd.n1088 vdd.n1087 585
R14236 vdd.n1083 vdd.n1082 585
R14237 vdd.n1154 vdd.n1153 585
R14238 vdd.n1152 vdd.n1119 585
R14239 vdd.n1151 vdd.n1150 585
R14240 vdd.n1122 vdd.n1120 585
R14241 vdd.n1145 vdd.n1144 585
R14242 vdd.n1143 vdd.n1142 585
R14243 vdd.n1126 vdd.n1125 585
R14244 vdd.n1137 vdd.n1136 585
R14245 vdd.n1135 vdd.n1134 585
R14246 vdd.n1130 vdd.n1129 585
R14247 vdd.n1017 vdd.n1016 585
R14248 vdd.n1015 vdd.n982 585
R14249 vdd.n1014 vdd.n1013 585
R14250 vdd.n985 vdd.n983 585
R14251 vdd.n1008 vdd.n1007 585
R14252 vdd.n1006 vdd.n1005 585
R14253 vdd.n989 vdd.n988 585
R14254 vdd.n1000 vdd.n999 585
R14255 vdd.n998 vdd.n997 585
R14256 vdd.n993 vdd.n992 585
R14257 vdd.n1064 vdd.n1063 585
R14258 vdd.n1062 vdd.n1029 585
R14259 vdd.n1061 vdd.n1060 585
R14260 vdd.n1032 vdd.n1030 585
R14261 vdd.n1055 vdd.n1054 585
R14262 vdd.n1053 vdd.n1052 585
R14263 vdd.n1036 vdd.n1035 585
R14264 vdd.n1047 vdd.n1046 585
R14265 vdd.n1045 vdd.n1044 585
R14266 vdd.n1040 vdd.n1039 585
R14267 vdd.n928 vdd.n927 585
R14268 vdd.n926 vdd.n893 585
R14269 vdd.n925 vdd.n924 585
R14270 vdd.n896 vdd.n894 585
R14271 vdd.n919 vdd.n918 585
R14272 vdd.n917 vdd.n916 585
R14273 vdd.n900 vdd.n899 585
R14274 vdd.n911 vdd.n910 585
R14275 vdd.n909 vdd.n908 585
R14276 vdd.n904 vdd.n903 585
R14277 vdd.n975 vdd.n974 585
R14278 vdd.n973 vdd.n940 585
R14279 vdd.n972 vdd.n971 585
R14280 vdd.n943 vdd.n941 585
R14281 vdd.n966 vdd.n965 585
R14282 vdd.n964 vdd.n963 585
R14283 vdd.n947 vdd.n946 585
R14284 vdd.n958 vdd.n957 585
R14285 vdd.n956 vdd.n955 585
R14286 vdd.n951 vdd.n950 585
R14287 vdd.n3024 vdd.n330 515.122
R14288 vdd.n2906 vdd.n328 515.122
R14289 vdd.n515 vdd.n478 515.122
R14290 vdd.n2842 vdd.n479 515.122
R14291 vdd.n1942 vdd.n865 515.122
R14292 vdd.n1945 vdd.n1944 515.122
R14293 vdd.n1227 vdd.n1191 515.122
R14294 vdd.n1423 vdd.n1192 515.122
R14295 vdd.n269 vdd.t121 329.043
R14296 vdd.n222 vdd.t132 329.043
R14297 vdd.n179 vdd.t117 329.043
R14298 vdd.n132 vdd.t127 329.043
R14299 vdd.n90 vdd.t158 329.043
R14300 vdd.n43 vdd.t100 329.043
R14301 vdd.n1084 vdd.t156 329.043
R14302 vdd.n1131 vdd.t142 329.043
R14303 vdd.n994 vdd.t148 329.043
R14304 vdd.n1041 vdd.t135 329.043
R14305 vdd.n905 vdd.t98 329.043
R14306 vdd.n952 vdd.t157 329.043
R14307 vdd.n1320 vdd.t35 319.788
R14308 vdd.n1358 vdd.t81 319.788
R14309 vdd.n1254 vdd.t84 319.788
R14310 vdd.n1947 vdd.t30 319.788
R14311 vdd.n1584 vdd.t41 319.788
R14312 vdd.n1544 vdd.t48 319.788
R14313 vdd.n2908 vdd.t92 319.788
R14314 vdd.n405 vdd.t45 319.788
R14315 vdd.n365 vdd.t51 319.788
R14316 vdd.n557 vdd.t24 319.788
R14317 vdd.n2804 vdd.t27 319.788
R14318 vdd.n2711 vdd.t90 319.788
R14319 vdd.n1321 vdd.t34 303.69
R14320 vdd.n1359 vdd.t80 303.69
R14321 vdd.n1255 vdd.t83 303.69
R14322 vdd.n1948 vdd.t31 303.69
R14323 vdd.n1585 vdd.t42 303.69
R14324 vdd.n1545 vdd.t49 303.69
R14325 vdd.n2909 vdd.t93 303.69
R14326 vdd.n406 vdd.t46 303.69
R14327 vdd.n366 vdd.t52 303.69
R14328 vdd.n558 vdd.t23 303.69
R14329 vdd.n2805 vdd.t26 303.69
R14330 vdd.n2712 vdd.t89 303.69
R14331 vdd.n2479 vdd.n703 297.074
R14332 vdd.n2672 vdd.n599 297.074
R14333 vdd.n2609 vdd.n596 297.074
R14334 vdd.n2402 vdd.n704 297.074
R14335 vdd.n2217 vdd.n744 297.074
R14336 vdd.n2148 vdd.n2147 297.074
R14337 vdd.n1894 vdd.n840 297.074
R14338 vdd.n1990 vdd.n838 297.074
R14339 vdd.n2588 vdd.n597 297.074
R14340 vdd.n2675 vdd.n2674 297.074
R14341 vdd.n2251 vdd.n705 297.074
R14342 vdd.n2477 vdd.n706 297.074
R14343 vdd.n2145 vdd.n753 297.074
R14344 vdd.n751 vdd.n726 297.074
R14345 vdd.n1831 vdd.n841 297.074
R14346 vdd.n1988 vdd.n842 297.074
R14347 vdd.n2590 vdd.n597 185
R14348 vdd.n2673 vdd.n597 185
R14349 vdd.n2592 vdd.n2591 185
R14350 vdd.n2591 vdd.n595 185
R14351 vdd.n2593 vdd.n629 185
R14352 vdd.n2603 vdd.n629 185
R14353 vdd.n2594 vdd.n638 185
R14354 vdd.n638 vdd.n636 185
R14355 vdd.n2596 vdd.n2595 185
R14356 vdd.n2597 vdd.n2596 185
R14357 vdd.n2549 vdd.n637 185
R14358 vdd.n637 vdd.n633 185
R14359 vdd.n2548 vdd.n2547 185
R14360 vdd.n2547 vdd.n2546 185
R14361 vdd.n640 vdd.n639 185
R14362 vdd.n641 vdd.n640 185
R14363 vdd.n2539 vdd.n2538 185
R14364 vdd.n2540 vdd.n2539 185
R14365 vdd.n2535 vdd.n650 185
R14366 vdd.n650 vdd.n647 185
R14367 vdd.n2534 vdd.n2533 185
R14368 vdd.n2533 vdd.n2532 185
R14369 vdd.n652 vdd.n651 185
R14370 vdd.n660 vdd.n652 185
R14371 vdd.n2525 vdd.n2524 185
R14372 vdd.n2526 vdd.n2525 185
R14373 vdd.n2523 vdd.n661 185
R14374 vdd.n2374 vdd.n661 185
R14375 vdd.n2522 vdd.n2521 185
R14376 vdd.n2521 vdd.n2520 185
R14377 vdd.n663 vdd.n662 185
R14378 vdd.n664 vdd.n663 185
R14379 vdd.n2513 vdd.n2512 185
R14380 vdd.n2514 vdd.n2513 185
R14381 vdd.n2511 vdd.n673 185
R14382 vdd.n673 vdd.n670 185
R14383 vdd.n2510 vdd.n2509 185
R14384 vdd.n2509 vdd.n2508 185
R14385 vdd.n675 vdd.n674 185
R14386 vdd.n683 vdd.n675 185
R14387 vdd.n2501 vdd.n2500 185
R14388 vdd.n2502 vdd.n2501 185
R14389 vdd.n2499 vdd.n684 185
R14390 vdd.n690 vdd.n684 185
R14391 vdd.n2498 vdd.n2497 185
R14392 vdd.n2497 vdd.n2496 185
R14393 vdd.n686 vdd.n685 185
R14394 vdd.n687 vdd.n686 185
R14395 vdd.n2489 vdd.n2488 185
R14396 vdd.n2490 vdd.n2489 185
R14397 vdd.n2487 vdd.n696 185
R14398 vdd.n2395 vdd.n696 185
R14399 vdd.n2486 vdd.n2485 185
R14400 vdd.n2485 vdd.n2484 185
R14401 vdd.n698 vdd.n697 185
R14402 vdd.t196 vdd.n698 185
R14403 vdd.n2477 vdd.n2476 185
R14404 vdd.n2478 vdd.n2477 185
R14405 vdd.n2475 vdd.n706 185
R14406 vdd.n2474 vdd.n2473 185
R14407 vdd.n708 vdd.n707 185
R14408 vdd.n2260 vdd.n2259 185
R14409 vdd.n2262 vdd.n2261 185
R14410 vdd.n2264 vdd.n2263 185
R14411 vdd.n2266 vdd.n2265 185
R14412 vdd.n2268 vdd.n2267 185
R14413 vdd.n2270 vdd.n2269 185
R14414 vdd.n2272 vdd.n2271 185
R14415 vdd.n2274 vdd.n2273 185
R14416 vdd.n2276 vdd.n2275 185
R14417 vdd.n2278 vdd.n2277 185
R14418 vdd.n2280 vdd.n2279 185
R14419 vdd.n2282 vdd.n2281 185
R14420 vdd.n2284 vdd.n2283 185
R14421 vdd.n2286 vdd.n2285 185
R14422 vdd.n2288 vdd.n2287 185
R14423 vdd.n2290 vdd.n2289 185
R14424 vdd.n2292 vdd.n2291 185
R14425 vdd.n2294 vdd.n2293 185
R14426 vdd.n2296 vdd.n2295 185
R14427 vdd.n2298 vdd.n2297 185
R14428 vdd.n2300 vdd.n2299 185
R14429 vdd.n2302 vdd.n2301 185
R14430 vdd.n2304 vdd.n2303 185
R14431 vdd.n2306 vdd.n2305 185
R14432 vdd.n2308 vdd.n2307 185
R14433 vdd.n2310 vdd.n2309 185
R14434 vdd.n2312 vdd.n2311 185
R14435 vdd.n2314 vdd.n2313 185
R14436 vdd.n2316 vdd.n2315 185
R14437 vdd.n2318 vdd.n2317 185
R14438 vdd.n2320 vdd.n2319 185
R14439 vdd.n2321 vdd.n2251 185
R14440 vdd.n2471 vdd.n2251 185
R14441 vdd.n2676 vdd.n2675 185
R14442 vdd.n2677 vdd.n588 185
R14443 vdd.n2679 vdd.n2678 185
R14444 vdd.n2681 vdd.n586 185
R14445 vdd.n2683 vdd.n2682 185
R14446 vdd.n2684 vdd.n585 185
R14447 vdd.n2686 vdd.n2685 185
R14448 vdd.n2688 vdd.n583 185
R14449 vdd.n2690 vdd.n2689 185
R14450 vdd.n2691 vdd.n582 185
R14451 vdd.n2693 vdd.n2692 185
R14452 vdd.n2695 vdd.n580 185
R14453 vdd.n2697 vdd.n2696 185
R14454 vdd.n2698 vdd.n579 185
R14455 vdd.n2700 vdd.n2699 185
R14456 vdd.n2702 vdd.n578 185
R14457 vdd.n2703 vdd.n576 185
R14458 vdd.n2706 vdd.n2705 185
R14459 vdd.n577 vdd.n575 185
R14460 vdd.n2562 vdd.n2561 185
R14461 vdd.n2564 vdd.n2563 185
R14462 vdd.n2566 vdd.n2558 185
R14463 vdd.n2568 vdd.n2567 185
R14464 vdd.n2569 vdd.n2557 185
R14465 vdd.n2571 vdd.n2570 185
R14466 vdd.n2573 vdd.n2555 185
R14467 vdd.n2575 vdd.n2574 185
R14468 vdd.n2576 vdd.n2554 185
R14469 vdd.n2578 vdd.n2577 185
R14470 vdd.n2580 vdd.n2552 185
R14471 vdd.n2582 vdd.n2581 185
R14472 vdd.n2583 vdd.n2551 185
R14473 vdd.n2585 vdd.n2584 185
R14474 vdd.n2587 vdd.n2550 185
R14475 vdd.n2589 vdd.n2588 185
R14476 vdd.n2588 vdd.n484 185
R14477 vdd.n2674 vdd.n592 185
R14478 vdd.n2674 vdd.n2673 185
R14479 vdd.n2326 vdd.n594 185
R14480 vdd.n595 vdd.n594 185
R14481 vdd.n2327 vdd.n628 185
R14482 vdd.n2603 vdd.n628 185
R14483 vdd.n2329 vdd.n2328 185
R14484 vdd.n2328 vdd.n636 185
R14485 vdd.n2330 vdd.n635 185
R14486 vdd.n2597 vdd.n635 185
R14487 vdd.n2332 vdd.n2331 185
R14488 vdd.n2331 vdd.n633 185
R14489 vdd.n2333 vdd.n643 185
R14490 vdd.n2546 vdd.n643 185
R14491 vdd.n2335 vdd.n2334 185
R14492 vdd.n2334 vdd.n641 185
R14493 vdd.n2336 vdd.n649 185
R14494 vdd.n2540 vdd.n649 185
R14495 vdd.n2338 vdd.n2337 185
R14496 vdd.n2337 vdd.n647 185
R14497 vdd.n2339 vdd.n654 185
R14498 vdd.n2532 vdd.n654 185
R14499 vdd.n2341 vdd.n2340 185
R14500 vdd.n2340 vdd.n660 185
R14501 vdd.n2342 vdd.n659 185
R14502 vdd.n2526 vdd.n659 185
R14503 vdd.n2376 vdd.n2375 185
R14504 vdd.n2375 vdd.n2374 185
R14505 vdd.n2377 vdd.n666 185
R14506 vdd.n2520 vdd.n666 185
R14507 vdd.n2379 vdd.n2378 185
R14508 vdd.n2378 vdd.n664 185
R14509 vdd.n2380 vdd.n672 185
R14510 vdd.n2514 vdd.n672 185
R14511 vdd.n2382 vdd.n2381 185
R14512 vdd.n2381 vdd.n670 185
R14513 vdd.n2383 vdd.n677 185
R14514 vdd.n2508 vdd.n677 185
R14515 vdd.n2385 vdd.n2384 185
R14516 vdd.n2384 vdd.n683 185
R14517 vdd.n2386 vdd.n682 185
R14518 vdd.n2502 vdd.n682 185
R14519 vdd.n2388 vdd.n2387 185
R14520 vdd.n2387 vdd.n690 185
R14521 vdd.n2389 vdd.n689 185
R14522 vdd.n2496 vdd.n689 185
R14523 vdd.n2391 vdd.n2390 185
R14524 vdd.n2390 vdd.n687 185
R14525 vdd.n2392 vdd.n695 185
R14526 vdd.n2490 vdd.n695 185
R14527 vdd.n2394 vdd.n2393 185
R14528 vdd.n2395 vdd.n2394 185
R14529 vdd.n2325 vdd.n700 185
R14530 vdd.n2484 vdd.n700 185
R14531 vdd.n2324 vdd.n2323 185
R14532 vdd.n2323 vdd.t196 185
R14533 vdd.n2322 vdd.n705 185
R14534 vdd.n2478 vdd.n705 185
R14535 vdd.n1942 vdd.n1941 185
R14536 vdd.n1943 vdd.n1942 185
R14537 vdd.n866 vdd.n864 185
R14538 vdd.n1508 vdd.n864 185
R14539 vdd.n1511 vdd.n1510 185
R14540 vdd.n1510 vdd.n1509 185
R14541 vdd.n869 vdd.n868 185
R14542 vdd.n870 vdd.n869 185
R14543 vdd.n1497 vdd.n1496 185
R14544 vdd.n1498 vdd.n1497 185
R14545 vdd.n878 vdd.n877 185
R14546 vdd.n1489 vdd.n877 185
R14547 vdd.n1492 vdd.n1491 185
R14548 vdd.n1491 vdd.n1490 185
R14549 vdd.n881 vdd.n880 185
R14550 vdd.n888 vdd.n881 185
R14551 vdd.n1480 vdd.n1479 185
R14552 vdd.n1481 vdd.n1480 185
R14553 vdd.n890 vdd.n889 185
R14554 vdd.n889 vdd.n887 185
R14555 vdd.n1475 vdd.n1474 185
R14556 vdd.n1474 vdd.n1473 185
R14557 vdd.n1163 vdd.n1162 185
R14558 vdd.n1164 vdd.n1163 185
R14559 vdd.n1464 vdd.n1463 185
R14560 vdd.n1465 vdd.n1464 185
R14561 vdd.n1171 vdd.n1170 185
R14562 vdd.n1455 vdd.n1170 185
R14563 vdd.n1458 vdd.n1457 185
R14564 vdd.n1457 vdd.n1456 185
R14565 vdd.n1174 vdd.n1173 185
R14566 vdd.n1180 vdd.n1174 185
R14567 vdd.n1446 vdd.n1445 185
R14568 vdd.n1447 vdd.n1446 185
R14569 vdd.n1182 vdd.n1181 185
R14570 vdd.n1438 vdd.n1181 185
R14571 vdd.n1441 vdd.n1440 185
R14572 vdd.n1440 vdd.n1439 185
R14573 vdd.n1185 vdd.n1184 185
R14574 vdd.n1186 vdd.n1185 185
R14575 vdd.n1429 vdd.n1428 185
R14576 vdd.n1430 vdd.n1429 185
R14577 vdd.n1193 vdd.n1192 185
R14578 vdd.n1228 vdd.n1192 185
R14579 vdd.n1424 vdd.n1423 185
R14580 vdd.n1196 vdd.n1195 185
R14581 vdd.n1420 vdd.n1419 185
R14582 vdd.n1421 vdd.n1420 185
R14583 vdd.n1230 vdd.n1229 185
R14584 vdd.n1415 vdd.n1232 185
R14585 vdd.n1414 vdd.n1233 185
R14586 vdd.n1413 vdd.n1234 185
R14587 vdd.n1236 vdd.n1235 185
R14588 vdd.n1409 vdd.n1238 185
R14589 vdd.n1408 vdd.n1239 185
R14590 vdd.n1407 vdd.n1240 185
R14591 vdd.n1242 vdd.n1241 185
R14592 vdd.n1403 vdd.n1244 185
R14593 vdd.n1402 vdd.n1245 185
R14594 vdd.n1401 vdd.n1246 185
R14595 vdd.n1248 vdd.n1247 185
R14596 vdd.n1397 vdd.n1250 185
R14597 vdd.n1396 vdd.n1251 185
R14598 vdd.n1395 vdd.n1252 185
R14599 vdd.n1256 vdd.n1253 185
R14600 vdd.n1391 vdd.n1258 185
R14601 vdd.n1390 vdd.n1259 185
R14602 vdd.n1389 vdd.n1260 185
R14603 vdd.n1262 vdd.n1261 185
R14604 vdd.n1385 vdd.n1264 185
R14605 vdd.n1384 vdd.n1265 185
R14606 vdd.n1383 vdd.n1266 185
R14607 vdd.n1268 vdd.n1267 185
R14608 vdd.n1379 vdd.n1270 185
R14609 vdd.n1378 vdd.n1271 185
R14610 vdd.n1377 vdd.n1272 185
R14611 vdd.n1274 vdd.n1273 185
R14612 vdd.n1373 vdd.n1276 185
R14613 vdd.n1372 vdd.n1277 185
R14614 vdd.n1371 vdd.n1278 185
R14615 vdd.n1280 vdd.n1279 185
R14616 vdd.n1367 vdd.n1282 185
R14617 vdd.n1366 vdd.n1283 185
R14618 vdd.n1365 vdd.n1284 185
R14619 vdd.n1286 vdd.n1285 185
R14620 vdd.n1361 vdd.n1288 185
R14621 vdd.n1360 vdd.n1357 185
R14622 vdd.n1356 vdd.n1289 185
R14623 vdd.n1291 vdd.n1290 185
R14624 vdd.n1352 vdd.n1293 185
R14625 vdd.n1351 vdd.n1294 185
R14626 vdd.n1350 vdd.n1295 185
R14627 vdd.n1297 vdd.n1296 185
R14628 vdd.n1346 vdd.n1299 185
R14629 vdd.n1345 vdd.n1300 185
R14630 vdd.n1344 vdd.n1301 185
R14631 vdd.n1303 vdd.n1302 185
R14632 vdd.n1340 vdd.n1305 185
R14633 vdd.n1339 vdd.n1306 185
R14634 vdd.n1338 vdd.n1307 185
R14635 vdd.n1309 vdd.n1308 185
R14636 vdd.n1334 vdd.n1311 185
R14637 vdd.n1333 vdd.n1312 185
R14638 vdd.n1332 vdd.n1313 185
R14639 vdd.n1315 vdd.n1314 185
R14640 vdd.n1328 vdd.n1317 185
R14641 vdd.n1327 vdd.n1318 185
R14642 vdd.n1326 vdd.n1319 185
R14643 vdd.n1323 vdd.n1227 185
R14644 vdd.n1421 vdd.n1227 185
R14645 vdd.n1946 vdd.n1945 185
R14646 vdd.n1950 vdd.n859 185
R14647 vdd.n1613 vdd.n858 185
R14648 vdd.n1616 vdd.n1615 185
R14649 vdd.n1618 vdd.n1617 185
R14650 vdd.n1621 vdd.n1620 185
R14651 vdd.n1623 vdd.n1622 185
R14652 vdd.n1625 vdd.n1611 185
R14653 vdd.n1627 vdd.n1626 185
R14654 vdd.n1628 vdd.n1605 185
R14655 vdd.n1630 vdd.n1629 185
R14656 vdd.n1632 vdd.n1603 185
R14657 vdd.n1634 vdd.n1633 185
R14658 vdd.n1635 vdd.n1598 185
R14659 vdd.n1637 vdd.n1636 185
R14660 vdd.n1639 vdd.n1596 185
R14661 vdd.n1641 vdd.n1640 185
R14662 vdd.n1642 vdd.n1592 185
R14663 vdd.n1644 vdd.n1643 185
R14664 vdd.n1646 vdd.n1589 185
R14665 vdd.n1648 vdd.n1647 185
R14666 vdd.n1590 vdd.n1583 185
R14667 vdd.n1652 vdd.n1587 185
R14668 vdd.n1653 vdd.n1579 185
R14669 vdd.n1655 vdd.n1654 185
R14670 vdd.n1657 vdd.n1577 185
R14671 vdd.n1659 vdd.n1658 185
R14672 vdd.n1660 vdd.n1572 185
R14673 vdd.n1662 vdd.n1661 185
R14674 vdd.n1664 vdd.n1570 185
R14675 vdd.n1666 vdd.n1665 185
R14676 vdd.n1667 vdd.n1565 185
R14677 vdd.n1669 vdd.n1668 185
R14678 vdd.n1671 vdd.n1563 185
R14679 vdd.n1673 vdd.n1672 185
R14680 vdd.n1674 vdd.n1558 185
R14681 vdd.n1676 vdd.n1675 185
R14682 vdd.n1678 vdd.n1556 185
R14683 vdd.n1680 vdd.n1679 185
R14684 vdd.n1681 vdd.n1552 185
R14685 vdd.n1683 vdd.n1682 185
R14686 vdd.n1685 vdd.n1549 185
R14687 vdd.n1687 vdd.n1686 185
R14688 vdd.n1550 vdd.n1543 185
R14689 vdd.n1691 vdd.n1547 185
R14690 vdd.n1692 vdd.n1539 185
R14691 vdd.n1694 vdd.n1693 185
R14692 vdd.n1696 vdd.n1537 185
R14693 vdd.n1698 vdd.n1697 185
R14694 vdd.n1699 vdd.n1532 185
R14695 vdd.n1701 vdd.n1700 185
R14696 vdd.n1703 vdd.n1530 185
R14697 vdd.n1705 vdd.n1704 185
R14698 vdd.n1706 vdd.n1525 185
R14699 vdd.n1708 vdd.n1707 185
R14700 vdd.n1710 vdd.n1524 185
R14701 vdd.n1711 vdd.n1521 185
R14702 vdd.n1714 vdd.n1713 185
R14703 vdd.n1523 vdd.n1519 185
R14704 vdd.n1931 vdd.n1517 185
R14705 vdd.n1933 vdd.n1932 185
R14706 vdd.n1935 vdd.n1515 185
R14707 vdd.n1937 vdd.n1936 185
R14708 vdd.n1938 vdd.n865 185
R14709 vdd.n1944 vdd.n862 185
R14710 vdd.n1944 vdd.n1943 185
R14711 vdd.n873 vdd.n861 185
R14712 vdd.n1508 vdd.n861 185
R14713 vdd.n1507 vdd.n1506 185
R14714 vdd.n1509 vdd.n1507 185
R14715 vdd.n872 vdd.n871 185
R14716 vdd.n871 vdd.n870 185
R14717 vdd.n1500 vdd.n1499 185
R14718 vdd.n1499 vdd.n1498 185
R14719 vdd.n876 vdd.n875 185
R14720 vdd.n1489 vdd.n876 185
R14721 vdd.n1488 vdd.n1487 185
R14722 vdd.n1490 vdd.n1488 185
R14723 vdd.n883 vdd.n882 185
R14724 vdd.n888 vdd.n882 185
R14725 vdd.n1483 vdd.n1482 185
R14726 vdd.n1482 vdd.n1481 185
R14727 vdd.n886 vdd.n885 185
R14728 vdd.n887 vdd.n886 185
R14729 vdd.n1472 vdd.n1471 185
R14730 vdd.n1473 vdd.n1472 185
R14731 vdd.n1166 vdd.n1165 185
R14732 vdd.n1165 vdd.n1164 185
R14733 vdd.n1467 vdd.n1466 185
R14734 vdd.n1466 vdd.n1465 185
R14735 vdd.n1169 vdd.n1168 185
R14736 vdd.n1455 vdd.n1169 185
R14737 vdd.n1454 vdd.n1453 185
R14738 vdd.n1456 vdd.n1454 185
R14739 vdd.n1176 vdd.n1175 185
R14740 vdd.n1180 vdd.n1175 185
R14741 vdd.n1449 vdd.n1448 185
R14742 vdd.n1448 vdd.n1447 185
R14743 vdd.n1179 vdd.n1178 185
R14744 vdd.n1438 vdd.n1179 185
R14745 vdd.n1437 vdd.n1436 185
R14746 vdd.n1439 vdd.n1437 185
R14747 vdd.n1188 vdd.n1187 185
R14748 vdd.n1187 vdd.n1186 185
R14749 vdd.n1432 vdd.n1431 185
R14750 vdd.n1431 vdd.n1430 185
R14751 vdd.n1191 vdd.n1190 185
R14752 vdd.n1228 vdd.n1191 185
R14753 vdd.n746 vdd.n744 185
R14754 vdd.n2146 vdd.n744 185
R14755 vdd.n2068 vdd.n763 185
R14756 vdd.n763 vdd.t19 185
R14757 vdd.n2070 vdd.n2069 185
R14758 vdd.n2071 vdd.n2070 185
R14759 vdd.n2067 vdd.n762 185
R14760 vdd.n1770 vdd.n762 185
R14761 vdd.n2066 vdd.n2065 185
R14762 vdd.n2065 vdd.n2064 185
R14763 vdd.n765 vdd.n764 185
R14764 vdd.n766 vdd.n765 185
R14765 vdd.n2055 vdd.n2054 185
R14766 vdd.n2056 vdd.n2055 185
R14767 vdd.n2053 vdd.n776 185
R14768 vdd.n776 vdd.n773 185
R14769 vdd.n2052 vdd.n2051 185
R14770 vdd.n2051 vdd.n2050 185
R14771 vdd.n778 vdd.n777 185
R14772 vdd.n779 vdd.n778 185
R14773 vdd.n2043 vdd.n2042 185
R14774 vdd.n2044 vdd.n2043 185
R14775 vdd.n2041 vdd.n787 185
R14776 vdd.n792 vdd.n787 185
R14777 vdd.n2040 vdd.n2039 185
R14778 vdd.n2039 vdd.n2038 185
R14779 vdd.n789 vdd.n788 185
R14780 vdd.n798 vdd.n789 185
R14781 vdd.n2031 vdd.n2030 185
R14782 vdd.n2032 vdd.n2031 185
R14783 vdd.n2029 vdd.n799 185
R14784 vdd.n1871 vdd.n799 185
R14785 vdd.n2028 vdd.n2027 185
R14786 vdd.n2027 vdd.n2026 185
R14787 vdd.n801 vdd.n800 185
R14788 vdd.n802 vdd.n801 185
R14789 vdd.n2019 vdd.n2018 185
R14790 vdd.n2020 vdd.n2019 185
R14791 vdd.n2017 vdd.n811 185
R14792 vdd.n811 vdd.n808 185
R14793 vdd.n2016 vdd.n2015 185
R14794 vdd.n2015 vdd.n2014 185
R14795 vdd.n813 vdd.n812 185
R14796 vdd.n823 vdd.n813 185
R14797 vdd.n2006 vdd.n2005 185
R14798 vdd.n2007 vdd.n2006 185
R14799 vdd.n2004 vdd.n824 185
R14800 vdd.n824 vdd.n820 185
R14801 vdd.n2003 vdd.n2002 185
R14802 vdd.n2002 vdd.n2001 185
R14803 vdd.n826 vdd.n825 185
R14804 vdd.n827 vdd.n826 185
R14805 vdd.n1994 vdd.n1993 185
R14806 vdd.n1995 vdd.n1994 185
R14807 vdd.n1992 vdd.n836 185
R14808 vdd.n836 vdd.n833 185
R14809 vdd.n1991 vdd.n1990 185
R14810 vdd.n1990 vdd.n1989 185
R14811 vdd.n838 vdd.n837 185
R14812 vdd.n1726 vdd.n1725 185
R14813 vdd.n1727 vdd.n1723 185
R14814 vdd.n1723 vdd.n839 185
R14815 vdd.n1729 vdd.n1728 185
R14816 vdd.n1731 vdd.n1722 185
R14817 vdd.n1734 vdd.n1733 185
R14818 vdd.n1735 vdd.n1721 185
R14819 vdd.n1737 vdd.n1736 185
R14820 vdd.n1739 vdd.n1720 185
R14821 vdd.n1742 vdd.n1741 185
R14822 vdd.n1743 vdd.n1719 185
R14823 vdd.n1745 vdd.n1744 185
R14824 vdd.n1747 vdd.n1718 185
R14825 vdd.n1750 vdd.n1749 185
R14826 vdd.n1751 vdd.n1717 185
R14827 vdd.n1753 vdd.n1752 185
R14828 vdd.n1755 vdd.n1716 185
R14829 vdd.n1928 vdd.n1756 185
R14830 vdd.n1927 vdd.n1926 185
R14831 vdd.n1924 vdd.n1757 185
R14832 vdd.n1922 vdd.n1921 185
R14833 vdd.n1920 vdd.n1758 185
R14834 vdd.n1919 vdd.n1918 185
R14835 vdd.n1916 vdd.n1759 185
R14836 vdd.n1914 vdd.n1913 185
R14837 vdd.n1912 vdd.n1760 185
R14838 vdd.n1911 vdd.n1910 185
R14839 vdd.n1908 vdd.n1761 185
R14840 vdd.n1906 vdd.n1905 185
R14841 vdd.n1904 vdd.n1762 185
R14842 vdd.n1903 vdd.n1902 185
R14843 vdd.n1900 vdd.n1763 185
R14844 vdd.n1898 vdd.n1897 185
R14845 vdd.n1896 vdd.n1764 185
R14846 vdd.n1895 vdd.n1894 185
R14847 vdd.n2149 vdd.n2148 185
R14848 vdd.n2151 vdd.n2150 185
R14849 vdd.n2153 vdd.n2152 185
R14850 vdd.n2156 vdd.n2155 185
R14851 vdd.n2158 vdd.n2157 185
R14852 vdd.n2160 vdd.n2159 185
R14853 vdd.n2162 vdd.n2161 185
R14854 vdd.n2164 vdd.n2163 185
R14855 vdd.n2166 vdd.n2165 185
R14856 vdd.n2168 vdd.n2167 185
R14857 vdd.n2170 vdd.n2169 185
R14858 vdd.n2172 vdd.n2171 185
R14859 vdd.n2174 vdd.n2173 185
R14860 vdd.n2176 vdd.n2175 185
R14861 vdd.n2178 vdd.n2177 185
R14862 vdd.n2180 vdd.n2179 185
R14863 vdd.n2182 vdd.n2181 185
R14864 vdd.n2184 vdd.n2183 185
R14865 vdd.n2186 vdd.n2185 185
R14866 vdd.n2188 vdd.n2187 185
R14867 vdd.n2190 vdd.n2189 185
R14868 vdd.n2192 vdd.n2191 185
R14869 vdd.n2194 vdd.n2193 185
R14870 vdd.n2196 vdd.n2195 185
R14871 vdd.n2198 vdd.n2197 185
R14872 vdd.n2200 vdd.n2199 185
R14873 vdd.n2202 vdd.n2201 185
R14874 vdd.n2204 vdd.n2203 185
R14875 vdd.n2206 vdd.n2205 185
R14876 vdd.n2208 vdd.n2207 185
R14877 vdd.n2210 vdd.n2209 185
R14878 vdd.n2212 vdd.n2211 185
R14879 vdd.n2214 vdd.n2213 185
R14880 vdd.n2215 vdd.n745 185
R14881 vdd.n2217 vdd.n2216 185
R14882 vdd.n2218 vdd.n2217 185
R14883 vdd.n2147 vdd.n749 185
R14884 vdd.n2147 vdd.n2146 185
R14885 vdd.n1768 vdd.n750 185
R14886 vdd.t19 vdd.n750 185
R14887 vdd.n1769 vdd.n760 185
R14888 vdd.n2071 vdd.n760 185
R14889 vdd.n1772 vdd.n1771 185
R14890 vdd.n1771 vdd.n1770 185
R14891 vdd.n1773 vdd.n767 185
R14892 vdd.n2064 vdd.n767 185
R14893 vdd.n1775 vdd.n1774 185
R14894 vdd.n1774 vdd.n766 185
R14895 vdd.n1776 vdd.n774 185
R14896 vdd.n2056 vdd.n774 185
R14897 vdd.n1778 vdd.n1777 185
R14898 vdd.n1777 vdd.n773 185
R14899 vdd.n1779 vdd.n780 185
R14900 vdd.n2050 vdd.n780 185
R14901 vdd.n1781 vdd.n1780 185
R14902 vdd.n1780 vdd.n779 185
R14903 vdd.n1782 vdd.n785 185
R14904 vdd.n2044 vdd.n785 185
R14905 vdd.n1784 vdd.n1783 185
R14906 vdd.n1783 vdd.n792 185
R14907 vdd.n1785 vdd.n790 185
R14908 vdd.n2038 vdd.n790 185
R14909 vdd.n1787 vdd.n1786 185
R14910 vdd.n1786 vdd.n798 185
R14911 vdd.n1788 vdd.n796 185
R14912 vdd.n2032 vdd.n796 185
R14913 vdd.n1873 vdd.n1872 185
R14914 vdd.n1872 vdd.n1871 185
R14915 vdd.n1874 vdd.n803 185
R14916 vdd.n2026 vdd.n803 185
R14917 vdd.n1876 vdd.n1875 185
R14918 vdd.n1875 vdd.n802 185
R14919 vdd.n1877 vdd.n809 185
R14920 vdd.n2020 vdd.n809 185
R14921 vdd.n1879 vdd.n1878 185
R14922 vdd.n1878 vdd.n808 185
R14923 vdd.n1880 vdd.n814 185
R14924 vdd.n2014 vdd.n814 185
R14925 vdd.n1882 vdd.n1881 185
R14926 vdd.n1881 vdd.n823 185
R14927 vdd.n1883 vdd.n821 185
R14928 vdd.n2007 vdd.n821 185
R14929 vdd.n1885 vdd.n1884 185
R14930 vdd.n1884 vdd.n820 185
R14931 vdd.n1886 vdd.n828 185
R14932 vdd.n2001 vdd.n828 185
R14933 vdd.n1888 vdd.n1887 185
R14934 vdd.n1887 vdd.n827 185
R14935 vdd.n1889 vdd.n834 185
R14936 vdd.n1995 vdd.n834 185
R14937 vdd.n1891 vdd.n1890 185
R14938 vdd.n1890 vdd.n833 185
R14939 vdd.n1892 vdd.n840 185
R14940 vdd.n1989 vdd.n840 185
R14941 vdd.n3024 vdd.n3023 185
R14942 vdd.n3025 vdd.n3024 185
R14943 vdd.n325 vdd.n324 185
R14944 vdd.n3026 vdd.n325 185
R14945 vdd.n3029 vdd.n3028 185
R14946 vdd.n3028 vdd.n3027 185
R14947 vdd.n3030 vdd.n319 185
R14948 vdd.n319 vdd.n318 185
R14949 vdd.n3032 vdd.n3031 185
R14950 vdd.n3033 vdd.n3032 185
R14951 vdd.n314 vdd.n313 185
R14952 vdd.n3034 vdd.n314 185
R14953 vdd.n3037 vdd.n3036 185
R14954 vdd.n3036 vdd.n3035 185
R14955 vdd.n3038 vdd.n309 185
R14956 vdd.n309 vdd.n308 185
R14957 vdd.n3040 vdd.n3039 185
R14958 vdd.n3041 vdd.n3040 185
R14959 vdd.n303 vdd.n301 185
R14960 vdd.n3042 vdd.n303 185
R14961 vdd.n3045 vdd.n3044 185
R14962 vdd.n3044 vdd.n3043 185
R14963 vdd.n302 vdd.n300 185
R14964 vdd.n304 vdd.n302 185
R14965 vdd.n2881 vdd.n2880 185
R14966 vdd.n2882 vdd.n2881 185
R14967 vdd.n458 vdd.n457 185
R14968 vdd.n457 vdd.n456 185
R14969 vdd.n2876 vdd.n2875 185
R14970 vdd.n2875 vdd.n2874 185
R14971 vdd.n461 vdd.n460 185
R14972 vdd.n467 vdd.n461 185
R14973 vdd.n2865 vdd.n2864 185
R14974 vdd.n2866 vdd.n2865 185
R14975 vdd.n469 vdd.n468 185
R14976 vdd.n2857 vdd.n468 185
R14977 vdd.n2860 vdd.n2859 185
R14978 vdd.n2859 vdd.n2858 185
R14979 vdd.n472 vdd.n471 185
R14980 vdd.n473 vdd.n472 185
R14981 vdd.n2848 vdd.n2847 185
R14982 vdd.n2849 vdd.n2848 185
R14983 vdd.n480 vdd.n479 185
R14984 vdd.n516 vdd.n479 185
R14985 vdd.n2843 vdd.n2842 185
R14986 vdd.n483 vdd.n482 185
R14987 vdd.n2839 vdd.n2838 185
R14988 vdd.n2840 vdd.n2839 185
R14989 vdd.n518 vdd.n517 185
R14990 vdd.n522 vdd.n521 185
R14991 vdd.n2834 vdd.n523 185
R14992 vdd.n2833 vdd.n2832 185
R14993 vdd.n2831 vdd.n2830 185
R14994 vdd.n2829 vdd.n2828 185
R14995 vdd.n2827 vdd.n2826 185
R14996 vdd.n2825 vdd.n2824 185
R14997 vdd.n2823 vdd.n2822 185
R14998 vdd.n2821 vdd.n2820 185
R14999 vdd.n2819 vdd.n2818 185
R15000 vdd.n2817 vdd.n2816 185
R15001 vdd.n2815 vdd.n2814 185
R15002 vdd.n2813 vdd.n2812 185
R15003 vdd.n2811 vdd.n2810 185
R15004 vdd.n2809 vdd.n2808 185
R15005 vdd.n2807 vdd.n2806 185
R15006 vdd.n2798 vdd.n536 185
R15007 vdd.n2800 vdd.n2799 185
R15008 vdd.n2797 vdd.n2796 185
R15009 vdd.n2795 vdd.n2794 185
R15010 vdd.n2793 vdd.n2792 185
R15011 vdd.n2791 vdd.n2790 185
R15012 vdd.n2789 vdd.n2788 185
R15013 vdd.n2787 vdd.n2786 185
R15014 vdd.n2785 vdd.n2784 185
R15015 vdd.n2783 vdd.n2782 185
R15016 vdd.n2781 vdd.n2780 185
R15017 vdd.n2779 vdd.n2778 185
R15018 vdd.n2777 vdd.n2776 185
R15019 vdd.n2775 vdd.n2774 185
R15020 vdd.n2773 vdd.n2772 185
R15021 vdd.n2771 vdd.n2770 185
R15022 vdd.n2769 vdd.n2768 185
R15023 vdd.n2767 vdd.n2766 185
R15024 vdd.n2765 vdd.n2764 185
R15025 vdd.n2763 vdd.n2762 185
R15026 vdd.n2761 vdd.n2760 185
R15027 vdd.n2759 vdd.n2758 185
R15028 vdd.n2752 vdd.n556 185
R15029 vdd.n2754 vdd.n2753 185
R15030 vdd.n2751 vdd.n2750 185
R15031 vdd.n2749 vdd.n2748 185
R15032 vdd.n2747 vdd.n2746 185
R15033 vdd.n2745 vdd.n2744 185
R15034 vdd.n2743 vdd.n2742 185
R15035 vdd.n2741 vdd.n2740 185
R15036 vdd.n2739 vdd.n2738 185
R15037 vdd.n2737 vdd.n2736 185
R15038 vdd.n2735 vdd.n2734 185
R15039 vdd.n2733 vdd.n2732 185
R15040 vdd.n2731 vdd.n2730 185
R15041 vdd.n2729 vdd.n2728 185
R15042 vdd.n2727 vdd.n2726 185
R15043 vdd.n2725 vdd.n2724 185
R15044 vdd.n2723 vdd.n2722 185
R15045 vdd.n2721 vdd.n2720 185
R15046 vdd.n2719 vdd.n2718 185
R15047 vdd.n2717 vdd.n2716 185
R15048 vdd.n2715 vdd.n2714 185
R15049 vdd.n2710 vdd.n515 185
R15050 vdd.n2840 vdd.n515 185
R15051 vdd.n2907 vdd.n2906 185
R15052 vdd.n2911 vdd.n440 185
R15053 vdd.n2913 vdd.n2912 185
R15054 vdd.n2915 vdd.n438 185
R15055 vdd.n2917 vdd.n2916 185
R15056 vdd.n2918 vdd.n433 185
R15057 vdd.n2920 vdd.n2919 185
R15058 vdd.n2922 vdd.n431 185
R15059 vdd.n2924 vdd.n2923 185
R15060 vdd.n2925 vdd.n426 185
R15061 vdd.n2927 vdd.n2926 185
R15062 vdd.n2929 vdd.n424 185
R15063 vdd.n2931 vdd.n2930 185
R15064 vdd.n2932 vdd.n419 185
R15065 vdd.n2934 vdd.n2933 185
R15066 vdd.n2936 vdd.n417 185
R15067 vdd.n2938 vdd.n2937 185
R15068 vdd.n2939 vdd.n413 185
R15069 vdd.n2941 vdd.n2940 185
R15070 vdd.n2943 vdd.n410 185
R15071 vdd.n2945 vdd.n2944 185
R15072 vdd.n411 vdd.n404 185
R15073 vdd.n2949 vdd.n408 185
R15074 vdd.n2950 vdd.n400 185
R15075 vdd.n2952 vdd.n2951 185
R15076 vdd.n2954 vdd.n398 185
R15077 vdd.n2956 vdd.n2955 185
R15078 vdd.n2957 vdd.n393 185
R15079 vdd.n2959 vdd.n2958 185
R15080 vdd.n2961 vdd.n391 185
R15081 vdd.n2963 vdd.n2962 185
R15082 vdd.n2964 vdd.n386 185
R15083 vdd.n2966 vdd.n2965 185
R15084 vdd.n2968 vdd.n384 185
R15085 vdd.n2970 vdd.n2969 185
R15086 vdd.n2971 vdd.n379 185
R15087 vdd.n2973 vdd.n2972 185
R15088 vdd.n2975 vdd.n377 185
R15089 vdd.n2977 vdd.n2976 185
R15090 vdd.n2978 vdd.n373 185
R15091 vdd.n2980 vdd.n2979 185
R15092 vdd.n2982 vdd.n370 185
R15093 vdd.n2984 vdd.n2983 185
R15094 vdd.n371 vdd.n364 185
R15095 vdd.n2988 vdd.n368 185
R15096 vdd.n2989 vdd.n360 185
R15097 vdd.n2991 vdd.n2990 185
R15098 vdd.n2993 vdd.n358 185
R15099 vdd.n2995 vdd.n2994 185
R15100 vdd.n2996 vdd.n353 185
R15101 vdd.n2998 vdd.n2997 185
R15102 vdd.n3000 vdd.n351 185
R15103 vdd.n3002 vdd.n3001 185
R15104 vdd.n3003 vdd.n346 185
R15105 vdd.n3005 vdd.n3004 185
R15106 vdd.n3007 vdd.n344 185
R15107 vdd.n3009 vdd.n3008 185
R15108 vdd.n3010 vdd.n338 185
R15109 vdd.n3012 vdd.n3011 185
R15110 vdd.n3014 vdd.n337 185
R15111 vdd.n3015 vdd.n336 185
R15112 vdd.n3018 vdd.n3017 185
R15113 vdd.n3019 vdd.n334 185
R15114 vdd.n3020 vdd.n330 185
R15115 vdd.n2902 vdd.n328 185
R15116 vdd.n3025 vdd.n328 185
R15117 vdd.n2901 vdd.n327 185
R15118 vdd.n3026 vdd.n327 185
R15119 vdd.n2900 vdd.n326 185
R15120 vdd.n3027 vdd.n326 185
R15121 vdd.n446 vdd.n445 185
R15122 vdd.n445 vdd.n318 185
R15123 vdd.n2896 vdd.n317 185
R15124 vdd.n3033 vdd.n317 185
R15125 vdd.n2895 vdd.n316 185
R15126 vdd.n3034 vdd.n316 185
R15127 vdd.n2894 vdd.n315 185
R15128 vdd.n3035 vdd.n315 185
R15129 vdd.n449 vdd.n448 185
R15130 vdd.n448 vdd.n308 185
R15131 vdd.n2890 vdd.n307 185
R15132 vdd.n3041 vdd.n307 185
R15133 vdd.n2889 vdd.n306 185
R15134 vdd.n3042 vdd.n306 185
R15135 vdd.n2888 vdd.n305 185
R15136 vdd.n3043 vdd.n305 185
R15137 vdd.n455 vdd.n451 185
R15138 vdd.n455 vdd.n304 185
R15139 vdd.n2884 vdd.n2883 185
R15140 vdd.n2883 vdd.n2882 185
R15141 vdd.n454 vdd.n453 185
R15142 vdd.n456 vdd.n454 185
R15143 vdd.n2873 vdd.n2872 185
R15144 vdd.n2874 vdd.n2873 185
R15145 vdd.n463 vdd.n462 185
R15146 vdd.n467 vdd.n462 185
R15147 vdd.n2868 vdd.n2867 185
R15148 vdd.n2867 vdd.n2866 185
R15149 vdd.n466 vdd.n465 185
R15150 vdd.n2857 vdd.n466 185
R15151 vdd.n2856 vdd.n2855 185
R15152 vdd.n2858 vdd.n2856 185
R15153 vdd.n475 vdd.n474 185
R15154 vdd.n474 vdd.n473 185
R15155 vdd.n2851 vdd.n2850 185
R15156 vdd.n2850 vdd.n2849 185
R15157 vdd.n478 vdd.n477 185
R15158 vdd.n516 vdd.n478 185
R15159 vdd.n703 vdd.n702 185
R15160 vdd.n2469 vdd.n2468 185
R15161 vdd.n2467 vdd.n2252 185
R15162 vdd.n2471 vdd.n2252 185
R15163 vdd.n2466 vdd.n2465 185
R15164 vdd.n2464 vdd.n2463 185
R15165 vdd.n2462 vdd.n2461 185
R15166 vdd.n2460 vdd.n2459 185
R15167 vdd.n2458 vdd.n2457 185
R15168 vdd.n2456 vdd.n2455 185
R15169 vdd.n2454 vdd.n2453 185
R15170 vdd.n2452 vdd.n2451 185
R15171 vdd.n2450 vdd.n2449 185
R15172 vdd.n2448 vdd.n2447 185
R15173 vdd.n2446 vdd.n2445 185
R15174 vdd.n2444 vdd.n2443 185
R15175 vdd.n2442 vdd.n2441 185
R15176 vdd.n2440 vdd.n2439 185
R15177 vdd.n2438 vdd.n2437 185
R15178 vdd.n2436 vdd.n2435 185
R15179 vdd.n2434 vdd.n2433 185
R15180 vdd.n2432 vdd.n2431 185
R15181 vdd.n2430 vdd.n2429 185
R15182 vdd.n2428 vdd.n2427 185
R15183 vdd.n2426 vdd.n2425 185
R15184 vdd.n2424 vdd.n2423 185
R15185 vdd.n2422 vdd.n2421 185
R15186 vdd.n2420 vdd.n2419 185
R15187 vdd.n2418 vdd.n2417 185
R15188 vdd.n2416 vdd.n2415 185
R15189 vdd.n2414 vdd.n2413 185
R15190 vdd.n2412 vdd.n2411 185
R15191 vdd.n2410 vdd.n2409 185
R15192 vdd.n2407 vdd.n2406 185
R15193 vdd.n2405 vdd.n2404 185
R15194 vdd.n2403 vdd.n2402 185
R15195 vdd.n2609 vdd.n2608 185
R15196 vdd.n2611 vdd.n624 185
R15197 vdd.n2613 vdd.n2612 185
R15198 vdd.n2615 vdd.n621 185
R15199 vdd.n2617 vdd.n2616 185
R15200 vdd.n2619 vdd.n619 185
R15201 vdd.n2621 vdd.n2620 185
R15202 vdd.n2622 vdd.n618 185
R15203 vdd.n2624 vdd.n2623 185
R15204 vdd.n2626 vdd.n616 185
R15205 vdd.n2628 vdd.n2627 185
R15206 vdd.n2629 vdd.n615 185
R15207 vdd.n2631 vdd.n2630 185
R15208 vdd.n2633 vdd.n613 185
R15209 vdd.n2635 vdd.n2634 185
R15210 vdd.n2636 vdd.n612 185
R15211 vdd.n2638 vdd.n2637 185
R15212 vdd.n2640 vdd.n520 185
R15213 vdd.n2642 vdd.n2641 185
R15214 vdd.n2644 vdd.n610 185
R15215 vdd.n2646 vdd.n2645 185
R15216 vdd.n2647 vdd.n609 185
R15217 vdd.n2649 vdd.n2648 185
R15218 vdd.n2651 vdd.n607 185
R15219 vdd.n2653 vdd.n2652 185
R15220 vdd.n2654 vdd.n606 185
R15221 vdd.n2656 vdd.n2655 185
R15222 vdd.n2658 vdd.n604 185
R15223 vdd.n2660 vdd.n2659 185
R15224 vdd.n2661 vdd.n603 185
R15225 vdd.n2663 vdd.n2662 185
R15226 vdd.n2665 vdd.n602 185
R15227 vdd.n2666 vdd.n601 185
R15228 vdd.n2669 vdd.n2668 185
R15229 vdd.n2670 vdd.n599 185
R15230 vdd.n599 vdd.n484 185
R15231 vdd.n2607 vdd.n596 185
R15232 vdd.n2673 vdd.n596 185
R15233 vdd.n2606 vdd.n2605 185
R15234 vdd.n2605 vdd.n595 185
R15235 vdd.n2604 vdd.n626 185
R15236 vdd.n2604 vdd.n2603 185
R15237 vdd.n2358 vdd.n627 185
R15238 vdd.n636 vdd.n627 185
R15239 vdd.n2359 vdd.n634 185
R15240 vdd.n2597 vdd.n634 185
R15241 vdd.n2361 vdd.n2360 185
R15242 vdd.n2360 vdd.n633 185
R15243 vdd.n2362 vdd.n642 185
R15244 vdd.n2546 vdd.n642 185
R15245 vdd.n2364 vdd.n2363 185
R15246 vdd.n2363 vdd.n641 185
R15247 vdd.n2365 vdd.n648 185
R15248 vdd.n2540 vdd.n648 185
R15249 vdd.n2367 vdd.n2366 185
R15250 vdd.n2366 vdd.n647 185
R15251 vdd.n2368 vdd.n653 185
R15252 vdd.n2532 vdd.n653 185
R15253 vdd.n2370 vdd.n2369 185
R15254 vdd.n2369 vdd.n660 185
R15255 vdd.n2371 vdd.n658 185
R15256 vdd.n2526 vdd.n658 185
R15257 vdd.n2373 vdd.n2372 185
R15258 vdd.n2374 vdd.n2373 185
R15259 vdd.n2357 vdd.n665 185
R15260 vdd.n2520 vdd.n665 185
R15261 vdd.n2356 vdd.n2355 185
R15262 vdd.n2355 vdd.n664 185
R15263 vdd.n2354 vdd.n671 185
R15264 vdd.n2514 vdd.n671 185
R15265 vdd.n2353 vdd.n2352 185
R15266 vdd.n2352 vdd.n670 185
R15267 vdd.n2351 vdd.n676 185
R15268 vdd.n2508 vdd.n676 185
R15269 vdd.n2350 vdd.n2349 185
R15270 vdd.n2349 vdd.n683 185
R15271 vdd.n2348 vdd.n681 185
R15272 vdd.n2502 vdd.n681 185
R15273 vdd.n2347 vdd.n2346 185
R15274 vdd.n2346 vdd.n690 185
R15275 vdd.n2345 vdd.n688 185
R15276 vdd.n2496 vdd.n688 185
R15277 vdd.n2344 vdd.n2343 185
R15278 vdd.n2343 vdd.n687 185
R15279 vdd.n2255 vdd.n694 185
R15280 vdd.n2490 vdd.n694 185
R15281 vdd.n2397 vdd.n2396 185
R15282 vdd.n2396 vdd.n2395 185
R15283 vdd.n2398 vdd.n699 185
R15284 vdd.n2484 vdd.n699 185
R15285 vdd.n2400 vdd.n2399 185
R15286 vdd.n2399 vdd.t196 185
R15287 vdd.n2401 vdd.n704 185
R15288 vdd.n2478 vdd.n704 185
R15289 vdd.n2480 vdd.n2479 185
R15290 vdd.n2479 vdd.n2478 185
R15291 vdd.n2481 vdd.n701 185
R15292 vdd.n701 vdd.t196 185
R15293 vdd.n2483 vdd.n2482 185
R15294 vdd.n2484 vdd.n2483 185
R15295 vdd.n693 vdd.n692 185
R15296 vdd.n2395 vdd.n693 185
R15297 vdd.n2492 vdd.n2491 185
R15298 vdd.n2491 vdd.n2490 185
R15299 vdd.n2493 vdd.n691 185
R15300 vdd.n691 vdd.n687 185
R15301 vdd.n2495 vdd.n2494 185
R15302 vdd.n2496 vdd.n2495 185
R15303 vdd.n680 vdd.n679 185
R15304 vdd.n690 vdd.n680 185
R15305 vdd.n2504 vdd.n2503 185
R15306 vdd.n2503 vdd.n2502 185
R15307 vdd.n2505 vdd.n678 185
R15308 vdd.n683 vdd.n678 185
R15309 vdd.n2507 vdd.n2506 185
R15310 vdd.n2508 vdd.n2507 185
R15311 vdd.n669 vdd.n668 185
R15312 vdd.n670 vdd.n669 185
R15313 vdd.n2516 vdd.n2515 185
R15314 vdd.n2515 vdd.n2514 185
R15315 vdd.n2517 vdd.n667 185
R15316 vdd.n667 vdd.n664 185
R15317 vdd.n2519 vdd.n2518 185
R15318 vdd.n2520 vdd.n2519 185
R15319 vdd.n657 vdd.n656 185
R15320 vdd.n2374 vdd.n657 185
R15321 vdd.n2528 vdd.n2527 185
R15322 vdd.n2527 vdd.n2526 185
R15323 vdd.n2529 vdd.n655 185
R15324 vdd.n660 vdd.n655 185
R15325 vdd.n2531 vdd.n2530 185
R15326 vdd.n2532 vdd.n2531 185
R15327 vdd.n646 vdd.n645 185
R15328 vdd.n647 vdd.n646 185
R15329 vdd.n2542 vdd.n2541 185
R15330 vdd.n2541 vdd.n2540 185
R15331 vdd.n2543 vdd.n644 185
R15332 vdd.n644 vdd.n641 185
R15333 vdd.n2545 vdd.n2544 185
R15334 vdd.n2546 vdd.n2545 185
R15335 vdd.n632 vdd.n631 185
R15336 vdd.n633 vdd.n632 185
R15337 vdd.n2599 vdd.n2598 185
R15338 vdd.n2598 vdd.n2597 185
R15339 vdd.n2600 vdd.n630 185
R15340 vdd.n636 vdd.n630 185
R15341 vdd.n2602 vdd.n2601 185
R15342 vdd.n2603 vdd.n2602 185
R15343 vdd.n600 vdd.n598 185
R15344 vdd.n598 vdd.n595 185
R15345 vdd.n2672 vdd.n2671 185
R15346 vdd.n2673 vdd.n2672 185
R15347 vdd.n2145 vdd.n2144 185
R15348 vdd.n2146 vdd.n2145 185
R15349 vdd.n754 vdd.n752 185
R15350 vdd.n752 vdd.t19 185
R15351 vdd.n2060 vdd.n761 185
R15352 vdd.n2071 vdd.n761 185
R15353 vdd.n2061 vdd.n770 185
R15354 vdd.n1770 vdd.n770 185
R15355 vdd.n2063 vdd.n2062 185
R15356 vdd.n2064 vdd.n2063 185
R15357 vdd.n2059 vdd.n769 185
R15358 vdd.n769 vdd.n766 185
R15359 vdd.n2058 vdd.n2057 185
R15360 vdd.n2057 vdd.n2056 185
R15361 vdd.n772 vdd.n771 185
R15362 vdd.n773 vdd.n772 185
R15363 vdd.n2049 vdd.n2048 185
R15364 vdd.n2050 vdd.n2049 185
R15365 vdd.n2047 vdd.n782 185
R15366 vdd.n782 vdd.n779 185
R15367 vdd.n2046 vdd.n2045 185
R15368 vdd.n2045 vdd.n2044 185
R15369 vdd.n784 vdd.n783 185
R15370 vdd.n792 vdd.n784 185
R15371 vdd.n2037 vdd.n2036 185
R15372 vdd.n2038 vdd.n2037 185
R15373 vdd.n2035 vdd.n793 185
R15374 vdd.n798 vdd.n793 185
R15375 vdd.n2034 vdd.n2033 185
R15376 vdd.n2033 vdd.n2032 185
R15377 vdd.n795 vdd.n794 185
R15378 vdd.n1871 vdd.n795 185
R15379 vdd.n2025 vdd.n2024 185
R15380 vdd.n2026 vdd.n2025 185
R15381 vdd.n2023 vdd.n805 185
R15382 vdd.n805 vdd.n802 185
R15383 vdd.n2022 vdd.n2021 185
R15384 vdd.n2021 vdd.n2020 185
R15385 vdd.n807 vdd.n806 185
R15386 vdd.n808 vdd.n807 185
R15387 vdd.n2013 vdd.n2012 185
R15388 vdd.n2014 vdd.n2013 185
R15389 vdd.n2010 vdd.n816 185
R15390 vdd.n823 vdd.n816 185
R15391 vdd.n2009 vdd.n2008 185
R15392 vdd.n2008 vdd.n2007 185
R15393 vdd.n819 vdd.n818 185
R15394 vdd.n820 vdd.n819 185
R15395 vdd.n2000 vdd.n1999 185
R15396 vdd.n2001 vdd.n2000 185
R15397 vdd.n1998 vdd.n830 185
R15398 vdd.n830 vdd.n827 185
R15399 vdd.n1997 vdd.n1996 185
R15400 vdd.n1996 vdd.n1995 185
R15401 vdd.n832 vdd.n831 185
R15402 vdd.n833 vdd.n832 185
R15403 vdd.n1988 vdd.n1987 185
R15404 vdd.n1989 vdd.n1988 185
R15405 vdd.n2076 vdd.n726 185
R15406 vdd.n2218 vdd.n726 185
R15407 vdd.n2078 vdd.n2077 185
R15408 vdd.n2080 vdd.n2079 185
R15409 vdd.n2082 vdd.n2081 185
R15410 vdd.n2084 vdd.n2083 185
R15411 vdd.n2086 vdd.n2085 185
R15412 vdd.n2088 vdd.n2087 185
R15413 vdd.n2090 vdd.n2089 185
R15414 vdd.n2092 vdd.n2091 185
R15415 vdd.n2094 vdd.n2093 185
R15416 vdd.n2096 vdd.n2095 185
R15417 vdd.n2098 vdd.n2097 185
R15418 vdd.n2100 vdd.n2099 185
R15419 vdd.n2102 vdd.n2101 185
R15420 vdd.n2104 vdd.n2103 185
R15421 vdd.n2106 vdd.n2105 185
R15422 vdd.n2108 vdd.n2107 185
R15423 vdd.n2110 vdd.n2109 185
R15424 vdd.n2112 vdd.n2111 185
R15425 vdd.n2114 vdd.n2113 185
R15426 vdd.n2116 vdd.n2115 185
R15427 vdd.n2118 vdd.n2117 185
R15428 vdd.n2120 vdd.n2119 185
R15429 vdd.n2122 vdd.n2121 185
R15430 vdd.n2124 vdd.n2123 185
R15431 vdd.n2126 vdd.n2125 185
R15432 vdd.n2128 vdd.n2127 185
R15433 vdd.n2130 vdd.n2129 185
R15434 vdd.n2132 vdd.n2131 185
R15435 vdd.n2134 vdd.n2133 185
R15436 vdd.n2136 vdd.n2135 185
R15437 vdd.n2138 vdd.n2137 185
R15438 vdd.n2140 vdd.n2139 185
R15439 vdd.n2142 vdd.n2141 185
R15440 vdd.n2143 vdd.n753 185
R15441 vdd.n2075 vdd.n751 185
R15442 vdd.n2146 vdd.n751 185
R15443 vdd.n2074 vdd.n2073 185
R15444 vdd.n2073 vdd.t19 185
R15445 vdd.n2072 vdd.n758 185
R15446 vdd.n2072 vdd.n2071 185
R15447 vdd.n1852 vdd.n759 185
R15448 vdd.n1770 vdd.n759 185
R15449 vdd.n1853 vdd.n768 185
R15450 vdd.n2064 vdd.n768 185
R15451 vdd.n1855 vdd.n1854 185
R15452 vdd.n1854 vdd.n766 185
R15453 vdd.n1856 vdd.n775 185
R15454 vdd.n2056 vdd.n775 185
R15455 vdd.n1858 vdd.n1857 185
R15456 vdd.n1857 vdd.n773 185
R15457 vdd.n1859 vdd.n781 185
R15458 vdd.n2050 vdd.n781 185
R15459 vdd.n1861 vdd.n1860 185
R15460 vdd.n1860 vdd.n779 185
R15461 vdd.n1862 vdd.n786 185
R15462 vdd.n2044 vdd.n786 185
R15463 vdd.n1864 vdd.n1863 185
R15464 vdd.n1863 vdd.n792 185
R15465 vdd.n1865 vdd.n791 185
R15466 vdd.n2038 vdd.n791 185
R15467 vdd.n1867 vdd.n1866 185
R15468 vdd.n1866 vdd.n798 185
R15469 vdd.n1868 vdd.n797 185
R15470 vdd.n2032 vdd.n797 185
R15471 vdd.n1870 vdd.n1869 185
R15472 vdd.n1871 vdd.n1870 185
R15473 vdd.n1851 vdd.n804 185
R15474 vdd.n2026 vdd.n804 185
R15475 vdd.n1850 vdd.n1849 185
R15476 vdd.n1849 vdd.n802 185
R15477 vdd.n1848 vdd.n810 185
R15478 vdd.n2020 vdd.n810 185
R15479 vdd.n1847 vdd.n1846 185
R15480 vdd.n1846 vdd.n808 185
R15481 vdd.n1845 vdd.n815 185
R15482 vdd.n2014 vdd.n815 185
R15483 vdd.n1844 vdd.n1843 185
R15484 vdd.n1843 vdd.n823 185
R15485 vdd.n1842 vdd.n822 185
R15486 vdd.n2007 vdd.n822 185
R15487 vdd.n1841 vdd.n1840 185
R15488 vdd.n1840 vdd.n820 185
R15489 vdd.n1839 vdd.n829 185
R15490 vdd.n2001 vdd.n829 185
R15491 vdd.n1838 vdd.n1837 185
R15492 vdd.n1837 vdd.n827 185
R15493 vdd.n1836 vdd.n835 185
R15494 vdd.n1995 vdd.n835 185
R15495 vdd.n1835 vdd.n1834 185
R15496 vdd.n1834 vdd.n833 185
R15497 vdd.n1833 vdd.n841 185
R15498 vdd.n1989 vdd.n841 185
R15499 vdd.n1986 vdd.n842 185
R15500 vdd.n1985 vdd.n1984 185
R15501 vdd.n1982 vdd.n843 185
R15502 vdd.n1980 vdd.n1979 185
R15503 vdd.n1978 vdd.n844 185
R15504 vdd.n1977 vdd.n1976 185
R15505 vdd.n1974 vdd.n845 185
R15506 vdd.n1972 vdd.n1971 185
R15507 vdd.n1970 vdd.n846 185
R15508 vdd.n1969 vdd.n1968 185
R15509 vdd.n1966 vdd.n847 185
R15510 vdd.n1964 vdd.n1963 185
R15511 vdd.n1962 vdd.n848 185
R15512 vdd.n1961 vdd.n1960 185
R15513 vdd.n1958 vdd.n849 185
R15514 vdd.n1956 vdd.n1955 185
R15515 vdd.n1954 vdd.n850 185
R15516 vdd.n1953 vdd.n852 185
R15517 vdd.n1798 vdd.n853 185
R15518 vdd.n1801 vdd.n1800 185
R15519 vdd.n1803 vdd.n1802 185
R15520 vdd.n1805 vdd.n1797 185
R15521 vdd.n1808 vdd.n1807 185
R15522 vdd.n1809 vdd.n1796 185
R15523 vdd.n1811 vdd.n1810 185
R15524 vdd.n1813 vdd.n1795 185
R15525 vdd.n1816 vdd.n1815 185
R15526 vdd.n1817 vdd.n1794 185
R15527 vdd.n1819 vdd.n1818 185
R15528 vdd.n1821 vdd.n1793 185
R15529 vdd.n1824 vdd.n1823 185
R15530 vdd.n1825 vdd.n1790 185
R15531 vdd.n1828 vdd.n1827 185
R15532 vdd.n1830 vdd.n1789 185
R15533 vdd.n1832 vdd.n1831 185
R15534 vdd.n1831 vdd.n839 185
R15535 vdd.n291 vdd.n290 171.744
R15536 vdd.n290 vdd.n289 171.744
R15537 vdd.n289 vdd.n258 171.744
R15538 vdd.n282 vdd.n258 171.744
R15539 vdd.n282 vdd.n281 171.744
R15540 vdd.n281 vdd.n263 171.744
R15541 vdd.n274 vdd.n263 171.744
R15542 vdd.n274 vdd.n273 171.744
R15543 vdd.n273 vdd.n267 171.744
R15544 vdd.n244 vdd.n243 171.744
R15545 vdd.n243 vdd.n242 171.744
R15546 vdd.n242 vdd.n211 171.744
R15547 vdd.n235 vdd.n211 171.744
R15548 vdd.n235 vdd.n234 171.744
R15549 vdd.n234 vdd.n216 171.744
R15550 vdd.n227 vdd.n216 171.744
R15551 vdd.n227 vdd.n226 171.744
R15552 vdd.n226 vdd.n220 171.744
R15553 vdd.n201 vdd.n200 171.744
R15554 vdd.n200 vdd.n199 171.744
R15555 vdd.n199 vdd.n168 171.744
R15556 vdd.n192 vdd.n168 171.744
R15557 vdd.n192 vdd.n191 171.744
R15558 vdd.n191 vdd.n173 171.744
R15559 vdd.n184 vdd.n173 171.744
R15560 vdd.n184 vdd.n183 171.744
R15561 vdd.n183 vdd.n177 171.744
R15562 vdd.n154 vdd.n153 171.744
R15563 vdd.n153 vdd.n152 171.744
R15564 vdd.n152 vdd.n121 171.744
R15565 vdd.n145 vdd.n121 171.744
R15566 vdd.n145 vdd.n144 171.744
R15567 vdd.n144 vdd.n126 171.744
R15568 vdd.n137 vdd.n126 171.744
R15569 vdd.n137 vdd.n136 171.744
R15570 vdd.n136 vdd.n130 171.744
R15571 vdd.n112 vdd.n111 171.744
R15572 vdd.n111 vdd.n110 171.744
R15573 vdd.n110 vdd.n79 171.744
R15574 vdd.n103 vdd.n79 171.744
R15575 vdd.n103 vdd.n102 171.744
R15576 vdd.n102 vdd.n84 171.744
R15577 vdd.n95 vdd.n84 171.744
R15578 vdd.n95 vdd.n94 171.744
R15579 vdd.n94 vdd.n88 171.744
R15580 vdd.n65 vdd.n64 171.744
R15581 vdd.n64 vdd.n63 171.744
R15582 vdd.n63 vdd.n32 171.744
R15583 vdd.n56 vdd.n32 171.744
R15584 vdd.n56 vdd.n55 171.744
R15585 vdd.n55 vdd.n37 171.744
R15586 vdd.n48 vdd.n37 171.744
R15587 vdd.n48 vdd.n47 171.744
R15588 vdd.n47 vdd.n41 171.744
R15589 vdd.n1106 vdd.n1105 171.744
R15590 vdd.n1105 vdd.n1104 171.744
R15591 vdd.n1104 vdd.n1073 171.744
R15592 vdd.n1097 vdd.n1073 171.744
R15593 vdd.n1097 vdd.n1096 171.744
R15594 vdd.n1096 vdd.n1078 171.744
R15595 vdd.n1089 vdd.n1078 171.744
R15596 vdd.n1089 vdd.n1088 171.744
R15597 vdd.n1088 vdd.n1082 171.744
R15598 vdd.n1153 vdd.n1152 171.744
R15599 vdd.n1152 vdd.n1151 171.744
R15600 vdd.n1151 vdd.n1120 171.744
R15601 vdd.n1144 vdd.n1120 171.744
R15602 vdd.n1144 vdd.n1143 171.744
R15603 vdd.n1143 vdd.n1125 171.744
R15604 vdd.n1136 vdd.n1125 171.744
R15605 vdd.n1136 vdd.n1135 171.744
R15606 vdd.n1135 vdd.n1129 171.744
R15607 vdd.n1016 vdd.n1015 171.744
R15608 vdd.n1015 vdd.n1014 171.744
R15609 vdd.n1014 vdd.n983 171.744
R15610 vdd.n1007 vdd.n983 171.744
R15611 vdd.n1007 vdd.n1006 171.744
R15612 vdd.n1006 vdd.n988 171.744
R15613 vdd.n999 vdd.n988 171.744
R15614 vdd.n999 vdd.n998 171.744
R15615 vdd.n998 vdd.n992 171.744
R15616 vdd.n1063 vdd.n1062 171.744
R15617 vdd.n1062 vdd.n1061 171.744
R15618 vdd.n1061 vdd.n1030 171.744
R15619 vdd.n1054 vdd.n1030 171.744
R15620 vdd.n1054 vdd.n1053 171.744
R15621 vdd.n1053 vdd.n1035 171.744
R15622 vdd.n1046 vdd.n1035 171.744
R15623 vdd.n1046 vdd.n1045 171.744
R15624 vdd.n1045 vdd.n1039 171.744
R15625 vdd.n927 vdd.n926 171.744
R15626 vdd.n926 vdd.n925 171.744
R15627 vdd.n925 vdd.n894 171.744
R15628 vdd.n918 vdd.n894 171.744
R15629 vdd.n918 vdd.n917 171.744
R15630 vdd.n917 vdd.n899 171.744
R15631 vdd.n910 vdd.n899 171.744
R15632 vdd.n910 vdd.n909 171.744
R15633 vdd.n909 vdd.n903 171.744
R15634 vdd.n974 vdd.n973 171.744
R15635 vdd.n973 vdd.n972 171.744
R15636 vdd.n972 vdd.n941 171.744
R15637 vdd.n965 vdd.n941 171.744
R15638 vdd.n965 vdd.n964 171.744
R15639 vdd.n964 vdd.n946 171.744
R15640 vdd.n957 vdd.n946 171.744
R15641 vdd.n957 vdd.n956 171.744
R15642 vdd.n956 vdd.n950 171.744
R15643 vdd.n3017 vdd.n334 146.341
R15644 vdd.n3015 vdd.n3014 146.341
R15645 vdd.n3012 vdd.n338 146.341
R15646 vdd.n3008 vdd.n3007 146.341
R15647 vdd.n3005 vdd.n346 146.341
R15648 vdd.n3001 vdd.n3000 146.341
R15649 vdd.n2998 vdd.n353 146.341
R15650 vdd.n2994 vdd.n2993 146.341
R15651 vdd.n2991 vdd.n360 146.341
R15652 vdd.n371 vdd.n368 146.341
R15653 vdd.n2983 vdd.n2982 146.341
R15654 vdd.n2980 vdd.n373 146.341
R15655 vdd.n2976 vdd.n2975 146.341
R15656 vdd.n2973 vdd.n379 146.341
R15657 vdd.n2969 vdd.n2968 146.341
R15658 vdd.n2966 vdd.n386 146.341
R15659 vdd.n2962 vdd.n2961 146.341
R15660 vdd.n2959 vdd.n393 146.341
R15661 vdd.n2955 vdd.n2954 146.341
R15662 vdd.n2952 vdd.n400 146.341
R15663 vdd.n411 vdd.n408 146.341
R15664 vdd.n2944 vdd.n2943 146.341
R15665 vdd.n2941 vdd.n413 146.341
R15666 vdd.n2937 vdd.n2936 146.341
R15667 vdd.n2934 vdd.n419 146.341
R15668 vdd.n2930 vdd.n2929 146.341
R15669 vdd.n2927 vdd.n426 146.341
R15670 vdd.n2923 vdd.n2922 146.341
R15671 vdd.n2920 vdd.n433 146.341
R15672 vdd.n2916 vdd.n2915 146.341
R15673 vdd.n2913 vdd.n440 146.341
R15674 vdd.n2850 vdd.n478 146.341
R15675 vdd.n2850 vdd.n474 146.341
R15676 vdd.n2856 vdd.n474 146.341
R15677 vdd.n2856 vdd.n466 146.341
R15678 vdd.n2867 vdd.n466 146.341
R15679 vdd.n2867 vdd.n462 146.341
R15680 vdd.n2873 vdd.n462 146.341
R15681 vdd.n2873 vdd.n454 146.341
R15682 vdd.n2883 vdd.n454 146.341
R15683 vdd.n2883 vdd.n455 146.341
R15684 vdd.n455 vdd.n305 146.341
R15685 vdd.n306 vdd.n305 146.341
R15686 vdd.n307 vdd.n306 146.341
R15687 vdd.n448 vdd.n307 146.341
R15688 vdd.n448 vdd.n315 146.341
R15689 vdd.n316 vdd.n315 146.341
R15690 vdd.n317 vdd.n316 146.341
R15691 vdd.n445 vdd.n317 146.341
R15692 vdd.n445 vdd.n326 146.341
R15693 vdd.n327 vdd.n326 146.341
R15694 vdd.n328 vdd.n327 146.341
R15695 vdd.n2839 vdd.n483 146.341
R15696 vdd.n2839 vdd.n517 146.341
R15697 vdd.n523 vdd.n522 146.341
R15698 vdd.n2832 vdd.n2831 146.341
R15699 vdd.n2828 vdd.n2827 146.341
R15700 vdd.n2824 vdd.n2823 146.341
R15701 vdd.n2820 vdd.n2819 146.341
R15702 vdd.n2816 vdd.n2815 146.341
R15703 vdd.n2812 vdd.n2811 146.341
R15704 vdd.n2808 vdd.n2807 146.341
R15705 vdd.n2799 vdd.n2798 146.341
R15706 vdd.n2796 vdd.n2795 146.341
R15707 vdd.n2792 vdd.n2791 146.341
R15708 vdd.n2788 vdd.n2787 146.341
R15709 vdd.n2784 vdd.n2783 146.341
R15710 vdd.n2780 vdd.n2779 146.341
R15711 vdd.n2776 vdd.n2775 146.341
R15712 vdd.n2772 vdd.n2771 146.341
R15713 vdd.n2768 vdd.n2767 146.341
R15714 vdd.n2764 vdd.n2763 146.341
R15715 vdd.n2760 vdd.n2759 146.341
R15716 vdd.n2753 vdd.n2752 146.341
R15717 vdd.n2750 vdd.n2749 146.341
R15718 vdd.n2746 vdd.n2745 146.341
R15719 vdd.n2742 vdd.n2741 146.341
R15720 vdd.n2738 vdd.n2737 146.341
R15721 vdd.n2734 vdd.n2733 146.341
R15722 vdd.n2730 vdd.n2729 146.341
R15723 vdd.n2726 vdd.n2725 146.341
R15724 vdd.n2722 vdd.n2721 146.341
R15725 vdd.n2718 vdd.n2717 146.341
R15726 vdd.n2714 vdd.n515 146.341
R15727 vdd.n2848 vdd.n479 146.341
R15728 vdd.n2848 vdd.n472 146.341
R15729 vdd.n2859 vdd.n472 146.341
R15730 vdd.n2859 vdd.n468 146.341
R15731 vdd.n2865 vdd.n468 146.341
R15732 vdd.n2865 vdd.n461 146.341
R15733 vdd.n2875 vdd.n461 146.341
R15734 vdd.n2875 vdd.n457 146.341
R15735 vdd.n2881 vdd.n457 146.341
R15736 vdd.n2881 vdd.n302 146.341
R15737 vdd.n3044 vdd.n302 146.341
R15738 vdd.n3044 vdd.n303 146.341
R15739 vdd.n3040 vdd.n303 146.341
R15740 vdd.n3040 vdd.n309 146.341
R15741 vdd.n3036 vdd.n309 146.341
R15742 vdd.n3036 vdd.n314 146.341
R15743 vdd.n3032 vdd.n314 146.341
R15744 vdd.n3032 vdd.n319 146.341
R15745 vdd.n3028 vdd.n319 146.341
R15746 vdd.n3028 vdd.n325 146.341
R15747 vdd.n3024 vdd.n325 146.341
R15748 vdd.n1936 vdd.n1935 146.341
R15749 vdd.n1933 vdd.n1517 146.341
R15750 vdd.n1713 vdd.n1523 146.341
R15751 vdd.n1711 vdd.n1710 146.341
R15752 vdd.n1708 vdd.n1525 146.341
R15753 vdd.n1704 vdd.n1703 146.341
R15754 vdd.n1701 vdd.n1532 146.341
R15755 vdd.n1697 vdd.n1696 146.341
R15756 vdd.n1694 vdd.n1539 146.341
R15757 vdd.n1550 vdd.n1547 146.341
R15758 vdd.n1686 vdd.n1685 146.341
R15759 vdd.n1683 vdd.n1552 146.341
R15760 vdd.n1679 vdd.n1678 146.341
R15761 vdd.n1676 vdd.n1558 146.341
R15762 vdd.n1672 vdd.n1671 146.341
R15763 vdd.n1669 vdd.n1565 146.341
R15764 vdd.n1665 vdd.n1664 146.341
R15765 vdd.n1662 vdd.n1572 146.341
R15766 vdd.n1658 vdd.n1657 146.341
R15767 vdd.n1655 vdd.n1579 146.341
R15768 vdd.n1590 vdd.n1587 146.341
R15769 vdd.n1647 vdd.n1646 146.341
R15770 vdd.n1644 vdd.n1592 146.341
R15771 vdd.n1640 vdd.n1639 146.341
R15772 vdd.n1637 vdd.n1598 146.341
R15773 vdd.n1633 vdd.n1632 146.341
R15774 vdd.n1630 vdd.n1605 146.341
R15775 vdd.n1626 vdd.n1625 146.341
R15776 vdd.n1623 vdd.n1620 146.341
R15777 vdd.n1618 vdd.n1615 146.341
R15778 vdd.n1613 vdd.n859 146.341
R15779 vdd.n1431 vdd.n1191 146.341
R15780 vdd.n1431 vdd.n1187 146.341
R15781 vdd.n1437 vdd.n1187 146.341
R15782 vdd.n1437 vdd.n1179 146.341
R15783 vdd.n1448 vdd.n1179 146.341
R15784 vdd.n1448 vdd.n1175 146.341
R15785 vdd.n1454 vdd.n1175 146.341
R15786 vdd.n1454 vdd.n1169 146.341
R15787 vdd.n1466 vdd.n1169 146.341
R15788 vdd.n1466 vdd.n1165 146.341
R15789 vdd.n1472 vdd.n1165 146.341
R15790 vdd.n1472 vdd.n886 146.341
R15791 vdd.n1482 vdd.n886 146.341
R15792 vdd.n1482 vdd.n882 146.341
R15793 vdd.n1488 vdd.n882 146.341
R15794 vdd.n1488 vdd.n876 146.341
R15795 vdd.n1499 vdd.n876 146.341
R15796 vdd.n1499 vdd.n871 146.341
R15797 vdd.n1507 vdd.n871 146.341
R15798 vdd.n1507 vdd.n861 146.341
R15799 vdd.n1944 vdd.n861 146.341
R15800 vdd.n1420 vdd.n1196 146.341
R15801 vdd.n1420 vdd.n1229 146.341
R15802 vdd.n1233 vdd.n1232 146.341
R15803 vdd.n1235 vdd.n1234 146.341
R15804 vdd.n1239 vdd.n1238 146.341
R15805 vdd.n1241 vdd.n1240 146.341
R15806 vdd.n1245 vdd.n1244 146.341
R15807 vdd.n1247 vdd.n1246 146.341
R15808 vdd.n1251 vdd.n1250 146.341
R15809 vdd.n1253 vdd.n1252 146.341
R15810 vdd.n1259 vdd.n1258 146.341
R15811 vdd.n1261 vdd.n1260 146.341
R15812 vdd.n1265 vdd.n1264 146.341
R15813 vdd.n1267 vdd.n1266 146.341
R15814 vdd.n1271 vdd.n1270 146.341
R15815 vdd.n1273 vdd.n1272 146.341
R15816 vdd.n1277 vdd.n1276 146.341
R15817 vdd.n1279 vdd.n1278 146.341
R15818 vdd.n1283 vdd.n1282 146.341
R15819 vdd.n1285 vdd.n1284 146.341
R15820 vdd.n1357 vdd.n1288 146.341
R15821 vdd.n1290 vdd.n1289 146.341
R15822 vdd.n1294 vdd.n1293 146.341
R15823 vdd.n1296 vdd.n1295 146.341
R15824 vdd.n1300 vdd.n1299 146.341
R15825 vdd.n1302 vdd.n1301 146.341
R15826 vdd.n1306 vdd.n1305 146.341
R15827 vdd.n1308 vdd.n1307 146.341
R15828 vdd.n1312 vdd.n1311 146.341
R15829 vdd.n1314 vdd.n1313 146.341
R15830 vdd.n1318 vdd.n1317 146.341
R15831 vdd.n1319 vdd.n1227 146.341
R15832 vdd.n1429 vdd.n1192 146.341
R15833 vdd.n1429 vdd.n1185 146.341
R15834 vdd.n1440 vdd.n1185 146.341
R15835 vdd.n1440 vdd.n1181 146.341
R15836 vdd.n1446 vdd.n1181 146.341
R15837 vdd.n1446 vdd.n1174 146.341
R15838 vdd.n1457 vdd.n1174 146.341
R15839 vdd.n1457 vdd.n1170 146.341
R15840 vdd.n1464 vdd.n1170 146.341
R15841 vdd.n1464 vdd.n1163 146.341
R15842 vdd.n1474 vdd.n1163 146.341
R15843 vdd.n1474 vdd.n889 146.341
R15844 vdd.n1480 vdd.n889 146.341
R15845 vdd.n1480 vdd.n881 146.341
R15846 vdd.n1491 vdd.n881 146.341
R15847 vdd.n1491 vdd.n877 146.341
R15848 vdd.n1497 vdd.n877 146.341
R15849 vdd.n1497 vdd.n869 146.341
R15850 vdd.n1510 vdd.n869 146.341
R15851 vdd.n1510 vdd.n864 146.341
R15852 vdd.n1942 vdd.n864 146.341
R15853 vdd.n863 vdd.n839 141.707
R15854 vdd.n2840 vdd.n484 141.707
R15855 vdd.n1791 vdd.t71 127.284
R15856 vdd.n755 vdd.t55 127.284
R15857 vdd.n1765 vdd.t96 127.284
R15858 vdd.n747 vdd.t86 127.284
R15859 vdd.n2536 vdd.t38 127.284
R15860 vdd.n2536 vdd.t39 127.284
R15861 vdd.n2256 vdd.t78 127.284
R15862 vdd.n622 vdd.t59 127.284
R15863 vdd.n2253 vdd.t64 127.284
R15864 vdd.n589 vdd.t66 127.284
R15865 vdd.n817 vdd.t74 127.284
R15866 vdd.n817 vdd.t75 127.284
R15867 vdd.n22 vdd.n20 117.314
R15868 vdd.n17 vdd.n15 117.314
R15869 vdd.n27 vdd.n26 116.927
R15870 vdd.n24 vdd.n23 116.927
R15871 vdd.n22 vdd.n21 116.927
R15872 vdd.n17 vdd.n16 116.927
R15873 vdd.n19 vdd.n18 116.927
R15874 vdd.n27 vdd.n25 116.927
R15875 vdd.n1792 vdd.t70 111.188
R15876 vdd.n756 vdd.t56 111.188
R15877 vdd.n1766 vdd.t95 111.188
R15878 vdd.n748 vdd.t87 111.188
R15879 vdd.n2257 vdd.t77 111.188
R15880 vdd.n623 vdd.t60 111.188
R15881 vdd.n2254 vdd.t63 111.188
R15882 vdd.n590 vdd.t67 111.188
R15883 vdd.n2479 vdd.n701 99.5127
R15884 vdd.n2483 vdd.n701 99.5127
R15885 vdd.n2483 vdd.n693 99.5127
R15886 vdd.n2491 vdd.n693 99.5127
R15887 vdd.n2491 vdd.n691 99.5127
R15888 vdd.n2495 vdd.n691 99.5127
R15889 vdd.n2495 vdd.n680 99.5127
R15890 vdd.n2503 vdd.n680 99.5127
R15891 vdd.n2503 vdd.n678 99.5127
R15892 vdd.n2507 vdd.n678 99.5127
R15893 vdd.n2507 vdd.n669 99.5127
R15894 vdd.n2515 vdd.n669 99.5127
R15895 vdd.n2515 vdd.n667 99.5127
R15896 vdd.n2519 vdd.n667 99.5127
R15897 vdd.n2519 vdd.n657 99.5127
R15898 vdd.n2527 vdd.n657 99.5127
R15899 vdd.n2527 vdd.n655 99.5127
R15900 vdd.n2531 vdd.n655 99.5127
R15901 vdd.n2531 vdd.n646 99.5127
R15902 vdd.n2541 vdd.n646 99.5127
R15903 vdd.n2541 vdd.n644 99.5127
R15904 vdd.n2545 vdd.n644 99.5127
R15905 vdd.n2545 vdd.n632 99.5127
R15906 vdd.n2598 vdd.n632 99.5127
R15907 vdd.n2598 vdd.n630 99.5127
R15908 vdd.n2602 vdd.n630 99.5127
R15909 vdd.n2602 vdd.n598 99.5127
R15910 vdd.n2672 vdd.n598 99.5127
R15911 vdd.n2668 vdd.n599 99.5127
R15912 vdd.n2666 vdd.n2665 99.5127
R15913 vdd.n2663 vdd.n603 99.5127
R15914 vdd.n2659 vdd.n2658 99.5127
R15915 vdd.n2656 vdd.n606 99.5127
R15916 vdd.n2652 vdd.n2651 99.5127
R15917 vdd.n2649 vdd.n609 99.5127
R15918 vdd.n2645 vdd.n2644 99.5127
R15919 vdd.n2642 vdd.n2640 99.5127
R15920 vdd.n2638 vdd.n612 99.5127
R15921 vdd.n2634 vdd.n2633 99.5127
R15922 vdd.n2631 vdd.n615 99.5127
R15923 vdd.n2627 vdd.n2626 99.5127
R15924 vdd.n2624 vdd.n618 99.5127
R15925 vdd.n2620 vdd.n2619 99.5127
R15926 vdd.n2617 vdd.n621 99.5127
R15927 vdd.n2612 vdd.n2611 99.5127
R15928 vdd.n2399 vdd.n704 99.5127
R15929 vdd.n2399 vdd.n699 99.5127
R15930 vdd.n2396 vdd.n699 99.5127
R15931 vdd.n2396 vdd.n694 99.5127
R15932 vdd.n2343 vdd.n694 99.5127
R15933 vdd.n2343 vdd.n688 99.5127
R15934 vdd.n2346 vdd.n688 99.5127
R15935 vdd.n2346 vdd.n681 99.5127
R15936 vdd.n2349 vdd.n681 99.5127
R15937 vdd.n2349 vdd.n676 99.5127
R15938 vdd.n2352 vdd.n676 99.5127
R15939 vdd.n2352 vdd.n671 99.5127
R15940 vdd.n2355 vdd.n671 99.5127
R15941 vdd.n2355 vdd.n665 99.5127
R15942 vdd.n2373 vdd.n665 99.5127
R15943 vdd.n2373 vdd.n658 99.5127
R15944 vdd.n2369 vdd.n658 99.5127
R15945 vdd.n2369 vdd.n653 99.5127
R15946 vdd.n2366 vdd.n653 99.5127
R15947 vdd.n2366 vdd.n648 99.5127
R15948 vdd.n2363 vdd.n648 99.5127
R15949 vdd.n2363 vdd.n642 99.5127
R15950 vdd.n2360 vdd.n642 99.5127
R15951 vdd.n2360 vdd.n634 99.5127
R15952 vdd.n634 vdd.n627 99.5127
R15953 vdd.n2604 vdd.n627 99.5127
R15954 vdd.n2605 vdd.n2604 99.5127
R15955 vdd.n2605 vdd.n596 99.5127
R15956 vdd.n2469 vdd.n2252 99.5127
R15957 vdd.n2465 vdd.n2252 99.5127
R15958 vdd.n2463 vdd.n2462 99.5127
R15959 vdd.n2459 vdd.n2458 99.5127
R15960 vdd.n2455 vdd.n2454 99.5127
R15961 vdd.n2451 vdd.n2450 99.5127
R15962 vdd.n2447 vdd.n2446 99.5127
R15963 vdd.n2443 vdd.n2442 99.5127
R15964 vdd.n2439 vdd.n2438 99.5127
R15965 vdd.n2435 vdd.n2434 99.5127
R15966 vdd.n2431 vdd.n2430 99.5127
R15967 vdd.n2427 vdd.n2426 99.5127
R15968 vdd.n2423 vdd.n2422 99.5127
R15969 vdd.n2419 vdd.n2418 99.5127
R15970 vdd.n2415 vdd.n2414 99.5127
R15971 vdd.n2411 vdd.n2410 99.5127
R15972 vdd.n2406 vdd.n2405 99.5127
R15973 vdd.n2217 vdd.n745 99.5127
R15974 vdd.n2213 vdd.n2212 99.5127
R15975 vdd.n2209 vdd.n2208 99.5127
R15976 vdd.n2205 vdd.n2204 99.5127
R15977 vdd.n2201 vdd.n2200 99.5127
R15978 vdd.n2197 vdd.n2196 99.5127
R15979 vdd.n2193 vdd.n2192 99.5127
R15980 vdd.n2189 vdd.n2188 99.5127
R15981 vdd.n2185 vdd.n2184 99.5127
R15982 vdd.n2181 vdd.n2180 99.5127
R15983 vdd.n2177 vdd.n2176 99.5127
R15984 vdd.n2173 vdd.n2172 99.5127
R15985 vdd.n2169 vdd.n2168 99.5127
R15986 vdd.n2165 vdd.n2164 99.5127
R15987 vdd.n2161 vdd.n2160 99.5127
R15988 vdd.n2157 vdd.n2156 99.5127
R15989 vdd.n2152 vdd.n2151 99.5127
R15990 vdd.n1890 vdd.n840 99.5127
R15991 vdd.n1890 vdd.n834 99.5127
R15992 vdd.n1887 vdd.n834 99.5127
R15993 vdd.n1887 vdd.n828 99.5127
R15994 vdd.n1884 vdd.n828 99.5127
R15995 vdd.n1884 vdd.n821 99.5127
R15996 vdd.n1881 vdd.n821 99.5127
R15997 vdd.n1881 vdd.n814 99.5127
R15998 vdd.n1878 vdd.n814 99.5127
R15999 vdd.n1878 vdd.n809 99.5127
R16000 vdd.n1875 vdd.n809 99.5127
R16001 vdd.n1875 vdd.n803 99.5127
R16002 vdd.n1872 vdd.n803 99.5127
R16003 vdd.n1872 vdd.n796 99.5127
R16004 vdd.n1786 vdd.n796 99.5127
R16005 vdd.n1786 vdd.n790 99.5127
R16006 vdd.n1783 vdd.n790 99.5127
R16007 vdd.n1783 vdd.n785 99.5127
R16008 vdd.n1780 vdd.n785 99.5127
R16009 vdd.n1780 vdd.n780 99.5127
R16010 vdd.n1777 vdd.n780 99.5127
R16011 vdd.n1777 vdd.n774 99.5127
R16012 vdd.n1774 vdd.n774 99.5127
R16013 vdd.n1774 vdd.n767 99.5127
R16014 vdd.n1771 vdd.n767 99.5127
R16015 vdd.n1771 vdd.n760 99.5127
R16016 vdd.n760 vdd.n750 99.5127
R16017 vdd.n2147 vdd.n750 99.5127
R16018 vdd.n1725 vdd.n1723 99.5127
R16019 vdd.n1729 vdd.n1723 99.5127
R16020 vdd.n1733 vdd.n1731 99.5127
R16021 vdd.n1737 vdd.n1721 99.5127
R16022 vdd.n1741 vdd.n1739 99.5127
R16023 vdd.n1745 vdd.n1719 99.5127
R16024 vdd.n1749 vdd.n1747 99.5127
R16025 vdd.n1753 vdd.n1717 99.5127
R16026 vdd.n1756 vdd.n1755 99.5127
R16027 vdd.n1926 vdd.n1924 99.5127
R16028 vdd.n1922 vdd.n1758 99.5127
R16029 vdd.n1918 vdd.n1916 99.5127
R16030 vdd.n1914 vdd.n1760 99.5127
R16031 vdd.n1910 vdd.n1908 99.5127
R16032 vdd.n1906 vdd.n1762 99.5127
R16033 vdd.n1902 vdd.n1900 99.5127
R16034 vdd.n1898 vdd.n1764 99.5127
R16035 vdd.n1990 vdd.n836 99.5127
R16036 vdd.n1994 vdd.n836 99.5127
R16037 vdd.n1994 vdd.n826 99.5127
R16038 vdd.n2002 vdd.n826 99.5127
R16039 vdd.n2002 vdd.n824 99.5127
R16040 vdd.n2006 vdd.n824 99.5127
R16041 vdd.n2006 vdd.n813 99.5127
R16042 vdd.n2015 vdd.n813 99.5127
R16043 vdd.n2015 vdd.n811 99.5127
R16044 vdd.n2019 vdd.n811 99.5127
R16045 vdd.n2019 vdd.n801 99.5127
R16046 vdd.n2027 vdd.n801 99.5127
R16047 vdd.n2027 vdd.n799 99.5127
R16048 vdd.n2031 vdd.n799 99.5127
R16049 vdd.n2031 vdd.n789 99.5127
R16050 vdd.n2039 vdd.n789 99.5127
R16051 vdd.n2039 vdd.n787 99.5127
R16052 vdd.n2043 vdd.n787 99.5127
R16053 vdd.n2043 vdd.n778 99.5127
R16054 vdd.n2051 vdd.n778 99.5127
R16055 vdd.n2051 vdd.n776 99.5127
R16056 vdd.n2055 vdd.n776 99.5127
R16057 vdd.n2055 vdd.n765 99.5127
R16058 vdd.n2065 vdd.n765 99.5127
R16059 vdd.n2065 vdd.n762 99.5127
R16060 vdd.n2070 vdd.n762 99.5127
R16061 vdd.n2070 vdd.n763 99.5127
R16062 vdd.n763 vdd.n744 99.5127
R16063 vdd.n2588 vdd.n2587 99.5127
R16064 vdd.n2585 vdd.n2551 99.5127
R16065 vdd.n2581 vdd.n2580 99.5127
R16066 vdd.n2578 vdd.n2554 99.5127
R16067 vdd.n2574 vdd.n2573 99.5127
R16068 vdd.n2571 vdd.n2557 99.5127
R16069 vdd.n2567 vdd.n2566 99.5127
R16070 vdd.n2564 vdd.n2561 99.5127
R16071 vdd.n2705 vdd.n577 99.5127
R16072 vdd.n2703 vdd.n2702 99.5127
R16073 vdd.n2700 vdd.n579 99.5127
R16074 vdd.n2696 vdd.n2695 99.5127
R16075 vdd.n2693 vdd.n582 99.5127
R16076 vdd.n2689 vdd.n2688 99.5127
R16077 vdd.n2686 vdd.n585 99.5127
R16078 vdd.n2682 vdd.n2681 99.5127
R16079 vdd.n2679 vdd.n588 99.5127
R16080 vdd.n2323 vdd.n705 99.5127
R16081 vdd.n2323 vdd.n700 99.5127
R16082 vdd.n2394 vdd.n700 99.5127
R16083 vdd.n2394 vdd.n695 99.5127
R16084 vdd.n2390 vdd.n695 99.5127
R16085 vdd.n2390 vdd.n689 99.5127
R16086 vdd.n2387 vdd.n689 99.5127
R16087 vdd.n2387 vdd.n682 99.5127
R16088 vdd.n2384 vdd.n682 99.5127
R16089 vdd.n2384 vdd.n677 99.5127
R16090 vdd.n2381 vdd.n677 99.5127
R16091 vdd.n2381 vdd.n672 99.5127
R16092 vdd.n2378 vdd.n672 99.5127
R16093 vdd.n2378 vdd.n666 99.5127
R16094 vdd.n2375 vdd.n666 99.5127
R16095 vdd.n2375 vdd.n659 99.5127
R16096 vdd.n2340 vdd.n659 99.5127
R16097 vdd.n2340 vdd.n654 99.5127
R16098 vdd.n2337 vdd.n654 99.5127
R16099 vdd.n2337 vdd.n649 99.5127
R16100 vdd.n2334 vdd.n649 99.5127
R16101 vdd.n2334 vdd.n643 99.5127
R16102 vdd.n2331 vdd.n643 99.5127
R16103 vdd.n2331 vdd.n635 99.5127
R16104 vdd.n2328 vdd.n635 99.5127
R16105 vdd.n2328 vdd.n628 99.5127
R16106 vdd.n628 vdd.n594 99.5127
R16107 vdd.n2674 vdd.n594 99.5127
R16108 vdd.n2473 vdd.n708 99.5127
R16109 vdd.n2261 vdd.n2260 99.5127
R16110 vdd.n2265 vdd.n2264 99.5127
R16111 vdd.n2269 vdd.n2268 99.5127
R16112 vdd.n2273 vdd.n2272 99.5127
R16113 vdd.n2277 vdd.n2276 99.5127
R16114 vdd.n2281 vdd.n2280 99.5127
R16115 vdd.n2285 vdd.n2284 99.5127
R16116 vdd.n2289 vdd.n2288 99.5127
R16117 vdd.n2293 vdd.n2292 99.5127
R16118 vdd.n2297 vdd.n2296 99.5127
R16119 vdd.n2301 vdd.n2300 99.5127
R16120 vdd.n2305 vdd.n2304 99.5127
R16121 vdd.n2309 vdd.n2308 99.5127
R16122 vdd.n2313 vdd.n2312 99.5127
R16123 vdd.n2317 vdd.n2316 99.5127
R16124 vdd.n2319 vdd.n2251 99.5127
R16125 vdd.n2477 vdd.n698 99.5127
R16126 vdd.n2485 vdd.n698 99.5127
R16127 vdd.n2485 vdd.n696 99.5127
R16128 vdd.n2489 vdd.n696 99.5127
R16129 vdd.n2489 vdd.n686 99.5127
R16130 vdd.n2497 vdd.n686 99.5127
R16131 vdd.n2497 vdd.n684 99.5127
R16132 vdd.n2501 vdd.n684 99.5127
R16133 vdd.n2501 vdd.n675 99.5127
R16134 vdd.n2509 vdd.n675 99.5127
R16135 vdd.n2509 vdd.n673 99.5127
R16136 vdd.n2513 vdd.n673 99.5127
R16137 vdd.n2513 vdd.n663 99.5127
R16138 vdd.n2521 vdd.n663 99.5127
R16139 vdd.n2521 vdd.n661 99.5127
R16140 vdd.n2525 vdd.n661 99.5127
R16141 vdd.n2525 vdd.n652 99.5127
R16142 vdd.n2533 vdd.n652 99.5127
R16143 vdd.n2533 vdd.n650 99.5127
R16144 vdd.n2539 vdd.n650 99.5127
R16145 vdd.n2539 vdd.n640 99.5127
R16146 vdd.n2547 vdd.n640 99.5127
R16147 vdd.n2547 vdd.n637 99.5127
R16148 vdd.n2596 vdd.n637 99.5127
R16149 vdd.n2596 vdd.n638 99.5127
R16150 vdd.n638 vdd.n629 99.5127
R16151 vdd.n2591 vdd.n629 99.5127
R16152 vdd.n2591 vdd.n597 99.5127
R16153 vdd.n2141 vdd.n2140 99.5127
R16154 vdd.n2137 vdd.n2136 99.5127
R16155 vdd.n2133 vdd.n2132 99.5127
R16156 vdd.n2129 vdd.n2128 99.5127
R16157 vdd.n2125 vdd.n2124 99.5127
R16158 vdd.n2121 vdd.n2120 99.5127
R16159 vdd.n2117 vdd.n2116 99.5127
R16160 vdd.n2113 vdd.n2112 99.5127
R16161 vdd.n2109 vdd.n2108 99.5127
R16162 vdd.n2105 vdd.n2104 99.5127
R16163 vdd.n2101 vdd.n2100 99.5127
R16164 vdd.n2097 vdd.n2096 99.5127
R16165 vdd.n2093 vdd.n2092 99.5127
R16166 vdd.n2089 vdd.n2088 99.5127
R16167 vdd.n2085 vdd.n2084 99.5127
R16168 vdd.n2081 vdd.n2080 99.5127
R16169 vdd.n2077 vdd.n726 99.5127
R16170 vdd.n1834 vdd.n841 99.5127
R16171 vdd.n1834 vdd.n835 99.5127
R16172 vdd.n1837 vdd.n835 99.5127
R16173 vdd.n1837 vdd.n829 99.5127
R16174 vdd.n1840 vdd.n829 99.5127
R16175 vdd.n1840 vdd.n822 99.5127
R16176 vdd.n1843 vdd.n822 99.5127
R16177 vdd.n1843 vdd.n815 99.5127
R16178 vdd.n1846 vdd.n815 99.5127
R16179 vdd.n1846 vdd.n810 99.5127
R16180 vdd.n1849 vdd.n810 99.5127
R16181 vdd.n1849 vdd.n804 99.5127
R16182 vdd.n1870 vdd.n804 99.5127
R16183 vdd.n1870 vdd.n797 99.5127
R16184 vdd.n1866 vdd.n797 99.5127
R16185 vdd.n1866 vdd.n791 99.5127
R16186 vdd.n1863 vdd.n791 99.5127
R16187 vdd.n1863 vdd.n786 99.5127
R16188 vdd.n1860 vdd.n786 99.5127
R16189 vdd.n1860 vdd.n781 99.5127
R16190 vdd.n1857 vdd.n781 99.5127
R16191 vdd.n1857 vdd.n775 99.5127
R16192 vdd.n1854 vdd.n775 99.5127
R16193 vdd.n1854 vdd.n768 99.5127
R16194 vdd.n768 vdd.n759 99.5127
R16195 vdd.n2072 vdd.n759 99.5127
R16196 vdd.n2073 vdd.n2072 99.5127
R16197 vdd.n2073 vdd.n751 99.5127
R16198 vdd.n1984 vdd.n1982 99.5127
R16199 vdd.n1980 vdd.n844 99.5127
R16200 vdd.n1976 vdd.n1974 99.5127
R16201 vdd.n1972 vdd.n846 99.5127
R16202 vdd.n1968 vdd.n1966 99.5127
R16203 vdd.n1964 vdd.n848 99.5127
R16204 vdd.n1960 vdd.n1958 99.5127
R16205 vdd.n1956 vdd.n850 99.5127
R16206 vdd.n1798 vdd.n852 99.5127
R16207 vdd.n1803 vdd.n1800 99.5127
R16208 vdd.n1807 vdd.n1805 99.5127
R16209 vdd.n1811 vdd.n1796 99.5127
R16210 vdd.n1815 vdd.n1813 99.5127
R16211 vdd.n1819 vdd.n1794 99.5127
R16212 vdd.n1823 vdd.n1821 99.5127
R16213 vdd.n1828 vdd.n1790 99.5127
R16214 vdd.n1831 vdd.n1830 99.5127
R16215 vdd.n1988 vdd.n832 99.5127
R16216 vdd.n1996 vdd.n832 99.5127
R16217 vdd.n1996 vdd.n830 99.5127
R16218 vdd.n2000 vdd.n830 99.5127
R16219 vdd.n2000 vdd.n819 99.5127
R16220 vdd.n2008 vdd.n819 99.5127
R16221 vdd.n2008 vdd.n816 99.5127
R16222 vdd.n2013 vdd.n816 99.5127
R16223 vdd.n2013 vdd.n807 99.5127
R16224 vdd.n2021 vdd.n807 99.5127
R16225 vdd.n2021 vdd.n805 99.5127
R16226 vdd.n2025 vdd.n805 99.5127
R16227 vdd.n2025 vdd.n795 99.5127
R16228 vdd.n2033 vdd.n795 99.5127
R16229 vdd.n2033 vdd.n793 99.5127
R16230 vdd.n2037 vdd.n793 99.5127
R16231 vdd.n2037 vdd.n784 99.5127
R16232 vdd.n2045 vdd.n784 99.5127
R16233 vdd.n2045 vdd.n782 99.5127
R16234 vdd.n2049 vdd.n782 99.5127
R16235 vdd.n2049 vdd.n772 99.5127
R16236 vdd.n2057 vdd.n772 99.5127
R16237 vdd.n2057 vdd.n769 99.5127
R16238 vdd.n2063 vdd.n769 99.5127
R16239 vdd.n2063 vdd.n770 99.5127
R16240 vdd.n770 vdd.n761 99.5127
R16241 vdd.n761 vdd.n752 99.5127
R16242 vdd.n2145 vdd.n752 99.5127
R16243 vdd.n9 vdd.n7 98.9633
R16244 vdd.n2 vdd.n0 98.9633
R16245 vdd.n9 vdd.n8 98.6055
R16246 vdd.n11 vdd.n10 98.6055
R16247 vdd.n13 vdd.n12 98.6055
R16248 vdd.n6 vdd.n5 98.6055
R16249 vdd.n4 vdd.n3 98.6055
R16250 vdd.n2 vdd.n1 98.6055
R16251 vdd.t121 vdd.n267 85.8723
R16252 vdd.t132 vdd.n220 85.8723
R16253 vdd.t117 vdd.n177 85.8723
R16254 vdd.t127 vdd.n130 85.8723
R16255 vdd.t158 vdd.n88 85.8723
R16256 vdd.t100 vdd.n41 85.8723
R16257 vdd.t156 vdd.n1082 85.8723
R16258 vdd.t142 vdd.n1129 85.8723
R16259 vdd.t148 vdd.n992 85.8723
R16260 vdd.t135 vdd.n1039 85.8723
R16261 vdd.t98 vdd.n903 85.8723
R16262 vdd.t157 vdd.n950 85.8723
R16263 vdd.n2537 vdd.n2536 78.546
R16264 vdd.n2011 vdd.n817 78.546
R16265 vdd.n254 vdd.n253 75.1835
R16266 vdd.n252 vdd.n251 75.1835
R16267 vdd.n250 vdd.n249 75.1835
R16268 vdd.n164 vdd.n163 75.1835
R16269 vdd.n162 vdd.n161 75.1835
R16270 vdd.n160 vdd.n159 75.1835
R16271 vdd.n75 vdd.n74 75.1835
R16272 vdd.n73 vdd.n72 75.1835
R16273 vdd.n71 vdd.n70 75.1835
R16274 vdd.n1112 vdd.n1111 75.1835
R16275 vdd.n1114 vdd.n1113 75.1835
R16276 vdd.n1116 vdd.n1115 75.1835
R16277 vdd.n1022 vdd.n1021 75.1835
R16278 vdd.n1024 vdd.n1023 75.1835
R16279 vdd.n1026 vdd.n1025 75.1835
R16280 vdd.n933 vdd.n932 75.1835
R16281 vdd.n935 vdd.n934 75.1835
R16282 vdd.n937 vdd.n936 75.1835
R16283 vdd.n2472 vdd.n2471 72.8958
R16284 vdd.n2471 vdd.n2235 72.8958
R16285 vdd.n2471 vdd.n2236 72.8958
R16286 vdd.n2471 vdd.n2237 72.8958
R16287 vdd.n2471 vdd.n2238 72.8958
R16288 vdd.n2471 vdd.n2239 72.8958
R16289 vdd.n2471 vdd.n2240 72.8958
R16290 vdd.n2471 vdd.n2241 72.8958
R16291 vdd.n2471 vdd.n2242 72.8958
R16292 vdd.n2471 vdd.n2243 72.8958
R16293 vdd.n2471 vdd.n2244 72.8958
R16294 vdd.n2471 vdd.n2245 72.8958
R16295 vdd.n2471 vdd.n2246 72.8958
R16296 vdd.n2471 vdd.n2247 72.8958
R16297 vdd.n2471 vdd.n2248 72.8958
R16298 vdd.n2471 vdd.n2249 72.8958
R16299 vdd.n2471 vdd.n2250 72.8958
R16300 vdd.n593 vdd.n484 72.8958
R16301 vdd.n2680 vdd.n484 72.8958
R16302 vdd.n587 vdd.n484 72.8958
R16303 vdd.n2687 vdd.n484 72.8958
R16304 vdd.n584 vdd.n484 72.8958
R16305 vdd.n2694 vdd.n484 72.8958
R16306 vdd.n581 vdd.n484 72.8958
R16307 vdd.n2701 vdd.n484 72.8958
R16308 vdd.n2704 vdd.n484 72.8958
R16309 vdd.n2560 vdd.n484 72.8958
R16310 vdd.n2565 vdd.n484 72.8958
R16311 vdd.n2559 vdd.n484 72.8958
R16312 vdd.n2572 vdd.n484 72.8958
R16313 vdd.n2556 vdd.n484 72.8958
R16314 vdd.n2579 vdd.n484 72.8958
R16315 vdd.n2553 vdd.n484 72.8958
R16316 vdd.n2586 vdd.n484 72.8958
R16317 vdd.n1724 vdd.n839 72.8958
R16318 vdd.n1730 vdd.n839 72.8958
R16319 vdd.n1732 vdd.n839 72.8958
R16320 vdd.n1738 vdd.n839 72.8958
R16321 vdd.n1740 vdd.n839 72.8958
R16322 vdd.n1746 vdd.n839 72.8958
R16323 vdd.n1748 vdd.n839 72.8958
R16324 vdd.n1754 vdd.n839 72.8958
R16325 vdd.n1925 vdd.n839 72.8958
R16326 vdd.n1923 vdd.n839 72.8958
R16327 vdd.n1917 vdd.n839 72.8958
R16328 vdd.n1915 vdd.n839 72.8958
R16329 vdd.n1909 vdd.n839 72.8958
R16330 vdd.n1907 vdd.n839 72.8958
R16331 vdd.n1901 vdd.n839 72.8958
R16332 vdd.n1899 vdd.n839 72.8958
R16333 vdd.n1893 vdd.n839 72.8958
R16334 vdd.n2218 vdd.n727 72.8958
R16335 vdd.n2218 vdd.n728 72.8958
R16336 vdd.n2218 vdd.n729 72.8958
R16337 vdd.n2218 vdd.n730 72.8958
R16338 vdd.n2218 vdd.n731 72.8958
R16339 vdd.n2218 vdd.n732 72.8958
R16340 vdd.n2218 vdd.n733 72.8958
R16341 vdd.n2218 vdd.n734 72.8958
R16342 vdd.n2218 vdd.n735 72.8958
R16343 vdd.n2218 vdd.n736 72.8958
R16344 vdd.n2218 vdd.n737 72.8958
R16345 vdd.n2218 vdd.n738 72.8958
R16346 vdd.n2218 vdd.n739 72.8958
R16347 vdd.n2218 vdd.n740 72.8958
R16348 vdd.n2218 vdd.n741 72.8958
R16349 vdd.n2218 vdd.n742 72.8958
R16350 vdd.n2218 vdd.n743 72.8958
R16351 vdd.n2471 vdd.n2470 72.8958
R16352 vdd.n2471 vdd.n2219 72.8958
R16353 vdd.n2471 vdd.n2220 72.8958
R16354 vdd.n2471 vdd.n2221 72.8958
R16355 vdd.n2471 vdd.n2222 72.8958
R16356 vdd.n2471 vdd.n2223 72.8958
R16357 vdd.n2471 vdd.n2224 72.8958
R16358 vdd.n2471 vdd.n2225 72.8958
R16359 vdd.n2471 vdd.n2226 72.8958
R16360 vdd.n2471 vdd.n2227 72.8958
R16361 vdd.n2471 vdd.n2228 72.8958
R16362 vdd.n2471 vdd.n2229 72.8958
R16363 vdd.n2471 vdd.n2230 72.8958
R16364 vdd.n2471 vdd.n2231 72.8958
R16365 vdd.n2471 vdd.n2232 72.8958
R16366 vdd.n2471 vdd.n2233 72.8958
R16367 vdd.n2471 vdd.n2234 72.8958
R16368 vdd.n2610 vdd.n484 72.8958
R16369 vdd.n625 vdd.n484 72.8958
R16370 vdd.n2618 vdd.n484 72.8958
R16371 vdd.n620 vdd.n484 72.8958
R16372 vdd.n2625 vdd.n484 72.8958
R16373 vdd.n617 vdd.n484 72.8958
R16374 vdd.n2632 vdd.n484 72.8958
R16375 vdd.n614 vdd.n484 72.8958
R16376 vdd.n2639 vdd.n484 72.8958
R16377 vdd.n2643 vdd.n484 72.8958
R16378 vdd.n611 vdd.n484 72.8958
R16379 vdd.n2650 vdd.n484 72.8958
R16380 vdd.n608 vdd.n484 72.8958
R16381 vdd.n2657 vdd.n484 72.8958
R16382 vdd.n605 vdd.n484 72.8958
R16383 vdd.n2664 vdd.n484 72.8958
R16384 vdd.n2667 vdd.n484 72.8958
R16385 vdd.n2218 vdd.n725 72.8958
R16386 vdd.n2218 vdd.n724 72.8958
R16387 vdd.n2218 vdd.n723 72.8958
R16388 vdd.n2218 vdd.n722 72.8958
R16389 vdd.n2218 vdd.n721 72.8958
R16390 vdd.n2218 vdd.n720 72.8958
R16391 vdd.n2218 vdd.n719 72.8958
R16392 vdd.n2218 vdd.n718 72.8958
R16393 vdd.n2218 vdd.n717 72.8958
R16394 vdd.n2218 vdd.n716 72.8958
R16395 vdd.n2218 vdd.n715 72.8958
R16396 vdd.n2218 vdd.n714 72.8958
R16397 vdd.n2218 vdd.n713 72.8958
R16398 vdd.n2218 vdd.n712 72.8958
R16399 vdd.n2218 vdd.n711 72.8958
R16400 vdd.n2218 vdd.n710 72.8958
R16401 vdd.n2218 vdd.n709 72.8958
R16402 vdd.n1983 vdd.n839 72.8958
R16403 vdd.n1981 vdd.n839 72.8958
R16404 vdd.n1975 vdd.n839 72.8958
R16405 vdd.n1973 vdd.n839 72.8958
R16406 vdd.n1967 vdd.n839 72.8958
R16407 vdd.n1965 vdd.n839 72.8958
R16408 vdd.n1959 vdd.n839 72.8958
R16409 vdd.n1957 vdd.n839 72.8958
R16410 vdd.n851 vdd.n839 72.8958
R16411 vdd.n1799 vdd.n839 72.8958
R16412 vdd.n1804 vdd.n839 72.8958
R16413 vdd.n1806 vdd.n839 72.8958
R16414 vdd.n1812 vdd.n839 72.8958
R16415 vdd.n1814 vdd.n839 72.8958
R16416 vdd.n1820 vdd.n839 72.8958
R16417 vdd.n1822 vdd.n839 72.8958
R16418 vdd.n1829 vdd.n839 72.8958
R16419 vdd.n1422 vdd.n1421 66.2847
R16420 vdd.n1421 vdd.n1197 66.2847
R16421 vdd.n1421 vdd.n1198 66.2847
R16422 vdd.n1421 vdd.n1199 66.2847
R16423 vdd.n1421 vdd.n1200 66.2847
R16424 vdd.n1421 vdd.n1201 66.2847
R16425 vdd.n1421 vdd.n1202 66.2847
R16426 vdd.n1421 vdd.n1203 66.2847
R16427 vdd.n1421 vdd.n1204 66.2847
R16428 vdd.n1421 vdd.n1205 66.2847
R16429 vdd.n1421 vdd.n1206 66.2847
R16430 vdd.n1421 vdd.n1207 66.2847
R16431 vdd.n1421 vdd.n1208 66.2847
R16432 vdd.n1421 vdd.n1209 66.2847
R16433 vdd.n1421 vdd.n1210 66.2847
R16434 vdd.n1421 vdd.n1211 66.2847
R16435 vdd.n1421 vdd.n1212 66.2847
R16436 vdd.n1421 vdd.n1213 66.2847
R16437 vdd.n1421 vdd.n1214 66.2847
R16438 vdd.n1421 vdd.n1215 66.2847
R16439 vdd.n1421 vdd.n1216 66.2847
R16440 vdd.n1421 vdd.n1217 66.2847
R16441 vdd.n1421 vdd.n1218 66.2847
R16442 vdd.n1421 vdd.n1219 66.2847
R16443 vdd.n1421 vdd.n1220 66.2847
R16444 vdd.n1421 vdd.n1221 66.2847
R16445 vdd.n1421 vdd.n1222 66.2847
R16446 vdd.n1421 vdd.n1223 66.2847
R16447 vdd.n1421 vdd.n1224 66.2847
R16448 vdd.n1421 vdd.n1225 66.2847
R16449 vdd.n1421 vdd.n1226 66.2847
R16450 vdd.n863 vdd.n860 66.2847
R16451 vdd.n1614 vdd.n863 66.2847
R16452 vdd.n1619 vdd.n863 66.2847
R16453 vdd.n1624 vdd.n863 66.2847
R16454 vdd.n1612 vdd.n863 66.2847
R16455 vdd.n1631 vdd.n863 66.2847
R16456 vdd.n1604 vdd.n863 66.2847
R16457 vdd.n1638 vdd.n863 66.2847
R16458 vdd.n1597 vdd.n863 66.2847
R16459 vdd.n1645 vdd.n863 66.2847
R16460 vdd.n1591 vdd.n863 66.2847
R16461 vdd.n1586 vdd.n863 66.2847
R16462 vdd.n1656 vdd.n863 66.2847
R16463 vdd.n1578 vdd.n863 66.2847
R16464 vdd.n1663 vdd.n863 66.2847
R16465 vdd.n1571 vdd.n863 66.2847
R16466 vdd.n1670 vdd.n863 66.2847
R16467 vdd.n1564 vdd.n863 66.2847
R16468 vdd.n1677 vdd.n863 66.2847
R16469 vdd.n1557 vdd.n863 66.2847
R16470 vdd.n1684 vdd.n863 66.2847
R16471 vdd.n1551 vdd.n863 66.2847
R16472 vdd.n1546 vdd.n863 66.2847
R16473 vdd.n1695 vdd.n863 66.2847
R16474 vdd.n1538 vdd.n863 66.2847
R16475 vdd.n1702 vdd.n863 66.2847
R16476 vdd.n1531 vdd.n863 66.2847
R16477 vdd.n1709 vdd.n863 66.2847
R16478 vdd.n1712 vdd.n863 66.2847
R16479 vdd.n1522 vdd.n863 66.2847
R16480 vdd.n1934 vdd.n863 66.2847
R16481 vdd.n1516 vdd.n863 66.2847
R16482 vdd.n2841 vdd.n2840 66.2847
R16483 vdd.n2840 vdd.n485 66.2847
R16484 vdd.n2840 vdd.n486 66.2847
R16485 vdd.n2840 vdd.n487 66.2847
R16486 vdd.n2840 vdd.n488 66.2847
R16487 vdd.n2840 vdd.n489 66.2847
R16488 vdd.n2840 vdd.n490 66.2847
R16489 vdd.n2840 vdd.n491 66.2847
R16490 vdd.n2840 vdd.n492 66.2847
R16491 vdd.n2840 vdd.n493 66.2847
R16492 vdd.n2840 vdd.n494 66.2847
R16493 vdd.n2840 vdd.n495 66.2847
R16494 vdd.n2840 vdd.n496 66.2847
R16495 vdd.n2840 vdd.n497 66.2847
R16496 vdd.n2840 vdd.n498 66.2847
R16497 vdd.n2840 vdd.n499 66.2847
R16498 vdd.n2840 vdd.n500 66.2847
R16499 vdd.n2840 vdd.n501 66.2847
R16500 vdd.n2840 vdd.n502 66.2847
R16501 vdd.n2840 vdd.n503 66.2847
R16502 vdd.n2840 vdd.n504 66.2847
R16503 vdd.n2840 vdd.n505 66.2847
R16504 vdd.n2840 vdd.n506 66.2847
R16505 vdd.n2840 vdd.n507 66.2847
R16506 vdd.n2840 vdd.n508 66.2847
R16507 vdd.n2840 vdd.n509 66.2847
R16508 vdd.n2840 vdd.n510 66.2847
R16509 vdd.n2840 vdd.n511 66.2847
R16510 vdd.n2840 vdd.n512 66.2847
R16511 vdd.n2840 vdd.n513 66.2847
R16512 vdd.n2840 vdd.n514 66.2847
R16513 vdd.n2905 vdd.n329 66.2847
R16514 vdd.n2914 vdd.n329 66.2847
R16515 vdd.n439 vdd.n329 66.2847
R16516 vdd.n2921 vdd.n329 66.2847
R16517 vdd.n432 vdd.n329 66.2847
R16518 vdd.n2928 vdd.n329 66.2847
R16519 vdd.n425 vdd.n329 66.2847
R16520 vdd.n2935 vdd.n329 66.2847
R16521 vdd.n418 vdd.n329 66.2847
R16522 vdd.n2942 vdd.n329 66.2847
R16523 vdd.n412 vdd.n329 66.2847
R16524 vdd.n407 vdd.n329 66.2847
R16525 vdd.n2953 vdd.n329 66.2847
R16526 vdd.n399 vdd.n329 66.2847
R16527 vdd.n2960 vdd.n329 66.2847
R16528 vdd.n392 vdd.n329 66.2847
R16529 vdd.n2967 vdd.n329 66.2847
R16530 vdd.n385 vdd.n329 66.2847
R16531 vdd.n2974 vdd.n329 66.2847
R16532 vdd.n378 vdd.n329 66.2847
R16533 vdd.n2981 vdd.n329 66.2847
R16534 vdd.n372 vdd.n329 66.2847
R16535 vdd.n367 vdd.n329 66.2847
R16536 vdd.n2992 vdd.n329 66.2847
R16537 vdd.n359 vdd.n329 66.2847
R16538 vdd.n2999 vdd.n329 66.2847
R16539 vdd.n352 vdd.n329 66.2847
R16540 vdd.n3006 vdd.n329 66.2847
R16541 vdd.n345 vdd.n329 66.2847
R16542 vdd.n3013 vdd.n329 66.2847
R16543 vdd.n3016 vdd.n329 66.2847
R16544 vdd.n333 vdd.n329 66.2847
R16545 vdd.n334 vdd.n333 52.4337
R16546 vdd.n3016 vdd.n3015 52.4337
R16547 vdd.n3013 vdd.n3012 52.4337
R16548 vdd.n3008 vdd.n345 52.4337
R16549 vdd.n3006 vdd.n3005 52.4337
R16550 vdd.n3001 vdd.n352 52.4337
R16551 vdd.n2999 vdd.n2998 52.4337
R16552 vdd.n2994 vdd.n359 52.4337
R16553 vdd.n2992 vdd.n2991 52.4337
R16554 vdd.n368 vdd.n367 52.4337
R16555 vdd.n2983 vdd.n372 52.4337
R16556 vdd.n2981 vdd.n2980 52.4337
R16557 vdd.n2976 vdd.n378 52.4337
R16558 vdd.n2974 vdd.n2973 52.4337
R16559 vdd.n2969 vdd.n385 52.4337
R16560 vdd.n2967 vdd.n2966 52.4337
R16561 vdd.n2962 vdd.n392 52.4337
R16562 vdd.n2960 vdd.n2959 52.4337
R16563 vdd.n2955 vdd.n399 52.4337
R16564 vdd.n2953 vdd.n2952 52.4337
R16565 vdd.n408 vdd.n407 52.4337
R16566 vdd.n2944 vdd.n412 52.4337
R16567 vdd.n2942 vdd.n2941 52.4337
R16568 vdd.n2937 vdd.n418 52.4337
R16569 vdd.n2935 vdd.n2934 52.4337
R16570 vdd.n2930 vdd.n425 52.4337
R16571 vdd.n2928 vdd.n2927 52.4337
R16572 vdd.n2923 vdd.n432 52.4337
R16573 vdd.n2921 vdd.n2920 52.4337
R16574 vdd.n2916 vdd.n439 52.4337
R16575 vdd.n2914 vdd.n2913 52.4337
R16576 vdd.n2906 vdd.n2905 52.4337
R16577 vdd.n2842 vdd.n2841 52.4337
R16578 vdd.n517 vdd.n485 52.4337
R16579 vdd.n523 vdd.n486 52.4337
R16580 vdd.n2831 vdd.n487 52.4337
R16581 vdd.n2827 vdd.n488 52.4337
R16582 vdd.n2823 vdd.n489 52.4337
R16583 vdd.n2819 vdd.n490 52.4337
R16584 vdd.n2815 vdd.n491 52.4337
R16585 vdd.n2811 vdd.n492 52.4337
R16586 vdd.n2807 vdd.n493 52.4337
R16587 vdd.n2799 vdd.n494 52.4337
R16588 vdd.n2795 vdd.n495 52.4337
R16589 vdd.n2791 vdd.n496 52.4337
R16590 vdd.n2787 vdd.n497 52.4337
R16591 vdd.n2783 vdd.n498 52.4337
R16592 vdd.n2779 vdd.n499 52.4337
R16593 vdd.n2775 vdd.n500 52.4337
R16594 vdd.n2771 vdd.n501 52.4337
R16595 vdd.n2767 vdd.n502 52.4337
R16596 vdd.n2763 vdd.n503 52.4337
R16597 vdd.n2759 vdd.n504 52.4337
R16598 vdd.n2753 vdd.n505 52.4337
R16599 vdd.n2749 vdd.n506 52.4337
R16600 vdd.n2745 vdd.n507 52.4337
R16601 vdd.n2741 vdd.n508 52.4337
R16602 vdd.n2737 vdd.n509 52.4337
R16603 vdd.n2733 vdd.n510 52.4337
R16604 vdd.n2729 vdd.n511 52.4337
R16605 vdd.n2725 vdd.n512 52.4337
R16606 vdd.n2721 vdd.n513 52.4337
R16607 vdd.n2717 vdd.n514 52.4337
R16608 vdd.n1936 vdd.n1516 52.4337
R16609 vdd.n1934 vdd.n1933 52.4337
R16610 vdd.n1523 vdd.n1522 52.4337
R16611 vdd.n1712 vdd.n1711 52.4337
R16612 vdd.n1709 vdd.n1708 52.4337
R16613 vdd.n1704 vdd.n1531 52.4337
R16614 vdd.n1702 vdd.n1701 52.4337
R16615 vdd.n1697 vdd.n1538 52.4337
R16616 vdd.n1695 vdd.n1694 52.4337
R16617 vdd.n1547 vdd.n1546 52.4337
R16618 vdd.n1686 vdd.n1551 52.4337
R16619 vdd.n1684 vdd.n1683 52.4337
R16620 vdd.n1679 vdd.n1557 52.4337
R16621 vdd.n1677 vdd.n1676 52.4337
R16622 vdd.n1672 vdd.n1564 52.4337
R16623 vdd.n1670 vdd.n1669 52.4337
R16624 vdd.n1665 vdd.n1571 52.4337
R16625 vdd.n1663 vdd.n1662 52.4337
R16626 vdd.n1658 vdd.n1578 52.4337
R16627 vdd.n1656 vdd.n1655 52.4337
R16628 vdd.n1587 vdd.n1586 52.4337
R16629 vdd.n1647 vdd.n1591 52.4337
R16630 vdd.n1645 vdd.n1644 52.4337
R16631 vdd.n1640 vdd.n1597 52.4337
R16632 vdd.n1638 vdd.n1637 52.4337
R16633 vdd.n1633 vdd.n1604 52.4337
R16634 vdd.n1631 vdd.n1630 52.4337
R16635 vdd.n1626 vdd.n1612 52.4337
R16636 vdd.n1624 vdd.n1623 52.4337
R16637 vdd.n1619 vdd.n1618 52.4337
R16638 vdd.n1614 vdd.n1613 52.4337
R16639 vdd.n1945 vdd.n860 52.4337
R16640 vdd.n1423 vdd.n1422 52.4337
R16641 vdd.n1229 vdd.n1197 52.4337
R16642 vdd.n1233 vdd.n1198 52.4337
R16643 vdd.n1235 vdd.n1199 52.4337
R16644 vdd.n1239 vdd.n1200 52.4337
R16645 vdd.n1241 vdd.n1201 52.4337
R16646 vdd.n1245 vdd.n1202 52.4337
R16647 vdd.n1247 vdd.n1203 52.4337
R16648 vdd.n1251 vdd.n1204 52.4337
R16649 vdd.n1253 vdd.n1205 52.4337
R16650 vdd.n1259 vdd.n1206 52.4337
R16651 vdd.n1261 vdd.n1207 52.4337
R16652 vdd.n1265 vdd.n1208 52.4337
R16653 vdd.n1267 vdd.n1209 52.4337
R16654 vdd.n1271 vdd.n1210 52.4337
R16655 vdd.n1273 vdd.n1211 52.4337
R16656 vdd.n1277 vdd.n1212 52.4337
R16657 vdd.n1279 vdd.n1213 52.4337
R16658 vdd.n1283 vdd.n1214 52.4337
R16659 vdd.n1285 vdd.n1215 52.4337
R16660 vdd.n1357 vdd.n1216 52.4337
R16661 vdd.n1290 vdd.n1217 52.4337
R16662 vdd.n1294 vdd.n1218 52.4337
R16663 vdd.n1296 vdd.n1219 52.4337
R16664 vdd.n1300 vdd.n1220 52.4337
R16665 vdd.n1302 vdd.n1221 52.4337
R16666 vdd.n1306 vdd.n1222 52.4337
R16667 vdd.n1308 vdd.n1223 52.4337
R16668 vdd.n1312 vdd.n1224 52.4337
R16669 vdd.n1314 vdd.n1225 52.4337
R16670 vdd.n1318 vdd.n1226 52.4337
R16671 vdd.n1422 vdd.n1196 52.4337
R16672 vdd.n1232 vdd.n1197 52.4337
R16673 vdd.n1234 vdd.n1198 52.4337
R16674 vdd.n1238 vdd.n1199 52.4337
R16675 vdd.n1240 vdd.n1200 52.4337
R16676 vdd.n1244 vdd.n1201 52.4337
R16677 vdd.n1246 vdd.n1202 52.4337
R16678 vdd.n1250 vdd.n1203 52.4337
R16679 vdd.n1252 vdd.n1204 52.4337
R16680 vdd.n1258 vdd.n1205 52.4337
R16681 vdd.n1260 vdd.n1206 52.4337
R16682 vdd.n1264 vdd.n1207 52.4337
R16683 vdd.n1266 vdd.n1208 52.4337
R16684 vdd.n1270 vdd.n1209 52.4337
R16685 vdd.n1272 vdd.n1210 52.4337
R16686 vdd.n1276 vdd.n1211 52.4337
R16687 vdd.n1278 vdd.n1212 52.4337
R16688 vdd.n1282 vdd.n1213 52.4337
R16689 vdd.n1284 vdd.n1214 52.4337
R16690 vdd.n1288 vdd.n1215 52.4337
R16691 vdd.n1289 vdd.n1216 52.4337
R16692 vdd.n1293 vdd.n1217 52.4337
R16693 vdd.n1295 vdd.n1218 52.4337
R16694 vdd.n1299 vdd.n1219 52.4337
R16695 vdd.n1301 vdd.n1220 52.4337
R16696 vdd.n1305 vdd.n1221 52.4337
R16697 vdd.n1307 vdd.n1222 52.4337
R16698 vdd.n1311 vdd.n1223 52.4337
R16699 vdd.n1313 vdd.n1224 52.4337
R16700 vdd.n1317 vdd.n1225 52.4337
R16701 vdd.n1319 vdd.n1226 52.4337
R16702 vdd.n860 vdd.n859 52.4337
R16703 vdd.n1615 vdd.n1614 52.4337
R16704 vdd.n1620 vdd.n1619 52.4337
R16705 vdd.n1625 vdd.n1624 52.4337
R16706 vdd.n1612 vdd.n1605 52.4337
R16707 vdd.n1632 vdd.n1631 52.4337
R16708 vdd.n1604 vdd.n1598 52.4337
R16709 vdd.n1639 vdd.n1638 52.4337
R16710 vdd.n1597 vdd.n1592 52.4337
R16711 vdd.n1646 vdd.n1645 52.4337
R16712 vdd.n1591 vdd.n1590 52.4337
R16713 vdd.n1586 vdd.n1579 52.4337
R16714 vdd.n1657 vdd.n1656 52.4337
R16715 vdd.n1578 vdd.n1572 52.4337
R16716 vdd.n1664 vdd.n1663 52.4337
R16717 vdd.n1571 vdd.n1565 52.4337
R16718 vdd.n1671 vdd.n1670 52.4337
R16719 vdd.n1564 vdd.n1558 52.4337
R16720 vdd.n1678 vdd.n1677 52.4337
R16721 vdd.n1557 vdd.n1552 52.4337
R16722 vdd.n1685 vdd.n1684 52.4337
R16723 vdd.n1551 vdd.n1550 52.4337
R16724 vdd.n1546 vdd.n1539 52.4337
R16725 vdd.n1696 vdd.n1695 52.4337
R16726 vdd.n1538 vdd.n1532 52.4337
R16727 vdd.n1703 vdd.n1702 52.4337
R16728 vdd.n1531 vdd.n1525 52.4337
R16729 vdd.n1710 vdd.n1709 52.4337
R16730 vdd.n1713 vdd.n1712 52.4337
R16731 vdd.n1522 vdd.n1517 52.4337
R16732 vdd.n1935 vdd.n1934 52.4337
R16733 vdd.n1516 vdd.n865 52.4337
R16734 vdd.n2841 vdd.n483 52.4337
R16735 vdd.n522 vdd.n485 52.4337
R16736 vdd.n2832 vdd.n486 52.4337
R16737 vdd.n2828 vdd.n487 52.4337
R16738 vdd.n2824 vdd.n488 52.4337
R16739 vdd.n2820 vdd.n489 52.4337
R16740 vdd.n2816 vdd.n490 52.4337
R16741 vdd.n2812 vdd.n491 52.4337
R16742 vdd.n2808 vdd.n492 52.4337
R16743 vdd.n2798 vdd.n493 52.4337
R16744 vdd.n2796 vdd.n494 52.4337
R16745 vdd.n2792 vdd.n495 52.4337
R16746 vdd.n2788 vdd.n496 52.4337
R16747 vdd.n2784 vdd.n497 52.4337
R16748 vdd.n2780 vdd.n498 52.4337
R16749 vdd.n2776 vdd.n499 52.4337
R16750 vdd.n2772 vdd.n500 52.4337
R16751 vdd.n2768 vdd.n501 52.4337
R16752 vdd.n2764 vdd.n502 52.4337
R16753 vdd.n2760 vdd.n503 52.4337
R16754 vdd.n2752 vdd.n504 52.4337
R16755 vdd.n2750 vdd.n505 52.4337
R16756 vdd.n2746 vdd.n506 52.4337
R16757 vdd.n2742 vdd.n507 52.4337
R16758 vdd.n2738 vdd.n508 52.4337
R16759 vdd.n2734 vdd.n509 52.4337
R16760 vdd.n2730 vdd.n510 52.4337
R16761 vdd.n2726 vdd.n511 52.4337
R16762 vdd.n2722 vdd.n512 52.4337
R16763 vdd.n2718 vdd.n513 52.4337
R16764 vdd.n2714 vdd.n514 52.4337
R16765 vdd.n2905 vdd.n440 52.4337
R16766 vdd.n2915 vdd.n2914 52.4337
R16767 vdd.n439 vdd.n433 52.4337
R16768 vdd.n2922 vdd.n2921 52.4337
R16769 vdd.n432 vdd.n426 52.4337
R16770 vdd.n2929 vdd.n2928 52.4337
R16771 vdd.n425 vdd.n419 52.4337
R16772 vdd.n2936 vdd.n2935 52.4337
R16773 vdd.n418 vdd.n413 52.4337
R16774 vdd.n2943 vdd.n2942 52.4337
R16775 vdd.n412 vdd.n411 52.4337
R16776 vdd.n407 vdd.n400 52.4337
R16777 vdd.n2954 vdd.n2953 52.4337
R16778 vdd.n399 vdd.n393 52.4337
R16779 vdd.n2961 vdd.n2960 52.4337
R16780 vdd.n392 vdd.n386 52.4337
R16781 vdd.n2968 vdd.n2967 52.4337
R16782 vdd.n385 vdd.n379 52.4337
R16783 vdd.n2975 vdd.n2974 52.4337
R16784 vdd.n378 vdd.n373 52.4337
R16785 vdd.n2982 vdd.n2981 52.4337
R16786 vdd.n372 vdd.n371 52.4337
R16787 vdd.n367 vdd.n360 52.4337
R16788 vdd.n2993 vdd.n2992 52.4337
R16789 vdd.n359 vdd.n353 52.4337
R16790 vdd.n3000 vdd.n2999 52.4337
R16791 vdd.n352 vdd.n346 52.4337
R16792 vdd.n3007 vdd.n3006 52.4337
R16793 vdd.n345 vdd.n338 52.4337
R16794 vdd.n3014 vdd.n3013 52.4337
R16795 vdd.n3017 vdd.n3016 52.4337
R16796 vdd.n333 vdd.n330 52.4337
R16797 vdd.t5 vdd.t12 51.4683
R16798 vdd.n250 vdd.n248 42.0461
R16799 vdd.n160 vdd.n158 42.0461
R16800 vdd.n71 vdd.n69 42.0461
R16801 vdd.n1112 vdd.n1110 42.0461
R16802 vdd.n1022 vdd.n1020 42.0461
R16803 vdd.n933 vdd.n931 42.0461
R16804 vdd.n296 vdd.n295 41.6884
R16805 vdd.n206 vdd.n205 41.6884
R16806 vdd.n117 vdd.n116 41.6884
R16807 vdd.n1158 vdd.n1157 41.6884
R16808 vdd.n1068 vdd.n1067 41.6884
R16809 vdd.n979 vdd.n978 41.6884
R16810 vdd.n1322 vdd.n1321 41.1157
R16811 vdd.n1360 vdd.n1359 41.1157
R16812 vdd.n1256 vdd.n1255 41.1157
R16813 vdd.n2910 vdd.n2909 41.1157
R16814 vdd.n2949 vdd.n406 41.1157
R16815 vdd.n2988 vdd.n366 41.1157
R16816 vdd.n2667 vdd.n2666 39.2114
R16817 vdd.n2664 vdd.n2663 39.2114
R16818 vdd.n2659 vdd.n605 39.2114
R16819 vdd.n2657 vdd.n2656 39.2114
R16820 vdd.n2652 vdd.n608 39.2114
R16821 vdd.n2650 vdd.n2649 39.2114
R16822 vdd.n2645 vdd.n611 39.2114
R16823 vdd.n2643 vdd.n2642 39.2114
R16824 vdd.n2639 vdd.n2638 39.2114
R16825 vdd.n2634 vdd.n614 39.2114
R16826 vdd.n2632 vdd.n2631 39.2114
R16827 vdd.n2627 vdd.n617 39.2114
R16828 vdd.n2625 vdd.n2624 39.2114
R16829 vdd.n2620 vdd.n620 39.2114
R16830 vdd.n2618 vdd.n2617 39.2114
R16831 vdd.n2612 vdd.n625 39.2114
R16832 vdd.n2610 vdd.n2609 39.2114
R16833 vdd.n2470 vdd.n703 39.2114
R16834 vdd.n2465 vdd.n2219 39.2114
R16835 vdd.n2462 vdd.n2220 39.2114
R16836 vdd.n2458 vdd.n2221 39.2114
R16837 vdd.n2454 vdd.n2222 39.2114
R16838 vdd.n2450 vdd.n2223 39.2114
R16839 vdd.n2446 vdd.n2224 39.2114
R16840 vdd.n2442 vdd.n2225 39.2114
R16841 vdd.n2438 vdd.n2226 39.2114
R16842 vdd.n2434 vdd.n2227 39.2114
R16843 vdd.n2430 vdd.n2228 39.2114
R16844 vdd.n2426 vdd.n2229 39.2114
R16845 vdd.n2422 vdd.n2230 39.2114
R16846 vdd.n2418 vdd.n2231 39.2114
R16847 vdd.n2414 vdd.n2232 39.2114
R16848 vdd.n2410 vdd.n2233 39.2114
R16849 vdd.n2405 vdd.n2234 39.2114
R16850 vdd.n2213 vdd.n743 39.2114
R16851 vdd.n2209 vdd.n742 39.2114
R16852 vdd.n2205 vdd.n741 39.2114
R16853 vdd.n2201 vdd.n740 39.2114
R16854 vdd.n2197 vdd.n739 39.2114
R16855 vdd.n2193 vdd.n738 39.2114
R16856 vdd.n2189 vdd.n737 39.2114
R16857 vdd.n2185 vdd.n736 39.2114
R16858 vdd.n2181 vdd.n735 39.2114
R16859 vdd.n2177 vdd.n734 39.2114
R16860 vdd.n2173 vdd.n733 39.2114
R16861 vdd.n2169 vdd.n732 39.2114
R16862 vdd.n2165 vdd.n731 39.2114
R16863 vdd.n2161 vdd.n730 39.2114
R16864 vdd.n2157 vdd.n729 39.2114
R16865 vdd.n2152 vdd.n728 39.2114
R16866 vdd.n2148 vdd.n727 39.2114
R16867 vdd.n1724 vdd.n838 39.2114
R16868 vdd.n1730 vdd.n1729 39.2114
R16869 vdd.n1733 vdd.n1732 39.2114
R16870 vdd.n1738 vdd.n1737 39.2114
R16871 vdd.n1741 vdd.n1740 39.2114
R16872 vdd.n1746 vdd.n1745 39.2114
R16873 vdd.n1749 vdd.n1748 39.2114
R16874 vdd.n1754 vdd.n1753 39.2114
R16875 vdd.n1925 vdd.n1756 39.2114
R16876 vdd.n1924 vdd.n1923 39.2114
R16877 vdd.n1917 vdd.n1758 39.2114
R16878 vdd.n1916 vdd.n1915 39.2114
R16879 vdd.n1909 vdd.n1760 39.2114
R16880 vdd.n1908 vdd.n1907 39.2114
R16881 vdd.n1901 vdd.n1762 39.2114
R16882 vdd.n1900 vdd.n1899 39.2114
R16883 vdd.n1893 vdd.n1764 39.2114
R16884 vdd.n2586 vdd.n2585 39.2114
R16885 vdd.n2581 vdd.n2553 39.2114
R16886 vdd.n2579 vdd.n2578 39.2114
R16887 vdd.n2574 vdd.n2556 39.2114
R16888 vdd.n2572 vdd.n2571 39.2114
R16889 vdd.n2567 vdd.n2559 39.2114
R16890 vdd.n2565 vdd.n2564 39.2114
R16891 vdd.n2560 vdd.n577 39.2114
R16892 vdd.n2704 vdd.n2703 39.2114
R16893 vdd.n2701 vdd.n2700 39.2114
R16894 vdd.n2696 vdd.n581 39.2114
R16895 vdd.n2694 vdd.n2693 39.2114
R16896 vdd.n2689 vdd.n584 39.2114
R16897 vdd.n2687 vdd.n2686 39.2114
R16898 vdd.n2682 vdd.n587 39.2114
R16899 vdd.n2680 vdd.n2679 39.2114
R16900 vdd.n2675 vdd.n593 39.2114
R16901 vdd.n2472 vdd.n706 39.2114
R16902 vdd.n2235 vdd.n708 39.2114
R16903 vdd.n2261 vdd.n2236 39.2114
R16904 vdd.n2265 vdd.n2237 39.2114
R16905 vdd.n2269 vdd.n2238 39.2114
R16906 vdd.n2273 vdd.n2239 39.2114
R16907 vdd.n2277 vdd.n2240 39.2114
R16908 vdd.n2281 vdd.n2241 39.2114
R16909 vdd.n2285 vdd.n2242 39.2114
R16910 vdd.n2289 vdd.n2243 39.2114
R16911 vdd.n2293 vdd.n2244 39.2114
R16912 vdd.n2297 vdd.n2245 39.2114
R16913 vdd.n2301 vdd.n2246 39.2114
R16914 vdd.n2305 vdd.n2247 39.2114
R16915 vdd.n2309 vdd.n2248 39.2114
R16916 vdd.n2313 vdd.n2249 39.2114
R16917 vdd.n2317 vdd.n2250 39.2114
R16918 vdd.n2473 vdd.n2472 39.2114
R16919 vdd.n2260 vdd.n2235 39.2114
R16920 vdd.n2264 vdd.n2236 39.2114
R16921 vdd.n2268 vdd.n2237 39.2114
R16922 vdd.n2272 vdd.n2238 39.2114
R16923 vdd.n2276 vdd.n2239 39.2114
R16924 vdd.n2280 vdd.n2240 39.2114
R16925 vdd.n2284 vdd.n2241 39.2114
R16926 vdd.n2288 vdd.n2242 39.2114
R16927 vdd.n2292 vdd.n2243 39.2114
R16928 vdd.n2296 vdd.n2244 39.2114
R16929 vdd.n2300 vdd.n2245 39.2114
R16930 vdd.n2304 vdd.n2246 39.2114
R16931 vdd.n2308 vdd.n2247 39.2114
R16932 vdd.n2312 vdd.n2248 39.2114
R16933 vdd.n2316 vdd.n2249 39.2114
R16934 vdd.n2319 vdd.n2250 39.2114
R16935 vdd.n593 vdd.n588 39.2114
R16936 vdd.n2681 vdd.n2680 39.2114
R16937 vdd.n587 vdd.n585 39.2114
R16938 vdd.n2688 vdd.n2687 39.2114
R16939 vdd.n584 vdd.n582 39.2114
R16940 vdd.n2695 vdd.n2694 39.2114
R16941 vdd.n581 vdd.n579 39.2114
R16942 vdd.n2702 vdd.n2701 39.2114
R16943 vdd.n2705 vdd.n2704 39.2114
R16944 vdd.n2561 vdd.n2560 39.2114
R16945 vdd.n2566 vdd.n2565 39.2114
R16946 vdd.n2559 vdd.n2557 39.2114
R16947 vdd.n2573 vdd.n2572 39.2114
R16948 vdd.n2556 vdd.n2554 39.2114
R16949 vdd.n2580 vdd.n2579 39.2114
R16950 vdd.n2553 vdd.n2551 39.2114
R16951 vdd.n2587 vdd.n2586 39.2114
R16952 vdd.n1725 vdd.n1724 39.2114
R16953 vdd.n1731 vdd.n1730 39.2114
R16954 vdd.n1732 vdd.n1721 39.2114
R16955 vdd.n1739 vdd.n1738 39.2114
R16956 vdd.n1740 vdd.n1719 39.2114
R16957 vdd.n1747 vdd.n1746 39.2114
R16958 vdd.n1748 vdd.n1717 39.2114
R16959 vdd.n1755 vdd.n1754 39.2114
R16960 vdd.n1926 vdd.n1925 39.2114
R16961 vdd.n1923 vdd.n1922 39.2114
R16962 vdd.n1918 vdd.n1917 39.2114
R16963 vdd.n1915 vdd.n1914 39.2114
R16964 vdd.n1910 vdd.n1909 39.2114
R16965 vdd.n1907 vdd.n1906 39.2114
R16966 vdd.n1902 vdd.n1901 39.2114
R16967 vdd.n1899 vdd.n1898 39.2114
R16968 vdd.n1894 vdd.n1893 39.2114
R16969 vdd.n2151 vdd.n727 39.2114
R16970 vdd.n2156 vdd.n728 39.2114
R16971 vdd.n2160 vdd.n729 39.2114
R16972 vdd.n2164 vdd.n730 39.2114
R16973 vdd.n2168 vdd.n731 39.2114
R16974 vdd.n2172 vdd.n732 39.2114
R16975 vdd.n2176 vdd.n733 39.2114
R16976 vdd.n2180 vdd.n734 39.2114
R16977 vdd.n2184 vdd.n735 39.2114
R16978 vdd.n2188 vdd.n736 39.2114
R16979 vdd.n2192 vdd.n737 39.2114
R16980 vdd.n2196 vdd.n738 39.2114
R16981 vdd.n2200 vdd.n739 39.2114
R16982 vdd.n2204 vdd.n740 39.2114
R16983 vdd.n2208 vdd.n741 39.2114
R16984 vdd.n2212 vdd.n742 39.2114
R16985 vdd.n745 vdd.n743 39.2114
R16986 vdd.n2470 vdd.n2469 39.2114
R16987 vdd.n2463 vdd.n2219 39.2114
R16988 vdd.n2459 vdd.n2220 39.2114
R16989 vdd.n2455 vdd.n2221 39.2114
R16990 vdd.n2451 vdd.n2222 39.2114
R16991 vdd.n2447 vdd.n2223 39.2114
R16992 vdd.n2443 vdd.n2224 39.2114
R16993 vdd.n2439 vdd.n2225 39.2114
R16994 vdd.n2435 vdd.n2226 39.2114
R16995 vdd.n2431 vdd.n2227 39.2114
R16996 vdd.n2427 vdd.n2228 39.2114
R16997 vdd.n2423 vdd.n2229 39.2114
R16998 vdd.n2419 vdd.n2230 39.2114
R16999 vdd.n2415 vdd.n2231 39.2114
R17000 vdd.n2411 vdd.n2232 39.2114
R17001 vdd.n2406 vdd.n2233 39.2114
R17002 vdd.n2402 vdd.n2234 39.2114
R17003 vdd.n2611 vdd.n2610 39.2114
R17004 vdd.n625 vdd.n621 39.2114
R17005 vdd.n2619 vdd.n2618 39.2114
R17006 vdd.n620 vdd.n618 39.2114
R17007 vdd.n2626 vdd.n2625 39.2114
R17008 vdd.n617 vdd.n615 39.2114
R17009 vdd.n2633 vdd.n2632 39.2114
R17010 vdd.n614 vdd.n612 39.2114
R17011 vdd.n2640 vdd.n2639 39.2114
R17012 vdd.n2644 vdd.n2643 39.2114
R17013 vdd.n611 vdd.n609 39.2114
R17014 vdd.n2651 vdd.n2650 39.2114
R17015 vdd.n608 vdd.n606 39.2114
R17016 vdd.n2658 vdd.n2657 39.2114
R17017 vdd.n605 vdd.n603 39.2114
R17018 vdd.n2665 vdd.n2664 39.2114
R17019 vdd.n2668 vdd.n2667 39.2114
R17020 vdd.n753 vdd.n709 39.2114
R17021 vdd.n2140 vdd.n710 39.2114
R17022 vdd.n2136 vdd.n711 39.2114
R17023 vdd.n2132 vdd.n712 39.2114
R17024 vdd.n2128 vdd.n713 39.2114
R17025 vdd.n2124 vdd.n714 39.2114
R17026 vdd.n2120 vdd.n715 39.2114
R17027 vdd.n2116 vdd.n716 39.2114
R17028 vdd.n2112 vdd.n717 39.2114
R17029 vdd.n2108 vdd.n718 39.2114
R17030 vdd.n2104 vdd.n719 39.2114
R17031 vdd.n2100 vdd.n720 39.2114
R17032 vdd.n2096 vdd.n721 39.2114
R17033 vdd.n2092 vdd.n722 39.2114
R17034 vdd.n2088 vdd.n723 39.2114
R17035 vdd.n2084 vdd.n724 39.2114
R17036 vdd.n2080 vdd.n725 39.2114
R17037 vdd.n1983 vdd.n842 39.2114
R17038 vdd.n1982 vdd.n1981 39.2114
R17039 vdd.n1975 vdd.n844 39.2114
R17040 vdd.n1974 vdd.n1973 39.2114
R17041 vdd.n1967 vdd.n846 39.2114
R17042 vdd.n1966 vdd.n1965 39.2114
R17043 vdd.n1959 vdd.n848 39.2114
R17044 vdd.n1958 vdd.n1957 39.2114
R17045 vdd.n851 vdd.n850 39.2114
R17046 vdd.n1799 vdd.n1798 39.2114
R17047 vdd.n1804 vdd.n1803 39.2114
R17048 vdd.n1807 vdd.n1806 39.2114
R17049 vdd.n1812 vdd.n1811 39.2114
R17050 vdd.n1815 vdd.n1814 39.2114
R17051 vdd.n1820 vdd.n1819 39.2114
R17052 vdd.n1823 vdd.n1822 39.2114
R17053 vdd.n1829 vdd.n1828 39.2114
R17054 vdd.n2077 vdd.n725 39.2114
R17055 vdd.n2081 vdd.n724 39.2114
R17056 vdd.n2085 vdd.n723 39.2114
R17057 vdd.n2089 vdd.n722 39.2114
R17058 vdd.n2093 vdd.n721 39.2114
R17059 vdd.n2097 vdd.n720 39.2114
R17060 vdd.n2101 vdd.n719 39.2114
R17061 vdd.n2105 vdd.n718 39.2114
R17062 vdd.n2109 vdd.n717 39.2114
R17063 vdd.n2113 vdd.n716 39.2114
R17064 vdd.n2117 vdd.n715 39.2114
R17065 vdd.n2121 vdd.n714 39.2114
R17066 vdd.n2125 vdd.n713 39.2114
R17067 vdd.n2129 vdd.n712 39.2114
R17068 vdd.n2133 vdd.n711 39.2114
R17069 vdd.n2137 vdd.n710 39.2114
R17070 vdd.n2141 vdd.n709 39.2114
R17071 vdd.n1984 vdd.n1983 39.2114
R17072 vdd.n1981 vdd.n1980 39.2114
R17073 vdd.n1976 vdd.n1975 39.2114
R17074 vdd.n1973 vdd.n1972 39.2114
R17075 vdd.n1968 vdd.n1967 39.2114
R17076 vdd.n1965 vdd.n1964 39.2114
R17077 vdd.n1960 vdd.n1959 39.2114
R17078 vdd.n1957 vdd.n1956 39.2114
R17079 vdd.n852 vdd.n851 39.2114
R17080 vdd.n1800 vdd.n1799 39.2114
R17081 vdd.n1805 vdd.n1804 39.2114
R17082 vdd.n1806 vdd.n1796 39.2114
R17083 vdd.n1813 vdd.n1812 39.2114
R17084 vdd.n1814 vdd.n1794 39.2114
R17085 vdd.n1821 vdd.n1820 39.2114
R17086 vdd.n1822 vdd.n1790 39.2114
R17087 vdd.n1830 vdd.n1829 39.2114
R17088 vdd.n1949 vdd.n1948 37.2369
R17089 vdd.n1652 vdd.n1585 37.2369
R17090 vdd.n1691 vdd.n1545 37.2369
R17091 vdd.n2758 vdd.n558 37.2369
R17092 vdd.n2806 vdd.n2805 37.2369
R17093 vdd.n2713 vdd.n2712 37.2369
R17094 vdd.n1991 vdd.n837 31.6883
R17095 vdd.n2216 vdd.n746 31.6883
R17096 vdd.n2149 vdd.n749 31.6883
R17097 vdd.n1895 vdd.n1892 31.6883
R17098 vdd.n2403 vdd.n2401 31.6883
R17099 vdd.n2608 vdd.n2607 31.6883
R17100 vdd.n2480 vdd.n702 31.6883
R17101 vdd.n2671 vdd.n2670 31.6883
R17102 vdd.n2590 vdd.n2589 31.6883
R17103 vdd.n2676 vdd.n592 31.6883
R17104 vdd.n2322 vdd.n2321 31.6883
R17105 vdd.n2476 vdd.n2475 31.6883
R17106 vdd.n1987 vdd.n1986 31.6883
R17107 vdd.n2144 vdd.n2143 31.6883
R17108 vdd.n2076 vdd.n2075 31.6883
R17109 vdd.n1833 vdd.n1832 31.6883
R17110 vdd.n1826 vdd.n1792 30.449
R17111 vdd.n757 vdd.n756 30.449
R17112 vdd.n1767 vdd.n1766 30.449
R17113 vdd.n2154 vdd.n748 30.449
R17114 vdd.n2258 vdd.n2257 30.449
R17115 vdd.n2614 vdd.n623 30.449
R17116 vdd.n2408 vdd.n2254 30.449
R17117 vdd.n591 vdd.n590 30.449
R17118 vdd.n1421 vdd.n1228 22.6735
R17119 vdd.n1943 vdd.n863 22.6735
R17120 vdd.n2840 vdd.n516 22.6735
R17121 vdd.n3025 vdd.n329 22.6735
R17122 vdd.n1432 vdd.n1190 19.3944
R17123 vdd.n1432 vdd.n1188 19.3944
R17124 vdd.n1436 vdd.n1188 19.3944
R17125 vdd.n1436 vdd.n1178 19.3944
R17126 vdd.n1449 vdd.n1178 19.3944
R17127 vdd.n1449 vdd.n1176 19.3944
R17128 vdd.n1453 vdd.n1176 19.3944
R17129 vdd.n1453 vdd.n1168 19.3944
R17130 vdd.n1467 vdd.n1168 19.3944
R17131 vdd.n1467 vdd.n1166 19.3944
R17132 vdd.n1471 vdd.n1166 19.3944
R17133 vdd.n1471 vdd.n885 19.3944
R17134 vdd.n1483 vdd.n885 19.3944
R17135 vdd.n1483 vdd.n883 19.3944
R17136 vdd.n1487 vdd.n883 19.3944
R17137 vdd.n1487 vdd.n875 19.3944
R17138 vdd.n1500 vdd.n875 19.3944
R17139 vdd.n1500 vdd.n872 19.3944
R17140 vdd.n1506 vdd.n872 19.3944
R17141 vdd.n1506 vdd.n873 19.3944
R17142 vdd.n873 vdd.n862 19.3944
R17143 vdd.n1356 vdd.n1291 19.3944
R17144 vdd.n1352 vdd.n1291 19.3944
R17145 vdd.n1352 vdd.n1351 19.3944
R17146 vdd.n1351 vdd.n1350 19.3944
R17147 vdd.n1350 vdd.n1297 19.3944
R17148 vdd.n1346 vdd.n1297 19.3944
R17149 vdd.n1346 vdd.n1345 19.3944
R17150 vdd.n1345 vdd.n1344 19.3944
R17151 vdd.n1344 vdd.n1303 19.3944
R17152 vdd.n1340 vdd.n1303 19.3944
R17153 vdd.n1340 vdd.n1339 19.3944
R17154 vdd.n1339 vdd.n1338 19.3944
R17155 vdd.n1338 vdd.n1309 19.3944
R17156 vdd.n1334 vdd.n1309 19.3944
R17157 vdd.n1334 vdd.n1333 19.3944
R17158 vdd.n1333 vdd.n1332 19.3944
R17159 vdd.n1332 vdd.n1315 19.3944
R17160 vdd.n1328 vdd.n1315 19.3944
R17161 vdd.n1328 vdd.n1327 19.3944
R17162 vdd.n1327 vdd.n1326 19.3944
R17163 vdd.n1391 vdd.n1390 19.3944
R17164 vdd.n1390 vdd.n1389 19.3944
R17165 vdd.n1389 vdd.n1262 19.3944
R17166 vdd.n1385 vdd.n1262 19.3944
R17167 vdd.n1385 vdd.n1384 19.3944
R17168 vdd.n1384 vdd.n1383 19.3944
R17169 vdd.n1383 vdd.n1268 19.3944
R17170 vdd.n1379 vdd.n1268 19.3944
R17171 vdd.n1379 vdd.n1378 19.3944
R17172 vdd.n1378 vdd.n1377 19.3944
R17173 vdd.n1377 vdd.n1274 19.3944
R17174 vdd.n1373 vdd.n1274 19.3944
R17175 vdd.n1373 vdd.n1372 19.3944
R17176 vdd.n1372 vdd.n1371 19.3944
R17177 vdd.n1371 vdd.n1280 19.3944
R17178 vdd.n1367 vdd.n1280 19.3944
R17179 vdd.n1367 vdd.n1366 19.3944
R17180 vdd.n1366 vdd.n1365 19.3944
R17181 vdd.n1365 vdd.n1286 19.3944
R17182 vdd.n1361 vdd.n1286 19.3944
R17183 vdd.n1424 vdd.n1195 19.3944
R17184 vdd.n1419 vdd.n1195 19.3944
R17185 vdd.n1419 vdd.n1230 19.3944
R17186 vdd.n1415 vdd.n1230 19.3944
R17187 vdd.n1415 vdd.n1414 19.3944
R17188 vdd.n1414 vdd.n1413 19.3944
R17189 vdd.n1413 vdd.n1236 19.3944
R17190 vdd.n1409 vdd.n1236 19.3944
R17191 vdd.n1409 vdd.n1408 19.3944
R17192 vdd.n1408 vdd.n1407 19.3944
R17193 vdd.n1407 vdd.n1242 19.3944
R17194 vdd.n1403 vdd.n1242 19.3944
R17195 vdd.n1403 vdd.n1402 19.3944
R17196 vdd.n1402 vdd.n1401 19.3944
R17197 vdd.n1401 vdd.n1248 19.3944
R17198 vdd.n1397 vdd.n1248 19.3944
R17199 vdd.n1397 vdd.n1396 19.3944
R17200 vdd.n1396 vdd.n1395 19.3944
R17201 vdd.n1648 vdd.n1583 19.3944
R17202 vdd.n1648 vdd.n1589 19.3944
R17203 vdd.n1643 vdd.n1589 19.3944
R17204 vdd.n1643 vdd.n1642 19.3944
R17205 vdd.n1642 vdd.n1641 19.3944
R17206 vdd.n1641 vdd.n1596 19.3944
R17207 vdd.n1636 vdd.n1596 19.3944
R17208 vdd.n1636 vdd.n1635 19.3944
R17209 vdd.n1635 vdd.n1634 19.3944
R17210 vdd.n1634 vdd.n1603 19.3944
R17211 vdd.n1629 vdd.n1603 19.3944
R17212 vdd.n1629 vdd.n1628 19.3944
R17213 vdd.n1628 vdd.n1627 19.3944
R17214 vdd.n1627 vdd.n1611 19.3944
R17215 vdd.n1622 vdd.n1611 19.3944
R17216 vdd.n1622 vdd.n1621 19.3944
R17217 vdd.n1617 vdd.n1616 19.3944
R17218 vdd.n1950 vdd.n858 19.3944
R17219 vdd.n1687 vdd.n1543 19.3944
R17220 vdd.n1687 vdd.n1549 19.3944
R17221 vdd.n1682 vdd.n1549 19.3944
R17222 vdd.n1682 vdd.n1681 19.3944
R17223 vdd.n1681 vdd.n1680 19.3944
R17224 vdd.n1680 vdd.n1556 19.3944
R17225 vdd.n1675 vdd.n1556 19.3944
R17226 vdd.n1675 vdd.n1674 19.3944
R17227 vdd.n1674 vdd.n1673 19.3944
R17228 vdd.n1673 vdd.n1563 19.3944
R17229 vdd.n1668 vdd.n1563 19.3944
R17230 vdd.n1668 vdd.n1667 19.3944
R17231 vdd.n1667 vdd.n1666 19.3944
R17232 vdd.n1666 vdd.n1570 19.3944
R17233 vdd.n1661 vdd.n1570 19.3944
R17234 vdd.n1661 vdd.n1660 19.3944
R17235 vdd.n1660 vdd.n1659 19.3944
R17236 vdd.n1659 vdd.n1577 19.3944
R17237 vdd.n1654 vdd.n1577 19.3944
R17238 vdd.n1654 vdd.n1653 19.3944
R17239 vdd.n1938 vdd.n1937 19.3944
R17240 vdd.n1937 vdd.n1515 19.3944
R17241 vdd.n1932 vdd.n1931 19.3944
R17242 vdd.n1714 vdd.n1519 19.3944
R17243 vdd.n1714 vdd.n1521 19.3944
R17244 vdd.n1524 vdd.n1521 19.3944
R17245 vdd.n1707 vdd.n1524 19.3944
R17246 vdd.n1707 vdd.n1706 19.3944
R17247 vdd.n1706 vdd.n1705 19.3944
R17248 vdd.n1705 vdd.n1530 19.3944
R17249 vdd.n1700 vdd.n1530 19.3944
R17250 vdd.n1700 vdd.n1699 19.3944
R17251 vdd.n1699 vdd.n1698 19.3944
R17252 vdd.n1698 vdd.n1537 19.3944
R17253 vdd.n1693 vdd.n1537 19.3944
R17254 vdd.n1693 vdd.n1692 19.3944
R17255 vdd.n1428 vdd.n1193 19.3944
R17256 vdd.n1428 vdd.n1184 19.3944
R17257 vdd.n1441 vdd.n1184 19.3944
R17258 vdd.n1441 vdd.n1182 19.3944
R17259 vdd.n1445 vdd.n1182 19.3944
R17260 vdd.n1445 vdd.n1173 19.3944
R17261 vdd.n1458 vdd.n1173 19.3944
R17262 vdd.n1458 vdd.n1171 19.3944
R17263 vdd.n1463 vdd.n1171 19.3944
R17264 vdd.n1463 vdd.n1162 19.3944
R17265 vdd.n1475 vdd.n1162 19.3944
R17266 vdd.n1475 vdd.n890 19.3944
R17267 vdd.n1479 vdd.n890 19.3944
R17268 vdd.n1479 vdd.n880 19.3944
R17269 vdd.n1492 vdd.n880 19.3944
R17270 vdd.n1492 vdd.n878 19.3944
R17271 vdd.n1496 vdd.n878 19.3944
R17272 vdd.n1496 vdd.n868 19.3944
R17273 vdd.n1511 vdd.n868 19.3944
R17274 vdd.n1511 vdd.n866 19.3944
R17275 vdd.n1941 vdd.n866 19.3944
R17276 vdd.n2851 vdd.n477 19.3944
R17277 vdd.n2851 vdd.n475 19.3944
R17278 vdd.n2855 vdd.n475 19.3944
R17279 vdd.n2855 vdd.n465 19.3944
R17280 vdd.n2868 vdd.n465 19.3944
R17281 vdd.n2868 vdd.n463 19.3944
R17282 vdd.n2872 vdd.n463 19.3944
R17283 vdd.n2872 vdd.n453 19.3944
R17284 vdd.n2884 vdd.n453 19.3944
R17285 vdd.n2884 vdd.n451 19.3944
R17286 vdd.n2888 vdd.n451 19.3944
R17287 vdd.n2889 vdd.n2888 19.3944
R17288 vdd.n2890 vdd.n2889 19.3944
R17289 vdd.n2890 vdd.n449 19.3944
R17290 vdd.n2894 vdd.n449 19.3944
R17291 vdd.n2895 vdd.n2894 19.3944
R17292 vdd.n2896 vdd.n2895 19.3944
R17293 vdd.n2896 vdd.n446 19.3944
R17294 vdd.n2900 vdd.n446 19.3944
R17295 vdd.n2901 vdd.n2900 19.3944
R17296 vdd.n2902 vdd.n2901 19.3944
R17297 vdd.n2945 vdd.n404 19.3944
R17298 vdd.n2945 vdd.n410 19.3944
R17299 vdd.n2940 vdd.n410 19.3944
R17300 vdd.n2940 vdd.n2939 19.3944
R17301 vdd.n2939 vdd.n2938 19.3944
R17302 vdd.n2938 vdd.n417 19.3944
R17303 vdd.n2933 vdd.n417 19.3944
R17304 vdd.n2933 vdd.n2932 19.3944
R17305 vdd.n2932 vdd.n2931 19.3944
R17306 vdd.n2931 vdd.n424 19.3944
R17307 vdd.n2926 vdd.n424 19.3944
R17308 vdd.n2926 vdd.n2925 19.3944
R17309 vdd.n2925 vdd.n2924 19.3944
R17310 vdd.n2924 vdd.n431 19.3944
R17311 vdd.n2919 vdd.n431 19.3944
R17312 vdd.n2919 vdd.n2918 19.3944
R17313 vdd.n2918 vdd.n2917 19.3944
R17314 vdd.n2917 vdd.n438 19.3944
R17315 vdd.n2912 vdd.n438 19.3944
R17316 vdd.n2912 vdd.n2911 19.3944
R17317 vdd.n2984 vdd.n364 19.3944
R17318 vdd.n2984 vdd.n370 19.3944
R17319 vdd.n2979 vdd.n370 19.3944
R17320 vdd.n2979 vdd.n2978 19.3944
R17321 vdd.n2978 vdd.n2977 19.3944
R17322 vdd.n2977 vdd.n377 19.3944
R17323 vdd.n2972 vdd.n377 19.3944
R17324 vdd.n2972 vdd.n2971 19.3944
R17325 vdd.n2971 vdd.n2970 19.3944
R17326 vdd.n2970 vdd.n384 19.3944
R17327 vdd.n2965 vdd.n384 19.3944
R17328 vdd.n2965 vdd.n2964 19.3944
R17329 vdd.n2964 vdd.n2963 19.3944
R17330 vdd.n2963 vdd.n391 19.3944
R17331 vdd.n2958 vdd.n391 19.3944
R17332 vdd.n2958 vdd.n2957 19.3944
R17333 vdd.n2957 vdd.n2956 19.3944
R17334 vdd.n2956 vdd.n398 19.3944
R17335 vdd.n2951 vdd.n398 19.3944
R17336 vdd.n2951 vdd.n2950 19.3944
R17337 vdd.n3020 vdd.n3019 19.3944
R17338 vdd.n3019 vdd.n3018 19.3944
R17339 vdd.n3018 vdd.n336 19.3944
R17340 vdd.n337 vdd.n336 19.3944
R17341 vdd.n3011 vdd.n337 19.3944
R17342 vdd.n3011 vdd.n3010 19.3944
R17343 vdd.n3010 vdd.n3009 19.3944
R17344 vdd.n3009 vdd.n344 19.3944
R17345 vdd.n3004 vdd.n344 19.3944
R17346 vdd.n3004 vdd.n3003 19.3944
R17347 vdd.n3003 vdd.n3002 19.3944
R17348 vdd.n3002 vdd.n351 19.3944
R17349 vdd.n2997 vdd.n351 19.3944
R17350 vdd.n2997 vdd.n2996 19.3944
R17351 vdd.n2996 vdd.n2995 19.3944
R17352 vdd.n2995 vdd.n358 19.3944
R17353 vdd.n2990 vdd.n358 19.3944
R17354 vdd.n2990 vdd.n2989 19.3944
R17355 vdd.n2847 vdd.n480 19.3944
R17356 vdd.n2847 vdd.n471 19.3944
R17357 vdd.n2860 vdd.n471 19.3944
R17358 vdd.n2860 vdd.n469 19.3944
R17359 vdd.n2864 vdd.n469 19.3944
R17360 vdd.n2864 vdd.n460 19.3944
R17361 vdd.n2876 vdd.n460 19.3944
R17362 vdd.n2876 vdd.n458 19.3944
R17363 vdd.n2880 vdd.n458 19.3944
R17364 vdd.n2880 vdd.n300 19.3944
R17365 vdd.n3045 vdd.n300 19.3944
R17366 vdd.n3045 vdd.n301 19.3944
R17367 vdd.n3039 vdd.n301 19.3944
R17368 vdd.n3039 vdd.n3038 19.3944
R17369 vdd.n3038 vdd.n3037 19.3944
R17370 vdd.n3037 vdd.n313 19.3944
R17371 vdd.n3031 vdd.n313 19.3944
R17372 vdd.n3031 vdd.n3030 19.3944
R17373 vdd.n3030 vdd.n3029 19.3944
R17374 vdd.n3029 vdd.n324 19.3944
R17375 vdd.n3023 vdd.n324 19.3944
R17376 vdd.n2800 vdd.n536 19.3944
R17377 vdd.n2800 vdd.n2797 19.3944
R17378 vdd.n2797 vdd.n2794 19.3944
R17379 vdd.n2794 vdd.n2793 19.3944
R17380 vdd.n2793 vdd.n2790 19.3944
R17381 vdd.n2790 vdd.n2789 19.3944
R17382 vdd.n2789 vdd.n2786 19.3944
R17383 vdd.n2786 vdd.n2785 19.3944
R17384 vdd.n2785 vdd.n2782 19.3944
R17385 vdd.n2782 vdd.n2781 19.3944
R17386 vdd.n2781 vdd.n2778 19.3944
R17387 vdd.n2778 vdd.n2777 19.3944
R17388 vdd.n2777 vdd.n2774 19.3944
R17389 vdd.n2774 vdd.n2773 19.3944
R17390 vdd.n2773 vdd.n2770 19.3944
R17391 vdd.n2770 vdd.n2769 19.3944
R17392 vdd.n2769 vdd.n2766 19.3944
R17393 vdd.n2766 vdd.n2765 19.3944
R17394 vdd.n2765 vdd.n2762 19.3944
R17395 vdd.n2762 vdd.n2761 19.3944
R17396 vdd.n2843 vdd.n482 19.3944
R17397 vdd.n2838 vdd.n482 19.3944
R17398 vdd.n521 vdd.n518 19.3944
R17399 vdd.n2834 vdd.n2833 19.3944
R17400 vdd.n2833 vdd.n2830 19.3944
R17401 vdd.n2830 vdd.n2829 19.3944
R17402 vdd.n2829 vdd.n2826 19.3944
R17403 vdd.n2826 vdd.n2825 19.3944
R17404 vdd.n2825 vdd.n2822 19.3944
R17405 vdd.n2822 vdd.n2821 19.3944
R17406 vdd.n2821 vdd.n2818 19.3944
R17407 vdd.n2818 vdd.n2817 19.3944
R17408 vdd.n2817 vdd.n2814 19.3944
R17409 vdd.n2814 vdd.n2813 19.3944
R17410 vdd.n2813 vdd.n2810 19.3944
R17411 vdd.n2810 vdd.n2809 19.3944
R17412 vdd.n2754 vdd.n556 19.3944
R17413 vdd.n2754 vdd.n2751 19.3944
R17414 vdd.n2751 vdd.n2748 19.3944
R17415 vdd.n2748 vdd.n2747 19.3944
R17416 vdd.n2747 vdd.n2744 19.3944
R17417 vdd.n2744 vdd.n2743 19.3944
R17418 vdd.n2743 vdd.n2740 19.3944
R17419 vdd.n2740 vdd.n2739 19.3944
R17420 vdd.n2739 vdd.n2736 19.3944
R17421 vdd.n2736 vdd.n2735 19.3944
R17422 vdd.n2735 vdd.n2732 19.3944
R17423 vdd.n2732 vdd.n2731 19.3944
R17424 vdd.n2731 vdd.n2728 19.3944
R17425 vdd.n2728 vdd.n2727 19.3944
R17426 vdd.n2727 vdd.n2724 19.3944
R17427 vdd.n2724 vdd.n2723 19.3944
R17428 vdd.n2720 vdd.n2719 19.3944
R17429 vdd.n2716 vdd.n2715 19.3944
R17430 vdd.n1360 vdd.n1356 19.0066
R17431 vdd.n1652 vdd.n1583 19.0066
R17432 vdd.n2949 vdd.n404 19.0066
R17433 vdd.n2758 vdd.n556 19.0066
R17434 vdd.n1792 vdd.n1791 16.0975
R17435 vdd.n756 vdd.n755 16.0975
R17436 vdd.n1321 vdd.n1320 16.0975
R17437 vdd.n1359 vdd.n1358 16.0975
R17438 vdd.n1255 vdd.n1254 16.0975
R17439 vdd.n1948 vdd.n1947 16.0975
R17440 vdd.n1585 vdd.n1584 16.0975
R17441 vdd.n1545 vdd.n1544 16.0975
R17442 vdd.n1766 vdd.n1765 16.0975
R17443 vdd.n748 vdd.n747 16.0975
R17444 vdd.n2257 vdd.n2256 16.0975
R17445 vdd.n2909 vdd.n2908 16.0975
R17446 vdd.n406 vdd.n405 16.0975
R17447 vdd.n366 vdd.n365 16.0975
R17448 vdd.n558 vdd.n557 16.0975
R17449 vdd.n2805 vdd.n2804 16.0975
R17450 vdd.n623 vdd.n622 16.0975
R17451 vdd.n2254 vdd.n2253 16.0975
R17452 vdd.n2712 vdd.n2711 16.0975
R17453 vdd.n590 vdd.n589 16.0975
R17454 vdd.t12 vdd.n2218 15.4182
R17455 vdd.n2471 vdd.t5 15.4182
R17456 vdd.n28 vdd.n27 14.5238
R17457 vdd.n1989 vdd.n839 14.5112
R17458 vdd.n2673 vdd.n484 14.5112
R17459 vdd.n292 vdd.n257 13.1884
R17460 vdd.n245 vdd.n210 13.1884
R17461 vdd.n202 vdd.n167 13.1884
R17462 vdd.n155 vdd.n120 13.1884
R17463 vdd.n113 vdd.n78 13.1884
R17464 vdd.n66 vdd.n31 13.1884
R17465 vdd.n1107 vdd.n1072 13.1884
R17466 vdd.n1154 vdd.n1119 13.1884
R17467 vdd.n1017 vdd.n982 13.1884
R17468 vdd.n1064 vdd.n1029 13.1884
R17469 vdd.n928 vdd.n893 13.1884
R17470 vdd.n975 vdd.n940 13.1884
R17471 vdd.n1391 vdd.n1256 12.9944
R17472 vdd.n1395 vdd.n1256 12.9944
R17473 vdd.n1691 vdd.n1543 12.9944
R17474 vdd.n1692 vdd.n1691 12.9944
R17475 vdd.n2988 vdd.n364 12.9944
R17476 vdd.n2989 vdd.n2988 12.9944
R17477 vdd.n2806 vdd.n536 12.9944
R17478 vdd.n2809 vdd.n2806 12.9944
R17479 vdd.n293 vdd.n255 12.8005
R17480 vdd.n288 vdd.n259 12.8005
R17481 vdd.n246 vdd.n208 12.8005
R17482 vdd.n241 vdd.n212 12.8005
R17483 vdd.n203 vdd.n165 12.8005
R17484 vdd.n198 vdd.n169 12.8005
R17485 vdd.n156 vdd.n118 12.8005
R17486 vdd.n151 vdd.n122 12.8005
R17487 vdd.n114 vdd.n76 12.8005
R17488 vdd.n109 vdd.n80 12.8005
R17489 vdd.n67 vdd.n29 12.8005
R17490 vdd.n62 vdd.n33 12.8005
R17491 vdd.n1108 vdd.n1070 12.8005
R17492 vdd.n1103 vdd.n1074 12.8005
R17493 vdd.n1155 vdd.n1117 12.8005
R17494 vdd.n1150 vdd.n1121 12.8005
R17495 vdd.n1018 vdd.n980 12.8005
R17496 vdd.n1013 vdd.n984 12.8005
R17497 vdd.n1065 vdd.n1027 12.8005
R17498 vdd.n1060 vdd.n1031 12.8005
R17499 vdd.n929 vdd.n891 12.8005
R17500 vdd.n924 vdd.n895 12.8005
R17501 vdd.n976 vdd.n938 12.8005
R17502 vdd.n971 vdd.n942 12.8005
R17503 vdd.n287 vdd.n260 12.0247
R17504 vdd.n240 vdd.n213 12.0247
R17505 vdd.n197 vdd.n170 12.0247
R17506 vdd.n150 vdd.n123 12.0247
R17507 vdd.n108 vdd.n81 12.0247
R17508 vdd.n61 vdd.n34 12.0247
R17509 vdd.n1102 vdd.n1075 12.0247
R17510 vdd.n1149 vdd.n1122 12.0247
R17511 vdd.n1012 vdd.n985 12.0247
R17512 vdd.n1059 vdd.n1032 12.0247
R17513 vdd.n923 vdd.n896 12.0247
R17514 vdd.n970 vdd.n943 12.0247
R17515 vdd.n1430 vdd.n1186 11.337
R17516 vdd.n1439 vdd.n1186 11.337
R17517 vdd.n1439 vdd.n1438 11.337
R17518 vdd.n1447 vdd.n1180 11.337
R17519 vdd.n1456 vdd.n1455 11.337
R17520 vdd.n1473 vdd.n1164 11.337
R17521 vdd.n1481 vdd.n887 11.337
R17522 vdd.n1490 vdd.n1489 11.337
R17523 vdd.n1498 vdd.n870 11.337
R17524 vdd.n1509 vdd.n870 11.337
R17525 vdd.n1509 vdd.n1508 11.337
R17526 vdd.n2849 vdd.n473 11.337
R17527 vdd.n2858 vdd.n473 11.337
R17528 vdd.n2858 vdd.n2857 11.337
R17529 vdd.n2866 vdd.n467 11.337
R17530 vdd.n2882 vdd.n456 11.337
R17531 vdd.n3043 vdd.n304 11.337
R17532 vdd.n3041 vdd.n308 11.337
R17533 vdd.n3035 vdd.n3034 11.337
R17534 vdd.n3033 vdd.n318 11.337
R17535 vdd.n3027 vdd.n318 11.337
R17536 vdd.n3027 vdd.n3026 11.337
R17537 vdd.n284 vdd.n283 11.249
R17538 vdd.n237 vdd.n236 11.249
R17539 vdd.n194 vdd.n193 11.249
R17540 vdd.n147 vdd.n146 11.249
R17541 vdd.n105 vdd.n104 11.249
R17542 vdd.n58 vdd.n57 11.249
R17543 vdd.n1099 vdd.n1098 11.249
R17544 vdd.n1146 vdd.n1145 11.249
R17545 vdd.n1009 vdd.n1008 11.249
R17546 vdd.n1056 vdd.n1055 11.249
R17547 vdd.n920 vdd.n919 11.249
R17548 vdd.n967 vdd.n966 11.249
R17549 vdd.n2146 vdd.t15 11.1103
R17550 vdd.n2478 vdd.t198 11.1103
R17551 vdd.n1228 vdd.t33 10.7702
R17552 vdd.t44 vdd.n3025 10.7702
R17553 vdd.n269 vdd.n268 10.7238
R17554 vdd.n222 vdd.n221 10.7238
R17555 vdd.n179 vdd.n178 10.7238
R17556 vdd.n132 vdd.n131 10.7238
R17557 vdd.n90 vdd.n89 10.7238
R17558 vdd.n43 vdd.n42 10.7238
R17559 vdd.n1084 vdd.n1083 10.7238
R17560 vdd.n1131 vdd.n1130 10.7238
R17561 vdd.n994 vdd.n993 10.7238
R17562 vdd.n1041 vdd.n1040 10.7238
R17563 vdd.n905 vdd.n904 10.7238
R17564 vdd.n952 vdd.n951 10.7238
R17565 vdd.n1992 vdd.n1991 10.6151
R17566 vdd.n1993 vdd.n1992 10.6151
R17567 vdd.n1993 vdd.n825 10.6151
R17568 vdd.n2003 vdd.n825 10.6151
R17569 vdd.n2004 vdd.n2003 10.6151
R17570 vdd.n2005 vdd.n2004 10.6151
R17571 vdd.n2005 vdd.n812 10.6151
R17572 vdd.n2016 vdd.n812 10.6151
R17573 vdd.n2017 vdd.n2016 10.6151
R17574 vdd.n2018 vdd.n2017 10.6151
R17575 vdd.n2018 vdd.n800 10.6151
R17576 vdd.n2028 vdd.n800 10.6151
R17577 vdd.n2029 vdd.n2028 10.6151
R17578 vdd.n2030 vdd.n2029 10.6151
R17579 vdd.n2030 vdd.n788 10.6151
R17580 vdd.n2040 vdd.n788 10.6151
R17581 vdd.n2041 vdd.n2040 10.6151
R17582 vdd.n2042 vdd.n2041 10.6151
R17583 vdd.n2042 vdd.n777 10.6151
R17584 vdd.n2052 vdd.n777 10.6151
R17585 vdd.n2053 vdd.n2052 10.6151
R17586 vdd.n2054 vdd.n2053 10.6151
R17587 vdd.n2054 vdd.n764 10.6151
R17588 vdd.n2066 vdd.n764 10.6151
R17589 vdd.n2067 vdd.n2066 10.6151
R17590 vdd.n2069 vdd.n2067 10.6151
R17591 vdd.n2069 vdd.n2068 10.6151
R17592 vdd.n2068 vdd.n746 10.6151
R17593 vdd.n2216 vdd.n2215 10.6151
R17594 vdd.n2215 vdd.n2214 10.6151
R17595 vdd.n2214 vdd.n2211 10.6151
R17596 vdd.n2211 vdd.n2210 10.6151
R17597 vdd.n2210 vdd.n2207 10.6151
R17598 vdd.n2207 vdd.n2206 10.6151
R17599 vdd.n2206 vdd.n2203 10.6151
R17600 vdd.n2203 vdd.n2202 10.6151
R17601 vdd.n2202 vdd.n2199 10.6151
R17602 vdd.n2199 vdd.n2198 10.6151
R17603 vdd.n2198 vdd.n2195 10.6151
R17604 vdd.n2195 vdd.n2194 10.6151
R17605 vdd.n2194 vdd.n2191 10.6151
R17606 vdd.n2191 vdd.n2190 10.6151
R17607 vdd.n2190 vdd.n2187 10.6151
R17608 vdd.n2187 vdd.n2186 10.6151
R17609 vdd.n2186 vdd.n2183 10.6151
R17610 vdd.n2183 vdd.n2182 10.6151
R17611 vdd.n2182 vdd.n2179 10.6151
R17612 vdd.n2179 vdd.n2178 10.6151
R17613 vdd.n2178 vdd.n2175 10.6151
R17614 vdd.n2175 vdd.n2174 10.6151
R17615 vdd.n2174 vdd.n2171 10.6151
R17616 vdd.n2171 vdd.n2170 10.6151
R17617 vdd.n2170 vdd.n2167 10.6151
R17618 vdd.n2167 vdd.n2166 10.6151
R17619 vdd.n2166 vdd.n2163 10.6151
R17620 vdd.n2163 vdd.n2162 10.6151
R17621 vdd.n2162 vdd.n2159 10.6151
R17622 vdd.n2159 vdd.n2158 10.6151
R17623 vdd.n2158 vdd.n2155 10.6151
R17624 vdd.n2153 vdd.n2150 10.6151
R17625 vdd.n2150 vdd.n2149 10.6151
R17626 vdd.n1892 vdd.n1891 10.6151
R17627 vdd.n1891 vdd.n1889 10.6151
R17628 vdd.n1889 vdd.n1888 10.6151
R17629 vdd.n1888 vdd.n1886 10.6151
R17630 vdd.n1886 vdd.n1885 10.6151
R17631 vdd.n1885 vdd.n1883 10.6151
R17632 vdd.n1883 vdd.n1882 10.6151
R17633 vdd.n1882 vdd.n1880 10.6151
R17634 vdd.n1880 vdd.n1879 10.6151
R17635 vdd.n1879 vdd.n1877 10.6151
R17636 vdd.n1877 vdd.n1876 10.6151
R17637 vdd.n1876 vdd.n1874 10.6151
R17638 vdd.n1874 vdd.n1873 10.6151
R17639 vdd.n1873 vdd.n1788 10.6151
R17640 vdd.n1788 vdd.n1787 10.6151
R17641 vdd.n1787 vdd.n1785 10.6151
R17642 vdd.n1785 vdd.n1784 10.6151
R17643 vdd.n1784 vdd.n1782 10.6151
R17644 vdd.n1782 vdd.n1781 10.6151
R17645 vdd.n1781 vdd.n1779 10.6151
R17646 vdd.n1779 vdd.n1778 10.6151
R17647 vdd.n1778 vdd.n1776 10.6151
R17648 vdd.n1776 vdd.n1775 10.6151
R17649 vdd.n1775 vdd.n1773 10.6151
R17650 vdd.n1773 vdd.n1772 10.6151
R17651 vdd.n1772 vdd.n1769 10.6151
R17652 vdd.n1769 vdd.n1768 10.6151
R17653 vdd.n1768 vdd.n749 10.6151
R17654 vdd.n1726 vdd.n837 10.6151
R17655 vdd.n1727 vdd.n1726 10.6151
R17656 vdd.n1728 vdd.n1727 10.6151
R17657 vdd.n1728 vdd.n1722 10.6151
R17658 vdd.n1734 vdd.n1722 10.6151
R17659 vdd.n1735 vdd.n1734 10.6151
R17660 vdd.n1736 vdd.n1735 10.6151
R17661 vdd.n1736 vdd.n1720 10.6151
R17662 vdd.n1742 vdd.n1720 10.6151
R17663 vdd.n1743 vdd.n1742 10.6151
R17664 vdd.n1744 vdd.n1743 10.6151
R17665 vdd.n1744 vdd.n1718 10.6151
R17666 vdd.n1750 vdd.n1718 10.6151
R17667 vdd.n1751 vdd.n1750 10.6151
R17668 vdd.n1752 vdd.n1751 10.6151
R17669 vdd.n1752 vdd.n1716 10.6151
R17670 vdd.n1928 vdd.n1716 10.6151
R17671 vdd.n1928 vdd.n1927 10.6151
R17672 vdd.n1927 vdd.n1757 10.6151
R17673 vdd.n1921 vdd.n1757 10.6151
R17674 vdd.n1921 vdd.n1920 10.6151
R17675 vdd.n1920 vdd.n1919 10.6151
R17676 vdd.n1919 vdd.n1759 10.6151
R17677 vdd.n1913 vdd.n1759 10.6151
R17678 vdd.n1913 vdd.n1912 10.6151
R17679 vdd.n1912 vdd.n1911 10.6151
R17680 vdd.n1911 vdd.n1761 10.6151
R17681 vdd.n1905 vdd.n1761 10.6151
R17682 vdd.n1905 vdd.n1904 10.6151
R17683 vdd.n1904 vdd.n1903 10.6151
R17684 vdd.n1903 vdd.n1763 10.6151
R17685 vdd.n1897 vdd.n1896 10.6151
R17686 vdd.n1896 vdd.n1895 10.6151
R17687 vdd.n2401 vdd.n2400 10.6151
R17688 vdd.n2400 vdd.n2398 10.6151
R17689 vdd.n2398 vdd.n2397 10.6151
R17690 vdd.n2397 vdd.n2255 10.6151
R17691 vdd.n2344 vdd.n2255 10.6151
R17692 vdd.n2345 vdd.n2344 10.6151
R17693 vdd.n2347 vdd.n2345 10.6151
R17694 vdd.n2348 vdd.n2347 10.6151
R17695 vdd.n2350 vdd.n2348 10.6151
R17696 vdd.n2351 vdd.n2350 10.6151
R17697 vdd.n2353 vdd.n2351 10.6151
R17698 vdd.n2354 vdd.n2353 10.6151
R17699 vdd.n2356 vdd.n2354 10.6151
R17700 vdd.n2357 vdd.n2356 10.6151
R17701 vdd.n2372 vdd.n2357 10.6151
R17702 vdd.n2372 vdd.n2371 10.6151
R17703 vdd.n2371 vdd.n2370 10.6151
R17704 vdd.n2370 vdd.n2368 10.6151
R17705 vdd.n2368 vdd.n2367 10.6151
R17706 vdd.n2367 vdd.n2365 10.6151
R17707 vdd.n2365 vdd.n2364 10.6151
R17708 vdd.n2364 vdd.n2362 10.6151
R17709 vdd.n2362 vdd.n2361 10.6151
R17710 vdd.n2361 vdd.n2359 10.6151
R17711 vdd.n2359 vdd.n2358 10.6151
R17712 vdd.n2358 vdd.n626 10.6151
R17713 vdd.n2606 vdd.n626 10.6151
R17714 vdd.n2607 vdd.n2606 10.6151
R17715 vdd.n2468 vdd.n702 10.6151
R17716 vdd.n2468 vdd.n2467 10.6151
R17717 vdd.n2467 vdd.n2466 10.6151
R17718 vdd.n2466 vdd.n2464 10.6151
R17719 vdd.n2464 vdd.n2461 10.6151
R17720 vdd.n2461 vdd.n2460 10.6151
R17721 vdd.n2460 vdd.n2457 10.6151
R17722 vdd.n2457 vdd.n2456 10.6151
R17723 vdd.n2456 vdd.n2453 10.6151
R17724 vdd.n2453 vdd.n2452 10.6151
R17725 vdd.n2452 vdd.n2449 10.6151
R17726 vdd.n2449 vdd.n2448 10.6151
R17727 vdd.n2448 vdd.n2445 10.6151
R17728 vdd.n2445 vdd.n2444 10.6151
R17729 vdd.n2444 vdd.n2441 10.6151
R17730 vdd.n2441 vdd.n2440 10.6151
R17731 vdd.n2440 vdd.n2437 10.6151
R17732 vdd.n2437 vdd.n2436 10.6151
R17733 vdd.n2436 vdd.n2433 10.6151
R17734 vdd.n2433 vdd.n2432 10.6151
R17735 vdd.n2432 vdd.n2429 10.6151
R17736 vdd.n2429 vdd.n2428 10.6151
R17737 vdd.n2428 vdd.n2425 10.6151
R17738 vdd.n2425 vdd.n2424 10.6151
R17739 vdd.n2424 vdd.n2421 10.6151
R17740 vdd.n2421 vdd.n2420 10.6151
R17741 vdd.n2420 vdd.n2417 10.6151
R17742 vdd.n2417 vdd.n2416 10.6151
R17743 vdd.n2416 vdd.n2413 10.6151
R17744 vdd.n2413 vdd.n2412 10.6151
R17745 vdd.n2412 vdd.n2409 10.6151
R17746 vdd.n2407 vdd.n2404 10.6151
R17747 vdd.n2404 vdd.n2403 10.6151
R17748 vdd.n2481 vdd.n2480 10.6151
R17749 vdd.n2482 vdd.n2481 10.6151
R17750 vdd.n2482 vdd.n692 10.6151
R17751 vdd.n2492 vdd.n692 10.6151
R17752 vdd.n2493 vdd.n2492 10.6151
R17753 vdd.n2494 vdd.n2493 10.6151
R17754 vdd.n2494 vdd.n679 10.6151
R17755 vdd.n2504 vdd.n679 10.6151
R17756 vdd.n2505 vdd.n2504 10.6151
R17757 vdd.n2506 vdd.n2505 10.6151
R17758 vdd.n2506 vdd.n668 10.6151
R17759 vdd.n2516 vdd.n668 10.6151
R17760 vdd.n2517 vdd.n2516 10.6151
R17761 vdd.n2518 vdd.n2517 10.6151
R17762 vdd.n2518 vdd.n656 10.6151
R17763 vdd.n2528 vdd.n656 10.6151
R17764 vdd.n2529 vdd.n2528 10.6151
R17765 vdd.n2530 vdd.n2529 10.6151
R17766 vdd.n2530 vdd.n645 10.6151
R17767 vdd.n2542 vdd.n645 10.6151
R17768 vdd.n2543 vdd.n2542 10.6151
R17769 vdd.n2544 vdd.n2543 10.6151
R17770 vdd.n2544 vdd.n631 10.6151
R17771 vdd.n2599 vdd.n631 10.6151
R17772 vdd.n2600 vdd.n2599 10.6151
R17773 vdd.n2601 vdd.n2600 10.6151
R17774 vdd.n2601 vdd.n600 10.6151
R17775 vdd.n2671 vdd.n600 10.6151
R17776 vdd.n2670 vdd.n2669 10.6151
R17777 vdd.n2669 vdd.n601 10.6151
R17778 vdd.n602 vdd.n601 10.6151
R17779 vdd.n2662 vdd.n602 10.6151
R17780 vdd.n2662 vdd.n2661 10.6151
R17781 vdd.n2661 vdd.n2660 10.6151
R17782 vdd.n2660 vdd.n604 10.6151
R17783 vdd.n2655 vdd.n604 10.6151
R17784 vdd.n2655 vdd.n2654 10.6151
R17785 vdd.n2654 vdd.n2653 10.6151
R17786 vdd.n2653 vdd.n607 10.6151
R17787 vdd.n2648 vdd.n607 10.6151
R17788 vdd.n2648 vdd.n2647 10.6151
R17789 vdd.n2647 vdd.n2646 10.6151
R17790 vdd.n2646 vdd.n610 10.6151
R17791 vdd.n2641 vdd.n610 10.6151
R17792 vdd.n2641 vdd.n520 10.6151
R17793 vdd.n2637 vdd.n520 10.6151
R17794 vdd.n2637 vdd.n2636 10.6151
R17795 vdd.n2636 vdd.n2635 10.6151
R17796 vdd.n2635 vdd.n613 10.6151
R17797 vdd.n2630 vdd.n613 10.6151
R17798 vdd.n2630 vdd.n2629 10.6151
R17799 vdd.n2629 vdd.n2628 10.6151
R17800 vdd.n2628 vdd.n616 10.6151
R17801 vdd.n2623 vdd.n616 10.6151
R17802 vdd.n2623 vdd.n2622 10.6151
R17803 vdd.n2622 vdd.n2621 10.6151
R17804 vdd.n2621 vdd.n619 10.6151
R17805 vdd.n2616 vdd.n619 10.6151
R17806 vdd.n2616 vdd.n2615 10.6151
R17807 vdd.n2613 vdd.n624 10.6151
R17808 vdd.n2608 vdd.n624 10.6151
R17809 vdd.n2589 vdd.n2550 10.6151
R17810 vdd.n2584 vdd.n2550 10.6151
R17811 vdd.n2584 vdd.n2583 10.6151
R17812 vdd.n2583 vdd.n2582 10.6151
R17813 vdd.n2582 vdd.n2552 10.6151
R17814 vdd.n2577 vdd.n2552 10.6151
R17815 vdd.n2577 vdd.n2576 10.6151
R17816 vdd.n2576 vdd.n2575 10.6151
R17817 vdd.n2575 vdd.n2555 10.6151
R17818 vdd.n2570 vdd.n2555 10.6151
R17819 vdd.n2570 vdd.n2569 10.6151
R17820 vdd.n2569 vdd.n2568 10.6151
R17821 vdd.n2568 vdd.n2558 10.6151
R17822 vdd.n2563 vdd.n2558 10.6151
R17823 vdd.n2563 vdd.n2562 10.6151
R17824 vdd.n2562 vdd.n575 10.6151
R17825 vdd.n2706 vdd.n575 10.6151
R17826 vdd.n2706 vdd.n576 10.6151
R17827 vdd.n578 vdd.n576 10.6151
R17828 vdd.n2699 vdd.n578 10.6151
R17829 vdd.n2699 vdd.n2698 10.6151
R17830 vdd.n2698 vdd.n2697 10.6151
R17831 vdd.n2697 vdd.n580 10.6151
R17832 vdd.n2692 vdd.n580 10.6151
R17833 vdd.n2692 vdd.n2691 10.6151
R17834 vdd.n2691 vdd.n2690 10.6151
R17835 vdd.n2690 vdd.n583 10.6151
R17836 vdd.n2685 vdd.n583 10.6151
R17837 vdd.n2685 vdd.n2684 10.6151
R17838 vdd.n2684 vdd.n2683 10.6151
R17839 vdd.n2683 vdd.n586 10.6151
R17840 vdd.n2678 vdd.n2677 10.6151
R17841 vdd.n2677 vdd.n2676 10.6151
R17842 vdd.n2324 vdd.n2322 10.6151
R17843 vdd.n2325 vdd.n2324 10.6151
R17844 vdd.n2393 vdd.n2325 10.6151
R17845 vdd.n2393 vdd.n2392 10.6151
R17846 vdd.n2392 vdd.n2391 10.6151
R17847 vdd.n2391 vdd.n2389 10.6151
R17848 vdd.n2389 vdd.n2388 10.6151
R17849 vdd.n2388 vdd.n2386 10.6151
R17850 vdd.n2386 vdd.n2385 10.6151
R17851 vdd.n2385 vdd.n2383 10.6151
R17852 vdd.n2383 vdd.n2382 10.6151
R17853 vdd.n2382 vdd.n2380 10.6151
R17854 vdd.n2380 vdd.n2379 10.6151
R17855 vdd.n2379 vdd.n2377 10.6151
R17856 vdd.n2377 vdd.n2376 10.6151
R17857 vdd.n2376 vdd.n2342 10.6151
R17858 vdd.n2342 vdd.n2341 10.6151
R17859 vdd.n2341 vdd.n2339 10.6151
R17860 vdd.n2339 vdd.n2338 10.6151
R17861 vdd.n2338 vdd.n2336 10.6151
R17862 vdd.n2336 vdd.n2335 10.6151
R17863 vdd.n2335 vdd.n2333 10.6151
R17864 vdd.n2333 vdd.n2332 10.6151
R17865 vdd.n2332 vdd.n2330 10.6151
R17866 vdd.n2330 vdd.n2329 10.6151
R17867 vdd.n2329 vdd.n2327 10.6151
R17868 vdd.n2327 vdd.n2326 10.6151
R17869 vdd.n2326 vdd.n592 10.6151
R17870 vdd.n2475 vdd.n2474 10.6151
R17871 vdd.n2474 vdd.n707 10.6151
R17872 vdd.n2259 vdd.n707 10.6151
R17873 vdd.n2262 vdd.n2259 10.6151
R17874 vdd.n2263 vdd.n2262 10.6151
R17875 vdd.n2266 vdd.n2263 10.6151
R17876 vdd.n2267 vdd.n2266 10.6151
R17877 vdd.n2270 vdd.n2267 10.6151
R17878 vdd.n2271 vdd.n2270 10.6151
R17879 vdd.n2274 vdd.n2271 10.6151
R17880 vdd.n2275 vdd.n2274 10.6151
R17881 vdd.n2278 vdd.n2275 10.6151
R17882 vdd.n2279 vdd.n2278 10.6151
R17883 vdd.n2282 vdd.n2279 10.6151
R17884 vdd.n2283 vdd.n2282 10.6151
R17885 vdd.n2286 vdd.n2283 10.6151
R17886 vdd.n2287 vdd.n2286 10.6151
R17887 vdd.n2290 vdd.n2287 10.6151
R17888 vdd.n2291 vdd.n2290 10.6151
R17889 vdd.n2294 vdd.n2291 10.6151
R17890 vdd.n2295 vdd.n2294 10.6151
R17891 vdd.n2298 vdd.n2295 10.6151
R17892 vdd.n2299 vdd.n2298 10.6151
R17893 vdd.n2302 vdd.n2299 10.6151
R17894 vdd.n2303 vdd.n2302 10.6151
R17895 vdd.n2306 vdd.n2303 10.6151
R17896 vdd.n2307 vdd.n2306 10.6151
R17897 vdd.n2310 vdd.n2307 10.6151
R17898 vdd.n2311 vdd.n2310 10.6151
R17899 vdd.n2314 vdd.n2311 10.6151
R17900 vdd.n2315 vdd.n2314 10.6151
R17901 vdd.n2320 vdd.n2318 10.6151
R17902 vdd.n2321 vdd.n2320 10.6151
R17903 vdd.n2476 vdd.n697 10.6151
R17904 vdd.n2486 vdd.n697 10.6151
R17905 vdd.n2487 vdd.n2486 10.6151
R17906 vdd.n2488 vdd.n2487 10.6151
R17907 vdd.n2488 vdd.n685 10.6151
R17908 vdd.n2498 vdd.n685 10.6151
R17909 vdd.n2499 vdd.n2498 10.6151
R17910 vdd.n2500 vdd.n2499 10.6151
R17911 vdd.n2500 vdd.n674 10.6151
R17912 vdd.n2510 vdd.n674 10.6151
R17913 vdd.n2511 vdd.n2510 10.6151
R17914 vdd.n2512 vdd.n2511 10.6151
R17915 vdd.n2512 vdd.n662 10.6151
R17916 vdd.n2522 vdd.n662 10.6151
R17917 vdd.n2523 vdd.n2522 10.6151
R17918 vdd.n2524 vdd.n2523 10.6151
R17919 vdd.n2524 vdd.n651 10.6151
R17920 vdd.n2534 vdd.n651 10.6151
R17921 vdd.n2535 vdd.n2534 10.6151
R17922 vdd.n2538 vdd.n2535 10.6151
R17923 vdd.n2548 vdd.n639 10.6151
R17924 vdd.n2549 vdd.n2548 10.6151
R17925 vdd.n2595 vdd.n2549 10.6151
R17926 vdd.n2595 vdd.n2594 10.6151
R17927 vdd.n2594 vdd.n2593 10.6151
R17928 vdd.n2593 vdd.n2592 10.6151
R17929 vdd.n2592 vdd.n2590 10.6151
R17930 vdd.n1987 vdd.n831 10.6151
R17931 vdd.n1997 vdd.n831 10.6151
R17932 vdd.n1998 vdd.n1997 10.6151
R17933 vdd.n1999 vdd.n1998 10.6151
R17934 vdd.n1999 vdd.n818 10.6151
R17935 vdd.n2009 vdd.n818 10.6151
R17936 vdd.n2010 vdd.n2009 10.6151
R17937 vdd.n2012 vdd.n806 10.6151
R17938 vdd.n2022 vdd.n806 10.6151
R17939 vdd.n2023 vdd.n2022 10.6151
R17940 vdd.n2024 vdd.n2023 10.6151
R17941 vdd.n2024 vdd.n794 10.6151
R17942 vdd.n2034 vdd.n794 10.6151
R17943 vdd.n2035 vdd.n2034 10.6151
R17944 vdd.n2036 vdd.n2035 10.6151
R17945 vdd.n2036 vdd.n783 10.6151
R17946 vdd.n2046 vdd.n783 10.6151
R17947 vdd.n2047 vdd.n2046 10.6151
R17948 vdd.n2048 vdd.n2047 10.6151
R17949 vdd.n2048 vdd.n771 10.6151
R17950 vdd.n2058 vdd.n771 10.6151
R17951 vdd.n2059 vdd.n2058 10.6151
R17952 vdd.n2062 vdd.n2059 10.6151
R17953 vdd.n2062 vdd.n2061 10.6151
R17954 vdd.n2061 vdd.n2060 10.6151
R17955 vdd.n2060 vdd.n754 10.6151
R17956 vdd.n2144 vdd.n754 10.6151
R17957 vdd.n2143 vdd.n2142 10.6151
R17958 vdd.n2142 vdd.n2139 10.6151
R17959 vdd.n2139 vdd.n2138 10.6151
R17960 vdd.n2138 vdd.n2135 10.6151
R17961 vdd.n2135 vdd.n2134 10.6151
R17962 vdd.n2134 vdd.n2131 10.6151
R17963 vdd.n2131 vdd.n2130 10.6151
R17964 vdd.n2130 vdd.n2127 10.6151
R17965 vdd.n2127 vdd.n2126 10.6151
R17966 vdd.n2126 vdd.n2123 10.6151
R17967 vdd.n2123 vdd.n2122 10.6151
R17968 vdd.n2122 vdd.n2119 10.6151
R17969 vdd.n2119 vdd.n2118 10.6151
R17970 vdd.n2118 vdd.n2115 10.6151
R17971 vdd.n2115 vdd.n2114 10.6151
R17972 vdd.n2114 vdd.n2111 10.6151
R17973 vdd.n2111 vdd.n2110 10.6151
R17974 vdd.n2110 vdd.n2107 10.6151
R17975 vdd.n2107 vdd.n2106 10.6151
R17976 vdd.n2106 vdd.n2103 10.6151
R17977 vdd.n2103 vdd.n2102 10.6151
R17978 vdd.n2102 vdd.n2099 10.6151
R17979 vdd.n2099 vdd.n2098 10.6151
R17980 vdd.n2098 vdd.n2095 10.6151
R17981 vdd.n2095 vdd.n2094 10.6151
R17982 vdd.n2094 vdd.n2091 10.6151
R17983 vdd.n2091 vdd.n2090 10.6151
R17984 vdd.n2090 vdd.n2087 10.6151
R17985 vdd.n2087 vdd.n2086 10.6151
R17986 vdd.n2086 vdd.n2083 10.6151
R17987 vdd.n2083 vdd.n2082 10.6151
R17988 vdd.n2079 vdd.n2078 10.6151
R17989 vdd.n2078 vdd.n2076 10.6151
R17990 vdd.n1835 vdd.n1833 10.6151
R17991 vdd.n1836 vdd.n1835 10.6151
R17992 vdd.n1838 vdd.n1836 10.6151
R17993 vdd.n1839 vdd.n1838 10.6151
R17994 vdd.n1841 vdd.n1839 10.6151
R17995 vdd.n1842 vdd.n1841 10.6151
R17996 vdd.n1844 vdd.n1842 10.6151
R17997 vdd.n1845 vdd.n1844 10.6151
R17998 vdd.n1847 vdd.n1845 10.6151
R17999 vdd.n1848 vdd.n1847 10.6151
R18000 vdd.n1850 vdd.n1848 10.6151
R18001 vdd.n1851 vdd.n1850 10.6151
R18002 vdd.n1869 vdd.n1851 10.6151
R18003 vdd.n1869 vdd.n1868 10.6151
R18004 vdd.n1868 vdd.n1867 10.6151
R18005 vdd.n1867 vdd.n1865 10.6151
R18006 vdd.n1865 vdd.n1864 10.6151
R18007 vdd.n1864 vdd.n1862 10.6151
R18008 vdd.n1862 vdd.n1861 10.6151
R18009 vdd.n1861 vdd.n1859 10.6151
R18010 vdd.n1859 vdd.n1858 10.6151
R18011 vdd.n1858 vdd.n1856 10.6151
R18012 vdd.n1856 vdd.n1855 10.6151
R18013 vdd.n1855 vdd.n1853 10.6151
R18014 vdd.n1853 vdd.n1852 10.6151
R18015 vdd.n1852 vdd.n758 10.6151
R18016 vdd.n2074 vdd.n758 10.6151
R18017 vdd.n2075 vdd.n2074 10.6151
R18018 vdd.n1986 vdd.n1985 10.6151
R18019 vdd.n1985 vdd.n843 10.6151
R18020 vdd.n1979 vdd.n843 10.6151
R18021 vdd.n1979 vdd.n1978 10.6151
R18022 vdd.n1978 vdd.n1977 10.6151
R18023 vdd.n1977 vdd.n845 10.6151
R18024 vdd.n1971 vdd.n845 10.6151
R18025 vdd.n1971 vdd.n1970 10.6151
R18026 vdd.n1970 vdd.n1969 10.6151
R18027 vdd.n1969 vdd.n847 10.6151
R18028 vdd.n1963 vdd.n847 10.6151
R18029 vdd.n1963 vdd.n1962 10.6151
R18030 vdd.n1962 vdd.n1961 10.6151
R18031 vdd.n1961 vdd.n849 10.6151
R18032 vdd.n1955 vdd.n849 10.6151
R18033 vdd.n1955 vdd.n1954 10.6151
R18034 vdd.n1954 vdd.n1953 10.6151
R18035 vdd.n1953 vdd.n853 10.6151
R18036 vdd.n1801 vdd.n853 10.6151
R18037 vdd.n1802 vdd.n1801 10.6151
R18038 vdd.n1802 vdd.n1797 10.6151
R18039 vdd.n1808 vdd.n1797 10.6151
R18040 vdd.n1809 vdd.n1808 10.6151
R18041 vdd.n1810 vdd.n1809 10.6151
R18042 vdd.n1810 vdd.n1795 10.6151
R18043 vdd.n1816 vdd.n1795 10.6151
R18044 vdd.n1817 vdd.n1816 10.6151
R18045 vdd.n1818 vdd.n1817 10.6151
R18046 vdd.n1818 vdd.n1793 10.6151
R18047 vdd.n1824 vdd.n1793 10.6151
R18048 vdd.n1825 vdd.n1824 10.6151
R18049 vdd.n1827 vdd.n1789 10.6151
R18050 vdd.n1832 vdd.n1789 10.6151
R18051 vdd.n280 vdd.n262 10.4732
R18052 vdd.n233 vdd.n215 10.4732
R18053 vdd.n190 vdd.n172 10.4732
R18054 vdd.n143 vdd.n125 10.4732
R18055 vdd.n101 vdd.n83 10.4732
R18056 vdd.n54 vdd.n36 10.4732
R18057 vdd.n1095 vdd.n1077 10.4732
R18058 vdd.n1142 vdd.n1124 10.4732
R18059 vdd.n1005 vdd.n987 10.4732
R18060 vdd.n1052 vdd.n1034 10.4732
R18061 vdd.n916 vdd.n898 10.4732
R18062 vdd.n963 vdd.n945 10.4732
R18063 vdd.t105 vdd.n888 10.3167
R18064 vdd.n2874 vdd.t125 10.3167
R18065 vdd.n1465 vdd.t101 10.09
R18066 vdd.n3042 vdd.t138 10.09
R18067 vdd.n279 vdd.n264 9.69747
R18068 vdd.n232 vdd.n217 9.69747
R18069 vdd.n189 vdd.n174 9.69747
R18070 vdd.n142 vdd.n127 9.69747
R18071 vdd.n100 vdd.n85 9.69747
R18072 vdd.n53 vdd.n38 9.69747
R18073 vdd.n1094 vdd.n1079 9.69747
R18074 vdd.n1141 vdd.n1126 9.69747
R18075 vdd.n1004 vdd.n989 9.69747
R18076 vdd.n1051 vdd.n1036 9.69747
R18077 vdd.n915 vdd.n900 9.69747
R18078 vdd.n962 vdd.n947 9.69747
R18079 vdd.n1929 vdd.n1928 9.67831
R18080 vdd.n2836 vdd.n520 9.67831
R18081 vdd.n2707 vdd.n2706 9.67831
R18082 vdd.n1953 vdd.n1952 9.67831
R18083 vdd.n295 vdd.n294 9.45567
R18084 vdd.n248 vdd.n247 9.45567
R18085 vdd.n205 vdd.n204 9.45567
R18086 vdd.n158 vdd.n157 9.45567
R18087 vdd.n116 vdd.n115 9.45567
R18088 vdd.n69 vdd.n68 9.45567
R18089 vdd.n1110 vdd.n1109 9.45567
R18090 vdd.n1157 vdd.n1156 9.45567
R18091 vdd.n1020 vdd.n1019 9.45567
R18092 vdd.n1067 vdd.n1066 9.45567
R18093 vdd.n931 vdd.n930 9.45567
R18094 vdd.n978 vdd.n977 9.45567
R18095 vdd.n1689 vdd.n1543 9.3005
R18096 vdd.n1688 vdd.n1687 9.3005
R18097 vdd.n1549 vdd.n1548 9.3005
R18098 vdd.n1682 vdd.n1553 9.3005
R18099 vdd.n1681 vdd.n1554 9.3005
R18100 vdd.n1680 vdd.n1555 9.3005
R18101 vdd.n1559 vdd.n1556 9.3005
R18102 vdd.n1675 vdd.n1560 9.3005
R18103 vdd.n1674 vdd.n1561 9.3005
R18104 vdd.n1673 vdd.n1562 9.3005
R18105 vdd.n1566 vdd.n1563 9.3005
R18106 vdd.n1668 vdd.n1567 9.3005
R18107 vdd.n1667 vdd.n1568 9.3005
R18108 vdd.n1666 vdd.n1569 9.3005
R18109 vdd.n1573 vdd.n1570 9.3005
R18110 vdd.n1661 vdd.n1574 9.3005
R18111 vdd.n1660 vdd.n1575 9.3005
R18112 vdd.n1659 vdd.n1576 9.3005
R18113 vdd.n1580 vdd.n1577 9.3005
R18114 vdd.n1654 vdd.n1581 9.3005
R18115 vdd.n1653 vdd.n1582 9.3005
R18116 vdd.n1652 vdd.n1651 9.3005
R18117 vdd.n1650 vdd.n1583 9.3005
R18118 vdd.n1649 vdd.n1648 9.3005
R18119 vdd.n1589 vdd.n1588 9.3005
R18120 vdd.n1643 vdd.n1593 9.3005
R18121 vdd.n1642 vdd.n1594 9.3005
R18122 vdd.n1641 vdd.n1595 9.3005
R18123 vdd.n1599 vdd.n1596 9.3005
R18124 vdd.n1636 vdd.n1600 9.3005
R18125 vdd.n1635 vdd.n1601 9.3005
R18126 vdd.n1634 vdd.n1602 9.3005
R18127 vdd.n1606 vdd.n1603 9.3005
R18128 vdd.n1629 vdd.n1607 9.3005
R18129 vdd.n1628 vdd.n1608 9.3005
R18130 vdd.n1627 vdd.n1609 9.3005
R18131 vdd.n1611 vdd.n1610 9.3005
R18132 vdd.n1622 vdd.n854 9.3005
R18133 vdd.n1691 vdd.n1690 9.3005
R18134 vdd.n1715 vdd.n1714 9.3005
R18135 vdd.n1521 vdd.n1520 9.3005
R18136 vdd.n1526 vdd.n1524 9.3005
R18137 vdd.n1707 vdd.n1527 9.3005
R18138 vdd.n1706 vdd.n1528 9.3005
R18139 vdd.n1705 vdd.n1529 9.3005
R18140 vdd.n1533 vdd.n1530 9.3005
R18141 vdd.n1700 vdd.n1534 9.3005
R18142 vdd.n1699 vdd.n1535 9.3005
R18143 vdd.n1698 vdd.n1536 9.3005
R18144 vdd.n1540 vdd.n1537 9.3005
R18145 vdd.n1693 vdd.n1541 9.3005
R18146 vdd.n1692 vdd.n1542 9.3005
R18147 vdd.n1937 vdd.n1514 9.3005
R18148 vdd.n1939 vdd.n1938 9.3005
R18149 vdd.n1476 vdd.n1475 9.3005
R18150 vdd.n1477 vdd.n890 9.3005
R18151 vdd.n1479 vdd.n1478 9.3005
R18152 vdd.n880 vdd.n879 9.3005
R18153 vdd.n1493 vdd.n1492 9.3005
R18154 vdd.n1494 vdd.n878 9.3005
R18155 vdd.n1496 vdd.n1495 9.3005
R18156 vdd.n868 vdd.n867 9.3005
R18157 vdd.n1512 vdd.n1511 9.3005
R18158 vdd.n1513 vdd.n866 9.3005
R18159 vdd.n1941 vdd.n1940 9.3005
R18160 vdd.n271 vdd.n270 9.3005
R18161 vdd.n266 vdd.n265 9.3005
R18162 vdd.n277 vdd.n276 9.3005
R18163 vdd.n279 vdd.n278 9.3005
R18164 vdd.n262 vdd.n261 9.3005
R18165 vdd.n285 vdd.n284 9.3005
R18166 vdd.n287 vdd.n286 9.3005
R18167 vdd.n259 vdd.n256 9.3005
R18168 vdd.n294 vdd.n293 9.3005
R18169 vdd.n224 vdd.n223 9.3005
R18170 vdd.n219 vdd.n218 9.3005
R18171 vdd.n230 vdd.n229 9.3005
R18172 vdd.n232 vdd.n231 9.3005
R18173 vdd.n215 vdd.n214 9.3005
R18174 vdd.n238 vdd.n237 9.3005
R18175 vdd.n240 vdd.n239 9.3005
R18176 vdd.n212 vdd.n209 9.3005
R18177 vdd.n247 vdd.n246 9.3005
R18178 vdd.n181 vdd.n180 9.3005
R18179 vdd.n176 vdd.n175 9.3005
R18180 vdd.n187 vdd.n186 9.3005
R18181 vdd.n189 vdd.n188 9.3005
R18182 vdd.n172 vdd.n171 9.3005
R18183 vdd.n195 vdd.n194 9.3005
R18184 vdd.n197 vdd.n196 9.3005
R18185 vdd.n169 vdd.n166 9.3005
R18186 vdd.n204 vdd.n203 9.3005
R18187 vdd.n134 vdd.n133 9.3005
R18188 vdd.n129 vdd.n128 9.3005
R18189 vdd.n140 vdd.n139 9.3005
R18190 vdd.n142 vdd.n141 9.3005
R18191 vdd.n125 vdd.n124 9.3005
R18192 vdd.n148 vdd.n147 9.3005
R18193 vdd.n150 vdd.n149 9.3005
R18194 vdd.n122 vdd.n119 9.3005
R18195 vdd.n157 vdd.n156 9.3005
R18196 vdd.n92 vdd.n91 9.3005
R18197 vdd.n87 vdd.n86 9.3005
R18198 vdd.n98 vdd.n97 9.3005
R18199 vdd.n100 vdd.n99 9.3005
R18200 vdd.n83 vdd.n82 9.3005
R18201 vdd.n106 vdd.n105 9.3005
R18202 vdd.n108 vdd.n107 9.3005
R18203 vdd.n80 vdd.n77 9.3005
R18204 vdd.n115 vdd.n114 9.3005
R18205 vdd.n45 vdd.n44 9.3005
R18206 vdd.n40 vdd.n39 9.3005
R18207 vdd.n51 vdd.n50 9.3005
R18208 vdd.n53 vdd.n52 9.3005
R18209 vdd.n36 vdd.n35 9.3005
R18210 vdd.n59 vdd.n58 9.3005
R18211 vdd.n61 vdd.n60 9.3005
R18212 vdd.n33 vdd.n30 9.3005
R18213 vdd.n68 vdd.n67 9.3005
R18214 vdd.n2758 vdd.n2757 9.3005
R18215 vdd.n2761 vdd.n555 9.3005
R18216 vdd.n2762 vdd.n554 9.3005
R18217 vdd.n2765 vdd.n553 9.3005
R18218 vdd.n2766 vdd.n552 9.3005
R18219 vdd.n2769 vdd.n551 9.3005
R18220 vdd.n2770 vdd.n550 9.3005
R18221 vdd.n2773 vdd.n549 9.3005
R18222 vdd.n2774 vdd.n548 9.3005
R18223 vdd.n2777 vdd.n547 9.3005
R18224 vdd.n2778 vdd.n546 9.3005
R18225 vdd.n2781 vdd.n545 9.3005
R18226 vdd.n2782 vdd.n544 9.3005
R18227 vdd.n2785 vdd.n543 9.3005
R18228 vdd.n2786 vdd.n542 9.3005
R18229 vdd.n2789 vdd.n541 9.3005
R18230 vdd.n2790 vdd.n540 9.3005
R18231 vdd.n2793 vdd.n539 9.3005
R18232 vdd.n2794 vdd.n538 9.3005
R18233 vdd.n2797 vdd.n537 9.3005
R18234 vdd.n2801 vdd.n2800 9.3005
R18235 vdd.n2802 vdd.n536 9.3005
R18236 vdd.n2806 vdd.n2803 9.3005
R18237 vdd.n2809 vdd.n535 9.3005
R18238 vdd.n2810 vdd.n534 9.3005
R18239 vdd.n2813 vdd.n533 9.3005
R18240 vdd.n2814 vdd.n532 9.3005
R18241 vdd.n2817 vdd.n531 9.3005
R18242 vdd.n2818 vdd.n530 9.3005
R18243 vdd.n2821 vdd.n529 9.3005
R18244 vdd.n2822 vdd.n528 9.3005
R18245 vdd.n2825 vdd.n527 9.3005
R18246 vdd.n2826 vdd.n526 9.3005
R18247 vdd.n2829 vdd.n525 9.3005
R18248 vdd.n2830 vdd.n524 9.3005
R18249 vdd.n2833 vdd.n519 9.3005
R18250 vdd.n482 vdd.n481 9.3005
R18251 vdd.n2844 vdd.n2843 9.3005
R18252 vdd.n2847 vdd.n2846 9.3005
R18253 vdd.n471 vdd.n470 9.3005
R18254 vdd.n2861 vdd.n2860 9.3005
R18255 vdd.n2862 vdd.n469 9.3005
R18256 vdd.n2864 vdd.n2863 9.3005
R18257 vdd.n460 vdd.n459 9.3005
R18258 vdd.n2877 vdd.n2876 9.3005
R18259 vdd.n2878 vdd.n458 9.3005
R18260 vdd.n2880 vdd.n2879 9.3005
R18261 vdd.n300 vdd.n298 9.3005
R18262 vdd.n2845 vdd.n480 9.3005
R18263 vdd.n3046 vdd.n3045 9.3005
R18264 vdd.n301 vdd.n299 9.3005
R18265 vdd.n3039 vdd.n310 9.3005
R18266 vdd.n3038 vdd.n311 9.3005
R18267 vdd.n3037 vdd.n312 9.3005
R18268 vdd.n320 vdd.n313 9.3005
R18269 vdd.n3031 vdd.n321 9.3005
R18270 vdd.n3030 vdd.n322 9.3005
R18271 vdd.n3029 vdd.n323 9.3005
R18272 vdd.n331 vdd.n324 9.3005
R18273 vdd.n3023 vdd.n3022 9.3005
R18274 vdd.n3019 vdd.n332 9.3005
R18275 vdd.n3018 vdd.n335 9.3005
R18276 vdd.n339 vdd.n336 9.3005
R18277 vdd.n340 vdd.n337 9.3005
R18278 vdd.n3011 vdd.n341 9.3005
R18279 vdd.n3010 vdd.n342 9.3005
R18280 vdd.n3009 vdd.n343 9.3005
R18281 vdd.n347 vdd.n344 9.3005
R18282 vdd.n3004 vdd.n348 9.3005
R18283 vdd.n3003 vdd.n349 9.3005
R18284 vdd.n3002 vdd.n350 9.3005
R18285 vdd.n354 vdd.n351 9.3005
R18286 vdd.n2997 vdd.n355 9.3005
R18287 vdd.n2996 vdd.n356 9.3005
R18288 vdd.n2995 vdd.n357 9.3005
R18289 vdd.n361 vdd.n358 9.3005
R18290 vdd.n2990 vdd.n362 9.3005
R18291 vdd.n2989 vdd.n363 9.3005
R18292 vdd.n2988 vdd.n2987 9.3005
R18293 vdd.n2986 vdd.n364 9.3005
R18294 vdd.n2985 vdd.n2984 9.3005
R18295 vdd.n370 vdd.n369 9.3005
R18296 vdd.n2979 vdd.n374 9.3005
R18297 vdd.n2978 vdd.n375 9.3005
R18298 vdd.n2977 vdd.n376 9.3005
R18299 vdd.n380 vdd.n377 9.3005
R18300 vdd.n2972 vdd.n381 9.3005
R18301 vdd.n2971 vdd.n382 9.3005
R18302 vdd.n2970 vdd.n383 9.3005
R18303 vdd.n387 vdd.n384 9.3005
R18304 vdd.n2965 vdd.n388 9.3005
R18305 vdd.n2964 vdd.n389 9.3005
R18306 vdd.n2963 vdd.n390 9.3005
R18307 vdd.n394 vdd.n391 9.3005
R18308 vdd.n2958 vdd.n395 9.3005
R18309 vdd.n2957 vdd.n396 9.3005
R18310 vdd.n2956 vdd.n397 9.3005
R18311 vdd.n401 vdd.n398 9.3005
R18312 vdd.n2951 vdd.n402 9.3005
R18313 vdd.n2950 vdd.n403 9.3005
R18314 vdd.n2949 vdd.n2948 9.3005
R18315 vdd.n2947 vdd.n404 9.3005
R18316 vdd.n2946 vdd.n2945 9.3005
R18317 vdd.n410 vdd.n409 9.3005
R18318 vdd.n2940 vdd.n414 9.3005
R18319 vdd.n2939 vdd.n415 9.3005
R18320 vdd.n2938 vdd.n416 9.3005
R18321 vdd.n420 vdd.n417 9.3005
R18322 vdd.n2933 vdd.n421 9.3005
R18323 vdd.n2932 vdd.n422 9.3005
R18324 vdd.n2931 vdd.n423 9.3005
R18325 vdd.n427 vdd.n424 9.3005
R18326 vdd.n2926 vdd.n428 9.3005
R18327 vdd.n2925 vdd.n429 9.3005
R18328 vdd.n2924 vdd.n430 9.3005
R18329 vdd.n434 vdd.n431 9.3005
R18330 vdd.n2919 vdd.n435 9.3005
R18331 vdd.n2918 vdd.n436 9.3005
R18332 vdd.n2917 vdd.n437 9.3005
R18333 vdd.n441 vdd.n438 9.3005
R18334 vdd.n2912 vdd.n442 9.3005
R18335 vdd.n2911 vdd.n443 9.3005
R18336 vdd.n2907 vdd.n2904 9.3005
R18337 vdd.n3021 vdd.n3020 9.3005
R18338 vdd.n2852 vdd.n2851 9.3005
R18339 vdd.n2853 vdd.n475 9.3005
R18340 vdd.n2855 vdd.n2854 9.3005
R18341 vdd.n465 vdd.n464 9.3005
R18342 vdd.n2869 vdd.n2868 9.3005
R18343 vdd.n2870 vdd.n463 9.3005
R18344 vdd.n2872 vdd.n2871 9.3005
R18345 vdd.n453 vdd.n452 9.3005
R18346 vdd.n2885 vdd.n2884 9.3005
R18347 vdd.n2886 vdd.n451 9.3005
R18348 vdd.n2888 vdd.n2887 9.3005
R18349 vdd.n2889 vdd.n450 9.3005
R18350 vdd.n2891 vdd.n2890 9.3005
R18351 vdd.n2892 vdd.n449 9.3005
R18352 vdd.n2894 vdd.n2893 9.3005
R18353 vdd.n2895 vdd.n447 9.3005
R18354 vdd.n2897 vdd.n2896 9.3005
R18355 vdd.n2898 vdd.n446 9.3005
R18356 vdd.n2900 vdd.n2899 9.3005
R18357 vdd.n2901 vdd.n444 9.3005
R18358 vdd.n2903 vdd.n2902 9.3005
R18359 vdd.n477 vdd.n476 9.3005
R18360 vdd.n2710 vdd.n2709 9.3005
R18361 vdd.n2715 vdd.n2708 9.3005
R18362 vdd.n2724 vdd.n572 9.3005
R18363 vdd.n2727 vdd.n571 9.3005
R18364 vdd.n2728 vdd.n570 9.3005
R18365 vdd.n2731 vdd.n569 9.3005
R18366 vdd.n2732 vdd.n568 9.3005
R18367 vdd.n2735 vdd.n567 9.3005
R18368 vdd.n2736 vdd.n566 9.3005
R18369 vdd.n2739 vdd.n565 9.3005
R18370 vdd.n2740 vdd.n564 9.3005
R18371 vdd.n2743 vdd.n563 9.3005
R18372 vdd.n2744 vdd.n562 9.3005
R18373 vdd.n2747 vdd.n561 9.3005
R18374 vdd.n2748 vdd.n560 9.3005
R18375 vdd.n2751 vdd.n559 9.3005
R18376 vdd.n2755 vdd.n2754 9.3005
R18377 vdd.n2756 vdd.n556 9.3005
R18378 vdd.n1951 vdd.n1950 9.3005
R18379 vdd.n1946 vdd.n857 9.3005
R18380 vdd.n1433 vdd.n1432 9.3005
R18381 vdd.n1434 vdd.n1188 9.3005
R18382 vdd.n1436 vdd.n1435 9.3005
R18383 vdd.n1178 vdd.n1177 9.3005
R18384 vdd.n1450 vdd.n1449 9.3005
R18385 vdd.n1451 vdd.n1176 9.3005
R18386 vdd.n1453 vdd.n1452 9.3005
R18387 vdd.n1168 vdd.n1167 9.3005
R18388 vdd.n1468 vdd.n1467 9.3005
R18389 vdd.n1469 vdd.n1166 9.3005
R18390 vdd.n1471 vdd.n1470 9.3005
R18391 vdd.n885 vdd.n884 9.3005
R18392 vdd.n1484 vdd.n1483 9.3005
R18393 vdd.n1485 vdd.n883 9.3005
R18394 vdd.n1487 vdd.n1486 9.3005
R18395 vdd.n875 vdd.n874 9.3005
R18396 vdd.n1501 vdd.n1500 9.3005
R18397 vdd.n1502 vdd.n872 9.3005
R18398 vdd.n1506 vdd.n1505 9.3005
R18399 vdd.n1504 vdd.n873 9.3005
R18400 vdd.n1503 vdd.n862 9.3005
R18401 vdd.n1190 vdd.n1189 9.3005
R18402 vdd.n1326 vdd.n1325 9.3005
R18403 vdd.n1327 vdd.n1316 9.3005
R18404 vdd.n1329 vdd.n1328 9.3005
R18405 vdd.n1330 vdd.n1315 9.3005
R18406 vdd.n1332 vdd.n1331 9.3005
R18407 vdd.n1333 vdd.n1310 9.3005
R18408 vdd.n1335 vdd.n1334 9.3005
R18409 vdd.n1336 vdd.n1309 9.3005
R18410 vdd.n1338 vdd.n1337 9.3005
R18411 vdd.n1339 vdd.n1304 9.3005
R18412 vdd.n1341 vdd.n1340 9.3005
R18413 vdd.n1342 vdd.n1303 9.3005
R18414 vdd.n1344 vdd.n1343 9.3005
R18415 vdd.n1345 vdd.n1298 9.3005
R18416 vdd.n1347 vdd.n1346 9.3005
R18417 vdd.n1348 vdd.n1297 9.3005
R18418 vdd.n1350 vdd.n1349 9.3005
R18419 vdd.n1351 vdd.n1292 9.3005
R18420 vdd.n1353 vdd.n1352 9.3005
R18421 vdd.n1354 vdd.n1291 9.3005
R18422 vdd.n1356 vdd.n1355 9.3005
R18423 vdd.n1360 vdd.n1287 9.3005
R18424 vdd.n1362 vdd.n1361 9.3005
R18425 vdd.n1363 vdd.n1286 9.3005
R18426 vdd.n1365 vdd.n1364 9.3005
R18427 vdd.n1366 vdd.n1281 9.3005
R18428 vdd.n1368 vdd.n1367 9.3005
R18429 vdd.n1369 vdd.n1280 9.3005
R18430 vdd.n1371 vdd.n1370 9.3005
R18431 vdd.n1372 vdd.n1275 9.3005
R18432 vdd.n1374 vdd.n1373 9.3005
R18433 vdd.n1375 vdd.n1274 9.3005
R18434 vdd.n1377 vdd.n1376 9.3005
R18435 vdd.n1378 vdd.n1269 9.3005
R18436 vdd.n1380 vdd.n1379 9.3005
R18437 vdd.n1381 vdd.n1268 9.3005
R18438 vdd.n1383 vdd.n1382 9.3005
R18439 vdd.n1384 vdd.n1263 9.3005
R18440 vdd.n1386 vdd.n1385 9.3005
R18441 vdd.n1387 vdd.n1262 9.3005
R18442 vdd.n1389 vdd.n1388 9.3005
R18443 vdd.n1390 vdd.n1257 9.3005
R18444 vdd.n1392 vdd.n1391 9.3005
R18445 vdd.n1393 vdd.n1256 9.3005
R18446 vdd.n1395 vdd.n1394 9.3005
R18447 vdd.n1396 vdd.n1249 9.3005
R18448 vdd.n1398 vdd.n1397 9.3005
R18449 vdd.n1399 vdd.n1248 9.3005
R18450 vdd.n1401 vdd.n1400 9.3005
R18451 vdd.n1402 vdd.n1243 9.3005
R18452 vdd.n1404 vdd.n1403 9.3005
R18453 vdd.n1405 vdd.n1242 9.3005
R18454 vdd.n1407 vdd.n1406 9.3005
R18455 vdd.n1408 vdd.n1237 9.3005
R18456 vdd.n1410 vdd.n1409 9.3005
R18457 vdd.n1411 vdd.n1236 9.3005
R18458 vdd.n1413 vdd.n1412 9.3005
R18459 vdd.n1414 vdd.n1231 9.3005
R18460 vdd.n1416 vdd.n1415 9.3005
R18461 vdd.n1417 vdd.n1230 9.3005
R18462 vdd.n1419 vdd.n1418 9.3005
R18463 vdd.n1195 vdd.n1194 9.3005
R18464 vdd.n1425 vdd.n1424 9.3005
R18465 vdd.n1324 vdd.n1323 9.3005
R18466 vdd.n1428 vdd.n1427 9.3005
R18467 vdd.n1184 vdd.n1183 9.3005
R18468 vdd.n1442 vdd.n1441 9.3005
R18469 vdd.n1443 vdd.n1182 9.3005
R18470 vdd.n1445 vdd.n1444 9.3005
R18471 vdd.n1173 vdd.n1172 9.3005
R18472 vdd.n1459 vdd.n1458 9.3005
R18473 vdd.n1460 vdd.n1171 9.3005
R18474 vdd.n1463 vdd.n1462 9.3005
R18475 vdd.n1461 vdd.n1162 9.3005
R18476 vdd.n1426 vdd.n1193 9.3005
R18477 vdd.n1086 vdd.n1085 9.3005
R18478 vdd.n1081 vdd.n1080 9.3005
R18479 vdd.n1092 vdd.n1091 9.3005
R18480 vdd.n1094 vdd.n1093 9.3005
R18481 vdd.n1077 vdd.n1076 9.3005
R18482 vdd.n1100 vdd.n1099 9.3005
R18483 vdd.n1102 vdd.n1101 9.3005
R18484 vdd.n1074 vdd.n1071 9.3005
R18485 vdd.n1109 vdd.n1108 9.3005
R18486 vdd.n1133 vdd.n1132 9.3005
R18487 vdd.n1128 vdd.n1127 9.3005
R18488 vdd.n1139 vdd.n1138 9.3005
R18489 vdd.n1141 vdd.n1140 9.3005
R18490 vdd.n1124 vdd.n1123 9.3005
R18491 vdd.n1147 vdd.n1146 9.3005
R18492 vdd.n1149 vdd.n1148 9.3005
R18493 vdd.n1121 vdd.n1118 9.3005
R18494 vdd.n1156 vdd.n1155 9.3005
R18495 vdd.n996 vdd.n995 9.3005
R18496 vdd.n991 vdd.n990 9.3005
R18497 vdd.n1002 vdd.n1001 9.3005
R18498 vdd.n1004 vdd.n1003 9.3005
R18499 vdd.n987 vdd.n986 9.3005
R18500 vdd.n1010 vdd.n1009 9.3005
R18501 vdd.n1012 vdd.n1011 9.3005
R18502 vdd.n984 vdd.n981 9.3005
R18503 vdd.n1019 vdd.n1018 9.3005
R18504 vdd.n1043 vdd.n1042 9.3005
R18505 vdd.n1038 vdd.n1037 9.3005
R18506 vdd.n1049 vdd.n1048 9.3005
R18507 vdd.n1051 vdd.n1050 9.3005
R18508 vdd.n1034 vdd.n1033 9.3005
R18509 vdd.n1057 vdd.n1056 9.3005
R18510 vdd.n1059 vdd.n1058 9.3005
R18511 vdd.n1031 vdd.n1028 9.3005
R18512 vdd.n1066 vdd.n1065 9.3005
R18513 vdd.n907 vdd.n906 9.3005
R18514 vdd.n902 vdd.n901 9.3005
R18515 vdd.n913 vdd.n912 9.3005
R18516 vdd.n915 vdd.n914 9.3005
R18517 vdd.n898 vdd.n897 9.3005
R18518 vdd.n921 vdd.n920 9.3005
R18519 vdd.n923 vdd.n922 9.3005
R18520 vdd.n895 vdd.n892 9.3005
R18521 vdd.n930 vdd.n929 9.3005
R18522 vdd.n954 vdd.n953 9.3005
R18523 vdd.n949 vdd.n948 9.3005
R18524 vdd.n960 vdd.n959 9.3005
R18525 vdd.n962 vdd.n961 9.3005
R18526 vdd.n945 vdd.n944 9.3005
R18527 vdd.n968 vdd.n967 9.3005
R18528 vdd.n970 vdd.n969 9.3005
R18529 vdd.n942 vdd.n939 9.3005
R18530 vdd.n977 vdd.n976 9.3005
R18531 vdd.n1438 vdd.t134 8.95635
R18532 vdd.t116 vdd.n3033 8.95635
R18533 vdd.n276 vdd.n275 8.92171
R18534 vdd.n229 vdd.n228 8.92171
R18535 vdd.n186 vdd.n185 8.92171
R18536 vdd.n139 vdd.n138 8.92171
R18537 vdd.n97 vdd.n96 8.92171
R18538 vdd.n50 vdd.n49 8.92171
R18539 vdd.n1091 vdd.n1090 8.92171
R18540 vdd.n1138 vdd.n1137 8.92171
R18541 vdd.n1001 vdd.n1000 8.92171
R18542 vdd.n1048 vdd.n1047 8.92171
R18543 vdd.n912 vdd.n911 8.92171
R18544 vdd.n959 vdd.n958 8.92171
R18545 vdd.n207 vdd.n117 8.81535
R18546 vdd.n1069 vdd.n979 8.81535
R18547 vdd.n1465 vdd.t112 8.72962
R18548 vdd.t114 vdd.n3042 8.72962
R18549 vdd.n888 vdd.t150 8.50289
R18550 vdd.n1943 vdd.t29 8.50289
R18551 vdd.n516 vdd.t22 8.50289
R18552 vdd.n2874 vdd.t128 8.50289
R18553 vdd.n28 vdd.n14 8.42249
R18554 vdd.n3048 vdd.n3047 8.16225
R18555 vdd.n1161 vdd.n1160 8.16225
R18556 vdd.n272 vdd.n266 8.14595
R18557 vdd.n225 vdd.n219 8.14595
R18558 vdd.n182 vdd.n176 8.14595
R18559 vdd.n135 vdd.n129 8.14595
R18560 vdd.n93 vdd.n87 8.14595
R18561 vdd.n46 vdd.n40 8.14595
R18562 vdd.n1087 vdd.n1081 8.14595
R18563 vdd.n1134 vdd.n1128 8.14595
R18564 vdd.n997 vdd.n991 8.14595
R18565 vdd.n1044 vdd.n1038 8.14595
R18566 vdd.n908 vdd.n902 8.14595
R18567 vdd.n955 vdd.n949 8.14595
R18568 vdd.n2537 vdd.n639 8.11757
R18569 vdd.n2011 vdd.n2010 8.11757
R18570 vdd.n1989 vdd.n833 7.70933
R18571 vdd.n1995 vdd.n833 7.70933
R18572 vdd.n2001 vdd.n827 7.70933
R18573 vdd.n2001 vdd.n820 7.70933
R18574 vdd.n2007 vdd.n820 7.70933
R18575 vdd.n2007 vdd.n823 7.70933
R18576 vdd.n2014 vdd.n808 7.70933
R18577 vdd.n2020 vdd.n808 7.70933
R18578 vdd.n2026 vdd.n802 7.70933
R18579 vdd.n2032 vdd.n798 7.70933
R18580 vdd.n2038 vdd.n792 7.70933
R18581 vdd.n2050 vdd.n779 7.70933
R18582 vdd.n2056 vdd.n773 7.70933
R18583 vdd.n2056 vdd.n766 7.70933
R18584 vdd.n2064 vdd.n766 7.70933
R18585 vdd.n2071 vdd.t19 7.70933
R18586 vdd.n2146 vdd.t19 7.70933
R18587 vdd.n2478 vdd.t196 7.70933
R18588 vdd.n2484 vdd.t196 7.70933
R18589 vdd.n2490 vdd.n687 7.70933
R18590 vdd.n2496 vdd.n687 7.70933
R18591 vdd.n2496 vdd.n690 7.70933
R18592 vdd.n2502 vdd.n683 7.70933
R18593 vdd.n2514 vdd.n670 7.70933
R18594 vdd.n2520 vdd.n664 7.70933
R18595 vdd.n2526 vdd.n660 7.70933
R18596 vdd.n2532 vdd.n647 7.70933
R18597 vdd.n2540 vdd.n647 7.70933
R18598 vdd.n2546 vdd.n641 7.70933
R18599 vdd.n2546 vdd.n633 7.70933
R18600 vdd.n2597 vdd.n633 7.70933
R18601 vdd.n2597 vdd.n636 7.70933
R18602 vdd.n2603 vdd.n595 7.70933
R18603 vdd.n2673 vdd.n595 7.70933
R18604 vdd.n271 vdd.n268 7.3702
R18605 vdd.n224 vdd.n221 7.3702
R18606 vdd.n181 vdd.n178 7.3702
R18607 vdd.n134 vdd.n131 7.3702
R18608 vdd.n92 vdd.n89 7.3702
R18609 vdd.n45 vdd.n42 7.3702
R18610 vdd.n1086 vdd.n1083 7.3702
R18611 vdd.n1133 vdd.n1130 7.3702
R18612 vdd.n996 vdd.n993 7.3702
R18613 vdd.n1043 vdd.n1040 7.3702
R18614 vdd.n907 vdd.n904 7.3702
R18615 vdd.n954 vdd.n951 7.3702
R18616 vdd.n1361 vdd.n1360 6.98232
R18617 vdd.n1653 vdd.n1652 6.98232
R18618 vdd.n2950 vdd.n2949 6.98232
R18619 vdd.n2761 vdd.n2758 6.98232
R18620 vdd.n1498 vdd.t97 6.68904
R18621 vdd.n2857 vdd.t99 6.68904
R18622 vdd.t136 vdd.n887 6.46231
R18623 vdd.n2882 vdd.t103 6.46231
R18624 vdd.n1456 vdd.t118 6.23558
R18625 vdd.t107 vdd.n308 6.23558
R18626 vdd.n3048 vdd.n297 6.22547
R18627 vdd.n1160 vdd.n1159 6.22547
R18628 vdd.n2026 vdd.t177 6.00885
R18629 vdd.n2526 vdd.t14 6.00885
R18630 vdd.n823 vdd.t73 5.89549
R18631 vdd.t37 vdd.n641 5.89549
R18632 vdd.n272 vdd.n271 5.81868
R18633 vdd.n225 vdd.n224 5.81868
R18634 vdd.n182 vdd.n181 5.81868
R18635 vdd.n135 vdd.n134 5.81868
R18636 vdd.n93 vdd.n92 5.81868
R18637 vdd.n46 vdd.n45 5.81868
R18638 vdd.n1087 vdd.n1086 5.81868
R18639 vdd.n1134 vdd.n1133 5.81868
R18640 vdd.n997 vdd.n996 5.81868
R18641 vdd.n1044 vdd.n1043 5.81868
R18642 vdd.n908 vdd.n907 5.81868
R18643 vdd.n955 vdd.n954 5.81868
R18644 vdd.t69 vdd.n827 5.78212
R18645 vdd.n1770 vdd.t54 5.78212
R18646 vdd.n2395 vdd.t62 5.78212
R18647 vdd.n636 vdd.t58 5.78212
R18648 vdd.n2154 vdd.n2153 5.77611
R18649 vdd.n1897 vdd.n1767 5.77611
R18650 vdd.n2408 vdd.n2407 5.77611
R18651 vdd.n2614 vdd.n2613 5.77611
R18652 vdd.n2678 vdd.n591 5.77611
R18653 vdd.n2318 vdd.n2258 5.77611
R18654 vdd.n2079 vdd.n757 5.77611
R18655 vdd.n1827 vdd.n1826 5.77611
R18656 vdd.n1323 vdd.n1322 5.62474
R18657 vdd.n1949 vdd.n1946 5.62474
R18658 vdd.n2910 vdd.n2907 5.62474
R18659 vdd.n2713 vdd.n2710 5.62474
R18660 vdd.t186 vdd.n779 5.44203
R18661 vdd.n683 vdd.t17 5.44203
R18662 vdd.n1180 vdd.t118 5.10193
R18663 vdd.t190 vdd.n802 5.10193
R18664 vdd.n792 vdd.t193 5.10193
R18665 vdd.t0 vdd.n670 5.10193
R18666 vdd.n660 vdd.t10 5.10193
R18667 vdd.n3035 vdd.t107 5.10193
R18668 vdd.n275 vdd.n266 5.04292
R18669 vdd.n228 vdd.n219 5.04292
R18670 vdd.n185 vdd.n176 5.04292
R18671 vdd.n138 vdd.n129 5.04292
R18672 vdd.n96 vdd.n87 5.04292
R18673 vdd.n49 vdd.n40 5.04292
R18674 vdd.n1090 vdd.n1081 5.04292
R18675 vdd.n1137 vdd.n1128 5.04292
R18676 vdd.n1000 vdd.n991 5.04292
R18677 vdd.n1047 vdd.n1038 5.04292
R18678 vdd.n911 vdd.n902 5.04292
R18679 vdd.n958 vdd.n949 5.04292
R18680 vdd.n1473 vdd.t136 4.8752
R18681 vdd.t1 vdd.t8 4.8752
R18682 vdd.t4 vdd.t194 4.8752
R18683 vdd.t191 vdd.t181 4.8752
R18684 vdd.t188 vdd.t11 4.8752
R18685 vdd.t103 vdd.n304 4.8752
R18686 vdd.n2155 vdd.n2154 4.83952
R18687 vdd.n1767 vdd.n1763 4.83952
R18688 vdd.n2409 vdd.n2408 4.83952
R18689 vdd.n2615 vdd.n2614 4.83952
R18690 vdd.n591 vdd.n586 4.83952
R18691 vdd.n2315 vdd.n2258 4.83952
R18692 vdd.n2082 vdd.n757 4.83952
R18693 vdd.n1826 vdd.n1825 4.83952
R18694 vdd.n1621 vdd.n855 4.74817
R18695 vdd.n1616 vdd.n856 4.74817
R18696 vdd.n1518 vdd.n1515 4.74817
R18697 vdd.n1930 vdd.n1519 4.74817
R18698 vdd.n1932 vdd.n1518 4.74817
R18699 vdd.n1931 vdd.n1930 4.74817
R18700 vdd.n2838 vdd.n2837 4.74817
R18701 vdd.n2835 vdd.n2834 4.74817
R18702 vdd.n2835 vdd.n521 4.74817
R18703 vdd.n2837 vdd.n518 4.74817
R18704 vdd.n2720 vdd.n573 4.74817
R18705 vdd.n2716 vdd.n574 4.74817
R18706 vdd.n2719 vdd.n574 4.74817
R18707 vdd.n2723 vdd.n573 4.74817
R18708 vdd.n1617 vdd.n855 4.74817
R18709 vdd.n858 vdd.n856 4.74817
R18710 vdd.n297 vdd.n296 4.7074
R18711 vdd.n207 vdd.n206 4.7074
R18712 vdd.n1159 vdd.n1158 4.7074
R18713 vdd.n1069 vdd.n1068 4.7074
R18714 vdd.n1489 vdd.t97 4.64847
R18715 vdd.n2866 vdd.t99 4.64847
R18716 vdd.n2032 vdd.t2 4.53511
R18717 vdd.n2520 vdd.t184 4.53511
R18718 vdd.n2064 vdd.t182 4.30838
R18719 vdd.n2490 vdd.t179 4.30838
R18720 vdd.n276 vdd.n264 4.26717
R18721 vdd.n229 vdd.n217 4.26717
R18722 vdd.n186 vdd.n174 4.26717
R18723 vdd.n139 vdd.n127 4.26717
R18724 vdd.n97 vdd.n85 4.26717
R18725 vdd.n50 vdd.n38 4.26717
R18726 vdd.n1091 vdd.n1079 4.26717
R18727 vdd.n1138 vdd.n1126 4.26717
R18728 vdd.n1001 vdd.n989 4.26717
R18729 vdd.n1048 vdd.n1036 4.26717
R18730 vdd.n912 vdd.n900 4.26717
R18731 vdd.n959 vdd.n947 4.26717
R18732 vdd.n297 vdd.n207 4.10845
R18733 vdd.n1159 vdd.n1069 4.10845
R18734 vdd.n253 vdd.t144 4.06363
R18735 vdd.n253 vdd.t108 4.06363
R18736 vdd.n251 vdd.t110 4.06363
R18737 vdd.n251 vdd.t131 4.06363
R18738 vdd.n249 vdd.t133 4.06363
R18739 vdd.n249 vdd.t149 4.06363
R18740 vdd.n163 vdd.t139 4.06363
R18741 vdd.n163 vdd.t160 4.06363
R18742 vdd.n161 vdd.t104 4.06363
R18743 vdd.n161 vdd.t123 4.06363
R18744 vdd.n159 vdd.t129 4.06363
R18745 vdd.n159 vdd.t140 4.06363
R18746 vdd.n74 vdd.t145 4.06363
R18747 vdd.n74 vdd.t120 4.06363
R18748 vdd.n72 vdd.t159 4.06363
R18749 vdd.n72 vdd.t115 4.06363
R18750 vdd.n70 vdd.t152 4.06363
R18751 vdd.n70 vdd.t126 4.06363
R18752 vdd.n1111 vdd.t111 4.06363
R18753 vdd.n1111 vdd.t155 4.06363
R18754 vdd.n1113 vdd.t154 4.06363
R18755 vdd.n1113 vdd.t143 4.06363
R18756 vdd.n1115 vdd.t130 4.06363
R18757 vdd.n1115 vdd.t109 4.06363
R18758 vdd.n1021 vdd.t106 4.06363
R18759 vdd.n1021 vdd.t151 4.06363
R18760 vdd.n1023 vdd.t146 4.06363
R18761 vdd.n1023 vdd.t137 4.06363
R18762 vdd.n1025 vdd.t122 4.06363
R18763 vdd.n1025 vdd.t102 4.06363
R18764 vdd.n932 vdd.t124 4.06363
R18765 vdd.n932 vdd.t153 4.06363
R18766 vdd.n934 vdd.t113 4.06363
R18767 vdd.n934 vdd.t141 4.06363
R18768 vdd.n936 vdd.t119 4.06363
R18769 vdd.n936 vdd.t147 4.06363
R18770 vdd.n26 vdd.t162 3.9605
R18771 vdd.n26 vdd.t163 3.9605
R18772 vdd.n23 vdd.t175 3.9605
R18773 vdd.n23 vdd.t169 3.9605
R18774 vdd.n21 vdd.t173 3.9605
R18775 vdd.n21 vdd.t161 3.9605
R18776 vdd.n20 vdd.t166 3.9605
R18777 vdd.n20 vdd.t165 3.9605
R18778 vdd.n15 vdd.t168 3.9605
R18779 vdd.n15 vdd.t167 3.9605
R18780 vdd.n16 vdd.t170 3.9605
R18781 vdd.n16 vdd.t176 3.9605
R18782 vdd.n18 vdd.t174 3.9605
R18783 vdd.n18 vdd.t164 3.9605
R18784 vdd.n25 vdd.t172 3.9605
R18785 vdd.n25 vdd.t171 3.9605
R18786 vdd.n7 vdd.t189 3.61217
R18787 vdd.n7 vdd.t185 3.61217
R18788 vdd.n8 vdd.t192 3.61217
R18789 vdd.n8 vdd.t18 3.61217
R18790 vdd.n10 vdd.t197 3.61217
R18791 vdd.n10 vdd.t180 3.61217
R18792 vdd.n12 vdd.t6 3.61217
R18793 vdd.n12 vdd.t199 3.61217
R18794 vdd.n5 vdd.t16 3.61217
R18795 vdd.n5 vdd.t13 3.61217
R18796 vdd.n3 vdd.t183 3.61217
R18797 vdd.n3 vdd.t20 3.61217
R18798 vdd.n1 vdd.t187 3.61217
R18799 vdd.n1 vdd.t195 3.61217
R18800 vdd.n0 vdd.t3 3.61217
R18801 vdd.n0 vdd.t9 3.61217
R18802 vdd.n280 vdd.n279 3.49141
R18803 vdd.n233 vdd.n232 3.49141
R18804 vdd.n190 vdd.n189 3.49141
R18805 vdd.n143 vdd.n142 3.49141
R18806 vdd.n101 vdd.n100 3.49141
R18807 vdd.n54 vdd.n53 3.49141
R18808 vdd.n1095 vdd.n1094 3.49141
R18809 vdd.n1142 vdd.n1141 3.49141
R18810 vdd.n1005 vdd.n1004 3.49141
R18811 vdd.n1052 vdd.n1051 3.49141
R18812 vdd.n916 vdd.n915 3.49141
R18813 vdd.n963 vdd.n962 3.49141
R18814 vdd.n1770 vdd.t182 3.40145
R18815 vdd.n2218 vdd.t15 3.40145
R18816 vdd.n2471 vdd.t198 3.40145
R18817 vdd.n2395 vdd.t179 3.40145
R18818 vdd.n1871 vdd.t2 3.17472
R18819 vdd.n2374 vdd.t184 3.17472
R18820 vdd.n1490 vdd.t150 2.83463
R18821 vdd.n1508 vdd.t29 2.83463
R18822 vdd.n2849 vdd.t22 2.83463
R18823 vdd.n467 vdd.t128 2.83463
R18824 vdd.n283 vdd.n262 2.71565
R18825 vdd.n236 vdd.n215 2.71565
R18826 vdd.n193 vdd.n172 2.71565
R18827 vdd.n146 vdd.n125 2.71565
R18828 vdd.n104 vdd.n83 2.71565
R18829 vdd.n57 vdd.n36 2.71565
R18830 vdd.n1098 vdd.n1077 2.71565
R18831 vdd.n1145 vdd.n1124 2.71565
R18832 vdd.n1008 vdd.n987 2.71565
R18833 vdd.n1055 vdd.n1034 2.71565
R18834 vdd.n919 vdd.n898 2.71565
R18835 vdd.n966 vdd.n945 2.71565
R18836 vdd.t112 vdd.n1164 2.6079
R18837 vdd.n2020 vdd.t190 2.6079
R18838 vdd.n2044 vdd.t193 2.6079
R18839 vdd.n2508 vdd.t0 2.6079
R18840 vdd.n2532 vdd.t10 2.6079
R18841 vdd.n3043 vdd.t114 2.6079
R18842 vdd.n2538 vdd.n2537 2.49806
R18843 vdd.n2012 vdd.n2011 2.49806
R18844 vdd.n270 vdd.n269 2.4129
R18845 vdd.n223 vdd.n222 2.4129
R18846 vdd.n180 vdd.n179 2.4129
R18847 vdd.n133 vdd.n132 2.4129
R18848 vdd.n91 vdd.n90 2.4129
R18849 vdd.n44 vdd.n43 2.4129
R18850 vdd.n1085 vdd.n1084 2.4129
R18851 vdd.n1132 vdd.n1131 2.4129
R18852 vdd.n995 vdd.n994 2.4129
R18853 vdd.n1042 vdd.n1041 2.4129
R18854 vdd.n906 vdd.n905 2.4129
R18855 vdd.n953 vdd.n952 2.4129
R18856 vdd.n1447 vdd.t134 2.38117
R18857 vdd.n3034 vdd.t116 2.38117
R18858 vdd.n1929 vdd.n1518 2.27742
R18859 vdd.n1930 vdd.n1929 2.27742
R18860 vdd.n2836 vdd.n2835 2.27742
R18861 vdd.n2837 vdd.n2836 2.27742
R18862 vdd.n2707 vdd.n574 2.27742
R18863 vdd.n2707 vdd.n573 2.27742
R18864 vdd.n1952 vdd.n855 2.27742
R18865 vdd.n1952 vdd.n856 2.27742
R18866 vdd.n2044 vdd.t186 2.2678
R18867 vdd.n2508 vdd.t17 2.2678
R18868 vdd.t194 vdd.n773 2.04107
R18869 vdd.n690 vdd.t191 2.04107
R18870 vdd.n284 vdd.n260 1.93989
R18871 vdd.n237 vdd.n213 1.93989
R18872 vdd.n194 vdd.n170 1.93989
R18873 vdd.n147 vdd.n123 1.93989
R18874 vdd.n105 vdd.n81 1.93989
R18875 vdd.n58 vdd.n34 1.93989
R18876 vdd.n1099 vdd.n1075 1.93989
R18877 vdd.n1146 vdd.n1122 1.93989
R18878 vdd.n1009 vdd.n985 1.93989
R18879 vdd.n1056 vdd.n1032 1.93989
R18880 vdd.n920 vdd.n896 1.93989
R18881 vdd.n967 vdd.n943 1.93989
R18882 vdd.n1995 vdd.t69 1.92771
R18883 vdd.n2071 vdd.t54 1.92771
R18884 vdd.n2484 vdd.t62 1.92771
R18885 vdd.n2603 vdd.t58 1.92771
R18886 vdd.n1871 vdd.t177 1.70098
R18887 vdd.n798 vdd.t1 1.70098
R18888 vdd.t11 vdd.n664 1.70098
R18889 vdd.n2374 vdd.t14 1.70098
R18890 vdd.n1455 vdd.t101 1.24752
R18891 vdd.t138 vdd.n3041 1.24752
R18892 vdd.n295 vdd.n255 1.16414
R18893 vdd.n288 vdd.n287 1.16414
R18894 vdd.n248 vdd.n208 1.16414
R18895 vdd.n241 vdd.n240 1.16414
R18896 vdd.n205 vdd.n165 1.16414
R18897 vdd.n198 vdd.n197 1.16414
R18898 vdd.n158 vdd.n118 1.16414
R18899 vdd.n151 vdd.n150 1.16414
R18900 vdd.n116 vdd.n76 1.16414
R18901 vdd.n109 vdd.n108 1.16414
R18902 vdd.n69 vdd.n29 1.16414
R18903 vdd.n62 vdd.n61 1.16414
R18904 vdd.n1110 vdd.n1070 1.16414
R18905 vdd.n1103 vdd.n1102 1.16414
R18906 vdd.n1157 vdd.n1117 1.16414
R18907 vdd.n1150 vdd.n1149 1.16414
R18908 vdd.n1020 vdd.n980 1.16414
R18909 vdd.n1013 vdd.n1012 1.16414
R18910 vdd.n1067 vdd.n1027 1.16414
R18911 vdd.n1060 vdd.n1059 1.16414
R18912 vdd.n931 vdd.n891 1.16414
R18913 vdd.n924 vdd.n923 1.16414
R18914 vdd.n978 vdd.n938 1.16414
R18915 vdd.n971 vdd.n970 1.16414
R18916 vdd.n2038 vdd.t8 1.13415
R18917 vdd.n2514 vdd.t188 1.13415
R18918 vdd.n1481 vdd.t105 1.02079
R18919 vdd.t73 vdd.t178 1.02079
R18920 vdd.t7 vdd.t37 1.02079
R18921 vdd.t125 vdd.n456 1.02079
R18922 vdd.n1326 vdd.n1322 0.970197
R18923 vdd.n1950 vdd.n1949 0.970197
R18924 vdd.n2911 vdd.n2910 0.970197
R18925 vdd.n2715 vdd.n2713 0.970197
R18926 vdd.n2014 vdd.t178 0.794056
R18927 vdd.n2050 vdd.t4 0.794056
R18928 vdd.n2502 vdd.t181 0.794056
R18929 vdd.n2540 vdd.t7 0.794056
R18930 vdd.n1160 vdd.n28 0.74827
R18931 vdd vdd.n3048 0.740437
R18932 vdd.n1430 vdd.t33 0.567326
R18933 vdd.n3026 vdd.t44 0.567326
R18934 vdd.n1940 vdd.n1939 0.537085
R18935 vdd.n2845 vdd.n2844 0.537085
R18936 vdd.n3022 vdd.n3021 0.537085
R18937 vdd.n2904 vdd.n2903 0.537085
R18938 vdd.n2709 vdd.n476 0.537085
R18939 vdd.n1503 vdd.n857 0.537085
R18940 vdd.n1324 vdd.n1189 0.537085
R18941 vdd.n1426 vdd.n1425 0.537085
R18942 vdd.n4 vdd.n2 0.459552
R18943 vdd.n11 vdd.n9 0.459552
R18944 vdd.n293 vdd.n292 0.388379
R18945 vdd.n259 vdd.n257 0.388379
R18946 vdd.n246 vdd.n245 0.388379
R18947 vdd.n212 vdd.n210 0.388379
R18948 vdd.n203 vdd.n202 0.388379
R18949 vdd.n169 vdd.n167 0.388379
R18950 vdd.n156 vdd.n155 0.388379
R18951 vdd.n122 vdd.n120 0.388379
R18952 vdd.n114 vdd.n113 0.388379
R18953 vdd.n80 vdd.n78 0.388379
R18954 vdd.n67 vdd.n66 0.388379
R18955 vdd.n33 vdd.n31 0.388379
R18956 vdd.n1108 vdd.n1107 0.388379
R18957 vdd.n1074 vdd.n1072 0.388379
R18958 vdd.n1155 vdd.n1154 0.388379
R18959 vdd.n1121 vdd.n1119 0.388379
R18960 vdd.n1018 vdd.n1017 0.388379
R18961 vdd.n984 vdd.n982 0.388379
R18962 vdd.n1065 vdd.n1064 0.388379
R18963 vdd.n1031 vdd.n1029 0.388379
R18964 vdd.n929 vdd.n928 0.388379
R18965 vdd.n895 vdd.n893 0.388379
R18966 vdd.n976 vdd.n975 0.388379
R18967 vdd.n942 vdd.n940 0.388379
R18968 vdd.n19 vdd.n17 0.387128
R18969 vdd.n24 vdd.n22 0.387128
R18970 vdd.n6 vdd.n4 0.358259
R18971 vdd.n13 vdd.n11 0.358259
R18972 vdd.n252 vdd.n250 0.358259
R18973 vdd.n254 vdd.n252 0.358259
R18974 vdd.n296 vdd.n254 0.358259
R18975 vdd.n162 vdd.n160 0.358259
R18976 vdd.n164 vdd.n162 0.358259
R18977 vdd.n206 vdd.n164 0.358259
R18978 vdd.n73 vdd.n71 0.358259
R18979 vdd.n75 vdd.n73 0.358259
R18980 vdd.n117 vdd.n75 0.358259
R18981 vdd.n1158 vdd.n1116 0.358259
R18982 vdd.n1116 vdd.n1114 0.358259
R18983 vdd.n1114 vdd.n1112 0.358259
R18984 vdd.n1068 vdd.n1026 0.358259
R18985 vdd.n1026 vdd.n1024 0.358259
R18986 vdd.n1024 vdd.n1022 0.358259
R18987 vdd.n979 vdd.n937 0.358259
R18988 vdd.n937 vdd.n935 0.358259
R18989 vdd.n935 vdd.n933 0.358259
R18990 vdd.n14 vdd.n6 0.334552
R18991 vdd.n14 vdd.n13 0.334552
R18992 vdd.n27 vdd.n19 0.21707
R18993 vdd.n27 vdd.n24 0.21707
R18994 vdd.n294 vdd.n256 0.155672
R18995 vdd.n286 vdd.n256 0.155672
R18996 vdd.n286 vdd.n285 0.155672
R18997 vdd.n285 vdd.n261 0.155672
R18998 vdd.n278 vdd.n261 0.155672
R18999 vdd.n278 vdd.n277 0.155672
R19000 vdd.n277 vdd.n265 0.155672
R19001 vdd.n270 vdd.n265 0.155672
R19002 vdd.n247 vdd.n209 0.155672
R19003 vdd.n239 vdd.n209 0.155672
R19004 vdd.n239 vdd.n238 0.155672
R19005 vdd.n238 vdd.n214 0.155672
R19006 vdd.n231 vdd.n214 0.155672
R19007 vdd.n231 vdd.n230 0.155672
R19008 vdd.n230 vdd.n218 0.155672
R19009 vdd.n223 vdd.n218 0.155672
R19010 vdd.n204 vdd.n166 0.155672
R19011 vdd.n196 vdd.n166 0.155672
R19012 vdd.n196 vdd.n195 0.155672
R19013 vdd.n195 vdd.n171 0.155672
R19014 vdd.n188 vdd.n171 0.155672
R19015 vdd.n188 vdd.n187 0.155672
R19016 vdd.n187 vdd.n175 0.155672
R19017 vdd.n180 vdd.n175 0.155672
R19018 vdd.n157 vdd.n119 0.155672
R19019 vdd.n149 vdd.n119 0.155672
R19020 vdd.n149 vdd.n148 0.155672
R19021 vdd.n148 vdd.n124 0.155672
R19022 vdd.n141 vdd.n124 0.155672
R19023 vdd.n141 vdd.n140 0.155672
R19024 vdd.n140 vdd.n128 0.155672
R19025 vdd.n133 vdd.n128 0.155672
R19026 vdd.n115 vdd.n77 0.155672
R19027 vdd.n107 vdd.n77 0.155672
R19028 vdd.n107 vdd.n106 0.155672
R19029 vdd.n106 vdd.n82 0.155672
R19030 vdd.n99 vdd.n82 0.155672
R19031 vdd.n99 vdd.n98 0.155672
R19032 vdd.n98 vdd.n86 0.155672
R19033 vdd.n91 vdd.n86 0.155672
R19034 vdd.n68 vdd.n30 0.155672
R19035 vdd.n60 vdd.n30 0.155672
R19036 vdd.n60 vdd.n59 0.155672
R19037 vdd.n59 vdd.n35 0.155672
R19038 vdd.n52 vdd.n35 0.155672
R19039 vdd.n52 vdd.n51 0.155672
R19040 vdd.n51 vdd.n39 0.155672
R19041 vdd.n44 vdd.n39 0.155672
R19042 vdd.n1109 vdd.n1071 0.155672
R19043 vdd.n1101 vdd.n1071 0.155672
R19044 vdd.n1101 vdd.n1100 0.155672
R19045 vdd.n1100 vdd.n1076 0.155672
R19046 vdd.n1093 vdd.n1076 0.155672
R19047 vdd.n1093 vdd.n1092 0.155672
R19048 vdd.n1092 vdd.n1080 0.155672
R19049 vdd.n1085 vdd.n1080 0.155672
R19050 vdd.n1156 vdd.n1118 0.155672
R19051 vdd.n1148 vdd.n1118 0.155672
R19052 vdd.n1148 vdd.n1147 0.155672
R19053 vdd.n1147 vdd.n1123 0.155672
R19054 vdd.n1140 vdd.n1123 0.155672
R19055 vdd.n1140 vdd.n1139 0.155672
R19056 vdd.n1139 vdd.n1127 0.155672
R19057 vdd.n1132 vdd.n1127 0.155672
R19058 vdd.n1019 vdd.n981 0.155672
R19059 vdd.n1011 vdd.n981 0.155672
R19060 vdd.n1011 vdd.n1010 0.155672
R19061 vdd.n1010 vdd.n986 0.155672
R19062 vdd.n1003 vdd.n986 0.155672
R19063 vdd.n1003 vdd.n1002 0.155672
R19064 vdd.n1002 vdd.n990 0.155672
R19065 vdd.n995 vdd.n990 0.155672
R19066 vdd.n1066 vdd.n1028 0.155672
R19067 vdd.n1058 vdd.n1028 0.155672
R19068 vdd.n1058 vdd.n1057 0.155672
R19069 vdd.n1057 vdd.n1033 0.155672
R19070 vdd.n1050 vdd.n1033 0.155672
R19071 vdd.n1050 vdd.n1049 0.155672
R19072 vdd.n1049 vdd.n1037 0.155672
R19073 vdd.n1042 vdd.n1037 0.155672
R19074 vdd.n930 vdd.n892 0.155672
R19075 vdd.n922 vdd.n892 0.155672
R19076 vdd.n922 vdd.n921 0.155672
R19077 vdd.n921 vdd.n897 0.155672
R19078 vdd.n914 vdd.n897 0.155672
R19079 vdd.n914 vdd.n913 0.155672
R19080 vdd.n913 vdd.n901 0.155672
R19081 vdd.n906 vdd.n901 0.155672
R19082 vdd.n977 vdd.n939 0.155672
R19083 vdd.n969 vdd.n939 0.155672
R19084 vdd.n969 vdd.n968 0.155672
R19085 vdd.n968 vdd.n944 0.155672
R19086 vdd.n961 vdd.n944 0.155672
R19087 vdd.n961 vdd.n960 0.155672
R19088 vdd.n960 vdd.n948 0.155672
R19089 vdd.n953 vdd.n948 0.155672
R19090 vdd.n1715 vdd.n1520 0.152939
R19091 vdd.n1526 vdd.n1520 0.152939
R19092 vdd.n1527 vdd.n1526 0.152939
R19093 vdd.n1528 vdd.n1527 0.152939
R19094 vdd.n1529 vdd.n1528 0.152939
R19095 vdd.n1533 vdd.n1529 0.152939
R19096 vdd.n1534 vdd.n1533 0.152939
R19097 vdd.n1535 vdd.n1534 0.152939
R19098 vdd.n1536 vdd.n1535 0.152939
R19099 vdd.n1540 vdd.n1536 0.152939
R19100 vdd.n1541 vdd.n1540 0.152939
R19101 vdd.n1542 vdd.n1541 0.152939
R19102 vdd.n1690 vdd.n1542 0.152939
R19103 vdd.n1690 vdd.n1689 0.152939
R19104 vdd.n1689 vdd.n1688 0.152939
R19105 vdd.n1688 vdd.n1548 0.152939
R19106 vdd.n1553 vdd.n1548 0.152939
R19107 vdd.n1554 vdd.n1553 0.152939
R19108 vdd.n1555 vdd.n1554 0.152939
R19109 vdd.n1559 vdd.n1555 0.152939
R19110 vdd.n1560 vdd.n1559 0.152939
R19111 vdd.n1561 vdd.n1560 0.152939
R19112 vdd.n1562 vdd.n1561 0.152939
R19113 vdd.n1566 vdd.n1562 0.152939
R19114 vdd.n1567 vdd.n1566 0.152939
R19115 vdd.n1568 vdd.n1567 0.152939
R19116 vdd.n1569 vdd.n1568 0.152939
R19117 vdd.n1573 vdd.n1569 0.152939
R19118 vdd.n1574 vdd.n1573 0.152939
R19119 vdd.n1575 vdd.n1574 0.152939
R19120 vdd.n1576 vdd.n1575 0.152939
R19121 vdd.n1580 vdd.n1576 0.152939
R19122 vdd.n1581 vdd.n1580 0.152939
R19123 vdd.n1582 vdd.n1581 0.152939
R19124 vdd.n1651 vdd.n1582 0.152939
R19125 vdd.n1651 vdd.n1650 0.152939
R19126 vdd.n1650 vdd.n1649 0.152939
R19127 vdd.n1649 vdd.n1588 0.152939
R19128 vdd.n1593 vdd.n1588 0.152939
R19129 vdd.n1594 vdd.n1593 0.152939
R19130 vdd.n1595 vdd.n1594 0.152939
R19131 vdd.n1599 vdd.n1595 0.152939
R19132 vdd.n1600 vdd.n1599 0.152939
R19133 vdd.n1601 vdd.n1600 0.152939
R19134 vdd.n1602 vdd.n1601 0.152939
R19135 vdd.n1606 vdd.n1602 0.152939
R19136 vdd.n1607 vdd.n1606 0.152939
R19137 vdd.n1608 vdd.n1607 0.152939
R19138 vdd.n1609 vdd.n1608 0.152939
R19139 vdd.n1610 vdd.n1609 0.152939
R19140 vdd.n1610 vdd.n854 0.152939
R19141 vdd.n1939 vdd.n1514 0.152939
R19142 vdd.n1477 vdd.n1476 0.152939
R19143 vdd.n1478 vdd.n1477 0.152939
R19144 vdd.n1478 vdd.n879 0.152939
R19145 vdd.n1493 vdd.n879 0.152939
R19146 vdd.n1494 vdd.n1493 0.152939
R19147 vdd.n1495 vdd.n1494 0.152939
R19148 vdd.n1495 vdd.n867 0.152939
R19149 vdd.n1512 vdd.n867 0.152939
R19150 vdd.n1513 vdd.n1512 0.152939
R19151 vdd.n1940 vdd.n1513 0.152939
R19152 vdd.n524 vdd.n519 0.152939
R19153 vdd.n525 vdd.n524 0.152939
R19154 vdd.n526 vdd.n525 0.152939
R19155 vdd.n527 vdd.n526 0.152939
R19156 vdd.n528 vdd.n527 0.152939
R19157 vdd.n529 vdd.n528 0.152939
R19158 vdd.n530 vdd.n529 0.152939
R19159 vdd.n531 vdd.n530 0.152939
R19160 vdd.n532 vdd.n531 0.152939
R19161 vdd.n533 vdd.n532 0.152939
R19162 vdd.n534 vdd.n533 0.152939
R19163 vdd.n535 vdd.n534 0.152939
R19164 vdd.n2803 vdd.n535 0.152939
R19165 vdd.n2803 vdd.n2802 0.152939
R19166 vdd.n2802 vdd.n2801 0.152939
R19167 vdd.n2801 vdd.n537 0.152939
R19168 vdd.n538 vdd.n537 0.152939
R19169 vdd.n539 vdd.n538 0.152939
R19170 vdd.n540 vdd.n539 0.152939
R19171 vdd.n541 vdd.n540 0.152939
R19172 vdd.n542 vdd.n541 0.152939
R19173 vdd.n543 vdd.n542 0.152939
R19174 vdd.n544 vdd.n543 0.152939
R19175 vdd.n545 vdd.n544 0.152939
R19176 vdd.n546 vdd.n545 0.152939
R19177 vdd.n547 vdd.n546 0.152939
R19178 vdd.n548 vdd.n547 0.152939
R19179 vdd.n549 vdd.n548 0.152939
R19180 vdd.n550 vdd.n549 0.152939
R19181 vdd.n551 vdd.n550 0.152939
R19182 vdd.n552 vdd.n551 0.152939
R19183 vdd.n553 vdd.n552 0.152939
R19184 vdd.n554 vdd.n553 0.152939
R19185 vdd.n555 vdd.n554 0.152939
R19186 vdd.n2757 vdd.n555 0.152939
R19187 vdd.n2757 vdd.n2756 0.152939
R19188 vdd.n2756 vdd.n2755 0.152939
R19189 vdd.n2755 vdd.n559 0.152939
R19190 vdd.n560 vdd.n559 0.152939
R19191 vdd.n561 vdd.n560 0.152939
R19192 vdd.n562 vdd.n561 0.152939
R19193 vdd.n563 vdd.n562 0.152939
R19194 vdd.n564 vdd.n563 0.152939
R19195 vdd.n565 vdd.n564 0.152939
R19196 vdd.n566 vdd.n565 0.152939
R19197 vdd.n567 vdd.n566 0.152939
R19198 vdd.n568 vdd.n567 0.152939
R19199 vdd.n569 vdd.n568 0.152939
R19200 vdd.n570 vdd.n569 0.152939
R19201 vdd.n571 vdd.n570 0.152939
R19202 vdd.n572 vdd.n571 0.152939
R19203 vdd.n2844 vdd.n481 0.152939
R19204 vdd.n2846 vdd.n2845 0.152939
R19205 vdd.n2846 vdd.n470 0.152939
R19206 vdd.n2861 vdd.n470 0.152939
R19207 vdd.n2862 vdd.n2861 0.152939
R19208 vdd.n2863 vdd.n2862 0.152939
R19209 vdd.n2863 vdd.n459 0.152939
R19210 vdd.n2877 vdd.n459 0.152939
R19211 vdd.n2878 vdd.n2877 0.152939
R19212 vdd.n2879 vdd.n2878 0.152939
R19213 vdd.n2879 vdd.n298 0.152939
R19214 vdd.n3046 vdd.n299 0.152939
R19215 vdd.n310 vdd.n299 0.152939
R19216 vdd.n311 vdd.n310 0.152939
R19217 vdd.n312 vdd.n311 0.152939
R19218 vdd.n320 vdd.n312 0.152939
R19219 vdd.n321 vdd.n320 0.152939
R19220 vdd.n322 vdd.n321 0.152939
R19221 vdd.n323 vdd.n322 0.152939
R19222 vdd.n331 vdd.n323 0.152939
R19223 vdd.n3022 vdd.n331 0.152939
R19224 vdd.n3021 vdd.n332 0.152939
R19225 vdd.n335 vdd.n332 0.152939
R19226 vdd.n339 vdd.n335 0.152939
R19227 vdd.n340 vdd.n339 0.152939
R19228 vdd.n341 vdd.n340 0.152939
R19229 vdd.n342 vdd.n341 0.152939
R19230 vdd.n343 vdd.n342 0.152939
R19231 vdd.n347 vdd.n343 0.152939
R19232 vdd.n348 vdd.n347 0.152939
R19233 vdd.n349 vdd.n348 0.152939
R19234 vdd.n350 vdd.n349 0.152939
R19235 vdd.n354 vdd.n350 0.152939
R19236 vdd.n355 vdd.n354 0.152939
R19237 vdd.n356 vdd.n355 0.152939
R19238 vdd.n357 vdd.n356 0.152939
R19239 vdd.n361 vdd.n357 0.152939
R19240 vdd.n362 vdd.n361 0.152939
R19241 vdd.n363 vdd.n362 0.152939
R19242 vdd.n2987 vdd.n363 0.152939
R19243 vdd.n2987 vdd.n2986 0.152939
R19244 vdd.n2986 vdd.n2985 0.152939
R19245 vdd.n2985 vdd.n369 0.152939
R19246 vdd.n374 vdd.n369 0.152939
R19247 vdd.n375 vdd.n374 0.152939
R19248 vdd.n376 vdd.n375 0.152939
R19249 vdd.n380 vdd.n376 0.152939
R19250 vdd.n381 vdd.n380 0.152939
R19251 vdd.n382 vdd.n381 0.152939
R19252 vdd.n383 vdd.n382 0.152939
R19253 vdd.n387 vdd.n383 0.152939
R19254 vdd.n388 vdd.n387 0.152939
R19255 vdd.n389 vdd.n388 0.152939
R19256 vdd.n390 vdd.n389 0.152939
R19257 vdd.n394 vdd.n390 0.152939
R19258 vdd.n395 vdd.n394 0.152939
R19259 vdd.n396 vdd.n395 0.152939
R19260 vdd.n397 vdd.n396 0.152939
R19261 vdd.n401 vdd.n397 0.152939
R19262 vdd.n402 vdd.n401 0.152939
R19263 vdd.n403 vdd.n402 0.152939
R19264 vdd.n2948 vdd.n403 0.152939
R19265 vdd.n2948 vdd.n2947 0.152939
R19266 vdd.n2947 vdd.n2946 0.152939
R19267 vdd.n2946 vdd.n409 0.152939
R19268 vdd.n414 vdd.n409 0.152939
R19269 vdd.n415 vdd.n414 0.152939
R19270 vdd.n416 vdd.n415 0.152939
R19271 vdd.n420 vdd.n416 0.152939
R19272 vdd.n421 vdd.n420 0.152939
R19273 vdd.n422 vdd.n421 0.152939
R19274 vdd.n423 vdd.n422 0.152939
R19275 vdd.n427 vdd.n423 0.152939
R19276 vdd.n428 vdd.n427 0.152939
R19277 vdd.n429 vdd.n428 0.152939
R19278 vdd.n430 vdd.n429 0.152939
R19279 vdd.n434 vdd.n430 0.152939
R19280 vdd.n435 vdd.n434 0.152939
R19281 vdd.n436 vdd.n435 0.152939
R19282 vdd.n437 vdd.n436 0.152939
R19283 vdd.n441 vdd.n437 0.152939
R19284 vdd.n442 vdd.n441 0.152939
R19285 vdd.n443 vdd.n442 0.152939
R19286 vdd.n2904 vdd.n443 0.152939
R19287 vdd.n2852 vdd.n476 0.152939
R19288 vdd.n2853 vdd.n2852 0.152939
R19289 vdd.n2854 vdd.n2853 0.152939
R19290 vdd.n2854 vdd.n464 0.152939
R19291 vdd.n2869 vdd.n464 0.152939
R19292 vdd.n2870 vdd.n2869 0.152939
R19293 vdd.n2871 vdd.n2870 0.152939
R19294 vdd.n2871 vdd.n452 0.152939
R19295 vdd.n2885 vdd.n452 0.152939
R19296 vdd.n2886 vdd.n2885 0.152939
R19297 vdd.n2887 vdd.n2886 0.152939
R19298 vdd.n2887 vdd.n450 0.152939
R19299 vdd.n2891 vdd.n450 0.152939
R19300 vdd.n2892 vdd.n2891 0.152939
R19301 vdd.n2893 vdd.n2892 0.152939
R19302 vdd.n2893 vdd.n447 0.152939
R19303 vdd.n2897 vdd.n447 0.152939
R19304 vdd.n2898 vdd.n2897 0.152939
R19305 vdd.n2899 vdd.n2898 0.152939
R19306 vdd.n2899 vdd.n444 0.152939
R19307 vdd.n2903 vdd.n444 0.152939
R19308 vdd.n2709 vdd.n2708 0.152939
R19309 vdd.n1951 vdd.n857 0.152939
R19310 vdd.n1433 vdd.n1189 0.152939
R19311 vdd.n1434 vdd.n1433 0.152939
R19312 vdd.n1435 vdd.n1434 0.152939
R19313 vdd.n1435 vdd.n1177 0.152939
R19314 vdd.n1450 vdd.n1177 0.152939
R19315 vdd.n1451 vdd.n1450 0.152939
R19316 vdd.n1452 vdd.n1451 0.152939
R19317 vdd.n1452 vdd.n1167 0.152939
R19318 vdd.n1468 vdd.n1167 0.152939
R19319 vdd.n1469 vdd.n1468 0.152939
R19320 vdd.n1470 vdd.n1469 0.152939
R19321 vdd.n1470 vdd.n884 0.152939
R19322 vdd.n1484 vdd.n884 0.152939
R19323 vdd.n1485 vdd.n1484 0.152939
R19324 vdd.n1486 vdd.n1485 0.152939
R19325 vdd.n1486 vdd.n874 0.152939
R19326 vdd.n1501 vdd.n874 0.152939
R19327 vdd.n1502 vdd.n1501 0.152939
R19328 vdd.n1505 vdd.n1502 0.152939
R19329 vdd.n1505 vdd.n1504 0.152939
R19330 vdd.n1504 vdd.n1503 0.152939
R19331 vdd.n1425 vdd.n1194 0.152939
R19332 vdd.n1418 vdd.n1194 0.152939
R19333 vdd.n1418 vdd.n1417 0.152939
R19334 vdd.n1417 vdd.n1416 0.152939
R19335 vdd.n1416 vdd.n1231 0.152939
R19336 vdd.n1412 vdd.n1231 0.152939
R19337 vdd.n1412 vdd.n1411 0.152939
R19338 vdd.n1411 vdd.n1410 0.152939
R19339 vdd.n1410 vdd.n1237 0.152939
R19340 vdd.n1406 vdd.n1237 0.152939
R19341 vdd.n1406 vdd.n1405 0.152939
R19342 vdd.n1405 vdd.n1404 0.152939
R19343 vdd.n1404 vdd.n1243 0.152939
R19344 vdd.n1400 vdd.n1243 0.152939
R19345 vdd.n1400 vdd.n1399 0.152939
R19346 vdd.n1399 vdd.n1398 0.152939
R19347 vdd.n1398 vdd.n1249 0.152939
R19348 vdd.n1394 vdd.n1249 0.152939
R19349 vdd.n1394 vdd.n1393 0.152939
R19350 vdd.n1393 vdd.n1392 0.152939
R19351 vdd.n1392 vdd.n1257 0.152939
R19352 vdd.n1388 vdd.n1257 0.152939
R19353 vdd.n1388 vdd.n1387 0.152939
R19354 vdd.n1387 vdd.n1386 0.152939
R19355 vdd.n1386 vdd.n1263 0.152939
R19356 vdd.n1382 vdd.n1263 0.152939
R19357 vdd.n1382 vdd.n1381 0.152939
R19358 vdd.n1381 vdd.n1380 0.152939
R19359 vdd.n1380 vdd.n1269 0.152939
R19360 vdd.n1376 vdd.n1269 0.152939
R19361 vdd.n1376 vdd.n1375 0.152939
R19362 vdd.n1375 vdd.n1374 0.152939
R19363 vdd.n1374 vdd.n1275 0.152939
R19364 vdd.n1370 vdd.n1275 0.152939
R19365 vdd.n1370 vdd.n1369 0.152939
R19366 vdd.n1369 vdd.n1368 0.152939
R19367 vdd.n1368 vdd.n1281 0.152939
R19368 vdd.n1364 vdd.n1281 0.152939
R19369 vdd.n1364 vdd.n1363 0.152939
R19370 vdd.n1363 vdd.n1362 0.152939
R19371 vdd.n1362 vdd.n1287 0.152939
R19372 vdd.n1355 vdd.n1287 0.152939
R19373 vdd.n1355 vdd.n1354 0.152939
R19374 vdd.n1354 vdd.n1353 0.152939
R19375 vdd.n1353 vdd.n1292 0.152939
R19376 vdd.n1349 vdd.n1292 0.152939
R19377 vdd.n1349 vdd.n1348 0.152939
R19378 vdd.n1348 vdd.n1347 0.152939
R19379 vdd.n1347 vdd.n1298 0.152939
R19380 vdd.n1343 vdd.n1298 0.152939
R19381 vdd.n1343 vdd.n1342 0.152939
R19382 vdd.n1342 vdd.n1341 0.152939
R19383 vdd.n1341 vdd.n1304 0.152939
R19384 vdd.n1337 vdd.n1304 0.152939
R19385 vdd.n1337 vdd.n1336 0.152939
R19386 vdd.n1336 vdd.n1335 0.152939
R19387 vdd.n1335 vdd.n1310 0.152939
R19388 vdd.n1331 vdd.n1310 0.152939
R19389 vdd.n1331 vdd.n1330 0.152939
R19390 vdd.n1330 vdd.n1329 0.152939
R19391 vdd.n1329 vdd.n1316 0.152939
R19392 vdd.n1325 vdd.n1316 0.152939
R19393 vdd.n1325 vdd.n1324 0.152939
R19394 vdd.n1427 vdd.n1426 0.152939
R19395 vdd.n1427 vdd.n1183 0.152939
R19396 vdd.n1442 vdd.n1183 0.152939
R19397 vdd.n1443 vdd.n1442 0.152939
R19398 vdd.n1444 vdd.n1443 0.152939
R19399 vdd.n1444 vdd.n1172 0.152939
R19400 vdd.n1459 vdd.n1172 0.152939
R19401 vdd.n1460 vdd.n1459 0.152939
R19402 vdd.n1462 vdd.n1460 0.152939
R19403 vdd.n1462 vdd.n1461 0.152939
R19404 vdd.n1929 vdd.n1514 0.110256
R19405 vdd.n2836 vdd.n481 0.110256
R19406 vdd.n2708 vdd.n2707 0.110256
R19407 vdd.n1952 vdd.n1951 0.110256
R19408 vdd.n1476 vdd.n1161 0.0695946
R19409 vdd.n3047 vdd.n298 0.0695946
R19410 vdd.n3047 vdd.n3046 0.0695946
R19411 vdd.n1461 vdd.n1161 0.0695946
R19412 vdd.n1929 vdd.n1715 0.0431829
R19413 vdd.n1952 vdd.n854 0.0431829
R19414 vdd.n2836 vdd.n519 0.0431829
R19415 vdd.n2707 vdd.n572 0.0431829
R19416 vdd vdd.n28 0.00833333
R19417 a_n2848_n452.n5 a_n2848_n452.t75 539.01
R19418 a_n2848_n452.n97 a_n2848_n452.t58 512.366
R19419 a_n2848_n452.n96 a_n2848_n452.t62 512.366
R19420 a_n2848_n452.n70 a_n2848_n452.t52 512.366
R19421 a_n2848_n452.n95 a_n2848_n452.t67 512.366
R19422 a_n2848_n452.n1 a_n2848_n452.t32 533.058
R19423 a_n2848_n452.n101 a_n2848_n452.t38 512.366
R19424 a_n2848_n452.n100 a_n2848_n452.t20 512.366
R19425 a_n2848_n452.n69 a_n2848_n452.t18 512.366
R19426 a_n2848_n452.n98 a_n2848_n452.t30 512.366
R19427 a_n2848_n452.n19 a_n2848_n452.t22 539.01
R19428 a_n2848_n452.n78 a_n2848_n452.t28 512.366
R19429 a_n2848_n452.n79 a_n2848_n452.t40 512.366
R19430 a_n2848_n452.n73 a_n2848_n452.t24 512.366
R19431 a_n2848_n452.n80 a_n2848_n452.t34 512.366
R19432 a_n2848_n452.n23 a_n2848_n452.t70 539.01
R19433 a_n2848_n452.n75 a_n2848_n452.t71 512.366
R19434 a_n2848_n452.n76 a_n2848_n452.t50 512.366
R19435 a_n2848_n452.n74 a_n2848_n452.t56 512.366
R19436 a_n2848_n452.n77 a_n2848_n452.t65 512.366
R19437 a_n2848_n452.n92 a_n2848_n452.t64 512.366
R19438 a_n2848_n452.n82 a_n2848_n452.t55 512.366
R19439 a_n2848_n452.n93 a_n2848_n452.t49 512.366
R19440 a_n2848_n452.n90 a_n2848_n452.t72 512.366
R19441 a_n2848_n452.n83 a_n2848_n452.t61 512.366
R19442 a_n2848_n452.n91 a_n2848_n452.t60 512.366
R19443 a_n2848_n452.n88 a_n2848_n452.t68 512.366
R19444 a_n2848_n452.n84 a_n2848_n452.t53 512.366
R19445 a_n2848_n452.n89 a_n2848_n452.t54 512.366
R19446 a_n2848_n452.n86 a_n2848_n452.t57 512.366
R19447 a_n2848_n452.n85 a_n2848_n452.t66 512.366
R19448 a_n2848_n452.n87 a_n2848_n452.t48 512.366
R19449 a_n2848_n452.n50 a_n2848_n452.n3 70.3058
R19450 a_n2848_n452.n47 a_n2848_n452.n6 70.3058
R19451 a_n2848_n452.n16 a_n2848_n452.n37 70.3058
R19452 a_n2848_n452.n20 a_n2848_n452.n34 70.3058
R19453 a_n2848_n452.n33 a_n2848_n452.n21 70.1674
R19454 a_n2848_n452.n33 a_n2848_n452.n74 20.9683
R19455 a_n2848_n452.n21 a_n2848_n452.n32 75.0448
R19456 a_n2848_n452.n76 a_n2848_n452.n32 11.2134
R19457 a_n2848_n452.n22 a_n2848_n452.n23 44.8194
R19458 a_n2848_n452.n36 a_n2848_n452.n17 70.1674
R19459 a_n2848_n452.n36 a_n2848_n452.n73 20.9683
R19460 a_n2848_n452.n17 a_n2848_n452.n35 75.0448
R19461 a_n2848_n452.n79 a_n2848_n452.n35 11.2134
R19462 a_n2848_n452.n18 a_n2848_n452.n19 44.8194
R19463 a_n2848_n452.n7 a_n2848_n452.n45 70.1674
R19464 a_n2848_n452.n9 a_n2848_n452.n43 70.1674
R19465 a_n2848_n452.n11 a_n2848_n452.n41 70.1674
R19466 a_n2848_n452.n14 a_n2848_n452.n39 70.1674
R19467 a_n2848_n452.n87 a_n2848_n452.n39 20.9683
R19468 a_n2848_n452.n38 a_n2848_n452.n15 75.0448
R19469 a_n2848_n452.n38 a_n2848_n452.n85 11.2134
R19470 a_n2848_n452.n15 a_n2848_n452.n86 161.3
R19471 a_n2848_n452.n89 a_n2848_n452.n41 20.9683
R19472 a_n2848_n452.n40 a_n2848_n452.n12 75.0448
R19473 a_n2848_n452.n40 a_n2848_n452.n84 11.2134
R19474 a_n2848_n452.n12 a_n2848_n452.n88 161.3
R19475 a_n2848_n452.n91 a_n2848_n452.n43 20.9683
R19476 a_n2848_n452.n42 a_n2848_n452.n10 75.0448
R19477 a_n2848_n452.n42 a_n2848_n452.n83 11.2134
R19478 a_n2848_n452.n10 a_n2848_n452.n90 161.3
R19479 a_n2848_n452.n93 a_n2848_n452.n45 20.9683
R19480 a_n2848_n452.n44 a_n2848_n452.n8 75.0448
R19481 a_n2848_n452.n44 a_n2848_n452.n82 11.2134
R19482 a_n2848_n452.n8 a_n2848_n452.n92 161.3
R19483 a_n2848_n452.n6 a_n2848_n452.n46 70.1674
R19484 a_n2848_n452.n46 a_n2848_n452.n69 20.9683
R19485 a_n2848_n452.n99 a_n2848_n452.n0 161.3
R19486 a_n2848_n452.n4 a_n2848_n452.n49 70.1674
R19487 a_n2848_n452.n49 a_n2848_n452.n70 20.9683
R19488 a_n2848_n452.n48 a_n2848_n452.n4 75.0448
R19489 a_n2848_n452.n96 a_n2848_n452.n48 11.2134
R19490 a_n2848_n452.n2 a_n2848_n452.n5 44.8194
R19491 a_n2848_n452.n100 a_n2848_n452.n51 20.9683
R19492 a_n2848_n452.n51 a_n2848_n452.n0 70.1674
R19493 a_n2848_n452.n0 a_n2848_n452.n1 70.3058
R19494 a_n2848_n452.n67 a_n2848_n452.n65 81.4626
R19495 a_n2848_n452.n58 a_n2848_n452.n56 81.4626
R19496 a_n2848_n452.n54 a_n2848_n452.n52 81.4626
R19497 a_n2848_n452.n67 a_n2848_n452.n66 80.9324
R19498 a_n2848_n452.n31 a_n2848_n452.n68 80.9324
R19499 a_n2848_n452.n30 a_n2848_n452.n64 80.9324
R19500 a_n2848_n452.n63 a_n2848_n452.n62 80.9324
R19501 a_n2848_n452.n61 a_n2848_n452.n60 80.9324
R19502 a_n2848_n452.n58 a_n2848_n452.n57 80.9324
R19503 a_n2848_n452.n29 a_n2848_n452.n59 80.9324
R19504 a_n2848_n452.n28 a_n2848_n452.n55 80.9324
R19505 a_n2848_n452.n54 a_n2848_n452.n53 80.9324
R19506 a_n2848_n452.n27 a_n2848_n452.t27 74.6477
R19507 a_n2848_n452.n24 a_n2848_n452.t23 74.6477
R19508 a_n2848_n452.n26 a_n2848_n452.t33 74.2899
R19509 a_n2848_n452.n25 a_n2848_n452.t37 74.2897
R19510 a_n2848_n452.n27 a_n2848_n452.n103 70.6783
R19511 a_n2848_n452.n25 a_n2848_n452.n72 70.6783
R19512 a_n2848_n452.n24 a_n2848_n452.n71 70.6783
R19513 a_n2848_n452.n104 a_n2848_n452.n27 70.6782
R19514 a_n2848_n452.n97 a_n2848_n452.n96 48.2005
R19515 a_n2848_n452.n95 a_n2848_n452.n49 20.9683
R19516 a_n2848_n452.n101 a_n2848_n452.n51 20.9683
R19517 a_n2848_n452.n98 a_n2848_n452.n46 20.9683
R19518 a_n2848_n452.n79 a_n2848_n452.n78 48.2005
R19519 a_n2848_n452.n80 a_n2848_n452.n36 20.9683
R19520 a_n2848_n452.n76 a_n2848_n452.n75 48.2005
R19521 a_n2848_n452.n77 a_n2848_n452.n33 20.9683
R19522 a_n2848_n452.n92 a_n2848_n452.n82 48.2005
R19523 a_n2848_n452.t69 a_n2848_n452.n45 533.335
R19524 a_n2848_n452.n90 a_n2848_n452.n83 48.2005
R19525 a_n2848_n452.t74 a_n2848_n452.n43 533.335
R19526 a_n2848_n452.n88 a_n2848_n452.n84 48.2005
R19527 a_n2848_n452.t63 a_n2848_n452.n41 533.335
R19528 a_n2848_n452.n86 a_n2848_n452.n85 48.2005
R19529 a_n2848_n452.t59 a_n2848_n452.n39 533.335
R19530 a_n2848_n452.n50 a_n2848_n452.t73 533.058
R19531 a_n2848_n452.n47 a_n2848_n452.t26 533.058
R19532 a_n2848_n452.t36 a_n2848_n452.n37 533.058
R19533 a_n2848_n452.t51 a_n2848_n452.n34 533.058
R19534 a_n2848_n452.n61 a_n2848_n452.n29 33.585
R19535 a_n2848_n452.n48 a_n2848_n452.n70 35.3134
R19536 a_n2848_n452.n100 a_n2848_n452.n99 24.1005
R19537 a_n2848_n452.n99 a_n2848_n452.n69 24.1005
R19538 a_n2848_n452.n73 a_n2848_n452.n35 35.3134
R19539 a_n2848_n452.n74 a_n2848_n452.n32 35.3134
R19540 a_n2848_n452.n93 a_n2848_n452.n44 35.3134
R19541 a_n2848_n452.n91 a_n2848_n452.n42 35.3134
R19542 a_n2848_n452.n89 a_n2848_n452.n40 35.3134
R19543 a_n2848_n452.n87 a_n2848_n452.n38 35.3134
R19544 a_n2848_n452.n0 a_n2848_n452.n31 23.891
R19545 a_n2848_n452.n22 a_n2848_n452.n13 12.046
R19546 a_n2848_n452.n3 a_n2848_n452.n94 11.8414
R19547 a_n2848_n452.n102 a_n2848_n452.n0 10.5365
R19548 a_n2848_n452.n81 a_n2848_n452.n25 9.50122
R19549 a_n2848_n452.n15 a_n2848_n452.n13 7.47588
R19550 a_n2848_n452.n94 a_n2848_n452.n7 7.47588
R19551 a_n2848_n452.n81 a_n2848_n452.n16 6.70126
R19552 a_n2848_n452.n26 a_n2848_n452.n102 5.65783
R19553 a_n2848_n452.n94 a_n2848_n452.n81 5.3452
R19554 a_n2848_n452.n18 a_n2848_n452.n20 3.95126
R19555 a_n2848_n452.n6 a_n2848_n452.n2 3.95126
R19556 a_n2848_n452.n103 a_n2848_n452.t39 3.61217
R19557 a_n2848_n452.n103 a_n2848_n452.t21 3.61217
R19558 a_n2848_n452.n72 a_n2848_n452.t25 3.61217
R19559 a_n2848_n452.n72 a_n2848_n452.t35 3.61217
R19560 a_n2848_n452.n71 a_n2848_n452.t29 3.61217
R19561 a_n2848_n452.n71 a_n2848_n452.t41 3.61217
R19562 a_n2848_n452.t19 a_n2848_n452.n104 3.61217
R19563 a_n2848_n452.n104 a_n2848_n452.t31 3.61217
R19564 a_n2848_n452.n65 a_n2848_n452.t5 2.82907
R19565 a_n2848_n452.n65 a_n2848_n452.t45 2.82907
R19566 a_n2848_n452.n66 a_n2848_n452.t14 2.82907
R19567 a_n2848_n452.n66 a_n2848_n452.t0 2.82907
R19568 a_n2848_n452.n68 a_n2848_n452.t2 2.82907
R19569 a_n2848_n452.n68 a_n2848_n452.t7 2.82907
R19570 a_n2848_n452.n64 a_n2848_n452.t9 2.82907
R19571 a_n2848_n452.n64 a_n2848_n452.t13 2.82907
R19572 a_n2848_n452.n62 a_n2848_n452.t10 2.82907
R19573 a_n2848_n452.n62 a_n2848_n452.t43 2.82907
R19574 a_n2848_n452.n60 a_n2848_n452.t4 2.82907
R19575 a_n2848_n452.n60 a_n2848_n452.t42 2.82907
R19576 a_n2848_n452.n56 a_n2848_n452.t17 2.82907
R19577 a_n2848_n452.n56 a_n2848_n452.t44 2.82907
R19578 a_n2848_n452.n57 a_n2848_n452.t15 2.82907
R19579 a_n2848_n452.n57 a_n2848_n452.t3 2.82907
R19580 a_n2848_n452.n59 a_n2848_n452.t16 2.82907
R19581 a_n2848_n452.n59 a_n2848_n452.t6 2.82907
R19582 a_n2848_n452.n55 a_n2848_n452.t46 2.82907
R19583 a_n2848_n452.n55 a_n2848_n452.t47 2.82907
R19584 a_n2848_n452.n53 a_n2848_n452.t1 2.82907
R19585 a_n2848_n452.n53 a_n2848_n452.t8 2.82907
R19586 a_n2848_n452.n52 a_n2848_n452.t11 2.82907
R19587 a_n2848_n452.n52 a_n2848_n452.t12 2.82907
R19588 a_n2848_n452.n102 a_n2848_n452.n13 1.30542
R19589 a_n2848_n452.n10 a_n2848_n452.n11 1.04595
R19590 a_n2848_n452.n5 a_n2848_n452.n97 13.657
R19591 a_n2848_n452.n95 a_n2848_n452.n50 21.4216
R19592 a_n2848_n452.n1 a_n2848_n452.n101 21.4216
R19593 a_n2848_n452.n98 a_n2848_n452.n47 21.4216
R19594 a_n2848_n452.n78 a_n2848_n452.n19 13.657
R19595 a_n2848_n452.n37 a_n2848_n452.n80 21.4216
R19596 a_n2848_n452.n75 a_n2848_n452.n23 13.657
R19597 a_n2848_n452.n34 a_n2848_n452.n77 21.4216
R19598 a_n2848_n452.n0 a_n2848_n452.n6 1.47777
R19599 a_n2848_n452.n22 a_n2848_n452.n21 0.758076
R19600 a_n2848_n452.n21 a_n2848_n452.n20 0.758076
R19601 a_n2848_n452.n18 a_n2848_n452.n17 0.758076
R19602 a_n2848_n452.n17 a_n2848_n452.n16 0.758076
R19603 a_n2848_n452.n15 a_n2848_n452.n14 0.758076
R19604 a_n2848_n452.n12 a_n2848_n452.n11 0.758076
R19605 a_n2848_n452.n10 a_n2848_n452.n9 0.758076
R19606 a_n2848_n452.n8 a_n2848_n452.n7 0.758076
R19607 a_n2848_n452.n4 a_n2848_n452.n2 0.758076
R19608 a_n2848_n452.n4 a_n2848_n452.n3 0.758076
R19609 a_n2848_n452.n27 a_n2848_n452.n26 0.716017
R19610 a_n2848_n452.n25 a_n2848_n452.n24 0.716017
R19611 a_n2848_n452.n12 a_n2848_n452.n14 0.67853
R19612 a_n2848_n452.n8 a_n2848_n452.n9 0.67853
R19613 a_n2848_n452.n28 a_n2848_n452.n54 0.530672
R19614 a_n2848_n452.n29 a_n2848_n452.n58 0.530672
R19615 a_n2848_n452.n63 a_n2848_n452.n61 0.530672
R19616 a_n2848_n452.n30 a_n2848_n452.n63 0.530672
R19617 a_n2848_n452.n31 a_n2848_n452.n67 0.530672
R19618 a_n2848_n452.n31 a_n2848_n452.n30 0.530672
R19619 a_n2848_n452.n29 a_n2848_n452.n28 0.530672
R19620 a_n1986_8322.n6 a_n1986_8322.t6 74.6477
R19621 a_n1986_8322.n1 a_n1986_8322.t13 74.6477
R19622 a_n1986_8322.t22 a_n1986_8322.n18 74.6476
R19623 a_n1986_8322.n14 a_n1986_8322.t15 74.2899
R19624 a_n1986_8322.n7 a_n1986_8322.t4 74.2899
R19625 a_n1986_8322.n8 a_n1986_8322.t7 74.2899
R19626 a_n1986_8322.n11 a_n1986_8322.t8 74.2899
R19627 a_n1986_8322.n4 a_n1986_8322.t12 74.2899
R19628 a_n1986_8322.n18 a_n1986_8322.n17 70.6783
R19629 a_n1986_8322.n16 a_n1986_8322.n15 70.6783
R19630 a_n1986_8322.n6 a_n1986_8322.n5 70.6783
R19631 a_n1986_8322.n10 a_n1986_8322.n9 70.6783
R19632 a_n1986_8322.n1 a_n1986_8322.n0 70.6783
R19633 a_n1986_8322.n3 a_n1986_8322.n2 70.6783
R19634 a_n1986_8322.n12 a_n1986_8322.n4 22.7556
R19635 a_n1986_8322.n13 a_n1986_8322.t2 9.7972
R19636 a_n1986_8322.n12 a_n1986_8322.n11 6.2408
R19637 a_n1986_8322.n14 a_n1986_8322.n13 5.83671
R19638 a_n1986_8322.n13 a_n1986_8322.n12 5.3452
R19639 a_n1986_8322.n17 a_n1986_8322.t20 3.61217
R19640 a_n1986_8322.n17 a_n1986_8322.t17 3.61217
R19641 a_n1986_8322.n15 a_n1986_8322.t14 3.61217
R19642 a_n1986_8322.n15 a_n1986_8322.t23 3.61217
R19643 a_n1986_8322.n5 a_n1986_8322.t10 3.61217
R19644 a_n1986_8322.n5 a_n1986_8322.t9 3.61217
R19645 a_n1986_8322.n9 a_n1986_8322.t5 3.61217
R19646 a_n1986_8322.n9 a_n1986_8322.t11 3.61217
R19647 a_n1986_8322.n0 a_n1986_8322.t21 3.61217
R19648 a_n1986_8322.n0 a_n1986_8322.t16 3.61217
R19649 a_n1986_8322.n2 a_n1986_8322.t19 3.61217
R19650 a_n1986_8322.n2 a_n1986_8322.t18 3.61217
R19651 a_n1986_8322.n11 a_n1986_8322.n10 0.358259
R19652 a_n1986_8322.n10 a_n1986_8322.n8 0.358259
R19653 a_n1986_8322.n7 a_n1986_8322.n6 0.358259
R19654 a_n1986_8322.n4 a_n1986_8322.n3 0.358259
R19655 a_n1986_8322.n3 a_n1986_8322.n1 0.358259
R19656 a_n1986_8322.n16 a_n1986_8322.n14 0.358259
R19657 a_n1986_8322.n18 a_n1986_8322.n16 0.358259
R19658 a_n1986_8322.n8 a_n1986_8322.n7 0.101793
R19659 a_n1986_8322.t3 a_n1986_8322.t0 0.0788333
R19660 a_n1986_8322.t1 a_n1986_8322.t3 0.0631667
R19661 a_n1986_8322.t2 a_n1986_8322.t1 0.0471944
R19662 a_n1986_8322.t2 a_n1986_8322.t0 0.0453889
R19663 a_n1808_13878.n16 a_n1808_13878.n0 98.9633
R19664 a_n1808_13878.n3 a_n1808_13878.n1 98.7517
R19665 a_n1808_13878.n5 a_n1808_13878.n4 98.6055
R19666 a_n1808_13878.n3 a_n1808_13878.n2 98.6055
R19667 a_n1808_13878.n17 a_n1808_13878.n16 98.6054
R19668 a_n1808_13878.n15 a_n1808_13878.n14 98.6054
R19669 a_n1808_13878.n7 a_n1808_13878.t1 74.6477
R19670 a_n1808_13878.n12 a_n1808_13878.t2 74.2899
R19671 a_n1808_13878.n9 a_n1808_13878.t3 74.2899
R19672 a_n1808_13878.n8 a_n1808_13878.t0 74.2899
R19673 a_n1808_13878.n11 a_n1808_13878.n10 70.6783
R19674 a_n1808_13878.n7 a_n1808_13878.n6 70.6783
R19675 a_n1808_13878.n13 a_n1808_13878.n5 13.5694
R19676 a_n1808_13878.n15 a_n1808_13878.n13 11.5762
R19677 a_n1808_13878.n13 a_n1808_13878.n12 6.2408
R19678 a_n1808_13878.n14 a_n1808_13878.t15 3.61217
R19679 a_n1808_13878.n14 a_n1808_13878.t16 3.61217
R19680 a_n1808_13878.n0 a_n1808_13878.t13 3.61217
R19681 a_n1808_13878.n0 a_n1808_13878.t17 3.61217
R19682 a_n1808_13878.n10 a_n1808_13878.t6 3.61217
R19683 a_n1808_13878.n10 a_n1808_13878.t7 3.61217
R19684 a_n1808_13878.n6 a_n1808_13878.t4 3.61217
R19685 a_n1808_13878.n6 a_n1808_13878.t5 3.61217
R19686 a_n1808_13878.n4 a_n1808_13878.t12 3.61217
R19687 a_n1808_13878.n4 a_n1808_13878.t19 3.61217
R19688 a_n1808_13878.n2 a_n1808_13878.t14 3.61217
R19689 a_n1808_13878.n2 a_n1808_13878.t9 3.61217
R19690 a_n1808_13878.n1 a_n1808_13878.t8 3.61217
R19691 a_n1808_13878.n1 a_n1808_13878.t10 3.61217
R19692 a_n1808_13878.t18 a_n1808_13878.n17 3.61217
R19693 a_n1808_13878.n17 a_n1808_13878.t11 3.61217
R19694 a_n1808_13878.n8 a_n1808_13878.n7 0.358259
R19695 a_n1808_13878.n11 a_n1808_13878.n9 0.358259
R19696 a_n1808_13878.n12 a_n1808_13878.n11 0.358259
R19697 a_n1808_13878.n16 a_n1808_13878.n15 0.358259
R19698 a_n1808_13878.n5 a_n1808_13878.n3 0.146627
R19699 a_n1808_13878.n9 a_n1808_13878.n8 0.101793
R19700 plus.n76 plus.t11 250.337
R19701 plus.n15 plus.t14 250.337
R19702 plus.n124 plus.t1 243.97
R19703 plus.n120 plus.t24 231.093
R19704 plus.n59 plus.t20 231.093
R19705 plus.n124 plus.n123 223.454
R19706 plus.n126 plus.n125 223.454
R19707 plus.n77 plus.t5 187.445
R19708 plus.n74 plus.t22 187.445
R19709 plus.n72 plus.t21 187.445
R19710 plus.n89 plus.t16 187.445
R19711 plus.n95 plus.t17 187.445
R19712 plus.n68 plus.t13 187.445
R19713 plus.n66 plus.t15 187.445
R19714 plus.n107 plus.t10 187.445
R19715 plus.n113 plus.t26 187.445
R19716 plus.n62 plus.t28 187.445
R19717 plus.n1 plus.t23 187.445
R19718 plus.n52 plus.t6 187.445
R19719 plus.n46 plus.t12 187.445
R19720 plus.n5 plus.t8 187.445
R19721 plus.n7 plus.t7 187.445
R19722 plus.n34 plus.t19 187.445
R19723 plus.n28 plus.t18 187.445
R19724 plus.n11 plus.t27 187.445
R19725 plus.n13 plus.t25 187.445
R19726 plus.n16 plus.t9 187.445
R19727 plus.n121 plus.n120 161.3
R19728 plus.n119 plus.n61 161.3
R19729 plus.n118 plus.n117 161.3
R19730 plus.n116 plus.n115 161.3
R19731 plus.n114 plus.n63 161.3
R19732 plus.n112 plus.n111 161.3
R19733 plus.n110 plus.n64 161.3
R19734 plus.n109 plus.n108 161.3
R19735 plus.n106 plus.n65 161.3
R19736 plus.n105 plus.n104 161.3
R19737 plus.n103 plus.n102 161.3
R19738 plus.n101 plus.n67 161.3
R19739 plus.n100 plus.n99 161.3
R19740 plus.n98 plus.n97 161.3
R19741 plus.n96 plus.n69 161.3
R19742 plus.n94 plus.n93 161.3
R19743 plus.n92 plus.n70 161.3
R19744 plus.n91 plus.n90 161.3
R19745 plus.n88 plus.n71 161.3
R19746 plus.n87 plus.n86 161.3
R19747 plus.n85 plus.n84 161.3
R19748 plus.n83 plus.n73 161.3
R19749 plus.n82 plus.n81 161.3
R19750 plus.n80 plus.n79 161.3
R19751 plus.n78 plus.n75 161.3
R19752 plus.n17 plus.n14 161.3
R19753 plus.n19 plus.n18 161.3
R19754 plus.n21 plus.n20 161.3
R19755 plus.n22 plus.n12 161.3
R19756 plus.n24 plus.n23 161.3
R19757 plus.n26 plus.n25 161.3
R19758 plus.n27 plus.n10 161.3
R19759 plus.n30 plus.n29 161.3
R19760 plus.n31 plus.n9 161.3
R19761 plus.n33 plus.n32 161.3
R19762 plus.n35 plus.n8 161.3
R19763 plus.n37 plus.n36 161.3
R19764 plus.n39 plus.n38 161.3
R19765 plus.n40 plus.n6 161.3
R19766 plus.n42 plus.n41 161.3
R19767 plus.n44 plus.n43 161.3
R19768 plus.n45 plus.n4 161.3
R19769 plus.n48 plus.n47 161.3
R19770 plus.n49 plus.n3 161.3
R19771 plus.n51 plus.n50 161.3
R19772 plus.n53 plus.n2 161.3
R19773 plus.n55 plus.n54 161.3
R19774 plus.n57 plus.n56 161.3
R19775 plus.n58 plus.n0 161.3
R19776 plus.n60 plus.n59 161.3
R19777 plus.n88 plus.n87 56.5617
R19778 plus.n97 plus.n96 56.5617
R19779 plus.n106 plus.n105 56.5617
R19780 plus.n45 plus.n44 56.5617
R19781 plus.n36 plus.n35 56.5617
R19782 plus.n27 plus.n26 56.5617
R19783 plus.n79 plus.n78 56.5617
R19784 plus.n115 plus.n114 56.5617
R19785 plus.n54 plus.n53 56.5617
R19786 plus.n18 plus.n17 56.5617
R19787 plus.n119 plus.n118 50.2647
R19788 plus.n58 plus.n57 50.2647
R19789 plus.n84 plus.n83 46.3896
R19790 plus.n108 plus.n64 46.3896
R19791 plus.n47 plus.n3 46.3896
R19792 plus.n23 plus.n22 46.3896
R19793 plus.n76 plus.n75 43.1929
R19794 plus.n15 plus.n14 43.1929
R19795 plus.n94 plus.n70 42.5146
R19796 plus.n101 plus.n100 42.5146
R19797 plus.n40 plus.n39 42.5146
R19798 plus.n33 plus.n9 42.5146
R19799 plus.n77 plus.n76 40.6041
R19800 plus.n16 plus.n15 40.6041
R19801 plus.n90 plus.n70 38.6395
R19802 plus.n102 plus.n101 38.6395
R19803 plus.n41 plus.n40 38.6395
R19804 plus.n29 plus.n9 38.6395
R19805 plus.n122 plus.n121 35.2031
R19806 plus.n83 plus.n82 34.7644
R19807 plus.n112 plus.n64 34.7644
R19808 plus.n51 plus.n3 34.7644
R19809 plus.n22 plus.n21 34.7644
R19810 plus.n79 plus.n74 21.8872
R19811 plus.n114 plus.n113 21.8872
R19812 plus.n53 plus.n52 21.8872
R19813 plus.n18 plus.n13 21.8872
R19814 plus.n89 plus.n88 19.9199
R19815 plus.n105 plus.n66 19.9199
R19816 plus.n44 plus.n5 19.9199
R19817 plus.n28 plus.n27 19.9199
R19818 plus.n123 plus.t2 19.8005
R19819 plus.n123 plus.t4 19.8005
R19820 plus.n125 plus.t3 19.8005
R19821 plus.n125 plus.t0 19.8005
R19822 plus.n96 plus.n95 17.9525
R19823 plus.n97 plus.n68 17.9525
R19824 plus.n36 plus.n7 17.9525
R19825 plus.n35 plus.n34 17.9525
R19826 plus.n87 plus.n72 15.9852
R19827 plus.n107 plus.n106 15.9852
R19828 plus.n46 plus.n45 15.9852
R19829 plus.n26 plus.n11 15.9852
R19830 plus plus.n127 14.4034
R19831 plus.n78 plus.n77 14.0178
R19832 plus.n115 plus.n62 14.0178
R19833 plus.n54 plus.n1 14.0178
R19834 plus.n17 plus.n16 14.0178
R19835 plus.n122 plus.n60 11.9342
R19836 plus.n118 plus.n62 10.575
R19837 plus.n57 plus.n1 10.575
R19838 plus.n120 plus.n119 9.49444
R19839 plus.n59 plus.n58 9.49444
R19840 plus.n84 plus.n72 8.60764
R19841 plus.n108 plus.n107 8.60764
R19842 plus.n47 plus.n46 8.60764
R19843 plus.n23 plus.n11 8.60764
R19844 plus.n95 plus.n94 6.6403
R19845 plus.n100 plus.n68 6.6403
R19846 plus.n39 plus.n7 6.6403
R19847 plus.n34 plus.n33 6.6403
R19848 plus.n127 plus.n126 5.40567
R19849 plus.n90 plus.n89 4.67295
R19850 plus.n102 plus.n66 4.67295
R19851 plus.n41 plus.n5 4.67295
R19852 plus.n29 plus.n28 4.67295
R19853 plus.n82 plus.n74 2.7056
R19854 plus.n113 plus.n112 2.7056
R19855 plus.n52 plus.n51 2.7056
R19856 plus.n21 plus.n13 2.7056
R19857 plus.n127 plus.n122 1.188
R19858 plus.n126 plus.n124 0.716017
R19859 plus.n80 plus.n75 0.189894
R19860 plus.n81 plus.n80 0.189894
R19861 plus.n81 plus.n73 0.189894
R19862 plus.n85 plus.n73 0.189894
R19863 plus.n86 plus.n85 0.189894
R19864 plus.n86 plus.n71 0.189894
R19865 plus.n91 plus.n71 0.189894
R19866 plus.n92 plus.n91 0.189894
R19867 plus.n93 plus.n92 0.189894
R19868 plus.n93 plus.n69 0.189894
R19869 plus.n98 plus.n69 0.189894
R19870 plus.n99 plus.n98 0.189894
R19871 plus.n99 plus.n67 0.189894
R19872 plus.n103 plus.n67 0.189894
R19873 plus.n104 plus.n103 0.189894
R19874 plus.n104 plus.n65 0.189894
R19875 plus.n109 plus.n65 0.189894
R19876 plus.n110 plus.n109 0.189894
R19877 plus.n111 plus.n110 0.189894
R19878 plus.n111 plus.n63 0.189894
R19879 plus.n116 plus.n63 0.189894
R19880 plus.n117 plus.n116 0.189894
R19881 plus.n117 plus.n61 0.189894
R19882 plus.n121 plus.n61 0.189894
R19883 plus.n60 plus.n0 0.189894
R19884 plus.n56 plus.n0 0.189894
R19885 plus.n56 plus.n55 0.189894
R19886 plus.n55 plus.n2 0.189894
R19887 plus.n50 plus.n2 0.189894
R19888 plus.n50 plus.n49 0.189894
R19889 plus.n49 plus.n48 0.189894
R19890 plus.n48 plus.n4 0.189894
R19891 plus.n43 plus.n4 0.189894
R19892 plus.n43 plus.n42 0.189894
R19893 plus.n42 plus.n6 0.189894
R19894 plus.n38 plus.n6 0.189894
R19895 plus.n38 plus.n37 0.189894
R19896 plus.n37 plus.n8 0.189894
R19897 plus.n32 plus.n8 0.189894
R19898 plus.n32 plus.n31 0.189894
R19899 plus.n31 plus.n30 0.189894
R19900 plus.n30 plus.n10 0.189894
R19901 plus.n25 plus.n10 0.189894
R19902 plus.n25 plus.n24 0.189894
R19903 plus.n24 plus.n12 0.189894
R19904 plus.n20 plus.n12 0.189894
R19905 plus.n20 plus.n19 0.189894
R19906 plus.n19 plus.n14 0.189894
R19907 a_n3106_n452.n1 a_n3106_n452.t10 214.321
R19908 a_n3106_n452.n14 a_n3106_n452.t9 214.321
R19909 a_n3106_n452.n15 a_n3106_n452.t49 214.321
R19910 a_n3106_n452.n16 a_n3106_n452.t48 214.321
R19911 a_n3106_n452.n17 a_n3106_n452.t41 214.321
R19912 a_n3106_n452.n18 a_n3106_n452.t11 214.321
R19913 a_n3106_n452.n19 a_n3106_n452.t16 214.321
R19914 a_n3106_n452.n20 a_n3106_n452.t15 214.321
R19915 a_n3106_n452.n0 a_n3106_n452.t34 55.8337
R19916 a_n3106_n452.n2 a_n3106_n452.t53 55.8337
R19917 a_n3106_n452.n13 a_n3106_n452.t4 55.8337
R19918 a_n3106_n452.n47 a_n3106_n452.t21 55.8335
R19919 a_n3106_n452.n45 a_n3106_n452.t52 55.8335
R19920 a_n3106_n452.n34 a_n3106_n452.t14 55.8335
R19921 a_n3106_n452.n33 a_n3106_n452.t31 55.8335
R19922 a_n3106_n452.n22 a_n3106_n452.t25 55.8335
R19923 a_n3106_n452.n49 a_n3106_n452.n48 53.0052
R19924 a_n3106_n452.n51 a_n3106_n452.n50 53.0052
R19925 a_n3106_n452.n53 a_n3106_n452.n52 53.0052
R19926 a_n3106_n452.n55 a_n3106_n452.n54 53.0052
R19927 a_n3106_n452.n4 a_n3106_n452.n3 53.0052
R19928 a_n3106_n452.n6 a_n3106_n452.n5 53.0052
R19929 a_n3106_n452.n8 a_n3106_n452.n7 53.0052
R19930 a_n3106_n452.n10 a_n3106_n452.n9 53.0052
R19931 a_n3106_n452.n12 a_n3106_n452.n11 53.0052
R19932 a_n3106_n452.n44 a_n3106_n452.n43 53.0051
R19933 a_n3106_n452.n42 a_n3106_n452.n41 53.0051
R19934 a_n3106_n452.n40 a_n3106_n452.n39 53.0051
R19935 a_n3106_n452.n38 a_n3106_n452.n37 53.0051
R19936 a_n3106_n452.n36 a_n3106_n452.n35 53.0051
R19937 a_n3106_n452.n32 a_n3106_n452.n31 53.0051
R19938 a_n3106_n452.n30 a_n3106_n452.n29 53.0051
R19939 a_n3106_n452.n28 a_n3106_n452.n27 53.0051
R19940 a_n3106_n452.n26 a_n3106_n452.n25 53.0051
R19941 a_n3106_n452.n24 a_n3106_n452.n23 53.0051
R19942 a_n3106_n452.n57 a_n3106_n452.n56 53.0051
R19943 a_n3106_n452.n21 a_n3106_n452.n13 12.2417
R19944 a_n3106_n452.n47 a_n3106_n452.n46 12.2417
R19945 a_n3106_n452.n22 a_n3106_n452.n21 5.16214
R19946 a_n3106_n452.n46 a_n3106_n452.n45 5.16214
R19947 a_n3106_n452.n48 a_n3106_n452.t19 2.82907
R19948 a_n3106_n452.n48 a_n3106_n452.t17 2.82907
R19949 a_n3106_n452.n50 a_n3106_n452.t30 2.82907
R19950 a_n3106_n452.n50 a_n3106_n452.t35 2.82907
R19951 a_n3106_n452.n52 a_n3106_n452.t28 2.82907
R19952 a_n3106_n452.n52 a_n3106_n452.t32 2.82907
R19953 a_n3106_n452.n54 a_n3106_n452.t24 2.82907
R19954 a_n3106_n452.n54 a_n3106_n452.t29 2.82907
R19955 a_n3106_n452.n3 a_n3106_n452.t0 2.82907
R19956 a_n3106_n452.n3 a_n3106_n452.t5 2.82907
R19957 a_n3106_n452.n5 a_n3106_n452.t7 2.82907
R19958 a_n3106_n452.n5 a_n3106_n452.t44 2.82907
R19959 a_n3106_n452.n7 a_n3106_n452.t43 2.82907
R19960 a_n3106_n452.n7 a_n3106_n452.t2 2.82907
R19961 a_n3106_n452.n9 a_n3106_n452.t51 2.82907
R19962 a_n3106_n452.n9 a_n3106_n452.t12 2.82907
R19963 a_n3106_n452.n11 a_n3106_n452.t50 2.82907
R19964 a_n3106_n452.n11 a_n3106_n452.t13 2.82907
R19965 a_n3106_n452.n43 a_n3106_n452.t3 2.82907
R19966 a_n3106_n452.n43 a_n3106_n452.t47 2.82907
R19967 a_n3106_n452.n41 a_n3106_n452.t6 2.82907
R19968 a_n3106_n452.n41 a_n3106_n452.t45 2.82907
R19969 a_n3106_n452.n39 a_n3106_n452.t55 2.82907
R19970 a_n3106_n452.n39 a_n3106_n452.t46 2.82907
R19971 a_n3106_n452.n37 a_n3106_n452.t8 2.82907
R19972 a_n3106_n452.n37 a_n3106_n452.t54 2.82907
R19973 a_n3106_n452.n35 a_n3106_n452.t42 2.82907
R19974 a_n3106_n452.n35 a_n3106_n452.t1 2.82907
R19975 a_n3106_n452.n31 a_n3106_n452.t20 2.82907
R19976 a_n3106_n452.n31 a_n3106_n452.t36 2.82907
R19977 a_n3106_n452.n29 a_n3106_n452.t27 2.82907
R19978 a_n3106_n452.n29 a_n3106_n452.t18 2.82907
R19979 a_n3106_n452.n27 a_n3106_n452.t38 2.82907
R19980 a_n3106_n452.n27 a_n3106_n452.t26 2.82907
R19981 a_n3106_n452.n25 a_n3106_n452.t33 2.82907
R19982 a_n3106_n452.n25 a_n3106_n452.t37 2.82907
R19983 a_n3106_n452.n23 a_n3106_n452.t22 2.82907
R19984 a_n3106_n452.n23 a_n3106_n452.t39 2.82907
R19985 a_n3106_n452.t40 a_n3106_n452.n57 2.82907
R19986 a_n3106_n452.n57 a_n3106_n452.t23 2.82907
R19987 a_n3106_n452.n46 a_n3106_n452.n1 2.54197
R19988 a_n3106_n452.n21 a_n3106_n452.n20 2.0129
R19989 a_n3106_n452.n20 a_n3106_n452.n19 0.672012
R19990 a_n3106_n452.n19 a_n3106_n452.n18 0.672012
R19991 a_n3106_n452.n18 a_n3106_n452.n17 0.672012
R19992 a_n3106_n452.n17 a_n3106_n452.n16 0.672012
R19993 a_n3106_n452.n16 a_n3106_n452.n15 0.672012
R19994 a_n3106_n452.n15 a_n3106_n452.n14 0.672012
R19995 a_n3106_n452.n14 a_n3106_n452.n1 0.672012
R19996 a_n3106_n452.n24 a_n3106_n452.n22 0.530672
R19997 a_n3106_n452.n26 a_n3106_n452.n24 0.530672
R19998 a_n3106_n452.n28 a_n3106_n452.n26 0.530672
R19999 a_n3106_n452.n30 a_n3106_n452.n28 0.530672
R20000 a_n3106_n452.n32 a_n3106_n452.n30 0.530672
R20001 a_n3106_n452.n33 a_n3106_n452.n32 0.530672
R20002 a_n3106_n452.n36 a_n3106_n452.n34 0.530672
R20003 a_n3106_n452.n38 a_n3106_n452.n36 0.530672
R20004 a_n3106_n452.n40 a_n3106_n452.n38 0.530672
R20005 a_n3106_n452.n42 a_n3106_n452.n40 0.530672
R20006 a_n3106_n452.n44 a_n3106_n452.n42 0.530672
R20007 a_n3106_n452.n45 a_n3106_n452.n44 0.530672
R20008 a_n3106_n452.n13 a_n3106_n452.n12 0.530672
R20009 a_n3106_n452.n12 a_n3106_n452.n10 0.530672
R20010 a_n3106_n452.n10 a_n3106_n452.n8 0.530672
R20011 a_n3106_n452.n8 a_n3106_n452.n6 0.530672
R20012 a_n3106_n452.n6 a_n3106_n452.n4 0.530672
R20013 a_n3106_n452.n4 a_n3106_n452.n2 0.530672
R20014 a_n3106_n452.n56 a_n3106_n452.n0 0.530672
R20015 a_n3106_n452.n56 a_n3106_n452.n55 0.530672
R20016 a_n3106_n452.n55 a_n3106_n452.n53 0.530672
R20017 a_n3106_n452.n53 a_n3106_n452.n51 0.530672
R20018 a_n3106_n452.n51 a_n3106_n452.n49 0.530672
R20019 a_n3106_n452.n49 a_n3106_n452.n47 0.530672
R20020 a_n3106_n452.n34 a_n3106_n452.n33 0.235414
R20021 a_n3106_n452.n2 a_n3106_n452.n0 0.235414
R20022 outputibias.n27 outputibias.n1 289.615
R20023 outputibias.n58 outputibias.n32 289.615
R20024 outputibias.n90 outputibias.n64 289.615
R20025 outputibias.n122 outputibias.n96 289.615
R20026 outputibias.n28 outputibias.n27 185
R20027 outputibias.n26 outputibias.n25 185
R20028 outputibias.n5 outputibias.n4 185
R20029 outputibias.n20 outputibias.n19 185
R20030 outputibias.n18 outputibias.n17 185
R20031 outputibias.n9 outputibias.n8 185
R20032 outputibias.n12 outputibias.n11 185
R20033 outputibias.n59 outputibias.n58 185
R20034 outputibias.n57 outputibias.n56 185
R20035 outputibias.n36 outputibias.n35 185
R20036 outputibias.n51 outputibias.n50 185
R20037 outputibias.n49 outputibias.n48 185
R20038 outputibias.n40 outputibias.n39 185
R20039 outputibias.n43 outputibias.n42 185
R20040 outputibias.n91 outputibias.n90 185
R20041 outputibias.n89 outputibias.n88 185
R20042 outputibias.n68 outputibias.n67 185
R20043 outputibias.n83 outputibias.n82 185
R20044 outputibias.n81 outputibias.n80 185
R20045 outputibias.n72 outputibias.n71 185
R20046 outputibias.n75 outputibias.n74 185
R20047 outputibias.n123 outputibias.n122 185
R20048 outputibias.n121 outputibias.n120 185
R20049 outputibias.n100 outputibias.n99 185
R20050 outputibias.n115 outputibias.n114 185
R20051 outputibias.n113 outputibias.n112 185
R20052 outputibias.n104 outputibias.n103 185
R20053 outputibias.n107 outputibias.n106 185
R20054 outputibias.n0 outputibias.t8 178.945
R20055 outputibias.n133 outputibias.t10 177.018
R20056 outputibias.n132 outputibias.t11 177.018
R20057 outputibias.n0 outputibias.t9 177.018
R20058 outputibias.t5 outputibias.n10 147.661
R20059 outputibias.t7 outputibias.n41 147.661
R20060 outputibias.t1 outputibias.n73 147.661
R20061 outputibias.t3 outputibias.n105 147.661
R20062 outputibias.n128 outputibias.t4 132.363
R20063 outputibias.n128 outputibias.t6 130.436
R20064 outputibias.n129 outputibias.t0 130.436
R20065 outputibias.n130 outputibias.t2 130.436
R20066 outputibias.n27 outputibias.n26 104.615
R20067 outputibias.n26 outputibias.n4 104.615
R20068 outputibias.n19 outputibias.n4 104.615
R20069 outputibias.n19 outputibias.n18 104.615
R20070 outputibias.n18 outputibias.n8 104.615
R20071 outputibias.n11 outputibias.n8 104.615
R20072 outputibias.n58 outputibias.n57 104.615
R20073 outputibias.n57 outputibias.n35 104.615
R20074 outputibias.n50 outputibias.n35 104.615
R20075 outputibias.n50 outputibias.n49 104.615
R20076 outputibias.n49 outputibias.n39 104.615
R20077 outputibias.n42 outputibias.n39 104.615
R20078 outputibias.n90 outputibias.n89 104.615
R20079 outputibias.n89 outputibias.n67 104.615
R20080 outputibias.n82 outputibias.n67 104.615
R20081 outputibias.n82 outputibias.n81 104.615
R20082 outputibias.n81 outputibias.n71 104.615
R20083 outputibias.n74 outputibias.n71 104.615
R20084 outputibias.n122 outputibias.n121 104.615
R20085 outputibias.n121 outputibias.n99 104.615
R20086 outputibias.n114 outputibias.n99 104.615
R20087 outputibias.n114 outputibias.n113 104.615
R20088 outputibias.n113 outputibias.n103 104.615
R20089 outputibias.n106 outputibias.n103 104.615
R20090 outputibias.n63 outputibias.n31 95.6354
R20091 outputibias.n63 outputibias.n62 94.6732
R20092 outputibias.n95 outputibias.n94 94.6732
R20093 outputibias.n127 outputibias.n126 94.6732
R20094 outputibias.n11 outputibias.t5 52.3082
R20095 outputibias.n42 outputibias.t7 52.3082
R20096 outputibias.n74 outputibias.t1 52.3082
R20097 outputibias.n106 outputibias.t3 52.3082
R20098 outputibias.n12 outputibias.n10 15.6674
R20099 outputibias.n43 outputibias.n41 15.6674
R20100 outputibias.n75 outputibias.n73 15.6674
R20101 outputibias.n107 outputibias.n105 15.6674
R20102 outputibias.n13 outputibias.n9 12.8005
R20103 outputibias.n44 outputibias.n40 12.8005
R20104 outputibias.n76 outputibias.n72 12.8005
R20105 outputibias.n108 outputibias.n104 12.8005
R20106 outputibias.n17 outputibias.n16 12.0247
R20107 outputibias.n48 outputibias.n47 12.0247
R20108 outputibias.n80 outputibias.n79 12.0247
R20109 outputibias.n112 outputibias.n111 12.0247
R20110 outputibias.n20 outputibias.n7 11.249
R20111 outputibias.n51 outputibias.n38 11.249
R20112 outputibias.n83 outputibias.n70 11.249
R20113 outputibias.n115 outputibias.n102 11.249
R20114 outputibias.n21 outputibias.n5 10.4732
R20115 outputibias.n52 outputibias.n36 10.4732
R20116 outputibias.n84 outputibias.n68 10.4732
R20117 outputibias.n116 outputibias.n100 10.4732
R20118 outputibias.n25 outputibias.n24 9.69747
R20119 outputibias.n56 outputibias.n55 9.69747
R20120 outputibias.n88 outputibias.n87 9.69747
R20121 outputibias.n120 outputibias.n119 9.69747
R20122 outputibias.n31 outputibias.n30 9.45567
R20123 outputibias.n62 outputibias.n61 9.45567
R20124 outputibias.n94 outputibias.n93 9.45567
R20125 outputibias.n126 outputibias.n125 9.45567
R20126 outputibias.n30 outputibias.n29 9.3005
R20127 outputibias.n3 outputibias.n2 9.3005
R20128 outputibias.n24 outputibias.n23 9.3005
R20129 outputibias.n22 outputibias.n21 9.3005
R20130 outputibias.n7 outputibias.n6 9.3005
R20131 outputibias.n16 outputibias.n15 9.3005
R20132 outputibias.n14 outputibias.n13 9.3005
R20133 outputibias.n61 outputibias.n60 9.3005
R20134 outputibias.n34 outputibias.n33 9.3005
R20135 outputibias.n55 outputibias.n54 9.3005
R20136 outputibias.n53 outputibias.n52 9.3005
R20137 outputibias.n38 outputibias.n37 9.3005
R20138 outputibias.n47 outputibias.n46 9.3005
R20139 outputibias.n45 outputibias.n44 9.3005
R20140 outputibias.n93 outputibias.n92 9.3005
R20141 outputibias.n66 outputibias.n65 9.3005
R20142 outputibias.n87 outputibias.n86 9.3005
R20143 outputibias.n85 outputibias.n84 9.3005
R20144 outputibias.n70 outputibias.n69 9.3005
R20145 outputibias.n79 outputibias.n78 9.3005
R20146 outputibias.n77 outputibias.n76 9.3005
R20147 outputibias.n125 outputibias.n124 9.3005
R20148 outputibias.n98 outputibias.n97 9.3005
R20149 outputibias.n119 outputibias.n118 9.3005
R20150 outputibias.n117 outputibias.n116 9.3005
R20151 outputibias.n102 outputibias.n101 9.3005
R20152 outputibias.n111 outputibias.n110 9.3005
R20153 outputibias.n109 outputibias.n108 9.3005
R20154 outputibias.n28 outputibias.n3 8.92171
R20155 outputibias.n59 outputibias.n34 8.92171
R20156 outputibias.n91 outputibias.n66 8.92171
R20157 outputibias.n123 outputibias.n98 8.92171
R20158 outputibias.n29 outputibias.n1 8.14595
R20159 outputibias.n60 outputibias.n32 8.14595
R20160 outputibias.n92 outputibias.n64 8.14595
R20161 outputibias.n124 outputibias.n96 8.14595
R20162 outputibias.n31 outputibias.n1 5.81868
R20163 outputibias.n62 outputibias.n32 5.81868
R20164 outputibias.n94 outputibias.n64 5.81868
R20165 outputibias.n126 outputibias.n96 5.81868
R20166 outputibias.n131 outputibias.n130 5.20947
R20167 outputibias.n29 outputibias.n28 5.04292
R20168 outputibias.n60 outputibias.n59 5.04292
R20169 outputibias.n92 outputibias.n91 5.04292
R20170 outputibias.n124 outputibias.n123 5.04292
R20171 outputibias.n131 outputibias.n127 4.42209
R20172 outputibias.n14 outputibias.n10 4.38594
R20173 outputibias.n45 outputibias.n41 4.38594
R20174 outputibias.n77 outputibias.n73 4.38594
R20175 outputibias.n109 outputibias.n105 4.38594
R20176 outputibias.n132 outputibias.n131 4.28454
R20177 outputibias.n25 outputibias.n3 4.26717
R20178 outputibias.n56 outputibias.n34 4.26717
R20179 outputibias.n88 outputibias.n66 4.26717
R20180 outputibias.n120 outputibias.n98 4.26717
R20181 outputibias.n24 outputibias.n5 3.49141
R20182 outputibias.n55 outputibias.n36 3.49141
R20183 outputibias.n87 outputibias.n68 3.49141
R20184 outputibias.n119 outputibias.n100 3.49141
R20185 outputibias.n21 outputibias.n20 2.71565
R20186 outputibias.n52 outputibias.n51 2.71565
R20187 outputibias.n84 outputibias.n83 2.71565
R20188 outputibias.n116 outputibias.n115 2.71565
R20189 outputibias.n17 outputibias.n7 1.93989
R20190 outputibias.n48 outputibias.n38 1.93989
R20191 outputibias.n80 outputibias.n70 1.93989
R20192 outputibias.n112 outputibias.n102 1.93989
R20193 outputibias.n130 outputibias.n129 1.9266
R20194 outputibias.n129 outputibias.n128 1.9266
R20195 outputibias.n133 outputibias.n132 1.92658
R20196 outputibias.n134 outputibias.n133 1.29913
R20197 outputibias.n16 outputibias.n9 1.16414
R20198 outputibias.n47 outputibias.n40 1.16414
R20199 outputibias.n79 outputibias.n72 1.16414
R20200 outputibias.n111 outputibias.n104 1.16414
R20201 outputibias.n127 outputibias.n95 0.962709
R20202 outputibias.n95 outputibias.n63 0.962709
R20203 outputibias.n13 outputibias.n12 0.388379
R20204 outputibias.n44 outputibias.n43 0.388379
R20205 outputibias.n76 outputibias.n75 0.388379
R20206 outputibias.n108 outputibias.n107 0.388379
R20207 outputibias.n134 outputibias.n0 0.337251
R20208 outputibias outputibias.n134 0.302375
R20209 outputibias.n30 outputibias.n2 0.155672
R20210 outputibias.n23 outputibias.n2 0.155672
R20211 outputibias.n23 outputibias.n22 0.155672
R20212 outputibias.n22 outputibias.n6 0.155672
R20213 outputibias.n15 outputibias.n6 0.155672
R20214 outputibias.n15 outputibias.n14 0.155672
R20215 outputibias.n61 outputibias.n33 0.155672
R20216 outputibias.n54 outputibias.n33 0.155672
R20217 outputibias.n54 outputibias.n53 0.155672
R20218 outputibias.n53 outputibias.n37 0.155672
R20219 outputibias.n46 outputibias.n37 0.155672
R20220 outputibias.n46 outputibias.n45 0.155672
R20221 outputibias.n93 outputibias.n65 0.155672
R20222 outputibias.n86 outputibias.n65 0.155672
R20223 outputibias.n86 outputibias.n85 0.155672
R20224 outputibias.n85 outputibias.n69 0.155672
R20225 outputibias.n78 outputibias.n69 0.155672
R20226 outputibias.n78 outputibias.n77 0.155672
R20227 outputibias.n125 outputibias.n97 0.155672
R20228 outputibias.n118 outputibias.n97 0.155672
R20229 outputibias.n118 outputibias.n117 0.155672
R20230 outputibias.n117 outputibias.n101 0.155672
R20231 outputibias.n110 outputibias.n101 0.155672
R20232 outputibias.n110 outputibias.n109 0.155672
R20233 output.n41 output.n15 289.615
R20234 output.n72 output.n46 289.615
R20235 output.n104 output.n78 289.615
R20236 output.n136 output.n110 289.615
R20237 output.n77 output.n45 197.26
R20238 output.n77 output.n76 196.298
R20239 output.n109 output.n108 196.298
R20240 output.n141 output.n140 196.298
R20241 output.n42 output.n41 185
R20242 output.n40 output.n39 185
R20243 output.n19 output.n18 185
R20244 output.n34 output.n33 185
R20245 output.n32 output.n31 185
R20246 output.n23 output.n22 185
R20247 output.n26 output.n25 185
R20248 output.n73 output.n72 185
R20249 output.n71 output.n70 185
R20250 output.n50 output.n49 185
R20251 output.n65 output.n64 185
R20252 output.n63 output.n62 185
R20253 output.n54 output.n53 185
R20254 output.n57 output.n56 185
R20255 output.n105 output.n104 185
R20256 output.n103 output.n102 185
R20257 output.n82 output.n81 185
R20258 output.n97 output.n96 185
R20259 output.n95 output.n94 185
R20260 output.n86 output.n85 185
R20261 output.n89 output.n88 185
R20262 output.n137 output.n136 185
R20263 output.n135 output.n134 185
R20264 output.n114 output.n113 185
R20265 output.n129 output.n128 185
R20266 output.n127 output.n126 185
R20267 output.n118 output.n117 185
R20268 output.n121 output.n120 185
R20269 output.t19 output.n24 147.661
R20270 output.t18 output.n55 147.661
R20271 output.t17 output.n87 147.661
R20272 output.t16 output.n119 147.661
R20273 output.n41 output.n40 104.615
R20274 output.n40 output.n18 104.615
R20275 output.n33 output.n18 104.615
R20276 output.n33 output.n32 104.615
R20277 output.n32 output.n22 104.615
R20278 output.n25 output.n22 104.615
R20279 output.n72 output.n71 104.615
R20280 output.n71 output.n49 104.615
R20281 output.n64 output.n49 104.615
R20282 output.n64 output.n63 104.615
R20283 output.n63 output.n53 104.615
R20284 output.n56 output.n53 104.615
R20285 output.n104 output.n103 104.615
R20286 output.n103 output.n81 104.615
R20287 output.n96 output.n81 104.615
R20288 output.n96 output.n95 104.615
R20289 output.n95 output.n85 104.615
R20290 output.n88 output.n85 104.615
R20291 output.n136 output.n135 104.615
R20292 output.n135 output.n113 104.615
R20293 output.n128 output.n113 104.615
R20294 output.n128 output.n127 104.615
R20295 output.n127 output.n117 104.615
R20296 output.n120 output.n117 104.615
R20297 output.n1 output.t15 77.056
R20298 output.n14 output.t0 76.6694
R20299 output.n1 output.n0 72.7095
R20300 output.n3 output.n2 72.7095
R20301 output.n5 output.n4 72.7095
R20302 output.n7 output.n6 72.7095
R20303 output.n9 output.n8 72.7095
R20304 output.n11 output.n10 72.7095
R20305 output.n13 output.n12 72.7095
R20306 output.n25 output.t19 52.3082
R20307 output.n56 output.t18 52.3082
R20308 output.n88 output.t17 52.3082
R20309 output.n120 output.t16 52.3082
R20310 output.n26 output.n24 15.6674
R20311 output.n57 output.n55 15.6674
R20312 output.n89 output.n87 15.6674
R20313 output.n121 output.n119 15.6674
R20314 output.n27 output.n23 12.8005
R20315 output.n58 output.n54 12.8005
R20316 output.n90 output.n86 12.8005
R20317 output.n122 output.n118 12.8005
R20318 output.n31 output.n30 12.0247
R20319 output.n62 output.n61 12.0247
R20320 output.n94 output.n93 12.0247
R20321 output.n126 output.n125 12.0247
R20322 output.n34 output.n21 11.249
R20323 output.n65 output.n52 11.249
R20324 output.n97 output.n84 11.249
R20325 output.n129 output.n116 11.249
R20326 output.n35 output.n19 10.4732
R20327 output.n66 output.n50 10.4732
R20328 output.n98 output.n82 10.4732
R20329 output.n130 output.n114 10.4732
R20330 output.n39 output.n38 9.69747
R20331 output.n70 output.n69 9.69747
R20332 output.n102 output.n101 9.69747
R20333 output.n134 output.n133 9.69747
R20334 output.n45 output.n44 9.45567
R20335 output.n76 output.n75 9.45567
R20336 output.n108 output.n107 9.45567
R20337 output.n140 output.n139 9.45567
R20338 output.n44 output.n43 9.3005
R20339 output.n17 output.n16 9.3005
R20340 output.n38 output.n37 9.3005
R20341 output.n36 output.n35 9.3005
R20342 output.n21 output.n20 9.3005
R20343 output.n30 output.n29 9.3005
R20344 output.n28 output.n27 9.3005
R20345 output.n75 output.n74 9.3005
R20346 output.n48 output.n47 9.3005
R20347 output.n69 output.n68 9.3005
R20348 output.n67 output.n66 9.3005
R20349 output.n52 output.n51 9.3005
R20350 output.n61 output.n60 9.3005
R20351 output.n59 output.n58 9.3005
R20352 output.n107 output.n106 9.3005
R20353 output.n80 output.n79 9.3005
R20354 output.n101 output.n100 9.3005
R20355 output.n99 output.n98 9.3005
R20356 output.n84 output.n83 9.3005
R20357 output.n93 output.n92 9.3005
R20358 output.n91 output.n90 9.3005
R20359 output.n139 output.n138 9.3005
R20360 output.n112 output.n111 9.3005
R20361 output.n133 output.n132 9.3005
R20362 output.n131 output.n130 9.3005
R20363 output.n116 output.n115 9.3005
R20364 output.n125 output.n124 9.3005
R20365 output.n123 output.n122 9.3005
R20366 output.n42 output.n17 8.92171
R20367 output.n73 output.n48 8.92171
R20368 output.n105 output.n80 8.92171
R20369 output.n137 output.n112 8.92171
R20370 output output.n141 8.15037
R20371 output.n43 output.n15 8.14595
R20372 output.n74 output.n46 8.14595
R20373 output.n106 output.n78 8.14595
R20374 output.n138 output.n110 8.14595
R20375 output.n45 output.n15 5.81868
R20376 output.n76 output.n46 5.81868
R20377 output.n108 output.n78 5.81868
R20378 output.n140 output.n110 5.81868
R20379 output.n43 output.n42 5.04292
R20380 output.n74 output.n73 5.04292
R20381 output.n106 output.n105 5.04292
R20382 output.n138 output.n137 5.04292
R20383 output.n28 output.n24 4.38594
R20384 output.n59 output.n55 4.38594
R20385 output.n91 output.n87 4.38594
R20386 output.n123 output.n119 4.38594
R20387 output.n39 output.n17 4.26717
R20388 output.n70 output.n48 4.26717
R20389 output.n102 output.n80 4.26717
R20390 output.n134 output.n112 4.26717
R20391 output.n0 output.t5 3.9605
R20392 output.n0 output.t9 3.9605
R20393 output.n2 output.t12 3.9605
R20394 output.n2 output.t1 3.9605
R20395 output.n4 output.t2 3.9605
R20396 output.n4 output.t7 3.9605
R20397 output.n6 output.t11 3.9605
R20398 output.n6 output.t3 3.9605
R20399 output.n8 output.t6 3.9605
R20400 output.n8 output.t4 3.9605
R20401 output.n10 output.t10 3.9605
R20402 output.n10 output.t13 3.9605
R20403 output.n12 output.t14 3.9605
R20404 output.n12 output.t8 3.9605
R20405 output.n38 output.n19 3.49141
R20406 output.n69 output.n50 3.49141
R20407 output.n101 output.n82 3.49141
R20408 output.n133 output.n114 3.49141
R20409 output.n35 output.n34 2.71565
R20410 output.n66 output.n65 2.71565
R20411 output.n98 output.n97 2.71565
R20412 output.n130 output.n129 2.71565
R20413 output.n31 output.n21 1.93989
R20414 output.n62 output.n52 1.93989
R20415 output.n94 output.n84 1.93989
R20416 output.n126 output.n116 1.93989
R20417 output.n30 output.n23 1.16414
R20418 output.n61 output.n54 1.16414
R20419 output.n93 output.n86 1.16414
R20420 output.n125 output.n118 1.16414
R20421 output.n141 output.n109 0.962709
R20422 output.n109 output.n77 0.962709
R20423 output.n27 output.n26 0.388379
R20424 output.n58 output.n57 0.388379
R20425 output.n90 output.n89 0.388379
R20426 output.n122 output.n121 0.388379
R20427 output.n14 output.n13 0.387128
R20428 output.n13 output.n11 0.387128
R20429 output.n11 output.n9 0.387128
R20430 output.n9 output.n7 0.387128
R20431 output.n7 output.n5 0.387128
R20432 output.n5 output.n3 0.387128
R20433 output.n3 output.n1 0.387128
R20434 output.n44 output.n16 0.155672
R20435 output.n37 output.n16 0.155672
R20436 output.n37 output.n36 0.155672
R20437 output.n36 output.n20 0.155672
R20438 output.n29 output.n20 0.155672
R20439 output.n29 output.n28 0.155672
R20440 output.n75 output.n47 0.155672
R20441 output.n68 output.n47 0.155672
R20442 output.n68 output.n67 0.155672
R20443 output.n67 output.n51 0.155672
R20444 output.n60 output.n51 0.155672
R20445 output.n60 output.n59 0.155672
R20446 output.n107 output.n79 0.155672
R20447 output.n100 output.n79 0.155672
R20448 output.n100 output.n99 0.155672
R20449 output.n99 output.n83 0.155672
R20450 output.n92 output.n83 0.155672
R20451 output.n92 output.n91 0.155672
R20452 output.n139 output.n111 0.155672
R20453 output.n132 output.n111 0.155672
R20454 output.n132 output.n131 0.155672
R20455 output.n131 output.n115 0.155672
R20456 output.n124 output.n115 0.155672
R20457 output.n124 output.n123 0.155672
R20458 output output.n14 0.126227
R20459 minus.n76 minus.t28 250.337
R20460 minus.n15 minus.t20 250.337
R20461 minus.n126 minus.t1 243.255
R20462 minus.n120 minus.t8 231.093
R20463 minus.n59 minus.t10 231.093
R20464 minus.n125 minus.n123 224.169
R20465 minus.n125 minus.n124 223.454
R20466 minus.n62 minus.t12 187.445
R20467 minus.n113 minus.t18 187.445
R20468 minus.n107 minus.t25 187.445
R20469 minus.n66 minus.t22 187.445
R20470 minus.n68 minus.t19 187.445
R20471 minus.n95 minus.t7 187.445
R20472 minus.n89 minus.t6 187.445
R20473 minus.n72 minus.t16 187.445
R20474 minus.n74 minus.t15 187.445
R20475 minus.n77 minus.t23 187.445
R20476 minus.n16 minus.t14 187.445
R20477 minus.n13 minus.t9 187.445
R20478 minus.n11 minus.t5 187.445
R20479 minus.n28 minus.t26 187.445
R20480 minus.n34 minus.t27 187.445
R20481 minus.n7 minus.t21 187.445
R20482 minus.n5 minus.t24 187.445
R20483 minus.n46 minus.t17 187.445
R20484 minus.n52 minus.t11 187.445
R20485 minus.n1 minus.t13 187.445
R20486 minus.n78 minus.n75 161.3
R20487 minus.n80 minus.n79 161.3
R20488 minus.n82 minus.n81 161.3
R20489 minus.n83 minus.n73 161.3
R20490 minus.n85 minus.n84 161.3
R20491 minus.n87 minus.n86 161.3
R20492 minus.n88 minus.n71 161.3
R20493 minus.n91 minus.n90 161.3
R20494 minus.n92 minus.n70 161.3
R20495 minus.n94 minus.n93 161.3
R20496 minus.n96 minus.n69 161.3
R20497 minus.n98 minus.n97 161.3
R20498 minus.n100 minus.n99 161.3
R20499 minus.n101 minus.n67 161.3
R20500 minus.n103 minus.n102 161.3
R20501 minus.n105 minus.n104 161.3
R20502 minus.n106 minus.n65 161.3
R20503 minus.n109 minus.n108 161.3
R20504 minus.n110 minus.n64 161.3
R20505 minus.n112 minus.n111 161.3
R20506 minus.n114 minus.n63 161.3
R20507 minus.n116 minus.n115 161.3
R20508 minus.n118 minus.n117 161.3
R20509 minus.n119 minus.n61 161.3
R20510 minus.n121 minus.n120 161.3
R20511 minus.n60 minus.n59 161.3
R20512 minus.n58 minus.n0 161.3
R20513 minus.n57 minus.n56 161.3
R20514 minus.n55 minus.n54 161.3
R20515 minus.n53 minus.n2 161.3
R20516 minus.n51 minus.n50 161.3
R20517 minus.n49 minus.n3 161.3
R20518 minus.n48 minus.n47 161.3
R20519 minus.n45 minus.n4 161.3
R20520 minus.n44 minus.n43 161.3
R20521 minus.n42 minus.n41 161.3
R20522 minus.n40 minus.n6 161.3
R20523 minus.n39 minus.n38 161.3
R20524 minus.n37 minus.n36 161.3
R20525 minus.n35 minus.n8 161.3
R20526 minus.n33 minus.n32 161.3
R20527 minus.n31 minus.n9 161.3
R20528 minus.n30 minus.n29 161.3
R20529 minus.n27 minus.n10 161.3
R20530 minus.n26 minus.n25 161.3
R20531 minus.n24 minus.n23 161.3
R20532 minus.n22 minus.n12 161.3
R20533 minus.n21 minus.n20 161.3
R20534 minus.n19 minus.n18 161.3
R20535 minus.n17 minus.n14 161.3
R20536 minus.n106 minus.n105 56.5617
R20537 minus.n97 minus.n96 56.5617
R20538 minus.n88 minus.n87 56.5617
R20539 minus.n27 minus.n26 56.5617
R20540 minus.n36 minus.n35 56.5617
R20541 minus.n45 minus.n44 56.5617
R20542 minus.n115 minus.n114 56.5617
R20543 minus.n79 minus.n78 56.5617
R20544 minus.n18 minus.n17 56.5617
R20545 minus.n54 minus.n53 56.5617
R20546 minus.n119 minus.n118 50.2647
R20547 minus.n58 minus.n57 50.2647
R20548 minus.n108 minus.n64 46.3896
R20549 minus.n84 minus.n83 46.3896
R20550 minus.n23 minus.n22 46.3896
R20551 minus.n47 minus.n3 46.3896
R20552 minus.n76 minus.n75 43.1929
R20553 minus.n15 minus.n14 43.1929
R20554 minus.n101 minus.n100 42.5146
R20555 minus.n94 minus.n70 42.5146
R20556 minus.n33 minus.n9 42.5146
R20557 minus.n40 minus.n39 42.5146
R20558 minus.n77 minus.n76 40.6041
R20559 minus.n16 minus.n15 40.6041
R20560 minus.n102 minus.n101 38.6395
R20561 minus.n90 minus.n70 38.6395
R20562 minus.n29 minus.n9 38.6395
R20563 minus.n41 minus.n40 38.6395
R20564 minus.n122 minus.n121 35.4191
R20565 minus.n112 minus.n64 34.7644
R20566 minus.n83 minus.n82 34.7644
R20567 minus.n22 minus.n21 34.7644
R20568 minus.n51 minus.n3 34.7644
R20569 minus.n114 minus.n113 21.8872
R20570 minus.n79 minus.n74 21.8872
R20571 minus.n18 minus.n13 21.8872
R20572 minus.n53 minus.n52 21.8872
R20573 minus.n105 minus.n66 19.9199
R20574 minus.n89 minus.n88 19.9199
R20575 minus.n28 minus.n27 19.9199
R20576 minus.n44 minus.n5 19.9199
R20577 minus.n124 minus.t0 19.8005
R20578 minus.n124 minus.t2 19.8005
R20579 minus.n123 minus.t4 19.8005
R20580 minus.n123 minus.t3 19.8005
R20581 minus.n97 minus.n68 17.9525
R20582 minus.n96 minus.n95 17.9525
R20583 minus.n35 minus.n34 17.9525
R20584 minus.n36 minus.n7 17.9525
R20585 minus.n107 minus.n106 15.9852
R20586 minus.n87 minus.n72 15.9852
R20587 minus.n26 minus.n11 15.9852
R20588 minus.n46 minus.n45 15.9852
R20589 minus.n115 minus.n62 14.0178
R20590 minus.n78 minus.n77 14.0178
R20591 minus.n17 minus.n16 14.0178
R20592 minus.n54 minus.n1 14.0178
R20593 minus.n122 minus.n60 12.1501
R20594 minus minus.n127 10.9162
R20595 minus.n118 minus.n62 10.575
R20596 minus.n57 minus.n1 10.575
R20597 minus.n120 minus.n119 9.49444
R20598 minus.n59 minus.n58 9.49444
R20599 minus.n108 minus.n107 8.60764
R20600 minus.n84 minus.n72 8.60764
R20601 minus.n23 minus.n11 8.60764
R20602 minus.n47 minus.n46 8.60764
R20603 minus.n100 minus.n68 6.6403
R20604 minus.n95 minus.n94 6.6403
R20605 minus.n34 minus.n33 6.6403
R20606 minus.n39 minus.n7 6.6403
R20607 minus.n127 minus.n126 4.80222
R20608 minus.n102 minus.n66 4.67295
R20609 minus.n90 minus.n89 4.67295
R20610 minus.n29 minus.n28 4.67295
R20611 minus.n41 minus.n5 4.67295
R20612 minus.n113 minus.n112 2.7056
R20613 minus.n82 minus.n74 2.7056
R20614 minus.n21 minus.n13 2.7056
R20615 minus.n52 minus.n51 2.7056
R20616 minus.n127 minus.n122 0.972091
R20617 minus.n126 minus.n125 0.716017
R20618 minus.n121 minus.n61 0.189894
R20619 minus.n117 minus.n61 0.189894
R20620 minus.n117 minus.n116 0.189894
R20621 minus.n116 minus.n63 0.189894
R20622 minus.n111 minus.n63 0.189894
R20623 minus.n111 minus.n110 0.189894
R20624 minus.n110 minus.n109 0.189894
R20625 minus.n109 minus.n65 0.189894
R20626 minus.n104 minus.n65 0.189894
R20627 minus.n104 minus.n103 0.189894
R20628 minus.n103 minus.n67 0.189894
R20629 minus.n99 minus.n67 0.189894
R20630 minus.n99 minus.n98 0.189894
R20631 minus.n98 minus.n69 0.189894
R20632 minus.n93 minus.n69 0.189894
R20633 minus.n93 minus.n92 0.189894
R20634 minus.n92 minus.n91 0.189894
R20635 minus.n91 minus.n71 0.189894
R20636 minus.n86 minus.n71 0.189894
R20637 minus.n86 minus.n85 0.189894
R20638 minus.n85 minus.n73 0.189894
R20639 minus.n81 minus.n73 0.189894
R20640 minus.n81 minus.n80 0.189894
R20641 minus.n80 minus.n75 0.189894
R20642 minus.n19 minus.n14 0.189894
R20643 minus.n20 minus.n19 0.189894
R20644 minus.n20 minus.n12 0.189894
R20645 minus.n24 minus.n12 0.189894
R20646 minus.n25 minus.n24 0.189894
R20647 minus.n25 minus.n10 0.189894
R20648 minus.n30 minus.n10 0.189894
R20649 minus.n31 minus.n30 0.189894
R20650 minus.n32 minus.n31 0.189894
R20651 minus.n32 minus.n8 0.189894
R20652 minus.n37 minus.n8 0.189894
R20653 minus.n38 minus.n37 0.189894
R20654 minus.n38 minus.n6 0.189894
R20655 minus.n42 minus.n6 0.189894
R20656 minus.n43 minus.n42 0.189894
R20657 minus.n43 minus.n4 0.189894
R20658 minus.n48 minus.n4 0.189894
R20659 minus.n49 minus.n48 0.189894
R20660 minus.n50 minus.n49 0.189894
R20661 minus.n50 minus.n2 0.189894
R20662 minus.n55 minus.n2 0.189894
R20663 minus.n56 minus.n55 0.189894
R20664 minus.n56 minus.n0 0.189894
R20665 minus.n60 minus.n0 0.189894
R20666 diffpairibias.n0 diffpairibias.t18 436.822
R20667 diffpairibias.n21 diffpairibias.t19 435.479
R20668 diffpairibias.n20 diffpairibias.t16 435.479
R20669 diffpairibias.n19 diffpairibias.t17 435.479
R20670 diffpairibias.n18 diffpairibias.t21 435.479
R20671 diffpairibias.n0 diffpairibias.t22 435.479
R20672 diffpairibias.n1 diffpairibias.t20 435.479
R20673 diffpairibias.n2 diffpairibias.t23 435.479
R20674 diffpairibias.n10 diffpairibias.t0 377.536
R20675 diffpairibias.n10 diffpairibias.t8 376.193
R20676 diffpairibias.n11 diffpairibias.t10 376.193
R20677 diffpairibias.n12 diffpairibias.t6 376.193
R20678 diffpairibias.n13 diffpairibias.t2 376.193
R20679 diffpairibias.n14 diffpairibias.t12 376.193
R20680 diffpairibias.n15 diffpairibias.t4 376.193
R20681 diffpairibias.n16 diffpairibias.t14 376.193
R20682 diffpairibias.n3 diffpairibias.t1 113.368
R20683 diffpairibias.n3 diffpairibias.t9 112.698
R20684 diffpairibias.n4 diffpairibias.t11 112.698
R20685 diffpairibias.n5 diffpairibias.t7 112.698
R20686 diffpairibias.n6 diffpairibias.t3 112.698
R20687 diffpairibias.n7 diffpairibias.t13 112.698
R20688 diffpairibias.n8 diffpairibias.t5 112.698
R20689 diffpairibias.n9 diffpairibias.t15 112.698
R20690 diffpairibias.n17 diffpairibias.n16 4.77242
R20691 diffpairibias.n17 diffpairibias.n9 4.30807
R20692 diffpairibias.n18 diffpairibias.n17 4.13945
R20693 diffpairibias.n16 diffpairibias.n15 1.34352
R20694 diffpairibias.n15 diffpairibias.n14 1.34352
R20695 diffpairibias.n14 diffpairibias.n13 1.34352
R20696 diffpairibias.n13 diffpairibias.n12 1.34352
R20697 diffpairibias.n12 diffpairibias.n11 1.34352
R20698 diffpairibias.n11 diffpairibias.n10 1.34352
R20699 diffpairibias.n2 diffpairibias.n1 1.34352
R20700 diffpairibias.n1 diffpairibias.n0 1.34352
R20701 diffpairibias.n19 diffpairibias.n18 1.34352
R20702 diffpairibias.n20 diffpairibias.n19 1.34352
R20703 diffpairibias.n21 diffpairibias.n20 1.34352
R20704 diffpairibias.n22 diffpairibias.n21 0.862419
R20705 diffpairibias diffpairibias.n22 0.684875
R20706 diffpairibias.n9 diffpairibias.n8 0.672012
R20707 diffpairibias.n8 diffpairibias.n7 0.672012
R20708 diffpairibias.n7 diffpairibias.n6 0.672012
R20709 diffpairibias.n6 diffpairibias.n5 0.672012
R20710 diffpairibias.n5 diffpairibias.n4 0.672012
R20711 diffpairibias.n4 diffpairibias.n3 0.672012
R20712 diffpairibias.n22 diffpairibias.n2 0.190907
C0 output outputibias 2.34152f
C1 vdd output 7.23429f
C2 CSoutput output 6.13571f
C3 CSoutput outputibias 0.032386f
C4 vdd CSoutput 67.66129f
C5 minus diffpairibias 5.39e-19
C6 commonsourceibias output 0.006808f
C7 CSoutput minus 2.25384f
C8 vdd plus 0.072837f
C9 commonsourceibias outputibias 0.003832f
C10 plus diffpairibias 4.4e-19
C11 vdd commonsourceibias 0.004218f
C12 CSoutput plus 0.874948f
C13 commonsourceibias diffpairibias 0.052851f
C14 CSoutput commonsourceibias 29.0223f
C15 minus plus 9.674179f
C16 minus commonsourceibias 0.515369f
C17 plus commonsourceibias 0.498793f
C18 diffpairibias gnd 48.95304f
C19 outputibias gnd 32.465668f
C20 output gnd 15.47879f
C21 commonsourceibias gnd 0.118072p
C22 plus gnd 37.554802f
C23 minus gnd 28.665808f
C24 CSoutput gnd 88.6703f
C25 vdd gnd 0.34557p
C26 diffpairibias.t18 gnd 0.087401f
C27 diffpairibias.t22 gnd 0.087239f
C28 diffpairibias.n0 gnd 0.102784f
C29 diffpairibias.t20 gnd 0.087239f
C30 diffpairibias.n1 gnd 0.050171f
C31 diffpairibias.t23 gnd 0.087239f
C32 diffpairibias.n2 gnd 0.039841f
C33 diffpairibias.t1 gnd 0.083757f
C34 diffpairibias.t9 gnd 0.083392f
C35 diffpairibias.n3 gnd 0.131682f
C36 diffpairibias.t11 gnd 0.083392f
C37 diffpairibias.n4 gnd 0.07027f
C38 diffpairibias.t7 gnd 0.083392f
C39 diffpairibias.n5 gnd 0.07027f
C40 diffpairibias.t3 gnd 0.083392f
C41 diffpairibias.n6 gnd 0.07027f
C42 diffpairibias.t13 gnd 0.083392f
C43 diffpairibias.n7 gnd 0.07027f
C44 diffpairibias.t5 gnd 0.083392f
C45 diffpairibias.n8 gnd 0.07027f
C46 diffpairibias.t15 gnd 0.083392f
C47 diffpairibias.n9 gnd 0.099771f
C48 diffpairibias.t0 gnd 0.08427f
C49 diffpairibias.t8 gnd 0.084123f
C50 diffpairibias.n10 gnd 0.091784f
C51 diffpairibias.t10 gnd 0.084123f
C52 diffpairibias.n11 gnd 0.050681f
C53 diffpairibias.t6 gnd 0.084123f
C54 diffpairibias.n12 gnd 0.050681f
C55 diffpairibias.t2 gnd 0.084123f
C56 diffpairibias.n13 gnd 0.050681f
C57 diffpairibias.t12 gnd 0.084123f
C58 diffpairibias.n14 gnd 0.050681f
C59 diffpairibias.t4 gnd 0.084123f
C60 diffpairibias.n15 gnd 0.050681f
C61 diffpairibias.t14 gnd 0.084123f
C62 diffpairibias.n16 gnd 0.059977f
C63 diffpairibias.n17 gnd 0.226448f
C64 diffpairibias.t21 gnd 0.087239f
C65 diffpairibias.n18 gnd 0.050181f
C66 diffpairibias.t17 gnd 0.087239f
C67 diffpairibias.n19 gnd 0.050171f
C68 diffpairibias.t16 gnd 0.087239f
C69 diffpairibias.n20 gnd 0.050171f
C70 diffpairibias.t19 gnd 0.087239f
C71 diffpairibias.n21 gnd 0.045859f
C72 diffpairibias.n22 gnd 0.046268f
C73 minus.n0 gnd 0.031832f
C74 minus.t13 gnd 0.535246f
C75 minus.n1 gnd 0.216477f
C76 minus.n2 gnd 0.031832f
C77 minus.t11 gnd 0.535246f
C78 minus.n3 gnd 0.027201f
C79 minus.n4 gnd 0.031832f
C80 minus.t17 gnd 0.535246f
C81 minus.t24 gnd 0.535246f
C82 minus.n5 gnd 0.216477f
C83 minus.n6 gnd 0.031832f
C84 minus.t21 gnd 0.535246f
C85 minus.n7 gnd 0.216477f
C86 minus.n8 gnd 0.031832f
C87 minus.t27 gnd 0.535246f
C88 minus.n9 gnd 0.025872f
C89 minus.n10 gnd 0.031832f
C90 minus.t26 gnd 0.535246f
C91 minus.t5 gnd 0.535246f
C92 minus.n11 gnd 0.216477f
C93 minus.n12 gnd 0.031832f
C94 minus.t9 gnd 0.535246f
C95 minus.n13 gnd 0.216477f
C96 minus.n14 gnd 0.135091f
C97 minus.t14 gnd 0.535246f
C98 minus.t20 gnd 0.59877f
C99 minus.n15 gnd 0.253084f
C100 minus.n16 gnd 0.247907f
C101 minus.n17 gnd 0.040787f
C102 minus.n18 gnd 0.036021f
C103 minus.n19 gnd 0.031832f
C104 minus.n20 gnd 0.031832f
C105 minus.n21 gnd 0.038039f
C106 minus.n22 gnd 0.027201f
C107 minus.n23 gnd 0.041457f
C108 minus.n24 gnd 0.031832f
C109 minus.n25 gnd 0.031832f
C110 minus.n26 gnd 0.039596f
C111 minus.n27 gnd 0.037213f
C112 minus.n28 gnd 0.216477f
C113 minus.n29 gnd 0.039874f
C114 minus.n30 gnd 0.031832f
C115 minus.n31 gnd 0.031832f
C116 minus.n32 gnd 0.031832f
C117 minus.n33 gnd 0.04095f
C118 minus.n34 gnd 0.216477f
C119 minus.n35 gnd 0.038404f
C120 minus.n36 gnd 0.038404f
C121 minus.n37 gnd 0.031832f
C122 minus.n38 gnd 0.031832f
C123 minus.n39 gnd 0.04095f
C124 minus.n40 gnd 0.025872f
C125 minus.n41 gnd 0.039874f
C126 minus.n42 gnd 0.031832f
C127 minus.n43 gnd 0.031832f
C128 minus.n44 gnd 0.037213f
C129 minus.n45 gnd 0.039596f
C130 minus.n46 gnd 0.216477f
C131 minus.n47 gnd 0.041457f
C132 minus.n48 gnd 0.031832f
C133 minus.n49 gnd 0.031832f
C134 minus.n50 gnd 0.031832f
C135 minus.n51 gnd 0.038039f
C136 minus.n52 gnd 0.216477f
C137 minus.n53 gnd 0.036021f
C138 minus.n54 gnd 0.040787f
C139 minus.n55 gnd 0.031832f
C140 minus.n56 gnd 0.031832f
C141 minus.n57 gnd 0.041526f
C142 minus.n58 gnd 0.011569f
C143 minus.t10 gnd 0.578869f
C144 minus.n59 gnd 0.250644f
C145 minus.n60 gnd 0.372897f
C146 minus.n61 gnd 0.031832f
C147 minus.t8 gnd 0.578869f
C148 minus.t12 gnd 0.535246f
C149 minus.n62 gnd 0.216477f
C150 minus.n63 gnd 0.031832f
C151 minus.t18 gnd 0.535246f
C152 minus.n64 gnd 0.027201f
C153 minus.n65 gnd 0.031832f
C154 minus.t25 gnd 0.535246f
C155 minus.t22 gnd 0.535246f
C156 minus.n66 gnd 0.216477f
C157 minus.n67 gnd 0.031832f
C158 minus.t19 gnd 0.535246f
C159 minus.n68 gnd 0.216477f
C160 minus.n69 gnd 0.031832f
C161 minus.t7 gnd 0.535246f
C162 minus.n70 gnd 0.025872f
C163 minus.n71 gnd 0.031832f
C164 minus.t6 gnd 0.535246f
C165 minus.t16 gnd 0.535246f
C166 minus.n72 gnd 0.216477f
C167 minus.n73 gnd 0.031832f
C168 minus.t15 gnd 0.535246f
C169 minus.n74 gnd 0.216477f
C170 minus.n75 gnd 0.135091f
C171 minus.t23 gnd 0.535246f
C172 minus.t28 gnd 0.59877f
C173 minus.n76 gnd 0.253084f
C174 minus.n77 gnd 0.247907f
C175 minus.n78 gnd 0.040787f
C176 minus.n79 gnd 0.036021f
C177 minus.n80 gnd 0.031832f
C178 minus.n81 gnd 0.031832f
C179 minus.n82 gnd 0.038039f
C180 minus.n83 gnd 0.027201f
C181 minus.n84 gnd 0.041457f
C182 minus.n85 gnd 0.031832f
C183 minus.n86 gnd 0.031832f
C184 minus.n87 gnd 0.039596f
C185 minus.n88 gnd 0.037213f
C186 minus.n89 gnd 0.216477f
C187 minus.n90 gnd 0.039874f
C188 minus.n91 gnd 0.031832f
C189 minus.n92 gnd 0.031832f
C190 minus.n93 gnd 0.031832f
C191 minus.n94 gnd 0.04095f
C192 minus.n95 gnd 0.216477f
C193 minus.n96 gnd 0.038404f
C194 minus.n97 gnd 0.038404f
C195 minus.n98 gnd 0.031832f
C196 minus.n99 gnd 0.031832f
C197 minus.n100 gnd 0.04095f
C198 minus.n101 gnd 0.025872f
C199 minus.n102 gnd 0.039874f
C200 minus.n103 gnd 0.031832f
C201 minus.n104 gnd 0.031832f
C202 minus.n105 gnd 0.037213f
C203 minus.n106 gnd 0.039596f
C204 minus.n107 gnd 0.216477f
C205 minus.n108 gnd 0.041457f
C206 minus.n109 gnd 0.031832f
C207 minus.n110 gnd 0.031832f
C208 minus.n111 gnd 0.031832f
C209 minus.n112 gnd 0.038039f
C210 minus.n113 gnd 0.216477f
C211 minus.n114 gnd 0.036021f
C212 minus.n115 gnd 0.040787f
C213 minus.n116 gnd 0.031832f
C214 minus.n117 gnd 0.031832f
C215 minus.n118 gnd 0.041526f
C216 minus.n119 gnd 0.011569f
C217 minus.n120 gnd 0.250644f
C218 minus.n121 gnd 1.16121f
C219 minus.n122 gnd 1.70573f
C220 minus.t4 gnd 0.009813f
C221 minus.t3 gnd 0.009813f
C222 minus.n123 gnd 0.032267f
C223 minus.t0 gnd 0.009813f
C224 minus.t2 gnd 0.009813f
C225 minus.n124 gnd 0.031825f
C226 minus.n125 gnd 0.271609f
C227 minus.t1 gnd 0.054617f
C228 minus.n126 gnd 0.148215f
C229 minus.n127 gnd 1.6183f
C230 output.t15 gnd 0.464308f
C231 output.t5 gnd 0.044422f
C232 output.t9 gnd 0.044422f
C233 output.n0 gnd 0.364624f
C234 output.n1 gnd 0.614102f
C235 output.t12 gnd 0.044422f
C236 output.t1 gnd 0.044422f
C237 output.n2 gnd 0.364624f
C238 output.n3 gnd 0.350265f
C239 output.t2 gnd 0.044422f
C240 output.t7 gnd 0.044422f
C241 output.n4 gnd 0.364624f
C242 output.n5 gnd 0.350265f
C243 output.t11 gnd 0.044422f
C244 output.t3 gnd 0.044422f
C245 output.n6 gnd 0.364624f
C246 output.n7 gnd 0.350265f
C247 output.t6 gnd 0.044422f
C248 output.t4 gnd 0.044422f
C249 output.n8 gnd 0.364624f
C250 output.n9 gnd 0.350265f
C251 output.t10 gnd 0.044422f
C252 output.t13 gnd 0.044422f
C253 output.n10 gnd 0.364624f
C254 output.n11 gnd 0.350265f
C255 output.t14 gnd 0.044422f
C256 output.t8 gnd 0.044422f
C257 output.n12 gnd 0.364624f
C258 output.n13 gnd 0.350265f
C259 output.t0 gnd 0.462979f
C260 output.n14 gnd 0.28994f
C261 output.n15 gnd 0.015803f
C262 output.n16 gnd 0.011243f
C263 output.n17 gnd 0.006041f
C264 output.n18 gnd 0.01428f
C265 output.n19 gnd 0.006397f
C266 output.n20 gnd 0.011243f
C267 output.n21 gnd 0.006041f
C268 output.n22 gnd 0.01428f
C269 output.n23 gnd 0.006397f
C270 output.n24 gnd 0.048111f
C271 output.t19 gnd 0.023274f
C272 output.n25 gnd 0.01071f
C273 output.n26 gnd 0.008435f
C274 output.n27 gnd 0.006041f
C275 output.n28 gnd 0.267512f
C276 output.n29 gnd 0.011243f
C277 output.n30 gnd 0.006041f
C278 output.n31 gnd 0.006397f
C279 output.n32 gnd 0.01428f
C280 output.n33 gnd 0.01428f
C281 output.n34 gnd 0.006397f
C282 output.n35 gnd 0.006041f
C283 output.n36 gnd 0.011243f
C284 output.n37 gnd 0.011243f
C285 output.n38 gnd 0.006041f
C286 output.n39 gnd 0.006397f
C287 output.n40 gnd 0.01428f
C288 output.n41 gnd 0.030913f
C289 output.n42 gnd 0.006397f
C290 output.n43 gnd 0.006041f
C291 output.n44 gnd 0.025987f
C292 output.n45 gnd 0.097665f
C293 output.n46 gnd 0.015803f
C294 output.n47 gnd 0.011243f
C295 output.n48 gnd 0.006041f
C296 output.n49 gnd 0.01428f
C297 output.n50 gnd 0.006397f
C298 output.n51 gnd 0.011243f
C299 output.n52 gnd 0.006041f
C300 output.n53 gnd 0.01428f
C301 output.n54 gnd 0.006397f
C302 output.n55 gnd 0.048111f
C303 output.t18 gnd 0.023274f
C304 output.n56 gnd 0.01071f
C305 output.n57 gnd 0.008435f
C306 output.n58 gnd 0.006041f
C307 output.n59 gnd 0.267512f
C308 output.n60 gnd 0.011243f
C309 output.n61 gnd 0.006041f
C310 output.n62 gnd 0.006397f
C311 output.n63 gnd 0.01428f
C312 output.n64 gnd 0.01428f
C313 output.n65 gnd 0.006397f
C314 output.n66 gnd 0.006041f
C315 output.n67 gnd 0.011243f
C316 output.n68 gnd 0.011243f
C317 output.n69 gnd 0.006041f
C318 output.n70 gnd 0.006397f
C319 output.n71 gnd 0.01428f
C320 output.n72 gnd 0.030913f
C321 output.n73 gnd 0.006397f
C322 output.n74 gnd 0.006041f
C323 output.n75 gnd 0.025987f
C324 output.n76 gnd 0.09306f
C325 output.n77 gnd 1.65264f
C326 output.n78 gnd 0.015803f
C327 output.n79 gnd 0.011243f
C328 output.n80 gnd 0.006041f
C329 output.n81 gnd 0.01428f
C330 output.n82 gnd 0.006397f
C331 output.n83 gnd 0.011243f
C332 output.n84 gnd 0.006041f
C333 output.n85 gnd 0.01428f
C334 output.n86 gnd 0.006397f
C335 output.n87 gnd 0.048111f
C336 output.t17 gnd 0.023274f
C337 output.n88 gnd 0.01071f
C338 output.n89 gnd 0.008435f
C339 output.n90 gnd 0.006041f
C340 output.n91 gnd 0.267512f
C341 output.n92 gnd 0.011243f
C342 output.n93 gnd 0.006041f
C343 output.n94 gnd 0.006397f
C344 output.n95 gnd 0.01428f
C345 output.n96 gnd 0.01428f
C346 output.n97 gnd 0.006397f
C347 output.n98 gnd 0.006041f
C348 output.n99 gnd 0.011243f
C349 output.n100 gnd 0.011243f
C350 output.n101 gnd 0.006041f
C351 output.n102 gnd 0.006397f
C352 output.n103 gnd 0.01428f
C353 output.n104 gnd 0.030913f
C354 output.n105 gnd 0.006397f
C355 output.n106 gnd 0.006041f
C356 output.n107 gnd 0.025987f
C357 output.n108 gnd 0.09306f
C358 output.n109 gnd 0.713089f
C359 output.n110 gnd 0.015803f
C360 output.n111 gnd 0.011243f
C361 output.n112 gnd 0.006041f
C362 output.n113 gnd 0.01428f
C363 output.n114 gnd 0.006397f
C364 output.n115 gnd 0.011243f
C365 output.n116 gnd 0.006041f
C366 output.n117 gnd 0.01428f
C367 output.n118 gnd 0.006397f
C368 output.n119 gnd 0.048111f
C369 output.t16 gnd 0.023274f
C370 output.n120 gnd 0.01071f
C371 output.n121 gnd 0.008435f
C372 output.n122 gnd 0.006041f
C373 output.n123 gnd 0.267512f
C374 output.n124 gnd 0.011243f
C375 output.n125 gnd 0.006041f
C376 output.n126 gnd 0.006397f
C377 output.n127 gnd 0.01428f
C378 output.n128 gnd 0.01428f
C379 output.n129 gnd 0.006397f
C380 output.n130 gnd 0.006041f
C381 output.n131 gnd 0.011243f
C382 output.n132 gnd 0.011243f
C383 output.n133 gnd 0.006041f
C384 output.n134 gnd 0.006397f
C385 output.n135 gnd 0.01428f
C386 output.n136 gnd 0.030913f
C387 output.n137 gnd 0.006397f
C388 output.n138 gnd 0.006041f
C389 output.n139 gnd 0.025987f
C390 output.n140 gnd 0.09306f
C391 output.n141 gnd 1.67353f
C392 outputibias.t9 gnd 0.11477f
C393 outputibias.t8 gnd 0.115567f
C394 outputibias.n0 gnd 0.130108f
C395 outputibias.n1 gnd 0.001372f
C396 outputibias.n2 gnd 9.76e-19
C397 outputibias.n3 gnd 5.24e-19
C398 outputibias.n4 gnd 0.001239f
C399 outputibias.n5 gnd 5.55e-19
C400 outputibias.n6 gnd 9.76e-19
C401 outputibias.n7 gnd 5.24e-19
C402 outputibias.n8 gnd 0.001239f
C403 outputibias.n9 gnd 5.55e-19
C404 outputibias.n10 gnd 0.004176f
C405 outputibias.t5 gnd 0.00202f
C406 outputibias.n11 gnd 9.3e-19
C407 outputibias.n12 gnd 7.32e-19
C408 outputibias.n13 gnd 5.24e-19
C409 outputibias.n14 gnd 0.02322f
C410 outputibias.n15 gnd 9.76e-19
C411 outputibias.n16 gnd 5.24e-19
C412 outputibias.n17 gnd 5.55e-19
C413 outputibias.n18 gnd 0.001239f
C414 outputibias.n19 gnd 0.001239f
C415 outputibias.n20 gnd 5.55e-19
C416 outputibias.n21 gnd 5.24e-19
C417 outputibias.n22 gnd 9.76e-19
C418 outputibias.n23 gnd 9.76e-19
C419 outputibias.n24 gnd 5.24e-19
C420 outputibias.n25 gnd 5.55e-19
C421 outputibias.n26 gnd 0.001239f
C422 outputibias.n27 gnd 0.002683f
C423 outputibias.n28 gnd 5.55e-19
C424 outputibias.n29 gnd 5.24e-19
C425 outputibias.n30 gnd 0.002256f
C426 outputibias.n31 gnd 0.005781f
C427 outputibias.n32 gnd 0.001372f
C428 outputibias.n33 gnd 9.76e-19
C429 outputibias.n34 gnd 5.24e-19
C430 outputibias.n35 gnd 0.001239f
C431 outputibias.n36 gnd 5.55e-19
C432 outputibias.n37 gnd 9.76e-19
C433 outputibias.n38 gnd 5.24e-19
C434 outputibias.n39 gnd 0.001239f
C435 outputibias.n40 gnd 5.55e-19
C436 outputibias.n41 gnd 0.004176f
C437 outputibias.t7 gnd 0.00202f
C438 outputibias.n42 gnd 9.3e-19
C439 outputibias.n43 gnd 7.32e-19
C440 outputibias.n44 gnd 5.24e-19
C441 outputibias.n45 gnd 0.02322f
C442 outputibias.n46 gnd 9.76e-19
C443 outputibias.n47 gnd 5.24e-19
C444 outputibias.n48 gnd 5.55e-19
C445 outputibias.n49 gnd 0.001239f
C446 outputibias.n50 gnd 0.001239f
C447 outputibias.n51 gnd 5.55e-19
C448 outputibias.n52 gnd 5.24e-19
C449 outputibias.n53 gnd 9.76e-19
C450 outputibias.n54 gnd 9.76e-19
C451 outputibias.n55 gnd 5.24e-19
C452 outputibias.n56 gnd 5.55e-19
C453 outputibias.n57 gnd 0.001239f
C454 outputibias.n58 gnd 0.002683f
C455 outputibias.n59 gnd 5.55e-19
C456 outputibias.n60 gnd 5.24e-19
C457 outputibias.n61 gnd 0.002256f
C458 outputibias.n62 gnd 0.005197f
C459 outputibias.n63 gnd 0.121892f
C460 outputibias.n64 gnd 0.001372f
C461 outputibias.n65 gnd 9.76e-19
C462 outputibias.n66 gnd 5.24e-19
C463 outputibias.n67 gnd 0.001239f
C464 outputibias.n68 gnd 5.55e-19
C465 outputibias.n69 gnd 9.76e-19
C466 outputibias.n70 gnd 5.24e-19
C467 outputibias.n71 gnd 0.001239f
C468 outputibias.n72 gnd 5.55e-19
C469 outputibias.n73 gnd 0.004176f
C470 outputibias.t1 gnd 0.00202f
C471 outputibias.n74 gnd 9.3e-19
C472 outputibias.n75 gnd 7.32e-19
C473 outputibias.n76 gnd 5.24e-19
C474 outputibias.n77 gnd 0.02322f
C475 outputibias.n78 gnd 9.76e-19
C476 outputibias.n79 gnd 5.24e-19
C477 outputibias.n80 gnd 5.55e-19
C478 outputibias.n81 gnd 0.001239f
C479 outputibias.n82 gnd 0.001239f
C480 outputibias.n83 gnd 5.55e-19
C481 outputibias.n84 gnd 5.24e-19
C482 outputibias.n85 gnd 9.76e-19
C483 outputibias.n86 gnd 9.76e-19
C484 outputibias.n87 gnd 5.24e-19
C485 outputibias.n88 gnd 5.55e-19
C486 outputibias.n89 gnd 0.001239f
C487 outputibias.n90 gnd 0.002683f
C488 outputibias.n91 gnd 5.55e-19
C489 outputibias.n92 gnd 5.24e-19
C490 outputibias.n93 gnd 0.002256f
C491 outputibias.n94 gnd 0.005197f
C492 outputibias.n95 gnd 0.064513f
C493 outputibias.n96 gnd 0.001372f
C494 outputibias.n97 gnd 9.76e-19
C495 outputibias.n98 gnd 5.24e-19
C496 outputibias.n99 gnd 0.001239f
C497 outputibias.n100 gnd 5.55e-19
C498 outputibias.n101 gnd 9.76e-19
C499 outputibias.n102 gnd 5.24e-19
C500 outputibias.n103 gnd 0.001239f
C501 outputibias.n104 gnd 5.55e-19
C502 outputibias.n105 gnd 0.004176f
C503 outputibias.t3 gnd 0.00202f
C504 outputibias.n106 gnd 9.3e-19
C505 outputibias.n107 gnd 7.32e-19
C506 outputibias.n108 gnd 5.24e-19
C507 outputibias.n109 gnd 0.02322f
C508 outputibias.n110 gnd 9.76e-19
C509 outputibias.n111 gnd 5.24e-19
C510 outputibias.n112 gnd 5.55e-19
C511 outputibias.n113 gnd 0.001239f
C512 outputibias.n114 gnd 0.001239f
C513 outputibias.n115 gnd 5.55e-19
C514 outputibias.n116 gnd 5.24e-19
C515 outputibias.n117 gnd 9.76e-19
C516 outputibias.n118 gnd 9.76e-19
C517 outputibias.n119 gnd 5.24e-19
C518 outputibias.n120 gnd 5.55e-19
C519 outputibias.n121 gnd 0.001239f
C520 outputibias.n122 gnd 0.002683f
C521 outputibias.n123 gnd 5.55e-19
C522 outputibias.n124 gnd 5.24e-19
C523 outputibias.n125 gnd 0.002256f
C524 outputibias.n126 gnd 0.005197f
C525 outputibias.n127 gnd 0.084814f
C526 outputibias.t2 gnd 0.108319f
C527 outputibias.t0 gnd 0.108319f
C528 outputibias.t6 gnd 0.108319f
C529 outputibias.t4 gnd 0.109238f
C530 outputibias.n128 gnd 0.134674f
C531 outputibias.n129 gnd 0.07244f
C532 outputibias.n130 gnd 0.079818f
C533 outputibias.n131 gnd 0.164901f
C534 outputibias.t11 gnd 0.11477f
C535 outputibias.n132 gnd 0.067481f
C536 outputibias.t10 gnd 0.11477f
C537 outputibias.n133 gnd 0.065115f
C538 outputibias.n134 gnd 0.029159f
C539 a_n3106_n452.t23 gnd 0.10001f
C540 a_n3106_n452.t34 gnd 1.03942f
C541 a_n3106_n452.n0 gnd 0.392946f
C542 a_n3106_n452.t10 gnd 1.29145f
C543 a_n3106_n452.n1 gnd 1.22854f
C544 a_n3106_n452.t53 gnd 1.03942f
C545 a_n3106_n452.n2 gnd 0.392946f
C546 a_n3106_n452.t0 gnd 0.10001f
C547 a_n3106_n452.t5 gnd 0.10001f
C548 a_n3106_n452.n3 gnd 0.816794f
C549 a_n3106_n452.n4 gnd 0.411618f
C550 a_n3106_n452.t7 gnd 0.10001f
C551 a_n3106_n452.t44 gnd 0.10001f
C552 a_n3106_n452.n5 gnd 0.816794f
C553 a_n3106_n452.n6 gnd 0.411618f
C554 a_n3106_n452.t43 gnd 0.10001f
C555 a_n3106_n452.t2 gnd 0.10001f
C556 a_n3106_n452.n7 gnd 0.816794f
C557 a_n3106_n452.n8 gnd 0.411618f
C558 a_n3106_n452.t51 gnd 0.10001f
C559 a_n3106_n452.t12 gnd 0.10001f
C560 a_n3106_n452.n9 gnd 0.816794f
C561 a_n3106_n452.n10 gnd 0.411618f
C562 a_n3106_n452.t50 gnd 0.10001f
C563 a_n3106_n452.t13 gnd 0.10001f
C564 a_n3106_n452.n11 gnd 0.816794f
C565 a_n3106_n452.n12 gnd 0.411618f
C566 a_n3106_n452.t4 gnd 1.03942f
C567 a_n3106_n452.n13 gnd 0.972974f
C568 a_n3106_n452.t9 gnd 1.29145f
C569 a_n3106_n452.n14 gnd 0.909591f
C570 a_n3106_n452.t49 gnd 1.29145f
C571 a_n3106_n452.n15 gnd 0.909591f
C572 a_n3106_n452.t48 gnd 1.29145f
C573 a_n3106_n452.n16 gnd 0.909591f
C574 a_n3106_n452.t41 gnd 1.29145f
C575 a_n3106_n452.n17 gnd 0.909591f
C576 a_n3106_n452.t11 gnd 1.29145f
C577 a_n3106_n452.n18 gnd 0.909591f
C578 a_n3106_n452.t16 gnd 1.29145f
C579 a_n3106_n452.n19 gnd 0.909591f
C580 a_n3106_n452.t15 gnd 1.29145f
C581 a_n3106_n452.n20 gnd 0.789472f
C582 a_n3106_n452.n21 gnd 0.948419f
C583 a_n3106_n452.t25 gnd 1.03941f
C584 a_n3106_n452.n22 gnd 0.645631f
C585 a_n3106_n452.t22 gnd 0.10001f
C586 a_n3106_n452.t39 gnd 0.10001f
C587 a_n3106_n452.n23 gnd 0.816793f
C588 a_n3106_n452.n24 gnd 0.41162f
C589 a_n3106_n452.t33 gnd 0.10001f
C590 a_n3106_n452.t37 gnd 0.10001f
C591 a_n3106_n452.n25 gnd 0.816793f
C592 a_n3106_n452.n26 gnd 0.41162f
C593 a_n3106_n452.t38 gnd 0.10001f
C594 a_n3106_n452.t26 gnd 0.10001f
C595 a_n3106_n452.n27 gnd 0.816793f
C596 a_n3106_n452.n28 gnd 0.41162f
C597 a_n3106_n452.t27 gnd 0.10001f
C598 a_n3106_n452.t18 gnd 0.10001f
C599 a_n3106_n452.n29 gnd 0.816793f
C600 a_n3106_n452.n30 gnd 0.41162f
C601 a_n3106_n452.t20 gnd 0.10001f
C602 a_n3106_n452.t36 gnd 0.10001f
C603 a_n3106_n452.n31 gnd 0.816793f
C604 a_n3106_n452.n32 gnd 0.41162f
C605 a_n3106_n452.t31 gnd 1.03941f
C606 a_n3106_n452.n33 gnd 0.39295f
C607 a_n3106_n452.t14 gnd 1.03941f
C608 a_n3106_n452.n34 gnd 0.39295f
C609 a_n3106_n452.t42 gnd 0.10001f
C610 a_n3106_n452.t1 gnd 0.10001f
C611 a_n3106_n452.n35 gnd 0.816793f
C612 a_n3106_n452.n36 gnd 0.41162f
C613 a_n3106_n452.t8 gnd 0.10001f
C614 a_n3106_n452.t54 gnd 0.10001f
C615 a_n3106_n452.n37 gnd 0.816793f
C616 a_n3106_n452.n38 gnd 0.41162f
C617 a_n3106_n452.t55 gnd 0.10001f
C618 a_n3106_n452.t46 gnd 0.10001f
C619 a_n3106_n452.n39 gnd 0.816793f
C620 a_n3106_n452.n40 gnd 0.41162f
C621 a_n3106_n452.t6 gnd 0.10001f
C622 a_n3106_n452.t45 gnd 0.10001f
C623 a_n3106_n452.n41 gnd 0.816793f
C624 a_n3106_n452.n42 gnd 0.41162f
C625 a_n3106_n452.t3 gnd 0.10001f
C626 a_n3106_n452.t47 gnd 0.10001f
C627 a_n3106_n452.n43 gnd 0.816793f
C628 a_n3106_n452.n44 gnd 0.41162f
C629 a_n3106_n452.t52 gnd 1.03941f
C630 a_n3106_n452.n45 gnd 0.645631f
C631 a_n3106_n452.n46 gnd 1.05146f
C632 a_n3106_n452.t21 gnd 1.03941f
C633 a_n3106_n452.n47 gnd 0.972978f
C634 a_n3106_n452.t19 gnd 0.10001f
C635 a_n3106_n452.t17 gnd 0.10001f
C636 a_n3106_n452.n48 gnd 0.816794f
C637 a_n3106_n452.n49 gnd 0.411618f
C638 a_n3106_n452.t30 gnd 0.10001f
C639 a_n3106_n452.t35 gnd 0.10001f
C640 a_n3106_n452.n50 gnd 0.816794f
C641 a_n3106_n452.n51 gnd 0.411618f
C642 a_n3106_n452.t28 gnd 0.10001f
C643 a_n3106_n452.t32 gnd 0.10001f
C644 a_n3106_n452.n52 gnd 0.816794f
C645 a_n3106_n452.n53 gnd 0.411618f
C646 a_n3106_n452.t24 gnd 0.10001f
C647 a_n3106_n452.t29 gnd 0.10001f
C648 a_n3106_n452.n54 gnd 0.816794f
C649 a_n3106_n452.n55 gnd 0.411618f
C650 a_n3106_n452.n56 gnd 0.411617f
C651 a_n3106_n452.n57 gnd 0.816796f
C652 a_n3106_n452.t40 gnd 0.10001f
C653 plus.n0 gnd 0.023652f
C654 plus.t20 gnd 0.430126f
C655 plus.t23 gnd 0.397712f
C656 plus.n1 gnd 0.160852f
C657 plus.n2 gnd 0.023652f
C658 plus.t6 gnd 0.397712f
C659 plus.n3 gnd 0.020211f
C660 plus.n4 gnd 0.023652f
C661 plus.t12 gnd 0.397712f
C662 plus.t8 gnd 0.397712f
C663 plus.n5 gnd 0.160852f
C664 plus.n6 gnd 0.023652f
C665 plus.t7 gnd 0.397712f
C666 plus.n7 gnd 0.160852f
C667 plus.n8 gnd 0.023652f
C668 plus.t19 gnd 0.397712f
C669 plus.n9 gnd 0.019224f
C670 plus.n10 gnd 0.023652f
C671 plus.t18 gnd 0.397712f
C672 plus.t27 gnd 0.397712f
C673 plus.n11 gnd 0.160852f
C674 plus.n12 gnd 0.023652f
C675 plus.t25 gnd 0.397712f
C676 plus.n13 gnd 0.160852f
C677 plus.n14 gnd 0.100378f
C678 plus.t9 gnd 0.397712f
C679 plus.t14 gnd 0.444913f
C680 plus.n15 gnd 0.188053f
C681 plus.n16 gnd 0.184206f
C682 plus.n17 gnd 0.030307f
C683 plus.n18 gnd 0.026765f
C684 plus.n19 gnd 0.023652f
C685 plus.n20 gnd 0.023652f
C686 plus.n21 gnd 0.028265f
C687 plus.n22 gnd 0.020211f
C688 plus.n23 gnd 0.030804f
C689 plus.n24 gnd 0.023652f
C690 plus.n25 gnd 0.023652f
C691 plus.n26 gnd 0.029422f
C692 plus.n27 gnd 0.027651f
C693 plus.n28 gnd 0.160852f
C694 plus.n29 gnd 0.029629f
C695 plus.n30 gnd 0.023652f
C696 plus.n31 gnd 0.023652f
C697 plus.n32 gnd 0.023652f
C698 plus.n33 gnd 0.030428f
C699 plus.n34 gnd 0.160852f
C700 plus.n35 gnd 0.028536f
C701 plus.n36 gnd 0.028536f
C702 plus.n37 gnd 0.023652f
C703 plus.n38 gnd 0.023652f
C704 plus.n39 gnd 0.030428f
C705 plus.n40 gnd 0.019224f
C706 plus.n41 gnd 0.029629f
C707 plus.n42 gnd 0.023652f
C708 plus.n43 gnd 0.023652f
C709 plus.n44 gnd 0.027651f
C710 plus.n45 gnd 0.029422f
C711 plus.n46 gnd 0.160852f
C712 plus.n47 gnd 0.030804f
C713 plus.n48 gnd 0.023652f
C714 plus.n49 gnd 0.023652f
C715 plus.n50 gnd 0.023652f
C716 plus.n51 gnd 0.028265f
C717 plus.n52 gnd 0.160852f
C718 plus.n53 gnd 0.026765f
C719 plus.n54 gnd 0.030307f
C720 plus.n55 gnd 0.023652f
C721 plus.n56 gnd 0.023652f
C722 plus.n57 gnd 0.030855f
C723 plus.n58 gnd 0.008596f
C724 plus.n59 gnd 0.18624f
C725 plus.n60 gnd 0.270994f
C726 plus.n61 gnd 0.023652f
C727 plus.t28 gnd 0.397712f
C728 plus.n62 gnd 0.160852f
C729 plus.n63 gnd 0.023652f
C730 plus.t26 gnd 0.397712f
C731 plus.n64 gnd 0.020211f
C732 plus.n65 gnd 0.023652f
C733 plus.t10 gnd 0.397712f
C734 plus.t15 gnd 0.397712f
C735 plus.n66 gnd 0.160852f
C736 plus.n67 gnd 0.023652f
C737 plus.t13 gnd 0.397712f
C738 plus.n68 gnd 0.160852f
C739 plus.n69 gnd 0.023652f
C740 plus.t17 gnd 0.397712f
C741 plus.n70 gnd 0.019224f
C742 plus.n71 gnd 0.023652f
C743 plus.t16 gnd 0.397712f
C744 plus.t21 gnd 0.397712f
C745 plus.n72 gnd 0.160852f
C746 plus.n73 gnd 0.023652f
C747 plus.t22 gnd 0.397712f
C748 plus.n74 gnd 0.160852f
C749 plus.n75 gnd 0.100378f
C750 plus.t5 gnd 0.397712f
C751 plus.t11 gnd 0.444913f
C752 plus.n76 gnd 0.188053f
C753 plus.n77 gnd 0.184206f
C754 plus.n78 gnd 0.030307f
C755 plus.n79 gnd 0.026765f
C756 plus.n80 gnd 0.023652f
C757 plus.n81 gnd 0.023652f
C758 plus.n82 gnd 0.028265f
C759 plus.n83 gnd 0.020211f
C760 plus.n84 gnd 0.030804f
C761 plus.n85 gnd 0.023652f
C762 plus.n86 gnd 0.023652f
C763 plus.n87 gnd 0.029422f
C764 plus.n88 gnd 0.027651f
C765 plus.n89 gnd 0.160852f
C766 plus.n90 gnd 0.029629f
C767 plus.n91 gnd 0.023652f
C768 plus.n92 gnd 0.023652f
C769 plus.n93 gnd 0.023652f
C770 plus.n94 gnd 0.030428f
C771 plus.n95 gnd 0.160852f
C772 plus.n96 gnd 0.028536f
C773 plus.n97 gnd 0.028536f
C774 plus.n98 gnd 0.023652f
C775 plus.n99 gnd 0.023652f
C776 plus.n100 gnd 0.030428f
C777 plus.n101 gnd 0.019224f
C778 plus.n102 gnd 0.029629f
C779 plus.n103 gnd 0.023652f
C780 plus.n104 gnd 0.023652f
C781 plus.n105 gnd 0.027651f
C782 plus.n106 gnd 0.029422f
C783 plus.n107 gnd 0.160852f
C784 plus.n108 gnd 0.030804f
C785 plus.n109 gnd 0.023652f
C786 plus.n110 gnd 0.023652f
C787 plus.n111 gnd 0.023652f
C788 plus.n112 gnd 0.028265f
C789 plus.n113 gnd 0.160852f
C790 plus.n114 gnd 0.026765f
C791 plus.n115 gnd 0.030307f
C792 plus.n116 gnd 0.023652f
C793 plus.n117 gnd 0.023652f
C794 plus.n118 gnd 0.030855f
C795 plus.n119 gnd 0.008596f
C796 plus.t24 gnd 0.430126f
C797 plus.n120 gnd 0.18624f
C798 plus.n121 gnd 0.853371f
C799 plus.n122 gnd 1.25804f
C800 plus.t1 gnd 0.040831f
C801 plus.t2 gnd 0.007291f
C802 plus.t4 gnd 0.007291f
C803 plus.n123 gnd 0.023647f
C804 plus.n124 gnd 0.183575f
C805 plus.t3 gnd 0.007291f
C806 plus.t0 gnd 0.007291f
C807 plus.n125 gnd 0.023647f
C808 plus.n126 gnd 0.137795f
C809 plus.n127 gnd 2.64316f
C810 a_n1808_13878.t11 gnd 0.185683f
C811 a_n1808_13878.t13 gnd 0.185683f
C812 a_n1808_13878.t17 gnd 0.185683f
C813 a_n1808_13878.n0 gnd 1.46451f
C814 a_n1808_13878.t8 gnd 0.185683f
C815 a_n1808_13878.t10 gnd 0.185683f
C816 a_n1808_13878.n1 gnd 1.46364f
C817 a_n1808_13878.t14 gnd 0.185683f
C818 a_n1808_13878.t9 gnd 0.185683f
C819 a_n1808_13878.n2 gnd 1.46209f
C820 a_n1808_13878.n3 gnd 2.04299f
C821 a_n1808_13878.t12 gnd 0.185683f
C822 a_n1808_13878.t19 gnd 0.185683f
C823 a_n1808_13878.n4 gnd 1.46209f
C824 a_n1808_13878.n5 gnd 3.70273f
C825 a_n1808_13878.t1 gnd 1.73864f
C826 a_n1808_13878.t4 gnd 0.185683f
C827 a_n1808_13878.t5 gnd 0.185683f
C828 a_n1808_13878.n6 gnd 1.30795f
C829 a_n1808_13878.n7 gnd 1.46144f
C830 a_n1808_13878.t0 gnd 1.73518f
C831 a_n1808_13878.n8 gnd 0.735417f
C832 a_n1808_13878.t3 gnd 1.73518f
C833 a_n1808_13878.n9 gnd 0.735417f
C834 a_n1808_13878.t6 gnd 0.185683f
C835 a_n1808_13878.t7 gnd 0.185683f
C836 a_n1808_13878.n10 gnd 1.30795f
C837 a_n1808_13878.n11 gnd 0.742539f
C838 a_n1808_13878.t2 gnd 1.73518f
C839 a_n1808_13878.n12 gnd 1.73174f
C840 a_n1808_13878.n13 gnd 2.52099f
C841 a_n1808_13878.t15 gnd 0.185683f
C842 a_n1808_13878.t16 gnd 0.185683f
C843 a_n1808_13878.n14 gnd 1.46209f
C844 a_n1808_13878.n15 gnd 1.80499f
C845 a_n1808_13878.n16 gnd 1.31424f
C846 a_n1808_13878.n17 gnd 1.46209f
C847 a_n1808_13878.t18 gnd 0.185683f
C848 a_n1986_8322.t0 gnd 38.672398f
C849 a_n1986_8322.t2 gnd 27.512402f
C850 a_n1986_8322.t3 gnd 19.268198f
C851 a_n1986_8322.t1 gnd 38.672398f
C852 a_n1986_8322.t13 gnd 0.875792f
C853 a_n1986_8322.t21 gnd 0.093533f
C854 a_n1986_8322.t16 gnd 0.093533f
C855 a_n1986_8322.n0 gnd 0.658844f
C856 a_n1986_8322.n1 gnd 0.736161f
C857 a_n1986_8322.t19 gnd 0.093533f
C858 a_n1986_8322.t18 gnd 0.093533f
C859 a_n1986_8322.n2 gnd 0.658844f
C860 a_n1986_8322.n3 gnd 0.374034f
C861 a_n1986_8322.t12 gnd 0.874048f
C862 a_n1986_8322.n4 gnd 1.39896f
C863 a_n1986_8322.t6 gnd 0.875792f
C864 a_n1986_8322.t10 gnd 0.093533f
C865 a_n1986_8322.t9 gnd 0.093533f
C866 a_n1986_8322.n5 gnd 0.658844f
C867 a_n1986_8322.n6 gnd 0.736161f
C868 a_n1986_8322.t4 gnd 0.874048f
C869 a_n1986_8322.n7 gnd 0.370446f
C870 a_n1986_8322.t7 gnd 0.874048f
C871 a_n1986_8322.n8 gnd 0.370446f
C872 a_n1986_8322.t5 gnd 0.093533f
C873 a_n1986_8322.t11 gnd 0.093533f
C874 a_n1986_8322.n9 gnd 0.658844f
C875 a_n1986_8322.n10 gnd 0.374034f
C876 a_n1986_8322.t8 gnd 0.874048f
C877 a_n1986_8322.n11 gnd 0.872317f
C878 a_n1986_8322.n12 gnd 1.59071f
C879 a_n1986_8322.n13 gnd 3.20172f
C880 a_n1986_8322.t15 gnd 0.874048f
C881 a_n1986_8322.n14 gnd 0.76652f
C882 a_n1986_8322.t14 gnd 0.093533f
C883 a_n1986_8322.t23 gnd 0.093533f
C884 a_n1986_8322.n15 gnd 0.658844f
C885 a_n1986_8322.n16 gnd 0.374034f
C886 a_n1986_8322.t20 gnd 0.093533f
C887 a_n1986_8322.t17 gnd 0.093533f
C888 a_n1986_8322.n17 gnd 0.658844f
C889 a_n1986_8322.n18 gnd 0.736159f
C890 a_n1986_8322.t22 gnd 0.875794f
C891 a_n2848_n452.n0 gnd 3.415f
C892 a_n2848_n452.n1 gnd 0.285666f
C893 a_n2848_n452.n2 gnd 0.492471f
C894 a_n2848_n452.n3 gnd 0.664435f
C895 a_n2848_n452.n4 gnd 0.215942f
C896 a_n2848_n452.n5 gnd 0.282512f
C897 a_n2848_n452.n6 gnd 0.546457f
C898 a_n2848_n452.n7 gnd 0.526038f
C899 a_n2848_n452.n8 gnd 0.204894f
C900 a_n2848_n452.n9 gnd 0.150908f
C901 a_n2848_n452.n10 gnd 0.23718f
C902 a_n2848_n452.n11 gnd 0.183194f
C903 a_n2848_n452.n12 gnd 0.204894f
C904 a_n2848_n452.n13 gnd 1.0063f
C905 a_n2848_n452.n14 gnd 0.150908f
C906 a_n2848_n452.n15 gnd 0.580023f
C907 a_n2848_n452.n16 gnd 0.432289f
C908 a_n2848_n452.n17 gnd 0.215942f
C909 a_n2848_n452.n18 gnd 0.492471f
C910 a_n2848_n452.n19 gnd 0.282512f
C911 a_n2848_n452.n20 gnd 0.438486f
C912 a_n2848_n452.n21 gnd 0.215942f
C913 a_n2848_n452.n22 gnd 0.731534f
C914 a_n2848_n452.n23 gnd 0.282512f
C915 a_n2848_n452.n24 gnd 1.17886f
C916 a_n2848_n452.n25 gnd 1.91568f
C917 a_n2848_n452.n26 gnd 1.14458f
C918 a_n2848_n452.n27 gnd 1.77783f
C919 a_n2848_n452.n28 gnd 0.377489f
C920 a_n2848_n452.n29 gnd 3.11576f
C921 a_n2848_n452.n30 gnd 0.377488f
C922 a_n2848_n452.n31 gnd 3.20158f
C923 a_n2848_n452.n32 gnd 0.008361f
C924 a_n2848_n452.n34 gnd 0.285666f
C925 a_n2848_n452.n35 gnd 0.008361f
C926 a_n2848_n452.n37 gnd 0.285666f
C927 a_n2848_n452.n38 gnd 0.008361f
C928 a_n2848_n452.n39 gnd 0.28526f
C929 a_n2848_n452.n40 gnd 0.008361f
C930 a_n2848_n452.n41 gnd 0.28526f
C931 a_n2848_n452.n42 gnd 0.008361f
C932 a_n2848_n452.n43 gnd 0.28526f
C933 a_n2848_n452.n44 gnd 0.008361f
C934 a_n2848_n452.n45 gnd 0.28526f
C935 a_n2848_n452.n47 gnd 0.285666f
C936 a_n2848_n452.n48 gnd 0.008361f
C937 a_n2848_n452.n50 gnd 0.285666f
C938 a_n2848_n452.t31 gnd 0.14978f
C939 a_n2848_n452.t32 gnd 0.708223f
C940 a_n2848_n452.t38 gnd 0.696704f
C941 a_n2848_n452.t20 gnd 0.696704f
C942 a_n2848_n452.t11 gnd 0.116496f
C943 a_n2848_n452.t12 gnd 0.116496f
C944 a_n2848_n452.n52 gnd 1.03243f
C945 a_n2848_n452.t1 gnd 0.116496f
C946 a_n2848_n452.t8 gnd 0.116496f
C947 a_n2848_n452.n53 gnd 1.02939f
C948 a_n2848_n452.n54 gnd 0.912816f
C949 a_n2848_n452.t46 gnd 0.116496f
C950 a_n2848_n452.t47 gnd 0.116496f
C951 a_n2848_n452.n55 gnd 1.02939f
C952 a_n2848_n452.t17 gnd 0.116496f
C953 a_n2848_n452.t44 gnd 0.116496f
C954 a_n2848_n452.n56 gnd 1.03243f
C955 a_n2848_n452.t15 gnd 0.116496f
C956 a_n2848_n452.t3 gnd 0.116496f
C957 a_n2848_n452.n57 gnd 1.02939f
C958 a_n2848_n452.n58 gnd 0.912816f
C959 a_n2848_n452.t16 gnd 0.116496f
C960 a_n2848_n452.t6 gnd 0.116496f
C961 a_n2848_n452.n59 gnd 1.02939f
C962 a_n2848_n452.t4 gnd 0.116496f
C963 a_n2848_n452.t42 gnd 0.116496f
C964 a_n2848_n452.n60 gnd 1.0294f
C965 a_n2848_n452.n61 gnd 3.15028f
C966 a_n2848_n452.t10 gnd 0.116496f
C967 a_n2848_n452.t43 gnd 0.116496f
C968 a_n2848_n452.n62 gnd 1.0294f
C969 a_n2848_n452.n63 gnd 0.449442f
C970 a_n2848_n452.t9 gnd 0.116496f
C971 a_n2848_n452.t13 gnd 0.116496f
C972 a_n2848_n452.n64 gnd 1.0294f
C973 a_n2848_n452.t5 gnd 0.116496f
C974 a_n2848_n452.t45 gnd 0.116496f
C975 a_n2848_n452.n65 gnd 1.03243f
C976 a_n2848_n452.t14 gnd 0.116496f
C977 a_n2848_n452.t0 gnd 0.116496f
C978 a_n2848_n452.n66 gnd 1.0294f
C979 a_n2848_n452.n67 gnd 0.912814f
C980 a_n2848_n452.t2 gnd 0.116496f
C981 a_n2848_n452.t7 gnd 0.116496f
C982 a_n2848_n452.n68 gnd 1.0294f
C983 a_n2848_n452.t18 gnd 0.696704f
C984 a_n2848_n452.n69 gnd 0.302425f
C985 a_n2848_n452.t30 gnd 0.696704f
C986 a_n2848_n452.t26 gnd 0.708223f
C987 a_n2848_n452.t75 gnd 0.711378f
C988 a_n2848_n452.t58 gnd 0.696704f
C989 a_n2848_n452.t62 gnd 0.696704f
C990 a_n2848_n452.t52 gnd 0.696704f
C991 a_n2848_n452.n70 gnd 0.306315f
C992 a_n2848_n452.t67 gnd 0.696704f
C993 a_n2848_n452.t73 gnd 0.708223f
C994 a_n2848_n452.t23 gnd 1.40246f
C995 a_n2848_n452.t29 gnd 0.14978f
C996 a_n2848_n452.t41 gnd 0.14978f
C997 a_n2848_n452.n71 gnd 1.05505f
C998 a_n2848_n452.t25 gnd 0.14978f
C999 a_n2848_n452.t35 gnd 0.14978f
C1000 a_n2848_n452.n72 gnd 1.05505f
C1001 a_n2848_n452.t37 gnd 1.39967f
C1002 a_n2848_n452.t24 gnd 0.696704f
C1003 a_n2848_n452.n73 gnd 0.306315f
C1004 a_n2848_n452.t34 gnd 0.696704f
C1005 a_n2848_n452.t28 gnd 0.696704f
C1006 a_n2848_n452.t56 gnd 0.696704f
C1007 a_n2848_n452.n74 gnd 0.306315f
C1008 a_n2848_n452.t65 gnd 0.696704f
C1009 a_n2848_n452.t71 gnd 0.696704f
C1010 a_n2848_n452.t70 gnd 0.711378f
C1011 a_n2848_n452.n75 gnd 0.308932f
C1012 a_n2848_n452.t50 gnd 0.696704f
C1013 a_n2848_n452.n76 gnd 0.302425f
C1014 a_n2848_n452.n77 gnd 0.308933f
C1015 a_n2848_n452.t51 gnd 0.708223f
C1016 a_n2848_n452.t22 gnd 0.711378f
C1017 a_n2848_n452.n78 gnd 0.308932f
C1018 a_n2848_n452.t40 gnd 0.696704f
C1019 a_n2848_n452.n79 gnd 0.302425f
C1020 a_n2848_n452.n80 gnd 0.308933f
C1021 a_n2848_n452.t36 gnd 0.708223f
C1022 a_n2848_n452.n81 gnd 1.13204f
C1023 a_n2848_n452.t55 gnd 0.696704f
C1024 a_n2848_n452.n82 gnd 0.302425f
C1025 a_n2848_n452.t61 gnd 0.696704f
C1026 a_n2848_n452.n83 gnd 0.302425f
C1027 a_n2848_n452.t53 gnd 0.696704f
C1028 a_n2848_n452.n84 gnd 0.302425f
C1029 a_n2848_n452.t66 gnd 0.696704f
C1030 a_n2848_n452.n85 gnd 0.302425f
C1031 a_n2848_n452.t57 gnd 0.696704f
C1032 a_n2848_n452.n86 gnd 0.296933f
C1033 a_n2848_n452.t48 gnd 0.696704f
C1034 a_n2848_n452.n87 gnd 0.306315f
C1035 a_n2848_n452.t59 gnd 0.708378f
C1036 a_n2848_n452.t68 gnd 0.696704f
C1037 a_n2848_n452.n88 gnd 0.296933f
C1038 a_n2848_n452.t54 gnd 0.696704f
C1039 a_n2848_n452.n89 gnd 0.306315f
C1040 a_n2848_n452.t63 gnd 0.708378f
C1041 a_n2848_n452.t72 gnd 0.696704f
C1042 a_n2848_n452.n90 gnd 0.296933f
C1043 a_n2848_n452.t60 gnd 0.696704f
C1044 a_n2848_n452.n91 gnd 0.306315f
C1045 a_n2848_n452.t74 gnd 0.708378f
C1046 a_n2848_n452.t64 gnd 0.696704f
C1047 a_n2848_n452.n92 gnd 0.296933f
C1048 a_n2848_n452.t49 gnd 0.696704f
C1049 a_n2848_n452.n93 gnd 0.306315f
C1050 a_n2848_n452.t69 gnd 0.708378f
C1051 a_n2848_n452.n94 gnd 1.33845f
C1052 a_n2848_n452.n95 gnd 0.308933f
C1053 a_n2848_n452.n96 gnd 0.302425f
C1054 a_n2848_n452.n97 gnd 0.308932f
C1055 a_n2848_n452.n98 gnd 0.308933f
C1056 a_n2848_n452.n99 gnd 0.01225f
C1057 a_n2848_n452.n100 gnd 0.302425f
C1058 a_n2848_n452.n101 gnd 0.308933f
C1059 a_n2848_n452.n102 gnd 0.786935f
C1060 a_n2848_n452.t33 gnd 1.39967f
C1061 a_n2848_n452.t39 gnd 0.14978f
C1062 a_n2848_n452.t21 gnd 0.14978f
C1063 a_n2848_n452.n103 gnd 1.05505f
C1064 a_n2848_n452.t27 gnd 1.40246f
C1065 a_n2848_n452.n104 gnd 1.05505f
C1066 a_n2848_n452.t19 gnd 0.14978f
C1067 vdd.t3 gnd 0.032757f
C1068 vdd.t9 gnd 0.032757f
C1069 vdd.n0 gnd 0.258361f
C1070 vdd.t187 gnd 0.032757f
C1071 vdd.t195 gnd 0.032757f
C1072 vdd.n1 gnd 0.257935f
C1073 vdd.n2 gnd 0.237865f
C1074 vdd.t183 gnd 0.032757f
C1075 vdd.t20 gnd 0.032757f
C1076 vdd.n3 gnd 0.257935f
C1077 vdd.n4 gnd 0.120297f
C1078 vdd.t16 gnd 0.032757f
C1079 vdd.t13 gnd 0.032757f
C1080 vdd.n5 gnd 0.257935f
C1081 vdd.n6 gnd 0.112877f
C1082 vdd.t189 gnd 0.032757f
C1083 vdd.t185 gnd 0.032757f
C1084 vdd.n7 gnd 0.258361f
C1085 vdd.t192 gnd 0.032757f
C1086 vdd.t18 gnd 0.032757f
C1087 vdd.n8 gnd 0.257935f
C1088 vdd.n9 gnd 0.237865f
C1089 vdd.t197 gnd 0.032757f
C1090 vdd.t180 gnd 0.032757f
C1091 vdd.n10 gnd 0.257935f
C1092 vdd.n11 gnd 0.120297f
C1093 vdd.t6 gnd 0.032757f
C1094 vdd.t199 gnd 0.032757f
C1095 vdd.n12 gnd 0.257935f
C1096 vdd.n13 gnd 0.112877f
C1097 vdd.n14 gnd 0.079802f
C1098 vdd.t168 gnd 0.018198f
C1099 vdd.t167 gnd 0.018198f
C1100 vdd.n15 gnd 0.167509f
C1101 vdd.t170 gnd 0.018198f
C1102 vdd.t176 gnd 0.018198f
C1103 vdd.n16 gnd 0.167019f
C1104 vdd.n17 gnd 0.290665f
C1105 vdd.t174 gnd 0.018198f
C1106 vdd.t164 gnd 0.018198f
C1107 vdd.n18 gnd 0.167019f
C1108 vdd.n19 gnd 0.120252f
C1109 vdd.t166 gnd 0.018198f
C1110 vdd.t165 gnd 0.018198f
C1111 vdd.n20 gnd 0.167509f
C1112 vdd.t173 gnd 0.018198f
C1113 vdd.t161 gnd 0.018198f
C1114 vdd.n21 gnd 0.167019f
C1115 vdd.n22 gnd 0.290665f
C1116 vdd.t175 gnd 0.018198f
C1117 vdd.t169 gnd 0.018198f
C1118 vdd.n23 gnd 0.167019f
C1119 vdd.n24 gnd 0.120252f
C1120 vdd.t172 gnd 0.018198f
C1121 vdd.t171 gnd 0.018198f
C1122 vdd.n25 gnd 0.167019f
C1123 vdd.t162 gnd 0.018198f
C1124 vdd.t163 gnd 0.018198f
C1125 vdd.n26 gnd 0.167019f
C1126 vdd.n27 gnd 19.0415f
C1127 vdd.n28 gnd 6.84325f
C1128 vdd.n29 gnd 0.004963f
C1129 vdd.n30 gnd 0.004606f
C1130 vdd.n31 gnd 0.002548f
C1131 vdd.n32 gnd 0.00585f
C1132 vdd.n33 gnd 0.002475f
C1133 vdd.n34 gnd 0.002621f
C1134 vdd.n35 gnd 0.004606f
C1135 vdd.n36 gnd 0.002475f
C1136 vdd.n37 gnd 0.00585f
C1137 vdd.n38 gnd 0.002621f
C1138 vdd.n39 gnd 0.004606f
C1139 vdd.n40 gnd 0.002475f
C1140 vdd.n41 gnd 0.004387f
C1141 vdd.n42 gnd 0.004401f
C1142 vdd.t100 gnd 0.012568f
C1143 vdd.n43 gnd 0.027964f
C1144 vdd.n44 gnd 0.145531f
C1145 vdd.n45 gnd 0.002475f
C1146 vdd.n46 gnd 0.002621f
C1147 vdd.n47 gnd 0.00585f
C1148 vdd.n48 gnd 0.00585f
C1149 vdd.n49 gnd 0.002621f
C1150 vdd.n50 gnd 0.002475f
C1151 vdd.n51 gnd 0.004606f
C1152 vdd.n52 gnd 0.004606f
C1153 vdd.n53 gnd 0.002475f
C1154 vdd.n54 gnd 0.002621f
C1155 vdd.n55 gnd 0.00585f
C1156 vdd.n56 gnd 0.00585f
C1157 vdd.n57 gnd 0.002621f
C1158 vdd.n58 gnd 0.002475f
C1159 vdd.n59 gnd 0.004606f
C1160 vdd.n60 gnd 0.004606f
C1161 vdd.n61 gnd 0.002475f
C1162 vdd.n62 gnd 0.002621f
C1163 vdd.n63 gnd 0.00585f
C1164 vdd.n64 gnd 0.00585f
C1165 vdd.n65 gnd 0.01383f
C1166 vdd.n66 gnd 0.002548f
C1167 vdd.n67 gnd 0.002475f
C1168 vdd.n68 gnd 0.011905f
C1169 vdd.n69 gnd 0.008311f
C1170 vdd.t152 gnd 0.029117f
C1171 vdd.t126 gnd 0.029117f
C1172 vdd.n70 gnd 0.200115f
C1173 vdd.n71 gnd 0.15736f
C1174 vdd.t159 gnd 0.029117f
C1175 vdd.t115 gnd 0.029117f
C1176 vdd.n72 gnd 0.200115f
C1177 vdd.n73 gnd 0.126989f
C1178 vdd.t145 gnd 0.029117f
C1179 vdd.t120 gnd 0.029117f
C1180 vdd.n74 gnd 0.200115f
C1181 vdd.n75 gnd 0.126989f
C1182 vdd.n76 gnd 0.004963f
C1183 vdd.n77 gnd 0.004606f
C1184 vdd.n78 gnd 0.002548f
C1185 vdd.n79 gnd 0.00585f
C1186 vdd.n80 gnd 0.002475f
C1187 vdd.n81 gnd 0.002621f
C1188 vdd.n82 gnd 0.004606f
C1189 vdd.n83 gnd 0.002475f
C1190 vdd.n84 gnd 0.00585f
C1191 vdd.n85 gnd 0.002621f
C1192 vdd.n86 gnd 0.004606f
C1193 vdd.n87 gnd 0.002475f
C1194 vdd.n88 gnd 0.004387f
C1195 vdd.n89 gnd 0.004401f
C1196 vdd.t158 gnd 0.012568f
C1197 vdd.n90 gnd 0.027964f
C1198 vdd.n91 gnd 0.145531f
C1199 vdd.n92 gnd 0.002475f
C1200 vdd.n93 gnd 0.002621f
C1201 vdd.n94 gnd 0.00585f
C1202 vdd.n95 gnd 0.00585f
C1203 vdd.n96 gnd 0.002621f
C1204 vdd.n97 gnd 0.002475f
C1205 vdd.n98 gnd 0.004606f
C1206 vdd.n99 gnd 0.004606f
C1207 vdd.n100 gnd 0.002475f
C1208 vdd.n101 gnd 0.002621f
C1209 vdd.n102 gnd 0.00585f
C1210 vdd.n103 gnd 0.00585f
C1211 vdd.n104 gnd 0.002621f
C1212 vdd.n105 gnd 0.002475f
C1213 vdd.n106 gnd 0.004606f
C1214 vdd.n107 gnd 0.004606f
C1215 vdd.n108 gnd 0.002475f
C1216 vdd.n109 gnd 0.002621f
C1217 vdd.n110 gnd 0.00585f
C1218 vdd.n111 gnd 0.00585f
C1219 vdd.n112 gnd 0.01383f
C1220 vdd.n113 gnd 0.002548f
C1221 vdd.n114 gnd 0.002475f
C1222 vdd.n115 gnd 0.011905f
C1223 vdd.n116 gnd 0.00805f
C1224 vdd.n117 gnd 0.09448f
C1225 vdd.n118 gnd 0.004963f
C1226 vdd.n119 gnd 0.004606f
C1227 vdd.n120 gnd 0.002548f
C1228 vdd.n121 gnd 0.00585f
C1229 vdd.n122 gnd 0.002475f
C1230 vdd.n123 gnd 0.002621f
C1231 vdd.n124 gnd 0.004606f
C1232 vdd.n125 gnd 0.002475f
C1233 vdd.n126 gnd 0.00585f
C1234 vdd.n127 gnd 0.002621f
C1235 vdd.n128 gnd 0.004606f
C1236 vdd.n129 gnd 0.002475f
C1237 vdd.n130 gnd 0.004387f
C1238 vdd.n131 gnd 0.004401f
C1239 vdd.t127 gnd 0.012568f
C1240 vdd.n132 gnd 0.027964f
C1241 vdd.n133 gnd 0.145531f
C1242 vdd.n134 gnd 0.002475f
C1243 vdd.n135 gnd 0.002621f
C1244 vdd.n136 gnd 0.00585f
C1245 vdd.n137 gnd 0.00585f
C1246 vdd.n138 gnd 0.002621f
C1247 vdd.n139 gnd 0.002475f
C1248 vdd.n140 gnd 0.004606f
C1249 vdd.n141 gnd 0.004606f
C1250 vdd.n142 gnd 0.002475f
C1251 vdd.n143 gnd 0.002621f
C1252 vdd.n144 gnd 0.00585f
C1253 vdd.n145 gnd 0.00585f
C1254 vdd.n146 gnd 0.002621f
C1255 vdd.n147 gnd 0.002475f
C1256 vdd.n148 gnd 0.004606f
C1257 vdd.n149 gnd 0.004606f
C1258 vdd.n150 gnd 0.002475f
C1259 vdd.n151 gnd 0.002621f
C1260 vdd.n152 gnd 0.00585f
C1261 vdd.n153 gnd 0.00585f
C1262 vdd.n154 gnd 0.01383f
C1263 vdd.n155 gnd 0.002548f
C1264 vdd.n156 gnd 0.002475f
C1265 vdd.n157 gnd 0.011905f
C1266 vdd.n158 gnd 0.008311f
C1267 vdd.t129 gnd 0.029117f
C1268 vdd.t140 gnd 0.029117f
C1269 vdd.n159 gnd 0.200115f
C1270 vdd.n160 gnd 0.15736f
C1271 vdd.t104 gnd 0.029117f
C1272 vdd.t123 gnd 0.029117f
C1273 vdd.n161 gnd 0.200115f
C1274 vdd.n162 gnd 0.126989f
C1275 vdd.t139 gnd 0.029117f
C1276 vdd.t160 gnd 0.029117f
C1277 vdd.n163 gnd 0.200115f
C1278 vdd.n164 gnd 0.126989f
C1279 vdd.n165 gnd 0.004963f
C1280 vdd.n166 gnd 0.004606f
C1281 vdd.n167 gnd 0.002548f
C1282 vdd.n168 gnd 0.00585f
C1283 vdd.n169 gnd 0.002475f
C1284 vdd.n170 gnd 0.002621f
C1285 vdd.n171 gnd 0.004606f
C1286 vdd.n172 gnd 0.002475f
C1287 vdd.n173 gnd 0.00585f
C1288 vdd.n174 gnd 0.002621f
C1289 vdd.n175 gnd 0.004606f
C1290 vdd.n176 gnd 0.002475f
C1291 vdd.n177 gnd 0.004387f
C1292 vdd.n178 gnd 0.004401f
C1293 vdd.t117 gnd 0.012568f
C1294 vdd.n179 gnd 0.027964f
C1295 vdd.n180 gnd 0.145531f
C1296 vdd.n181 gnd 0.002475f
C1297 vdd.n182 gnd 0.002621f
C1298 vdd.n183 gnd 0.00585f
C1299 vdd.n184 gnd 0.00585f
C1300 vdd.n185 gnd 0.002621f
C1301 vdd.n186 gnd 0.002475f
C1302 vdd.n187 gnd 0.004606f
C1303 vdd.n188 gnd 0.004606f
C1304 vdd.n189 gnd 0.002475f
C1305 vdd.n190 gnd 0.002621f
C1306 vdd.n191 gnd 0.00585f
C1307 vdd.n192 gnd 0.00585f
C1308 vdd.n193 gnd 0.002621f
C1309 vdd.n194 gnd 0.002475f
C1310 vdd.n195 gnd 0.004606f
C1311 vdd.n196 gnd 0.004606f
C1312 vdd.n197 gnd 0.002475f
C1313 vdd.n198 gnd 0.002621f
C1314 vdd.n199 gnd 0.00585f
C1315 vdd.n200 gnd 0.00585f
C1316 vdd.n201 gnd 0.01383f
C1317 vdd.n202 gnd 0.002548f
C1318 vdd.n203 gnd 0.002475f
C1319 vdd.n204 gnd 0.011905f
C1320 vdd.n205 gnd 0.00805f
C1321 vdd.n206 gnd 0.056206f
C1322 vdd.n207 gnd 0.202526f
C1323 vdd.n208 gnd 0.004963f
C1324 vdd.n209 gnd 0.004606f
C1325 vdd.n210 gnd 0.002548f
C1326 vdd.n211 gnd 0.00585f
C1327 vdd.n212 gnd 0.002475f
C1328 vdd.n213 gnd 0.002621f
C1329 vdd.n214 gnd 0.004606f
C1330 vdd.n215 gnd 0.002475f
C1331 vdd.n216 gnd 0.00585f
C1332 vdd.n217 gnd 0.002621f
C1333 vdd.n218 gnd 0.004606f
C1334 vdd.n219 gnd 0.002475f
C1335 vdd.n220 gnd 0.004387f
C1336 vdd.n221 gnd 0.004401f
C1337 vdd.t132 gnd 0.012568f
C1338 vdd.n222 gnd 0.027964f
C1339 vdd.n223 gnd 0.145531f
C1340 vdd.n224 gnd 0.002475f
C1341 vdd.n225 gnd 0.002621f
C1342 vdd.n226 gnd 0.00585f
C1343 vdd.n227 gnd 0.00585f
C1344 vdd.n228 gnd 0.002621f
C1345 vdd.n229 gnd 0.002475f
C1346 vdd.n230 gnd 0.004606f
C1347 vdd.n231 gnd 0.004606f
C1348 vdd.n232 gnd 0.002475f
C1349 vdd.n233 gnd 0.002621f
C1350 vdd.n234 gnd 0.00585f
C1351 vdd.n235 gnd 0.00585f
C1352 vdd.n236 gnd 0.002621f
C1353 vdd.n237 gnd 0.002475f
C1354 vdd.n238 gnd 0.004606f
C1355 vdd.n239 gnd 0.004606f
C1356 vdd.n240 gnd 0.002475f
C1357 vdd.n241 gnd 0.002621f
C1358 vdd.n242 gnd 0.00585f
C1359 vdd.n243 gnd 0.00585f
C1360 vdd.n244 gnd 0.01383f
C1361 vdd.n245 gnd 0.002548f
C1362 vdd.n246 gnd 0.002475f
C1363 vdd.n247 gnd 0.011905f
C1364 vdd.n248 gnd 0.008311f
C1365 vdd.t133 gnd 0.029117f
C1366 vdd.t149 gnd 0.029117f
C1367 vdd.n249 gnd 0.200115f
C1368 vdd.n250 gnd 0.15736f
C1369 vdd.t110 gnd 0.029117f
C1370 vdd.t131 gnd 0.029117f
C1371 vdd.n251 gnd 0.200115f
C1372 vdd.n252 gnd 0.126989f
C1373 vdd.t144 gnd 0.029117f
C1374 vdd.t108 gnd 0.029117f
C1375 vdd.n253 gnd 0.200115f
C1376 vdd.n254 gnd 0.126989f
C1377 vdd.n255 gnd 0.004963f
C1378 vdd.n256 gnd 0.004606f
C1379 vdd.n257 gnd 0.002548f
C1380 vdd.n258 gnd 0.00585f
C1381 vdd.n259 gnd 0.002475f
C1382 vdd.n260 gnd 0.002621f
C1383 vdd.n261 gnd 0.004606f
C1384 vdd.n262 gnd 0.002475f
C1385 vdd.n263 gnd 0.00585f
C1386 vdd.n264 gnd 0.002621f
C1387 vdd.n265 gnd 0.004606f
C1388 vdd.n266 gnd 0.002475f
C1389 vdd.n267 gnd 0.004387f
C1390 vdd.n268 gnd 0.004401f
C1391 vdd.t121 gnd 0.012568f
C1392 vdd.n269 gnd 0.027964f
C1393 vdd.n270 gnd 0.145531f
C1394 vdd.n271 gnd 0.002475f
C1395 vdd.n272 gnd 0.002621f
C1396 vdd.n273 gnd 0.00585f
C1397 vdd.n274 gnd 0.00585f
C1398 vdd.n275 gnd 0.002621f
C1399 vdd.n276 gnd 0.002475f
C1400 vdd.n277 gnd 0.004606f
C1401 vdd.n278 gnd 0.004606f
C1402 vdd.n279 gnd 0.002475f
C1403 vdd.n280 gnd 0.002621f
C1404 vdd.n281 gnd 0.00585f
C1405 vdd.n282 gnd 0.00585f
C1406 vdd.n283 gnd 0.002621f
C1407 vdd.n284 gnd 0.002475f
C1408 vdd.n285 gnd 0.004606f
C1409 vdd.n286 gnd 0.004606f
C1410 vdd.n287 gnd 0.002475f
C1411 vdd.n288 gnd 0.002621f
C1412 vdd.n289 gnd 0.00585f
C1413 vdd.n290 gnd 0.00585f
C1414 vdd.n291 gnd 0.01383f
C1415 vdd.n292 gnd 0.002548f
C1416 vdd.n293 gnd 0.002475f
C1417 vdd.n294 gnd 0.011905f
C1418 vdd.n295 gnd 0.00805f
C1419 vdd.n296 gnd 0.056206f
C1420 vdd.n297 gnd 0.21921f
C1421 vdd.n298 gnd 0.006951f
C1422 vdd.n299 gnd 0.009044f
C1423 vdd.n300 gnd 0.007279f
C1424 vdd.n301 gnd 0.007279f
C1425 vdd.n302 gnd 0.009044f
C1426 vdd.n303 gnd 0.009044f
C1427 vdd.n304 gnd 0.660846f
C1428 vdd.n305 gnd 0.009044f
C1429 vdd.n306 gnd 0.009044f
C1430 vdd.n307 gnd 0.009044f
C1431 vdd.n308 gnd 0.716301f
C1432 vdd.n309 gnd 0.009044f
C1433 vdd.n310 gnd 0.009044f
C1434 vdd.n311 gnd 0.009044f
C1435 vdd.n312 gnd 0.009044f
C1436 vdd.n313 gnd 0.007279f
C1437 vdd.n314 gnd 0.009044f
C1438 vdd.t107 gnd 0.46213f
C1439 vdd.n315 gnd 0.009044f
C1440 vdd.n316 gnd 0.009044f
C1441 vdd.n317 gnd 0.009044f
C1442 vdd.n318 gnd 0.92426f
C1443 vdd.n319 gnd 0.009044f
C1444 vdd.n320 gnd 0.009044f
C1445 vdd.n321 gnd 0.009044f
C1446 vdd.n322 gnd 0.009044f
C1447 vdd.n323 gnd 0.009044f
C1448 vdd.n324 gnd 0.007279f
C1449 vdd.n325 gnd 0.009044f
C1450 vdd.n326 gnd 0.009044f
C1451 vdd.n327 gnd 0.009044f
C1452 vdd.n328 gnd 0.022041f
C1453 vdd.n329 gnd 2.20898f
C1454 vdd.n330 gnd 0.022546f
C1455 vdd.n331 gnd 0.009044f
C1456 vdd.n332 gnd 0.009044f
C1457 vdd.n334 gnd 0.009044f
C1458 vdd.n335 gnd 0.009044f
C1459 vdd.n336 gnd 0.007279f
C1460 vdd.n337 gnd 0.007279f
C1461 vdd.n338 gnd 0.009044f
C1462 vdd.n339 gnd 0.009044f
C1463 vdd.n340 gnd 0.009044f
C1464 vdd.n341 gnd 0.009044f
C1465 vdd.n342 gnd 0.009044f
C1466 vdd.n343 gnd 0.009044f
C1467 vdd.n344 gnd 0.007279f
C1468 vdd.n346 gnd 0.009044f
C1469 vdd.n347 gnd 0.009044f
C1470 vdd.n348 gnd 0.009044f
C1471 vdd.n349 gnd 0.009044f
C1472 vdd.n350 gnd 0.009044f
C1473 vdd.n351 gnd 0.007279f
C1474 vdd.n353 gnd 0.009044f
C1475 vdd.n354 gnd 0.009044f
C1476 vdd.n355 gnd 0.009044f
C1477 vdd.n356 gnd 0.009044f
C1478 vdd.n357 gnd 0.009044f
C1479 vdd.n358 gnd 0.007279f
C1480 vdd.n360 gnd 0.009044f
C1481 vdd.n361 gnd 0.009044f
C1482 vdd.n362 gnd 0.009044f
C1483 vdd.n363 gnd 0.009044f
C1484 vdd.n364 gnd 0.006078f
C1485 vdd.t52 gnd 0.111266f
C1486 vdd.t51 gnd 0.118912f
C1487 vdd.t50 gnd 0.145312f
C1488 vdd.n365 gnd 0.186269f
C1489 vdd.n366 gnd 0.157227f
C1490 vdd.n368 gnd 0.009044f
C1491 vdd.n369 gnd 0.009044f
C1492 vdd.n370 gnd 0.007279f
C1493 vdd.n371 gnd 0.009044f
C1494 vdd.n373 gnd 0.009044f
C1495 vdd.n374 gnd 0.009044f
C1496 vdd.n375 gnd 0.009044f
C1497 vdd.n376 gnd 0.009044f
C1498 vdd.n377 gnd 0.007279f
C1499 vdd.n379 gnd 0.009044f
C1500 vdd.n380 gnd 0.009044f
C1501 vdd.n381 gnd 0.009044f
C1502 vdd.n382 gnd 0.009044f
C1503 vdd.n383 gnd 0.009044f
C1504 vdd.n384 gnd 0.007279f
C1505 vdd.n386 gnd 0.009044f
C1506 vdd.n387 gnd 0.009044f
C1507 vdd.n388 gnd 0.009044f
C1508 vdd.n389 gnd 0.009044f
C1509 vdd.n390 gnd 0.009044f
C1510 vdd.n391 gnd 0.007279f
C1511 vdd.n393 gnd 0.009044f
C1512 vdd.n394 gnd 0.009044f
C1513 vdd.n395 gnd 0.009044f
C1514 vdd.n396 gnd 0.009044f
C1515 vdd.n397 gnd 0.009044f
C1516 vdd.n398 gnd 0.007279f
C1517 vdd.n400 gnd 0.009044f
C1518 vdd.n401 gnd 0.009044f
C1519 vdd.n402 gnd 0.009044f
C1520 vdd.n403 gnd 0.009044f
C1521 vdd.n404 gnd 0.007207f
C1522 vdd.t46 gnd 0.111266f
C1523 vdd.t45 gnd 0.118912f
C1524 vdd.t43 gnd 0.145312f
C1525 vdd.n405 gnd 0.186269f
C1526 vdd.n406 gnd 0.157227f
C1527 vdd.n408 gnd 0.009044f
C1528 vdd.n409 gnd 0.009044f
C1529 vdd.n410 gnd 0.007279f
C1530 vdd.n411 gnd 0.009044f
C1531 vdd.n413 gnd 0.009044f
C1532 vdd.n414 gnd 0.009044f
C1533 vdd.n415 gnd 0.009044f
C1534 vdd.n416 gnd 0.009044f
C1535 vdd.n417 gnd 0.007279f
C1536 vdd.n419 gnd 0.009044f
C1537 vdd.n420 gnd 0.009044f
C1538 vdd.n421 gnd 0.009044f
C1539 vdd.n422 gnd 0.009044f
C1540 vdd.n423 gnd 0.009044f
C1541 vdd.n424 gnd 0.007279f
C1542 vdd.n426 gnd 0.009044f
C1543 vdd.n427 gnd 0.009044f
C1544 vdd.n428 gnd 0.009044f
C1545 vdd.n429 gnd 0.009044f
C1546 vdd.n430 gnd 0.009044f
C1547 vdd.n431 gnd 0.007279f
C1548 vdd.n433 gnd 0.009044f
C1549 vdd.n434 gnd 0.009044f
C1550 vdd.n435 gnd 0.009044f
C1551 vdd.n436 gnd 0.009044f
C1552 vdd.n437 gnd 0.009044f
C1553 vdd.n438 gnd 0.007279f
C1554 vdd.n440 gnd 0.009044f
C1555 vdd.n441 gnd 0.009044f
C1556 vdd.n442 gnd 0.009044f
C1557 vdd.n443 gnd 0.009044f
C1558 vdd.n444 gnd 0.009044f
C1559 vdd.n445 gnd 0.009044f
C1560 vdd.n446 gnd 0.007279f
C1561 vdd.n447 gnd 0.009044f
C1562 vdd.n448 gnd 0.009044f
C1563 vdd.n449 gnd 0.007279f
C1564 vdd.n450 gnd 0.009044f
C1565 vdd.n451 gnd 0.007279f
C1566 vdd.n452 gnd 0.009044f
C1567 vdd.n453 gnd 0.007279f
C1568 vdd.n454 gnd 0.009044f
C1569 vdd.n455 gnd 0.009044f
C1570 vdd.n456 gnd 0.503722f
C1571 vdd.t103 gnd 0.46213f
C1572 vdd.n457 gnd 0.009044f
C1573 vdd.n458 gnd 0.007279f
C1574 vdd.n459 gnd 0.009044f
C1575 vdd.n460 gnd 0.007279f
C1576 vdd.n461 gnd 0.009044f
C1577 vdd.t128 gnd 0.46213f
C1578 vdd.n462 gnd 0.009044f
C1579 vdd.n463 gnd 0.007279f
C1580 vdd.n464 gnd 0.009044f
C1581 vdd.n465 gnd 0.007279f
C1582 vdd.n466 gnd 0.009044f
C1583 vdd.t99 gnd 0.46213f
C1584 vdd.n467 gnd 0.577662f
C1585 vdd.n468 gnd 0.009044f
C1586 vdd.n469 gnd 0.007279f
C1587 vdd.n470 gnd 0.009044f
C1588 vdd.n471 gnd 0.007279f
C1589 vdd.n472 gnd 0.009044f
C1590 vdd.n473 gnd 0.92426f
C1591 vdd.n474 gnd 0.009044f
C1592 vdd.n475 gnd 0.007279f
C1593 vdd.n476 gnd 0.022041f
C1594 vdd.n477 gnd 0.006042f
C1595 vdd.n478 gnd 0.022041f
C1596 vdd.t22 gnd 0.46213f
C1597 vdd.n479 gnd 0.022041f
C1598 vdd.n480 gnd 0.006042f
C1599 vdd.n481 gnd 0.007778f
C1600 vdd.n482 gnd 0.007279f
C1601 vdd.n483 gnd 0.009044f
C1602 vdd.n484 gnd 6.36815f
C1603 vdd.n515 gnd 0.022546f
C1604 vdd.n516 gnd 1.27086f
C1605 vdd.n517 gnd 0.009044f
C1606 vdd.n518 gnd 0.007279f
C1607 vdd.n519 gnd 0.005788f
C1608 vdd.n520 gnd 0.014779f
C1609 vdd.n521 gnd 0.007279f
C1610 vdd.n522 gnd 0.009044f
C1611 vdd.n523 gnd 0.009044f
C1612 vdd.n524 gnd 0.009044f
C1613 vdd.n525 gnd 0.009044f
C1614 vdd.n526 gnd 0.009044f
C1615 vdd.n527 gnd 0.009044f
C1616 vdd.n528 gnd 0.009044f
C1617 vdd.n529 gnd 0.009044f
C1618 vdd.n530 gnd 0.009044f
C1619 vdd.n531 gnd 0.009044f
C1620 vdd.n532 gnd 0.009044f
C1621 vdd.n533 gnd 0.009044f
C1622 vdd.n534 gnd 0.009044f
C1623 vdd.n535 gnd 0.009044f
C1624 vdd.n536 gnd 0.006078f
C1625 vdd.n537 gnd 0.009044f
C1626 vdd.n538 gnd 0.009044f
C1627 vdd.n539 gnd 0.009044f
C1628 vdd.n540 gnd 0.009044f
C1629 vdd.n541 gnd 0.009044f
C1630 vdd.n542 gnd 0.009044f
C1631 vdd.n543 gnd 0.009044f
C1632 vdd.n544 gnd 0.009044f
C1633 vdd.n545 gnd 0.009044f
C1634 vdd.n546 gnd 0.009044f
C1635 vdd.n547 gnd 0.009044f
C1636 vdd.n548 gnd 0.009044f
C1637 vdd.n549 gnd 0.009044f
C1638 vdd.n550 gnd 0.009044f
C1639 vdd.n551 gnd 0.009044f
C1640 vdd.n552 gnd 0.009044f
C1641 vdd.n553 gnd 0.009044f
C1642 vdd.n554 gnd 0.009044f
C1643 vdd.n555 gnd 0.009044f
C1644 vdd.n556 gnd 0.007207f
C1645 vdd.t23 gnd 0.111266f
C1646 vdd.t24 gnd 0.118912f
C1647 vdd.t21 gnd 0.145312f
C1648 vdd.n557 gnd 0.186269f
C1649 vdd.n558 gnd 0.1565f
C1650 vdd.n559 gnd 0.009044f
C1651 vdd.n560 gnd 0.009044f
C1652 vdd.n561 gnd 0.009044f
C1653 vdd.n562 gnd 0.009044f
C1654 vdd.n563 gnd 0.009044f
C1655 vdd.n564 gnd 0.009044f
C1656 vdd.n565 gnd 0.009044f
C1657 vdd.n566 gnd 0.009044f
C1658 vdd.n567 gnd 0.009044f
C1659 vdd.n568 gnd 0.009044f
C1660 vdd.n569 gnd 0.009044f
C1661 vdd.n570 gnd 0.009044f
C1662 vdd.n571 gnd 0.009044f
C1663 vdd.n572 gnd 0.005788f
C1664 vdd.n575 gnd 0.00615f
C1665 vdd.n576 gnd 0.00615f
C1666 vdd.n577 gnd 0.00615f
C1667 vdd.n578 gnd 0.00615f
C1668 vdd.n579 gnd 0.00615f
C1669 vdd.n580 gnd 0.00615f
C1670 vdd.n582 gnd 0.00615f
C1671 vdd.n583 gnd 0.00615f
C1672 vdd.n585 gnd 0.00615f
C1673 vdd.n586 gnd 0.004477f
C1674 vdd.n588 gnd 0.00615f
C1675 vdd.t67 gnd 0.248519f
C1676 vdd.t66 gnd 0.25439f
C1677 vdd.t65 gnd 0.162243f
C1678 vdd.n589 gnd 0.087683f
C1679 vdd.n590 gnd 0.049737f
C1680 vdd.n591 gnd 0.008789f
C1681 vdd.n592 gnd 0.014374f
C1682 vdd.n594 gnd 0.00615f
C1683 vdd.n595 gnd 0.628497f
C1684 vdd.n596 gnd 0.013625f
C1685 vdd.n597 gnd 0.013625f
C1686 vdd.n598 gnd 0.00615f
C1687 vdd.n599 gnd 0.014593f
C1688 vdd.n600 gnd 0.00615f
C1689 vdd.n601 gnd 0.00615f
C1690 vdd.n602 gnd 0.00615f
C1691 vdd.n603 gnd 0.00615f
C1692 vdd.n604 gnd 0.00615f
C1693 vdd.n606 gnd 0.00615f
C1694 vdd.n607 gnd 0.00615f
C1695 vdd.n609 gnd 0.00615f
C1696 vdd.n610 gnd 0.00615f
C1697 vdd.n612 gnd 0.00615f
C1698 vdd.n613 gnd 0.00615f
C1699 vdd.n615 gnd 0.00615f
C1700 vdd.n616 gnd 0.00615f
C1701 vdd.n618 gnd 0.00615f
C1702 vdd.n619 gnd 0.00615f
C1703 vdd.n621 gnd 0.00615f
C1704 vdd.t60 gnd 0.248519f
C1705 vdd.t59 gnd 0.25439f
C1706 vdd.t57 gnd 0.162243f
C1707 vdd.n622 gnd 0.087683f
C1708 vdd.n623 gnd 0.049737f
C1709 vdd.n624 gnd 0.00615f
C1710 vdd.n626 gnd 0.00615f
C1711 vdd.n627 gnd 0.00615f
C1712 vdd.t58 gnd 0.314248f
C1713 vdd.n628 gnd 0.00615f
C1714 vdd.n629 gnd 0.00615f
C1715 vdd.n630 gnd 0.00615f
C1716 vdd.n631 gnd 0.00615f
C1717 vdd.n632 gnd 0.00615f
C1718 vdd.n633 gnd 0.628497f
C1719 vdd.n634 gnd 0.00615f
C1720 vdd.n635 gnd 0.00615f
C1721 vdd.n636 gnd 0.549935f
C1722 vdd.n637 gnd 0.00615f
C1723 vdd.n638 gnd 0.00615f
C1724 vdd.n639 gnd 0.005426f
C1725 vdd.n640 gnd 0.00615f
C1726 vdd.n641 gnd 0.554556f
C1727 vdd.n642 gnd 0.00615f
C1728 vdd.n643 gnd 0.00615f
C1729 vdd.n644 gnd 0.00615f
C1730 vdd.n645 gnd 0.00615f
C1731 vdd.n646 gnd 0.00615f
C1732 vdd.n647 gnd 0.628497f
C1733 vdd.n648 gnd 0.00615f
C1734 vdd.n649 gnd 0.00615f
C1735 vdd.t37 gnd 0.281899f
C1736 vdd.t7 gnd 0.073941f
C1737 vdd.n650 gnd 0.00615f
C1738 vdd.n651 gnd 0.00615f
C1739 vdd.n652 gnd 0.00615f
C1740 vdd.t10 gnd 0.314248f
C1741 vdd.n653 gnd 0.00615f
C1742 vdd.n654 gnd 0.00615f
C1743 vdd.n655 gnd 0.00615f
C1744 vdd.n656 gnd 0.00615f
C1745 vdd.n657 gnd 0.00615f
C1746 vdd.t14 gnd 0.314248f
C1747 vdd.n658 gnd 0.00615f
C1748 vdd.n659 gnd 0.00615f
C1749 vdd.n660 gnd 0.522207f
C1750 vdd.n661 gnd 0.00615f
C1751 vdd.n662 gnd 0.00615f
C1752 vdd.n663 gnd 0.00615f
C1753 vdd.n664 gnd 0.383568f
C1754 vdd.n665 gnd 0.00615f
C1755 vdd.n666 gnd 0.00615f
C1756 vdd.t184 gnd 0.314248f
C1757 vdd.n667 gnd 0.00615f
C1758 vdd.n668 gnd 0.00615f
C1759 vdd.n669 gnd 0.00615f
C1760 vdd.n670 gnd 0.522207f
C1761 vdd.n671 gnd 0.00615f
C1762 vdd.n672 gnd 0.00615f
C1763 vdd.t11 gnd 0.268035f
C1764 vdd.t188 gnd 0.244929f
C1765 vdd.n673 gnd 0.00615f
C1766 vdd.n674 gnd 0.00615f
C1767 vdd.n675 gnd 0.00615f
C1768 vdd.t17 gnd 0.314248f
C1769 vdd.n676 gnd 0.00615f
C1770 vdd.n677 gnd 0.00615f
C1771 vdd.t0 gnd 0.314248f
C1772 vdd.n678 gnd 0.00615f
C1773 vdd.n679 gnd 0.00615f
C1774 vdd.n680 gnd 0.00615f
C1775 vdd.t181 gnd 0.231065f
C1776 vdd.n681 gnd 0.00615f
C1777 vdd.n682 gnd 0.00615f
C1778 vdd.n683 gnd 0.536071f
C1779 vdd.n684 gnd 0.00615f
C1780 vdd.n685 gnd 0.00615f
C1781 vdd.n686 gnd 0.00615f
C1782 vdd.n687 gnd 0.628497f
C1783 vdd.n688 gnd 0.00615f
C1784 vdd.n689 gnd 0.00615f
C1785 vdd.t191 gnd 0.281899f
C1786 vdd.n690 gnd 0.397432f
C1787 vdd.n691 gnd 0.00615f
C1788 vdd.n692 gnd 0.00615f
C1789 vdd.n693 gnd 0.00615f
C1790 vdd.t179 gnd 0.314248f
C1791 vdd.n694 gnd 0.00615f
C1792 vdd.n695 gnd 0.00615f
C1793 vdd.n696 gnd 0.00615f
C1794 vdd.n697 gnd 0.00615f
C1795 vdd.n698 gnd 0.00615f
C1796 vdd.t196 gnd 0.628497f
C1797 vdd.n699 gnd 0.00615f
C1798 vdd.n700 gnd 0.00615f
C1799 vdd.t62 gnd 0.314248f
C1800 vdd.n701 gnd 0.00615f
C1801 vdd.n702 gnd 0.014593f
C1802 vdd.n703 gnd 0.014593f
C1803 vdd.t198 gnd 0.591526f
C1804 vdd.n704 gnd 0.013625f
C1805 vdd.n705 gnd 0.013625f
C1806 vdd.n706 gnd 0.014593f
C1807 vdd.n707 gnd 0.00615f
C1808 vdd.n708 gnd 0.00615f
C1809 vdd.t15 gnd 0.591526f
C1810 vdd.n726 gnd 0.014593f
C1811 vdd.n744 gnd 0.013625f
C1812 vdd.n745 gnd 0.00615f
C1813 vdd.n746 gnd 0.013625f
C1814 vdd.t87 gnd 0.248519f
C1815 vdd.t86 gnd 0.25439f
C1816 vdd.t85 gnd 0.162243f
C1817 vdd.n747 gnd 0.087683f
C1818 vdd.n748 gnd 0.049737f
C1819 vdd.n749 gnd 0.014374f
C1820 vdd.n750 gnd 0.00615f
C1821 vdd.t19 gnd 0.628497f
C1822 vdd.n751 gnd 0.013625f
C1823 vdd.n752 gnd 0.00615f
C1824 vdd.n753 gnd 0.014593f
C1825 vdd.n754 gnd 0.00615f
C1826 vdd.t56 gnd 0.248519f
C1827 vdd.t55 gnd 0.25439f
C1828 vdd.t53 gnd 0.162243f
C1829 vdd.n755 gnd 0.087683f
C1830 vdd.n756 gnd 0.049737f
C1831 vdd.n757 gnd 0.008789f
C1832 vdd.n758 gnd 0.00615f
C1833 vdd.n759 gnd 0.00615f
C1834 vdd.t54 gnd 0.314248f
C1835 vdd.n760 gnd 0.00615f
C1836 vdd.n761 gnd 0.00615f
C1837 vdd.n762 gnd 0.00615f
C1838 vdd.n763 gnd 0.00615f
C1839 vdd.n764 gnd 0.00615f
C1840 vdd.n765 gnd 0.00615f
C1841 vdd.n766 gnd 0.628497f
C1842 vdd.n767 gnd 0.00615f
C1843 vdd.n768 gnd 0.00615f
C1844 vdd.t182 gnd 0.314248f
C1845 vdd.n769 gnd 0.00615f
C1846 vdd.n770 gnd 0.00615f
C1847 vdd.n771 gnd 0.00615f
C1848 vdd.n772 gnd 0.00615f
C1849 vdd.n773 gnd 0.397432f
C1850 vdd.n774 gnd 0.00615f
C1851 vdd.n775 gnd 0.00615f
C1852 vdd.n776 gnd 0.00615f
C1853 vdd.n777 gnd 0.00615f
C1854 vdd.n778 gnd 0.00615f
C1855 vdd.n779 gnd 0.536071f
C1856 vdd.n780 gnd 0.00615f
C1857 vdd.n781 gnd 0.00615f
C1858 vdd.t194 gnd 0.281899f
C1859 vdd.t4 gnd 0.231065f
C1860 vdd.n782 gnd 0.00615f
C1861 vdd.n783 gnd 0.00615f
C1862 vdd.n784 gnd 0.00615f
C1863 vdd.t193 gnd 0.314248f
C1864 vdd.n785 gnd 0.00615f
C1865 vdd.n786 gnd 0.00615f
C1866 vdd.t186 gnd 0.314248f
C1867 vdd.n787 gnd 0.00615f
C1868 vdd.n788 gnd 0.00615f
C1869 vdd.n789 gnd 0.00615f
C1870 vdd.t8 gnd 0.244929f
C1871 vdd.n790 gnd 0.00615f
C1872 vdd.n791 gnd 0.00615f
C1873 vdd.n792 gnd 0.522207f
C1874 vdd.n793 gnd 0.00615f
C1875 vdd.n794 gnd 0.00615f
C1876 vdd.n795 gnd 0.00615f
C1877 vdd.t2 gnd 0.314248f
C1878 vdd.n796 gnd 0.00615f
C1879 vdd.n797 gnd 0.00615f
C1880 vdd.t1 gnd 0.268035f
C1881 vdd.n798 gnd 0.383568f
C1882 vdd.n799 gnd 0.00615f
C1883 vdd.n800 gnd 0.00615f
C1884 vdd.n801 gnd 0.00615f
C1885 vdd.n802 gnd 0.522207f
C1886 vdd.n803 gnd 0.00615f
C1887 vdd.n804 gnd 0.00615f
C1888 vdd.t177 gnd 0.314248f
C1889 vdd.n805 gnd 0.00615f
C1890 vdd.n806 gnd 0.00615f
C1891 vdd.n807 gnd 0.00615f
C1892 vdd.n808 gnd 0.628497f
C1893 vdd.n809 gnd 0.00615f
C1894 vdd.n810 gnd 0.00615f
C1895 vdd.t190 gnd 0.314248f
C1896 vdd.n811 gnd 0.00615f
C1897 vdd.n812 gnd 0.00615f
C1898 vdd.n813 gnd 0.00615f
C1899 vdd.t178 gnd 0.073941f
C1900 vdd.n814 gnd 0.00615f
C1901 vdd.n815 gnd 0.00615f
C1902 vdd.n816 gnd 0.00615f
C1903 vdd.t74 gnd 0.25439f
C1904 vdd.t72 gnd 0.162243f
C1905 vdd.t75 gnd 0.25439f
C1906 vdd.n817 gnd 0.142978f
C1907 vdd.n818 gnd 0.00615f
C1908 vdd.n819 gnd 0.00615f
C1909 vdd.n820 gnd 0.628497f
C1910 vdd.n821 gnd 0.00615f
C1911 vdd.n822 gnd 0.00615f
C1912 vdd.t73 gnd 0.281899f
C1913 vdd.n823 gnd 0.554556f
C1914 vdd.n824 gnd 0.00615f
C1915 vdd.n825 gnd 0.00615f
C1916 vdd.n826 gnd 0.00615f
C1917 vdd.n827 gnd 0.549935f
C1918 vdd.n828 gnd 0.00615f
C1919 vdd.n829 gnd 0.00615f
C1920 vdd.n830 gnd 0.00615f
C1921 vdd.n831 gnd 0.00615f
C1922 vdd.n832 gnd 0.00615f
C1923 vdd.n833 gnd 0.628497f
C1924 vdd.n834 gnd 0.00615f
C1925 vdd.n835 gnd 0.00615f
C1926 vdd.t69 gnd 0.314248f
C1927 vdd.n836 gnd 0.00615f
C1928 vdd.n837 gnd 0.014593f
C1929 vdd.n838 gnd 0.014593f
C1930 vdd.n839 gnd 6.36815f
C1931 vdd.n840 gnd 0.013625f
C1932 vdd.n841 gnd 0.013625f
C1933 vdd.n842 gnd 0.014593f
C1934 vdd.n843 gnd 0.00615f
C1935 vdd.n844 gnd 0.00615f
C1936 vdd.n845 gnd 0.00615f
C1937 vdd.n846 gnd 0.00615f
C1938 vdd.n847 gnd 0.00615f
C1939 vdd.n848 gnd 0.00615f
C1940 vdd.n849 gnd 0.00615f
C1941 vdd.n850 gnd 0.00615f
C1942 vdd.n852 gnd 0.00615f
C1943 vdd.n853 gnd 0.00615f
C1944 vdd.n854 gnd 0.005788f
C1945 vdd.n857 gnd 0.022546f
C1946 vdd.n858 gnd 0.007279f
C1947 vdd.n859 gnd 0.009044f
C1948 vdd.n861 gnd 0.009044f
C1949 vdd.n862 gnd 0.006042f
C1950 vdd.t29 gnd 0.46213f
C1951 vdd.n863 gnd 6.70088f
C1952 vdd.n864 gnd 0.009044f
C1953 vdd.n865 gnd 0.022546f
C1954 vdd.n866 gnd 0.007279f
C1955 vdd.n867 gnd 0.009044f
C1956 vdd.n868 gnd 0.007279f
C1957 vdd.n869 gnd 0.009044f
C1958 vdd.n870 gnd 0.92426f
C1959 vdd.n871 gnd 0.009044f
C1960 vdd.n872 gnd 0.007279f
C1961 vdd.n873 gnd 0.007279f
C1962 vdd.n874 gnd 0.009044f
C1963 vdd.n875 gnd 0.007279f
C1964 vdd.n876 gnd 0.009044f
C1965 vdd.t97 gnd 0.46213f
C1966 vdd.n877 gnd 0.009044f
C1967 vdd.n878 gnd 0.007279f
C1968 vdd.n879 gnd 0.009044f
C1969 vdd.n880 gnd 0.007279f
C1970 vdd.n881 gnd 0.009044f
C1971 vdd.t150 gnd 0.46213f
C1972 vdd.n882 gnd 0.009044f
C1973 vdd.n883 gnd 0.007279f
C1974 vdd.n884 gnd 0.009044f
C1975 vdd.n885 gnd 0.007279f
C1976 vdd.n886 gnd 0.009044f
C1977 vdd.n887 gnd 0.725544f
C1978 vdd.n888 gnd 0.767136f
C1979 vdd.t105 gnd 0.46213f
C1980 vdd.n889 gnd 0.009044f
C1981 vdd.n890 gnd 0.007279f
C1982 vdd.n891 gnd 0.004963f
C1983 vdd.n892 gnd 0.004606f
C1984 vdd.n893 gnd 0.002548f
C1985 vdd.n894 gnd 0.00585f
C1986 vdd.n895 gnd 0.002475f
C1987 vdd.n896 gnd 0.002621f
C1988 vdd.n897 gnd 0.004606f
C1989 vdd.n898 gnd 0.002475f
C1990 vdd.n899 gnd 0.00585f
C1991 vdd.n900 gnd 0.002621f
C1992 vdd.n901 gnd 0.004606f
C1993 vdd.n902 gnd 0.002475f
C1994 vdd.n903 gnd 0.004387f
C1995 vdd.n904 gnd 0.004401f
C1996 vdd.t98 gnd 0.012568f
C1997 vdd.n905 gnd 0.027964f
C1998 vdd.n906 gnd 0.145531f
C1999 vdd.n907 gnd 0.002475f
C2000 vdd.n908 gnd 0.002621f
C2001 vdd.n909 gnd 0.00585f
C2002 vdd.n910 gnd 0.00585f
C2003 vdd.n911 gnd 0.002621f
C2004 vdd.n912 gnd 0.002475f
C2005 vdd.n913 gnd 0.004606f
C2006 vdd.n914 gnd 0.004606f
C2007 vdd.n915 gnd 0.002475f
C2008 vdd.n916 gnd 0.002621f
C2009 vdd.n917 gnd 0.00585f
C2010 vdd.n918 gnd 0.00585f
C2011 vdd.n919 gnd 0.002621f
C2012 vdd.n920 gnd 0.002475f
C2013 vdd.n921 gnd 0.004606f
C2014 vdd.n922 gnd 0.004606f
C2015 vdd.n923 gnd 0.002475f
C2016 vdd.n924 gnd 0.002621f
C2017 vdd.n925 gnd 0.00585f
C2018 vdd.n926 gnd 0.00585f
C2019 vdd.n927 gnd 0.01383f
C2020 vdd.n928 gnd 0.002548f
C2021 vdd.n929 gnd 0.002475f
C2022 vdd.n930 gnd 0.011905f
C2023 vdd.n931 gnd 0.008311f
C2024 vdd.t124 gnd 0.029117f
C2025 vdd.t153 gnd 0.029117f
C2026 vdd.n932 gnd 0.200115f
C2027 vdd.n933 gnd 0.15736f
C2028 vdd.t113 gnd 0.029117f
C2029 vdd.t141 gnd 0.029117f
C2030 vdd.n934 gnd 0.200115f
C2031 vdd.n935 gnd 0.126989f
C2032 vdd.t119 gnd 0.029117f
C2033 vdd.t147 gnd 0.029117f
C2034 vdd.n936 gnd 0.200115f
C2035 vdd.n937 gnd 0.126989f
C2036 vdd.n938 gnd 0.004963f
C2037 vdd.n939 gnd 0.004606f
C2038 vdd.n940 gnd 0.002548f
C2039 vdd.n941 gnd 0.00585f
C2040 vdd.n942 gnd 0.002475f
C2041 vdd.n943 gnd 0.002621f
C2042 vdd.n944 gnd 0.004606f
C2043 vdd.n945 gnd 0.002475f
C2044 vdd.n946 gnd 0.00585f
C2045 vdd.n947 gnd 0.002621f
C2046 vdd.n948 gnd 0.004606f
C2047 vdd.n949 gnd 0.002475f
C2048 vdd.n950 gnd 0.004387f
C2049 vdd.n951 gnd 0.004401f
C2050 vdd.t157 gnd 0.012568f
C2051 vdd.n952 gnd 0.027964f
C2052 vdd.n953 gnd 0.145531f
C2053 vdd.n954 gnd 0.002475f
C2054 vdd.n955 gnd 0.002621f
C2055 vdd.n956 gnd 0.00585f
C2056 vdd.n957 gnd 0.00585f
C2057 vdd.n958 gnd 0.002621f
C2058 vdd.n959 gnd 0.002475f
C2059 vdd.n960 gnd 0.004606f
C2060 vdd.n961 gnd 0.004606f
C2061 vdd.n962 gnd 0.002475f
C2062 vdd.n963 gnd 0.002621f
C2063 vdd.n964 gnd 0.00585f
C2064 vdd.n965 gnd 0.00585f
C2065 vdd.n966 gnd 0.002621f
C2066 vdd.n967 gnd 0.002475f
C2067 vdd.n968 gnd 0.004606f
C2068 vdd.n969 gnd 0.004606f
C2069 vdd.n970 gnd 0.002475f
C2070 vdd.n971 gnd 0.002621f
C2071 vdd.n972 gnd 0.00585f
C2072 vdd.n973 gnd 0.00585f
C2073 vdd.n974 gnd 0.01383f
C2074 vdd.n975 gnd 0.002548f
C2075 vdd.n976 gnd 0.002475f
C2076 vdd.n977 gnd 0.011905f
C2077 vdd.n978 gnd 0.00805f
C2078 vdd.n979 gnd 0.09448f
C2079 vdd.n980 gnd 0.004963f
C2080 vdd.n981 gnd 0.004606f
C2081 vdd.n982 gnd 0.002548f
C2082 vdd.n983 gnd 0.00585f
C2083 vdd.n984 gnd 0.002475f
C2084 vdd.n985 gnd 0.002621f
C2085 vdd.n986 gnd 0.004606f
C2086 vdd.n987 gnd 0.002475f
C2087 vdd.n988 gnd 0.00585f
C2088 vdd.n989 gnd 0.002621f
C2089 vdd.n990 gnd 0.004606f
C2090 vdd.n991 gnd 0.002475f
C2091 vdd.n992 gnd 0.004387f
C2092 vdd.n993 gnd 0.004401f
C2093 vdd.t148 gnd 0.012568f
C2094 vdd.n994 gnd 0.027964f
C2095 vdd.n995 gnd 0.145531f
C2096 vdd.n996 gnd 0.002475f
C2097 vdd.n997 gnd 0.002621f
C2098 vdd.n998 gnd 0.00585f
C2099 vdd.n999 gnd 0.00585f
C2100 vdd.n1000 gnd 0.002621f
C2101 vdd.n1001 gnd 0.002475f
C2102 vdd.n1002 gnd 0.004606f
C2103 vdd.n1003 gnd 0.004606f
C2104 vdd.n1004 gnd 0.002475f
C2105 vdd.n1005 gnd 0.002621f
C2106 vdd.n1006 gnd 0.00585f
C2107 vdd.n1007 gnd 0.00585f
C2108 vdd.n1008 gnd 0.002621f
C2109 vdd.n1009 gnd 0.002475f
C2110 vdd.n1010 gnd 0.004606f
C2111 vdd.n1011 gnd 0.004606f
C2112 vdd.n1012 gnd 0.002475f
C2113 vdd.n1013 gnd 0.002621f
C2114 vdd.n1014 gnd 0.00585f
C2115 vdd.n1015 gnd 0.00585f
C2116 vdd.n1016 gnd 0.01383f
C2117 vdd.n1017 gnd 0.002548f
C2118 vdd.n1018 gnd 0.002475f
C2119 vdd.n1019 gnd 0.011905f
C2120 vdd.n1020 gnd 0.008311f
C2121 vdd.t106 gnd 0.029117f
C2122 vdd.t151 gnd 0.029117f
C2123 vdd.n1021 gnd 0.200115f
C2124 vdd.n1022 gnd 0.15736f
C2125 vdd.t146 gnd 0.029117f
C2126 vdd.t137 gnd 0.029117f
C2127 vdd.n1023 gnd 0.200115f
C2128 vdd.n1024 gnd 0.126989f
C2129 vdd.t122 gnd 0.029117f
C2130 vdd.t102 gnd 0.029117f
C2131 vdd.n1025 gnd 0.200115f
C2132 vdd.n1026 gnd 0.126989f
C2133 vdd.n1027 gnd 0.004963f
C2134 vdd.n1028 gnd 0.004606f
C2135 vdd.n1029 gnd 0.002548f
C2136 vdd.n1030 gnd 0.00585f
C2137 vdd.n1031 gnd 0.002475f
C2138 vdd.n1032 gnd 0.002621f
C2139 vdd.n1033 gnd 0.004606f
C2140 vdd.n1034 gnd 0.002475f
C2141 vdd.n1035 gnd 0.00585f
C2142 vdd.n1036 gnd 0.002621f
C2143 vdd.n1037 gnd 0.004606f
C2144 vdd.n1038 gnd 0.002475f
C2145 vdd.n1039 gnd 0.004387f
C2146 vdd.n1040 gnd 0.004401f
C2147 vdd.t135 gnd 0.012568f
C2148 vdd.n1041 gnd 0.027964f
C2149 vdd.n1042 gnd 0.145531f
C2150 vdd.n1043 gnd 0.002475f
C2151 vdd.n1044 gnd 0.002621f
C2152 vdd.n1045 gnd 0.00585f
C2153 vdd.n1046 gnd 0.00585f
C2154 vdd.n1047 gnd 0.002621f
C2155 vdd.n1048 gnd 0.002475f
C2156 vdd.n1049 gnd 0.004606f
C2157 vdd.n1050 gnd 0.004606f
C2158 vdd.n1051 gnd 0.002475f
C2159 vdd.n1052 gnd 0.002621f
C2160 vdd.n1053 gnd 0.00585f
C2161 vdd.n1054 gnd 0.00585f
C2162 vdd.n1055 gnd 0.002621f
C2163 vdd.n1056 gnd 0.002475f
C2164 vdd.n1057 gnd 0.004606f
C2165 vdd.n1058 gnd 0.004606f
C2166 vdd.n1059 gnd 0.002475f
C2167 vdd.n1060 gnd 0.002621f
C2168 vdd.n1061 gnd 0.00585f
C2169 vdd.n1062 gnd 0.00585f
C2170 vdd.n1063 gnd 0.01383f
C2171 vdd.n1064 gnd 0.002548f
C2172 vdd.n1065 gnd 0.002475f
C2173 vdd.n1066 gnd 0.011905f
C2174 vdd.n1067 gnd 0.00805f
C2175 vdd.n1068 gnd 0.056206f
C2176 vdd.n1069 gnd 0.202526f
C2177 vdd.n1070 gnd 0.004963f
C2178 vdd.n1071 gnd 0.004606f
C2179 vdd.n1072 gnd 0.002548f
C2180 vdd.n1073 gnd 0.00585f
C2181 vdd.n1074 gnd 0.002475f
C2182 vdd.n1075 gnd 0.002621f
C2183 vdd.n1076 gnd 0.004606f
C2184 vdd.n1077 gnd 0.002475f
C2185 vdd.n1078 gnd 0.00585f
C2186 vdd.n1079 gnd 0.002621f
C2187 vdd.n1080 gnd 0.004606f
C2188 vdd.n1081 gnd 0.002475f
C2189 vdd.n1082 gnd 0.004387f
C2190 vdd.n1083 gnd 0.004401f
C2191 vdd.t156 gnd 0.012568f
C2192 vdd.n1084 gnd 0.027964f
C2193 vdd.n1085 gnd 0.145531f
C2194 vdd.n1086 gnd 0.002475f
C2195 vdd.n1087 gnd 0.002621f
C2196 vdd.n1088 gnd 0.00585f
C2197 vdd.n1089 gnd 0.00585f
C2198 vdd.n1090 gnd 0.002621f
C2199 vdd.n1091 gnd 0.002475f
C2200 vdd.n1092 gnd 0.004606f
C2201 vdd.n1093 gnd 0.004606f
C2202 vdd.n1094 gnd 0.002475f
C2203 vdd.n1095 gnd 0.002621f
C2204 vdd.n1096 gnd 0.00585f
C2205 vdd.n1097 gnd 0.00585f
C2206 vdd.n1098 gnd 0.002621f
C2207 vdd.n1099 gnd 0.002475f
C2208 vdd.n1100 gnd 0.004606f
C2209 vdd.n1101 gnd 0.004606f
C2210 vdd.n1102 gnd 0.002475f
C2211 vdd.n1103 gnd 0.002621f
C2212 vdd.n1104 gnd 0.00585f
C2213 vdd.n1105 gnd 0.00585f
C2214 vdd.n1106 gnd 0.01383f
C2215 vdd.n1107 gnd 0.002548f
C2216 vdd.n1108 gnd 0.002475f
C2217 vdd.n1109 gnd 0.011905f
C2218 vdd.n1110 gnd 0.008311f
C2219 vdd.t111 gnd 0.029117f
C2220 vdd.t155 gnd 0.029117f
C2221 vdd.n1111 gnd 0.200115f
C2222 vdd.n1112 gnd 0.15736f
C2223 vdd.t154 gnd 0.029117f
C2224 vdd.t143 gnd 0.029117f
C2225 vdd.n1113 gnd 0.200115f
C2226 vdd.n1114 gnd 0.126989f
C2227 vdd.t130 gnd 0.029117f
C2228 vdd.t109 gnd 0.029117f
C2229 vdd.n1115 gnd 0.200115f
C2230 vdd.n1116 gnd 0.126989f
C2231 vdd.n1117 gnd 0.004963f
C2232 vdd.n1118 gnd 0.004606f
C2233 vdd.n1119 gnd 0.002548f
C2234 vdd.n1120 gnd 0.00585f
C2235 vdd.n1121 gnd 0.002475f
C2236 vdd.n1122 gnd 0.002621f
C2237 vdd.n1123 gnd 0.004606f
C2238 vdd.n1124 gnd 0.002475f
C2239 vdd.n1125 gnd 0.00585f
C2240 vdd.n1126 gnd 0.002621f
C2241 vdd.n1127 gnd 0.004606f
C2242 vdd.n1128 gnd 0.002475f
C2243 vdd.n1129 gnd 0.004387f
C2244 vdd.n1130 gnd 0.004401f
C2245 vdd.t142 gnd 0.012568f
C2246 vdd.n1131 gnd 0.027964f
C2247 vdd.n1132 gnd 0.145531f
C2248 vdd.n1133 gnd 0.002475f
C2249 vdd.n1134 gnd 0.002621f
C2250 vdd.n1135 gnd 0.00585f
C2251 vdd.n1136 gnd 0.00585f
C2252 vdd.n1137 gnd 0.002621f
C2253 vdd.n1138 gnd 0.002475f
C2254 vdd.n1139 gnd 0.004606f
C2255 vdd.n1140 gnd 0.004606f
C2256 vdd.n1141 gnd 0.002475f
C2257 vdd.n1142 gnd 0.002621f
C2258 vdd.n1143 gnd 0.00585f
C2259 vdd.n1144 gnd 0.00585f
C2260 vdd.n1145 gnd 0.002621f
C2261 vdd.n1146 gnd 0.002475f
C2262 vdd.n1147 gnd 0.004606f
C2263 vdd.n1148 gnd 0.004606f
C2264 vdd.n1149 gnd 0.002475f
C2265 vdd.n1150 gnd 0.002621f
C2266 vdd.n1151 gnd 0.00585f
C2267 vdd.n1152 gnd 0.00585f
C2268 vdd.n1153 gnd 0.01383f
C2269 vdd.n1154 gnd 0.002548f
C2270 vdd.n1155 gnd 0.002475f
C2271 vdd.n1156 gnd 0.011905f
C2272 vdd.n1157 gnd 0.00805f
C2273 vdd.n1158 gnd 0.056206f
C2274 vdd.n1159 gnd 0.21921f
C2275 vdd.n1160 gnd 1.8423f
C2276 vdd.n1161 gnd 0.533453f
C2277 vdd.n1162 gnd 0.007279f
C2278 vdd.n1163 gnd 0.009044f
C2279 vdd.n1164 gnd 0.56842f
C2280 vdd.n1165 gnd 0.009044f
C2281 vdd.n1166 gnd 0.007279f
C2282 vdd.n1167 gnd 0.009044f
C2283 vdd.n1168 gnd 0.007279f
C2284 vdd.n1169 gnd 0.009044f
C2285 vdd.t101 gnd 0.46213f
C2286 vdd.t112 gnd 0.46213f
C2287 vdd.n1170 gnd 0.009044f
C2288 vdd.n1171 gnd 0.007279f
C2289 vdd.n1172 gnd 0.009044f
C2290 vdd.n1173 gnd 0.007279f
C2291 vdd.n1174 gnd 0.009044f
C2292 vdd.t118 gnd 0.46213f
C2293 vdd.n1175 gnd 0.009044f
C2294 vdd.n1176 gnd 0.007279f
C2295 vdd.n1177 gnd 0.009044f
C2296 vdd.n1178 gnd 0.007279f
C2297 vdd.n1179 gnd 0.009044f
C2298 vdd.t134 gnd 0.46213f
C2299 vdd.n1180 gnd 0.670088f
C2300 vdd.n1181 gnd 0.009044f
C2301 vdd.n1182 gnd 0.007279f
C2302 vdd.n1183 gnd 0.009044f
C2303 vdd.n1184 gnd 0.007279f
C2304 vdd.n1185 gnd 0.009044f
C2305 vdd.n1186 gnd 0.92426f
C2306 vdd.n1187 gnd 0.009044f
C2307 vdd.n1188 gnd 0.007279f
C2308 vdd.n1189 gnd 0.022041f
C2309 vdd.n1190 gnd 0.006042f
C2310 vdd.n1191 gnd 0.022041f
C2311 vdd.t33 gnd 0.46213f
C2312 vdd.n1192 gnd 0.022041f
C2313 vdd.n1193 gnd 0.006042f
C2314 vdd.n1194 gnd 0.009044f
C2315 vdd.n1195 gnd 0.007279f
C2316 vdd.n1196 gnd 0.009044f
C2317 vdd.n1227 gnd 0.022546f
C2318 vdd.n1228 gnd 1.36328f
C2319 vdd.n1229 gnd 0.009044f
C2320 vdd.n1230 gnd 0.007279f
C2321 vdd.n1231 gnd 0.009044f
C2322 vdd.n1232 gnd 0.009044f
C2323 vdd.n1233 gnd 0.009044f
C2324 vdd.n1234 gnd 0.009044f
C2325 vdd.n1235 gnd 0.009044f
C2326 vdd.n1236 gnd 0.007279f
C2327 vdd.n1237 gnd 0.009044f
C2328 vdd.n1238 gnd 0.009044f
C2329 vdd.n1239 gnd 0.009044f
C2330 vdd.n1240 gnd 0.009044f
C2331 vdd.n1241 gnd 0.009044f
C2332 vdd.n1242 gnd 0.007279f
C2333 vdd.n1243 gnd 0.009044f
C2334 vdd.n1244 gnd 0.009044f
C2335 vdd.n1245 gnd 0.009044f
C2336 vdd.n1246 gnd 0.009044f
C2337 vdd.n1247 gnd 0.009044f
C2338 vdd.n1248 gnd 0.007279f
C2339 vdd.n1249 gnd 0.009044f
C2340 vdd.n1250 gnd 0.009044f
C2341 vdd.n1251 gnd 0.009044f
C2342 vdd.n1252 gnd 0.009044f
C2343 vdd.n1253 gnd 0.009044f
C2344 vdd.t83 gnd 0.111266f
C2345 vdd.t84 gnd 0.118912f
C2346 vdd.t82 gnd 0.145312f
C2347 vdd.n1254 gnd 0.186269f
C2348 vdd.n1255 gnd 0.157227f
C2349 vdd.n1256 gnd 0.015578f
C2350 vdd.n1257 gnd 0.009044f
C2351 vdd.n1258 gnd 0.009044f
C2352 vdd.n1259 gnd 0.009044f
C2353 vdd.n1260 gnd 0.009044f
C2354 vdd.n1261 gnd 0.009044f
C2355 vdd.n1262 gnd 0.007279f
C2356 vdd.n1263 gnd 0.009044f
C2357 vdd.n1264 gnd 0.009044f
C2358 vdd.n1265 gnd 0.009044f
C2359 vdd.n1266 gnd 0.009044f
C2360 vdd.n1267 gnd 0.009044f
C2361 vdd.n1268 gnd 0.007279f
C2362 vdd.n1269 gnd 0.009044f
C2363 vdd.n1270 gnd 0.009044f
C2364 vdd.n1271 gnd 0.009044f
C2365 vdd.n1272 gnd 0.009044f
C2366 vdd.n1273 gnd 0.009044f
C2367 vdd.n1274 gnd 0.007279f
C2368 vdd.n1275 gnd 0.009044f
C2369 vdd.n1276 gnd 0.009044f
C2370 vdd.n1277 gnd 0.009044f
C2371 vdd.n1278 gnd 0.009044f
C2372 vdd.n1279 gnd 0.009044f
C2373 vdd.n1280 gnd 0.007279f
C2374 vdd.n1281 gnd 0.009044f
C2375 vdd.n1282 gnd 0.009044f
C2376 vdd.n1283 gnd 0.009044f
C2377 vdd.n1284 gnd 0.009044f
C2378 vdd.n1285 gnd 0.009044f
C2379 vdd.n1286 gnd 0.007279f
C2380 vdd.n1287 gnd 0.009044f
C2381 vdd.n1288 gnd 0.009044f
C2382 vdd.n1289 gnd 0.009044f
C2383 vdd.n1290 gnd 0.009044f
C2384 vdd.n1291 gnd 0.007279f
C2385 vdd.n1292 gnd 0.009044f
C2386 vdd.n1293 gnd 0.009044f
C2387 vdd.n1294 gnd 0.009044f
C2388 vdd.n1295 gnd 0.009044f
C2389 vdd.n1296 gnd 0.009044f
C2390 vdd.n1297 gnd 0.007279f
C2391 vdd.n1298 gnd 0.009044f
C2392 vdd.n1299 gnd 0.009044f
C2393 vdd.n1300 gnd 0.009044f
C2394 vdd.n1301 gnd 0.009044f
C2395 vdd.n1302 gnd 0.009044f
C2396 vdd.n1303 gnd 0.007279f
C2397 vdd.n1304 gnd 0.009044f
C2398 vdd.n1305 gnd 0.009044f
C2399 vdd.n1306 gnd 0.009044f
C2400 vdd.n1307 gnd 0.009044f
C2401 vdd.n1308 gnd 0.009044f
C2402 vdd.n1309 gnd 0.007279f
C2403 vdd.n1310 gnd 0.009044f
C2404 vdd.n1311 gnd 0.009044f
C2405 vdd.n1312 gnd 0.009044f
C2406 vdd.n1313 gnd 0.009044f
C2407 vdd.n1314 gnd 0.009044f
C2408 vdd.n1315 gnd 0.007279f
C2409 vdd.n1316 gnd 0.009044f
C2410 vdd.n1317 gnd 0.009044f
C2411 vdd.n1318 gnd 0.009044f
C2412 vdd.n1319 gnd 0.009044f
C2413 vdd.t34 gnd 0.111266f
C2414 vdd.t35 gnd 0.118912f
C2415 vdd.t32 gnd 0.145312f
C2416 vdd.n1320 gnd 0.186269f
C2417 vdd.n1321 gnd 0.157227f
C2418 vdd.n1322 gnd 0.011938f
C2419 vdd.n1323 gnd 0.003458f
C2420 vdd.n1324 gnd 0.022546f
C2421 vdd.n1325 gnd 0.009044f
C2422 vdd.n1326 gnd 0.003822f
C2423 vdd.n1327 gnd 0.007279f
C2424 vdd.n1328 gnd 0.007279f
C2425 vdd.n1329 gnd 0.009044f
C2426 vdd.n1330 gnd 0.009044f
C2427 vdd.n1331 gnd 0.009044f
C2428 vdd.n1332 gnd 0.007279f
C2429 vdd.n1333 gnd 0.007279f
C2430 vdd.n1334 gnd 0.007279f
C2431 vdd.n1335 gnd 0.009044f
C2432 vdd.n1336 gnd 0.009044f
C2433 vdd.n1337 gnd 0.009044f
C2434 vdd.n1338 gnd 0.007279f
C2435 vdd.n1339 gnd 0.007279f
C2436 vdd.n1340 gnd 0.007279f
C2437 vdd.n1341 gnd 0.009044f
C2438 vdd.n1342 gnd 0.009044f
C2439 vdd.n1343 gnd 0.009044f
C2440 vdd.n1344 gnd 0.007279f
C2441 vdd.n1345 gnd 0.007279f
C2442 vdd.n1346 gnd 0.007279f
C2443 vdd.n1347 gnd 0.009044f
C2444 vdd.n1348 gnd 0.009044f
C2445 vdd.n1349 gnd 0.009044f
C2446 vdd.n1350 gnd 0.007279f
C2447 vdd.n1351 gnd 0.007279f
C2448 vdd.n1352 gnd 0.007279f
C2449 vdd.n1353 gnd 0.009044f
C2450 vdd.n1354 gnd 0.009044f
C2451 vdd.n1355 gnd 0.009044f
C2452 vdd.n1356 gnd 0.007207f
C2453 vdd.n1357 gnd 0.009044f
C2454 vdd.t80 gnd 0.111266f
C2455 vdd.t81 gnd 0.118912f
C2456 vdd.t79 gnd 0.145312f
C2457 vdd.n1358 gnd 0.186269f
C2458 vdd.n1359 gnd 0.157227f
C2459 vdd.n1360 gnd 0.015578f
C2460 vdd.n1361 gnd 0.00495f
C2461 vdd.n1362 gnd 0.009044f
C2462 vdd.n1363 gnd 0.009044f
C2463 vdd.n1364 gnd 0.009044f
C2464 vdd.n1365 gnd 0.007279f
C2465 vdd.n1366 gnd 0.007279f
C2466 vdd.n1367 gnd 0.007279f
C2467 vdd.n1368 gnd 0.009044f
C2468 vdd.n1369 gnd 0.009044f
C2469 vdd.n1370 gnd 0.009044f
C2470 vdd.n1371 gnd 0.007279f
C2471 vdd.n1372 gnd 0.007279f
C2472 vdd.n1373 gnd 0.007279f
C2473 vdd.n1374 gnd 0.009044f
C2474 vdd.n1375 gnd 0.009044f
C2475 vdd.n1376 gnd 0.009044f
C2476 vdd.n1377 gnd 0.007279f
C2477 vdd.n1378 gnd 0.007279f
C2478 vdd.n1379 gnd 0.007279f
C2479 vdd.n1380 gnd 0.009044f
C2480 vdd.n1381 gnd 0.009044f
C2481 vdd.n1382 gnd 0.009044f
C2482 vdd.n1383 gnd 0.007279f
C2483 vdd.n1384 gnd 0.007279f
C2484 vdd.n1385 gnd 0.007279f
C2485 vdd.n1386 gnd 0.009044f
C2486 vdd.n1387 gnd 0.009044f
C2487 vdd.n1388 gnd 0.009044f
C2488 vdd.n1389 gnd 0.007279f
C2489 vdd.n1390 gnd 0.007279f
C2490 vdd.n1391 gnd 0.006078f
C2491 vdd.n1392 gnd 0.009044f
C2492 vdd.n1393 gnd 0.009044f
C2493 vdd.n1394 gnd 0.009044f
C2494 vdd.n1395 gnd 0.006078f
C2495 vdd.n1396 gnd 0.007279f
C2496 vdd.n1397 gnd 0.007279f
C2497 vdd.n1398 gnd 0.009044f
C2498 vdd.n1399 gnd 0.009044f
C2499 vdd.n1400 gnd 0.009044f
C2500 vdd.n1401 gnd 0.007279f
C2501 vdd.n1402 gnd 0.007279f
C2502 vdd.n1403 gnd 0.007279f
C2503 vdd.n1404 gnd 0.009044f
C2504 vdd.n1405 gnd 0.009044f
C2505 vdd.n1406 gnd 0.009044f
C2506 vdd.n1407 gnd 0.007279f
C2507 vdd.n1408 gnd 0.007279f
C2508 vdd.n1409 gnd 0.007279f
C2509 vdd.n1410 gnd 0.009044f
C2510 vdd.n1411 gnd 0.009044f
C2511 vdd.n1412 gnd 0.009044f
C2512 vdd.n1413 gnd 0.007279f
C2513 vdd.n1414 gnd 0.007279f
C2514 vdd.n1415 gnd 0.007279f
C2515 vdd.n1416 gnd 0.009044f
C2516 vdd.n1417 gnd 0.009044f
C2517 vdd.n1418 gnd 0.009044f
C2518 vdd.n1419 gnd 0.007279f
C2519 vdd.n1420 gnd 0.009044f
C2520 vdd.n1421 gnd 2.20898f
C2521 vdd.n1423 gnd 0.022546f
C2522 vdd.n1424 gnd 0.006042f
C2523 vdd.n1425 gnd 0.022546f
C2524 vdd.n1426 gnd 0.022041f
C2525 vdd.n1427 gnd 0.009044f
C2526 vdd.n1428 gnd 0.007279f
C2527 vdd.n1429 gnd 0.009044f
C2528 vdd.n1430 gnd 0.485236f
C2529 vdd.n1431 gnd 0.009044f
C2530 vdd.n1432 gnd 0.007279f
C2531 vdd.n1433 gnd 0.009044f
C2532 vdd.n1434 gnd 0.009044f
C2533 vdd.n1435 gnd 0.009044f
C2534 vdd.n1436 gnd 0.007279f
C2535 vdd.n1437 gnd 0.009044f
C2536 vdd.n1438 gnd 0.827213f
C2537 vdd.n1439 gnd 0.92426f
C2538 vdd.n1440 gnd 0.009044f
C2539 vdd.n1441 gnd 0.007279f
C2540 vdd.n1442 gnd 0.009044f
C2541 vdd.n1443 gnd 0.009044f
C2542 vdd.n1444 gnd 0.009044f
C2543 vdd.n1445 gnd 0.007279f
C2544 vdd.n1446 gnd 0.009044f
C2545 vdd.n1447 gnd 0.559177f
C2546 vdd.n1448 gnd 0.009044f
C2547 vdd.n1449 gnd 0.007279f
C2548 vdd.n1450 gnd 0.009044f
C2549 vdd.n1451 gnd 0.009044f
C2550 vdd.n1452 gnd 0.009044f
C2551 vdd.n1453 gnd 0.007279f
C2552 vdd.n1454 gnd 0.009044f
C2553 vdd.n1455 gnd 0.512964f
C2554 vdd.n1456 gnd 0.716301f
C2555 vdd.n1457 gnd 0.009044f
C2556 vdd.n1458 gnd 0.007279f
C2557 vdd.n1459 gnd 0.009044f
C2558 vdd.n1460 gnd 0.009044f
C2559 vdd.n1461 gnd 0.006951f
C2560 vdd.n1462 gnd 0.009044f
C2561 vdd.n1463 gnd 0.007279f
C2562 vdd.n1464 gnd 0.009044f
C2563 vdd.n1465 gnd 0.767136f
C2564 vdd.n1466 gnd 0.009044f
C2565 vdd.n1467 gnd 0.007279f
C2566 vdd.n1468 gnd 0.009044f
C2567 vdd.n1469 gnd 0.009044f
C2568 vdd.n1470 gnd 0.009044f
C2569 vdd.n1471 gnd 0.007279f
C2570 vdd.n1472 gnd 0.009044f
C2571 vdd.t136 gnd 0.46213f
C2572 vdd.n1473 gnd 0.660846f
C2573 vdd.n1474 gnd 0.009044f
C2574 vdd.n1475 gnd 0.007279f
C2575 vdd.n1476 gnd 0.006951f
C2576 vdd.n1477 gnd 0.009044f
C2577 vdd.n1478 gnd 0.009044f
C2578 vdd.n1479 gnd 0.007279f
C2579 vdd.n1480 gnd 0.009044f
C2580 vdd.n1481 gnd 0.503722f
C2581 vdd.n1482 gnd 0.009044f
C2582 vdd.n1483 gnd 0.007279f
C2583 vdd.n1484 gnd 0.009044f
C2584 vdd.n1485 gnd 0.009044f
C2585 vdd.n1486 gnd 0.009044f
C2586 vdd.n1487 gnd 0.007279f
C2587 vdd.n1488 gnd 0.009044f
C2588 vdd.n1489 gnd 0.651603f
C2589 vdd.n1490 gnd 0.577662f
C2590 vdd.n1491 gnd 0.009044f
C2591 vdd.n1492 gnd 0.007279f
C2592 vdd.n1493 gnd 0.009044f
C2593 vdd.n1494 gnd 0.009044f
C2594 vdd.n1495 gnd 0.009044f
C2595 vdd.n1496 gnd 0.007279f
C2596 vdd.n1497 gnd 0.009044f
C2597 vdd.n1498 gnd 0.734786f
C2598 vdd.n1499 gnd 0.009044f
C2599 vdd.n1500 gnd 0.007279f
C2600 vdd.n1501 gnd 0.009044f
C2601 vdd.n1502 gnd 0.009044f
C2602 vdd.n1503 gnd 0.022041f
C2603 vdd.n1504 gnd 0.009044f
C2604 vdd.n1505 gnd 0.009044f
C2605 vdd.n1506 gnd 0.007279f
C2606 vdd.n1507 gnd 0.009044f
C2607 vdd.n1508 gnd 0.577662f
C2608 vdd.n1509 gnd 0.92426f
C2609 vdd.n1510 gnd 0.009044f
C2610 vdd.n1511 gnd 0.007279f
C2611 vdd.n1512 gnd 0.009044f
C2612 vdd.n1513 gnd 0.009044f
C2613 vdd.n1514 gnd 0.007778f
C2614 vdd.n1515 gnd 0.007279f
C2615 vdd.n1517 gnd 0.009044f
C2616 vdd.n1519 gnd 0.007279f
C2617 vdd.n1520 gnd 0.009044f
C2618 vdd.n1521 gnd 0.007279f
C2619 vdd.n1523 gnd 0.009044f
C2620 vdd.n1524 gnd 0.007279f
C2621 vdd.n1525 gnd 0.009044f
C2622 vdd.n1526 gnd 0.009044f
C2623 vdd.n1527 gnd 0.009044f
C2624 vdd.n1528 gnd 0.009044f
C2625 vdd.n1529 gnd 0.009044f
C2626 vdd.n1530 gnd 0.007279f
C2627 vdd.n1532 gnd 0.009044f
C2628 vdd.n1533 gnd 0.009044f
C2629 vdd.n1534 gnd 0.009044f
C2630 vdd.n1535 gnd 0.009044f
C2631 vdd.n1536 gnd 0.009044f
C2632 vdd.n1537 gnd 0.007279f
C2633 vdd.n1539 gnd 0.009044f
C2634 vdd.n1540 gnd 0.009044f
C2635 vdd.n1541 gnd 0.009044f
C2636 vdd.n1542 gnd 0.009044f
C2637 vdd.n1543 gnd 0.006078f
C2638 vdd.t49 gnd 0.111266f
C2639 vdd.t48 gnd 0.118912f
C2640 vdd.t47 gnd 0.145312f
C2641 vdd.n1544 gnd 0.186269f
C2642 vdd.n1545 gnd 0.1565f
C2643 vdd.n1547 gnd 0.009044f
C2644 vdd.n1548 gnd 0.009044f
C2645 vdd.n1549 gnd 0.007279f
C2646 vdd.n1550 gnd 0.009044f
C2647 vdd.n1552 gnd 0.009044f
C2648 vdd.n1553 gnd 0.009044f
C2649 vdd.n1554 gnd 0.009044f
C2650 vdd.n1555 gnd 0.009044f
C2651 vdd.n1556 gnd 0.007279f
C2652 vdd.n1558 gnd 0.009044f
C2653 vdd.n1559 gnd 0.009044f
C2654 vdd.n1560 gnd 0.009044f
C2655 vdd.n1561 gnd 0.009044f
C2656 vdd.n1562 gnd 0.009044f
C2657 vdd.n1563 gnd 0.007279f
C2658 vdd.n1565 gnd 0.009044f
C2659 vdd.n1566 gnd 0.009044f
C2660 vdd.n1567 gnd 0.009044f
C2661 vdd.n1568 gnd 0.009044f
C2662 vdd.n1569 gnd 0.009044f
C2663 vdd.n1570 gnd 0.007279f
C2664 vdd.n1572 gnd 0.009044f
C2665 vdd.n1573 gnd 0.009044f
C2666 vdd.n1574 gnd 0.009044f
C2667 vdd.n1575 gnd 0.009044f
C2668 vdd.n1576 gnd 0.009044f
C2669 vdd.n1577 gnd 0.007279f
C2670 vdd.n1579 gnd 0.009044f
C2671 vdd.n1580 gnd 0.009044f
C2672 vdd.n1581 gnd 0.009044f
C2673 vdd.n1582 gnd 0.009044f
C2674 vdd.n1583 gnd 0.007207f
C2675 vdd.t42 gnd 0.111266f
C2676 vdd.t41 gnd 0.118912f
C2677 vdd.t40 gnd 0.145312f
C2678 vdd.n1584 gnd 0.186269f
C2679 vdd.n1585 gnd 0.1565f
C2680 vdd.n1587 gnd 0.009044f
C2681 vdd.n1588 gnd 0.009044f
C2682 vdd.n1589 gnd 0.007279f
C2683 vdd.n1590 gnd 0.009044f
C2684 vdd.n1592 gnd 0.009044f
C2685 vdd.n1593 gnd 0.009044f
C2686 vdd.n1594 gnd 0.009044f
C2687 vdd.n1595 gnd 0.009044f
C2688 vdd.n1596 gnd 0.007279f
C2689 vdd.n1598 gnd 0.009044f
C2690 vdd.n1599 gnd 0.009044f
C2691 vdd.n1600 gnd 0.009044f
C2692 vdd.n1601 gnd 0.009044f
C2693 vdd.n1602 gnd 0.009044f
C2694 vdd.n1603 gnd 0.007279f
C2695 vdd.n1605 gnd 0.009044f
C2696 vdd.n1606 gnd 0.009044f
C2697 vdd.n1607 gnd 0.009044f
C2698 vdd.n1608 gnd 0.009044f
C2699 vdd.n1609 gnd 0.009044f
C2700 vdd.n1610 gnd 0.009044f
C2701 vdd.n1611 gnd 0.007279f
C2702 vdd.n1613 gnd 0.009044f
C2703 vdd.n1615 gnd 0.009044f
C2704 vdd.n1616 gnd 0.007279f
C2705 vdd.n1617 gnd 0.007279f
C2706 vdd.n1618 gnd 0.009044f
C2707 vdd.n1620 gnd 0.009044f
C2708 vdd.n1621 gnd 0.007279f
C2709 vdd.n1622 gnd 0.007279f
C2710 vdd.n1623 gnd 0.009044f
C2711 vdd.n1625 gnd 0.009044f
C2712 vdd.n1626 gnd 0.009044f
C2713 vdd.n1627 gnd 0.007279f
C2714 vdd.n1628 gnd 0.007279f
C2715 vdd.n1629 gnd 0.007279f
C2716 vdd.n1630 gnd 0.009044f
C2717 vdd.n1632 gnd 0.009044f
C2718 vdd.n1633 gnd 0.009044f
C2719 vdd.n1634 gnd 0.007279f
C2720 vdd.n1635 gnd 0.007279f
C2721 vdd.n1636 gnd 0.007279f
C2722 vdd.n1637 gnd 0.009044f
C2723 vdd.n1639 gnd 0.009044f
C2724 vdd.n1640 gnd 0.009044f
C2725 vdd.n1641 gnd 0.007279f
C2726 vdd.n1642 gnd 0.007279f
C2727 vdd.n1643 gnd 0.007279f
C2728 vdd.n1644 gnd 0.009044f
C2729 vdd.n1646 gnd 0.009044f
C2730 vdd.n1647 gnd 0.009044f
C2731 vdd.n1648 gnd 0.007279f
C2732 vdd.n1649 gnd 0.009044f
C2733 vdd.n1650 gnd 0.009044f
C2734 vdd.n1651 gnd 0.009044f
C2735 vdd.n1652 gnd 0.01485f
C2736 vdd.n1653 gnd 0.00495f
C2737 vdd.n1654 gnd 0.007279f
C2738 vdd.n1655 gnd 0.009044f
C2739 vdd.n1657 gnd 0.009044f
C2740 vdd.n1658 gnd 0.009044f
C2741 vdd.n1659 gnd 0.007279f
C2742 vdd.n1660 gnd 0.007279f
C2743 vdd.n1661 gnd 0.007279f
C2744 vdd.n1662 gnd 0.009044f
C2745 vdd.n1664 gnd 0.009044f
C2746 vdd.n1665 gnd 0.009044f
C2747 vdd.n1666 gnd 0.007279f
C2748 vdd.n1667 gnd 0.007279f
C2749 vdd.n1668 gnd 0.007279f
C2750 vdd.n1669 gnd 0.009044f
C2751 vdd.n1671 gnd 0.009044f
C2752 vdd.n1672 gnd 0.009044f
C2753 vdd.n1673 gnd 0.007279f
C2754 vdd.n1674 gnd 0.007279f
C2755 vdd.n1675 gnd 0.007279f
C2756 vdd.n1676 gnd 0.009044f
C2757 vdd.n1678 gnd 0.009044f
C2758 vdd.n1679 gnd 0.009044f
C2759 vdd.n1680 gnd 0.007279f
C2760 vdd.n1681 gnd 0.007279f
C2761 vdd.n1682 gnd 0.007279f
C2762 vdd.n1683 gnd 0.009044f
C2763 vdd.n1685 gnd 0.009044f
C2764 vdd.n1686 gnd 0.009044f
C2765 vdd.n1687 gnd 0.007279f
C2766 vdd.n1688 gnd 0.009044f
C2767 vdd.n1689 gnd 0.009044f
C2768 vdd.n1690 gnd 0.009044f
C2769 vdd.n1691 gnd 0.01485f
C2770 vdd.n1692 gnd 0.006078f
C2771 vdd.n1693 gnd 0.007279f
C2772 vdd.n1694 gnd 0.009044f
C2773 vdd.n1696 gnd 0.009044f
C2774 vdd.n1697 gnd 0.009044f
C2775 vdd.n1698 gnd 0.007279f
C2776 vdd.n1699 gnd 0.007279f
C2777 vdd.n1700 gnd 0.007279f
C2778 vdd.n1701 gnd 0.009044f
C2779 vdd.n1703 gnd 0.009044f
C2780 vdd.n1704 gnd 0.009044f
C2781 vdd.n1705 gnd 0.007279f
C2782 vdd.n1706 gnd 0.007279f
C2783 vdd.n1707 gnd 0.007279f
C2784 vdd.n1708 gnd 0.009044f
C2785 vdd.n1710 gnd 0.009044f
C2786 vdd.n1711 gnd 0.009044f
C2787 vdd.n1713 gnd 0.009044f
C2788 vdd.n1714 gnd 0.007279f
C2789 vdd.n1715 gnd 0.005788f
C2790 vdd.n1716 gnd 0.00615f
C2791 vdd.n1717 gnd 0.00615f
C2792 vdd.n1718 gnd 0.00615f
C2793 vdd.n1719 gnd 0.00615f
C2794 vdd.n1720 gnd 0.00615f
C2795 vdd.n1721 gnd 0.00615f
C2796 vdd.n1722 gnd 0.00615f
C2797 vdd.n1723 gnd 0.00615f
C2798 vdd.n1725 gnd 0.00615f
C2799 vdd.n1726 gnd 0.00615f
C2800 vdd.n1727 gnd 0.00615f
C2801 vdd.n1728 gnd 0.00615f
C2802 vdd.n1729 gnd 0.00615f
C2803 vdd.n1731 gnd 0.00615f
C2804 vdd.n1733 gnd 0.00615f
C2805 vdd.n1734 gnd 0.00615f
C2806 vdd.n1735 gnd 0.00615f
C2807 vdd.n1736 gnd 0.00615f
C2808 vdd.n1737 gnd 0.00615f
C2809 vdd.n1739 gnd 0.00615f
C2810 vdd.n1741 gnd 0.00615f
C2811 vdd.n1742 gnd 0.00615f
C2812 vdd.n1743 gnd 0.00615f
C2813 vdd.n1744 gnd 0.00615f
C2814 vdd.n1745 gnd 0.00615f
C2815 vdd.n1747 gnd 0.00615f
C2816 vdd.n1749 gnd 0.00615f
C2817 vdd.n1750 gnd 0.00615f
C2818 vdd.n1751 gnd 0.00615f
C2819 vdd.n1752 gnd 0.00615f
C2820 vdd.n1753 gnd 0.00615f
C2821 vdd.n1755 gnd 0.00615f
C2822 vdd.n1756 gnd 0.00615f
C2823 vdd.n1757 gnd 0.00615f
C2824 vdd.n1758 gnd 0.00615f
C2825 vdd.n1759 gnd 0.00615f
C2826 vdd.n1760 gnd 0.00615f
C2827 vdd.n1761 gnd 0.00615f
C2828 vdd.n1762 gnd 0.00615f
C2829 vdd.n1763 gnd 0.004477f
C2830 vdd.n1764 gnd 0.00615f
C2831 vdd.t95 gnd 0.248519f
C2832 vdd.t96 gnd 0.25439f
C2833 vdd.t94 gnd 0.162243f
C2834 vdd.n1765 gnd 0.087683f
C2835 vdd.n1766 gnd 0.049737f
C2836 vdd.n1767 gnd 0.008789f
C2837 vdd.n1768 gnd 0.00615f
C2838 vdd.n1769 gnd 0.00615f
C2839 vdd.n1770 gnd 0.374325f
C2840 vdd.n1771 gnd 0.00615f
C2841 vdd.n1772 gnd 0.00615f
C2842 vdd.n1773 gnd 0.00615f
C2843 vdd.n1774 gnd 0.00615f
C2844 vdd.n1775 gnd 0.00615f
C2845 vdd.n1776 gnd 0.00615f
C2846 vdd.n1777 gnd 0.00615f
C2847 vdd.n1778 gnd 0.00615f
C2848 vdd.n1779 gnd 0.00615f
C2849 vdd.n1780 gnd 0.00615f
C2850 vdd.n1781 gnd 0.00615f
C2851 vdd.n1782 gnd 0.00615f
C2852 vdd.n1783 gnd 0.00615f
C2853 vdd.n1784 gnd 0.00615f
C2854 vdd.n1785 gnd 0.00615f
C2855 vdd.n1786 gnd 0.00615f
C2856 vdd.n1787 gnd 0.00615f
C2857 vdd.n1788 gnd 0.00615f
C2858 vdd.n1789 gnd 0.00615f
C2859 vdd.n1790 gnd 0.00615f
C2860 vdd.t70 gnd 0.248519f
C2861 vdd.t71 gnd 0.25439f
C2862 vdd.t68 gnd 0.162243f
C2863 vdd.n1791 gnd 0.087683f
C2864 vdd.n1792 gnd 0.049737f
C2865 vdd.n1793 gnd 0.00615f
C2866 vdd.n1794 gnd 0.00615f
C2867 vdd.n1795 gnd 0.00615f
C2868 vdd.n1796 gnd 0.00615f
C2869 vdd.n1797 gnd 0.00615f
C2870 vdd.n1798 gnd 0.00615f
C2871 vdd.n1800 gnd 0.00615f
C2872 vdd.n1801 gnd 0.00615f
C2873 vdd.n1802 gnd 0.00615f
C2874 vdd.n1803 gnd 0.00615f
C2875 vdd.n1805 gnd 0.00615f
C2876 vdd.n1807 gnd 0.00615f
C2877 vdd.n1808 gnd 0.00615f
C2878 vdd.n1809 gnd 0.00615f
C2879 vdd.n1810 gnd 0.00615f
C2880 vdd.n1811 gnd 0.00615f
C2881 vdd.n1813 gnd 0.00615f
C2882 vdd.n1815 gnd 0.00615f
C2883 vdd.n1816 gnd 0.00615f
C2884 vdd.n1817 gnd 0.00615f
C2885 vdd.n1818 gnd 0.00615f
C2886 vdd.n1819 gnd 0.00615f
C2887 vdd.n1821 gnd 0.00615f
C2888 vdd.n1823 gnd 0.00615f
C2889 vdd.n1824 gnd 0.00615f
C2890 vdd.n1825 gnd 0.004477f
C2891 vdd.n1826 gnd 0.008789f
C2892 vdd.n1827 gnd 0.004748f
C2893 vdd.n1828 gnd 0.00615f
C2894 vdd.n1830 gnd 0.00615f
C2895 vdd.n1831 gnd 0.014593f
C2896 vdd.n1832 gnd 0.014593f
C2897 vdd.n1833 gnd 0.013625f
C2898 vdd.n1834 gnd 0.00615f
C2899 vdd.n1835 gnd 0.00615f
C2900 vdd.n1836 gnd 0.00615f
C2901 vdd.n1837 gnd 0.00615f
C2902 vdd.n1838 gnd 0.00615f
C2903 vdd.n1839 gnd 0.00615f
C2904 vdd.n1840 gnd 0.00615f
C2905 vdd.n1841 gnd 0.00615f
C2906 vdd.n1842 gnd 0.00615f
C2907 vdd.n1843 gnd 0.00615f
C2908 vdd.n1844 gnd 0.00615f
C2909 vdd.n1845 gnd 0.00615f
C2910 vdd.n1846 gnd 0.00615f
C2911 vdd.n1847 gnd 0.00615f
C2912 vdd.n1848 gnd 0.00615f
C2913 vdd.n1849 gnd 0.00615f
C2914 vdd.n1850 gnd 0.00615f
C2915 vdd.n1851 gnd 0.00615f
C2916 vdd.n1852 gnd 0.00615f
C2917 vdd.n1853 gnd 0.00615f
C2918 vdd.n1854 gnd 0.00615f
C2919 vdd.n1855 gnd 0.00615f
C2920 vdd.n1856 gnd 0.00615f
C2921 vdd.n1857 gnd 0.00615f
C2922 vdd.n1858 gnd 0.00615f
C2923 vdd.n1859 gnd 0.00615f
C2924 vdd.n1860 gnd 0.00615f
C2925 vdd.n1861 gnd 0.00615f
C2926 vdd.n1862 gnd 0.00615f
C2927 vdd.n1863 gnd 0.00615f
C2928 vdd.n1864 gnd 0.00615f
C2929 vdd.n1865 gnd 0.00615f
C2930 vdd.n1866 gnd 0.00615f
C2931 vdd.n1867 gnd 0.00615f
C2932 vdd.n1868 gnd 0.00615f
C2933 vdd.n1869 gnd 0.00615f
C2934 vdd.n1870 gnd 0.00615f
C2935 vdd.n1871 gnd 0.198716f
C2936 vdd.n1872 gnd 0.00615f
C2937 vdd.n1873 gnd 0.00615f
C2938 vdd.n1874 gnd 0.00615f
C2939 vdd.n1875 gnd 0.00615f
C2940 vdd.n1876 gnd 0.00615f
C2941 vdd.n1877 gnd 0.00615f
C2942 vdd.n1878 gnd 0.00615f
C2943 vdd.n1879 gnd 0.00615f
C2944 vdd.n1880 gnd 0.00615f
C2945 vdd.n1881 gnd 0.00615f
C2946 vdd.n1882 gnd 0.00615f
C2947 vdd.n1883 gnd 0.00615f
C2948 vdd.n1884 gnd 0.00615f
C2949 vdd.n1885 gnd 0.00615f
C2950 vdd.n1886 gnd 0.00615f
C2951 vdd.n1887 gnd 0.00615f
C2952 vdd.n1888 gnd 0.00615f
C2953 vdd.n1889 gnd 0.00615f
C2954 vdd.n1890 gnd 0.00615f
C2955 vdd.n1891 gnd 0.00615f
C2956 vdd.n1892 gnd 0.013625f
C2957 vdd.n1894 gnd 0.014593f
C2958 vdd.n1895 gnd 0.014593f
C2959 vdd.n1896 gnd 0.00615f
C2960 vdd.n1897 gnd 0.004748f
C2961 vdd.n1898 gnd 0.00615f
C2962 vdd.n1900 gnd 0.00615f
C2963 vdd.n1902 gnd 0.00615f
C2964 vdd.n1903 gnd 0.00615f
C2965 vdd.n1904 gnd 0.00615f
C2966 vdd.n1905 gnd 0.00615f
C2967 vdd.n1906 gnd 0.00615f
C2968 vdd.n1908 gnd 0.00615f
C2969 vdd.n1910 gnd 0.00615f
C2970 vdd.n1911 gnd 0.00615f
C2971 vdd.n1912 gnd 0.00615f
C2972 vdd.n1913 gnd 0.00615f
C2973 vdd.n1914 gnd 0.00615f
C2974 vdd.n1916 gnd 0.00615f
C2975 vdd.n1918 gnd 0.00615f
C2976 vdd.n1919 gnd 0.00615f
C2977 vdd.n1920 gnd 0.00615f
C2978 vdd.n1921 gnd 0.00615f
C2979 vdd.n1922 gnd 0.00615f
C2980 vdd.n1924 gnd 0.00615f
C2981 vdd.n1926 gnd 0.00615f
C2982 vdd.n1927 gnd 0.00615f
C2983 vdd.n1928 gnd 0.018344f
C2984 vdd.n1929 gnd 0.543796f
C2985 vdd.n1931 gnd 0.007279f
C2986 vdd.n1932 gnd 0.007279f
C2987 vdd.n1933 gnd 0.009044f
C2988 vdd.n1935 gnd 0.009044f
C2989 vdd.n1936 gnd 0.009044f
C2990 vdd.n1937 gnd 0.007279f
C2991 vdd.n1938 gnd 0.006042f
C2992 vdd.n1939 gnd 0.022546f
C2993 vdd.n1940 gnd 0.022041f
C2994 vdd.n1941 gnd 0.006042f
C2995 vdd.n1942 gnd 0.022041f
C2996 vdd.n1943 gnd 1.27086f
C2997 vdd.n1944 gnd 0.022041f
C2998 vdd.n1945 gnd 0.022546f
C2999 vdd.n1946 gnd 0.003458f
C3000 vdd.t31 gnd 0.111266f
C3001 vdd.t30 gnd 0.118912f
C3002 vdd.t28 gnd 0.145312f
C3003 vdd.n1947 gnd 0.186269f
C3004 vdd.n1948 gnd 0.1565f
C3005 vdd.n1949 gnd 0.01121f
C3006 vdd.n1950 gnd 0.003822f
C3007 vdd.n1951 gnd 0.007778f
C3008 vdd.n1952 gnd 0.543796f
C3009 vdd.n1953 gnd 0.018344f
C3010 vdd.n1954 gnd 0.00615f
C3011 vdd.n1955 gnd 0.00615f
C3012 vdd.n1956 gnd 0.00615f
C3013 vdd.n1958 gnd 0.00615f
C3014 vdd.n1960 gnd 0.00615f
C3015 vdd.n1961 gnd 0.00615f
C3016 vdd.n1962 gnd 0.00615f
C3017 vdd.n1963 gnd 0.00615f
C3018 vdd.n1964 gnd 0.00615f
C3019 vdd.n1966 gnd 0.00615f
C3020 vdd.n1968 gnd 0.00615f
C3021 vdd.n1969 gnd 0.00615f
C3022 vdd.n1970 gnd 0.00615f
C3023 vdd.n1971 gnd 0.00615f
C3024 vdd.n1972 gnd 0.00615f
C3025 vdd.n1974 gnd 0.00615f
C3026 vdd.n1976 gnd 0.00615f
C3027 vdd.n1977 gnd 0.00615f
C3028 vdd.n1978 gnd 0.00615f
C3029 vdd.n1979 gnd 0.00615f
C3030 vdd.n1980 gnd 0.00615f
C3031 vdd.n1982 gnd 0.00615f
C3032 vdd.n1984 gnd 0.00615f
C3033 vdd.n1985 gnd 0.00615f
C3034 vdd.n1986 gnd 0.014593f
C3035 vdd.n1987 gnd 0.013625f
C3036 vdd.n1988 gnd 0.013625f
C3037 vdd.n1989 gnd 0.905775f
C3038 vdd.n1990 gnd 0.013625f
C3039 vdd.n1991 gnd 0.013625f
C3040 vdd.n1992 gnd 0.00615f
C3041 vdd.n1993 gnd 0.00615f
C3042 vdd.n1994 gnd 0.00615f
C3043 vdd.n1995 gnd 0.39281f
C3044 vdd.n1996 gnd 0.00615f
C3045 vdd.n1997 gnd 0.00615f
C3046 vdd.n1998 gnd 0.00615f
C3047 vdd.n1999 gnd 0.00615f
C3048 vdd.n2000 gnd 0.00615f
C3049 vdd.n2001 gnd 0.628497f
C3050 vdd.n2002 gnd 0.00615f
C3051 vdd.n2003 gnd 0.00615f
C3052 vdd.n2004 gnd 0.00615f
C3053 vdd.n2005 gnd 0.00615f
C3054 vdd.n2006 gnd 0.00615f
C3055 vdd.n2007 gnd 0.628497f
C3056 vdd.n2008 gnd 0.00615f
C3057 vdd.n2009 gnd 0.00615f
C3058 vdd.n2010 gnd 0.005426f
C3059 vdd.n2011 gnd 0.017816f
C3060 vdd.n2012 gnd 0.003799f
C3061 vdd.n2013 gnd 0.00615f
C3062 vdd.n2014 gnd 0.346597f
C3063 vdd.n2015 gnd 0.00615f
C3064 vdd.n2016 gnd 0.00615f
C3065 vdd.n2017 gnd 0.00615f
C3066 vdd.n2018 gnd 0.00615f
C3067 vdd.n2019 gnd 0.00615f
C3068 vdd.n2020 gnd 0.420538f
C3069 vdd.n2021 gnd 0.00615f
C3070 vdd.n2022 gnd 0.00615f
C3071 vdd.n2023 gnd 0.00615f
C3072 vdd.n2024 gnd 0.00615f
C3073 vdd.n2025 gnd 0.00615f
C3074 vdd.n2026 gnd 0.559177f
C3075 vdd.n2027 gnd 0.00615f
C3076 vdd.n2028 gnd 0.00615f
C3077 vdd.n2029 gnd 0.00615f
C3078 vdd.n2030 gnd 0.00615f
C3079 vdd.n2031 gnd 0.00615f
C3080 vdd.n2032 gnd 0.4991f
C3081 vdd.n2033 gnd 0.00615f
C3082 vdd.n2034 gnd 0.00615f
C3083 vdd.n2035 gnd 0.00615f
C3084 vdd.n2036 gnd 0.00615f
C3085 vdd.n2037 gnd 0.00615f
C3086 vdd.n2038 gnd 0.360461f
C3087 vdd.n2039 gnd 0.00615f
C3088 vdd.n2040 gnd 0.00615f
C3089 vdd.n2041 gnd 0.00615f
C3090 vdd.n2042 gnd 0.00615f
C3091 vdd.n2043 gnd 0.00615f
C3092 vdd.n2044 gnd 0.198716f
C3093 vdd.n2045 gnd 0.00615f
C3094 vdd.n2046 gnd 0.00615f
C3095 vdd.n2047 gnd 0.00615f
C3096 vdd.n2048 gnd 0.00615f
C3097 vdd.n2049 gnd 0.00615f
C3098 vdd.n2050 gnd 0.346597f
C3099 vdd.n2051 gnd 0.00615f
C3100 vdd.n2052 gnd 0.00615f
C3101 vdd.n2053 gnd 0.00615f
C3102 vdd.n2054 gnd 0.00615f
C3103 vdd.n2055 gnd 0.00615f
C3104 vdd.n2056 gnd 0.628497f
C3105 vdd.n2057 gnd 0.00615f
C3106 vdd.n2058 gnd 0.00615f
C3107 vdd.n2059 gnd 0.00615f
C3108 vdd.n2060 gnd 0.00615f
C3109 vdd.n2061 gnd 0.00615f
C3110 vdd.n2062 gnd 0.00615f
C3111 vdd.n2063 gnd 0.00615f
C3112 vdd.n2064 gnd 0.489858f
C3113 vdd.n2065 gnd 0.00615f
C3114 vdd.n2066 gnd 0.00615f
C3115 vdd.n2067 gnd 0.00615f
C3116 vdd.n2068 gnd 0.00615f
C3117 vdd.n2069 gnd 0.00615f
C3118 vdd.n2070 gnd 0.00615f
C3119 vdd.n2071 gnd 0.39281f
C3120 vdd.n2072 gnd 0.00615f
C3121 vdd.n2073 gnd 0.00615f
C3122 vdd.n2074 gnd 0.00615f
C3123 vdd.n2075 gnd 0.014374f
C3124 vdd.n2076 gnd 0.013844f
C3125 vdd.n2077 gnd 0.00615f
C3126 vdd.n2078 gnd 0.00615f
C3127 vdd.n2079 gnd 0.004748f
C3128 vdd.n2080 gnd 0.00615f
C3129 vdd.n2081 gnd 0.00615f
C3130 vdd.n2082 gnd 0.004477f
C3131 vdd.n2083 gnd 0.00615f
C3132 vdd.n2084 gnd 0.00615f
C3133 vdd.n2085 gnd 0.00615f
C3134 vdd.n2086 gnd 0.00615f
C3135 vdd.n2087 gnd 0.00615f
C3136 vdd.n2088 gnd 0.00615f
C3137 vdd.n2089 gnd 0.00615f
C3138 vdd.n2090 gnd 0.00615f
C3139 vdd.n2091 gnd 0.00615f
C3140 vdd.n2092 gnd 0.00615f
C3141 vdd.n2093 gnd 0.00615f
C3142 vdd.n2094 gnd 0.00615f
C3143 vdd.n2095 gnd 0.00615f
C3144 vdd.n2096 gnd 0.00615f
C3145 vdd.n2097 gnd 0.00615f
C3146 vdd.n2098 gnd 0.00615f
C3147 vdd.n2099 gnd 0.00615f
C3148 vdd.n2100 gnd 0.00615f
C3149 vdd.n2101 gnd 0.00615f
C3150 vdd.n2102 gnd 0.00615f
C3151 vdd.n2103 gnd 0.00615f
C3152 vdd.n2104 gnd 0.00615f
C3153 vdd.n2105 gnd 0.00615f
C3154 vdd.n2106 gnd 0.00615f
C3155 vdd.n2107 gnd 0.00615f
C3156 vdd.n2108 gnd 0.00615f
C3157 vdd.n2109 gnd 0.00615f
C3158 vdd.n2110 gnd 0.00615f
C3159 vdd.n2111 gnd 0.00615f
C3160 vdd.n2112 gnd 0.00615f
C3161 vdd.n2113 gnd 0.00615f
C3162 vdd.n2114 gnd 0.00615f
C3163 vdd.n2115 gnd 0.00615f
C3164 vdd.n2116 gnd 0.00615f
C3165 vdd.n2117 gnd 0.00615f
C3166 vdd.n2118 gnd 0.00615f
C3167 vdd.n2119 gnd 0.00615f
C3168 vdd.n2120 gnd 0.00615f
C3169 vdd.n2121 gnd 0.00615f
C3170 vdd.n2122 gnd 0.00615f
C3171 vdd.n2123 gnd 0.00615f
C3172 vdd.n2124 gnd 0.00615f
C3173 vdd.n2125 gnd 0.00615f
C3174 vdd.n2126 gnd 0.00615f
C3175 vdd.n2127 gnd 0.00615f
C3176 vdd.n2128 gnd 0.00615f
C3177 vdd.n2129 gnd 0.00615f
C3178 vdd.n2130 gnd 0.00615f
C3179 vdd.n2131 gnd 0.00615f
C3180 vdd.n2132 gnd 0.00615f
C3181 vdd.n2133 gnd 0.00615f
C3182 vdd.n2134 gnd 0.00615f
C3183 vdd.n2135 gnd 0.00615f
C3184 vdd.n2136 gnd 0.00615f
C3185 vdd.n2137 gnd 0.00615f
C3186 vdd.n2138 gnd 0.00615f
C3187 vdd.n2139 gnd 0.00615f
C3188 vdd.n2140 gnd 0.00615f
C3189 vdd.n2141 gnd 0.00615f
C3190 vdd.n2142 gnd 0.00615f
C3191 vdd.n2143 gnd 0.014593f
C3192 vdd.n2144 gnd 0.013625f
C3193 vdd.n2145 gnd 0.013625f
C3194 vdd.n2146 gnd 0.767136f
C3195 vdd.n2147 gnd 0.013625f
C3196 vdd.n2148 gnd 0.014593f
C3197 vdd.n2149 gnd 0.013844f
C3198 vdd.n2150 gnd 0.00615f
C3199 vdd.n2151 gnd 0.00615f
C3200 vdd.n2152 gnd 0.00615f
C3201 vdd.n2153 gnd 0.004748f
C3202 vdd.n2154 gnd 0.008789f
C3203 vdd.n2155 gnd 0.004477f
C3204 vdd.n2156 gnd 0.00615f
C3205 vdd.n2157 gnd 0.00615f
C3206 vdd.n2158 gnd 0.00615f
C3207 vdd.n2159 gnd 0.00615f
C3208 vdd.n2160 gnd 0.00615f
C3209 vdd.n2161 gnd 0.00615f
C3210 vdd.n2162 gnd 0.00615f
C3211 vdd.n2163 gnd 0.00615f
C3212 vdd.n2164 gnd 0.00615f
C3213 vdd.n2165 gnd 0.00615f
C3214 vdd.n2166 gnd 0.00615f
C3215 vdd.n2167 gnd 0.00615f
C3216 vdd.n2168 gnd 0.00615f
C3217 vdd.n2169 gnd 0.00615f
C3218 vdd.n2170 gnd 0.00615f
C3219 vdd.n2171 gnd 0.00615f
C3220 vdd.n2172 gnd 0.00615f
C3221 vdd.n2173 gnd 0.00615f
C3222 vdd.n2174 gnd 0.00615f
C3223 vdd.n2175 gnd 0.00615f
C3224 vdd.n2176 gnd 0.00615f
C3225 vdd.n2177 gnd 0.00615f
C3226 vdd.n2178 gnd 0.00615f
C3227 vdd.n2179 gnd 0.00615f
C3228 vdd.n2180 gnd 0.00615f
C3229 vdd.n2181 gnd 0.00615f
C3230 vdd.n2182 gnd 0.00615f
C3231 vdd.n2183 gnd 0.00615f
C3232 vdd.n2184 gnd 0.00615f
C3233 vdd.n2185 gnd 0.00615f
C3234 vdd.n2186 gnd 0.00615f
C3235 vdd.n2187 gnd 0.00615f
C3236 vdd.n2188 gnd 0.00615f
C3237 vdd.n2189 gnd 0.00615f
C3238 vdd.n2190 gnd 0.00615f
C3239 vdd.n2191 gnd 0.00615f
C3240 vdd.n2192 gnd 0.00615f
C3241 vdd.n2193 gnd 0.00615f
C3242 vdd.n2194 gnd 0.00615f
C3243 vdd.n2195 gnd 0.00615f
C3244 vdd.n2196 gnd 0.00615f
C3245 vdd.n2197 gnd 0.00615f
C3246 vdd.n2198 gnd 0.00615f
C3247 vdd.n2199 gnd 0.00615f
C3248 vdd.n2200 gnd 0.00615f
C3249 vdd.n2201 gnd 0.00615f
C3250 vdd.n2202 gnd 0.00615f
C3251 vdd.n2203 gnd 0.00615f
C3252 vdd.n2204 gnd 0.00615f
C3253 vdd.n2205 gnd 0.00615f
C3254 vdd.n2206 gnd 0.00615f
C3255 vdd.n2207 gnd 0.00615f
C3256 vdd.n2208 gnd 0.00615f
C3257 vdd.n2209 gnd 0.00615f
C3258 vdd.n2210 gnd 0.00615f
C3259 vdd.n2211 gnd 0.00615f
C3260 vdd.n2212 gnd 0.00615f
C3261 vdd.n2213 gnd 0.00615f
C3262 vdd.n2214 gnd 0.00615f
C3263 vdd.n2215 gnd 0.00615f
C3264 vdd.n2216 gnd 0.014593f
C3265 vdd.n2217 gnd 0.014593f
C3266 vdd.n2218 gnd 0.767136f
C3267 vdd.t12 gnd 2.72657f
C3268 vdd.t5 gnd 2.72657f
C3269 vdd.n2251 gnd 0.014593f
C3270 vdd.n2252 gnd 0.00615f
C3271 vdd.t63 gnd 0.248519f
C3272 vdd.t64 gnd 0.25439f
C3273 vdd.t61 gnd 0.162243f
C3274 vdd.n2253 gnd 0.087683f
C3275 vdd.n2254 gnd 0.049737f
C3276 vdd.n2255 gnd 0.00615f
C3277 vdd.t77 gnd 0.248519f
C3278 vdd.t78 gnd 0.25439f
C3279 vdd.t76 gnd 0.162243f
C3280 vdd.n2256 gnd 0.087683f
C3281 vdd.n2257 gnd 0.049737f
C3282 vdd.n2258 gnd 0.008789f
C3283 vdd.n2259 gnd 0.00615f
C3284 vdd.n2260 gnd 0.00615f
C3285 vdd.n2261 gnd 0.00615f
C3286 vdd.n2262 gnd 0.00615f
C3287 vdd.n2263 gnd 0.00615f
C3288 vdd.n2264 gnd 0.00615f
C3289 vdd.n2265 gnd 0.00615f
C3290 vdd.n2266 gnd 0.00615f
C3291 vdd.n2267 gnd 0.00615f
C3292 vdd.n2268 gnd 0.00615f
C3293 vdd.n2269 gnd 0.00615f
C3294 vdd.n2270 gnd 0.00615f
C3295 vdd.n2271 gnd 0.00615f
C3296 vdd.n2272 gnd 0.00615f
C3297 vdd.n2273 gnd 0.00615f
C3298 vdd.n2274 gnd 0.00615f
C3299 vdd.n2275 gnd 0.00615f
C3300 vdd.n2276 gnd 0.00615f
C3301 vdd.n2277 gnd 0.00615f
C3302 vdd.n2278 gnd 0.00615f
C3303 vdd.n2279 gnd 0.00615f
C3304 vdd.n2280 gnd 0.00615f
C3305 vdd.n2281 gnd 0.00615f
C3306 vdd.n2282 gnd 0.00615f
C3307 vdd.n2283 gnd 0.00615f
C3308 vdd.n2284 gnd 0.00615f
C3309 vdd.n2285 gnd 0.00615f
C3310 vdd.n2286 gnd 0.00615f
C3311 vdd.n2287 gnd 0.00615f
C3312 vdd.n2288 gnd 0.00615f
C3313 vdd.n2289 gnd 0.00615f
C3314 vdd.n2290 gnd 0.00615f
C3315 vdd.n2291 gnd 0.00615f
C3316 vdd.n2292 gnd 0.00615f
C3317 vdd.n2293 gnd 0.00615f
C3318 vdd.n2294 gnd 0.00615f
C3319 vdd.n2295 gnd 0.00615f
C3320 vdd.n2296 gnd 0.00615f
C3321 vdd.n2297 gnd 0.00615f
C3322 vdd.n2298 gnd 0.00615f
C3323 vdd.n2299 gnd 0.00615f
C3324 vdd.n2300 gnd 0.00615f
C3325 vdd.n2301 gnd 0.00615f
C3326 vdd.n2302 gnd 0.00615f
C3327 vdd.n2303 gnd 0.00615f
C3328 vdd.n2304 gnd 0.00615f
C3329 vdd.n2305 gnd 0.00615f
C3330 vdd.n2306 gnd 0.00615f
C3331 vdd.n2307 gnd 0.00615f
C3332 vdd.n2308 gnd 0.00615f
C3333 vdd.n2309 gnd 0.00615f
C3334 vdd.n2310 gnd 0.00615f
C3335 vdd.n2311 gnd 0.00615f
C3336 vdd.n2312 gnd 0.00615f
C3337 vdd.n2313 gnd 0.00615f
C3338 vdd.n2314 gnd 0.00615f
C3339 vdd.n2315 gnd 0.004477f
C3340 vdd.n2316 gnd 0.00615f
C3341 vdd.n2317 gnd 0.00615f
C3342 vdd.n2318 gnd 0.004748f
C3343 vdd.n2319 gnd 0.00615f
C3344 vdd.n2320 gnd 0.00615f
C3345 vdd.n2321 gnd 0.014593f
C3346 vdd.n2322 gnd 0.013625f
C3347 vdd.n2323 gnd 0.00615f
C3348 vdd.n2324 gnd 0.00615f
C3349 vdd.n2325 gnd 0.00615f
C3350 vdd.n2326 gnd 0.00615f
C3351 vdd.n2327 gnd 0.00615f
C3352 vdd.n2328 gnd 0.00615f
C3353 vdd.n2329 gnd 0.00615f
C3354 vdd.n2330 gnd 0.00615f
C3355 vdd.n2331 gnd 0.00615f
C3356 vdd.n2332 gnd 0.00615f
C3357 vdd.n2333 gnd 0.00615f
C3358 vdd.n2334 gnd 0.00615f
C3359 vdd.n2335 gnd 0.00615f
C3360 vdd.n2336 gnd 0.00615f
C3361 vdd.n2337 gnd 0.00615f
C3362 vdd.n2338 gnd 0.00615f
C3363 vdd.n2339 gnd 0.00615f
C3364 vdd.n2340 gnd 0.00615f
C3365 vdd.n2341 gnd 0.00615f
C3366 vdd.n2342 gnd 0.00615f
C3367 vdd.n2343 gnd 0.00615f
C3368 vdd.n2344 gnd 0.00615f
C3369 vdd.n2345 gnd 0.00615f
C3370 vdd.n2346 gnd 0.00615f
C3371 vdd.n2347 gnd 0.00615f
C3372 vdd.n2348 gnd 0.00615f
C3373 vdd.n2349 gnd 0.00615f
C3374 vdd.n2350 gnd 0.00615f
C3375 vdd.n2351 gnd 0.00615f
C3376 vdd.n2352 gnd 0.00615f
C3377 vdd.n2353 gnd 0.00615f
C3378 vdd.n2354 gnd 0.00615f
C3379 vdd.n2355 gnd 0.00615f
C3380 vdd.n2356 gnd 0.00615f
C3381 vdd.n2357 gnd 0.00615f
C3382 vdd.n2358 gnd 0.00615f
C3383 vdd.n2359 gnd 0.00615f
C3384 vdd.n2360 gnd 0.00615f
C3385 vdd.n2361 gnd 0.00615f
C3386 vdd.n2362 gnd 0.00615f
C3387 vdd.n2363 gnd 0.00615f
C3388 vdd.n2364 gnd 0.00615f
C3389 vdd.n2365 gnd 0.00615f
C3390 vdd.n2366 gnd 0.00615f
C3391 vdd.n2367 gnd 0.00615f
C3392 vdd.n2368 gnd 0.00615f
C3393 vdd.n2369 gnd 0.00615f
C3394 vdd.n2370 gnd 0.00615f
C3395 vdd.n2371 gnd 0.00615f
C3396 vdd.n2372 gnd 0.00615f
C3397 vdd.n2373 gnd 0.00615f
C3398 vdd.n2374 gnd 0.198716f
C3399 vdd.n2375 gnd 0.00615f
C3400 vdd.n2376 gnd 0.00615f
C3401 vdd.n2377 gnd 0.00615f
C3402 vdd.n2378 gnd 0.00615f
C3403 vdd.n2379 gnd 0.00615f
C3404 vdd.n2380 gnd 0.00615f
C3405 vdd.n2381 gnd 0.00615f
C3406 vdd.n2382 gnd 0.00615f
C3407 vdd.n2383 gnd 0.00615f
C3408 vdd.n2384 gnd 0.00615f
C3409 vdd.n2385 gnd 0.00615f
C3410 vdd.n2386 gnd 0.00615f
C3411 vdd.n2387 gnd 0.00615f
C3412 vdd.n2388 gnd 0.00615f
C3413 vdd.n2389 gnd 0.00615f
C3414 vdd.n2390 gnd 0.00615f
C3415 vdd.n2391 gnd 0.00615f
C3416 vdd.n2392 gnd 0.00615f
C3417 vdd.n2393 gnd 0.00615f
C3418 vdd.n2394 gnd 0.00615f
C3419 vdd.n2395 gnd 0.374325f
C3420 vdd.n2396 gnd 0.00615f
C3421 vdd.n2397 gnd 0.00615f
C3422 vdd.n2398 gnd 0.00615f
C3423 vdd.n2399 gnd 0.00615f
C3424 vdd.n2400 gnd 0.00615f
C3425 vdd.n2401 gnd 0.013625f
C3426 vdd.n2402 gnd 0.014593f
C3427 vdd.n2403 gnd 0.014593f
C3428 vdd.n2404 gnd 0.00615f
C3429 vdd.n2405 gnd 0.00615f
C3430 vdd.n2406 gnd 0.00615f
C3431 vdd.n2407 gnd 0.004748f
C3432 vdd.n2408 gnd 0.008789f
C3433 vdd.n2409 gnd 0.004477f
C3434 vdd.n2410 gnd 0.00615f
C3435 vdd.n2411 gnd 0.00615f
C3436 vdd.n2412 gnd 0.00615f
C3437 vdd.n2413 gnd 0.00615f
C3438 vdd.n2414 gnd 0.00615f
C3439 vdd.n2415 gnd 0.00615f
C3440 vdd.n2416 gnd 0.00615f
C3441 vdd.n2417 gnd 0.00615f
C3442 vdd.n2418 gnd 0.00615f
C3443 vdd.n2419 gnd 0.00615f
C3444 vdd.n2420 gnd 0.00615f
C3445 vdd.n2421 gnd 0.00615f
C3446 vdd.n2422 gnd 0.00615f
C3447 vdd.n2423 gnd 0.00615f
C3448 vdd.n2424 gnd 0.00615f
C3449 vdd.n2425 gnd 0.00615f
C3450 vdd.n2426 gnd 0.00615f
C3451 vdd.n2427 gnd 0.00615f
C3452 vdd.n2428 gnd 0.00615f
C3453 vdd.n2429 gnd 0.00615f
C3454 vdd.n2430 gnd 0.00615f
C3455 vdd.n2431 gnd 0.00615f
C3456 vdd.n2432 gnd 0.00615f
C3457 vdd.n2433 gnd 0.00615f
C3458 vdd.n2434 gnd 0.00615f
C3459 vdd.n2435 gnd 0.00615f
C3460 vdd.n2436 gnd 0.00615f
C3461 vdd.n2437 gnd 0.00615f
C3462 vdd.n2438 gnd 0.00615f
C3463 vdd.n2439 gnd 0.00615f
C3464 vdd.n2440 gnd 0.00615f
C3465 vdd.n2441 gnd 0.00615f
C3466 vdd.n2442 gnd 0.00615f
C3467 vdd.n2443 gnd 0.00615f
C3468 vdd.n2444 gnd 0.00615f
C3469 vdd.n2445 gnd 0.00615f
C3470 vdd.n2446 gnd 0.00615f
C3471 vdd.n2447 gnd 0.00615f
C3472 vdd.n2448 gnd 0.00615f
C3473 vdd.n2449 gnd 0.00615f
C3474 vdd.n2450 gnd 0.00615f
C3475 vdd.n2451 gnd 0.00615f
C3476 vdd.n2452 gnd 0.00615f
C3477 vdd.n2453 gnd 0.00615f
C3478 vdd.n2454 gnd 0.00615f
C3479 vdd.n2455 gnd 0.00615f
C3480 vdd.n2456 gnd 0.00615f
C3481 vdd.n2457 gnd 0.00615f
C3482 vdd.n2458 gnd 0.00615f
C3483 vdd.n2459 gnd 0.00615f
C3484 vdd.n2460 gnd 0.00615f
C3485 vdd.n2461 gnd 0.00615f
C3486 vdd.n2462 gnd 0.00615f
C3487 vdd.n2463 gnd 0.00615f
C3488 vdd.n2464 gnd 0.00615f
C3489 vdd.n2465 gnd 0.00615f
C3490 vdd.n2466 gnd 0.00615f
C3491 vdd.n2467 gnd 0.00615f
C3492 vdd.n2468 gnd 0.00615f
C3493 vdd.n2469 gnd 0.00615f
C3494 vdd.n2471 gnd 0.767136f
C3495 vdd.n2473 gnd 0.00615f
C3496 vdd.n2474 gnd 0.00615f
C3497 vdd.n2475 gnd 0.014593f
C3498 vdd.n2476 gnd 0.013625f
C3499 vdd.n2477 gnd 0.013625f
C3500 vdd.n2478 gnd 0.767136f
C3501 vdd.n2479 gnd 0.013625f
C3502 vdd.n2480 gnd 0.013625f
C3503 vdd.n2481 gnd 0.00615f
C3504 vdd.n2482 gnd 0.00615f
C3505 vdd.n2483 gnd 0.00615f
C3506 vdd.n2484 gnd 0.39281f
C3507 vdd.n2485 gnd 0.00615f
C3508 vdd.n2486 gnd 0.00615f
C3509 vdd.n2487 gnd 0.00615f
C3510 vdd.n2488 gnd 0.00615f
C3511 vdd.n2489 gnd 0.00615f
C3512 vdd.n2490 gnd 0.489858f
C3513 vdd.n2491 gnd 0.00615f
C3514 vdd.n2492 gnd 0.00615f
C3515 vdd.n2493 gnd 0.00615f
C3516 vdd.n2494 gnd 0.00615f
C3517 vdd.n2495 gnd 0.00615f
C3518 vdd.n2496 gnd 0.628497f
C3519 vdd.n2497 gnd 0.00615f
C3520 vdd.n2498 gnd 0.00615f
C3521 vdd.n2499 gnd 0.00615f
C3522 vdd.n2500 gnd 0.00615f
C3523 vdd.n2501 gnd 0.00615f
C3524 vdd.n2502 gnd 0.346597f
C3525 vdd.n2503 gnd 0.00615f
C3526 vdd.n2504 gnd 0.00615f
C3527 vdd.n2505 gnd 0.00615f
C3528 vdd.n2506 gnd 0.00615f
C3529 vdd.n2507 gnd 0.00615f
C3530 vdd.n2508 gnd 0.198716f
C3531 vdd.n2509 gnd 0.00615f
C3532 vdd.n2510 gnd 0.00615f
C3533 vdd.n2511 gnd 0.00615f
C3534 vdd.n2512 gnd 0.00615f
C3535 vdd.n2513 gnd 0.00615f
C3536 vdd.n2514 gnd 0.360461f
C3537 vdd.n2515 gnd 0.00615f
C3538 vdd.n2516 gnd 0.00615f
C3539 vdd.n2517 gnd 0.00615f
C3540 vdd.n2518 gnd 0.00615f
C3541 vdd.n2519 gnd 0.00615f
C3542 vdd.n2520 gnd 0.4991f
C3543 vdd.n2521 gnd 0.00615f
C3544 vdd.n2522 gnd 0.00615f
C3545 vdd.n2523 gnd 0.00615f
C3546 vdd.n2524 gnd 0.00615f
C3547 vdd.n2525 gnd 0.00615f
C3548 vdd.n2526 gnd 0.559177f
C3549 vdd.n2527 gnd 0.00615f
C3550 vdd.n2528 gnd 0.00615f
C3551 vdd.n2529 gnd 0.00615f
C3552 vdd.n2530 gnd 0.00615f
C3553 vdd.n2531 gnd 0.00615f
C3554 vdd.n2532 gnd 0.420538f
C3555 vdd.n2533 gnd 0.00615f
C3556 vdd.n2534 gnd 0.00615f
C3557 vdd.n2535 gnd 0.00615f
C3558 vdd.t38 gnd 0.25439f
C3559 vdd.t36 gnd 0.162243f
C3560 vdd.t39 gnd 0.25439f
C3561 vdd.n2536 gnd 0.142978f
C3562 vdd.n2537 gnd 0.017816f
C3563 vdd.n2538 gnd 0.003799f
C3564 vdd.n2539 gnd 0.00615f
C3565 vdd.n2540 gnd 0.346597f
C3566 vdd.n2541 gnd 0.00615f
C3567 vdd.n2542 gnd 0.00615f
C3568 vdd.n2543 gnd 0.00615f
C3569 vdd.n2544 gnd 0.00615f
C3570 vdd.n2545 gnd 0.00615f
C3571 vdd.n2546 gnd 0.628497f
C3572 vdd.n2547 gnd 0.00615f
C3573 vdd.n2548 gnd 0.00615f
C3574 vdd.n2549 gnd 0.00615f
C3575 vdd.n2550 gnd 0.00615f
C3576 vdd.n2551 gnd 0.00615f
C3577 vdd.n2552 gnd 0.00615f
C3578 vdd.n2554 gnd 0.00615f
C3579 vdd.n2555 gnd 0.00615f
C3580 vdd.n2557 gnd 0.00615f
C3581 vdd.n2558 gnd 0.00615f
C3582 vdd.n2561 gnd 0.00615f
C3583 vdd.n2562 gnd 0.00615f
C3584 vdd.n2563 gnd 0.00615f
C3585 vdd.n2564 gnd 0.00615f
C3586 vdd.n2566 gnd 0.00615f
C3587 vdd.n2567 gnd 0.00615f
C3588 vdd.n2568 gnd 0.00615f
C3589 vdd.n2569 gnd 0.00615f
C3590 vdd.n2570 gnd 0.00615f
C3591 vdd.n2571 gnd 0.00615f
C3592 vdd.n2573 gnd 0.00615f
C3593 vdd.n2574 gnd 0.00615f
C3594 vdd.n2575 gnd 0.00615f
C3595 vdd.n2576 gnd 0.00615f
C3596 vdd.n2577 gnd 0.00615f
C3597 vdd.n2578 gnd 0.00615f
C3598 vdd.n2580 gnd 0.00615f
C3599 vdd.n2581 gnd 0.00615f
C3600 vdd.n2582 gnd 0.00615f
C3601 vdd.n2583 gnd 0.00615f
C3602 vdd.n2584 gnd 0.00615f
C3603 vdd.n2585 gnd 0.00615f
C3604 vdd.n2587 gnd 0.00615f
C3605 vdd.n2588 gnd 0.014593f
C3606 vdd.n2589 gnd 0.014593f
C3607 vdd.n2590 gnd 0.013625f
C3608 vdd.n2591 gnd 0.00615f
C3609 vdd.n2592 gnd 0.00615f
C3610 vdd.n2593 gnd 0.00615f
C3611 vdd.n2594 gnd 0.00615f
C3612 vdd.n2595 gnd 0.00615f
C3613 vdd.n2596 gnd 0.00615f
C3614 vdd.n2597 gnd 0.628497f
C3615 vdd.n2598 gnd 0.00615f
C3616 vdd.n2599 gnd 0.00615f
C3617 vdd.n2600 gnd 0.00615f
C3618 vdd.n2601 gnd 0.00615f
C3619 vdd.n2602 gnd 0.00615f
C3620 vdd.n2603 gnd 0.39281f
C3621 vdd.n2604 gnd 0.00615f
C3622 vdd.n2605 gnd 0.00615f
C3623 vdd.n2606 gnd 0.00615f
C3624 vdd.n2607 gnd 0.014374f
C3625 vdd.n2608 gnd 0.013844f
C3626 vdd.n2609 gnd 0.014593f
C3627 vdd.n2611 gnd 0.00615f
C3628 vdd.n2612 gnd 0.00615f
C3629 vdd.n2613 gnd 0.004748f
C3630 vdd.n2614 gnd 0.008789f
C3631 vdd.n2615 gnd 0.004477f
C3632 vdd.n2616 gnd 0.00615f
C3633 vdd.n2617 gnd 0.00615f
C3634 vdd.n2619 gnd 0.00615f
C3635 vdd.n2620 gnd 0.00615f
C3636 vdd.n2621 gnd 0.00615f
C3637 vdd.n2622 gnd 0.00615f
C3638 vdd.n2623 gnd 0.00615f
C3639 vdd.n2624 gnd 0.00615f
C3640 vdd.n2626 gnd 0.00615f
C3641 vdd.n2627 gnd 0.00615f
C3642 vdd.n2628 gnd 0.00615f
C3643 vdd.n2629 gnd 0.00615f
C3644 vdd.n2630 gnd 0.00615f
C3645 vdd.n2631 gnd 0.00615f
C3646 vdd.n2633 gnd 0.00615f
C3647 vdd.n2634 gnd 0.00615f
C3648 vdd.n2635 gnd 0.00615f
C3649 vdd.n2636 gnd 0.00615f
C3650 vdd.n2637 gnd 0.00615f
C3651 vdd.n2638 gnd 0.00615f
C3652 vdd.n2640 gnd 0.00615f
C3653 vdd.n2641 gnd 0.00615f
C3654 vdd.n2642 gnd 0.00615f
C3655 vdd.n2644 gnd 0.00615f
C3656 vdd.n2645 gnd 0.00615f
C3657 vdd.n2646 gnd 0.00615f
C3658 vdd.n2647 gnd 0.00615f
C3659 vdd.n2648 gnd 0.00615f
C3660 vdd.n2649 gnd 0.00615f
C3661 vdd.n2651 gnd 0.00615f
C3662 vdd.n2652 gnd 0.00615f
C3663 vdd.n2653 gnd 0.00615f
C3664 vdd.n2654 gnd 0.00615f
C3665 vdd.n2655 gnd 0.00615f
C3666 vdd.n2656 gnd 0.00615f
C3667 vdd.n2658 gnd 0.00615f
C3668 vdd.n2659 gnd 0.00615f
C3669 vdd.n2660 gnd 0.00615f
C3670 vdd.n2661 gnd 0.00615f
C3671 vdd.n2662 gnd 0.00615f
C3672 vdd.n2663 gnd 0.00615f
C3673 vdd.n2665 gnd 0.00615f
C3674 vdd.n2666 gnd 0.00615f
C3675 vdd.n2668 gnd 0.00615f
C3676 vdd.n2669 gnd 0.00615f
C3677 vdd.n2670 gnd 0.014593f
C3678 vdd.n2671 gnd 0.013625f
C3679 vdd.n2672 gnd 0.013625f
C3680 vdd.n2673 gnd 0.905775f
C3681 vdd.n2674 gnd 0.013625f
C3682 vdd.n2675 gnd 0.014593f
C3683 vdd.n2676 gnd 0.013844f
C3684 vdd.n2677 gnd 0.00615f
C3685 vdd.n2678 gnd 0.004748f
C3686 vdd.n2679 gnd 0.00615f
C3687 vdd.n2681 gnd 0.00615f
C3688 vdd.n2682 gnd 0.00615f
C3689 vdd.n2683 gnd 0.00615f
C3690 vdd.n2684 gnd 0.00615f
C3691 vdd.n2685 gnd 0.00615f
C3692 vdd.n2686 gnd 0.00615f
C3693 vdd.n2688 gnd 0.00615f
C3694 vdd.n2689 gnd 0.00615f
C3695 vdd.n2690 gnd 0.00615f
C3696 vdd.n2691 gnd 0.00615f
C3697 vdd.n2692 gnd 0.00615f
C3698 vdd.n2693 gnd 0.00615f
C3699 vdd.n2695 gnd 0.00615f
C3700 vdd.n2696 gnd 0.00615f
C3701 vdd.n2697 gnd 0.00615f
C3702 vdd.n2698 gnd 0.00615f
C3703 vdd.n2699 gnd 0.00615f
C3704 vdd.n2700 gnd 0.00615f
C3705 vdd.n2702 gnd 0.00615f
C3706 vdd.n2703 gnd 0.00615f
C3707 vdd.n2705 gnd 0.00615f
C3708 vdd.n2706 gnd 0.014779f
C3709 vdd.n2707 gnd 0.547361f
C3710 vdd.n2708 gnd 0.007778f
C3711 vdd.n2709 gnd 0.022546f
C3712 vdd.n2710 gnd 0.003458f
C3713 vdd.t89 gnd 0.111266f
C3714 vdd.t90 gnd 0.118912f
C3715 vdd.t88 gnd 0.145312f
C3716 vdd.n2711 gnd 0.186269f
C3717 vdd.n2712 gnd 0.1565f
C3718 vdd.n2713 gnd 0.01121f
C3719 vdd.n2714 gnd 0.009044f
C3720 vdd.n2715 gnd 0.003822f
C3721 vdd.n2716 gnd 0.007279f
C3722 vdd.n2717 gnd 0.009044f
C3723 vdd.n2718 gnd 0.009044f
C3724 vdd.n2719 gnd 0.007279f
C3725 vdd.n2720 gnd 0.007279f
C3726 vdd.n2721 gnd 0.009044f
C3727 vdd.n2722 gnd 0.009044f
C3728 vdd.n2723 gnd 0.007279f
C3729 vdd.n2724 gnd 0.007279f
C3730 vdd.n2725 gnd 0.009044f
C3731 vdd.n2726 gnd 0.009044f
C3732 vdd.n2727 gnd 0.007279f
C3733 vdd.n2728 gnd 0.007279f
C3734 vdd.n2729 gnd 0.009044f
C3735 vdd.n2730 gnd 0.009044f
C3736 vdd.n2731 gnd 0.007279f
C3737 vdd.n2732 gnd 0.007279f
C3738 vdd.n2733 gnd 0.009044f
C3739 vdd.n2734 gnd 0.009044f
C3740 vdd.n2735 gnd 0.007279f
C3741 vdd.n2736 gnd 0.007279f
C3742 vdd.n2737 gnd 0.009044f
C3743 vdd.n2738 gnd 0.009044f
C3744 vdd.n2739 gnd 0.007279f
C3745 vdd.n2740 gnd 0.007279f
C3746 vdd.n2741 gnd 0.009044f
C3747 vdd.n2742 gnd 0.009044f
C3748 vdd.n2743 gnd 0.007279f
C3749 vdd.n2744 gnd 0.007279f
C3750 vdd.n2745 gnd 0.009044f
C3751 vdd.n2746 gnd 0.009044f
C3752 vdd.n2747 gnd 0.007279f
C3753 vdd.n2748 gnd 0.007279f
C3754 vdd.n2749 gnd 0.009044f
C3755 vdd.n2750 gnd 0.009044f
C3756 vdd.n2751 gnd 0.007279f
C3757 vdd.n2752 gnd 0.009044f
C3758 vdd.n2753 gnd 0.009044f
C3759 vdd.n2754 gnd 0.007279f
C3760 vdd.n2755 gnd 0.009044f
C3761 vdd.n2756 gnd 0.009044f
C3762 vdd.n2757 gnd 0.009044f
C3763 vdd.n2758 gnd 0.01485f
C3764 vdd.n2759 gnd 0.009044f
C3765 vdd.n2760 gnd 0.009044f
C3766 vdd.n2761 gnd 0.00495f
C3767 vdd.n2762 gnd 0.007279f
C3768 vdd.n2763 gnd 0.009044f
C3769 vdd.n2764 gnd 0.009044f
C3770 vdd.n2765 gnd 0.007279f
C3771 vdd.n2766 gnd 0.007279f
C3772 vdd.n2767 gnd 0.009044f
C3773 vdd.n2768 gnd 0.009044f
C3774 vdd.n2769 gnd 0.007279f
C3775 vdd.n2770 gnd 0.007279f
C3776 vdd.n2771 gnd 0.009044f
C3777 vdd.n2772 gnd 0.009044f
C3778 vdd.n2773 gnd 0.007279f
C3779 vdd.n2774 gnd 0.007279f
C3780 vdd.n2775 gnd 0.009044f
C3781 vdd.n2776 gnd 0.009044f
C3782 vdd.n2777 gnd 0.007279f
C3783 vdd.n2778 gnd 0.007279f
C3784 vdd.n2779 gnd 0.009044f
C3785 vdd.n2780 gnd 0.009044f
C3786 vdd.n2781 gnd 0.007279f
C3787 vdd.n2782 gnd 0.007279f
C3788 vdd.n2783 gnd 0.009044f
C3789 vdd.n2784 gnd 0.009044f
C3790 vdd.n2785 gnd 0.007279f
C3791 vdd.n2786 gnd 0.007279f
C3792 vdd.n2787 gnd 0.009044f
C3793 vdd.n2788 gnd 0.009044f
C3794 vdd.n2789 gnd 0.007279f
C3795 vdd.n2790 gnd 0.007279f
C3796 vdd.n2791 gnd 0.009044f
C3797 vdd.n2792 gnd 0.009044f
C3798 vdd.n2793 gnd 0.007279f
C3799 vdd.n2794 gnd 0.007279f
C3800 vdd.n2795 gnd 0.009044f
C3801 vdd.n2796 gnd 0.009044f
C3802 vdd.n2797 gnd 0.007279f
C3803 vdd.n2798 gnd 0.009044f
C3804 vdd.n2799 gnd 0.009044f
C3805 vdd.n2800 gnd 0.007279f
C3806 vdd.n2801 gnd 0.009044f
C3807 vdd.n2802 gnd 0.009044f
C3808 vdd.n2803 gnd 0.009044f
C3809 vdd.t26 gnd 0.111266f
C3810 vdd.t27 gnd 0.118912f
C3811 vdd.t25 gnd 0.145312f
C3812 vdd.n2804 gnd 0.186269f
C3813 vdd.n2805 gnd 0.1565f
C3814 vdd.n2806 gnd 0.01485f
C3815 vdd.n2807 gnd 0.009044f
C3816 vdd.n2808 gnd 0.009044f
C3817 vdd.n2809 gnd 0.006078f
C3818 vdd.n2810 gnd 0.007279f
C3819 vdd.n2811 gnd 0.009044f
C3820 vdd.n2812 gnd 0.009044f
C3821 vdd.n2813 gnd 0.007279f
C3822 vdd.n2814 gnd 0.007279f
C3823 vdd.n2815 gnd 0.009044f
C3824 vdd.n2816 gnd 0.009044f
C3825 vdd.n2817 gnd 0.007279f
C3826 vdd.n2818 gnd 0.007279f
C3827 vdd.n2819 gnd 0.009044f
C3828 vdd.n2820 gnd 0.009044f
C3829 vdd.n2821 gnd 0.007279f
C3830 vdd.n2822 gnd 0.007279f
C3831 vdd.n2823 gnd 0.009044f
C3832 vdd.n2824 gnd 0.009044f
C3833 vdd.n2825 gnd 0.007279f
C3834 vdd.n2826 gnd 0.007279f
C3835 vdd.n2827 gnd 0.009044f
C3836 vdd.n2828 gnd 0.009044f
C3837 vdd.n2829 gnd 0.007279f
C3838 vdd.n2830 gnd 0.007279f
C3839 vdd.n2831 gnd 0.009044f
C3840 vdd.n2832 gnd 0.009044f
C3841 vdd.n2833 gnd 0.007279f
C3842 vdd.n2834 gnd 0.007279f
C3843 vdd.n2836 gnd 0.547361f
C3844 vdd.n2838 gnd 0.007279f
C3845 vdd.n2839 gnd 0.009044f
C3846 vdd.n2840 gnd 6.70088f
C3847 vdd.n2842 gnd 0.022546f
C3848 vdd.n2843 gnd 0.006042f
C3849 vdd.n2844 gnd 0.022546f
C3850 vdd.n2845 gnd 0.022041f
C3851 vdd.n2846 gnd 0.009044f
C3852 vdd.n2847 gnd 0.007279f
C3853 vdd.n2848 gnd 0.009044f
C3854 vdd.n2849 gnd 0.577662f
C3855 vdd.n2850 gnd 0.009044f
C3856 vdd.n2851 gnd 0.007279f
C3857 vdd.n2852 gnd 0.009044f
C3858 vdd.n2853 gnd 0.009044f
C3859 vdd.n2854 gnd 0.009044f
C3860 vdd.n2855 gnd 0.007279f
C3861 vdd.n2856 gnd 0.009044f
C3862 vdd.n2857 gnd 0.734786f
C3863 vdd.n2858 gnd 0.92426f
C3864 vdd.n2859 gnd 0.009044f
C3865 vdd.n2860 gnd 0.007279f
C3866 vdd.n2861 gnd 0.009044f
C3867 vdd.n2862 gnd 0.009044f
C3868 vdd.n2863 gnd 0.009044f
C3869 vdd.n2864 gnd 0.007279f
C3870 vdd.n2865 gnd 0.009044f
C3871 vdd.n2866 gnd 0.651603f
C3872 vdd.n2867 gnd 0.009044f
C3873 vdd.n2868 gnd 0.007279f
C3874 vdd.n2869 gnd 0.009044f
C3875 vdd.n2870 gnd 0.009044f
C3876 vdd.n2871 gnd 0.009044f
C3877 vdd.n2872 gnd 0.007279f
C3878 vdd.n2873 gnd 0.009044f
C3879 vdd.t125 gnd 0.46213f
C3880 vdd.n2874 gnd 0.767136f
C3881 vdd.n2875 gnd 0.009044f
C3882 vdd.n2876 gnd 0.007279f
C3883 vdd.n2877 gnd 0.009044f
C3884 vdd.n2878 gnd 0.009044f
C3885 vdd.n2879 gnd 0.009044f
C3886 vdd.n2880 gnd 0.007279f
C3887 vdd.n2881 gnd 0.009044f
C3888 vdd.n2882 gnd 0.725544f
C3889 vdd.n2883 gnd 0.009044f
C3890 vdd.n2884 gnd 0.007279f
C3891 vdd.n2885 gnd 0.009044f
C3892 vdd.n2886 gnd 0.009044f
C3893 vdd.n2887 gnd 0.009044f
C3894 vdd.n2888 gnd 0.007279f
C3895 vdd.n2889 gnd 0.007279f
C3896 vdd.n2890 gnd 0.007279f
C3897 vdd.n2891 gnd 0.009044f
C3898 vdd.n2892 gnd 0.009044f
C3899 vdd.n2893 gnd 0.009044f
C3900 vdd.n2894 gnd 0.007279f
C3901 vdd.n2895 gnd 0.007279f
C3902 vdd.n2896 gnd 0.007279f
C3903 vdd.n2897 gnd 0.009044f
C3904 vdd.n2898 gnd 0.009044f
C3905 vdd.n2899 gnd 0.009044f
C3906 vdd.n2900 gnd 0.007279f
C3907 vdd.n2901 gnd 0.007279f
C3908 vdd.n2902 gnd 0.006042f
C3909 vdd.n2903 gnd 0.022041f
C3910 vdd.n2904 gnd 0.022546f
C3911 vdd.n2906 gnd 0.022546f
C3912 vdd.n2907 gnd 0.003458f
C3913 vdd.t93 gnd 0.111266f
C3914 vdd.t92 gnd 0.118912f
C3915 vdd.t91 gnd 0.145312f
C3916 vdd.n2908 gnd 0.186269f
C3917 vdd.n2909 gnd 0.157227f
C3918 vdd.n2910 gnd 0.011938f
C3919 vdd.n2911 gnd 0.003822f
C3920 vdd.n2912 gnd 0.007279f
C3921 vdd.n2913 gnd 0.009044f
C3922 vdd.n2915 gnd 0.009044f
C3923 vdd.n2916 gnd 0.009044f
C3924 vdd.n2917 gnd 0.007279f
C3925 vdd.n2918 gnd 0.007279f
C3926 vdd.n2919 gnd 0.007279f
C3927 vdd.n2920 gnd 0.009044f
C3928 vdd.n2922 gnd 0.009044f
C3929 vdd.n2923 gnd 0.009044f
C3930 vdd.n2924 gnd 0.007279f
C3931 vdd.n2925 gnd 0.007279f
C3932 vdd.n2926 gnd 0.007279f
C3933 vdd.n2927 gnd 0.009044f
C3934 vdd.n2929 gnd 0.009044f
C3935 vdd.n2930 gnd 0.009044f
C3936 vdd.n2931 gnd 0.007279f
C3937 vdd.n2932 gnd 0.007279f
C3938 vdd.n2933 gnd 0.007279f
C3939 vdd.n2934 gnd 0.009044f
C3940 vdd.n2936 gnd 0.009044f
C3941 vdd.n2937 gnd 0.009044f
C3942 vdd.n2938 gnd 0.007279f
C3943 vdd.n2939 gnd 0.007279f
C3944 vdd.n2940 gnd 0.007279f
C3945 vdd.n2941 gnd 0.009044f
C3946 vdd.n2943 gnd 0.009044f
C3947 vdd.n2944 gnd 0.009044f
C3948 vdd.n2945 gnd 0.007279f
C3949 vdd.n2946 gnd 0.009044f
C3950 vdd.n2947 gnd 0.009044f
C3951 vdd.n2948 gnd 0.009044f
C3952 vdd.n2949 gnd 0.015578f
C3953 vdd.n2950 gnd 0.00495f
C3954 vdd.n2951 gnd 0.007279f
C3955 vdd.n2952 gnd 0.009044f
C3956 vdd.n2954 gnd 0.009044f
C3957 vdd.n2955 gnd 0.009044f
C3958 vdd.n2956 gnd 0.007279f
C3959 vdd.n2957 gnd 0.007279f
C3960 vdd.n2958 gnd 0.007279f
C3961 vdd.n2959 gnd 0.009044f
C3962 vdd.n2961 gnd 0.009044f
C3963 vdd.n2962 gnd 0.009044f
C3964 vdd.n2963 gnd 0.007279f
C3965 vdd.n2964 gnd 0.007279f
C3966 vdd.n2965 gnd 0.007279f
C3967 vdd.n2966 gnd 0.009044f
C3968 vdd.n2968 gnd 0.009044f
C3969 vdd.n2969 gnd 0.009044f
C3970 vdd.n2970 gnd 0.007279f
C3971 vdd.n2971 gnd 0.007279f
C3972 vdd.n2972 gnd 0.007279f
C3973 vdd.n2973 gnd 0.009044f
C3974 vdd.n2975 gnd 0.009044f
C3975 vdd.n2976 gnd 0.009044f
C3976 vdd.n2977 gnd 0.007279f
C3977 vdd.n2978 gnd 0.007279f
C3978 vdd.n2979 gnd 0.007279f
C3979 vdd.n2980 gnd 0.009044f
C3980 vdd.n2982 gnd 0.009044f
C3981 vdd.n2983 gnd 0.009044f
C3982 vdd.n2984 gnd 0.007279f
C3983 vdd.n2985 gnd 0.009044f
C3984 vdd.n2986 gnd 0.009044f
C3985 vdd.n2987 gnd 0.009044f
C3986 vdd.n2988 gnd 0.015578f
C3987 vdd.n2989 gnd 0.006078f
C3988 vdd.n2990 gnd 0.007279f
C3989 vdd.n2991 gnd 0.009044f
C3990 vdd.n2993 gnd 0.009044f
C3991 vdd.n2994 gnd 0.009044f
C3992 vdd.n2995 gnd 0.007279f
C3993 vdd.n2996 gnd 0.007279f
C3994 vdd.n2997 gnd 0.007279f
C3995 vdd.n2998 gnd 0.009044f
C3996 vdd.n3000 gnd 0.009044f
C3997 vdd.n3001 gnd 0.009044f
C3998 vdd.n3002 gnd 0.007279f
C3999 vdd.n3003 gnd 0.007279f
C4000 vdd.n3004 gnd 0.007279f
C4001 vdd.n3005 gnd 0.009044f
C4002 vdd.n3007 gnd 0.009044f
C4003 vdd.n3008 gnd 0.009044f
C4004 vdd.n3009 gnd 0.007279f
C4005 vdd.n3010 gnd 0.007279f
C4006 vdd.n3011 gnd 0.007279f
C4007 vdd.n3012 gnd 0.009044f
C4008 vdd.n3014 gnd 0.009044f
C4009 vdd.n3015 gnd 0.009044f
C4010 vdd.n3017 gnd 0.009044f
C4011 vdd.n3018 gnd 0.007279f
C4012 vdd.n3019 gnd 0.007279f
C4013 vdd.n3020 gnd 0.006042f
C4014 vdd.n3021 gnd 0.022546f
C4015 vdd.n3022 gnd 0.022041f
C4016 vdd.n3023 gnd 0.006042f
C4017 vdd.n3024 gnd 0.022041f
C4018 vdd.n3025 gnd 1.36328f
C4019 vdd.t44 gnd 0.46213f
C4020 vdd.n3026 gnd 0.485236f
C4021 vdd.n3027 gnd 0.92426f
C4022 vdd.n3028 gnd 0.009044f
C4023 vdd.n3029 gnd 0.007279f
C4024 vdd.n3030 gnd 0.007279f
C4025 vdd.n3031 gnd 0.007279f
C4026 vdd.n3032 gnd 0.009044f
C4027 vdd.n3033 gnd 0.827213f
C4028 vdd.t116 gnd 0.46213f
C4029 vdd.n3034 gnd 0.559177f
C4030 vdd.n3035 gnd 0.670088f
C4031 vdd.n3036 gnd 0.009044f
C4032 vdd.n3037 gnd 0.007279f
C4033 vdd.n3038 gnd 0.007279f
C4034 vdd.n3039 gnd 0.007279f
C4035 vdd.n3040 gnd 0.009044f
C4036 vdd.n3041 gnd 0.512964f
C4037 vdd.t138 gnd 0.46213f
C4038 vdd.n3042 gnd 0.767136f
C4039 vdd.t114 gnd 0.46213f
C4040 vdd.n3043 gnd 0.56842f
C4041 vdd.n3044 gnd 0.009044f
C4042 vdd.n3045 gnd 0.007279f
C4043 vdd.n3046 gnd 0.006951f
C4044 vdd.n3047 gnd 0.533453f
C4045 vdd.n3048 gnd 1.83173f
C4046 a_n5644_8799.n0 gnd 0.207505f
C4047 a_n5644_8799.n1 gnd 0.286067f
C4048 a_n5644_8799.n2 gnd 0.217042f
C4049 a_n5644_8799.n3 gnd 0.207505f
C4050 a_n5644_8799.n4 gnd 0.286067f
C4051 a_n5644_8799.n5 gnd 0.217042f
C4052 a_n5644_8799.n6 gnd 0.207505f
C4053 a_n5644_8799.n7 gnd 0.450817f
C4054 a_n5644_8799.n8 gnd 0.217042f
C4055 a_n5644_8799.n9 gnd 0.207505f
C4056 a_n5644_8799.n10 gnd 0.320795f
C4057 a_n5644_8799.n11 gnd 0.182314f
C4058 a_n5644_8799.n12 gnd 0.207505f
C4059 a_n5644_8799.n13 gnd 0.320795f
C4060 a_n5644_8799.n14 gnd 0.182314f
C4061 a_n5644_8799.n15 gnd 0.207505f
C4062 a_n5644_8799.n16 gnd 0.320795f
C4063 a_n5644_8799.n17 gnd 0.347064f
C4064 a_n5644_8799.n18 gnd 2.78717f
C4065 a_n5644_8799.n19 gnd 4.02361f
C4066 a_n5644_8799.n20 gnd 0.362739f
C4067 a_n5644_8799.n21 gnd 3.04009f
C4068 a_n5644_8799.n22 gnd 0.362738f
C4069 a_n5644_8799.n23 gnd 0.854945f
C4070 a_n5644_8799.n24 gnd 0.249816f
C4071 a_n5644_8799.n25 gnd 0.004664f
C4072 a_n5644_8799.n26 gnd 0.010087f
C4073 a_n5644_8799.n27 gnd 0.010087f
C4074 a_n5644_8799.n28 gnd 0.004664f
C4075 a_n5644_8799.n29 gnd 0.249816f
C4076 a_n5644_8799.n30 gnd 0.004664f
C4077 a_n5644_8799.n31 gnd 0.010087f
C4078 a_n5644_8799.n32 gnd 0.010087f
C4079 a_n5644_8799.n33 gnd 0.004664f
C4080 a_n5644_8799.n34 gnd 0.249816f
C4081 a_n5644_8799.n35 gnd 0.004664f
C4082 a_n5644_8799.n36 gnd 0.010087f
C4083 a_n5644_8799.n37 gnd 0.010087f
C4084 a_n5644_8799.n38 gnd 0.004664f
C4085 a_n5644_8799.n39 gnd 0.004664f
C4086 a_n5644_8799.n40 gnd 0.010087f
C4087 a_n5644_8799.n41 gnd 0.010087f
C4088 a_n5644_8799.n42 gnd 0.004664f
C4089 a_n5644_8799.n43 gnd 0.249816f
C4090 a_n5644_8799.n44 gnd 0.004664f
C4091 a_n5644_8799.n45 gnd 0.010087f
C4092 a_n5644_8799.n46 gnd 0.010087f
C4093 a_n5644_8799.n47 gnd 0.004664f
C4094 a_n5644_8799.n48 gnd 0.249816f
C4095 a_n5644_8799.n49 gnd 0.004664f
C4096 a_n5644_8799.n50 gnd 0.010087f
C4097 a_n5644_8799.n51 gnd 0.010087f
C4098 a_n5644_8799.n52 gnd 0.004664f
C4099 a_n5644_8799.n53 gnd 0.249816f
C4100 a_n5644_8799.t15 gnd 0.143928f
C4101 a_n5644_8799.t21 gnd 0.143928f
C4102 a_n5644_8799.t30 gnd 0.143928f
C4103 a_n5644_8799.n54 gnd 1.13518f
C4104 a_n5644_8799.t8 gnd 0.143928f
C4105 a_n5644_8799.t10 gnd 0.143928f
C4106 a_n5644_8799.n55 gnd 1.13331f
C4107 a_n5644_8799.t7 gnd 0.143928f
C4108 a_n5644_8799.t6 gnd 0.143928f
C4109 a_n5644_8799.n56 gnd 1.13331f
C4110 a_n5644_8799.t18 gnd 0.111944f
C4111 a_n5644_8799.t24 gnd 0.111944f
C4112 a_n5644_8799.n57 gnd 0.992092f
C4113 a_n5644_8799.t35 gnd 0.111944f
C4114 a_n5644_8799.t23 gnd 0.111944f
C4115 a_n5644_8799.n58 gnd 0.989175f
C4116 a_n5644_8799.n59 gnd 0.877149f
C4117 a_n5644_8799.t20 gnd 0.111944f
C4118 a_n5644_8799.t19 gnd 0.111944f
C4119 a_n5644_8799.n60 gnd 0.989175f
C4120 a_n5644_8799.t25 gnd 0.111944f
C4121 a_n5644_8799.t31 gnd 0.111944f
C4122 a_n5644_8799.n61 gnd 0.992091f
C4123 a_n5644_8799.t2 gnd 0.111944f
C4124 a_n5644_8799.t29 gnd 0.111944f
C4125 a_n5644_8799.n62 gnd 0.989174f
C4126 a_n5644_8799.n63 gnd 0.877151f
C4127 a_n5644_8799.t13 gnd 0.111944f
C4128 a_n5644_8799.t22 gnd 0.111944f
C4129 a_n5644_8799.n64 gnd 0.989174f
C4130 a_n5644_8799.t14 gnd 0.111944f
C4131 a_n5644_8799.t3 gnd 0.111944f
C4132 a_n5644_8799.n65 gnd 0.992091f
C4133 a_n5644_8799.t4 gnd 0.111944f
C4134 a_n5644_8799.t34 gnd 0.111944f
C4135 a_n5644_8799.n66 gnd 0.989174f
C4136 a_n5644_8799.n67 gnd 0.877151f
C4137 a_n5644_8799.t11 gnd 0.111944f
C4138 a_n5644_8799.t17 gnd 0.111944f
C4139 a_n5644_8799.n68 gnd 0.989174f
C4140 a_n5644_8799.t33 gnd 0.111944f
C4141 a_n5644_8799.t32 gnd 0.111944f
C4142 a_n5644_8799.n69 gnd 0.989175f
C4143 a_n5644_8799.n70 gnd 3.08572f
C4144 a_n5644_8799.t0 gnd 0.111944f
C4145 a_n5644_8799.t12 gnd 0.111944f
C4146 a_n5644_8799.n71 gnd 0.989175f
C4147 a_n5644_8799.n72 gnd 0.431882f
C4148 a_n5644_8799.t1 gnd 0.111944f
C4149 a_n5644_8799.t9 gnd 0.111944f
C4150 a_n5644_8799.n73 gnd 0.989175f
C4151 a_n5644_8799.t75 gnd 0.596792f
C4152 a_n5644_8799.n74 gnd 0.268224f
C4153 a_n5644_8799.t42 gnd 0.596792f
C4154 a_n5644_8799.t62 gnd 0.596792f
C4155 a_n5644_8799.t53 gnd 0.608087f
C4156 a_n5644_8799.n75 gnd 0.250184f
C4157 a_n5644_8799.n76 gnd 0.270608f
C4158 a_n5644_8799.t77 gnd 0.596792f
C4159 a_n5644_8799.n77 gnd 0.268224f
C4160 a_n5644_8799.n78 gnd 0.26382f
C4161 a_n5644_8799.t52 gnd 0.596792f
C4162 a_n5644_8799.n79 gnd 0.26382f
C4163 a_n5644_8799.t41 gnd 0.596792f
C4164 a_n5644_8799.n80 gnd 0.270608f
C4165 a_n5644_8799.t40 gnd 0.608077f
C4166 a_n5644_8799.t79 gnd 0.596792f
C4167 a_n5644_8799.n81 gnd 0.268224f
C4168 a_n5644_8799.t49 gnd 0.596792f
C4169 a_n5644_8799.t68 gnd 0.596792f
C4170 a_n5644_8799.t58 gnd 0.608087f
C4171 a_n5644_8799.n82 gnd 0.250184f
C4172 a_n5644_8799.n83 gnd 0.270608f
C4173 a_n5644_8799.t81 gnd 0.596792f
C4174 a_n5644_8799.n84 gnd 0.268224f
C4175 a_n5644_8799.n85 gnd 0.26382f
C4176 a_n5644_8799.t57 gnd 0.596792f
C4177 a_n5644_8799.n86 gnd 0.26382f
C4178 a_n5644_8799.t45 gnd 0.596792f
C4179 a_n5644_8799.n87 gnd 0.270608f
C4180 a_n5644_8799.t47 gnd 0.608077f
C4181 a_n5644_8799.n88 gnd 0.897554f
C4182 a_n5644_8799.t66 gnd 0.596792f
C4183 a_n5644_8799.n89 gnd 0.268224f
C4184 a_n5644_8799.t74 gnd 0.596792f
C4185 a_n5644_8799.t71 gnd 0.596792f
C4186 a_n5644_8799.t39 gnd 0.608087f
C4187 a_n5644_8799.n90 gnd 0.250184f
C4188 a_n5644_8799.n91 gnd 0.270608f
C4189 a_n5644_8799.t48 gnd 0.596792f
C4190 a_n5644_8799.n92 gnd 0.268224f
C4191 a_n5644_8799.n93 gnd 0.26382f
C4192 a_n5644_8799.t54 gnd 0.596792f
C4193 a_n5644_8799.n94 gnd 0.26382f
C4194 a_n5644_8799.t43 gnd 0.596792f
C4195 a_n5644_8799.n95 gnd 0.270608f
C4196 a_n5644_8799.t83 gnd 0.608077f
C4197 a_n5644_8799.n96 gnd 1.53678f
C4198 a_n5644_8799.t60 gnd 0.608077f
C4199 a_n5644_8799.t59 gnd 0.596792f
C4200 a_n5644_8799.t46 gnd 0.596792f
C4201 a_n5644_8799.n97 gnd 0.268224f
C4202 a_n5644_8799.t76 gnd 0.596792f
C4203 a_n5644_8799.t61 gnd 0.596792f
C4204 a_n5644_8799.t51 gnd 0.596792f
C4205 a_n5644_8799.n98 gnd 0.268224f
C4206 a_n5644_8799.t69 gnd 0.608087f
C4207 a_n5644_8799.n99 gnd 0.250184f
C4208 a_n5644_8799.t78 gnd 0.596792f
C4209 a_n5644_8799.n100 gnd 0.270608f
C4210 a_n5644_8799.n101 gnd 0.26382f
C4211 a_n5644_8799.n102 gnd 0.26382f
C4212 a_n5644_8799.n103 gnd 0.270608f
C4213 a_n5644_8799.t64 gnd 0.608077f
C4214 a_n5644_8799.t63 gnd 0.596792f
C4215 a_n5644_8799.t55 gnd 0.596792f
C4216 a_n5644_8799.n104 gnd 0.268224f
C4217 a_n5644_8799.t80 gnd 0.596792f
C4218 a_n5644_8799.t67 gnd 0.596792f
C4219 a_n5644_8799.t56 gnd 0.596792f
C4220 a_n5644_8799.n105 gnd 0.268224f
C4221 a_n5644_8799.t72 gnd 0.608087f
C4222 a_n5644_8799.n106 gnd 0.250184f
C4223 a_n5644_8799.t36 gnd 0.596792f
C4224 a_n5644_8799.n107 gnd 0.270608f
C4225 a_n5644_8799.n108 gnd 0.26382f
C4226 a_n5644_8799.n109 gnd 0.26382f
C4227 a_n5644_8799.n110 gnd 0.270608f
C4228 a_n5644_8799.n111 gnd 0.897554f
C4229 a_n5644_8799.t82 gnd 0.608077f
C4230 a_n5644_8799.t44 gnd 0.596792f
C4231 a_n5644_8799.t65 gnd 0.596792f
C4232 a_n5644_8799.n112 gnd 0.268224f
C4233 a_n5644_8799.t37 gnd 0.596792f
C4234 a_n5644_8799.t73 gnd 0.596792f
C4235 a_n5644_8799.t50 gnd 0.596792f
C4236 a_n5644_8799.n113 gnd 0.268224f
C4237 a_n5644_8799.t38 gnd 0.608087f
C4238 a_n5644_8799.n114 gnd 0.250184f
C4239 a_n5644_8799.t70 gnd 0.596792f
C4240 a_n5644_8799.n115 gnd 0.270608f
C4241 a_n5644_8799.n116 gnd 0.26382f
C4242 a_n5644_8799.n117 gnd 0.26382f
C4243 a_n5644_8799.n118 gnd 0.270608f
C4244 a_n5644_8799.n119 gnd 1.0844f
C4245 a_n5644_8799.n120 gnd 12.1892f
C4246 a_n5644_8799.n121 gnd 4.36765f
C4247 a_n5644_8799.n122 gnd 5.66677f
C4248 a_n5644_8799.t26 gnd 0.143928f
C4249 a_n5644_8799.t27 gnd 0.143928f
C4250 a_n5644_8799.n123 gnd 1.13331f
C4251 a_n5644_8799.t28 gnd 0.143928f
C4252 a_n5644_8799.t16 gnd 0.143928f
C4253 a_n5644_8799.n124 gnd 1.13518f
C4254 a_n5644_8799.n125 gnd 1.13331f
C4255 a_n5644_8799.t5 gnd 0.143928f
C4256 CSoutput.n0 gnd 0.036216f
C4257 CSoutput.t106 gnd 0.239559f
C4258 CSoutput.n1 gnd 0.108173f
C4259 CSoutput.n2 gnd 0.036216f
C4260 CSoutput.t111 gnd 0.239559f
C4261 CSoutput.n3 gnd 0.028704f
C4262 CSoutput.n4 gnd 0.036216f
C4263 CSoutput.t100 gnd 0.239559f
C4264 CSoutput.n5 gnd 0.024752f
C4265 CSoutput.n6 gnd 0.036216f
C4266 CSoutput.t108 gnd 0.239559f
C4267 CSoutput.t114 gnd 0.239559f
C4268 CSoutput.n7 gnd 0.106994f
C4269 CSoutput.n8 gnd 0.036216f
C4270 CSoutput.t113 gnd 0.239559f
C4271 CSoutput.n9 gnd 0.023599f
C4272 CSoutput.n10 gnd 0.036216f
C4273 CSoutput.t101 gnd 0.239559f
C4274 CSoutput.t112 gnd 0.239559f
C4275 CSoutput.n11 gnd 0.106994f
C4276 CSoutput.n12 gnd 0.036216f
C4277 CSoutput.t110 gnd 0.239559f
C4278 CSoutput.n13 gnd 0.024752f
C4279 CSoutput.n14 gnd 0.036216f
C4280 CSoutput.t99 gnd 0.239559f
C4281 CSoutput.t103 gnd 0.239559f
C4282 CSoutput.n15 gnd 0.106994f
C4283 CSoutput.n16 gnd 0.036216f
C4284 CSoutput.t107 gnd 0.239559f
C4285 CSoutput.n17 gnd 0.026436f
C4286 CSoutput.t117 gnd 0.286279f
C4287 CSoutput.t97 gnd 0.239559f
C4288 CSoutput.n18 gnd 0.13659f
C4289 CSoutput.n19 gnd 0.132539f
C4290 CSoutput.n20 gnd 0.153761f
C4291 CSoutput.n21 gnd 0.036216f
C4292 CSoutput.n22 gnd 0.030226f
C4293 CSoutput.n23 gnd 0.106994f
C4294 CSoutput.n24 gnd 0.029137f
C4295 CSoutput.n25 gnd 0.028704f
C4296 CSoutput.n26 gnd 0.036216f
C4297 CSoutput.n27 gnd 0.036216f
C4298 CSoutput.n28 gnd 0.029994f
C4299 CSoutput.n29 gnd 0.025465f
C4300 CSoutput.n30 gnd 0.109376f
C4301 CSoutput.n31 gnd 0.025816f
C4302 CSoutput.n32 gnd 0.036216f
C4303 CSoutput.n33 gnd 0.036216f
C4304 CSoutput.n34 gnd 0.036216f
C4305 CSoutput.n35 gnd 0.029674f
C4306 CSoutput.n36 gnd 0.106994f
C4307 CSoutput.n37 gnd 0.028379f
C4308 CSoutput.n38 gnd 0.029462f
C4309 CSoutput.n39 gnd 0.036216f
C4310 CSoutput.n40 gnd 0.036216f
C4311 CSoutput.n41 gnd 0.03022f
C4312 CSoutput.n42 gnd 0.027621f
C4313 CSoutput.n43 gnd 0.106994f
C4314 CSoutput.n44 gnd 0.028321f
C4315 CSoutput.n45 gnd 0.036216f
C4316 CSoutput.n46 gnd 0.036216f
C4317 CSoutput.n47 gnd 0.036216f
C4318 CSoutput.n48 gnd 0.028321f
C4319 CSoutput.n49 gnd 0.106994f
C4320 CSoutput.n50 gnd 0.027621f
C4321 CSoutput.n51 gnd 0.03022f
C4322 CSoutput.n52 gnd 0.036216f
C4323 CSoutput.n53 gnd 0.036216f
C4324 CSoutput.n54 gnd 0.029462f
C4325 CSoutput.n55 gnd 0.028379f
C4326 CSoutput.n56 gnd 0.106994f
C4327 CSoutput.n57 gnd 0.029674f
C4328 CSoutput.n58 gnd 0.036216f
C4329 CSoutput.n59 gnd 0.036216f
C4330 CSoutput.n60 gnd 0.036216f
C4331 CSoutput.n61 gnd 0.025816f
C4332 CSoutput.n62 gnd 0.109376f
C4333 CSoutput.n63 gnd 0.025465f
C4334 CSoutput.t116 gnd 0.239559f
C4335 CSoutput.n64 gnd 0.106994f
C4336 CSoutput.n65 gnd 0.029994f
C4337 CSoutput.n66 gnd 0.036216f
C4338 CSoutput.n67 gnd 0.036216f
C4339 CSoutput.n68 gnd 0.036216f
C4340 CSoutput.n69 gnd 0.029137f
C4341 CSoutput.n70 gnd 0.106994f
C4342 CSoutput.n71 gnd 0.030226f
C4343 CSoutput.n72 gnd 0.026436f
C4344 CSoutput.n73 gnd 0.036216f
C4345 CSoutput.n74 gnd 0.036216f
C4346 CSoutput.n75 gnd 0.027416f
C4347 CSoutput.n76 gnd 0.016282f
C4348 CSoutput.t96 gnd 0.269161f
C4349 CSoutput.n77 gnd 0.133709f
C4350 CSoutput.n78 gnd 0.572127f
C4351 CSoutput.t84 gnd 0.045174f
C4352 CSoutput.t93 gnd 0.045174f
C4353 CSoutput.n79 gnd 0.349752f
C4354 CSoutput.t77 gnd 0.045174f
C4355 CSoutput.t82 gnd 0.045174f
C4356 CSoutput.n80 gnd 0.349128f
C4357 CSoutput.n81 gnd 0.354365f
C4358 CSoutput.t72 gnd 0.045174f
C4359 CSoutput.t85 gnd 0.045174f
C4360 CSoutput.n82 gnd 0.349128f
C4361 CSoutput.n83 gnd 0.174616f
C4362 CSoutput.t10 gnd 0.045174f
C4363 CSoutput.t80 gnd 0.045174f
C4364 CSoutput.n84 gnd 0.349128f
C4365 CSoutput.n85 gnd 0.320205f
C4366 CSoutput.t76 gnd 0.045174f
C4367 CSoutput.t9 gnd 0.045174f
C4368 CSoutput.n86 gnd 0.349752f
C4369 CSoutput.t73 gnd 0.045174f
C4370 CSoutput.t88 gnd 0.045174f
C4371 CSoutput.n87 gnd 0.349128f
C4372 CSoutput.n88 gnd 0.354365f
C4373 CSoutput.t83 gnd 0.045174f
C4374 CSoutput.t79 gnd 0.045174f
C4375 CSoutput.n89 gnd 0.349128f
C4376 CSoutput.n90 gnd 0.174616f
C4377 CSoutput.t5 gnd 0.045174f
C4378 CSoutput.t69 gnd 0.045174f
C4379 CSoutput.n91 gnd 0.349128f
C4380 CSoutput.n92 gnd 0.260396f
C4381 CSoutput.n93 gnd 0.328358f
C4382 CSoutput.t0 gnd 0.045174f
C4383 CSoutput.t14 gnd 0.045174f
C4384 CSoutput.n94 gnd 0.349752f
C4385 CSoutput.t11 gnd 0.045174f
C4386 CSoutput.t17 gnd 0.045174f
C4387 CSoutput.n95 gnd 0.349128f
C4388 CSoutput.n96 gnd 0.354365f
C4389 CSoutput.t2 gnd 0.045174f
C4390 CSoutput.t94 gnd 0.045174f
C4391 CSoutput.n97 gnd 0.349128f
C4392 CSoutput.n98 gnd 0.174616f
C4393 CSoutput.t87 gnd 0.045174f
C4394 CSoutput.t92 gnd 0.045174f
C4395 CSoutput.n99 gnd 0.349128f
C4396 CSoutput.n100 gnd 0.260396f
C4397 CSoutput.n101 gnd 0.36702f
C4398 CSoutput.n102 gnd 6.17074f
C4399 CSoutput.n104 gnd 0.640649f
C4400 CSoutput.n105 gnd 0.480487f
C4401 CSoutput.n106 gnd 0.640649f
C4402 CSoutput.n107 gnd 0.640649f
C4403 CSoutput.n108 gnd 1.72482f
C4404 CSoutput.n109 gnd 0.640649f
C4405 CSoutput.n110 gnd 0.640649f
C4406 CSoutput.t115 gnd 0.800811f
C4407 CSoutput.n111 gnd 0.640649f
C4408 CSoutput.n112 gnd 0.640649f
C4409 CSoutput.n116 gnd 0.640649f
C4410 CSoutput.n120 gnd 0.640649f
C4411 CSoutput.n121 gnd 0.640649f
C4412 CSoutput.n123 gnd 0.640649f
C4413 CSoutput.n128 gnd 0.640649f
C4414 CSoutput.n130 gnd 0.640649f
C4415 CSoutput.n131 gnd 0.640649f
C4416 CSoutput.n133 gnd 0.640649f
C4417 CSoutput.n134 gnd 0.640649f
C4418 CSoutput.n136 gnd 0.640649f
C4419 CSoutput.t104 gnd 10.7052f
C4420 CSoutput.n138 gnd 0.640649f
C4421 CSoutput.n139 gnd 0.480487f
C4422 CSoutput.n140 gnd 0.640649f
C4423 CSoutput.n141 gnd 0.640649f
C4424 CSoutput.n142 gnd 1.72482f
C4425 CSoutput.n143 gnd 0.640649f
C4426 CSoutput.n144 gnd 0.640649f
C4427 CSoutput.t102 gnd 0.800811f
C4428 CSoutput.n145 gnd 0.640649f
C4429 CSoutput.n146 gnd 0.640649f
C4430 CSoutput.n150 gnd 0.640649f
C4431 CSoutput.n154 gnd 0.640649f
C4432 CSoutput.n155 gnd 0.640649f
C4433 CSoutput.n157 gnd 0.640649f
C4434 CSoutput.n162 gnd 0.640649f
C4435 CSoutput.n164 gnd 0.640649f
C4436 CSoutput.n165 gnd 0.640649f
C4437 CSoutput.n167 gnd 0.640649f
C4438 CSoutput.n168 gnd 0.640649f
C4439 CSoutput.n170 gnd 0.640649f
C4440 CSoutput.n171 gnd 0.480487f
C4441 CSoutput.n173 gnd 0.640649f
C4442 CSoutput.n174 gnd 0.480487f
C4443 CSoutput.n175 gnd 0.640649f
C4444 CSoutput.n176 gnd 0.640649f
C4445 CSoutput.n177 gnd 1.72482f
C4446 CSoutput.n178 gnd 0.640649f
C4447 CSoutput.n179 gnd 0.640649f
C4448 CSoutput.t98 gnd 0.800811f
C4449 CSoutput.n180 gnd 0.640649f
C4450 CSoutput.n181 gnd 1.72482f
C4451 CSoutput.n183 gnd 0.640649f
C4452 CSoutput.n184 gnd 0.640649f
C4453 CSoutput.n186 gnd 0.640649f
C4454 CSoutput.n187 gnd 0.640649f
C4455 CSoutput.t105 gnd 10.5307f
C4456 CSoutput.t109 gnd 10.7052f
C4457 CSoutput.n193 gnd 2.00981f
C4458 CSoutput.n194 gnd 8.18723f
C4459 CSoutput.n195 gnd 8.52982f
C4460 CSoutput.n200 gnd 2.17717f
C4461 CSoutput.n206 gnd 0.640649f
C4462 CSoutput.n208 gnd 0.640649f
C4463 CSoutput.n210 gnd 0.640649f
C4464 CSoutput.n212 gnd 0.640649f
C4465 CSoutput.n214 gnd 0.640649f
C4466 CSoutput.n220 gnd 0.640649f
C4467 CSoutput.n227 gnd 1.17534f
C4468 CSoutput.n228 gnd 1.17534f
C4469 CSoutput.n229 gnd 0.640649f
C4470 CSoutput.n230 gnd 0.640649f
C4471 CSoutput.n232 gnd 0.480487f
C4472 CSoutput.n233 gnd 0.411494f
C4473 CSoutput.n235 gnd 0.480487f
C4474 CSoutput.n236 gnd 0.411494f
C4475 CSoutput.n237 gnd 0.480487f
C4476 CSoutput.n239 gnd 0.640649f
C4477 CSoutput.n241 gnd 1.72482f
C4478 CSoutput.n242 gnd 2.00981f
C4479 CSoutput.n243 gnd 7.53015f
C4480 CSoutput.n245 gnd 0.480487f
C4481 CSoutput.n246 gnd 1.23632f
C4482 CSoutput.n247 gnd 0.480487f
C4483 CSoutput.n249 gnd 0.640649f
C4484 CSoutput.n251 gnd 1.72482f
C4485 CSoutput.n252 gnd 3.75694f
C4486 CSoutput.t89 gnd 0.045174f
C4487 CSoutput.t6 gnd 0.045174f
C4488 CSoutput.n253 gnd 0.349752f
C4489 CSoutput.t12 gnd 0.045174f
C4490 CSoutput.t90 gnd 0.045174f
C4491 CSoutput.n254 gnd 0.349128f
C4492 CSoutput.n255 gnd 0.354365f
C4493 CSoutput.t8 gnd 0.045174f
C4494 CSoutput.t74 gnd 0.045174f
C4495 CSoutput.n256 gnd 0.349128f
C4496 CSoutput.n257 gnd 0.174616f
C4497 CSoutput.t71 gnd 0.045174f
C4498 CSoutput.t68 gnd 0.045174f
C4499 CSoutput.n258 gnd 0.349128f
C4500 CSoutput.n259 gnd 0.320205f
C4501 CSoutput.t18 gnd 0.045174f
C4502 CSoutput.t91 gnd 0.045174f
C4503 CSoutput.n260 gnd 0.349752f
C4504 CSoutput.t86 gnd 0.045174f
C4505 CSoutput.t19 gnd 0.045174f
C4506 CSoutput.n261 gnd 0.349128f
C4507 CSoutput.n262 gnd 0.354365f
C4508 CSoutput.t70 gnd 0.045174f
C4509 CSoutput.t95 gnd 0.045174f
C4510 CSoutput.n263 gnd 0.349128f
C4511 CSoutput.n264 gnd 0.174616f
C4512 CSoutput.t1 gnd 0.045174f
C4513 CSoutput.t4 gnd 0.045174f
C4514 CSoutput.n265 gnd 0.349128f
C4515 CSoutput.n266 gnd 0.260396f
C4516 CSoutput.n267 gnd 0.328358f
C4517 CSoutput.t13 gnd 0.045174f
C4518 CSoutput.t15 gnd 0.045174f
C4519 CSoutput.n268 gnd 0.349752f
C4520 CSoutput.t75 gnd 0.045174f
C4521 CSoutput.t16 gnd 0.045174f
C4522 CSoutput.n269 gnd 0.349128f
C4523 CSoutput.n270 gnd 0.354365f
C4524 CSoutput.t81 gnd 0.045174f
C4525 CSoutput.t3 gnd 0.045174f
C4526 CSoutput.n271 gnd 0.349128f
C4527 CSoutput.n272 gnd 0.174616f
C4528 CSoutput.t78 gnd 0.045174f
C4529 CSoutput.t7 gnd 0.045174f
C4530 CSoutput.n273 gnd 0.349127f
C4531 CSoutput.n274 gnd 0.260397f
C4532 CSoutput.n275 gnd 0.36702f
C4533 CSoutput.n276 gnd 9.063099f
C4534 CSoutput.t44 gnd 0.039527f
C4535 CSoutput.t34 gnd 0.039527f
C4536 CSoutput.n277 gnd 0.350445f
C4537 CSoutput.t60 gnd 0.039527f
C4538 CSoutput.t62 gnd 0.039527f
C4539 CSoutput.n278 gnd 0.349276f
C4540 CSoutput.n279 gnd 0.32546f
C4541 CSoutput.t39 gnd 0.039527f
C4542 CSoutput.t29 gnd 0.039527f
C4543 CSoutput.n280 gnd 0.349276f
C4544 CSoutput.n281 gnd 0.160437f
C4545 CSoutput.t65 gnd 0.039527f
C4546 CSoutput.t46 gnd 0.039527f
C4547 CSoutput.n282 gnd 0.349276f
C4548 CSoutput.n283 gnd 0.160437f
C4549 CSoutput.t48 gnd 0.039527f
C4550 CSoutput.t37 gnd 0.039527f
C4551 CSoutput.n284 gnd 0.349276f
C4552 CSoutput.n285 gnd 0.160437f
C4553 CSoutput.t51 gnd 0.039527f
C4554 CSoutput.t53 gnd 0.039527f
C4555 CSoutput.n286 gnd 0.349276f
C4556 CSoutput.n287 gnd 0.295878f
C4557 CSoutput.t54 gnd 0.039527f
C4558 CSoutput.t43 gnd 0.039527f
C4559 CSoutput.n288 gnd 0.350445f
C4560 CSoutput.t66 gnd 0.039527f
C4561 CSoutput.t20 gnd 0.039527f
C4562 CSoutput.n289 gnd 0.349276f
C4563 CSoutput.n290 gnd 0.32546f
C4564 CSoutput.t49 gnd 0.039527f
C4565 CSoutput.t38 gnd 0.039527f
C4566 CSoutput.n291 gnd 0.349276f
C4567 CSoutput.n292 gnd 0.160437f
C4568 CSoutput.t24 gnd 0.039527f
C4569 CSoutput.t55 gnd 0.039527f
C4570 CSoutput.n293 gnd 0.349276f
C4571 CSoutput.n294 gnd 0.160437f
C4572 CSoutput.t57 gnd 0.039527f
C4573 CSoutput.t47 gnd 0.039527f
C4574 CSoutput.n295 gnd 0.349276f
C4575 CSoutput.n296 gnd 0.160437f
C4576 CSoutput.t58 gnd 0.039527f
C4577 CSoutput.t61 gnd 0.039527f
C4578 CSoutput.n297 gnd 0.349276f
C4579 CSoutput.n298 gnd 0.243577f
C4580 CSoutput.n299 gnd 0.452585f
C4581 CSoutput.n300 gnd 9.567129f
C4582 CSoutput.t23 gnd 0.039527f
C4583 CSoutput.t31 gnd 0.039527f
C4584 CSoutput.n301 gnd 0.350445f
C4585 CSoutput.t52 gnd 0.039527f
C4586 CSoutput.t64 gnd 0.039527f
C4587 CSoutput.n302 gnd 0.349276f
C4588 CSoutput.n303 gnd 0.32546f
C4589 CSoutput.t67 gnd 0.039527f
C4590 CSoutput.t27 gnd 0.039527f
C4591 CSoutput.n304 gnd 0.349276f
C4592 CSoutput.n305 gnd 0.160437f
C4593 CSoutput.t32 gnd 0.039527f
C4594 CSoutput.t21 gnd 0.039527f
C4595 CSoutput.n306 gnd 0.349276f
C4596 CSoutput.n307 gnd 0.160437f
C4597 CSoutput.t25 gnd 0.039527f
C4598 CSoutput.t35 gnd 0.039527f
C4599 CSoutput.n308 gnd 0.349276f
C4600 CSoutput.n309 gnd 0.160437f
C4601 CSoutput.t40 gnd 0.039527f
C4602 CSoutput.t56 gnd 0.039527f
C4603 CSoutput.n310 gnd 0.349276f
C4604 CSoutput.n311 gnd 0.295878f
C4605 CSoutput.t30 gnd 0.039527f
C4606 CSoutput.t42 gnd 0.039527f
C4607 CSoutput.n312 gnd 0.350445f
C4608 CSoutput.t59 gnd 0.039527f
C4609 CSoutput.t22 gnd 0.039527f
C4610 CSoutput.n313 gnd 0.349276f
C4611 CSoutput.n314 gnd 0.32546f
C4612 CSoutput.t26 gnd 0.039527f
C4613 CSoutput.t36 gnd 0.039527f
C4614 CSoutput.n315 gnd 0.349276f
C4615 CSoutput.n316 gnd 0.160437f
C4616 CSoutput.t41 gnd 0.039527f
C4617 CSoutput.t28 gnd 0.039527f
C4618 CSoutput.n317 gnd 0.349276f
C4619 CSoutput.n318 gnd 0.160437f
C4620 CSoutput.t33 gnd 0.039527f
C4621 CSoutput.t45 gnd 0.039527f
C4622 CSoutput.n319 gnd 0.349276f
C4623 CSoutput.n320 gnd 0.160437f
C4624 CSoutput.t50 gnd 0.039527f
C4625 CSoutput.t63 gnd 0.039527f
C4626 CSoutput.n321 gnd 0.349276f
C4627 CSoutput.n322 gnd 0.243577f
C4628 CSoutput.n323 gnd 0.452585f
C4629 CSoutput.n324 gnd 5.271f
C4630 CSoutput.n325 gnd 11.7115f
C4631 commonsourceibias.n0 gnd 0.010301f
C4632 commonsourceibias.t71 gnd 0.155981f
C4633 commonsourceibias.t81 gnd 0.144227f
C4634 commonsourceibias.n1 gnd 0.057546f
C4635 commonsourceibias.n2 gnd 0.00772f
C4636 commonsourceibias.t55 gnd 0.144227f
C4637 commonsourceibias.n3 gnd 0.006245f
C4638 commonsourceibias.n4 gnd 0.00772f
C4639 commonsourceibias.t53 gnd 0.144227f
C4640 commonsourceibias.n5 gnd 0.007453f
C4641 commonsourceibias.n6 gnd 0.00772f
C4642 commonsourceibias.t76 gnd 0.144227f
C4643 commonsourceibias.n7 gnd 0.057546f
C4644 commonsourceibias.t86 gnd 0.144227f
C4645 commonsourceibias.n8 gnd 0.006235f
C4646 commonsourceibias.n9 gnd 0.010301f
C4647 commonsourceibias.t32 gnd 0.155981f
C4648 commonsourceibias.t14 gnd 0.144227f
C4649 commonsourceibias.n10 gnd 0.057546f
C4650 commonsourceibias.n11 gnd 0.00772f
C4651 commonsourceibias.t24 gnd 0.144227f
C4652 commonsourceibias.n12 gnd 0.006245f
C4653 commonsourceibias.n13 gnd 0.00772f
C4654 commonsourceibias.t30 gnd 0.144227f
C4655 commonsourceibias.n14 gnd 0.007453f
C4656 commonsourceibias.n15 gnd 0.00772f
C4657 commonsourceibias.t20 gnd 0.144227f
C4658 commonsourceibias.n16 gnd 0.057546f
C4659 commonsourceibias.t36 gnd 0.144227f
C4660 commonsourceibias.n17 gnd 0.006235f
C4661 commonsourceibias.n18 gnd 0.00772f
C4662 commonsourceibias.t44 gnd 0.144227f
C4663 commonsourceibias.t26 gnd 0.144227f
C4664 commonsourceibias.n19 gnd 0.057546f
C4665 commonsourceibias.n20 gnd 0.00772f
C4666 commonsourceibias.t34 gnd 0.144227f
C4667 commonsourceibias.n21 gnd 0.057546f
C4668 commonsourceibias.n22 gnd 0.00772f
C4669 commonsourceibias.t10 gnd 0.144227f
C4670 commonsourceibias.n23 gnd 0.057546f
C4671 commonsourceibias.n24 gnd 0.038863f
C4672 commonsourceibias.t40 gnd 0.144227f
C4673 commonsourceibias.t46 gnd 0.162743f
C4674 commonsourceibias.n25 gnd 0.066782f
C4675 commonsourceibias.n26 gnd 0.069137f
C4676 commonsourceibias.n27 gnd 0.009515f
C4677 commonsourceibias.n28 gnd 0.010526f
C4678 commonsourceibias.n29 gnd 0.00772f
C4679 commonsourceibias.n30 gnd 0.00772f
C4680 commonsourceibias.n31 gnd 0.010457f
C4681 commonsourceibias.n32 gnd 0.006245f
C4682 commonsourceibias.n33 gnd 0.010587f
C4683 commonsourceibias.n34 gnd 0.00772f
C4684 commonsourceibias.n35 gnd 0.00772f
C4685 commonsourceibias.n36 gnd 0.010651f
C4686 commonsourceibias.n37 gnd 0.009185f
C4687 commonsourceibias.n38 gnd 0.007453f
C4688 commonsourceibias.n39 gnd 0.00772f
C4689 commonsourceibias.n40 gnd 0.00772f
C4690 commonsourceibias.n41 gnd 0.009442f
C4691 commonsourceibias.n42 gnd 0.010598f
C4692 commonsourceibias.n43 gnd 0.057546f
C4693 commonsourceibias.n44 gnd 0.010527f
C4694 commonsourceibias.n45 gnd 0.00772f
C4695 commonsourceibias.n46 gnd 0.00772f
C4696 commonsourceibias.n47 gnd 0.00772f
C4697 commonsourceibias.n48 gnd 0.010527f
C4698 commonsourceibias.n49 gnd 0.057546f
C4699 commonsourceibias.n50 gnd 0.010598f
C4700 commonsourceibias.n51 gnd 0.009442f
C4701 commonsourceibias.n52 gnd 0.00772f
C4702 commonsourceibias.n53 gnd 0.00772f
C4703 commonsourceibias.n54 gnd 0.00772f
C4704 commonsourceibias.n55 gnd 0.009185f
C4705 commonsourceibias.n56 gnd 0.010651f
C4706 commonsourceibias.n57 gnd 0.057546f
C4707 commonsourceibias.n58 gnd 0.010587f
C4708 commonsourceibias.n59 gnd 0.00772f
C4709 commonsourceibias.n60 gnd 0.00772f
C4710 commonsourceibias.n61 gnd 0.00772f
C4711 commonsourceibias.n62 gnd 0.010457f
C4712 commonsourceibias.n63 gnd 0.057546f
C4713 commonsourceibias.n64 gnd 0.010526f
C4714 commonsourceibias.n65 gnd 0.009515f
C4715 commonsourceibias.n66 gnd 0.00772f
C4716 commonsourceibias.n67 gnd 0.00772f
C4717 commonsourceibias.n68 gnd 0.007831f
C4718 commonsourceibias.n69 gnd 0.008096f
C4719 commonsourceibias.n70 gnd 0.068855f
C4720 commonsourceibias.n71 gnd 0.076384f
C4721 commonsourceibias.t33 gnd 0.016658f
C4722 commonsourceibias.t15 gnd 0.016658f
C4723 commonsourceibias.n72 gnd 0.147197f
C4724 commonsourceibias.n73 gnd 0.12719f
C4725 commonsourceibias.t25 gnd 0.016658f
C4726 commonsourceibias.t31 gnd 0.016658f
C4727 commonsourceibias.n74 gnd 0.147197f
C4728 commonsourceibias.n75 gnd 0.067614f
C4729 commonsourceibias.t21 gnd 0.016658f
C4730 commonsourceibias.t37 gnd 0.016658f
C4731 commonsourceibias.n76 gnd 0.147197f
C4732 commonsourceibias.n77 gnd 0.056488f
C4733 commonsourceibias.t41 gnd 0.016658f
C4734 commonsourceibias.t47 gnd 0.016658f
C4735 commonsourceibias.n78 gnd 0.14769f
C4736 commonsourceibias.t35 gnd 0.016658f
C4737 commonsourceibias.t11 gnd 0.016658f
C4738 commonsourceibias.n79 gnd 0.147197f
C4739 commonsourceibias.n80 gnd 0.13716f
C4740 commonsourceibias.t45 gnd 0.016658f
C4741 commonsourceibias.t27 gnd 0.016658f
C4742 commonsourceibias.n81 gnd 0.147197f
C4743 commonsourceibias.n82 gnd 0.056488f
C4744 commonsourceibias.n83 gnd 0.068401f
C4745 commonsourceibias.n84 gnd 0.00772f
C4746 commonsourceibias.t50 gnd 0.144227f
C4747 commonsourceibias.t69 gnd 0.144227f
C4748 commonsourceibias.n85 gnd 0.057546f
C4749 commonsourceibias.n86 gnd 0.00772f
C4750 commonsourceibias.t67 gnd 0.144227f
C4751 commonsourceibias.n87 gnd 0.057546f
C4752 commonsourceibias.n88 gnd 0.00772f
C4753 commonsourceibias.t78 gnd 0.144227f
C4754 commonsourceibias.n89 gnd 0.057546f
C4755 commonsourceibias.n90 gnd 0.038863f
C4756 commonsourceibias.t64 gnd 0.144227f
C4757 commonsourceibias.t62 gnd 0.162743f
C4758 commonsourceibias.n91 gnd 0.066782f
C4759 commonsourceibias.n92 gnd 0.069137f
C4760 commonsourceibias.n93 gnd 0.009515f
C4761 commonsourceibias.n94 gnd 0.010526f
C4762 commonsourceibias.n95 gnd 0.00772f
C4763 commonsourceibias.n96 gnd 0.00772f
C4764 commonsourceibias.n97 gnd 0.010457f
C4765 commonsourceibias.n98 gnd 0.006245f
C4766 commonsourceibias.n99 gnd 0.010587f
C4767 commonsourceibias.n100 gnd 0.00772f
C4768 commonsourceibias.n101 gnd 0.00772f
C4769 commonsourceibias.n102 gnd 0.010651f
C4770 commonsourceibias.n103 gnd 0.009185f
C4771 commonsourceibias.n104 gnd 0.007453f
C4772 commonsourceibias.n105 gnd 0.00772f
C4773 commonsourceibias.n106 gnd 0.00772f
C4774 commonsourceibias.n107 gnd 0.009442f
C4775 commonsourceibias.n108 gnd 0.010598f
C4776 commonsourceibias.n109 gnd 0.057546f
C4777 commonsourceibias.n110 gnd 0.010527f
C4778 commonsourceibias.n111 gnd 0.007683f
C4779 commonsourceibias.n112 gnd 0.055804f
C4780 commonsourceibias.n113 gnd 0.007683f
C4781 commonsourceibias.n114 gnd 0.010527f
C4782 commonsourceibias.n115 gnd 0.057546f
C4783 commonsourceibias.n116 gnd 0.010598f
C4784 commonsourceibias.n117 gnd 0.009442f
C4785 commonsourceibias.n118 gnd 0.00772f
C4786 commonsourceibias.n119 gnd 0.00772f
C4787 commonsourceibias.n120 gnd 0.00772f
C4788 commonsourceibias.n121 gnd 0.009185f
C4789 commonsourceibias.n122 gnd 0.010651f
C4790 commonsourceibias.n123 gnd 0.057546f
C4791 commonsourceibias.n124 gnd 0.010587f
C4792 commonsourceibias.n125 gnd 0.00772f
C4793 commonsourceibias.n126 gnd 0.00772f
C4794 commonsourceibias.n127 gnd 0.00772f
C4795 commonsourceibias.n128 gnd 0.010457f
C4796 commonsourceibias.n129 gnd 0.057546f
C4797 commonsourceibias.n130 gnd 0.010526f
C4798 commonsourceibias.n131 gnd 0.009515f
C4799 commonsourceibias.n132 gnd 0.00772f
C4800 commonsourceibias.n133 gnd 0.00772f
C4801 commonsourceibias.n134 gnd 0.007831f
C4802 commonsourceibias.n135 gnd 0.008096f
C4803 commonsourceibias.n136 gnd 0.068855f
C4804 commonsourceibias.n137 gnd 0.04456f
C4805 commonsourceibias.n138 gnd 0.010301f
C4806 commonsourceibias.t72 gnd 0.144227f
C4807 commonsourceibias.n139 gnd 0.057546f
C4808 commonsourceibias.n140 gnd 0.00772f
C4809 commonsourceibias.t49 gnd 0.144227f
C4810 commonsourceibias.n141 gnd 0.006245f
C4811 commonsourceibias.n142 gnd 0.00772f
C4812 commonsourceibias.t95 gnd 0.144227f
C4813 commonsourceibias.n143 gnd 0.007453f
C4814 commonsourceibias.n144 gnd 0.00772f
C4815 commonsourceibias.t66 gnd 0.144227f
C4816 commonsourceibias.n145 gnd 0.057546f
C4817 commonsourceibias.t77 gnd 0.144227f
C4818 commonsourceibias.n146 gnd 0.006235f
C4819 commonsourceibias.n147 gnd 0.00772f
C4820 commonsourceibias.t91 gnd 0.144227f
C4821 commonsourceibias.t60 gnd 0.144227f
C4822 commonsourceibias.n148 gnd 0.057546f
C4823 commonsourceibias.n149 gnd 0.00772f
C4824 commonsourceibias.t58 gnd 0.144227f
C4825 commonsourceibias.n150 gnd 0.057546f
C4826 commonsourceibias.n151 gnd 0.00772f
C4827 commonsourceibias.t68 gnd 0.144227f
C4828 commonsourceibias.n152 gnd 0.057546f
C4829 commonsourceibias.n153 gnd 0.038863f
C4830 commonsourceibias.t57 gnd 0.144227f
C4831 commonsourceibias.t54 gnd 0.162743f
C4832 commonsourceibias.n154 gnd 0.066782f
C4833 commonsourceibias.n155 gnd 0.069137f
C4834 commonsourceibias.n156 gnd 0.009515f
C4835 commonsourceibias.n157 gnd 0.010526f
C4836 commonsourceibias.n158 gnd 0.00772f
C4837 commonsourceibias.n159 gnd 0.00772f
C4838 commonsourceibias.n160 gnd 0.010457f
C4839 commonsourceibias.n161 gnd 0.006245f
C4840 commonsourceibias.n162 gnd 0.010587f
C4841 commonsourceibias.n163 gnd 0.00772f
C4842 commonsourceibias.n164 gnd 0.00772f
C4843 commonsourceibias.n165 gnd 0.010651f
C4844 commonsourceibias.n166 gnd 0.009185f
C4845 commonsourceibias.n167 gnd 0.007453f
C4846 commonsourceibias.n168 gnd 0.00772f
C4847 commonsourceibias.n169 gnd 0.00772f
C4848 commonsourceibias.n170 gnd 0.009442f
C4849 commonsourceibias.n171 gnd 0.010598f
C4850 commonsourceibias.n172 gnd 0.057546f
C4851 commonsourceibias.n173 gnd 0.010527f
C4852 commonsourceibias.n174 gnd 0.00772f
C4853 commonsourceibias.n175 gnd 0.00772f
C4854 commonsourceibias.n176 gnd 0.00772f
C4855 commonsourceibias.n177 gnd 0.010527f
C4856 commonsourceibias.n178 gnd 0.057546f
C4857 commonsourceibias.n179 gnd 0.010598f
C4858 commonsourceibias.n180 gnd 0.009442f
C4859 commonsourceibias.n181 gnd 0.00772f
C4860 commonsourceibias.n182 gnd 0.00772f
C4861 commonsourceibias.n183 gnd 0.00772f
C4862 commonsourceibias.n184 gnd 0.009185f
C4863 commonsourceibias.n185 gnd 0.010651f
C4864 commonsourceibias.n186 gnd 0.057546f
C4865 commonsourceibias.n187 gnd 0.010587f
C4866 commonsourceibias.n188 gnd 0.00772f
C4867 commonsourceibias.n189 gnd 0.00772f
C4868 commonsourceibias.n190 gnd 0.00772f
C4869 commonsourceibias.n191 gnd 0.010457f
C4870 commonsourceibias.n192 gnd 0.057546f
C4871 commonsourceibias.n193 gnd 0.010526f
C4872 commonsourceibias.n194 gnd 0.009515f
C4873 commonsourceibias.n195 gnd 0.00772f
C4874 commonsourceibias.n196 gnd 0.00772f
C4875 commonsourceibias.n197 gnd 0.007831f
C4876 commonsourceibias.n198 gnd 0.008096f
C4877 commonsourceibias.t61 gnd 0.155981f
C4878 commonsourceibias.n199 gnd 0.068855f
C4879 commonsourceibias.n200 gnd 0.023432f
C4880 commonsourceibias.n201 gnd 0.388694f
C4881 commonsourceibias.n202 gnd 0.010301f
C4882 commonsourceibias.t84 gnd 0.155981f
C4883 commonsourceibias.t92 gnd 0.144227f
C4884 commonsourceibias.n203 gnd 0.057546f
C4885 commonsourceibias.n204 gnd 0.00772f
C4886 commonsourceibias.t51 gnd 0.144227f
C4887 commonsourceibias.n205 gnd 0.006245f
C4888 commonsourceibias.n206 gnd 0.00772f
C4889 commonsourceibias.t63 gnd 0.144227f
C4890 commonsourceibias.n207 gnd 0.007453f
C4891 commonsourceibias.n208 gnd 0.00772f
C4892 commonsourceibias.t48 gnd 0.144227f
C4893 commonsourceibias.n209 gnd 0.006235f
C4894 commonsourceibias.n210 gnd 0.00772f
C4895 commonsourceibias.t94 gnd 0.144227f
C4896 commonsourceibias.t83 gnd 0.144227f
C4897 commonsourceibias.n211 gnd 0.057546f
C4898 commonsourceibias.n212 gnd 0.00772f
C4899 commonsourceibias.t80 gnd 0.144227f
C4900 commonsourceibias.n213 gnd 0.057546f
C4901 commonsourceibias.n214 gnd 0.00772f
C4902 commonsourceibias.t90 gnd 0.144227f
C4903 commonsourceibias.n215 gnd 0.057546f
C4904 commonsourceibias.n216 gnd 0.038863f
C4905 commonsourceibias.t59 gnd 0.144227f
C4906 commonsourceibias.t75 gnd 0.162743f
C4907 commonsourceibias.n217 gnd 0.066782f
C4908 commonsourceibias.n218 gnd 0.069137f
C4909 commonsourceibias.n219 gnd 0.009515f
C4910 commonsourceibias.n220 gnd 0.010526f
C4911 commonsourceibias.n221 gnd 0.00772f
C4912 commonsourceibias.n222 gnd 0.00772f
C4913 commonsourceibias.n223 gnd 0.010457f
C4914 commonsourceibias.n224 gnd 0.006245f
C4915 commonsourceibias.n225 gnd 0.010587f
C4916 commonsourceibias.n226 gnd 0.00772f
C4917 commonsourceibias.n227 gnd 0.00772f
C4918 commonsourceibias.n228 gnd 0.010651f
C4919 commonsourceibias.n229 gnd 0.009185f
C4920 commonsourceibias.n230 gnd 0.007453f
C4921 commonsourceibias.n231 gnd 0.00772f
C4922 commonsourceibias.n232 gnd 0.00772f
C4923 commonsourceibias.n233 gnd 0.009442f
C4924 commonsourceibias.n234 gnd 0.010598f
C4925 commonsourceibias.n235 gnd 0.057546f
C4926 commonsourceibias.n236 gnd 0.010527f
C4927 commonsourceibias.n237 gnd 0.007683f
C4928 commonsourceibias.t17 gnd 0.016658f
C4929 commonsourceibias.t9 gnd 0.016658f
C4930 commonsourceibias.n238 gnd 0.14769f
C4931 commonsourceibias.t19 gnd 0.016658f
C4932 commonsourceibias.t5 gnd 0.016658f
C4933 commonsourceibias.n239 gnd 0.147197f
C4934 commonsourceibias.n240 gnd 0.13716f
C4935 commonsourceibias.t43 gnd 0.016658f
C4936 commonsourceibias.t13 gnd 0.016658f
C4937 commonsourceibias.n241 gnd 0.147197f
C4938 commonsourceibias.n242 gnd 0.056488f
C4939 commonsourceibias.n243 gnd 0.010301f
C4940 commonsourceibias.t22 gnd 0.144227f
C4941 commonsourceibias.n244 gnd 0.057546f
C4942 commonsourceibias.n245 gnd 0.00772f
C4943 commonsourceibias.t38 gnd 0.144227f
C4944 commonsourceibias.n246 gnd 0.006245f
C4945 commonsourceibias.n247 gnd 0.00772f
C4946 commonsourceibias.t0 gnd 0.144227f
C4947 commonsourceibias.n248 gnd 0.007453f
C4948 commonsourceibias.n249 gnd 0.00772f
C4949 commonsourceibias.t6 gnd 0.144227f
C4950 commonsourceibias.n250 gnd 0.006235f
C4951 commonsourceibias.n251 gnd 0.00772f
C4952 commonsourceibias.t12 gnd 0.144227f
C4953 commonsourceibias.t42 gnd 0.144227f
C4954 commonsourceibias.n252 gnd 0.057546f
C4955 commonsourceibias.n253 gnd 0.00772f
C4956 commonsourceibias.t4 gnd 0.144227f
C4957 commonsourceibias.n254 gnd 0.057546f
C4958 commonsourceibias.n255 gnd 0.00772f
C4959 commonsourceibias.t18 gnd 0.144227f
C4960 commonsourceibias.n256 gnd 0.057546f
C4961 commonsourceibias.n257 gnd 0.038863f
C4962 commonsourceibias.t8 gnd 0.144227f
C4963 commonsourceibias.t16 gnd 0.162743f
C4964 commonsourceibias.n258 gnd 0.066782f
C4965 commonsourceibias.n259 gnd 0.069137f
C4966 commonsourceibias.n260 gnd 0.009515f
C4967 commonsourceibias.n261 gnd 0.010526f
C4968 commonsourceibias.n262 gnd 0.00772f
C4969 commonsourceibias.n263 gnd 0.00772f
C4970 commonsourceibias.n264 gnd 0.010457f
C4971 commonsourceibias.n265 gnd 0.006245f
C4972 commonsourceibias.n266 gnd 0.010587f
C4973 commonsourceibias.n267 gnd 0.00772f
C4974 commonsourceibias.n268 gnd 0.00772f
C4975 commonsourceibias.n269 gnd 0.010651f
C4976 commonsourceibias.n270 gnd 0.009185f
C4977 commonsourceibias.n271 gnd 0.007453f
C4978 commonsourceibias.n272 gnd 0.00772f
C4979 commonsourceibias.n273 gnd 0.00772f
C4980 commonsourceibias.n274 gnd 0.009442f
C4981 commonsourceibias.n275 gnd 0.010598f
C4982 commonsourceibias.n276 gnd 0.057546f
C4983 commonsourceibias.n277 gnd 0.010527f
C4984 commonsourceibias.n278 gnd 0.00772f
C4985 commonsourceibias.n279 gnd 0.00772f
C4986 commonsourceibias.n280 gnd 0.00772f
C4987 commonsourceibias.n281 gnd 0.010527f
C4988 commonsourceibias.n282 gnd 0.057546f
C4989 commonsourceibias.n283 gnd 0.010598f
C4990 commonsourceibias.t28 gnd 0.144227f
C4991 commonsourceibias.n284 gnd 0.057546f
C4992 commonsourceibias.n285 gnd 0.009442f
C4993 commonsourceibias.n286 gnd 0.00772f
C4994 commonsourceibias.n287 gnd 0.00772f
C4995 commonsourceibias.n288 gnd 0.00772f
C4996 commonsourceibias.n289 gnd 0.009185f
C4997 commonsourceibias.n290 gnd 0.010651f
C4998 commonsourceibias.n291 gnd 0.057546f
C4999 commonsourceibias.n292 gnd 0.010587f
C5000 commonsourceibias.n293 gnd 0.00772f
C5001 commonsourceibias.n294 gnd 0.00772f
C5002 commonsourceibias.n295 gnd 0.00772f
C5003 commonsourceibias.n296 gnd 0.010457f
C5004 commonsourceibias.n297 gnd 0.057546f
C5005 commonsourceibias.n298 gnd 0.010526f
C5006 commonsourceibias.n299 gnd 0.009515f
C5007 commonsourceibias.n300 gnd 0.00772f
C5008 commonsourceibias.n301 gnd 0.00772f
C5009 commonsourceibias.n302 gnd 0.007831f
C5010 commonsourceibias.n303 gnd 0.008096f
C5011 commonsourceibias.t2 gnd 0.155981f
C5012 commonsourceibias.n304 gnd 0.068855f
C5013 commonsourceibias.n305 gnd 0.076384f
C5014 commonsourceibias.t23 gnd 0.016658f
C5015 commonsourceibias.t3 gnd 0.016658f
C5016 commonsourceibias.n306 gnd 0.147197f
C5017 commonsourceibias.n307 gnd 0.12719f
C5018 commonsourceibias.t1 gnd 0.016658f
C5019 commonsourceibias.t39 gnd 0.016658f
C5020 commonsourceibias.n308 gnd 0.147197f
C5021 commonsourceibias.n309 gnd 0.067614f
C5022 commonsourceibias.t7 gnd 0.016658f
C5023 commonsourceibias.t29 gnd 0.016658f
C5024 commonsourceibias.n310 gnd 0.147197f
C5025 commonsourceibias.n311 gnd 0.056488f
C5026 commonsourceibias.n312 gnd 0.068401f
C5027 commonsourceibias.n313 gnd 0.055804f
C5028 commonsourceibias.n314 gnd 0.007683f
C5029 commonsourceibias.n315 gnd 0.010527f
C5030 commonsourceibias.n316 gnd 0.057546f
C5031 commonsourceibias.n317 gnd 0.010598f
C5032 commonsourceibias.t88 gnd 0.144227f
C5033 commonsourceibias.n318 gnd 0.057546f
C5034 commonsourceibias.n319 gnd 0.009442f
C5035 commonsourceibias.n320 gnd 0.00772f
C5036 commonsourceibias.n321 gnd 0.00772f
C5037 commonsourceibias.n322 gnd 0.00772f
C5038 commonsourceibias.n323 gnd 0.009185f
C5039 commonsourceibias.n324 gnd 0.010651f
C5040 commonsourceibias.n325 gnd 0.057546f
C5041 commonsourceibias.n326 gnd 0.010587f
C5042 commonsourceibias.n327 gnd 0.00772f
C5043 commonsourceibias.n328 gnd 0.00772f
C5044 commonsourceibias.n329 gnd 0.00772f
C5045 commonsourceibias.n330 gnd 0.010457f
C5046 commonsourceibias.n331 gnd 0.057546f
C5047 commonsourceibias.n332 gnd 0.010526f
C5048 commonsourceibias.n333 gnd 0.009515f
C5049 commonsourceibias.n334 gnd 0.00772f
C5050 commonsourceibias.n335 gnd 0.00772f
C5051 commonsourceibias.n336 gnd 0.007831f
C5052 commonsourceibias.n337 gnd 0.008096f
C5053 commonsourceibias.n338 gnd 0.068855f
C5054 commonsourceibias.n339 gnd 0.04456f
C5055 commonsourceibias.n340 gnd 0.010301f
C5056 commonsourceibias.t85 gnd 0.144227f
C5057 commonsourceibias.n341 gnd 0.057546f
C5058 commonsourceibias.n342 gnd 0.00772f
C5059 commonsourceibias.t93 gnd 0.144227f
C5060 commonsourceibias.n343 gnd 0.006245f
C5061 commonsourceibias.n344 gnd 0.00772f
C5062 commonsourceibias.t56 gnd 0.144227f
C5063 commonsourceibias.n345 gnd 0.007453f
C5064 commonsourceibias.n346 gnd 0.00772f
C5065 commonsourceibias.t89 gnd 0.144227f
C5066 commonsourceibias.n347 gnd 0.006235f
C5067 commonsourceibias.n348 gnd 0.00772f
C5068 commonsourceibias.t87 gnd 0.144227f
C5069 commonsourceibias.t74 gnd 0.144227f
C5070 commonsourceibias.n349 gnd 0.057546f
C5071 commonsourceibias.n350 gnd 0.00772f
C5072 commonsourceibias.t70 gnd 0.144227f
C5073 commonsourceibias.n351 gnd 0.057546f
C5074 commonsourceibias.n352 gnd 0.00772f
C5075 commonsourceibias.t82 gnd 0.144227f
C5076 commonsourceibias.n353 gnd 0.057546f
C5077 commonsourceibias.n354 gnd 0.038863f
C5078 commonsourceibias.t52 gnd 0.144227f
C5079 commonsourceibias.t65 gnd 0.162743f
C5080 commonsourceibias.n355 gnd 0.066782f
C5081 commonsourceibias.n356 gnd 0.069137f
C5082 commonsourceibias.n357 gnd 0.009515f
C5083 commonsourceibias.n358 gnd 0.010526f
C5084 commonsourceibias.n359 gnd 0.00772f
C5085 commonsourceibias.n360 gnd 0.00772f
C5086 commonsourceibias.n361 gnd 0.010457f
C5087 commonsourceibias.n362 gnd 0.006245f
C5088 commonsourceibias.n363 gnd 0.010587f
C5089 commonsourceibias.n364 gnd 0.00772f
C5090 commonsourceibias.n365 gnd 0.00772f
C5091 commonsourceibias.n366 gnd 0.010651f
C5092 commonsourceibias.n367 gnd 0.009185f
C5093 commonsourceibias.n368 gnd 0.007453f
C5094 commonsourceibias.n369 gnd 0.00772f
C5095 commonsourceibias.n370 gnd 0.00772f
C5096 commonsourceibias.n371 gnd 0.009442f
C5097 commonsourceibias.n372 gnd 0.010598f
C5098 commonsourceibias.n373 gnd 0.057546f
C5099 commonsourceibias.n374 gnd 0.010527f
C5100 commonsourceibias.n375 gnd 0.00772f
C5101 commonsourceibias.n376 gnd 0.00772f
C5102 commonsourceibias.n377 gnd 0.00772f
C5103 commonsourceibias.n378 gnd 0.010527f
C5104 commonsourceibias.n379 gnd 0.057546f
C5105 commonsourceibias.n380 gnd 0.010598f
C5106 commonsourceibias.t79 gnd 0.144227f
C5107 commonsourceibias.n381 gnd 0.057546f
C5108 commonsourceibias.n382 gnd 0.009442f
C5109 commonsourceibias.n383 gnd 0.00772f
C5110 commonsourceibias.n384 gnd 0.00772f
C5111 commonsourceibias.n385 gnd 0.00772f
C5112 commonsourceibias.n386 gnd 0.009185f
C5113 commonsourceibias.n387 gnd 0.010651f
C5114 commonsourceibias.n388 gnd 0.057546f
C5115 commonsourceibias.n389 gnd 0.010587f
C5116 commonsourceibias.n390 gnd 0.00772f
C5117 commonsourceibias.n391 gnd 0.00772f
C5118 commonsourceibias.n392 gnd 0.00772f
C5119 commonsourceibias.n393 gnd 0.010457f
C5120 commonsourceibias.n394 gnd 0.057546f
C5121 commonsourceibias.n395 gnd 0.010526f
C5122 commonsourceibias.n396 gnd 0.009515f
C5123 commonsourceibias.n397 gnd 0.00772f
C5124 commonsourceibias.n398 gnd 0.00772f
C5125 commonsourceibias.n399 gnd 0.007831f
C5126 commonsourceibias.n400 gnd 0.008096f
C5127 commonsourceibias.t73 gnd 0.155981f
C5128 commonsourceibias.n401 gnd 0.068855f
C5129 commonsourceibias.n402 gnd 0.023432f
C5130 commonsourceibias.n403 gnd 0.212991f
C5131 commonsourceibias.n404 gnd 4.01312f
.ends

