* NGSPICE file created from opamp.ext - technology: sky130A

.subckt opamp output vdd plus minus commonsourceibias outputibias diffpairibias gnd CSoutput
Cload output gnd 0.0p
X0 gnd.t200 gnd.t197 gnd.t199 gnd.t198 sky130_fd_pr__nfet_01v8 ad=2.34 pd=12.78 as=0 ps=0 w=6 l=2
X1 commonsourceibias.t47 commonsourceibias.t46 gnd.t290 gnd.t11 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=2.73 ps=14.78 w=7 l=1
X2 gnd.t273 commonsourceibias.t48 CSoutput.t49 gnd.t0 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X3 gnd.t196 gnd.t194 gnd.t195 gnd.t171 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=0 ps=0 w=7 l=1
X4 vdd.t161 vdd.t159 vdd.t160 vdd.t147 sky130_fd_pr__pfet_01v8_lvt ad=3.12 pd=16.78 as=0 ps=0 w=8 l=0.5
X5 vdd.t172 a_n6308_8799.t36 CSoutput.t86 vdd.t63 sky130_fd_pr__pfet_01v8_lvt ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X6 a_n1986_8322.t23 a_n1986_13878.t48 vdd.t13 vdd.t12 sky130_fd_pr__pfet_01v8_lvt ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X7 a_n1808_13878.t19 a_n1986_13878.t16 a_n1986_13878.t17 vdd.t180 sky130_fd_pr__pfet_01v8_lvt ad=1.485 pd=9.33 as=3.51 ps=18.78 w=9 l=0.5
X8 output.t19 outputibias.t8 gnd.t217 gnd.t216 sky130_fd_pr__nfet_01v8 ad=2.34 pd=12.78 as=2.34 ps=12.78 w=6 l=2
X9 gnd.t72 commonsourceibias.t49 CSoutput.t48 gnd.t46 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X10 vdd.t45 CSoutput.t120 output.t15 gnd.t51 sky130_fd_pr__nfet_01v8_lvt ad=0.825 pd=5.33 as=1.95 ps=10.78 w=5 l=1
X11 a_n1986_13878.t5 a_n1986_13878.t4 a_n1808_13878.t18 vdd.t175 sky130_fd_pr__pfet_01v8_lvt ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X12 a_n1808_13878.t17 a_n1986_13878.t8 a_n1986_13878.t9 vdd.t21 sky130_fd_pr__pfet_01v8_lvt ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X13 vdd.t158 vdd.t156 vdd.t157 vdd.t130 sky130_fd_pr__pfet_01v8_lvt ad=3.51 pd=18.78 as=0 ps=0 w=9 l=0.5
X14 CSoutput.t87 a_n6308_8799.t37 vdd.t173 vdd.t66 sky130_fd_pr__pfet_01v8_lvt ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X15 a_n1808_13878.t7 a_n1986_13878.t49 vdd.t15 vdd.t14 sky130_fd_pr__pfet_01v8_lvt ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X16 vdd.t155 vdd.t153 vdd.t154 vdd.t147 sky130_fd_pr__pfet_01v8_lvt ad=3.12 pd=16.78 as=0 ps=0 w=8 l=0.5
X17 vdd.t152 vdd.t150 vdd.t151 vdd.t98 sky130_fd_pr__pfet_01v8_lvt ad=3.12 pd=16.78 as=0 ps=0 w=8 l=0.5
X18 gnd.t92 commonsourceibias.t44 commonsourceibias.t45 gnd.t61 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X19 vdd.t39 CSoutput.t121 output.t14 gnd.t52 sky130_fd_pr__nfet_01v8_lvt ad=0.825 pd=5.33 as=0.825 ps=5.33 w=5 l=1
X20 CSoutput.t74 a_n6308_8799.t38 vdd.t71 vdd.t0 sky130_fd_pr__pfet_01v8_lvt ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X21 gnd.t62 commonsourceibias.t50 CSoutput.t47 gnd.t61 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X22 gnd.t193 gnd.t191 gnd.t192 gnd.t142 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=0 ps=0 w=7 l=0.5
X23 outputibias.t7 outputibias.t6 gnd.t21 gnd.t20 sky130_fd_pr__nfet_01v8 ad=2.34 pd=12.78 as=2.34 ps=12.78 w=6 l=2
X24 CSoutput.t75 a_n6308_8799.t39 vdd.t73 vdd.t72 sky130_fd_pr__pfet_01v8_lvt ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X25 minus.t4 gnd.t188 gnd.t190 gnd.t189 sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.5
X26 gnd.t187 gnd.t186 plus.t4 gnd.t142 sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.5
X27 a_n6308_8799.t29 plus.t5 a_n2903_n3924.t25 gnd.t234 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.5
X28 gnd.t185 gnd.t183 gnd.t184 gnd.t138 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=0 ps=0 w=7 l=0.5
X29 a_n1986_8322.t15 a_n1986_13878.t50 a_n6308_8799.t20 vdd.t85 sky130_fd_pr__pfet_01v8_lvt ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X30 gnd.t261 commonsourceibias.t42 commonsourceibias.t43 gnd.t206 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X31 a_n6308_8799.t12 plus.t6 a_n2903_n3924.t24 gnd.t89 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.5
X32 CSoutput.t46 commonsourceibias.t51 gnd.t58 gnd.t4 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X33 CSoutput.t122 a_n1986_8322.t0 sky130_fd_pr__cap_mim_m3_1 l=12 w=12
X34 gnd.t29 commonsourceibias.t40 commonsourceibias.t41 gnd.t22 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X35 CSoutput.t72 a_n6308_8799.t40 vdd.t68 vdd.t60 sky130_fd_pr__pfet_01v8_lvt ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X36 vdd.t70 a_n6308_8799.t41 CSoutput.t73 vdd.t69 sky130_fd_pr__pfet_01v8_lvt ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X37 a_n6308_8799.t21 a_n1986_13878.t51 a_n1986_8322.t14 vdd.t180 sky130_fd_pr__pfet_01v8_lvt ad=1.485 pd=9.33 as=3.51 ps=18.78 w=9 l=0.5
X38 CSoutput.t52 a_n6308_8799.t42 vdd.t9 vdd.t8 sky130_fd_pr__pfet_01v8_lvt ad=1.32 pd=8.33 as=3.12 ps=16.78 w=8 l=0.5
X39 vdd.t11 a_n6308_8799.t43 CSoutput.t53 vdd.t10 sky130_fd_pr__pfet_01v8_lvt ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X40 a_n2903_n3924.t54 minus.t5 a_n1986_13878.t47 gnd.t33 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.5
X41 CSoutput.t45 commonsourceibias.t52 gnd.t215 gnd.t68 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X42 a_n2903_n3924.t1 diffpairibias.t16 gnd.t10 gnd.t9 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=2.73 ps=14.78 w=7 l=1
X43 vdd.t149 vdd.t146 vdd.t148 vdd.t147 sky130_fd_pr__pfet_01v8_lvt ad=3.12 pd=16.78 as=0 ps=0 w=8 l=0.5
X44 a_n1986_13878.t44 minus.t6 a_n2903_n3924.t53 gnd.t209 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.5
X45 a_n2903_n3924.t23 plus.t7 a_n6308_8799.t5 gnd.t59 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.5
X46 output.t13 CSoutput.t123 vdd.t40 gnd.t224 sky130_fd_pr__nfet_01v8_lvt ad=0.825 pd=5.33 as=0.825 ps=5.33 w=5 l=1
X47 vdd.t50 CSoutput.t124 output.t12 gnd.t225 sky130_fd_pr__nfet_01v8_lvt ad=0.825 pd=5.33 as=0.825 ps=5.33 w=5 l=1
X48 CSoutput.t44 commonsourceibias.t53 gnd.t65 gnd.t64 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X49 a_n2903_n3924.t22 plus.t8 a_n6308_8799.t23 gnd.t219 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.5
X50 a_n2903_n3924.t52 minus.t7 a_n1986_13878.t39 gnd.t241 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.5
X51 CSoutput.t110 a_n6308_8799.t44 vdd.t222 vdd.t32 sky130_fd_pr__pfet_01v8_lvt ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X52 CSoutput.t111 a_n6308_8799.t45 vdd.t223 vdd.t66 sky130_fd_pr__pfet_01v8_lvt ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X53 vdd.t145 vdd.t143 vdd.t144 vdd.t87 sky130_fd_pr__pfet_01v8_lvt ad=3.12 pd=16.78 as=0 ps=0 w=8 l=0.5
X54 CSoutput.t43 commonsourceibias.t54 gnd.t12 gnd.t11 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=2.73 ps=14.78 w=7 l=1
X55 CSoutput.t114 a_n6308_8799.t46 vdd.t226 vdd.t72 sky130_fd_pr__pfet_01v8_lvt ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X56 a_n2903_n3924.t51 minus.t8 a_n1986_13878.t38 gnd.t240 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.5
X57 a_n1808_13878.t16 a_n1986_13878.t22 a_n1986_13878.t23 vdd.t79 sky130_fd_pr__pfet_01v8_lvt ad=1.485 pd=9.33 as=3.51 ps=18.78 w=9 l=0.5
X58 vdd.t227 a_n6308_8799.t47 CSoutput.t115 vdd.t10 sky130_fd_pr__pfet_01v8_lvt ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X59 diffpairibias.t15 diffpairibias.t14 gnd.t283 gnd.t282 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=2.73 ps=14.78 w=7 l=1
X60 a_n1986_13878.t15 a_n1986_13878.t14 a_n1808_13878.t15 vdd.t192 sky130_fd_pr__pfet_01v8_lvt ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X61 CSoutput.t62 a_n6308_8799.t48 vdd.t35 vdd.t34 sky130_fd_pr__pfet_01v8_lvt ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X62 gnd.t182 gnd.t180 gnd.t181 gnd.t171 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=0 ps=0 w=7 l=1
X63 vdd.t142 vdd.t140 vdd.t141 vdd.t115 sky130_fd_pr__pfet_01v8_lvt ad=3.51 pd=18.78 as=0 ps=0 w=9 l=0.5
X64 gnd.t179 gnd.t177 plus.t3 gnd.t178 sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.39 ps=2.78 w=1 l=0.5
X65 a_n1986_13878.t37 minus.t9 a_n2903_n3924.t50 gnd.t26 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=2.73 ps=14.78 w=7 l=0.5
X66 gnd.t47 commonsourceibias.t55 CSoutput.t42 gnd.t46 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X67 gnd.t28 commonsourceibias.t56 CSoutput.t41 gnd.t27 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X68 diffpairibias.t13 diffpairibias.t12 gnd.t37 gnd.t36 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=2.73 ps=14.78 w=7 l=1
X69 gnd.t287 commonsourceibias.t57 CSoutput.t40 gnd.t22 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X70 commonsourceibias.t39 commonsourceibias.t38 gnd.t90 gnd.t4 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X71 vdd.t36 a_n6308_8799.t49 CSoutput.t63 vdd.t10 sky130_fd_pr__pfet_01v8_lvt ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X72 vdd.t43 CSoutput.t125 output.t11 gnd.t75 sky130_fd_pr__nfet_01v8_lvt ad=0.825 pd=5.33 as=0.825 ps=5.33 w=5 l=1
X73 vdd.t218 a_n6308_8799.t50 CSoutput.t108 vdd.t213 sky130_fd_pr__pfet_01v8_lvt ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X74 CSoutput.t109 a_n6308_8799.t51 vdd.t219 vdd.t8 sky130_fd_pr__pfet_01v8_lvt ad=1.32 pd=8.33 as=3.12 ps=16.78 w=8 l=0.5
X75 plus.t2 gnd.t174 gnd.t176 gnd.t175 sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.5
X76 vdd.t31 a_n6308_8799.t52 CSoutput.t60 vdd.t2 sky130_fd_pr__pfet_01v8_lvt ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X77 gnd.t280 commonsourceibias.t58 CSoutput.t39 gnd.t83 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X78 a_n6308_8799.t26 plus.t9 a_n2903_n3924.t21 gnd.t232 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.5
X79 commonsourceibias.t37 commonsourceibias.t36 gnd.t208 gnd.t16 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X80 CSoutput.t61 a_n6308_8799.t53 vdd.t33 vdd.t32 sky130_fd_pr__pfet_01v8_lvt ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X81 CSoutput.t92 a_n6308_8799.t54 vdd.t190 vdd.t189 sky130_fd_pr__pfet_01v8_lvt ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X82 a_n2903_n3924.t26 diffpairibias.t17 gnd.t35 gnd.t34 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=2.73 ps=14.78 w=7 l=1
X83 gnd.t211 commonsourceibias.t34 commonsourceibias.t35 gnd.t83 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X84 CSoutput.t93 a_n6308_8799.t55 vdd.t191 vdd.t189 sky130_fd_pr__pfet_01v8_lvt ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X85 a_n2903_n3924.t49 minus.t10 a_n1986_13878.t36 gnd.t239 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.5
X86 vdd.t216 a_n6308_8799.t56 CSoutput.t106 vdd.t29 sky130_fd_pr__pfet_01v8_lvt ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X87 a_n2903_n3924.t20 plus.t10 a_n6308_8799.t24 gnd.t220 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.5
X88 a_n1986_13878.t43 minus.t11 a_n2903_n3924.t48 gnd.t93 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.5
X89 gnd.t88 commonsourceibias.t32 commonsourceibias.t33 gnd.t87 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=1.155 ps=7.33 w=7 l=1
X90 commonsourceibias.t31 commonsourceibias.t30 gnd.t267 gnd.t64 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X91 a_n1986_13878.t7 a_n1986_13878.t6 a_n1808_13878.t14 vdd.t85 sky130_fd_pr__pfet_01v8_lvt ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X92 outputibias.t5 outputibias.t4 gnd.t289 gnd.t288 sky130_fd_pr__nfet_01v8 ad=2.34 pd=12.78 as=2.34 ps=12.78 w=6 l=2
X93 a_n1986_13878.t19 a_n1986_13878.t18 a_n1808_13878.t13 vdd.t76 sky130_fd_pr__pfet_01v8_lvt ad=3.51 pd=18.78 as=1.485 ps=9.33 w=9 l=0.5
X94 vdd.t217 a_n6308_8799.t57 CSoutput.t107 vdd.t69 sky130_fd_pr__pfet_01v8_lvt ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X95 vdd.t28 a_n6308_8799.t58 CSoutput.t58 vdd.t24 sky130_fd_pr__pfet_01v8_lvt ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X96 a_n6308_8799.t22 a_n1986_13878.t52 a_n1986_8322.t13 vdd.t181 sky130_fd_pr__pfet_01v8_lvt ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X97 CSoutput.t38 commonsourceibias.t59 gnd.t91 gnd.t68 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X98 vdd.t30 a_n6308_8799.t59 CSoutput.t59 vdd.t29 sky130_fd_pr__pfet_01v8_lvt ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X99 a_n2903_n3924.t47 minus.t12 a_n1986_13878.t45 gnd.t60 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=1.155 ps=7.33 w=7 l=0.5
X100 CSoutput.t37 commonsourceibias.t60 gnd.t245 gnd.t18 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X101 vdd.t187 a_n6308_8799.t60 CSoutput.t90 vdd.t186 sky130_fd_pr__pfet_01v8_lvt ad=3.12 pd=16.78 as=1.32 ps=8.33 w=8 l=0.5
X102 gnd.t250 commonsourceibias.t61 CSoutput.t36 gnd.t87 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=1.155 ps=7.33 w=7 l=1
X103 gnd.t173 gnd.t170 gnd.t172 gnd.t171 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=0 ps=0 w=7 l=1
X104 commonsourceibias.t29 commonsourceibias.t28 gnd.t86 gnd.t81 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X105 CSoutput.t91 a_n6308_8799.t61 vdd.t188 vdd.t166 sky130_fd_pr__pfet_01v8_lvt ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X106 CSoutput.t35 commonsourceibias.t62 gnd.t259 gnd.t11 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=2.73 ps=14.78 w=7 l=1
X107 CSoutput.t126 a_n1986_8322.t1 sky130_fd_pr__cap_mim_m3_1 l=12 w=12
X108 outputibias.t3 outputibias.t2 gnd.t279 gnd.t278 sky130_fd_pr__nfet_01v8 ad=2.34 pd=12.78 as=2.34 ps=12.78 w=6 l=2
X109 vdd.t214 a_n6308_8799.t62 CSoutput.t104 vdd.t213 sky130_fd_pr__pfet_01v8_lvt ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X110 vdd.t139 vdd.t137 vdd.t138 vdd.t123 sky130_fd_pr__pfet_01v8_lvt ad=3.51 pd=18.78 as=0 ps=0 w=9 l=0.5
X111 vdd.t136 vdd.t133 vdd.t135 vdd.t134 sky130_fd_pr__pfet_01v8_lvt ad=3.51 pd=18.78 as=0 ps=0 w=9 l=0.5
X112 a_n1986_13878.t46 minus.t13 a_n2903_n3924.t46 gnd.t80 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.5
X113 a_n2903_n3924.t30 diffpairibias.t18 gnd.t238 gnd.t237 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=2.73 ps=14.78 w=7 l=1
X114 vdd.t132 vdd.t129 vdd.t131 vdd.t130 sky130_fd_pr__pfet_01v8_lvt ad=3.51 pd=18.78 as=0 ps=0 w=9 l=0.5
X115 commonsourceibias.t27 commonsourceibias.t26 gnd.t19 gnd.t18 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X116 vdd.t183 a_n1986_13878.t53 a_n1986_8322.t22 vdd.t182 sky130_fd_pr__pfet_01v8_lvt ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X117 vdd.t128 vdd.t126 vdd.t127 vdd.t119 sky130_fd_pr__pfet_01v8_lvt ad=3.51 pd=18.78 as=0 ps=0 w=9 l=0.5
X118 gnd.t169 gnd.t167 minus.t3 gnd.t168 sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.39 ps=2.78 w=1 l=0.5
X119 a_n2903_n3924.t19 plus.t11 a_n6308_8799.t4 gnd.t50 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.5
X120 CSoutput.t105 a_n6308_8799.t63 vdd.t215 vdd.t189 sky130_fd_pr__pfet_01v8_lvt ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X121 a_n1986_8322.t21 a_n1986_13878.t54 vdd.t18 vdd.t17 sky130_fd_pr__pfet_01v8_lvt ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X122 vdd.t170 a_n6308_8799.t64 CSoutput.t84 vdd.t29 sky130_fd_pr__pfet_01v8_lvt ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X123 gnd.t55 commonsourceibias.t24 commonsourceibias.t25 gnd.t46 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X124 gnd.t246 commonsourceibias.t63 CSoutput.t34 gnd.t27 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X125 vdd.t20 a_n1986_13878.t55 a_n1808_13878.t6 vdd.t19 sky130_fd_pr__pfet_01v8_lvt ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X126 gnd.t23 commonsourceibias.t64 CSoutput.t33 gnd.t22 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X127 a_n1986_13878.t40 minus.t14 a_n2903_n3924.t45 gnd.t242 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.5
X128 a_n6308_8799.t2 plus.t12 a_n2903_n3924.t18 gnd.t32 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=2.73 ps=14.78 w=7 l=0.5
X129 gnd.t25 commonsourceibias.t65 CSoutput.t32 gnd.t24 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=1.155 ps=7.33 w=7 l=1
X130 vdd.t125 vdd.t122 vdd.t124 vdd.t123 sky130_fd_pr__pfet_01v8_lvt ad=3.51 pd=18.78 as=0 ps=0 w=9 l=0.5
X131 diffpairibias.t11 diffpairibias.t10 gnd.t272 gnd.t271 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=2.73 ps=14.78 w=7 l=1
X132 vdd.t44 CSoutput.t127 output.t10 gnd.t76 sky130_fd_pr__nfet_01v8_lvt ad=0.825 pd=5.33 as=0.825 ps=5.33 w=5 l=1
X133 vdd.t121 vdd.t118 vdd.t120 vdd.t119 sky130_fd_pr__pfet_01v8_lvt ad=3.51 pd=18.78 as=0 ps=0 w=9 l=0.5
X134 vdd.t171 a_n6308_8799.t65 CSoutput.t85 vdd.t69 sky130_fd_pr__pfet_01v8_lvt ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X135 gnd.t85 commonsourceibias.t66 CSoutput.t31 gnd.t70 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X136 outputibias.t1 outputibias.t0 gnd.t214 gnd.t213 sky130_fd_pr__nfet_01v8 ad=2.34 pd=12.78 as=2.34 ps=12.78 w=6 l=2
X137 a_n6308_8799.t28 a_n1986_13878.t56 a_n1986_8322.t12 vdd.t37 sky130_fd_pr__pfet_01v8_lvt ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X138 a_n1986_8322.t20 a_n1986_13878.t57 vdd.t221 vdd.t220 sky130_fd_pr__pfet_01v8_lvt ad=3.51 pd=18.78 as=1.485 ps=9.33 w=9 l=0.5
X139 vdd.t117 vdd.t114 vdd.t116 vdd.t115 sky130_fd_pr__pfet_01v8_lvt ad=3.51 pd=18.78 as=0 ps=0 w=9 l=0.5
X140 gnd.t84 commonsourceibias.t67 CSoutput.t30 gnd.t83 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X141 vdd.t201 a_n6308_8799.t66 CSoutput.t102 vdd.t186 sky130_fd_pr__pfet_01v8_lvt ad=3.12 pd=16.78 as=1.32 ps=8.33 w=8 l=0.5
X142 a_n1986_13878.t13 a_n1986_13878.t12 a_n1808_13878.t12 vdd.t38 sky130_fd_pr__pfet_01v8_lvt ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X143 a_n2903_n3924.t44 minus.t15 a_n1986_13878.t30 gnd.t210 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=1.155 ps=7.33 w=7 l=0.5
X144 a_n2903_n3924.t43 minus.t16 a_n1986_13878.t33 gnd.t236 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.5
X145 a_n6308_8799.t0 plus.t13 a_n2903_n3924.t17 gnd.t6 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.5
X146 CSoutput.t128 a_n1986_8322.t3 sky130_fd_pr__cap_mim_m3_1 l=12 w=12
X147 CSoutput.t103 a_n6308_8799.t67 vdd.t202 vdd.t166 sky130_fd_pr__pfet_01v8_lvt ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X148 a_n6308_8799.t16 a_n1986_13878.t58 a_n1986_8322.t11 vdd.t21 sky130_fd_pr__pfet_01v8_lvt ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X149 CSoutput.t29 commonsourceibias.t68 gnd.t264 gnd.t73 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X150 a_n1986_13878.t32 minus.t17 a_n2903_n3924.t42 gnd.t235 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.5
X151 CSoutput.t129 a_n1986_8322.t2 sky130_fd_pr__cap_mim_m3_1 l=12 w=12
X152 a_n1808_13878.t11 a_n1986_13878.t10 a_n1986_13878.t11 vdd.t181 sky130_fd_pr__pfet_01v8_lvt ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X153 vdd.t179 a_n1986_13878.t59 a_n1986_8322.t19 vdd.t178 sky130_fd_pr__pfet_01v8_lvt ad=1.485 pd=9.33 as=3.51 ps=18.78 w=9 l=0.5
X154 gnd.t166 gnd.t163 gnd.t165 gnd.t164 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=0 ps=0 w=7 l=1
X155 a_n2903_n3924.t0 diffpairibias.t19 gnd.t8 gnd.t7 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=2.73 ps=14.78 w=7 l=1
X156 CSoutput.t82 a_n6308_8799.t68 vdd.t168 vdd.t34 sky130_fd_pr__pfet_01v8_lvt ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X157 CSoutput.t28 commonsourceibias.t69 gnd.t256 gnd.t18 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X158 a_n1986_13878.t29 minus.t18 a_n2903_n3924.t41 gnd.t234 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.5
X159 CSoutput.t27 commonsourceibias.t70 gnd.t257 gnd.t56 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X160 a_n2903_n3924.t29 diffpairibias.t20 gnd.t231 gnd.t230 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=2.73 ps=14.78 w=7 l=1
X161 vdd.t169 a_n6308_8799.t69 CSoutput.t83 vdd.t82 sky130_fd_pr__pfet_01v8_lvt ad=3.12 pd=16.78 as=1.32 ps=8.33 w=8 l=0.5
X162 gnd.t249 commonsourceibias.t71 CSoutput.t26 gnd.t87 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=1.155 ps=7.33 w=7 l=1
X163 gnd.t162 gnd.t160 minus.t2 gnd.t161 sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.5
X164 CSoutput.t25 commonsourceibias.t72 gnd.t281 gnd.t44 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X165 vdd.t65 a_n6308_8799.t70 CSoutput.t70 vdd.t57 sky130_fd_pr__pfet_01v8_lvt ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X166 a_n1986_13878.t35 minus.t19 a_n2903_n3924.t40 gnd.t89 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.5
X167 gnd.t159 gnd.t157 gnd.t158 gnd.t117 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=0 ps=0 w=7 l=1
X168 diffpairibias.t9 diffpairibias.t8 gnd.t204 gnd.t203 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=2.73 ps=14.78 w=7 l=1
X169 CSoutput.t71 a_n6308_8799.t71 vdd.t67 vdd.t66 sky130_fd_pr__pfet_01v8_lvt ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X170 a_n2903_n3924.t16 plus.t14 a_n6308_8799.t3 gnd.t33 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.5
X171 CSoutput.t100 a_n6308_8799.t72 vdd.t199 vdd.t26 sky130_fd_pr__pfet_01v8_lvt ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X172 CSoutput.t24 commonsourceibias.t73 gnd.t223 gnd.t222 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=2.73 ps=14.78 w=7 l=1
X173 gnd.t207 commonsourceibias.t74 CSoutput.t23 gnd.t206 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X174 vdd.t113 vdd.t111 vdd.t112 vdd.t94 sky130_fd_pr__pfet_01v8_lvt ad=3.12 pd=16.78 as=0 ps=0 w=8 l=0.5
X175 a_n1808_13878.t5 a_n1986_13878.t60 vdd.t210 vdd.t209 sky130_fd_pr__pfet_01v8_lvt ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X176 vdd.t212 a_n1986_13878.t61 a_n1808_13878.t4 vdd.t211 sky130_fd_pr__pfet_01v8_lvt ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X177 a_n2903_n3924.t39 minus.t20 a_n1986_13878.t42 gnd.t219 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.5
X178 a_n2903_n3924.t15 plus.t15 a_n6308_8799.t32 gnd.t241 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.5
X179 gnd.t212 commonsourceibias.t22 commonsourceibias.t23 gnd.t2 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X180 gnd.t40 commonsourceibias.t75 CSoutput.t22 gnd.t24 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=1.155 ps=7.33 w=7 l=1
X181 output.t9 CSoutput.t130 vdd.t41 gnd.t79 sky130_fd_pr__nfet_01v8_lvt ad=0.825 pd=5.33 as=0.825 ps=5.33 w=5 l=1
X182 a_n6308_8799.t33 plus.t16 a_n2903_n3924.t14 gnd.t233 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.5
X183 a_n2903_n3924.t38 minus.t21 a_n1986_13878.t41 gnd.t77 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.5
X184 gnd.t255 commonsourceibias.t76 CSoutput.t21 gnd.t70 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X185 diffpairibias.t7 diffpairibias.t6 gnd.t275 gnd.t274 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=2.73 ps=14.78 w=7 l=1
X186 CSoutput.t101 a_n6308_8799.t73 vdd.t200 vdd.t34 sky130_fd_pr__pfet_01v8_lvt ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X187 gnd.t71 commonsourceibias.t20 commonsourceibias.t21 gnd.t70 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X188 output.t8 CSoutput.t131 vdd.t54 gnd.t53 sky130_fd_pr__nfet_01v8_lvt ad=0.825 pd=5.33 as=0.825 ps=5.33 w=5 l=1
X189 vdd.t224 a_n6308_8799.t74 CSoutput.t112 vdd.t82 sky130_fd_pr__pfet_01v8_lvt ad=3.12 pd=16.78 as=1.32 ps=8.33 w=8 l=0.5
X190 CSoutput.t20 commonsourceibias.t77 gnd.t266 gnd.t16 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X191 gnd.t156 gnd.t154 gnd.t155 gnd.t117 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=0 ps=0 w=7 l=1
X192 gnd.t150 gnd.t148 gnd.t149 gnd.t95 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=0 ps=0 w=7 l=1
X193 a_n1986_8322.t10 a_n1986_13878.t62 a_n6308_8799.t15 vdd.t175 sky130_fd_pr__pfet_01v8_lvt ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X194 CSoutput.t19 commonsourceibias.t78 gnd.t74 gnd.t73 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X195 vdd.t225 a_n6308_8799.t75 CSoutput.t113 vdd.t213 sky130_fd_pr__pfet_01v8_lvt ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X196 CSoutput.t116 a_n6308_8799.t76 vdd.t228 vdd.t6 sky130_fd_pr__pfet_01v8_lvt ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X197 vdd.t229 a_n6308_8799.t77 CSoutput.t117 vdd.t57 sky130_fd_pr__pfet_01v8_lvt ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X198 vdd.t177 a_n1986_13878.t63 a_n1986_8322.t18 vdd.t176 sky130_fd_pr__pfet_01v8_lvt ad=1.485 pd=9.33 as=3.51 ps=18.78 w=9 l=0.5
X199 plus.t1 gnd.t151 gnd.t153 gnd.t152 sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.5
X200 gnd.t147 gnd.t145 minus.t1 gnd.t146 sky130_fd_pr__nfet_01v8 ad=0.39 pd=2.78 as=0.165 ps=1.33 w=1 l=0.5
X201 gnd.t144 gnd.t141 gnd.t143 gnd.t142 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=0 ps=0 w=7 l=0.5
X202 gnd.t39 commonsourceibias.t18 commonsourceibias.t19 gnd.t38 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X203 a_n1808_13878.t3 a_n1986_13878.t64 vdd.t81 vdd.t80 sky130_fd_pr__pfet_01v8_lvt ad=3.51 pd=18.78 as=1.485 ps=9.33 w=9 l=0.5
X204 gnd.t140 gnd.t137 gnd.t139 gnd.t138 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=0 ps=0 w=7 l=0.5
X205 gnd.t136 gnd.t133 gnd.t135 gnd.t134 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=0 ps=0 w=7 l=1
X206 CSoutput.t18 commonsourceibias.t79 gnd.t260 gnd.t81 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X207 a_n2903_n3924.t27 diffpairibias.t21 gnd.t202 gnd.t201 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=2.73 ps=14.78 w=7 l=1
X208 vdd.t25 a_n6308_8799.t78 CSoutput.t56 vdd.t24 sky130_fd_pr__pfet_01v8_lvt ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X209 vdd.t110 vdd.t108 vdd.t109 vdd.t98 sky130_fd_pr__pfet_01v8_lvt ad=3.12 pd=16.78 as=0 ps=0 w=8 l=0.5
X210 CSoutput.t57 a_n6308_8799.t79 vdd.t27 vdd.t26 sky130_fd_pr__pfet_01v8_lvt ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X211 CSoutput.t17 commonsourceibias.t80 gnd.t57 gnd.t56 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X212 output.t7 CSoutput.t132 vdd.t49 gnd.t54 sky130_fd_pr__nfet_01v8_lvt ad=0.825 pd=5.33 as=0.825 ps=5.33 w=5 l=1
X213 CSoutput.t68 a_n6308_8799.t80 vdd.t62 vdd.t60 sky130_fd_pr__pfet_01v8_lvt ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X214 CSoutput.t133 a_n1986_8322.t1 sky130_fd_pr__cap_mim_m3_1 l=12 w=12
X215 vdd.t107 vdd.t105 vdd.t106 vdd.t94 sky130_fd_pr__pfet_01v8_lvt ad=3.12 pd=16.78 as=0 ps=0 w=8 l=0.5
X216 CSoutput.t16 commonsourceibias.t81 gnd.t78 gnd.t44 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X217 gnd.t132 gnd.t129 gnd.t131 gnd.t130 sky130_fd_pr__nfet_01v8_lvt ad=1.95 pd=10.78 as=0 ps=0 w=5 l=1
X218 a_n1986_8322.t9 a_n1986_13878.t65 a_n6308_8799.t9 vdd.t38 sky130_fd_pr__pfet_01v8_lvt ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X219 vdd.t208 a_n1986_13878.t66 a_n1986_8322.t17 vdd.t207 sky130_fd_pr__pfet_01v8_lvt ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X220 vdd.t64 a_n6308_8799.t81 CSoutput.t69 vdd.t63 sky130_fd_pr__pfet_01v8_lvt ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X221 CSoutput.t98 a_n6308_8799.t82 vdd.t197 vdd.t26 sky130_fd_pr__pfet_01v8_lvt ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X222 gnd.t268 commonsourceibias.t82 CSoutput.t15 gnd.t38 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X223 output.t18 outputibias.t9 gnd.t31 gnd.t30 sky130_fd_pr__nfet_01v8 ad=2.34 pd=12.78 as=2.34 ps=12.78 w=6 l=2
X224 CSoutput.t99 a_n6308_8799.t83 vdd.t198 vdd.t4 sky130_fd_pr__pfet_01v8_lvt ad=1.32 pd=8.33 as=3.12 ps=16.78 w=8 l=0.5
X225 a_n2903_n3924.t13 plus.t17 a_n6308_8799.t34 gnd.t239 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.5
X226 gnd.t128 gnd.t126 gnd.t127 gnd.t113 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=0 ps=0 w=7 l=1
X227 vdd.t42 CSoutput.t134 output.t6 gnd.t13 sky130_fd_pr__nfet_01v8_lvt ad=0.825 pd=5.33 as=0.825 ps=5.33 w=5 l=1
X228 vdd.t195 a_n6308_8799.t84 CSoutput.t96 vdd.t163 sky130_fd_pr__pfet_01v8_lvt ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X229 vdd.t196 a_n6308_8799.t85 CSoutput.t97 vdd.t55 sky130_fd_pr__pfet_01v8_lvt ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X230 a_n2903_n3924.t37 minus.t22 a_n1986_13878.t34 gnd.t220 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.5
X231 a_n6308_8799.t17 plus.t18 a_n2903_n3924.t12 gnd.t93 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.5
X232 gnd.t125 gnd.t123 gnd.t124 gnd.t113 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=0 ps=0 w=7 l=1
X233 output.t17 outputibias.t10 gnd.t252 gnd.t251 sky130_fd_pr__nfet_01v8 ad=2.34 pd=12.78 as=2.34 ps=12.78 w=6 l=2
X234 diffpairibias.t5 diffpairibias.t4 gnd.t277 gnd.t276 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=2.73 ps=14.78 w=7 l=1
X235 vdd.t104 vdd.t101 vdd.t103 vdd.t102 sky130_fd_pr__pfet_01v8_lvt ad=3.51 pd=18.78 as=0 ps=0 w=9 l=0.5
X236 a_n6308_8799.t18 plus.t19 a_n2903_n3924.t11 gnd.t209 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.5
X237 a_n2903_n3924.t36 minus.t23 a_n1986_13878.t27 gnd.t59 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.5
X238 a_n1808_13878.t10 a_n1986_13878.t2 a_n1986_13878.t3 vdd.t16 sky130_fd_pr__pfet_01v8_lvt ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X239 gnd.t254 commonsourceibias.t83 CSoutput.t14 gnd.t206 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X240 CSoutput.t13 commonsourceibias.t84 gnd.t286 gnd.t222 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=2.73 ps=14.78 w=7 l=1
X241 a_n1986_8322.t8 a_n1986_13878.t67 a_n6308_8799.t25 vdd.t192 sky130_fd_pr__pfet_01v8_lvt ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X242 gnd.t244 commonsourceibias.t85 CSoutput.t12 gnd.t2 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X243 gnd.t43 commonsourceibias.t16 commonsourceibias.t17 gnd.t24 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=1.155 ps=7.33 w=7 l=1
X244 vdd.t165 a_n6308_8799.t86 CSoutput.t80 vdd.t163 sky130_fd_pr__pfet_01v8_lvt ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X245 CSoutput.t81 a_n6308_8799.t87 vdd.t167 vdd.t166 sky130_fd_pr__pfet_01v8_lvt ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X246 a_n2903_n3924.t10 plus.t20 a_n6308_8799.t30 gnd.t240 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.5
X247 gnd.t108 gnd.t105 gnd.t107 gnd.t106 sky130_fd_pr__nfet_01v8 ad=2.34 pd=12.78 as=0 ps=0 w=6 l=2
X248 vdd.t53 CSoutput.t135 output.t5 gnd.t14 sky130_fd_pr__nfet_01v8_lvt ad=0.825 pd=5.33 as=0.825 ps=5.33 w=5 l=1
X249 output.t4 CSoutput.t136 vdd.t46 gnd.t15 sky130_fd_pr__nfet_01v8_lvt ad=0.825 pd=5.33 as=0.825 ps=5.33 w=5 l=1
X250 vdd.t59 a_n6308_8799.t88 CSoutput.t66 vdd.t24 sky130_fd_pr__pfet_01v8_lvt ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X251 CSoutput.t67 a_n6308_8799.t89 vdd.t61 vdd.t60 sky130_fd_pr__pfet_01v8_lvt ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X252 a_n1986_8322.t16 a_n1986_13878.t68 vdd.t204 vdd.t203 sky130_fd_pr__pfet_01v8_lvt ad=3.51 pd=18.78 as=1.485 ps=9.33 w=9 l=0.5
X253 vdd.t100 vdd.t97 vdd.t99 vdd.t98 sky130_fd_pr__pfet_01v8_lvt ad=3.12 pd=16.78 as=0 ps=0 w=8 l=0.5
X254 gnd.t122 gnd.t120 gnd.t121 gnd.t95 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=0 ps=0 w=7 l=1
X255 CSoutput.t11 commonsourceibias.t86 gnd.t17 gnd.t16 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X256 a_n6308_8799.t1 plus.t21 a_n2903_n3924.t9 gnd.t26 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=2.73 ps=14.78 w=7 l=0.5
X257 CSoutput.t10 commonsourceibias.t87 gnd.t221 gnd.t66 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X258 gnd.t119 gnd.t116 gnd.t118 gnd.t117 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=0 ps=0 w=7 l=1
X259 a_n2903_n3924.t35 minus.t24 a_n1986_13878.t26 gnd.t50 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.5
X260 output.t3 CSoutput.t137 vdd.t48 gnd.t41 sky130_fd_pr__nfet_01v8_lvt ad=0.825 pd=5.33 as=0.825 ps=5.33 w=5 l=1
X261 vdd.t206 a_n1986_13878.t69 a_n1808_13878.t2 vdd.t205 sky130_fd_pr__pfet_01v8_lvt ad=1.485 pd=9.33 as=3.51 ps=18.78 w=9 l=0.5
X262 CSoutput.t78 a_n6308_8799.t90 vdd.t162 vdd.t4 sky130_fd_pr__pfet_01v8_lvt ad=1.32 pd=8.33 as=3.12 ps=16.78 w=8 l=0.5
X263 vdd.t164 a_n6308_8799.t91 CSoutput.t79 vdd.t163 sky130_fd_pr__pfet_01v8_lvt ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X264 vdd.t56 a_n6308_8799.t92 CSoutput.t64 vdd.t55 sky130_fd_pr__pfet_01v8_lvt ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X265 vdd.t96 vdd.t93 vdd.t95 vdd.t94 sky130_fd_pr__pfet_01v8_lvt ad=3.12 pd=16.78 as=0 ps=0 w=8 l=0.5
X266 a_n1986_8322.t7 a_n1986_13878.t70 a_n6308_8799.t13 vdd.t174 sky130_fd_pr__pfet_01v8_lvt ad=3.51 pd=18.78 as=1.485 ps=9.33 w=9 l=0.5
X267 a_n6308_8799.t35 plus.t22 a_n2903_n3924.t8 gnd.t242 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.5
X268 output.t16 outputibias.t11 gnd.t263 gnd.t262 sky130_fd_pr__nfet_01v8 ad=2.34 pd=12.78 as=2.34 ps=12.78 w=6 l=2
X269 vdd.t92 vdd.t90 vdd.t91 vdd.t87 sky130_fd_pr__pfet_01v8_lvt ad=3.12 pd=16.78 as=0 ps=0 w=8 l=0.5
X270 a_n6308_8799.t14 a_n1986_13878.t71 a_n1986_8322.t6 vdd.t16 sky130_fd_pr__pfet_01v8_lvt ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X271 a_n1808_13878.t1 a_n1986_13878.t72 vdd.t78 vdd.t77 sky130_fd_pr__pfet_01v8_lvt ad=3.51 pd=18.78 as=1.485 ps=9.33 w=9 l=0.5
X272 vdd.t58 a_n6308_8799.t93 CSoutput.t65 vdd.t57 sky130_fd_pr__pfet_01v8_lvt ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X273 CSoutput.t94 a_n6308_8799.t94 vdd.t193 vdd.t32 sky130_fd_pr__pfet_01v8_lvt ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X274 CSoutput.t9 commonsourceibias.t88 gnd.t82 gnd.t81 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X275 a_n1986_13878.t25 minus.t25 a_n2903_n3924.t34 gnd.t232 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.5
X276 commonsourceibias.t15 commonsourceibias.t14 gnd.t45 gnd.t44 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X277 gnd.t1 commonsourceibias.t89 CSoutput.t8 gnd.t0 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X278 vdd.t47 CSoutput.t138 output.t2 gnd.t42 sky130_fd_pr__nfet_01v8_lvt ad=0.825 pd=5.33 as=0.825 ps=5.33 w=5 l=1
X279 a_n2903_n3924.t7 plus.t23 a_n6308_8799.t19 gnd.t210 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=1.155 ps=7.33 w=7 l=0.5
X280 gnd.t63 commonsourceibias.t90 CSoutput.t7 gnd.t38 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X281 a_n6308_8799.t31 plus.t24 a_n2903_n3924.t6 gnd.t235 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.5
X282 CSoutput.t95 a_n6308_8799.t95 vdd.t194 vdd.t6 sky130_fd_pr__pfet_01v8_lvt ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X283 a_n1808_13878.t9 a_n1986_13878.t20 a_n1986_13878.t21 vdd.t37 sky130_fd_pr__pfet_01v8_lvt ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X284 gnd.t115 gnd.t112 gnd.t114 gnd.t113 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=0 ps=0 w=7 l=1
X285 a_n2903_n3924.t55 diffpairibias.t22 gnd.t270 gnd.t269 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=2.73 ps=14.78 w=7 l=1
X286 gnd.t205 commonsourceibias.t91 CSoutput.t6 gnd.t61 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X287 commonsourceibias.t13 commonsourceibias.t12 gnd.t67 gnd.t66 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X288 a_n2903_n3924.t5 plus.t25 a_n6308_8799.t6 gnd.t60 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=1.155 ps=7.33 w=7 l=0.5
X289 CSoutput.t54 a_n6308_8799.t96 vdd.t22 vdd.t0 sky130_fd_pr__pfet_01v8_lvt ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X290 vdd.t23 a_n6308_8799.t97 CSoutput.t55 vdd.t2 sky130_fd_pr__pfet_01v8_lvt ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X291 diffpairibias.t3 diffpairibias.t2 gnd.t285 gnd.t284 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=2.73 ps=14.78 w=7 l=1
X292 a_n6308_8799.t8 a_n1986_13878.t73 a_n1986_8322.t5 vdd.t79 sky130_fd_pr__pfet_01v8_lvt ad=1.485 pd=9.33 as=3.51 ps=18.78 w=9 l=0.5
X293 a_n1986_13878.t1 a_n1986_13878.t0 a_n1808_13878.t8 vdd.t174 sky130_fd_pr__pfet_01v8_lvt ad=3.51 pd=18.78 as=1.485 ps=9.33 w=9 l=0.5
X294 vdd.t230 a_n6308_8799.t98 CSoutput.t118 vdd.t63 sky130_fd_pr__pfet_01v8_lvt ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X295 commonsourceibias.t11 commonsourceibias.t10 gnd.t265 gnd.t73 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X296 gnd.t3 commonsourceibias.t92 CSoutput.t5 gnd.t2 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X297 vdd.t89 vdd.t86 vdd.t88 vdd.t87 sky130_fd_pr__pfet_01v8_lvt ad=3.12 pd=16.78 as=0 ps=0 w=8 l=0.5
X298 vdd.t231 a_n6308_8799.t99 CSoutput.t119 vdd.t186 sky130_fd_pr__pfet_01v8_lvt ad=3.12 pd=16.78 as=1.32 ps=8.33 w=8 l=0.5
X299 gnd.t111 gnd.t109 plus.t0 gnd.t110 sky130_fd_pr__nfet_01v8 ad=0.39 pd=2.78 as=0.165 ps=1.33 w=1 l=0.5
X300 a_n6308_8799.t11 plus.t26 a_n2903_n3924.t4 gnd.t80 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.5
X301 CSoutput.t139 a_n1986_8322.t0 sky130_fd_pr__cap_mim_m3_1 l=12 w=12
X302 diffpairibias.t1 diffpairibias.t0 gnd.t229 gnd.t228 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=2.73 ps=14.78 w=7 l=1
X303 CSoutput.t50 a_n6308_8799.t100 vdd.t5 vdd.t4 sky130_fd_pr__pfet_01v8_lvt ad=1.32 pd=8.33 as=3.12 ps=16.78 w=8 l=0.5
X304 minus.t0 gnd.t102 gnd.t104 gnd.t103 sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.5
X305 CSoutput.t4 commonsourceibias.t93 gnd.t5 gnd.t4 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X306 gnd.t101 gnd.t98 gnd.t100 gnd.t99 sky130_fd_pr__nfet_01v8_lvt ad=1.95 pd=10.78 as=0 ps=0 w=5 l=1
X307 output.t1 CSoutput.t140 vdd.t51 gnd.t48 sky130_fd_pr__nfet_01v8_lvt ad=0.825 pd=5.33 as=0.825 ps=5.33 w=5 l=1
X308 gnd.t97 gnd.t94 gnd.t96 gnd.t95 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=0 ps=0 w=7 l=1
X309 CSoutput.t3 commonsourceibias.t94 gnd.t258 gnd.t66 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X310 commonsourceibias.t9 commonsourceibias.t8 gnd.t69 gnd.t68 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X311 vdd.t75 a_n1986_13878.t74 a_n1808_13878.t0 vdd.t74 sky130_fd_pr__pfet_01v8_lvt ad=1.485 pd=9.33 as=3.51 ps=18.78 w=9 l=0.5
X312 CSoutput.t51 a_n6308_8799.t101 vdd.t7 vdd.t6 sky130_fd_pr__pfet_01v8_lvt ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X313 CSoutput.t2 commonsourceibias.t95 gnd.t218 gnd.t64 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X314 a_n1986_13878.t24 minus.t26 a_n2903_n3924.t33 gnd.t32 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=2.73 ps=14.78 w=7 l=0.5
X315 output.t0 CSoutput.t141 vdd.t52 gnd.t49 sky130_fd_pr__nfet_01v8_lvt ad=1.95 pd=10.78 as=0.825 ps=5.33 w=5 l=1
X316 CSoutput.t88 a_n6308_8799.t102 vdd.t184 vdd.t72 sky130_fd_pr__pfet_01v8_lvt ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X317 vdd.t185 a_n6308_8799.t103 CSoutput.t89 vdd.t55 sky130_fd_pr__pfet_01v8_lvt ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X318 gnd.t248 commonsourceibias.t6 commonsourceibias.t7 gnd.t0 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X319 commonsourceibias.t5 commonsourceibias.t4 gnd.t247 gnd.t56 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X320 CSoutput.t0 a_n6308_8799.t104 vdd.t1 vdd.t0 sky130_fd_pr__pfet_01v8_lvt ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X321 a_n1986_13878.t28 minus.t27 a_n2903_n3924.t32 gnd.t233 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.5
X322 a_n2903_n3924.t3 plus.t27 a_n6308_8799.t10 gnd.t77 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.5
X323 vdd.t3 a_n6308_8799.t105 CSoutput.t1 vdd.t2 sky130_fd_pr__pfet_01v8_lvt ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X324 a_n1986_8322.t4 a_n1986_13878.t75 a_n6308_8799.t7 vdd.t76 sky130_fd_pr__pfet_01v8_lvt ad=3.51 pd=18.78 as=1.485 ps=9.33 w=9 l=0.5
X325 commonsourceibias.t3 commonsourceibias.t2 gnd.t243 gnd.t222 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=2.73 ps=14.78 w=7 l=1
X326 vdd.t83 a_n6308_8799.t106 CSoutput.t76 vdd.t82 sky130_fd_pr__pfet_01v8_lvt ad=3.12 pd=16.78 as=1.32 ps=8.33 w=8 l=0.5
X327 CSoutput.t77 a_n6308_8799.t107 vdd.t84 vdd.t8 sky130_fd_pr__pfet_01v8_lvt ad=1.32 pd=8.33 as=3.12 ps=16.78 w=8 l=0.5
X328 a_n2903_n3924.t2 plus.t28 a_n6308_8799.t27 gnd.t236 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.5
X329 a_n1986_13878.t31 minus.t28 a_n2903_n3924.t31 gnd.t6 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.5
X330 gnd.t253 commonsourceibias.t0 commonsourceibias.t1 gnd.t27 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X331 a_n2903_n3924.t28 diffpairibias.t23 gnd.t227 gnd.t226 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=2.73 ps=14.78 w=7 l=1
R0 gnd.n6348 gnd.n383 1323.14
R1 gnd.n4407 gnd.n4406 939.716
R2 gnd.n6643 gnd.n84 838.452
R3 gnd.n6806 gnd.n80 838.452
R4 gnd.n3452 gnd.n1214 838.452
R5 gnd.n3371 gnd.n1216 838.452
R6 gnd.n4200 gnd.n1083 838.452
R7 gnd.n2627 gnd.n1081 838.452
R8 gnd.n2085 gnd.n829 838.452
R9 gnd.n2148 gnd.n2086 838.452
R10 gnd.n6804 gnd.n86 819.232
R11 gnd.n154 gnd.n82 819.232
R12 gnd.n3807 gnd.n1213 819.232
R13 gnd.n4053 gnd.n1217 819.232
R14 gnd.n4202 gnd.n1078 819.232
R15 gnd.n1994 gnd.n1080 819.232
R16 gnd.n4328 gnd.n4327 819.232
R17 gnd.n4404 gnd.n833 819.232
R18 gnd.n2673 gnd.n1088 771.183
R19 gnd.n4071 gnd.n1191 771.183
R20 gnd.n2677 gnd.n1844 771.183
R21 gnd.n3485 gnd.n1193 771.183
R22 gnd.n5800 gnd.n798 766.379
R23 gnd.n5716 gnd.n800 766.379
R24 gnd.n4916 gnd.n4819 766.379
R25 gnd.n4912 gnd.n4817 766.379
R26 gnd.n5797 gnd.n4409 756.769
R27 gnd.n5766 gnd.n801 756.769
R28 gnd.n5083 gnd.n4726 756.769
R29 gnd.n5081 gnd.n4729 756.769
R30 gnd.n5990 gnd.n596 689.5
R31 gnd.n6347 gnd.n384 689.5
R32 gnd.n6561 gnd.n6559 689.5
R33 gnd.n2046 gnd.n764 689.5
R34 gnd.n599 gnd.n596 585
R35 gnd.n5988 gnd.n596 585
R36 gnd.n5986 gnd.n5985 585
R37 gnd.n5987 gnd.n5986 585
R38 gnd.n5984 gnd.n598 585
R39 gnd.n598 gnd.n597 585
R40 gnd.n5983 gnd.n5982 585
R41 gnd.n5982 gnd.n5981 585
R42 gnd.n604 gnd.n603 585
R43 gnd.n5980 gnd.n604 585
R44 gnd.n5978 gnd.n5977 585
R45 gnd.n5979 gnd.n5978 585
R46 gnd.n5976 gnd.n606 585
R47 gnd.n606 gnd.n605 585
R48 gnd.n5975 gnd.n5974 585
R49 gnd.n5974 gnd.n5973 585
R50 gnd.n612 gnd.n611 585
R51 gnd.n5972 gnd.n612 585
R52 gnd.n5970 gnd.n5969 585
R53 gnd.n5971 gnd.n5970 585
R54 gnd.n5968 gnd.n614 585
R55 gnd.n614 gnd.n613 585
R56 gnd.n5967 gnd.n5966 585
R57 gnd.n5966 gnd.n5965 585
R58 gnd.n620 gnd.n619 585
R59 gnd.n5964 gnd.n620 585
R60 gnd.n5962 gnd.n5961 585
R61 gnd.n5963 gnd.n5962 585
R62 gnd.n5960 gnd.n622 585
R63 gnd.n622 gnd.n621 585
R64 gnd.n5959 gnd.n5958 585
R65 gnd.n5958 gnd.n5957 585
R66 gnd.n628 gnd.n627 585
R67 gnd.n5956 gnd.n628 585
R68 gnd.n5954 gnd.n5953 585
R69 gnd.n5955 gnd.n5954 585
R70 gnd.n5952 gnd.n630 585
R71 gnd.n630 gnd.n629 585
R72 gnd.n5951 gnd.n5950 585
R73 gnd.n5950 gnd.n5949 585
R74 gnd.n636 gnd.n635 585
R75 gnd.n5948 gnd.n636 585
R76 gnd.n5946 gnd.n5945 585
R77 gnd.n5947 gnd.n5946 585
R78 gnd.n5944 gnd.n638 585
R79 gnd.n638 gnd.n637 585
R80 gnd.n5943 gnd.n5942 585
R81 gnd.n5942 gnd.n5941 585
R82 gnd.n644 gnd.n643 585
R83 gnd.n5940 gnd.n644 585
R84 gnd.n5938 gnd.n5937 585
R85 gnd.n5939 gnd.n5938 585
R86 gnd.n5936 gnd.n646 585
R87 gnd.n646 gnd.n645 585
R88 gnd.n5935 gnd.n5934 585
R89 gnd.n5934 gnd.n5933 585
R90 gnd.n652 gnd.n651 585
R91 gnd.n5932 gnd.n652 585
R92 gnd.n5930 gnd.n5929 585
R93 gnd.n5931 gnd.n5930 585
R94 gnd.n5928 gnd.n654 585
R95 gnd.n654 gnd.n653 585
R96 gnd.n5927 gnd.n5926 585
R97 gnd.n5926 gnd.n5925 585
R98 gnd.n660 gnd.n659 585
R99 gnd.n5924 gnd.n660 585
R100 gnd.n5922 gnd.n5921 585
R101 gnd.n5923 gnd.n5922 585
R102 gnd.n5920 gnd.n662 585
R103 gnd.n662 gnd.n661 585
R104 gnd.n5919 gnd.n5918 585
R105 gnd.n5918 gnd.n5917 585
R106 gnd.n668 gnd.n667 585
R107 gnd.n5916 gnd.n668 585
R108 gnd.n5914 gnd.n5913 585
R109 gnd.n5915 gnd.n5914 585
R110 gnd.n5912 gnd.n670 585
R111 gnd.n670 gnd.n669 585
R112 gnd.n5911 gnd.n5910 585
R113 gnd.n5910 gnd.n5909 585
R114 gnd.n676 gnd.n675 585
R115 gnd.n5908 gnd.n676 585
R116 gnd.n5906 gnd.n5905 585
R117 gnd.n5907 gnd.n5906 585
R118 gnd.n5904 gnd.n678 585
R119 gnd.n678 gnd.n677 585
R120 gnd.n5903 gnd.n5902 585
R121 gnd.n5902 gnd.n5901 585
R122 gnd.n684 gnd.n683 585
R123 gnd.n5900 gnd.n684 585
R124 gnd.n5898 gnd.n5897 585
R125 gnd.n5899 gnd.n5898 585
R126 gnd.n5896 gnd.n686 585
R127 gnd.n686 gnd.n685 585
R128 gnd.n5895 gnd.n5894 585
R129 gnd.n5894 gnd.n5893 585
R130 gnd.n692 gnd.n691 585
R131 gnd.n5892 gnd.n692 585
R132 gnd.n5890 gnd.n5889 585
R133 gnd.n5891 gnd.n5890 585
R134 gnd.n5888 gnd.n694 585
R135 gnd.n694 gnd.n693 585
R136 gnd.n5887 gnd.n5886 585
R137 gnd.n5886 gnd.n5885 585
R138 gnd.n700 gnd.n699 585
R139 gnd.n5884 gnd.n700 585
R140 gnd.n5882 gnd.n5881 585
R141 gnd.n5883 gnd.n5882 585
R142 gnd.n5880 gnd.n702 585
R143 gnd.n702 gnd.n701 585
R144 gnd.n5879 gnd.n5878 585
R145 gnd.n5878 gnd.n5877 585
R146 gnd.n708 gnd.n707 585
R147 gnd.n5876 gnd.n708 585
R148 gnd.n5874 gnd.n5873 585
R149 gnd.n5875 gnd.n5874 585
R150 gnd.n5872 gnd.n710 585
R151 gnd.n710 gnd.n709 585
R152 gnd.n5871 gnd.n5870 585
R153 gnd.n5870 gnd.n5869 585
R154 gnd.n716 gnd.n715 585
R155 gnd.n5868 gnd.n716 585
R156 gnd.n5866 gnd.n5865 585
R157 gnd.n5867 gnd.n5866 585
R158 gnd.n5864 gnd.n718 585
R159 gnd.n718 gnd.n717 585
R160 gnd.n5863 gnd.n5862 585
R161 gnd.n5862 gnd.n5861 585
R162 gnd.n724 gnd.n723 585
R163 gnd.n5860 gnd.n724 585
R164 gnd.n5858 gnd.n5857 585
R165 gnd.n5859 gnd.n5858 585
R166 gnd.n5856 gnd.n726 585
R167 gnd.n726 gnd.n725 585
R168 gnd.n5855 gnd.n5854 585
R169 gnd.n5854 gnd.n5853 585
R170 gnd.n732 gnd.n731 585
R171 gnd.n5852 gnd.n732 585
R172 gnd.n5850 gnd.n5849 585
R173 gnd.n5851 gnd.n5850 585
R174 gnd.n5848 gnd.n734 585
R175 gnd.n734 gnd.n733 585
R176 gnd.n5847 gnd.n5846 585
R177 gnd.n5846 gnd.n5845 585
R178 gnd.n740 gnd.n739 585
R179 gnd.n5844 gnd.n740 585
R180 gnd.n5842 gnd.n5841 585
R181 gnd.n5843 gnd.n5842 585
R182 gnd.n5840 gnd.n742 585
R183 gnd.n742 gnd.n741 585
R184 gnd.n5839 gnd.n5838 585
R185 gnd.n5838 gnd.n5837 585
R186 gnd.n748 gnd.n747 585
R187 gnd.n5836 gnd.n748 585
R188 gnd.n5834 gnd.n5833 585
R189 gnd.n5835 gnd.n5834 585
R190 gnd.n5832 gnd.n750 585
R191 gnd.n750 gnd.n749 585
R192 gnd.n5831 gnd.n5830 585
R193 gnd.n5830 gnd.n5829 585
R194 gnd.n756 gnd.n755 585
R195 gnd.n5828 gnd.n756 585
R196 gnd.n5826 gnd.n5825 585
R197 gnd.n5827 gnd.n5826 585
R198 gnd.n5824 gnd.n758 585
R199 gnd.n758 gnd.n757 585
R200 gnd.n5823 gnd.n5822 585
R201 gnd.n5822 gnd.n5821 585
R202 gnd.n5991 gnd.n5990 585
R203 gnd.n5990 gnd.n5989 585
R204 gnd.n594 gnd.n593 585
R205 gnd.n593 gnd.n592 585
R206 gnd.n5996 gnd.n5995 585
R207 gnd.n5997 gnd.n5996 585
R208 gnd.n591 gnd.n590 585
R209 gnd.n5998 gnd.n591 585
R210 gnd.n6001 gnd.n6000 585
R211 gnd.n6000 gnd.n5999 585
R212 gnd.n588 gnd.n587 585
R213 gnd.n587 gnd.n586 585
R214 gnd.n6006 gnd.n6005 585
R215 gnd.n6007 gnd.n6006 585
R216 gnd.n585 gnd.n584 585
R217 gnd.n6008 gnd.n585 585
R218 gnd.n6011 gnd.n6010 585
R219 gnd.n6010 gnd.n6009 585
R220 gnd.n582 gnd.n581 585
R221 gnd.n581 gnd.n580 585
R222 gnd.n6016 gnd.n6015 585
R223 gnd.n6017 gnd.n6016 585
R224 gnd.n579 gnd.n578 585
R225 gnd.n6018 gnd.n579 585
R226 gnd.n6021 gnd.n6020 585
R227 gnd.n6020 gnd.n6019 585
R228 gnd.n576 gnd.n575 585
R229 gnd.n575 gnd.n574 585
R230 gnd.n6026 gnd.n6025 585
R231 gnd.n6027 gnd.n6026 585
R232 gnd.n573 gnd.n572 585
R233 gnd.n6028 gnd.n573 585
R234 gnd.n6031 gnd.n6030 585
R235 gnd.n6030 gnd.n6029 585
R236 gnd.n570 gnd.n569 585
R237 gnd.n569 gnd.n568 585
R238 gnd.n6036 gnd.n6035 585
R239 gnd.n6037 gnd.n6036 585
R240 gnd.n567 gnd.n566 585
R241 gnd.n6038 gnd.n567 585
R242 gnd.n6041 gnd.n6040 585
R243 gnd.n6040 gnd.n6039 585
R244 gnd.n564 gnd.n563 585
R245 gnd.n563 gnd.n562 585
R246 gnd.n6046 gnd.n6045 585
R247 gnd.n6047 gnd.n6046 585
R248 gnd.n561 gnd.n560 585
R249 gnd.n6048 gnd.n561 585
R250 gnd.n6051 gnd.n6050 585
R251 gnd.n6050 gnd.n6049 585
R252 gnd.n558 gnd.n557 585
R253 gnd.n557 gnd.n556 585
R254 gnd.n6056 gnd.n6055 585
R255 gnd.n6057 gnd.n6056 585
R256 gnd.n555 gnd.n554 585
R257 gnd.n6058 gnd.n555 585
R258 gnd.n6061 gnd.n6060 585
R259 gnd.n6060 gnd.n6059 585
R260 gnd.n552 gnd.n551 585
R261 gnd.n551 gnd.n550 585
R262 gnd.n6066 gnd.n6065 585
R263 gnd.n6067 gnd.n6066 585
R264 gnd.n549 gnd.n548 585
R265 gnd.n6068 gnd.n549 585
R266 gnd.n6071 gnd.n6070 585
R267 gnd.n6070 gnd.n6069 585
R268 gnd.n546 gnd.n545 585
R269 gnd.n545 gnd.n544 585
R270 gnd.n6076 gnd.n6075 585
R271 gnd.n6077 gnd.n6076 585
R272 gnd.n543 gnd.n542 585
R273 gnd.n6078 gnd.n543 585
R274 gnd.n6081 gnd.n6080 585
R275 gnd.n6080 gnd.n6079 585
R276 gnd.n540 gnd.n539 585
R277 gnd.n539 gnd.n538 585
R278 gnd.n6086 gnd.n6085 585
R279 gnd.n6087 gnd.n6086 585
R280 gnd.n537 gnd.n536 585
R281 gnd.n6088 gnd.n537 585
R282 gnd.n6091 gnd.n6090 585
R283 gnd.n6090 gnd.n6089 585
R284 gnd.n534 gnd.n533 585
R285 gnd.n533 gnd.n532 585
R286 gnd.n6096 gnd.n6095 585
R287 gnd.n6097 gnd.n6096 585
R288 gnd.n531 gnd.n530 585
R289 gnd.n6098 gnd.n531 585
R290 gnd.n6101 gnd.n6100 585
R291 gnd.n6100 gnd.n6099 585
R292 gnd.n528 gnd.n527 585
R293 gnd.n527 gnd.n526 585
R294 gnd.n6106 gnd.n6105 585
R295 gnd.n6107 gnd.n6106 585
R296 gnd.n525 gnd.n524 585
R297 gnd.n6108 gnd.n525 585
R298 gnd.n6111 gnd.n6110 585
R299 gnd.n6110 gnd.n6109 585
R300 gnd.n522 gnd.n521 585
R301 gnd.n521 gnd.n520 585
R302 gnd.n6116 gnd.n6115 585
R303 gnd.n6117 gnd.n6116 585
R304 gnd.n519 gnd.n518 585
R305 gnd.n6118 gnd.n519 585
R306 gnd.n6121 gnd.n6120 585
R307 gnd.n6120 gnd.n6119 585
R308 gnd.n516 gnd.n515 585
R309 gnd.n515 gnd.n514 585
R310 gnd.n6126 gnd.n6125 585
R311 gnd.n6127 gnd.n6126 585
R312 gnd.n513 gnd.n512 585
R313 gnd.n6128 gnd.n513 585
R314 gnd.n6131 gnd.n6130 585
R315 gnd.n6130 gnd.n6129 585
R316 gnd.n510 gnd.n509 585
R317 gnd.n509 gnd.n508 585
R318 gnd.n6136 gnd.n6135 585
R319 gnd.n6137 gnd.n6136 585
R320 gnd.n507 gnd.n506 585
R321 gnd.n6138 gnd.n507 585
R322 gnd.n6141 gnd.n6140 585
R323 gnd.n6140 gnd.n6139 585
R324 gnd.n504 gnd.n503 585
R325 gnd.n503 gnd.n502 585
R326 gnd.n6146 gnd.n6145 585
R327 gnd.n6147 gnd.n6146 585
R328 gnd.n501 gnd.n500 585
R329 gnd.n6148 gnd.n501 585
R330 gnd.n6151 gnd.n6150 585
R331 gnd.n6150 gnd.n6149 585
R332 gnd.n498 gnd.n497 585
R333 gnd.n497 gnd.n496 585
R334 gnd.n6156 gnd.n6155 585
R335 gnd.n6157 gnd.n6156 585
R336 gnd.n495 gnd.n494 585
R337 gnd.n6158 gnd.n495 585
R338 gnd.n6161 gnd.n6160 585
R339 gnd.n6160 gnd.n6159 585
R340 gnd.n492 gnd.n491 585
R341 gnd.n491 gnd.n490 585
R342 gnd.n6166 gnd.n6165 585
R343 gnd.n6167 gnd.n6166 585
R344 gnd.n489 gnd.n488 585
R345 gnd.n6168 gnd.n489 585
R346 gnd.n6171 gnd.n6170 585
R347 gnd.n6170 gnd.n6169 585
R348 gnd.n486 gnd.n485 585
R349 gnd.n485 gnd.n484 585
R350 gnd.n6176 gnd.n6175 585
R351 gnd.n6177 gnd.n6176 585
R352 gnd.n483 gnd.n482 585
R353 gnd.n6178 gnd.n483 585
R354 gnd.n6181 gnd.n6180 585
R355 gnd.n6180 gnd.n6179 585
R356 gnd.n480 gnd.n479 585
R357 gnd.n479 gnd.n478 585
R358 gnd.n6186 gnd.n6185 585
R359 gnd.n6187 gnd.n6186 585
R360 gnd.n477 gnd.n476 585
R361 gnd.n6188 gnd.n477 585
R362 gnd.n6191 gnd.n6190 585
R363 gnd.n6190 gnd.n6189 585
R364 gnd.n474 gnd.n473 585
R365 gnd.n473 gnd.n472 585
R366 gnd.n6196 gnd.n6195 585
R367 gnd.n6197 gnd.n6196 585
R368 gnd.n471 gnd.n470 585
R369 gnd.n6198 gnd.n471 585
R370 gnd.n6201 gnd.n6200 585
R371 gnd.n6200 gnd.n6199 585
R372 gnd.n468 gnd.n467 585
R373 gnd.n467 gnd.n466 585
R374 gnd.n6206 gnd.n6205 585
R375 gnd.n6207 gnd.n6206 585
R376 gnd.n465 gnd.n464 585
R377 gnd.n6208 gnd.n465 585
R378 gnd.n6211 gnd.n6210 585
R379 gnd.n6210 gnd.n6209 585
R380 gnd.n462 gnd.n461 585
R381 gnd.n461 gnd.n460 585
R382 gnd.n6216 gnd.n6215 585
R383 gnd.n6217 gnd.n6216 585
R384 gnd.n459 gnd.n458 585
R385 gnd.n6218 gnd.n459 585
R386 gnd.n6221 gnd.n6220 585
R387 gnd.n6220 gnd.n6219 585
R388 gnd.n456 gnd.n455 585
R389 gnd.n455 gnd.n454 585
R390 gnd.n6226 gnd.n6225 585
R391 gnd.n6227 gnd.n6226 585
R392 gnd.n453 gnd.n452 585
R393 gnd.n6228 gnd.n453 585
R394 gnd.n6231 gnd.n6230 585
R395 gnd.n6230 gnd.n6229 585
R396 gnd.n450 gnd.n449 585
R397 gnd.n449 gnd.n448 585
R398 gnd.n6236 gnd.n6235 585
R399 gnd.n6237 gnd.n6236 585
R400 gnd.n447 gnd.n446 585
R401 gnd.n6238 gnd.n447 585
R402 gnd.n6241 gnd.n6240 585
R403 gnd.n6240 gnd.n6239 585
R404 gnd.n444 gnd.n443 585
R405 gnd.n443 gnd.n442 585
R406 gnd.n6246 gnd.n6245 585
R407 gnd.n6247 gnd.n6246 585
R408 gnd.n441 gnd.n440 585
R409 gnd.n6248 gnd.n441 585
R410 gnd.n6251 gnd.n6250 585
R411 gnd.n6250 gnd.n6249 585
R412 gnd.n438 gnd.n437 585
R413 gnd.n437 gnd.n436 585
R414 gnd.n6256 gnd.n6255 585
R415 gnd.n6257 gnd.n6256 585
R416 gnd.n435 gnd.n434 585
R417 gnd.n6258 gnd.n435 585
R418 gnd.n6261 gnd.n6260 585
R419 gnd.n6260 gnd.n6259 585
R420 gnd.n432 gnd.n431 585
R421 gnd.n431 gnd.n430 585
R422 gnd.n6266 gnd.n6265 585
R423 gnd.n6267 gnd.n6266 585
R424 gnd.n429 gnd.n428 585
R425 gnd.n6268 gnd.n429 585
R426 gnd.n6271 gnd.n6270 585
R427 gnd.n6270 gnd.n6269 585
R428 gnd.n426 gnd.n425 585
R429 gnd.n425 gnd.n424 585
R430 gnd.n6276 gnd.n6275 585
R431 gnd.n6277 gnd.n6276 585
R432 gnd.n423 gnd.n422 585
R433 gnd.n6278 gnd.n423 585
R434 gnd.n6281 gnd.n6280 585
R435 gnd.n6280 gnd.n6279 585
R436 gnd.n420 gnd.n419 585
R437 gnd.n419 gnd.n418 585
R438 gnd.n6286 gnd.n6285 585
R439 gnd.n6287 gnd.n6286 585
R440 gnd.n417 gnd.n416 585
R441 gnd.n6288 gnd.n417 585
R442 gnd.n6291 gnd.n6290 585
R443 gnd.n6290 gnd.n6289 585
R444 gnd.n414 gnd.n413 585
R445 gnd.n413 gnd.n412 585
R446 gnd.n6296 gnd.n6295 585
R447 gnd.n6297 gnd.n6296 585
R448 gnd.n411 gnd.n410 585
R449 gnd.n6298 gnd.n411 585
R450 gnd.n6301 gnd.n6300 585
R451 gnd.n6300 gnd.n6299 585
R452 gnd.n408 gnd.n407 585
R453 gnd.n407 gnd.n406 585
R454 gnd.n6306 gnd.n6305 585
R455 gnd.n6307 gnd.n6306 585
R456 gnd.n405 gnd.n404 585
R457 gnd.n6308 gnd.n405 585
R458 gnd.n6311 gnd.n6310 585
R459 gnd.n6310 gnd.n6309 585
R460 gnd.n402 gnd.n401 585
R461 gnd.n401 gnd.n400 585
R462 gnd.n6316 gnd.n6315 585
R463 gnd.n6317 gnd.n6316 585
R464 gnd.n399 gnd.n398 585
R465 gnd.n6318 gnd.n399 585
R466 gnd.n6321 gnd.n6320 585
R467 gnd.n6320 gnd.n6319 585
R468 gnd.n396 gnd.n395 585
R469 gnd.n395 gnd.n394 585
R470 gnd.n6326 gnd.n6325 585
R471 gnd.n6327 gnd.n6326 585
R472 gnd.n393 gnd.n392 585
R473 gnd.n6328 gnd.n393 585
R474 gnd.n6331 gnd.n6330 585
R475 gnd.n6330 gnd.n6329 585
R476 gnd.n390 gnd.n389 585
R477 gnd.n389 gnd.n388 585
R478 gnd.n6337 gnd.n6336 585
R479 gnd.n6338 gnd.n6337 585
R480 gnd.n387 gnd.n386 585
R481 gnd.n6339 gnd.n387 585
R482 gnd.n6342 gnd.n6341 585
R483 gnd.n6341 gnd.n6340 585
R484 gnd.n6343 gnd.n384 585
R485 gnd.n384 gnd.n383 585
R486 gnd.n259 gnd.n258 585
R487 gnd.n6550 gnd.n258 585
R488 gnd.n6553 gnd.n6552 585
R489 gnd.n6552 gnd.n6551 585
R490 gnd.n262 gnd.n261 585
R491 gnd.n6549 gnd.n262 585
R492 gnd.n6547 gnd.n6546 585
R493 gnd.n6548 gnd.n6547 585
R494 gnd.n265 gnd.n264 585
R495 gnd.n264 gnd.n263 585
R496 gnd.n6542 gnd.n6541 585
R497 gnd.n6541 gnd.n6540 585
R498 gnd.n268 gnd.n267 585
R499 gnd.n6539 gnd.n268 585
R500 gnd.n6537 gnd.n6536 585
R501 gnd.n6538 gnd.n6537 585
R502 gnd.n271 gnd.n270 585
R503 gnd.n270 gnd.n269 585
R504 gnd.n6532 gnd.n6531 585
R505 gnd.n6531 gnd.n6530 585
R506 gnd.n274 gnd.n273 585
R507 gnd.n6529 gnd.n274 585
R508 gnd.n6527 gnd.n6526 585
R509 gnd.n6528 gnd.n6527 585
R510 gnd.n277 gnd.n276 585
R511 gnd.n276 gnd.n275 585
R512 gnd.n6522 gnd.n6521 585
R513 gnd.n6521 gnd.n6520 585
R514 gnd.n280 gnd.n279 585
R515 gnd.n6519 gnd.n280 585
R516 gnd.n6517 gnd.n6516 585
R517 gnd.n6518 gnd.n6517 585
R518 gnd.n283 gnd.n282 585
R519 gnd.n282 gnd.n281 585
R520 gnd.n6512 gnd.n6511 585
R521 gnd.n6511 gnd.n6510 585
R522 gnd.n286 gnd.n285 585
R523 gnd.n6509 gnd.n286 585
R524 gnd.n6507 gnd.n6506 585
R525 gnd.n6508 gnd.n6507 585
R526 gnd.n289 gnd.n288 585
R527 gnd.n288 gnd.n287 585
R528 gnd.n6502 gnd.n6501 585
R529 gnd.n6501 gnd.n6500 585
R530 gnd.n292 gnd.n291 585
R531 gnd.n6499 gnd.n292 585
R532 gnd.n6497 gnd.n6496 585
R533 gnd.n6498 gnd.n6497 585
R534 gnd.n295 gnd.n294 585
R535 gnd.n294 gnd.n293 585
R536 gnd.n6492 gnd.n6491 585
R537 gnd.n6491 gnd.n6490 585
R538 gnd.n298 gnd.n297 585
R539 gnd.n6489 gnd.n298 585
R540 gnd.n6487 gnd.n6486 585
R541 gnd.n6488 gnd.n6487 585
R542 gnd.n301 gnd.n300 585
R543 gnd.n300 gnd.n299 585
R544 gnd.n6482 gnd.n6481 585
R545 gnd.n6481 gnd.n6480 585
R546 gnd.n304 gnd.n303 585
R547 gnd.n6479 gnd.n304 585
R548 gnd.n6477 gnd.n6476 585
R549 gnd.n6478 gnd.n6477 585
R550 gnd.n307 gnd.n306 585
R551 gnd.n306 gnd.n305 585
R552 gnd.n6472 gnd.n6471 585
R553 gnd.n6471 gnd.n6470 585
R554 gnd.n310 gnd.n309 585
R555 gnd.n6469 gnd.n310 585
R556 gnd.n6467 gnd.n6466 585
R557 gnd.n6468 gnd.n6467 585
R558 gnd.n313 gnd.n312 585
R559 gnd.n312 gnd.n311 585
R560 gnd.n6462 gnd.n6461 585
R561 gnd.n6461 gnd.n6460 585
R562 gnd.n316 gnd.n315 585
R563 gnd.n6459 gnd.n316 585
R564 gnd.n6457 gnd.n6456 585
R565 gnd.n6458 gnd.n6457 585
R566 gnd.n319 gnd.n318 585
R567 gnd.n318 gnd.n317 585
R568 gnd.n6452 gnd.n6451 585
R569 gnd.n6451 gnd.n6450 585
R570 gnd.n322 gnd.n321 585
R571 gnd.n6449 gnd.n322 585
R572 gnd.n6447 gnd.n6446 585
R573 gnd.n6448 gnd.n6447 585
R574 gnd.n325 gnd.n324 585
R575 gnd.n324 gnd.n323 585
R576 gnd.n6442 gnd.n6441 585
R577 gnd.n6441 gnd.n6440 585
R578 gnd.n328 gnd.n327 585
R579 gnd.n6439 gnd.n328 585
R580 gnd.n6437 gnd.n6436 585
R581 gnd.n6438 gnd.n6437 585
R582 gnd.n331 gnd.n330 585
R583 gnd.n330 gnd.n329 585
R584 gnd.n6432 gnd.n6431 585
R585 gnd.n6431 gnd.n6430 585
R586 gnd.n334 gnd.n333 585
R587 gnd.n6429 gnd.n334 585
R588 gnd.n6427 gnd.n6426 585
R589 gnd.n6428 gnd.n6427 585
R590 gnd.n337 gnd.n336 585
R591 gnd.n336 gnd.n335 585
R592 gnd.n6422 gnd.n6421 585
R593 gnd.n6421 gnd.n6420 585
R594 gnd.n340 gnd.n339 585
R595 gnd.n6419 gnd.n340 585
R596 gnd.n6417 gnd.n6416 585
R597 gnd.n6418 gnd.n6417 585
R598 gnd.n343 gnd.n342 585
R599 gnd.n342 gnd.n341 585
R600 gnd.n6412 gnd.n6411 585
R601 gnd.n6411 gnd.n6410 585
R602 gnd.n346 gnd.n345 585
R603 gnd.n6409 gnd.n346 585
R604 gnd.n6407 gnd.n6406 585
R605 gnd.n6408 gnd.n6407 585
R606 gnd.n349 gnd.n348 585
R607 gnd.n348 gnd.n347 585
R608 gnd.n6402 gnd.n6401 585
R609 gnd.n6401 gnd.n6400 585
R610 gnd.n352 gnd.n351 585
R611 gnd.n6399 gnd.n352 585
R612 gnd.n6397 gnd.n6396 585
R613 gnd.n6398 gnd.n6397 585
R614 gnd.n355 gnd.n354 585
R615 gnd.n354 gnd.n353 585
R616 gnd.n6392 gnd.n6391 585
R617 gnd.n6391 gnd.n6390 585
R618 gnd.n358 gnd.n357 585
R619 gnd.n6389 gnd.n358 585
R620 gnd.n6387 gnd.n6386 585
R621 gnd.n6388 gnd.n6387 585
R622 gnd.n361 gnd.n360 585
R623 gnd.n360 gnd.n359 585
R624 gnd.n6382 gnd.n6381 585
R625 gnd.n6381 gnd.n6380 585
R626 gnd.n364 gnd.n363 585
R627 gnd.n6379 gnd.n364 585
R628 gnd.n6377 gnd.n6376 585
R629 gnd.n6378 gnd.n6377 585
R630 gnd.n367 gnd.n366 585
R631 gnd.n366 gnd.n365 585
R632 gnd.n6372 gnd.n6371 585
R633 gnd.n6371 gnd.n6370 585
R634 gnd.n370 gnd.n369 585
R635 gnd.n6369 gnd.n370 585
R636 gnd.n6367 gnd.n6366 585
R637 gnd.n6368 gnd.n6367 585
R638 gnd.n373 gnd.n372 585
R639 gnd.n372 gnd.n371 585
R640 gnd.n6362 gnd.n6361 585
R641 gnd.n6361 gnd.n6360 585
R642 gnd.n376 gnd.n375 585
R643 gnd.n6359 gnd.n376 585
R644 gnd.n6357 gnd.n6356 585
R645 gnd.n6358 gnd.n6357 585
R646 gnd.n379 gnd.n378 585
R647 gnd.n378 gnd.n377 585
R648 gnd.n6352 gnd.n6351 585
R649 gnd.n6351 gnd.n6350 585
R650 gnd.n382 gnd.n381 585
R651 gnd.n6349 gnd.n382 585
R652 gnd.n6347 gnd.n6346 585
R653 gnd.n6348 gnd.n6347 585
R654 gnd.n4200 gnd.n4199 585
R655 gnd.n4201 gnd.n4200 585
R656 gnd.n1068 gnd.n1067 585
R657 gnd.n2418 gnd.n1068 585
R658 gnd.n4209 gnd.n4208 585
R659 gnd.n4208 gnd.n4207 585
R660 gnd.n4210 gnd.n1062 585
R661 gnd.n2378 gnd.n1062 585
R662 gnd.n4212 gnd.n4211 585
R663 gnd.n4213 gnd.n4212 585
R664 gnd.n1047 gnd.n1046 585
R665 gnd.n2369 gnd.n1047 585
R666 gnd.n4221 gnd.n4220 585
R667 gnd.n4220 gnd.n4219 585
R668 gnd.n4222 gnd.n1041 585
R669 gnd.n2361 gnd.n1041 585
R670 gnd.n4224 gnd.n4223 585
R671 gnd.n4225 gnd.n4224 585
R672 gnd.n1025 gnd.n1024 585
R673 gnd.n2286 gnd.n1025 585
R674 gnd.n4233 gnd.n4232 585
R675 gnd.n4232 gnd.n4231 585
R676 gnd.n4234 gnd.n1019 585
R677 gnd.n2274 gnd.n1019 585
R678 gnd.n4236 gnd.n4235 585
R679 gnd.n4237 gnd.n4236 585
R680 gnd.n1005 gnd.n1004 585
R681 gnd.n2269 gnd.n1005 585
R682 gnd.n4245 gnd.n4244 585
R683 gnd.n4244 gnd.n4243 585
R684 gnd.n4246 gnd.n999 585
R685 gnd.n2300 gnd.n999 585
R686 gnd.n4248 gnd.n4247 585
R687 gnd.n4249 gnd.n4248 585
R688 gnd.n986 gnd.n985 585
R689 gnd.n2261 gnd.n986 585
R690 gnd.n4258 gnd.n4257 585
R691 gnd.n4257 gnd.n4256 585
R692 gnd.n4259 gnd.n981 585
R693 gnd.n2253 gnd.n981 585
R694 gnd.n4261 gnd.n4260 585
R695 gnd.n4262 gnd.n4261 585
R696 gnd.n970 gnd.n969 585
R697 gnd.n2244 gnd.n970 585
R698 gnd.n4271 gnd.n4270 585
R699 gnd.n4270 gnd.n4269 585
R700 gnd.n4272 gnd.n962 585
R701 gnd.n962 gnd.n960 585
R702 gnd.n4274 gnd.n4273 585
R703 gnd.n4275 gnd.n4274 585
R704 gnd.n963 gnd.n961 585
R705 gnd.n2233 gnd.n961 585
R706 gnd.n946 gnd.n945 585
R707 gnd.n949 gnd.n946 585
R708 gnd.n4285 gnd.n4284 585
R709 gnd.n4284 gnd.n4283 585
R710 gnd.n4286 gnd.n940 585
R711 gnd.n940 gnd.n939 585
R712 gnd.n4288 gnd.n4287 585
R713 gnd.n4289 gnd.n4288 585
R714 gnd.n925 gnd.n924 585
R715 gnd.n936 gnd.n925 585
R716 gnd.n4297 gnd.n4296 585
R717 gnd.n4296 gnd.n4295 585
R718 gnd.n4298 gnd.n919 585
R719 gnd.n926 gnd.n919 585
R720 gnd.n4300 gnd.n4299 585
R721 gnd.n4301 gnd.n4300 585
R722 gnd.n906 gnd.n905 585
R723 gnd.n909 gnd.n906 585
R724 gnd.n4309 gnd.n4308 585
R725 gnd.n4308 gnd.n4307 585
R726 gnd.n4310 gnd.n900 585
R727 gnd.n900 gnd.n898 585
R728 gnd.n4312 gnd.n4311 585
R729 gnd.n4313 gnd.n4312 585
R730 gnd.n901 gnd.n899 585
R731 gnd.n899 gnd.n886 585
R732 gnd.n2153 gnd.n887 585
R733 gnd.n4319 gnd.n887 585
R734 gnd.n2089 gnd.n2087 585
R735 gnd.n2087 gnd.n884 585
R736 gnd.n2158 gnd.n2157 585
R737 gnd.n2165 gnd.n2158 585
R738 gnd.n2088 gnd.n2086 585
R739 gnd.n2086 gnd.n830 585
R740 gnd.n2149 gnd.n2148 585
R741 gnd.n2147 gnd.n2146 585
R742 gnd.n2145 gnd.n2144 585
R743 gnd.n2143 gnd.n2142 585
R744 gnd.n2141 gnd.n2140 585
R745 gnd.n2139 gnd.n2138 585
R746 gnd.n2137 gnd.n2136 585
R747 gnd.n2135 gnd.n2134 585
R748 gnd.n2133 gnd.n2132 585
R749 gnd.n2131 gnd.n2130 585
R750 gnd.n2129 gnd.n2128 585
R751 gnd.n2127 gnd.n2126 585
R752 gnd.n2125 gnd.n2124 585
R753 gnd.n2123 gnd.n2122 585
R754 gnd.n2121 gnd.n2120 585
R755 gnd.n2119 gnd.n2118 585
R756 gnd.n2117 gnd.n2116 585
R757 gnd.n2108 gnd.n2105 585
R758 gnd.n2112 gnd.n829 585
R759 gnd.n4406 gnd.n829 585
R760 gnd.n2628 gnd.n2627 585
R761 gnd.n1917 gnd.n1909 585
R762 gnd.n2635 gnd.n1906 585
R763 gnd.n2636 gnd.n1905 585
R764 gnd.n1931 gnd.n1899 585
R765 gnd.n2643 gnd.n1898 585
R766 gnd.n2644 gnd.n1897 585
R767 gnd.n1929 gnd.n1889 585
R768 gnd.n2651 gnd.n1888 585
R769 gnd.n2652 gnd.n1887 585
R770 gnd.n1926 gnd.n1881 585
R771 gnd.n2659 gnd.n1880 585
R772 gnd.n2660 gnd.n1879 585
R773 gnd.n1924 gnd.n1872 585
R774 gnd.n2667 gnd.n1871 585
R775 gnd.n2668 gnd.n1870 585
R776 gnd.n1921 gnd.n1869 585
R777 gnd.n1920 gnd.n1919 585
R778 gnd.n1085 gnd.n1083 585
R779 gnd.n2625 gnd.n1083 585
R780 gnd.n2001 gnd.n1081 585
R781 gnd.n4201 gnd.n1081 585
R782 gnd.n2417 gnd.n2416 585
R783 gnd.n2418 gnd.n2417 585
R784 gnd.n2000 gnd.n1071 585
R785 gnd.n4207 gnd.n1071 585
R786 gnd.n2380 gnd.n2379 585
R787 gnd.n2379 gnd.n2378 585
R788 gnd.n2003 gnd.n1060 585
R789 gnd.n4213 gnd.n1060 585
R790 gnd.n2368 gnd.n2367 585
R791 gnd.n2369 gnd.n2368 585
R792 gnd.n2007 gnd.n1049 585
R793 gnd.n4219 gnd.n1049 585
R794 gnd.n2363 gnd.n2362 585
R795 gnd.n2362 gnd.n2361 585
R796 gnd.n2009 gnd.n1039 585
R797 gnd.n4225 gnd.n1039 585
R798 gnd.n2288 gnd.n2287 585
R799 gnd.n2287 gnd.n2286 585
R800 gnd.n2029 gnd.n1028 585
R801 gnd.n4231 gnd.n1028 585
R802 gnd.n2292 gnd.n2028 585
R803 gnd.n2274 gnd.n2028 585
R804 gnd.n2293 gnd.n1018 585
R805 gnd.n4237 gnd.n1018 585
R806 gnd.n2294 gnd.n2027 585
R807 gnd.n2269 gnd.n2027 585
R808 gnd.n2024 gnd.n1007 585
R809 gnd.n4243 gnd.n1007 585
R810 gnd.n2299 gnd.n2298 585
R811 gnd.n2300 gnd.n2299 585
R812 gnd.n2023 gnd.n997 585
R813 gnd.n4249 gnd.n997 585
R814 gnd.n2260 gnd.n2259 585
R815 gnd.n2261 gnd.n2260 585
R816 gnd.n2036 gnd.n989 585
R817 gnd.n4256 gnd.n989 585
R818 gnd.n2255 gnd.n2254 585
R819 gnd.n2254 gnd.n2253 585
R820 gnd.n2038 gnd.n980 585
R821 gnd.n4262 gnd.n980 585
R822 gnd.n2243 gnd.n2242 585
R823 gnd.n2244 gnd.n2243 585
R824 gnd.n2071 gnd.n972 585
R825 gnd.n4269 gnd.n972 585
R826 gnd.n2238 gnd.n2237 585
R827 gnd.n2237 gnd.n960 585
R828 gnd.n2236 gnd.n959 585
R829 gnd.n4275 gnd.n959 585
R830 gnd.n2235 gnd.n2234 585
R831 gnd.n2234 gnd.n2233 585
R832 gnd.n2194 gnd.n2073 585
R833 gnd.n2194 gnd.n949 585
R834 gnd.n2190 gnd.n948 585
R835 gnd.n4283 gnd.n948 585
R836 gnd.n2189 gnd.n2188 585
R837 gnd.n2188 gnd.n939 585
R838 gnd.n2187 gnd.n938 585
R839 gnd.n4289 gnd.n938 585
R840 gnd.n2076 gnd.n2075 585
R841 gnd.n2075 gnd.n936 585
R842 gnd.n2183 gnd.n928 585
R843 gnd.n4295 gnd.n928 585
R844 gnd.n2182 gnd.n2181 585
R845 gnd.n2181 gnd.n926 585
R846 gnd.n2180 gnd.n918 585
R847 gnd.n4301 gnd.n918 585
R848 gnd.n2079 gnd.n2078 585
R849 gnd.n2078 gnd.n909 585
R850 gnd.n2176 gnd.n908 585
R851 gnd.n4307 gnd.n908 585
R852 gnd.n2175 gnd.n2174 585
R853 gnd.n2174 gnd.n898 585
R854 gnd.n2173 gnd.n897 585
R855 gnd.n4313 gnd.n897 585
R856 gnd.n2082 gnd.n2081 585
R857 gnd.n2081 gnd.n886 585
R858 gnd.n2169 gnd.n885 585
R859 gnd.n4319 gnd.n885 585
R860 gnd.n2168 gnd.n2167 585
R861 gnd.n2167 gnd.n884 585
R862 gnd.n2166 gnd.n2084 585
R863 gnd.n2166 gnd.n2165 585
R864 gnd.n2110 gnd.n2085 585
R865 gnd.n2085 gnd.n830 585
R866 gnd.n6709 gnd.n84 585
R867 gnd.n6805 gnd.n84 585
R868 gnd.n6710 gnd.n6641 585
R869 gnd.n6641 gnd.n81 585
R870 gnd.n6711 gnd.n163 585
R871 gnd.n6725 gnd.n163 585
R872 gnd.n175 gnd.n173 585
R873 gnd.n173 gnd.n161 585
R874 gnd.n6716 gnd.n6715 585
R875 gnd.n6717 gnd.n6716 585
R876 gnd.n174 gnd.n172 585
R877 gnd.n172 gnd.n170 585
R878 gnd.n6637 gnd.n6636 585
R879 gnd.n6636 gnd.n6635 585
R880 gnd.n178 gnd.n177 585
R881 gnd.n188 gnd.n178 585
R882 gnd.n6626 gnd.n6625 585
R883 gnd.n6627 gnd.n6626 585
R884 gnd.n190 gnd.n189 585
R885 gnd.n189 gnd.n186 585
R886 gnd.n6621 gnd.n6620 585
R887 gnd.n6620 gnd.n6619 585
R888 gnd.n193 gnd.n192 585
R889 gnd.n194 gnd.n193 585
R890 gnd.n6610 gnd.n6609 585
R891 gnd.n6611 gnd.n6610 585
R892 gnd.n205 gnd.n204 585
R893 gnd.n204 gnd.n202 585
R894 gnd.n6605 gnd.n6604 585
R895 gnd.n6604 gnd.n6603 585
R896 gnd.n208 gnd.n207 585
R897 gnd.n224 gnd.n208 585
R898 gnd.n6594 gnd.n6593 585
R899 gnd.n6595 gnd.n6594 585
R900 gnd.n226 gnd.n225 585
R901 gnd.n225 gnd.n222 585
R902 gnd.n6589 gnd.n6588 585
R903 gnd.n6588 gnd.n6587 585
R904 gnd.n229 gnd.n228 585
R905 gnd.n230 gnd.n229 585
R906 gnd.n6580 gnd.n6579 585
R907 gnd.n6581 gnd.n6580 585
R908 gnd.n239 gnd.n238 585
R909 gnd.n3890 gnd.n238 585
R910 gnd.n6575 gnd.n6574 585
R911 gnd.n6574 gnd.n6573 585
R912 gnd.n243 gnd.n242 585
R913 gnd.n6568 gnd.n243 585
R914 gnd.n4022 gnd.n4020 585
R915 gnd.n4020 gnd.n4019 585
R916 gnd.n4023 gnd.n1250 585
R917 gnd.n3896 gnd.n1250 585
R918 gnd.n4024 gnd.n1249 585
R919 gnd.n4010 gnd.n1249 585
R920 gnd.n1273 gnd.n1247 585
R921 gnd.n1274 gnd.n1273 585
R922 gnd.n4028 gnd.n1246 585
R923 gnd.n4004 gnd.n1246 585
R924 gnd.n4029 gnd.n1245 585
R925 gnd.n3985 gnd.n1245 585
R926 gnd.n4030 gnd.n1244 585
R927 gnd.n1281 gnd.n1244 585
R928 gnd.n1292 gnd.n1242 585
R929 gnd.n3976 gnd.n1292 585
R930 gnd.n4034 gnd.n1241 585
R931 gnd.n1302 gnd.n1241 585
R932 gnd.n4035 gnd.n1240 585
R933 gnd.n3965 gnd.n1240 585
R934 gnd.n4036 gnd.n1239 585
R935 gnd.n3953 gnd.n1239 585
R936 gnd.n1309 gnd.n1237 585
R937 gnd.n1310 gnd.n1309 585
R938 gnd.n4040 gnd.n1236 585
R939 gnd.n3944 gnd.n1236 585
R940 gnd.n4041 gnd.n1235 585
R941 gnd.n3916 gnd.n1235 585
R942 gnd.n4042 gnd.n1234 585
R943 gnd.n3934 gnd.n1234 585
R944 gnd.n1231 gnd.n1229 585
R945 gnd.n3823 gnd.n1229 585
R946 gnd.n4047 gnd.n4046 585
R947 gnd.n4048 gnd.n4047 585
R948 gnd.n1230 gnd.n1228 585
R949 gnd.n3814 gnd.n1228 585
R950 gnd.n3367 gnd.n1216 585
R951 gnd.n4054 gnd.n1216 585
R952 gnd.n3371 gnd.n3370 585
R953 gnd.n3373 gnd.n3364 585
R954 gnd.n3376 gnd.n3375 585
R955 gnd.n3357 gnd.n3356 585
R956 gnd.n3390 gnd.n3389 585
R957 gnd.n3392 gnd.n3355 585
R958 gnd.n3395 gnd.n3394 585
R959 gnd.n3348 gnd.n3347 585
R960 gnd.n3409 gnd.n3408 585
R961 gnd.n3411 gnd.n3346 585
R962 gnd.n3414 gnd.n3413 585
R963 gnd.n3339 gnd.n3338 585
R964 gnd.n3428 gnd.n3427 585
R965 gnd.n3430 gnd.n3337 585
R966 gnd.n3433 gnd.n3432 585
R967 gnd.n3330 gnd.n3329 585
R968 gnd.n3449 gnd.n3448 585
R969 gnd.n3451 gnd.n3328 585
R970 gnd.n3453 gnd.n3452 585
R971 gnd.n3452 gnd.n1204 585
R972 gnd.n6680 gnd.n80 585
R973 gnd.n6681 gnd.n6679 585
R974 gnd.n6682 gnd.n6675 585
R975 gnd.n6673 gnd.n6671 585
R976 gnd.n6686 gnd.n6670 585
R977 gnd.n6687 gnd.n6668 585
R978 gnd.n6688 gnd.n6667 585
R979 gnd.n6665 gnd.n6663 585
R980 gnd.n6692 gnd.n6662 585
R981 gnd.n6693 gnd.n6660 585
R982 gnd.n6694 gnd.n6659 585
R983 gnd.n6657 gnd.n6655 585
R984 gnd.n6698 gnd.n6654 585
R985 gnd.n6699 gnd.n6652 585
R986 gnd.n6700 gnd.n6651 585
R987 gnd.n6649 gnd.n6647 585
R988 gnd.n6704 gnd.n6646 585
R989 gnd.n6705 gnd.n6644 585
R990 gnd.n6706 gnd.n6643 585
R991 gnd.n6643 gnd.n83 585
R992 gnd.n6807 gnd.n6806 585
R993 gnd.n6806 gnd.n6805 585
R994 gnd.n79 gnd.n77 585
R995 gnd.n81 gnd.n79 585
R996 gnd.n6811 gnd.n76 585
R997 gnd.n6725 gnd.n76 585
R998 gnd.n6812 gnd.n75 585
R999 gnd.n161 gnd.n75 585
R1000 gnd.n6813 gnd.n74 585
R1001 gnd.n6717 gnd.n74 585
R1002 gnd.n169 gnd.n72 585
R1003 gnd.n170 gnd.n169 585
R1004 gnd.n6817 gnd.n71 585
R1005 gnd.n6635 gnd.n71 585
R1006 gnd.n6818 gnd.n70 585
R1007 gnd.n188 gnd.n70 585
R1008 gnd.n6819 gnd.n69 585
R1009 gnd.n6627 gnd.n69 585
R1010 gnd.n185 gnd.n67 585
R1011 gnd.n186 gnd.n185 585
R1012 gnd.n6823 gnd.n66 585
R1013 gnd.n6619 gnd.n66 585
R1014 gnd.n6824 gnd.n65 585
R1015 gnd.n194 gnd.n65 585
R1016 gnd.n6825 gnd.n64 585
R1017 gnd.n6611 gnd.n64 585
R1018 gnd.n201 gnd.n62 585
R1019 gnd.n202 gnd.n201 585
R1020 gnd.n6829 gnd.n61 585
R1021 gnd.n6603 gnd.n61 585
R1022 gnd.n6830 gnd.n60 585
R1023 gnd.n224 gnd.n60 585
R1024 gnd.n6831 gnd.n59 585
R1025 gnd.n6595 gnd.n59 585
R1026 gnd.n221 gnd.n57 585
R1027 gnd.n222 gnd.n221 585
R1028 gnd.n6835 gnd.n56 585
R1029 gnd.n6587 gnd.n56 585
R1030 gnd.n6836 gnd.n55 585
R1031 gnd.n230 gnd.n55 585
R1032 gnd.n6837 gnd.n54 585
R1033 gnd.n6581 gnd.n54 585
R1034 gnd.n3889 gnd.n52 585
R1035 gnd.n3890 gnd.n3889 585
R1036 gnd.n1255 gnd.n245 585
R1037 gnd.n6573 gnd.n245 585
R1038 gnd.n1256 gnd.n250 585
R1039 gnd.n6568 gnd.n250 585
R1040 gnd.n4018 gnd.n4017 585
R1041 gnd.n4019 gnd.n4018 585
R1042 gnd.n1254 gnd.n1253 585
R1043 gnd.n3896 gnd.n1253 585
R1044 gnd.n4012 gnd.n4011 585
R1045 gnd.n4011 gnd.n4010 585
R1046 gnd.n1259 gnd.n1258 585
R1047 gnd.n1274 gnd.n1259 585
R1048 gnd.n1285 gnd.n1272 585
R1049 gnd.n4004 gnd.n1272 585
R1050 gnd.n3984 gnd.n3983 585
R1051 gnd.n3985 gnd.n3984 585
R1052 gnd.n1284 gnd.n1283 585
R1053 gnd.n1283 gnd.n1281 585
R1054 gnd.n3978 gnd.n3977 585
R1055 gnd.n3977 gnd.n3976 585
R1056 gnd.n1288 gnd.n1287 585
R1057 gnd.n1302 gnd.n1288 585
R1058 gnd.n1314 gnd.n1301 585
R1059 gnd.n3965 gnd.n1301 585
R1060 gnd.n3952 gnd.n3951 585
R1061 gnd.n3953 gnd.n3952 585
R1062 gnd.n1313 gnd.n1312 585
R1063 gnd.n1312 gnd.n1310 585
R1064 gnd.n3946 gnd.n3945 585
R1065 gnd.n3945 gnd.n3944 585
R1066 gnd.n1317 gnd.n1316 585
R1067 gnd.n3916 gnd.n1317 585
R1068 gnd.n1332 gnd.n1327 585
R1069 gnd.n3934 gnd.n1327 585
R1070 gnd.n3822 gnd.n3821 585
R1071 gnd.n3823 gnd.n3822 585
R1072 gnd.n1331 gnd.n1226 585
R1073 gnd.n4048 gnd.n1226 585
R1074 gnd.n3816 gnd.n3815 585
R1075 gnd.n3815 gnd.n3814 585
R1076 gnd.n1334 gnd.n1214 585
R1077 gnd.n4054 gnd.n1214 585
R1078 gnd.n5801 gnd.n5800 585
R1079 gnd.n5800 gnd.n5799 585
R1080 gnd.n5802 gnd.n793 585
R1081 gnd.n5709 gnd.n793 585
R1082 gnd.n5804 gnd.n5803 585
R1083 gnd.n5805 gnd.n5804 585
R1084 gnd.n794 gnd.n792 585
R1085 gnd.n792 gnd.n788 585
R1086 gnd.n775 gnd.n774 585
R1087 gnd.n779 gnd.n775 585
R1088 gnd.n5815 gnd.n5814 585
R1089 gnd.n5814 gnd.n5813 585
R1090 gnd.n5816 gnd.n769 585
R1091 gnd.n5698 gnd.n769 585
R1092 gnd.n5818 gnd.n5817 585
R1093 gnd.n5819 gnd.n5818 585
R1094 gnd.n770 gnd.n768 585
R1095 gnd.n5692 gnd.n768 585
R1096 gnd.n5673 gnd.n4510 585
R1097 gnd.n4510 gnd.n4509 585
R1098 gnd.n5675 gnd.n5674 585
R1099 gnd.n5676 gnd.n5675 585
R1100 gnd.n4511 gnd.n4508 585
R1101 gnd.n4508 gnd.n4504 585
R1102 gnd.n5380 gnd.n5379 585
R1103 gnd.n5379 gnd.n5378 585
R1104 gnd.n4518 gnd.n4517 585
R1105 gnd.n4527 gnd.n4518 585
R1106 gnd.n5369 gnd.n5368 585
R1107 gnd.n5368 gnd.n5367 585
R1108 gnd.n4525 gnd.n4524 585
R1109 gnd.n5355 gnd.n4525 585
R1110 gnd.n5330 gnd.n4542 585
R1111 gnd.n5323 gnd.n4542 585
R1112 gnd.n5332 gnd.n5331 585
R1113 gnd.n5333 gnd.n5332 585
R1114 gnd.n4543 gnd.n4541 585
R1115 gnd.n4551 gnd.n4541 585
R1116 gnd.n5306 gnd.n4563 585
R1117 gnd.n4563 gnd.n4550 585
R1118 gnd.n5308 gnd.n5307 585
R1119 gnd.n5309 gnd.n5308 585
R1120 gnd.n4564 gnd.n4562 585
R1121 gnd.n4562 gnd.n4558 585
R1122 gnd.n5294 gnd.n5293 585
R1123 gnd.n5293 gnd.n5292 585
R1124 gnd.n4569 gnd.n4568 585
R1125 gnd.n4573 gnd.n4569 585
R1126 gnd.n5278 gnd.n5277 585
R1127 gnd.n5279 gnd.n5278 585
R1128 gnd.n4583 gnd.n4582 585
R1129 gnd.n5269 gnd.n4582 585
R1130 gnd.n5243 gnd.n4598 585
R1131 gnd.n4598 gnd.n4590 585
R1132 gnd.n5245 gnd.n5244 585
R1133 gnd.n5246 gnd.n5245 585
R1134 gnd.n4599 gnd.n4597 585
R1135 gnd.n4603 gnd.n4597 585
R1136 gnd.n5224 gnd.n5223 585
R1137 gnd.n5225 gnd.n5224 585
R1138 gnd.n4615 gnd.n4614 585
R1139 gnd.n4614 gnd.n4610 585
R1140 gnd.n5214 gnd.n5213 585
R1141 gnd.n5215 gnd.n5214 585
R1142 gnd.n4623 gnd.n4622 585
R1143 gnd.n4627 gnd.n4622 585
R1144 gnd.n5192 gnd.n4639 585
R1145 gnd.n4983 gnd.n4639 585
R1146 gnd.n5194 gnd.n5193 585
R1147 gnd.n5195 gnd.n5194 585
R1148 gnd.n4640 gnd.n4638 585
R1149 gnd.n4638 gnd.n4634 585
R1150 gnd.n5183 gnd.n5182 585
R1151 gnd.n5184 gnd.n5183 585
R1152 gnd.n4648 gnd.n4647 585
R1153 gnd.n4653 gnd.n4647 585
R1154 gnd.n5161 gnd.n4665 585
R1155 gnd.n4665 gnd.n4652 585
R1156 gnd.n5163 gnd.n5162 585
R1157 gnd.n5164 gnd.n5163 585
R1158 gnd.n4666 gnd.n4664 585
R1159 gnd.n4664 gnd.n4660 585
R1160 gnd.n5152 gnd.n5151 585
R1161 gnd.n5153 gnd.n5152 585
R1162 gnd.n4674 gnd.n4673 585
R1163 gnd.n5036 gnd.n4673 585
R1164 gnd.n5130 gnd.n4690 585
R1165 gnd.n4690 gnd.n4678 585
R1166 gnd.n5132 gnd.n5131 585
R1167 gnd.n5133 gnd.n5132 585
R1168 gnd.n4691 gnd.n4689 585
R1169 gnd.n4689 gnd.n4685 585
R1170 gnd.n5121 gnd.n5120 585
R1171 gnd.n5122 gnd.n5121 585
R1172 gnd.n4698 gnd.n4697 585
R1173 gnd.n4703 gnd.n4697 585
R1174 gnd.n5099 gnd.n4716 585
R1175 gnd.n4716 gnd.n4702 585
R1176 gnd.n5101 gnd.n5100 585
R1177 gnd.n5102 gnd.n5101 585
R1178 gnd.n4717 gnd.n4715 585
R1179 gnd.n4715 gnd.n4711 585
R1180 gnd.n5090 gnd.n5089 585
R1181 gnd.n5091 gnd.n5090 585
R1182 gnd.n4724 gnd.n4723 585
R1183 gnd.n4728 gnd.n4723 585
R1184 gnd.n5067 gnd.n4745 585
R1185 gnd.n4745 gnd.n4727 585
R1186 gnd.n5069 gnd.n5068 585
R1187 gnd.n5070 gnd.n5069 585
R1188 gnd.n4746 gnd.n4744 585
R1189 gnd.n4744 gnd.n4735 585
R1190 gnd.n5062 gnd.n5061 585
R1191 gnd.n5061 gnd.n5060 585
R1192 gnd.n4793 gnd.n4792 585
R1193 gnd.n4794 gnd.n4793 585
R1194 gnd.n4947 gnd.n4946 585
R1195 gnd.n4948 gnd.n4947 585
R1196 gnd.n4803 gnd.n4802 585
R1197 gnd.n4802 gnd.n4801 585
R1198 gnd.n4942 gnd.n4941 585
R1199 gnd.n4941 gnd.n4940 585
R1200 gnd.n4806 gnd.n4805 585
R1201 gnd.n4807 gnd.n4806 585
R1202 gnd.n4931 gnd.n4930 585
R1203 gnd.n4932 gnd.n4931 585
R1204 gnd.n4814 gnd.n4813 585
R1205 gnd.n4923 gnd.n4813 585
R1206 gnd.n4926 gnd.n4925 585
R1207 gnd.n4925 gnd.n4924 585
R1208 gnd.n4817 gnd.n4816 585
R1209 gnd.n4818 gnd.n4817 585
R1210 gnd.n4912 gnd.n4911 585
R1211 gnd.n4910 gnd.n4836 585
R1212 gnd.n4909 gnd.n4835 585
R1213 gnd.n4914 gnd.n4835 585
R1214 gnd.n4908 gnd.n4907 585
R1215 gnd.n4906 gnd.n4905 585
R1216 gnd.n4904 gnd.n4903 585
R1217 gnd.n4902 gnd.n4901 585
R1218 gnd.n4900 gnd.n4899 585
R1219 gnd.n4898 gnd.n4897 585
R1220 gnd.n4896 gnd.n4895 585
R1221 gnd.n4894 gnd.n4893 585
R1222 gnd.n4892 gnd.n4891 585
R1223 gnd.n4890 gnd.n4889 585
R1224 gnd.n4888 gnd.n4887 585
R1225 gnd.n4886 gnd.n4885 585
R1226 gnd.n4884 gnd.n4883 585
R1227 gnd.n4882 gnd.n4881 585
R1228 gnd.n4880 gnd.n4879 585
R1229 gnd.n4878 gnd.n4877 585
R1230 gnd.n4876 gnd.n4875 585
R1231 gnd.n4874 gnd.n4873 585
R1232 gnd.n4872 gnd.n4871 585
R1233 gnd.n4870 gnd.n4869 585
R1234 gnd.n4868 gnd.n4867 585
R1235 gnd.n4866 gnd.n4865 585
R1236 gnd.n4823 gnd.n4822 585
R1237 gnd.n4917 gnd.n4916 585
R1238 gnd.n5717 gnd.n5716 585
R1239 gnd.n5718 gnd.n4486 585
R1240 gnd.n5720 gnd.n5719 585
R1241 gnd.n5722 gnd.n4485 585
R1242 gnd.n5724 gnd.n5723 585
R1243 gnd.n5725 gnd.n4476 585
R1244 gnd.n5727 gnd.n5726 585
R1245 gnd.n5729 gnd.n4474 585
R1246 gnd.n5731 gnd.n5730 585
R1247 gnd.n5732 gnd.n4469 585
R1248 gnd.n5734 gnd.n5733 585
R1249 gnd.n5736 gnd.n4467 585
R1250 gnd.n5738 gnd.n5737 585
R1251 gnd.n5739 gnd.n4462 585
R1252 gnd.n5741 gnd.n5740 585
R1253 gnd.n5743 gnd.n4460 585
R1254 gnd.n5745 gnd.n5744 585
R1255 gnd.n5746 gnd.n4455 585
R1256 gnd.n5748 gnd.n5747 585
R1257 gnd.n5750 gnd.n4453 585
R1258 gnd.n5752 gnd.n5751 585
R1259 gnd.n5753 gnd.n4448 585
R1260 gnd.n5755 gnd.n5754 585
R1261 gnd.n5757 gnd.n4446 585
R1262 gnd.n5759 gnd.n5758 585
R1263 gnd.n5760 gnd.n4444 585
R1264 gnd.n5761 gnd.n798 585
R1265 gnd.n4407 gnd.n798 585
R1266 gnd.n5712 gnd.n800 585
R1267 gnd.n5799 gnd.n800 585
R1268 gnd.n5711 gnd.n5710 585
R1269 gnd.n5710 gnd.n5709 585
R1270 gnd.n5708 gnd.n790 585
R1271 gnd.n5805 gnd.n790 585
R1272 gnd.n5702 gnd.n4491 585
R1273 gnd.n5702 gnd.n788 585
R1274 gnd.n5704 gnd.n5703 585
R1275 gnd.n5703 gnd.n779 585
R1276 gnd.n5701 gnd.n777 585
R1277 gnd.n5813 gnd.n777 585
R1278 gnd.n5700 gnd.n5699 585
R1279 gnd.n5699 gnd.n5698 585
R1280 gnd.n4493 gnd.n766 585
R1281 gnd.n5819 gnd.n766 585
R1282 gnd.n5694 gnd.n5693 585
R1283 gnd.n5693 gnd.n5692 585
R1284 gnd.n4496 gnd.n4495 585
R1285 gnd.n4509 gnd.n4496 585
R1286 gnd.n5344 gnd.n4506 585
R1287 gnd.n5676 gnd.n4506 585
R1288 gnd.n5346 gnd.n5345 585
R1289 gnd.n5345 gnd.n4504 585
R1290 gnd.n5347 gnd.n4520 585
R1291 gnd.n5378 gnd.n4520 585
R1292 gnd.n5349 gnd.n5348 585
R1293 gnd.n5348 gnd.n4527 585
R1294 gnd.n5350 gnd.n4526 585
R1295 gnd.n5367 gnd.n4526 585
R1296 gnd.n5352 gnd.n5351 585
R1297 gnd.n5355 gnd.n5352 585
R1298 gnd.n4536 gnd.n4535 585
R1299 gnd.n5323 gnd.n4535 585
R1300 gnd.n5335 gnd.n5334 585
R1301 gnd.n5334 gnd.n5333 585
R1302 gnd.n4539 gnd.n4538 585
R1303 gnd.n4551 gnd.n4539 585
R1304 gnd.n5259 gnd.n5258 585
R1305 gnd.n5258 gnd.n4550 585
R1306 gnd.n5260 gnd.n4560 585
R1307 gnd.n5309 gnd.n4560 585
R1308 gnd.n5262 gnd.n5261 585
R1309 gnd.n5261 gnd.n4558 585
R1310 gnd.n5263 gnd.n4570 585
R1311 gnd.n5292 gnd.n4570 585
R1312 gnd.n5265 gnd.n5264 585
R1313 gnd.n5264 gnd.n4573 585
R1314 gnd.n5266 gnd.n4580 585
R1315 gnd.n5279 gnd.n4580 585
R1316 gnd.n5268 gnd.n5267 585
R1317 gnd.n5269 gnd.n5268 585
R1318 gnd.n4592 gnd.n4591 585
R1319 gnd.n4591 gnd.n4590 585
R1320 gnd.n5248 gnd.n5247 585
R1321 gnd.n5247 gnd.n5246 585
R1322 gnd.n4595 gnd.n4594 585
R1323 gnd.n4603 gnd.n4595 585
R1324 gnd.n4975 gnd.n4612 585
R1325 gnd.n5225 gnd.n4612 585
R1326 gnd.n4978 gnd.n4977 585
R1327 gnd.n4977 gnd.n4610 585
R1328 gnd.n4979 gnd.n4621 585
R1329 gnd.n5215 gnd.n4621 585
R1330 gnd.n4982 gnd.n4981 585
R1331 gnd.n4982 gnd.n4627 585
R1332 gnd.n4985 gnd.n4984 585
R1333 gnd.n4984 gnd.n4983 585
R1334 gnd.n4986 gnd.n4636 585
R1335 gnd.n5195 gnd.n4636 585
R1336 gnd.n4974 gnd.n4973 585
R1337 gnd.n4973 gnd.n4634 585
R1338 gnd.n5026 gnd.n4646 585
R1339 gnd.n5184 gnd.n4646 585
R1340 gnd.n5028 gnd.n5027 585
R1341 gnd.n5028 gnd.n4653 585
R1342 gnd.n5030 gnd.n5029 585
R1343 gnd.n5029 gnd.n4652 585
R1344 gnd.n5031 gnd.n4662 585
R1345 gnd.n5164 gnd.n4662 585
R1346 gnd.n5033 gnd.n5032 585
R1347 gnd.n5032 gnd.n4660 585
R1348 gnd.n5034 gnd.n4672 585
R1349 gnd.n5153 gnd.n4672 585
R1350 gnd.n5037 gnd.n5035 585
R1351 gnd.n5037 gnd.n5036 585
R1352 gnd.n5039 gnd.n5038 585
R1353 gnd.n5038 gnd.n4678 585
R1354 gnd.n5040 gnd.n4687 585
R1355 gnd.n5133 gnd.n4687 585
R1356 gnd.n5042 gnd.n5041 585
R1357 gnd.n5041 gnd.n4685 585
R1358 gnd.n5043 gnd.n4696 585
R1359 gnd.n5122 gnd.n4696 585
R1360 gnd.n5045 gnd.n5044 585
R1361 gnd.n5045 gnd.n4703 585
R1362 gnd.n5047 gnd.n5046 585
R1363 gnd.n5046 gnd.n4702 585
R1364 gnd.n5048 gnd.n4713 585
R1365 gnd.n5102 gnd.n4713 585
R1366 gnd.n5050 gnd.n5049 585
R1367 gnd.n5049 gnd.n4711 585
R1368 gnd.n5051 gnd.n4722 585
R1369 gnd.n5091 gnd.n4722 585
R1370 gnd.n5053 gnd.n5052 585
R1371 gnd.n5053 gnd.n4728 585
R1372 gnd.n5055 gnd.n5054 585
R1373 gnd.n5054 gnd.n4727 585
R1374 gnd.n5056 gnd.n4743 585
R1375 gnd.n5070 gnd.n4743 585
R1376 gnd.n5057 gnd.n4796 585
R1377 gnd.n4796 gnd.n4735 585
R1378 gnd.n5059 gnd.n5058 585
R1379 gnd.n5060 gnd.n5059 585
R1380 gnd.n4797 gnd.n4795 585
R1381 gnd.n4795 gnd.n4794 585
R1382 gnd.n4950 gnd.n4949 585
R1383 gnd.n4949 gnd.n4948 585
R1384 gnd.n4800 gnd.n4799 585
R1385 gnd.n4801 gnd.n4800 585
R1386 gnd.n4939 gnd.n4938 585
R1387 gnd.n4940 gnd.n4939 585
R1388 gnd.n4809 gnd.n4808 585
R1389 gnd.n4808 gnd.n4807 585
R1390 gnd.n4934 gnd.n4933 585
R1391 gnd.n4933 gnd.n4932 585
R1392 gnd.n4812 gnd.n4811 585
R1393 gnd.n4923 gnd.n4812 585
R1394 gnd.n4922 gnd.n4921 585
R1395 gnd.n4924 gnd.n4922 585
R1396 gnd.n4820 gnd.n4819 585
R1397 gnd.n4819 gnd.n4818 585
R1398 gnd.n5797 gnd.n5796 585
R1399 gnd.n5798 gnd.n5797 585
R1400 gnd.n4410 gnd.n4408 585
R1401 gnd.n4408 gnd.n799 585
R1402 gnd.n787 gnd.n786 585
R1403 gnd.n791 gnd.n787 585
R1404 gnd.n5808 gnd.n5807 585
R1405 gnd.n5807 gnd.n5806 585
R1406 gnd.n5809 gnd.n781 585
R1407 gnd.n5661 gnd.n781 585
R1408 gnd.n5811 gnd.n5810 585
R1409 gnd.n5812 gnd.n5811 585
R1410 gnd.n782 gnd.n780 585
R1411 gnd.n780 gnd.n776 585
R1412 gnd.n5687 gnd.n5686 585
R1413 gnd.n5686 gnd.n767 585
R1414 gnd.n5688 gnd.n4499 585
R1415 gnd.n4499 gnd.n765 585
R1416 gnd.n5690 gnd.n5689 585
R1417 gnd.n5691 gnd.n5690 585
R1418 gnd.n4500 gnd.n4498 585
R1419 gnd.n4507 gnd.n4498 585
R1420 gnd.n5679 gnd.n5678 585
R1421 gnd.n5678 gnd.n5677 585
R1422 gnd.n4503 gnd.n4502 585
R1423 gnd.n5377 gnd.n4503 585
R1424 gnd.n5363 gnd.n4529 585
R1425 gnd.n4529 gnd.n4519 585
R1426 gnd.n5365 gnd.n5364 585
R1427 gnd.n5366 gnd.n5365 585
R1428 gnd.n4530 gnd.n4528 585
R1429 gnd.n5354 gnd.n4528 585
R1430 gnd.n5358 gnd.n5357 585
R1431 gnd.n5357 gnd.n5356 585
R1432 gnd.n4533 gnd.n4532 585
R1433 gnd.n5324 gnd.n4533 585
R1434 gnd.n5317 gnd.n4553 585
R1435 gnd.n4553 gnd.n4540 585
R1436 gnd.n5319 gnd.n5318 585
R1437 gnd.n5320 gnd.n5319 585
R1438 gnd.n4554 gnd.n4552 585
R1439 gnd.n4561 gnd.n4552 585
R1440 gnd.n5312 gnd.n5311 585
R1441 gnd.n5311 gnd.n5310 585
R1442 gnd.n4557 gnd.n4556 585
R1443 gnd.n5291 gnd.n4557 585
R1444 gnd.n5287 gnd.n5286 585
R1445 gnd.n5288 gnd.n5287 585
R1446 gnd.n4575 gnd.n4574 585
R1447 gnd.n4581 gnd.n4574 585
R1448 gnd.n5282 gnd.n5281 585
R1449 gnd.n5281 gnd.n5280 585
R1450 gnd.n4578 gnd.n4577 585
R1451 gnd.n5270 gnd.n4578 585
R1452 gnd.n5233 gnd.n4605 585
R1453 gnd.n4605 gnd.n4596 585
R1454 gnd.n5235 gnd.n5234 585
R1455 gnd.n5236 gnd.n5235 585
R1456 gnd.n4606 gnd.n4604 585
R1457 gnd.n4613 gnd.n4604 585
R1458 gnd.n5228 gnd.n5227 585
R1459 gnd.n5227 gnd.n5226 585
R1460 gnd.n4609 gnd.n4608 585
R1461 gnd.n5216 gnd.n4609 585
R1462 gnd.n5203 gnd.n4629 585
R1463 gnd.n4629 gnd.n4620 585
R1464 gnd.n5205 gnd.n5204 585
R1465 gnd.n5206 gnd.n5205 585
R1466 gnd.n4630 gnd.n4628 585
R1467 gnd.n4637 gnd.n4628 585
R1468 gnd.n5198 gnd.n5197 585
R1469 gnd.n5197 gnd.n5196 585
R1470 gnd.n4633 gnd.n4632 585
R1471 gnd.n5185 gnd.n4633 585
R1472 gnd.n5172 gnd.n4655 585
R1473 gnd.n4655 gnd.n4645 585
R1474 gnd.n5174 gnd.n5173 585
R1475 gnd.n5175 gnd.n5174 585
R1476 gnd.n4656 gnd.n4654 585
R1477 gnd.n4663 gnd.n4654 585
R1478 gnd.n5167 gnd.n5166 585
R1479 gnd.n5166 gnd.n5165 585
R1480 gnd.n4659 gnd.n4658 585
R1481 gnd.n5154 gnd.n4659 585
R1482 gnd.n5141 gnd.n4680 585
R1483 gnd.n4680 gnd.n4671 585
R1484 gnd.n5143 gnd.n5142 585
R1485 gnd.n5144 gnd.n5143 585
R1486 gnd.n4681 gnd.n4679 585
R1487 gnd.n4688 gnd.n4679 585
R1488 gnd.n5136 gnd.n5135 585
R1489 gnd.n5135 gnd.n5134 585
R1490 gnd.n4684 gnd.n4683 585
R1491 gnd.n5123 gnd.n4684 585
R1492 gnd.n5110 gnd.n4706 585
R1493 gnd.n4706 gnd.n4705 585
R1494 gnd.n5112 gnd.n5111 585
R1495 gnd.n5113 gnd.n5112 585
R1496 gnd.n4707 gnd.n4704 585
R1497 gnd.n4714 gnd.n4704 585
R1498 gnd.n5105 gnd.n5104 585
R1499 gnd.n5104 gnd.n5103 585
R1500 gnd.n4710 gnd.n4709 585
R1501 gnd.n5092 gnd.n4710 585
R1502 gnd.n5079 gnd.n4731 585
R1503 gnd.n4731 gnd.n4730 585
R1504 gnd.n5081 gnd.n5080 585
R1505 gnd.n5082 gnd.n5081 585
R1506 gnd.n5075 gnd.n4729 585
R1507 gnd.n5074 gnd.n5073 585
R1508 gnd.n4734 gnd.n4733 585
R1509 gnd.n5071 gnd.n4734 585
R1510 gnd.n4756 gnd.n4755 585
R1511 gnd.n4759 gnd.n4758 585
R1512 gnd.n4757 gnd.n4752 585
R1513 gnd.n4764 gnd.n4763 585
R1514 gnd.n4766 gnd.n4765 585
R1515 gnd.n4769 gnd.n4768 585
R1516 gnd.n4767 gnd.n4750 585
R1517 gnd.n4774 gnd.n4773 585
R1518 gnd.n4776 gnd.n4775 585
R1519 gnd.n4779 gnd.n4778 585
R1520 gnd.n4777 gnd.n4748 585
R1521 gnd.n4784 gnd.n4783 585
R1522 gnd.n4788 gnd.n4785 585
R1523 gnd.n4789 gnd.n4726 585
R1524 gnd.n5766 gnd.n5765 585
R1525 gnd.n5768 gnd.n4439 585
R1526 gnd.n5770 gnd.n5769 585
R1527 gnd.n5771 gnd.n4432 585
R1528 gnd.n5773 gnd.n5772 585
R1529 gnd.n5775 gnd.n4430 585
R1530 gnd.n5777 gnd.n5776 585
R1531 gnd.n5778 gnd.n4425 585
R1532 gnd.n5780 gnd.n5779 585
R1533 gnd.n5782 gnd.n4423 585
R1534 gnd.n5784 gnd.n5783 585
R1535 gnd.n5785 gnd.n4418 585
R1536 gnd.n5787 gnd.n5786 585
R1537 gnd.n5789 gnd.n4416 585
R1538 gnd.n5791 gnd.n5790 585
R1539 gnd.n5792 gnd.n4414 585
R1540 gnd.n5793 gnd.n4409 585
R1541 gnd.n4409 gnd.n4407 585
R1542 gnd.n5655 gnd.n801 585
R1543 gnd.n5798 gnd.n801 585
R1544 gnd.n5657 gnd.n5656 585
R1545 gnd.n5657 gnd.n799 585
R1546 gnd.n5659 gnd.n5658 585
R1547 gnd.n5658 gnd.n791 585
R1548 gnd.n5660 gnd.n789 585
R1549 gnd.n5806 gnd.n789 585
R1550 gnd.n5663 gnd.n5662 585
R1551 gnd.n5662 gnd.n5661 585
R1552 gnd.n5664 gnd.n778 585
R1553 gnd.n5812 gnd.n778 585
R1554 gnd.n5666 gnd.n5665 585
R1555 gnd.n5666 gnd.n776 585
R1556 gnd.n5667 gnd.n5390 585
R1557 gnd.n5667 gnd.n767 585
R1558 gnd.n5669 gnd.n5668 585
R1559 gnd.n5668 gnd.n765 585
R1560 gnd.n5670 gnd.n4497 585
R1561 gnd.n5691 gnd.n4497 585
R1562 gnd.n5387 gnd.n5386 585
R1563 gnd.n5386 gnd.n4507 585
R1564 gnd.n5385 gnd.n4505 585
R1565 gnd.n5677 gnd.n4505 585
R1566 gnd.n5376 gnd.n4515 585
R1567 gnd.n5377 gnd.n5376 585
R1568 gnd.n5375 gnd.n5374 585
R1569 gnd.n5375 gnd.n4519 585
R1570 gnd.n5373 gnd.n4521 585
R1571 gnd.n5366 gnd.n4521 585
R1572 gnd.n5353 gnd.n4522 585
R1573 gnd.n5354 gnd.n5353 585
R1574 gnd.n5327 gnd.n4534 585
R1575 gnd.n5356 gnd.n4534 585
R1576 gnd.n5326 gnd.n5325 585
R1577 gnd.n5325 gnd.n5324 585
R1578 gnd.n5322 gnd.n4547 585
R1579 gnd.n5322 gnd.n4540 585
R1580 gnd.n5321 gnd.n4549 585
R1581 gnd.n5321 gnd.n5320 585
R1582 gnd.n5300 gnd.n4548 585
R1583 gnd.n4561 gnd.n4548 585
R1584 gnd.n5299 gnd.n4559 585
R1585 gnd.n5310 gnd.n4559 585
R1586 gnd.n5290 gnd.n4566 585
R1587 gnd.n5291 gnd.n5290 585
R1588 gnd.n5289 gnd.n4572 585
R1589 gnd.n5289 gnd.n5288 585
R1590 gnd.n5274 gnd.n4571 585
R1591 gnd.n4581 gnd.n4571 585
R1592 gnd.n5273 gnd.n4579 585
R1593 gnd.n5280 gnd.n4579 585
R1594 gnd.n5272 gnd.n5271 585
R1595 gnd.n5271 gnd.n5270 585
R1596 gnd.n4589 gnd.n4586 585
R1597 gnd.n4596 gnd.n4589 585
R1598 gnd.n5238 gnd.n5237 585
R1599 gnd.n5237 gnd.n5236 585
R1600 gnd.n4602 gnd.n4601 585
R1601 gnd.n4613 gnd.n4602 585
R1602 gnd.n5219 gnd.n4611 585
R1603 gnd.n5226 gnd.n4611 585
R1604 gnd.n5218 gnd.n5217 585
R1605 gnd.n5217 gnd.n5216 585
R1606 gnd.n4619 gnd.n4617 585
R1607 gnd.n4620 gnd.n4619 585
R1608 gnd.n5208 gnd.n5207 585
R1609 gnd.n5207 gnd.n5206 585
R1610 gnd.n4626 gnd.n4625 585
R1611 gnd.n4637 gnd.n4626 585
R1612 gnd.n5188 gnd.n4635 585
R1613 gnd.n5196 gnd.n4635 585
R1614 gnd.n5187 gnd.n5186 585
R1615 gnd.n5186 gnd.n5185 585
R1616 gnd.n4644 gnd.n4642 585
R1617 gnd.n4645 gnd.n4644 585
R1618 gnd.n5177 gnd.n5176 585
R1619 gnd.n5176 gnd.n5175 585
R1620 gnd.n4651 gnd.n4650 585
R1621 gnd.n4663 gnd.n4651 585
R1622 gnd.n5157 gnd.n4661 585
R1623 gnd.n5165 gnd.n4661 585
R1624 gnd.n5156 gnd.n5155 585
R1625 gnd.n5155 gnd.n5154 585
R1626 gnd.n4670 gnd.n4668 585
R1627 gnd.n4671 gnd.n4670 585
R1628 gnd.n5146 gnd.n5145 585
R1629 gnd.n5145 gnd.n5144 585
R1630 gnd.n4677 gnd.n4676 585
R1631 gnd.n4688 gnd.n4677 585
R1632 gnd.n5126 gnd.n4686 585
R1633 gnd.n5134 gnd.n4686 585
R1634 gnd.n5125 gnd.n5124 585
R1635 gnd.n5124 gnd.n5123 585
R1636 gnd.n4695 gnd.n4693 585
R1637 gnd.n4705 gnd.n4695 585
R1638 gnd.n5115 gnd.n5114 585
R1639 gnd.n5114 gnd.n5113 585
R1640 gnd.n4701 gnd.n4700 585
R1641 gnd.n4714 gnd.n4701 585
R1642 gnd.n5095 gnd.n4712 585
R1643 gnd.n5103 gnd.n4712 585
R1644 gnd.n5094 gnd.n5093 585
R1645 gnd.n5093 gnd.n5092 585
R1646 gnd.n4721 gnd.n4719 585
R1647 gnd.n4730 gnd.n4721 585
R1648 gnd.n5084 gnd.n5083 585
R1649 gnd.n5083 gnd.n5082 585
R1650 gnd.n4203 gnd.n4202 585
R1651 gnd.n4202 gnd.n4201 585
R1652 gnd.n4204 gnd.n1073 585
R1653 gnd.n2418 gnd.n1073 585
R1654 gnd.n4206 gnd.n4205 585
R1655 gnd.n4207 gnd.n4206 585
R1656 gnd.n1057 gnd.n1056 585
R1657 gnd.n2378 gnd.n1057 585
R1658 gnd.n4215 gnd.n4214 585
R1659 gnd.n4214 gnd.n4213 585
R1660 gnd.n4216 gnd.n1051 585
R1661 gnd.n2369 gnd.n1051 585
R1662 gnd.n4218 gnd.n4217 585
R1663 gnd.n4219 gnd.n4218 585
R1664 gnd.n1036 gnd.n1035 585
R1665 gnd.n2361 gnd.n1036 585
R1666 gnd.n4227 gnd.n4226 585
R1667 gnd.n4226 gnd.n4225 585
R1668 gnd.n4228 gnd.n1030 585
R1669 gnd.n2286 gnd.n1030 585
R1670 gnd.n4230 gnd.n4229 585
R1671 gnd.n4231 gnd.n4230 585
R1672 gnd.n1015 gnd.n1014 585
R1673 gnd.n2274 gnd.n1015 585
R1674 gnd.n4239 gnd.n4238 585
R1675 gnd.n4238 gnd.n4237 585
R1676 gnd.n4240 gnd.n1009 585
R1677 gnd.n2269 gnd.n1009 585
R1678 gnd.n4242 gnd.n4241 585
R1679 gnd.n4243 gnd.n4242 585
R1680 gnd.n994 gnd.n993 585
R1681 gnd.n2300 gnd.n994 585
R1682 gnd.n4251 gnd.n4250 585
R1683 gnd.n4250 gnd.n4249 585
R1684 gnd.n4252 gnd.n991 585
R1685 gnd.n2261 gnd.n991 585
R1686 gnd.n4255 gnd.n4254 585
R1687 gnd.n4256 gnd.n4255 585
R1688 gnd.n992 gnd.n977 585
R1689 gnd.n2253 gnd.n977 585
R1690 gnd.n4264 gnd.n4263 585
R1691 gnd.n4263 gnd.n4262 585
R1692 gnd.n4265 gnd.n974 585
R1693 gnd.n2244 gnd.n974 585
R1694 gnd.n4268 gnd.n4267 585
R1695 gnd.n4269 gnd.n4268 585
R1696 gnd.n975 gnd.n956 585
R1697 gnd.n960 gnd.n956 585
R1698 gnd.n4277 gnd.n4276 585
R1699 gnd.n4276 gnd.n4275 585
R1700 gnd.n4278 gnd.n954 585
R1701 gnd.n2233 gnd.n954 585
R1702 gnd.n4280 gnd.n950 585
R1703 gnd.n950 gnd.n949 585
R1704 gnd.n4282 gnd.n4281 585
R1705 gnd.n4283 gnd.n4282 585
R1706 gnd.n935 gnd.n934 585
R1707 gnd.n939 gnd.n935 585
R1708 gnd.n4291 gnd.n4290 585
R1709 gnd.n4290 gnd.n4289 585
R1710 gnd.n4292 gnd.n929 585
R1711 gnd.n936 gnd.n929 585
R1712 gnd.n4294 gnd.n4293 585
R1713 gnd.n4295 gnd.n4294 585
R1714 gnd.n916 gnd.n915 585
R1715 gnd.n926 gnd.n916 585
R1716 gnd.n4303 gnd.n4302 585
R1717 gnd.n4302 gnd.n4301 585
R1718 gnd.n4304 gnd.n910 585
R1719 gnd.n910 gnd.n909 585
R1720 gnd.n4306 gnd.n4305 585
R1721 gnd.n4307 gnd.n4306 585
R1722 gnd.n895 gnd.n894 585
R1723 gnd.n898 gnd.n895 585
R1724 gnd.n4315 gnd.n4314 585
R1725 gnd.n4314 gnd.n4313 585
R1726 gnd.n4316 gnd.n889 585
R1727 gnd.n889 gnd.n886 585
R1728 gnd.n4318 gnd.n4317 585
R1729 gnd.n4319 gnd.n4318 585
R1730 gnd.n890 gnd.n888 585
R1731 gnd.n888 gnd.n884 585
R1732 gnd.n2164 gnd.n2163 585
R1733 gnd.n2165 gnd.n2164 585
R1734 gnd.n2159 gnd.n833 585
R1735 gnd.n833 gnd.n830 585
R1736 gnd.n4404 gnd.n4403 585
R1737 gnd.n4402 gnd.n832 585
R1738 gnd.n4401 gnd.n831 585
R1739 gnd.n4406 gnd.n831 585
R1740 gnd.n4400 gnd.n4399 585
R1741 gnd.n4398 gnd.n4397 585
R1742 gnd.n4396 gnd.n4395 585
R1743 gnd.n4394 gnd.n4393 585
R1744 gnd.n4392 gnd.n4391 585
R1745 gnd.n4390 gnd.n4389 585
R1746 gnd.n4388 gnd.n4387 585
R1747 gnd.n4386 gnd.n4385 585
R1748 gnd.n4384 gnd.n4383 585
R1749 gnd.n4382 gnd.n4381 585
R1750 gnd.n4380 gnd.n4379 585
R1751 gnd.n4378 gnd.n4377 585
R1752 gnd.n4376 gnd.n4375 585
R1753 gnd.n4374 gnd.n4373 585
R1754 gnd.n4372 gnd.n4371 585
R1755 gnd.n4369 gnd.n4368 585
R1756 gnd.n4367 gnd.n4366 585
R1757 gnd.n4365 gnd.n4364 585
R1758 gnd.n4363 gnd.n4362 585
R1759 gnd.n4361 gnd.n4360 585
R1760 gnd.n4359 gnd.n4358 585
R1761 gnd.n4357 gnd.n4356 585
R1762 gnd.n4355 gnd.n4354 585
R1763 gnd.n4353 gnd.n4352 585
R1764 gnd.n4351 gnd.n4350 585
R1765 gnd.n4349 gnd.n4348 585
R1766 gnd.n4347 gnd.n4346 585
R1767 gnd.n4345 gnd.n4344 585
R1768 gnd.n4343 gnd.n4342 585
R1769 gnd.n4341 gnd.n4340 585
R1770 gnd.n4339 gnd.n4338 585
R1771 gnd.n4337 gnd.n4336 585
R1772 gnd.n4335 gnd.n4334 585
R1773 gnd.n4333 gnd.n872 585
R1774 gnd.n876 gnd.n873 585
R1775 gnd.n4329 gnd.n4328 585
R1776 gnd.n1995 gnd.n1994 585
R1777 gnd.n2426 gnd.n2425 585
R1778 gnd.n2428 gnd.n2427 585
R1779 gnd.n2430 gnd.n2429 585
R1780 gnd.n2432 gnd.n2431 585
R1781 gnd.n2434 gnd.n2433 585
R1782 gnd.n2436 gnd.n2435 585
R1783 gnd.n2438 gnd.n2437 585
R1784 gnd.n2440 gnd.n2439 585
R1785 gnd.n2442 gnd.n2441 585
R1786 gnd.n2444 gnd.n2443 585
R1787 gnd.n2446 gnd.n2445 585
R1788 gnd.n2448 gnd.n2447 585
R1789 gnd.n2450 gnd.n2449 585
R1790 gnd.n2452 gnd.n2451 585
R1791 gnd.n2454 gnd.n2453 585
R1792 gnd.n2456 gnd.n2455 585
R1793 gnd.n2458 gnd.n2457 585
R1794 gnd.n2460 gnd.n2459 585
R1795 gnd.n2463 gnd.n2462 585
R1796 gnd.n2461 gnd.n1973 585
R1797 gnd.n2598 gnd.n2597 585
R1798 gnd.n2600 gnd.n2599 585
R1799 gnd.n2602 gnd.n2601 585
R1800 gnd.n2604 gnd.n2603 585
R1801 gnd.n2606 gnd.n2605 585
R1802 gnd.n2608 gnd.n2607 585
R1803 gnd.n2610 gnd.n2609 585
R1804 gnd.n2612 gnd.n2611 585
R1805 gnd.n2614 gnd.n2613 585
R1806 gnd.n2616 gnd.n2615 585
R1807 gnd.n2618 gnd.n2617 585
R1808 gnd.n2620 gnd.n2619 585
R1809 gnd.n2621 gnd.n1954 585
R1810 gnd.n2623 gnd.n2622 585
R1811 gnd.n1955 gnd.n1953 585
R1812 gnd.n1956 gnd.n1078 585
R1813 gnd.n2625 gnd.n1078 585
R1814 gnd.n2421 gnd.n1080 585
R1815 gnd.n4201 gnd.n1080 585
R1816 gnd.n2420 gnd.n2419 585
R1817 gnd.n2419 gnd.n2418 585
R1818 gnd.n1999 gnd.n1070 585
R1819 gnd.n4207 gnd.n1070 585
R1820 gnd.n2377 gnd.n2376 585
R1821 gnd.n2378 gnd.n2377 585
R1822 gnd.n2004 gnd.n1059 585
R1823 gnd.n4213 gnd.n1059 585
R1824 gnd.n2371 gnd.n2370 585
R1825 gnd.n2370 gnd.n2369 585
R1826 gnd.n2006 gnd.n1048 585
R1827 gnd.n4219 gnd.n1048 585
R1828 gnd.n2282 gnd.n2010 585
R1829 gnd.n2361 gnd.n2010 585
R1830 gnd.n2283 gnd.n1038 585
R1831 gnd.n4225 gnd.n1038 585
R1832 gnd.n2285 gnd.n2284 585
R1833 gnd.n2286 gnd.n2285 585
R1834 gnd.n2030 gnd.n1027 585
R1835 gnd.n4231 gnd.n1027 585
R1836 gnd.n2276 gnd.n2275 585
R1837 gnd.n2275 gnd.n2274 585
R1838 gnd.n2272 gnd.n1017 585
R1839 gnd.n4237 gnd.n1017 585
R1840 gnd.n2271 gnd.n2270 585
R1841 gnd.n2270 gnd.n2269 585
R1842 gnd.n2032 gnd.n1006 585
R1843 gnd.n4243 gnd.n1006 585
R1844 gnd.n2265 gnd.n2022 585
R1845 gnd.n2300 gnd.n2022 585
R1846 gnd.n2264 gnd.n996 585
R1847 gnd.n4249 gnd.n996 585
R1848 gnd.n2263 gnd.n2262 585
R1849 gnd.n2262 gnd.n2261 585
R1850 gnd.n2034 gnd.n988 585
R1851 gnd.n4256 gnd.n988 585
R1852 gnd.n2252 gnd.n2251 585
R1853 gnd.n2253 gnd.n2252 585
R1854 gnd.n2067 gnd.n979 585
R1855 gnd.n4262 gnd.n979 585
R1856 gnd.n2246 gnd.n2245 585
R1857 gnd.n2245 gnd.n2244 585
R1858 gnd.n2070 gnd.n971 585
R1859 gnd.n4269 gnd.n971 585
R1860 gnd.n2229 gnd.n2228 585
R1861 gnd.n2228 gnd.n960 585
R1862 gnd.n2230 gnd.n958 585
R1863 gnd.n4275 gnd.n958 585
R1864 gnd.n2232 gnd.n2231 585
R1865 gnd.n2233 gnd.n2232 585
R1866 gnd.n2196 gnd.n2195 585
R1867 gnd.n2195 gnd.n949 585
R1868 gnd.n2222 gnd.n947 585
R1869 gnd.n4283 gnd.n947 585
R1870 gnd.n2221 gnd.n2220 585
R1871 gnd.n2220 gnd.n939 585
R1872 gnd.n2219 gnd.n937 585
R1873 gnd.n4289 gnd.n937 585
R1874 gnd.n2199 gnd.n2198 585
R1875 gnd.n2198 gnd.n936 585
R1876 gnd.n2215 gnd.n927 585
R1877 gnd.n4295 gnd.n927 585
R1878 gnd.n2214 gnd.n2213 585
R1879 gnd.n2213 gnd.n926 585
R1880 gnd.n2212 gnd.n917 585
R1881 gnd.n4301 gnd.n917 585
R1882 gnd.n2202 gnd.n2201 585
R1883 gnd.n2201 gnd.n909 585
R1884 gnd.n2208 gnd.n907 585
R1885 gnd.n4307 gnd.n907 585
R1886 gnd.n2207 gnd.n2206 585
R1887 gnd.n2206 gnd.n898 585
R1888 gnd.n2205 gnd.n896 585
R1889 gnd.n4313 gnd.n896 585
R1890 gnd.n883 gnd.n881 585
R1891 gnd.n886 gnd.n883 585
R1892 gnd.n4321 gnd.n4320 585
R1893 gnd.n4320 gnd.n4319 585
R1894 gnd.n882 gnd.n879 585
R1895 gnd.n884 gnd.n882 585
R1896 gnd.n4325 gnd.n878 585
R1897 gnd.n2165 gnd.n878 585
R1898 gnd.n4327 gnd.n4326 585
R1899 gnd.n4327 gnd.n830 585
R1900 gnd.n6804 gnd.n6803 585
R1901 gnd.n6805 gnd.n6804 585
R1902 gnd.n87 gnd.n85 585
R1903 gnd.n85 gnd.n81 585
R1904 gnd.n6724 gnd.n6723 585
R1905 gnd.n6725 gnd.n6724 585
R1906 gnd.n165 gnd.n164 585
R1907 gnd.n164 gnd.n161 585
R1908 gnd.n6719 gnd.n6718 585
R1909 gnd.n6718 gnd.n6717 585
R1910 gnd.n168 gnd.n167 585
R1911 gnd.n170 gnd.n168 585
R1912 gnd.n6634 gnd.n6633 585
R1913 gnd.n6635 gnd.n6634 585
R1914 gnd.n181 gnd.n180 585
R1915 gnd.n188 gnd.n180 585
R1916 gnd.n6629 gnd.n6628 585
R1917 gnd.n6628 gnd.n6627 585
R1918 gnd.n184 gnd.n183 585
R1919 gnd.n186 gnd.n184 585
R1920 gnd.n6618 gnd.n6617 585
R1921 gnd.n6619 gnd.n6618 585
R1922 gnd.n197 gnd.n196 585
R1923 gnd.n196 gnd.n194 585
R1924 gnd.n6613 gnd.n6612 585
R1925 gnd.n6612 gnd.n6611 585
R1926 gnd.n200 gnd.n199 585
R1927 gnd.n202 gnd.n200 585
R1928 gnd.n6602 gnd.n6601 585
R1929 gnd.n6603 gnd.n6602 585
R1930 gnd.n211 gnd.n210 585
R1931 gnd.n224 gnd.n210 585
R1932 gnd.n6597 gnd.n6596 585
R1933 gnd.n6596 gnd.n6595 585
R1934 gnd.n220 gnd.n219 585
R1935 gnd.n222 gnd.n220 585
R1936 gnd.n6586 gnd.n6585 585
R1937 gnd.n6587 gnd.n6586 585
R1938 gnd.n6584 gnd.n6583 585
R1939 gnd.n6583 gnd.n230 585
R1940 gnd.n6582 gnd.n235 585
R1941 gnd.n6582 gnd.n6581 585
R1942 gnd.n234 gnd.n233 585
R1943 gnd.n3890 gnd.n233 585
R1944 gnd.n6572 gnd.n6571 585
R1945 gnd.n6573 gnd.n6572 585
R1946 gnd.n6570 gnd.n6569 585
R1947 gnd.n6569 gnd.n6568 585
R1948 gnd.n1264 gnd.n247 585
R1949 gnd.n4019 gnd.n247 585
R1950 gnd.n1266 gnd.n1265 585
R1951 gnd.n3896 gnd.n1266 585
R1952 gnd.n4009 gnd.n4008 585
R1953 gnd.n4010 gnd.n4009 585
R1954 gnd.n4007 gnd.n1263 585
R1955 gnd.n1274 gnd.n1263 585
R1956 gnd.n4006 gnd.n4005 585
R1957 gnd.n4005 gnd.n4004 585
R1958 gnd.n1269 gnd.n1267 585
R1959 gnd.n3985 gnd.n1269 585
R1960 gnd.n3973 gnd.n1294 585
R1961 gnd.n1294 gnd.n1281 585
R1962 gnd.n3975 gnd.n3974 585
R1963 gnd.n3976 gnd.n3975 585
R1964 gnd.n1295 gnd.n1293 585
R1965 gnd.n1302 gnd.n1293 585
R1966 gnd.n3967 gnd.n3966 585
R1967 gnd.n3966 gnd.n3965 585
R1968 gnd.n1298 gnd.n1297 585
R1969 gnd.n3953 gnd.n1298 585
R1970 gnd.n3941 gnd.n1322 585
R1971 gnd.n1322 gnd.n1310 585
R1972 gnd.n3943 gnd.n3942 585
R1973 gnd.n3944 gnd.n3943 585
R1974 gnd.n1323 gnd.n1321 585
R1975 gnd.n3916 gnd.n1321 585
R1976 gnd.n3936 gnd.n3935 585
R1977 gnd.n3935 gnd.n3934 585
R1978 gnd.n1223 gnd.n1222 585
R1979 gnd.n3823 gnd.n1223 585
R1980 gnd.n4050 gnd.n4049 585
R1981 gnd.n4049 gnd.n4048 585
R1982 gnd.n4051 gnd.n1218 585
R1983 gnd.n3814 gnd.n1218 585
R1984 gnd.n4053 gnd.n4052 585
R1985 gnd.n4054 gnd.n4053 585
R1986 gnd.n3713 gnd.n1217 585
R1987 gnd.n3718 gnd.n3716 585
R1988 gnd.n3719 gnd.n3712 585
R1989 gnd.n3719 gnd.n1204 585
R1990 gnd.n3722 gnd.n3721 585
R1991 gnd.n3710 gnd.n3709 585
R1992 gnd.n3727 gnd.n3726 585
R1993 gnd.n3729 gnd.n3708 585
R1994 gnd.n3732 gnd.n3731 585
R1995 gnd.n3706 gnd.n3705 585
R1996 gnd.n3737 gnd.n3736 585
R1997 gnd.n3739 gnd.n3704 585
R1998 gnd.n3742 gnd.n3741 585
R1999 gnd.n3702 gnd.n3701 585
R2000 gnd.n3748 gnd.n3747 585
R2001 gnd.n3750 gnd.n3700 585
R2002 gnd.n3751 gnd.n1360 585
R2003 gnd.n1358 gnd.n1357 585
R2004 gnd.n3761 gnd.n3760 585
R2005 gnd.n3763 gnd.n1356 585
R2006 gnd.n3766 gnd.n3765 585
R2007 gnd.n1354 gnd.n1353 585
R2008 gnd.n3771 gnd.n3770 585
R2009 gnd.n3773 gnd.n1352 585
R2010 gnd.n3776 gnd.n3775 585
R2011 gnd.n1350 gnd.n1349 585
R2012 gnd.n3781 gnd.n3780 585
R2013 gnd.n3783 gnd.n1348 585
R2014 gnd.n3786 gnd.n3785 585
R2015 gnd.n1346 gnd.n1345 585
R2016 gnd.n3791 gnd.n3790 585
R2017 gnd.n3793 gnd.n1344 585
R2018 gnd.n3796 gnd.n3795 585
R2019 gnd.n1342 gnd.n1341 585
R2020 gnd.n3802 gnd.n3801 585
R2021 gnd.n3804 gnd.n1340 585
R2022 gnd.n3805 gnd.n1339 585
R2023 gnd.n3808 gnd.n3807 585
R2024 gnd.n155 gnd.n154 585
R2025 gnd.n6733 gnd.n150 585
R2026 gnd.n6735 gnd.n6734 585
R2027 gnd.n6737 gnd.n148 585
R2028 gnd.n6739 gnd.n6738 585
R2029 gnd.n6740 gnd.n143 585
R2030 gnd.n6742 gnd.n6741 585
R2031 gnd.n6744 gnd.n141 585
R2032 gnd.n6746 gnd.n6745 585
R2033 gnd.n6747 gnd.n136 585
R2034 gnd.n6749 gnd.n6748 585
R2035 gnd.n6751 gnd.n134 585
R2036 gnd.n6753 gnd.n6752 585
R2037 gnd.n6754 gnd.n129 585
R2038 gnd.n6756 gnd.n6755 585
R2039 gnd.n6758 gnd.n127 585
R2040 gnd.n6760 gnd.n6759 585
R2041 gnd.n6761 gnd.n122 585
R2042 gnd.n6763 gnd.n6762 585
R2043 gnd.n6765 gnd.n120 585
R2044 gnd.n6767 gnd.n6766 585
R2045 gnd.n6771 gnd.n115 585
R2046 gnd.n6773 gnd.n6772 585
R2047 gnd.n6775 gnd.n113 585
R2048 gnd.n6777 gnd.n6776 585
R2049 gnd.n6778 gnd.n108 585
R2050 gnd.n6780 gnd.n6779 585
R2051 gnd.n6782 gnd.n106 585
R2052 gnd.n6784 gnd.n6783 585
R2053 gnd.n6785 gnd.n101 585
R2054 gnd.n6787 gnd.n6786 585
R2055 gnd.n6789 gnd.n99 585
R2056 gnd.n6791 gnd.n6790 585
R2057 gnd.n6792 gnd.n94 585
R2058 gnd.n6794 gnd.n6793 585
R2059 gnd.n6796 gnd.n92 585
R2060 gnd.n6798 gnd.n6797 585
R2061 gnd.n6799 gnd.n90 585
R2062 gnd.n6800 gnd.n86 585
R2063 gnd.n86 gnd.n83 585
R2064 gnd.n6729 gnd.n82 585
R2065 gnd.n6805 gnd.n82 585
R2066 gnd.n6728 gnd.n6727 585
R2067 gnd.n6727 gnd.n81 585
R2068 gnd.n6726 gnd.n159 585
R2069 gnd.n6726 gnd.n6725 585
R2070 gnd.n3863 gnd.n160 585
R2071 gnd.n161 gnd.n160 585
R2072 gnd.n3864 gnd.n171 585
R2073 gnd.n6717 gnd.n171 585
R2074 gnd.n3866 gnd.n3865 585
R2075 gnd.n3865 gnd.n170 585
R2076 gnd.n3867 gnd.n179 585
R2077 gnd.n6635 gnd.n179 585
R2078 gnd.n3869 gnd.n3868 585
R2079 gnd.n3868 gnd.n188 585
R2080 gnd.n3870 gnd.n187 585
R2081 gnd.n6627 gnd.n187 585
R2082 gnd.n3872 gnd.n3871 585
R2083 gnd.n3871 gnd.n186 585
R2084 gnd.n3873 gnd.n195 585
R2085 gnd.n6619 gnd.n195 585
R2086 gnd.n3875 gnd.n3874 585
R2087 gnd.n3874 gnd.n194 585
R2088 gnd.n3876 gnd.n203 585
R2089 gnd.n6611 gnd.n203 585
R2090 gnd.n3878 gnd.n3877 585
R2091 gnd.n3877 gnd.n202 585
R2092 gnd.n3879 gnd.n209 585
R2093 gnd.n6603 gnd.n209 585
R2094 gnd.n3881 gnd.n3880 585
R2095 gnd.n3880 gnd.n224 585
R2096 gnd.n3882 gnd.n223 585
R2097 gnd.n6595 gnd.n223 585
R2098 gnd.n3884 gnd.n3883 585
R2099 gnd.n3883 gnd.n222 585
R2100 gnd.n3885 gnd.n231 585
R2101 gnd.n6587 gnd.n231 585
R2102 gnd.n3887 gnd.n3886 585
R2103 gnd.n3886 gnd.n230 585
R2104 gnd.n3888 gnd.n237 585
R2105 gnd.n6581 gnd.n237 585
R2106 gnd.n3892 gnd.n3891 585
R2107 gnd.n3891 gnd.n3890 585
R2108 gnd.n3893 gnd.n244 585
R2109 gnd.n6573 gnd.n244 585
R2110 gnd.n3894 gnd.n249 585
R2111 gnd.n6568 gnd.n249 585
R2112 gnd.n3895 gnd.n1252 585
R2113 gnd.n4019 gnd.n1252 585
R2114 gnd.n3898 gnd.n3897 585
R2115 gnd.n3897 gnd.n3896 585
R2116 gnd.n3899 gnd.n1261 585
R2117 gnd.n4010 gnd.n1261 585
R2118 gnd.n3901 gnd.n3900 585
R2119 gnd.n3900 gnd.n1274 585
R2120 gnd.n3902 gnd.n1271 585
R2121 gnd.n4004 gnd.n1271 585
R2122 gnd.n3903 gnd.n1282 585
R2123 gnd.n3985 gnd.n1282 585
R2124 gnd.n3905 gnd.n3904 585
R2125 gnd.n3904 gnd.n1281 585
R2126 gnd.n3906 gnd.n1290 585
R2127 gnd.n3976 gnd.n1290 585
R2128 gnd.n3908 gnd.n3907 585
R2129 gnd.n3907 gnd.n1302 585
R2130 gnd.n3909 gnd.n1300 585
R2131 gnd.n3965 gnd.n1300 585
R2132 gnd.n3910 gnd.n1311 585
R2133 gnd.n3953 gnd.n1311 585
R2134 gnd.n3912 gnd.n3911 585
R2135 gnd.n3911 gnd.n1310 585
R2136 gnd.n3913 gnd.n1319 585
R2137 gnd.n3944 gnd.n1319 585
R2138 gnd.n3915 gnd.n3914 585
R2139 gnd.n3916 gnd.n3915 585
R2140 gnd.n1328 gnd.n1326 585
R2141 gnd.n3934 gnd.n1326 585
R2142 gnd.n3825 gnd.n3824 585
R2143 gnd.n3824 gnd.n3823 585
R2144 gnd.n1330 gnd.n1225 585
R2145 gnd.n4048 gnd.n1225 585
R2146 gnd.n3813 gnd.n3812 585
R2147 gnd.n3814 gnd.n3813 585
R2148 gnd.n1335 gnd.n1213 585
R2149 gnd.n4054 gnd.n1213 585
R2150 gnd.n3627 gnd.n3626 585
R2151 gnd.n3628 gnd.n3627 585
R2152 gnd.n3541 gnd.n1404 585
R2153 gnd.n1411 gnd.n1404 585
R2154 gnd.n3540 gnd.n3539 585
R2155 gnd.n3539 gnd.n3538 585
R2156 gnd.n1407 gnd.n1406 585
R2157 gnd.t161 gnd.n1407 585
R2158 gnd.n3278 gnd.n1472 585
R2159 gnd.n1472 gnd.n1471 585
R2160 gnd.n3280 gnd.n3279 585
R2161 gnd.n3281 gnd.n3280 585
R2162 gnd.n3277 gnd.n1470 585
R2163 gnd.n1478 gnd.n1470 585
R2164 gnd.n3276 gnd.n3275 585
R2165 gnd.n3275 gnd.n3274 585
R2166 gnd.n1474 gnd.n1473 585
R2167 gnd.n3141 gnd.n1474 585
R2168 gnd.n3256 gnd.n3255 585
R2169 gnd.n3257 gnd.n3256 585
R2170 gnd.n3254 gnd.n1490 585
R2171 gnd.n1490 gnd.n1486 585
R2172 gnd.n3253 gnd.n3252 585
R2173 gnd.n3252 gnd.n3251 585
R2174 gnd.n1492 gnd.n1491 585
R2175 gnd.n3149 gnd.n1492 585
R2176 gnd.n3231 gnd.n3230 585
R2177 gnd.n3232 gnd.n3231 585
R2178 gnd.n3229 gnd.n1504 585
R2179 gnd.n1504 gnd.n1501 585
R2180 gnd.n3228 gnd.n3227 585
R2181 gnd.n3227 gnd.n3226 585
R2182 gnd.n1506 gnd.n1505 585
R2183 gnd.n3157 gnd.n1506 585
R2184 gnd.n3213 gnd.n3212 585
R2185 gnd.n3214 gnd.n3213 585
R2186 gnd.n3211 gnd.n1516 585
R2187 gnd.n3206 gnd.n1516 585
R2188 gnd.n3210 gnd.n3209 585
R2189 gnd.n3209 gnd.n3208 585
R2190 gnd.n1518 gnd.n1517 585
R2191 gnd.n3164 gnd.n1518 585
R2192 gnd.n3182 gnd.n3181 585
R2193 gnd.n3181 gnd.n1530 585
R2194 gnd.n3183 gnd.n1539 585
R2195 gnd.n3169 gnd.n1539 585
R2196 gnd.n3185 gnd.n3184 585
R2197 gnd.n3186 gnd.n3185 585
R2198 gnd.n3180 gnd.n1538 585
R2199 gnd.n3175 gnd.n1538 585
R2200 gnd.n3179 gnd.n3178 585
R2201 gnd.n3178 gnd.n3177 585
R2202 gnd.n1541 gnd.n1540 585
R2203 gnd.n3135 gnd.n1541 585
R2204 gnd.n3121 gnd.n1559 585
R2205 gnd.n1559 gnd.n1558 585
R2206 gnd.n3123 gnd.n3122 585
R2207 gnd.n3124 gnd.n3123 585
R2208 gnd.n3120 gnd.n1557 585
R2209 gnd.n1557 gnd.n1553 585
R2210 gnd.n3119 gnd.n3118 585
R2211 gnd.n3118 gnd.n3117 585
R2212 gnd.n1561 gnd.n1560 585
R2213 gnd.n3055 gnd.n1561 585
R2214 gnd.n3096 gnd.n3095 585
R2215 gnd.n3097 gnd.n3096 585
R2216 gnd.n3094 gnd.n1573 585
R2217 gnd.n1573 gnd.n1570 585
R2218 gnd.n3093 gnd.n3092 585
R2219 gnd.n3092 gnd.n3091 585
R2220 gnd.n1575 gnd.n1574 585
R2221 gnd.n3063 gnd.n1575 585
R2222 gnd.n3078 gnd.n3077 585
R2223 gnd.n3079 gnd.n3078 585
R2224 gnd.n3076 gnd.n1586 585
R2225 gnd.n3069 gnd.n1586 585
R2226 gnd.n3075 gnd.n3074 585
R2227 gnd.n3074 gnd.n3073 585
R2228 gnd.n1588 gnd.n1587 585
R2229 gnd.n3045 gnd.n1588 585
R2230 gnd.n3031 gnd.n3030 585
R2231 gnd.n3030 gnd.n1594 585
R2232 gnd.n3032 gnd.n1603 585
R2233 gnd.n2964 gnd.n1603 585
R2234 gnd.n3034 gnd.n3033 585
R2235 gnd.n3035 gnd.n3034 585
R2236 gnd.n3029 gnd.n1602 585
R2237 gnd.n3024 gnd.n1602 585
R2238 gnd.n3028 gnd.n3027 585
R2239 gnd.n3027 gnd.n3026 585
R2240 gnd.n1605 gnd.n1604 585
R2241 gnd.n1617 gnd.n1605 585
R2242 gnd.n2988 gnd.n2987 585
R2243 gnd.n2987 gnd.n1616 585
R2244 gnd.n2989 gnd.n1627 585
R2245 gnd.n2975 gnd.n1627 585
R2246 gnd.n2991 gnd.n2990 585
R2247 gnd.n2992 gnd.n2991 585
R2248 gnd.n2986 gnd.n1626 585
R2249 gnd.n2981 gnd.n1626 585
R2250 gnd.n2985 gnd.n2984 585
R2251 gnd.n2984 gnd.n2983 585
R2252 gnd.n1629 gnd.n1628 585
R2253 gnd.n2958 gnd.n1629 585
R2254 gnd.n2944 gnd.n1644 585
R2255 gnd.n2922 gnd.n1644 585
R2256 gnd.n2946 gnd.n2945 585
R2257 gnd.n2947 gnd.n2946 585
R2258 gnd.n2943 gnd.n1643 585
R2259 gnd.n2937 gnd.n1643 585
R2260 gnd.n2942 gnd.n2941 585
R2261 gnd.n2941 gnd.n2940 585
R2262 gnd.n1646 gnd.n1645 585
R2263 gnd.n2930 gnd.n1646 585
R2264 gnd.n2906 gnd.n1663 585
R2265 gnd.n1663 gnd.n1662 585
R2266 gnd.n2908 gnd.n2907 585
R2267 gnd.n2909 gnd.n2908 585
R2268 gnd.n2905 gnd.n1660 585
R2269 gnd.n1660 gnd.n1657 585
R2270 gnd.n2904 gnd.n2903 585
R2271 gnd.n2903 gnd.n2902 585
R2272 gnd.n1665 gnd.n1664 585
R2273 gnd.n2769 gnd.n1665 585
R2274 gnd.n2886 gnd.n2885 585
R2275 gnd.n2887 gnd.n2886 585
R2276 gnd.n2884 gnd.n1678 585
R2277 gnd.n2879 gnd.n1678 585
R2278 gnd.n2883 gnd.n2882 585
R2279 gnd.n2882 gnd.n2881 585
R2280 gnd.n1680 gnd.n1679 585
R2281 gnd.n2867 gnd.n1680 585
R2282 gnd.n2854 gnd.n1702 585
R2283 gnd.n1702 gnd.n1690 585
R2284 gnd.n2856 gnd.n2855 585
R2285 gnd.n2857 gnd.n2856 585
R2286 gnd.n2853 gnd.n1701 585
R2287 gnd.n1701 gnd.n1697 585
R2288 gnd.n2852 gnd.n2851 585
R2289 gnd.n2851 gnd.n2850 585
R2290 gnd.n1704 gnd.n1703 585
R2291 gnd.n2783 gnd.n1704 585
R2292 gnd.n2839 gnd.n2838 585
R2293 gnd.n2840 gnd.n2839 585
R2294 gnd.n2837 gnd.n1715 585
R2295 gnd.n1715 gnd.n1712 585
R2296 gnd.n2836 gnd.n2835 585
R2297 gnd.n2835 gnd.n2834 585
R2298 gnd.n1717 gnd.n1716 585
R2299 gnd.n2791 gnd.n1717 585
R2300 gnd.n2821 gnd.n2820 585
R2301 gnd.n2822 gnd.n2821 585
R2302 gnd.n2819 gnd.n1729 585
R2303 gnd.n1733 gnd.n1729 585
R2304 gnd.n2818 gnd.n2817 585
R2305 gnd.n2817 gnd.n2816 585
R2306 gnd.n1731 gnd.n1730 585
R2307 gnd.n2801 gnd.n1731 585
R2308 gnd.n2758 gnd.n1747 585
R2309 gnd.n1747 gnd.n1740 585
R2310 gnd.n2760 gnd.n2759 585
R2311 gnd.n2761 gnd.n2760 585
R2312 gnd.n2756 gnd.n1746 585
R2313 gnd.n2755 gnd.n2754 585
R2314 gnd.n1769 gnd.n1768 585
R2315 gnd.n2752 gnd.n1769 585
R2316 gnd.n2535 gnd.n2534 585
R2317 gnd.n2537 gnd.n2536 585
R2318 gnd.n2539 gnd.n2538 585
R2319 gnd.n2541 gnd.n2540 585
R2320 gnd.n2543 gnd.n2542 585
R2321 gnd.n2545 gnd.n2544 585
R2322 gnd.n2547 gnd.n2546 585
R2323 gnd.n2549 gnd.n2548 585
R2324 gnd.n2551 gnd.n2550 585
R2325 gnd.n2553 gnd.n2552 585
R2326 gnd.n2555 gnd.n2554 585
R2327 gnd.n2557 gnd.n2556 585
R2328 gnd.n2559 gnd.n2558 585
R2329 gnd.n2561 gnd.n2560 585
R2330 gnd.n2563 gnd.n2562 585
R2331 gnd.n2565 gnd.n2564 585
R2332 gnd.n2567 gnd.n2566 585
R2333 gnd.n2569 gnd.n2568 585
R2334 gnd.n2571 gnd.n2570 585
R2335 gnd.n2573 gnd.n2572 585
R2336 gnd.n2575 gnd.n2574 585
R2337 gnd.n2577 gnd.n2576 585
R2338 gnd.n2579 gnd.n2578 585
R2339 gnd.n2581 gnd.n2580 585
R2340 gnd.n2583 gnd.n2582 585
R2341 gnd.n2585 gnd.n2584 585
R2342 gnd.n2587 gnd.n2586 585
R2343 gnd.n2589 gnd.n2588 585
R2344 gnd.n2591 gnd.n2590 585
R2345 gnd.n2595 gnd.n2594 585
R2346 gnd.n2593 gnd.n2530 585
R2347 gnd.n2529 gnd.n2528 585
R2348 gnd.n2527 gnd.n2526 585
R2349 gnd.n2524 gnd.n2523 585
R2350 gnd.n2522 gnd.n2521 585
R2351 gnd.n2520 gnd.n2519 585
R2352 gnd.n2518 gnd.n2517 585
R2353 gnd.n2516 gnd.n2515 585
R2354 gnd.n2514 gnd.n2513 585
R2355 gnd.n2512 gnd.n2511 585
R2356 gnd.n2510 gnd.n2509 585
R2357 gnd.n2508 gnd.n2507 585
R2358 gnd.n2506 gnd.n2505 585
R2359 gnd.n2504 gnd.n2503 585
R2360 gnd.n2502 gnd.n2501 585
R2361 gnd.n2500 gnd.n2499 585
R2362 gnd.n2498 gnd.n2497 585
R2363 gnd.n2496 gnd.n2495 585
R2364 gnd.n2494 gnd.n2493 585
R2365 gnd.n2492 gnd.n2491 585
R2366 gnd.n2490 gnd.n2489 585
R2367 gnd.n2488 gnd.n2487 585
R2368 gnd.n2486 gnd.n2485 585
R2369 gnd.n2484 gnd.n2483 585
R2370 gnd.n2482 gnd.n2481 585
R2371 gnd.n2480 gnd.n2479 585
R2372 gnd.n2478 gnd.n2477 585
R2373 gnd.n2476 gnd.n2475 585
R2374 gnd.n2474 gnd.n2473 585
R2375 gnd.n2472 gnd.n2471 585
R2376 gnd.n2470 gnd.n2469 585
R2377 gnd.n1744 gnd.n1743 585
R2378 gnd.n3631 gnd.n3630 585
R2379 gnd.n3633 gnd.n3632 585
R2380 gnd.n3635 gnd.n3634 585
R2381 gnd.n3637 gnd.n3636 585
R2382 gnd.n3639 gnd.n3638 585
R2383 gnd.n3641 gnd.n3640 585
R2384 gnd.n3643 gnd.n3642 585
R2385 gnd.n3645 gnd.n3644 585
R2386 gnd.n3647 gnd.n3646 585
R2387 gnd.n3649 gnd.n3648 585
R2388 gnd.n3651 gnd.n3650 585
R2389 gnd.n3653 gnd.n3652 585
R2390 gnd.n3655 gnd.n3654 585
R2391 gnd.n3657 gnd.n3656 585
R2392 gnd.n3659 gnd.n3658 585
R2393 gnd.n3661 gnd.n3660 585
R2394 gnd.n3663 gnd.n3662 585
R2395 gnd.n3665 gnd.n3664 585
R2396 gnd.n3667 gnd.n3666 585
R2397 gnd.n3669 gnd.n3668 585
R2398 gnd.n3671 gnd.n3670 585
R2399 gnd.n3673 gnd.n3672 585
R2400 gnd.n3675 gnd.n3674 585
R2401 gnd.n3677 gnd.n3676 585
R2402 gnd.n3679 gnd.n3678 585
R2403 gnd.n3681 gnd.n3680 585
R2404 gnd.n3683 gnd.n3682 585
R2405 gnd.n3685 gnd.n3684 585
R2406 gnd.n3687 gnd.n3686 585
R2407 gnd.n3689 gnd.n1397 585
R2408 gnd.n3691 gnd.n3690 585
R2409 gnd.n3693 gnd.n1361 585
R2410 gnd.n3695 gnd.n3694 585
R2411 gnd.n3698 gnd.n3697 585
R2412 gnd.n1364 gnd.n1362 585
R2413 gnd.n3564 gnd.n3563 585
R2414 gnd.n3566 gnd.n3565 585
R2415 gnd.n3569 gnd.n3568 585
R2416 gnd.n3571 gnd.n3570 585
R2417 gnd.n3573 gnd.n3572 585
R2418 gnd.n3575 gnd.n3574 585
R2419 gnd.n3577 gnd.n3576 585
R2420 gnd.n3579 gnd.n3578 585
R2421 gnd.n3581 gnd.n3580 585
R2422 gnd.n3583 gnd.n3582 585
R2423 gnd.n3585 gnd.n3584 585
R2424 gnd.n3587 gnd.n3586 585
R2425 gnd.n3589 gnd.n3588 585
R2426 gnd.n3591 gnd.n3590 585
R2427 gnd.n3593 gnd.n3592 585
R2428 gnd.n3595 gnd.n3594 585
R2429 gnd.n3597 gnd.n3596 585
R2430 gnd.n3599 gnd.n3598 585
R2431 gnd.n3601 gnd.n3600 585
R2432 gnd.n3603 gnd.n3602 585
R2433 gnd.n3605 gnd.n3604 585
R2434 gnd.n3607 gnd.n3606 585
R2435 gnd.n3609 gnd.n3608 585
R2436 gnd.n3611 gnd.n3610 585
R2437 gnd.n3613 gnd.n3612 585
R2438 gnd.n3615 gnd.n3614 585
R2439 gnd.n3617 gnd.n3616 585
R2440 gnd.n3619 gnd.n3618 585
R2441 gnd.n3621 gnd.n3620 585
R2442 gnd.n3623 gnd.n3622 585
R2443 gnd.n3624 gnd.n1405 585
R2444 gnd.n3629 gnd.n1400 585
R2445 gnd.n3629 gnd.n3628 585
R2446 gnd.n3285 gnd.n1401 585
R2447 gnd.n1411 gnd.n1401 585
R2448 gnd.n3286 gnd.n1409 585
R2449 gnd.n3538 gnd.n1409 585
R2450 gnd.n3288 gnd.n3287 585
R2451 gnd.t161 gnd.n3288 585
R2452 gnd.n3284 gnd.n1466 585
R2453 gnd.n1471 gnd.n1466 585
R2454 gnd.n3283 gnd.n3282 585
R2455 gnd.n3282 gnd.n3281 585
R2456 gnd.n1468 gnd.n1467 585
R2457 gnd.n1478 gnd.n1468 585
R2458 gnd.n3140 gnd.n1477 585
R2459 gnd.n3274 gnd.n1477 585
R2460 gnd.n3143 gnd.n3142 585
R2461 gnd.n3142 gnd.n3141 585
R2462 gnd.n3144 gnd.n1488 585
R2463 gnd.n3257 gnd.n1488 585
R2464 gnd.n3146 gnd.n3145 585
R2465 gnd.n3145 gnd.n1486 585
R2466 gnd.n3147 gnd.n1494 585
R2467 gnd.n3251 gnd.n1494 585
R2468 gnd.n3151 gnd.n3150 585
R2469 gnd.n3150 gnd.n3149 585
R2470 gnd.n3152 gnd.n1502 585
R2471 gnd.n3232 gnd.n1502 585
R2472 gnd.n3154 gnd.n3153 585
R2473 gnd.n3153 gnd.n1501 585
R2474 gnd.n3155 gnd.n1507 585
R2475 gnd.n3226 gnd.n1507 585
R2476 gnd.n3159 gnd.n3158 585
R2477 gnd.n3158 gnd.n3157 585
R2478 gnd.n3160 gnd.n1514 585
R2479 gnd.n3214 gnd.n1514 585
R2480 gnd.n3161 gnd.n1522 585
R2481 gnd.n3206 gnd.n1522 585
R2482 gnd.n3162 gnd.n1521 585
R2483 gnd.n3208 gnd.n1521 585
R2484 gnd.n3165 gnd.n3163 585
R2485 gnd.n3165 gnd.n3164 585
R2486 gnd.n3166 gnd.n3139 585
R2487 gnd.n3166 gnd.n1530 585
R2488 gnd.n3171 gnd.n3170 585
R2489 gnd.n3170 gnd.n3169 585
R2490 gnd.n3172 gnd.n1537 585
R2491 gnd.n3186 gnd.n1537 585
R2492 gnd.n3174 gnd.n3173 585
R2493 gnd.n3175 gnd.n3174 585
R2494 gnd.n3138 gnd.n1544 585
R2495 gnd.n3177 gnd.n1544 585
R2496 gnd.n3137 gnd.n3136 585
R2497 gnd.n3136 gnd.n3135 585
R2498 gnd.n1546 gnd.n1545 585
R2499 gnd.n1558 gnd.n1546 585
R2500 gnd.n3049 gnd.n1555 585
R2501 gnd.n3124 gnd.n1555 585
R2502 gnd.n3051 gnd.n3050 585
R2503 gnd.n3050 gnd.n1553 585
R2504 gnd.n3052 gnd.n1563 585
R2505 gnd.n3117 gnd.n1563 585
R2506 gnd.n3057 gnd.n3056 585
R2507 gnd.n3056 gnd.n3055 585
R2508 gnd.n3058 gnd.n1571 585
R2509 gnd.n3097 gnd.n1571 585
R2510 gnd.n3060 gnd.n3059 585
R2511 gnd.n3059 gnd.n1570 585
R2512 gnd.n3061 gnd.n1577 585
R2513 gnd.n3091 gnd.n1577 585
R2514 gnd.n3065 gnd.n3064 585
R2515 gnd.n3064 gnd.n3063 585
R2516 gnd.n3066 gnd.n1584 585
R2517 gnd.n3079 gnd.n1584 585
R2518 gnd.n3068 gnd.n3067 585
R2519 gnd.n3069 gnd.n3068 585
R2520 gnd.n3048 gnd.n1590 585
R2521 gnd.n3073 gnd.n1590 585
R2522 gnd.n3047 gnd.n3046 585
R2523 gnd.n3046 gnd.n3045 585
R2524 gnd.n1593 gnd.n1592 585
R2525 gnd.n1594 gnd.n1593 585
R2526 gnd.n2966 gnd.n2965 585
R2527 gnd.n2965 gnd.n2964 585
R2528 gnd.n2967 gnd.n1600 585
R2529 gnd.n3035 gnd.n1600 585
R2530 gnd.n2968 gnd.n1608 585
R2531 gnd.n3024 gnd.n1608 585
R2532 gnd.n2969 gnd.n1607 585
R2533 gnd.n3026 gnd.n1607 585
R2534 gnd.n2971 gnd.n2970 585
R2535 gnd.n2971 gnd.n1617 585
R2536 gnd.n2972 gnd.n2962 585
R2537 gnd.n2972 gnd.n1616 585
R2538 gnd.n2977 gnd.n2976 585
R2539 gnd.n2976 gnd.n2975 585
R2540 gnd.n2978 gnd.n1625 585
R2541 gnd.n2992 gnd.n1625 585
R2542 gnd.n2980 gnd.n2979 585
R2543 gnd.n2981 gnd.n2980 585
R2544 gnd.n2961 gnd.n1630 585
R2545 gnd.n2983 gnd.n1630 585
R2546 gnd.n2960 gnd.n2959 585
R2547 gnd.n2959 gnd.n2958 585
R2548 gnd.n1632 gnd.n1631 585
R2549 gnd.n2922 gnd.n1632 585
R2550 gnd.n2934 gnd.n1642 585
R2551 gnd.n2947 gnd.n1642 585
R2552 gnd.n2936 gnd.n2935 585
R2553 gnd.n2937 gnd.n2936 585
R2554 gnd.n2933 gnd.n1647 585
R2555 gnd.n2940 gnd.n1647 585
R2556 gnd.n2932 gnd.n2931 585
R2557 gnd.n2931 gnd.n2930 585
R2558 gnd.n1649 gnd.n1648 585
R2559 gnd.n1662 gnd.n1649 585
R2560 gnd.n2765 gnd.n1658 585
R2561 gnd.n2909 gnd.n1658 585
R2562 gnd.n2767 gnd.n2766 585
R2563 gnd.n2766 gnd.n1657 585
R2564 gnd.n2768 gnd.n1668 585
R2565 gnd.n2902 gnd.n1668 585
R2566 gnd.n2771 gnd.n2770 585
R2567 gnd.n2770 gnd.n2769 585
R2568 gnd.n2772 gnd.n1676 585
R2569 gnd.n2887 gnd.n1676 585
R2570 gnd.n2773 gnd.n1683 585
R2571 gnd.n2879 gnd.n1683 585
R2572 gnd.n2774 gnd.n1682 585
R2573 gnd.n2881 gnd.n1682 585
R2574 gnd.n2775 gnd.n1691 585
R2575 gnd.n2867 gnd.n1691 585
R2576 gnd.n2777 gnd.n2776 585
R2577 gnd.n2776 gnd.n1690 585
R2578 gnd.n2778 gnd.n1698 585
R2579 gnd.n2857 gnd.n1698 585
R2580 gnd.n2780 gnd.n2779 585
R2581 gnd.n2779 gnd.n1697 585
R2582 gnd.n2781 gnd.n1706 585
R2583 gnd.n2850 gnd.n1706 585
R2584 gnd.n2785 gnd.n2784 585
R2585 gnd.n2784 gnd.n2783 585
R2586 gnd.n2786 gnd.n1713 585
R2587 gnd.n2840 gnd.n1713 585
R2588 gnd.n2788 gnd.n2787 585
R2589 gnd.n2787 gnd.n1712 585
R2590 gnd.n2789 gnd.n1719 585
R2591 gnd.n2834 gnd.n1719 585
R2592 gnd.n2793 gnd.n2792 585
R2593 gnd.n2792 gnd.n2791 585
R2594 gnd.n2794 gnd.n1727 585
R2595 gnd.n2822 gnd.n1727 585
R2596 gnd.n2796 gnd.n2795 585
R2597 gnd.n2795 gnd.n1733 585
R2598 gnd.n2797 gnd.n1732 585
R2599 gnd.n2816 gnd.n1732 585
R2600 gnd.n2799 gnd.n2798 585
R2601 gnd.n2801 gnd.n2799 585
R2602 gnd.n2764 gnd.n1742 585
R2603 gnd.n1742 gnd.n1740 585
R2604 gnd.n2763 gnd.n2762 585
R2605 gnd.n2762 gnd.n2761 585
R2606 gnd.n764 gnd.n763 585
R2607 gnd.n957 gnd.n764 585
R2608 gnd.n6559 gnd.n6558 585
R2609 gnd.n6559 gnd.n232 585
R2610 gnd.n6561 gnd.n257 585
R2611 gnd.n6561 gnd.n6560 585
R2612 gnd.n6563 gnd.n6562 585
R2613 gnd.n6562 gnd.n236 585
R2614 gnd.n6564 gnd.n252 585
R2615 gnd.n252 gnd.n246 585
R2616 gnd.n6566 gnd.n6565 585
R2617 gnd.n6567 gnd.n6566 585
R2618 gnd.n253 gnd.n251 585
R2619 gnd.n251 gnd.n248 585
R2620 gnd.n3995 gnd.n3994 585
R2621 gnd.n3994 gnd.n1251 585
R2622 gnd.n3999 gnd.n3993 585
R2623 gnd.n3993 gnd.n1262 585
R2624 gnd.n4000 gnd.n1276 585
R2625 gnd.n1276 gnd.n1260 585
R2626 gnd.n4002 gnd.n4001 585
R2627 gnd.n4003 gnd.n4002 585
R2628 gnd.n1277 gnd.n1275 585
R2629 gnd.n1275 gnd.n1270 585
R2630 gnd.n3988 gnd.n3987 585
R2631 gnd.n3987 gnd.n3986 585
R2632 gnd.n1280 gnd.n1279 585
R2633 gnd.n1291 gnd.n1280 585
R2634 gnd.n3961 gnd.n1304 585
R2635 gnd.n1304 gnd.n1289 585
R2636 gnd.n3963 gnd.n3962 585
R2637 gnd.n3964 gnd.n3963 585
R2638 gnd.n1305 gnd.n1303 585
R2639 gnd.n1303 gnd.n1299 585
R2640 gnd.n3956 gnd.n3955 585
R2641 gnd.n3955 gnd.n3954 585
R2642 gnd.n1308 gnd.n1307 585
R2643 gnd.n1320 gnd.n1308 585
R2644 gnd.n3930 gnd.n3918 585
R2645 gnd.n3918 gnd.n1318 585
R2646 gnd.n3932 gnd.n3931 585
R2647 gnd.n3933 gnd.n3932 585
R2648 gnd.n3919 gnd.n3917 585
R2649 gnd.n3917 gnd.n1325 585
R2650 gnd.n3925 gnd.n3924 585
R2651 gnd.n3924 gnd.n1227 585
R2652 gnd.n3923 gnd.n3922 585
R2653 gnd.n3923 gnd.n1224 585
R2654 gnd.n1211 gnd.n1210 585
R2655 gnd.n1215 gnd.n1211 585
R2656 gnd.n4057 gnd.n4056 585
R2657 gnd.n4056 gnd.n4055 585
R2658 gnd.n4058 gnd.n1205 585
R2659 gnd.n1212 gnd.n1205 585
R2660 gnd.n4060 gnd.n4059 585
R2661 gnd.n4061 gnd.n4060 585
R2662 gnd.n1202 gnd.n1201 585
R2663 gnd.n4062 gnd.n1202 585
R2664 gnd.n4065 gnd.n4064 585
R2665 gnd.n4064 gnd.n4063 585
R2666 gnd.n4066 gnd.n1196 585
R2667 gnd.n1196 gnd.n1194 585
R2668 gnd.n4068 gnd.n4067 585
R2669 gnd.n4069 gnd.n4068 585
R2670 gnd.n1197 gnd.n1195 585
R2671 gnd.n1195 gnd.n1192 585
R2672 gnd.n3499 gnd.n3494 585
R2673 gnd.n3494 gnd.n3493 585
R2674 gnd.n3501 gnd.n3500 585
R2675 gnd.n3502 gnd.n3501 585
R2676 gnd.n1440 gnd.n1439 585
R2677 gnd.n3505 gnd.n1440 585
R2678 gnd.n3509 gnd.n3508 585
R2679 gnd.n3508 gnd.n3507 585
R2680 gnd.n3510 gnd.n1434 585
R2681 gnd.n1450 gnd.n1434 585
R2682 gnd.n3512 gnd.n3511 585
R2683 gnd.n3513 gnd.n3512 585
R2684 gnd.n1429 gnd.n1428 585
R2685 gnd.n3516 gnd.n1429 585
R2686 gnd.n3520 gnd.n3519 585
R2687 gnd.n3519 gnd.n3518 585
R2688 gnd.n3521 gnd.n1423 585
R2689 gnd.n1430 gnd.n1423 585
R2690 gnd.n3523 gnd.n3522 585
R2691 gnd.n3524 gnd.n3523 585
R2692 gnd.n1419 gnd.n1418 585
R2693 gnd.n3527 gnd.n1419 585
R2694 gnd.n3531 gnd.n3530 585
R2695 gnd.n3530 gnd.n3529 585
R2696 gnd.n3532 gnd.n1413 585
R2697 gnd.n1413 gnd.n1403 585
R2698 gnd.n3534 gnd.n3533 585
R2699 gnd.n3535 gnd.n3534 585
R2700 gnd.n1414 gnd.n1412 585
R2701 gnd.n1412 gnd.n1408 585
R2702 gnd.n3269 gnd.n3268 585
R2703 gnd.n3268 gnd.n1465 585
R2704 gnd.n3270 gnd.n1481 585
R2705 gnd.n1481 gnd.t189 585
R2706 gnd.n3272 gnd.n3271 585
R2707 gnd.n3273 gnd.n3272 585
R2708 gnd.n1482 gnd.n1480 585
R2709 gnd.n1489 gnd.n1480 585
R2710 gnd.n3261 gnd.n3260 585
R2711 gnd.n3260 gnd.n3259 585
R2712 gnd.n1485 gnd.n1484 585
R2713 gnd.n1493 gnd.n1485 585
R2714 gnd.n3222 gnd.n1509 585
R2715 gnd.n1509 gnd.n1503 585
R2716 gnd.n3224 gnd.n3223 585
R2717 gnd.n3225 gnd.n3224 585
R2718 gnd.n1510 gnd.n1508 585
R2719 gnd.n3156 gnd.n1508 585
R2720 gnd.n3217 gnd.n3216 585
R2721 gnd.n3216 gnd.n3215 585
R2722 gnd.n1513 gnd.n1512 585
R2723 gnd.n3207 gnd.n1513 585
R2724 gnd.n3194 gnd.n3193 585
R2725 gnd.n3195 gnd.n3194 585
R2726 gnd.n1532 gnd.n1531 585
R2727 gnd.n3168 gnd.n1531 585
R2728 gnd.n3189 gnd.n3188 585
R2729 gnd.n3188 gnd.n3187 585
R2730 gnd.n1535 gnd.n1534 585
R2731 gnd.n3176 gnd.n1535 585
R2732 gnd.n3133 gnd.n3132 585
R2733 gnd.n3134 gnd.n3133 585
R2734 gnd.n1549 gnd.n1548 585
R2735 gnd.n1556 gnd.n1548 585
R2736 gnd.n3128 gnd.n3127 585
R2737 gnd.n3127 gnd.n3126 585
R2738 gnd.n1552 gnd.n1551 585
R2739 gnd.n1562 gnd.n1552 585
R2740 gnd.n3087 gnd.n1579 585
R2741 gnd.n1579 gnd.n1572 585
R2742 gnd.n3089 gnd.n3088 585
R2743 gnd.n3090 gnd.n3089 585
R2744 gnd.n1580 gnd.n1578 585
R2745 gnd.n3062 gnd.n1578 585
R2746 gnd.n3082 gnd.n3081 585
R2747 gnd.n3081 gnd.n3080 585
R2748 gnd.n1583 gnd.n1582 585
R2749 gnd.n3072 gnd.n1583 585
R2750 gnd.n3043 gnd.n3042 585
R2751 gnd.n3044 gnd.n3043 585
R2752 gnd.n1596 gnd.n1595 585
R2753 gnd.n2963 gnd.n1595 585
R2754 gnd.n3038 gnd.n3037 585
R2755 gnd.n3037 gnd.n3036 585
R2756 gnd.n1599 gnd.n1598 585
R2757 gnd.n3025 gnd.n1599 585
R2758 gnd.n3000 gnd.n2999 585
R2759 gnd.n3001 gnd.n3000 585
R2760 gnd.n1619 gnd.n1618 585
R2761 gnd.n2974 gnd.n1618 585
R2762 gnd.n2995 gnd.n2994 585
R2763 gnd.n2994 gnd.n2993 585
R2764 gnd.n1622 gnd.n1621 585
R2765 gnd.n2982 gnd.n1622 585
R2766 gnd.n2920 gnd.n2919 585
R2767 gnd.n2920 gnd.n1633 585
R2768 gnd.n2925 gnd.n2924 585
R2769 gnd.n2924 gnd.n2923 585
R2770 gnd.n2926 gnd.n1652 585
R2771 gnd.n1652 gnd.n1641 585
R2772 gnd.n2928 gnd.n2927 585
R2773 gnd.n2929 gnd.n2928 585
R2774 gnd.n1653 gnd.n1651 585
R2775 gnd.n1661 gnd.n1651 585
R2776 gnd.n2912 gnd.n2911 585
R2777 gnd.n2911 gnd.n2910 585
R2778 gnd.n1656 gnd.n1655 585
R2779 gnd.n2901 gnd.n1656 585
R2780 gnd.n2875 gnd.n1685 585
R2781 gnd.n1685 gnd.n1677 585
R2782 gnd.n2877 gnd.n2876 585
R2783 gnd.n2878 gnd.n2877 585
R2784 gnd.n1686 gnd.n1684 585
R2785 gnd.n1684 gnd.n1681 585
R2786 gnd.n2870 gnd.n2869 585
R2787 gnd.n2869 gnd.n2868 585
R2788 gnd.n1689 gnd.n1688 585
R2789 gnd.n2858 gnd.n1689 585
R2790 gnd.n2848 gnd.n2847 585
R2791 gnd.n2849 gnd.n2848 585
R2792 gnd.n1708 gnd.n1707 585
R2793 gnd.n2782 gnd.n1707 585
R2794 gnd.n2843 gnd.n2842 585
R2795 gnd.n2842 gnd.n2841 585
R2796 gnd.n1711 gnd.n1710 585
R2797 gnd.n1718 gnd.n1711 585
R2798 gnd.n2811 gnd.n1735 585
R2799 gnd.n1735 gnd.n1728 585
R2800 gnd.n2813 gnd.n2812 585
R2801 gnd.n2814 gnd.n2813 585
R2802 gnd.n1736 gnd.n1734 585
R2803 gnd.n2800 gnd.n1734 585
R2804 gnd.n2806 gnd.n2805 585
R2805 gnd.n2805 gnd.n2804 585
R2806 gnd.n1739 gnd.n1738 585
R2807 gnd.n2750 gnd.n1739 585
R2808 gnd.n2734 gnd.n1812 585
R2809 gnd.n1812 gnd.n1770 585
R2810 gnd.n2736 gnd.n2735 585
R2811 gnd.n2737 gnd.n2736 585
R2812 gnd.n1813 gnd.n1811 585
R2813 gnd.n2725 gnd.n1811 585
R2814 gnd.n2729 gnd.n2728 585
R2815 gnd.n2728 gnd.n2727 585
R2816 gnd.n1816 gnd.n1815 585
R2817 gnd.n1817 gnd.n1816 585
R2818 gnd.n2713 gnd.n2712 585
R2819 gnd.n2714 gnd.n2713 585
R2820 gnd.n1826 gnd.n1825 585
R2821 gnd.n1825 gnd.n1823 585
R2822 gnd.n2708 gnd.n2707 585
R2823 gnd.n2707 gnd.n2706 585
R2824 gnd.n1829 gnd.n1828 585
R2825 gnd.n1830 gnd.n1829 585
R2826 gnd.n2693 gnd.n2692 585
R2827 gnd.n2694 gnd.n2693 585
R2828 gnd.n1839 gnd.n1838 585
R2829 gnd.n1838 gnd.n1836 585
R2830 gnd.n2688 gnd.n2687 585
R2831 gnd.n2687 gnd.n2686 585
R2832 gnd.n1842 gnd.n1841 585
R2833 gnd.n1843 gnd.n1842 585
R2834 gnd.n2338 gnd.n2334 585
R2835 gnd.n2334 gnd.n2333 585
R2836 gnd.n2340 gnd.n2339 585
R2837 gnd.n2340 gnd.n1862 585
R2838 gnd.n2341 gnd.n2331 585
R2839 gnd.n2341 gnd.n1849 585
R2840 gnd.n2344 gnd.n2343 585
R2841 gnd.n2343 gnd.n2342 585
R2842 gnd.n2345 gnd.n2326 585
R2843 gnd.n2326 gnd.n1934 585
R2844 gnd.n2347 gnd.n2346 585
R2845 gnd.n2347 gnd.n1918 585
R2846 gnd.n2348 gnd.n2325 585
R2847 gnd.n2348 gnd.n1082 585
R2848 gnd.n2350 gnd.n2349 585
R2849 gnd.n2349 gnd.n1079 585
R2850 gnd.n2351 gnd.n2320 585
R2851 gnd.n2320 gnd.n1072 585
R2852 gnd.n2353 gnd.n2352 585
R2853 gnd.n2353 gnd.n1069 585
R2854 gnd.n2354 gnd.n2319 585
R2855 gnd.n2354 gnd.n1061 585
R2856 gnd.n2356 gnd.n2355 585
R2857 gnd.n2355 gnd.n1058 585
R2858 gnd.n2357 gnd.n2012 585
R2859 gnd.n2012 gnd.n1050 585
R2860 gnd.n2359 gnd.n2358 585
R2861 gnd.n2360 gnd.n2359 585
R2862 gnd.n2013 gnd.n2011 585
R2863 gnd.n2011 gnd.n1040 585
R2864 gnd.n2313 gnd.n2312 585
R2865 gnd.n2312 gnd.n1037 585
R2866 gnd.n2311 gnd.n2015 585
R2867 gnd.n2311 gnd.n1029 585
R2868 gnd.n2310 gnd.n2309 585
R2869 gnd.n2310 gnd.n1026 585
R2870 gnd.n2017 gnd.n2016 585
R2871 gnd.n2273 gnd.n2016 585
R2872 gnd.n2305 gnd.n2304 585
R2873 gnd.n2304 gnd.n1016 585
R2874 gnd.n2303 gnd.n2019 585
R2875 gnd.n2303 gnd.n1008 585
R2876 gnd.n2302 gnd.n2021 585
R2877 gnd.n2302 gnd.n2301 585
R2878 gnd.n2058 gnd.n2020 585
R2879 gnd.n2020 gnd.n998 585
R2880 gnd.n2060 gnd.n2059 585
R2881 gnd.n2060 gnd.n995 585
R2882 gnd.n2062 gnd.n2061 585
R2883 gnd.n2061 gnd.n990 585
R2884 gnd.n2063 gnd.n2040 585
R2885 gnd.n2040 gnd.n987 585
R2886 gnd.n2065 gnd.n2064 585
R2887 gnd.n2066 gnd.n2065 585
R2888 gnd.n2041 gnd.n2039 585
R2889 gnd.n2039 gnd.n978 585
R2890 gnd.n2048 gnd.n2047 585
R2891 gnd.n2047 gnd.n973 585
R2892 gnd.n2046 gnd.n2044 585
R2893 gnd.n2046 gnd.n2045 585
R2894 gnd.n4072 gnd.n4071 585
R2895 gnd.n4071 gnd.n4070 585
R2896 gnd.n4073 gnd.n1189 585
R2897 gnd.n3492 gnd.n1189 585
R2898 gnd.n4074 gnd.n1188 585
R2899 gnd.n1444 gnd.n1188 585
R2900 gnd.n3503 gnd.n1186 585
R2901 gnd.n3504 gnd.n3503 585
R2902 gnd.n4078 gnd.n1185 585
R2903 gnd.n3506 gnd.n1185 585
R2904 gnd.n4079 gnd.n1184 585
R2905 gnd.n1441 gnd.n1184 585
R2906 gnd.n4080 gnd.n1183 585
R2907 gnd.n1451 gnd.n1183 585
R2908 gnd.n3514 gnd.n1181 585
R2909 gnd.n3515 gnd.n3514 585
R2910 gnd.n4084 gnd.n1180 585
R2911 gnd.n3517 gnd.n1180 585
R2912 gnd.n4085 gnd.n1179 585
R2913 gnd.n1431 gnd.n1179 585
R2914 gnd.n4086 gnd.n1178 585
R2915 gnd.n1422 gnd.n1178 585
R2916 gnd.n3525 gnd.n1176 585
R2917 gnd.n3526 gnd.n3525 585
R2918 gnd.n4090 gnd.n1175 585
R2919 gnd.n3528 gnd.n1175 585
R2920 gnd.n4091 gnd.n1174 585
R2921 gnd.n1365 gnd.n1174 585
R2922 gnd.n4092 gnd.n1173 585
R2923 gnd.n1402 gnd.n1173 585
R2924 gnd.n3536 gnd.n1171 585
R2925 gnd.n3537 gnd.n3536 585
R2926 gnd.n4096 gnd.n1170 585
R2927 gnd.n3289 gnd.n1170 585
R2928 gnd.n4097 gnd.n1169 585
R2929 gnd.n1469 gnd.n1169 585
R2930 gnd.n4098 gnd.n1168 585
R2931 gnd.n1479 gnd.n1168 585
R2932 gnd.n1475 gnd.n1166 585
R2933 gnd.n1476 gnd.n1475 585
R2934 gnd.n4102 gnd.n1165 585
R2935 gnd.n3258 gnd.n1165 585
R2936 gnd.n4103 gnd.n1164 585
R2937 gnd.n3250 gnd.n1164 585
R2938 gnd.n4104 gnd.n1163 585
R2939 gnd.n3148 gnd.n1163 585
R2940 gnd.n3233 gnd.n1161 585
R2941 gnd.n3234 gnd.n3233 585
R2942 gnd.n4108 gnd.n1160 585
R2943 gnd.n3226 gnd.n1160 585
R2944 gnd.n4109 gnd.n1159 585
R2945 gnd.n1515 gnd.n1159 585
R2946 gnd.n4110 gnd.n1158 585
R2947 gnd.n3205 gnd.n1158 585
R2948 gnd.n1519 gnd.n1156 585
R2949 gnd.n1520 gnd.n1519 585
R2950 gnd.n4114 gnd.n1155 585
R2951 gnd.n3196 gnd.n1155 585
R2952 gnd.n4115 gnd.n1154 585
R2953 gnd.n3167 gnd.n1154 585
R2954 gnd.n4116 gnd.n1153 585
R2955 gnd.n1536 gnd.n1153 585
R2956 gnd.n1542 gnd.n1151 585
R2957 gnd.n1543 gnd.n1542 585
R2958 gnd.n4120 gnd.n1150 585
R2959 gnd.n1547 gnd.n1150 585
R2960 gnd.n4121 gnd.n1149 585
R2961 gnd.n3125 gnd.n1149 585
R2962 gnd.n4122 gnd.n1148 585
R2963 gnd.n3116 gnd.n1148 585
R2964 gnd.n3053 gnd.n1146 585
R2965 gnd.n3054 gnd.n3053 585
R2966 gnd.n4126 gnd.n1145 585
R2967 gnd.n3098 gnd.n1145 585
R2968 gnd.n4127 gnd.n1144 585
R2969 gnd.n1576 gnd.n1144 585
R2970 gnd.n4128 gnd.n1143 585
R2971 gnd.n1585 gnd.n1143 585
R2972 gnd.n3070 gnd.n1141 585
R2973 gnd.n3071 gnd.n3070 585
R2974 gnd.n4132 gnd.n1140 585
R2975 gnd.n1589 gnd.n1140 585
R2976 gnd.n4133 gnd.n1139 585
R2977 gnd.n1594 gnd.n1139 585
R2978 gnd.n4134 gnd.n1138 585
R2979 gnd.n1601 gnd.n1138 585
R2980 gnd.n3022 gnd.n1136 585
R2981 gnd.n3023 gnd.n3022 585
R2982 gnd.n4138 gnd.n1135 585
R2983 gnd.n1606 gnd.n1135 585
R2984 gnd.n4139 gnd.n1134 585
R2985 gnd.n3002 gnd.n1134 585
R2986 gnd.n4140 gnd.n1133 585
R2987 gnd.n2973 gnd.n1133 585
R2988 gnd.n1623 gnd.n1131 585
R2989 gnd.n1624 gnd.n1623 585
R2990 gnd.n4144 gnd.n1130 585
R2991 gnd.n2957 gnd.n1130 585
R2992 gnd.n4145 gnd.n1129 585
R2993 gnd.n2921 gnd.n1129 585
R2994 gnd.n4146 gnd.n1128 585
R2995 gnd.n2948 gnd.n1128 585
R2996 gnd.n2938 gnd.n1126 585
R2997 gnd.n2939 gnd.n2938 585
R2998 gnd.n4150 gnd.n1125 585
R2999 gnd.n1650 gnd.n1125 585
R3000 gnd.n4151 gnd.n1124 585
R3001 gnd.n1659 gnd.n1124 585
R3002 gnd.n4152 gnd.n1123 585
R3003 gnd.n2900 gnd.n1123 585
R3004 gnd.n1666 gnd.n1121 585
R3005 gnd.n1667 gnd.n1666 585
R3006 gnd.n4156 gnd.n1120 585
R3007 gnd.n2888 gnd.n1120 585
R3008 gnd.n4157 gnd.n1119 585
R3009 gnd.n2880 gnd.n1119 585
R3010 gnd.n4158 gnd.n1118 585
R3011 gnd.n2867 gnd.n1118 585
R3012 gnd.n1699 gnd.n1116 585
R3013 gnd.n1700 gnd.n1699 585
R3014 gnd.n4162 gnd.n1115 585
R3015 gnd.n2859 gnd.n1115 585
R3016 gnd.n4163 gnd.n1114 585
R3017 gnd.n1705 gnd.n1114 585
R3018 gnd.n4164 gnd.n1113 585
R3019 gnd.n1714 gnd.n1113 585
R3020 gnd.n2832 gnd.n1111 585
R3021 gnd.n2833 gnd.n2832 585
R3022 gnd.n4168 gnd.n1110 585
R3023 gnd.n2790 gnd.n1110 585
R3024 gnd.n4169 gnd.n1109 585
R3025 gnd.n2823 gnd.n1109 585
R3026 gnd.n4170 gnd.n1108 585
R3027 gnd.n2815 gnd.n1108 585
R3028 gnd.n2802 gnd.n1106 585
R3029 gnd.n2803 gnd.n2802 585
R3030 gnd.n4174 gnd.n1105 585
R3031 gnd.n1745 gnd.n1105 585
R3032 gnd.n4175 gnd.n1104 585
R3033 gnd.n2751 gnd.n1104 585
R3034 gnd.n4176 gnd.n1103 585
R3035 gnd.n1810 gnd.n1103 585
R3036 gnd.n2738 gnd.n1101 585
R3037 gnd.n2739 gnd.n2738 585
R3038 gnd.n4180 gnd.n1100 585
R3039 gnd.n2726 gnd.n1100 585
R3040 gnd.n4181 gnd.n1099 585
R3041 gnd.n2724 gnd.n1099 585
R3042 gnd.n4182 gnd.n1098 585
R3043 gnd.n1824 gnd.n1098 585
R3044 gnd.n2715 gnd.n1096 585
R3045 gnd.n2716 gnd.n2715 585
R3046 gnd.n4186 gnd.n1095 585
R3047 gnd.n2705 gnd.n1095 585
R3048 gnd.n4187 gnd.n1094 585
R3049 gnd.n2704 gnd.n1094 585
R3050 gnd.n4188 gnd.n1093 585
R3051 gnd.n1837 gnd.n1093 585
R3052 gnd.n2695 gnd.n1091 585
R3053 gnd.n2696 gnd.n2695 585
R3054 gnd.n4192 gnd.n1090 585
R3055 gnd.n2685 gnd.n1090 585
R3056 gnd.n4193 gnd.n1089 585
R3057 gnd.n2684 gnd.n1089 585
R3058 gnd.n4194 gnd.n1088 585
R3059 gnd.n2332 gnd.n1088 585
R3060 gnd.n2673 gnd.n2672 585
R3061 gnd.n2671 gnd.n1864 585
R3062 gnd.n1866 gnd.n1863 585
R3063 gnd.n2675 gnd.n1863 585
R3064 gnd.n2664 gnd.n1874 585
R3065 gnd.n2663 gnd.n1875 585
R3066 gnd.n1877 gnd.n1876 585
R3067 gnd.n2656 gnd.n1883 585
R3068 gnd.n2655 gnd.n1884 585
R3069 gnd.n1891 gnd.n1885 585
R3070 gnd.n2648 gnd.n1892 585
R3071 gnd.n2647 gnd.n1893 585
R3072 gnd.n1895 gnd.n1894 585
R3073 gnd.n2640 gnd.n1901 585
R3074 gnd.n2639 gnd.n1902 585
R3075 gnd.n1911 gnd.n1903 585
R3076 gnd.n2632 gnd.n1912 585
R3077 gnd.n2631 gnd.n1913 585
R3078 gnd.n1915 gnd.n1914 585
R3079 gnd.n2411 gnd.n2384 585
R3080 gnd.n2410 gnd.n2385 585
R3081 gnd.n2409 gnd.n2386 585
R3082 gnd.n2388 gnd.n2387 585
R3083 gnd.n2405 gnd.n2390 585
R3084 gnd.n2404 gnd.n2391 585
R3085 gnd.n2403 gnd.n2392 585
R3086 gnd.n2400 gnd.n2397 585
R3087 gnd.n2399 gnd.n2398 585
R3088 gnd.n1848 gnd.n1847 585
R3089 gnd.n2678 gnd.n2677 585
R3090 gnd.n1447 gnd.n1193 585
R3091 gnd.n4070 gnd.n1193 585
R3092 gnd.n3491 gnd.n3490 585
R3093 gnd.n3492 gnd.n3491 585
R3094 gnd.n1446 gnd.n1445 585
R3095 gnd.n1445 gnd.n1444 585
R3096 gnd.n3310 gnd.n1443 585
R3097 gnd.n3504 gnd.n1443 585
R3098 gnd.n3309 gnd.n1442 585
R3099 gnd.n3506 gnd.n1442 585
R3100 gnd.n3308 gnd.n1453 585
R3101 gnd.n1453 gnd.n1441 585
R3102 gnd.n1452 gnd.n1449 585
R3103 gnd.n1452 gnd.n1451 585
R3104 gnd.n3304 gnd.n1433 585
R3105 gnd.n3515 gnd.n1433 585
R3106 gnd.n3303 gnd.n1432 585
R3107 gnd.n3517 gnd.n1432 585
R3108 gnd.n3302 gnd.n1457 585
R3109 gnd.n1457 gnd.n1431 585
R3110 gnd.n1456 gnd.n1455 585
R3111 gnd.n1456 gnd.n1422 585
R3112 gnd.n3298 gnd.n1421 585
R3113 gnd.n3526 gnd.n1421 585
R3114 gnd.n3297 gnd.n1420 585
R3115 gnd.n3528 gnd.n1420 585
R3116 gnd.n3296 gnd.n1461 585
R3117 gnd.n1461 gnd.n1365 585
R3118 gnd.n1460 gnd.n1459 585
R3119 gnd.n1460 gnd.n1402 585
R3120 gnd.n3292 gnd.n1410 585
R3121 gnd.n3537 gnd.n1410 585
R3122 gnd.n3291 gnd.n3290 585
R3123 gnd.n3290 gnd.n3289 585
R3124 gnd.n1464 gnd.n1463 585
R3125 gnd.n1469 gnd.n1464 585
R3126 gnd.n3243 gnd.n3242 585
R3127 gnd.n3242 gnd.n1479 585
R3128 gnd.n3244 gnd.n3241 585
R3129 gnd.n3241 gnd.n1476 585
R3130 gnd.n1497 gnd.n1487 585
R3131 gnd.n3258 gnd.n1487 585
R3132 gnd.n3249 gnd.n3248 585
R3133 gnd.n3250 gnd.n3249 585
R3134 gnd.n1496 gnd.n1495 585
R3135 gnd.n3148 gnd.n1495 585
R3136 gnd.n3236 gnd.n3235 585
R3137 gnd.n3235 gnd.n3234 585
R3138 gnd.n1500 gnd.n1499 585
R3139 gnd.n3226 gnd.n1500 585
R3140 gnd.n1526 gnd.n1524 585
R3141 gnd.n1524 gnd.n1515 585
R3142 gnd.n3204 gnd.n3203 585
R3143 gnd.n3205 gnd.n3204 585
R3144 gnd.n1525 gnd.n1523 585
R3145 gnd.n1523 gnd.n1520 585
R3146 gnd.n3198 gnd.n3197 585
R3147 gnd.n3197 gnd.n3196 585
R3148 gnd.n1529 gnd.n1528 585
R3149 gnd.n3167 gnd.n1529 585
R3150 gnd.n3108 gnd.n3106 585
R3151 gnd.n3106 gnd.n1536 585
R3152 gnd.n3109 gnd.n3105 585
R3153 gnd.n3105 gnd.n1543 585
R3154 gnd.n3110 gnd.n3104 585
R3155 gnd.n3104 gnd.n1547 585
R3156 gnd.n1566 gnd.n1554 585
R3157 gnd.n3125 gnd.n1554 585
R3158 gnd.n3115 gnd.n3114 585
R3159 gnd.n3116 gnd.n3115 585
R3160 gnd.n1565 gnd.n1564 585
R3161 gnd.n3054 gnd.n1564 585
R3162 gnd.n3100 gnd.n3099 585
R3163 gnd.n3099 gnd.n3098 585
R3164 gnd.n1569 gnd.n1568 585
R3165 gnd.n1576 gnd.n1569 585
R3166 gnd.n3011 gnd.n3010 585
R3167 gnd.n3010 gnd.n1585 585
R3168 gnd.n3014 gnd.n1591 585
R3169 gnd.n3071 gnd.n1591 585
R3170 gnd.n3015 gnd.n3009 585
R3171 gnd.n3009 gnd.n1589 585
R3172 gnd.n3016 gnd.n3008 585
R3173 gnd.n3008 gnd.n1594 585
R3174 gnd.n1612 gnd.n1610 585
R3175 gnd.n1610 gnd.n1601 585
R3176 gnd.n3021 gnd.n3020 585
R3177 gnd.n3023 gnd.n3021 585
R3178 gnd.n1611 gnd.n1609 585
R3179 gnd.n1609 gnd.n1606 585
R3180 gnd.n3004 gnd.n3003 585
R3181 gnd.n3003 gnd.n3002 585
R3182 gnd.n1615 gnd.n1614 585
R3183 gnd.n2973 gnd.n1615 585
R3184 gnd.n1637 gnd.n1635 585
R3185 gnd.n1635 gnd.n1624 585
R3186 gnd.n2956 gnd.n2955 585
R3187 gnd.n2957 gnd.n2956 585
R3188 gnd.n1636 gnd.n1634 585
R3189 gnd.n2921 gnd.n1634 585
R3190 gnd.n2950 gnd.n2949 585
R3191 gnd.n2949 gnd.n2948 585
R3192 gnd.n1640 gnd.n1639 585
R3193 gnd.n2939 gnd.n1640 585
R3194 gnd.n2894 gnd.n2893 585
R3195 gnd.n2893 gnd.n1650 585
R3196 gnd.n1672 gnd.n1670 585
R3197 gnd.n1670 gnd.n1659 585
R3198 gnd.n2899 gnd.n2898 585
R3199 gnd.n2900 gnd.n2899 585
R3200 gnd.n1671 gnd.n1669 585
R3201 gnd.n1669 gnd.n1667 585
R3202 gnd.n2890 gnd.n2889 585
R3203 gnd.n2889 gnd.n2888 585
R3204 gnd.n1675 gnd.n1674 585
R3205 gnd.n2880 gnd.n1675 585
R3206 gnd.n2866 gnd.n2865 585
R3207 gnd.n2867 gnd.n2866 585
R3208 gnd.n1693 gnd.n1692 585
R3209 gnd.n1700 gnd.n1692 585
R3210 gnd.n2861 gnd.n2860 585
R3211 gnd.n2860 gnd.n2859 585
R3212 gnd.n1696 gnd.n1695 585
R3213 gnd.n1705 gnd.n1696 585
R3214 gnd.n1723 gnd.n1721 585
R3215 gnd.n1721 gnd.n1714 585
R3216 gnd.n2831 gnd.n2830 585
R3217 gnd.n2833 gnd.n2831 585
R3218 gnd.n1722 gnd.n1720 585
R3219 gnd.n2790 gnd.n1720 585
R3220 gnd.n2825 gnd.n2824 585
R3221 gnd.n2824 gnd.n2823 585
R3222 gnd.n1726 gnd.n1725 585
R3223 gnd.n2815 gnd.n1726 585
R3224 gnd.n2744 gnd.n1741 585
R3225 gnd.n2803 gnd.n1741 585
R3226 gnd.n1806 gnd.n1804 585
R3227 gnd.n1804 gnd.n1745 585
R3228 gnd.n2749 gnd.n2748 585
R3229 gnd.n2751 gnd.n2749 585
R3230 gnd.n1805 gnd.n1803 585
R3231 gnd.n1810 gnd.n1803 585
R3232 gnd.n2741 gnd.n2740 585
R3233 gnd.n2740 gnd.n2739 585
R3234 gnd.n1809 gnd.n1808 585
R3235 gnd.n2726 gnd.n1809 585
R3236 gnd.n2723 gnd.n2722 585
R3237 gnd.n2724 gnd.n2723 585
R3238 gnd.n1819 gnd.n1818 585
R3239 gnd.n1824 gnd.n1818 585
R3240 gnd.n2718 gnd.n2717 585
R3241 gnd.n2717 gnd.n2716 585
R3242 gnd.n1822 gnd.n1821 585
R3243 gnd.n2705 gnd.n1822 585
R3244 gnd.n2703 gnd.n2702 585
R3245 gnd.n2704 gnd.n2703 585
R3246 gnd.n1832 gnd.n1831 585
R3247 gnd.n1837 gnd.n1831 585
R3248 gnd.n2698 gnd.n2697 585
R3249 gnd.n2697 gnd.n2696 585
R3250 gnd.n1835 gnd.n1834 585
R3251 gnd.n2685 gnd.n1835 585
R3252 gnd.n2683 gnd.n2682 585
R3253 gnd.n2684 gnd.n2683 585
R3254 gnd.n1845 gnd.n1844 585
R3255 gnd.n2332 gnd.n1844 585
R3256 gnd.n3486 gnd.n3485 585
R3257 gnd.n3485 gnd.n1203 585
R3258 gnd.n3484 gnd.n3314 585
R3259 gnd.n3482 gnd.n3481 585
R3260 gnd.n3316 gnd.n3315 585
R3261 gnd.n3477 gnd.n3473 585
R3262 gnd.n3471 gnd.n3318 585
R3263 gnd.n3469 gnd.n3468 585
R3264 gnd.n3320 gnd.n3319 585
R3265 gnd.n3464 gnd.n3463 585
R3266 gnd.n3461 gnd.n3322 585
R3267 gnd.n3459 gnd.n3458 585
R3268 gnd.n3324 gnd.n3323 585
R3269 gnd.n3444 gnd.n3443 585
R3270 gnd.n3445 gnd.n3441 585
R3271 gnd.n3439 gnd.n3333 585
R3272 gnd.n3438 gnd.n3437 585
R3273 gnd.n3422 gnd.n3335 585
R3274 gnd.n3424 gnd.n3423 585
R3275 gnd.n3420 gnd.n3342 585
R3276 gnd.n3419 gnd.n3418 585
R3277 gnd.n3403 gnd.n3344 585
R3278 gnd.n3405 gnd.n3404 585
R3279 gnd.n3401 gnd.n3351 585
R3280 gnd.n3400 gnd.n3399 585
R3281 gnd.n3384 gnd.n3353 585
R3282 gnd.n3386 gnd.n3385 585
R3283 gnd.n3382 gnd.n3360 585
R3284 gnd.n3381 gnd.n3380 585
R3285 gnd.n3362 gnd.n1191 585
R3286 gnd.n2467 gnd.t191 543.808
R3287 gnd.n1398 gnd.t183 543.808
R3288 gnd.n2531 gnd.t141 543.808
R3289 gnd.n3561 gnd.t137 543.808
R3290 gnd.n3627 gnd.n1405 458.866
R3291 gnd.n3630 gnd.n3629 458.866
R3292 gnd.n2762 gnd.n1744 458.866
R3293 gnd.n2760 gnd.n1746 458.866
R3294 gnd.n5989 gnd.n5988 422.406
R3295 gnd.n2393 gnd.t163 371.625
R3296 gnd.n6676 gnd.t148 371.625
R3297 gnd.n3326 gnd.t126 371.625
R3298 gnd.n1907 gnd.t157 371.625
R3299 gnd.n3754 gnd.t123 371.625
R3300 gnd.n1337 gnd.t112 371.625
R3301 gnd.n156 gnd.t94 371.625
R3302 gnd.n6768 gnd.t120 371.625
R3303 gnd.n852 gnd.t194 371.625
R3304 gnd.n874 gnd.t180 371.625
R3305 gnd.n2106 gnd.t170 371.625
R3306 gnd.n1996 gnd.t116 371.625
R3307 gnd.n1974 gnd.t154 371.625
R3308 gnd.n3474 gnd.t133 371.625
R3309 gnd.n4786 gnd.t98 323.425
R3310 gnd.n4437 gnd.t129 323.425
R3311 gnd.n5641 gnd.n5615 289.615
R3312 gnd.n5609 gnd.n5583 289.615
R3313 gnd.n5577 gnd.n5551 289.615
R3314 gnd.n5546 gnd.n5520 289.615
R3315 gnd.n5514 gnd.n5488 289.615
R3316 gnd.n5482 gnd.n5456 289.615
R3317 gnd.n5450 gnd.n5424 289.615
R3318 gnd.n5419 gnd.n5393 289.615
R3319 gnd.n4860 gnd.t197 279.217
R3320 gnd.n4481 gnd.t105 279.217
R3321 gnd.n1754 gnd.t111 260.649
R3322 gnd.n3553 gnd.t147 260.649
R3323 gnd.n2753 gnd.n2752 256.663
R3324 gnd.n2752 gnd.n1771 256.663
R3325 gnd.n2752 gnd.n1772 256.663
R3326 gnd.n2752 gnd.n1773 256.663
R3327 gnd.n2752 gnd.n1774 256.663
R3328 gnd.n2752 gnd.n1775 256.663
R3329 gnd.n2752 gnd.n1776 256.663
R3330 gnd.n2752 gnd.n1777 256.663
R3331 gnd.n2752 gnd.n1778 256.663
R3332 gnd.n2752 gnd.n1779 256.663
R3333 gnd.n2752 gnd.n1780 256.663
R3334 gnd.n2752 gnd.n1781 256.663
R3335 gnd.n2752 gnd.n1782 256.663
R3336 gnd.n2752 gnd.n1783 256.663
R3337 gnd.n2752 gnd.n1784 256.663
R3338 gnd.n2752 gnd.n1785 256.663
R3339 gnd.n2595 gnd.n2592 256.663
R3340 gnd.n2752 gnd.n1786 256.663
R3341 gnd.n2752 gnd.n1787 256.663
R3342 gnd.n2752 gnd.n1788 256.663
R3343 gnd.n2752 gnd.n1789 256.663
R3344 gnd.n2752 gnd.n1790 256.663
R3345 gnd.n2752 gnd.n1791 256.663
R3346 gnd.n2752 gnd.n1792 256.663
R3347 gnd.n2752 gnd.n1793 256.663
R3348 gnd.n2752 gnd.n1794 256.663
R3349 gnd.n2752 gnd.n1795 256.663
R3350 gnd.n2752 gnd.n1796 256.663
R3351 gnd.n2752 gnd.n1797 256.663
R3352 gnd.n2752 gnd.n1798 256.663
R3353 gnd.n2752 gnd.n1799 256.663
R3354 gnd.n2752 gnd.n1800 256.663
R3355 gnd.n2752 gnd.n1801 256.663
R3356 gnd.n2752 gnd.n1802 256.663
R3357 gnd.n3695 gnd.n1382 256.663
R3358 gnd.n3695 gnd.n1383 256.663
R3359 gnd.n3695 gnd.n1384 256.663
R3360 gnd.n3695 gnd.n1385 256.663
R3361 gnd.n3695 gnd.n1386 256.663
R3362 gnd.n3695 gnd.n1387 256.663
R3363 gnd.n3695 gnd.n1388 256.663
R3364 gnd.n3695 gnd.n1389 256.663
R3365 gnd.n3695 gnd.n1390 256.663
R3366 gnd.n3695 gnd.n1391 256.663
R3367 gnd.n3695 gnd.n1392 256.663
R3368 gnd.n3695 gnd.n1393 256.663
R3369 gnd.n3695 gnd.n1394 256.663
R3370 gnd.n3695 gnd.n1395 256.663
R3371 gnd.n3695 gnd.n1396 256.663
R3372 gnd.n3695 gnd.n3692 256.663
R3373 gnd.n3698 gnd.n1363 256.663
R3374 gnd.n3696 gnd.n3695 256.663
R3375 gnd.n3695 gnd.n1381 256.663
R3376 gnd.n3695 gnd.n1380 256.663
R3377 gnd.n3695 gnd.n1379 256.663
R3378 gnd.n3695 gnd.n1378 256.663
R3379 gnd.n3695 gnd.n1377 256.663
R3380 gnd.n3695 gnd.n1376 256.663
R3381 gnd.n3695 gnd.n1375 256.663
R3382 gnd.n3695 gnd.n1374 256.663
R3383 gnd.n3695 gnd.n1373 256.663
R3384 gnd.n3695 gnd.n1372 256.663
R3385 gnd.n3695 gnd.n1371 256.663
R3386 gnd.n3695 gnd.n1370 256.663
R3387 gnd.n3695 gnd.n1369 256.663
R3388 gnd.n3695 gnd.n1368 256.663
R3389 gnd.n3695 gnd.n1367 256.663
R3390 gnd.n3695 gnd.n1366 256.663
R3391 gnd.n4406 gnd.n820 242.672
R3392 gnd.n4406 gnd.n821 242.672
R3393 gnd.n4406 gnd.n822 242.672
R3394 gnd.n4406 gnd.n823 242.672
R3395 gnd.n4406 gnd.n824 242.672
R3396 gnd.n4406 gnd.n825 242.672
R3397 gnd.n4406 gnd.n826 242.672
R3398 gnd.n4406 gnd.n827 242.672
R3399 gnd.n4406 gnd.n828 242.672
R3400 gnd.n2626 gnd.n2625 242.672
R3401 gnd.n2625 gnd.n1933 242.672
R3402 gnd.n2625 gnd.n1932 242.672
R3403 gnd.n2625 gnd.n1930 242.672
R3404 gnd.n2625 gnd.n1928 242.672
R3405 gnd.n2625 gnd.n1927 242.672
R3406 gnd.n2625 gnd.n1925 242.672
R3407 gnd.n2625 gnd.n1923 242.672
R3408 gnd.n2625 gnd.n1922 242.672
R3409 gnd.n3372 gnd.n1204 242.672
R3410 gnd.n3374 gnd.n1204 242.672
R3411 gnd.n3391 gnd.n1204 242.672
R3412 gnd.n3393 gnd.n1204 242.672
R3413 gnd.n3410 gnd.n1204 242.672
R3414 gnd.n3412 gnd.n1204 242.672
R3415 gnd.n3429 gnd.n1204 242.672
R3416 gnd.n3431 gnd.n1204 242.672
R3417 gnd.n3450 gnd.n1204 242.672
R3418 gnd.n6678 gnd.n83 242.672
R3419 gnd.n6674 gnd.n83 242.672
R3420 gnd.n6669 gnd.n83 242.672
R3421 gnd.n6666 gnd.n83 242.672
R3422 gnd.n6661 gnd.n83 242.672
R3423 gnd.n6658 gnd.n83 242.672
R3424 gnd.n6653 gnd.n83 242.672
R3425 gnd.n6650 gnd.n83 242.672
R3426 gnd.n6645 gnd.n83 242.672
R3427 gnd.n4914 gnd.n4913 242.672
R3428 gnd.n4914 gnd.n4824 242.672
R3429 gnd.n4914 gnd.n4825 242.672
R3430 gnd.n4914 gnd.n4826 242.672
R3431 gnd.n4914 gnd.n4827 242.672
R3432 gnd.n4914 gnd.n4828 242.672
R3433 gnd.n4914 gnd.n4829 242.672
R3434 gnd.n4914 gnd.n4830 242.672
R3435 gnd.n4914 gnd.n4831 242.672
R3436 gnd.n4914 gnd.n4832 242.672
R3437 gnd.n4914 gnd.n4833 242.672
R3438 gnd.n4914 gnd.n4834 242.672
R3439 gnd.n4915 gnd.n4914 242.672
R3440 gnd.n5715 gnd.n4407 242.672
R3441 gnd.n5721 gnd.n4407 242.672
R3442 gnd.n4484 gnd.n4407 242.672
R3443 gnd.n5728 gnd.n4407 242.672
R3444 gnd.n4475 gnd.n4407 242.672
R3445 gnd.n5735 gnd.n4407 242.672
R3446 gnd.n4468 gnd.n4407 242.672
R3447 gnd.n5742 gnd.n4407 242.672
R3448 gnd.n4461 gnd.n4407 242.672
R3449 gnd.n5749 gnd.n4407 242.672
R3450 gnd.n4454 gnd.n4407 242.672
R3451 gnd.n5756 gnd.n4407 242.672
R3452 gnd.n4447 gnd.n4407 242.672
R3453 gnd.n5072 gnd.n5071 242.672
R3454 gnd.n5071 gnd.n4736 242.672
R3455 gnd.n5071 gnd.n4737 242.672
R3456 gnd.n5071 gnd.n4738 242.672
R3457 gnd.n5071 gnd.n4739 242.672
R3458 gnd.n5071 gnd.n4740 242.672
R3459 gnd.n5071 gnd.n4741 242.672
R3460 gnd.n5071 gnd.n4742 242.672
R3461 gnd.n5767 gnd.n4407 242.672
R3462 gnd.n4440 gnd.n4407 242.672
R3463 gnd.n5774 gnd.n4407 242.672
R3464 gnd.n4431 gnd.n4407 242.672
R3465 gnd.n5781 gnd.n4407 242.672
R3466 gnd.n4424 gnd.n4407 242.672
R3467 gnd.n5788 gnd.n4407 242.672
R3468 gnd.n4417 gnd.n4407 242.672
R3469 gnd.n4406 gnd.n4405 242.672
R3470 gnd.n4406 gnd.n802 242.672
R3471 gnd.n4406 gnd.n803 242.672
R3472 gnd.n4406 gnd.n804 242.672
R3473 gnd.n4406 gnd.n805 242.672
R3474 gnd.n4406 gnd.n806 242.672
R3475 gnd.n4406 gnd.n807 242.672
R3476 gnd.n4406 gnd.n808 242.672
R3477 gnd.n4406 gnd.n809 242.672
R3478 gnd.n4406 gnd.n810 242.672
R3479 gnd.n4406 gnd.n811 242.672
R3480 gnd.n4406 gnd.n812 242.672
R3481 gnd.n4406 gnd.n813 242.672
R3482 gnd.n4406 gnd.n814 242.672
R3483 gnd.n4406 gnd.n815 242.672
R3484 gnd.n4406 gnd.n816 242.672
R3485 gnd.n4406 gnd.n817 242.672
R3486 gnd.n4406 gnd.n818 242.672
R3487 gnd.n4406 gnd.n819 242.672
R3488 gnd.n2625 gnd.n1935 242.672
R3489 gnd.n2625 gnd.n1936 242.672
R3490 gnd.n2625 gnd.n1937 242.672
R3491 gnd.n2625 gnd.n1938 242.672
R3492 gnd.n2625 gnd.n1939 242.672
R3493 gnd.n2625 gnd.n1940 242.672
R3494 gnd.n2625 gnd.n1941 242.672
R3495 gnd.n2625 gnd.n1942 242.672
R3496 gnd.n2625 gnd.n1943 242.672
R3497 gnd.n2625 gnd.n1944 242.672
R3498 gnd.n2625 gnd.n1945 242.672
R3499 gnd.n2596 gnd.n1976 242.672
R3500 gnd.n2625 gnd.n1946 242.672
R3501 gnd.n2625 gnd.n1947 242.672
R3502 gnd.n2625 gnd.n1948 242.672
R3503 gnd.n2625 gnd.n1949 242.672
R3504 gnd.n2625 gnd.n1950 242.672
R3505 gnd.n2625 gnd.n1951 242.672
R3506 gnd.n2625 gnd.n1952 242.672
R3507 gnd.n2625 gnd.n2624 242.672
R3508 gnd.n3717 gnd.n1204 242.672
R3509 gnd.n3720 gnd.n1204 242.672
R3510 gnd.n3728 gnd.n1204 242.672
R3511 gnd.n3730 gnd.n1204 242.672
R3512 gnd.n3738 gnd.n1204 242.672
R3513 gnd.n3740 gnd.n1204 242.672
R3514 gnd.n3749 gnd.n1204 242.672
R3515 gnd.n3752 gnd.n1204 242.672
R3516 gnd.n3756 gnd.n3753 242.672
R3517 gnd.n3699 gnd.n1204 242.672
R3518 gnd.n3762 gnd.n1204 242.672
R3519 gnd.n3764 gnd.n1204 242.672
R3520 gnd.n3772 gnd.n1204 242.672
R3521 gnd.n3774 gnd.n1204 242.672
R3522 gnd.n3782 gnd.n1204 242.672
R3523 gnd.n3784 gnd.n1204 242.672
R3524 gnd.n3792 gnd.n1204 242.672
R3525 gnd.n3794 gnd.n1204 242.672
R3526 gnd.n3803 gnd.n1204 242.672
R3527 gnd.n3806 gnd.n1204 242.672
R3528 gnd.n153 gnd.n83 242.672
R3529 gnd.n6736 gnd.n83 242.672
R3530 gnd.n149 gnd.n83 242.672
R3531 gnd.n6743 gnd.n83 242.672
R3532 gnd.n142 gnd.n83 242.672
R3533 gnd.n6750 gnd.n83 242.672
R3534 gnd.n135 gnd.n83 242.672
R3535 gnd.n6757 gnd.n83 242.672
R3536 gnd.n128 gnd.n83 242.672
R3537 gnd.n6764 gnd.n83 242.672
R3538 gnd.n121 gnd.n83 242.672
R3539 gnd.n6774 gnd.n83 242.672
R3540 gnd.n114 gnd.n83 242.672
R3541 gnd.n6781 gnd.n83 242.672
R3542 gnd.n107 gnd.n83 242.672
R3543 gnd.n6788 gnd.n83 242.672
R3544 gnd.n100 gnd.n83 242.672
R3545 gnd.n6795 gnd.n83 242.672
R3546 gnd.n93 gnd.n83 242.672
R3547 gnd.n2675 gnd.n2674 242.672
R3548 gnd.n2675 gnd.n1850 242.672
R3549 gnd.n2675 gnd.n1851 242.672
R3550 gnd.n2675 gnd.n1852 242.672
R3551 gnd.n2675 gnd.n1853 242.672
R3552 gnd.n2675 gnd.n1854 242.672
R3553 gnd.n2675 gnd.n1855 242.672
R3554 gnd.n2675 gnd.n1856 242.672
R3555 gnd.n2675 gnd.n1857 242.672
R3556 gnd.n2675 gnd.n1858 242.672
R3557 gnd.n2675 gnd.n1859 242.672
R3558 gnd.n2675 gnd.n1860 242.672
R3559 gnd.n2675 gnd.n1861 242.672
R3560 gnd.n2676 gnd.n2675 242.672
R3561 gnd.n3483 gnd.n1203 242.672
R3562 gnd.n3472 gnd.n1203 242.672
R3563 gnd.n3470 gnd.n1203 242.672
R3564 gnd.n3462 gnd.n1203 242.672
R3565 gnd.n3460 gnd.n1203 242.672
R3566 gnd.n3442 gnd.n1203 242.672
R3567 gnd.n3440 gnd.n1203 242.672
R3568 gnd.n3334 gnd.n1203 242.672
R3569 gnd.n3421 gnd.n1203 242.672
R3570 gnd.n3343 gnd.n1203 242.672
R3571 gnd.n3402 gnd.n1203 242.672
R3572 gnd.n3352 gnd.n1203 242.672
R3573 gnd.n3383 gnd.n1203 242.672
R3574 gnd.n3361 gnd.n1203 242.672
R3575 gnd.n90 gnd.n86 240.244
R3576 gnd.n6797 gnd.n6796 240.244
R3577 gnd.n6794 gnd.n94 240.244
R3578 gnd.n6790 gnd.n6789 240.244
R3579 gnd.n6787 gnd.n101 240.244
R3580 gnd.n6783 gnd.n6782 240.244
R3581 gnd.n6780 gnd.n108 240.244
R3582 gnd.n6776 gnd.n6775 240.244
R3583 gnd.n6773 gnd.n115 240.244
R3584 gnd.n6766 gnd.n6765 240.244
R3585 gnd.n6763 gnd.n122 240.244
R3586 gnd.n6759 gnd.n6758 240.244
R3587 gnd.n6756 gnd.n129 240.244
R3588 gnd.n6752 gnd.n6751 240.244
R3589 gnd.n6749 gnd.n136 240.244
R3590 gnd.n6745 gnd.n6744 240.244
R3591 gnd.n6742 gnd.n143 240.244
R3592 gnd.n6738 gnd.n6737 240.244
R3593 gnd.n6735 gnd.n150 240.244
R3594 gnd.n3813 gnd.n1213 240.244
R3595 gnd.n3813 gnd.n1225 240.244
R3596 gnd.n3824 gnd.n1225 240.244
R3597 gnd.n3824 gnd.n1326 240.244
R3598 gnd.n3915 gnd.n1326 240.244
R3599 gnd.n3915 gnd.n1319 240.244
R3600 gnd.n3911 gnd.n1319 240.244
R3601 gnd.n3911 gnd.n1311 240.244
R3602 gnd.n1311 gnd.n1300 240.244
R3603 gnd.n3907 gnd.n1300 240.244
R3604 gnd.n3907 gnd.n1290 240.244
R3605 gnd.n3904 gnd.n1290 240.244
R3606 gnd.n3904 gnd.n1282 240.244
R3607 gnd.n1282 gnd.n1271 240.244
R3608 gnd.n3900 gnd.n1271 240.244
R3609 gnd.n3900 gnd.n1261 240.244
R3610 gnd.n3897 gnd.n1261 240.244
R3611 gnd.n3897 gnd.n1252 240.244
R3612 gnd.n1252 gnd.n249 240.244
R3613 gnd.n249 gnd.n244 240.244
R3614 gnd.n3891 gnd.n244 240.244
R3615 gnd.n3891 gnd.n237 240.244
R3616 gnd.n3886 gnd.n237 240.244
R3617 gnd.n3886 gnd.n231 240.244
R3618 gnd.n3883 gnd.n231 240.244
R3619 gnd.n3883 gnd.n223 240.244
R3620 gnd.n3880 gnd.n223 240.244
R3621 gnd.n3880 gnd.n209 240.244
R3622 gnd.n3877 gnd.n209 240.244
R3623 gnd.n3877 gnd.n203 240.244
R3624 gnd.n3874 gnd.n203 240.244
R3625 gnd.n3874 gnd.n195 240.244
R3626 gnd.n3871 gnd.n195 240.244
R3627 gnd.n3871 gnd.n187 240.244
R3628 gnd.n3868 gnd.n187 240.244
R3629 gnd.n3868 gnd.n179 240.244
R3630 gnd.n3865 gnd.n179 240.244
R3631 gnd.n3865 gnd.n171 240.244
R3632 gnd.n171 gnd.n160 240.244
R3633 gnd.n6726 gnd.n160 240.244
R3634 gnd.n6727 gnd.n6726 240.244
R3635 gnd.n6727 gnd.n82 240.244
R3636 gnd.n3719 gnd.n3718 240.244
R3637 gnd.n3721 gnd.n3719 240.244
R3638 gnd.n3727 gnd.n3709 240.244
R3639 gnd.n3731 gnd.n3729 240.244
R3640 gnd.n3737 gnd.n3705 240.244
R3641 gnd.n3741 gnd.n3739 240.244
R3642 gnd.n3748 gnd.n3701 240.244
R3643 gnd.n3751 gnd.n3750 240.244
R3644 gnd.n3761 gnd.n1357 240.244
R3645 gnd.n3765 gnd.n3763 240.244
R3646 gnd.n3771 gnd.n1353 240.244
R3647 gnd.n3775 gnd.n3773 240.244
R3648 gnd.n3781 gnd.n1349 240.244
R3649 gnd.n3785 gnd.n3783 240.244
R3650 gnd.n3791 gnd.n1345 240.244
R3651 gnd.n3795 gnd.n3793 240.244
R3652 gnd.n3802 gnd.n1341 240.244
R3653 gnd.n3805 gnd.n3804 240.244
R3654 gnd.n4053 gnd.n1218 240.244
R3655 gnd.n4049 gnd.n1218 240.244
R3656 gnd.n4049 gnd.n1223 240.244
R3657 gnd.n3935 gnd.n1223 240.244
R3658 gnd.n3935 gnd.n1321 240.244
R3659 gnd.n3943 gnd.n1321 240.244
R3660 gnd.n3943 gnd.n1322 240.244
R3661 gnd.n1322 gnd.n1298 240.244
R3662 gnd.n3966 gnd.n1298 240.244
R3663 gnd.n3966 gnd.n1293 240.244
R3664 gnd.n3975 gnd.n1293 240.244
R3665 gnd.n3975 gnd.n1294 240.244
R3666 gnd.n1294 gnd.n1269 240.244
R3667 gnd.n4005 gnd.n1269 240.244
R3668 gnd.n4005 gnd.n1263 240.244
R3669 gnd.n4009 gnd.n1263 240.244
R3670 gnd.n4009 gnd.n1266 240.244
R3671 gnd.n1266 gnd.n247 240.244
R3672 gnd.n6569 gnd.n247 240.244
R3673 gnd.n6572 gnd.n6569 240.244
R3674 gnd.n6572 gnd.n233 240.244
R3675 gnd.n6582 gnd.n233 240.244
R3676 gnd.n6583 gnd.n6582 240.244
R3677 gnd.n6586 gnd.n6583 240.244
R3678 gnd.n6586 gnd.n220 240.244
R3679 gnd.n6596 gnd.n220 240.244
R3680 gnd.n6596 gnd.n210 240.244
R3681 gnd.n6602 gnd.n210 240.244
R3682 gnd.n6602 gnd.n200 240.244
R3683 gnd.n6612 gnd.n200 240.244
R3684 gnd.n6612 gnd.n196 240.244
R3685 gnd.n6618 gnd.n196 240.244
R3686 gnd.n6618 gnd.n184 240.244
R3687 gnd.n6628 gnd.n184 240.244
R3688 gnd.n6628 gnd.n180 240.244
R3689 gnd.n6634 gnd.n180 240.244
R3690 gnd.n6634 gnd.n168 240.244
R3691 gnd.n6718 gnd.n168 240.244
R3692 gnd.n6718 gnd.n164 240.244
R3693 gnd.n6724 gnd.n164 240.244
R3694 gnd.n6724 gnd.n85 240.244
R3695 gnd.n6804 gnd.n85 240.244
R3696 gnd.n1953 gnd.n1078 240.244
R3697 gnd.n2623 gnd.n1954 240.244
R3698 gnd.n2619 gnd.n2618 240.244
R3699 gnd.n2615 gnd.n2614 240.244
R3700 gnd.n2611 gnd.n2610 240.244
R3701 gnd.n2607 gnd.n2606 240.244
R3702 gnd.n2603 gnd.n2602 240.244
R3703 gnd.n2599 gnd.n2598 240.244
R3704 gnd.n2462 gnd.n2461 240.244
R3705 gnd.n2459 gnd.n2458 240.244
R3706 gnd.n2455 gnd.n2454 240.244
R3707 gnd.n2451 gnd.n2450 240.244
R3708 gnd.n2447 gnd.n2446 240.244
R3709 gnd.n2443 gnd.n2442 240.244
R3710 gnd.n2439 gnd.n2438 240.244
R3711 gnd.n2435 gnd.n2434 240.244
R3712 gnd.n2431 gnd.n2430 240.244
R3713 gnd.n2427 gnd.n2426 240.244
R3714 gnd.n4327 gnd.n878 240.244
R3715 gnd.n882 gnd.n878 240.244
R3716 gnd.n4320 gnd.n882 240.244
R3717 gnd.n4320 gnd.n883 240.244
R3718 gnd.n896 gnd.n883 240.244
R3719 gnd.n2206 gnd.n896 240.244
R3720 gnd.n2206 gnd.n907 240.244
R3721 gnd.n2201 gnd.n907 240.244
R3722 gnd.n2201 gnd.n917 240.244
R3723 gnd.n2213 gnd.n917 240.244
R3724 gnd.n2213 gnd.n927 240.244
R3725 gnd.n2198 gnd.n927 240.244
R3726 gnd.n2198 gnd.n937 240.244
R3727 gnd.n2220 gnd.n937 240.244
R3728 gnd.n2220 gnd.n947 240.244
R3729 gnd.n2195 gnd.n947 240.244
R3730 gnd.n2232 gnd.n2195 240.244
R3731 gnd.n2232 gnd.n958 240.244
R3732 gnd.n2228 gnd.n958 240.244
R3733 gnd.n2228 gnd.n971 240.244
R3734 gnd.n2245 gnd.n971 240.244
R3735 gnd.n2245 gnd.n979 240.244
R3736 gnd.n2252 gnd.n979 240.244
R3737 gnd.n2252 gnd.n988 240.244
R3738 gnd.n2262 gnd.n988 240.244
R3739 gnd.n2262 gnd.n996 240.244
R3740 gnd.n2022 gnd.n996 240.244
R3741 gnd.n2022 gnd.n1006 240.244
R3742 gnd.n2270 gnd.n1006 240.244
R3743 gnd.n2270 gnd.n1017 240.244
R3744 gnd.n2275 gnd.n1017 240.244
R3745 gnd.n2275 gnd.n1027 240.244
R3746 gnd.n2285 gnd.n1027 240.244
R3747 gnd.n2285 gnd.n1038 240.244
R3748 gnd.n2010 gnd.n1038 240.244
R3749 gnd.n2010 gnd.n1048 240.244
R3750 gnd.n2370 gnd.n1048 240.244
R3751 gnd.n2370 gnd.n1059 240.244
R3752 gnd.n2377 gnd.n1059 240.244
R3753 gnd.n2377 gnd.n1070 240.244
R3754 gnd.n2419 gnd.n1070 240.244
R3755 gnd.n2419 gnd.n1080 240.244
R3756 gnd.n832 gnd.n831 240.244
R3757 gnd.n4399 gnd.n831 240.244
R3758 gnd.n4397 gnd.n4396 240.244
R3759 gnd.n4393 gnd.n4392 240.244
R3760 gnd.n4389 gnd.n4388 240.244
R3761 gnd.n4385 gnd.n4384 240.244
R3762 gnd.n4381 gnd.n4380 240.244
R3763 gnd.n4377 gnd.n4376 240.244
R3764 gnd.n4373 gnd.n4372 240.244
R3765 gnd.n4368 gnd.n4367 240.244
R3766 gnd.n4364 gnd.n4363 240.244
R3767 gnd.n4360 gnd.n4359 240.244
R3768 gnd.n4356 gnd.n4355 240.244
R3769 gnd.n4352 gnd.n4351 240.244
R3770 gnd.n4348 gnd.n4347 240.244
R3771 gnd.n4344 gnd.n4343 240.244
R3772 gnd.n4340 gnd.n4339 240.244
R3773 gnd.n4336 gnd.n4335 240.244
R3774 gnd.n873 gnd.n872 240.244
R3775 gnd.n2164 gnd.n833 240.244
R3776 gnd.n2164 gnd.n888 240.244
R3777 gnd.n4318 gnd.n888 240.244
R3778 gnd.n4318 gnd.n889 240.244
R3779 gnd.n4314 gnd.n889 240.244
R3780 gnd.n4314 gnd.n895 240.244
R3781 gnd.n4306 gnd.n895 240.244
R3782 gnd.n4306 gnd.n910 240.244
R3783 gnd.n4302 gnd.n910 240.244
R3784 gnd.n4302 gnd.n916 240.244
R3785 gnd.n4294 gnd.n916 240.244
R3786 gnd.n4294 gnd.n929 240.244
R3787 gnd.n4290 gnd.n929 240.244
R3788 gnd.n4290 gnd.n935 240.244
R3789 gnd.n4282 gnd.n935 240.244
R3790 gnd.n4282 gnd.n950 240.244
R3791 gnd.n954 gnd.n950 240.244
R3792 gnd.n4276 gnd.n954 240.244
R3793 gnd.n4276 gnd.n956 240.244
R3794 gnd.n4268 gnd.n956 240.244
R3795 gnd.n4268 gnd.n974 240.244
R3796 gnd.n4263 gnd.n974 240.244
R3797 gnd.n4263 gnd.n977 240.244
R3798 gnd.n4255 gnd.n977 240.244
R3799 gnd.n4255 gnd.n991 240.244
R3800 gnd.n4250 gnd.n991 240.244
R3801 gnd.n4250 gnd.n994 240.244
R3802 gnd.n4242 gnd.n994 240.244
R3803 gnd.n4242 gnd.n1009 240.244
R3804 gnd.n4238 gnd.n1009 240.244
R3805 gnd.n4238 gnd.n1015 240.244
R3806 gnd.n4230 gnd.n1015 240.244
R3807 gnd.n4230 gnd.n1030 240.244
R3808 gnd.n4226 gnd.n1030 240.244
R3809 gnd.n4226 gnd.n1036 240.244
R3810 gnd.n4218 gnd.n1036 240.244
R3811 gnd.n4218 gnd.n1051 240.244
R3812 gnd.n4214 gnd.n1051 240.244
R3813 gnd.n4214 gnd.n1057 240.244
R3814 gnd.n4206 gnd.n1057 240.244
R3815 gnd.n4206 gnd.n1073 240.244
R3816 gnd.n4202 gnd.n1073 240.244
R3817 gnd.n4414 gnd.n4409 240.244
R3818 gnd.n5790 gnd.n5789 240.244
R3819 gnd.n5787 gnd.n4418 240.244
R3820 gnd.n5783 gnd.n5782 240.244
R3821 gnd.n5780 gnd.n4425 240.244
R3822 gnd.n5776 gnd.n5775 240.244
R3823 gnd.n5773 gnd.n4432 240.244
R3824 gnd.n5769 gnd.n5768 240.244
R3825 gnd.n5083 gnd.n4721 240.244
R3826 gnd.n5093 gnd.n4721 240.244
R3827 gnd.n5093 gnd.n4712 240.244
R3828 gnd.n4712 gnd.n4701 240.244
R3829 gnd.n5114 gnd.n4701 240.244
R3830 gnd.n5114 gnd.n4695 240.244
R3831 gnd.n5124 gnd.n4695 240.244
R3832 gnd.n5124 gnd.n4686 240.244
R3833 gnd.n4686 gnd.n4677 240.244
R3834 gnd.n5145 gnd.n4677 240.244
R3835 gnd.n5145 gnd.n4670 240.244
R3836 gnd.n5155 gnd.n4670 240.244
R3837 gnd.n5155 gnd.n4661 240.244
R3838 gnd.n4661 gnd.n4651 240.244
R3839 gnd.n5176 gnd.n4651 240.244
R3840 gnd.n5176 gnd.n4644 240.244
R3841 gnd.n5186 gnd.n4644 240.244
R3842 gnd.n5186 gnd.n4635 240.244
R3843 gnd.n4635 gnd.n4626 240.244
R3844 gnd.n5207 gnd.n4626 240.244
R3845 gnd.n5207 gnd.n4619 240.244
R3846 gnd.n5217 gnd.n4619 240.244
R3847 gnd.n5217 gnd.n4611 240.244
R3848 gnd.n4611 gnd.n4602 240.244
R3849 gnd.n5237 gnd.n4602 240.244
R3850 gnd.n5237 gnd.n4589 240.244
R3851 gnd.n5271 gnd.n4589 240.244
R3852 gnd.n5271 gnd.n4579 240.244
R3853 gnd.n4579 gnd.n4571 240.244
R3854 gnd.n5289 gnd.n4571 240.244
R3855 gnd.n5290 gnd.n5289 240.244
R3856 gnd.n5290 gnd.n4559 240.244
R3857 gnd.n4559 gnd.n4548 240.244
R3858 gnd.n5321 gnd.n4548 240.244
R3859 gnd.n5322 gnd.n5321 240.244
R3860 gnd.n5325 gnd.n5322 240.244
R3861 gnd.n5325 gnd.n4534 240.244
R3862 gnd.n5353 gnd.n4534 240.244
R3863 gnd.n5353 gnd.n4521 240.244
R3864 gnd.n5375 gnd.n4521 240.244
R3865 gnd.n5376 gnd.n5375 240.244
R3866 gnd.n5376 gnd.n4505 240.244
R3867 gnd.n5386 gnd.n4505 240.244
R3868 gnd.n5386 gnd.n4497 240.244
R3869 gnd.n5668 gnd.n4497 240.244
R3870 gnd.n5668 gnd.n5667 240.244
R3871 gnd.n5667 gnd.n5666 240.244
R3872 gnd.n5666 gnd.n778 240.244
R3873 gnd.n5662 gnd.n778 240.244
R3874 gnd.n5662 gnd.n789 240.244
R3875 gnd.n5658 gnd.n789 240.244
R3876 gnd.n5658 gnd.n5657 240.244
R3877 gnd.n5657 gnd.n801 240.244
R3878 gnd.n5073 gnd.n4734 240.244
R3879 gnd.n4755 gnd.n4734 240.244
R3880 gnd.n4758 gnd.n4757 240.244
R3881 gnd.n4765 gnd.n4764 240.244
R3882 gnd.n4768 gnd.n4767 240.244
R3883 gnd.n4775 gnd.n4774 240.244
R3884 gnd.n4778 gnd.n4777 240.244
R3885 gnd.n4785 gnd.n4784 240.244
R3886 gnd.n5081 gnd.n4731 240.244
R3887 gnd.n4731 gnd.n4710 240.244
R3888 gnd.n5104 gnd.n4710 240.244
R3889 gnd.n5104 gnd.n4704 240.244
R3890 gnd.n5112 gnd.n4704 240.244
R3891 gnd.n5112 gnd.n4706 240.244
R3892 gnd.n4706 gnd.n4684 240.244
R3893 gnd.n5135 gnd.n4684 240.244
R3894 gnd.n5135 gnd.n4679 240.244
R3895 gnd.n5143 gnd.n4679 240.244
R3896 gnd.n5143 gnd.n4680 240.244
R3897 gnd.n4680 gnd.n4659 240.244
R3898 gnd.n5166 gnd.n4659 240.244
R3899 gnd.n5166 gnd.n4654 240.244
R3900 gnd.n5174 gnd.n4654 240.244
R3901 gnd.n5174 gnd.n4655 240.244
R3902 gnd.n4655 gnd.n4633 240.244
R3903 gnd.n5197 gnd.n4633 240.244
R3904 gnd.n5197 gnd.n4628 240.244
R3905 gnd.n5205 gnd.n4628 240.244
R3906 gnd.n5205 gnd.n4629 240.244
R3907 gnd.n4629 gnd.n4609 240.244
R3908 gnd.n5227 gnd.n4609 240.244
R3909 gnd.n5227 gnd.n4604 240.244
R3910 gnd.n5235 gnd.n4604 240.244
R3911 gnd.n5235 gnd.n4605 240.244
R3912 gnd.n4605 gnd.n4578 240.244
R3913 gnd.n5281 gnd.n4578 240.244
R3914 gnd.n5281 gnd.n4574 240.244
R3915 gnd.n5287 gnd.n4574 240.244
R3916 gnd.n5287 gnd.n4557 240.244
R3917 gnd.n5311 gnd.n4557 240.244
R3918 gnd.n5311 gnd.n4552 240.244
R3919 gnd.n5319 gnd.n4552 240.244
R3920 gnd.n5319 gnd.n4553 240.244
R3921 gnd.n4553 gnd.n4533 240.244
R3922 gnd.n5357 gnd.n4533 240.244
R3923 gnd.n5357 gnd.n4528 240.244
R3924 gnd.n5365 gnd.n4528 240.244
R3925 gnd.n5365 gnd.n4529 240.244
R3926 gnd.n4529 gnd.n4503 240.244
R3927 gnd.n5678 gnd.n4503 240.244
R3928 gnd.n5678 gnd.n4498 240.244
R3929 gnd.n5690 gnd.n4498 240.244
R3930 gnd.n5690 gnd.n4499 240.244
R3931 gnd.n5686 gnd.n4499 240.244
R3932 gnd.n5686 gnd.n780 240.244
R3933 gnd.n5811 gnd.n780 240.244
R3934 gnd.n5811 gnd.n781 240.244
R3935 gnd.n5807 gnd.n781 240.244
R3936 gnd.n5807 gnd.n787 240.244
R3937 gnd.n4408 gnd.n787 240.244
R3938 gnd.n5797 gnd.n4408 240.244
R3939 gnd.n4444 gnd.n798 240.244
R3940 gnd.n5758 gnd.n5757 240.244
R3941 gnd.n5755 gnd.n4448 240.244
R3942 gnd.n5751 gnd.n5750 240.244
R3943 gnd.n5748 gnd.n4455 240.244
R3944 gnd.n5744 gnd.n5743 240.244
R3945 gnd.n5741 gnd.n4462 240.244
R3946 gnd.n5737 gnd.n5736 240.244
R3947 gnd.n5734 gnd.n4469 240.244
R3948 gnd.n5730 gnd.n5729 240.244
R3949 gnd.n5727 gnd.n4476 240.244
R3950 gnd.n5723 gnd.n5722 240.244
R3951 gnd.n5720 gnd.n4486 240.244
R3952 gnd.n4922 gnd.n4819 240.244
R3953 gnd.n4922 gnd.n4812 240.244
R3954 gnd.n4933 gnd.n4812 240.244
R3955 gnd.n4933 gnd.n4808 240.244
R3956 gnd.n4939 gnd.n4808 240.244
R3957 gnd.n4939 gnd.n4800 240.244
R3958 gnd.n4949 gnd.n4800 240.244
R3959 gnd.n4949 gnd.n4795 240.244
R3960 gnd.n5059 gnd.n4795 240.244
R3961 gnd.n5059 gnd.n4796 240.244
R3962 gnd.n4796 gnd.n4743 240.244
R3963 gnd.n5054 gnd.n4743 240.244
R3964 gnd.n5054 gnd.n5053 240.244
R3965 gnd.n5053 gnd.n4722 240.244
R3966 gnd.n5049 gnd.n4722 240.244
R3967 gnd.n5049 gnd.n4713 240.244
R3968 gnd.n5046 gnd.n4713 240.244
R3969 gnd.n5046 gnd.n5045 240.244
R3970 gnd.n5045 gnd.n4696 240.244
R3971 gnd.n5041 gnd.n4696 240.244
R3972 gnd.n5041 gnd.n4687 240.244
R3973 gnd.n5038 gnd.n4687 240.244
R3974 gnd.n5038 gnd.n5037 240.244
R3975 gnd.n5037 gnd.n4672 240.244
R3976 gnd.n5032 gnd.n4672 240.244
R3977 gnd.n5032 gnd.n4662 240.244
R3978 gnd.n5029 gnd.n4662 240.244
R3979 gnd.n5029 gnd.n5028 240.244
R3980 gnd.n5028 gnd.n4646 240.244
R3981 gnd.n4973 gnd.n4646 240.244
R3982 gnd.n4973 gnd.n4636 240.244
R3983 gnd.n4984 gnd.n4636 240.244
R3984 gnd.n4984 gnd.n4982 240.244
R3985 gnd.n4982 gnd.n4621 240.244
R3986 gnd.n4977 gnd.n4621 240.244
R3987 gnd.n4977 gnd.n4612 240.244
R3988 gnd.n4612 gnd.n4595 240.244
R3989 gnd.n5247 gnd.n4595 240.244
R3990 gnd.n5247 gnd.n4591 240.244
R3991 gnd.n5268 gnd.n4591 240.244
R3992 gnd.n5268 gnd.n4580 240.244
R3993 gnd.n5264 gnd.n4580 240.244
R3994 gnd.n5264 gnd.n4570 240.244
R3995 gnd.n5261 gnd.n4570 240.244
R3996 gnd.n5261 gnd.n4560 240.244
R3997 gnd.n5258 gnd.n4560 240.244
R3998 gnd.n5258 gnd.n4539 240.244
R3999 gnd.n5334 gnd.n4539 240.244
R4000 gnd.n5334 gnd.n4535 240.244
R4001 gnd.n5352 gnd.n4535 240.244
R4002 gnd.n5352 gnd.n4526 240.244
R4003 gnd.n5348 gnd.n4526 240.244
R4004 gnd.n5348 gnd.n4520 240.244
R4005 gnd.n5345 gnd.n4520 240.244
R4006 gnd.n5345 gnd.n4506 240.244
R4007 gnd.n4506 gnd.n4496 240.244
R4008 gnd.n5693 gnd.n4496 240.244
R4009 gnd.n5693 gnd.n766 240.244
R4010 gnd.n5699 gnd.n766 240.244
R4011 gnd.n5699 gnd.n777 240.244
R4012 gnd.n5703 gnd.n777 240.244
R4013 gnd.n5703 gnd.n5702 240.244
R4014 gnd.n5702 gnd.n790 240.244
R4015 gnd.n5710 gnd.n790 240.244
R4016 gnd.n5710 gnd.n800 240.244
R4017 gnd.n4836 gnd.n4835 240.244
R4018 gnd.n4907 gnd.n4835 240.244
R4019 gnd.n4905 gnd.n4904 240.244
R4020 gnd.n4901 gnd.n4900 240.244
R4021 gnd.n4897 gnd.n4896 240.244
R4022 gnd.n4893 gnd.n4892 240.244
R4023 gnd.n4889 gnd.n4888 240.244
R4024 gnd.n4885 gnd.n4884 240.244
R4025 gnd.n4881 gnd.n4880 240.244
R4026 gnd.n4877 gnd.n4876 240.244
R4027 gnd.n4873 gnd.n4872 240.244
R4028 gnd.n4869 gnd.n4868 240.244
R4029 gnd.n4865 gnd.n4823 240.244
R4030 gnd.n4925 gnd.n4817 240.244
R4031 gnd.n4925 gnd.n4813 240.244
R4032 gnd.n4931 gnd.n4813 240.244
R4033 gnd.n4931 gnd.n4806 240.244
R4034 gnd.n4941 gnd.n4806 240.244
R4035 gnd.n4941 gnd.n4802 240.244
R4036 gnd.n4947 gnd.n4802 240.244
R4037 gnd.n4947 gnd.n4793 240.244
R4038 gnd.n5061 gnd.n4793 240.244
R4039 gnd.n5061 gnd.n4744 240.244
R4040 gnd.n5069 gnd.n4744 240.244
R4041 gnd.n5069 gnd.n4745 240.244
R4042 gnd.n4745 gnd.n4723 240.244
R4043 gnd.n5090 gnd.n4723 240.244
R4044 gnd.n5090 gnd.n4715 240.244
R4045 gnd.n5101 gnd.n4715 240.244
R4046 gnd.n5101 gnd.n4716 240.244
R4047 gnd.n4716 gnd.n4697 240.244
R4048 gnd.n5121 gnd.n4697 240.244
R4049 gnd.n5121 gnd.n4689 240.244
R4050 gnd.n5132 gnd.n4689 240.244
R4051 gnd.n5132 gnd.n4690 240.244
R4052 gnd.n4690 gnd.n4673 240.244
R4053 gnd.n5152 gnd.n4673 240.244
R4054 gnd.n5152 gnd.n4664 240.244
R4055 gnd.n5163 gnd.n4664 240.244
R4056 gnd.n5163 gnd.n4665 240.244
R4057 gnd.n4665 gnd.n4647 240.244
R4058 gnd.n5183 gnd.n4647 240.244
R4059 gnd.n5183 gnd.n4638 240.244
R4060 gnd.n5194 gnd.n4638 240.244
R4061 gnd.n5194 gnd.n4639 240.244
R4062 gnd.n4639 gnd.n4622 240.244
R4063 gnd.n5214 gnd.n4622 240.244
R4064 gnd.n5214 gnd.n4614 240.244
R4065 gnd.n5224 gnd.n4614 240.244
R4066 gnd.n5224 gnd.n4597 240.244
R4067 gnd.n5245 gnd.n4597 240.244
R4068 gnd.n5245 gnd.n4598 240.244
R4069 gnd.n4598 gnd.n4582 240.244
R4070 gnd.n5278 gnd.n4582 240.244
R4071 gnd.n5278 gnd.n4569 240.244
R4072 gnd.n5293 gnd.n4569 240.244
R4073 gnd.n5293 gnd.n4562 240.244
R4074 gnd.n5308 gnd.n4562 240.244
R4075 gnd.n5308 gnd.n4563 240.244
R4076 gnd.n4563 gnd.n4541 240.244
R4077 gnd.n5332 gnd.n4541 240.244
R4078 gnd.n5332 gnd.n4542 240.244
R4079 gnd.n4542 gnd.n4525 240.244
R4080 gnd.n5368 gnd.n4525 240.244
R4081 gnd.n5368 gnd.n4518 240.244
R4082 gnd.n5379 gnd.n4518 240.244
R4083 gnd.n5379 gnd.n4508 240.244
R4084 gnd.n5675 gnd.n4508 240.244
R4085 gnd.n5675 gnd.n4510 240.244
R4086 gnd.n4510 gnd.n768 240.244
R4087 gnd.n5818 gnd.n768 240.244
R4088 gnd.n5818 gnd.n769 240.244
R4089 gnd.n5814 gnd.n769 240.244
R4090 gnd.n5814 gnd.n775 240.244
R4091 gnd.n792 gnd.n775 240.244
R4092 gnd.n5804 gnd.n792 240.244
R4093 gnd.n5804 gnd.n793 240.244
R4094 gnd.n5800 gnd.n793 240.244
R4095 gnd.n6644 gnd.n6643 240.244
R4096 gnd.n6649 gnd.n6646 240.244
R4097 gnd.n6652 gnd.n6651 240.244
R4098 gnd.n6657 gnd.n6654 240.244
R4099 gnd.n6660 gnd.n6659 240.244
R4100 gnd.n6665 gnd.n6662 240.244
R4101 gnd.n6668 gnd.n6667 240.244
R4102 gnd.n6673 gnd.n6670 240.244
R4103 gnd.n6679 gnd.n6675 240.244
R4104 gnd.n3815 gnd.n1214 240.244
R4105 gnd.n3815 gnd.n1226 240.244
R4106 gnd.n3822 gnd.n1226 240.244
R4107 gnd.n3822 gnd.n1327 240.244
R4108 gnd.n1327 gnd.n1317 240.244
R4109 gnd.n3945 gnd.n1317 240.244
R4110 gnd.n3945 gnd.n1312 240.244
R4111 gnd.n3952 gnd.n1312 240.244
R4112 gnd.n3952 gnd.n1301 240.244
R4113 gnd.n1301 gnd.n1288 240.244
R4114 gnd.n3977 gnd.n1288 240.244
R4115 gnd.n3977 gnd.n1283 240.244
R4116 gnd.n3984 gnd.n1283 240.244
R4117 gnd.n3984 gnd.n1272 240.244
R4118 gnd.n1272 gnd.n1259 240.244
R4119 gnd.n4011 gnd.n1259 240.244
R4120 gnd.n4011 gnd.n1253 240.244
R4121 gnd.n4018 gnd.n1253 240.244
R4122 gnd.n4018 gnd.n250 240.244
R4123 gnd.n250 gnd.n245 240.244
R4124 gnd.n3889 gnd.n245 240.244
R4125 gnd.n3889 gnd.n54 240.244
R4126 gnd.n55 gnd.n54 240.244
R4127 gnd.n56 gnd.n55 240.244
R4128 gnd.n221 gnd.n56 240.244
R4129 gnd.n221 gnd.n59 240.244
R4130 gnd.n60 gnd.n59 240.244
R4131 gnd.n61 gnd.n60 240.244
R4132 gnd.n201 gnd.n61 240.244
R4133 gnd.n201 gnd.n64 240.244
R4134 gnd.n65 gnd.n64 240.244
R4135 gnd.n66 gnd.n65 240.244
R4136 gnd.n185 gnd.n66 240.244
R4137 gnd.n185 gnd.n69 240.244
R4138 gnd.n70 gnd.n69 240.244
R4139 gnd.n71 gnd.n70 240.244
R4140 gnd.n169 gnd.n71 240.244
R4141 gnd.n169 gnd.n74 240.244
R4142 gnd.n75 gnd.n74 240.244
R4143 gnd.n76 gnd.n75 240.244
R4144 gnd.n79 gnd.n76 240.244
R4145 gnd.n6806 gnd.n79 240.244
R4146 gnd.n3375 gnd.n3373 240.244
R4147 gnd.n3390 gnd.n3356 240.244
R4148 gnd.n3394 gnd.n3392 240.244
R4149 gnd.n3409 gnd.n3347 240.244
R4150 gnd.n3413 gnd.n3411 240.244
R4151 gnd.n3428 gnd.n3338 240.244
R4152 gnd.n3432 gnd.n3430 240.244
R4153 gnd.n3449 gnd.n3329 240.244
R4154 gnd.n3452 gnd.n3451 240.244
R4155 gnd.n1228 gnd.n1216 240.244
R4156 gnd.n4047 gnd.n1228 240.244
R4157 gnd.n4047 gnd.n1229 240.244
R4158 gnd.n1234 gnd.n1229 240.244
R4159 gnd.n1235 gnd.n1234 240.244
R4160 gnd.n1236 gnd.n1235 240.244
R4161 gnd.n1309 gnd.n1236 240.244
R4162 gnd.n1309 gnd.n1239 240.244
R4163 gnd.n1240 gnd.n1239 240.244
R4164 gnd.n1241 gnd.n1240 240.244
R4165 gnd.n1292 gnd.n1241 240.244
R4166 gnd.n1292 gnd.n1244 240.244
R4167 gnd.n1245 gnd.n1244 240.244
R4168 gnd.n1246 gnd.n1245 240.244
R4169 gnd.n1273 gnd.n1246 240.244
R4170 gnd.n1273 gnd.n1249 240.244
R4171 gnd.n1250 gnd.n1249 240.244
R4172 gnd.n4020 gnd.n1250 240.244
R4173 gnd.n4020 gnd.n243 240.244
R4174 gnd.n6574 gnd.n243 240.244
R4175 gnd.n6574 gnd.n238 240.244
R4176 gnd.n6580 gnd.n238 240.244
R4177 gnd.n6580 gnd.n229 240.244
R4178 gnd.n6588 gnd.n229 240.244
R4179 gnd.n6588 gnd.n225 240.244
R4180 gnd.n6594 gnd.n225 240.244
R4181 gnd.n6594 gnd.n208 240.244
R4182 gnd.n6604 gnd.n208 240.244
R4183 gnd.n6604 gnd.n204 240.244
R4184 gnd.n6610 gnd.n204 240.244
R4185 gnd.n6610 gnd.n193 240.244
R4186 gnd.n6620 gnd.n193 240.244
R4187 gnd.n6620 gnd.n189 240.244
R4188 gnd.n6626 gnd.n189 240.244
R4189 gnd.n6626 gnd.n178 240.244
R4190 gnd.n6636 gnd.n178 240.244
R4191 gnd.n6636 gnd.n172 240.244
R4192 gnd.n6716 gnd.n172 240.244
R4193 gnd.n6716 gnd.n173 240.244
R4194 gnd.n173 gnd.n163 240.244
R4195 gnd.n6641 gnd.n163 240.244
R4196 gnd.n6641 gnd.n84 240.244
R4197 gnd.n1920 gnd.n1083 240.244
R4198 gnd.n1921 gnd.n1870 240.244
R4199 gnd.n1924 gnd.n1871 240.244
R4200 gnd.n1880 gnd.n1879 240.244
R4201 gnd.n1926 gnd.n1887 240.244
R4202 gnd.n1929 gnd.n1888 240.244
R4203 gnd.n1898 gnd.n1897 240.244
R4204 gnd.n1931 gnd.n1905 240.244
R4205 gnd.n1917 gnd.n1906 240.244
R4206 gnd.n2166 gnd.n2085 240.244
R4207 gnd.n2167 gnd.n2166 240.244
R4208 gnd.n2167 gnd.n885 240.244
R4209 gnd.n2081 gnd.n885 240.244
R4210 gnd.n2081 gnd.n897 240.244
R4211 gnd.n2174 gnd.n897 240.244
R4212 gnd.n2174 gnd.n908 240.244
R4213 gnd.n2078 gnd.n908 240.244
R4214 gnd.n2078 gnd.n918 240.244
R4215 gnd.n2181 gnd.n918 240.244
R4216 gnd.n2181 gnd.n928 240.244
R4217 gnd.n2075 gnd.n928 240.244
R4218 gnd.n2075 gnd.n938 240.244
R4219 gnd.n2188 gnd.n938 240.244
R4220 gnd.n2188 gnd.n948 240.244
R4221 gnd.n2194 gnd.n948 240.244
R4222 gnd.n2234 gnd.n2194 240.244
R4223 gnd.n2234 gnd.n959 240.244
R4224 gnd.n2237 gnd.n959 240.244
R4225 gnd.n2237 gnd.n972 240.244
R4226 gnd.n2243 gnd.n972 240.244
R4227 gnd.n2243 gnd.n980 240.244
R4228 gnd.n2254 gnd.n980 240.244
R4229 gnd.n2254 gnd.n989 240.244
R4230 gnd.n2260 gnd.n989 240.244
R4231 gnd.n2260 gnd.n997 240.244
R4232 gnd.n2299 gnd.n997 240.244
R4233 gnd.n2299 gnd.n1007 240.244
R4234 gnd.n2027 gnd.n1007 240.244
R4235 gnd.n2027 gnd.n1018 240.244
R4236 gnd.n2028 gnd.n1018 240.244
R4237 gnd.n2028 gnd.n1028 240.244
R4238 gnd.n2287 gnd.n1028 240.244
R4239 gnd.n2287 gnd.n1039 240.244
R4240 gnd.n2362 gnd.n1039 240.244
R4241 gnd.n2362 gnd.n1049 240.244
R4242 gnd.n2368 gnd.n1049 240.244
R4243 gnd.n2368 gnd.n1060 240.244
R4244 gnd.n2379 gnd.n1060 240.244
R4245 gnd.n2379 gnd.n1071 240.244
R4246 gnd.n2417 gnd.n1071 240.244
R4247 gnd.n2417 gnd.n1081 240.244
R4248 gnd.n2146 gnd.n2145 240.244
R4249 gnd.n2142 gnd.n2141 240.244
R4250 gnd.n2138 gnd.n2137 240.244
R4251 gnd.n2134 gnd.n2133 240.244
R4252 gnd.n2130 gnd.n2129 240.244
R4253 gnd.n2126 gnd.n2125 240.244
R4254 gnd.n2122 gnd.n2121 240.244
R4255 gnd.n2118 gnd.n2117 240.244
R4256 gnd.n2105 gnd.n829 240.244
R4257 gnd.n2158 gnd.n2086 240.244
R4258 gnd.n2158 gnd.n2087 240.244
R4259 gnd.n2087 gnd.n887 240.244
R4260 gnd.n899 gnd.n887 240.244
R4261 gnd.n4312 gnd.n899 240.244
R4262 gnd.n4312 gnd.n900 240.244
R4263 gnd.n4308 gnd.n900 240.244
R4264 gnd.n4308 gnd.n906 240.244
R4265 gnd.n4300 gnd.n906 240.244
R4266 gnd.n4300 gnd.n919 240.244
R4267 gnd.n4296 gnd.n919 240.244
R4268 gnd.n4296 gnd.n925 240.244
R4269 gnd.n4288 gnd.n925 240.244
R4270 gnd.n4288 gnd.n940 240.244
R4271 gnd.n4284 gnd.n940 240.244
R4272 gnd.n4284 gnd.n946 240.244
R4273 gnd.n961 gnd.n946 240.244
R4274 gnd.n4274 gnd.n961 240.244
R4275 gnd.n4274 gnd.n962 240.244
R4276 gnd.n4270 gnd.n962 240.244
R4277 gnd.n4270 gnd.n970 240.244
R4278 gnd.n4261 gnd.n970 240.244
R4279 gnd.n4261 gnd.n981 240.244
R4280 gnd.n4257 gnd.n981 240.244
R4281 gnd.n4257 gnd.n986 240.244
R4282 gnd.n4248 gnd.n986 240.244
R4283 gnd.n4248 gnd.n999 240.244
R4284 gnd.n4244 gnd.n999 240.244
R4285 gnd.n4244 gnd.n1005 240.244
R4286 gnd.n4236 gnd.n1005 240.244
R4287 gnd.n4236 gnd.n1019 240.244
R4288 gnd.n4232 gnd.n1019 240.244
R4289 gnd.n4232 gnd.n1025 240.244
R4290 gnd.n4224 gnd.n1025 240.244
R4291 gnd.n4224 gnd.n1041 240.244
R4292 gnd.n4220 gnd.n1041 240.244
R4293 gnd.n4220 gnd.n1047 240.244
R4294 gnd.n4212 gnd.n1047 240.244
R4295 gnd.n4212 gnd.n1062 240.244
R4296 gnd.n4208 gnd.n1062 240.244
R4297 gnd.n4208 gnd.n1068 240.244
R4298 gnd.n4200 gnd.n1068 240.244
R4299 gnd.n5990 gnd.n593 240.244
R4300 gnd.n5996 gnd.n593 240.244
R4301 gnd.n5996 gnd.n591 240.244
R4302 gnd.n6000 gnd.n591 240.244
R4303 gnd.n6000 gnd.n587 240.244
R4304 gnd.n6006 gnd.n587 240.244
R4305 gnd.n6006 gnd.n585 240.244
R4306 gnd.n6010 gnd.n585 240.244
R4307 gnd.n6010 gnd.n581 240.244
R4308 gnd.n6016 gnd.n581 240.244
R4309 gnd.n6016 gnd.n579 240.244
R4310 gnd.n6020 gnd.n579 240.244
R4311 gnd.n6020 gnd.n575 240.244
R4312 gnd.n6026 gnd.n575 240.244
R4313 gnd.n6026 gnd.n573 240.244
R4314 gnd.n6030 gnd.n573 240.244
R4315 gnd.n6030 gnd.n569 240.244
R4316 gnd.n6036 gnd.n569 240.244
R4317 gnd.n6036 gnd.n567 240.244
R4318 gnd.n6040 gnd.n567 240.244
R4319 gnd.n6040 gnd.n563 240.244
R4320 gnd.n6046 gnd.n563 240.244
R4321 gnd.n6046 gnd.n561 240.244
R4322 gnd.n6050 gnd.n561 240.244
R4323 gnd.n6050 gnd.n557 240.244
R4324 gnd.n6056 gnd.n557 240.244
R4325 gnd.n6056 gnd.n555 240.244
R4326 gnd.n6060 gnd.n555 240.244
R4327 gnd.n6060 gnd.n551 240.244
R4328 gnd.n6066 gnd.n551 240.244
R4329 gnd.n6066 gnd.n549 240.244
R4330 gnd.n6070 gnd.n549 240.244
R4331 gnd.n6070 gnd.n545 240.244
R4332 gnd.n6076 gnd.n545 240.244
R4333 gnd.n6076 gnd.n543 240.244
R4334 gnd.n6080 gnd.n543 240.244
R4335 gnd.n6080 gnd.n539 240.244
R4336 gnd.n6086 gnd.n539 240.244
R4337 gnd.n6086 gnd.n537 240.244
R4338 gnd.n6090 gnd.n537 240.244
R4339 gnd.n6090 gnd.n533 240.244
R4340 gnd.n6096 gnd.n533 240.244
R4341 gnd.n6096 gnd.n531 240.244
R4342 gnd.n6100 gnd.n531 240.244
R4343 gnd.n6100 gnd.n527 240.244
R4344 gnd.n6106 gnd.n527 240.244
R4345 gnd.n6106 gnd.n525 240.244
R4346 gnd.n6110 gnd.n525 240.244
R4347 gnd.n6110 gnd.n521 240.244
R4348 gnd.n6116 gnd.n521 240.244
R4349 gnd.n6116 gnd.n519 240.244
R4350 gnd.n6120 gnd.n519 240.244
R4351 gnd.n6120 gnd.n515 240.244
R4352 gnd.n6126 gnd.n515 240.244
R4353 gnd.n6126 gnd.n513 240.244
R4354 gnd.n6130 gnd.n513 240.244
R4355 gnd.n6130 gnd.n509 240.244
R4356 gnd.n6136 gnd.n509 240.244
R4357 gnd.n6136 gnd.n507 240.244
R4358 gnd.n6140 gnd.n507 240.244
R4359 gnd.n6140 gnd.n503 240.244
R4360 gnd.n6146 gnd.n503 240.244
R4361 gnd.n6146 gnd.n501 240.244
R4362 gnd.n6150 gnd.n501 240.244
R4363 gnd.n6150 gnd.n497 240.244
R4364 gnd.n6156 gnd.n497 240.244
R4365 gnd.n6156 gnd.n495 240.244
R4366 gnd.n6160 gnd.n495 240.244
R4367 gnd.n6160 gnd.n491 240.244
R4368 gnd.n6166 gnd.n491 240.244
R4369 gnd.n6166 gnd.n489 240.244
R4370 gnd.n6170 gnd.n489 240.244
R4371 gnd.n6170 gnd.n485 240.244
R4372 gnd.n6176 gnd.n485 240.244
R4373 gnd.n6176 gnd.n483 240.244
R4374 gnd.n6180 gnd.n483 240.244
R4375 gnd.n6180 gnd.n479 240.244
R4376 gnd.n6186 gnd.n479 240.244
R4377 gnd.n6186 gnd.n477 240.244
R4378 gnd.n6190 gnd.n477 240.244
R4379 gnd.n6190 gnd.n473 240.244
R4380 gnd.n6196 gnd.n473 240.244
R4381 gnd.n6196 gnd.n471 240.244
R4382 gnd.n6200 gnd.n471 240.244
R4383 gnd.n6200 gnd.n467 240.244
R4384 gnd.n6206 gnd.n467 240.244
R4385 gnd.n6206 gnd.n465 240.244
R4386 gnd.n6210 gnd.n465 240.244
R4387 gnd.n6210 gnd.n461 240.244
R4388 gnd.n6216 gnd.n461 240.244
R4389 gnd.n6216 gnd.n459 240.244
R4390 gnd.n6220 gnd.n459 240.244
R4391 gnd.n6220 gnd.n455 240.244
R4392 gnd.n6226 gnd.n455 240.244
R4393 gnd.n6226 gnd.n453 240.244
R4394 gnd.n6230 gnd.n453 240.244
R4395 gnd.n6230 gnd.n449 240.244
R4396 gnd.n6236 gnd.n449 240.244
R4397 gnd.n6236 gnd.n447 240.244
R4398 gnd.n6240 gnd.n447 240.244
R4399 gnd.n6240 gnd.n443 240.244
R4400 gnd.n6246 gnd.n443 240.244
R4401 gnd.n6246 gnd.n441 240.244
R4402 gnd.n6250 gnd.n441 240.244
R4403 gnd.n6250 gnd.n437 240.244
R4404 gnd.n6256 gnd.n437 240.244
R4405 gnd.n6256 gnd.n435 240.244
R4406 gnd.n6260 gnd.n435 240.244
R4407 gnd.n6260 gnd.n431 240.244
R4408 gnd.n6266 gnd.n431 240.244
R4409 gnd.n6266 gnd.n429 240.244
R4410 gnd.n6270 gnd.n429 240.244
R4411 gnd.n6270 gnd.n425 240.244
R4412 gnd.n6276 gnd.n425 240.244
R4413 gnd.n6276 gnd.n423 240.244
R4414 gnd.n6280 gnd.n423 240.244
R4415 gnd.n6280 gnd.n419 240.244
R4416 gnd.n6286 gnd.n419 240.244
R4417 gnd.n6286 gnd.n417 240.244
R4418 gnd.n6290 gnd.n417 240.244
R4419 gnd.n6290 gnd.n413 240.244
R4420 gnd.n6296 gnd.n413 240.244
R4421 gnd.n6296 gnd.n411 240.244
R4422 gnd.n6300 gnd.n411 240.244
R4423 gnd.n6300 gnd.n407 240.244
R4424 gnd.n6306 gnd.n407 240.244
R4425 gnd.n6306 gnd.n405 240.244
R4426 gnd.n6310 gnd.n405 240.244
R4427 gnd.n6310 gnd.n401 240.244
R4428 gnd.n6316 gnd.n401 240.244
R4429 gnd.n6316 gnd.n399 240.244
R4430 gnd.n6320 gnd.n399 240.244
R4431 gnd.n6320 gnd.n395 240.244
R4432 gnd.n6326 gnd.n395 240.244
R4433 gnd.n6326 gnd.n393 240.244
R4434 gnd.n6330 gnd.n393 240.244
R4435 gnd.n6330 gnd.n389 240.244
R4436 gnd.n6337 gnd.n389 240.244
R4437 gnd.n6337 gnd.n387 240.244
R4438 gnd.n6341 gnd.n387 240.244
R4439 gnd.n6341 gnd.n384 240.244
R4440 gnd.n6347 gnd.n382 240.244
R4441 gnd.n6351 gnd.n382 240.244
R4442 gnd.n6351 gnd.n378 240.244
R4443 gnd.n6357 gnd.n378 240.244
R4444 gnd.n6357 gnd.n376 240.244
R4445 gnd.n6361 gnd.n376 240.244
R4446 gnd.n6361 gnd.n372 240.244
R4447 gnd.n6367 gnd.n372 240.244
R4448 gnd.n6367 gnd.n370 240.244
R4449 gnd.n6371 gnd.n370 240.244
R4450 gnd.n6371 gnd.n366 240.244
R4451 gnd.n6377 gnd.n366 240.244
R4452 gnd.n6377 gnd.n364 240.244
R4453 gnd.n6381 gnd.n364 240.244
R4454 gnd.n6381 gnd.n360 240.244
R4455 gnd.n6387 gnd.n360 240.244
R4456 gnd.n6387 gnd.n358 240.244
R4457 gnd.n6391 gnd.n358 240.244
R4458 gnd.n6391 gnd.n354 240.244
R4459 gnd.n6397 gnd.n354 240.244
R4460 gnd.n6397 gnd.n352 240.244
R4461 gnd.n6401 gnd.n352 240.244
R4462 gnd.n6401 gnd.n348 240.244
R4463 gnd.n6407 gnd.n348 240.244
R4464 gnd.n6407 gnd.n346 240.244
R4465 gnd.n6411 gnd.n346 240.244
R4466 gnd.n6411 gnd.n342 240.244
R4467 gnd.n6417 gnd.n342 240.244
R4468 gnd.n6417 gnd.n340 240.244
R4469 gnd.n6421 gnd.n340 240.244
R4470 gnd.n6421 gnd.n336 240.244
R4471 gnd.n6427 gnd.n336 240.244
R4472 gnd.n6427 gnd.n334 240.244
R4473 gnd.n6431 gnd.n334 240.244
R4474 gnd.n6431 gnd.n330 240.244
R4475 gnd.n6437 gnd.n330 240.244
R4476 gnd.n6437 gnd.n328 240.244
R4477 gnd.n6441 gnd.n328 240.244
R4478 gnd.n6441 gnd.n324 240.244
R4479 gnd.n6447 gnd.n324 240.244
R4480 gnd.n6447 gnd.n322 240.244
R4481 gnd.n6451 gnd.n322 240.244
R4482 gnd.n6451 gnd.n318 240.244
R4483 gnd.n6457 gnd.n318 240.244
R4484 gnd.n6457 gnd.n316 240.244
R4485 gnd.n6461 gnd.n316 240.244
R4486 gnd.n6461 gnd.n312 240.244
R4487 gnd.n6467 gnd.n312 240.244
R4488 gnd.n6467 gnd.n310 240.244
R4489 gnd.n6471 gnd.n310 240.244
R4490 gnd.n6471 gnd.n306 240.244
R4491 gnd.n6477 gnd.n306 240.244
R4492 gnd.n6477 gnd.n304 240.244
R4493 gnd.n6481 gnd.n304 240.244
R4494 gnd.n6481 gnd.n300 240.244
R4495 gnd.n6487 gnd.n300 240.244
R4496 gnd.n6487 gnd.n298 240.244
R4497 gnd.n6491 gnd.n298 240.244
R4498 gnd.n6491 gnd.n294 240.244
R4499 gnd.n6497 gnd.n294 240.244
R4500 gnd.n6497 gnd.n292 240.244
R4501 gnd.n6501 gnd.n292 240.244
R4502 gnd.n6501 gnd.n288 240.244
R4503 gnd.n6507 gnd.n288 240.244
R4504 gnd.n6507 gnd.n286 240.244
R4505 gnd.n6511 gnd.n286 240.244
R4506 gnd.n6511 gnd.n282 240.244
R4507 gnd.n6517 gnd.n282 240.244
R4508 gnd.n6517 gnd.n280 240.244
R4509 gnd.n6521 gnd.n280 240.244
R4510 gnd.n6521 gnd.n276 240.244
R4511 gnd.n6527 gnd.n276 240.244
R4512 gnd.n6527 gnd.n274 240.244
R4513 gnd.n6531 gnd.n274 240.244
R4514 gnd.n6531 gnd.n270 240.244
R4515 gnd.n6537 gnd.n270 240.244
R4516 gnd.n6537 gnd.n268 240.244
R4517 gnd.n6541 gnd.n268 240.244
R4518 gnd.n6541 gnd.n264 240.244
R4519 gnd.n6547 gnd.n264 240.244
R4520 gnd.n6547 gnd.n262 240.244
R4521 gnd.n6552 gnd.n262 240.244
R4522 gnd.n6552 gnd.n258 240.244
R4523 gnd.n6559 gnd.n258 240.244
R4524 gnd.n2047 gnd.n2046 240.244
R4525 gnd.n2047 gnd.n2039 240.244
R4526 gnd.n2065 gnd.n2039 240.244
R4527 gnd.n2065 gnd.n2040 240.244
R4528 gnd.n2061 gnd.n2040 240.244
R4529 gnd.n2061 gnd.n2060 240.244
R4530 gnd.n2060 gnd.n2020 240.244
R4531 gnd.n2302 gnd.n2020 240.244
R4532 gnd.n2303 gnd.n2302 240.244
R4533 gnd.n2304 gnd.n2303 240.244
R4534 gnd.n2304 gnd.n2016 240.244
R4535 gnd.n2310 gnd.n2016 240.244
R4536 gnd.n2311 gnd.n2310 240.244
R4537 gnd.n2312 gnd.n2311 240.244
R4538 gnd.n2312 gnd.n2011 240.244
R4539 gnd.n2359 gnd.n2011 240.244
R4540 gnd.n2359 gnd.n2012 240.244
R4541 gnd.n2355 gnd.n2012 240.244
R4542 gnd.n2355 gnd.n2354 240.244
R4543 gnd.n2354 gnd.n2353 240.244
R4544 gnd.n2353 gnd.n2320 240.244
R4545 gnd.n2349 gnd.n2320 240.244
R4546 gnd.n2349 gnd.n2348 240.244
R4547 gnd.n2348 gnd.n2347 240.244
R4548 gnd.n2347 gnd.n2326 240.244
R4549 gnd.n2343 gnd.n2326 240.244
R4550 gnd.n2343 gnd.n2341 240.244
R4551 gnd.n2341 gnd.n2340 240.244
R4552 gnd.n2340 gnd.n2334 240.244
R4553 gnd.n2334 gnd.n1842 240.244
R4554 gnd.n2687 gnd.n1842 240.244
R4555 gnd.n2687 gnd.n1838 240.244
R4556 gnd.n2693 gnd.n1838 240.244
R4557 gnd.n2693 gnd.n1829 240.244
R4558 gnd.n2707 gnd.n1829 240.244
R4559 gnd.n2707 gnd.n1825 240.244
R4560 gnd.n2713 gnd.n1825 240.244
R4561 gnd.n2713 gnd.n1816 240.244
R4562 gnd.n2728 gnd.n1816 240.244
R4563 gnd.n2728 gnd.n1811 240.244
R4564 gnd.n2736 gnd.n1811 240.244
R4565 gnd.n2736 gnd.n1812 240.244
R4566 gnd.n1812 gnd.n1739 240.244
R4567 gnd.n2805 gnd.n1739 240.244
R4568 gnd.n2805 gnd.n1734 240.244
R4569 gnd.n2813 gnd.n1734 240.244
R4570 gnd.n2813 gnd.n1735 240.244
R4571 gnd.n1735 gnd.n1711 240.244
R4572 gnd.n2842 gnd.n1711 240.244
R4573 gnd.n2842 gnd.n1707 240.244
R4574 gnd.n2848 gnd.n1707 240.244
R4575 gnd.n2848 gnd.n1689 240.244
R4576 gnd.n2869 gnd.n1689 240.244
R4577 gnd.n2869 gnd.n1684 240.244
R4578 gnd.n2877 gnd.n1684 240.244
R4579 gnd.n2877 gnd.n1685 240.244
R4580 gnd.n1685 gnd.n1656 240.244
R4581 gnd.n2911 gnd.n1656 240.244
R4582 gnd.n2911 gnd.n1651 240.244
R4583 gnd.n2928 gnd.n1651 240.244
R4584 gnd.n2928 gnd.n1652 240.244
R4585 gnd.n2924 gnd.n1652 240.244
R4586 gnd.n2924 gnd.n2920 240.244
R4587 gnd.n2920 gnd.n1622 240.244
R4588 gnd.n2994 gnd.n1622 240.244
R4589 gnd.n2994 gnd.n1618 240.244
R4590 gnd.n3000 gnd.n1618 240.244
R4591 gnd.n3000 gnd.n1599 240.244
R4592 gnd.n3037 gnd.n1599 240.244
R4593 gnd.n3037 gnd.n1595 240.244
R4594 gnd.n3043 gnd.n1595 240.244
R4595 gnd.n3043 gnd.n1583 240.244
R4596 gnd.n3081 gnd.n1583 240.244
R4597 gnd.n3081 gnd.n1578 240.244
R4598 gnd.n3089 gnd.n1578 240.244
R4599 gnd.n3089 gnd.n1579 240.244
R4600 gnd.n1579 gnd.n1552 240.244
R4601 gnd.n3127 gnd.n1552 240.244
R4602 gnd.n3127 gnd.n1548 240.244
R4603 gnd.n3133 gnd.n1548 240.244
R4604 gnd.n3133 gnd.n1535 240.244
R4605 gnd.n3188 gnd.n1535 240.244
R4606 gnd.n3188 gnd.n1531 240.244
R4607 gnd.n3194 gnd.n1531 240.244
R4608 gnd.n3194 gnd.n1513 240.244
R4609 gnd.n3216 gnd.n1513 240.244
R4610 gnd.n3216 gnd.n1508 240.244
R4611 gnd.n3224 gnd.n1508 240.244
R4612 gnd.n3224 gnd.n1509 240.244
R4613 gnd.n1509 gnd.n1485 240.244
R4614 gnd.n3260 gnd.n1485 240.244
R4615 gnd.n3260 gnd.n1480 240.244
R4616 gnd.n3272 gnd.n1480 240.244
R4617 gnd.n3272 gnd.n1481 240.244
R4618 gnd.n3268 gnd.n1481 240.244
R4619 gnd.n3268 gnd.n1412 240.244
R4620 gnd.n3534 gnd.n1412 240.244
R4621 gnd.n3534 gnd.n1413 240.244
R4622 gnd.n3530 gnd.n1413 240.244
R4623 gnd.n3530 gnd.n1419 240.244
R4624 gnd.n3523 gnd.n1419 240.244
R4625 gnd.n3523 gnd.n1423 240.244
R4626 gnd.n3519 gnd.n1423 240.244
R4627 gnd.n3519 gnd.n1429 240.244
R4628 gnd.n3512 gnd.n1429 240.244
R4629 gnd.n3512 gnd.n1434 240.244
R4630 gnd.n3508 gnd.n1434 240.244
R4631 gnd.n3508 gnd.n1440 240.244
R4632 gnd.n3501 gnd.n1440 240.244
R4633 gnd.n3501 gnd.n3494 240.244
R4634 gnd.n3494 gnd.n1195 240.244
R4635 gnd.n4068 gnd.n1195 240.244
R4636 gnd.n4068 gnd.n1196 240.244
R4637 gnd.n4064 gnd.n1196 240.244
R4638 gnd.n4064 gnd.n1202 240.244
R4639 gnd.n4060 gnd.n1202 240.244
R4640 gnd.n4060 gnd.n1205 240.244
R4641 gnd.n4056 gnd.n1205 240.244
R4642 gnd.n4056 gnd.n1211 240.244
R4643 gnd.n3923 gnd.n1211 240.244
R4644 gnd.n3924 gnd.n3923 240.244
R4645 gnd.n3924 gnd.n3917 240.244
R4646 gnd.n3932 gnd.n3917 240.244
R4647 gnd.n3932 gnd.n3918 240.244
R4648 gnd.n3918 gnd.n1308 240.244
R4649 gnd.n3955 gnd.n1308 240.244
R4650 gnd.n3955 gnd.n1303 240.244
R4651 gnd.n3963 gnd.n1303 240.244
R4652 gnd.n3963 gnd.n1304 240.244
R4653 gnd.n1304 gnd.n1280 240.244
R4654 gnd.n3987 gnd.n1280 240.244
R4655 gnd.n3987 gnd.n1275 240.244
R4656 gnd.n4002 gnd.n1275 240.244
R4657 gnd.n4002 gnd.n1276 240.244
R4658 gnd.n3993 gnd.n1276 240.244
R4659 gnd.n3994 gnd.n3993 240.244
R4660 gnd.n3994 gnd.n251 240.244
R4661 gnd.n6566 gnd.n251 240.244
R4662 gnd.n6566 gnd.n252 240.244
R4663 gnd.n6562 gnd.n252 240.244
R4664 gnd.n6562 gnd.n6561 240.244
R4665 gnd.n5986 gnd.n596 240.244
R4666 gnd.n5986 gnd.n598 240.244
R4667 gnd.n5982 gnd.n598 240.244
R4668 gnd.n5982 gnd.n604 240.244
R4669 gnd.n5978 gnd.n604 240.244
R4670 gnd.n5978 gnd.n606 240.244
R4671 gnd.n5974 gnd.n606 240.244
R4672 gnd.n5974 gnd.n612 240.244
R4673 gnd.n5970 gnd.n612 240.244
R4674 gnd.n5970 gnd.n614 240.244
R4675 gnd.n5966 gnd.n614 240.244
R4676 gnd.n5966 gnd.n620 240.244
R4677 gnd.n5962 gnd.n620 240.244
R4678 gnd.n5962 gnd.n622 240.244
R4679 gnd.n5958 gnd.n622 240.244
R4680 gnd.n5958 gnd.n628 240.244
R4681 gnd.n5954 gnd.n628 240.244
R4682 gnd.n5954 gnd.n630 240.244
R4683 gnd.n5950 gnd.n630 240.244
R4684 gnd.n5950 gnd.n636 240.244
R4685 gnd.n5946 gnd.n636 240.244
R4686 gnd.n5946 gnd.n638 240.244
R4687 gnd.n5942 gnd.n638 240.244
R4688 gnd.n5942 gnd.n644 240.244
R4689 gnd.n5938 gnd.n644 240.244
R4690 gnd.n5938 gnd.n646 240.244
R4691 gnd.n5934 gnd.n646 240.244
R4692 gnd.n5934 gnd.n652 240.244
R4693 gnd.n5930 gnd.n652 240.244
R4694 gnd.n5930 gnd.n654 240.244
R4695 gnd.n5926 gnd.n654 240.244
R4696 gnd.n5926 gnd.n660 240.244
R4697 gnd.n5922 gnd.n660 240.244
R4698 gnd.n5922 gnd.n662 240.244
R4699 gnd.n5918 gnd.n662 240.244
R4700 gnd.n5918 gnd.n668 240.244
R4701 gnd.n5914 gnd.n668 240.244
R4702 gnd.n5914 gnd.n670 240.244
R4703 gnd.n5910 gnd.n670 240.244
R4704 gnd.n5910 gnd.n676 240.244
R4705 gnd.n5906 gnd.n676 240.244
R4706 gnd.n5906 gnd.n678 240.244
R4707 gnd.n5902 gnd.n678 240.244
R4708 gnd.n5902 gnd.n684 240.244
R4709 gnd.n5898 gnd.n684 240.244
R4710 gnd.n5898 gnd.n686 240.244
R4711 gnd.n5894 gnd.n686 240.244
R4712 gnd.n5894 gnd.n692 240.244
R4713 gnd.n5890 gnd.n692 240.244
R4714 gnd.n5890 gnd.n694 240.244
R4715 gnd.n5886 gnd.n694 240.244
R4716 gnd.n5886 gnd.n700 240.244
R4717 gnd.n5882 gnd.n700 240.244
R4718 gnd.n5882 gnd.n702 240.244
R4719 gnd.n5878 gnd.n702 240.244
R4720 gnd.n5878 gnd.n708 240.244
R4721 gnd.n5874 gnd.n708 240.244
R4722 gnd.n5874 gnd.n710 240.244
R4723 gnd.n5870 gnd.n710 240.244
R4724 gnd.n5870 gnd.n716 240.244
R4725 gnd.n5866 gnd.n716 240.244
R4726 gnd.n5866 gnd.n718 240.244
R4727 gnd.n5862 gnd.n718 240.244
R4728 gnd.n5862 gnd.n724 240.244
R4729 gnd.n5858 gnd.n724 240.244
R4730 gnd.n5858 gnd.n726 240.244
R4731 gnd.n5854 gnd.n726 240.244
R4732 gnd.n5854 gnd.n732 240.244
R4733 gnd.n5850 gnd.n732 240.244
R4734 gnd.n5850 gnd.n734 240.244
R4735 gnd.n5846 gnd.n734 240.244
R4736 gnd.n5846 gnd.n740 240.244
R4737 gnd.n5842 gnd.n740 240.244
R4738 gnd.n5842 gnd.n742 240.244
R4739 gnd.n5838 gnd.n742 240.244
R4740 gnd.n5838 gnd.n748 240.244
R4741 gnd.n5834 gnd.n748 240.244
R4742 gnd.n5834 gnd.n750 240.244
R4743 gnd.n5830 gnd.n750 240.244
R4744 gnd.n5830 gnd.n756 240.244
R4745 gnd.n5826 gnd.n756 240.244
R4746 gnd.n5826 gnd.n758 240.244
R4747 gnd.n5822 gnd.n758 240.244
R4748 gnd.n5822 gnd.n764 240.244
R4749 gnd.n1089 gnd.n1088 240.244
R4750 gnd.n1090 gnd.n1089 240.244
R4751 gnd.n2695 gnd.n1090 240.244
R4752 gnd.n2695 gnd.n1093 240.244
R4753 gnd.n1094 gnd.n1093 240.244
R4754 gnd.n1095 gnd.n1094 240.244
R4755 gnd.n2715 gnd.n1095 240.244
R4756 gnd.n2715 gnd.n1098 240.244
R4757 gnd.n1099 gnd.n1098 240.244
R4758 gnd.n1100 gnd.n1099 240.244
R4759 gnd.n2738 gnd.n1100 240.244
R4760 gnd.n2738 gnd.n1103 240.244
R4761 gnd.n1104 gnd.n1103 240.244
R4762 gnd.n1105 gnd.n1104 240.244
R4763 gnd.n2802 gnd.n1105 240.244
R4764 gnd.n2802 gnd.n1108 240.244
R4765 gnd.n1109 gnd.n1108 240.244
R4766 gnd.n1110 gnd.n1109 240.244
R4767 gnd.n2832 gnd.n1110 240.244
R4768 gnd.n2832 gnd.n1113 240.244
R4769 gnd.n1114 gnd.n1113 240.244
R4770 gnd.n1115 gnd.n1114 240.244
R4771 gnd.n1699 gnd.n1115 240.244
R4772 gnd.n1699 gnd.n1118 240.244
R4773 gnd.n1119 gnd.n1118 240.244
R4774 gnd.n1120 gnd.n1119 240.244
R4775 gnd.n1666 gnd.n1120 240.244
R4776 gnd.n1666 gnd.n1123 240.244
R4777 gnd.n1124 gnd.n1123 240.244
R4778 gnd.n1125 gnd.n1124 240.244
R4779 gnd.n2938 gnd.n1125 240.244
R4780 gnd.n2938 gnd.n1128 240.244
R4781 gnd.n1129 gnd.n1128 240.244
R4782 gnd.n1130 gnd.n1129 240.244
R4783 gnd.n1623 gnd.n1130 240.244
R4784 gnd.n1623 gnd.n1133 240.244
R4785 gnd.n1134 gnd.n1133 240.244
R4786 gnd.n1135 gnd.n1134 240.244
R4787 gnd.n3022 gnd.n1135 240.244
R4788 gnd.n3022 gnd.n1138 240.244
R4789 gnd.n1139 gnd.n1138 240.244
R4790 gnd.n1140 gnd.n1139 240.244
R4791 gnd.n3070 gnd.n1140 240.244
R4792 gnd.n3070 gnd.n1143 240.244
R4793 gnd.n1144 gnd.n1143 240.244
R4794 gnd.n1145 gnd.n1144 240.244
R4795 gnd.n3053 gnd.n1145 240.244
R4796 gnd.n3053 gnd.n1148 240.244
R4797 gnd.n1149 gnd.n1148 240.244
R4798 gnd.n1150 gnd.n1149 240.244
R4799 gnd.n1542 gnd.n1150 240.244
R4800 gnd.n1542 gnd.n1153 240.244
R4801 gnd.n1154 gnd.n1153 240.244
R4802 gnd.n1155 gnd.n1154 240.244
R4803 gnd.n1519 gnd.n1155 240.244
R4804 gnd.n1519 gnd.n1158 240.244
R4805 gnd.n1159 gnd.n1158 240.244
R4806 gnd.n1160 gnd.n1159 240.244
R4807 gnd.n3233 gnd.n1160 240.244
R4808 gnd.n3233 gnd.n1163 240.244
R4809 gnd.n1164 gnd.n1163 240.244
R4810 gnd.n1165 gnd.n1164 240.244
R4811 gnd.n1475 gnd.n1165 240.244
R4812 gnd.n1475 gnd.n1168 240.244
R4813 gnd.n1169 gnd.n1168 240.244
R4814 gnd.n1170 gnd.n1169 240.244
R4815 gnd.n3536 gnd.n1170 240.244
R4816 gnd.n3536 gnd.n1173 240.244
R4817 gnd.n1174 gnd.n1173 240.244
R4818 gnd.n1175 gnd.n1174 240.244
R4819 gnd.n3525 gnd.n1175 240.244
R4820 gnd.n3525 gnd.n1178 240.244
R4821 gnd.n1179 gnd.n1178 240.244
R4822 gnd.n1180 gnd.n1179 240.244
R4823 gnd.n3514 gnd.n1180 240.244
R4824 gnd.n3514 gnd.n1183 240.244
R4825 gnd.n1184 gnd.n1183 240.244
R4826 gnd.n1185 gnd.n1184 240.244
R4827 gnd.n3503 gnd.n1185 240.244
R4828 gnd.n3503 gnd.n1188 240.244
R4829 gnd.n1189 gnd.n1188 240.244
R4830 gnd.n4071 gnd.n1189 240.244
R4831 gnd.n1864 gnd.n1863 240.244
R4832 gnd.n1874 gnd.n1863 240.244
R4833 gnd.n1876 gnd.n1875 240.244
R4834 gnd.n1884 gnd.n1883 240.244
R4835 gnd.n1892 gnd.n1891 240.244
R4836 gnd.n1894 gnd.n1893 240.244
R4837 gnd.n1902 gnd.n1901 240.244
R4838 gnd.n1912 gnd.n1911 240.244
R4839 gnd.n1914 gnd.n1913 240.244
R4840 gnd.n2385 gnd.n2384 240.244
R4841 gnd.n2387 gnd.n2386 240.244
R4842 gnd.n2391 gnd.n2390 240.244
R4843 gnd.n2397 gnd.n2392 240.244
R4844 gnd.n2398 gnd.n1848 240.244
R4845 gnd.n2683 gnd.n1844 240.244
R4846 gnd.n2683 gnd.n1835 240.244
R4847 gnd.n2697 gnd.n1835 240.244
R4848 gnd.n2697 gnd.n1831 240.244
R4849 gnd.n2703 gnd.n1831 240.244
R4850 gnd.n2703 gnd.n1822 240.244
R4851 gnd.n2717 gnd.n1822 240.244
R4852 gnd.n2717 gnd.n1818 240.244
R4853 gnd.n2723 gnd.n1818 240.244
R4854 gnd.n2723 gnd.n1809 240.244
R4855 gnd.n2740 gnd.n1809 240.244
R4856 gnd.n2740 gnd.n1803 240.244
R4857 gnd.n2749 gnd.n1803 240.244
R4858 gnd.n2749 gnd.n1804 240.244
R4859 gnd.n1804 gnd.n1741 240.244
R4860 gnd.n1741 gnd.n1726 240.244
R4861 gnd.n2824 gnd.n1726 240.244
R4862 gnd.n2824 gnd.n1720 240.244
R4863 gnd.n2831 gnd.n1720 240.244
R4864 gnd.n2831 gnd.n1721 240.244
R4865 gnd.n1721 gnd.n1696 240.244
R4866 gnd.n2860 gnd.n1696 240.244
R4867 gnd.n2860 gnd.n1692 240.244
R4868 gnd.n2866 gnd.n1692 240.244
R4869 gnd.n2866 gnd.n1675 240.244
R4870 gnd.n2889 gnd.n1675 240.244
R4871 gnd.n2889 gnd.n1669 240.244
R4872 gnd.n2899 gnd.n1669 240.244
R4873 gnd.n2899 gnd.n1670 240.244
R4874 gnd.n2893 gnd.n1670 240.244
R4875 gnd.n2893 gnd.n1640 240.244
R4876 gnd.n2949 gnd.n1640 240.244
R4877 gnd.n2949 gnd.n1634 240.244
R4878 gnd.n2956 gnd.n1634 240.244
R4879 gnd.n2956 gnd.n1635 240.244
R4880 gnd.n1635 gnd.n1615 240.244
R4881 gnd.n3003 gnd.n1615 240.244
R4882 gnd.n3003 gnd.n1609 240.244
R4883 gnd.n3021 gnd.n1609 240.244
R4884 gnd.n3021 gnd.n1610 240.244
R4885 gnd.n3008 gnd.n1610 240.244
R4886 gnd.n3009 gnd.n3008 240.244
R4887 gnd.n3009 gnd.n1591 240.244
R4888 gnd.n3010 gnd.n1591 240.244
R4889 gnd.n3010 gnd.n1569 240.244
R4890 gnd.n3099 gnd.n1569 240.244
R4891 gnd.n3099 gnd.n1564 240.244
R4892 gnd.n3115 gnd.n1564 240.244
R4893 gnd.n3115 gnd.n1554 240.244
R4894 gnd.n3104 gnd.n1554 240.244
R4895 gnd.n3105 gnd.n3104 240.244
R4896 gnd.n3106 gnd.n3105 240.244
R4897 gnd.n3106 gnd.n1529 240.244
R4898 gnd.n3197 gnd.n1529 240.244
R4899 gnd.n3197 gnd.n1523 240.244
R4900 gnd.n3204 gnd.n1523 240.244
R4901 gnd.n3204 gnd.n1524 240.244
R4902 gnd.n1524 gnd.n1500 240.244
R4903 gnd.n3235 gnd.n1500 240.244
R4904 gnd.n3235 gnd.n1495 240.244
R4905 gnd.n3249 gnd.n1495 240.244
R4906 gnd.n3249 gnd.n1487 240.244
R4907 gnd.n3241 gnd.n1487 240.244
R4908 gnd.n3242 gnd.n3241 240.244
R4909 gnd.n3242 gnd.n1464 240.244
R4910 gnd.n3290 gnd.n1464 240.244
R4911 gnd.n3290 gnd.n1410 240.244
R4912 gnd.n1460 gnd.n1410 240.244
R4913 gnd.n1461 gnd.n1460 240.244
R4914 gnd.n1461 gnd.n1420 240.244
R4915 gnd.n1421 gnd.n1420 240.244
R4916 gnd.n1456 gnd.n1421 240.244
R4917 gnd.n1457 gnd.n1456 240.244
R4918 gnd.n1457 gnd.n1432 240.244
R4919 gnd.n1433 gnd.n1432 240.244
R4920 gnd.n1452 gnd.n1433 240.244
R4921 gnd.n1453 gnd.n1452 240.244
R4922 gnd.n1453 gnd.n1442 240.244
R4923 gnd.n1443 gnd.n1442 240.244
R4924 gnd.n1445 gnd.n1443 240.244
R4925 gnd.n3491 gnd.n1445 240.244
R4926 gnd.n3491 gnd.n1193 240.244
R4927 gnd.n3382 gnd.n3381 240.244
R4928 gnd.n3385 gnd.n3384 240.244
R4929 gnd.n3401 gnd.n3400 240.244
R4930 gnd.n3404 gnd.n3403 240.244
R4931 gnd.n3420 gnd.n3419 240.244
R4932 gnd.n3423 gnd.n3422 240.244
R4933 gnd.n3439 gnd.n3438 240.244
R4934 gnd.n3443 gnd.n3441 240.244
R4935 gnd.n3459 gnd.n3323 240.244
R4936 gnd.n3463 gnd.n3461 240.244
R4937 gnd.n3469 gnd.n3319 240.244
R4938 gnd.n3473 gnd.n3471 240.244
R4939 gnd.n3482 gnd.n3315 240.244
R4940 gnd.n3485 gnd.n3484 240.244
R4941 gnd.n1754 gnd.n1753 240.132
R4942 gnd.n3553 gnd.n3552 240.132
R4943 gnd.n5989 gnd.n592 225.874
R4944 gnd.n5997 gnd.n592 225.874
R4945 gnd.n5998 gnd.n5997 225.874
R4946 gnd.n5999 gnd.n5998 225.874
R4947 gnd.n5999 gnd.n586 225.874
R4948 gnd.n6007 gnd.n586 225.874
R4949 gnd.n6008 gnd.n6007 225.874
R4950 gnd.n6009 gnd.n6008 225.874
R4951 gnd.n6009 gnd.n580 225.874
R4952 gnd.n6017 gnd.n580 225.874
R4953 gnd.n6018 gnd.n6017 225.874
R4954 gnd.n6019 gnd.n6018 225.874
R4955 gnd.n6019 gnd.n574 225.874
R4956 gnd.n6027 gnd.n574 225.874
R4957 gnd.n6028 gnd.n6027 225.874
R4958 gnd.n6029 gnd.n6028 225.874
R4959 gnd.n6029 gnd.n568 225.874
R4960 gnd.n6037 gnd.n568 225.874
R4961 gnd.n6038 gnd.n6037 225.874
R4962 gnd.n6039 gnd.n6038 225.874
R4963 gnd.n6039 gnd.n562 225.874
R4964 gnd.n6047 gnd.n562 225.874
R4965 gnd.n6048 gnd.n6047 225.874
R4966 gnd.n6049 gnd.n6048 225.874
R4967 gnd.n6049 gnd.n556 225.874
R4968 gnd.n6057 gnd.n556 225.874
R4969 gnd.n6058 gnd.n6057 225.874
R4970 gnd.n6059 gnd.n6058 225.874
R4971 gnd.n6059 gnd.n550 225.874
R4972 gnd.n6067 gnd.n550 225.874
R4973 gnd.n6068 gnd.n6067 225.874
R4974 gnd.n6069 gnd.n6068 225.874
R4975 gnd.n6069 gnd.n544 225.874
R4976 gnd.n6077 gnd.n544 225.874
R4977 gnd.n6078 gnd.n6077 225.874
R4978 gnd.n6079 gnd.n6078 225.874
R4979 gnd.n6079 gnd.n538 225.874
R4980 gnd.n6087 gnd.n538 225.874
R4981 gnd.n6088 gnd.n6087 225.874
R4982 gnd.n6089 gnd.n6088 225.874
R4983 gnd.n6089 gnd.n532 225.874
R4984 gnd.n6097 gnd.n532 225.874
R4985 gnd.n6098 gnd.n6097 225.874
R4986 gnd.n6099 gnd.n6098 225.874
R4987 gnd.n6099 gnd.n526 225.874
R4988 gnd.n6107 gnd.n526 225.874
R4989 gnd.n6108 gnd.n6107 225.874
R4990 gnd.n6109 gnd.n6108 225.874
R4991 gnd.n6109 gnd.n520 225.874
R4992 gnd.n6117 gnd.n520 225.874
R4993 gnd.n6118 gnd.n6117 225.874
R4994 gnd.n6119 gnd.n6118 225.874
R4995 gnd.n6119 gnd.n514 225.874
R4996 gnd.n6127 gnd.n514 225.874
R4997 gnd.n6128 gnd.n6127 225.874
R4998 gnd.n6129 gnd.n6128 225.874
R4999 gnd.n6129 gnd.n508 225.874
R5000 gnd.n6137 gnd.n508 225.874
R5001 gnd.n6138 gnd.n6137 225.874
R5002 gnd.n6139 gnd.n6138 225.874
R5003 gnd.n6139 gnd.n502 225.874
R5004 gnd.n6147 gnd.n502 225.874
R5005 gnd.n6148 gnd.n6147 225.874
R5006 gnd.n6149 gnd.n6148 225.874
R5007 gnd.n6149 gnd.n496 225.874
R5008 gnd.n6157 gnd.n496 225.874
R5009 gnd.n6158 gnd.n6157 225.874
R5010 gnd.n6159 gnd.n6158 225.874
R5011 gnd.n6159 gnd.n490 225.874
R5012 gnd.n6167 gnd.n490 225.874
R5013 gnd.n6168 gnd.n6167 225.874
R5014 gnd.n6169 gnd.n6168 225.874
R5015 gnd.n6169 gnd.n484 225.874
R5016 gnd.n6177 gnd.n484 225.874
R5017 gnd.n6178 gnd.n6177 225.874
R5018 gnd.n6179 gnd.n6178 225.874
R5019 gnd.n6179 gnd.n478 225.874
R5020 gnd.n6187 gnd.n478 225.874
R5021 gnd.n6188 gnd.n6187 225.874
R5022 gnd.n6189 gnd.n6188 225.874
R5023 gnd.n6189 gnd.n472 225.874
R5024 gnd.n6197 gnd.n472 225.874
R5025 gnd.n6198 gnd.n6197 225.874
R5026 gnd.n6199 gnd.n6198 225.874
R5027 gnd.n6199 gnd.n466 225.874
R5028 gnd.n6207 gnd.n466 225.874
R5029 gnd.n6208 gnd.n6207 225.874
R5030 gnd.n6209 gnd.n6208 225.874
R5031 gnd.n6209 gnd.n460 225.874
R5032 gnd.n6217 gnd.n460 225.874
R5033 gnd.n6218 gnd.n6217 225.874
R5034 gnd.n6219 gnd.n6218 225.874
R5035 gnd.n6219 gnd.n454 225.874
R5036 gnd.n6227 gnd.n454 225.874
R5037 gnd.n6228 gnd.n6227 225.874
R5038 gnd.n6229 gnd.n6228 225.874
R5039 gnd.n6229 gnd.n448 225.874
R5040 gnd.n6237 gnd.n448 225.874
R5041 gnd.n6238 gnd.n6237 225.874
R5042 gnd.n6239 gnd.n6238 225.874
R5043 gnd.n6239 gnd.n442 225.874
R5044 gnd.n6247 gnd.n442 225.874
R5045 gnd.n6248 gnd.n6247 225.874
R5046 gnd.n6249 gnd.n6248 225.874
R5047 gnd.n6249 gnd.n436 225.874
R5048 gnd.n6257 gnd.n436 225.874
R5049 gnd.n6258 gnd.n6257 225.874
R5050 gnd.n6259 gnd.n6258 225.874
R5051 gnd.n6259 gnd.n430 225.874
R5052 gnd.n6267 gnd.n430 225.874
R5053 gnd.n6268 gnd.n6267 225.874
R5054 gnd.n6269 gnd.n6268 225.874
R5055 gnd.n6269 gnd.n424 225.874
R5056 gnd.n6277 gnd.n424 225.874
R5057 gnd.n6278 gnd.n6277 225.874
R5058 gnd.n6279 gnd.n6278 225.874
R5059 gnd.n6279 gnd.n418 225.874
R5060 gnd.n6287 gnd.n418 225.874
R5061 gnd.n6288 gnd.n6287 225.874
R5062 gnd.n6289 gnd.n6288 225.874
R5063 gnd.n6289 gnd.n412 225.874
R5064 gnd.n6297 gnd.n412 225.874
R5065 gnd.n6298 gnd.n6297 225.874
R5066 gnd.n6299 gnd.n6298 225.874
R5067 gnd.n6299 gnd.n406 225.874
R5068 gnd.n6307 gnd.n406 225.874
R5069 gnd.n6308 gnd.n6307 225.874
R5070 gnd.n6309 gnd.n6308 225.874
R5071 gnd.n6309 gnd.n400 225.874
R5072 gnd.n6317 gnd.n400 225.874
R5073 gnd.n6318 gnd.n6317 225.874
R5074 gnd.n6319 gnd.n6318 225.874
R5075 gnd.n6319 gnd.n394 225.874
R5076 gnd.n6327 gnd.n394 225.874
R5077 gnd.n6328 gnd.n6327 225.874
R5078 gnd.n6329 gnd.n6328 225.874
R5079 gnd.n6329 gnd.n388 225.874
R5080 gnd.n6338 gnd.n388 225.874
R5081 gnd.n6339 gnd.n6338 225.874
R5082 gnd.n6340 gnd.n6339 225.874
R5083 gnd.n6340 gnd.n383 225.874
R5084 gnd.n4860 gnd.t200 224.174
R5085 gnd.n4481 gnd.t107 224.174
R5086 gnd.n3753 gnd.n3752 199.319
R5087 gnd.n3753 gnd.n3699 199.319
R5088 gnd.n1976 gnd.n1946 199.319
R5089 gnd.n1976 gnd.n1945 199.319
R5090 gnd.n1755 gnd.n1752 186.49
R5091 gnd.n3554 gnd.n3551 186.49
R5092 gnd.n5642 gnd.n5641 185
R5093 gnd.n5640 gnd.n5639 185
R5094 gnd.n5619 gnd.n5618 185
R5095 gnd.n5634 gnd.n5633 185
R5096 gnd.n5632 gnd.n5631 185
R5097 gnd.n5623 gnd.n5622 185
R5098 gnd.n5626 gnd.n5625 185
R5099 gnd.n5610 gnd.n5609 185
R5100 gnd.n5608 gnd.n5607 185
R5101 gnd.n5587 gnd.n5586 185
R5102 gnd.n5602 gnd.n5601 185
R5103 gnd.n5600 gnd.n5599 185
R5104 gnd.n5591 gnd.n5590 185
R5105 gnd.n5594 gnd.n5593 185
R5106 gnd.n5578 gnd.n5577 185
R5107 gnd.n5576 gnd.n5575 185
R5108 gnd.n5555 gnd.n5554 185
R5109 gnd.n5570 gnd.n5569 185
R5110 gnd.n5568 gnd.n5567 185
R5111 gnd.n5559 gnd.n5558 185
R5112 gnd.n5562 gnd.n5561 185
R5113 gnd.n5547 gnd.n5546 185
R5114 gnd.n5545 gnd.n5544 185
R5115 gnd.n5524 gnd.n5523 185
R5116 gnd.n5539 gnd.n5538 185
R5117 gnd.n5537 gnd.n5536 185
R5118 gnd.n5528 gnd.n5527 185
R5119 gnd.n5531 gnd.n5530 185
R5120 gnd.n5515 gnd.n5514 185
R5121 gnd.n5513 gnd.n5512 185
R5122 gnd.n5492 gnd.n5491 185
R5123 gnd.n5507 gnd.n5506 185
R5124 gnd.n5505 gnd.n5504 185
R5125 gnd.n5496 gnd.n5495 185
R5126 gnd.n5499 gnd.n5498 185
R5127 gnd.n5483 gnd.n5482 185
R5128 gnd.n5481 gnd.n5480 185
R5129 gnd.n5460 gnd.n5459 185
R5130 gnd.n5475 gnd.n5474 185
R5131 gnd.n5473 gnd.n5472 185
R5132 gnd.n5464 gnd.n5463 185
R5133 gnd.n5467 gnd.n5466 185
R5134 gnd.n5451 gnd.n5450 185
R5135 gnd.n5449 gnd.n5448 185
R5136 gnd.n5428 gnd.n5427 185
R5137 gnd.n5443 gnd.n5442 185
R5138 gnd.n5441 gnd.n5440 185
R5139 gnd.n5432 gnd.n5431 185
R5140 gnd.n5435 gnd.n5434 185
R5141 gnd.n5420 gnd.n5419 185
R5142 gnd.n5418 gnd.n5417 185
R5143 gnd.n5397 gnd.n5396 185
R5144 gnd.n5412 gnd.n5411 185
R5145 gnd.n5410 gnd.n5409 185
R5146 gnd.n5401 gnd.n5400 185
R5147 gnd.n5404 gnd.n5403 185
R5148 gnd.n4861 gnd.t199 178.987
R5149 gnd.n4482 gnd.t108 178.987
R5150 gnd.n1 gnd.t202 170.774
R5151 gnd.n7 gnd.t238 170.103
R5152 gnd.n6 gnd.t270 170.103
R5153 gnd.n5 gnd.t231 170.103
R5154 gnd.n4 gnd.t227 170.103
R5155 gnd.n3 gnd.t8 170.103
R5156 gnd.n2 gnd.t10 170.103
R5157 gnd.n1 gnd.t35 170.103
R5158 gnd.n3622 gnd.n3621 163.367
R5159 gnd.n3618 gnd.n3617 163.367
R5160 gnd.n3614 gnd.n3613 163.367
R5161 gnd.n3610 gnd.n3609 163.367
R5162 gnd.n3606 gnd.n3605 163.367
R5163 gnd.n3602 gnd.n3601 163.367
R5164 gnd.n3598 gnd.n3597 163.367
R5165 gnd.n3594 gnd.n3593 163.367
R5166 gnd.n3590 gnd.n3589 163.367
R5167 gnd.n3586 gnd.n3585 163.367
R5168 gnd.n3582 gnd.n3581 163.367
R5169 gnd.n3578 gnd.n3577 163.367
R5170 gnd.n3574 gnd.n3573 163.367
R5171 gnd.n3570 gnd.n3569 163.367
R5172 gnd.n3565 gnd.n3564 163.367
R5173 gnd.n3697 gnd.n1364 163.367
R5174 gnd.n3694 gnd.n3693 163.367
R5175 gnd.n3691 gnd.n1397 163.367
R5176 gnd.n3686 gnd.n3685 163.367
R5177 gnd.n3682 gnd.n3681 163.367
R5178 gnd.n3678 gnd.n3677 163.367
R5179 gnd.n3674 gnd.n3673 163.367
R5180 gnd.n3670 gnd.n3669 163.367
R5181 gnd.n3666 gnd.n3665 163.367
R5182 gnd.n3662 gnd.n3661 163.367
R5183 gnd.n3658 gnd.n3657 163.367
R5184 gnd.n3654 gnd.n3653 163.367
R5185 gnd.n3650 gnd.n3649 163.367
R5186 gnd.n3646 gnd.n3645 163.367
R5187 gnd.n3642 gnd.n3641 163.367
R5188 gnd.n3638 gnd.n3637 163.367
R5189 gnd.n3634 gnd.n3633 163.367
R5190 gnd.n2762 gnd.n1742 163.367
R5191 gnd.n2799 gnd.n1742 163.367
R5192 gnd.n2799 gnd.n1732 163.367
R5193 gnd.n2795 gnd.n1732 163.367
R5194 gnd.n2795 gnd.n1727 163.367
R5195 gnd.n2792 gnd.n1727 163.367
R5196 gnd.n2792 gnd.n1719 163.367
R5197 gnd.n2787 gnd.n1719 163.367
R5198 gnd.n2787 gnd.n1713 163.367
R5199 gnd.n2784 gnd.n1713 163.367
R5200 gnd.n2784 gnd.n1706 163.367
R5201 gnd.n2779 gnd.n1706 163.367
R5202 gnd.n2779 gnd.n1698 163.367
R5203 gnd.n2776 gnd.n1698 163.367
R5204 gnd.n2776 gnd.n1691 163.367
R5205 gnd.n1691 gnd.n1682 163.367
R5206 gnd.n1683 gnd.n1682 163.367
R5207 gnd.n1683 gnd.n1676 163.367
R5208 gnd.n2770 gnd.n1676 163.367
R5209 gnd.n2770 gnd.n1668 163.367
R5210 gnd.n2766 gnd.n1668 163.367
R5211 gnd.n2766 gnd.n1658 163.367
R5212 gnd.n1658 gnd.n1649 163.367
R5213 gnd.n2931 gnd.n1649 163.367
R5214 gnd.n2931 gnd.n1647 163.367
R5215 gnd.n2936 gnd.n1647 163.367
R5216 gnd.n2936 gnd.n1642 163.367
R5217 gnd.n1642 gnd.n1632 163.367
R5218 gnd.n2959 gnd.n1632 163.367
R5219 gnd.n2959 gnd.n1630 163.367
R5220 gnd.n2980 gnd.n1630 163.367
R5221 gnd.n2980 gnd.n1625 163.367
R5222 gnd.n2976 gnd.n1625 163.367
R5223 gnd.n2976 gnd.n2972 163.367
R5224 gnd.n2972 gnd.n2971 163.367
R5225 gnd.n2971 gnd.n1607 163.367
R5226 gnd.n1608 gnd.n1607 163.367
R5227 gnd.n1608 gnd.n1600 163.367
R5228 gnd.n2965 gnd.n1600 163.367
R5229 gnd.n2965 gnd.n1593 163.367
R5230 gnd.n3046 gnd.n1593 163.367
R5231 gnd.n3046 gnd.n1590 163.367
R5232 gnd.n3068 gnd.n1590 163.367
R5233 gnd.n3068 gnd.n1584 163.367
R5234 gnd.n3064 gnd.n1584 163.367
R5235 gnd.n3064 gnd.n1577 163.367
R5236 gnd.n3059 gnd.n1577 163.367
R5237 gnd.n3059 gnd.n1571 163.367
R5238 gnd.n3056 gnd.n1571 163.367
R5239 gnd.n3056 gnd.n1563 163.367
R5240 gnd.n3050 gnd.n1563 163.367
R5241 gnd.n3050 gnd.n1555 163.367
R5242 gnd.n1555 gnd.n1546 163.367
R5243 gnd.n3136 gnd.n1546 163.367
R5244 gnd.n3136 gnd.n1544 163.367
R5245 gnd.n3174 gnd.n1544 163.367
R5246 gnd.n3174 gnd.n1537 163.367
R5247 gnd.n3170 gnd.n1537 163.367
R5248 gnd.n3170 gnd.n3166 163.367
R5249 gnd.n3166 gnd.n3165 163.367
R5250 gnd.n3165 gnd.n1521 163.367
R5251 gnd.n1522 gnd.n1521 163.367
R5252 gnd.n1522 gnd.n1514 163.367
R5253 gnd.n3158 gnd.n1514 163.367
R5254 gnd.n3158 gnd.n1507 163.367
R5255 gnd.n3153 gnd.n1507 163.367
R5256 gnd.n3153 gnd.n1502 163.367
R5257 gnd.n3150 gnd.n1502 163.367
R5258 gnd.n3150 gnd.n1494 163.367
R5259 gnd.n3145 gnd.n1494 163.367
R5260 gnd.n3145 gnd.n1488 163.367
R5261 gnd.n3142 gnd.n1488 163.367
R5262 gnd.n3142 gnd.n1477 163.367
R5263 gnd.n1477 gnd.n1468 163.367
R5264 gnd.n3282 gnd.n1468 163.367
R5265 gnd.n3282 gnd.n1466 163.367
R5266 gnd.n3288 gnd.n1466 163.367
R5267 gnd.n3288 gnd.n1409 163.367
R5268 gnd.n1409 gnd.n1401 163.367
R5269 gnd.n3629 gnd.n1401 163.367
R5270 gnd.n2754 gnd.n1769 163.367
R5271 gnd.n2534 gnd.n1769 163.367
R5272 gnd.n2538 gnd.n2537 163.367
R5273 gnd.n2542 gnd.n2541 163.367
R5274 gnd.n2546 gnd.n2545 163.367
R5275 gnd.n2550 gnd.n2549 163.367
R5276 gnd.n2554 gnd.n2553 163.367
R5277 gnd.n2558 gnd.n2557 163.367
R5278 gnd.n2562 gnd.n2561 163.367
R5279 gnd.n2566 gnd.n2565 163.367
R5280 gnd.n2570 gnd.n2569 163.367
R5281 gnd.n2574 gnd.n2573 163.367
R5282 gnd.n2578 gnd.n2577 163.367
R5283 gnd.n2582 gnd.n2581 163.367
R5284 gnd.n2586 gnd.n2585 163.367
R5285 gnd.n2590 gnd.n2589 163.367
R5286 gnd.n2594 gnd.n2593 163.367
R5287 gnd.n2528 gnd.n2527 163.367
R5288 gnd.n2523 gnd.n2522 163.367
R5289 gnd.n2519 gnd.n2518 163.367
R5290 gnd.n2515 gnd.n2514 163.367
R5291 gnd.n2511 gnd.n2510 163.367
R5292 gnd.n2507 gnd.n2506 163.367
R5293 gnd.n2503 gnd.n2502 163.367
R5294 gnd.n2499 gnd.n2498 163.367
R5295 gnd.n2495 gnd.n2494 163.367
R5296 gnd.n2491 gnd.n2490 163.367
R5297 gnd.n2487 gnd.n2486 163.367
R5298 gnd.n2483 gnd.n2482 163.367
R5299 gnd.n2479 gnd.n2478 163.367
R5300 gnd.n2475 gnd.n2474 163.367
R5301 gnd.n2471 gnd.n2470 163.367
R5302 gnd.n2760 gnd.n1747 163.367
R5303 gnd.n1747 gnd.n1731 163.367
R5304 gnd.n2817 gnd.n1731 163.367
R5305 gnd.n2817 gnd.n1729 163.367
R5306 gnd.n2821 gnd.n1729 163.367
R5307 gnd.n2821 gnd.n1717 163.367
R5308 gnd.n2835 gnd.n1717 163.367
R5309 gnd.n2835 gnd.n1715 163.367
R5310 gnd.n2839 gnd.n1715 163.367
R5311 gnd.n2839 gnd.n1704 163.367
R5312 gnd.n2851 gnd.n1704 163.367
R5313 gnd.n2851 gnd.n1701 163.367
R5314 gnd.n2856 gnd.n1701 163.367
R5315 gnd.n2856 gnd.n1702 163.367
R5316 gnd.n1702 gnd.n1680 163.367
R5317 gnd.n2882 gnd.n1680 163.367
R5318 gnd.n2882 gnd.n1678 163.367
R5319 gnd.n2886 gnd.n1678 163.367
R5320 gnd.n2886 gnd.n1665 163.367
R5321 gnd.n2903 gnd.n1665 163.367
R5322 gnd.n2903 gnd.n1660 163.367
R5323 gnd.n2908 gnd.n1660 163.367
R5324 gnd.n2908 gnd.n1663 163.367
R5325 gnd.n1663 gnd.n1646 163.367
R5326 gnd.n2941 gnd.n1646 163.367
R5327 gnd.n2941 gnd.n1643 163.367
R5328 gnd.n2946 gnd.n1643 163.367
R5329 gnd.n2946 gnd.n1644 163.367
R5330 gnd.n1644 gnd.n1629 163.367
R5331 gnd.n2984 gnd.n1629 163.367
R5332 gnd.n2984 gnd.n1626 163.367
R5333 gnd.n2991 gnd.n1626 163.367
R5334 gnd.n2991 gnd.n1627 163.367
R5335 gnd.n2987 gnd.n1627 163.367
R5336 gnd.n2987 gnd.n1605 163.367
R5337 gnd.n3027 gnd.n1605 163.367
R5338 gnd.n3027 gnd.n1602 163.367
R5339 gnd.n3034 gnd.n1602 163.367
R5340 gnd.n3034 gnd.n1603 163.367
R5341 gnd.n3030 gnd.n1603 163.367
R5342 gnd.n3030 gnd.n1588 163.367
R5343 gnd.n3074 gnd.n1588 163.367
R5344 gnd.n3074 gnd.n1586 163.367
R5345 gnd.n3078 gnd.n1586 163.367
R5346 gnd.n3078 gnd.n1575 163.367
R5347 gnd.n3092 gnd.n1575 163.367
R5348 gnd.n3092 gnd.n1573 163.367
R5349 gnd.n3096 gnd.n1573 163.367
R5350 gnd.n3096 gnd.n1561 163.367
R5351 gnd.n3118 gnd.n1561 163.367
R5352 gnd.n3118 gnd.n1557 163.367
R5353 gnd.n3123 gnd.n1557 163.367
R5354 gnd.n3123 gnd.n1559 163.367
R5355 gnd.n1559 gnd.n1541 163.367
R5356 gnd.n3178 gnd.n1541 163.367
R5357 gnd.n3178 gnd.n1538 163.367
R5358 gnd.n3185 gnd.n1538 163.367
R5359 gnd.n3185 gnd.n1539 163.367
R5360 gnd.n3181 gnd.n1539 163.367
R5361 gnd.n3181 gnd.n1518 163.367
R5362 gnd.n3209 gnd.n1518 163.367
R5363 gnd.n3209 gnd.n1516 163.367
R5364 gnd.n3213 gnd.n1516 163.367
R5365 gnd.n3213 gnd.n1506 163.367
R5366 gnd.n3227 gnd.n1506 163.367
R5367 gnd.n3227 gnd.n1504 163.367
R5368 gnd.n3231 gnd.n1504 163.367
R5369 gnd.n3231 gnd.n1492 163.367
R5370 gnd.n3252 gnd.n1492 163.367
R5371 gnd.n3252 gnd.n1490 163.367
R5372 gnd.n3256 gnd.n1490 163.367
R5373 gnd.n3256 gnd.n1474 163.367
R5374 gnd.n3275 gnd.n1474 163.367
R5375 gnd.n3275 gnd.n1470 163.367
R5376 gnd.n3280 gnd.n1470 163.367
R5377 gnd.n3280 gnd.n1472 163.367
R5378 gnd.n1472 gnd.n1407 163.367
R5379 gnd.n3539 gnd.n1407 163.367
R5380 gnd.n3539 gnd.n1404 163.367
R5381 gnd.n3627 gnd.n1404 163.367
R5382 gnd.n3560 gnd.n3559 156.462
R5383 gnd.n5582 gnd.n5550 153.042
R5384 gnd.n5646 gnd.n5645 152.079
R5385 gnd.n5614 gnd.n5613 152.079
R5386 gnd.n5582 gnd.n5581 152.079
R5387 gnd.n1760 gnd.n1759 152
R5388 gnd.n1761 gnd.n1750 152
R5389 gnd.n1763 gnd.n1762 152
R5390 gnd.n1765 gnd.n1748 152
R5391 gnd.n1767 gnd.n1766 152
R5392 gnd.n3558 gnd.n3542 152
R5393 gnd.n3550 gnd.n3543 152
R5394 gnd.n3549 gnd.n3548 152
R5395 gnd.n3547 gnd.n3544 152
R5396 gnd.n3545 gnd.t145 150.546
R5397 gnd.t217 gnd.n5624 147.661
R5398 gnd.t31 gnd.n5592 147.661
R5399 gnd.t252 gnd.n5560 147.661
R5400 gnd.t263 gnd.n5529 147.661
R5401 gnd.t289 gnd.n5497 147.661
R5402 gnd.t21 gnd.n5465 147.661
R5403 gnd.t214 gnd.n5433 147.661
R5404 gnd.t279 gnd.n5402 147.661
R5405 gnd.n3696 gnd.n1363 143.351
R5406 gnd.n2592 gnd.n1785 143.351
R5407 gnd.n2592 gnd.n1786 143.351
R5408 gnd.n1757 gnd.t177 130.484
R5409 gnd.n6349 gnd.n6348 127.204
R5410 gnd.n6350 gnd.n6349 127.204
R5411 gnd.n6350 gnd.n377 127.204
R5412 gnd.n6358 gnd.n377 127.204
R5413 gnd.n6359 gnd.n6358 127.204
R5414 gnd.n6360 gnd.n6359 127.204
R5415 gnd.n6360 gnd.n371 127.204
R5416 gnd.n6368 gnd.n371 127.204
R5417 gnd.n6369 gnd.n6368 127.204
R5418 gnd.n6370 gnd.n6369 127.204
R5419 gnd.n6370 gnd.n365 127.204
R5420 gnd.n6378 gnd.n365 127.204
R5421 gnd.n6379 gnd.n6378 127.204
R5422 gnd.n6380 gnd.n6379 127.204
R5423 gnd.n6380 gnd.n359 127.204
R5424 gnd.n6388 gnd.n359 127.204
R5425 gnd.n6389 gnd.n6388 127.204
R5426 gnd.n6390 gnd.n6389 127.204
R5427 gnd.n6390 gnd.n353 127.204
R5428 gnd.n6398 gnd.n353 127.204
R5429 gnd.n6399 gnd.n6398 127.204
R5430 gnd.n6400 gnd.n6399 127.204
R5431 gnd.n6400 gnd.n347 127.204
R5432 gnd.n6408 gnd.n347 127.204
R5433 gnd.n6409 gnd.n6408 127.204
R5434 gnd.n6410 gnd.n6409 127.204
R5435 gnd.n6410 gnd.n341 127.204
R5436 gnd.n6418 gnd.n341 127.204
R5437 gnd.n6419 gnd.n6418 127.204
R5438 gnd.n6420 gnd.n6419 127.204
R5439 gnd.n6420 gnd.n335 127.204
R5440 gnd.n6428 gnd.n335 127.204
R5441 gnd.n6429 gnd.n6428 127.204
R5442 gnd.n6430 gnd.n6429 127.204
R5443 gnd.n6430 gnd.n329 127.204
R5444 gnd.n6438 gnd.n329 127.204
R5445 gnd.n6439 gnd.n6438 127.204
R5446 gnd.n6440 gnd.n6439 127.204
R5447 gnd.n6440 gnd.n323 127.204
R5448 gnd.n6448 gnd.n323 127.204
R5449 gnd.n6449 gnd.n6448 127.204
R5450 gnd.n6450 gnd.n6449 127.204
R5451 gnd.n6450 gnd.n317 127.204
R5452 gnd.n6458 gnd.n317 127.204
R5453 gnd.n6459 gnd.n6458 127.204
R5454 gnd.n6460 gnd.n6459 127.204
R5455 gnd.n6460 gnd.n311 127.204
R5456 gnd.n6468 gnd.n311 127.204
R5457 gnd.n6469 gnd.n6468 127.204
R5458 gnd.n6470 gnd.n6469 127.204
R5459 gnd.n6470 gnd.n305 127.204
R5460 gnd.n6478 gnd.n305 127.204
R5461 gnd.n6479 gnd.n6478 127.204
R5462 gnd.n6480 gnd.n6479 127.204
R5463 gnd.n6480 gnd.n299 127.204
R5464 gnd.n6488 gnd.n299 127.204
R5465 gnd.n6489 gnd.n6488 127.204
R5466 gnd.n6490 gnd.n6489 127.204
R5467 gnd.n6490 gnd.n293 127.204
R5468 gnd.n6498 gnd.n293 127.204
R5469 gnd.n6499 gnd.n6498 127.204
R5470 gnd.n6500 gnd.n6499 127.204
R5471 gnd.n6500 gnd.n287 127.204
R5472 gnd.n6508 gnd.n287 127.204
R5473 gnd.n6509 gnd.n6508 127.204
R5474 gnd.n6510 gnd.n6509 127.204
R5475 gnd.n6510 gnd.n281 127.204
R5476 gnd.n6518 gnd.n281 127.204
R5477 gnd.n6519 gnd.n6518 127.204
R5478 gnd.n6520 gnd.n6519 127.204
R5479 gnd.n6520 gnd.n275 127.204
R5480 gnd.n6528 gnd.n275 127.204
R5481 gnd.n6529 gnd.n6528 127.204
R5482 gnd.n6530 gnd.n6529 127.204
R5483 gnd.n6530 gnd.n269 127.204
R5484 gnd.n6538 gnd.n269 127.204
R5485 gnd.n6539 gnd.n6538 127.204
R5486 gnd.n6540 gnd.n6539 127.204
R5487 gnd.n6540 gnd.n263 127.204
R5488 gnd.n6548 gnd.n263 127.204
R5489 gnd.n6549 gnd.n6548 127.204
R5490 gnd.n6551 gnd.n6549 127.204
R5491 gnd.n6551 gnd.n6550 127.204
R5492 gnd.n1766 gnd.t109 126.766
R5493 gnd.n1764 gnd.t174 126.766
R5494 gnd.n1750 gnd.t186 126.766
R5495 gnd.n1758 gnd.t151 126.766
R5496 gnd.n3546 gnd.t188 126.766
R5497 gnd.n3548 gnd.t160 126.766
R5498 gnd.n3557 gnd.t102 126.766
R5499 gnd.n3559 gnd.t167 126.766
R5500 gnd.n3756 gnd.n3698 112.192
R5501 gnd.n2596 gnd.n2595 112.192
R5502 gnd.n5641 gnd.n5640 104.615
R5503 gnd.n5640 gnd.n5618 104.615
R5504 gnd.n5633 gnd.n5618 104.615
R5505 gnd.n5633 gnd.n5632 104.615
R5506 gnd.n5632 gnd.n5622 104.615
R5507 gnd.n5625 gnd.n5622 104.615
R5508 gnd.n5609 gnd.n5608 104.615
R5509 gnd.n5608 gnd.n5586 104.615
R5510 gnd.n5601 gnd.n5586 104.615
R5511 gnd.n5601 gnd.n5600 104.615
R5512 gnd.n5600 gnd.n5590 104.615
R5513 gnd.n5593 gnd.n5590 104.615
R5514 gnd.n5577 gnd.n5576 104.615
R5515 gnd.n5576 gnd.n5554 104.615
R5516 gnd.n5569 gnd.n5554 104.615
R5517 gnd.n5569 gnd.n5568 104.615
R5518 gnd.n5568 gnd.n5558 104.615
R5519 gnd.n5561 gnd.n5558 104.615
R5520 gnd.n5546 gnd.n5545 104.615
R5521 gnd.n5545 gnd.n5523 104.615
R5522 gnd.n5538 gnd.n5523 104.615
R5523 gnd.n5538 gnd.n5537 104.615
R5524 gnd.n5537 gnd.n5527 104.615
R5525 gnd.n5530 gnd.n5527 104.615
R5526 gnd.n5514 gnd.n5513 104.615
R5527 gnd.n5513 gnd.n5491 104.615
R5528 gnd.n5506 gnd.n5491 104.615
R5529 gnd.n5506 gnd.n5505 104.615
R5530 gnd.n5505 gnd.n5495 104.615
R5531 gnd.n5498 gnd.n5495 104.615
R5532 gnd.n5482 gnd.n5481 104.615
R5533 gnd.n5481 gnd.n5459 104.615
R5534 gnd.n5474 gnd.n5459 104.615
R5535 gnd.n5474 gnd.n5473 104.615
R5536 gnd.n5473 gnd.n5463 104.615
R5537 gnd.n5466 gnd.n5463 104.615
R5538 gnd.n5450 gnd.n5449 104.615
R5539 gnd.n5449 gnd.n5427 104.615
R5540 gnd.n5442 gnd.n5427 104.615
R5541 gnd.n5442 gnd.n5441 104.615
R5542 gnd.n5441 gnd.n5431 104.615
R5543 gnd.n5434 gnd.n5431 104.615
R5544 gnd.n5419 gnd.n5418 104.615
R5545 gnd.n5418 gnd.n5396 104.615
R5546 gnd.n5411 gnd.n5396 104.615
R5547 gnd.n5411 gnd.n5410 104.615
R5548 gnd.n5410 gnd.n5400 104.615
R5549 gnd.n5403 gnd.n5400 104.615
R5550 gnd.n4786 gnd.t101 100.632
R5551 gnd.n4437 gnd.t131 100.632
R5552 gnd.n6797 gnd.n93 99.6594
R5553 gnd.n6795 gnd.n6794 99.6594
R5554 gnd.n6790 gnd.n100 99.6594
R5555 gnd.n6788 gnd.n6787 99.6594
R5556 gnd.n6783 gnd.n107 99.6594
R5557 gnd.n6781 gnd.n6780 99.6594
R5558 gnd.n6776 gnd.n114 99.6594
R5559 gnd.n6774 gnd.n6773 99.6594
R5560 gnd.n6766 gnd.n121 99.6594
R5561 gnd.n6764 gnd.n6763 99.6594
R5562 gnd.n6759 gnd.n128 99.6594
R5563 gnd.n6757 gnd.n6756 99.6594
R5564 gnd.n6752 gnd.n135 99.6594
R5565 gnd.n6750 gnd.n6749 99.6594
R5566 gnd.n6745 gnd.n142 99.6594
R5567 gnd.n6743 gnd.n6742 99.6594
R5568 gnd.n6738 gnd.n149 99.6594
R5569 gnd.n6736 gnd.n6735 99.6594
R5570 gnd.n154 gnd.n153 99.6594
R5571 gnd.n3717 gnd.n1217 99.6594
R5572 gnd.n3721 gnd.n3720 99.6594
R5573 gnd.n3728 gnd.n3727 99.6594
R5574 gnd.n3731 gnd.n3730 99.6594
R5575 gnd.n3738 gnd.n3737 99.6594
R5576 gnd.n3741 gnd.n3740 99.6594
R5577 gnd.n3749 gnd.n3748 99.6594
R5578 gnd.n3752 gnd.n3751 99.6594
R5579 gnd.n3762 gnd.n3761 99.6594
R5580 gnd.n3765 gnd.n3764 99.6594
R5581 gnd.n3772 gnd.n3771 99.6594
R5582 gnd.n3775 gnd.n3774 99.6594
R5583 gnd.n3782 gnd.n3781 99.6594
R5584 gnd.n3785 gnd.n3784 99.6594
R5585 gnd.n3792 gnd.n3791 99.6594
R5586 gnd.n3795 gnd.n3794 99.6594
R5587 gnd.n3803 gnd.n3802 99.6594
R5588 gnd.n3806 gnd.n3805 99.6594
R5589 gnd.n2624 gnd.n2623 99.6594
R5590 gnd.n2619 gnd.n1952 99.6594
R5591 gnd.n2615 gnd.n1951 99.6594
R5592 gnd.n2611 gnd.n1950 99.6594
R5593 gnd.n2607 gnd.n1949 99.6594
R5594 gnd.n2603 gnd.n1948 99.6594
R5595 gnd.n2599 gnd.n1947 99.6594
R5596 gnd.n2461 gnd.n1945 99.6594
R5597 gnd.n2459 gnd.n1944 99.6594
R5598 gnd.n2455 gnd.n1943 99.6594
R5599 gnd.n2451 gnd.n1942 99.6594
R5600 gnd.n2447 gnd.n1941 99.6594
R5601 gnd.n2443 gnd.n1940 99.6594
R5602 gnd.n2439 gnd.n1939 99.6594
R5603 gnd.n2435 gnd.n1938 99.6594
R5604 gnd.n2431 gnd.n1937 99.6594
R5605 gnd.n2427 gnd.n1936 99.6594
R5606 gnd.n1994 gnd.n1935 99.6594
R5607 gnd.n4405 gnd.n4404 99.6594
R5608 gnd.n4399 gnd.n802 99.6594
R5609 gnd.n4396 gnd.n803 99.6594
R5610 gnd.n4392 gnd.n804 99.6594
R5611 gnd.n4388 gnd.n805 99.6594
R5612 gnd.n4384 gnd.n806 99.6594
R5613 gnd.n4380 gnd.n807 99.6594
R5614 gnd.n4376 gnd.n808 99.6594
R5615 gnd.n4372 gnd.n809 99.6594
R5616 gnd.n4367 gnd.n810 99.6594
R5617 gnd.n4363 gnd.n811 99.6594
R5618 gnd.n4359 gnd.n812 99.6594
R5619 gnd.n4355 gnd.n813 99.6594
R5620 gnd.n4351 gnd.n814 99.6594
R5621 gnd.n4347 gnd.n815 99.6594
R5622 gnd.n4343 gnd.n816 99.6594
R5623 gnd.n4339 gnd.n817 99.6594
R5624 gnd.n4335 gnd.n818 99.6594
R5625 gnd.n873 gnd.n819 99.6594
R5626 gnd.n5790 gnd.n4417 99.6594
R5627 gnd.n5788 gnd.n5787 99.6594
R5628 gnd.n5783 gnd.n4424 99.6594
R5629 gnd.n5781 gnd.n5780 99.6594
R5630 gnd.n5776 gnd.n4431 99.6594
R5631 gnd.n5774 gnd.n5773 99.6594
R5632 gnd.n5769 gnd.n4440 99.6594
R5633 gnd.n5767 gnd.n5766 99.6594
R5634 gnd.n5072 gnd.n4729 99.6594
R5635 gnd.n4755 gnd.n4736 99.6594
R5636 gnd.n4757 gnd.n4737 99.6594
R5637 gnd.n4765 gnd.n4738 99.6594
R5638 gnd.n4767 gnd.n4739 99.6594
R5639 gnd.n4775 gnd.n4740 99.6594
R5640 gnd.n4777 gnd.n4741 99.6594
R5641 gnd.n4785 gnd.n4742 99.6594
R5642 gnd.n5758 gnd.n4447 99.6594
R5643 gnd.n5756 gnd.n5755 99.6594
R5644 gnd.n5751 gnd.n4454 99.6594
R5645 gnd.n5749 gnd.n5748 99.6594
R5646 gnd.n5744 gnd.n4461 99.6594
R5647 gnd.n5742 gnd.n5741 99.6594
R5648 gnd.n5737 gnd.n4468 99.6594
R5649 gnd.n5735 gnd.n5734 99.6594
R5650 gnd.n5730 gnd.n4475 99.6594
R5651 gnd.n5728 gnd.n5727 99.6594
R5652 gnd.n5723 gnd.n4484 99.6594
R5653 gnd.n5721 gnd.n5720 99.6594
R5654 gnd.n5716 gnd.n5715 99.6594
R5655 gnd.n4913 gnd.n4912 99.6594
R5656 gnd.n4907 gnd.n4824 99.6594
R5657 gnd.n4904 gnd.n4825 99.6594
R5658 gnd.n4900 gnd.n4826 99.6594
R5659 gnd.n4896 gnd.n4827 99.6594
R5660 gnd.n4892 gnd.n4828 99.6594
R5661 gnd.n4888 gnd.n4829 99.6594
R5662 gnd.n4884 gnd.n4830 99.6594
R5663 gnd.n4880 gnd.n4831 99.6594
R5664 gnd.n4876 gnd.n4832 99.6594
R5665 gnd.n4872 gnd.n4833 99.6594
R5666 gnd.n4868 gnd.n4834 99.6594
R5667 gnd.n4915 gnd.n4823 99.6594
R5668 gnd.n6646 gnd.n6645 99.6594
R5669 gnd.n6651 gnd.n6650 99.6594
R5670 gnd.n6654 gnd.n6653 99.6594
R5671 gnd.n6659 gnd.n6658 99.6594
R5672 gnd.n6662 gnd.n6661 99.6594
R5673 gnd.n6667 gnd.n6666 99.6594
R5674 gnd.n6670 gnd.n6669 99.6594
R5675 gnd.n6675 gnd.n6674 99.6594
R5676 gnd.n6678 gnd.n80 99.6594
R5677 gnd.n3372 gnd.n3371 99.6594
R5678 gnd.n3375 gnd.n3374 99.6594
R5679 gnd.n3391 gnd.n3390 99.6594
R5680 gnd.n3394 gnd.n3393 99.6594
R5681 gnd.n3410 gnd.n3409 99.6594
R5682 gnd.n3413 gnd.n3412 99.6594
R5683 gnd.n3429 gnd.n3428 99.6594
R5684 gnd.n3432 gnd.n3431 99.6594
R5685 gnd.n3450 gnd.n3449 99.6594
R5686 gnd.n1922 gnd.n1921 99.6594
R5687 gnd.n1923 gnd.n1871 99.6594
R5688 gnd.n1925 gnd.n1879 99.6594
R5689 gnd.n1927 gnd.n1926 99.6594
R5690 gnd.n1928 gnd.n1888 99.6594
R5691 gnd.n1930 gnd.n1897 99.6594
R5692 gnd.n1932 gnd.n1931 99.6594
R5693 gnd.n1933 gnd.n1906 99.6594
R5694 gnd.n2627 gnd.n2626 99.6594
R5695 gnd.n2148 gnd.n820 99.6594
R5696 gnd.n2145 gnd.n821 99.6594
R5697 gnd.n2141 gnd.n822 99.6594
R5698 gnd.n2137 gnd.n823 99.6594
R5699 gnd.n2133 gnd.n824 99.6594
R5700 gnd.n2129 gnd.n825 99.6594
R5701 gnd.n2125 gnd.n826 99.6594
R5702 gnd.n2121 gnd.n827 99.6594
R5703 gnd.n2117 gnd.n828 99.6594
R5704 gnd.n2146 gnd.n820 99.6594
R5705 gnd.n2142 gnd.n821 99.6594
R5706 gnd.n2138 gnd.n822 99.6594
R5707 gnd.n2134 gnd.n823 99.6594
R5708 gnd.n2130 gnd.n824 99.6594
R5709 gnd.n2126 gnd.n825 99.6594
R5710 gnd.n2122 gnd.n826 99.6594
R5711 gnd.n2118 gnd.n827 99.6594
R5712 gnd.n2105 gnd.n828 99.6594
R5713 gnd.n2626 gnd.n1917 99.6594
R5714 gnd.n1933 gnd.n1905 99.6594
R5715 gnd.n1932 gnd.n1898 99.6594
R5716 gnd.n1930 gnd.n1929 99.6594
R5717 gnd.n1928 gnd.n1887 99.6594
R5718 gnd.n1927 gnd.n1880 99.6594
R5719 gnd.n1925 gnd.n1924 99.6594
R5720 gnd.n1923 gnd.n1870 99.6594
R5721 gnd.n1922 gnd.n1920 99.6594
R5722 gnd.n3373 gnd.n3372 99.6594
R5723 gnd.n3374 gnd.n3356 99.6594
R5724 gnd.n3392 gnd.n3391 99.6594
R5725 gnd.n3393 gnd.n3347 99.6594
R5726 gnd.n3411 gnd.n3410 99.6594
R5727 gnd.n3412 gnd.n3338 99.6594
R5728 gnd.n3430 gnd.n3429 99.6594
R5729 gnd.n3431 gnd.n3329 99.6594
R5730 gnd.n3451 gnd.n3450 99.6594
R5731 gnd.n6679 gnd.n6678 99.6594
R5732 gnd.n6674 gnd.n6673 99.6594
R5733 gnd.n6669 gnd.n6668 99.6594
R5734 gnd.n6666 gnd.n6665 99.6594
R5735 gnd.n6661 gnd.n6660 99.6594
R5736 gnd.n6658 gnd.n6657 99.6594
R5737 gnd.n6653 gnd.n6652 99.6594
R5738 gnd.n6650 gnd.n6649 99.6594
R5739 gnd.n6645 gnd.n6644 99.6594
R5740 gnd.n4913 gnd.n4836 99.6594
R5741 gnd.n4905 gnd.n4824 99.6594
R5742 gnd.n4901 gnd.n4825 99.6594
R5743 gnd.n4897 gnd.n4826 99.6594
R5744 gnd.n4893 gnd.n4827 99.6594
R5745 gnd.n4889 gnd.n4828 99.6594
R5746 gnd.n4885 gnd.n4829 99.6594
R5747 gnd.n4881 gnd.n4830 99.6594
R5748 gnd.n4877 gnd.n4831 99.6594
R5749 gnd.n4873 gnd.n4832 99.6594
R5750 gnd.n4869 gnd.n4833 99.6594
R5751 gnd.n4865 gnd.n4834 99.6594
R5752 gnd.n4916 gnd.n4915 99.6594
R5753 gnd.n5715 gnd.n4486 99.6594
R5754 gnd.n5722 gnd.n5721 99.6594
R5755 gnd.n4484 gnd.n4476 99.6594
R5756 gnd.n5729 gnd.n5728 99.6594
R5757 gnd.n4475 gnd.n4469 99.6594
R5758 gnd.n5736 gnd.n5735 99.6594
R5759 gnd.n4468 gnd.n4462 99.6594
R5760 gnd.n5743 gnd.n5742 99.6594
R5761 gnd.n4461 gnd.n4455 99.6594
R5762 gnd.n5750 gnd.n5749 99.6594
R5763 gnd.n4454 gnd.n4448 99.6594
R5764 gnd.n5757 gnd.n5756 99.6594
R5765 gnd.n4447 gnd.n4444 99.6594
R5766 gnd.n5073 gnd.n5072 99.6594
R5767 gnd.n4758 gnd.n4736 99.6594
R5768 gnd.n4764 gnd.n4737 99.6594
R5769 gnd.n4768 gnd.n4738 99.6594
R5770 gnd.n4774 gnd.n4739 99.6594
R5771 gnd.n4778 gnd.n4740 99.6594
R5772 gnd.n4784 gnd.n4741 99.6594
R5773 gnd.n4742 gnd.n4726 99.6594
R5774 gnd.n5768 gnd.n5767 99.6594
R5775 gnd.n4440 gnd.n4432 99.6594
R5776 gnd.n5775 gnd.n5774 99.6594
R5777 gnd.n4431 gnd.n4425 99.6594
R5778 gnd.n5782 gnd.n5781 99.6594
R5779 gnd.n4424 gnd.n4418 99.6594
R5780 gnd.n5789 gnd.n5788 99.6594
R5781 gnd.n4417 gnd.n4414 99.6594
R5782 gnd.n4405 gnd.n832 99.6594
R5783 gnd.n4397 gnd.n802 99.6594
R5784 gnd.n4393 gnd.n803 99.6594
R5785 gnd.n4389 gnd.n804 99.6594
R5786 gnd.n4385 gnd.n805 99.6594
R5787 gnd.n4381 gnd.n806 99.6594
R5788 gnd.n4377 gnd.n807 99.6594
R5789 gnd.n4373 gnd.n808 99.6594
R5790 gnd.n4368 gnd.n809 99.6594
R5791 gnd.n4364 gnd.n810 99.6594
R5792 gnd.n4360 gnd.n811 99.6594
R5793 gnd.n4356 gnd.n812 99.6594
R5794 gnd.n4352 gnd.n813 99.6594
R5795 gnd.n4348 gnd.n814 99.6594
R5796 gnd.n4344 gnd.n815 99.6594
R5797 gnd.n4340 gnd.n816 99.6594
R5798 gnd.n4336 gnd.n817 99.6594
R5799 gnd.n872 gnd.n818 99.6594
R5800 gnd.n4328 gnd.n819 99.6594
R5801 gnd.n2426 gnd.n1935 99.6594
R5802 gnd.n2430 gnd.n1936 99.6594
R5803 gnd.n2434 gnd.n1937 99.6594
R5804 gnd.n2438 gnd.n1938 99.6594
R5805 gnd.n2442 gnd.n1939 99.6594
R5806 gnd.n2446 gnd.n1940 99.6594
R5807 gnd.n2450 gnd.n1941 99.6594
R5808 gnd.n2454 gnd.n1942 99.6594
R5809 gnd.n2458 gnd.n1943 99.6594
R5810 gnd.n2462 gnd.n1944 99.6594
R5811 gnd.n2598 gnd.n1946 99.6594
R5812 gnd.n2602 gnd.n1947 99.6594
R5813 gnd.n2606 gnd.n1948 99.6594
R5814 gnd.n2610 gnd.n1949 99.6594
R5815 gnd.n2614 gnd.n1950 99.6594
R5816 gnd.n2618 gnd.n1951 99.6594
R5817 gnd.n1954 gnd.n1952 99.6594
R5818 gnd.n2624 gnd.n1953 99.6594
R5819 gnd.n3718 gnd.n3717 99.6594
R5820 gnd.n3720 gnd.n3709 99.6594
R5821 gnd.n3729 gnd.n3728 99.6594
R5822 gnd.n3730 gnd.n3705 99.6594
R5823 gnd.n3739 gnd.n3738 99.6594
R5824 gnd.n3740 gnd.n3701 99.6594
R5825 gnd.n3750 gnd.n3749 99.6594
R5826 gnd.n3699 gnd.n1357 99.6594
R5827 gnd.n3763 gnd.n3762 99.6594
R5828 gnd.n3764 gnd.n1353 99.6594
R5829 gnd.n3773 gnd.n3772 99.6594
R5830 gnd.n3774 gnd.n1349 99.6594
R5831 gnd.n3783 gnd.n3782 99.6594
R5832 gnd.n3784 gnd.n1345 99.6594
R5833 gnd.n3793 gnd.n3792 99.6594
R5834 gnd.n3794 gnd.n1341 99.6594
R5835 gnd.n3804 gnd.n3803 99.6594
R5836 gnd.n3807 gnd.n3806 99.6594
R5837 gnd.n153 gnd.n150 99.6594
R5838 gnd.n6737 gnd.n6736 99.6594
R5839 gnd.n149 gnd.n143 99.6594
R5840 gnd.n6744 gnd.n6743 99.6594
R5841 gnd.n142 gnd.n136 99.6594
R5842 gnd.n6751 gnd.n6750 99.6594
R5843 gnd.n135 gnd.n129 99.6594
R5844 gnd.n6758 gnd.n6757 99.6594
R5845 gnd.n128 gnd.n122 99.6594
R5846 gnd.n6765 gnd.n6764 99.6594
R5847 gnd.n121 gnd.n115 99.6594
R5848 gnd.n6775 gnd.n6774 99.6594
R5849 gnd.n114 gnd.n108 99.6594
R5850 gnd.n6782 gnd.n6781 99.6594
R5851 gnd.n107 gnd.n101 99.6594
R5852 gnd.n6789 gnd.n6788 99.6594
R5853 gnd.n100 gnd.n94 99.6594
R5854 gnd.n6796 gnd.n6795 99.6594
R5855 gnd.n93 gnd.n90 99.6594
R5856 gnd.n2674 gnd.n2673 99.6594
R5857 gnd.n1874 gnd.n1850 99.6594
R5858 gnd.n1876 gnd.n1851 99.6594
R5859 gnd.n1884 gnd.n1852 99.6594
R5860 gnd.n1892 gnd.n1853 99.6594
R5861 gnd.n1894 gnd.n1854 99.6594
R5862 gnd.n1902 gnd.n1855 99.6594
R5863 gnd.n1912 gnd.n1856 99.6594
R5864 gnd.n1914 gnd.n1857 99.6594
R5865 gnd.n2385 gnd.n1858 99.6594
R5866 gnd.n2387 gnd.n1859 99.6594
R5867 gnd.n2391 gnd.n1860 99.6594
R5868 gnd.n2397 gnd.n1861 99.6594
R5869 gnd.n2676 gnd.n1848 99.6594
R5870 gnd.n2674 gnd.n1864 99.6594
R5871 gnd.n1875 gnd.n1850 99.6594
R5872 gnd.n1883 gnd.n1851 99.6594
R5873 gnd.n1891 gnd.n1852 99.6594
R5874 gnd.n1893 gnd.n1853 99.6594
R5875 gnd.n1901 gnd.n1854 99.6594
R5876 gnd.n1911 gnd.n1855 99.6594
R5877 gnd.n1913 gnd.n1856 99.6594
R5878 gnd.n2384 gnd.n1857 99.6594
R5879 gnd.n2386 gnd.n1858 99.6594
R5880 gnd.n2390 gnd.n1859 99.6594
R5881 gnd.n2392 gnd.n1860 99.6594
R5882 gnd.n2398 gnd.n1861 99.6594
R5883 gnd.n2677 gnd.n2676 99.6594
R5884 gnd.n3381 gnd.n3361 99.6594
R5885 gnd.n3385 gnd.n3383 99.6594
R5886 gnd.n3400 gnd.n3352 99.6594
R5887 gnd.n3404 gnd.n3402 99.6594
R5888 gnd.n3419 gnd.n3343 99.6594
R5889 gnd.n3423 gnd.n3421 99.6594
R5890 gnd.n3438 gnd.n3334 99.6594
R5891 gnd.n3441 gnd.n3440 99.6594
R5892 gnd.n3442 gnd.n3323 99.6594
R5893 gnd.n3461 gnd.n3460 99.6594
R5894 gnd.n3462 gnd.n3319 99.6594
R5895 gnd.n3471 gnd.n3470 99.6594
R5896 gnd.n3472 gnd.n3315 99.6594
R5897 gnd.n3484 gnd.n3483 99.6594
R5898 gnd.n3483 gnd.n3482 99.6594
R5899 gnd.n3473 gnd.n3472 99.6594
R5900 gnd.n3470 gnd.n3469 99.6594
R5901 gnd.n3463 gnd.n3462 99.6594
R5902 gnd.n3460 gnd.n3459 99.6594
R5903 gnd.n3443 gnd.n3442 99.6594
R5904 gnd.n3440 gnd.n3439 99.6594
R5905 gnd.n3422 gnd.n3334 99.6594
R5906 gnd.n3421 gnd.n3420 99.6594
R5907 gnd.n3403 gnd.n3343 99.6594
R5908 gnd.n3402 gnd.n3401 99.6594
R5909 gnd.n3384 gnd.n3352 99.6594
R5910 gnd.n3383 gnd.n3382 99.6594
R5911 gnd.n3361 gnd.n1191 99.6594
R5912 gnd.n2393 gnd.t166 98.63
R5913 gnd.n6676 gnd.t149 98.63
R5914 gnd.n3326 gnd.t128 98.63
R5915 gnd.n1907 gnd.t158 98.63
R5916 gnd.n3754 gnd.t125 98.63
R5917 gnd.n1337 gnd.t115 98.63
R5918 gnd.n156 gnd.t96 98.63
R5919 gnd.n6768 gnd.t121 98.63
R5920 gnd.n852 gnd.t196 98.63
R5921 gnd.n874 gnd.t182 98.63
R5922 gnd.n2106 gnd.t173 98.63
R5923 gnd.n1996 gnd.t118 98.63
R5924 gnd.n1974 gnd.t155 98.63
R5925 gnd.n3474 gnd.t135 98.63
R5926 gnd.n2467 gnd.t193 88.9408
R5927 gnd.n1398 gnd.t184 88.9408
R5928 gnd.n2531 gnd.t144 88.933
R5929 gnd.n3561 gnd.t139 88.933
R5930 gnd.n1757 gnd.n1756 81.8399
R5931 gnd.n6550 gnd.n162 76.3231
R5932 gnd.n4787 gnd.t100 74.8376
R5933 gnd.n4438 gnd.t132 74.8376
R5934 gnd.n2468 gnd.t192 72.8438
R5935 gnd.n1399 gnd.t185 72.8438
R5936 gnd.n1758 gnd.n1751 72.8411
R5937 gnd.n1764 gnd.n1749 72.8411
R5938 gnd.n3557 gnd.n3556 72.8411
R5939 gnd.n2394 gnd.t165 72.836
R5940 gnd.n2532 gnd.t143 72.836
R5941 gnd.n3562 gnd.t140 72.836
R5942 gnd.n6677 gnd.t150 72.836
R5943 gnd.n3327 gnd.t127 72.836
R5944 gnd.n1908 gnd.t159 72.836
R5945 gnd.n3755 gnd.t124 72.836
R5946 gnd.n1338 gnd.t114 72.836
R5947 gnd.n157 gnd.t97 72.836
R5948 gnd.n6769 gnd.t122 72.836
R5949 gnd.n853 gnd.t195 72.836
R5950 gnd.n875 gnd.t181 72.836
R5951 gnd.n2107 gnd.t172 72.836
R5952 gnd.n1997 gnd.t119 72.836
R5953 gnd.n1975 gnd.t156 72.836
R5954 gnd.n3475 gnd.t136 72.836
R5955 gnd.n3622 gnd.n1366 71.676
R5956 gnd.n3618 gnd.n1367 71.676
R5957 gnd.n3614 gnd.n1368 71.676
R5958 gnd.n3610 gnd.n1369 71.676
R5959 gnd.n3606 gnd.n1370 71.676
R5960 gnd.n3602 gnd.n1371 71.676
R5961 gnd.n3598 gnd.n1372 71.676
R5962 gnd.n3594 gnd.n1373 71.676
R5963 gnd.n3590 gnd.n1374 71.676
R5964 gnd.n3586 gnd.n1375 71.676
R5965 gnd.n3582 gnd.n1376 71.676
R5966 gnd.n3578 gnd.n1377 71.676
R5967 gnd.n3574 gnd.n1378 71.676
R5968 gnd.n3570 gnd.n1379 71.676
R5969 gnd.n3565 gnd.n1380 71.676
R5970 gnd.n1381 gnd.n1364 71.676
R5971 gnd.n3694 gnd.n1363 71.676
R5972 gnd.n3692 gnd.n3691 71.676
R5973 gnd.n3686 gnd.n1396 71.676
R5974 gnd.n3682 gnd.n1395 71.676
R5975 gnd.n3678 gnd.n1394 71.676
R5976 gnd.n3674 gnd.n1393 71.676
R5977 gnd.n3670 gnd.n1392 71.676
R5978 gnd.n3666 gnd.n1391 71.676
R5979 gnd.n3662 gnd.n1390 71.676
R5980 gnd.n3658 gnd.n1389 71.676
R5981 gnd.n3654 gnd.n1388 71.676
R5982 gnd.n3650 gnd.n1387 71.676
R5983 gnd.n3646 gnd.n1386 71.676
R5984 gnd.n3642 gnd.n1385 71.676
R5985 gnd.n3638 gnd.n1384 71.676
R5986 gnd.n3634 gnd.n1383 71.676
R5987 gnd.n3630 gnd.n1382 71.676
R5988 gnd.n2753 gnd.n1746 71.676
R5989 gnd.n2534 gnd.n1771 71.676
R5990 gnd.n2538 gnd.n1772 71.676
R5991 gnd.n2542 gnd.n1773 71.676
R5992 gnd.n2546 gnd.n1774 71.676
R5993 gnd.n2550 gnd.n1775 71.676
R5994 gnd.n2554 gnd.n1776 71.676
R5995 gnd.n2558 gnd.n1777 71.676
R5996 gnd.n2562 gnd.n1778 71.676
R5997 gnd.n2566 gnd.n1779 71.676
R5998 gnd.n2570 gnd.n1780 71.676
R5999 gnd.n2574 gnd.n1781 71.676
R6000 gnd.n2578 gnd.n1782 71.676
R6001 gnd.n2582 gnd.n1783 71.676
R6002 gnd.n2586 gnd.n1784 71.676
R6003 gnd.n2590 gnd.n1785 71.676
R6004 gnd.n2593 gnd.n1787 71.676
R6005 gnd.n2527 gnd.n1788 71.676
R6006 gnd.n2522 gnd.n1789 71.676
R6007 gnd.n2518 gnd.n1790 71.676
R6008 gnd.n2514 gnd.n1791 71.676
R6009 gnd.n2510 gnd.n1792 71.676
R6010 gnd.n2506 gnd.n1793 71.676
R6011 gnd.n2502 gnd.n1794 71.676
R6012 gnd.n2498 gnd.n1795 71.676
R6013 gnd.n2494 gnd.n1796 71.676
R6014 gnd.n2490 gnd.n1797 71.676
R6015 gnd.n2486 gnd.n1798 71.676
R6016 gnd.n2482 gnd.n1799 71.676
R6017 gnd.n2478 gnd.n1800 71.676
R6018 gnd.n2474 gnd.n1801 71.676
R6019 gnd.n2470 gnd.n1802 71.676
R6020 gnd.n2754 gnd.n2753 71.676
R6021 gnd.n2537 gnd.n1771 71.676
R6022 gnd.n2541 gnd.n1772 71.676
R6023 gnd.n2545 gnd.n1773 71.676
R6024 gnd.n2549 gnd.n1774 71.676
R6025 gnd.n2553 gnd.n1775 71.676
R6026 gnd.n2557 gnd.n1776 71.676
R6027 gnd.n2561 gnd.n1777 71.676
R6028 gnd.n2565 gnd.n1778 71.676
R6029 gnd.n2569 gnd.n1779 71.676
R6030 gnd.n2573 gnd.n1780 71.676
R6031 gnd.n2577 gnd.n1781 71.676
R6032 gnd.n2581 gnd.n1782 71.676
R6033 gnd.n2585 gnd.n1783 71.676
R6034 gnd.n2589 gnd.n1784 71.676
R6035 gnd.n2594 gnd.n1786 71.676
R6036 gnd.n2528 gnd.n1787 71.676
R6037 gnd.n2523 gnd.n1788 71.676
R6038 gnd.n2519 gnd.n1789 71.676
R6039 gnd.n2515 gnd.n1790 71.676
R6040 gnd.n2511 gnd.n1791 71.676
R6041 gnd.n2507 gnd.n1792 71.676
R6042 gnd.n2503 gnd.n1793 71.676
R6043 gnd.n2499 gnd.n1794 71.676
R6044 gnd.n2495 gnd.n1795 71.676
R6045 gnd.n2491 gnd.n1796 71.676
R6046 gnd.n2487 gnd.n1797 71.676
R6047 gnd.n2483 gnd.n1798 71.676
R6048 gnd.n2479 gnd.n1799 71.676
R6049 gnd.n2475 gnd.n1800 71.676
R6050 gnd.n2471 gnd.n1801 71.676
R6051 gnd.n1802 gnd.n1744 71.676
R6052 gnd.n3633 gnd.n1382 71.676
R6053 gnd.n3637 gnd.n1383 71.676
R6054 gnd.n3641 gnd.n1384 71.676
R6055 gnd.n3645 gnd.n1385 71.676
R6056 gnd.n3649 gnd.n1386 71.676
R6057 gnd.n3653 gnd.n1387 71.676
R6058 gnd.n3657 gnd.n1388 71.676
R6059 gnd.n3661 gnd.n1389 71.676
R6060 gnd.n3665 gnd.n1390 71.676
R6061 gnd.n3669 gnd.n1391 71.676
R6062 gnd.n3673 gnd.n1392 71.676
R6063 gnd.n3677 gnd.n1393 71.676
R6064 gnd.n3681 gnd.n1394 71.676
R6065 gnd.n3685 gnd.n1395 71.676
R6066 gnd.n1397 gnd.n1396 71.676
R6067 gnd.n3693 gnd.n3692 71.676
R6068 gnd.n3697 gnd.n3696 71.676
R6069 gnd.n3564 gnd.n1381 71.676
R6070 gnd.n3569 gnd.n1380 71.676
R6071 gnd.n3573 gnd.n1379 71.676
R6072 gnd.n3577 gnd.n1378 71.676
R6073 gnd.n3581 gnd.n1377 71.676
R6074 gnd.n3585 gnd.n1376 71.676
R6075 gnd.n3589 gnd.n1375 71.676
R6076 gnd.n3593 gnd.n1374 71.676
R6077 gnd.n3597 gnd.n1373 71.676
R6078 gnd.n3601 gnd.n1372 71.676
R6079 gnd.n3605 gnd.n1371 71.676
R6080 gnd.n3609 gnd.n1370 71.676
R6081 gnd.n3613 gnd.n1369 71.676
R6082 gnd.n3617 gnd.n1368 71.676
R6083 gnd.n3621 gnd.n1367 71.676
R6084 gnd.n1405 gnd.n1366 71.676
R6085 gnd.n8 gnd.t283 69.1507
R6086 gnd.n14 gnd.t229 68.4792
R6087 gnd.n13 gnd.t204 68.4792
R6088 gnd.n12 gnd.t272 68.4792
R6089 gnd.n11 gnd.t275 68.4792
R6090 gnd.n10 gnd.t285 68.4792
R6091 gnd.n9 gnd.t37 68.4792
R6092 gnd.n8 gnd.t277 68.4792
R6093 gnd.n4914 gnd.n4818 64.369
R6094 gnd.n4406 gnd.n830 63.0944
R6095 gnd.n6805 gnd.n83 63.0944
R6096 gnd.n2525 gnd.n2468 59.5399
R6097 gnd.n3688 gnd.n1399 59.5399
R6098 gnd.n2533 gnd.n2532 59.5399
R6099 gnd.n3567 gnd.n3562 59.5399
R6100 gnd.n2757 gnd.n1767 59.1804
R6101 gnd.n5798 gnd.n4407 57.3586
R6102 gnd.n5012 gnd.t243 56.607
R6103 gnd.n40 gnd.t88 56.607
R6104 gnd.n4989 gnd.t223 56.407
R6105 gnd.n5000 gnd.t286 56.407
R6106 gnd.n17 gnd.t250 56.407
R6107 gnd.n28 gnd.t249 56.407
R6108 gnd.n5021 gnd.t43 55.8337
R6109 gnd.n4998 gnd.t25 55.8337
R6110 gnd.n5009 gnd.t40 55.8337
R6111 gnd.n49 gnd.t290 55.8337
R6112 gnd.n26 gnd.t12 55.8337
R6113 gnd.n37 gnd.t259 55.8337
R6114 gnd.n1755 gnd.n1754 54.358
R6115 gnd.n3554 gnd.n3553 54.358
R6116 gnd.n5012 gnd.n5011 53.0052
R6117 gnd.n5014 gnd.n5013 53.0052
R6118 gnd.n5016 gnd.n5015 53.0052
R6119 gnd.n5018 gnd.n5017 53.0052
R6120 gnd.n5020 gnd.n5019 53.0052
R6121 gnd.n4989 gnd.n4988 53.0052
R6122 gnd.n4991 gnd.n4990 53.0052
R6123 gnd.n4993 gnd.n4992 53.0052
R6124 gnd.n4995 gnd.n4994 53.0052
R6125 gnd.n4997 gnd.n4996 53.0052
R6126 gnd.n5000 gnd.n4999 53.0052
R6127 gnd.n5002 gnd.n5001 53.0052
R6128 gnd.n5004 gnd.n5003 53.0052
R6129 gnd.n5006 gnd.n5005 53.0052
R6130 gnd.n5008 gnd.n5007 53.0052
R6131 gnd.n48 gnd.n47 53.0052
R6132 gnd.n46 gnd.n45 53.0052
R6133 gnd.n44 gnd.n43 53.0052
R6134 gnd.n42 gnd.n41 53.0052
R6135 gnd.n40 gnd.n39 53.0052
R6136 gnd.n25 gnd.n24 53.0052
R6137 gnd.n23 gnd.n22 53.0052
R6138 gnd.n21 gnd.n20 53.0052
R6139 gnd.n19 gnd.n18 53.0052
R6140 gnd.n17 gnd.n16 53.0052
R6141 gnd.n36 gnd.n35 53.0052
R6142 gnd.n34 gnd.n33 53.0052
R6143 gnd.n32 gnd.n31 53.0052
R6144 gnd.n30 gnd.n29 53.0052
R6145 gnd.n28 gnd.n27 53.0052
R6146 gnd.n3545 gnd.n3544 52.4801
R6147 gnd.n5625 gnd.t217 52.3082
R6148 gnd.n5593 gnd.t31 52.3082
R6149 gnd.n5561 gnd.t252 52.3082
R6150 gnd.n5530 gnd.t263 52.3082
R6151 gnd.n5498 gnd.t289 52.3082
R6152 gnd.n5466 gnd.t21 52.3082
R6153 gnd.n5434 gnd.t214 52.3082
R6154 gnd.n5403 gnd.t279 52.3082
R6155 gnd.n5455 gnd.n5423 51.4173
R6156 gnd.n5519 gnd.n5518 50.455
R6157 gnd.n5487 gnd.n5486 50.455
R6158 gnd.n5455 gnd.n5454 50.455
R6159 gnd.n4861 gnd.n4860 45.1884
R6160 gnd.n4482 gnd.n4481 45.1884
R6161 gnd.n3625 gnd.n3560 44.3322
R6162 gnd.n1758 gnd.n1757 44.3189
R6163 gnd.n2395 gnd.n2394 42.2793
R6164 gnd.n4862 gnd.n4861 42.2793
R6165 gnd.n4483 gnd.n4482 42.2793
R6166 gnd.n4788 gnd.n4787 42.2793
R6167 gnd.n4439 gnd.n4438 42.2793
R6168 gnd.n6681 gnd.n6677 42.2793
R6169 gnd.n3328 gnd.n3327 42.2793
R6170 gnd.n1909 gnd.n1908 42.2793
R6171 gnd.n1339 gnd.n1338 42.2793
R6172 gnd.n6733 gnd.n157 42.2793
R6173 gnd.n6770 gnd.n6769 42.2793
R6174 gnd.n4370 gnd.n853 42.2793
R6175 gnd.n876 gnd.n875 42.2793
R6176 gnd.n2108 gnd.n2107 42.2793
R6177 gnd.n2425 gnd.n1997 42.2793
R6178 gnd.n3476 gnd.n3475 42.2793
R6179 gnd.n1756 gnd.n1755 41.6274
R6180 gnd.n3555 gnd.n3554 41.6274
R6181 gnd.n1765 gnd.n1764 40.8975
R6182 gnd.n3558 gnd.n3557 40.8975
R6183 gnd.n3756 gnd.n3755 36.9518
R6184 gnd.n2596 gnd.n1975 36.9518
R6185 gnd.n5988 gnd.n5987 36.5879
R6186 gnd.n5987 gnd.n597 36.5879
R6187 gnd.n5981 gnd.n597 36.5879
R6188 gnd.n5981 gnd.n5980 36.5879
R6189 gnd.n5980 gnd.n5979 36.5879
R6190 gnd.n5979 gnd.n605 36.5879
R6191 gnd.n5973 gnd.n605 36.5879
R6192 gnd.n5973 gnd.n5972 36.5879
R6193 gnd.n5972 gnd.n5971 36.5879
R6194 gnd.n5971 gnd.n613 36.5879
R6195 gnd.n5965 gnd.n613 36.5879
R6196 gnd.n5965 gnd.n5964 36.5879
R6197 gnd.n5964 gnd.n5963 36.5879
R6198 gnd.n5963 gnd.n621 36.5879
R6199 gnd.n5957 gnd.n621 36.5879
R6200 gnd.n5957 gnd.n5956 36.5879
R6201 gnd.n5956 gnd.n5955 36.5879
R6202 gnd.n5955 gnd.n629 36.5879
R6203 gnd.n5949 gnd.n629 36.5879
R6204 gnd.n5949 gnd.n5948 36.5879
R6205 gnd.n5948 gnd.n5947 36.5879
R6206 gnd.n5947 gnd.n637 36.5879
R6207 gnd.n5941 gnd.n637 36.5879
R6208 gnd.n5941 gnd.n5940 36.5879
R6209 gnd.n5940 gnd.n5939 36.5879
R6210 gnd.n5939 gnd.n645 36.5879
R6211 gnd.n5933 gnd.n645 36.5879
R6212 gnd.n5933 gnd.n5932 36.5879
R6213 gnd.n5932 gnd.n5931 36.5879
R6214 gnd.n5931 gnd.n653 36.5879
R6215 gnd.n5925 gnd.n653 36.5879
R6216 gnd.n5925 gnd.n5924 36.5879
R6217 gnd.n5924 gnd.n5923 36.5879
R6218 gnd.n5923 gnd.n661 36.5879
R6219 gnd.n5917 gnd.n661 36.5879
R6220 gnd.n5917 gnd.n5916 36.5879
R6221 gnd.n5916 gnd.n5915 36.5879
R6222 gnd.n5915 gnd.n669 36.5879
R6223 gnd.n5909 gnd.n669 36.5879
R6224 gnd.n5909 gnd.n5908 36.5879
R6225 gnd.n5908 gnd.n5907 36.5879
R6226 gnd.n5907 gnd.n677 36.5879
R6227 gnd.n5901 gnd.n677 36.5879
R6228 gnd.n5901 gnd.n5900 36.5879
R6229 gnd.n5900 gnd.n5899 36.5879
R6230 gnd.n5899 gnd.n685 36.5879
R6231 gnd.n5893 gnd.n685 36.5879
R6232 gnd.n5893 gnd.n5892 36.5879
R6233 gnd.n5892 gnd.n5891 36.5879
R6234 gnd.n5891 gnd.n693 36.5879
R6235 gnd.n5885 gnd.n693 36.5879
R6236 gnd.n5885 gnd.n5884 36.5879
R6237 gnd.n5884 gnd.n5883 36.5879
R6238 gnd.n5883 gnd.n701 36.5879
R6239 gnd.n5877 gnd.n701 36.5879
R6240 gnd.n5877 gnd.n5876 36.5879
R6241 gnd.n5876 gnd.n5875 36.5879
R6242 gnd.n5875 gnd.n709 36.5879
R6243 gnd.n5869 gnd.n709 36.5879
R6244 gnd.n5869 gnd.n5868 36.5879
R6245 gnd.n5868 gnd.n5867 36.5879
R6246 gnd.n5867 gnd.n717 36.5879
R6247 gnd.n5861 gnd.n717 36.5879
R6248 gnd.n5861 gnd.n5860 36.5879
R6249 gnd.n5860 gnd.n5859 36.5879
R6250 gnd.n5859 gnd.n725 36.5879
R6251 gnd.n5853 gnd.n725 36.5879
R6252 gnd.n5853 gnd.n5852 36.5879
R6253 gnd.n5852 gnd.n5851 36.5879
R6254 gnd.n5851 gnd.n733 36.5879
R6255 gnd.n5845 gnd.n733 36.5879
R6256 gnd.n5845 gnd.n5844 36.5879
R6257 gnd.n5844 gnd.n5843 36.5879
R6258 gnd.n5843 gnd.n741 36.5879
R6259 gnd.n5837 gnd.n741 36.5879
R6260 gnd.n5837 gnd.n5836 36.5879
R6261 gnd.n5836 gnd.n5835 36.5879
R6262 gnd.n5835 gnd.n749 36.5879
R6263 gnd.n5829 gnd.n749 36.5879
R6264 gnd.n5829 gnd.n5828 36.5879
R6265 gnd.n5828 gnd.n5827 36.5879
R6266 gnd.n5827 gnd.n757 36.5879
R6267 gnd.n5821 gnd.n757 36.5879
R6268 gnd.n1764 gnd.n1763 35.055
R6269 gnd.n1759 gnd.n1758 35.055
R6270 gnd.n3547 gnd.n3546 35.055
R6271 gnd.n3557 gnd.n3543 35.055
R6272 gnd.n4924 gnd.n4818 31.8661
R6273 gnd.n4924 gnd.n4923 31.8661
R6274 gnd.n4932 gnd.n4807 31.8661
R6275 gnd.n4940 gnd.n4807 31.8661
R6276 gnd.n4940 gnd.n4801 31.8661
R6277 gnd.n4948 gnd.n4801 31.8661
R6278 gnd.n4948 gnd.n4794 31.8661
R6279 gnd.n5060 gnd.n4794 31.8661
R6280 gnd.n5070 gnd.n4727 31.8661
R6281 gnd.n2165 gnd.n830 31.8661
R6282 gnd.n4319 gnd.n884 31.8661
R6283 gnd.n4319 gnd.n886 31.8661
R6284 gnd.n4313 gnd.n886 31.8661
R6285 gnd.n4313 gnd.n898 31.8661
R6286 gnd.n4307 gnd.n909 31.8661
R6287 gnd.n4301 gnd.n909 31.8661
R6288 gnd.n4295 gnd.n926 31.8661
R6289 gnd.n4289 gnd.n936 31.8661
R6290 gnd.n4289 gnd.n939 31.8661
R6291 gnd.n4283 gnd.n949 31.8661
R6292 gnd.n2233 gnd.n949 31.8661
R6293 gnd.n4275 gnd.n960 31.8661
R6294 gnd.n1918 gnd.n1082 31.8661
R6295 gnd.n2342 gnd.n1934 31.8661
R6296 gnd.n2342 gnd.n1849 31.8661
R6297 gnd.n2333 gnd.n1862 31.8661
R6298 gnd.n4069 gnd.n1194 31.8661
R6299 gnd.n4063 gnd.n4062 31.8661
R6300 gnd.n4062 gnd.n4061 31.8661
R6301 gnd.n4055 gnd.n1212 31.8661
R6302 gnd.n6587 gnd.n230 31.8661
R6303 gnd.n6595 gnd.n222 31.8661
R6304 gnd.n6595 gnd.n224 31.8661
R6305 gnd.n6603 gnd.n202 31.8661
R6306 gnd.n6611 gnd.n202 31.8661
R6307 gnd.n6619 gnd.n194 31.8661
R6308 gnd.n6627 gnd.n186 31.8661
R6309 gnd.n6627 gnd.n188 31.8661
R6310 gnd.n6635 gnd.n170 31.8661
R6311 gnd.n6717 gnd.n170 31.8661
R6312 gnd.n6717 gnd.n161 31.8661
R6313 gnd.n6725 gnd.n161 31.8661
R6314 gnd.n6805 gnd.n81 31.8661
R6315 gnd.n926 gnd.t68 30.9101
R6316 gnd.n6619 gnd.t22 30.9101
R6317 gnd.n3631 gnd.n1400 29.8151
R6318 gnd.n2763 gnd.n1743 29.8151
R6319 gnd.n2394 gnd.n2393 25.7944
R6320 gnd.n4787 gnd.n4786 25.7944
R6321 gnd.n4438 gnd.n4437 25.7944
R6322 gnd.n6677 gnd.n6676 25.7944
R6323 gnd.n3327 gnd.n3326 25.7944
R6324 gnd.n1908 gnd.n1907 25.7944
R6325 gnd.n3755 gnd.n3754 25.7944
R6326 gnd.n1338 gnd.n1337 25.7944
R6327 gnd.n157 gnd.n156 25.7944
R6328 gnd.n6769 gnd.n6768 25.7944
R6329 gnd.n853 gnd.n852 25.7944
R6330 gnd.n875 gnd.n874 25.7944
R6331 gnd.n2107 gnd.n2106 25.7944
R6332 gnd.n1997 gnd.n1996 25.7944
R6333 gnd.n1975 gnd.n1974 25.7944
R6334 gnd.n3475 gnd.n3474 25.7944
R6335 gnd.n5082 gnd.n4728 24.8557
R6336 gnd.n5092 gnd.n4711 24.8557
R6337 gnd.n4714 gnd.n4702 24.8557
R6338 gnd.n5113 gnd.n4703 24.8557
R6339 gnd.n5123 gnd.n4685 24.8557
R6340 gnd.n5134 gnd.n5133 24.8557
R6341 gnd.n5153 gnd.n4671 24.8557
R6342 gnd.n5154 gnd.n4660 24.8557
R6343 gnd.n5165 gnd.n5164 24.8557
R6344 gnd.n5175 gnd.n4653 24.8557
R6345 gnd.n5184 gnd.n4645 24.8557
R6346 gnd.n5196 gnd.n5195 24.8557
R6347 gnd.n4983 gnd.n4637 24.8557
R6348 gnd.n5206 gnd.n4627 24.8557
R6349 gnd.n5215 gnd.n4620 24.8557
R6350 gnd.n4613 gnd.n4603 24.8557
R6351 gnd.n4596 gnd.n4590 24.8557
R6352 gnd.n5270 gnd.n5269 24.8557
R6353 gnd.n5280 gnd.n5279 24.8557
R6354 gnd.n4581 gnd.n4573 24.8557
R6355 gnd.n5291 gnd.n4558 24.8557
R6356 gnd.n5310 gnd.n5309 24.8557
R6357 gnd.n5320 gnd.n4551 24.8557
R6358 gnd.n5333 gnd.n4540 24.8557
R6359 gnd.n5324 gnd.n5323 24.8557
R6360 gnd.n5356 gnd.n5355 24.8557
R6361 gnd.n5366 gnd.n4527 24.8557
R6362 gnd.n5378 gnd.n4519 24.8557
R6363 gnd.n5677 gnd.n5676 24.8557
R6364 gnd.n5692 gnd.n5691 24.8557
R6365 gnd.n5813 gnd.n776 24.8557
R6366 gnd.n5812 gnd.n779 24.8557
R6367 gnd.n5661 gnd.n788 24.8557
R6368 gnd.n5799 gnd.n799 24.8557
R6369 gnd.n5103 gnd.t278 23.2624
R6370 gnd.n4730 gnd.t99 22.6251
R6371 gnd.n4295 gnd.t38 21.9878
R6372 gnd.t73 gnd.n194 21.9878
R6373 gnd.n5821 gnd.n5820 21.9529
R6374 gnd.t262 gnd.n4735 21.3504
R6375 gnd.t206 gnd.n957 21.0318
R6376 gnd.n2244 gnd.n973 21.0318
R6377 gnd.n4262 gnd.n978 21.0318
R6378 gnd.n2253 gnd.n2066 21.0318
R6379 gnd.n4256 gnd.n987 21.0318
R6380 gnd.n4249 gnd.n995 21.0318
R6381 gnd.n2300 gnd.n998 21.0318
R6382 gnd.n2269 gnd.n1008 21.0318
R6383 gnd.n4237 gnd.n1016 21.0318
R6384 gnd.n2274 gnd.n2273 21.0318
R6385 gnd.n4231 gnd.n1026 21.0318
R6386 gnd.n4225 gnd.n1037 21.0318
R6387 gnd.n2361 gnd.n1040 21.0318
R6388 gnd.n2369 gnd.n1050 21.0318
R6389 gnd.n4213 gnd.n1058 21.0318
R6390 gnd.n2378 gnd.n1061 21.0318
R6391 gnd.n4207 gnd.n1069 21.0318
R6392 gnd.n4201 gnd.n1079 21.0318
R6393 gnd.n4054 gnd.n1215 21.0318
R6394 gnd.n4048 gnd.n1227 21.0318
R6395 gnd.n3823 gnd.n1325 21.0318
R6396 gnd.n3934 gnd.n3933 21.0318
R6397 gnd.n3916 gnd.n1318 21.0318
R6398 gnd.n3954 gnd.n1310 21.0318
R6399 gnd.n3953 gnd.n1299 21.0318
R6400 gnd.n1302 gnd.n1289 21.0318
R6401 gnd.n3976 gnd.n1291 21.0318
R6402 gnd.n3986 gnd.n1281 21.0318
R6403 gnd.n3985 gnd.n1270 21.0318
R6404 gnd.n1274 gnd.n1260 21.0318
R6405 gnd.n4010 gnd.n1262 21.0318
R6406 gnd.n4019 gnd.n248 21.0318
R6407 gnd.n6568 gnd.n6567 21.0318
R6408 gnd.n6573 gnd.n246 21.0318
R6409 gnd.n3890 gnd.n236 21.0318
R6410 gnd.n232 gnd.t18 21.0318
R6411 gnd.t14 gnd.n4504 20.7131
R6412 gnd.n4283 gnd.t56 20.7131
R6413 gnd.t81 gnd.n990 20.7131
R6414 gnd.t70 gnd.n1251 20.7131
R6415 gnd.n224 gnd.t83 20.7131
R6416 gnd.n2625 gnd.n1918 20.3945
R6417 gnd.n1212 gnd.n1204 20.3945
R6418 gnd.t54 gnd.n4550 20.0758
R6419 gnd.n4307 gnd.t24 20.0758
R6420 gnd.t2 gnd.n1029 20.0758
R6421 gnd.t44 gnd.n3964 20.0758
R6422 gnd.n188 gnd.t11 20.0758
R6423 gnd.n1752 gnd.t153 19.8005
R6424 gnd.n1752 gnd.t179 19.8005
R6425 gnd.n1753 gnd.t176 19.8005
R6426 gnd.n1753 gnd.t187 19.8005
R6427 gnd.n3551 gnd.t104 19.8005
R6428 gnd.n3551 gnd.t169 19.8005
R6429 gnd.n3552 gnd.t190 19.8005
R6430 gnd.n3552 gnd.t162 19.8005
R6431 gnd.n1749 gnd.n1748 19.5087
R6432 gnd.n1762 gnd.n1749 19.5087
R6433 gnd.n1760 gnd.n1751 19.5087
R6434 gnd.n3556 gnd.n3550 19.5087
R6435 gnd.n5246 gnd.t75 19.4385
R6436 gnd.n2682 gnd.n1845 19.3944
R6437 gnd.n2682 gnd.n1834 19.3944
R6438 gnd.n2698 gnd.n1834 19.3944
R6439 gnd.n2698 gnd.n1832 19.3944
R6440 gnd.n2702 gnd.n1832 19.3944
R6441 gnd.n2702 gnd.n1821 19.3944
R6442 gnd.n2718 gnd.n1821 19.3944
R6443 gnd.n2718 gnd.n1819 19.3944
R6444 gnd.n2722 gnd.n1819 19.3944
R6445 gnd.n2722 gnd.n1808 19.3944
R6446 gnd.n2741 gnd.n1808 19.3944
R6447 gnd.n2741 gnd.n1805 19.3944
R6448 gnd.n2748 gnd.n1805 19.3944
R6449 gnd.n2748 gnd.n1806 19.3944
R6450 gnd.n2744 gnd.n1806 19.3944
R6451 gnd.n2744 gnd.n1725 19.3944
R6452 gnd.n2825 gnd.n1725 19.3944
R6453 gnd.n2825 gnd.n1722 19.3944
R6454 gnd.n2830 gnd.n1722 19.3944
R6455 gnd.n2830 gnd.n1723 19.3944
R6456 gnd.n1723 gnd.n1695 19.3944
R6457 gnd.n2861 gnd.n1695 19.3944
R6458 gnd.n2861 gnd.n1693 19.3944
R6459 gnd.n2865 gnd.n1693 19.3944
R6460 gnd.n2865 gnd.n1674 19.3944
R6461 gnd.n2890 gnd.n1674 19.3944
R6462 gnd.n2890 gnd.n1671 19.3944
R6463 gnd.n2898 gnd.n1671 19.3944
R6464 gnd.n2898 gnd.n1672 19.3944
R6465 gnd.n2894 gnd.n1672 19.3944
R6466 gnd.n2894 gnd.n1639 19.3944
R6467 gnd.n2950 gnd.n1639 19.3944
R6468 gnd.n2950 gnd.n1636 19.3944
R6469 gnd.n2955 gnd.n1636 19.3944
R6470 gnd.n2955 gnd.n1637 19.3944
R6471 gnd.n1637 gnd.n1614 19.3944
R6472 gnd.n3004 gnd.n1614 19.3944
R6473 gnd.n3004 gnd.n1611 19.3944
R6474 gnd.n3020 gnd.n1611 19.3944
R6475 gnd.n3020 gnd.n1612 19.3944
R6476 gnd.n3016 gnd.n1612 19.3944
R6477 gnd.n3016 gnd.n3015 19.3944
R6478 gnd.n3015 gnd.n3014 19.3944
R6479 gnd.n3014 gnd.n3011 19.3944
R6480 gnd.n3011 gnd.n1568 19.3944
R6481 gnd.n3100 gnd.n1568 19.3944
R6482 gnd.n3100 gnd.n1565 19.3944
R6483 gnd.n3114 gnd.n1565 19.3944
R6484 gnd.n3114 gnd.n1566 19.3944
R6485 gnd.n3110 gnd.n1566 19.3944
R6486 gnd.n3110 gnd.n3109 19.3944
R6487 gnd.n3109 gnd.n3108 19.3944
R6488 gnd.n3108 gnd.n1528 19.3944
R6489 gnd.n3198 gnd.n1528 19.3944
R6490 gnd.n3198 gnd.n1525 19.3944
R6491 gnd.n3203 gnd.n1525 19.3944
R6492 gnd.n3203 gnd.n1526 19.3944
R6493 gnd.n1526 gnd.n1499 19.3944
R6494 gnd.n3236 gnd.n1499 19.3944
R6495 gnd.n3236 gnd.n1496 19.3944
R6496 gnd.n3248 gnd.n1496 19.3944
R6497 gnd.n3248 gnd.n1497 19.3944
R6498 gnd.n3244 gnd.n1497 19.3944
R6499 gnd.n3244 gnd.n3243 19.3944
R6500 gnd.n3243 gnd.n1463 19.3944
R6501 gnd.n3291 gnd.n1463 19.3944
R6502 gnd.n3292 gnd.n3291 19.3944
R6503 gnd.n3292 gnd.n1459 19.3944
R6504 gnd.n3296 gnd.n1459 19.3944
R6505 gnd.n3297 gnd.n3296 19.3944
R6506 gnd.n3298 gnd.n3297 19.3944
R6507 gnd.n3298 gnd.n1455 19.3944
R6508 gnd.n3302 gnd.n1455 19.3944
R6509 gnd.n3303 gnd.n3302 19.3944
R6510 gnd.n3304 gnd.n3303 19.3944
R6511 gnd.n3304 gnd.n1449 19.3944
R6512 gnd.n3308 gnd.n1449 19.3944
R6513 gnd.n3309 gnd.n3308 19.3944
R6514 gnd.n3310 gnd.n3309 19.3944
R6515 gnd.n3310 gnd.n1446 19.3944
R6516 gnd.n3490 gnd.n1446 19.3944
R6517 gnd.n3490 gnd.n1447 19.3944
R6518 gnd.n2400 gnd.n2399 19.3944
R6519 gnd.n2399 gnd.n1847 19.3944
R6520 gnd.n2678 gnd.n1847 19.3944
R6521 gnd.n2672 gnd.n2671 19.3944
R6522 gnd.n2671 gnd.n1866 19.3944
R6523 gnd.n2664 gnd.n1866 19.3944
R6524 gnd.n2664 gnd.n2663 19.3944
R6525 gnd.n2663 gnd.n1877 19.3944
R6526 gnd.n2656 gnd.n1877 19.3944
R6527 gnd.n2656 gnd.n2655 19.3944
R6528 gnd.n2655 gnd.n1885 19.3944
R6529 gnd.n2648 gnd.n1885 19.3944
R6530 gnd.n2648 gnd.n2647 19.3944
R6531 gnd.n2647 gnd.n1895 19.3944
R6532 gnd.n2640 gnd.n1895 19.3944
R6533 gnd.n2640 gnd.n2639 19.3944
R6534 gnd.n2639 gnd.n1903 19.3944
R6535 gnd.n2632 gnd.n1903 19.3944
R6536 gnd.n2632 gnd.n2631 19.3944
R6537 gnd.n2631 gnd.n1915 19.3944
R6538 gnd.n2411 gnd.n1915 19.3944
R6539 gnd.n2411 gnd.n2410 19.3944
R6540 gnd.n2410 gnd.n2409 19.3944
R6541 gnd.n2409 gnd.n2388 19.3944
R6542 gnd.n2405 gnd.n2388 19.3944
R6543 gnd.n2405 gnd.n2404 19.3944
R6544 gnd.n2404 gnd.n2403 19.3944
R6545 gnd.n4911 gnd.n4910 19.3944
R6546 gnd.n4910 gnd.n4909 19.3944
R6547 gnd.n4909 gnd.n4908 19.3944
R6548 gnd.n4908 gnd.n4906 19.3944
R6549 gnd.n4906 gnd.n4903 19.3944
R6550 gnd.n4903 gnd.n4902 19.3944
R6551 gnd.n4902 gnd.n4899 19.3944
R6552 gnd.n4899 gnd.n4898 19.3944
R6553 gnd.n4898 gnd.n4895 19.3944
R6554 gnd.n4895 gnd.n4894 19.3944
R6555 gnd.n4894 gnd.n4891 19.3944
R6556 gnd.n4891 gnd.n4890 19.3944
R6557 gnd.n4890 gnd.n4887 19.3944
R6558 gnd.n4887 gnd.n4886 19.3944
R6559 gnd.n4886 gnd.n4883 19.3944
R6560 gnd.n4883 gnd.n4882 19.3944
R6561 gnd.n4882 gnd.n4879 19.3944
R6562 gnd.n4879 gnd.n4878 19.3944
R6563 gnd.n4878 gnd.n4875 19.3944
R6564 gnd.n4875 gnd.n4874 19.3944
R6565 gnd.n4874 gnd.n4871 19.3944
R6566 gnd.n4871 gnd.n4870 19.3944
R6567 gnd.n4867 gnd.n4866 19.3944
R6568 gnd.n4866 gnd.n4822 19.3944
R6569 gnd.n4917 gnd.n4822 19.3944
R6570 gnd.n5719 gnd.n4485 19.3944
R6571 gnd.n5719 gnd.n5718 19.3944
R6572 gnd.n5718 gnd.n5717 19.3944
R6573 gnd.n5761 gnd.n5760 19.3944
R6574 gnd.n5760 gnd.n5759 19.3944
R6575 gnd.n5759 gnd.n4446 19.3944
R6576 gnd.n5754 gnd.n4446 19.3944
R6577 gnd.n5754 gnd.n5753 19.3944
R6578 gnd.n5753 gnd.n5752 19.3944
R6579 gnd.n5752 gnd.n4453 19.3944
R6580 gnd.n5747 gnd.n4453 19.3944
R6581 gnd.n5747 gnd.n5746 19.3944
R6582 gnd.n5746 gnd.n5745 19.3944
R6583 gnd.n5745 gnd.n4460 19.3944
R6584 gnd.n5740 gnd.n4460 19.3944
R6585 gnd.n5740 gnd.n5739 19.3944
R6586 gnd.n5739 gnd.n5738 19.3944
R6587 gnd.n5738 gnd.n4467 19.3944
R6588 gnd.n5733 gnd.n4467 19.3944
R6589 gnd.n5733 gnd.n5732 19.3944
R6590 gnd.n5732 gnd.n5731 19.3944
R6591 gnd.n5731 gnd.n4474 19.3944
R6592 gnd.n5726 gnd.n4474 19.3944
R6593 gnd.n5726 gnd.n5725 19.3944
R6594 gnd.n5725 gnd.n5724 19.3944
R6595 gnd.n5084 gnd.n4719 19.3944
R6596 gnd.n5094 gnd.n4719 19.3944
R6597 gnd.n5095 gnd.n5094 19.3944
R6598 gnd.n5095 gnd.n4700 19.3944
R6599 gnd.n5115 gnd.n4700 19.3944
R6600 gnd.n5115 gnd.n4693 19.3944
R6601 gnd.n5125 gnd.n4693 19.3944
R6602 gnd.n5126 gnd.n5125 19.3944
R6603 gnd.n5126 gnd.n4676 19.3944
R6604 gnd.n5146 gnd.n4676 19.3944
R6605 gnd.n5146 gnd.n4668 19.3944
R6606 gnd.n5156 gnd.n4668 19.3944
R6607 gnd.n5157 gnd.n5156 19.3944
R6608 gnd.n5157 gnd.n4650 19.3944
R6609 gnd.n5177 gnd.n4650 19.3944
R6610 gnd.n5177 gnd.n4642 19.3944
R6611 gnd.n5187 gnd.n4642 19.3944
R6612 gnd.n5188 gnd.n5187 19.3944
R6613 gnd.n5188 gnd.n4625 19.3944
R6614 gnd.n5208 gnd.n4625 19.3944
R6615 gnd.n5208 gnd.n4617 19.3944
R6616 gnd.n5218 gnd.n4617 19.3944
R6617 gnd.n5219 gnd.n5218 19.3944
R6618 gnd.n5219 gnd.n4601 19.3944
R6619 gnd.n5238 gnd.n4601 19.3944
R6620 gnd.n5238 gnd.n4586 19.3944
R6621 gnd.n5272 gnd.n4586 19.3944
R6622 gnd.n5273 gnd.n5272 19.3944
R6623 gnd.n5274 gnd.n5273 19.3944
R6624 gnd.n5274 gnd.n4572 19.3944
R6625 gnd.n4572 gnd.n4566 19.3944
R6626 gnd.n5299 gnd.n4566 19.3944
R6627 gnd.n5300 gnd.n5299 19.3944
R6628 gnd.n5300 gnd.n4549 19.3944
R6629 gnd.n4549 gnd.n4547 19.3944
R6630 gnd.n5326 gnd.n4547 19.3944
R6631 gnd.n5327 gnd.n5326 19.3944
R6632 gnd.n5327 gnd.n4522 19.3944
R6633 gnd.n5373 gnd.n4522 19.3944
R6634 gnd.n5374 gnd.n5373 19.3944
R6635 gnd.n5374 gnd.n4515 19.3944
R6636 gnd.n5385 gnd.n4515 19.3944
R6637 gnd.n5387 gnd.n5385 19.3944
R6638 gnd.n5670 gnd.n5387 19.3944
R6639 gnd.n5670 gnd.n5669 19.3944
R6640 gnd.n5669 gnd.n5390 19.3944
R6641 gnd.n5665 gnd.n5390 19.3944
R6642 gnd.n5665 gnd.n5664 19.3944
R6643 gnd.n5664 gnd.n5663 19.3944
R6644 gnd.n5663 gnd.n5660 19.3944
R6645 gnd.n5660 gnd.n5659 19.3944
R6646 gnd.n5659 gnd.n5656 19.3944
R6647 gnd.n5656 gnd.n5655 19.3944
R6648 gnd.n5075 gnd.n5074 19.3944
R6649 gnd.n5074 gnd.n4733 19.3944
R6650 gnd.n4756 gnd.n4733 19.3944
R6651 gnd.n4759 gnd.n4756 19.3944
R6652 gnd.n4759 gnd.n4752 19.3944
R6653 gnd.n4763 gnd.n4752 19.3944
R6654 gnd.n4766 gnd.n4763 19.3944
R6655 gnd.n4769 gnd.n4766 19.3944
R6656 gnd.n4769 gnd.n4750 19.3944
R6657 gnd.n4773 gnd.n4750 19.3944
R6658 gnd.n4776 gnd.n4773 19.3944
R6659 gnd.n4779 gnd.n4776 19.3944
R6660 gnd.n4779 gnd.n4748 19.3944
R6661 gnd.n4783 gnd.n4748 19.3944
R6662 gnd.n5080 gnd.n5079 19.3944
R6663 gnd.n5079 gnd.n4709 19.3944
R6664 gnd.n5105 gnd.n4709 19.3944
R6665 gnd.n5105 gnd.n4707 19.3944
R6666 gnd.n5111 gnd.n4707 19.3944
R6667 gnd.n5111 gnd.n5110 19.3944
R6668 gnd.n5110 gnd.n4683 19.3944
R6669 gnd.n5136 gnd.n4683 19.3944
R6670 gnd.n5136 gnd.n4681 19.3944
R6671 gnd.n5142 gnd.n4681 19.3944
R6672 gnd.n5142 gnd.n5141 19.3944
R6673 gnd.n5141 gnd.n4658 19.3944
R6674 gnd.n5167 gnd.n4658 19.3944
R6675 gnd.n5167 gnd.n4656 19.3944
R6676 gnd.n5173 gnd.n4656 19.3944
R6677 gnd.n5173 gnd.n5172 19.3944
R6678 gnd.n5172 gnd.n4632 19.3944
R6679 gnd.n5198 gnd.n4632 19.3944
R6680 gnd.n5198 gnd.n4630 19.3944
R6681 gnd.n5204 gnd.n4630 19.3944
R6682 gnd.n5204 gnd.n5203 19.3944
R6683 gnd.n5203 gnd.n4608 19.3944
R6684 gnd.n5228 gnd.n4608 19.3944
R6685 gnd.n5228 gnd.n4606 19.3944
R6686 gnd.n5234 gnd.n4606 19.3944
R6687 gnd.n5234 gnd.n5233 19.3944
R6688 gnd.n5233 gnd.n4577 19.3944
R6689 gnd.n5282 gnd.n4577 19.3944
R6690 gnd.n5282 gnd.n4575 19.3944
R6691 gnd.n5286 gnd.n4575 19.3944
R6692 gnd.n5286 gnd.n4556 19.3944
R6693 gnd.n5312 gnd.n4556 19.3944
R6694 gnd.n5312 gnd.n4554 19.3944
R6695 gnd.n5318 gnd.n4554 19.3944
R6696 gnd.n5318 gnd.n5317 19.3944
R6697 gnd.n5317 gnd.n4532 19.3944
R6698 gnd.n5358 gnd.n4532 19.3944
R6699 gnd.n5358 gnd.n4530 19.3944
R6700 gnd.n5364 gnd.n4530 19.3944
R6701 gnd.n5364 gnd.n5363 19.3944
R6702 gnd.n5363 gnd.n4502 19.3944
R6703 gnd.n5679 gnd.n4502 19.3944
R6704 gnd.n5679 gnd.n4500 19.3944
R6705 gnd.n5689 gnd.n4500 19.3944
R6706 gnd.n5689 gnd.n5688 19.3944
R6707 gnd.n5688 gnd.n5687 19.3944
R6708 gnd.n5687 gnd.n782 19.3944
R6709 gnd.n5810 gnd.n782 19.3944
R6710 gnd.n5810 gnd.n5809 19.3944
R6711 gnd.n5809 gnd.n5808 19.3944
R6712 gnd.n5808 gnd.n786 19.3944
R6713 gnd.n4410 gnd.n786 19.3944
R6714 gnd.n5796 gnd.n4410 19.3944
R6715 gnd.n5793 gnd.n5792 19.3944
R6716 gnd.n5792 gnd.n5791 19.3944
R6717 gnd.n5791 gnd.n4416 19.3944
R6718 gnd.n5786 gnd.n4416 19.3944
R6719 gnd.n5786 gnd.n5785 19.3944
R6720 gnd.n5785 gnd.n5784 19.3944
R6721 gnd.n5784 gnd.n4423 19.3944
R6722 gnd.n5779 gnd.n4423 19.3944
R6723 gnd.n5779 gnd.n5778 19.3944
R6724 gnd.n5778 gnd.n5777 19.3944
R6725 gnd.n5777 gnd.n4430 19.3944
R6726 gnd.n5772 gnd.n4430 19.3944
R6727 gnd.n5772 gnd.n5771 19.3944
R6728 gnd.n5771 gnd.n5770 19.3944
R6729 gnd.n4921 gnd.n4820 19.3944
R6730 gnd.n4921 gnd.n4811 19.3944
R6731 gnd.n4934 gnd.n4811 19.3944
R6732 gnd.n4934 gnd.n4809 19.3944
R6733 gnd.n4938 gnd.n4809 19.3944
R6734 gnd.n4938 gnd.n4799 19.3944
R6735 gnd.n4950 gnd.n4799 19.3944
R6736 gnd.n4950 gnd.n4797 19.3944
R6737 gnd.n5058 gnd.n4797 19.3944
R6738 gnd.n5058 gnd.n5057 19.3944
R6739 gnd.n5057 gnd.n5056 19.3944
R6740 gnd.n5056 gnd.n5055 19.3944
R6741 gnd.n5055 gnd.n5052 19.3944
R6742 gnd.n5052 gnd.n5051 19.3944
R6743 gnd.n5051 gnd.n5050 19.3944
R6744 gnd.n5050 gnd.n5048 19.3944
R6745 gnd.n5048 gnd.n5047 19.3944
R6746 gnd.n5047 gnd.n5044 19.3944
R6747 gnd.n5044 gnd.n5043 19.3944
R6748 gnd.n5043 gnd.n5042 19.3944
R6749 gnd.n5042 gnd.n5040 19.3944
R6750 gnd.n5040 gnd.n5039 19.3944
R6751 gnd.n5039 gnd.n5035 19.3944
R6752 gnd.n5035 gnd.n5034 19.3944
R6753 gnd.n5034 gnd.n5033 19.3944
R6754 gnd.n5033 gnd.n5031 19.3944
R6755 gnd.n5031 gnd.n5030 19.3944
R6756 gnd.n5030 gnd.n5027 19.3944
R6757 gnd.n5027 gnd.n5026 19.3944
R6758 gnd.n4986 gnd.n4974 19.3944
R6759 gnd.n4985 gnd.n4981 19.3944
R6760 gnd.n4979 gnd.n4978 19.3944
R6761 gnd.n4975 gnd.n4594 19.3944
R6762 gnd.n5248 gnd.n4594 19.3944
R6763 gnd.n5248 gnd.n4592 19.3944
R6764 gnd.n5267 gnd.n4592 19.3944
R6765 gnd.n5267 gnd.n5266 19.3944
R6766 gnd.n5266 gnd.n5265 19.3944
R6767 gnd.n5265 gnd.n5263 19.3944
R6768 gnd.n5263 gnd.n5262 19.3944
R6769 gnd.n5262 gnd.n5260 19.3944
R6770 gnd.n5260 gnd.n5259 19.3944
R6771 gnd.n5259 gnd.n4538 19.3944
R6772 gnd.n5335 gnd.n4538 19.3944
R6773 gnd.n5335 gnd.n4536 19.3944
R6774 gnd.n5351 gnd.n4536 19.3944
R6775 gnd.n5351 gnd.n5350 19.3944
R6776 gnd.n5350 gnd.n5349 19.3944
R6777 gnd.n5349 gnd.n5347 19.3944
R6778 gnd.n5347 gnd.n5346 19.3944
R6779 gnd.n5346 gnd.n5344 19.3944
R6780 gnd.n5344 gnd.n4495 19.3944
R6781 gnd.n5694 gnd.n4495 19.3944
R6782 gnd.n5694 gnd.n4493 19.3944
R6783 gnd.n5700 gnd.n4493 19.3944
R6784 gnd.n5701 gnd.n5700 19.3944
R6785 gnd.n5704 gnd.n5701 19.3944
R6786 gnd.n5704 gnd.n4491 19.3944
R6787 gnd.n5708 gnd.n4491 19.3944
R6788 gnd.n5711 gnd.n5708 19.3944
R6789 gnd.n5712 gnd.n5711 19.3944
R6790 gnd.n4926 gnd.n4816 19.3944
R6791 gnd.n4926 gnd.n4814 19.3944
R6792 gnd.n4930 gnd.n4814 19.3944
R6793 gnd.n4930 gnd.n4805 19.3944
R6794 gnd.n4942 gnd.n4805 19.3944
R6795 gnd.n4942 gnd.n4803 19.3944
R6796 gnd.n4946 gnd.n4803 19.3944
R6797 gnd.n4946 gnd.n4792 19.3944
R6798 gnd.n5062 gnd.n4792 19.3944
R6799 gnd.n5062 gnd.n4746 19.3944
R6800 gnd.n5068 gnd.n4746 19.3944
R6801 gnd.n5068 gnd.n5067 19.3944
R6802 gnd.n5067 gnd.n4724 19.3944
R6803 gnd.n5089 gnd.n4724 19.3944
R6804 gnd.n5089 gnd.n4717 19.3944
R6805 gnd.n5100 gnd.n4717 19.3944
R6806 gnd.n5100 gnd.n5099 19.3944
R6807 gnd.n5099 gnd.n4698 19.3944
R6808 gnd.n5120 gnd.n4698 19.3944
R6809 gnd.n5120 gnd.n4691 19.3944
R6810 gnd.n5131 gnd.n4691 19.3944
R6811 gnd.n5131 gnd.n5130 19.3944
R6812 gnd.n5130 gnd.n4674 19.3944
R6813 gnd.n5151 gnd.n4674 19.3944
R6814 gnd.n5151 gnd.n4666 19.3944
R6815 gnd.n5162 gnd.n4666 19.3944
R6816 gnd.n5162 gnd.n5161 19.3944
R6817 gnd.n5161 gnd.n4648 19.3944
R6818 gnd.n5182 gnd.n4648 19.3944
R6819 gnd.n5182 gnd.n4640 19.3944
R6820 gnd.n5193 gnd.n4640 19.3944
R6821 gnd.n5193 gnd.n5192 19.3944
R6822 gnd.n5192 gnd.n4623 19.3944
R6823 gnd.n5213 gnd.n4623 19.3944
R6824 gnd.n5213 gnd.n4615 19.3944
R6825 gnd.n5223 gnd.n4615 19.3944
R6826 gnd.n5223 gnd.n4599 19.3944
R6827 gnd.n5244 gnd.n4599 19.3944
R6828 gnd.n5244 gnd.n5243 19.3944
R6829 gnd.n5243 gnd.n4583 19.3944
R6830 gnd.n5277 gnd.n4583 19.3944
R6831 gnd.n5277 gnd.n4568 19.3944
R6832 gnd.n5294 gnd.n4568 19.3944
R6833 gnd.n5294 gnd.n4564 19.3944
R6834 gnd.n5307 gnd.n4564 19.3944
R6835 gnd.n5307 gnd.n5306 19.3944
R6836 gnd.n5306 gnd.n4543 19.3944
R6837 gnd.n5331 gnd.n4543 19.3944
R6838 gnd.n5331 gnd.n5330 19.3944
R6839 gnd.n5330 gnd.n4524 19.3944
R6840 gnd.n5369 gnd.n4524 19.3944
R6841 gnd.n5369 gnd.n4517 19.3944
R6842 gnd.n5380 gnd.n4517 19.3944
R6843 gnd.n5380 gnd.n4511 19.3944
R6844 gnd.n5674 gnd.n4511 19.3944
R6845 gnd.n5674 gnd.n5673 19.3944
R6846 gnd.n5673 gnd.n770 19.3944
R6847 gnd.n5817 gnd.n770 19.3944
R6848 gnd.n5817 gnd.n5816 19.3944
R6849 gnd.n5816 gnd.n5815 19.3944
R6850 gnd.n5815 gnd.n774 19.3944
R6851 gnd.n794 gnd.n774 19.3944
R6852 gnd.n5803 gnd.n794 19.3944
R6853 gnd.n5803 gnd.n5802 19.3944
R6854 gnd.n5802 gnd.n5801 19.3944
R6855 gnd.n3816 gnd.n1334 19.3944
R6856 gnd.n3816 gnd.n1331 19.3944
R6857 gnd.n3821 gnd.n1331 19.3944
R6858 gnd.n3821 gnd.n1332 19.3944
R6859 gnd.n1332 gnd.n1316 19.3944
R6860 gnd.n3946 gnd.n1316 19.3944
R6861 gnd.n3946 gnd.n1313 19.3944
R6862 gnd.n3951 gnd.n1313 19.3944
R6863 gnd.n3951 gnd.n1314 19.3944
R6864 gnd.n1314 gnd.n1287 19.3944
R6865 gnd.n3978 gnd.n1287 19.3944
R6866 gnd.n3978 gnd.n1284 19.3944
R6867 gnd.n3983 gnd.n1284 19.3944
R6868 gnd.n3983 gnd.n1285 19.3944
R6869 gnd.n1285 gnd.n1258 19.3944
R6870 gnd.n4012 gnd.n1258 19.3944
R6871 gnd.n4012 gnd.n1254 19.3944
R6872 gnd.n4017 gnd.n1254 19.3944
R6873 gnd.n4017 gnd.n1256 19.3944
R6874 gnd.n1256 gnd.n1255 19.3944
R6875 gnd.n1255 gnd.n52 19.3944
R6876 gnd.n6837 gnd.n52 19.3944
R6877 gnd.n6837 gnd.n6836 19.3944
R6878 gnd.n6836 gnd.n6835 19.3944
R6879 gnd.n6835 gnd.n57 19.3944
R6880 gnd.n6831 gnd.n57 19.3944
R6881 gnd.n6831 gnd.n6830 19.3944
R6882 gnd.n6830 gnd.n6829 19.3944
R6883 gnd.n6829 gnd.n62 19.3944
R6884 gnd.n6825 gnd.n62 19.3944
R6885 gnd.n6825 gnd.n6824 19.3944
R6886 gnd.n6824 gnd.n6823 19.3944
R6887 gnd.n6823 gnd.n67 19.3944
R6888 gnd.n6819 gnd.n67 19.3944
R6889 gnd.n6819 gnd.n6818 19.3944
R6890 gnd.n6818 gnd.n6817 19.3944
R6891 gnd.n6817 gnd.n72 19.3944
R6892 gnd.n6813 gnd.n72 19.3944
R6893 gnd.n6813 gnd.n6812 19.3944
R6894 gnd.n6812 gnd.n6811 19.3944
R6895 gnd.n6811 gnd.n77 19.3944
R6896 gnd.n6807 gnd.n77 19.3944
R6897 gnd.n6706 gnd.n6705 19.3944
R6898 gnd.n6705 gnd.n6704 19.3944
R6899 gnd.n6704 gnd.n6647 19.3944
R6900 gnd.n6700 gnd.n6647 19.3944
R6901 gnd.n6700 gnd.n6699 19.3944
R6902 gnd.n6699 gnd.n6698 19.3944
R6903 gnd.n6698 gnd.n6655 19.3944
R6904 gnd.n6694 gnd.n6655 19.3944
R6905 gnd.n6694 gnd.n6693 19.3944
R6906 gnd.n6693 gnd.n6692 19.3944
R6907 gnd.n6692 gnd.n6663 19.3944
R6908 gnd.n6688 gnd.n6663 19.3944
R6909 gnd.n6688 gnd.n6687 19.3944
R6910 gnd.n6687 gnd.n6686 19.3944
R6911 gnd.n6686 gnd.n6671 19.3944
R6912 gnd.n6682 gnd.n6671 19.3944
R6913 gnd.n3370 gnd.n3364 19.3944
R6914 gnd.n3376 gnd.n3364 19.3944
R6915 gnd.n3376 gnd.n3357 19.3944
R6916 gnd.n3389 gnd.n3357 19.3944
R6917 gnd.n3389 gnd.n3355 19.3944
R6918 gnd.n3395 gnd.n3355 19.3944
R6919 gnd.n3395 gnd.n3348 19.3944
R6920 gnd.n3408 gnd.n3348 19.3944
R6921 gnd.n3408 gnd.n3346 19.3944
R6922 gnd.n3414 gnd.n3346 19.3944
R6923 gnd.n3414 gnd.n3339 19.3944
R6924 gnd.n3427 gnd.n3339 19.3944
R6925 gnd.n3427 gnd.n3337 19.3944
R6926 gnd.n3433 gnd.n3337 19.3944
R6927 gnd.n3433 gnd.n3330 19.3944
R6928 gnd.n3448 gnd.n3330 19.3944
R6929 gnd.n3367 gnd.n1230 19.3944
R6930 gnd.n4046 gnd.n1230 19.3944
R6931 gnd.n4046 gnd.n1231 19.3944
R6932 gnd.n4042 gnd.n1231 19.3944
R6933 gnd.n4042 gnd.n4041 19.3944
R6934 gnd.n4041 gnd.n4040 19.3944
R6935 gnd.n4040 gnd.n1237 19.3944
R6936 gnd.n4036 gnd.n1237 19.3944
R6937 gnd.n4036 gnd.n4035 19.3944
R6938 gnd.n4035 gnd.n4034 19.3944
R6939 gnd.n4034 gnd.n1242 19.3944
R6940 gnd.n4030 gnd.n1242 19.3944
R6941 gnd.n4030 gnd.n4029 19.3944
R6942 gnd.n4029 gnd.n4028 19.3944
R6943 gnd.n4028 gnd.n1247 19.3944
R6944 gnd.n4024 gnd.n1247 19.3944
R6945 gnd.n4024 gnd.n4023 19.3944
R6946 gnd.n4023 gnd.n4022 19.3944
R6947 gnd.n4022 gnd.n242 19.3944
R6948 gnd.n6575 gnd.n242 19.3944
R6949 gnd.n6575 gnd.n239 19.3944
R6950 gnd.n6579 gnd.n239 19.3944
R6951 gnd.n6579 gnd.n228 19.3944
R6952 gnd.n6589 gnd.n228 19.3944
R6953 gnd.n6589 gnd.n226 19.3944
R6954 gnd.n6593 gnd.n226 19.3944
R6955 gnd.n6593 gnd.n207 19.3944
R6956 gnd.n6605 gnd.n207 19.3944
R6957 gnd.n6605 gnd.n205 19.3944
R6958 gnd.n6609 gnd.n205 19.3944
R6959 gnd.n6609 gnd.n192 19.3944
R6960 gnd.n6621 gnd.n192 19.3944
R6961 gnd.n6621 gnd.n190 19.3944
R6962 gnd.n6625 gnd.n190 19.3944
R6963 gnd.n6625 gnd.n177 19.3944
R6964 gnd.n6637 gnd.n177 19.3944
R6965 gnd.n6637 gnd.n174 19.3944
R6966 gnd.n6715 gnd.n174 19.3944
R6967 gnd.n6715 gnd.n175 19.3944
R6968 gnd.n6711 gnd.n175 19.3944
R6969 gnd.n6711 gnd.n6710 19.3944
R6970 gnd.n6710 gnd.n6709 19.3944
R6971 gnd.n1919 gnd.n1085 19.3944
R6972 gnd.n1919 gnd.n1869 19.3944
R6973 gnd.n2668 gnd.n1869 19.3944
R6974 gnd.n2668 gnd.n2667 19.3944
R6975 gnd.n2667 gnd.n1872 19.3944
R6976 gnd.n2660 gnd.n1872 19.3944
R6977 gnd.n2660 gnd.n2659 19.3944
R6978 gnd.n2659 gnd.n1881 19.3944
R6979 gnd.n2652 gnd.n1881 19.3944
R6980 gnd.n2652 gnd.n2651 19.3944
R6981 gnd.n2651 gnd.n1889 19.3944
R6982 gnd.n2644 gnd.n1889 19.3944
R6983 gnd.n2644 gnd.n2643 19.3944
R6984 gnd.n2643 gnd.n1899 19.3944
R6985 gnd.n2636 gnd.n1899 19.3944
R6986 gnd.n2636 gnd.n2635 19.3944
R6987 gnd.n2048 gnd.n2044 19.3944
R6988 gnd.n2048 gnd.n2041 19.3944
R6989 gnd.n2064 gnd.n2041 19.3944
R6990 gnd.n2064 gnd.n2063 19.3944
R6991 gnd.n2063 gnd.n2062 19.3944
R6992 gnd.n2062 gnd.n2059 19.3944
R6993 gnd.n2059 gnd.n2058 19.3944
R6994 gnd.n2058 gnd.n2021 19.3944
R6995 gnd.n2021 gnd.n2019 19.3944
R6996 gnd.n2305 gnd.n2019 19.3944
R6997 gnd.n2305 gnd.n2017 19.3944
R6998 gnd.n2309 gnd.n2017 19.3944
R6999 gnd.n2309 gnd.n2015 19.3944
R7000 gnd.n2313 gnd.n2015 19.3944
R7001 gnd.n2313 gnd.n2013 19.3944
R7002 gnd.n2358 gnd.n2013 19.3944
R7003 gnd.n2358 gnd.n2357 19.3944
R7004 gnd.n2357 gnd.n2356 19.3944
R7005 gnd.n2356 gnd.n2319 19.3944
R7006 gnd.n2352 gnd.n2319 19.3944
R7007 gnd.n2352 gnd.n2351 19.3944
R7008 gnd.n2351 gnd.n2350 19.3944
R7009 gnd.n2350 gnd.n2325 19.3944
R7010 gnd.n2346 gnd.n2325 19.3944
R7011 gnd.n2346 gnd.n2345 19.3944
R7012 gnd.n2345 gnd.n2344 19.3944
R7013 gnd.n2344 gnd.n2331 19.3944
R7014 gnd.n2339 gnd.n2331 19.3944
R7015 gnd.n2339 gnd.n2338 19.3944
R7016 gnd.n2338 gnd.n1841 19.3944
R7017 gnd.n2688 gnd.n1841 19.3944
R7018 gnd.n2688 gnd.n1839 19.3944
R7019 gnd.n2692 gnd.n1839 19.3944
R7020 gnd.n2692 gnd.n1828 19.3944
R7021 gnd.n2708 gnd.n1828 19.3944
R7022 gnd.n2708 gnd.n1826 19.3944
R7023 gnd.n2712 gnd.n1826 19.3944
R7024 gnd.n2712 gnd.n1815 19.3944
R7025 gnd.n2729 gnd.n1815 19.3944
R7026 gnd.n2729 gnd.n1813 19.3944
R7027 gnd.n2735 gnd.n1813 19.3944
R7028 gnd.n2735 gnd.n2734 19.3944
R7029 gnd.n2734 gnd.n1738 19.3944
R7030 gnd.n2806 gnd.n1738 19.3944
R7031 gnd.n2806 gnd.n1736 19.3944
R7032 gnd.n2812 gnd.n1736 19.3944
R7033 gnd.n2812 gnd.n2811 19.3944
R7034 gnd.n2811 gnd.n1710 19.3944
R7035 gnd.n2843 gnd.n1710 19.3944
R7036 gnd.n2843 gnd.n1708 19.3944
R7037 gnd.n2847 gnd.n1708 19.3944
R7038 gnd.n2847 gnd.n1688 19.3944
R7039 gnd.n2870 gnd.n1688 19.3944
R7040 gnd.n2870 gnd.n1686 19.3944
R7041 gnd.n2876 gnd.n1686 19.3944
R7042 gnd.n2876 gnd.n2875 19.3944
R7043 gnd.n2875 gnd.n1655 19.3944
R7044 gnd.n2912 gnd.n1655 19.3944
R7045 gnd.n2912 gnd.n1653 19.3944
R7046 gnd.n2927 gnd.n1653 19.3944
R7047 gnd.n2927 gnd.n2926 19.3944
R7048 gnd.n2926 gnd.n2925 19.3944
R7049 gnd.n2925 gnd.n2919 19.3944
R7050 gnd.n2919 gnd.n1621 19.3944
R7051 gnd.n2995 gnd.n1621 19.3944
R7052 gnd.n2995 gnd.n1619 19.3944
R7053 gnd.n2999 gnd.n1619 19.3944
R7054 gnd.n2999 gnd.n1598 19.3944
R7055 gnd.n3038 gnd.n1598 19.3944
R7056 gnd.n3038 gnd.n1596 19.3944
R7057 gnd.n3042 gnd.n1596 19.3944
R7058 gnd.n3042 gnd.n1582 19.3944
R7059 gnd.n3082 gnd.n1582 19.3944
R7060 gnd.n3082 gnd.n1580 19.3944
R7061 gnd.n3088 gnd.n1580 19.3944
R7062 gnd.n3088 gnd.n3087 19.3944
R7063 gnd.n3087 gnd.n1551 19.3944
R7064 gnd.n3128 gnd.n1551 19.3944
R7065 gnd.n3128 gnd.n1549 19.3944
R7066 gnd.n3132 gnd.n1549 19.3944
R7067 gnd.n3132 gnd.n1534 19.3944
R7068 gnd.n3189 gnd.n1534 19.3944
R7069 gnd.n3189 gnd.n1532 19.3944
R7070 gnd.n3193 gnd.n1532 19.3944
R7071 gnd.n3193 gnd.n1512 19.3944
R7072 gnd.n3217 gnd.n1512 19.3944
R7073 gnd.n3217 gnd.n1510 19.3944
R7074 gnd.n3223 gnd.n1510 19.3944
R7075 gnd.n3223 gnd.n3222 19.3944
R7076 gnd.n3222 gnd.n1484 19.3944
R7077 gnd.n3261 gnd.n1484 19.3944
R7078 gnd.n3261 gnd.n1482 19.3944
R7079 gnd.n3271 gnd.n1482 19.3944
R7080 gnd.n3271 gnd.n3270 19.3944
R7081 gnd.n3270 gnd.n3269 19.3944
R7082 gnd.n3269 gnd.n1414 19.3944
R7083 gnd.n3533 gnd.n1414 19.3944
R7084 gnd.n3533 gnd.n3532 19.3944
R7085 gnd.n3532 gnd.n3531 19.3944
R7086 gnd.n3531 gnd.n1418 19.3944
R7087 gnd.n3522 gnd.n1418 19.3944
R7088 gnd.n3522 gnd.n3521 19.3944
R7089 gnd.n3521 gnd.n3520 19.3944
R7090 gnd.n3520 gnd.n1428 19.3944
R7091 gnd.n3511 gnd.n1428 19.3944
R7092 gnd.n3511 gnd.n3510 19.3944
R7093 gnd.n3510 gnd.n3509 19.3944
R7094 gnd.n3509 gnd.n1439 19.3944
R7095 gnd.n3500 gnd.n1439 19.3944
R7096 gnd.n3500 gnd.n3499 19.3944
R7097 gnd.n3499 gnd.n1197 19.3944
R7098 gnd.n4067 gnd.n1197 19.3944
R7099 gnd.n4067 gnd.n4066 19.3944
R7100 gnd.n4066 gnd.n4065 19.3944
R7101 gnd.n4065 gnd.n1201 19.3944
R7102 gnd.n4059 gnd.n1201 19.3944
R7103 gnd.n4059 gnd.n4058 19.3944
R7104 gnd.n4058 gnd.n4057 19.3944
R7105 gnd.n4057 gnd.n1210 19.3944
R7106 gnd.n3922 gnd.n1210 19.3944
R7107 gnd.n3925 gnd.n3922 19.3944
R7108 gnd.n3925 gnd.n3919 19.3944
R7109 gnd.n3931 gnd.n3919 19.3944
R7110 gnd.n3931 gnd.n3930 19.3944
R7111 gnd.n3930 gnd.n1307 19.3944
R7112 gnd.n3956 gnd.n1307 19.3944
R7113 gnd.n3956 gnd.n1305 19.3944
R7114 gnd.n3962 gnd.n1305 19.3944
R7115 gnd.n3962 gnd.n3961 19.3944
R7116 gnd.n3961 gnd.n1279 19.3944
R7117 gnd.n3988 gnd.n1279 19.3944
R7118 gnd.n3988 gnd.n1277 19.3944
R7119 gnd.n4001 gnd.n1277 19.3944
R7120 gnd.n4001 gnd.n4000 19.3944
R7121 gnd.n4000 gnd.n3999 19.3944
R7122 gnd.n3999 gnd.n3995 19.3944
R7123 gnd.n3995 gnd.n253 19.3944
R7124 gnd.n6565 gnd.n253 19.3944
R7125 gnd.n6565 gnd.n6564 19.3944
R7126 gnd.n6564 gnd.n6563 19.3944
R7127 gnd.n6563 gnd.n257 19.3944
R7128 gnd.n6346 gnd.n381 19.3944
R7129 gnd.n6352 gnd.n381 19.3944
R7130 gnd.n6352 gnd.n379 19.3944
R7131 gnd.n6356 gnd.n379 19.3944
R7132 gnd.n6356 gnd.n375 19.3944
R7133 gnd.n6362 gnd.n375 19.3944
R7134 gnd.n6362 gnd.n373 19.3944
R7135 gnd.n6366 gnd.n373 19.3944
R7136 gnd.n6366 gnd.n369 19.3944
R7137 gnd.n6372 gnd.n369 19.3944
R7138 gnd.n6372 gnd.n367 19.3944
R7139 gnd.n6376 gnd.n367 19.3944
R7140 gnd.n6376 gnd.n363 19.3944
R7141 gnd.n6382 gnd.n363 19.3944
R7142 gnd.n6382 gnd.n361 19.3944
R7143 gnd.n6386 gnd.n361 19.3944
R7144 gnd.n6386 gnd.n357 19.3944
R7145 gnd.n6392 gnd.n357 19.3944
R7146 gnd.n6392 gnd.n355 19.3944
R7147 gnd.n6396 gnd.n355 19.3944
R7148 gnd.n6396 gnd.n351 19.3944
R7149 gnd.n6402 gnd.n351 19.3944
R7150 gnd.n6402 gnd.n349 19.3944
R7151 gnd.n6406 gnd.n349 19.3944
R7152 gnd.n6406 gnd.n345 19.3944
R7153 gnd.n6412 gnd.n345 19.3944
R7154 gnd.n6412 gnd.n343 19.3944
R7155 gnd.n6416 gnd.n343 19.3944
R7156 gnd.n6416 gnd.n339 19.3944
R7157 gnd.n6422 gnd.n339 19.3944
R7158 gnd.n6422 gnd.n337 19.3944
R7159 gnd.n6426 gnd.n337 19.3944
R7160 gnd.n6426 gnd.n333 19.3944
R7161 gnd.n6432 gnd.n333 19.3944
R7162 gnd.n6432 gnd.n331 19.3944
R7163 gnd.n6436 gnd.n331 19.3944
R7164 gnd.n6436 gnd.n327 19.3944
R7165 gnd.n6442 gnd.n327 19.3944
R7166 gnd.n6442 gnd.n325 19.3944
R7167 gnd.n6446 gnd.n325 19.3944
R7168 gnd.n6446 gnd.n321 19.3944
R7169 gnd.n6452 gnd.n321 19.3944
R7170 gnd.n6452 gnd.n319 19.3944
R7171 gnd.n6456 gnd.n319 19.3944
R7172 gnd.n6456 gnd.n315 19.3944
R7173 gnd.n6462 gnd.n315 19.3944
R7174 gnd.n6462 gnd.n313 19.3944
R7175 gnd.n6466 gnd.n313 19.3944
R7176 gnd.n6466 gnd.n309 19.3944
R7177 gnd.n6472 gnd.n309 19.3944
R7178 gnd.n6472 gnd.n307 19.3944
R7179 gnd.n6476 gnd.n307 19.3944
R7180 gnd.n6476 gnd.n303 19.3944
R7181 gnd.n6482 gnd.n303 19.3944
R7182 gnd.n6482 gnd.n301 19.3944
R7183 gnd.n6486 gnd.n301 19.3944
R7184 gnd.n6486 gnd.n297 19.3944
R7185 gnd.n6492 gnd.n297 19.3944
R7186 gnd.n6492 gnd.n295 19.3944
R7187 gnd.n6496 gnd.n295 19.3944
R7188 gnd.n6496 gnd.n291 19.3944
R7189 gnd.n6502 gnd.n291 19.3944
R7190 gnd.n6502 gnd.n289 19.3944
R7191 gnd.n6506 gnd.n289 19.3944
R7192 gnd.n6506 gnd.n285 19.3944
R7193 gnd.n6512 gnd.n285 19.3944
R7194 gnd.n6512 gnd.n283 19.3944
R7195 gnd.n6516 gnd.n283 19.3944
R7196 gnd.n6516 gnd.n279 19.3944
R7197 gnd.n6522 gnd.n279 19.3944
R7198 gnd.n6522 gnd.n277 19.3944
R7199 gnd.n6526 gnd.n277 19.3944
R7200 gnd.n6526 gnd.n273 19.3944
R7201 gnd.n6532 gnd.n273 19.3944
R7202 gnd.n6532 gnd.n271 19.3944
R7203 gnd.n6536 gnd.n271 19.3944
R7204 gnd.n6536 gnd.n267 19.3944
R7205 gnd.n6542 gnd.n267 19.3944
R7206 gnd.n6542 gnd.n265 19.3944
R7207 gnd.n6546 gnd.n265 19.3944
R7208 gnd.n6546 gnd.n261 19.3944
R7209 gnd.n6553 gnd.n261 19.3944
R7210 gnd.n6553 gnd.n259 19.3944
R7211 gnd.n6558 gnd.n259 19.3944
R7212 gnd.n5991 gnd.n594 19.3944
R7213 gnd.n5995 gnd.n594 19.3944
R7214 gnd.n5995 gnd.n590 19.3944
R7215 gnd.n6001 gnd.n590 19.3944
R7216 gnd.n6001 gnd.n588 19.3944
R7217 gnd.n6005 gnd.n588 19.3944
R7218 gnd.n6005 gnd.n584 19.3944
R7219 gnd.n6011 gnd.n584 19.3944
R7220 gnd.n6011 gnd.n582 19.3944
R7221 gnd.n6015 gnd.n582 19.3944
R7222 gnd.n6015 gnd.n578 19.3944
R7223 gnd.n6021 gnd.n578 19.3944
R7224 gnd.n6021 gnd.n576 19.3944
R7225 gnd.n6025 gnd.n576 19.3944
R7226 gnd.n6025 gnd.n572 19.3944
R7227 gnd.n6031 gnd.n572 19.3944
R7228 gnd.n6031 gnd.n570 19.3944
R7229 gnd.n6035 gnd.n570 19.3944
R7230 gnd.n6035 gnd.n566 19.3944
R7231 gnd.n6041 gnd.n566 19.3944
R7232 gnd.n6041 gnd.n564 19.3944
R7233 gnd.n6045 gnd.n564 19.3944
R7234 gnd.n6045 gnd.n560 19.3944
R7235 gnd.n6051 gnd.n560 19.3944
R7236 gnd.n6051 gnd.n558 19.3944
R7237 gnd.n6055 gnd.n558 19.3944
R7238 gnd.n6055 gnd.n554 19.3944
R7239 gnd.n6061 gnd.n554 19.3944
R7240 gnd.n6061 gnd.n552 19.3944
R7241 gnd.n6065 gnd.n552 19.3944
R7242 gnd.n6065 gnd.n548 19.3944
R7243 gnd.n6071 gnd.n548 19.3944
R7244 gnd.n6071 gnd.n546 19.3944
R7245 gnd.n6075 gnd.n546 19.3944
R7246 gnd.n6075 gnd.n542 19.3944
R7247 gnd.n6081 gnd.n542 19.3944
R7248 gnd.n6081 gnd.n540 19.3944
R7249 gnd.n6085 gnd.n540 19.3944
R7250 gnd.n6085 gnd.n536 19.3944
R7251 gnd.n6091 gnd.n536 19.3944
R7252 gnd.n6091 gnd.n534 19.3944
R7253 gnd.n6095 gnd.n534 19.3944
R7254 gnd.n6095 gnd.n530 19.3944
R7255 gnd.n6101 gnd.n530 19.3944
R7256 gnd.n6101 gnd.n528 19.3944
R7257 gnd.n6105 gnd.n528 19.3944
R7258 gnd.n6105 gnd.n524 19.3944
R7259 gnd.n6111 gnd.n524 19.3944
R7260 gnd.n6111 gnd.n522 19.3944
R7261 gnd.n6115 gnd.n522 19.3944
R7262 gnd.n6115 gnd.n518 19.3944
R7263 gnd.n6121 gnd.n518 19.3944
R7264 gnd.n6121 gnd.n516 19.3944
R7265 gnd.n6125 gnd.n516 19.3944
R7266 gnd.n6125 gnd.n512 19.3944
R7267 gnd.n6131 gnd.n512 19.3944
R7268 gnd.n6131 gnd.n510 19.3944
R7269 gnd.n6135 gnd.n510 19.3944
R7270 gnd.n6135 gnd.n506 19.3944
R7271 gnd.n6141 gnd.n506 19.3944
R7272 gnd.n6141 gnd.n504 19.3944
R7273 gnd.n6145 gnd.n504 19.3944
R7274 gnd.n6145 gnd.n500 19.3944
R7275 gnd.n6151 gnd.n500 19.3944
R7276 gnd.n6151 gnd.n498 19.3944
R7277 gnd.n6155 gnd.n498 19.3944
R7278 gnd.n6155 gnd.n494 19.3944
R7279 gnd.n6161 gnd.n494 19.3944
R7280 gnd.n6161 gnd.n492 19.3944
R7281 gnd.n6165 gnd.n492 19.3944
R7282 gnd.n6165 gnd.n488 19.3944
R7283 gnd.n6171 gnd.n488 19.3944
R7284 gnd.n6171 gnd.n486 19.3944
R7285 gnd.n6175 gnd.n486 19.3944
R7286 gnd.n6175 gnd.n482 19.3944
R7287 gnd.n6181 gnd.n482 19.3944
R7288 gnd.n6181 gnd.n480 19.3944
R7289 gnd.n6185 gnd.n480 19.3944
R7290 gnd.n6185 gnd.n476 19.3944
R7291 gnd.n6191 gnd.n476 19.3944
R7292 gnd.n6191 gnd.n474 19.3944
R7293 gnd.n6195 gnd.n474 19.3944
R7294 gnd.n6195 gnd.n470 19.3944
R7295 gnd.n6201 gnd.n470 19.3944
R7296 gnd.n6201 gnd.n468 19.3944
R7297 gnd.n6205 gnd.n468 19.3944
R7298 gnd.n6205 gnd.n464 19.3944
R7299 gnd.n6211 gnd.n464 19.3944
R7300 gnd.n6211 gnd.n462 19.3944
R7301 gnd.n6215 gnd.n462 19.3944
R7302 gnd.n6215 gnd.n458 19.3944
R7303 gnd.n6221 gnd.n458 19.3944
R7304 gnd.n6221 gnd.n456 19.3944
R7305 gnd.n6225 gnd.n456 19.3944
R7306 gnd.n6225 gnd.n452 19.3944
R7307 gnd.n6231 gnd.n452 19.3944
R7308 gnd.n6231 gnd.n450 19.3944
R7309 gnd.n6235 gnd.n450 19.3944
R7310 gnd.n6235 gnd.n446 19.3944
R7311 gnd.n6241 gnd.n446 19.3944
R7312 gnd.n6241 gnd.n444 19.3944
R7313 gnd.n6245 gnd.n444 19.3944
R7314 gnd.n6245 gnd.n440 19.3944
R7315 gnd.n6251 gnd.n440 19.3944
R7316 gnd.n6251 gnd.n438 19.3944
R7317 gnd.n6255 gnd.n438 19.3944
R7318 gnd.n6255 gnd.n434 19.3944
R7319 gnd.n6261 gnd.n434 19.3944
R7320 gnd.n6261 gnd.n432 19.3944
R7321 gnd.n6265 gnd.n432 19.3944
R7322 gnd.n6265 gnd.n428 19.3944
R7323 gnd.n6271 gnd.n428 19.3944
R7324 gnd.n6271 gnd.n426 19.3944
R7325 gnd.n6275 gnd.n426 19.3944
R7326 gnd.n6275 gnd.n422 19.3944
R7327 gnd.n6281 gnd.n422 19.3944
R7328 gnd.n6281 gnd.n420 19.3944
R7329 gnd.n6285 gnd.n420 19.3944
R7330 gnd.n6285 gnd.n416 19.3944
R7331 gnd.n6291 gnd.n416 19.3944
R7332 gnd.n6291 gnd.n414 19.3944
R7333 gnd.n6295 gnd.n414 19.3944
R7334 gnd.n6295 gnd.n410 19.3944
R7335 gnd.n6301 gnd.n410 19.3944
R7336 gnd.n6301 gnd.n408 19.3944
R7337 gnd.n6305 gnd.n408 19.3944
R7338 gnd.n6305 gnd.n404 19.3944
R7339 gnd.n6311 gnd.n404 19.3944
R7340 gnd.n6311 gnd.n402 19.3944
R7341 gnd.n6315 gnd.n402 19.3944
R7342 gnd.n6315 gnd.n398 19.3944
R7343 gnd.n6321 gnd.n398 19.3944
R7344 gnd.n6321 gnd.n396 19.3944
R7345 gnd.n6325 gnd.n396 19.3944
R7346 gnd.n6325 gnd.n392 19.3944
R7347 gnd.n6331 gnd.n392 19.3944
R7348 gnd.n6331 gnd.n390 19.3944
R7349 gnd.n6336 gnd.n390 19.3944
R7350 gnd.n6336 gnd.n386 19.3944
R7351 gnd.n6342 gnd.n386 19.3944
R7352 gnd.n6343 gnd.n6342 19.3944
R7353 gnd.n3716 gnd.n3713 19.3944
R7354 gnd.n3716 gnd.n3712 19.3944
R7355 gnd.n3722 gnd.n3712 19.3944
R7356 gnd.n3722 gnd.n3710 19.3944
R7357 gnd.n3726 gnd.n3710 19.3944
R7358 gnd.n3726 gnd.n3708 19.3944
R7359 gnd.n3732 gnd.n3708 19.3944
R7360 gnd.n3732 gnd.n3706 19.3944
R7361 gnd.n3736 gnd.n3706 19.3944
R7362 gnd.n3736 gnd.n3704 19.3944
R7363 gnd.n3742 gnd.n3704 19.3944
R7364 gnd.n3742 gnd.n3702 19.3944
R7365 gnd.n3747 gnd.n3702 19.3944
R7366 gnd.n3747 gnd.n3700 19.3944
R7367 gnd.n3700 gnd.n1360 19.3944
R7368 gnd.n3760 gnd.n1358 19.3944
R7369 gnd.n3760 gnd.n1356 19.3944
R7370 gnd.n3766 gnd.n1356 19.3944
R7371 gnd.n3766 gnd.n1354 19.3944
R7372 gnd.n3770 gnd.n1354 19.3944
R7373 gnd.n3770 gnd.n1352 19.3944
R7374 gnd.n3776 gnd.n1352 19.3944
R7375 gnd.n3776 gnd.n1350 19.3944
R7376 gnd.n3780 gnd.n1350 19.3944
R7377 gnd.n3780 gnd.n1348 19.3944
R7378 gnd.n3786 gnd.n1348 19.3944
R7379 gnd.n3786 gnd.n1346 19.3944
R7380 gnd.n3790 gnd.n1346 19.3944
R7381 gnd.n3790 gnd.n1344 19.3944
R7382 gnd.n3796 gnd.n1344 19.3944
R7383 gnd.n3796 gnd.n1342 19.3944
R7384 gnd.n3801 gnd.n1342 19.3944
R7385 gnd.n3801 gnd.n1340 19.3944
R7386 gnd.n3812 gnd.n1335 19.3944
R7387 gnd.n3812 gnd.n1330 19.3944
R7388 gnd.n3825 gnd.n1330 19.3944
R7389 gnd.n3825 gnd.n1328 19.3944
R7390 gnd.n3914 gnd.n1328 19.3944
R7391 gnd.n3914 gnd.n3913 19.3944
R7392 gnd.n3913 gnd.n3912 19.3944
R7393 gnd.n3912 gnd.n3910 19.3944
R7394 gnd.n3910 gnd.n3909 19.3944
R7395 gnd.n3909 gnd.n3908 19.3944
R7396 gnd.n3908 gnd.n3906 19.3944
R7397 gnd.n3906 gnd.n3905 19.3944
R7398 gnd.n3905 gnd.n3903 19.3944
R7399 gnd.n3903 gnd.n3902 19.3944
R7400 gnd.n3902 gnd.n3901 19.3944
R7401 gnd.n3901 gnd.n3899 19.3944
R7402 gnd.n3899 gnd.n3898 19.3944
R7403 gnd.n3898 gnd.n3895 19.3944
R7404 gnd.n3895 gnd.n3894 19.3944
R7405 gnd.n3894 gnd.n3893 19.3944
R7406 gnd.n3893 gnd.n3892 19.3944
R7407 gnd.n3892 gnd.n3888 19.3944
R7408 gnd.n3888 gnd.n3887 19.3944
R7409 gnd.n3887 gnd.n3885 19.3944
R7410 gnd.n3885 gnd.n3884 19.3944
R7411 gnd.n3884 gnd.n3882 19.3944
R7412 gnd.n3882 gnd.n3881 19.3944
R7413 gnd.n3881 gnd.n3879 19.3944
R7414 gnd.n3879 gnd.n3878 19.3944
R7415 gnd.n3878 gnd.n3876 19.3944
R7416 gnd.n3876 gnd.n3875 19.3944
R7417 gnd.n3875 gnd.n3873 19.3944
R7418 gnd.n3873 gnd.n3872 19.3944
R7419 gnd.n3872 gnd.n3870 19.3944
R7420 gnd.n3870 gnd.n3869 19.3944
R7421 gnd.n3869 gnd.n3867 19.3944
R7422 gnd.n3867 gnd.n3866 19.3944
R7423 gnd.n3866 gnd.n3864 19.3944
R7424 gnd.n3864 gnd.n3863 19.3944
R7425 gnd.n3863 gnd.n159 19.3944
R7426 gnd.n6728 gnd.n159 19.3944
R7427 gnd.n6729 gnd.n6728 19.3944
R7428 gnd.n6767 gnd.n120 19.3944
R7429 gnd.n6762 gnd.n120 19.3944
R7430 gnd.n6762 gnd.n6761 19.3944
R7431 gnd.n6761 gnd.n6760 19.3944
R7432 gnd.n6760 gnd.n127 19.3944
R7433 gnd.n6755 gnd.n127 19.3944
R7434 gnd.n6755 gnd.n6754 19.3944
R7435 gnd.n6754 gnd.n6753 19.3944
R7436 gnd.n6753 gnd.n134 19.3944
R7437 gnd.n6748 gnd.n134 19.3944
R7438 gnd.n6748 gnd.n6747 19.3944
R7439 gnd.n6747 gnd.n6746 19.3944
R7440 gnd.n6746 gnd.n141 19.3944
R7441 gnd.n6741 gnd.n141 19.3944
R7442 gnd.n6741 gnd.n6740 19.3944
R7443 gnd.n6740 gnd.n6739 19.3944
R7444 gnd.n6739 gnd.n148 19.3944
R7445 gnd.n6734 gnd.n148 19.3944
R7446 gnd.n6800 gnd.n6799 19.3944
R7447 gnd.n6799 gnd.n6798 19.3944
R7448 gnd.n6798 gnd.n92 19.3944
R7449 gnd.n6793 gnd.n92 19.3944
R7450 gnd.n6793 gnd.n6792 19.3944
R7451 gnd.n6792 gnd.n6791 19.3944
R7452 gnd.n6791 gnd.n99 19.3944
R7453 gnd.n6786 gnd.n99 19.3944
R7454 gnd.n6786 gnd.n6785 19.3944
R7455 gnd.n6785 gnd.n6784 19.3944
R7456 gnd.n6784 gnd.n106 19.3944
R7457 gnd.n6779 gnd.n106 19.3944
R7458 gnd.n6779 gnd.n6778 19.3944
R7459 gnd.n6778 gnd.n6777 19.3944
R7460 gnd.n6777 gnd.n113 19.3944
R7461 gnd.n6772 gnd.n113 19.3944
R7462 gnd.n6772 gnd.n6771 19.3944
R7463 gnd.n4052 gnd.n4051 19.3944
R7464 gnd.n4051 gnd.n4050 19.3944
R7465 gnd.n4050 gnd.n1222 19.3944
R7466 gnd.n3936 gnd.n1222 19.3944
R7467 gnd.n3936 gnd.n1323 19.3944
R7468 gnd.n3942 gnd.n1323 19.3944
R7469 gnd.n3942 gnd.n3941 19.3944
R7470 gnd.n3941 gnd.n1297 19.3944
R7471 gnd.n3967 gnd.n1297 19.3944
R7472 gnd.n3967 gnd.n1295 19.3944
R7473 gnd.n3974 gnd.n1295 19.3944
R7474 gnd.n3974 gnd.n3973 19.3944
R7475 gnd.n3973 gnd.n1267 19.3944
R7476 gnd.n4006 gnd.n1267 19.3944
R7477 gnd.n4007 gnd.n4006 19.3944
R7478 gnd.n4008 gnd.n4007 19.3944
R7479 gnd.n1265 gnd.n1264 19.3944
R7480 gnd.n6571 gnd.n6570 19.3944
R7481 gnd.n235 gnd.n234 19.3944
R7482 gnd.n6585 gnd.n6584 19.3944
R7483 gnd.n6597 gnd.n219 19.3944
R7484 gnd.n6597 gnd.n211 19.3944
R7485 gnd.n6601 gnd.n211 19.3944
R7486 gnd.n6601 gnd.n199 19.3944
R7487 gnd.n6613 gnd.n199 19.3944
R7488 gnd.n6613 gnd.n197 19.3944
R7489 gnd.n6617 gnd.n197 19.3944
R7490 gnd.n6617 gnd.n183 19.3944
R7491 gnd.n6629 gnd.n183 19.3944
R7492 gnd.n6629 gnd.n181 19.3944
R7493 gnd.n6633 gnd.n181 19.3944
R7494 gnd.n6633 gnd.n167 19.3944
R7495 gnd.n6719 gnd.n167 19.3944
R7496 gnd.n6719 gnd.n165 19.3944
R7497 gnd.n6723 gnd.n165 19.3944
R7498 gnd.n6723 gnd.n87 19.3944
R7499 gnd.n6803 gnd.n87 19.3944
R7500 gnd.n4403 gnd.n4402 19.3944
R7501 gnd.n4402 gnd.n4401 19.3944
R7502 gnd.n4401 gnd.n4400 19.3944
R7503 gnd.n4400 gnd.n4398 19.3944
R7504 gnd.n4398 gnd.n4395 19.3944
R7505 gnd.n4395 gnd.n4394 19.3944
R7506 gnd.n4394 gnd.n4391 19.3944
R7507 gnd.n4391 gnd.n4390 19.3944
R7508 gnd.n4390 gnd.n4387 19.3944
R7509 gnd.n4387 gnd.n4386 19.3944
R7510 gnd.n4386 gnd.n4383 19.3944
R7511 gnd.n4383 gnd.n4382 19.3944
R7512 gnd.n4382 gnd.n4379 19.3944
R7513 gnd.n4379 gnd.n4378 19.3944
R7514 gnd.n4378 gnd.n4375 19.3944
R7515 gnd.n4375 gnd.n4374 19.3944
R7516 gnd.n4374 gnd.n4371 19.3944
R7517 gnd.n4369 gnd.n4366 19.3944
R7518 gnd.n4366 gnd.n4365 19.3944
R7519 gnd.n4365 gnd.n4362 19.3944
R7520 gnd.n4362 gnd.n4361 19.3944
R7521 gnd.n4361 gnd.n4358 19.3944
R7522 gnd.n4358 gnd.n4357 19.3944
R7523 gnd.n4357 gnd.n4354 19.3944
R7524 gnd.n4354 gnd.n4353 19.3944
R7525 gnd.n4353 gnd.n4350 19.3944
R7526 gnd.n4350 gnd.n4349 19.3944
R7527 gnd.n4349 gnd.n4346 19.3944
R7528 gnd.n4346 gnd.n4345 19.3944
R7529 gnd.n4345 gnd.n4342 19.3944
R7530 gnd.n4342 gnd.n4341 19.3944
R7531 gnd.n4341 gnd.n4338 19.3944
R7532 gnd.n4338 gnd.n4337 19.3944
R7533 gnd.n4337 gnd.n4334 19.3944
R7534 gnd.n4334 gnd.n4333 19.3944
R7535 gnd.n2157 gnd.n2088 19.3944
R7536 gnd.n2157 gnd.n2089 19.3944
R7537 gnd.n2153 gnd.n2089 19.3944
R7538 gnd.n2153 gnd.n901 19.3944
R7539 gnd.n4311 gnd.n901 19.3944
R7540 gnd.n4311 gnd.n4310 19.3944
R7541 gnd.n4310 gnd.n4309 19.3944
R7542 gnd.n4309 gnd.n905 19.3944
R7543 gnd.n4299 gnd.n905 19.3944
R7544 gnd.n4299 gnd.n4298 19.3944
R7545 gnd.n4298 gnd.n4297 19.3944
R7546 gnd.n4297 gnd.n924 19.3944
R7547 gnd.n4287 gnd.n924 19.3944
R7548 gnd.n4287 gnd.n4286 19.3944
R7549 gnd.n4286 gnd.n4285 19.3944
R7550 gnd.n4285 gnd.n945 19.3944
R7551 gnd.n963 gnd.n945 19.3944
R7552 gnd.n4273 gnd.n963 19.3944
R7553 gnd.n4273 gnd.n4272 19.3944
R7554 gnd.n4272 gnd.n4271 19.3944
R7555 gnd.n4271 gnd.n969 19.3944
R7556 gnd.n4260 gnd.n969 19.3944
R7557 gnd.n4260 gnd.n4259 19.3944
R7558 gnd.n4259 gnd.n4258 19.3944
R7559 gnd.n4258 gnd.n985 19.3944
R7560 gnd.n4247 gnd.n985 19.3944
R7561 gnd.n4247 gnd.n4246 19.3944
R7562 gnd.n4246 gnd.n4245 19.3944
R7563 gnd.n4245 gnd.n1004 19.3944
R7564 gnd.n4235 gnd.n1004 19.3944
R7565 gnd.n4235 gnd.n4234 19.3944
R7566 gnd.n4234 gnd.n4233 19.3944
R7567 gnd.n4233 gnd.n1024 19.3944
R7568 gnd.n4223 gnd.n1024 19.3944
R7569 gnd.n4223 gnd.n4222 19.3944
R7570 gnd.n4222 gnd.n4221 19.3944
R7571 gnd.n4221 gnd.n1046 19.3944
R7572 gnd.n4211 gnd.n1046 19.3944
R7573 gnd.n4211 gnd.n4210 19.3944
R7574 gnd.n4210 gnd.n4209 19.3944
R7575 gnd.n4209 gnd.n1067 19.3944
R7576 gnd.n4199 gnd.n1067 19.3944
R7577 gnd.n2149 gnd.n2147 19.3944
R7578 gnd.n2147 gnd.n2144 19.3944
R7579 gnd.n2144 gnd.n2143 19.3944
R7580 gnd.n2143 gnd.n2140 19.3944
R7581 gnd.n2140 gnd.n2139 19.3944
R7582 gnd.n2139 gnd.n2136 19.3944
R7583 gnd.n2136 gnd.n2135 19.3944
R7584 gnd.n2135 gnd.n2132 19.3944
R7585 gnd.n2132 gnd.n2131 19.3944
R7586 gnd.n2131 gnd.n2128 19.3944
R7587 gnd.n2128 gnd.n2127 19.3944
R7588 gnd.n2127 gnd.n2124 19.3944
R7589 gnd.n2124 gnd.n2123 19.3944
R7590 gnd.n2123 gnd.n2120 19.3944
R7591 gnd.n2120 gnd.n2119 19.3944
R7592 gnd.n2119 gnd.n2116 19.3944
R7593 gnd.n2110 gnd.n2084 19.3944
R7594 gnd.n2168 gnd.n2084 19.3944
R7595 gnd.n2169 gnd.n2168 19.3944
R7596 gnd.n2169 gnd.n2082 19.3944
R7597 gnd.n2173 gnd.n2082 19.3944
R7598 gnd.n2175 gnd.n2173 19.3944
R7599 gnd.n2176 gnd.n2175 19.3944
R7600 gnd.n2176 gnd.n2079 19.3944
R7601 gnd.n2180 gnd.n2079 19.3944
R7602 gnd.n2182 gnd.n2180 19.3944
R7603 gnd.n2183 gnd.n2182 19.3944
R7604 gnd.n2183 gnd.n2076 19.3944
R7605 gnd.n2187 gnd.n2076 19.3944
R7606 gnd.n2189 gnd.n2187 19.3944
R7607 gnd.n2190 gnd.n2189 19.3944
R7608 gnd.n2190 gnd.n2073 19.3944
R7609 gnd.n2235 gnd.n2073 19.3944
R7610 gnd.n2236 gnd.n2235 19.3944
R7611 gnd.n2238 gnd.n2236 19.3944
R7612 gnd.n2238 gnd.n2071 19.3944
R7613 gnd.n2242 gnd.n2071 19.3944
R7614 gnd.n2242 gnd.n2038 19.3944
R7615 gnd.n2255 gnd.n2038 19.3944
R7616 gnd.n2255 gnd.n2036 19.3944
R7617 gnd.n2259 gnd.n2036 19.3944
R7618 gnd.n2259 gnd.n2023 19.3944
R7619 gnd.n2298 gnd.n2023 19.3944
R7620 gnd.n2298 gnd.n2024 19.3944
R7621 gnd.n2294 gnd.n2024 19.3944
R7622 gnd.n2294 gnd.n2293 19.3944
R7623 gnd.n2293 gnd.n2292 19.3944
R7624 gnd.n2292 gnd.n2029 19.3944
R7625 gnd.n2288 gnd.n2029 19.3944
R7626 gnd.n2288 gnd.n2009 19.3944
R7627 gnd.n2363 gnd.n2009 19.3944
R7628 gnd.n2363 gnd.n2007 19.3944
R7629 gnd.n2367 gnd.n2007 19.3944
R7630 gnd.n2367 gnd.n2003 19.3944
R7631 gnd.n2380 gnd.n2003 19.3944
R7632 gnd.n2380 gnd.n2000 19.3944
R7633 gnd.n2416 gnd.n2000 19.3944
R7634 gnd.n2416 gnd.n2001 19.3944
R7635 gnd.n4326 gnd.n4325 19.3944
R7636 gnd.n4325 gnd.n879 19.3944
R7637 gnd.n4321 gnd.n879 19.3944
R7638 gnd.n4321 gnd.n881 19.3944
R7639 gnd.n2205 gnd.n881 19.3944
R7640 gnd.n2207 gnd.n2205 19.3944
R7641 gnd.n2208 gnd.n2207 19.3944
R7642 gnd.n2208 gnd.n2202 19.3944
R7643 gnd.n2212 gnd.n2202 19.3944
R7644 gnd.n2214 gnd.n2212 19.3944
R7645 gnd.n2215 gnd.n2214 19.3944
R7646 gnd.n2215 gnd.n2199 19.3944
R7647 gnd.n2219 gnd.n2199 19.3944
R7648 gnd.n2221 gnd.n2219 19.3944
R7649 gnd.n2222 gnd.n2221 19.3944
R7650 gnd.n2222 gnd.n2196 19.3944
R7651 gnd.n2231 gnd.n2196 19.3944
R7652 gnd.n2231 gnd.n2230 19.3944
R7653 gnd.n2230 gnd.n2229 19.3944
R7654 gnd.n2229 gnd.n2070 19.3944
R7655 gnd.n2246 gnd.n2070 19.3944
R7656 gnd.n2246 gnd.n2067 19.3944
R7657 gnd.n2251 gnd.n2067 19.3944
R7658 gnd.n2251 gnd.n2034 19.3944
R7659 gnd.n2263 gnd.n2034 19.3944
R7660 gnd.n2264 gnd.n2263 19.3944
R7661 gnd.n2265 gnd.n2264 19.3944
R7662 gnd.n2265 gnd.n2032 19.3944
R7663 gnd.n2271 gnd.n2032 19.3944
R7664 gnd.n2272 gnd.n2271 19.3944
R7665 gnd.n2276 gnd.n2272 19.3944
R7666 gnd.n2276 gnd.n2030 19.3944
R7667 gnd.n2284 gnd.n2030 19.3944
R7668 gnd.n2284 gnd.n2283 19.3944
R7669 gnd.n2283 gnd.n2282 19.3944
R7670 gnd.n2282 gnd.n2006 19.3944
R7671 gnd.n2371 gnd.n2006 19.3944
R7672 gnd.n2371 gnd.n2004 19.3944
R7673 gnd.n2376 gnd.n2004 19.3944
R7674 gnd.n2376 gnd.n1999 19.3944
R7675 gnd.n2420 gnd.n1999 19.3944
R7676 gnd.n2421 gnd.n2420 19.3944
R7677 gnd.n2463 gnd.n1973 19.3944
R7678 gnd.n2463 gnd.n2460 19.3944
R7679 gnd.n2460 gnd.n2457 19.3944
R7680 gnd.n2457 gnd.n2456 19.3944
R7681 gnd.n2456 gnd.n2453 19.3944
R7682 gnd.n2453 gnd.n2452 19.3944
R7683 gnd.n2452 gnd.n2449 19.3944
R7684 gnd.n2449 gnd.n2448 19.3944
R7685 gnd.n2448 gnd.n2445 19.3944
R7686 gnd.n2445 gnd.n2444 19.3944
R7687 gnd.n2444 gnd.n2441 19.3944
R7688 gnd.n2441 gnd.n2440 19.3944
R7689 gnd.n2440 gnd.n2437 19.3944
R7690 gnd.n2437 gnd.n2436 19.3944
R7691 gnd.n2436 gnd.n2433 19.3944
R7692 gnd.n2433 gnd.n2432 19.3944
R7693 gnd.n2432 gnd.n2429 19.3944
R7694 gnd.n2429 gnd.n2428 19.3944
R7695 gnd.n1956 gnd.n1955 19.3944
R7696 gnd.n2622 gnd.n1955 19.3944
R7697 gnd.n2622 gnd.n2621 19.3944
R7698 gnd.n2621 gnd.n2620 19.3944
R7699 gnd.n2620 gnd.n2617 19.3944
R7700 gnd.n2617 gnd.n2616 19.3944
R7701 gnd.n2616 gnd.n2613 19.3944
R7702 gnd.n2613 gnd.n2612 19.3944
R7703 gnd.n2612 gnd.n2609 19.3944
R7704 gnd.n2609 gnd.n2608 19.3944
R7705 gnd.n2608 gnd.n2605 19.3944
R7706 gnd.n2605 gnd.n2604 19.3944
R7707 gnd.n2604 gnd.n2601 19.3944
R7708 gnd.n2601 gnd.n2600 19.3944
R7709 gnd.n2600 gnd.n2597 19.3944
R7710 gnd.n2163 gnd.n2159 19.3944
R7711 gnd.n2163 gnd.n890 19.3944
R7712 gnd.n4317 gnd.n890 19.3944
R7713 gnd.n4317 gnd.n4316 19.3944
R7714 gnd.n4316 gnd.n4315 19.3944
R7715 gnd.n4315 gnd.n894 19.3944
R7716 gnd.n4305 gnd.n894 19.3944
R7717 gnd.n4305 gnd.n4304 19.3944
R7718 gnd.n4304 gnd.n4303 19.3944
R7719 gnd.n4303 gnd.n915 19.3944
R7720 gnd.n4293 gnd.n915 19.3944
R7721 gnd.n4293 gnd.n4292 19.3944
R7722 gnd.n4292 gnd.n4291 19.3944
R7723 gnd.n4291 gnd.n934 19.3944
R7724 gnd.n4281 gnd.n934 19.3944
R7725 gnd.n4281 gnd.n4280 19.3944
R7726 gnd.n4278 gnd.n4277 19.3944
R7727 gnd.n4267 gnd.n975 19.3944
R7728 gnd.n4265 gnd.n4264 19.3944
R7729 gnd.n4254 gnd.n992 19.3944
R7730 gnd.n4252 gnd.n4251 19.3944
R7731 gnd.n4251 gnd.n993 19.3944
R7732 gnd.n4241 gnd.n993 19.3944
R7733 gnd.n4241 gnd.n4240 19.3944
R7734 gnd.n4240 gnd.n4239 19.3944
R7735 gnd.n4239 gnd.n1014 19.3944
R7736 gnd.n4229 gnd.n1014 19.3944
R7737 gnd.n4229 gnd.n4228 19.3944
R7738 gnd.n4228 gnd.n4227 19.3944
R7739 gnd.n4227 gnd.n1035 19.3944
R7740 gnd.n4217 gnd.n1035 19.3944
R7741 gnd.n4217 gnd.n4216 19.3944
R7742 gnd.n4216 gnd.n4215 19.3944
R7743 gnd.n4215 gnd.n1056 19.3944
R7744 gnd.n4205 gnd.n1056 19.3944
R7745 gnd.n4205 gnd.n4204 19.3944
R7746 gnd.n4204 gnd.n4203 19.3944
R7747 gnd.n5985 gnd.n599 19.3944
R7748 gnd.n5985 gnd.n5984 19.3944
R7749 gnd.n5984 gnd.n5983 19.3944
R7750 gnd.n5983 gnd.n603 19.3944
R7751 gnd.n5977 gnd.n603 19.3944
R7752 gnd.n5977 gnd.n5976 19.3944
R7753 gnd.n5976 gnd.n5975 19.3944
R7754 gnd.n5975 gnd.n611 19.3944
R7755 gnd.n5969 gnd.n611 19.3944
R7756 gnd.n5969 gnd.n5968 19.3944
R7757 gnd.n5968 gnd.n5967 19.3944
R7758 gnd.n5967 gnd.n619 19.3944
R7759 gnd.n5961 gnd.n619 19.3944
R7760 gnd.n5961 gnd.n5960 19.3944
R7761 gnd.n5960 gnd.n5959 19.3944
R7762 gnd.n5959 gnd.n627 19.3944
R7763 gnd.n5953 gnd.n627 19.3944
R7764 gnd.n5953 gnd.n5952 19.3944
R7765 gnd.n5952 gnd.n5951 19.3944
R7766 gnd.n5951 gnd.n635 19.3944
R7767 gnd.n5945 gnd.n635 19.3944
R7768 gnd.n5945 gnd.n5944 19.3944
R7769 gnd.n5944 gnd.n5943 19.3944
R7770 gnd.n5943 gnd.n643 19.3944
R7771 gnd.n5937 gnd.n643 19.3944
R7772 gnd.n5937 gnd.n5936 19.3944
R7773 gnd.n5936 gnd.n5935 19.3944
R7774 gnd.n5935 gnd.n651 19.3944
R7775 gnd.n5929 gnd.n651 19.3944
R7776 gnd.n5929 gnd.n5928 19.3944
R7777 gnd.n5928 gnd.n5927 19.3944
R7778 gnd.n5927 gnd.n659 19.3944
R7779 gnd.n5921 gnd.n659 19.3944
R7780 gnd.n5921 gnd.n5920 19.3944
R7781 gnd.n5920 gnd.n5919 19.3944
R7782 gnd.n5919 gnd.n667 19.3944
R7783 gnd.n5913 gnd.n667 19.3944
R7784 gnd.n5913 gnd.n5912 19.3944
R7785 gnd.n5912 gnd.n5911 19.3944
R7786 gnd.n5911 gnd.n675 19.3944
R7787 gnd.n5905 gnd.n675 19.3944
R7788 gnd.n5905 gnd.n5904 19.3944
R7789 gnd.n5904 gnd.n5903 19.3944
R7790 gnd.n5903 gnd.n683 19.3944
R7791 gnd.n5897 gnd.n683 19.3944
R7792 gnd.n5897 gnd.n5896 19.3944
R7793 gnd.n5896 gnd.n5895 19.3944
R7794 gnd.n5895 gnd.n691 19.3944
R7795 gnd.n5889 gnd.n691 19.3944
R7796 gnd.n5889 gnd.n5888 19.3944
R7797 gnd.n5888 gnd.n5887 19.3944
R7798 gnd.n5887 gnd.n699 19.3944
R7799 gnd.n5881 gnd.n699 19.3944
R7800 gnd.n5881 gnd.n5880 19.3944
R7801 gnd.n5880 gnd.n5879 19.3944
R7802 gnd.n5879 gnd.n707 19.3944
R7803 gnd.n5873 gnd.n707 19.3944
R7804 gnd.n5873 gnd.n5872 19.3944
R7805 gnd.n5872 gnd.n5871 19.3944
R7806 gnd.n5871 gnd.n715 19.3944
R7807 gnd.n5865 gnd.n715 19.3944
R7808 gnd.n5865 gnd.n5864 19.3944
R7809 gnd.n5864 gnd.n5863 19.3944
R7810 gnd.n5863 gnd.n723 19.3944
R7811 gnd.n5857 gnd.n723 19.3944
R7812 gnd.n5857 gnd.n5856 19.3944
R7813 gnd.n5856 gnd.n5855 19.3944
R7814 gnd.n5855 gnd.n731 19.3944
R7815 gnd.n5849 gnd.n731 19.3944
R7816 gnd.n5849 gnd.n5848 19.3944
R7817 gnd.n5848 gnd.n5847 19.3944
R7818 gnd.n5847 gnd.n739 19.3944
R7819 gnd.n5841 gnd.n739 19.3944
R7820 gnd.n5841 gnd.n5840 19.3944
R7821 gnd.n5840 gnd.n5839 19.3944
R7822 gnd.n5839 gnd.n747 19.3944
R7823 gnd.n5833 gnd.n747 19.3944
R7824 gnd.n5833 gnd.n5832 19.3944
R7825 gnd.n5832 gnd.n5831 19.3944
R7826 gnd.n5831 gnd.n755 19.3944
R7827 gnd.n5825 gnd.n755 19.3944
R7828 gnd.n5825 gnd.n5824 19.3944
R7829 gnd.n5824 gnd.n5823 19.3944
R7830 gnd.n5823 gnd.n763 19.3944
R7831 gnd.n4194 gnd.n4193 19.3944
R7832 gnd.n4193 gnd.n4192 19.3944
R7833 gnd.n4192 gnd.n1091 19.3944
R7834 gnd.n4188 gnd.n1091 19.3944
R7835 gnd.n4188 gnd.n4187 19.3944
R7836 gnd.n4187 gnd.n4186 19.3944
R7837 gnd.n4186 gnd.n1096 19.3944
R7838 gnd.n4182 gnd.n1096 19.3944
R7839 gnd.n4182 gnd.n4181 19.3944
R7840 gnd.n4181 gnd.n4180 19.3944
R7841 gnd.n4180 gnd.n1101 19.3944
R7842 gnd.n4176 gnd.n1101 19.3944
R7843 gnd.n4176 gnd.n4175 19.3944
R7844 gnd.n4175 gnd.n4174 19.3944
R7845 gnd.n4174 gnd.n1106 19.3944
R7846 gnd.n4170 gnd.n1106 19.3944
R7847 gnd.n4170 gnd.n4169 19.3944
R7848 gnd.n4169 gnd.n4168 19.3944
R7849 gnd.n4168 gnd.n1111 19.3944
R7850 gnd.n4164 gnd.n1111 19.3944
R7851 gnd.n4164 gnd.n4163 19.3944
R7852 gnd.n4163 gnd.n4162 19.3944
R7853 gnd.n4162 gnd.n1116 19.3944
R7854 gnd.n4158 gnd.n1116 19.3944
R7855 gnd.n4158 gnd.n4157 19.3944
R7856 gnd.n4157 gnd.n4156 19.3944
R7857 gnd.n4156 gnd.n1121 19.3944
R7858 gnd.n4152 gnd.n1121 19.3944
R7859 gnd.n4152 gnd.n4151 19.3944
R7860 gnd.n4151 gnd.n4150 19.3944
R7861 gnd.n4150 gnd.n1126 19.3944
R7862 gnd.n4146 gnd.n1126 19.3944
R7863 gnd.n4146 gnd.n4145 19.3944
R7864 gnd.n4145 gnd.n4144 19.3944
R7865 gnd.n4144 gnd.n1131 19.3944
R7866 gnd.n4140 gnd.n1131 19.3944
R7867 gnd.n4140 gnd.n4139 19.3944
R7868 gnd.n4139 gnd.n4138 19.3944
R7869 gnd.n4138 gnd.n1136 19.3944
R7870 gnd.n4134 gnd.n1136 19.3944
R7871 gnd.n4134 gnd.n4133 19.3944
R7872 gnd.n4133 gnd.n4132 19.3944
R7873 gnd.n4132 gnd.n1141 19.3944
R7874 gnd.n4128 gnd.n1141 19.3944
R7875 gnd.n4128 gnd.n4127 19.3944
R7876 gnd.n4127 gnd.n4126 19.3944
R7877 gnd.n4126 gnd.n1146 19.3944
R7878 gnd.n4122 gnd.n1146 19.3944
R7879 gnd.n4122 gnd.n4121 19.3944
R7880 gnd.n4121 gnd.n4120 19.3944
R7881 gnd.n4120 gnd.n1151 19.3944
R7882 gnd.n4116 gnd.n1151 19.3944
R7883 gnd.n4116 gnd.n4115 19.3944
R7884 gnd.n4115 gnd.n4114 19.3944
R7885 gnd.n4114 gnd.n1156 19.3944
R7886 gnd.n4110 gnd.n1156 19.3944
R7887 gnd.n4110 gnd.n4109 19.3944
R7888 gnd.n4109 gnd.n4108 19.3944
R7889 gnd.n4108 gnd.n1161 19.3944
R7890 gnd.n4104 gnd.n1161 19.3944
R7891 gnd.n4104 gnd.n4103 19.3944
R7892 gnd.n4103 gnd.n4102 19.3944
R7893 gnd.n4102 gnd.n1166 19.3944
R7894 gnd.n4098 gnd.n1166 19.3944
R7895 gnd.n4098 gnd.n4097 19.3944
R7896 gnd.n4097 gnd.n4096 19.3944
R7897 gnd.n4096 gnd.n1171 19.3944
R7898 gnd.n4092 gnd.n1171 19.3944
R7899 gnd.n4092 gnd.n4091 19.3944
R7900 gnd.n4091 gnd.n4090 19.3944
R7901 gnd.n4090 gnd.n1176 19.3944
R7902 gnd.n4086 gnd.n1176 19.3944
R7903 gnd.n4086 gnd.n4085 19.3944
R7904 gnd.n4085 gnd.n4084 19.3944
R7905 gnd.n4084 gnd.n1181 19.3944
R7906 gnd.n4080 gnd.n1181 19.3944
R7907 gnd.n4080 gnd.n4079 19.3944
R7908 gnd.n4079 gnd.n4078 19.3944
R7909 gnd.n4078 gnd.n1186 19.3944
R7910 gnd.n4074 gnd.n1186 19.3944
R7911 gnd.n4074 gnd.n4073 19.3944
R7912 gnd.n4073 gnd.n4072 19.3944
R7913 gnd.n3481 gnd.n3316 19.3944
R7914 gnd.n3481 gnd.n3314 19.3944
R7915 gnd.n3486 gnd.n3314 19.3944
R7916 gnd.n3380 gnd.n3362 19.3944
R7917 gnd.n3380 gnd.n3360 19.3944
R7918 gnd.n3386 gnd.n3360 19.3944
R7919 gnd.n3386 gnd.n3353 19.3944
R7920 gnd.n3399 gnd.n3353 19.3944
R7921 gnd.n3399 gnd.n3351 19.3944
R7922 gnd.n3405 gnd.n3351 19.3944
R7923 gnd.n3405 gnd.n3344 19.3944
R7924 gnd.n3418 gnd.n3344 19.3944
R7925 gnd.n3418 gnd.n3342 19.3944
R7926 gnd.n3424 gnd.n3342 19.3944
R7927 gnd.n3424 gnd.n3335 19.3944
R7928 gnd.n3437 gnd.n3335 19.3944
R7929 gnd.n3437 gnd.n3333 19.3944
R7930 gnd.n3445 gnd.n3333 19.3944
R7931 gnd.n3445 gnd.n3444 19.3944
R7932 gnd.n3444 gnd.n3324 19.3944
R7933 gnd.n3458 gnd.n3324 19.3944
R7934 gnd.n3458 gnd.n3322 19.3944
R7935 gnd.n3464 gnd.n3322 19.3944
R7936 gnd.n3464 gnd.n3320 19.3944
R7937 gnd.n3468 gnd.n3320 19.3944
R7938 gnd.n3468 gnd.n3318 19.3944
R7939 gnd.n3477 gnd.n3318 19.3944
R7940 gnd.t224 gnd.n4634 18.8012
R7941 gnd.n5226 gnd.t30 18.8012
R7942 gnd.n5071 gnd.n5070 18.4825
R7943 gnd.n3756 gnd.n1360 18.4247
R7944 gnd.n2597 gnd.n2596 18.4247
R7945 gnd.n6682 gnd.n6681 18.2308
R7946 gnd.n3448 gnd.n3328 18.2308
R7947 gnd.n2635 gnd.n1909 18.2308
R7948 gnd.n2116 gnd.n2108 18.2308
R7949 gnd.t52 gnd.n4678 18.1639
R7950 gnd.n5820 gnd.n5819 17.8452
R7951 gnd.n2759 gnd.n2757 17.6395
R7952 gnd.n3626 gnd.n3625 17.6395
R7953 gnd.n4705 gnd.t49 17.5266
R7954 gnd.n4663 gnd.t76 16.8893
R7955 gnd.n2165 gnd.t171 16.8893
R7956 gnd.n2418 gnd.t117 16.8893
R7957 gnd.n3814 gnd.t113 16.8893
R7958 gnd.t95 gnd.n81 16.8893
R7959 gnd.n4932 gnd.t198 16.2519
R7960 gnd.n5216 gnd.t15 16.2519
R7961 gnd.n2468 gnd.n2467 16.0975
R7962 gnd.n1399 gnd.n1398 16.0975
R7963 gnd.n2532 gnd.n2531 16.0975
R7964 gnd.n3562 gnd.n3561 16.0975
R7965 gnd.n2675 gnd.n1849 15.9333
R7966 gnd.n2675 gnd.n1862 15.9333
R7967 gnd.n2333 gnd.n2332 15.9333
R7968 gnd.n2332 gnd.n1843 15.9333
R7969 gnd.n2684 gnd.n1843 15.9333
R7970 gnd.n2686 gnd.n2684 15.9333
R7971 gnd.n2685 gnd.n1836 15.9333
R7972 gnd.n2696 gnd.n1836 15.9333
R7973 gnd.n2696 gnd.n2694 15.9333
R7974 gnd.n2694 gnd.n1837 15.9333
R7975 gnd.n1837 gnd.n1830 15.9333
R7976 gnd.n2704 gnd.n1830 15.9333
R7977 gnd.n2706 gnd.n2704 15.9333
R7978 gnd.n2706 gnd.n2705 15.9333
R7979 gnd.n2716 gnd.n1823 15.9333
R7980 gnd.n2716 gnd.n2714 15.9333
R7981 gnd.n2714 gnd.n1824 15.9333
R7982 gnd.n1824 gnd.n1817 15.9333
R7983 gnd.n2724 gnd.n1817 15.9333
R7984 gnd.n2727 gnd.n2724 15.9333
R7985 gnd.n2727 gnd.n2726 15.9333
R7986 gnd.n2726 gnd.n2725 15.9333
R7987 gnd.n2739 gnd.n2737 15.9333
R7988 gnd.n2737 gnd.n1810 15.9333
R7989 gnd.n1810 gnd.n1770 15.9333
R7990 gnd.n2751 gnd.n2750 15.9333
R7991 gnd.n2804 gnd.n2803 15.9333
R7992 gnd.n2815 gnd.n2814 15.9333
R7993 gnd.n2790 gnd.n1718 15.9333
R7994 gnd.n2868 gnd.n2867 15.9333
R7995 gnd.n2901 gnd.n2900 15.9333
R7996 gnd.n1661 gnd.n1650 15.9333
R7997 gnd.n2948 gnd.n1641 15.9333
R7998 gnd.n2921 gnd.n1633 15.9333
R7999 gnd.n2993 gnd.n1624 15.9333
R8000 gnd.n2963 gnd.n1594 15.9333
R8001 gnd.n3044 gnd.n1594 15.9333
R8002 gnd.n3054 gnd.n1572 15.9333
R8003 gnd.n3126 gnd.n3125 15.9333
R8004 gnd.n3134 gnd.n1547 15.9333
R8005 gnd.n3187 gnd.n1536 15.9333
R8006 gnd.n3196 gnd.n3195 15.9333
R8007 gnd.n3226 gnd.n3225 15.9333
R8008 gnd.n3273 gnd.n1479 15.9333
R8009 gnd.n3289 gnd.n1465 15.9333
R8010 gnd.n3537 gnd.n3535 15.9333
R8011 gnd.n1403 gnd.n1365 15.9333
R8012 gnd.n3529 gnd.n3528 15.9333
R8013 gnd.n3528 gnd.n3527 15.9333
R8014 gnd.n3527 gnd.n3526 15.9333
R8015 gnd.n3524 gnd.n1422 15.9333
R8016 gnd.n1430 gnd.n1422 15.9333
R8017 gnd.n1431 gnd.n1430 15.9333
R8018 gnd.n3518 gnd.n1431 15.9333
R8019 gnd.n3518 gnd.n3517 15.9333
R8020 gnd.n3517 gnd.n3516 15.9333
R8021 gnd.n3516 gnd.n3515 15.9333
R8022 gnd.n3515 gnd.n3513 15.9333
R8023 gnd.n1451 gnd.n1450 15.9333
R8024 gnd.n1450 gnd.n1441 15.9333
R8025 gnd.n3507 gnd.n1441 15.9333
R8026 gnd.n3507 gnd.n3506 15.9333
R8027 gnd.n3506 gnd.n3505 15.9333
R8028 gnd.n3505 gnd.n3504 15.9333
R8029 gnd.n3504 gnd.n3502 15.9333
R8030 gnd.n3502 gnd.n1444 15.9333
R8031 gnd.n3493 gnd.n3492 15.9333
R8032 gnd.n3492 gnd.n1192 15.9333
R8033 gnd.n4070 gnd.n1192 15.9333
R8034 gnd.n4070 gnd.n4069 15.9333
R8035 gnd.n1203 gnd.n1194 15.9333
R8036 gnd.n4063 gnd.n1203 15.9333
R8037 gnd.n5626 gnd.n5624 15.6674
R8038 gnd.n5594 gnd.n5592 15.6674
R8039 gnd.n5562 gnd.n5560 15.6674
R8040 gnd.n5531 gnd.n5529 15.6674
R8041 gnd.n5499 gnd.n5497 15.6674
R8042 gnd.n5467 gnd.n5465 15.6674
R8043 gnd.n5435 gnd.n5433 15.6674
R8044 gnd.n5404 gnd.n5402 15.6674
R8045 gnd.n4923 gnd.t198 15.6146
R8046 gnd.t106 gnd.n5805 15.6146
R8047 gnd.n5709 gnd.t130 15.6146
R8048 gnd.t164 gnd.n2685 15.6146
R8049 gnd.t134 gnd.n1444 15.6146
R8050 gnd.n1745 gnd.n1740 15.296
R8051 gnd.n2859 gnd.t6 15.296
R8052 gnd.n2939 gnd.n2937 15.296
R8053 gnd.n2958 gnd.n2957 15.296
R8054 gnd.n3116 gnd.n1553 15.296
R8055 gnd.n3135 gnd.n1543 15.296
R8056 gnd.n3148 gnd.t236 15.296
R8057 gnd.n3546 gnd.n3545 15.0827
R8058 gnd.n1756 gnd.n1751 15.0481
R8059 gnd.n3556 gnd.n3555 15.0481
R8060 gnd.n5354 gnd.t48 14.9773
R8061 gnd.t171 gnd.n884 14.9773
R8062 gnd.n2725 gnd.t282 14.9773
R8063 gnd.t237 gnd.n3524 14.9773
R8064 gnd.n1733 gnd.t142 14.6587
R8065 gnd.n2849 gnd.n1697 14.6587
R8066 gnd.n2887 gnd.n1677 14.6587
R8067 gnd.n3207 gnd.n3206 14.6587
R8068 gnd.n3149 gnd.n1493 14.6587
R8069 gnd.n1471 gnd.t138 14.6587
R8070 gnd.t288 gnd.n4507 14.34
R8071 gnd.t51 gnd.n767 14.34
R8072 gnd.n3274 gnd.n1476 14.0214
R8073 gnd.n5036 gnd.t251 13.7027
R8074 gnd.n4789 gnd.n4788 13.5763
R8075 gnd.n5765 gnd.n4439 13.5763
R8076 gnd.n1340 gnd.n1339 13.5763
R8077 gnd.n6734 gnd.n6733 13.5763
R8078 gnd.n4333 gnd.n876 13.5763
R8079 gnd.n2428 gnd.n2425 13.5763
R8080 gnd.n5071 gnd.n4735 13.384
R8081 gnd.n2841 gnd.n2840 13.384
R8082 gnd.n2910 gnd.n1657 13.384
R8083 gnd.n2974 gnd.n1616 13.384
R8084 gnd.n3002 gnd.t241 13.384
R8085 gnd.n3036 gnd.t32 13.384
R8086 gnd.n3072 gnd.t60 13.384
R8087 gnd.t234 gnd.n1576 13.384
R8088 gnd.n3091 gnd.n3090 13.384
R8089 gnd.n3168 gnd.n1530 13.384
R8090 gnd.n3257 gnd.n1489 13.384
R8091 gnd.n1767 gnd.n1748 13.1884
R8092 gnd.n1762 gnd.n1761 13.1884
R8093 gnd.n1761 gnd.n1760 13.1884
R8094 gnd.n3549 gnd.n3544 13.1884
R8095 gnd.n3550 gnd.n3549 13.1884
R8096 gnd.n1763 gnd.n1750 13.146
R8097 gnd.n1759 gnd.n1750 13.146
R8098 gnd.n3548 gnd.n3547 13.146
R8099 gnd.n3548 gnd.n3543 13.146
R8100 gnd.n5627 gnd.n5623 12.8005
R8101 gnd.n5595 gnd.n5591 12.8005
R8102 gnd.n5563 gnd.n5559 12.8005
R8103 gnd.n5532 gnd.n5528 12.8005
R8104 gnd.n5500 gnd.n5496 12.8005
R8105 gnd.n5468 gnd.n5464 12.8005
R8106 gnd.n5436 gnd.n5432 12.8005
R8107 gnd.n5405 gnd.n5401 12.8005
R8108 gnd.n2902 gnd.n1667 12.7467
R8109 gnd.n1617 gnd.n1606 12.7467
R8110 gnd.n3063 gnd.n1585 12.7467
R8111 gnd.n3164 gnd.n1520 12.7467
R8112 gnd.n4788 gnd.n4783 12.4126
R8113 gnd.n5770 gnd.n4439 12.4126
R8114 gnd.n3808 gnd.n1339 12.4126
R8115 gnd.n6733 gnd.n155 12.4126
R8116 gnd.n4329 gnd.n876 12.4126
R8117 gnd.n2425 gnd.n1995 12.4126
R8118 gnd.n2757 gnd.n2756 12.1761
R8119 gnd.n3625 gnd.n3624 12.1761
R8120 gnd.n2791 gnd.n1728 12.1094
R8121 gnd.n2930 gnd.n2929 12.1094
R8122 gnd.n2982 gnd.n2981 12.1094
R8123 gnd.n3055 gnd.n1562 12.1094
R8124 gnd.n3176 gnd.n3175 12.1094
R8125 gnd.n1478 gnd.t189 12.1094
R8126 gnd.n5631 gnd.n5630 12.0247
R8127 gnd.n5599 gnd.n5598 12.0247
R8128 gnd.n5567 gnd.n5566 12.0247
R8129 gnd.n5536 gnd.n5535 12.0247
R8130 gnd.n5504 gnd.n5503 12.0247
R8131 gnd.n5472 gnd.n5471 12.0247
R8132 gnd.n5440 gnd.n5439 12.0247
R8133 gnd.n5409 gnd.n5408 12.0247
R8134 gnd.t24 gnd.n898 11.7908
R8135 gnd.n4219 gnd.t222 11.7908
R8136 gnd.n3944 gnd.t87 11.7908
R8137 gnd.n6635 gnd.t11 11.7908
R8138 gnd.n2625 gnd.n1934 11.4721
R8139 gnd.t152 gnd.n2833 11.4721
R8140 gnd.n2857 gnd.n1700 11.4721
R8141 gnd.t77 gnd.n1681 11.4721
R8142 gnd.n2880 gnd.n2879 11.4721
R8143 gnd.n3035 gnd.n1601 11.4721
R8144 gnd.n3073 gnd.n1589 11.4721
R8145 gnd.n3214 gnd.n1515 11.4721
R8146 gnd.n3156 gnd.t233 11.4721
R8147 gnd.n3234 gnd.n3232 11.4721
R8148 gnd.n4061 gnd.n1204 11.4721
R8149 gnd.n5634 gnd.n5621 11.249
R8150 gnd.n5602 gnd.n5589 11.249
R8151 gnd.n5570 gnd.n5557 11.249
R8152 gnd.n5539 gnd.n5526 11.249
R8153 gnd.n5507 gnd.n5494 11.249
R8154 gnd.n5475 gnd.n5462 11.249
R8155 gnd.n5443 gnd.n5430 11.249
R8156 gnd.n5412 gnd.n5399 11.249
R8157 gnd.n5144 gnd.t251 11.1535
R8158 gnd.t56 gnd.n939 11.1535
R8159 gnd.n4243 gnd.t27 11.1535
R8160 gnd.n2705 gnd.t201 11.1535
R8161 gnd.n1451 gnd.t228 11.1535
R8162 gnd.n4004 gnd.t64 11.1535
R8163 gnd.n6603 gnd.t83 11.1535
R8164 gnd.n2045 gnd.n960 10.8348
R8165 gnd.n4269 gnd.n973 10.8348
R8166 gnd.n2244 gnd.n978 10.8348
R8167 gnd.n2253 gnd.n987 10.8348
R8168 gnd.n4256 gnd.n990 10.8348
R8169 gnd.n2261 gnd.n995 10.8348
R8170 gnd.n4249 gnd.n998 10.8348
R8171 gnd.n2301 gnd.n2300 10.8348
R8172 gnd.n4243 gnd.n1008 10.8348
R8173 gnd.n2269 gnd.n1016 10.8348
R8174 gnd.n2274 gnd.n1026 10.8348
R8175 gnd.n4231 gnd.n1029 10.8348
R8176 gnd.n2286 gnd.n1037 10.8348
R8177 gnd.n4225 gnd.n1040 10.8348
R8178 gnd.n2361 gnd.n2360 10.8348
R8179 gnd.n4219 gnd.n1050 10.8348
R8180 gnd.n2369 gnd.n1058 10.8348
R8181 gnd.n4213 gnd.n1061 10.8348
R8182 gnd.n2378 gnd.n1069 10.8348
R8183 gnd.n4207 gnd.n1072 10.8348
R8184 gnd.n2418 gnd.n1079 10.8348
R8185 gnd.n4201 gnd.n1082 10.8348
R8186 gnd.n2923 gnd.n2922 10.8348
R8187 gnd.n3124 gnd.n1556 10.8348
R8188 gnd.n3538 gnd.n1408 10.8348
R8189 gnd.n4055 gnd.n4054 10.8348
R8190 gnd.n3814 gnd.n1215 10.8348
R8191 gnd.n4048 gnd.n1224 10.8348
R8192 gnd.n3823 gnd.n1227 10.8348
R8193 gnd.n3934 gnd.n1325 10.8348
R8194 gnd.n3933 gnd.n3916 10.8348
R8195 gnd.n3944 gnd.n1318 10.8348
R8196 gnd.n1320 gnd.n1310 10.8348
R8197 gnd.n3954 gnd.n3953 10.8348
R8198 gnd.n3965 gnd.n1299 10.8348
R8199 gnd.n3964 gnd.n1302 10.8348
R8200 gnd.n3976 gnd.n1289 10.8348
R8201 gnd.n3986 gnd.n3985 10.8348
R8202 gnd.n4004 gnd.n1270 10.8348
R8203 gnd.n4003 gnd.n1274 10.8348
R8204 gnd.n4010 gnd.n1260 10.8348
R8205 gnd.n3896 gnd.n1262 10.8348
R8206 gnd.n4019 gnd.n1251 10.8348
R8207 gnd.n6568 gnd.n248 10.8348
R8208 gnd.n3890 gnd.n246 10.8348
R8209 gnd.n6581 gnd.n236 10.8348
R8210 gnd.n6560 gnd.n230 10.8348
R8211 gnd.n3690 gnd.n1361 10.6151
R8212 gnd.n3690 gnd.n3689 10.6151
R8213 gnd.n3687 gnd.n3684 10.6151
R8214 gnd.n3684 gnd.n3683 10.6151
R8215 gnd.n3683 gnd.n3680 10.6151
R8216 gnd.n3680 gnd.n3679 10.6151
R8217 gnd.n3679 gnd.n3676 10.6151
R8218 gnd.n3676 gnd.n3675 10.6151
R8219 gnd.n3675 gnd.n3672 10.6151
R8220 gnd.n3672 gnd.n3671 10.6151
R8221 gnd.n3671 gnd.n3668 10.6151
R8222 gnd.n3668 gnd.n3667 10.6151
R8223 gnd.n3667 gnd.n3664 10.6151
R8224 gnd.n3664 gnd.n3663 10.6151
R8225 gnd.n3663 gnd.n3660 10.6151
R8226 gnd.n3660 gnd.n3659 10.6151
R8227 gnd.n3659 gnd.n3656 10.6151
R8228 gnd.n3656 gnd.n3655 10.6151
R8229 gnd.n3655 gnd.n3652 10.6151
R8230 gnd.n3652 gnd.n3651 10.6151
R8231 gnd.n3651 gnd.n3648 10.6151
R8232 gnd.n3648 gnd.n3647 10.6151
R8233 gnd.n3647 gnd.n3644 10.6151
R8234 gnd.n3644 gnd.n3643 10.6151
R8235 gnd.n3643 gnd.n3640 10.6151
R8236 gnd.n3640 gnd.n3639 10.6151
R8237 gnd.n3639 gnd.n3636 10.6151
R8238 gnd.n3636 gnd.n3635 10.6151
R8239 gnd.n3635 gnd.n3632 10.6151
R8240 gnd.n3632 gnd.n3631 10.6151
R8241 gnd.n2764 gnd.n2763 10.6151
R8242 gnd.n2798 gnd.n2764 10.6151
R8243 gnd.n2798 gnd.n2797 10.6151
R8244 gnd.n2797 gnd.n2796 10.6151
R8245 gnd.n2796 gnd.n2794 10.6151
R8246 gnd.n2794 gnd.n2793 10.6151
R8247 gnd.n2793 gnd.n2789 10.6151
R8248 gnd.n2789 gnd.n2788 10.6151
R8249 gnd.n2788 gnd.n2786 10.6151
R8250 gnd.n2786 gnd.n2785 10.6151
R8251 gnd.n2785 gnd.n2781 10.6151
R8252 gnd.n2781 gnd.n2780 10.6151
R8253 gnd.n2780 gnd.n2778 10.6151
R8254 gnd.n2778 gnd.n2777 10.6151
R8255 gnd.n2777 gnd.n2775 10.6151
R8256 gnd.n2775 gnd.n2774 10.6151
R8257 gnd.n2774 gnd.n2773 10.6151
R8258 gnd.n2773 gnd.n2772 10.6151
R8259 gnd.n2772 gnd.n2771 10.6151
R8260 gnd.n2771 gnd.n2768 10.6151
R8261 gnd.n2768 gnd.n2767 10.6151
R8262 gnd.n2767 gnd.n2765 10.6151
R8263 gnd.n2765 gnd.n1648 10.6151
R8264 gnd.n2932 gnd.n1648 10.6151
R8265 gnd.n2933 gnd.n2932 10.6151
R8266 gnd.n2935 gnd.n2933 10.6151
R8267 gnd.n2935 gnd.n2934 10.6151
R8268 gnd.n2934 gnd.n1631 10.6151
R8269 gnd.n2960 gnd.n1631 10.6151
R8270 gnd.n2961 gnd.n2960 10.6151
R8271 gnd.n2979 gnd.n2961 10.6151
R8272 gnd.n2979 gnd.n2978 10.6151
R8273 gnd.n2978 gnd.n2977 10.6151
R8274 gnd.n2977 gnd.n2962 10.6151
R8275 gnd.n2970 gnd.n2962 10.6151
R8276 gnd.n2970 gnd.n2969 10.6151
R8277 gnd.n2969 gnd.n2968 10.6151
R8278 gnd.n2968 gnd.n2967 10.6151
R8279 gnd.n2967 gnd.n2966 10.6151
R8280 gnd.n2966 gnd.n1592 10.6151
R8281 gnd.n3047 gnd.n1592 10.6151
R8282 gnd.n3048 gnd.n3047 10.6151
R8283 gnd.n3067 gnd.n3048 10.6151
R8284 gnd.n3067 gnd.n3066 10.6151
R8285 gnd.n3066 gnd.n3065 10.6151
R8286 gnd.n3065 gnd.n3061 10.6151
R8287 gnd.n3061 gnd.n3060 10.6151
R8288 gnd.n3060 gnd.n3058 10.6151
R8289 gnd.n3058 gnd.n3057 10.6151
R8290 gnd.n3057 gnd.n3052 10.6151
R8291 gnd.n3052 gnd.n3051 10.6151
R8292 gnd.n3051 gnd.n3049 10.6151
R8293 gnd.n3049 gnd.n1545 10.6151
R8294 gnd.n3137 gnd.n1545 10.6151
R8295 gnd.n3138 gnd.n3137 10.6151
R8296 gnd.n3173 gnd.n3138 10.6151
R8297 gnd.n3173 gnd.n3172 10.6151
R8298 gnd.n3172 gnd.n3171 10.6151
R8299 gnd.n3171 gnd.n3139 10.6151
R8300 gnd.n3163 gnd.n3139 10.6151
R8301 gnd.n3163 gnd.n3162 10.6151
R8302 gnd.n3162 gnd.n3161 10.6151
R8303 gnd.n3161 gnd.n3160 10.6151
R8304 gnd.n3160 gnd.n3159 10.6151
R8305 gnd.n3159 gnd.n3155 10.6151
R8306 gnd.n3155 gnd.n3154 10.6151
R8307 gnd.n3154 gnd.n3152 10.6151
R8308 gnd.n3152 gnd.n3151 10.6151
R8309 gnd.n3151 gnd.n3147 10.6151
R8310 gnd.n3147 gnd.n3146 10.6151
R8311 gnd.n3146 gnd.n3144 10.6151
R8312 gnd.n3144 gnd.n3143 10.6151
R8313 gnd.n3143 gnd.n3140 10.6151
R8314 gnd.n3140 gnd.n1467 10.6151
R8315 gnd.n3283 gnd.n1467 10.6151
R8316 gnd.n3284 gnd.n3283 10.6151
R8317 gnd.n3287 gnd.n3284 10.6151
R8318 gnd.n3287 gnd.n3286 10.6151
R8319 gnd.n3286 gnd.n3285 10.6151
R8320 gnd.n3285 gnd.n1400 10.6151
R8321 gnd.n2530 gnd.n2529 10.6151
R8322 gnd.n2529 gnd.n2526 10.6151
R8323 gnd.n2524 gnd.n2521 10.6151
R8324 gnd.n2521 gnd.n2520 10.6151
R8325 gnd.n2520 gnd.n2517 10.6151
R8326 gnd.n2517 gnd.n2516 10.6151
R8327 gnd.n2516 gnd.n2513 10.6151
R8328 gnd.n2513 gnd.n2512 10.6151
R8329 gnd.n2512 gnd.n2509 10.6151
R8330 gnd.n2509 gnd.n2508 10.6151
R8331 gnd.n2508 gnd.n2505 10.6151
R8332 gnd.n2505 gnd.n2504 10.6151
R8333 gnd.n2504 gnd.n2501 10.6151
R8334 gnd.n2501 gnd.n2500 10.6151
R8335 gnd.n2500 gnd.n2497 10.6151
R8336 gnd.n2497 gnd.n2496 10.6151
R8337 gnd.n2496 gnd.n2493 10.6151
R8338 gnd.n2493 gnd.n2492 10.6151
R8339 gnd.n2492 gnd.n2489 10.6151
R8340 gnd.n2489 gnd.n2488 10.6151
R8341 gnd.n2488 gnd.n2485 10.6151
R8342 gnd.n2485 gnd.n2484 10.6151
R8343 gnd.n2484 gnd.n2481 10.6151
R8344 gnd.n2481 gnd.n2480 10.6151
R8345 gnd.n2480 gnd.n2477 10.6151
R8346 gnd.n2477 gnd.n2476 10.6151
R8347 gnd.n2476 gnd.n2473 10.6151
R8348 gnd.n2473 gnd.n2472 10.6151
R8349 gnd.n2472 gnd.n2469 10.6151
R8350 gnd.n2469 gnd.n1743 10.6151
R8351 gnd.n2756 gnd.n2755 10.6151
R8352 gnd.n2755 gnd.n1768 10.6151
R8353 gnd.n2535 gnd.n1768 10.6151
R8354 gnd.n2536 gnd.n2535 10.6151
R8355 gnd.n2539 gnd.n2536 10.6151
R8356 gnd.n2540 gnd.n2539 10.6151
R8357 gnd.n2543 gnd.n2540 10.6151
R8358 gnd.n2544 gnd.n2543 10.6151
R8359 gnd.n2547 gnd.n2544 10.6151
R8360 gnd.n2548 gnd.n2547 10.6151
R8361 gnd.n2551 gnd.n2548 10.6151
R8362 gnd.n2552 gnd.n2551 10.6151
R8363 gnd.n2555 gnd.n2552 10.6151
R8364 gnd.n2556 gnd.n2555 10.6151
R8365 gnd.n2559 gnd.n2556 10.6151
R8366 gnd.n2560 gnd.n2559 10.6151
R8367 gnd.n2563 gnd.n2560 10.6151
R8368 gnd.n2564 gnd.n2563 10.6151
R8369 gnd.n2567 gnd.n2564 10.6151
R8370 gnd.n2568 gnd.n2567 10.6151
R8371 gnd.n2571 gnd.n2568 10.6151
R8372 gnd.n2572 gnd.n2571 10.6151
R8373 gnd.n2575 gnd.n2572 10.6151
R8374 gnd.n2576 gnd.n2575 10.6151
R8375 gnd.n2579 gnd.n2576 10.6151
R8376 gnd.n2580 gnd.n2579 10.6151
R8377 gnd.n2583 gnd.n2580 10.6151
R8378 gnd.n2584 gnd.n2583 10.6151
R8379 gnd.n2588 gnd.n2587 10.6151
R8380 gnd.n2591 gnd.n2588 10.6151
R8381 gnd.n3624 gnd.n3623 10.6151
R8382 gnd.n3623 gnd.n3620 10.6151
R8383 gnd.n3620 gnd.n3619 10.6151
R8384 gnd.n3619 gnd.n3616 10.6151
R8385 gnd.n3616 gnd.n3615 10.6151
R8386 gnd.n3615 gnd.n3612 10.6151
R8387 gnd.n3612 gnd.n3611 10.6151
R8388 gnd.n3611 gnd.n3608 10.6151
R8389 gnd.n3608 gnd.n3607 10.6151
R8390 gnd.n3607 gnd.n3604 10.6151
R8391 gnd.n3604 gnd.n3603 10.6151
R8392 gnd.n3603 gnd.n3600 10.6151
R8393 gnd.n3600 gnd.n3599 10.6151
R8394 gnd.n3599 gnd.n3596 10.6151
R8395 gnd.n3596 gnd.n3595 10.6151
R8396 gnd.n3595 gnd.n3592 10.6151
R8397 gnd.n3592 gnd.n3591 10.6151
R8398 gnd.n3591 gnd.n3588 10.6151
R8399 gnd.n3588 gnd.n3587 10.6151
R8400 gnd.n3587 gnd.n3584 10.6151
R8401 gnd.n3584 gnd.n3583 10.6151
R8402 gnd.n3583 gnd.n3580 10.6151
R8403 gnd.n3580 gnd.n3579 10.6151
R8404 gnd.n3579 gnd.n3576 10.6151
R8405 gnd.n3576 gnd.n3575 10.6151
R8406 gnd.n3575 gnd.n3572 10.6151
R8407 gnd.n3572 gnd.n3571 10.6151
R8408 gnd.n3571 gnd.n3568 10.6151
R8409 gnd.n3566 gnd.n3563 10.6151
R8410 gnd.n3563 gnd.n1362 10.6151
R8411 gnd.n2759 gnd.n2758 10.6151
R8412 gnd.n2758 gnd.n1730 10.6151
R8413 gnd.n2818 gnd.n1730 10.6151
R8414 gnd.n2819 gnd.n2818 10.6151
R8415 gnd.n2820 gnd.n2819 10.6151
R8416 gnd.n2820 gnd.n1716 10.6151
R8417 gnd.n2836 gnd.n1716 10.6151
R8418 gnd.n2837 gnd.n2836 10.6151
R8419 gnd.n2838 gnd.n2837 10.6151
R8420 gnd.n2838 gnd.n1703 10.6151
R8421 gnd.n2852 gnd.n1703 10.6151
R8422 gnd.n2853 gnd.n2852 10.6151
R8423 gnd.n2855 gnd.n2853 10.6151
R8424 gnd.n2855 gnd.n2854 10.6151
R8425 gnd.n2854 gnd.n1679 10.6151
R8426 gnd.n2883 gnd.n1679 10.6151
R8427 gnd.n2884 gnd.n2883 10.6151
R8428 gnd.n2885 gnd.n2884 10.6151
R8429 gnd.n2885 gnd.n1664 10.6151
R8430 gnd.n2904 gnd.n1664 10.6151
R8431 gnd.n2905 gnd.n2904 10.6151
R8432 gnd.n2907 gnd.n2905 10.6151
R8433 gnd.n2907 gnd.n2906 10.6151
R8434 gnd.n2906 gnd.n1645 10.6151
R8435 gnd.n2942 gnd.n1645 10.6151
R8436 gnd.n2943 gnd.n2942 10.6151
R8437 gnd.n2945 gnd.n2943 10.6151
R8438 gnd.n2945 gnd.n2944 10.6151
R8439 gnd.n2944 gnd.n1628 10.6151
R8440 gnd.n2985 gnd.n1628 10.6151
R8441 gnd.n2986 gnd.n2985 10.6151
R8442 gnd.n2990 gnd.n2986 10.6151
R8443 gnd.n2990 gnd.n2989 10.6151
R8444 gnd.n2989 gnd.n2988 10.6151
R8445 gnd.n2988 gnd.n1604 10.6151
R8446 gnd.n3028 gnd.n1604 10.6151
R8447 gnd.n3029 gnd.n3028 10.6151
R8448 gnd.n3033 gnd.n3029 10.6151
R8449 gnd.n3033 gnd.n3032 10.6151
R8450 gnd.n3032 gnd.n3031 10.6151
R8451 gnd.n3031 gnd.n1587 10.6151
R8452 gnd.n3075 gnd.n1587 10.6151
R8453 gnd.n3076 gnd.n3075 10.6151
R8454 gnd.n3077 gnd.n3076 10.6151
R8455 gnd.n3077 gnd.n1574 10.6151
R8456 gnd.n3093 gnd.n1574 10.6151
R8457 gnd.n3094 gnd.n3093 10.6151
R8458 gnd.n3095 gnd.n3094 10.6151
R8459 gnd.n3095 gnd.n1560 10.6151
R8460 gnd.n3119 gnd.n1560 10.6151
R8461 gnd.n3120 gnd.n3119 10.6151
R8462 gnd.n3122 gnd.n3120 10.6151
R8463 gnd.n3122 gnd.n3121 10.6151
R8464 gnd.n3121 gnd.n1540 10.6151
R8465 gnd.n3179 gnd.n1540 10.6151
R8466 gnd.n3180 gnd.n3179 10.6151
R8467 gnd.n3184 gnd.n3180 10.6151
R8468 gnd.n3184 gnd.n3183 10.6151
R8469 gnd.n3183 gnd.n3182 10.6151
R8470 gnd.n3182 gnd.n1517 10.6151
R8471 gnd.n3210 gnd.n1517 10.6151
R8472 gnd.n3211 gnd.n3210 10.6151
R8473 gnd.n3212 gnd.n3211 10.6151
R8474 gnd.n3212 gnd.n1505 10.6151
R8475 gnd.n3228 gnd.n1505 10.6151
R8476 gnd.n3229 gnd.n3228 10.6151
R8477 gnd.n3230 gnd.n3229 10.6151
R8478 gnd.n3230 gnd.n1491 10.6151
R8479 gnd.n3253 gnd.n1491 10.6151
R8480 gnd.n3254 gnd.n3253 10.6151
R8481 gnd.n3255 gnd.n3254 10.6151
R8482 gnd.n3255 gnd.n1473 10.6151
R8483 gnd.n3276 gnd.n1473 10.6151
R8484 gnd.n3277 gnd.n3276 10.6151
R8485 gnd.n3279 gnd.n3277 10.6151
R8486 gnd.n3279 gnd.n3278 10.6151
R8487 gnd.n3278 gnd.n1406 10.6151
R8488 gnd.n3540 gnd.n1406 10.6151
R8489 gnd.n3541 gnd.n3540 10.6151
R8490 gnd.n3626 gnd.n3541 10.6151
R8491 gnd.n5060 gnd.t262 10.5161
R8492 gnd.n4509 gnd.t288 10.5161
R8493 gnd.n5698 gnd.t51 10.5161
R8494 gnd.n4275 gnd.n957 10.5161
R8495 gnd.n2045 gnd.t66 10.5161
R8496 gnd.n4269 gnd.t66 10.5161
R8497 gnd.n4262 gnd.t0 10.5161
R8498 gnd.n2752 gnd.n2751 10.5161
R8499 gnd.n3695 gnd.n1365 10.5161
R8500 gnd.n6573 gnd.t16 10.5161
R8501 gnd.n6581 gnd.t61 10.5161
R8502 gnd.n6560 gnd.t61 10.5161
R8503 gnd.n6587 gnd.n232 10.5161
R8504 gnd.n5635 gnd.n5619 10.4732
R8505 gnd.n5603 gnd.n5587 10.4732
R8506 gnd.n5571 gnd.n5555 10.4732
R8507 gnd.n5540 gnd.n5524 10.4732
R8508 gnd.n5508 gnd.n5492 10.4732
R8509 gnd.n5476 gnd.n5460 10.4732
R8510 gnd.n5444 gnd.n5428 10.4732
R8511 gnd.n5413 gnd.n5397 10.4732
R8512 gnd.n1700 gnd.n1690 10.1975
R8513 gnd.n1662 gnd.t93 10.1975
R8514 gnd.n2964 gnd.n1601 10.1975
R8515 gnd.n3045 gnd.n1589 10.1975
R8516 gnd.n3186 gnd.t220 10.1975
R8517 gnd.n3234 gnd.n1501 10.1975
R8518 gnd.n5367 gnd.t48 9.87883
R8519 gnd.n936 gnd.t38 9.87883
R8520 gnd.n2301 gnd.t27 9.87883
R8521 gnd.n4237 gnd.t4 9.87883
R8522 gnd.t46 gnd.n1281 9.87883
R8523 gnd.t64 gnd.n4003 9.87883
R8524 gnd.n6611 gnd.t73 9.87883
R8525 gnd.n5639 gnd.n5638 9.69747
R8526 gnd.n5607 gnd.n5606 9.69747
R8527 gnd.n5575 gnd.n5574 9.69747
R8528 gnd.n5544 gnd.n5543 9.69747
R8529 gnd.n5512 gnd.n5511 9.69747
R8530 gnd.n5480 gnd.n5479 9.69747
R8531 gnd.n5448 gnd.n5447 9.69747
R8532 gnd.n5417 gnd.n5416 9.69747
R8533 gnd.n6840 gnd.n50 9.6512
R8534 gnd.n2822 gnd.n1728 9.56018
R8535 gnd.n2878 gnd.t242 9.56018
R8536 gnd.n2983 gnd.n2982 9.56018
R8537 gnd.n3117 gnd.n1562 9.56018
R8538 gnd.n3215 gnd.t219 9.56018
R8539 gnd.n3281 gnd.t189 9.56018
R8540 gnd.n1411 gnd.t103 9.56018
R8541 gnd.n3628 gnd.n1403 9.56018
R8542 gnd.n4197 gnd.n1085 9.45599
R8543 gnd.n3370 gnd.n3369 9.45599
R8544 gnd.n5645 gnd.n5644 9.45567
R8545 gnd.n5613 gnd.n5612 9.45567
R8546 gnd.n5581 gnd.n5580 9.45567
R8547 gnd.n5550 gnd.n5549 9.45567
R8548 gnd.n5518 gnd.n5517 9.45567
R8549 gnd.n5486 gnd.n5485 9.45567
R8550 gnd.n5454 gnd.n5453 9.45567
R8551 gnd.n5423 gnd.n5422 9.45567
R8552 gnd.n5023 gnd.n5022 9.39724
R8553 gnd.n5644 gnd.n5643 9.3005
R8554 gnd.n5617 gnd.n5616 9.3005
R8555 gnd.n5638 gnd.n5637 9.3005
R8556 gnd.n5636 gnd.n5635 9.3005
R8557 gnd.n5621 gnd.n5620 9.3005
R8558 gnd.n5630 gnd.n5629 9.3005
R8559 gnd.n5628 gnd.n5627 9.3005
R8560 gnd.n5612 gnd.n5611 9.3005
R8561 gnd.n5585 gnd.n5584 9.3005
R8562 gnd.n5606 gnd.n5605 9.3005
R8563 gnd.n5604 gnd.n5603 9.3005
R8564 gnd.n5589 gnd.n5588 9.3005
R8565 gnd.n5598 gnd.n5597 9.3005
R8566 gnd.n5596 gnd.n5595 9.3005
R8567 gnd.n5580 gnd.n5579 9.3005
R8568 gnd.n5553 gnd.n5552 9.3005
R8569 gnd.n5574 gnd.n5573 9.3005
R8570 gnd.n5572 gnd.n5571 9.3005
R8571 gnd.n5557 gnd.n5556 9.3005
R8572 gnd.n5566 gnd.n5565 9.3005
R8573 gnd.n5564 gnd.n5563 9.3005
R8574 gnd.n5549 gnd.n5548 9.3005
R8575 gnd.n5522 gnd.n5521 9.3005
R8576 gnd.n5543 gnd.n5542 9.3005
R8577 gnd.n5541 gnd.n5540 9.3005
R8578 gnd.n5526 gnd.n5525 9.3005
R8579 gnd.n5535 gnd.n5534 9.3005
R8580 gnd.n5533 gnd.n5532 9.3005
R8581 gnd.n5517 gnd.n5516 9.3005
R8582 gnd.n5490 gnd.n5489 9.3005
R8583 gnd.n5511 gnd.n5510 9.3005
R8584 gnd.n5509 gnd.n5508 9.3005
R8585 gnd.n5494 gnd.n5493 9.3005
R8586 gnd.n5503 gnd.n5502 9.3005
R8587 gnd.n5501 gnd.n5500 9.3005
R8588 gnd.n5485 gnd.n5484 9.3005
R8589 gnd.n5458 gnd.n5457 9.3005
R8590 gnd.n5479 gnd.n5478 9.3005
R8591 gnd.n5477 gnd.n5476 9.3005
R8592 gnd.n5462 gnd.n5461 9.3005
R8593 gnd.n5471 gnd.n5470 9.3005
R8594 gnd.n5469 gnd.n5468 9.3005
R8595 gnd.n5453 gnd.n5452 9.3005
R8596 gnd.n5426 gnd.n5425 9.3005
R8597 gnd.n5447 gnd.n5446 9.3005
R8598 gnd.n5445 gnd.n5444 9.3005
R8599 gnd.n5430 gnd.n5429 9.3005
R8600 gnd.n5439 gnd.n5438 9.3005
R8601 gnd.n5437 gnd.n5436 9.3005
R8602 gnd.n5422 gnd.n5421 9.3005
R8603 gnd.n5395 gnd.n5394 9.3005
R8604 gnd.n5416 gnd.n5415 9.3005
R8605 gnd.n5414 gnd.n5413 9.3005
R8606 gnd.n5399 gnd.n5398 9.3005
R8607 gnd.n5408 gnd.n5407 9.3005
R8608 gnd.n5406 gnd.n5405 9.3005
R8609 gnd.n5792 gnd.n4413 9.3005
R8610 gnd.n5791 gnd.n4415 9.3005
R8611 gnd.n4419 gnd.n4416 9.3005
R8612 gnd.n5786 gnd.n4420 9.3005
R8613 gnd.n5785 gnd.n4421 9.3005
R8614 gnd.n5784 gnd.n4422 9.3005
R8615 gnd.n4426 gnd.n4423 9.3005
R8616 gnd.n5779 gnd.n4427 9.3005
R8617 gnd.n5778 gnd.n4428 9.3005
R8618 gnd.n5777 gnd.n4429 9.3005
R8619 gnd.n4433 gnd.n4430 9.3005
R8620 gnd.n5772 gnd.n4434 9.3005
R8621 gnd.n5771 gnd.n4435 9.3005
R8622 gnd.n5770 gnd.n4436 9.3005
R8623 gnd.n4441 gnd.n4439 9.3005
R8624 gnd.n5765 gnd.n5764 9.3005
R8625 gnd.n5794 gnd.n5793 9.3005
R8626 gnd.n5079 gnd.n5078 9.3005
R8627 gnd.n4709 gnd.n4708 9.3005
R8628 gnd.n5106 gnd.n5105 9.3005
R8629 gnd.n5107 gnd.n4707 9.3005
R8630 gnd.n5111 gnd.n5108 9.3005
R8631 gnd.n5110 gnd.n5109 9.3005
R8632 gnd.n4683 gnd.n4682 9.3005
R8633 gnd.n5137 gnd.n5136 9.3005
R8634 gnd.n5138 gnd.n4681 9.3005
R8635 gnd.n5142 gnd.n5139 9.3005
R8636 gnd.n5141 gnd.n5140 9.3005
R8637 gnd.n4658 gnd.n4657 9.3005
R8638 gnd.n5168 gnd.n5167 9.3005
R8639 gnd.n5169 gnd.n4656 9.3005
R8640 gnd.n5173 gnd.n5170 9.3005
R8641 gnd.n5172 gnd.n5171 9.3005
R8642 gnd.n4632 gnd.n4631 9.3005
R8643 gnd.n5199 gnd.n5198 9.3005
R8644 gnd.n5200 gnd.n4630 9.3005
R8645 gnd.n5204 gnd.n5201 9.3005
R8646 gnd.n5203 gnd.n5202 9.3005
R8647 gnd.n4608 gnd.n4607 9.3005
R8648 gnd.n5229 gnd.n5228 9.3005
R8649 gnd.n5230 gnd.n4606 9.3005
R8650 gnd.n5234 gnd.n5231 9.3005
R8651 gnd.n5233 gnd.n5232 9.3005
R8652 gnd.n4577 gnd.n4576 9.3005
R8653 gnd.n5283 gnd.n5282 9.3005
R8654 gnd.n5284 gnd.n4575 9.3005
R8655 gnd.n5286 gnd.n5285 9.3005
R8656 gnd.n4556 gnd.n4555 9.3005
R8657 gnd.n5313 gnd.n5312 9.3005
R8658 gnd.n5314 gnd.n4554 9.3005
R8659 gnd.n5318 gnd.n5315 9.3005
R8660 gnd.n5317 gnd.n5316 9.3005
R8661 gnd.n4532 gnd.n4531 9.3005
R8662 gnd.n5359 gnd.n5358 9.3005
R8663 gnd.n5360 gnd.n4530 9.3005
R8664 gnd.n5364 gnd.n5361 9.3005
R8665 gnd.n5363 gnd.n5362 9.3005
R8666 gnd.n4502 gnd.n4501 9.3005
R8667 gnd.n5680 gnd.n5679 9.3005
R8668 gnd.n5681 gnd.n4500 9.3005
R8669 gnd.n5689 gnd.n5682 9.3005
R8670 gnd.n5688 gnd.n5683 9.3005
R8671 gnd.n5687 gnd.n5685 9.3005
R8672 gnd.n5684 gnd.n782 9.3005
R8673 gnd.n5810 gnd.n783 9.3005
R8674 gnd.n5809 gnd.n784 9.3005
R8675 gnd.n5808 gnd.n785 9.3005
R8676 gnd.n4411 gnd.n786 9.3005
R8677 gnd.n4412 gnd.n4410 9.3005
R8678 gnd.n5796 gnd.n5795 9.3005
R8679 gnd.n5080 gnd.n5077 9.3005
R8680 gnd.n4788 gnd.n4747 9.3005
R8681 gnd.n4783 gnd.n4782 9.3005
R8682 gnd.n4781 gnd.n4748 9.3005
R8683 gnd.n4780 gnd.n4779 9.3005
R8684 gnd.n4776 gnd.n4749 9.3005
R8685 gnd.n4773 gnd.n4772 9.3005
R8686 gnd.n4771 gnd.n4750 9.3005
R8687 gnd.n4770 gnd.n4769 9.3005
R8688 gnd.n4766 gnd.n4751 9.3005
R8689 gnd.n4763 gnd.n4762 9.3005
R8690 gnd.n4761 gnd.n4752 9.3005
R8691 gnd.n4760 gnd.n4759 9.3005
R8692 gnd.n4756 gnd.n4754 9.3005
R8693 gnd.n4753 gnd.n4733 9.3005
R8694 gnd.n5074 gnd.n4732 9.3005
R8695 gnd.n5076 gnd.n5075 9.3005
R8696 gnd.n4790 gnd.n4789 9.3005
R8697 gnd.n5087 gnd.n4719 9.3005
R8698 gnd.n5094 gnd.n4720 9.3005
R8699 gnd.n5096 gnd.n5095 9.3005
R8700 gnd.n5097 gnd.n4700 9.3005
R8701 gnd.n5116 gnd.n5115 9.3005
R8702 gnd.n5118 gnd.n4693 9.3005
R8703 gnd.n5125 gnd.n4694 9.3005
R8704 gnd.n5127 gnd.n5126 9.3005
R8705 gnd.n5128 gnd.n4676 9.3005
R8706 gnd.n5147 gnd.n5146 9.3005
R8707 gnd.n5149 gnd.n4668 9.3005
R8708 gnd.n5156 gnd.n4669 9.3005
R8709 gnd.n5158 gnd.n5157 9.3005
R8710 gnd.n5159 gnd.n4650 9.3005
R8711 gnd.n5178 gnd.n5177 9.3005
R8712 gnd.n5180 gnd.n4642 9.3005
R8713 gnd.n5187 gnd.n4643 9.3005
R8714 gnd.n5189 gnd.n5188 9.3005
R8715 gnd.n5190 gnd.n4625 9.3005
R8716 gnd.n5209 gnd.n5208 9.3005
R8717 gnd.n5211 gnd.n4617 9.3005
R8718 gnd.n5218 gnd.n4618 9.3005
R8719 gnd.n5220 gnd.n5219 9.3005
R8720 gnd.n5221 gnd.n4601 9.3005
R8721 gnd.n5239 gnd.n5238 9.3005
R8722 gnd.n5241 gnd.n4586 9.3005
R8723 gnd.n5272 gnd.n4588 9.3005
R8724 gnd.n5273 gnd.n4584 9.3005
R8725 gnd.n5275 gnd.n5274 9.3005
R8726 gnd.n4572 gnd.n4567 9.3005
R8727 gnd.n5296 gnd.n4566 9.3005
R8728 gnd.n5299 gnd.n5298 9.3005
R8729 gnd.n5301 gnd.n5300 9.3005
R8730 gnd.n5304 gnd.n4549 9.3005
R8731 gnd.n5302 gnd.n4547 9.3005
R8732 gnd.n5326 gnd.n4545 9.3005
R8733 gnd.n5328 gnd.n5327 9.3005
R8734 gnd.n4523 gnd.n4522 9.3005
R8735 gnd.n5373 gnd.n5372 9.3005
R8736 gnd.n5374 gnd.n4516 9.3005
R8737 gnd.n5382 gnd.n4515 9.3005
R8738 gnd.n5385 gnd.n5384 9.3005
R8739 gnd.n5387 gnd.n4513 9.3005
R8740 gnd.n5671 gnd.n5670 9.3005
R8741 gnd.n5669 gnd.n5388 9.3005
R8742 gnd.n5390 gnd.n5389 9.3005
R8743 gnd.n5665 gnd.n5391 9.3005
R8744 gnd.n5664 gnd.n5392 9.3005
R8745 gnd.n5663 gnd.n5650 9.3005
R8746 gnd.n5660 gnd.n5652 9.3005
R8747 gnd.n5659 gnd.n5653 9.3005
R8748 gnd.n5656 gnd.n5654 9.3005
R8749 gnd.n5655 gnd.n4442 9.3005
R8750 gnd.n5085 gnd.n5084 9.3005
R8751 gnd.n5760 gnd.n4443 9.3005
R8752 gnd.n5759 gnd.n4445 9.3005
R8753 gnd.n4449 gnd.n4446 9.3005
R8754 gnd.n5754 gnd.n4450 9.3005
R8755 gnd.n5753 gnd.n4451 9.3005
R8756 gnd.n5752 gnd.n4452 9.3005
R8757 gnd.n4456 gnd.n4453 9.3005
R8758 gnd.n5747 gnd.n4457 9.3005
R8759 gnd.n5746 gnd.n4458 9.3005
R8760 gnd.n5745 gnd.n4459 9.3005
R8761 gnd.n4463 gnd.n4460 9.3005
R8762 gnd.n5740 gnd.n4464 9.3005
R8763 gnd.n5739 gnd.n4465 9.3005
R8764 gnd.n5738 gnd.n4466 9.3005
R8765 gnd.n4470 gnd.n4467 9.3005
R8766 gnd.n5733 gnd.n4471 9.3005
R8767 gnd.n5732 gnd.n4472 9.3005
R8768 gnd.n5731 gnd.n4473 9.3005
R8769 gnd.n4477 gnd.n4474 9.3005
R8770 gnd.n5726 gnd.n4478 9.3005
R8771 gnd.n5725 gnd.n4479 9.3005
R8772 gnd.n5724 gnd.n4480 9.3005
R8773 gnd.n4487 gnd.n4485 9.3005
R8774 gnd.n5719 gnd.n4488 9.3005
R8775 gnd.n5718 gnd.n4489 9.3005
R8776 gnd.n5717 gnd.n5714 9.3005
R8777 gnd.n5762 gnd.n5761 9.3005
R8778 gnd.n4594 gnd.n4593 9.3005
R8779 gnd.n5249 gnd.n5248 9.3005
R8780 gnd.n5250 gnd.n4592 9.3005
R8781 gnd.n5267 gnd.n5251 9.3005
R8782 gnd.n5266 gnd.n5252 9.3005
R8783 gnd.n5265 gnd.n5253 9.3005
R8784 gnd.n5263 gnd.n5254 9.3005
R8785 gnd.n5262 gnd.n5255 9.3005
R8786 gnd.n5260 gnd.n5256 9.3005
R8787 gnd.n5259 gnd.n5257 9.3005
R8788 gnd.n4538 gnd.n4537 9.3005
R8789 gnd.n5336 gnd.n5335 9.3005
R8790 gnd.n5337 gnd.n4536 9.3005
R8791 gnd.n5351 gnd.n5338 9.3005
R8792 gnd.n5350 gnd.n5339 9.3005
R8793 gnd.n5349 gnd.n5340 9.3005
R8794 gnd.n5347 gnd.n5341 9.3005
R8795 gnd.n5346 gnd.n5342 9.3005
R8796 gnd.n5344 gnd.n5343 9.3005
R8797 gnd.n4495 gnd.n4494 9.3005
R8798 gnd.n5695 gnd.n5694 9.3005
R8799 gnd.n5696 gnd.n4493 9.3005
R8800 gnd.n5700 gnd.n5697 9.3005
R8801 gnd.n5701 gnd.n4492 9.3005
R8802 gnd.n5705 gnd.n5704 9.3005
R8803 gnd.n5706 gnd.n4491 9.3005
R8804 gnd.n5708 gnd.n5707 9.3005
R8805 gnd.n5711 gnd.n4490 9.3005
R8806 gnd.n5713 gnd.n5712 9.3005
R8807 gnd.n4921 gnd.n4920 9.3005
R8808 gnd.n4811 gnd.n4810 9.3005
R8809 gnd.n4935 gnd.n4934 9.3005
R8810 gnd.n4936 gnd.n4809 9.3005
R8811 gnd.n4938 gnd.n4937 9.3005
R8812 gnd.n4799 gnd.n4798 9.3005
R8813 gnd.n4951 gnd.n4950 9.3005
R8814 gnd.n4952 gnd.n4797 9.3005
R8815 gnd.n5058 gnd.n4953 9.3005
R8816 gnd.n5057 gnd.n4954 9.3005
R8817 gnd.n5056 gnd.n4955 9.3005
R8818 gnd.n5055 gnd.n4956 9.3005
R8819 gnd.n5052 gnd.n4957 9.3005
R8820 gnd.n5051 gnd.n4958 9.3005
R8821 gnd.n5050 gnd.n4959 9.3005
R8822 gnd.n5048 gnd.n4960 9.3005
R8823 gnd.n5047 gnd.n4961 9.3005
R8824 gnd.n5044 gnd.n4962 9.3005
R8825 gnd.n5043 gnd.n4963 9.3005
R8826 gnd.n5042 gnd.n4964 9.3005
R8827 gnd.n5040 gnd.n4965 9.3005
R8828 gnd.n5039 gnd.n4966 9.3005
R8829 gnd.n5035 gnd.n4967 9.3005
R8830 gnd.n5034 gnd.n4968 9.3005
R8831 gnd.n5033 gnd.n4969 9.3005
R8832 gnd.n5031 gnd.n4970 9.3005
R8833 gnd.n5030 gnd.n4971 9.3005
R8834 gnd.n5027 gnd.n4972 9.3005
R8835 gnd.n4919 gnd.n4820 9.3005
R8836 gnd.n4822 gnd.n4821 9.3005
R8837 gnd.n4866 gnd.n4864 9.3005
R8838 gnd.n4867 gnd.n4863 9.3005
R8839 gnd.n4870 gnd.n4859 9.3005
R8840 gnd.n4871 gnd.n4858 9.3005
R8841 gnd.n4874 gnd.n4857 9.3005
R8842 gnd.n4875 gnd.n4856 9.3005
R8843 gnd.n4878 gnd.n4855 9.3005
R8844 gnd.n4879 gnd.n4854 9.3005
R8845 gnd.n4882 gnd.n4853 9.3005
R8846 gnd.n4883 gnd.n4852 9.3005
R8847 gnd.n4886 gnd.n4851 9.3005
R8848 gnd.n4887 gnd.n4850 9.3005
R8849 gnd.n4890 gnd.n4849 9.3005
R8850 gnd.n4891 gnd.n4848 9.3005
R8851 gnd.n4894 gnd.n4847 9.3005
R8852 gnd.n4895 gnd.n4846 9.3005
R8853 gnd.n4898 gnd.n4845 9.3005
R8854 gnd.n4899 gnd.n4844 9.3005
R8855 gnd.n4902 gnd.n4843 9.3005
R8856 gnd.n4903 gnd.n4842 9.3005
R8857 gnd.n4906 gnd.n4841 9.3005
R8858 gnd.n4908 gnd.n4840 9.3005
R8859 gnd.n4909 gnd.n4839 9.3005
R8860 gnd.n4910 gnd.n4838 9.3005
R8861 gnd.n4911 gnd.n4837 9.3005
R8862 gnd.n4918 gnd.n4917 9.3005
R8863 gnd.n4927 gnd.n4926 9.3005
R8864 gnd.n4928 gnd.n4814 9.3005
R8865 gnd.n4930 gnd.n4929 9.3005
R8866 gnd.n4805 gnd.n4804 9.3005
R8867 gnd.n4943 gnd.n4942 9.3005
R8868 gnd.n4944 gnd.n4803 9.3005
R8869 gnd.n4946 gnd.n4945 9.3005
R8870 gnd.n4792 gnd.n4791 9.3005
R8871 gnd.n5063 gnd.n5062 9.3005
R8872 gnd.n5064 gnd.n4746 9.3005
R8873 gnd.n5068 gnd.n5066 9.3005
R8874 gnd.n5067 gnd.n4725 9.3005
R8875 gnd.n5086 gnd.n4724 9.3005
R8876 gnd.n5089 gnd.n5088 9.3005
R8877 gnd.n4718 gnd.n4717 9.3005
R8878 gnd.n5100 gnd.n5098 9.3005
R8879 gnd.n5099 gnd.n4699 9.3005
R8880 gnd.n5117 gnd.n4698 9.3005
R8881 gnd.n5120 gnd.n5119 9.3005
R8882 gnd.n4692 gnd.n4691 9.3005
R8883 gnd.n5131 gnd.n5129 9.3005
R8884 gnd.n5130 gnd.n4675 9.3005
R8885 gnd.n5148 gnd.n4674 9.3005
R8886 gnd.n5151 gnd.n5150 9.3005
R8887 gnd.n4667 gnd.n4666 9.3005
R8888 gnd.n5162 gnd.n5160 9.3005
R8889 gnd.n5161 gnd.n4649 9.3005
R8890 gnd.n5179 gnd.n4648 9.3005
R8891 gnd.n5182 gnd.n5181 9.3005
R8892 gnd.n4641 gnd.n4640 9.3005
R8893 gnd.n5193 gnd.n5191 9.3005
R8894 gnd.n5192 gnd.n4624 9.3005
R8895 gnd.n5210 gnd.n4623 9.3005
R8896 gnd.n5213 gnd.n5212 9.3005
R8897 gnd.n4616 gnd.n4615 9.3005
R8898 gnd.n5223 gnd.n5222 9.3005
R8899 gnd.n4600 gnd.n4599 9.3005
R8900 gnd.n5244 gnd.n5240 9.3005
R8901 gnd.n5243 gnd.n5242 9.3005
R8902 gnd.n4587 gnd.n4583 9.3005
R8903 gnd.n5277 gnd.n5276 9.3005
R8904 gnd.n4585 gnd.n4568 9.3005
R8905 gnd.n5295 gnd.n5294 9.3005
R8906 gnd.n5297 gnd.n4564 9.3005
R8907 gnd.n5307 gnd.n4565 9.3005
R8908 gnd.n5306 gnd.n5305 9.3005
R8909 gnd.n5303 gnd.n4543 9.3005
R8910 gnd.n5331 gnd.n4544 9.3005
R8911 gnd.n5330 gnd.n5329 9.3005
R8912 gnd.n4546 gnd.n4524 9.3005
R8913 gnd.n5370 gnd.n5369 9.3005
R8914 gnd.n5371 gnd.n4517 9.3005
R8915 gnd.n5381 gnd.n5380 9.3005
R8916 gnd.n5383 gnd.n4511 9.3005
R8917 gnd.n5674 gnd.n4512 9.3005
R8918 gnd.n5673 gnd.n5672 9.3005
R8919 gnd.n4514 gnd.n770 9.3005
R8920 gnd.n5817 gnd.n771 9.3005
R8921 gnd.n5816 gnd.n772 9.3005
R8922 gnd.n5815 gnd.n773 9.3005
R8923 gnd.n5649 gnd.n774 9.3005
R8924 gnd.n5651 gnd.n794 9.3005
R8925 gnd.n5803 gnd.n795 9.3005
R8926 gnd.n5802 gnd.n796 9.3005
R8927 gnd.n5801 gnd.n797 9.3005
R8928 gnd.n4816 gnd.n4815 9.3005
R8929 gnd.n5992 gnd.n5991 9.3005
R8930 gnd.n5993 gnd.n594 9.3005
R8931 gnd.n5995 gnd.n5994 9.3005
R8932 gnd.n590 gnd.n589 9.3005
R8933 gnd.n6002 gnd.n6001 9.3005
R8934 gnd.n6003 gnd.n588 9.3005
R8935 gnd.n6005 gnd.n6004 9.3005
R8936 gnd.n584 gnd.n583 9.3005
R8937 gnd.n6012 gnd.n6011 9.3005
R8938 gnd.n6013 gnd.n582 9.3005
R8939 gnd.n6015 gnd.n6014 9.3005
R8940 gnd.n578 gnd.n577 9.3005
R8941 gnd.n6022 gnd.n6021 9.3005
R8942 gnd.n6023 gnd.n576 9.3005
R8943 gnd.n6025 gnd.n6024 9.3005
R8944 gnd.n572 gnd.n571 9.3005
R8945 gnd.n6032 gnd.n6031 9.3005
R8946 gnd.n6033 gnd.n570 9.3005
R8947 gnd.n6035 gnd.n6034 9.3005
R8948 gnd.n566 gnd.n565 9.3005
R8949 gnd.n6042 gnd.n6041 9.3005
R8950 gnd.n6043 gnd.n564 9.3005
R8951 gnd.n6045 gnd.n6044 9.3005
R8952 gnd.n560 gnd.n559 9.3005
R8953 gnd.n6052 gnd.n6051 9.3005
R8954 gnd.n6053 gnd.n558 9.3005
R8955 gnd.n6055 gnd.n6054 9.3005
R8956 gnd.n554 gnd.n553 9.3005
R8957 gnd.n6062 gnd.n6061 9.3005
R8958 gnd.n6063 gnd.n552 9.3005
R8959 gnd.n6065 gnd.n6064 9.3005
R8960 gnd.n548 gnd.n547 9.3005
R8961 gnd.n6072 gnd.n6071 9.3005
R8962 gnd.n6073 gnd.n546 9.3005
R8963 gnd.n6075 gnd.n6074 9.3005
R8964 gnd.n542 gnd.n541 9.3005
R8965 gnd.n6082 gnd.n6081 9.3005
R8966 gnd.n6083 gnd.n540 9.3005
R8967 gnd.n6085 gnd.n6084 9.3005
R8968 gnd.n536 gnd.n535 9.3005
R8969 gnd.n6092 gnd.n6091 9.3005
R8970 gnd.n6093 gnd.n534 9.3005
R8971 gnd.n6095 gnd.n6094 9.3005
R8972 gnd.n530 gnd.n529 9.3005
R8973 gnd.n6102 gnd.n6101 9.3005
R8974 gnd.n6103 gnd.n528 9.3005
R8975 gnd.n6105 gnd.n6104 9.3005
R8976 gnd.n524 gnd.n523 9.3005
R8977 gnd.n6112 gnd.n6111 9.3005
R8978 gnd.n6113 gnd.n522 9.3005
R8979 gnd.n6115 gnd.n6114 9.3005
R8980 gnd.n518 gnd.n517 9.3005
R8981 gnd.n6122 gnd.n6121 9.3005
R8982 gnd.n6123 gnd.n516 9.3005
R8983 gnd.n6125 gnd.n6124 9.3005
R8984 gnd.n512 gnd.n511 9.3005
R8985 gnd.n6132 gnd.n6131 9.3005
R8986 gnd.n6133 gnd.n510 9.3005
R8987 gnd.n6135 gnd.n6134 9.3005
R8988 gnd.n506 gnd.n505 9.3005
R8989 gnd.n6142 gnd.n6141 9.3005
R8990 gnd.n6143 gnd.n504 9.3005
R8991 gnd.n6145 gnd.n6144 9.3005
R8992 gnd.n500 gnd.n499 9.3005
R8993 gnd.n6152 gnd.n6151 9.3005
R8994 gnd.n6153 gnd.n498 9.3005
R8995 gnd.n6155 gnd.n6154 9.3005
R8996 gnd.n494 gnd.n493 9.3005
R8997 gnd.n6162 gnd.n6161 9.3005
R8998 gnd.n6163 gnd.n492 9.3005
R8999 gnd.n6165 gnd.n6164 9.3005
R9000 gnd.n488 gnd.n487 9.3005
R9001 gnd.n6172 gnd.n6171 9.3005
R9002 gnd.n6173 gnd.n486 9.3005
R9003 gnd.n6175 gnd.n6174 9.3005
R9004 gnd.n482 gnd.n481 9.3005
R9005 gnd.n6182 gnd.n6181 9.3005
R9006 gnd.n6183 gnd.n480 9.3005
R9007 gnd.n6185 gnd.n6184 9.3005
R9008 gnd.n476 gnd.n475 9.3005
R9009 gnd.n6192 gnd.n6191 9.3005
R9010 gnd.n6193 gnd.n474 9.3005
R9011 gnd.n6195 gnd.n6194 9.3005
R9012 gnd.n470 gnd.n469 9.3005
R9013 gnd.n6202 gnd.n6201 9.3005
R9014 gnd.n6203 gnd.n468 9.3005
R9015 gnd.n6205 gnd.n6204 9.3005
R9016 gnd.n464 gnd.n463 9.3005
R9017 gnd.n6212 gnd.n6211 9.3005
R9018 gnd.n6213 gnd.n462 9.3005
R9019 gnd.n6215 gnd.n6214 9.3005
R9020 gnd.n458 gnd.n457 9.3005
R9021 gnd.n6222 gnd.n6221 9.3005
R9022 gnd.n6223 gnd.n456 9.3005
R9023 gnd.n6225 gnd.n6224 9.3005
R9024 gnd.n452 gnd.n451 9.3005
R9025 gnd.n6232 gnd.n6231 9.3005
R9026 gnd.n6233 gnd.n450 9.3005
R9027 gnd.n6235 gnd.n6234 9.3005
R9028 gnd.n446 gnd.n445 9.3005
R9029 gnd.n6242 gnd.n6241 9.3005
R9030 gnd.n6243 gnd.n444 9.3005
R9031 gnd.n6245 gnd.n6244 9.3005
R9032 gnd.n440 gnd.n439 9.3005
R9033 gnd.n6252 gnd.n6251 9.3005
R9034 gnd.n6253 gnd.n438 9.3005
R9035 gnd.n6255 gnd.n6254 9.3005
R9036 gnd.n434 gnd.n433 9.3005
R9037 gnd.n6262 gnd.n6261 9.3005
R9038 gnd.n6263 gnd.n432 9.3005
R9039 gnd.n6265 gnd.n6264 9.3005
R9040 gnd.n428 gnd.n427 9.3005
R9041 gnd.n6272 gnd.n6271 9.3005
R9042 gnd.n6273 gnd.n426 9.3005
R9043 gnd.n6275 gnd.n6274 9.3005
R9044 gnd.n422 gnd.n421 9.3005
R9045 gnd.n6282 gnd.n6281 9.3005
R9046 gnd.n6283 gnd.n420 9.3005
R9047 gnd.n6285 gnd.n6284 9.3005
R9048 gnd.n416 gnd.n415 9.3005
R9049 gnd.n6292 gnd.n6291 9.3005
R9050 gnd.n6293 gnd.n414 9.3005
R9051 gnd.n6295 gnd.n6294 9.3005
R9052 gnd.n410 gnd.n409 9.3005
R9053 gnd.n6302 gnd.n6301 9.3005
R9054 gnd.n6303 gnd.n408 9.3005
R9055 gnd.n6305 gnd.n6304 9.3005
R9056 gnd.n404 gnd.n403 9.3005
R9057 gnd.n6312 gnd.n6311 9.3005
R9058 gnd.n6313 gnd.n402 9.3005
R9059 gnd.n6315 gnd.n6314 9.3005
R9060 gnd.n398 gnd.n397 9.3005
R9061 gnd.n6322 gnd.n6321 9.3005
R9062 gnd.n6323 gnd.n396 9.3005
R9063 gnd.n6325 gnd.n6324 9.3005
R9064 gnd.n392 gnd.n391 9.3005
R9065 gnd.n6332 gnd.n6331 9.3005
R9066 gnd.n6333 gnd.n390 9.3005
R9067 gnd.n6336 gnd.n6335 9.3005
R9068 gnd.n6334 gnd.n386 9.3005
R9069 gnd.n6342 gnd.n385 9.3005
R9070 gnd.n6344 gnd.n6343 9.3005
R9071 gnd.n381 gnd.n380 9.3005
R9072 gnd.n6353 gnd.n6352 9.3005
R9073 gnd.n6354 gnd.n379 9.3005
R9074 gnd.n6356 gnd.n6355 9.3005
R9075 gnd.n375 gnd.n374 9.3005
R9076 gnd.n6363 gnd.n6362 9.3005
R9077 gnd.n6364 gnd.n373 9.3005
R9078 gnd.n6366 gnd.n6365 9.3005
R9079 gnd.n369 gnd.n368 9.3005
R9080 gnd.n6373 gnd.n6372 9.3005
R9081 gnd.n6374 gnd.n367 9.3005
R9082 gnd.n6376 gnd.n6375 9.3005
R9083 gnd.n363 gnd.n362 9.3005
R9084 gnd.n6383 gnd.n6382 9.3005
R9085 gnd.n6384 gnd.n361 9.3005
R9086 gnd.n6386 gnd.n6385 9.3005
R9087 gnd.n357 gnd.n356 9.3005
R9088 gnd.n6393 gnd.n6392 9.3005
R9089 gnd.n6394 gnd.n355 9.3005
R9090 gnd.n6396 gnd.n6395 9.3005
R9091 gnd.n351 gnd.n350 9.3005
R9092 gnd.n6403 gnd.n6402 9.3005
R9093 gnd.n6404 gnd.n349 9.3005
R9094 gnd.n6406 gnd.n6405 9.3005
R9095 gnd.n345 gnd.n344 9.3005
R9096 gnd.n6413 gnd.n6412 9.3005
R9097 gnd.n6414 gnd.n343 9.3005
R9098 gnd.n6416 gnd.n6415 9.3005
R9099 gnd.n339 gnd.n338 9.3005
R9100 gnd.n6423 gnd.n6422 9.3005
R9101 gnd.n6424 gnd.n337 9.3005
R9102 gnd.n6426 gnd.n6425 9.3005
R9103 gnd.n333 gnd.n332 9.3005
R9104 gnd.n6433 gnd.n6432 9.3005
R9105 gnd.n6434 gnd.n331 9.3005
R9106 gnd.n6436 gnd.n6435 9.3005
R9107 gnd.n327 gnd.n326 9.3005
R9108 gnd.n6443 gnd.n6442 9.3005
R9109 gnd.n6444 gnd.n325 9.3005
R9110 gnd.n6446 gnd.n6445 9.3005
R9111 gnd.n321 gnd.n320 9.3005
R9112 gnd.n6453 gnd.n6452 9.3005
R9113 gnd.n6454 gnd.n319 9.3005
R9114 gnd.n6456 gnd.n6455 9.3005
R9115 gnd.n315 gnd.n314 9.3005
R9116 gnd.n6463 gnd.n6462 9.3005
R9117 gnd.n6464 gnd.n313 9.3005
R9118 gnd.n6466 gnd.n6465 9.3005
R9119 gnd.n309 gnd.n308 9.3005
R9120 gnd.n6473 gnd.n6472 9.3005
R9121 gnd.n6474 gnd.n307 9.3005
R9122 gnd.n6476 gnd.n6475 9.3005
R9123 gnd.n303 gnd.n302 9.3005
R9124 gnd.n6483 gnd.n6482 9.3005
R9125 gnd.n6484 gnd.n301 9.3005
R9126 gnd.n6486 gnd.n6485 9.3005
R9127 gnd.n297 gnd.n296 9.3005
R9128 gnd.n6493 gnd.n6492 9.3005
R9129 gnd.n6494 gnd.n295 9.3005
R9130 gnd.n6496 gnd.n6495 9.3005
R9131 gnd.n291 gnd.n290 9.3005
R9132 gnd.n6503 gnd.n6502 9.3005
R9133 gnd.n6504 gnd.n289 9.3005
R9134 gnd.n6506 gnd.n6505 9.3005
R9135 gnd.n285 gnd.n284 9.3005
R9136 gnd.n6513 gnd.n6512 9.3005
R9137 gnd.n6514 gnd.n283 9.3005
R9138 gnd.n6516 gnd.n6515 9.3005
R9139 gnd.n279 gnd.n278 9.3005
R9140 gnd.n6523 gnd.n6522 9.3005
R9141 gnd.n6524 gnd.n277 9.3005
R9142 gnd.n6526 gnd.n6525 9.3005
R9143 gnd.n273 gnd.n272 9.3005
R9144 gnd.n6533 gnd.n6532 9.3005
R9145 gnd.n6534 gnd.n271 9.3005
R9146 gnd.n6536 gnd.n6535 9.3005
R9147 gnd.n267 gnd.n266 9.3005
R9148 gnd.n6543 gnd.n6542 9.3005
R9149 gnd.n6544 gnd.n265 9.3005
R9150 gnd.n6546 gnd.n6545 9.3005
R9151 gnd.n261 gnd.n260 9.3005
R9152 gnd.n6554 gnd.n6553 9.3005
R9153 gnd.n6555 gnd.n259 9.3005
R9154 gnd.n6558 gnd.n6557 9.3005
R9155 gnd.n6346 gnd.n6345 9.3005
R9156 gnd.n6799 gnd.n89 9.3005
R9157 gnd.n6798 gnd.n91 9.3005
R9158 gnd.n95 gnd.n92 9.3005
R9159 gnd.n6793 gnd.n96 9.3005
R9160 gnd.n6792 gnd.n97 9.3005
R9161 gnd.n6791 gnd.n98 9.3005
R9162 gnd.n102 gnd.n99 9.3005
R9163 gnd.n6786 gnd.n103 9.3005
R9164 gnd.n6785 gnd.n104 9.3005
R9165 gnd.n6784 gnd.n105 9.3005
R9166 gnd.n109 gnd.n106 9.3005
R9167 gnd.n6779 gnd.n110 9.3005
R9168 gnd.n6778 gnd.n111 9.3005
R9169 gnd.n6777 gnd.n112 9.3005
R9170 gnd.n116 gnd.n113 9.3005
R9171 gnd.n6772 gnd.n117 9.3005
R9172 gnd.n6771 gnd.n118 9.3005
R9173 gnd.n6767 gnd.n119 9.3005
R9174 gnd.n123 gnd.n120 9.3005
R9175 gnd.n6762 gnd.n124 9.3005
R9176 gnd.n6761 gnd.n125 9.3005
R9177 gnd.n6760 gnd.n126 9.3005
R9178 gnd.n130 gnd.n127 9.3005
R9179 gnd.n6755 gnd.n131 9.3005
R9180 gnd.n6754 gnd.n132 9.3005
R9181 gnd.n6753 gnd.n133 9.3005
R9182 gnd.n137 gnd.n134 9.3005
R9183 gnd.n6748 gnd.n138 9.3005
R9184 gnd.n6747 gnd.n139 9.3005
R9185 gnd.n6746 gnd.n140 9.3005
R9186 gnd.n144 gnd.n141 9.3005
R9187 gnd.n6741 gnd.n145 9.3005
R9188 gnd.n6740 gnd.n146 9.3005
R9189 gnd.n6739 gnd.n147 9.3005
R9190 gnd.n151 gnd.n148 9.3005
R9191 gnd.n6734 gnd.n152 9.3005
R9192 gnd.n6733 gnd.n6732 9.3005
R9193 gnd.n6731 gnd.n155 9.3005
R9194 gnd.n6801 gnd.n6800 9.3005
R9195 gnd.n3812 gnd.n3811 9.3005
R9196 gnd.n1330 gnd.n1329 9.3005
R9197 gnd.n3826 gnd.n3825 9.3005
R9198 gnd.n3827 gnd.n1328 9.3005
R9199 gnd.n3914 gnd.n3828 9.3005
R9200 gnd.n3913 gnd.n3829 9.3005
R9201 gnd.n3912 gnd.n3830 9.3005
R9202 gnd.n3910 gnd.n3831 9.3005
R9203 gnd.n3909 gnd.n3832 9.3005
R9204 gnd.n3908 gnd.n3833 9.3005
R9205 gnd.n3906 gnd.n3834 9.3005
R9206 gnd.n3905 gnd.n3835 9.3005
R9207 gnd.n3903 gnd.n3836 9.3005
R9208 gnd.n3902 gnd.n3837 9.3005
R9209 gnd.n3901 gnd.n3838 9.3005
R9210 gnd.n3899 gnd.n3839 9.3005
R9211 gnd.n3898 gnd.n3840 9.3005
R9212 gnd.n3895 gnd.n3841 9.3005
R9213 gnd.n3894 gnd.n3842 9.3005
R9214 gnd.n3893 gnd.n3843 9.3005
R9215 gnd.n3892 gnd.n240 9.3005
R9216 gnd.n3888 gnd.n3844 9.3005
R9217 gnd.n3887 gnd.n3845 9.3005
R9218 gnd.n3885 gnd.n3846 9.3005
R9219 gnd.n3884 gnd.n3847 9.3005
R9220 gnd.n3882 gnd.n3848 9.3005
R9221 gnd.n3881 gnd.n3849 9.3005
R9222 gnd.n3879 gnd.n3850 9.3005
R9223 gnd.n3878 gnd.n3851 9.3005
R9224 gnd.n3876 gnd.n3852 9.3005
R9225 gnd.n3875 gnd.n3853 9.3005
R9226 gnd.n3873 gnd.n3854 9.3005
R9227 gnd.n3872 gnd.n3855 9.3005
R9228 gnd.n3870 gnd.n3856 9.3005
R9229 gnd.n3869 gnd.n3857 9.3005
R9230 gnd.n3867 gnd.n3858 9.3005
R9231 gnd.n3866 gnd.n3859 9.3005
R9232 gnd.n3864 gnd.n3860 9.3005
R9233 gnd.n3863 gnd.n3862 9.3005
R9234 gnd.n3861 gnd.n159 9.3005
R9235 gnd.n6728 gnd.n158 9.3005
R9236 gnd.n6730 gnd.n6729 9.3005
R9237 gnd.n3810 gnd.n1335 9.3005
R9238 gnd.n3799 gnd.n1340 9.3005
R9239 gnd.n3801 gnd.n3800 9.3005
R9240 gnd.n3798 gnd.n1342 9.3005
R9241 gnd.n3797 gnd.n3796 9.3005
R9242 gnd.n1344 gnd.n1343 9.3005
R9243 gnd.n3790 gnd.n3789 9.3005
R9244 gnd.n3788 gnd.n1346 9.3005
R9245 gnd.n3787 gnd.n3786 9.3005
R9246 gnd.n1348 gnd.n1347 9.3005
R9247 gnd.n3780 gnd.n3779 9.3005
R9248 gnd.n3778 gnd.n1350 9.3005
R9249 gnd.n3777 gnd.n3776 9.3005
R9250 gnd.n1352 gnd.n1351 9.3005
R9251 gnd.n3770 gnd.n3769 9.3005
R9252 gnd.n3768 gnd.n1354 9.3005
R9253 gnd.n3767 gnd.n3766 9.3005
R9254 gnd.n1356 gnd.n1355 9.3005
R9255 gnd.n3760 gnd.n3759 9.3005
R9256 gnd.n3758 gnd.n1358 9.3005
R9257 gnd.n1360 gnd.n1359 9.3005
R9258 gnd.n3745 gnd.n3700 9.3005
R9259 gnd.n3747 gnd.n3746 9.3005
R9260 gnd.n3744 gnd.n3702 9.3005
R9261 gnd.n3743 gnd.n3742 9.3005
R9262 gnd.n3704 gnd.n3703 9.3005
R9263 gnd.n3736 gnd.n3735 9.3005
R9264 gnd.n3734 gnd.n3706 9.3005
R9265 gnd.n3733 gnd.n3732 9.3005
R9266 gnd.n3708 gnd.n3707 9.3005
R9267 gnd.n3726 gnd.n3725 9.3005
R9268 gnd.n3724 gnd.n3710 9.3005
R9269 gnd.n3723 gnd.n3722 9.3005
R9270 gnd.n3712 gnd.n3711 9.3005
R9271 gnd.n3716 gnd.n3715 9.3005
R9272 gnd.n3714 gnd.n3713 9.3005
R9273 gnd.n1339 gnd.n1336 9.3005
R9274 gnd.n3809 gnd.n3808 9.3005
R9275 gnd.n4051 gnd.n1220 9.3005
R9276 gnd.n4050 gnd.n1221 9.3005
R9277 gnd.n1324 gnd.n1222 9.3005
R9278 gnd.n3937 gnd.n3936 9.3005
R9279 gnd.n3938 gnd.n1323 9.3005
R9280 gnd.n3942 gnd.n3939 9.3005
R9281 gnd.n3941 gnd.n3940 9.3005
R9282 gnd.n1297 gnd.n1296 9.3005
R9283 gnd.n3968 gnd.n3967 9.3005
R9284 gnd.n3969 gnd.n1295 9.3005
R9285 gnd.n3974 gnd.n3970 9.3005
R9286 gnd.n3973 gnd.n3972 9.3005
R9287 gnd.n3971 gnd.n1267 9.3005
R9288 gnd.n4006 gnd.n1268 9.3005
R9289 gnd.n4007 gnd.n212 9.3005
R9290 gnd.n6599 gnd.n211 9.3005
R9291 gnd.n6601 gnd.n6600 9.3005
R9292 gnd.n199 gnd.n198 9.3005
R9293 gnd.n6614 gnd.n6613 9.3005
R9294 gnd.n6615 gnd.n197 9.3005
R9295 gnd.n6617 gnd.n6616 9.3005
R9296 gnd.n183 gnd.n182 9.3005
R9297 gnd.n6630 gnd.n6629 9.3005
R9298 gnd.n6631 gnd.n181 9.3005
R9299 gnd.n6633 gnd.n6632 9.3005
R9300 gnd.n167 gnd.n166 9.3005
R9301 gnd.n6720 gnd.n6719 9.3005
R9302 gnd.n6721 gnd.n165 9.3005
R9303 gnd.n6723 gnd.n6722 9.3005
R9304 gnd.n88 gnd.n87 9.3005
R9305 gnd.n6803 gnd.n6802 9.3005
R9306 gnd.n4052 gnd.n1219 9.3005
R9307 gnd.n6598 gnd.n6597 9.3005
R9308 gnd.n3999 gnd.n3998 9.3005
R9309 gnd.n3997 gnd.n3995 9.3005
R9310 gnd.n3996 gnd.n253 9.3005
R9311 gnd.n6565 gnd.n254 9.3005
R9312 gnd.n6564 gnd.n255 9.3005
R9313 gnd.n6563 gnd.n256 9.3005
R9314 gnd.n6556 gnd.n257 9.3005
R9315 gnd.n2058 gnd.n2057 9.3005
R9316 gnd.n2056 gnd.n2021 9.3005
R9317 gnd.n2019 gnd.n2018 9.3005
R9318 gnd.n2306 gnd.n2305 9.3005
R9319 gnd.n2307 gnd.n2017 9.3005
R9320 gnd.n2309 gnd.n2308 9.3005
R9321 gnd.n2015 gnd.n2014 9.3005
R9322 gnd.n2314 gnd.n2313 9.3005
R9323 gnd.n2315 gnd.n2013 9.3005
R9324 gnd.n2358 gnd.n2316 9.3005
R9325 gnd.n2357 gnd.n2317 9.3005
R9326 gnd.n2356 gnd.n2318 9.3005
R9327 gnd.n2321 gnd.n2319 9.3005
R9328 gnd.n2352 gnd.n2322 9.3005
R9329 gnd.n2351 gnd.n2323 9.3005
R9330 gnd.n2350 gnd.n2324 9.3005
R9331 gnd.n2327 gnd.n2325 9.3005
R9332 gnd.n2346 gnd.n2328 9.3005
R9333 gnd.n2345 gnd.n2329 9.3005
R9334 gnd.n2344 gnd.n2330 9.3005
R9335 gnd.n2335 gnd.n2331 9.3005
R9336 gnd.n2339 gnd.n2336 9.3005
R9337 gnd.n2338 gnd.n2337 9.3005
R9338 gnd.n1841 gnd.n1840 9.3005
R9339 gnd.n2689 gnd.n2688 9.3005
R9340 gnd.n2690 gnd.n1839 9.3005
R9341 gnd.n2692 gnd.n2691 9.3005
R9342 gnd.n1828 gnd.n1827 9.3005
R9343 gnd.n2709 gnd.n2708 9.3005
R9344 gnd.n2710 gnd.n1826 9.3005
R9345 gnd.n2712 gnd.n2711 9.3005
R9346 gnd.n1815 gnd.n1814 9.3005
R9347 gnd.n2730 gnd.n2729 9.3005
R9348 gnd.n2731 gnd.n1813 9.3005
R9349 gnd.n2735 gnd.n2732 9.3005
R9350 gnd.n2734 gnd.n2733 9.3005
R9351 gnd.n1738 gnd.n1737 9.3005
R9352 gnd.n2807 gnd.n2806 9.3005
R9353 gnd.n2808 gnd.n1736 9.3005
R9354 gnd.n2812 gnd.n2809 9.3005
R9355 gnd.n2811 gnd.n2810 9.3005
R9356 gnd.n1710 gnd.n1709 9.3005
R9357 gnd.n2844 gnd.n2843 9.3005
R9358 gnd.n2845 gnd.n1708 9.3005
R9359 gnd.n2847 gnd.n2846 9.3005
R9360 gnd.n1688 gnd.n1687 9.3005
R9361 gnd.n2871 gnd.n2870 9.3005
R9362 gnd.n2872 gnd.n1686 9.3005
R9363 gnd.n2876 gnd.n2873 9.3005
R9364 gnd.n2875 gnd.n2874 9.3005
R9365 gnd.n1655 gnd.n1654 9.3005
R9366 gnd.n2913 gnd.n2912 9.3005
R9367 gnd.n2914 gnd.n1653 9.3005
R9368 gnd.n2927 gnd.n2915 9.3005
R9369 gnd.n2926 gnd.n2916 9.3005
R9370 gnd.n2925 gnd.n2917 9.3005
R9371 gnd.n2919 gnd.n2918 9.3005
R9372 gnd.n1621 gnd.n1620 9.3005
R9373 gnd.n2996 gnd.n2995 9.3005
R9374 gnd.n2997 gnd.n1619 9.3005
R9375 gnd.n2999 gnd.n2998 9.3005
R9376 gnd.n1598 gnd.n1597 9.3005
R9377 gnd.n3039 gnd.n3038 9.3005
R9378 gnd.n3040 gnd.n1596 9.3005
R9379 gnd.n3042 gnd.n3041 9.3005
R9380 gnd.n1582 gnd.n1581 9.3005
R9381 gnd.n3083 gnd.n3082 9.3005
R9382 gnd.n3084 gnd.n1580 9.3005
R9383 gnd.n3088 gnd.n3085 9.3005
R9384 gnd.n3087 gnd.n3086 9.3005
R9385 gnd.n1551 gnd.n1550 9.3005
R9386 gnd.n3129 gnd.n3128 9.3005
R9387 gnd.n3130 gnd.n1549 9.3005
R9388 gnd.n3132 gnd.n3131 9.3005
R9389 gnd.n1534 gnd.n1533 9.3005
R9390 gnd.n3190 gnd.n3189 9.3005
R9391 gnd.n3191 gnd.n1532 9.3005
R9392 gnd.n3193 gnd.n3192 9.3005
R9393 gnd.n1512 gnd.n1511 9.3005
R9394 gnd.n3218 gnd.n3217 9.3005
R9395 gnd.n3219 gnd.n1510 9.3005
R9396 gnd.n3223 gnd.n3220 9.3005
R9397 gnd.n3222 gnd.n3221 9.3005
R9398 gnd.n1484 gnd.n1483 9.3005
R9399 gnd.n3262 gnd.n3261 9.3005
R9400 gnd.n3263 gnd.n1482 9.3005
R9401 gnd.n3271 gnd.n3264 9.3005
R9402 gnd.n3270 gnd.n3265 9.3005
R9403 gnd.n3269 gnd.n3267 9.3005
R9404 gnd.n3266 gnd.n1414 9.3005
R9405 gnd.n3533 gnd.n1415 9.3005
R9406 gnd.n3532 gnd.n1416 9.3005
R9407 gnd.n3531 gnd.n1417 9.3005
R9408 gnd.n1424 gnd.n1418 9.3005
R9409 gnd.n3522 gnd.n1425 9.3005
R9410 gnd.n3521 gnd.n1426 9.3005
R9411 gnd.n3520 gnd.n1427 9.3005
R9412 gnd.n1435 gnd.n1428 9.3005
R9413 gnd.n3511 gnd.n1436 9.3005
R9414 gnd.n3510 gnd.n1437 9.3005
R9415 gnd.n3509 gnd.n1438 9.3005
R9416 gnd.n3495 gnd.n1439 9.3005
R9417 gnd.n3500 gnd.n3496 9.3005
R9418 gnd.n3499 gnd.n3498 9.3005
R9419 gnd.n3497 gnd.n1197 9.3005
R9420 gnd.n4067 gnd.n1198 9.3005
R9421 gnd.n4066 gnd.n1199 9.3005
R9422 gnd.n4065 gnd.n1200 9.3005
R9423 gnd.n1206 gnd.n1201 9.3005
R9424 gnd.n4059 gnd.n1207 9.3005
R9425 gnd.n4058 gnd.n1208 9.3005
R9426 gnd.n4057 gnd.n1209 9.3005
R9427 gnd.n3920 gnd.n1210 9.3005
R9428 gnd.n3922 gnd.n3921 9.3005
R9429 gnd.n3926 gnd.n3925 9.3005
R9430 gnd.n3927 gnd.n3919 9.3005
R9431 gnd.n3931 gnd.n3928 9.3005
R9432 gnd.n3930 gnd.n3929 9.3005
R9433 gnd.n1307 gnd.n1306 9.3005
R9434 gnd.n3957 gnd.n3956 9.3005
R9435 gnd.n3958 gnd.n1305 9.3005
R9436 gnd.n3962 gnd.n3959 9.3005
R9437 gnd.n3961 gnd.n3960 9.3005
R9438 gnd.n1279 gnd.n1278 9.3005
R9439 gnd.n3989 gnd.n3988 9.3005
R9440 gnd.n3990 gnd.n1277 9.3005
R9441 gnd.n4001 gnd.n3991 9.3005
R9442 gnd.n4000 gnd.n3992 9.3005
R9443 gnd.n2242 gnd.n2241 9.3005
R9444 gnd.n2109 gnd.n2084 9.3005
R9445 gnd.n2168 gnd.n2083 9.3005
R9446 gnd.n2170 gnd.n2169 9.3005
R9447 gnd.n2171 gnd.n2082 9.3005
R9448 gnd.n2173 gnd.n2172 9.3005
R9449 gnd.n2175 gnd.n2080 9.3005
R9450 gnd.n2177 gnd.n2176 9.3005
R9451 gnd.n2178 gnd.n2079 9.3005
R9452 gnd.n2180 gnd.n2179 9.3005
R9453 gnd.n2182 gnd.n2077 9.3005
R9454 gnd.n2184 gnd.n2183 9.3005
R9455 gnd.n2185 gnd.n2076 9.3005
R9456 gnd.n2187 gnd.n2186 9.3005
R9457 gnd.n2189 gnd.n2074 9.3005
R9458 gnd.n2191 gnd.n2190 9.3005
R9459 gnd.n2192 gnd.n2073 9.3005
R9460 gnd.n2235 gnd.n2193 9.3005
R9461 gnd.n2236 gnd.n2072 9.3005
R9462 gnd.n2239 gnd.n2238 9.3005
R9463 gnd.n2240 gnd.n2071 9.3005
R9464 gnd.n2111 gnd.n2110 9.3005
R9465 gnd.n2116 gnd.n2115 9.3005
R9466 gnd.n2119 gnd.n2104 9.3005
R9467 gnd.n2120 gnd.n2103 9.3005
R9468 gnd.n2123 gnd.n2102 9.3005
R9469 gnd.n2124 gnd.n2101 9.3005
R9470 gnd.n2127 gnd.n2100 9.3005
R9471 gnd.n2128 gnd.n2099 9.3005
R9472 gnd.n2131 gnd.n2098 9.3005
R9473 gnd.n2132 gnd.n2097 9.3005
R9474 gnd.n2135 gnd.n2096 9.3005
R9475 gnd.n2136 gnd.n2095 9.3005
R9476 gnd.n2139 gnd.n2094 9.3005
R9477 gnd.n2140 gnd.n2093 9.3005
R9478 gnd.n2143 gnd.n2092 9.3005
R9479 gnd.n2144 gnd.n2091 9.3005
R9480 gnd.n2147 gnd.n2090 9.3005
R9481 gnd.n2150 gnd.n2149 9.3005
R9482 gnd.n2114 gnd.n2108 9.3005
R9483 gnd.n2113 gnd.n2112 9.3005
R9484 gnd.n2157 gnd.n2156 9.3005
R9485 gnd.n2155 gnd.n2089 9.3005
R9486 gnd.n2154 gnd.n2153 9.3005
R9487 gnd.n2152 gnd.n901 9.3005
R9488 gnd.n4311 gnd.n902 9.3005
R9489 gnd.n4310 gnd.n903 9.3005
R9490 gnd.n4309 gnd.n904 9.3005
R9491 gnd.n920 gnd.n905 9.3005
R9492 gnd.n4299 gnd.n921 9.3005
R9493 gnd.n4298 gnd.n922 9.3005
R9494 gnd.n4297 gnd.n923 9.3005
R9495 gnd.n941 gnd.n924 9.3005
R9496 gnd.n4287 gnd.n942 9.3005
R9497 gnd.n4286 gnd.n943 9.3005
R9498 gnd.n4285 gnd.n944 9.3005
R9499 gnd.n964 gnd.n945 9.3005
R9500 gnd.n965 gnd.n963 9.3005
R9501 gnd.n4273 gnd.n966 9.3005
R9502 gnd.n4272 gnd.n967 9.3005
R9503 gnd.n4271 gnd.n968 9.3005
R9504 gnd.n2068 gnd.n969 9.3005
R9505 gnd.n4260 gnd.n982 9.3005
R9506 gnd.n4259 gnd.n983 9.3005
R9507 gnd.n4258 gnd.n984 9.3005
R9508 gnd.n1000 gnd.n985 9.3005
R9509 gnd.n4247 gnd.n1001 9.3005
R9510 gnd.n4246 gnd.n1002 9.3005
R9511 gnd.n4245 gnd.n1003 9.3005
R9512 gnd.n1020 gnd.n1004 9.3005
R9513 gnd.n4235 gnd.n1021 9.3005
R9514 gnd.n4234 gnd.n1022 9.3005
R9515 gnd.n4233 gnd.n1023 9.3005
R9516 gnd.n1042 gnd.n1024 9.3005
R9517 gnd.n4223 gnd.n1043 9.3005
R9518 gnd.n4222 gnd.n1044 9.3005
R9519 gnd.n4221 gnd.n1045 9.3005
R9520 gnd.n1063 gnd.n1046 9.3005
R9521 gnd.n4211 gnd.n1064 9.3005
R9522 gnd.n4210 gnd.n1065 9.3005
R9523 gnd.n4209 gnd.n1066 9.3005
R9524 gnd.n1084 gnd.n1067 9.3005
R9525 gnd.n4199 gnd.n4198 9.3005
R9526 gnd.n2151 gnd.n2088 9.3005
R9527 gnd.n2597 gnd.n1972 9.3005
R9528 gnd.n2600 gnd.n1971 9.3005
R9529 gnd.n2601 gnd.n1970 9.3005
R9530 gnd.n2604 gnd.n1969 9.3005
R9531 gnd.n2605 gnd.n1968 9.3005
R9532 gnd.n2608 gnd.n1967 9.3005
R9533 gnd.n2609 gnd.n1966 9.3005
R9534 gnd.n2612 gnd.n1965 9.3005
R9535 gnd.n2613 gnd.n1964 9.3005
R9536 gnd.n2616 gnd.n1963 9.3005
R9537 gnd.n2617 gnd.n1962 9.3005
R9538 gnd.n2620 gnd.n1961 9.3005
R9539 gnd.n2621 gnd.n1960 9.3005
R9540 gnd.n2622 gnd.n1959 9.3005
R9541 gnd.n1958 gnd.n1955 9.3005
R9542 gnd.n1957 gnd.n1956 9.3005
R9543 gnd.n2464 gnd.n2463 9.3005
R9544 gnd.n2460 gnd.n1977 9.3005
R9545 gnd.n2457 gnd.n1978 9.3005
R9546 gnd.n2456 gnd.n1979 9.3005
R9547 gnd.n2453 gnd.n1980 9.3005
R9548 gnd.n2452 gnd.n1981 9.3005
R9549 gnd.n2449 gnd.n1982 9.3005
R9550 gnd.n2448 gnd.n1983 9.3005
R9551 gnd.n2445 gnd.n1984 9.3005
R9552 gnd.n2444 gnd.n1985 9.3005
R9553 gnd.n2441 gnd.n1986 9.3005
R9554 gnd.n2440 gnd.n1987 9.3005
R9555 gnd.n2437 gnd.n1988 9.3005
R9556 gnd.n2436 gnd.n1989 9.3005
R9557 gnd.n2433 gnd.n1990 9.3005
R9558 gnd.n2432 gnd.n1991 9.3005
R9559 gnd.n2429 gnd.n1992 9.3005
R9560 gnd.n2428 gnd.n1993 9.3005
R9561 gnd.n2425 gnd.n2424 9.3005
R9562 gnd.n2423 gnd.n1995 9.3005
R9563 gnd.n2465 gnd.n1973 9.3005
R9564 gnd.n4325 gnd.n4324 9.3005
R9565 gnd.n4323 gnd.n879 9.3005
R9566 gnd.n4322 gnd.n4321 9.3005
R9567 gnd.n881 gnd.n880 9.3005
R9568 gnd.n2205 gnd.n2204 9.3005
R9569 gnd.n2207 gnd.n2203 9.3005
R9570 gnd.n2209 gnd.n2208 9.3005
R9571 gnd.n2210 gnd.n2202 9.3005
R9572 gnd.n2212 gnd.n2211 9.3005
R9573 gnd.n2214 gnd.n2200 9.3005
R9574 gnd.n2216 gnd.n2215 9.3005
R9575 gnd.n2217 gnd.n2199 9.3005
R9576 gnd.n2219 gnd.n2218 9.3005
R9577 gnd.n2221 gnd.n2197 9.3005
R9578 gnd.n2223 gnd.n2222 9.3005
R9579 gnd.n2224 gnd.n2196 9.3005
R9580 gnd.n2231 gnd.n2225 9.3005
R9581 gnd.n2230 gnd.n2226 9.3005
R9582 gnd.n2229 gnd.n2227 9.3005
R9583 gnd.n2070 gnd.n2069 9.3005
R9584 gnd.n2247 gnd.n2246 9.3005
R9585 gnd.n2248 gnd.n2067 9.3005
R9586 gnd.n2251 gnd.n2250 9.3005
R9587 gnd.n2249 gnd.n2034 9.3005
R9588 gnd.n2263 gnd.n2035 9.3005
R9589 gnd.n2264 gnd.n2033 9.3005
R9590 gnd.n2266 gnd.n2265 9.3005
R9591 gnd.n2267 gnd.n2032 9.3005
R9592 gnd.n2271 gnd.n2268 9.3005
R9593 gnd.n2272 gnd.n2031 9.3005
R9594 gnd.n2277 gnd.n2276 9.3005
R9595 gnd.n2278 gnd.n2030 9.3005
R9596 gnd.n2284 gnd.n2279 9.3005
R9597 gnd.n2283 gnd.n2280 9.3005
R9598 gnd.n2282 gnd.n2281 9.3005
R9599 gnd.n2006 gnd.n2005 9.3005
R9600 gnd.n2372 gnd.n2371 9.3005
R9601 gnd.n2373 gnd.n2004 9.3005
R9602 gnd.n2376 gnd.n2375 9.3005
R9603 gnd.n2374 gnd.n1999 9.3005
R9604 gnd.n2420 gnd.n1998 9.3005
R9605 gnd.n2422 gnd.n2421 9.3005
R9606 gnd.n4326 gnd.n877 9.3005
R9607 gnd.n4333 gnd.n4332 9.3005
R9608 gnd.n4334 gnd.n871 9.3005
R9609 gnd.n4337 gnd.n870 9.3005
R9610 gnd.n4338 gnd.n869 9.3005
R9611 gnd.n4341 gnd.n868 9.3005
R9612 gnd.n4342 gnd.n867 9.3005
R9613 gnd.n4345 gnd.n866 9.3005
R9614 gnd.n4346 gnd.n865 9.3005
R9615 gnd.n4349 gnd.n864 9.3005
R9616 gnd.n4350 gnd.n863 9.3005
R9617 gnd.n4353 gnd.n862 9.3005
R9618 gnd.n4354 gnd.n861 9.3005
R9619 gnd.n4357 gnd.n860 9.3005
R9620 gnd.n4358 gnd.n859 9.3005
R9621 gnd.n4361 gnd.n858 9.3005
R9622 gnd.n4362 gnd.n857 9.3005
R9623 gnd.n4365 gnd.n856 9.3005
R9624 gnd.n4366 gnd.n855 9.3005
R9625 gnd.n4369 gnd.n854 9.3005
R9626 gnd.n4371 gnd.n851 9.3005
R9627 gnd.n4374 gnd.n850 9.3005
R9628 gnd.n4375 gnd.n849 9.3005
R9629 gnd.n4378 gnd.n848 9.3005
R9630 gnd.n4379 gnd.n847 9.3005
R9631 gnd.n4382 gnd.n846 9.3005
R9632 gnd.n4383 gnd.n845 9.3005
R9633 gnd.n4386 gnd.n844 9.3005
R9634 gnd.n4387 gnd.n843 9.3005
R9635 gnd.n4390 gnd.n842 9.3005
R9636 gnd.n4391 gnd.n841 9.3005
R9637 gnd.n4394 gnd.n840 9.3005
R9638 gnd.n4395 gnd.n839 9.3005
R9639 gnd.n4398 gnd.n838 9.3005
R9640 gnd.n4400 gnd.n837 9.3005
R9641 gnd.n4401 gnd.n836 9.3005
R9642 gnd.n4402 gnd.n835 9.3005
R9643 gnd.n4403 gnd.n834 9.3005
R9644 gnd.n4331 gnd.n876 9.3005
R9645 gnd.n4330 gnd.n4329 9.3005
R9646 gnd.n2163 gnd.n2162 9.3005
R9647 gnd.n2161 gnd.n890 9.3005
R9648 gnd.n4317 gnd.n891 9.3005
R9649 gnd.n4316 gnd.n892 9.3005
R9650 gnd.n4315 gnd.n893 9.3005
R9651 gnd.n911 gnd.n894 9.3005
R9652 gnd.n4305 gnd.n912 9.3005
R9653 gnd.n4304 gnd.n913 9.3005
R9654 gnd.n4303 gnd.n914 9.3005
R9655 gnd.n930 gnd.n915 9.3005
R9656 gnd.n4293 gnd.n931 9.3005
R9657 gnd.n4292 gnd.n932 9.3005
R9658 gnd.n4291 gnd.n933 9.3005
R9659 gnd.n951 gnd.n934 9.3005
R9660 gnd.n4281 gnd.n952 9.3005
R9661 gnd.n1010 gnd.n993 9.3005
R9662 gnd.n4241 gnd.n1011 9.3005
R9663 gnd.n4240 gnd.n1012 9.3005
R9664 gnd.n4239 gnd.n1013 9.3005
R9665 gnd.n1031 gnd.n1014 9.3005
R9666 gnd.n4229 gnd.n1032 9.3005
R9667 gnd.n4228 gnd.n1033 9.3005
R9668 gnd.n4227 gnd.n1034 9.3005
R9669 gnd.n1052 gnd.n1035 9.3005
R9670 gnd.n4217 gnd.n1053 9.3005
R9671 gnd.n4216 gnd.n1054 9.3005
R9672 gnd.n4215 gnd.n1055 9.3005
R9673 gnd.n1074 gnd.n1056 9.3005
R9674 gnd.n4205 gnd.n1075 9.3005
R9675 gnd.n4204 gnd.n1076 9.3005
R9676 gnd.n4203 gnd.n1077 9.3005
R9677 gnd.n2160 gnd.n2159 9.3005
R9678 gnd.n4251 gnd.n953 9.3005
R9679 gnd.n2049 gnd.n2048 9.3005
R9680 gnd.n2050 gnd.n2041 9.3005
R9681 gnd.n2064 gnd.n2052 9.3005
R9682 gnd.n2063 gnd.n2053 9.3005
R9683 gnd.n2062 gnd.n2054 9.3005
R9684 gnd.n2059 gnd.n2055 9.3005
R9685 gnd.n2044 gnd.n2043 9.3005
R9686 gnd.n5823 gnd.n762 9.3005
R9687 gnd.n5824 gnd.n761 9.3005
R9688 gnd.n5825 gnd.n760 9.3005
R9689 gnd.n759 gnd.n755 9.3005
R9690 gnd.n5831 gnd.n754 9.3005
R9691 gnd.n5832 gnd.n753 9.3005
R9692 gnd.n5833 gnd.n752 9.3005
R9693 gnd.n751 gnd.n747 9.3005
R9694 gnd.n5839 gnd.n746 9.3005
R9695 gnd.n5840 gnd.n745 9.3005
R9696 gnd.n5841 gnd.n744 9.3005
R9697 gnd.n743 gnd.n739 9.3005
R9698 gnd.n5847 gnd.n738 9.3005
R9699 gnd.n5848 gnd.n737 9.3005
R9700 gnd.n5849 gnd.n736 9.3005
R9701 gnd.n735 gnd.n731 9.3005
R9702 gnd.n5855 gnd.n730 9.3005
R9703 gnd.n5856 gnd.n729 9.3005
R9704 gnd.n5857 gnd.n728 9.3005
R9705 gnd.n727 gnd.n723 9.3005
R9706 gnd.n5863 gnd.n722 9.3005
R9707 gnd.n5864 gnd.n721 9.3005
R9708 gnd.n5865 gnd.n720 9.3005
R9709 gnd.n719 gnd.n715 9.3005
R9710 gnd.n5871 gnd.n714 9.3005
R9711 gnd.n5872 gnd.n713 9.3005
R9712 gnd.n5873 gnd.n712 9.3005
R9713 gnd.n711 gnd.n707 9.3005
R9714 gnd.n5879 gnd.n706 9.3005
R9715 gnd.n5880 gnd.n705 9.3005
R9716 gnd.n5881 gnd.n704 9.3005
R9717 gnd.n703 gnd.n699 9.3005
R9718 gnd.n5887 gnd.n698 9.3005
R9719 gnd.n5888 gnd.n697 9.3005
R9720 gnd.n5889 gnd.n696 9.3005
R9721 gnd.n695 gnd.n691 9.3005
R9722 gnd.n5895 gnd.n690 9.3005
R9723 gnd.n5896 gnd.n689 9.3005
R9724 gnd.n5897 gnd.n688 9.3005
R9725 gnd.n687 gnd.n683 9.3005
R9726 gnd.n5903 gnd.n682 9.3005
R9727 gnd.n5904 gnd.n681 9.3005
R9728 gnd.n5905 gnd.n680 9.3005
R9729 gnd.n679 gnd.n675 9.3005
R9730 gnd.n5911 gnd.n674 9.3005
R9731 gnd.n5912 gnd.n673 9.3005
R9732 gnd.n5913 gnd.n672 9.3005
R9733 gnd.n671 gnd.n667 9.3005
R9734 gnd.n5919 gnd.n666 9.3005
R9735 gnd.n5920 gnd.n665 9.3005
R9736 gnd.n5921 gnd.n664 9.3005
R9737 gnd.n663 gnd.n659 9.3005
R9738 gnd.n5927 gnd.n658 9.3005
R9739 gnd.n5928 gnd.n657 9.3005
R9740 gnd.n5929 gnd.n656 9.3005
R9741 gnd.n655 gnd.n651 9.3005
R9742 gnd.n5935 gnd.n650 9.3005
R9743 gnd.n5936 gnd.n649 9.3005
R9744 gnd.n5937 gnd.n648 9.3005
R9745 gnd.n647 gnd.n643 9.3005
R9746 gnd.n5943 gnd.n642 9.3005
R9747 gnd.n5944 gnd.n641 9.3005
R9748 gnd.n5945 gnd.n640 9.3005
R9749 gnd.n639 gnd.n635 9.3005
R9750 gnd.n5951 gnd.n634 9.3005
R9751 gnd.n5952 gnd.n633 9.3005
R9752 gnd.n5953 gnd.n632 9.3005
R9753 gnd.n631 gnd.n627 9.3005
R9754 gnd.n5959 gnd.n626 9.3005
R9755 gnd.n5960 gnd.n625 9.3005
R9756 gnd.n5961 gnd.n624 9.3005
R9757 gnd.n623 gnd.n619 9.3005
R9758 gnd.n5967 gnd.n618 9.3005
R9759 gnd.n5968 gnd.n617 9.3005
R9760 gnd.n5969 gnd.n616 9.3005
R9761 gnd.n615 gnd.n611 9.3005
R9762 gnd.n5975 gnd.n610 9.3005
R9763 gnd.n5976 gnd.n609 9.3005
R9764 gnd.n5977 gnd.n608 9.3005
R9765 gnd.n607 gnd.n603 9.3005
R9766 gnd.n5983 gnd.n602 9.3005
R9767 gnd.n5984 gnd.n601 9.3005
R9768 gnd.n5985 gnd.n600 9.3005
R9769 gnd.n599 gnd.n595 9.3005
R9770 gnd.n2042 gnd.n763 9.3005
R9771 gnd.n3380 gnd.n3379 9.3005
R9772 gnd.n3360 gnd.n3358 9.3005
R9773 gnd.n3387 gnd.n3386 9.3005
R9774 gnd.n3354 gnd.n3353 9.3005
R9775 gnd.n3399 gnd.n3398 9.3005
R9776 gnd.n3351 gnd.n3349 9.3005
R9777 gnd.n3406 gnd.n3405 9.3005
R9778 gnd.n3345 gnd.n3344 9.3005
R9779 gnd.n3418 gnd.n3417 9.3005
R9780 gnd.n3342 gnd.n3340 9.3005
R9781 gnd.n3425 gnd.n3424 9.3005
R9782 gnd.n3336 gnd.n3335 9.3005
R9783 gnd.n3437 gnd.n3436 9.3005
R9784 gnd.n3333 gnd.n3331 9.3005
R9785 gnd.n3446 gnd.n3445 9.3005
R9786 gnd.n3444 gnd.n3325 9.3005
R9787 gnd.n3455 gnd.n3324 9.3005
R9788 gnd.n3458 gnd.n3457 9.3005
R9789 gnd.n3363 gnd.n3362 9.3005
R9790 gnd.n3448 gnd.n3447 9.3005
R9791 gnd.n3435 gnd.n3330 9.3005
R9792 gnd.n3434 gnd.n3433 9.3005
R9793 gnd.n3341 gnd.n3337 9.3005
R9794 gnd.n3427 gnd.n3426 9.3005
R9795 gnd.n3416 gnd.n3339 9.3005
R9796 gnd.n3415 gnd.n3414 9.3005
R9797 gnd.n3350 gnd.n3346 9.3005
R9798 gnd.n3408 gnd.n3407 9.3005
R9799 gnd.n3397 gnd.n3348 9.3005
R9800 gnd.n3396 gnd.n3395 9.3005
R9801 gnd.n3359 gnd.n3355 9.3005
R9802 gnd.n3389 gnd.n3388 9.3005
R9803 gnd.n3378 gnd.n3357 9.3005
R9804 gnd.n3377 gnd.n3376 9.3005
R9805 gnd.n3365 gnd.n3364 9.3005
R9806 gnd.n3332 gnd.n3328 9.3005
R9807 gnd.n3454 gnd.n3453 9.3005
R9808 gnd.n3322 gnd.n3321 9.3005
R9809 gnd.n3465 gnd.n3464 9.3005
R9810 gnd.n3466 gnd.n3320 9.3005
R9811 gnd.n3468 gnd.n3467 9.3005
R9812 gnd.n3318 gnd.n3317 9.3005
R9813 gnd.n3478 gnd.n3477 9.3005
R9814 gnd.n3479 gnd.n3316 9.3005
R9815 gnd.n3481 gnd.n3480 9.3005
R9816 gnd.n3314 gnd.n3313 9.3005
R9817 gnd.n3487 gnd.n3486 9.3005
R9818 gnd.n2682 gnd.n2681 9.3005
R9819 gnd.n1834 gnd.n1833 9.3005
R9820 gnd.n2699 gnd.n2698 9.3005
R9821 gnd.n2700 gnd.n1832 9.3005
R9822 gnd.n2702 gnd.n2701 9.3005
R9823 gnd.n1821 gnd.n1820 9.3005
R9824 gnd.n2719 gnd.n2718 9.3005
R9825 gnd.n2720 gnd.n1819 9.3005
R9826 gnd.n2722 gnd.n2721 9.3005
R9827 gnd.n1808 gnd.n1807 9.3005
R9828 gnd.n2742 gnd.n2741 9.3005
R9829 gnd.n2743 gnd.n1805 9.3005
R9830 gnd.n2748 gnd.n2747 9.3005
R9831 gnd.n2746 gnd.n1806 9.3005
R9832 gnd.n2745 gnd.n2744 9.3005
R9833 gnd.n1725 gnd.n1724 9.3005
R9834 gnd.n2826 gnd.n2825 9.3005
R9835 gnd.n2827 gnd.n1722 9.3005
R9836 gnd.n2830 gnd.n2829 9.3005
R9837 gnd.n2828 gnd.n1723 9.3005
R9838 gnd.n1695 gnd.n1694 9.3005
R9839 gnd.n2862 gnd.n2861 9.3005
R9840 gnd.n2863 gnd.n1693 9.3005
R9841 gnd.n2865 gnd.n2864 9.3005
R9842 gnd.n1674 gnd.n1673 9.3005
R9843 gnd.n2891 gnd.n2890 9.3005
R9844 gnd.n2892 gnd.n1671 9.3005
R9845 gnd.n2898 gnd.n2897 9.3005
R9846 gnd.n2896 gnd.n1672 9.3005
R9847 gnd.n2895 gnd.n2894 9.3005
R9848 gnd.n1639 gnd.n1638 9.3005
R9849 gnd.n2951 gnd.n2950 9.3005
R9850 gnd.n2952 gnd.n1636 9.3005
R9851 gnd.n2955 gnd.n2954 9.3005
R9852 gnd.n2953 gnd.n1637 9.3005
R9853 gnd.n1614 gnd.n1613 9.3005
R9854 gnd.n3005 gnd.n3004 9.3005
R9855 gnd.n3006 gnd.n1611 9.3005
R9856 gnd.n3020 gnd.n3019 9.3005
R9857 gnd.n3018 gnd.n1612 9.3005
R9858 gnd.n3017 gnd.n3016 9.3005
R9859 gnd.n3015 gnd.n3007 9.3005
R9860 gnd.n3014 gnd.n3013 9.3005
R9861 gnd.n3012 gnd.n3011 9.3005
R9862 gnd.n1568 gnd.n1567 9.3005
R9863 gnd.n3101 gnd.n3100 9.3005
R9864 gnd.n3102 gnd.n1565 9.3005
R9865 gnd.n3114 gnd.n3113 9.3005
R9866 gnd.n3112 gnd.n1566 9.3005
R9867 gnd.n3111 gnd.n3110 9.3005
R9868 gnd.n3109 gnd.n3103 9.3005
R9869 gnd.n3108 gnd.n3107 9.3005
R9870 gnd.n1528 gnd.n1527 9.3005
R9871 gnd.n3199 gnd.n3198 9.3005
R9872 gnd.n3200 gnd.n1525 9.3005
R9873 gnd.n3203 gnd.n3202 9.3005
R9874 gnd.n3201 gnd.n1526 9.3005
R9875 gnd.n1499 gnd.n1498 9.3005
R9876 gnd.n3237 gnd.n3236 9.3005
R9877 gnd.n3238 gnd.n1496 9.3005
R9878 gnd.n3248 gnd.n3247 9.3005
R9879 gnd.n3246 gnd.n1497 9.3005
R9880 gnd.n3245 gnd.n3244 9.3005
R9881 gnd.n3243 gnd.n3240 9.3005
R9882 gnd.n3239 gnd.n1463 9.3005
R9883 gnd.n3291 gnd.n1462 9.3005
R9884 gnd.n3293 gnd.n3292 9.3005
R9885 gnd.n3294 gnd.n1459 9.3005
R9886 gnd.n3296 gnd.n3295 9.3005
R9887 gnd.n3297 gnd.n1458 9.3005
R9888 gnd.n3299 gnd.n3298 9.3005
R9889 gnd.n3300 gnd.n1455 9.3005
R9890 gnd.n3302 gnd.n3301 9.3005
R9891 gnd.n3303 gnd.n1454 9.3005
R9892 gnd.n3305 gnd.n3304 9.3005
R9893 gnd.n3306 gnd.n1449 9.3005
R9894 gnd.n3308 gnd.n3307 9.3005
R9895 gnd.n3309 gnd.n1448 9.3005
R9896 gnd.n3311 gnd.n3310 9.3005
R9897 gnd.n3312 gnd.n1446 9.3005
R9898 gnd.n3490 gnd.n3489 9.3005
R9899 gnd.n3488 gnd.n1447 9.3005
R9900 gnd.n2680 gnd.n1845 9.3005
R9901 gnd.n1847 gnd.n1846 9.3005
R9902 gnd.n2399 gnd.n2396 9.3005
R9903 gnd.n2401 gnd.n2400 9.3005
R9904 gnd.n2403 gnd.n2402 9.3005
R9905 gnd.n2404 gnd.n2389 9.3005
R9906 gnd.n2406 gnd.n2405 9.3005
R9907 gnd.n2407 gnd.n2388 9.3005
R9908 gnd.n2409 gnd.n2408 9.3005
R9909 gnd.n2410 gnd.n2383 9.3005
R9910 gnd.n2679 gnd.n2678 9.3005
R9911 gnd.n2038 gnd.n2037 9.3005
R9912 gnd.n2256 gnd.n2255 9.3005
R9913 gnd.n2257 gnd.n2036 9.3005
R9914 gnd.n2259 gnd.n2258 9.3005
R9915 gnd.n2025 gnd.n2023 9.3005
R9916 gnd.n2298 gnd.n2297 9.3005
R9917 gnd.n2296 gnd.n2024 9.3005
R9918 gnd.n2295 gnd.n2294 9.3005
R9919 gnd.n2293 gnd.n2026 9.3005
R9920 gnd.n2292 gnd.n2291 9.3005
R9921 gnd.n2290 gnd.n2029 9.3005
R9922 gnd.n2289 gnd.n2288 9.3005
R9923 gnd.n2009 gnd.n2008 9.3005
R9924 gnd.n2364 gnd.n2363 9.3005
R9925 gnd.n2365 gnd.n2007 9.3005
R9926 gnd.n2367 gnd.n2366 9.3005
R9927 gnd.n2003 gnd.n2002 9.3005
R9928 gnd.n2381 gnd.n2380 9.3005
R9929 gnd.n2382 gnd.n2000 9.3005
R9930 gnd.n2416 gnd.n2415 9.3005
R9931 gnd.n2414 gnd.n2001 9.3005
R9932 gnd.n2412 gnd.n2411 9.3005
R9933 gnd.n1916 gnd.n1915 9.3005
R9934 gnd.n2631 gnd.n2630 9.3005
R9935 gnd.n2633 gnd.n2632 9.3005
R9936 gnd.n1904 gnd.n1903 9.3005
R9937 gnd.n2639 gnd.n2638 9.3005
R9938 gnd.n2641 gnd.n2640 9.3005
R9939 gnd.n1896 gnd.n1895 9.3005
R9940 gnd.n2647 gnd.n2646 9.3005
R9941 gnd.n2649 gnd.n2648 9.3005
R9942 gnd.n1886 gnd.n1885 9.3005
R9943 gnd.n2655 gnd.n2654 9.3005
R9944 gnd.n2657 gnd.n2656 9.3005
R9945 gnd.n1878 gnd.n1877 9.3005
R9946 gnd.n2663 gnd.n2662 9.3005
R9947 gnd.n2665 gnd.n2664 9.3005
R9948 gnd.n1868 gnd.n1866 9.3005
R9949 gnd.n2671 gnd.n2670 9.3005
R9950 gnd.n2672 gnd.n1865 9.3005
R9951 gnd.n1919 gnd.n1086 9.3005
R9952 gnd.n1869 gnd.n1867 9.3005
R9953 gnd.n2669 gnd.n2668 9.3005
R9954 gnd.n2667 gnd.n2666 9.3005
R9955 gnd.n1873 gnd.n1872 9.3005
R9956 gnd.n2661 gnd.n2660 9.3005
R9957 gnd.n2659 gnd.n2658 9.3005
R9958 gnd.n1882 gnd.n1881 9.3005
R9959 gnd.n2653 gnd.n2652 9.3005
R9960 gnd.n2651 gnd.n2650 9.3005
R9961 gnd.n1890 gnd.n1889 9.3005
R9962 gnd.n2645 gnd.n2644 9.3005
R9963 gnd.n2643 gnd.n2642 9.3005
R9964 gnd.n1900 gnd.n1899 9.3005
R9965 gnd.n2637 gnd.n2636 9.3005
R9966 gnd.n2635 gnd.n2634 9.3005
R9967 gnd.n1910 gnd.n1909 9.3005
R9968 gnd.n2629 gnd.n2628 9.3005
R9969 gnd.n4193 gnd.n1087 9.3005
R9970 gnd.n4192 gnd.n4191 9.3005
R9971 gnd.n4190 gnd.n1091 9.3005
R9972 gnd.n4189 gnd.n4188 9.3005
R9973 gnd.n4187 gnd.n1092 9.3005
R9974 gnd.n4186 gnd.n4185 9.3005
R9975 gnd.n4184 gnd.n1096 9.3005
R9976 gnd.n4183 gnd.n4182 9.3005
R9977 gnd.n4181 gnd.n1097 9.3005
R9978 gnd.n4180 gnd.n4179 9.3005
R9979 gnd.n4178 gnd.n1101 9.3005
R9980 gnd.n4177 gnd.n4176 9.3005
R9981 gnd.n4175 gnd.n1102 9.3005
R9982 gnd.n4174 gnd.n4173 9.3005
R9983 gnd.n4172 gnd.n1106 9.3005
R9984 gnd.n4171 gnd.n4170 9.3005
R9985 gnd.n4169 gnd.n1107 9.3005
R9986 gnd.n4168 gnd.n4167 9.3005
R9987 gnd.n4166 gnd.n1111 9.3005
R9988 gnd.n4165 gnd.n4164 9.3005
R9989 gnd.n4163 gnd.n1112 9.3005
R9990 gnd.n4162 gnd.n4161 9.3005
R9991 gnd.n4160 gnd.n1116 9.3005
R9992 gnd.n4159 gnd.n4158 9.3005
R9993 gnd.n4157 gnd.n1117 9.3005
R9994 gnd.n4156 gnd.n4155 9.3005
R9995 gnd.n4154 gnd.n1121 9.3005
R9996 gnd.n4153 gnd.n4152 9.3005
R9997 gnd.n4151 gnd.n1122 9.3005
R9998 gnd.n4150 gnd.n4149 9.3005
R9999 gnd.n4148 gnd.n1126 9.3005
R10000 gnd.n4147 gnd.n4146 9.3005
R10001 gnd.n4145 gnd.n1127 9.3005
R10002 gnd.n4144 gnd.n4143 9.3005
R10003 gnd.n4142 gnd.n1131 9.3005
R10004 gnd.n4141 gnd.n4140 9.3005
R10005 gnd.n4139 gnd.n1132 9.3005
R10006 gnd.n4138 gnd.n4137 9.3005
R10007 gnd.n4136 gnd.n1136 9.3005
R10008 gnd.n4135 gnd.n4134 9.3005
R10009 gnd.n4133 gnd.n1137 9.3005
R10010 gnd.n4132 gnd.n4131 9.3005
R10011 gnd.n4130 gnd.n1141 9.3005
R10012 gnd.n4129 gnd.n4128 9.3005
R10013 gnd.n4127 gnd.n1142 9.3005
R10014 gnd.n4126 gnd.n4125 9.3005
R10015 gnd.n4124 gnd.n1146 9.3005
R10016 gnd.n4123 gnd.n4122 9.3005
R10017 gnd.n4121 gnd.n1147 9.3005
R10018 gnd.n4120 gnd.n4119 9.3005
R10019 gnd.n4118 gnd.n1151 9.3005
R10020 gnd.n4117 gnd.n4116 9.3005
R10021 gnd.n4115 gnd.n1152 9.3005
R10022 gnd.n4114 gnd.n4113 9.3005
R10023 gnd.n4112 gnd.n1156 9.3005
R10024 gnd.n4111 gnd.n4110 9.3005
R10025 gnd.n4109 gnd.n1157 9.3005
R10026 gnd.n4108 gnd.n4107 9.3005
R10027 gnd.n4106 gnd.n1161 9.3005
R10028 gnd.n4105 gnd.n4104 9.3005
R10029 gnd.n4103 gnd.n1162 9.3005
R10030 gnd.n4102 gnd.n4101 9.3005
R10031 gnd.n4100 gnd.n1166 9.3005
R10032 gnd.n4099 gnd.n4098 9.3005
R10033 gnd.n4097 gnd.n1167 9.3005
R10034 gnd.n4096 gnd.n4095 9.3005
R10035 gnd.n4094 gnd.n1171 9.3005
R10036 gnd.n4093 gnd.n4092 9.3005
R10037 gnd.n4091 gnd.n1172 9.3005
R10038 gnd.n4090 gnd.n4089 9.3005
R10039 gnd.n4088 gnd.n1176 9.3005
R10040 gnd.n4087 gnd.n4086 9.3005
R10041 gnd.n4085 gnd.n1177 9.3005
R10042 gnd.n4084 gnd.n4083 9.3005
R10043 gnd.n4082 gnd.n1181 9.3005
R10044 gnd.n4081 gnd.n4080 9.3005
R10045 gnd.n4079 gnd.n1182 9.3005
R10046 gnd.n4078 gnd.n4077 9.3005
R10047 gnd.n4076 gnd.n1186 9.3005
R10048 gnd.n4075 gnd.n4074 9.3005
R10049 gnd.n4073 gnd.n1187 9.3005
R10050 gnd.n4072 gnd.n1190 9.3005
R10051 gnd.n4195 gnd.n4194 9.3005
R10052 gnd.n1232 gnd.n1230 9.3005
R10053 gnd.n4046 gnd.n4045 9.3005
R10054 gnd.n4044 gnd.n1231 9.3005
R10055 gnd.n4043 gnd.n4042 9.3005
R10056 gnd.n4041 gnd.n1233 9.3005
R10057 gnd.n4040 gnd.n4039 9.3005
R10058 gnd.n4038 gnd.n1237 9.3005
R10059 gnd.n4037 gnd.n4036 9.3005
R10060 gnd.n4035 gnd.n1238 9.3005
R10061 gnd.n4034 gnd.n4033 9.3005
R10062 gnd.n4032 gnd.n1242 9.3005
R10063 gnd.n4031 gnd.n4030 9.3005
R10064 gnd.n4029 gnd.n1243 9.3005
R10065 gnd.n4028 gnd.n4027 9.3005
R10066 gnd.n4026 gnd.n1247 9.3005
R10067 gnd.n4025 gnd.n4024 9.3005
R10068 gnd.n4023 gnd.n1248 9.3005
R10069 gnd.n4022 gnd.n4021 9.3005
R10070 gnd.n242 gnd.n241 9.3005
R10071 gnd.n6576 gnd.n6575 9.3005
R10072 gnd.n6577 gnd.n239 9.3005
R10073 gnd.n6579 gnd.n6578 9.3005
R10074 gnd.n228 gnd.n227 9.3005
R10075 gnd.n6590 gnd.n6589 9.3005
R10076 gnd.n6591 gnd.n226 9.3005
R10077 gnd.n6593 gnd.n6592 9.3005
R10078 gnd.n207 gnd.n206 9.3005
R10079 gnd.n6606 gnd.n6605 9.3005
R10080 gnd.n6607 gnd.n205 9.3005
R10081 gnd.n6609 gnd.n6608 9.3005
R10082 gnd.n192 gnd.n191 9.3005
R10083 gnd.n6622 gnd.n6621 9.3005
R10084 gnd.n6623 gnd.n190 9.3005
R10085 gnd.n6625 gnd.n6624 9.3005
R10086 gnd.n177 gnd.n176 9.3005
R10087 gnd.n6638 gnd.n6637 9.3005
R10088 gnd.n6639 gnd.n174 9.3005
R10089 gnd.n6715 gnd.n6714 9.3005
R10090 gnd.n6713 gnd.n175 9.3005
R10091 gnd.n6712 gnd.n6711 9.3005
R10092 gnd.n6710 gnd.n6640 9.3005
R10093 gnd.n6709 gnd.n6708 9.3005
R10094 gnd.n3368 gnd.n3367 9.3005
R10095 gnd.n6705 gnd.n6642 9.3005
R10096 gnd.n6704 gnd.n6703 9.3005
R10097 gnd.n6702 gnd.n6647 9.3005
R10098 gnd.n6701 gnd.n6700 9.3005
R10099 gnd.n6699 gnd.n6648 9.3005
R10100 gnd.n6698 gnd.n6697 9.3005
R10101 gnd.n6696 gnd.n6655 9.3005
R10102 gnd.n6695 gnd.n6694 9.3005
R10103 gnd.n6693 gnd.n6656 9.3005
R10104 gnd.n6692 gnd.n6691 9.3005
R10105 gnd.n6690 gnd.n6663 9.3005
R10106 gnd.n6689 gnd.n6688 9.3005
R10107 gnd.n6687 gnd.n6664 9.3005
R10108 gnd.n6686 gnd.n6685 9.3005
R10109 gnd.n6684 gnd.n6671 9.3005
R10110 gnd.n6683 gnd.n6682 9.3005
R10111 gnd.n6681 gnd.n6672 9.3005
R10112 gnd.n6680 gnd.n78 9.3005
R10113 gnd.n6707 gnd.n6706 9.3005
R10114 gnd.n3817 gnd.n3816 9.3005
R10115 gnd.n3818 gnd.n1331 9.3005
R10116 gnd.n3821 gnd.n3820 9.3005
R10117 gnd.n3819 gnd.n1332 9.3005
R10118 gnd.n1316 gnd.n1315 9.3005
R10119 gnd.n3947 gnd.n3946 9.3005
R10120 gnd.n3948 gnd.n1313 9.3005
R10121 gnd.n3951 gnd.n3950 9.3005
R10122 gnd.n3949 gnd.n1314 9.3005
R10123 gnd.n1287 gnd.n1286 9.3005
R10124 gnd.n3979 gnd.n3978 9.3005
R10125 gnd.n3980 gnd.n1284 9.3005
R10126 gnd.n3983 gnd.n3982 9.3005
R10127 gnd.n3981 gnd.n1285 9.3005
R10128 gnd.n1258 gnd.n1257 9.3005
R10129 gnd.n4013 gnd.n4012 9.3005
R10130 gnd.n4014 gnd.n1254 9.3005
R10131 gnd.n4017 gnd.n4016 9.3005
R10132 gnd.n4015 gnd.n1256 9.3005
R10133 gnd.n1255 gnd.n51 9.3005
R10134 gnd.n6839 gnd.n52 9.3005
R10135 gnd.n6838 gnd.n6837 9.3005
R10136 gnd.n6836 gnd.n53 9.3005
R10137 gnd.n6835 gnd.n6834 9.3005
R10138 gnd.n6833 gnd.n57 9.3005
R10139 gnd.n6832 gnd.n6831 9.3005
R10140 gnd.n6830 gnd.n58 9.3005
R10141 gnd.n6829 gnd.n6828 9.3005
R10142 gnd.n6827 gnd.n62 9.3005
R10143 gnd.n6826 gnd.n6825 9.3005
R10144 gnd.n6824 gnd.n63 9.3005
R10145 gnd.n6823 gnd.n6822 9.3005
R10146 gnd.n6821 gnd.n67 9.3005
R10147 gnd.n6820 gnd.n6819 9.3005
R10148 gnd.n6818 gnd.n68 9.3005
R10149 gnd.n6817 gnd.n6816 9.3005
R10150 gnd.n6815 gnd.n72 9.3005
R10151 gnd.n6814 gnd.n6813 9.3005
R10152 gnd.n6812 gnd.n73 9.3005
R10153 gnd.n6811 gnd.n6810 9.3005
R10154 gnd.n6809 gnd.n77 9.3005
R10155 gnd.n6808 gnd.n6807 9.3005
R10156 gnd.n1334 gnd.n1333 9.3005
R10157 gnd.n5292 gnd.t42 9.24152
R10158 gnd.n5806 gnd.t106 9.24152
R10159 gnd.t130 gnd.n791 9.24152
R10160 gnd.n2360 gnd.t222 9.24152
R10161 gnd.n3259 gnd.t269 9.24152
R10162 gnd.t87 gnd.n1320 9.24152
R10163 gnd.t20 gnd.t42 8.92286
R10164 gnd.n2850 gnd.n1705 8.92286
R10165 gnd.n2769 gnd.n1667 8.92286
R10166 gnd.n2929 gnd.t33 8.92286
R10167 gnd.n2947 gnd.t235 8.92286
R10168 gnd.n3026 gnd.n1606 8.92286
R10169 gnd.n3079 gnd.n1585 8.92286
R10170 gnd.n1558 gnd.t50 8.92286
R10171 gnd.t89 gnd.n3176 8.92286
R10172 gnd.n3208 gnd.n1520 8.92286
R10173 gnd.n3251 gnd.n3250 8.92286
R10174 gnd.n5642 gnd.n5617 8.92171
R10175 gnd.n5610 gnd.n5585 8.92171
R10176 gnd.n5578 gnd.n5553 8.92171
R10177 gnd.n5547 gnd.n5522 8.92171
R10178 gnd.n5515 gnd.n5490 8.92171
R10179 gnd.n5483 gnd.n5458 8.92171
R10180 gnd.n5451 gnd.n5426 8.92171
R10181 gnd.n5420 gnd.n5395 8.92171
R10182 gnd.n3560 gnd.n3542 8.72777
R10183 gnd.t15 gnd.n4610 8.60421
R10184 gnd.t284 gnd.n3024 8.60421
R10185 gnd.n3069 gnd.t226 8.60421
R10186 gnd.n5010 gnd.n4998 8.43467
R10187 gnd.n38 gnd.n26 8.43467
R10188 gnd.n2241 gnd.n0 8.41456
R10189 gnd.n6840 gnd.n6839 8.41456
R10190 gnd.n2841 gnd.n1712 8.28555
R10191 gnd.n2910 gnd.n2909 8.28555
R10192 gnd.n2975 gnd.n2974 8.28555
R10193 gnd.n3090 gnd.n1570 8.28555
R10194 gnd.n3169 gnd.n3168 8.28555
R10195 gnd.n3141 gnd.n1489 8.28555
R10196 gnd.n5643 gnd.n5615 8.14595
R10197 gnd.n5611 gnd.n5583 8.14595
R10198 gnd.n5579 gnd.n5551 8.14595
R10199 gnd.n5548 gnd.n5520 8.14595
R10200 gnd.n5516 gnd.n5488 8.14595
R10201 gnd.n5484 gnd.n5456 8.14595
R10202 gnd.n5452 gnd.n5424 8.14595
R10203 gnd.n5421 gnd.n5393 8.14595
R10204 gnd.n5648 gnd.n5647 7.97301
R10205 gnd.t76 gnd.n4652 7.9669
R10206 gnd.n2816 gnd.t34 7.9669
R10207 gnd.t161 gnd.t203 7.9669
R10208 gnd.n162 gnd.t95 7.9669
R10209 gnd.n6681 gnd.n6680 7.75808
R10210 gnd.n3453 gnd.n3328 7.75808
R10211 gnd.n2628 gnd.n1909 7.75808
R10212 gnd.n2112 gnd.n2108 7.75808
R10213 gnd.n2833 gnd.n1712 7.64824
R10214 gnd.n2909 gnd.n1659 7.64824
R10215 gnd.n2973 gnd.t232 7.64824
R10216 gnd.n2975 gnd.n2973 7.64824
R10217 gnd.n3098 gnd.n1570 7.64824
R10218 gnd.n3098 gnd.t240 7.64824
R10219 gnd.n3169 gnd.n3167 7.64824
R10220 gnd.n5122 gnd.t49 7.32958
R10221 gnd.n1766 gnd.n1765 7.30353
R10222 gnd.n3559 gnd.n3558 7.30353
R10223 gnd.n5082 gnd.n4727 7.01093
R10224 gnd.n4730 gnd.n4728 7.01093
R10225 gnd.n5092 gnd.n5091 7.01093
R10226 gnd.n5103 gnd.n4711 7.01093
R10227 gnd.n5102 gnd.n4714 7.01093
R10228 gnd.n5113 gnd.n4702 7.01093
R10229 gnd.n4705 gnd.n4703 7.01093
R10230 gnd.n5123 gnd.n5122 7.01093
R10231 gnd.n5134 gnd.n4685 7.01093
R10232 gnd.n5133 gnd.n4688 7.01093
R10233 gnd.n5144 gnd.n4678 7.01093
R10234 gnd.n5036 gnd.n4671 7.01093
R10235 gnd.n5165 gnd.n4660 7.01093
R10236 gnd.n5164 gnd.n4663 7.01093
R10237 gnd.n5175 gnd.n4652 7.01093
R10238 gnd.n4653 gnd.n4645 7.01093
R10239 gnd.n5196 gnd.n4634 7.01093
R10240 gnd.n5195 gnd.n4637 7.01093
R10241 gnd.n4627 gnd.n4620 7.01093
R10242 gnd.n5216 gnd.n5215 7.01093
R10243 gnd.n5226 gnd.n4610 7.01093
R10244 gnd.n5225 gnd.n4613 7.01093
R10245 gnd.n5236 gnd.n4603 7.01093
R10246 gnd.n5246 gnd.n4596 7.01093
R10247 gnd.n5270 gnd.n4590 7.01093
R10248 gnd.n5279 gnd.n4581 7.01093
R10249 gnd.n5288 gnd.n4573 7.01093
R10250 gnd.n5292 gnd.n5291 7.01093
R10251 gnd.n5310 gnd.n4558 7.01093
R10252 gnd.n5309 gnd.n4561 7.01093
R10253 gnd.n5320 gnd.n4550 7.01093
R10254 gnd.n4551 gnd.n4540 7.01093
R10255 gnd.n5355 gnd.n5354 7.01093
R10256 gnd.n5367 gnd.n5366 7.01093
R10257 gnd.n4527 gnd.n4519 7.01093
R10258 gnd.n5378 gnd.n5377 7.01093
R10259 gnd.n5677 gnd.n4504 7.01093
R10260 gnd.n5676 gnd.n4507 7.01093
R10261 gnd.n5692 gnd.n765 7.01093
R10262 gnd.n5820 gnd.n765 7.01093
R10263 gnd.n5819 gnd.n767 7.01093
R10264 gnd.n5698 gnd.n776 7.01093
R10265 gnd.n5813 gnd.n5812 7.01093
R10266 gnd.n5661 gnd.n779 7.01093
R10267 gnd.n5806 gnd.n788 7.01093
R10268 gnd.n5805 gnd.n791 7.01093
R10269 gnd.n5709 gnd.n799 7.01093
R10270 gnd.n5799 gnd.n5798 7.01093
R10271 gnd.n2783 gnd.t210 7.01093
R10272 gnd.n2850 gnd.n2849 7.01093
R10273 gnd.n2769 gnd.n1677 7.01093
R10274 gnd.n3026 gnd.n3025 7.01093
R10275 gnd.n3080 gnd.n3079 7.01093
R10276 gnd.n3208 gnd.n3207 7.01093
R10277 gnd.n3251 gnd.n1493 7.01093
R10278 gnd.t26 gnd.n1486 7.01093
R10279 gnd.n6725 gnd.n162 7.01093
R10280 gnd.n4688 gnd.t52 6.69227
R10281 gnd.n5288 gnd.t20 6.69227
R10282 gnd.n5691 gnd.t79 6.69227
R10283 gnd.t276 gnd.n1714 6.69227
R10284 gnd.t269 gnd.n3258 6.69227
R10285 gnd.n3689 gnd.n3688 6.5566
R10286 gnd.n2526 gnd.n2525 6.5566
R10287 gnd.n2587 gnd.n2533 6.5566
R10288 gnd.n3567 gnd.n3566 6.5566
R10289 gnd.n2761 gnd.n1745 6.37362
R10290 gnd.n2823 gnd.n2822 6.37362
R10291 gnd.n2782 gnd.t178 6.37362
R10292 gnd.n2888 gnd.t242 6.37362
R10293 gnd.n2940 gnd.n2939 6.37362
R10294 gnd.n2992 gnd.t232 6.37362
R10295 gnd.t240 gnd.n3097 6.37362
R10296 gnd.n3177 gnd.n1543 6.37362
R10297 gnd.n3205 gnd.t219 6.37362
R10298 gnd.n3281 gnd.n1469 6.37362
R10299 gnd.n3628 gnd.n1402 6.37362
R10300 gnd.n2400 gnd.n2395 6.20656
R10301 gnd.n6770 gnd.n6767 6.20656
R10302 gnd.n4370 gnd.n4369 6.20656
R10303 gnd.n3476 gnd.n3316 6.20656
R10304 gnd.t213 gnd.n5184 6.05496
R10305 gnd.n5185 gnd.t224 6.05496
R10306 gnd.t30 gnd.n5225 6.05496
R10307 gnd.n5324 gnd.t225 6.05496
R10308 gnd.n3025 gnd.t284 6.05496
R10309 gnd.n3080 gnd.t226 6.05496
R10310 gnd.n5645 gnd.n5615 5.81868
R10311 gnd.n5613 gnd.n5583 5.81868
R10312 gnd.n5581 gnd.n5551 5.81868
R10313 gnd.n5550 gnd.n5520 5.81868
R10314 gnd.n5518 gnd.n5488 5.81868
R10315 gnd.n5486 gnd.n5456 5.81868
R10316 gnd.n5454 gnd.n5424 5.81868
R10317 gnd.n5423 gnd.n5393 5.81868
R10318 gnd.t175 gnd.n2800 5.73631
R10319 gnd.t210 gnd.n1705 5.73631
R10320 gnd.n2868 gnd.n1690 5.73631
R10321 gnd.n2881 gnd.n1681 5.73631
R10322 gnd.n2964 gnd.n2963 5.73631
R10323 gnd.n3045 gnd.n3044 5.73631
R10324 gnd.n3157 gnd.n3156 5.73631
R10325 gnd.n3225 gnd.n1501 5.73631
R10326 gnd.n3250 gnd.t26 5.73631
R10327 gnd.t103 gnd.n1402 5.73631
R10328 gnd.n3698 gnd.n1361 5.62001
R10329 gnd.n2595 gnd.n2530 5.62001
R10330 gnd.n2595 gnd.n2591 5.62001
R10331 gnd.n3698 gnd.n1362 5.62001
R10332 gnd.n4867 gnd.n4862 5.4308
R10333 gnd.n4485 gnd.n4483 5.4308
R10334 gnd.n5236 gnd.t75 5.41765
R10335 gnd.n5280 gnd.t41 5.41765
R10336 gnd.n5356 gnd.t216 5.41765
R10337 gnd.n2752 gnd.n1770 5.41765
R10338 gnd.t9 gnd.n2880 5.41765
R10339 gnd.t271 gnd.n1515 5.41765
R10340 gnd.n2750 gnd.t110 5.09899
R10341 gnd.n2803 gnd.n2801 5.09899
R10342 gnd.n2801 gnd.t175 5.09899
R10343 gnd.n2816 gnd.n2815 5.09899
R10344 gnd.n2948 gnd.n2947 5.09899
R10345 gnd.n2922 gnd.n2921 5.09899
R10346 gnd.n3125 gnd.n3124 5.09899
R10347 gnd.n1558 gnd.n1547 5.09899
R10348 gnd.t146 gnd.n1476 5.09899
R10349 gnd.n3289 gnd.t161 5.09899
R10350 gnd.n3538 gnd.n3537 5.09899
R10351 gnd.n5643 gnd.n5642 5.04292
R10352 gnd.n5611 gnd.n5610 5.04292
R10353 gnd.n5579 gnd.n5578 5.04292
R10354 gnd.n5548 gnd.n5547 5.04292
R10355 gnd.n5516 gnd.n5515 5.04292
R10356 gnd.n5484 gnd.n5483 5.04292
R10357 gnd.n5452 gnd.n5451 5.04292
R10358 gnd.n5421 gnd.n5420 5.04292
R10359 gnd.n5022 gnd.n5021 4.82753
R10360 gnd.n50 gnd.n49 4.82753
R10361 gnd.n5206 gnd.t13 4.78034
R10362 gnd.n4561 gnd.t54 4.78034
R10363 gnd.t201 gnd.n1823 4.78034
R10364 gnd.n2881 gnd.t9 4.78034
R10365 gnd.n3157 gnd.t271 4.78034
R10366 gnd.n3695 gnd.t168 4.78034
R10367 gnd.n3513 gnd.t228 4.78034
R10368 gnd.n5026 gnd.n5025 4.74817
R10369 gnd.n4987 gnd.n4985 4.74817
R10370 gnd.n4980 gnd.n4979 4.74817
R10371 gnd.n4976 gnd.n4975 4.74817
R10372 gnd.n5025 gnd.n4974 4.74817
R10373 gnd.n4987 gnd.n4986 4.74817
R10374 gnd.n4981 gnd.n4980 4.74817
R10375 gnd.n4978 gnd.n4976 4.74817
R10376 gnd.n1265 gnd.n218 4.74817
R10377 gnd.n6570 gnd.n217 4.74817
R10378 gnd.n234 gnd.n216 4.74817
R10379 gnd.n6584 gnd.n215 4.74817
R10380 gnd.n219 gnd.n214 4.74817
R10381 gnd.n4008 gnd.n218 4.74817
R10382 gnd.n1264 gnd.n217 4.74817
R10383 gnd.n6571 gnd.n216 4.74817
R10384 gnd.n235 gnd.n215 4.74817
R10385 gnd.n6585 gnd.n214 4.74817
R10386 gnd.n4279 gnd.n4278 4.74817
R10387 gnd.n975 gnd.n955 4.74817
R10388 gnd.n4266 gnd.n4265 4.74817
R10389 gnd.n992 gnd.n976 4.74817
R10390 gnd.n4253 gnd.n4252 4.74817
R10391 gnd.n4280 gnd.n4279 4.74817
R10392 gnd.n4277 gnd.n955 4.74817
R10393 gnd.n4267 gnd.n4266 4.74817
R10394 gnd.n4264 gnd.n976 4.74817
R10395 gnd.n4254 gnd.n4253 4.74817
R10396 gnd.n5010 gnd.n5009 4.7074
R10397 gnd.n38 gnd.n37 4.7074
R10398 gnd.n5022 gnd.n5010 4.65959
R10399 gnd.n50 gnd.n38 4.65959
R10400 gnd.n3757 gnd.n3756 4.6132
R10401 gnd.n2596 gnd.n2466 4.6132
R10402 gnd.n2761 gnd.t110 4.46168
R10403 gnd.n2858 gnd.n2857 4.46168
R10404 gnd.n2867 gnd.t77 4.46168
R10405 gnd.n2879 gnd.n2878 4.46168
R10406 gnd.n3036 gnd.n3035 4.46168
R10407 gnd.n3073 gnd.n3072 4.46168
R10408 gnd.n3215 gnd.n3214 4.46168
R10409 gnd.n3226 gnd.t233 4.46168
R10410 gnd.n3232 gnd.n1503 4.46168
R10411 gnd.n3555 gnd.n3542 4.46111
R10412 gnd.n5628 gnd.n5624 4.38594
R10413 gnd.n5596 gnd.n5592 4.38594
R10414 gnd.n5564 gnd.n5560 4.38594
R10415 gnd.n5533 gnd.n5529 4.38594
R10416 gnd.n5501 gnd.n5497 4.38594
R10417 gnd.n5469 gnd.n5465 4.38594
R10418 gnd.n5437 gnd.n5433 4.38594
R10419 gnd.n5406 gnd.n5402 4.38594
R10420 gnd.n5639 gnd.n5617 4.26717
R10421 gnd.n5607 gnd.n5585 4.26717
R10422 gnd.n5575 gnd.n5553 4.26717
R10423 gnd.n5544 gnd.n5522 4.26717
R10424 gnd.n5512 gnd.n5490 4.26717
R10425 gnd.n5480 gnd.n5458 4.26717
R10426 gnd.n5448 gnd.n5426 4.26717
R10427 gnd.n5417 gnd.n5395 4.26717
R10428 gnd.n5154 gnd.t53 4.14303
R10429 gnd.n5377 gnd.t14 4.14303
R10430 gnd.t117 gnd.n1072 4.14303
R10431 gnd.t113 gnd.n1224 4.14303
R10432 gnd.n5647 gnd.n5646 4.08274
R10433 gnd.n3688 gnd.n3687 4.05904
R10434 gnd.n2525 gnd.n2524 4.05904
R10435 gnd.n2584 gnd.n2533 4.05904
R10436 gnd.n3568 gnd.n3567 4.05904
R10437 gnd.n15 gnd.n7 3.99943
R10438 gnd.n2791 gnd.n2790 3.82437
R10439 gnd.t93 gnd.n1659 3.82437
R10440 gnd.n2930 gnd.n1650 3.82437
R10441 gnd.n2981 gnd.n1624 3.82437
R10442 gnd.n3055 gnd.n3054 3.82437
R10443 gnd.n3175 gnd.n1536 3.82437
R10444 gnd.n3167 gnd.t220 3.82437
R10445 gnd.n1479 gnd.n1478 3.82437
R10446 gnd.n5647 gnd.n5519 3.70378
R10447 gnd.n5024 gnd.n5023 3.65935
R10448 gnd.n15 gnd.n14 3.60163
R10449 gnd.n5638 gnd.n5619 3.49141
R10450 gnd.n5606 gnd.n5587 3.49141
R10451 gnd.n5574 gnd.n5555 3.49141
R10452 gnd.n5543 gnd.n5524 3.49141
R10453 gnd.n5511 gnd.n5492 3.49141
R10454 gnd.n5479 gnd.n5460 3.49141
R10455 gnd.n5447 gnd.n5428 3.49141
R10456 gnd.n5416 gnd.n5397 3.49141
R10457 gnd.n2783 gnd.n2782 3.18706
R10458 gnd.n2983 gnd.t239 3.18706
R10459 gnd.n3001 gnd.n1617 3.18706
R10460 gnd.n3063 gnd.n3062 3.18706
R10461 gnd.n3117 gnd.t80 3.18706
R10462 gnd.n3259 gnd.n1486 3.18706
R10463 gnd.t53 gnd.n5153 2.8684
R10464 gnd.n2800 gnd.t34 2.8684
R10465 gnd.t178 gnd.t276 2.8684
R10466 gnd.t203 gnd.n1408 2.8684
R10467 gnd.n5011 gnd.t90 2.82907
R10468 gnd.n5011 gnd.t212 2.82907
R10469 gnd.n5013 gnd.t86 2.82907
R10470 gnd.n5013 gnd.t253 2.82907
R10471 gnd.n5015 gnd.t67 2.82907
R10472 gnd.n5015 gnd.t248 2.82907
R10473 gnd.n5017 gnd.t247 2.82907
R10474 gnd.n5017 gnd.t261 2.82907
R10475 gnd.n5019 gnd.t69 2.82907
R10476 gnd.n5019 gnd.t39 2.82907
R10477 gnd.n4988 gnd.t5 2.82907
R10478 gnd.n4988 gnd.t244 2.82907
R10479 gnd.n4990 gnd.t260 2.82907
R10480 gnd.n4990 gnd.t28 2.82907
R10481 gnd.n4992 gnd.t221 2.82907
R10482 gnd.n4992 gnd.t1 2.82907
R10483 gnd.n4994 gnd.t257 2.82907
R10484 gnd.n4994 gnd.t207 2.82907
R10485 gnd.n4996 gnd.t215 2.82907
R10486 gnd.n4996 gnd.t268 2.82907
R10487 gnd.n4999 gnd.t58 2.82907
R10488 gnd.n4999 gnd.t3 2.82907
R10489 gnd.n5001 gnd.t82 2.82907
R10490 gnd.n5001 gnd.t246 2.82907
R10491 gnd.n5003 gnd.t258 2.82907
R10492 gnd.n5003 gnd.t273 2.82907
R10493 gnd.n5005 gnd.t57 2.82907
R10494 gnd.n5005 gnd.t254 2.82907
R10495 gnd.n5007 gnd.t91 2.82907
R10496 gnd.n5007 gnd.t63 2.82907
R10497 gnd.n47 gnd.t265 2.82907
R10498 gnd.n47 gnd.t29 2.82907
R10499 gnd.n45 gnd.t19 2.82907
R10500 gnd.n45 gnd.t211 2.82907
R10501 gnd.n43 gnd.t208 2.82907
R10502 gnd.n43 gnd.t92 2.82907
R10503 gnd.n41 gnd.t267 2.82907
R10504 gnd.n41 gnd.t71 2.82907
R10505 gnd.n39 gnd.t45 2.82907
R10506 gnd.n39 gnd.t55 2.82907
R10507 gnd.n24 gnd.t264 2.82907
R10508 gnd.n24 gnd.t287 2.82907
R10509 gnd.n22 gnd.t245 2.82907
R10510 gnd.n22 gnd.t280 2.82907
R10511 gnd.n20 gnd.t266 2.82907
R10512 gnd.n20 gnd.t205 2.82907
R10513 gnd.n18 gnd.t218 2.82907
R10514 gnd.n18 gnd.t85 2.82907
R10515 gnd.n16 gnd.t281 2.82907
R10516 gnd.n16 gnd.t72 2.82907
R10517 gnd.n35 gnd.t74 2.82907
R10518 gnd.n35 gnd.t23 2.82907
R10519 gnd.n33 gnd.t256 2.82907
R10520 gnd.n33 gnd.t84 2.82907
R10521 gnd.n31 gnd.t17 2.82907
R10522 gnd.n31 gnd.t62 2.82907
R10523 gnd.n29 gnd.t65 2.82907
R10524 gnd.n29 gnd.t255 2.82907
R10525 gnd.n27 gnd.t78 2.82907
R10526 gnd.n27 gnd.t47 2.82907
R10527 gnd.n5635 gnd.n5634 2.71565
R10528 gnd.n5603 gnd.n5602 2.71565
R10529 gnd.n5571 gnd.n5570 2.71565
R10530 gnd.n5540 gnd.n5539 2.71565
R10531 gnd.n5508 gnd.n5507 2.71565
R10532 gnd.n5476 gnd.n5475 2.71565
R10533 gnd.n5444 gnd.n5443 2.71565
R10534 gnd.n5413 gnd.n5412 2.71565
R10535 gnd.n2834 gnd.t152 2.54975
R10536 gnd.n2840 gnd.n1714 2.54975
R10537 gnd.n2900 gnd.n1657 2.54975
R10538 gnd.n3002 gnd.n1616 2.54975
R10539 gnd.t241 gnd.n3001 2.54975
R10540 gnd.n3023 gnd.t32 2.54975
R10541 gnd.t60 gnd.n3071 2.54975
R10542 gnd.n3062 gnd.t234 2.54975
R10543 gnd.n3091 gnd.n1576 2.54975
R10544 gnd.n3196 gnd.n1530 2.54975
R10545 gnd.n3258 gnd.n3257 2.54975
R10546 gnd.n3141 gnd.t146 2.54975
R10547 gnd.n5025 gnd.n5024 2.27742
R10548 gnd.n5024 gnd.n4987 2.27742
R10549 gnd.n5024 gnd.n4980 2.27742
R10550 gnd.n5024 gnd.n4976 2.27742
R10551 gnd.n6598 gnd.n218 2.27742
R10552 gnd.n6598 gnd.n217 2.27742
R10553 gnd.n6598 gnd.n216 2.27742
R10554 gnd.n6598 gnd.n215 2.27742
R10555 gnd.n6598 gnd.n214 2.27742
R10556 gnd.n4279 gnd.n953 2.27742
R10557 gnd.n955 gnd.n953 2.27742
R10558 gnd.n4266 gnd.n953 2.27742
R10559 gnd.n976 gnd.n953 2.27742
R10560 gnd.n4253 gnd.n953 2.27742
R10561 gnd.n5091 gnd.t99 2.23109
R10562 gnd.n4983 gnd.t13 2.23109
R10563 gnd.n2957 gnd.t7 2.23109
R10564 gnd.t274 gnd.n3116 2.23109
R10565 gnd.n5631 gnd.n5621 1.93989
R10566 gnd.n5599 gnd.n5589 1.93989
R10567 gnd.n5567 gnd.n5557 1.93989
R10568 gnd.n5536 gnd.n5526 1.93989
R10569 gnd.n5504 gnd.n5494 1.93989
R10570 gnd.n5472 gnd.n5462 1.93989
R10571 gnd.n5440 gnd.n5430 1.93989
R10572 gnd.n5409 gnd.n5399 1.93989
R10573 gnd.n2834 gnd.n1718 1.91244
R10574 gnd.n2902 gnd.t59 1.91244
R10575 gnd.n2923 gnd.t235 1.91244
R10576 gnd.n2993 gnd.n2992 1.91244
R10577 gnd.n3097 gnd.n1572 1.91244
R10578 gnd.t50 gnd.n1556 1.91244
R10579 gnd.n3164 gnd.t209 1.91244
R10580 gnd.n3274 gnd.n3273 1.91244
R10581 gnd.t278 gnd.n5102 1.59378
R10582 gnd.n5269 gnd.t41 1.59378
R10583 gnd.n5323 gnd.t216 1.59378
R10584 gnd.t36 gnd.n1661 1.59378
R10585 gnd.n3187 gnd.t230 1.59378
R10586 gnd.n2859 gnd.n1697 1.27512
R10587 gnd.n2888 gnd.n2887 1.27512
R10588 gnd.t59 gnd.n2901 1.27512
R10589 gnd.n3024 gnd.n3023 1.27512
R10590 gnd.n3071 gnd.n3069 1.27512
R10591 gnd.n3195 gnd.t209 1.27512
R10592 gnd.n3206 gnd.n3205 1.27512
R10593 gnd.n3149 gnd.n3148 1.27512
R10594 gnd.n4870 gnd.n4862 1.16414
R10595 gnd.n5724 gnd.n4483 1.16414
R10596 gnd.n5630 gnd.n5623 1.16414
R10597 gnd.n5598 gnd.n5591 1.16414
R10598 gnd.n5566 gnd.n5559 1.16414
R10599 gnd.n5535 gnd.n5528 1.16414
R10600 gnd.n5503 gnd.n5496 1.16414
R10601 gnd.n5471 gnd.n5464 1.16414
R10602 gnd.n5439 gnd.n5432 1.16414
R10603 gnd.n5408 gnd.n5401 1.16414
R10604 gnd.n3756 gnd.n1358 0.970197
R10605 gnd.n2596 gnd.n1973 0.970197
R10606 gnd.n5614 gnd.n5582 0.962709
R10607 gnd.n5646 gnd.n5614 0.962709
R10608 gnd.n5487 gnd.n5455 0.962709
R10609 gnd.n5519 gnd.n5487 0.962709
R10610 gnd.n5185 gnd.t213 0.956468
R10611 gnd.n5333 gnd.t225 0.956468
R10612 gnd.n4301 gnd.t68 0.956468
R10613 gnd.n2273 gnd.t4 0.956468
R10614 gnd.n2286 gnd.t2 0.956468
R10615 gnd.n2739 gnd.t282 0.956468
R10616 gnd.t7 gnd.t239 0.956468
R10617 gnd.t80 gnd.t274 0.956468
R10618 gnd.n3526 gnd.t237 0.956468
R10619 gnd.n3965 gnd.t44 0.956468
R10620 gnd.n1291 gnd.t46 0.956468
R10621 gnd.t22 gnd.n186 0.956468
R10622 gnd.n5018 gnd.n5016 0.773756
R10623 gnd.n46 gnd.n44 0.773756
R10624 gnd.n5021 gnd.n5020 0.773756
R10625 gnd.n5020 gnd.n5018 0.773756
R10626 gnd.n5016 gnd.n5014 0.773756
R10627 gnd.n5014 gnd.n5012 0.773756
R10628 gnd.n42 gnd.n40 0.773756
R10629 gnd.n44 gnd.n42 0.773756
R10630 gnd.n48 gnd.n46 0.773756
R10631 gnd.n49 gnd.n48 0.773756
R10632 gnd.n2 gnd.n1 0.672012
R10633 gnd.n3 gnd.n2 0.672012
R10634 gnd.n4 gnd.n3 0.672012
R10635 gnd.n5 gnd.n4 0.672012
R10636 gnd.n6 gnd.n5 0.672012
R10637 gnd.n7 gnd.n6 0.672012
R10638 gnd.n9 gnd.n8 0.672012
R10639 gnd.n10 gnd.n9 0.672012
R10640 gnd.n11 gnd.n10 0.672012
R10641 gnd.n12 gnd.n11 0.672012
R10642 gnd.n13 gnd.n12 0.672012
R10643 gnd.n14 gnd.n13 0.672012
R10644 gnd.n2804 gnd.n1740 0.637812
R10645 gnd.n2814 gnd.n1733 0.637812
R10646 gnd.n2823 gnd.t142 0.637812
R10647 gnd.t6 gnd.n2858 0.637812
R10648 gnd.n2940 gnd.t33 0.637812
R10649 gnd.n2937 gnd.n1641 0.637812
R10650 gnd.n2958 gnd.n1633 0.637812
R10651 gnd.n3126 gnd.n1553 0.637812
R10652 gnd.n3135 gnd.n3134 0.637812
R10653 gnd.n3177 gnd.t89 0.637812
R10654 gnd.t236 gnd.n1503 0.637812
R10655 gnd.t138 gnd.n1469 0.637812
R10656 gnd.n1471 gnd.n1465 0.637812
R10657 gnd.n3535 gnd.n1411 0.637812
R10658 gnd.n3529 gnd.t168 0.637812
R10659 gnd.n4998 gnd.n4997 0.573776
R10660 gnd.n4997 gnd.n4995 0.573776
R10661 gnd.n4995 gnd.n4993 0.573776
R10662 gnd.n4993 gnd.n4991 0.573776
R10663 gnd.n4991 gnd.n4989 0.573776
R10664 gnd.n5009 gnd.n5008 0.573776
R10665 gnd.n5008 gnd.n5006 0.573776
R10666 gnd.n5006 gnd.n5004 0.573776
R10667 gnd.n5004 gnd.n5002 0.573776
R10668 gnd.n5002 gnd.n5000 0.573776
R10669 gnd.n19 gnd.n17 0.573776
R10670 gnd.n21 gnd.n19 0.573776
R10671 gnd.n23 gnd.n21 0.573776
R10672 gnd.n25 gnd.n23 0.573776
R10673 gnd.n26 gnd.n25 0.573776
R10674 gnd.n30 gnd.n28 0.573776
R10675 gnd.n32 gnd.n30 0.573776
R10676 gnd.n34 gnd.n32 0.573776
R10677 gnd.n36 gnd.n34 0.573776
R10678 gnd.n37 gnd.n36 0.573776
R10679 gnd gnd.n0 0.551497
R10680 gnd.n6598 gnd.n213 0.5435
R10681 gnd.n2051 gnd.n953 0.5435
R10682 gnd.n2113 gnd.n2111 0.532512
R10683 gnd.n2151 gnd.n2150 0.532512
R10684 gnd.n6708 gnd.n6707 0.532512
R10685 gnd.n6808 gnd.n78 0.532512
R10686 gnd.n4196 gnd.n4195 0.523366
R10687 gnd.n3366 gnd.n1190 0.523366
R10688 gnd.n6802 gnd.n6801 0.520317
R10689 gnd.n6731 gnd.n6730 0.520317
R10690 gnd.n3810 gnd.n3809 0.520317
R10691 gnd.n3714 gnd.n1219 0.520317
R10692 gnd.n1957 gnd.n1077 0.520317
R10693 gnd.n2423 gnd.n2422 0.520317
R10694 gnd.n4330 gnd.n877 0.520317
R10695 gnd.n2160 gnd.n834 0.520317
R10696 gnd.n3488 gnd.n3487 0.489829
R10697 gnd.n2680 gnd.n2679 0.489829
R10698 gnd.n5714 gnd.n5713 0.486781
R10699 gnd.n4919 gnd.n4918 0.48678
R10700 gnd.n5795 gnd.n5794 0.480683
R10701 gnd.n5077 gnd.n5076 0.480683
R10702 gnd.n6841 gnd.n6840 0.470187
R10703 gnd.n5992 gnd.n595 0.438
R10704 gnd.n6345 gnd.n6344 0.438
R10705 gnd.n6557 gnd.n6556 0.438
R10706 gnd.n2043 gnd.n2042 0.438
R10707 gnd.n4198 gnd.n4197 0.432431
R10708 gnd.n3369 gnd.n3368 0.432431
R10709 gnd.n2403 gnd.n2395 0.388379
R10710 gnd.n5627 gnd.n5626 0.388379
R10711 gnd.n5595 gnd.n5594 0.388379
R10712 gnd.n5563 gnd.n5562 0.388379
R10713 gnd.n5532 gnd.n5531 0.388379
R10714 gnd.n5500 gnd.n5499 0.388379
R10715 gnd.n5468 gnd.n5467 0.388379
R10716 gnd.n5436 gnd.n5435 0.388379
R10717 gnd.n5405 gnd.n5404 0.388379
R10718 gnd.n6771 gnd.n6770 0.388379
R10719 gnd.n4371 gnd.n4370 0.388379
R10720 gnd.n3477 gnd.n3476 0.388379
R10721 gnd.n6841 gnd.n15 0.374463
R10722 gnd.n4509 gnd.t79 0.319156
R10723 gnd.n2233 gnd.t206 0.319156
R10724 gnd.n2066 gnd.t0 0.319156
R10725 gnd.n2261 gnd.t81 0.319156
R10726 gnd.n2686 gnd.t164 0.319156
R10727 gnd.n1662 gnd.t36 0.319156
R10728 gnd.t230 gnd.n3186 0.319156
R10729 gnd.n3493 gnd.t134 0.319156
R10730 gnd.n3896 gnd.t70 0.319156
R10731 gnd.n6567 gnd.t16 0.319156
R10732 gnd.t18 gnd.n222 0.319156
R10733 gnd.n4837 gnd.n4815 0.311721
R10734 gnd.n2414 gnd.n2413 0.302329
R10735 gnd.n3456 gnd.n1333 0.302329
R10736 gnd gnd.n6841 0.295112
R10737 gnd.n5764 gnd.n5763 0.268793
R10738 gnd.n5763 gnd.n5762 0.241354
R10739 gnd.n3757 gnd.n1359 0.229039
R10740 gnd.n3758 gnd.n3757 0.229039
R10741 gnd.n2466 gnd.n1972 0.229039
R10742 gnd.n2466 gnd.n2465 0.229039
R10743 gnd.n5065 gnd.n4790 0.206293
R10744 gnd.n5644 gnd.n5616 0.155672
R10745 gnd.n5637 gnd.n5616 0.155672
R10746 gnd.n5637 gnd.n5636 0.155672
R10747 gnd.n5636 gnd.n5620 0.155672
R10748 gnd.n5629 gnd.n5620 0.155672
R10749 gnd.n5629 gnd.n5628 0.155672
R10750 gnd.n5612 gnd.n5584 0.155672
R10751 gnd.n5605 gnd.n5584 0.155672
R10752 gnd.n5605 gnd.n5604 0.155672
R10753 gnd.n5604 gnd.n5588 0.155672
R10754 gnd.n5597 gnd.n5588 0.155672
R10755 gnd.n5597 gnd.n5596 0.155672
R10756 gnd.n5580 gnd.n5552 0.155672
R10757 gnd.n5573 gnd.n5552 0.155672
R10758 gnd.n5573 gnd.n5572 0.155672
R10759 gnd.n5572 gnd.n5556 0.155672
R10760 gnd.n5565 gnd.n5556 0.155672
R10761 gnd.n5565 gnd.n5564 0.155672
R10762 gnd.n5549 gnd.n5521 0.155672
R10763 gnd.n5542 gnd.n5521 0.155672
R10764 gnd.n5542 gnd.n5541 0.155672
R10765 gnd.n5541 gnd.n5525 0.155672
R10766 gnd.n5534 gnd.n5525 0.155672
R10767 gnd.n5534 gnd.n5533 0.155672
R10768 gnd.n5517 gnd.n5489 0.155672
R10769 gnd.n5510 gnd.n5489 0.155672
R10770 gnd.n5510 gnd.n5509 0.155672
R10771 gnd.n5509 gnd.n5493 0.155672
R10772 gnd.n5502 gnd.n5493 0.155672
R10773 gnd.n5502 gnd.n5501 0.155672
R10774 gnd.n5485 gnd.n5457 0.155672
R10775 gnd.n5478 gnd.n5457 0.155672
R10776 gnd.n5478 gnd.n5477 0.155672
R10777 gnd.n5477 gnd.n5461 0.155672
R10778 gnd.n5470 gnd.n5461 0.155672
R10779 gnd.n5470 gnd.n5469 0.155672
R10780 gnd.n5453 gnd.n5425 0.155672
R10781 gnd.n5446 gnd.n5425 0.155672
R10782 gnd.n5446 gnd.n5445 0.155672
R10783 gnd.n5445 gnd.n5429 0.155672
R10784 gnd.n5438 gnd.n5429 0.155672
R10785 gnd.n5438 gnd.n5437 0.155672
R10786 gnd.n5422 gnd.n5394 0.155672
R10787 gnd.n5415 gnd.n5394 0.155672
R10788 gnd.n5415 gnd.n5414 0.155672
R10789 gnd.n5414 gnd.n5398 0.155672
R10790 gnd.n5407 gnd.n5398 0.155672
R10791 gnd.n5407 gnd.n5406 0.155672
R10792 gnd.n5794 gnd.n4413 0.152939
R10793 gnd.n4415 gnd.n4413 0.152939
R10794 gnd.n4419 gnd.n4415 0.152939
R10795 gnd.n4420 gnd.n4419 0.152939
R10796 gnd.n4421 gnd.n4420 0.152939
R10797 gnd.n4422 gnd.n4421 0.152939
R10798 gnd.n4426 gnd.n4422 0.152939
R10799 gnd.n4427 gnd.n4426 0.152939
R10800 gnd.n4428 gnd.n4427 0.152939
R10801 gnd.n4429 gnd.n4428 0.152939
R10802 gnd.n4433 gnd.n4429 0.152939
R10803 gnd.n4434 gnd.n4433 0.152939
R10804 gnd.n4435 gnd.n4434 0.152939
R10805 gnd.n4436 gnd.n4435 0.152939
R10806 gnd.n4441 gnd.n4436 0.152939
R10807 gnd.n5764 gnd.n4441 0.152939
R10808 gnd.n5078 gnd.n5077 0.152939
R10809 gnd.n5078 gnd.n4708 0.152939
R10810 gnd.n5106 gnd.n4708 0.152939
R10811 gnd.n5107 gnd.n5106 0.152939
R10812 gnd.n5108 gnd.n5107 0.152939
R10813 gnd.n5109 gnd.n5108 0.152939
R10814 gnd.n5109 gnd.n4682 0.152939
R10815 gnd.n5137 gnd.n4682 0.152939
R10816 gnd.n5138 gnd.n5137 0.152939
R10817 gnd.n5139 gnd.n5138 0.152939
R10818 gnd.n5140 gnd.n5139 0.152939
R10819 gnd.n5140 gnd.n4657 0.152939
R10820 gnd.n5168 gnd.n4657 0.152939
R10821 gnd.n5169 gnd.n5168 0.152939
R10822 gnd.n5170 gnd.n5169 0.152939
R10823 gnd.n5171 gnd.n5170 0.152939
R10824 gnd.n5171 gnd.n4631 0.152939
R10825 gnd.n5199 gnd.n4631 0.152939
R10826 gnd.n5200 gnd.n5199 0.152939
R10827 gnd.n5201 gnd.n5200 0.152939
R10828 gnd.n5202 gnd.n5201 0.152939
R10829 gnd.n5202 gnd.n4607 0.152939
R10830 gnd.n5229 gnd.n4607 0.152939
R10831 gnd.n5230 gnd.n5229 0.152939
R10832 gnd.n5231 gnd.n5230 0.152939
R10833 gnd.n5232 gnd.n5231 0.152939
R10834 gnd.n5232 gnd.n4576 0.152939
R10835 gnd.n5283 gnd.n4576 0.152939
R10836 gnd.n5284 gnd.n5283 0.152939
R10837 gnd.n5285 gnd.n5284 0.152939
R10838 gnd.n5285 gnd.n4555 0.152939
R10839 gnd.n5313 gnd.n4555 0.152939
R10840 gnd.n5314 gnd.n5313 0.152939
R10841 gnd.n5315 gnd.n5314 0.152939
R10842 gnd.n5316 gnd.n5315 0.152939
R10843 gnd.n5316 gnd.n4531 0.152939
R10844 gnd.n5359 gnd.n4531 0.152939
R10845 gnd.n5360 gnd.n5359 0.152939
R10846 gnd.n5361 gnd.n5360 0.152939
R10847 gnd.n5362 gnd.n5361 0.152939
R10848 gnd.n5362 gnd.n4501 0.152939
R10849 gnd.n5680 gnd.n4501 0.152939
R10850 gnd.n5681 gnd.n5680 0.152939
R10851 gnd.n5682 gnd.n5681 0.152939
R10852 gnd.n5683 gnd.n5682 0.152939
R10853 gnd.n5685 gnd.n5683 0.152939
R10854 gnd.n5685 gnd.n5684 0.152939
R10855 gnd.n5684 gnd.n783 0.152939
R10856 gnd.n784 gnd.n783 0.152939
R10857 gnd.n785 gnd.n784 0.152939
R10858 gnd.n4411 gnd.n785 0.152939
R10859 gnd.n4412 gnd.n4411 0.152939
R10860 gnd.n5795 gnd.n4412 0.152939
R10861 gnd.n5076 gnd.n4732 0.152939
R10862 gnd.n4753 gnd.n4732 0.152939
R10863 gnd.n4754 gnd.n4753 0.152939
R10864 gnd.n4760 gnd.n4754 0.152939
R10865 gnd.n4761 gnd.n4760 0.152939
R10866 gnd.n4762 gnd.n4761 0.152939
R10867 gnd.n4762 gnd.n4751 0.152939
R10868 gnd.n4770 gnd.n4751 0.152939
R10869 gnd.n4771 gnd.n4770 0.152939
R10870 gnd.n4772 gnd.n4771 0.152939
R10871 gnd.n4772 gnd.n4749 0.152939
R10872 gnd.n4780 gnd.n4749 0.152939
R10873 gnd.n4781 gnd.n4780 0.152939
R10874 gnd.n4782 gnd.n4781 0.152939
R10875 gnd.n4782 gnd.n4747 0.152939
R10876 gnd.n4790 gnd.n4747 0.152939
R10877 gnd.n5762 gnd.n4443 0.152939
R10878 gnd.n4445 gnd.n4443 0.152939
R10879 gnd.n4449 gnd.n4445 0.152939
R10880 gnd.n4450 gnd.n4449 0.152939
R10881 gnd.n4451 gnd.n4450 0.152939
R10882 gnd.n4452 gnd.n4451 0.152939
R10883 gnd.n4456 gnd.n4452 0.152939
R10884 gnd.n4457 gnd.n4456 0.152939
R10885 gnd.n4458 gnd.n4457 0.152939
R10886 gnd.n4459 gnd.n4458 0.152939
R10887 gnd.n4463 gnd.n4459 0.152939
R10888 gnd.n4464 gnd.n4463 0.152939
R10889 gnd.n4465 gnd.n4464 0.152939
R10890 gnd.n4466 gnd.n4465 0.152939
R10891 gnd.n4470 gnd.n4466 0.152939
R10892 gnd.n4471 gnd.n4470 0.152939
R10893 gnd.n4472 gnd.n4471 0.152939
R10894 gnd.n4473 gnd.n4472 0.152939
R10895 gnd.n4477 gnd.n4473 0.152939
R10896 gnd.n4478 gnd.n4477 0.152939
R10897 gnd.n4479 gnd.n4478 0.152939
R10898 gnd.n4480 gnd.n4479 0.152939
R10899 gnd.n4487 gnd.n4480 0.152939
R10900 gnd.n4488 gnd.n4487 0.152939
R10901 gnd.n4489 gnd.n4488 0.152939
R10902 gnd.n5714 gnd.n4489 0.152939
R10903 gnd.n5249 gnd.n4593 0.152939
R10904 gnd.n5250 gnd.n5249 0.152939
R10905 gnd.n5251 gnd.n5250 0.152939
R10906 gnd.n5252 gnd.n5251 0.152939
R10907 gnd.n5253 gnd.n5252 0.152939
R10908 gnd.n5254 gnd.n5253 0.152939
R10909 gnd.n5255 gnd.n5254 0.152939
R10910 gnd.n5256 gnd.n5255 0.152939
R10911 gnd.n5257 gnd.n5256 0.152939
R10912 gnd.n5257 gnd.n4537 0.152939
R10913 gnd.n5336 gnd.n4537 0.152939
R10914 gnd.n5337 gnd.n5336 0.152939
R10915 gnd.n5338 gnd.n5337 0.152939
R10916 gnd.n5339 gnd.n5338 0.152939
R10917 gnd.n5340 gnd.n5339 0.152939
R10918 gnd.n5341 gnd.n5340 0.152939
R10919 gnd.n5342 gnd.n5341 0.152939
R10920 gnd.n5343 gnd.n5342 0.152939
R10921 gnd.n5343 gnd.n4494 0.152939
R10922 gnd.n5695 gnd.n4494 0.152939
R10923 gnd.n5696 gnd.n5695 0.152939
R10924 gnd.n5697 gnd.n5696 0.152939
R10925 gnd.n5697 gnd.n4492 0.152939
R10926 gnd.n5705 gnd.n4492 0.152939
R10927 gnd.n5706 gnd.n5705 0.152939
R10928 gnd.n5707 gnd.n5706 0.152939
R10929 gnd.n5707 gnd.n4490 0.152939
R10930 gnd.n5713 gnd.n4490 0.152939
R10931 gnd.n4920 gnd.n4919 0.152939
R10932 gnd.n4920 gnd.n4810 0.152939
R10933 gnd.n4935 gnd.n4810 0.152939
R10934 gnd.n4936 gnd.n4935 0.152939
R10935 gnd.n4937 gnd.n4936 0.152939
R10936 gnd.n4937 gnd.n4798 0.152939
R10937 gnd.n4951 gnd.n4798 0.152939
R10938 gnd.n4952 gnd.n4951 0.152939
R10939 gnd.n4953 gnd.n4952 0.152939
R10940 gnd.n4954 gnd.n4953 0.152939
R10941 gnd.n4955 gnd.n4954 0.152939
R10942 gnd.n4956 gnd.n4955 0.152939
R10943 gnd.n4957 gnd.n4956 0.152939
R10944 gnd.n4958 gnd.n4957 0.152939
R10945 gnd.n4959 gnd.n4958 0.152939
R10946 gnd.n4960 gnd.n4959 0.152939
R10947 gnd.n4961 gnd.n4960 0.152939
R10948 gnd.n4962 gnd.n4961 0.152939
R10949 gnd.n4963 gnd.n4962 0.152939
R10950 gnd.n4964 gnd.n4963 0.152939
R10951 gnd.n4965 gnd.n4964 0.152939
R10952 gnd.n4966 gnd.n4965 0.152939
R10953 gnd.n4967 gnd.n4966 0.152939
R10954 gnd.n4968 gnd.n4967 0.152939
R10955 gnd.n4969 gnd.n4968 0.152939
R10956 gnd.n4970 gnd.n4969 0.152939
R10957 gnd.n4971 gnd.n4970 0.152939
R10958 gnd.n4972 gnd.n4971 0.152939
R10959 gnd.n4838 gnd.n4837 0.152939
R10960 gnd.n4839 gnd.n4838 0.152939
R10961 gnd.n4840 gnd.n4839 0.152939
R10962 gnd.n4841 gnd.n4840 0.152939
R10963 gnd.n4842 gnd.n4841 0.152939
R10964 gnd.n4843 gnd.n4842 0.152939
R10965 gnd.n4844 gnd.n4843 0.152939
R10966 gnd.n4845 gnd.n4844 0.152939
R10967 gnd.n4846 gnd.n4845 0.152939
R10968 gnd.n4847 gnd.n4846 0.152939
R10969 gnd.n4848 gnd.n4847 0.152939
R10970 gnd.n4849 gnd.n4848 0.152939
R10971 gnd.n4850 gnd.n4849 0.152939
R10972 gnd.n4851 gnd.n4850 0.152939
R10973 gnd.n4852 gnd.n4851 0.152939
R10974 gnd.n4853 gnd.n4852 0.152939
R10975 gnd.n4854 gnd.n4853 0.152939
R10976 gnd.n4855 gnd.n4854 0.152939
R10977 gnd.n4856 gnd.n4855 0.152939
R10978 gnd.n4857 gnd.n4856 0.152939
R10979 gnd.n4858 gnd.n4857 0.152939
R10980 gnd.n4859 gnd.n4858 0.152939
R10981 gnd.n4863 gnd.n4859 0.152939
R10982 gnd.n4864 gnd.n4863 0.152939
R10983 gnd.n4864 gnd.n4821 0.152939
R10984 gnd.n4918 gnd.n4821 0.152939
R10985 gnd.n5993 gnd.n5992 0.152939
R10986 gnd.n5994 gnd.n5993 0.152939
R10987 gnd.n5994 gnd.n589 0.152939
R10988 gnd.n6002 gnd.n589 0.152939
R10989 gnd.n6003 gnd.n6002 0.152939
R10990 gnd.n6004 gnd.n6003 0.152939
R10991 gnd.n6004 gnd.n583 0.152939
R10992 gnd.n6012 gnd.n583 0.152939
R10993 gnd.n6013 gnd.n6012 0.152939
R10994 gnd.n6014 gnd.n6013 0.152939
R10995 gnd.n6014 gnd.n577 0.152939
R10996 gnd.n6022 gnd.n577 0.152939
R10997 gnd.n6023 gnd.n6022 0.152939
R10998 gnd.n6024 gnd.n6023 0.152939
R10999 gnd.n6024 gnd.n571 0.152939
R11000 gnd.n6032 gnd.n571 0.152939
R11001 gnd.n6033 gnd.n6032 0.152939
R11002 gnd.n6034 gnd.n6033 0.152939
R11003 gnd.n6034 gnd.n565 0.152939
R11004 gnd.n6042 gnd.n565 0.152939
R11005 gnd.n6043 gnd.n6042 0.152939
R11006 gnd.n6044 gnd.n6043 0.152939
R11007 gnd.n6044 gnd.n559 0.152939
R11008 gnd.n6052 gnd.n559 0.152939
R11009 gnd.n6053 gnd.n6052 0.152939
R11010 gnd.n6054 gnd.n6053 0.152939
R11011 gnd.n6054 gnd.n553 0.152939
R11012 gnd.n6062 gnd.n553 0.152939
R11013 gnd.n6063 gnd.n6062 0.152939
R11014 gnd.n6064 gnd.n6063 0.152939
R11015 gnd.n6064 gnd.n547 0.152939
R11016 gnd.n6072 gnd.n547 0.152939
R11017 gnd.n6073 gnd.n6072 0.152939
R11018 gnd.n6074 gnd.n6073 0.152939
R11019 gnd.n6074 gnd.n541 0.152939
R11020 gnd.n6082 gnd.n541 0.152939
R11021 gnd.n6083 gnd.n6082 0.152939
R11022 gnd.n6084 gnd.n6083 0.152939
R11023 gnd.n6084 gnd.n535 0.152939
R11024 gnd.n6092 gnd.n535 0.152939
R11025 gnd.n6093 gnd.n6092 0.152939
R11026 gnd.n6094 gnd.n6093 0.152939
R11027 gnd.n6094 gnd.n529 0.152939
R11028 gnd.n6102 gnd.n529 0.152939
R11029 gnd.n6103 gnd.n6102 0.152939
R11030 gnd.n6104 gnd.n6103 0.152939
R11031 gnd.n6104 gnd.n523 0.152939
R11032 gnd.n6112 gnd.n523 0.152939
R11033 gnd.n6113 gnd.n6112 0.152939
R11034 gnd.n6114 gnd.n6113 0.152939
R11035 gnd.n6114 gnd.n517 0.152939
R11036 gnd.n6122 gnd.n517 0.152939
R11037 gnd.n6123 gnd.n6122 0.152939
R11038 gnd.n6124 gnd.n6123 0.152939
R11039 gnd.n6124 gnd.n511 0.152939
R11040 gnd.n6132 gnd.n511 0.152939
R11041 gnd.n6133 gnd.n6132 0.152939
R11042 gnd.n6134 gnd.n6133 0.152939
R11043 gnd.n6134 gnd.n505 0.152939
R11044 gnd.n6142 gnd.n505 0.152939
R11045 gnd.n6143 gnd.n6142 0.152939
R11046 gnd.n6144 gnd.n6143 0.152939
R11047 gnd.n6144 gnd.n499 0.152939
R11048 gnd.n6152 gnd.n499 0.152939
R11049 gnd.n6153 gnd.n6152 0.152939
R11050 gnd.n6154 gnd.n6153 0.152939
R11051 gnd.n6154 gnd.n493 0.152939
R11052 gnd.n6162 gnd.n493 0.152939
R11053 gnd.n6163 gnd.n6162 0.152939
R11054 gnd.n6164 gnd.n6163 0.152939
R11055 gnd.n6164 gnd.n487 0.152939
R11056 gnd.n6172 gnd.n487 0.152939
R11057 gnd.n6173 gnd.n6172 0.152939
R11058 gnd.n6174 gnd.n6173 0.152939
R11059 gnd.n6174 gnd.n481 0.152939
R11060 gnd.n6182 gnd.n481 0.152939
R11061 gnd.n6183 gnd.n6182 0.152939
R11062 gnd.n6184 gnd.n6183 0.152939
R11063 gnd.n6184 gnd.n475 0.152939
R11064 gnd.n6192 gnd.n475 0.152939
R11065 gnd.n6193 gnd.n6192 0.152939
R11066 gnd.n6194 gnd.n6193 0.152939
R11067 gnd.n6194 gnd.n469 0.152939
R11068 gnd.n6202 gnd.n469 0.152939
R11069 gnd.n6203 gnd.n6202 0.152939
R11070 gnd.n6204 gnd.n6203 0.152939
R11071 gnd.n6204 gnd.n463 0.152939
R11072 gnd.n6212 gnd.n463 0.152939
R11073 gnd.n6213 gnd.n6212 0.152939
R11074 gnd.n6214 gnd.n6213 0.152939
R11075 gnd.n6214 gnd.n457 0.152939
R11076 gnd.n6222 gnd.n457 0.152939
R11077 gnd.n6223 gnd.n6222 0.152939
R11078 gnd.n6224 gnd.n6223 0.152939
R11079 gnd.n6224 gnd.n451 0.152939
R11080 gnd.n6232 gnd.n451 0.152939
R11081 gnd.n6233 gnd.n6232 0.152939
R11082 gnd.n6234 gnd.n6233 0.152939
R11083 gnd.n6234 gnd.n445 0.152939
R11084 gnd.n6242 gnd.n445 0.152939
R11085 gnd.n6243 gnd.n6242 0.152939
R11086 gnd.n6244 gnd.n6243 0.152939
R11087 gnd.n6244 gnd.n439 0.152939
R11088 gnd.n6252 gnd.n439 0.152939
R11089 gnd.n6253 gnd.n6252 0.152939
R11090 gnd.n6254 gnd.n6253 0.152939
R11091 gnd.n6254 gnd.n433 0.152939
R11092 gnd.n6262 gnd.n433 0.152939
R11093 gnd.n6263 gnd.n6262 0.152939
R11094 gnd.n6264 gnd.n6263 0.152939
R11095 gnd.n6264 gnd.n427 0.152939
R11096 gnd.n6272 gnd.n427 0.152939
R11097 gnd.n6273 gnd.n6272 0.152939
R11098 gnd.n6274 gnd.n6273 0.152939
R11099 gnd.n6274 gnd.n421 0.152939
R11100 gnd.n6282 gnd.n421 0.152939
R11101 gnd.n6283 gnd.n6282 0.152939
R11102 gnd.n6284 gnd.n6283 0.152939
R11103 gnd.n6284 gnd.n415 0.152939
R11104 gnd.n6292 gnd.n415 0.152939
R11105 gnd.n6293 gnd.n6292 0.152939
R11106 gnd.n6294 gnd.n6293 0.152939
R11107 gnd.n6294 gnd.n409 0.152939
R11108 gnd.n6302 gnd.n409 0.152939
R11109 gnd.n6303 gnd.n6302 0.152939
R11110 gnd.n6304 gnd.n6303 0.152939
R11111 gnd.n6304 gnd.n403 0.152939
R11112 gnd.n6312 gnd.n403 0.152939
R11113 gnd.n6313 gnd.n6312 0.152939
R11114 gnd.n6314 gnd.n6313 0.152939
R11115 gnd.n6314 gnd.n397 0.152939
R11116 gnd.n6322 gnd.n397 0.152939
R11117 gnd.n6323 gnd.n6322 0.152939
R11118 gnd.n6324 gnd.n6323 0.152939
R11119 gnd.n6324 gnd.n391 0.152939
R11120 gnd.n6332 gnd.n391 0.152939
R11121 gnd.n6333 gnd.n6332 0.152939
R11122 gnd.n6335 gnd.n6333 0.152939
R11123 gnd.n6335 gnd.n6334 0.152939
R11124 gnd.n6334 gnd.n385 0.152939
R11125 gnd.n6344 gnd.n385 0.152939
R11126 gnd.n6345 gnd.n380 0.152939
R11127 gnd.n6353 gnd.n380 0.152939
R11128 gnd.n6354 gnd.n6353 0.152939
R11129 gnd.n6355 gnd.n6354 0.152939
R11130 gnd.n6355 gnd.n374 0.152939
R11131 gnd.n6363 gnd.n374 0.152939
R11132 gnd.n6364 gnd.n6363 0.152939
R11133 gnd.n6365 gnd.n6364 0.152939
R11134 gnd.n6365 gnd.n368 0.152939
R11135 gnd.n6373 gnd.n368 0.152939
R11136 gnd.n6374 gnd.n6373 0.152939
R11137 gnd.n6375 gnd.n6374 0.152939
R11138 gnd.n6375 gnd.n362 0.152939
R11139 gnd.n6383 gnd.n362 0.152939
R11140 gnd.n6384 gnd.n6383 0.152939
R11141 gnd.n6385 gnd.n6384 0.152939
R11142 gnd.n6385 gnd.n356 0.152939
R11143 gnd.n6393 gnd.n356 0.152939
R11144 gnd.n6394 gnd.n6393 0.152939
R11145 gnd.n6395 gnd.n6394 0.152939
R11146 gnd.n6395 gnd.n350 0.152939
R11147 gnd.n6403 gnd.n350 0.152939
R11148 gnd.n6404 gnd.n6403 0.152939
R11149 gnd.n6405 gnd.n6404 0.152939
R11150 gnd.n6405 gnd.n344 0.152939
R11151 gnd.n6413 gnd.n344 0.152939
R11152 gnd.n6414 gnd.n6413 0.152939
R11153 gnd.n6415 gnd.n6414 0.152939
R11154 gnd.n6415 gnd.n338 0.152939
R11155 gnd.n6423 gnd.n338 0.152939
R11156 gnd.n6424 gnd.n6423 0.152939
R11157 gnd.n6425 gnd.n6424 0.152939
R11158 gnd.n6425 gnd.n332 0.152939
R11159 gnd.n6433 gnd.n332 0.152939
R11160 gnd.n6434 gnd.n6433 0.152939
R11161 gnd.n6435 gnd.n6434 0.152939
R11162 gnd.n6435 gnd.n326 0.152939
R11163 gnd.n6443 gnd.n326 0.152939
R11164 gnd.n6444 gnd.n6443 0.152939
R11165 gnd.n6445 gnd.n6444 0.152939
R11166 gnd.n6445 gnd.n320 0.152939
R11167 gnd.n6453 gnd.n320 0.152939
R11168 gnd.n6454 gnd.n6453 0.152939
R11169 gnd.n6455 gnd.n6454 0.152939
R11170 gnd.n6455 gnd.n314 0.152939
R11171 gnd.n6463 gnd.n314 0.152939
R11172 gnd.n6464 gnd.n6463 0.152939
R11173 gnd.n6465 gnd.n6464 0.152939
R11174 gnd.n6465 gnd.n308 0.152939
R11175 gnd.n6473 gnd.n308 0.152939
R11176 gnd.n6474 gnd.n6473 0.152939
R11177 gnd.n6475 gnd.n6474 0.152939
R11178 gnd.n6475 gnd.n302 0.152939
R11179 gnd.n6483 gnd.n302 0.152939
R11180 gnd.n6484 gnd.n6483 0.152939
R11181 gnd.n6485 gnd.n6484 0.152939
R11182 gnd.n6485 gnd.n296 0.152939
R11183 gnd.n6493 gnd.n296 0.152939
R11184 gnd.n6494 gnd.n6493 0.152939
R11185 gnd.n6495 gnd.n6494 0.152939
R11186 gnd.n6495 gnd.n290 0.152939
R11187 gnd.n6503 gnd.n290 0.152939
R11188 gnd.n6504 gnd.n6503 0.152939
R11189 gnd.n6505 gnd.n6504 0.152939
R11190 gnd.n6505 gnd.n284 0.152939
R11191 gnd.n6513 gnd.n284 0.152939
R11192 gnd.n6514 gnd.n6513 0.152939
R11193 gnd.n6515 gnd.n6514 0.152939
R11194 gnd.n6515 gnd.n278 0.152939
R11195 gnd.n6523 gnd.n278 0.152939
R11196 gnd.n6524 gnd.n6523 0.152939
R11197 gnd.n6525 gnd.n6524 0.152939
R11198 gnd.n6525 gnd.n272 0.152939
R11199 gnd.n6533 gnd.n272 0.152939
R11200 gnd.n6534 gnd.n6533 0.152939
R11201 gnd.n6535 gnd.n6534 0.152939
R11202 gnd.n6535 gnd.n266 0.152939
R11203 gnd.n6543 gnd.n266 0.152939
R11204 gnd.n6544 gnd.n6543 0.152939
R11205 gnd.n6545 gnd.n6544 0.152939
R11206 gnd.n6545 gnd.n260 0.152939
R11207 gnd.n6554 gnd.n260 0.152939
R11208 gnd.n6555 gnd.n6554 0.152939
R11209 gnd.n6557 gnd.n6555 0.152939
R11210 gnd.n6599 gnd.n6598 0.152939
R11211 gnd.n6600 gnd.n6599 0.152939
R11212 gnd.n6600 gnd.n198 0.152939
R11213 gnd.n6614 gnd.n198 0.152939
R11214 gnd.n6615 gnd.n6614 0.152939
R11215 gnd.n6616 gnd.n6615 0.152939
R11216 gnd.n6616 gnd.n182 0.152939
R11217 gnd.n6630 gnd.n182 0.152939
R11218 gnd.n6631 gnd.n6630 0.152939
R11219 gnd.n6632 gnd.n6631 0.152939
R11220 gnd.n6632 gnd.n166 0.152939
R11221 gnd.n6720 gnd.n166 0.152939
R11222 gnd.n6721 gnd.n6720 0.152939
R11223 gnd.n6722 gnd.n6721 0.152939
R11224 gnd.n6722 gnd.n88 0.152939
R11225 gnd.n6802 gnd.n88 0.152939
R11226 gnd.n6801 gnd.n89 0.152939
R11227 gnd.n91 gnd.n89 0.152939
R11228 gnd.n95 gnd.n91 0.152939
R11229 gnd.n96 gnd.n95 0.152939
R11230 gnd.n97 gnd.n96 0.152939
R11231 gnd.n98 gnd.n97 0.152939
R11232 gnd.n102 gnd.n98 0.152939
R11233 gnd.n103 gnd.n102 0.152939
R11234 gnd.n104 gnd.n103 0.152939
R11235 gnd.n105 gnd.n104 0.152939
R11236 gnd.n109 gnd.n105 0.152939
R11237 gnd.n110 gnd.n109 0.152939
R11238 gnd.n111 gnd.n110 0.152939
R11239 gnd.n112 gnd.n111 0.152939
R11240 gnd.n116 gnd.n112 0.152939
R11241 gnd.n117 gnd.n116 0.152939
R11242 gnd.n118 gnd.n117 0.152939
R11243 gnd.n119 gnd.n118 0.152939
R11244 gnd.n123 gnd.n119 0.152939
R11245 gnd.n124 gnd.n123 0.152939
R11246 gnd.n125 gnd.n124 0.152939
R11247 gnd.n126 gnd.n125 0.152939
R11248 gnd.n130 gnd.n126 0.152939
R11249 gnd.n131 gnd.n130 0.152939
R11250 gnd.n132 gnd.n131 0.152939
R11251 gnd.n133 gnd.n132 0.152939
R11252 gnd.n137 gnd.n133 0.152939
R11253 gnd.n138 gnd.n137 0.152939
R11254 gnd.n139 gnd.n138 0.152939
R11255 gnd.n140 gnd.n139 0.152939
R11256 gnd.n144 gnd.n140 0.152939
R11257 gnd.n145 gnd.n144 0.152939
R11258 gnd.n146 gnd.n145 0.152939
R11259 gnd.n147 gnd.n146 0.152939
R11260 gnd.n151 gnd.n147 0.152939
R11261 gnd.n152 gnd.n151 0.152939
R11262 gnd.n6732 gnd.n152 0.152939
R11263 gnd.n6732 gnd.n6731 0.152939
R11264 gnd.n3811 gnd.n3810 0.152939
R11265 gnd.n3811 gnd.n1329 0.152939
R11266 gnd.n3826 gnd.n1329 0.152939
R11267 gnd.n3827 gnd.n3826 0.152939
R11268 gnd.n3828 gnd.n3827 0.152939
R11269 gnd.n3829 gnd.n3828 0.152939
R11270 gnd.n3830 gnd.n3829 0.152939
R11271 gnd.n3831 gnd.n3830 0.152939
R11272 gnd.n3832 gnd.n3831 0.152939
R11273 gnd.n3833 gnd.n3832 0.152939
R11274 gnd.n3834 gnd.n3833 0.152939
R11275 gnd.n3835 gnd.n3834 0.152939
R11276 gnd.n3836 gnd.n3835 0.152939
R11277 gnd.n3837 gnd.n3836 0.152939
R11278 gnd.n3838 gnd.n3837 0.152939
R11279 gnd.n3839 gnd.n3838 0.152939
R11280 gnd.n3840 gnd.n3839 0.152939
R11281 gnd.n3841 gnd.n3840 0.152939
R11282 gnd.n3842 gnd.n3841 0.152939
R11283 gnd.n3843 gnd.n3842 0.152939
R11284 gnd.n3843 gnd.n240 0.152939
R11285 gnd.n3844 gnd.n240 0.152939
R11286 gnd.n3845 gnd.n3844 0.152939
R11287 gnd.n3846 gnd.n3845 0.152939
R11288 gnd.n3847 gnd.n3846 0.152939
R11289 gnd.n3848 gnd.n3847 0.152939
R11290 gnd.n3849 gnd.n3848 0.152939
R11291 gnd.n3850 gnd.n3849 0.152939
R11292 gnd.n3851 gnd.n3850 0.152939
R11293 gnd.n3852 gnd.n3851 0.152939
R11294 gnd.n3853 gnd.n3852 0.152939
R11295 gnd.n3854 gnd.n3853 0.152939
R11296 gnd.n3855 gnd.n3854 0.152939
R11297 gnd.n3856 gnd.n3855 0.152939
R11298 gnd.n3857 gnd.n3856 0.152939
R11299 gnd.n3858 gnd.n3857 0.152939
R11300 gnd.n3859 gnd.n3858 0.152939
R11301 gnd.n3860 gnd.n3859 0.152939
R11302 gnd.n3862 gnd.n3860 0.152939
R11303 gnd.n3862 gnd.n3861 0.152939
R11304 gnd.n3861 gnd.n158 0.152939
R11305 gnd.n6730 gnd.n158 0.152939
R11306 gnd.n3715 gnd.n3714 0.152939
R11307 gnd.n3715 gnd.n3711 0.152939
R11308 gnd.n3723 gnd.n3711 0.152939
R11309 gnd.n3724 gnd.n3723 0.152939
R11310 gnd.n3725 gnd.n3724 0.152939
R11311 gnd.n3725 gnd.n3707 0.152939
R11312 gnd.n3733 gnd.n3707 0.152939
R11313 gnd.n3734 gnd.n3733 0.152939
R11314 gnd.n3735 gnd.n3734 0.152939
R11315 gnd.n3735 gnd.n3703 0.152939
R11316 gnd.n3743 gnd.n3703 0.152939
R11317 gnd.n3744 gnd.n3743 0.152939
R11318 gnd.n3746 gnd.n3744 0.152939
R11319 gnd.n3746 gnd.n3745 0.152939
R11320 gnd.n3745 gnd.n1359 0.152939
R11321 gnd.n3759 gnd.n3758 0.152939
R11322 gnd.n3759 gnd.n1355 0.152939
R11323 gnd.n3767 gnd.n1355 0.152939
R11324 gnd.n3768 gnd.n3767 0.152939
R11325 gnd.n3769 gnd.n3768 0.152939
R11326 gnd.n3769 gnd.n1351 0.152939
R11327 gnd.n3777 gnd.n1351 0.152939
R11328 gnd.n3778 gnd.n3777 0.152939
R11329 gnd.n3779 gnd.n3778 0.152939
R11330 gnd.n3779 gnd.n1347 0.152939
R11331 gnd.n3787 gnd.n1347 0.152939
R11332 gnd.n3788 gnd.n3787 0.152939
R11333 gnd.n3789 gnd.n3788 0.152939
R11334 gnd.n3789 gnd.n1343 0.152939
R11335 gnd.n3797 gnd.n1343 0.152939
R11336 gnd.n3798 gnd.n3797 0.152939
R11337 gnd.n3800 gnd.n3798 0.152939
R11338 gnd.n3800 gnd.n3799 0.152939
R11339 gnd.n3799 gnd.n1336 0.152939
R11340 gnd.n3809 gnd.n1336 0.152939
R11341 gnd.n1220 gnd.n1219 0.152939
R11342 gnd.n1221 gnd.n1220 0.152939
R11343 gnd.n1324 gnd.n1221 0.152939
R11344 gnd.n3937 gnd.n1324 0.152939
R11345 gnd.n3938 gnd.n3937 0.152939
R11346 gnd.n3939 gnd.n3938 0.152939
R11347 gnd.n3940 gnd.n3939 0.152939
R11348 gnd.n3940 gnd.n1296 0.152939
R11349 gnd.n3968 gnd.n1296 0.152939
R11350 gnd.n3969 gnd.n3968 0.152939
R11351 gnd.n3970 gnd.n3969 0.152939
R11352 gnd.n3972 gnd.n3970 0.152939
R11353 gnd.n3972 gnd.n3971 0.152939
R11354 gnd.n3971 gnd.n1268 0.152939
R11355 gnd.n1268 gnd.n212 0.152939
R11356 gnd.n6598 gnd.n212 0.152939
R11357 gnd.n3998 gnd.n3992 0.152939
R11358 gnd.n3998 gnd.n3997 0.152939
R11359 gnd.n3997 gnd.n3996 0.152939
R11360 gnd.n3996 gnd.n254 0.152939
R11361 gnd.n256 gnd.n255 0.152939
R11362 gnd.n6556 gnd.n256 0.152939
R11363 gnd.n2057 gnd.n2055 0.152939
R11364 gnd.n2057 gnd.n2056 0.152939
R11365 gnd.n2056 gnd.n2018 0.152939
R11366 gnd.n2306 gnd.n2018 0.152939
R11367 gnd.n2307 gnd.n2306 0.152939
R11368 gnd.n2308 gnd.n2307 0.152939
R11369 gnd.n2308 gnd.n2014 0.152939
R11370 gnd.n2314 gnd.n2014 0.152939
R11371 gnd.n2315 gnd.n2314 0.152939
R11372 gnd.n2316 gnd.n2315 0.152939
R11373 gnd.n2317 gnd.n2316 0.152939
R11374 gnd.n2318 gnd.n2317 0.152939
R11375 gnd.n2321 gnd.n2318 0.152939
R11376 gnd.n2322 gnd.n2321 0.152939
R11377 gnd.n2323 gnd.n2322 0.152939
R11378 gnd.n2324 gnd.n2323 0.152939
R11379 gnd.n2327 gnd.n2324 0.152939
R11380 gnd.n2328 gnd.n2327 0.152939
R11381 gnd.n2329 gnd.n2328 0.152939
R11382 gnd.n2330 gnd.n2329 0.152939
R11383 gnd.n2335 gnd.n2330 0.152939
R11384 gnd.n2336 gnd.n2335 0.152939
R11385 gnd.n2337 gnd.n2336 0.152939
R11386 gnd.n2337 gnd.n1840 0.152939
R11387 gnd.n2689 gnd.n1840 0.152939
R11388 gnd.n2690 gnd.n2689 0.152939
R11389 gnd.n2691 gnd.n2690 0.152939
R11390 gnd.n2691 gnd.n1827 0.152939
R11391 gnd.n2709 gnd.n1827 0.152939
R11392 gnd.n2710 gnd.n2709 0.152939
R11393 gnd.n2711 gnd.n2710 0.152939
R11394 gnd.n2711 gnd.n1814 0.152939
R11395 gnd.n2730 gnd.n1814 0.152939
R11396 gnd.n2731 gnd.n2730 0.152939
R11397 gnd.n2732 gnd.n2731 0.152939
R11398 gnd.n2733 gnd.n2732 0.152939
R11399 gnd.n2733 gnd.n1737 0.152939
R11400 gnd.n2807 gnd.n1737 0.152939
R11401 gnd.n2808 gnd.n2807 0.152939
R11402 gnd.n2809 gnd.n2808 0.152939
R11403 gnd.n2810 gnd.n2809 0.152939
R11404 gnd.n2810 gnd.n1709 0.152939
R11405 gnd.n2844 gnd.n1709 0.152939
R11406 gnd.n2845 gnd.n2844 0.152939
R11407 gnd.n2846 gnd.n2845 0.152939
R11408 gnd.n2846 gnd.n1687 0.152939
R11409 gnd.n2871 gnd.n1687 0.152939
R11410 gnd.n2872 gnd.n2871 0.152939
R11411 gnd.n2873 gnd.n2872 0.152939
R11412 gnd.n2874 gnd.n2873 0.152939
R11413 gnd.n2874 gnd.n1654 0.152939
R11414 gnd.n2913 gnd.n1654 0.152939
R11415 gnd.n2914 gnd.n2913 0.152939
R11416 gnd.n2915 gnd.n2914 0.152939
R11417 gnd.n2916 gnd.n2915 0.152939
R11418 gnd.n2917 gnd.n2916 0.152939
R11419 gnd.n2918 gnd.n2917 0.152939
R11420 gnd.n2918 gnd.n1620 0.152939
R11421 gnd.n2996 gnd.n1620 0.152939
R11422 gnd.n2997 gnd.n2996 0.152939
R11423 gnd.n2998 gnd.n2997 0.152939
R11424 gnd.n2998 gnd.n1597 0.152939
R11425 gnd.n3039 gnd.n1597 0.152939
R11426 gnd.n3040 gnd.n3039 0.152939
R11427 gnd.n3041 gnd.n3040 0.152939
R11428 gnd.n3041 gnd.n1581 0.152939
R11429 gnd.n3083 gnd.n1581 0.152939
R11430 gnd.n3084 gnd.n3083 0.152939
R11431 gnd.n3085 gnd.n3084 0.152939
R11432 gnd.n3086 gnd.n3085 0.152939
R11433 gnd.n3086 gnd.n1550 0.152939
R11434 gnd.n3129 gnd.n1550 0.152939
R11435 gnd.n3130 gnd.n3129 0.152939
R11436 gnd.n3131 gnd.n3130 0.152939
R11437 gnd.n3131 gnd.n1533 0.152939
R11438 gnd.n3190 gnd.n1533 0.152939
R11439 gnd.n3191 gnd.n3190 0.152939
R11440 gnd.n3192 gnd.n3191 0.152939
R11441 gnd.n3192 gnd.n1511 0.152939
R11442 gnd.n3218 gnd.n1511 0.152939
R11443 gnd.n3219 gnd.n3218 0.152939
R11444 gnd.n3220 gnd.n3219 0.152939
R11445 gnd.n3221 gnd.n3220 0.152939
R11446 gnd.n3221 gnd.n1483 0.152939
R11447 gnd.n3262 gnd.n1483 0.152939
R11448 gnd.n3263 gnd.n3262 0.152939
R11449 gnd.n3264 gnd.n3263 0.152939
R11450 gnd.n3265 gnd.n3264 0.152939
R11451 gnd.n3267 gnd.n3265 0.152939
R11452 gnd.n3267 gnd.n3266 0.152939
R11453 gnd.n3266 gnd.n1415 0.152939
R11454 gnd.n1416 gnd.n1415 0.152939
R11455 gnd.n1417 gnd.n1416 0.152939
R11456 gnd.n1424 gnd.n1417 0.152939
R11457 gnd.n1425 gnd.n1424 0.152939
R11458 gnd.n1426 gnd.n1425 0.152939
R11459 gnd.n1427 gnd.n1426 0.152939
R11460 gnd.n1435 gnd.n1427 0.152939
R11461 gnd.n1436 gnd.n1435 0.152939
R11462 gnd.n1437 gnd.n1436 0.152939
R11463 gnd.n1438 gnd.n1437 0.152939
R11464 gnd.n3495 gnd.n1438 0.152939
R11465 gnd.n3496 gnd.n3495 0.152939
R11466 gnd.n3498 gnd.n3496 0.152939
R11467 gnd.n3498 gnd.n3497 0.152939
R11468 gnd.n3497 gnd.n1198 0.152939
R11469 gnd.n1199 gnd.n1198 0.152939
R11470 gnd.n1200 gnd.n1199 0.152939
R11471 gnd.n1206 gnd.n1200 0.152939
R11472 gnd.n1207 gnd.n1206 0.152939
R11473 gnd.n1208 gnd.n1207 0.152939
R11474 gnd.n1209 gnd.n1208 0.152939
R11475 gnd.n3920 gnd.n1209 0.152939
R11476 gnd.n3921 gnd.n3920 0.152939
R11477 gnd.n3926 gnd.n3921 0.152939
R11478 gnd.n3927 gnd.n3926 0.152939
R11479 gnd.n3928 gnd.n3927 0.152939
R11480 gnd.n3929 gnd.n3928 0.152939
R11481 gnd.n3929 gnd.n1306 0.152939
R11482 gnd.n3957 gnd.n1306 0.152939
R11483 gnd.n3958 gnd.n3957 0.152939
R11484 gnd.n3959 gnd.n3958 0.152939
R11485 gnd.n3960 gnd.n3959 0.152939
R11486 gnd.n3960 gnd.n1278 0.152939
R11487 gnd.n3989 gnd.n1278 0.152939
R11488 gnd.n3990 gnd.n3989 0.152939
R11489 gnd.n3991 gnd.n3990 0.152939
R11490 gnd.n3992 gnd.n3991 0.152939
R11491 gnd.n2111 gnd.n2109 0.152939
R11492 gnd.n2109 gnd.n2083 0.152939
R11493 gnd.n2170 gnd.n2083 0.152939
R11494 gnd.n2171 gnd.n2170 0.152939
R11495 gnd.n2172 gnd.n2171 0.152939
R11496 gnd.n2172 gnd.n2080 0.152939
R11497 gnd.n2177 gnd.n2080 0.152939
R11498 gnd.n2178 gnd.n2177 0.152939
R11499 gnd.n2179 gnd.n2178 0.152939
R11500 gnd.n2179 gnd.n2077 0.152939
R11501 gnd.n2184 gnd.n2077 0.152939
R11502 gnd.n2185 gnd.n2184 0.152939
R11503 gnd.n2186 gnd.n2185 0.152939
R11504 gnd.n2186 gnd.n2074 0.152939
R11505 gnd.n2191 gnd.n2074 0.152939
R11506 gnd.n2192 gnd.n2191 0.152939
R11507 gnd.n2193 gnd.n2192 0.152939
R11508 gnd.n2193 gnd.n2072 0.152939
R11509 gnd.n2239 gnd.n2072 0.152939
R11510 gnd.n2240 gnd.n2239 0.152939
R11511 gnd.n2150 gnd.n2090 0.152939
R11512 gnd.n2091 gnd.n2090 0.152939
R11513 gnd.n2092 gnd.n2091 0.152939
R11514 gnd.n2093 gnd.n2092 0.152939
R11515 gnd.n2094 gnd.n2093 0.152939
R11516 gnd.n2095 gnd.n2094 0.152939
R11517 gnd.n2096 gnd.n2095 0.152939
R11518 gnd.n2097 gnd.n2096 0.152939
R11519 gnd.n2098 gnd.n2097 0.152939
R11520 gnd.n2099 gnd.n2098 0.152939
R11521 gnd.n2100 gnd.n2099 0.152939
R11522 gnd.n2101 gnd.n2100 0.152939
R11523 gnd.n2102 gnd.n2101 0.152939
R11524 gnd.n2103 gnd.n2102 0.152939
R11525 gnd.n2104 gnd.n2103 0.152939
R11526 gnd.n2115 gnd.n2104 0.152939
R11527 gnd.n2115 gnd.n2114 0.152939
R11528 gnd.n2114 gnd.n2113 0.152939
R11529 gnd.n2156 gnd.n2151 0.152939
R11530 gnd.n2156 gnd.n2155 0.152939
R11531 gnd.n2155 gnd.n2154 0.152939
R11532 gnd.n2154 gnd.n2152 0.152939
R11533 gnd.n2152 gnd.n902 0.152939
R11534 gnd.n903 gnd.n902 0.152939
R11535 gnd.n904 gnd.n903 0.152939
R11536 gnd.n920 gnd.n904 0.152939
R11537 gnd.n921 gnd.n920 0.152939
R11538 gnd.n922 gnd.n921 0.152939
R11539 gnd.n923 gnd.n922 0.152939
R11540 gnd.n941 gnd.n923 0.152939
R11541 gnd.n942 gnd.n941 0.152939
R11542 gnd.n943 gnd.n942 0.152939
R11543 gnd.n944 gnd.n943 0.152939
R11544 gnd.n964 gnd.n944 0.152939
R11545 gnd.n965 gnd.n964 0.152939
R11546 gnd.n966 gnd.n965 0.152939
R11547 gnd.n967 gnd.n966 0.152939
R11548 gnd.n968 gnd.n967 0.152939
R11549 gnd.n2068 gnd.n968 0.152939
R11550 gnd.n2068 gnd.n982 0.152939
R11551 gnd.n983 gnd.n982 0.152939
R11552 gnd.n984 gnd.n983 0.152939
R11553 gnd.n1000 gnd.n984 0.152939
R11554 gnd.n1001 gnd.n1000 0.152939
R11555 gnd.n1002 gnd.n1001 0.152939
R11556 gnd.n1003 gnd.n1002 0.152939
R11557 gnd.n1020 gnd.n1003 0.152939
R11558 gnd.n1021 gnd.n1020 0.152939
R11559 gnd.n1022 gnd.n1021 0.152939
R11560 gnd.n1023 gnd.n1022 0.152939
R11561 gnd.n1042 gnd.n1023 0.152939
R11562 gnd.n1043 gnd.n1042 0.152939
R11563 gnd.n1044 gnd.n1043 0.152939
R11564 gnd.n1045 gnd.n1044 0.152939
R11565 gnd.n1063 gnd.n1045 0.152939
R11566 gnd.n1064 gnd.n1063 0.152939
R11567 gnd.n1065 gnd.n1064 0.152939
R11568 gnd.n1066 gnd.n1065 0.152939
R11569 gnd.n1084 gnd.n1066 0.152939
R11570 gnd.n4198 gnd.n1084 0.152939
R11571 gnd.n1010 gnd.n953 0.152939
R11572 gnd.n1011 gnd.n1010 0.152939
R11573 gnd.n1012 gnd.n1011 0.152939
R11574 gnd.n1013 gnd.n1012 0.152939
R11575 gnd.n1031 gnd.n1013 0.152939
R11576 gnd.n1032 gnd.n1031 0.152939
R11577 gnd.n1033 gnd.n1032 0.152939
R11578 gnd.n1034 gnd.n1033 0.152939
R11579 gnd.n1052 gnd.n1034 0.152939
R11580 gnd.n1053 gnd.n1052 0.152939
R11581 gnd.n1054 gnd.n1053 0.152939
R11582 gnd.n1055 gnd.n1054 0.152939
R11583 gnd.n1074 gnd.n1055 0.152939
R11584 gnd.n1075 gnd.n1074 0.152939
R11585 gnd.n1076 gnd.n1075 0.152939
R11586 gnd.n1077 gnd.n1076 0.152939
R11587 gnd.n1958 gnd.n1957 0.152939
R11588 gnd.n1959 gnd.n1958 0.152939
R11589 gnd.n1960 gnd.n1959 0.152939
R11590 gnd.n1961 gnd.n1960 0.152939
R11591 gnd.n1962 gnd.n1961 0.152939
R11592 gnd.n1963 gnd.n1962 0.152939
R11593 gnd.n1964 gnd.n1963 0.152939
R11594 gnd.n1965 gnd.n1964 0.152939
R11595 gnd.n1966 gnd.n1965 0.152939
R11596 gnd.n1967 gnd.n1966 0.152939
R11597 gnd.n1968 gnd.n1967 0.152939
R11598 gnd.n1969 gnd.n1968 0.152939
R11599 gnd.n1970 gnd.n1969 0.152939
R11600 gnd.n1971 gnd.n1970 0.152939
R11601 gnd.n1972 gnd.n1971 0.152939
R11602 gnd.n2465 gnd.n2464 0.152939
R11603 gnd.n2464 gnd.n1977 0.152939
R11604 gnd.n1978 gnd.n1977 0.152939
R11605 gnd.n1979 gnd.n1978 0.152939
R11606 gnd.n1980 gnd.n1979 0.152939
R11607 gnd.n1981 gnd.n1980 0.152939
R11608 gnd.n1982 gnd.n1981 0.152939
R11609 gnd.n1983 gnd.n1982 0.152939
R11610 gnd.n1984 gnd.n1983 0.152939
R11611 gnd.n1985 gnd.n1984 0.152939
R11612 gnd.n1986 gnd.n1985 0.152939
R11613 gnd.n1987 gnd.n1986 0.152939
R11614 gnd.n1988 gnd.n1987 0.152939
R11615 gnd.n1989 gnd.n1988 0.152939
R11616 gnd.n1990 gnd.n1989 0.152939
R11617 gnd.n1991 gnd.n1990 0.152939
R11618 gnd.n1992 gnd.n1991 0.152939
R11619 gnd.n1993 gnd.n1992 0.152939
R11620 gnd.n2424 gnd.n1993 0.152939
R11621 gnd.n2424 gnd.n2423 0.152939
R11622 gnd.n4324 gnd.n877 0.152939
R11623 gnd.n4324 gnd.n4323 0.152939
R11624 gnd.n4323 gnd.n4322 0.152939
R11625 gnd.n4322 gnd.n880 0.152939
R11626 gnd.n2204 gnd.n880 0.152939
R11627 gnd.n2204 gnd.n2203 0.152939
R11628 gnd.n2209 gnd.n2203 0.152939
R11629 gnd.n2210 gnd.n2209 0.152939
R11630 gnd.n2211 gnd.n2210 0.152939
R11631 gnd.n2211 gnd.n2200 0.152939
R11632 gnd.n2216 gnd.n2200 0.152939
R11633 gnd.n2217 gnd.n2216 0.152939
R11634 gnd.n2218 gnd.n2217 0.152939
R11635 gnd.n2218 gnd.n2197 0.152939
R11636 gnd.n2223 gnd.n2197 0.152939
R11637 gnd.n2224 gnd.n2223 0.152939
R11638 gnd.n2225 gnd.n2224 0.152939
R11639 gnd.n2226 gnd.n2225 0.152939
R11640 gnd.n2227 gnd.n2226 0.152939
R11641 gnd.n2227 gnd.n2069 0.152939
R11642 gnd.n2247 gnd.n2069 0.152939
R11643 gnd.n2248 gnd.n2247 0.152939
R11644 gnd.n2250 gnd.n2248 0.152939
R11645 gnd.n2250 gnd.n2249 0.152939
R11646 gnd.n2249 gnd.n2035 0.152939
R11647 gnd.n2035 gnd.n2033 0.152939
R11648 gnd.n2266 gnd.n2033 0.152939
R11649 gnd.n2267 gnd.n2266 0.152939
R11650 gnd.n2268 gnd.n2267 0.152939
R11651 gnd.n2268 gnd.n2031 0.152939
R11652 gnd.n2277 gnd.n2031 0.152939
R11653 gnd.n2278 gnd.n2277 0.152939
R11654 gnd.n2279 gnd.n2278 0.152939
R11655 gnd.n2280 gnd.n2279 0.152939
R11656 gnd.n2281 gnd.n2280 0.152939
R11657 gnd.n2281 gnd.n2005 0.152939
R11658 gnd.n2372 gnd.n2005 0.152939
R11659 gnd.n2373 gnd.n2372 0.152939
R11660 gnd.n2375 gnd.n2373 0.152939
R11661 gnd.n2375 gnd.n2374 0.152939
R11662 gnd.n2374 gnd.n1998 0.152939
R11663 gnd.n2422 gnd.n1998 0.152939
R11664 gnd.n835 gnd.n834 0.152939
R11665 gnd.n836 gnd.n835 0.152939
R11666 gnd.n837 gnd.n836 0.152939
R11667 gnd.n838 gnd.n837 0.152939
R11668 gnd.n839 gnd.n838 0.152939
R11669 gnd.n840 gnd.n839 0.152939
R11670 gnd.n841 gnd.n840 0.152939
R11671 gnd.n842 gnd.n841 0.152939
R11672 gnd.n843 gnd.n842 0.152939
R11673 gnd.n844 gnd.n843 0.152939
R11674 gnd.n845 gnd.n844 0.152939
R11675 gnd.n846 gnd.n845 0.152939
R11676 gnd.n847 gnd.n846 0.152939
R11677 gnd.n848 gnd.n847 0.152939
R11678 gnd.n849 gnd.n848 0.152939
R11679 gnd.n850 gnd.n849 0.152939
R11680 gnd.n851 gnd.n850 0.152939
R11681 gnd.n854 gnd.n851 0.152939
R11682 gnd.n855 gnd.n854 0.152939
R11683 gnd.n856 gnd.n855 0.152939
R11684 gnd.n857 gnd.n856 0.152939
R11685 gnd.n858 gnd.n857 0.152939
R11686 gnd.n859 gnd.n858 0.152939
R11687 gnd.n860 gnd.n859 0.152939
R11688 gnd.n861 gnd.n860 0.152939
R11689 gnd.n862 gnd.n861 0.152939
R11690 gnd.n863 gnd.n862 0.152939
R11691 gnd.n864 gnd.n863 0.152939
R11692 gnd.n865 gnd.n864 0.152939
R11693 gnd.n866 gnd.n865 0.152939
R11694 gnd.n867 gnd.n866 0.152939
R11695 gnd.n868 gnd.n867 0.152939
R11696 gnd.n869 gnd.n868 0.152939
R11697 gnd.n870 gnd.n869 0.152939
R11698 gnd.n871 gnd.n870 0.152939
R11699 gnd.n4332 gnd.n871 0.152939
R11700 gnd.n4332 gnd.n4331 0.152939
R11701 gnd.n4331 gnd.n4330 0.152939
R11702 gnd.n2162 gnd.n2160 0.152939
R11703 gnd.n2162 gnd.n2161 0.152939
R11704 gnd.n2161 gnd.n891 0.152939
R11705 gnd.n892 gnd.n891 0.152939
R11706 gnd.n893 gnd.n892 0.152939
R11707 gnd.n911 gnd.n893 0.152939
R11708 gnd.n912 gnd.n911 0.152939
R11709 gnd.n913 gnd.n912 0.152939
R11710 gnd.n914 gnd.n913 0.152939
R11711 gnd.n930 gnd.n914 0.152939
R11712 gnd.n931 gnd.n930 0.152939
R11713 gnd.n932 gnd.n931 0.152939
R11714 gnd.n933 gnd.n932 0.152939
R11715 gnd.n951 gnd.n933 0.152939
R11716 gnd.n952 gnd.n951 0.152939
R11717 gnd.n953 gnd.n952 0.152939
R11718 gnd.n2049 gnd.n2043 0.152939
R11719 gnd.n2050 gnd.n2049 0.152939
R11720 gnd.n2053 gnd.n2052 0.152939
R11721 gnd.n2054 gnd.n2053 0.152939
R11722 gnd.n2055 gnd.n2054 0.152939
R11723 gnd.n600 gnd.n595 0.152939
R11724 gnd.n601 gnd.n600 0.152939
R11725 gnd.n602 gnd.n601 0.152939
R11726 gnd.n607 gnd.n602 0.152939
R11727 gnd.n608 gnd.n607 0.152939
R11728 gnd.n609 gnd.n608 0.152939
R11729 gnd.n610 gnd.n609 0.152939
R11730 gnd.n615 gnd.n610 0.152939
R11731 gnd.n616 gnd.n615 0.152939
R11732 gnd.n617 gnd.n616 0.152939
R11733 gnd.n618 gnd.n617 0.152939
R11734 gnd.n623 gnd.n618 0.152939
R11735 gnd.n624 gnd.n623 0.152939
R11736 gnd.n625 gnd.n624 0.152939
R11737 gnd.n626 gnd.n625 0.152939
R11738 gnd.n631 gnd.n626 0.152939
R11739 gnd.n632 gnd.n631 0.152939
R11740 gnd.n633 gnd.n632 0.152939
R11741 gnd.n634 gnd.n633 0.152939
R11742 gnd.n639 gnd.n634 0.152939
R11743 gnd.n640 gnd.n639 0.152939
R11744 gnd.n641 gnd.n640 0.152939
R11745 gnd.n642 gnd.n641 0.152939
R11746 gnd.n647 gnd.n642 0.152939
R11747 gnd.n648 gnd.n647 0.152939
R11748 gnd.n649 gnd.n648 0.152939
R11749 gnd.n650 gnd.n649 0.152939
R11750 gnd.n655 gnd.n650 0.152939
R11751 gnd.n656 gnd.n655 0.152939
R11752 gnd.n657 gnd.n656 0.152939
R11753 gnd.n658 gnd.n657 0.152939
R11754 gnd.n663 gnd.n658 0.152939
R11755 gnd.n664 gnd.n663 0.152939
R11756 gnd.n665 gnd.n664 0.152939
R11757 gnd.n666 gnd.n665 0.152939
R11758 gnd.n671 gnd.n666 0.152939
R11759 gnd.n672 gnd.n671 0.152939
R11760 gnd.n673 gnd.n672 0.152939
R11761 gnd.n674 gnd.n673 0.152939
R11762 gnd.n679 gnd.n674 0.152939
R11763 gnd.n680 gnd.n679 0.152939
R11764 gnd.n681 gnd.n680 0.152939
R11765 gnd.n682 gnd.n681 0.152939
R11766 gnd.n687 gnd.n682 0.152939
R11767 gnd.n688 gnd.n687 0.152939
R11768 gnd.n689 gnd.n688 0.152939
R11769 gnd.n690 gnd.n689 0.152939
R11770 gnd.n695 gnd.n690 0.152939
R11771 gnd.n696 gnd.n695 0.152939
R11772 gnd.n697 gnd.n696 0.152939
R11773 gnd.n698 gnd.n697 0.152939
R11774 gnd.n703 gnd.n698 0.152939
R11775 gnd.n704 gnd.n703 0.152939
R11776 gnd.n705 gnd.n704 0.152939
R11777 gnd.n706 gnd.n705 0.152939
R11778 gnd.n711 gnd.n706 0.152939
R11779 gnd.n712 gnd.n711 0.152939
R11780 gnd.n713 gnd.n712 0.152939
R11781 gnd.n714 gnd.n713 0.152939
R11782 gnd.n719 gnd.n714 0.152939
R11783 gnd.n720 gnd.n719 0.152939
R11784 gnd.n721 gnd.n720 0.152939
R11785 gnd.n722 gnd.n721 0.152939
R11786 gnd.n727 gnd.n722 0.152939
R11787 gnd.n728 gnd.n727 0.152939
R11788 gnd.n729 gnd.n728 0.152939
R11789 gnd.n730 gnd.n729 0.152939
R11790 gnd.n735 gnd.n730 0.152939
R11791 gnd.n736 gnd.n735 0.152939
R11792 gnd.n737 gnd.n736 0.152939
R11793 gnd.n738 gnd.n737 0.152939
R11794 gnd.n743 gnd.n738 0.152939
R11795 gnd.n744 gnd.n743 0.152939
R11796 gnd.n745 gnd.n744 0.152939
R11797 gnd.n746 gnd.n745 0.152939
R11798 gnd.n751 gnd.n746 0.152939
R11799 gnd.n752 gnd.n751 0.152939
R11800 gnd.n753 gnd.n752 0.152939
R11801 gnd.n754 gnd.n753 0.152939
R11802 gnd.n759 gnd.n754 0.152939
R11803 gnd.n760 gnd.n759 0.152939
R11804 gnd.n761 gnd.n760 0.152939
R11805 gnd.n762 gnd.n761 0.152939
R11806 gnd.n2042 gnd.n762 0.152939
R11807 gnd.n3465 gnd.n3321 0.152939
R11808 gnd.n3466 gnd.n3465 0.152939
R11809 gnd.n3467 gnd.n3466 0.152939
R11810 gnd.n3467 gnd.n3317 0.152939
R11811 gnd.n3478 gnd.n3317 0.152939
R11812 gnd.n3479 gnd.n3478 0.152939
R11813 gnd.n3480 gnd.n3479 0.152939
R11814 gnd.n3480 gnd.n3313 0.152939
R11815 gnd.n3487 gnd.n3313 0.152939
R11816 gnd.n2681 gnd.n2680 0.152939
R11817 gnd.n2681 gnd.n1833 0.152939
R11818 gnd.n2699 gnd.n1833 0.152939
R11819 gnd.n2700 gnd.n2699 0.152939
R11820 gnd.n2701 gnd.n2700 0.152939
R11821 gnd.n2701 gnd.n1820 0.152939
R11822 gnd.n2719 gnd.n1820 0.152939
R11823 gnd.n2720 gnd.n2719 0.152939
R11824 gnd.n2721 gnd.n2720 0.152939
R11825 gnd.n2721 gnd.n1807 0.152939
R11826 gnd.n2742 gnd.n1807 0.152939
R11827 gnd.n2743 gnd.n2742 0.152939
R11828 gnd.n2747 gnd.n2743 0.152939
R11829 gnd.n2747 gnd.n2746 0.152939
R11830 gnd.n2746 gnd.n2745 0.152939
R11831 gnd.n2745 gnd.n1724 0.152939
R11832 gnd.n2826 gnd.n1724 0.152939
R11833 gnd.n2827 gnd.n2826 0.152939
R11834 gnd.n2829 gnd.n2827 0.152939
R11835 gnd.n2829 gnd.n2828 0.152939
R11836 gnd.n2828 gnd.n1694 0.152939
R11837 gnd.n2862 gnd.n1694 0.152939
R11838 gnd.n2863 gnd.n2862 0.152939
R11839 gnd.n2864 gnd.n2863 0.152939
R11840 gnd.n2864 gnd.n1673 0.152939
R11841 gnd.n2891 gnd.n1673 0.152939
R11842 gnd.n2892 gnd.n2891 0.152939
R11843 gnd.n2897 gnd.n2892 0.152939
R11844 gnd.n2897 gnd.n2896 0.152939
R11845 gnd.n2896 gnd.n2895 0.152939
R11846 gnd.n2895 gnd.n1638 0.152939
R11847 gnd.n2951 gnd.n1638 0.152939
R11848 gnd.n2952 gnd.n2951 0.152939
R11849 gnd.n2954 gnd.n2952 0.152939
R11850 gnd.n2954 gnd.n2953 0.152939
R11851 gnd.n2953 gnd.n1613 0.152939
R11852 gnd.n3005 gnd.n1613 0.152939
R11853 gnd.n3006 gnd.n3005 0.152939
R11854 gnd.n3019 gnd.n3006 0.152939
R11855 gnd.n3019 gnd.n3018 0.152939
R11856 gnd.n3018 gnd.n3017 0.152939
R11857 gnd.n3017 gnd.n3007 0.152939
R11858 gnd.n3013 gnd.n3007 0.152939
R11859 gnd.n3013 gnd.n3012 0.152939
R11860 gnd.n3012 gnd.n1567 0.152939
R11861 gnd.n3101 gnd.n1567 0.152939
R11862 gnd.n3102 gnd.n3101 0.152939
R11863 gnd.n3113 gnd.n3102 0.152939
R11864 gnd.n3113 gnd.n3112 0.152939
R11865 gnd.n3112 gnd.n3111 0.152939
R11866 gnd.n3111 gnd.n3103 0.152939
R11867 gnd.n3107 gnd.n3103 0.152939
R11868 gnd.n3107 gnd.n1527 0.152939
R11869 gnd.n3199 gnd.n1527 0.152939
R11870 gnd.n3200 gnd.n3199 0.152939
R11871 gnd.n3202 gnd.n3200 0.152939
R11872 gnd.n3202 gnd.n3201 0.152939
R11873 gnd.n3201 gnd.n1498 0.152939
R11874 gnd.n3237 gnd.n1498 0.152939
R11875 gnd.n3238 gnd.n3237 0.152939
R11876 gnd.n3247 gnd.n3238 0.152939
R11877 gnd.n3247 gnd.n3246 0.152939
R11878 gnd.n3246 gnd.n3245 0.152939
R11879 gnd.n3245 gnd.n3240 0.152939
R11880 gnd.n3240 gnd.n3239 0.152939
R11881 gnd.n3239 gnd.n1462 0.152939
R11882 gnd.n3293 gnd.n1462 0.152939
R11883 gnd.n3294 gnd.n3293 0.152939
R11884 gnd.n3295 gnd.n3294 0.152939
R11885 gnd.n3295 gnd.n1458 0.152939
R11886 gnd.n3299 gnd.n1458 0.152939
R11887 gnd.n3300 gnd.n3299 0.152939
R11888 gnd.n3301 gnd.n3300 0.152939
R11889 gnd.n3301 gnd.n1454 0.152939
R11890 gnd.n3305 gnd.n1454 0.152939
R11891 gnd.n3306 gnd.n3305 0.152939
R11892 gnd.n3307 gnd.n3306 0.152939
R11893 gnd.n3307 gnd.n1448 0.152939
R11894 gnd.n3311 gnd.n1448 0.152939
R11895 gnd.n3312 gnd.n3311 0.152939
R11896 gnd.n3489 gnd.n3312 0.152939
R11897 gnd.n3489 gnd.n3488 0.152939
R11898 gnd.n2408 gnd.n2383 0.152939
R11899 gnd.n2408 gnd.n2407 0.152939
R11900 gnd.n2407 gnd.n2406 0.152939
R11901 gnd.n2406 gnd.n2389 0.152939
R11902 gnd.n2402 gnd.n2389 0.152939
R11903 gnd.n2402 gnd.n2401 0.152939
R11904 gnd.n2401 gnd.n2396 0.152939
R11905 gnd.n2396 gnd.n1846 0.152939
R11906 gnd.n2679 gnd.n1846 0.152939
R11907 gnd.n2256 gnd.n2037 0.152939
R11908 gnd.n2257 gnd.n2256 0.152939
R11909 gnd.n2258 gnd.n2257 0.152939
R11910 gnd.n2258 gnd.n2025 0.152939
R11911 gnd.n2297 gnd.n2025 0.152939
R11912 gnd.n2297 gnd.n2296 0.152939
R11913 gnd.n2296 gnd.n2295 0.152939
R11914 gnd.n2295 gnd.n2026 0.152939
R11915 gnd.n2291 gnd.n2026 0.152939
R11916 gnd.n2291 gnd.n2290 0.152939
R11917 gnd.n2290 gnd.n2289 0.152939
R11918 gnd.n2289 gnd.n2008 0.152939
R11919 gnd.n2364 gnd.n2008 0.152939
R11920 gnd.n2365 gnd.n2364 0.152939
R11921 gnd.n2366 gnd.n2365 0.152939
R11922 gnd.n2366 gnd.n2002 0.152939
R11923 gnd.n2381 gnd.n2002 0.152939
R11924 gnd.n2382 gnd.n2381 0.152939
R11925 gnd.n2415 gnd.n2382 0.152939
R11926 gnd.n2415 gnd.n2414 0.152939
R11927 gnd.n4195 gnd.n1087 0.152939
R11928 gnd.n4191 gnd.n1087 0.152939
R11929 gnd.n4191 gnd.n4190 0.152939
R11930 gnd.n4190 gnd.n4189 0.152939
R11931 gnd.n4189 gnd.n1092 0.152939
R11932 gnd.n4185 gnd.n1092 0.152939
R11933 gnd.n4185 gnd.n4184 0.152939
R11934 gnd.n4184 gnd.n4183 0.152939
R11935 gnd.n4183 gnd.n1097 0.152939
R11936 gnd.n4179 gnd.n1097 0.152939
R11937 gnd.n4179 gnd.n4178 0.152939
R11938 gnd.n4178 gnd.n4177 0.152939
R11939 gnd.n4177 gnd.n1102 0.152939
R11940 gnd.n4173 gnd.n1102 0.152939
R11941 gnd.n4173 gnd.n4172 0.152939
R11942 gnd.n4172 gnd.n4171 0.152939
R11943 gnd.n4171 gnd.n1107 0.152939
R11944 gnd.n4167 gnd.n1107 0.152939
R11945 gnd.n4167 gnd.n4166 0.152939
R11946 gnd.n4166 gnd.n4165 0.152939
R11947 gnd.n4165 gnd.n1112 0.152939
R11948 gnd.n4161 gnd.n1112 0.152939
R11949 gnd.n4161 gnd.n4160 0.152939
R11950 gnd.n4160 gnd.n4159 0.152939
R11951 gnd.n4159 gnd.n1117 0.152939
R11952 gnd.n4155 gnd.n1117 0.152939
R11953 gnd.n4155 gnd.n4154 0.152939
R11954 gnd.n4154 gnd.n4153 0.152939
R11955 gnd.n4153 gnd.n1122 0.152939
R11956 gnd.n4149 gnd.n1122 0.152939
R11957 gnd.n4149 gnd.n4148 0.152939
R11958 gnd.n4148 gnd.n4147 0.152939
R11959 gnd.n4147 gnd.n1127 0.152939
R11960 gnd.n4143 gnd.n1127 0.152939
R11961 gnd.n4143 gnd.n4142 0.152939
R11962 gnd.n4142 gnd.n4141 0.152939
R11963 gnd.n4141 gnd.n1132 0.152939
R11964 gnd.n4137 gnd.n1132 0.152939
R11965 gnd.n4137 gnd.n4136 0.152939
R11966 gnd.n4136 gnd.n4135 0.152939
R11967 gnd.n4135 gnd.n1137 0.152939
R11968 gnd.n4131 gnd.n1137 0.152939
R11969 gnd.n4131 gnd.n4130 0.152939
R11970 gnd.n4130 gnd.n4129 0.152939
R11971 gnd.n4129 gnd.n1142 0.152939
R11972 gnd.n4125 gnd.n1142 0.152939
R11973 gnd.n4125 gnd.n4124 0.152939
R11974 gnd.n4124 gnd.n4123 0.152939
R11975 gnd.n4123 gnd.n1147 0.152939
R11976 gnd.n4119 gnd.n1147 0.152939
R11977 gnd.n4119 gnd.n4118 0.152939
R11978 gnd.n4118 gnd.n4117 0.152939
R11979 gnd.n4117 gnd.n1152 0.152939
R11980 gnd.n4113 gnd.n1152 0.152939
R11981 gnd.n4113 gnd.n4112 0.152939
R11982 gnd.n4112 gnd.n4111 0.152939
R11983 gnd.n4111 gnd.n1157 0.152939
R11984 gnd.n4107 gnd.n1157 0.152939
R11985 gnd.n4107 gnd.n4106 0.152939
R11986 gnd.n4106 gnd.n4105 0.152939
R11987 gnd.n4105 gnd.n1162 0.152939
R11988 gnd.n4101 gnd.n1162 0.152939
R11989 gnd.n4101 gnd.n4100 0.152939
R11990 gnd.n4100 gnd.n4099 0.152939
R11991 gnd.n4099 gnd.n1167 0.152939
R11992 gnd.n4095 gnd.n1167 0.152939
R11993 gnd.n4095 gnd.n4094 0.152939
R11994 gnd.n4094 gnd.n4093 0.152939
R11995 gnd.n4093 gnd.n1172 0.152939
R11996 gnd.n4089 gnd.n1172 0.152939
R11997 gnd.n4089 gnd.n4088 0.152939
R11998 gnd.n4088 gnd.n4087 0.152939
R11999 gnd.n4087 gnd.n1177 0.152939
R12000 gnd.n4083 gnd.n1177 0.152939
R12001 gnd.n4083 gnd.n4082 0.152939
R12002 gnd.n4082 gnd.n4081 0.152939
R12003 gnd.n4081 gnd.n1182 0.152939
R12004 gnd.n4077 gnd.n1182 0.152939
R12005 gnd.n4077 gnd.n4076 0.152939
R12006 gnd.n4076 gnd.n4075 0.152939
R12007 gnd.n4075 gnd.n1187 0.152939
R12008 gnd.n1190 gnd.n1187 0.152939
R12009 gnd.n3368 gnd.n1232 0.152939
R12010 gnd.n4045 gnd.n1232 0.152939
R12011 gnd.n4045 gnd.n4044 0.152939
R12012 gnd.n4044 gnd.n4043 0.152939
R12013 gnd.n4043 gnd.n1233 0.152939
R12014 gnd.n4039 gnd.n1233 0.152939
R12015 gnd.n4039 gnd.n4038 0.152939
R12016 gnd.n4038 gnd.n4037 0.152939
R12017 gnd.n4037 gnd.n1238 0.152939
R12018 gnd.n4033 gnd.n1238 0.152939
R12019 gnd.n4033 gnd.n4032 0.152939
R12020 gnd.n4032 gnd.n4031 0.152939
R12021 gnd.n4031 gnd.n1243 0.152939
R12022 gnd.n4027 gnd.n1243 0.152939
R12023 gnd.n4027 gnd.n4026 0.152939
R12024 gnd.n4026 gnd.n4025 0.152939
R12025 gnd.n4025 gnd.n1248 0.152939
R12026 gnd.n4021 gnd.n1248 0.152939
R12027 gnd.n4021 gnd.n241 0.152939
R12028 gnd.n6576 gnd.n241 0.152939
R12029 gnd.n6577 gnd.n6576 0.152939
R12030 gnd.n6578 gnd.n6577 0.152939
R12031 gnd.n6578 gnd.n227 0.152939
R12032 gnd.n6590 gnd.n227 0.152939
R12033 gnd.n6591 gnd.n6590 0.152939
R12034 gnd.n6592 gnd.n6591 0.152939
R12035 gnd.n6592 gnd.n206 0.152939
R12036 gnd.n6606 gnd.n206 0.152939
R12037 gnd.n6607 gnd.n6606 0.152939
R12038 gnd.n6608 gnd.n6607 0.152939
R12039 gnd.n6608 gnd.n191 0.152939
R12040 gnd.n6622 gnd.n191 0.152939
R12041 gnd.n6623 gnd.n6622 0.152939
R12042 gnd.n6624 gnd.n6623 0.152939
R12043 gnd.n6624 gnd.n176 0.152939
R12044 gnd.n6638 gnd.n176 0.152939
R12045 gnd.n6639 gnd.n6638 0.152939
R12046 gnd.n6714 gnd.n6639 0.152939
R12047 gnd.n6714 gnd.n6713 0.152939
R12048 gnd.n6713 gnd.n6712 0.152939
R12049 gnd.n6712 gnd.n6640 0.152939
R12050 gnd.n6708 gnd.n6640 0.152939
R12051 gnd.n6707 gnd.n6642 0.152939
R12052 gnd.n6703 gnd.n6642 0.152939
R12053 gnd.n6703 gnd.n6702 0.152939
R12054 gnd.n6702 gnd.n6701 0.152939
R12055 gnd.n6701 gnd.n6648 0.152939
R12056 gnd.n6697 gnd.n6648 0.152939
R12057 gnd.n6697 gnd.n6696 0.152939
R12058 gnd.n6696 gnd.n6695 0.152939
R12059 gnd.n6695 gnd.n6656 0.152939
R12060 gnd.n6691 gnd.n6656 0.152939
R12061 gnd.n6691 gnd.n6690 0.152939
R12062 gnd.n6690 gnd.n6689 0.152939
R12063 gnd.n6689 gnd.n6664 0.152939
R12064 gnd.n6685 gnd.n6664 0.152939
R12065 gnd.n6685 gnd.n6684 0.152939
R12066 gnd.n6684 gnd.n6683 0.152939
R12067 gnd.n6683 gnd.n6672 0.152939
R12068 gnd.n6672 gnd.n78 0.152939
R12069 gnd.n3817 gnd.n1333 0.152939
R12070 gnd.n3818 gnd.n3817 0.152939
R12071 gnd.n3820 gnd.n3818 0.152939
R12072 gnd.n3820 gnd.n3819 0.152939
R12073 gnd.n3819 gnd.n1315 0.152939
R12074 gnd.n3947 gnd.n1315 0.152939
R12075 gnd.n3948 gnd.n3947 0.152939
R12076 gnd.n3950 gnd.n3948 0.152939
R12077 gnd.n3950 gnd.n3949 0.152939
R12078 gnd.n3949 gnd.n1286 0.152939
R12079 gnd.n3979 gnd.n1286 0.152939
R12080 gnd.n3980 gnd.n3979 0.152939
R12081 gnd.n3982 gnd.n3980 0.152939
R12082 gnd.n3982 gnd.n3981 0.152939
R12083 gnd.n3981 gnd.n1257 0.152939
R12084 gnd.n4013 gnd.n1257 0.152939
R12085 gnd.n4014 gnd.n4013 0.152939
R12086 gnd.n4016 gnd.n4014 0.152939
R12087 gnd.n4016 gnd.n4015 0.152939
R12088 gnd.n4015 gnd.n51 0.152939
R12089 gnd.n6839 gnd.n51 0.152939
R12090 gnd.n6839 gnd.n6838 0.152939
R12091 gnd.n6838 gnd.n53 0.152939
R12092 gnd.n6834 gnd.n53 0.152939
R12093 gnd.n6834 gnd.n6833 0.152939
R12094 gnd.n6833 gnd.n6832 0.152939
R12095 gnd.n6832 gnd.n58 0.152939
R12096 gnd.n6828 gnd.n58 0.152939
R12097 gnd.n6828 gnd.n6827 0.152939
R12098 gnd.n6827 gnd.n6826 0.152939
R12099 gnd.n6826 gnd.n63 0.152939
R12100 gnd.n6822 gnd.n63 0.152939
R12101 gnd.n6822 gnd.n6821 0.152939
R12102 gnd.n6821 gnd.n6820 0.152939
R12103 gnd.n6820 gnd.n68 0.152939
R12104 gnd.n6816 gnd.n68 0.152939
R12105 gnd.n6816 gnd.n6815 0.152939
R12106 gnd.n6815 gnd.n6814 0.152939
R12107 gnd.n6814 gnd.n73 0.152939
R12108 gnd.n6810 gnd.n73 0.152939
R12109 gnd.n6810 gnd.n6809 0.152939
R12110 gnd.n6809 gnd.n6808 0.152939
R12111 gnd.n3456 gnd.n3321 0.151415
R12112 gnd.n2413 gnd.n2383 0.151415
R12113 gnd.n2241 gnd.n2240 0.145814
R12114 gnd.n2241 gnd.n2037 0.145814
R12115 gnd.n5023 gnd.n0 0.127478
R12116 gnd.n254 gnd.n213 0.108732
R12117 gnd.n2052 gnd.n2051 0.108732
R12118 gnd.n5024 gnd.n4593 0.0767195
R12119 gnd.n5024 gnd.n4972 0.0767195
R12120 gnd.n4197 gnd.n4196 0.063
R12121 gnd.n3369 gnd.n3366 0.063
R12122 gnd.n5763 gnd.n4442 0.0477147
R12123 gnd.n255 gnd.n213 0.0447073
R12124 gnd.n2051 gnd.n2050 0.0447073
R12125 gnd.n4927 gnd.n4815 0.0442063
R12126 gnd.n4928 gnd.n4927 0.0442063
R12127 gnd.n4929 gnd.n4928 0.0442063
R12128 gnd.n4929 gnd.n4804 0.0442063
R12129 gnd.n4943 gnd.n4804 0.0442063
R12130 gnd.n4944 gnd.n4943 0.0442063
R12131 gnd.n4945 gnd.n4944 0.0442063
R12132 gnd.n4945 gnd.n4791 0.0442063
R12133 gnd.n5063 gnd.n4791 0.0442063
R12134 gnd.n5064 gnd.n5063 0.0442063
R12135 gnd.n5066 gnd.n4725 0.0344674
R12136 gnd.n3457 gnd.n3455 0.0344674
R12137 gnd.n2412 gnd.n1916 0.0344674
R12138 gnd.n5086 gnd.n5085 0.0269946
R12139 gnd.n5088 gnd.n5087 0.0269946
R12140 gnd.n4720 gnd.n4718 0.0269946
R12141 gnd.n5098 gnd.n5096 0.0269946
R12142 gnd.n5097 gnd.n4699 0.0269946
R12143 gnd.n5117 gnd.n5116 0.0269946
R12144 gnd.n5119 gnd.n5118 0.0269946
R12145 gnd.n4694 gnd.n4692 0.0269946
R12146 gnd.n5129 gnd.n5127 0.0269946
R12147 gnd.n5128 gnd.n4675 0.0269946
R12148 gnd.n5148 gnd.n5147 0.0269946
R12149 gnd.n5150 gnd.n5149 0.0269946
R12150 gnd.n4669 gnd.n4667 0.0269946
R12151 gnd.n5160 gnd.n5158 0.0269946
R12152 gnd.n5159 gnd.n4649 0.0269946
R12153 gnd.n5179 gnd.n5178 0.0269946
R12154 gnd.n5181 gnd.n5180 0.0269946
R12155 gnd.n4643 gnd.n4641 0.0269946
R12156 gnd.n5191 gnd.n5189 0.0269946
R12157 gnd.n5190 gnd.n4624 0.0269946
R12158 gnd.n5210 gnd.n5209 0.0269946
R12159 gnd.n5212 gnd.n5211 0.0269946
R12160 gnd.n4618 gnd.n4616 0.0269946
R12161 gnd.n5222 gnd.n5220 0.0269946
R12162 gnd.n5221 gnd.n4600 0.0269946
R12163 gnd.n5240 gnd.n5239 0.0269946
R12164 gnd.n5242 gnd.n5241 0.0269946
R12165 gnd.n4588 gnd.n4587 0.0269946
R12166 gnd.n5276 gnd.n4584 0.0269946
R12167 gnd.n5275 gnd.n4585 0.0269946
R12168 gnd.n5295 gnd.n4567 0.0269946
R12169 gnd.n5297 gnd.n5296 0.0269946
R12170 gnd.n5298 gnd.n4565 0.0269946
R12171 gnd.n5305 gnd.n5301 0.0269946
R12172 gnd.n5304 gnd.n5303 0.0269946
R12173 gnd.n5302 gnd.n4544 0.0269946
R12174 gnd.n5329 gnd.n4545 0.0269946
R12175 gnd.n5328 gnd.n4546 0.0269946
R12176 gnd.n5370 gnd.n4523 0.0269946
R12177 gnd.n5372 gnd.n5371 0.0269946
R12178 gnd.n5381 gnd.n4516 0.0269946
R12179 gnd.n5383 gnd.n5382 0.0269946
R12180 gnd.n5384 gnd.n4512 0.0269946
R12181 gnd.n5672 gnd.n4513 0.0269946
R12182 gnd.n5671 gnd.n4514 0.0269946
R12183 gnd.n5388 gnd.n771 0.0269946
R12184 gnd.n5389 gnd.n772 0.0269946
R12185 gnd.n5391 gnd.n773 0.0269946
R12186 gnd.n5651 gnd.n5650 0.0269946
R12187 gnd.n5652 gnd.n795 0.0269946
R12188 gnd.n5653 gnd.n796 0.0269946
R12189 gnd.n5654 gnd.n797 0.0269946
R12190 gnd.n3366 gnd.n3365 0.0246168
R12191 gnd.n4196 gnd.n1086 0.0246168
R12192 gnd.n5066 gnd.n5065 0.0202011
R12193 gnd.n3365 gnd.n3363 0.0174837
R12194 gnd.n3377 gnd.n3363 0.0174837
R12195 gnd.n3379 gnd.n3377 0.0174837
R12196 gnd.n3379 gnd.n3378 0.0174837
R12197 gnd.n3378 gnd.n3358 0.0174837
R12198 gnd.n3388 gnd.n3358 0.0174837
R12199 gnd.n3388 gnd.n3387 0.0174837
R12200 gnd.n3387 gnd.n3359 0.0174837
R12201 gnd.n3359 gnd.n3354 0.0174837
R12202 gnd.n3396 gnd.n3354 0.0174837
R12203 gnd.n3398 gnd.n3396 0.0174837
R12204 gnd.n3398 gnd.n3397 0.0174837
R12205 gnd.n3397 gnd.n3349 0.0174837
R12206 gnd.n3407 gnd.n3349 0.0174837
R12207 gnd.n3407 gnd.n3406 0.0174837
R12208 gnd.n3406 gnd.n3350 0.0174837
R12209 gnd.n3350 gnd.n3345 0.0174837
R12210 gnd.n3415 gnd.n3345 0.0174837
R12211 gnd.n3417 gnd.n3415 0.0174837
R12212 gnd.n3417 gnd.n3416 0.0174837
R12213 gnd.n3416 gnd.n3340 0.0174837
R12214 gnd.n3426 gnd.n3340 0.0174837
R12215 gnd.n3426 gnd.n3425 0.0174837
R12216 gnd.n3425 gnd.n3341 0.0174837
R12217 gnd.n3341 gnd.n3336 0.0174837
R12218 gnd.n3434 gnd.n3336 0.0174837
R12219 gnd.n3436 gnd.n3434 0.0174837
R12220 gnd.n3436 gnd.n3435 0.0174837
R12221 gnd.n3435 gnd.n3331 0.0174837
R12222 gnd.n3447 gnd.n3331 0.0174837
R12223 gnd.n3447 gnd.n3446 0.0174837
R12224 gnd.n3446 gnd.n3332 0.0174837
R12225 gnd.n3332 gnd.n3325 0.0174837
R12226 gnd.n3454 gnd.n3325 0.0174837
R12227 gnd.n3455 gnd.n3454 0.0174837
R12228 gnd.n1865 gnd.n1086 0.0174837
R12229 gnd.n1867 gnd.n1865 0.0174837
R12230 gnd.n2670 gnd.n1867 0.0174837
R12231 gnd.n2670 gnd.n2669 0.0174837
R12232 gnd.n2669 gnd.n1868 0.0174837
R12233 gnd.n2666 gnd.n1868 0.0174837
R12234 gnd.n2666 gnd.n2665 0.0174837
R12235 gnd.n2665 gnd.n1873 0.0174837
R12236 gnd.n2662 gnd.n1873 0.0174837
R12237 gnd.n2662 gnd.n2661 0.0174837
R12238 gnd.n2661 gnd.n1878 0.0174837
R12239 gnd.n2658 gnd.n1878 0.0174837
R12240 gnd.n2658 gnd.n2657 0.0174837
R12241 gnd.n2657 gnd.n1882 0.0174837
R12242 gnd.n2654 gnd.n1882 0.0174837
R12243 gnd.n2654 gnd.n2653 0.0174837
R12244 gnd.n2653 gnd.n1886 0.0174837
R12245 gnd.n2650 gnd.n1886 0.0174837
R12246 gnd.n2650 gnd.n2649 0.0174837
R12247 gnd.n2649 gnd.n1890 0.0174837
R12248 gnd.n2646 gnd.n1890 0.0174837
R12249 gnd.n2646 gnd.n2645 0.0174837
R12250 gnd.n2645 gnd.n1896 0.0174837
R12251 gnd.n2642 gnd.n1896 0.0174837
R12252 gnd.n2642 gnd.n2641 0.0174837
R12253 gnd.n2641 gnd.n1900 0.0174837
R12254 gnd.n2638 gnd.n1900 0.0174837
R12255 gnd.n2638 gnd.n2637 0.0174837
R12256 gnd.n2637 gnd.n1904 0.0174837
R12257 gnd.n2634 gnd.n1904 0.0174837
R12258 gnd.n2634 gnd.n2633 0.0174837
R12259 gnd.n2633 gnd.n1910 0.0174837
R12260 gnd.n2630 gnd.n1910 0.0174837
R12261 gnd.n2630 gnd.n2629 0.0174837
R12262 gnd.n2629 gnd.n1916 0.0174837
R12263 gnd.n5065 gnd.n5064 0.0148637
R12264 gnd.n5648 gnd.n5392 0.0144266
R12265 gnd.n5649 gnd.n5648 0.0130679
R12266 gnd.n5085 gnd.n4725 0.00797283
R12267 gnd.n5087 gnd.n5086 0.00797283
R12268 gnd.n5088 gnd.n4720 0.00797283
R12269 gnd.n5096 gnd.n4718 0.00797283
R12270 gnd.n5098 gnd.n5097 0.00797283
R12271 gnd.n5116 gnd.n4699 0.00797283
R12272 gnd.n5118 gnd.n5117 0.00797283
R12273 gnd.n5119 gnd.n4694 0.00797283
R12274 gnd.n5127 gnd.n4692 0.00797283
R12275 gnd.n5129 gnd.n5128 0.00797283
R12276 gnd.n5147 gnd.n4675 0.00797283
R12277 gnd.n5149 gnd.n5148 0.00797283
R12278 gnd.n5150 gnd.n4669 0.00797283
R12279 gnd.n5158 gnd.n4667 0.00797283
R12280 gnd.n5160 gnd.n5159 0.00797283
R12281 gnd.n5178 gnd.n4649 0.00797283
R12282 gnd.n5180 gnd.n5179 0.00797283
R12283 gnd.n5181 gnd.n4643 0.00797283
R12284 gnd.n5189 gnd.n4641 0.00797283
R12285 gnd.n5191 gnd.n5190 0.00797283
R12286 gnd.n5209 gnd.n4624 0.00797283
R12287 gnd.n5211 gnd.n5210 0.00797283
R12288 gnd.n5212 gnd.n4618 0.00797283
R12289 gnd.n5220 gnd.n4616 0.00797283
R12290 gnd.n5222 gnd.n5221 0.00797283
R12291 gnd.n5239 gnd.n4600 0.00797283
R12292 gnd.n5241 gnd.n5240 0.00797283
R12293 gnd.n5242 gnd.n4588 0.00797283
R12294 gnd.n4587 gnd.n4584 0.00797283
R12295 gnd.n5276 gnd.n5275 0.00797283
R12296 gnd.n4585 gnd.n4567 0.00797283
R12297 gnd.n5296 gnd.n5295 0.00797283
R12298 gnd.n5298 gnd.n5297 0.00797283
R12299 gnd.n5301 gnd.n4565 0.00797283
R12300 gnd.n5305 gnd.n5304 0.00797283
R12301 gnd.n5303 gnd.n5302 0.00797283
R12302 gnd.n4545 gnd.n4544 0.00797283
R12303 gnd.n5329 gnd.n5328 0.00797283
R12304 gnd.n4546 gnd.n4523 0.00797283
R12305 gnd.n5372 gnd.n5370 0.00797283
R12306 gnd.n5371 gnd.n4516 0.00797283
R12307 gnd.n5382 gnd.n5381 0.00797283
R12308 gnd.n5384 gnd.n5383 0.00797283
R12309 gnd.n4513 gnd.n4512 0.00797283
R12310 gnd.n5672 gnd.n5671 0.00797283
R12311 gnd.n5388 gnd.n4514 0.00797283
R12312 gnd.n5389 gnd.n771 0.00797283
R12313 gnd.n5391 gnd.n772 0.00797283
R12314 gnd.n5392 gnd.n773 0.00797283
R12315 gnd.n5650 gnd.n5649 0.00797283
R12316 gnd.n5652 gnd.n5651 0.00797283
R12317 gnd.n5653 gnd.n795 0.00797283
R12318 gnd.n5654 gnd.n796 0.00797283
R12319 gnd.n4442 gnd.n797 0.00797283
R12320 gnd.n6577 gnd.n240 0.00614909
R12321 gnd.n2247 gnd.n2068 0.00614909
R12322 gnd.n3457 gnd.n3456 0.000839674
R12323 gnd.n2413 gnd.n2412 0.000839674
R12324 commonsourceibias.n25 commonsourceibias.t46 230.006
R12325 commonsourceibias.n91 commonsourceibias.t62 230.006
R12326 commonsourceibias.n154 commonsourceibias.t54 230.006
R12327 commonsourceibias.n258 commonsourceibias.t16 230.006
R12328 commonsourceibias.n217 commonsourceibias.t75 230.006
R12329 commonsourceibias.n355 commonsourceibias.t65 230.006
R12330 commonsourceibias.n70 commonsourceibias.t32 207.983
R12331 commonsourceibias.n136 commonsourceibias.t71 207.983
R12332 commonsourceibias.n199 commonsourceibias.t61 207.983
R12333 commonsourceibias.n304 commonsourceibias.t2 207.983
R12334 commonsourceibias.n338 commonsourceibias.t84 207.983
R12335 commonsourceibias.n401 commonsourceibias.t73 207.983
R12336 commonsourceibias.n10 commonsourceibias.t14 168.701
R12337 commonsourceibias.n63 commonsourceibias.t24 168.701
R12338 commonsourceibias.n57 commonsourceibias.t30 168.701
R12339 commonsourceibias.n16 commonsourceibias.t20 168.701
R12340 commonsourceibias.n49 commonsourceibias.t36 168.701
R12341 commonsourceibias.n43 commonsourceibias.t44 168.701
R12342 commonsourceibias.n19 commonsourceibias.t26 168.701
R12343 commonsourceibias.n21 commonsourceibias.t34 168.701
R12344 commonsourceibias.n23 commonsourceibias.t10 168.701
R12345 commonsourceibias.n26 commonsourceibias.t40 168.701
R12346 commonsourceibias.n1 commonsourceibias.t81 168.701
R12347 commonsourceibias.n129 commonsourceibias.t55 168.701
R12348 commonsourceibias.n123 commonsourceibias.t53 168.701
R12349 commonsourceibias.n7 commonsourceibias.t76 168.701
R12350 commonsourceibias.n115 commonsourceibias.t86 168.701
R12351 commonsourceibias.n109 commonsourceibias.t50 168.701
R12352 commonsourceibias.n85 commonsourceibias.t69 168.701
R12353 commonsourceibias.n87 commonsourceibias.t67 168.701
R12354 commonsourceibias.n89 commonsourceibias.t78 168.701
R12355 commonsourceibias.n92 commonsourceibias.t64 168.701
R12356 commonsourceibias.n155 commonsourceibias.t57 168.701
R12357 commonsourceibias.n152 commonsourceibias.t68 168.701
R12358 commonsourceibias.n150 commonsourceibias.t58 168.701
R12359 commonsourceibias.n148 commonsourceibias.t60 168.701
R12360 commonsourceibias.n172 commonsourceibias.t91 168.701
R12361 commonsourceibias.n178 commonsourceibias.t77 168.701
R12362 commonsourceibias.n145 commonsourceibias.t66 168.701
R12363 commonsourceibias.n186 commonsourceibias.t95 168.701
R12364 commonsourceibias.n192 commonsourceibias.t49 168.701
R12365 commonsourceibias.n139 commonsourceibias.t72 168.701
R12366 commonsourceibias.n259 commonsourceibias.t8 168.701
R12367 commonsourceibias.n256 commonsourceibias.t18 168.701
R12368 commonsourceibias.n254 commonsourceibias.t4 168.701
R12369 commonsourceibias.n252 commonsourceibias.t42 168.701
R12370 commonsourceibias.n276 commonsourceibias.t12 168.701
R12371 commonsourceibias.n282 commonsourceibias.t6 168.701
R12372 commonsourceibias.n284 commonsourceibias.t28 168.701
R12373 commonsourceibias.n291 commonsourceibias.t0 168.701
R12374 commonsourceibias.n297 commonsourceibias.t38 168.701
R12375 commonsourceibias.n244 commonsourceibias.t22 168.701
R12376 commonsourceibias.n203 commonsourceibias.t92 168.701
R12377 commonsourceibias.n331 commonsourceibias.t51 168.701
R12378 commonsourceibias.n325 commonsourceibias.t63 168.701
R12379 commonsourceibias.n318 commonsourceibias.t88 168.701
R12380 commonsourceibias.n316 commonsourceibias.t48 168.701
R12381 commonsourceibias.n218 commonsourceibias.t59 168.701
R12382 commonsourceibias.n215 commonsourceibias.t90 168.701
R12383 commonsourceibias.n213 commonsourceibias.t80 168.701
R12384 commonsourceibias.n211 commonsourceibias.t83 168.701
R12385 commonsourceibias.n235 commonsourceibias.t94 168.701
R12386 commonsourceibias.n356 commonsourceibias.t52 168.701
R12387 commonsourceibias.n353 commonsourceibias.t82 168.701
R12388 commonsourceibias.n351 commonsourceibias.t70 168.701
R12389 commonsourceibias.n349 commonsourceibias.t74 168.701
R12390 commonsourceibias.n373 commonsourceibias.t87 168.701
R12391 commonsourceibias.n379 commonsourceibias.t89 168.701
R12392 commonsourceibias.n381 commonsourceibias.t79 168.701
R12393 commonsourceibias.n388 commonsourceibias.t56 168.701
R12394 commonsourceibias.n394 commonsourceibias.t93 168.701
R12395 commonsourceibias.n341 commonsourceibias.t85 168.701
R12396 commonsourceibias.n27 commonsourceibias.n24 161.3
R12397 commonsourceibias.n29 commonsourceibias.n28 161.3
R12398 commonsourceibias.n31 commonsourceibias.n30 161.3
R12399 commonsourceibias.n32 commonsourceibias.n22 161.3
R12400 commonsourceibias.n34 commonsourceibias.n33 161.3
R12401 commonsourceibias.n36 commonsourceibias.n35 161.3
R12402 commonsourceibias.n37 commonsourceibias.n20 161.3
R12403 commonsourceibias.n39 commonsourceibias.n38 161.3
R12404 commonsourceibias.n41 commonsourceibias.n40 161.3
R12405 commonsourceibias.n42 commonsourceibias.n18 161.3
R12406 commonsourceibias.n45 commonsourceibias.n44 161.3
R12407 commonsourceibias.n46 commonsourceibias.n17 161.3
R12408 commonsourceibias.n48 commonsourceibias.n47 161.3
R12409 commonsourceibias.n50 commonsourceibias.n15 161.3
R12410 commonsourceibias.n52 commonsourceibias.n51 161.3
R12411 commonsourceibias.n53 commonsourceibias.n14 161.3
R12412 commonsourceibias.n55 commonsourceibias.n54 161.3
R12413 commonsourceibias.n56 commonsourceibias.n13 161.3
R12414 commonsourceibias.n59 commonsourceibias.n58 161.3
R12415 commonsourceibias.n60 commonsourceibias.n12 161.3
R12416 commonsourceibias.n62 commonsourceibias.n61 161.3
R12417 commonsourceibias.n64 commonsourceibias.n11 161.3
R12418 commonsourceibias.n66 commonsourceibias.n65 161.3
R12419 commonsourceibias.n68 commonsourceibias.n67 161.3
R12420 commonsourceibias.n69 commonsourceibias.n9 161.3
R12421 commonsourceibias.n93 commonsourceibias.n90 161.3
R12422 commonsourceibias.n95 commonsourceibias.n94 161.3
R12423 commonsourceibias.n97 commonsourceibias.n96 161.3
R12424 commonsourceibias.n98 commonsourceibias.n88 161.3
R12425 commonsourceibias.n100 commonsourceibias.n99 161.3
R12426 commonsourceibias.n102 commonsourceibias.n101 161.3
R12427 commonsourceibias.n103 commonsourceibias.n86 161.3
R12428 commonsourceibias.n105 commonsourceibias.n104 161.3
R12429 commonsourceibias.n107 commonsourceibias.n106 161.3
R12430 commonsourceibias.n108 commonsourceibias.n84 161.3
R12431 commonsourceibias.n111 commonsourceibias.n110 161.3
R12432 commonsourceibias.n112 commonsourceibias.n8 161.3
R12433 commonsourceibias.n114 commonsourceibias.n113 161.3
R12434 commonsourceibias.n116 commonsourceibias.n6 161.3
R12435 commonsourceibias.n118 commonsourceibias.n117 161.3
R12436 commonsourceibias.n119 commonsourceibias.n5 161.3
R12437 commonsourceibias.n121 commonsourceibias.n120 161.3
R12438 commonsourceibias.n122 commonsourceibias.n4 161.3
R12439 commonsourceibias.n125 commonsourceibias.n124 161.3
R12440 commonsourceibias.n126 commonsourceibias.n3 161.3
R12441 commonsourceibias.n128 commonsourceibias.n127 161.3
R12442 commonsourceibias.n130 commonsourceibias.n2 161.3
R12443 commonsourceibias.n132 commonsourceibias.n131 161.3
R12444 commonsourceibias.n134 commonsourceibias.n133 161.3
R12445 commonsourceibias.n135 commonsourceibias.n0 161.3
R12446 commonsourceibias.n198 commonsourceibias.n138 161.3
R12447 commonsourceibias.n197 commonsourceibias.n196 161.3
R12448 commonsourceibias.n195 commonsourceibias.n194 161.3
R12449 commonsourceibias.n193 commonsourceibias.n140 161.3
R12450 commonsourceibias.n191 commonsourceibias.n190 161.3
R12451 commonsourceibias.n189 commonsourceibias.n141 161.3
R12452 commonsourceibias.n188 commonsourceibias.n187 161.3
R12453 commonsourceibias.n185 commonsourceibias.n142 161.3
R12454 commonsourceibias.n184 commonsourceibias.n183 161.3
R12455 commonsourceibias.n182 commonsourceibias.n143 161.3
R12456 commonsourceibias.n181 commonsourceibias.n180 161.3
R12457 commonsourceibias.n179 commonsourceibias.n144 161.3
R12458 commonsourceibias.n177 commonsourceibias.n176 161.3
R12459 commonsourceibias.n175 commonsourceibias.n146 161.3
R12460 commonsourceibias.n174 commonsourceibias.n173 161.3
R12461 commonsourceibias.n171 commonsourceibias.n147 161.3
R12462 commonsourceibias.n170 commonsourceibias.n169 161.3
R12463 commonsourceibias.n168 commonsourceibias.n167 161.3
R12464 commonsourceibias.n166 commonsourceibias.n149 161.3
R12465 commonsourceibias.n165 commonsourceibias.n164 161.3
R12466 commonsourceibias.n163 commonsourceibias.n162 161.3
R12467 commonsourceibias.n161 commonsourceibias.n151 161.3
R12468 commonsourceibias.n160 commonsourceibias.n159 161.3
R12469 commonsourceibias.n158 commonsourceibias.n157 161.3
R12470 commonsourceibias.n156 commonsourceibias.n153 161.3
R12471 commonsourceibias.n303 commonsourceibias.n243 161.3
R12472 commonsourceibias.n302 commonsourceibias.n301 161.3
R12473 commonsourceibias.n300 commonsourceibias.n299 161.3
R12474 commonsourceibias.n298 commonsourceibias.n245 161.3
R12475 commonsourceibias.n296 commonsourceibias.n295 161.3
R12476 commonsourceibias.n294 commonsourceibias.n246 161.3
R12477 commonsourceibias.n293 commonsourceibias.n292 161.3
R12478 commonsourceibias.n290 commonsourceibias.n247 161.3
R12479 commonsourceibias.n289 commonsourceibias.n288 161.3
R12480 commonsourceibias.n287 commonsourceibias.n248 161.3
R12481 commonsourceibias.n286 commonsourceibias.n285 161.3
R12482 commonsourceibias.n283 commonsourceibias.n249 161.3
R12483 commonsourceibias.n281 commonsourceibias.n280 161.3
R12484 commonsourceibias.n279 commonsourceibias.n250 161.3
R12485 commonsourceibias.n278 commonsourceibias.n277 161.3
R12486 commonsourceibias.n275 commonsourceibias.n251 161.3
R12487 commonsourceibias.n274 commonsourceibias.n273 161.3
R12488 commonsourceibias.n272 commonsourceibias.n271 161.3
R12489 commonsourceibias.n270 commonsourceibias.n253 161.3
R12490 commonsourceibias.n269 commonsourceibias.n268 161.3
R12491 commonsourceibias.n267 commonsourceibias.n266 161.3
R12492 commonsourceibias.n265 commonsourceibias.n255 161.3
R12493 commonsourceibias.n264 commonsourceibias.n263 161.3
R12494 commonsourceibias.n262 commonsourceibias.n261 161.3
R12495 commonsourceibias.n260 commonsourceibias.n257 161.3
R12496 commonsourceibias.n237 commonsourceibias.n236 161.3
R12497 commonsourceibias.n234 commonsourceibias.n210 161.3
R12498 commonsourceibias.n233 commonsourceibias.n232 161.3
R12499 commonsourceibias.n231 commonsourceibias.n230 161.3
R12500 commonsourceibias.n229 commonsourceibias.n212 161.3
R12501 commonsourceibias.n228 commonsourceibias.n227 161.3
R12502 commonsourceibias.n226 commonsourceibias.n225 161.3
R12503 commonsourceibias.n224 commonsourceibias.n214 161.3
R12504 commonsourceibias.n223 commonsourceibias.n222 161.3
R12505 commonsourceibias.n221 commonsourceibias.n220 161.3
R12506 commonsourceibias.n219 commonsourceibias.n216 161.3
R12507 commonsourceibias.n313 commonsourceibias.n209 161.3
R12508 commonsourceibias.n337 commonsourceibias.n202 161.3
R12509 commonsourceibias.n336 commonsourceibias.n335 161.3
R12510 commonsourceibias.n334 commonsourceibias.n333 161.3
R12511 commonsourceibias.n332 commonsourceibias.n204 161.3
R12512 commonsourceibias.n330 commonsourceibias.n329 161.3
R12513 commonsourceibias.n328 commonsourceibias.n205 161.3
R12514 commonsourceibias.n327 commonsourceibias.n326 161.3
R12515 commonsourceibias.n324 commonsourceibias.n206 161.3
R12516 commonsourceibias.n323 commonsourceibias.n322 161.3
R12517 commonsourceibias.n321 commonsourceibias.n207 161.3
R12518 commonsourceibias.n320 commonsourceibias.n319 161.3
R12519 commonsourceibias.n317 commonsourceibias.n208 161.3
R12520 commonsourceibias.n315 commonsourceibias.n314 161.3
R12521 commonsourceibias.n400 commonsourceibias.n340 161.3
R12522 commonsourceibias.n399 commonsourceibias.n398 161.3
R12523 commonsourceibias.n397 commonsourceibias.n396 161.3
R12524 commonsourceibias.n395 commonsourceibias.n342 161.3
R12525 commonsourceibias.n393 commonsourceibias.n392 161.3
R12526 commonsourceibias.n391 commonsourceibias.n343 161.3
R12527 commonsourceibias.n390 commonsourceibias.n389 161.3
R12528 commonsourceibias.n387 commonsourceibias.n344 161.3
R12529 commonsourceibias.n386 commonsourceibias.n385 161.3
R12530 commonsourceibias.n384 commonsourceibias.n345 161.3
R12531 commonsourceibias.n383 commonsourceibias.n382 161.3
R12532 commonsourceibias.n380 commonsourceibias.n346 161.3
R12533 commonsourceibias.n378 commonsourceibias.n377 161.3
R12534 commonsourceibias.n376 commonsourceibias.n347 161.3
R12535 commonsourceibias.n375 commonsourceibias.n374 161.3
R12536 commonsourceibias.n372 commonsourceibias.n348 161.3
R12537 commonsourceibias.n371 commonsourceibias.n370 161.3
R12538 commonsourceibias.n369 commonsourceibias.n368 161.3
R12539 commonsourceibias.n367 commonsourceibias.n350 161.3
R12540 commonsourceibias.n366 commonsourceibias.n365 161.3
R12541 commonsourceibias.n364 commonsourceibias.n363 161.3
R12542 commonsourceibias.n362 commonsourceibias.n352 161.3
R12543 commonsourceibias.n361 commonsourceibias.n360 161.3
R12544 commonsourceibias.n359 commonsourceibias.n358 161.3
R12545 commonsourceibias.n357 commonsourceibias.n354 161.3
R12546 commonsourceibias.n80 commonsourceibias.n78 81.5057
R12547 commonsourceibias.n240 commonsourceibias.n238 81.5057
R12548 commonsourceibias.n80 commonsourceibias.n79 80.9324
R12549 commonsourceibias.n82 commonsourceibias.n81 80.9324
R12550 commonsourceibias.n77 commonsourceibias.n76 80.9324
R12551 commonsourceibias.n75 commonsourceibias.n74 80.9324
R12552 commonsourceibias.n73 commonsourceibias.n72 80.9324
R12553 commonsourceibias.n307 commonsourceibias.n306 80.9324
R12554 commonsourceibias.n309 commonsourceibias.n308 80.9324
R12555 commonsourceibias.n311 commonsourceibias.n310 80.9324
R12556 commonsourceibias.n242 commonsourceibias.n241 80.9324
R12557 commonsourceibias.n240 commonsourceibias.n239 80.9324
R12558 commonsourceibias.n71 commonsourceibias.n70 80.6037
R12559 commonsourceibias.n137 commonsourceibias.n136 80.6037
R12560 commonsourceibias.n200 commonsourceibias.n199 80.6037
R12561 commonsourceibias.n305 commonsourceibias.n304 80.6037
R12562 commonsourceibias.n339 commonsourceibias.n338 80.6037
R12563 commonsourceibias.n402 commonsourceibias.n401 80.6037
R12564 commonsourceibias.n65 commonsourceibias.n64 56.5617
R12565 commonsourceibias.n51 commonsourceibias.n50 56.5617
R12566 commonsourceibias.n42 commonsourceibias.n41 56.5617
R12567 commonsourceibias.n28 commonsourceibias.n27 56.5617
R12568 commonsourceibias.n131 commonsourceibias.n130 56.5617
R12569 commonsourceibias.n117 commonsourceibias.n116 56.5617
R12570 commonsourceibias.n108 commonsourceibias.n107 56.5617
R12571 commonsourceibias.n94 commonsourceibias.n93 56.5617
R12572 commonsourceibias.n157 commonsourceibias.n156 56.5617
R12573 commonsourceibias.n171 commonsourceibias.n170 56.5617
R12574 commonsourceibias.n180 commonsourceibias.n179 56.5617
R12575 commonsourceibias.n194 commonsourceibias.n193 56.5617
R12576 commonsourceibias.n261 commonsourceibias.n260 56.5617
R12577 commonsourceibias.n275 commonsourceibias.n274 56.5617
R12578 commonsourceibias.n285 commonsourceibias.n283 56.5617
R12579 commonsourceibias.n299 commonsourceibias.n298 56.5617
R12580 commonsourceibias.n333 commonsourceibias.n332 56.5617
R12581 commonsourceibias.n319 commonsourceibias.n317 56.5617
R12582 commonsourceibias.n220 commonsourceibias.n219 56.5617
R12583 commonsourceibias.n234 commonsourceibias.n233 56.5617
R12584 commonsourceibias.n358 commonsourceibias.n357 56.5617
R12585 commonsourceibias.n372 commonsourceibias.n371 56.5617
R12586 commonsourceibias.n382 commonsourceibias.n380 56.5617
R12587 commonsourceibias.n396 commonsourceibias.n395 56.5617
R12588 commonsourceibias.n56 commonsourceibias.n55 56.0773
R12589 commonsourceibias.n37 commonsourceibias.n36 56.0773
R12590 commonsourceibias.n122 commonsourceibias.n121 56.0773
R12591 commonsourceibias.n103 commonsourceibias.n102 56.0773
R12592 commonsourceibias.n166 commonsourceibias.n165 56.0773
R12593 commonsourceibias.n185 commonsourceibias.n184 56.0773
R12594 commonsourceibias.n270 commonsourceibias.n269 56.0773
R12595 commonsourceibias.n290 commonsourceibias.n289 56.0773
R12596 commonsourceibias.n324 commonsourceibias.n323 56.0773
R12597 commonsourceibias.n229 commonsourceibias.n228 56.0773
R12598 commonsourceibias.n367 commonsourceibias.n366 56.0773
R12599 commonsourceibias.n387 commonsourceibias.n386 56.0773
R12600 commonsourceibias.n70 commonsourceibias.n69 46.0096
R12601 commonsourceibias.n136 commonsourceibias.n135 46.0096
R12602 commonsourceibias.n199 commonsourceibias.n198 46.0096
R12603 commonsourceibias.n304 commonsourceibias.n303 46.0096
R12604 commonsourceibias.n338 commonsourceibias.n337 46.0096
R12605 commonsourceibias.n401 commonsourceibias.n400 46.0096
R12606 commonsourceibias.n58 commonsourceibias.n12 41.5458
R12607 commonsourceibias.n33 commonsourceibias.n32 41.5458
R12608 commonsourceibias.n124 commonsourceibias.n3 41.5458
R12609 commonsourceibias.n99 commonsourceibias.n98 41.5458
R12610 commonsourceibias.n162 commonsourceibias.n161 41.5458
R12611 commonsourceibias.n187 commonsourceibias.n141 41.5458
R12612 commonsourceibias.n266 commonsourceibias.n265 41.5458
R12613 commonsourceibias.n292 commonsourceibias.n246 41.5458
R12614 commonsourceibias.n326 commonsourceibias.n205 41.5458
R12615 commonsourceibias.n225 commonsourceibias.n224 41.5458
R12616 commonsourceibias.n363 commonsourceibias.n362 41.5458
R12617 commonsourceibias.n389 commonsourceibias.n343 41.5458
R12618 commonsourceibias.n48 commonsourceibias.n17 40.577
R12619 commonsourceibias.n44 commonsourceibias.n17 40.577
R12620 commonsourceibias.n114 commonsourceibias.n8 40.577
R12621 commonsourceibias.n110 commonsourceibias.n8 40.577
R12622 commonsourceibias.n173 commonsourceibias.n146 40.577
R12623 commonsourceibias.n177 commonsourceibias.n146 40.577
R12624 commonsourceibias.n277 commonsourceibias.n250 40.577
R12625 commonsourceibias.n281 commonsourceibias.n250 40.577
R12626 commonsourceibias.n315 commonsourceibias.n209 40.577
R12627 commonsourceibias.n236 commonsourceibias.n209 40.577
R12628 commonsourceibias.n374 commonsourceibias.n347 40.577
R12629 commonsourceibias.n378 commonsourceibias.n347 40.577
R12630 commonsourceibias.n62 commonsourceibias.n12 39.6083
R12631 commonsourceibias.n32 commonsourceibias.n31 39.6083
R12632 commonsourceibias.n128 commonsourceibias.n3 39.6083
R12633 commonsourceibias.n98 commonsourceibias.n97 39.6083
R12634 commonsourceibias.n161 commonsourceibias.n160 39.6083
R12635 commonsourceibias.n191 commonsourceibias.n141 39.6083
R12636 commonsourceibias.n265 commonsourceibias.n264 39.6083
R12637 commonsourceibias.n296 commonsourceibias.n246 39.6083
R12638 commonsourceibias.n330 commonsourceibias.n205 39.6083
R12639 commonsourceibias.n224 commonsourceibias.n223 39.6083
R12640 commonsourceibias.n362 commonsourceibias.n361 39.6083
R12641 commonsourceibias.n393 commonsourceibias.n343 39.6083
R12642 commonsourceibias.n26 commonsourceibias.n25 33.0515
R12643 commonsourceibias.n92 commonsourceibias.n91 33.0515
R12644 commonsourceibias.n155 commonsourceibias.n154 33.0515
R12645 commonsourceibias.n259 commonsourceibias.n258 33.0515
R12646 commonsourceibias.n218 commonsourceibias.n217 33.0515
R12647 commonsourceibias.n356 commonsourceibias.n355 33.0515
R12648 commonsourceibias.n25 commonsourceibias.n24 28.5514
R12649 commonsourceibias.n91 commonsourceibias.n90 28.5514
R12650 commonsourceibias.n154 commonsourceibias.n153 28.5514
R12651 commonsourceibias.n258 commonsourceibias.n257 28.5514
R12652 commonsourceibias.n217 commonsourceibias.n216 28.5514
R12653 commonsourceibias.n355 commonsourceibias.n354 28.5514
R12654 commonsourceibias.n69 commonsourceibias.n68 26.0455
R12655 commonsourceibias.n135 commonsourceibias.n134 26.0455
R12656 commonsourceibias.n198 commonsourceibias.n197 26.0455
R12657 commonsourceibias.n303 commonsourceibias.n302 26.0455
R12658 commonsourceibias.n337 commonsourceibias.n336 26.0455
R12659 commonsourceibias.n400 commonsourceibias.n399 26.0455
R12660 commonsourceibias.n55 commonsourceibias.n14 25.0767
R12661 commonsourceibias.n38 commonsourceibias.n37 25.0767
R12662 commonsourceibias.n121 commonsourceibias.n5 25.0767
R12663 commonsourceibias.n104 commonsourceibias.n103 25.0767
R12664 commonsourceibias.n167 commonsourceibias.n166 25.0767
R12665 commonsourceibias.n184 commonsourceibias.n143 25.0767
R12666 commonsourceibias.n271 commonsourceibias.n270 25.0767
R12667 commonsourceibias.n289 commonsourceibias.n248 25.0767
R12668 commonsourceibias.n323 commonsourceibias.n207 25.0767
R12669 commonsourceibias.n230 commonsourceibias.n229 25.0767
R12670 commonsourceibias.n368 commonsourceibias.n367 25.0767
R12671 commonsourceibias.n386 commonsourceibias.n345 25.0767
R12672 commonsourceibias.n51 commonsourceibias.n16 24.3464
R12673 commonsourceibias.n41 commonsourceibias.n19 24.3464
R12674 commonsourceibias.n117 commonsourceibias.n7 24.3464
R12675 commonsourceibias.n107 commonsourceibias.n85 24.3464
R12676 commonsourceibias.n170 commonsourceibias.n148 24.3464
R12677 commonsourceibias.n180 commonsourceibias.n145 24.3464
R12678 commonsourceibias.n274 commonsourceibias.n252 24.3464
R12679 commonsourceibias.n285 commonsourceibias.n284 24.3464
R12680 commonsourceibias.n319 commonsourceibias.n318 24.3464
R12681 commonsourceibias.n233 commonsourceibias.n211 24.3464
R12682 commonsourceibias.n371 commonsourceibias.n349 24.3464
R12683 commonsourceibias.n382 commonsourceibias.n381 24.3464
R12684 commonsourceibias.n65 commonsourceibias.n10 23.8546
R12685 commonsourceibias.n27 commonsourceibias.n26 23.8546
R12686 commonsourceibias.n131 commonsourceibias.n1 23.8546
R12687 commonsourceibias.n93 commonsourceibias.n92 23.8546
R12688 commonsourceibias.n156 commonsourceibias.n155 23.8546
R12689 commonsourceibias.n194 commonsourceibias.n139 23.8546
R12690 commonsourceibias.n260 commonsourceibias.n259 23.8546
R12691 commonsourceibias.n299 commonsourceibias.n244 23.8546
R12692 commonsourceibias.n333 commonsourceibias.n203 23.8546
R12693 commonsourceibias.n219 commonsourceibias.n218 23.8546
R12694 commonsourceibias.n357 commonsourceibias.n356 23.8546
R12695 commonsourceibias.n396 commonsourceibias.n341 23.8546
R12696 commonsourceibias.n64 commonsourceibias.n63 16.9689
R12697 commonsourceibias.n28 commonsourceibias.n23 16.9689
R12698 commonsourceibias.n130 commonsourceibias.n129 16.9689
R12699 commonsourceibias.n94 commonsourceibias.n89 16.9689
R12700 commonsourceibias.n157 commonsourceibias.n152 16.9689
R12701 commonsourceibias.n193 commonsourceibias.n192 16.9689
R12702 commonsourceibias.n261 commonsourceibias.n256 16.9689
R12703 commonsourceibias.n298 commonsourceibias.n297 16.9689
R12704 commonsourceibias.n332 commonsourceibias.n331 16.9689
R12705 commonsourceibias.n220 commonsourceibias.n215 16.9689
R12706 commonsourceibias.n358 commonsourceibias.n353 16.9689
R12707 commonsourceibias.n395 commonsourceibias.n394 16.9689
R12708 commonsourceibias.n50 commonsourceibias.n49 16.477
R12709 commonsourceibias.n43 commonsourceibias.n42 16.477
R12710 commonsourceibias.n116 commonsourceibias.n115 16.477
R12711 commonsourceibias.n109 commonsourceibias.n108 16.477
R12712 commonsourceibias.n172 commonsourceibias.n171 16.477
R12713 commonsourceibias.n179 commonsourceibias.n178 16.477
R12714 commonsourceibias.n276 commonsourceibias.n275 16.477
R12715 commonsourceibias.n283 commonsourceibias.n282 16.477
R12716 commonsourceibias.n317 commonsourceibias.n316 16.477
R12717 commonsourceibias.n235 commonsourceibias.n234 16.477
R12718 commonsourceibias.n373 commonsourceibias.n372 16.477
R12719 commonsourceibias.n380 commonsourceibias.n379 16.477
R12720 commonsourceibias.n57 commonsourceibias.n56 15.9852
R12721 commonsourceibias.n36 commonsourceibias.n21 15.9852
R12722 commonsourceibias.n123 commonsourceibias.n122 15.9852
R12723 commonsourceibias.n102 commonsourceibias.n87 15.9852
R12724 commonsourceibias.n165 commonsourceibias.n150 15.9852
R12725 commonsourceibias.n186 commonsourceibias.n185 15.9852
R12726 commonsourceibias.n269 commonsourceibias.n254 15.9852
R12727 commonsourceibias.n291 commonsourceibias.n290 15.9852
R12728 commonsourceibias.n325 commonsourceibias.n324 15.9852
R12729 commonsourceibias.n228 commonsourceibias.n213 15.9852
R12730 commonsourceibias.n366 commonsourceibias.n351 15.9852
R12731 commonsourceibias.n388 commonsourceibias.n387 15.9852
R12732 commonsourceibias.n73 commonsourceibias.n71 13.2057
R12733 commonsourceibias.n307 commonsourceibias.n305 13.2057
R12734 commonsourceibias.n404 commonsourceibias.n201 11.9876
R12735 commonsourceibias.n404 commonsourceibias.n403 10.3347
R12736 commonsourceibias.n112 commonsourceibias.n83 9.50363
R12737 commonsourceibias.n313 commonsourceibias.n312 9.50363
R12738 commonsourceibias.n201 commonsourceibias.n137 8.732
R12739 commonsourceibias.n403 commonsourceibias.n339 8.732
R12740 commonsourceibias.n58 commonsourceibias.n57 8.60764
R12741 commonsourceibias.n33 commonsourceibias.n21 8.60764
R12742 commonsourceibias.n124 commonsourceibias.n123 8.60764
R12743 commonsourceibias.n99 commonsourceibias.n87 8.60764
R12744 commonsourceibias.n162 commonsourceibias.n150 8.60764
R12745 commonsourceibias.n187 commonsourceibias.n186 8.60764
R12746 commonsourceibias.n266 commonsourceibias.n254 8.60764
R12747 commonsourceibias.n292 commonsourceibias.n291 8.60764
R12748 commonsourceibias.n326 commonsourceibias.n325 8.60764
R12749 commonsourceibias.n225 commonsourceibias.n213 8.60764
R12750 commonsourceibias.n363 commonsourceibias.n351 8.60764
R12751 commonsourceibias.n389 commonsourceibias.n388 8.60764
R12752 commonsourceibias.n49 commonsourceibias.n48 8.11581
R12753 commonsourceibias.n44 commonsourceibias.n43 8.11581
R12754 commonsourceibias.n115 commonsourceibias.n114 8.11581
R12755 commonsourceibias.n110 commonsourceibias.n109 8.11581
R12756 commonsourceibias.n173 commonsourceibias.n172 8.11581
R12757 commonsourceibias.n178 commonsourceibias.n177 8.11581
R12758 commonsourceibias.n277 commonsourceibias.n276 8.11581
R12759 commonsourceibias.n282 commonsourceibias.n281 8.11581
R12760 commonsourceibias.n316 commonsourceibias.n315 8.11581
R12761 commonsourceibias.n236 commonsourceibias.n235 8.11581
R12762 commonsourceibias.n374 commonsourceibias.n373 8.11581
R12763 commonsourceibias.n379 commonsourceibias.n378 8.11581
R12764 commonsourceibias.n63 commonsourceibias.n62 7.62397
R12765 commonsourceibias.n31 commonsourceibias.n23 7.62397
R12766 commonsourceibias.n129 commonsourceibias.n128 7.62397
R12767 commonsourceibias.n97 commonsourceibias.n89 7.62397
R12768 commonsourceibias.n160 commonsourceibias.n152 7.62397
R12769 commonsourceibias.n192 commonsourceibias.n191 7.62397
R12770 commonsourceibias.n264 commonsourceibias.n256 7.62397
R12771 commonsourceibias.n297 commonsourceibias.n296 7.62397
R12772 commonsourceibias.n331 commonsourceibias.n330 7.62397
R12773 commonsourceibias.n223 commonsourceibias.n215 7.62397
R12774 commonsourceibias.n361 commonsourceibias.n353 7.62397
R12775 commonsourceibias.n394 commonsourceibias.n393 7.62397
R12776 commonsourceibias.n201 commonsourceibias.n200 5.00473
R12777 commonsourceibias.n403 commonsourceibias.n402 5.00473
R12778 commonsourceibias commonsourceibias.n404 3.87639
R12779 commonsourceibias.n78 commonsourceibias.t41 2.82907
R12780 commonsourceibias.n78 commonsourceibias.t47 2.82907
R12781 commonsourceibias.n79 commonsourceibias.t35 2.82907
R12782 commonsourceibias.n79 commonsourceibias.t11 2.82907
R12783 commonsourceibias.n81 commonsourceibias.t45 2.82907
R12784 commonsourceibias.n81 commonsourceibias.t27 2.82907
R12785 commonsourceibias.n76 commonsourceibias.t21 2.82907
R12786 commonsourceibias.n76 commonsourceibias.t37 2.82907
R12787 commonsourceibias.n74 commonsourceibias.t25 2.82907
R12788 commonsourceibias.n74 commonsourceibias.t31 2.82907
R12789 commonsourceibias.n72 commonsourceibias.t33 2.82907
R12790 commonsourceibias.n72 commonsourceibias.t15 2.82907
R12791 commonsourceibias.n306 commonsourceibias.t23 2.82907
R12792 commonsourceibias.n306 commonsourceibias.t3 2.82907
R12793 commonsourceibias.n308 commonsourceibias.t1 2.82907
R12794 commonsourceibias.n308 commonsourceibias.t39 2.82907
R12795 commonsourceibias.n310 commonsourceibias.t7 2.82907
R12796 commonsourceibias.n310 commonsourceibias.t29 2.82907
R12797 commonsourceibias.n241 commonsourceibias.t43 2.82907
R12798 commonsourceibias.n241 commonsourceibias.t13 2.82907
R12799 commonsourceibias.n239 commonsourceibias.t19 2.82907
R12800 commonsourceibias.n239 commonsourceibias.t5 2.82907
R12801 commonsourceibias.n238 commonsourceibias.t17 2.82907
R12802 commonsourceibias.n238 commonsourceibias.t9 2.82907
R12803 commonsourceibias.n68 commonsourceibias.n10 0.738255
R12804 commonsourceibias.n134 commonsourceibias.n1 0.738255
R12805 commonsourceibias.n197 commonsourceibias.n139 0.738255
R12806 commonsourceibias.n302 commonsourceibias.n244 0.738255
R12807 commonsourceibias.n336 commonsourceibias.n203 0.738255
R12808 commonsourceibias.n399 commonsourceibias.n341 0.738255
R12809 commonsourceibias.n75 commonsourceibias.n73 0.573776
R12810 commonsourceibias.n77 commonsourceibias.n75 0.573776
R12811 commonsourceibias.n82 commonsourceibias.n80 0.573776
R12812 commonsourceibias.n242 commonsourceibias.n240 0.573776
R12813 commonsourceibias.n311 commonsourceibias.n309 0.573776
R12814 commonsourceibias.n309 commonsourceibias.n307 0.573776
R12815 commonsourceibias.n83 commonsourceibias.n77 0.287138
R12816 commonsourceibias.n83 commonsourceibias.n82 0.287138
R12817 commonsourceibias.n312 commonsourceibias.n242 0.287138
R12818 commonsourceibias.n312 commonsourceibias.n311 0.287138
R12819 commonsourceibias.n71 commonsourceibias.n9 0.285035
R12820 commonsourceibias.n137 commonsourceibias.n0 0.285035
R12821 commonsourceibias.n200 commonsourceibias.n138 0.285035
R12822 commonsourceibias.n305 commonsourceibias.n243 0.285035
R12823 commonsourceibias.n339 commonsourceibias.n202 0.285035
R12824 commonsourceibias.n402 commonsourceibias.n340 0.285035
R12825 commonsourceibias.n16 commonsourceibias.n14 0.246418
R12826 commonsourceibias.n38 commonsourceibias.n19 0.246418
R12827 commonsourceibias.n7 commonsourceibias.n5 0.246418
R12828 commonsourceibias.n104 commonsourceibias.n85 0.246418
R12829 commonsourceibias.n167 commonsourceibias.n148 0.246418
R12830 commonsourceibias.n145 commonsourceibias.n143 0.246418
R12831 commonsourceibias.n271 commonsourceibias.n252 0.246418
R12832 commonsourceibias.n284 commonsourceibias.n248 0.246418
R12833 commonsourceibias.n318 commonsourceibias.n207 0.246418
R12834 commonsourceibias.n230 commonsourceibias.n211 0.246418
R12835 commonsourceibias.n368 commonsourceibias.n349 0.246418
R12836 commonsourceibias.n381 commonsourceibias.n345 0.246418
R12837 commonsourceibias.n67 commonsourceibias.n9 0.189894
R12838 commonsourceibias.n67 commonsourceibias.n66 0.189894
R12839 commonsourceibias.n66 commonsourceibias.n11 0.189894
R12840 commonsourceibias.n61 commonsourceibias.n11 0.189894
R12841 commonsourceibias.n61 commonsourceibias.n60 0.189894
R12842 commonsourceibias.n60 commonsourceibias.n59 0.189894
R12843 commonsourceibias.n59 commonsourceibias.n13 0.189894
R12844 commonsourceibias.n54 commonsourceibias.n13 0.189894
R12845 commonsourceibias.n54 commonsourceibias.n53 0.189894
R12846 commonsourceibias.n53 commonsourceibias.n52 0.189894
R12847 commonsourceibias.n52 commonsourceibias.n15 0.189894
R12848 commonsourceibias.n47 commonsourceibias.n15 0.189894
R12849 commonsourceibias.n47 commonsourceibias.n46 0.189894
R12850 commonsourceibias.n46 commonsourceibias.n45 0.189894
R12851 commonsourceibias.n45 commonsourceibias.n18 0.189894
R12852 commonsourceibias.n40 commonsourceibias.n18 0.189894
R12853 commonsourceibias.n40 commonsourceibias.n39 0.189894
R12854 commonsourceibias.n39 commonsourceibias.n20 0.189894
R12855 commonsourceibias.n35 commonsourceibias.n20 0.189894
R12856 commonsourceibias.n35 commonsourceibias.n34 0.189894
R12857 commonsourceibias.n34 commonsourceibias.n22 0.189894
R12858 commonsourceibias.n30 commonsourceibias.n22 0.189894
R12859 commonsourceibias.n30 commonsourceibias.n29 0.189894
R12860 commonsourceibias.n29 commonsourceibias.n24 0.189894
R12861 commonsourceibias.n111 commonsourceibias.n84 0.189894
R12862 commonsourceibias.n106 commonsourceibias.n84 0.189894
R12863 commonsourceibias.n106 commonsourceibias.n105 0.189894
R12864 commonsourceibias.n105 commonsourceibias.n86 0.189894
R12865 commonsourceibias.n101 commonsourceibias.n86 0.189894
R12866 commonsourceibias.n101 commonsourceibias.n100 0.189894
R12867 commonsourceibias.n100 commonsourceibias.n88 0.189894
R12868 commonsourceibias.n96 commonsourceibias.n88 0.189894
R12869 commonsourceibias.n96 commonsourceibias.n95 0.189894
R12870 commonsourceibias.n95 commonsourceibias.n90 0.189894
R12871 commonsourceibias.n133 commonsourceibias.n0 0.189894
R12872 commonsourceibias.n133 commonsourceibias.n132 0.189894
R12873 commonsourceibias.n132 commonsourceibias.n2 0.189894
R12874 commonsourceibias.n127 commonsourceibias.n2 0.189894
R12875 commonsourceibias.n127 commonsourceibias.n126 0.189894
R12876 commonsourceibias.n126 commonsourceibias.n125 0.189894
R12877 commonsourceibias.n125 commonsourceibias.n4 0.189894
R12878 commonsourceibias.n120 commonsourceibias.n4 0.189894
R12879 commonsourceibias.n120 commonsourceibias.n119 0.189894
R12880 commonsourceibias.n119 commonsourceibias.n118 0.189894
R12881 commonsourceibias.n118 commonsourceibias.n6 0.189894
R12882 commonsourceibias.n113 commonsourceibias.n6 0.189894
R12883 commonsourceibias.n196 commonsourceibias.n138 0.189894
R12884 commonsourceibias.n196 commonsourceibias.n195 0.189894
R12885 commonsourceibias.n195 commonsourceibias.n140 0.189894
R12886 commonsourceibias.n190 commonsourceibias.n140 0.189894
R12887 commonsourceibias.n190 commonsourceibias.n189 0.189894
R12888 commonsourceibias.n189 commonsourceibias.n188 0.189894
R12889 commonsourceibias.n188 commonsourceibias.n142 0.189894
R12890 commonsourceibias.n183 commonsourceibias.n142 0.189894
R12891 commonsourceibias.n183 commonsourceibias.n182 0.189894
R12892 commonsourceibias.n182 commonsourceibias.n181 0.189894
R12893 commonsourceibias.n181 commonsourceibias.n144 0.189894
R12894 commonsourceibias.n176 commonsourceibias.n144 0.189894
R12895 commonsourceibias.n176 commonsourceibias.n175 0.189894
R12896 commonsourceibias.n175 commonsourceibias.n174 0.189894
R12897 commonsourceibias.n174 commonsourceibias.n147 0.189894
R12898 commonsourceibias.n169 commonsourceibias.n147 0.189894
R12899 commonsourceibias.n169 commonsourceibias.n168 0.189894
R12900 commonsourceibias.n168 commonsourceibias.n149 0.189894
R12901 commonsourceibias.n164 commonsourceibias.n149 0.189894
R12902 commonsourceibias.n164 commonsourceibias.n163 0.189894
R12903 commonsourceibias.n163 commonsourceibias.n151 0.189894
R12904 commonsourceibias.n159 commonsourceibias.n151 0.189894
R12905 commonsourceibias.n159 commonsourceibias.n158 0.189894
R12906 commonsourceibias.n158 commonsourceibias.n153 0.189894
R12907 commonsourceibias.n262 commonsourceibias.n257 0.189894
R12908 commonsourceibias.n263 commonsourceibias.n262 0.189894
R12909 commonsourceibias.n263 commonsourceibias.n255 0.189894
R12910 commonsourceibias.n267 commonsourceibias.n255 0.189894
R12911 commonsourceibias.n268 commonsourceibias.n267 0.189894
R12912 commonsourceibias.n268 commonsourceibias.n253 0.189894
R12913 commonsourceibias.n272 commonsourceibias.n253 0.189894
R12914 commonsourceibias.n273 commonsourceibias.n272 0.189894
R12915 commonsourceibias.n273 commonsourceibias.n251 0.189894
R12916 commonsourceibias.n278 commonsourceibias.n251 0.189894
R12917 commonsourceibias.n279 commonsourceibias.n278 0.189894
R12918 commonsourceibias.n280 commonsourceibias.n279 0.189894
R12919 commonsourceibias.n280 commonsourceibias.n249 0.189894
R12920 commonsourceibias.n286 commonsourceibias.n249 0.189894
R12921 commonsourceibias.n287 commonsourceibias.n286 0.189894
R12922 commonsourceibias.n288 commonsourceibias.n287 0.189894
R12923 commonsourceibias.n288 commonsourceibias.n247 0.189894
R12924 commonsourceibias.n293 commonsourceibias.n247 0.189894
R12925 commonsourceibias.n294 commonsourceibias.n293 0.189894
R12926 commonsourceibias.n295 commonsourceibias.n294 0.189894
R12927 commonsourceibias.n295 commonsourceibias.n245 0.189894
R12928 commonsourceibias.n300 commonsourceibias.n245 0.189894
R12929 commonsourceibias.n301 commonsourceibias.n300 0.189894
R12930 commonsourceibias.n301 commonsourceibias.n243 0.189894
R12931 commonsourceibias.n221 commonsourceibias.n216 0.189894
R12932 commonsourceibias.n222 commonsourceibias.n221 0.189894
R12933 commonsourceibias.n222 commonsourceibias.n214 0.189894
R12934 commonsourceibias.n226 commonsourceibias.n214 0.189894
R12935 commonsourceibias.n227 commonsourceibias.n226 0.189894
R12936 commonsourceibias.n227 commonsourceibias.n212 0.189894
R12937 commonsourceibias.n231 commonsourceibias.n212 0.189894
R12938 commonsourceibias.n232 commonsourceibias.n231 0.189894
R12939 commonsourceibias.n232 commonsourceibias.n210 0.189894
R12940 commonsourceibias.n237 commonsourceibias.n210 0.189894
R12941 commonsourceibias.n314 commonsourceibias.n208 0.189894
R12942 commonsourceibias.n320 commonsourceibias.n208 0.189894
R12943 commonsourceibias.n321 commonsourceibias.n320 0.189894
R12944 commonsourceibias.n322 commonsourceibias.n321 0.189894
R12945 commonsourceibias.n322 commonsourceibias.n206 0.189894
R12946 commonsourceibias.n327 commonsourceibias.n206 0.189894
R12947 commonsourceibias.n328 commonsourceibias.n327 0.189894
R12948 commonsourceibias.n329 commonsourceibias.n328 0.189894
R12949 commonsourceibias.n329 commonsourceibias.n204 0.189894
R12950 commonsourceibias.n334 commonsourceibias.n204 0.189894
R12951 commonsourceibias.n335 commonsourceibias.n334 0.189894
R12952 commonsourceibias.n335 commonsourceibias.n202 0.189894
R12953 commonsourceibias.n359 commonsourceibias.n354 0.189894
R12954 commonsourceibias.n360 commonsourceibias.n359 0.189894
R12955 commonsourceibias.n360 commonsourceibias.n352 0.189894
R12956 commonsourceibias.n364 commonsourceibias.n352 0.189894
R12957 commonsourceibias.n365 commonsourceibias.n364 0.189894
R12958 commonsourceibias.n365 commonsourceibias.n350 0.189894
R12959 commonsourceibias.n369 commonsourceibias.n350 0.189894
R12960 commonsourceibias.n370 commonsourceibias.n369 0.189894
R12961 commonsourceibias.n370 commonsourceibias.n348 0.189894
R12962 commonsourceibias.n375 commonsourceibias.n348 0.189894
R12963 commonsourceibias.n376 commonsourceibias.n375 0.189894
R12964 commonsourceibias.n377 commonsourceibias.n376 0.189894
R12965 commonsourceibias.n377 commonsourceibias.n346 0.189894
R12966 commonsourceibias.n383 commonsourceibias.n346 0.189894
R12967 commonsourceibias.n384 commonsourceibias.n383 0.189894
R12968 commonsourceibias.n385 commonsourceibias.n384 0.189894
R12969 commonsourceibias.n385 commonsourceibias.n344 0.189894
R12970 commonsourceibias.n390 commonsourceibias.n344 0.189894
R12971 commonsourceibias.n391 commonsourceibias.n390 0.189894
R12972 commonsourceibias.n392 commonsourceibias.n391 0.189894
R12973 commonsourceibias.n392 commonsourceibias.n342 0.189894
R12974 commonsourceibias.n397 commonsourceibias.n342 0.189894
R12975 commonsourceibias.n398 commonsourceibias.n397 0.189894
R12976 commonsourceibias.n398 commonsourceibias.n340 0.189894
R12977 commonsourceibias.n112 commonsourceibias.n111 0.170955
R12978 commonsourceibias.n113 commonsourceibias.n112 0.170955
R12979 commonsourceibias.n313 commonsourceibias.n237 0.170955
R12980 commonsourceibias.n314 commonsourceibias.n313 0.170955
R12981 CSoutput.n19 CSoutput.t141 184.661
R12982 CSoutput.n78 CSoutput.n77 165.8
R12983 CSoutput.n76 CSoutput.n0 165.8
R12984 CSoutput.n75 CSoutput.n74 165.8
R12985 CSoutput.n73 CSoutput.n72 165.8
R12986 CSoutput.n71 CSoutput.n2 165.8
R12987 CSoutput.n69 CSoutput.n68 165.8
R12988 CSoutput.n67 CSoutput.n3 165.8
R12989 CSoutput.n66 CSoutput.n65 165.8
R12990 CSoutput.n63 CSoutput.n4 165.8
R12991 CSoutput.n61 CSoutput.n60 165.8
R12992 CSoutput.n59 CSoutput.n5 165.8
R12993 CSoutput.n58 CSoutput.n57 165.8
R12994 CSoutput.n55 CSoutput.n6 165.8
R12995 CSoutput.n54 CSoutput.n53 165.8
R12996 CSoutput.n52 CSoutput.n51 165.8
R12997 CSoutput.n50 CSoutput.n8 165.8
R12998 CSoutput.n48 CSoutput.n47 165.8
R12999 CSoutput.n46 CSoutput.n9 165.8
R13000 CSoutput.n45 CSoutput.n44 165.8
R13001 CSoutput.n42 CSoutput.n10 165.8
R13002 CSoutput.n41 CSoutput.n40 165.8
R13003 CSoutput.n39 CSoutput.n38 165.8
R13004 CSoutput.n37 CSoutput.n12 165.8
R13005 CSoutput.n35 CSoutput.n34 165.8
R13006 CSoutput.n33 CSoutput.n13 165.8
R13007 CSoutput.n32 CSoutput.n31 165.8
R13008 CSoutput.n29 CSoutput.n14 165.8
R13009 CSoutput.n28 CSoutput.n27 165.8
R13010 CSoutput.n26 CSoutput.n25 165.8
R13011 CSoutput.n24 CSoutput.n16 165.8
R13012 CSoutput.n22 CSoutput.n21 165.8
R13013 CSoutput.n20 CSoutput.n17 165.8
R13014 CSoutput.n77 CSoutput.t120 162.194
R13015 CSoutput.n18 CSoutput.t121 120.501
R13016 CSoutput.n23 CSoutput.t131 120.501
R13017 CSoutput.n15 CSoutput.t127 120.501
R13018 CSoutput.n30 CSoutput.t123 120.501
R13019 CSoutput.n36 CSoutput.t134 120.501
R13020 CSoutput.n11 CSoutput.t136 120.501
R13021 CSoutput.n43 CSoutput.t125 120.501
R13022 CSoutput.n49 CSoutput.t137 120.501
R13023 CSoutput.n7 CSoutput.t138 120.501
R13024 CSoutput.n56 CSoutput.t132 120.501
R13025 CSoutput.n62 CSoutput.t124 120.501
R13026 CSoutput.n64 CSoutput.t140 120.501
R13027 CSoutput.n70 CSoutput.t135 120.501
R13028 CSoutput.n1 CSoutput.t130 120.501
R13029 CSoutput.n290 CSoutput.n288 103.469
R13030 CSoutput.n278 CSoutput.n276 103.469
R13031 CSoutput.n267 CSoutput.n265 103.469
R13032 CSoutput.n104 CSoutput.n102 103.469
R13033 CSoutput.n92 CSoutput.n90 103.469
R13034 CSoutput.n81 CSoutput.n79 103.469
R13035 CSoutput.n296 CSoutput.n295 103.111
R13036 CSoutput.n294 CSoutput.n293 103.111
R13037 CSoutput.n292 CSoutput.n291 103.111
R13038 CSoutput.n290 CSoutput.n289 103.111
R13039 CSoutput.n286 CSoutput.n285 103.111
R13040 CSoutput.n284 CSoutput.n283 103.111
R13041 CSoutput.n282 CSoutput.n281 103.111
R13042 CSoutput.n280 CSoutput.n279 103.111
R13043 CSoutput.n278 CSoutput.n277 103.111
R13044 CSoutput.n275 CSoutput.n274 103.111
R13045 CSoutput.n273 CSoutput.n272 103.111
R13046 CSoutput.n271 CSoutput.n270 103.111
R13047 CSoutput.n269 CSoutput.n268 103.111
R13048 CSoutput.n267 CSoutput.n266 103.111
R13049 CSoutput.n104 CSoutput.n103 103.111
R13050 CSoutput.n106 CSoutput.n105 103.111
R13051 CSoutput.n108 CSoutput.n107 103.111
R13052 CSoutput.n110 CSoutput.n109 103.111
R13053 CSoutput.n112 CSoutput.n111 103.111
R13054 CSoutput.n92 CSoutput.n91 103.111
R13055 CSoutput.n94 CSoutput.n93 103.111
R13056 CSoutput.n96 CSoutput.n95 103.111
R13057 CSoutput.n98 CSoutput.n97 103.111
R13058 CSoutput.n100 CSoutput.n99 103.111
R13059 CSoutput.n81 CSoutput.n80 103.111
R13060 CSoutput.n83 CSoutput.n82 103.111
R13061 CSoutput.n85 CSoutput.n84 103.111
R13062 CSoutput.n87 CSoutput.n86 103.111
R13063 CSoutput.n89 CSoutput.n88 103.111
R13064 CSoutput.n298 CSoutput.n297 103.111
R13065 CSoutput.n314 CSoutput.n312 81.5057
R13066 CSoutput.n303 CSoutput.n301 81.5057
R13067 CSoutput.n338 CSoutput.n336 81.5057
R13068 CSoutput.n327 CSoutput.n325 81.5057
R13069 CSoutput.n322 CSoutput.n321 80.9324
R13070 CSoutput.n320 CSoutput.n319 80.9324
R13071 CSoutput.n318 CSoutput.n317 80.9324
R13072 CSoutput.n316 CSoutput.n315 80.9324
R13073 CSoutput.n314 CSoutput.n313 80.9324
R13074 CSoutput.n311 CSoutput.n310 80.9324
R13075 CSoutput.n309 CSoutput.n308 80.9324
R13076 CSoutput.n307 CSoutput.n306 80.9324
R13077 CSoutput.n305 CSoutput.n304 80.9324
R13078 CSoutput.n303 CSoutput.n302 80.9324
R13079 CSoutput.n338 CSoutput.n337 80.9324
R13080 CSoutput.n340 CSoutput.n339 80.9324
R13081 CSoutput.n342 CSoutput.n341 80.9324
R13082 CSoutput.n344 CSoutput.n343 80.9324
R13083 CSoutput.n346 CSoutput.n345 80.9324
R13084 CSoutput.n327 CSoutput.n326 80.9324
R13085 CSoutput.n329 CSoutput.n328 80.9324
R13086 CSoutput.n331 CSoutput.n330 80.9324
R13087 CSoutput.n333 CSoutput.n332 80.9324
R13088 CSoutput.n335 CSoutput.n334 80.9324
R13089 CSoutput.n25 CSoutput.n24 48.1486
R13090 CSoutput.n69 CSoutput.n3 48.1486
R13091 CSoutput.n38 CSoutput.n37 48.1486
R13092 CSoutput.n42 CSoutput.n41 48.1486
R13093 CSoutput.n51 CSoutput.n50 48.1486
R13094 CSoutput.n55 CSoutput.n54 48.1486
R13095 CSoutput.n22 CSoutput.n17 46.462
R13096 CSoutput.n72 CSoutput.n71 46.462
R13097 CSoutput.n20 CSoutput.n19 44.9055
R13098 CSoutput.n29 CSoutput.n28 43.7635
R13099 CSoutput.n65 CSoutput.n63 43.7635
R13100 CSoutput.n35 CSoutput.n13 41.7396
R13101 CSoutput.n57 CSoutput.n5 41.7396
R13102 CSoutput.n44 CSoutput.n9 37.0171
R13103 CSoutput.n48 CSoutput.n9 37.0171
R13104 CSoutput.n76 CSoutput.n75 34.9932
R13105 CSoutput.n31 CSoutput.n13 32.2947
R13106 CSoutput.n61 CSoutput.n5 32.2947
R13107 CSoutput.n30 CSoutput.n29 29.6014
R13108 CSoutput.n63 CSoutput.n62 29.6014
R13109 CSoutput.n19 CSoutput.n18 28.4085
R13110 CSoutput.n18 CSoutput.n17 25.1176
R13111 CSoutput.n72 CSoutput.n1 25.1176
R13112 CSoutput.n43 CSoutput.n42 22.0922
R13113 CSoutput.n50 CSoutput.n49 22.0922
R13114 CSoutput.n77 CSoutput.n76 21.8586
R13115 CSoutput.n37 CSoutput.n36 18.9681
R13116 CSoutput.n56 CSoutput.n55 18.9681
R13117 CSoutput.n25 CSoutput.n15 17.6292
R13118 CSoutput.n64 CSoutput.n3 17.6292
R13119 CSoutput.n24 CSoutput.n23 15.844
R13120 CSoutput.n70 CSoutput.n69 15.844
R13121 CSoutput.n38 CSoutput.n11 14.5051
R13122 CSoutput.n54 CSoutput.n7 14.5051
R13123 CSoutput.n349 CSoutput.n78 11.6139
R13124 CSoutput.n41 CSoutput.n11 11.3811
R13125 CSoutput.n51 CSoutput.n7 11.3811
R13126 CSoutput.n23 CSoutput.n22 10.0422
R13127 CSoutput.n71 CSoutput.n70 10.0422
R13128 CSoutput.n287 CSoutput.n275 9.25285
R13129 CSoutput.n101 CSoutput.n89 9.25285
R13130 CSoutput.n323 CSoutput.n311 8.97993
R13131 CSoutput.n347 CSoutput.n335 8.97993
R13132 CSoutput.n324 CSoutput.n300 8.82427
R13133 CSoutput.n28 CSoutput.n15 8.25698
R13134 CSoutput.n65 CSoutput.n64 8.25698
R13135 CSoutput.n324 CSoutput.n323 7.89345
R13136 CSoutput.n348 CSoutput.n347 7.89345
R13137 CSoutput.n300 CSoutput.n299 7.12641
R13138 CSoutput.n114 CSoutput.n113 7.12641
R13139 CSoutput.n36 CSoutput.n35 6.91809
R13140 CSoutput.n57 CSoutput.n56 6.91809
R13141 CSoutput.n323 CSoutput.n322 5.25266
R13142 CSoutput.n347 CSoutput.n346 5.25266
R13143 CSoutput.n349 CSoutput.n114 5.23183
R13144 CSoutput.n299 CSoutput.n298 5.1449
R13145 CSoutput.n287 CSoutput.n286 5.1449
R13146 CSoutput.n113 CSoutput.n112 5.1449
R13147 CSoutput.n101 CSoutput.n100 5.1449
R13148 CSoutput.n205 CSoutput.n158 4.5005
R13149 CSoutput.n174 CSoutput.n158 4.5005
R13150 CSoutput.n169 CSoutput.n153 4.5005
R13151 CSoutput.n169 CSoutput.n155 4.5005
R13152 CSoutput.n169 CSoutput.n152 4.5005
R13153 CSoutput.n169 CSoutput.n156 4.5005
R13154 CSoutput.n169 CSoutput.n151 4.5005
R13155 CSoutput.n169 CSoutput.t126 4.5005
R13156 CSoutput.n169 CSoutput.n150 4.5005
R13157 CSoutput.n169 CSoutput.n157 4.5005
R13158 CSoutput.n169 CSoutput.n158 4.5005
R13159 CSoutput.n167 CSoutput.n153 4.5005
R13160 CSoutput.n167 CSoutput.n155 4.5005
R13161 CSoutput.n167 CSoutput.n152 4.5005
R13162 CSoutput.n167 CSoutput.n156 4.5005
R13163 CSoutput.n167 CSoutput.n151 4.5005
R13164 CSoutput.n167 CSoutput.t126 4.5005
R13165 CSoutput.n167 CSoutput.n150 4.5005
R13166 CSoutput.n167 CSoutput.n157 4.5005
R13167 CSoutput.n167 CSoutput.n158 4.5005
R13168 CSoutput.n166 CSoutput.n153 4.5005
R13169 CSoutput.n166 CSoutput.n155 4.5005
R13170 CSoutput.n166 CSoutput.n152 4.5005
R13171 CSoutput.n166 CSoutput.n156 4.5005
R13172 CSoutput.n166 CSoutput.n151 4.5005
R13173 CSoutput.n166 CSoutput.t126 4.5005
R13174 CSoutput.n166 CSoutput.n150 4.5005
R13175 CSoutput.n166 CSoutput.n157 4.5005
R13176 CSoutput.n166 CSoutput.n158 4.5005
R13177 CSoutput.n251 CSoutput.n153 4.5005
R13178 CSoutput.n251 CSoutput.n155 4.5005
R13179 CSoutput.n251 CSoutput.n152 4.5005
R13180 CSoutput.n251 CSoutput.n156 4.5005
R13181 CSoutput.n251 CSoutput.n151 4.5005
R13182 CSoutput.n251 CSoutput.t126 4.5005
R13183 CSoutput.n251 CSoutput.n150 4.5005
R13184 CSoutput.n251 CSoutput.n157 4.5005
R13185 CSoutput.n251 CSoutput.n158 4.5005
R13186 CSoutput.n249 CSoutput.n153 4.5005
R13187 CSoutput.n249 CSoutput.n155 4.5005
R13188 CSoutput.n249 CSoutput.n152 4.5005
R13189 CSoutput.n249 CSoutput.n156 4.5005
R13190 CSoutput.n249 CSoutput.n151 4.5005
R13191 CSoutput.n249 CSoutput.t126 4.5005
R13192 CSoutput.n249 CSoutput.n150 4.5005
R13193 CSoutput.n249 CSoutput.n157 4.5005
R13194 CSoutput.n247 CSoutput.n153 4.5005
R13195 CSoutput.n247 CSoutput.n155 4.5005
R13196 CSoutput.n247 CSoutput.n152 4.5005
R13197 CSoutput.n247 CSoutput.n156 4.5005
R13198 CSoutput.n247 CSoutput.n151 4.5005
R13199 CSoutput.n247 CSoutput.t126 4.5005
R13200 CSoutput.n247 CSoutput.n150 4.5005
R13201 CSoutput.n247 CSoutput.n157 4.5005
R13202 CSoutput.n177 CSoutput.n153 4.5005
R13203 CSoutput.n177 CSoutput.n155 4.5005
R13204 CSoutput.n177 CSoutput.n152 4.5005
R13205 CSoutput.n177 CSoutput.n156 4.5005
R13206 CSoutput.n177 CSoutput.n151 4.5005
R13207 CSoutput.n177 CSoutput.t126 4.5005
R13208 CSoutput.n177 CSoutput.n150 4.5005
R13209 CSoutput.n177 CSoutput.n157 4.5005
R13210 CSoutput.n177 CSoutput.n158 4.5005
R13211 CSoutput.n176 CSoutput.n153 4.5005
R13212 CSoutput.n176 CSoutput.n155 4.5005
R13213 CSoutput.n176 CSoutput.n152 4.5005
R13214 CSoutput.n176 CSoutput.n156 4.5005
R13215 CSoutput.n176 CSoutput.n151 4.5005
R13216 CSoutput.n176 CSoutput.t126 4.5005
R13217 CSoutput.n176 CSoutput.n150 4.5005
R13218 CSoutput.n176 CSoutput.n157 4.5005
R13219 CSoutput.n176 CSoutput.n158 4.5005
R13220 CSoutput.n180 CSoutput.n153 4.5005
R13221 CSoutput.n180 CSoutput.n155 4.5005
R13222 CSoutput.n180 CSoutput.n152 4.5005
R13223 CSoutput.n180 CSoutput.n156 4.5005
R13224 CSoutput.n180 CSoutput.n151 4.5005
R13225 CSoutput.n180 CSoutput.t126 4.5005
R13226 CSoutput.n180 CSoutput.n150 4.5005
R13227 CSoutput.n180 CSoutput.n157 4.5005
R13228 CSoutput.n180 CSoutput.n158 4.5005
R13229 CSoutput.n179 CSoutput.n153 4.5005
R13230 CSoutput.n179 CSoutput.n155 4.5005
R13231 CSoutput.n179 CSoutput.n152 4.5005
R13232 CSoutput.n179 CSoutput.n156 4.5005
R13233 CSoutput.n179 CSoutput.n151 4.5005
R13234 CSoutput.n179 CSoutput.t126 4.5005
R13235 CSoutput.n179 CSoutput.n150 4.5005
R13236 CSoutput.n179 CSoutput.n157 4.5005
R13237 CSoutput.n179 CSoutput.n158 4.5005
R13238 CSoutput.n162 CSoutput.n153 4.5005
R13239 CSoutput.n162 CSoutput.n155 4.5005
R13240 CSoutput.n162 CSoutput.n152 4.5005
R13241 CSoutput.n162 CSoutput.n156 4.5005
R13242 CSoutput.n162 CSoutput.n151 4.5005
R13243 CSoutput.n162 CSoutput.t126 4.5005
R13244 CSoutput.n162 CSoutput.n150 4.5005
R13245 CSoutput.n162 CSoutput.n157 4.5005
R13246 CSoutput.n162 CSoutput.n158 4.5005
R13247 CSoutput.n254 CSoutput.n153 4.5005
R13248 CSoutput.n254 CSoutput.n155 4.5005
R13249 CSoutput.n254 CSoutput.n152 4.5005
R13250 CSoutput.n254 CSoutput.n156 4.5005
R13251 CSoutput.n254 CSoutput.n151 4.5005
R13252 CSoutput.n254 CSoutput.t126 4.5005
R13253 CSoutput.n254 CSoutput.n150 4.5005
R13254 CSoutput.n254 CSoutput.n157 4.5005
R13255 CSoutput.n254 CSoutput.n158 4.5005
R13256 CSoutput.n241 CSoutput.n212 4.5005
R13257 CSoutput.n241 CSoutput.n218 4.5005
R13258 CSoutput.n199 CSoutput.n188 4.5005
R13259 CSoutput.n199 CSoutput.n190 4.5005
R13260 CSoutput.n199 CSoutput.n187 4.5005
R13261 CSoutput.n199 CSoutput.n191 4.5005
R13262 CSoutput.n199 CSoutput.n186 4.5005
R13263 CSoutput.n199 CSoutput.t122 4.5005
R13264 CSoutput.n199 CSoutput.n185 4.5005
R13265 CSoutput.n199 CSoutput.n192 4.5005
R13266 CSoutput.n241 CSoutput.n199 4.5005
R13267 CSoutput.n220 CSoutput.n188 4.5005
R13268 CSoutput.n220 CSoutput.n190 4.5005
R13269 CSoutput.n220 CSoutput.n187 4.5005
R13270 CSoutput.n220 CSoutput.n191 4.5005
R13271 CSoutput.n220 CSoutput.n186 4.5005
R13272 CSoutput.n220 CSoutput.t122 4.5005
R13273 CSoutput.n220 CSoutput.n185 4.5005
R13274 CSoutput.n220 CSoutput.n192 4.5005
R13275 CSoutput.n241 CSoutput.n220 4.5005
R13276 CSoutput.n198 CSoutput.n188 4.5005
R13277 CSoutput.n198 CSoutput.n190 4.5005
R13278 CSoutput.n198 CSoutput.n187 4.5005
R13279 CSoutput.n198 CSoutput.n191 4.5005
R13280 CSoutput.n198 CSoutput.n186 4.5005
R13281 CSoutput.n198 CSoutput.t122 4.5005
R13282 CSoutput.n198 CSoutput.n185 4.5005
R13283 CSoutput.n198 CSoutput.n192 4.5005
R13284 CSoutput.n241 CSoutput.n198 4.5005
R13285 CSoutput.n222 CSoutput.n188 4.5005
R13286 CSoutput.n222 CSoutput.n190 4.5005
R13287 CSoutput.n222 CSoutput.n187 4.5005
R13288 CSoutput.n222 CSoutput.n191 4.5005
R13289 CSoutput.n222 CSoutput.n186 4.5005
R13290 CSoutput.n222 CSoutput.t122 4.5005
R13291 CSoutput.n222 CSoutput.n185 4.5005
R13292 CSoutput.n222 CSoutput.n192 4.5005
R13293 CSoutput.n241 CSoutput.n222 4.5005
R13294 CSoutput.n188 CSoutput.n183 4.5005
R13295 CSoutput.n190 CSoutput.n183 4.5005
R13296 CSoutput.n187 CSoutput.n183 4.5005
R13297 CSoutput.n191 CSoutput.n183 4.5005
R13298 CSoutput.n186 CSoutput.n183 4.5005
R13299 CSoutput.t122 CSoutput.n183 4.5005
R13300 CSoutput.n185 CSoutput.n183 4.5005
R13301 CSoutput.n192 CSoutput.n183 4.5005
R13302 CSoutput.n244 CSoutput.n188 4.5005
R13303 CSoutput.n244 CSoutput.n190 4.5005
R13304 CSoutput.n244 CSoutput.n187 4.5005
R13305 CSoutput.n244 CSoutput.n191 4.5005
R13306 CSoutput.n244 CSoutput.n186 4.5005
R13307 CSoutput.n244 CSoutput.t122 4.5005
R13308 CSoutput.n244 CSoutput.n185 4.5005
R13309 CSoutput.n244 CSoutput.n192 4.5005
R13310 CSoutput.n242 CSoutput.n188 4.5005
R13311 CSoutput.n242 CSoutput.n190 4.5005
R13312 CSoutput.n242 CSoutput.n187 4.5005
R13313 CSoutput.n242 CSoutput.n191 4.5005
R13314 CSoutput.n242 CSoutput.n186 4.5005
R13315 CSoutput.n242 CSoutput.t122 4.5005
R13316 CSoutput.n242 CSoutput.n185 4.5005
R13317 CSoutput.n242 CSoutput.n192 4.5005
R13318 CSoutput.n242 CSoutput.n241 4.5005
R13319 CSoutput.n224 CSoutput.n188 4.5005
R13320 CSoutput.n224 CSoutput.n190 4.5005
R13321 CSoutput.n224 CSoutput.n187 4.5005
R13322 CSoutput.n224 CSoutput.n191 4.5005
R13323 CSoutput.n224 CSoutput.n186 4.5005
R13324 CSoutput.n224 CSoutput.t122 4.5005
R13325 CSoutput.n224 CSoutput.n185 4.5005
R13326 CSoutput.n224 CSoutput.n192 4.5005
R13327 CSoutput.n241 CSoutput.n224 4.5005
R13328 CSoutput.n196 CSoutput.n188 4.5005
R13329 CSoutput.n196 CSoutput.n190 4.5005
R13330 CSoutput.n196 CSoutput.n187 4.5005
R13331 CSoutput.n196 CSoutput.n191 4.5005
R13332 CSoutput.n196 CSoutput.n186 4.5005
R13333 CSoutput.n196 CSoutput.t122 4.5005
R13334 CSoutput.n196 CSoutput.n185 4.5005
R13335 CSoutput.n196 CSoutput.n192 4.5005
R13336 CSoutput.n241 CSoutput.n196 4.5005
R13337 CSoutput.n226 CSoutput.n188 4.5005
R13338 CSoutput.n226 CSoutput.n190 4.5005
R13339 CSoutput.n226 CSoutput.n187 4.5005
R13340 CSoutput.n226 CSoutput.n191 4.5005
R13341 CSoutput.n226 CSoutput.n186 4.5005
R13342 CSoutput.n226 CSoutput.t122 4.5005
R13343 CSoutput.n226 CSoutput.n185 4.5005
R13344 CSoutput.n226 CSoutput.n192 4.5005
R13345 CSoutput.n241 CSoutput.n226 4.5005
R13346 CSoutput.n195 CSoutput.n188 4.5005
R13347 CSoutput.n195 CSoutput.n190 4.5005
R13348 CSoutput.n195 CSoutput.n187 4.5005
R13349 CSoutput.n195 CSoutput.n191 4.5005
R13350 CSoutput.n195 CSoutput.n186 4.5005
R13351 CSoutput.n195 CSoutput.t122 4.5005
R13352 CSoutput.n195 CSoutput.n185 4.5005
R13353 CSoutput.n195 CSoutput.n192 4.5005
R13354 CSoutput.n241 CSoutput.n195 4.5005
R13355 CSoutput.n240 CSoutput.n188 4.5005
R13356 CSoutput.n240 CSoutput.n190 4.5005
R13357 CSoutput.n240 CSoutput.n187 4.5005
R13358 CSoutput.n240 CSoutput.n191 4.5005
R13359 CSoutput.n240 CSoutput.n186 4.5005
R13360 CSoutput.n240 CSoutput.t122 4.5005
R13361 CSoutput.n240 CSoutput.n185 4.5005
R13362 CSoutput.n240 CSoutput.n192 4.5005
R13363 CSoutput.n241 CSoutput.n240 4.5005
R13364 CSoutput.n239 CSoutput.n124 4.5005
R13365 CSoutput.n140 CSoutput.n124 4.5005
R13366 CSoutput.n135 CSoutput.n119 4.5005
R13367 CSoutput.n135 CSoutput.n121 4.5005
R13368 CSoutput.n135 CSoutput.n118 4.5005
R13369 CSoutput.n135 CSoutput.n122 4.5005
R13370 CSoutput.n135 CSoutput.n117 4.5005
R13371 CSoutput.n135 CSoutput.t139 4.5005
R13372 CSoutput.n135 CSoutput.n116 4.5005
R13373 CSoutput.n135 CSoutput.n123 4.5005
R13374 CSoutput.n135 CSoutput.n124 4.5005
R13375 CSoutput.n133 CSoutput.n119 4.5005
R13376 CSoutput.n133 CSoutput.n121 4.5005
R13377 CSoutput.n133 CSoutput.n118 4.5005
R13378 CSoutput.n133 CSoutput.n122 4.5005
R13379 CSoutput.n133 CSoutput.n117 4.5005
R13380 CSoutput.n133 CSoutput.t139 4.5005
R13381 CSoutput.n133 CSoutput.n116 4.5005
R13382 CSoutput.n133 CSoutput.n123 4.5005
R13383 CSoutput.n133 CSoutput.n124 4.5005
R13384 CSoutput.n132 CSoutput.n119 4.5005
R13385 CSoutput.n132 CSoutput.n121 4.5005
R13386 CSoutput.n132 CSoutput.n118 4.5005
R13387 CSoutput.n132 CSoutput.n122 4.5005
R13388 CSoutput.n132 CSoutput.n117 4.5005
R13389 CSoutput.n132 CSoutput.t139 4.5005
R13390 CSoutput.n132 CSoutput.n116 4.5005
R13391 CSoutput.n132 CSoutput.n123 4.5005
R13392 CSoutput.n132 CSoutput.n124 4.5005
R13393 CSoutput.n261 CSoutput.n119 4.5005
R13394 CSoutput.n261 CSoutput.n121 4.5005
R13395 CSoutput.n261 CSoutput.n118 4.5005
R13396 CSoutput.n261 CSoutput.n122 4.5005
R13397 CSoutput.n261 CSoutput.n117 4.5005
R13398 CSoutput.n261 CSoutput.t139 4.5005
R13399 CSoutput.n261 CSoutput.n116 4.5005
R13400 CSoutput.n261 CSoutput.n123 4.5005
R13401 CSoutput.n261 CSoutput.n124 4.5005
R13402 CSoutput.n259 CSoutput.n119 4.5005
R13403 CSoutput.n259 CSoutput.n121 4.5005
R13404 CSoutput.n259 CSoutput.n118 4.5005
R13405 CSoutput.n259 CSoutput.n122 4.5005
R13406 CSoutput.n259 CSoutput.n117 4.5005
R13407 CSoutput.n259 CSoutput.t139 4.5005
R13408 CSoutput.n259 CSoutput.n116 4.5005
R13409 CSoutput.n259 CSoutput.n123 4.5005
R13410 CSoutput.n257 CSoutput.n119 4.5005
R13411 CSoutput.n257 CSoutput.n121 4.5005
R13412 CSoutput.n257 CSoutput.n118 4.5005
R13413 CSoutput.n257 CSoutput.n122 4.5005
R13414 CSoutput.n257 CSoutput.n117 4.5005
R13415 CSoutput.n257 CSoutput.t139 4.5005
R13416 CSoutput.n257 CSoutput.n116 4.5005
R13417 CSoutput.n257 CSoutput.n123 4.5005
R13418 CSoutput.n143 CSoutput.n119 4.5005
R13419 CSoutput.n143 CSoutput.n121 4.5005
R13420 CSoutput.n143 CSoutput.n118 4.5005
R13421 CSoutput.n143 CSoutput.n122 4.5005
R13422 CSoutput.n143 CSoutput.n117 4.5005
R13423 CSoutput.n143 CSoutput.t139 4.5005
R13424 CSoutput.n143 CSoutput.n116 4.5005
R13425 CSoutput.n143 CSoutput.n123 4.5005
R13426 CSoutput.n143 CSoutput.n124 4.5005
R13427 CSoutput.n142 CSoutput.n119 4.5005
R13428 CSoutput.n142 CSoutput.n121 4.5005
R13429 CSoutput.n142 CSoutput.n118 4.5005
R13430 CSoutput.n142 CSoutput.n122 4.5005
R13431 CSoutput.n142 CSoutput.n117 4.5005
R13432 CSoutput.n142 CSoutput.t139 4.5005
R13433 CSoutput.n142 CSoutput.n116 4.5005
R13434 CSoutput.n142 CSoutput.n123 4.5005
R13435 CSoutput.n142 CSoutput.n124 4.5005
R13436 CSoutput.n146 CSoutput.n119 4.5005
R13437 CSoutput.n146 CSoutput.n121 4.5005
R13438 CSoutput.n146 CSoutput.n118 4.5005
R13439 CSoutput.n146 CSoutput.n122 4.5005
R13440 CSoutput.n146 CSoutput.n117 4.5005
R13441 CSoutput.n146 CSoutput.t139 4.5005
R13442 CSoutput.n146 CSoutput.n116 4.5005
R13443 CSoutput.n146 CSoutput.n123 4.5005
R13444 CSoutput.n146 CSoutput.n124 4.5005
R13445 CSoutput.n145 CSoutput.n119 4.5005
R13446 CSoutput.n145 CSoutput.n121 4.5005
R13447 CSoutput.n145 CSoutput.n118 4.5005
R13448 CSoutput.n145 CSoutput.n122 4.5005
R13449 CSoutput.n145 CSoutput.n117 4.5005
R13450 CSoutput.n145 CSoutput.t139 4.5005
R13451 CSoutput.n145 CSoutput.n116 4.5005
R13452 CSoutput.n145 CSoutput.n123 4.5005
R13453 CSoutput.n145 CSoutput.n124 4.5005
R13454 CSoutput.n128 CSoutput.n119 4.5005
R13455 CSoutput.n128 CSoutput.n121 4.5005
R13456 CSoutput.n128 CSoutput.n118 4.5005
R13457 CSoutput.n128 CSoutput.n122 4.5005
R13458 CSoutput.n128 CSoutput.n117 4.5005
R13459 CSoutput.n128 CSoutput.t139 4.5005
R13460 CSoutput.n128 CSoutput.n116 4.5005
R13461 CSoutput.n128 CSoutput.n123 4.5005
R13462 CSoutput.n128 CSoutput.n124 4.5005
R13463 CSoutput.n264 CSoutput.n119 4.5005
R13464 CSoutput.n264 CSoutput.n121 4.5005
R13465 CSoutput.n264 CSoutput.n118 4.5005
R13466 CSoutput.n264 CSoutput.n122 4.5005
R13467 CSoutput.n264 CSoutput.n117 4.5005
R13468 CSoutput.n264 CSoutput.t139 4.5005
R13469 CSoutput.n264 CSoutput.n116 4.5005
R13470 CSoutput.n264 CSoutput.n123 4.5005
R13471 CSoutput.n264 CSoutput.n124 4.5005
R13472 CSoutput.n299 CSoutput.n287 4.10845
R13473 CSoutput.n113 CSoutput.n101 4.10845
R13474 CSoutput.n297 CSoutput.t96 4.06363
R13475 CSoutput.n297 CSoutput.t99 4.06363
R13476 CSoutput.n295 CSoutput.t56 4.06363
R13477 CSoutput.n295 CSoutput.t75 4.06363
R13478 CSoutput.n293 CSoutput.t118 4.06363
R13479 CSoutput.n293 CSoutput.t68 4.06363
R13480 CSoutput.n291 CSoutput.t70 4.06363
R13481 CSoutput.n291 CSoutput.t93 4.06363
R13482 CSoutput.n289 CSoutput.t108 4.06363
R13483 CSoutput.n289 CSoutput.t54 4.06363
R13484 CSoutput.n288 CSoutput.t83 4.06363
R13485 CSoutput.n288 CSoutput.t82 4.06363
R13486 CSoutput.n285 CSoutput.t79 4.06363
R13487 CSoutput.n285 CSoutput.t78 4.06363
R13488 CSoutput.n283 CSoutput.t66 4.06363
R13489 CSoutput.n283 CSoutput.t114 4.06363
R13490 CSoutput.n281 CSoutput.t86 4.06363
R13491 CSoutput.n281 CSoutput.t67 4.06363
R13492 CSoutput.n279 CSoutput.t117 4.06363
R13493 CSoutput.n279 CSoutput.t105 4.06363
R13494 CSoutput.n277 CSoutput.t104 4.06363
R13495 CSoutput.n277 CSoutput.t0 4.06363
R13496 CSoutput.n276 CSoutput.t112 4.06363
R13497 CSoutput.n276 CSoutput.t101 4.06363
R13498 CSoutput.n274 CSoutput.t80 4.06363
R13499 CSoutput.n274 CSoutput.t50 4.06363
R13500 CSoutput.n272 CSoutput.t58 4.06363
R13501 CSoutput.n272 CSoutput.t88 4.06363
R13502 CSoutput.n270 CSoutput.t69 4.06363
R13503 CSoutput.n270 CSoutput.t72 4.06363
R13504 CSoutput.n268 CSoutput.t65 4.06363
R13505 CSoutput.n268 CSoutput.t92 4.06363
R13506 CSoutput.n266 CSoutput.t113 4.06363
R13507 CSoutput.n266 CSoutput.t74 4.06363
R13508 CSoutput.n265 CSoutput.t76 4.06363
R13509 CSoutput.n265 CSoutput.t62 4.06363
R13510 CSoutput.n102 CSoutput.t53 4.06363
R13511 CSoutput.n102 CSoutput.t52 4.06363
R13512 CSoutput.n103 CSoutput.t106 4.06363
R13513 CSoutput.n103 CSoutput.t95 4.06363
R13514 CSoutput.n105 CSoutput.t55 4.06363
R13515 CSoutput.n105 CSoutput.t110 4.06363
R13516 CSoutput.n107 CSoutput.t107 4.06363
R13517 CSoutput.n107 CSoutput.t100 4.06363
R13518 CSoutput.n109 CSoutput.t97 4.06363
R13519 CSoutput.n109 CSoutput.t87 4.06363
R13520 CSoutput.n111 CSoutput.t90 4.06363
R13521 CSoutput.n111 CSoutput.t91 4.06363
R13522 CSoutput.n90 CSoutput.t63 4.06363
R13523 CSoutput.n90 CSoutput.t109 4.06363
R13524 CSoutput.n91 CSoutput.t84 4.06363
R13525 CSoutput.n91 CSoutput.t51 4.06363
R13526 CSoutput.n93 CSoutput.t1 4.06363
R13527 CSoutput.n93 CSoutput.t61 4.06363
R13528 CSoutput.n95 CSoutput.t85 4.06363
R13529 CSoutput.n95 CSoutput.t57 4.06363
R13530 CSoutput.n97 CSoutput.t64 4.06363
R13531 CSoutput.n97 CSoutput.t111 4.06363
R13532 CSoutput.n99 CSoutput.t102 4.06363
R13533 CSoutput.n99 CSoutput.t103 4.06363
R13534 CSoutput.n79 CSoutput.t115 4.06363
R13535 CSoutput.n79 CSoutput.t77 4.06363
R13536 CSoutput.n80 CSoutput.t59 4.06363
R13537 CSoutput.n80 CSoutput.t116 4.06363
R13538 CSoutput.n82 CSoutput.t60 4.06363
R13539 CSoutput.n82 CSoutput.t94 4.06363
R13540 CSoutput.n84 CSoutput.t73 4.06363
R13541 CSoutput.n84 CSoutput.t98 4.06363
R13542 CSoutput.n86 CSoutput.t89 4.06363
R13543 CSoutput.n86 CSoutput.t71 4.06363
R13544 CSoutput.n88 CSoutput.t119 4.06363
R13545 CSoutput.n88 CSoutput.t81 4.06363
R13546 CSoutput.n44 CSoutput.n43 3.79402
R13547 CSoutput.n49 CSoutput.n48 3.79402
R13548 CSoutput.n349 CSoutput.n348 3.57343
R13549 CSoutput.n321 CSoutput.t40 2.82907
R13550 CSoutput.n321 CSoutput.t43 2.82907
R13551 CSoutput.n319 CSoutput.t39 2.82907
R13552 CSoutput.n319 CSoutput.t29 2.82907
R13553 CSoutput.n317 CSoutput.t6 2.82907
R13554 CSoutput.n317 CSoutput.t37 2.82907
R13555 CSoutput.n315 CSoutput.t31 2.82907
R13556 CSoutput.n315 CSoutput.t20 2.82907
R13557 CSoutput.n313 CSoutput.t48 2.82907
R13558 CSoutput.n313 CSoutput.t2 2.82907
R13559 CSoutput.n312 CSoutput.t36 2.82907
R13560 CSoutput.n312 CSoutput.t25 2.82907
R13561 CSoutput.n310 CSoutput.t33 2.82907
R13562 CSoutput.n310 CSoutput.t35 2.82907
R13563 CSoutput.n308 CSoutput.t30 2.82907
R13564 CSoutput.n308 CSoutput.t19 2.82907
R13565 CSoutput.n306 CSoutput.t47 2.82907
R13566 CSoutput.n306 CSoutput.t28 2.82907
R13567 CSoutput.n304 CSoutput.t21 2.82907
R13568 CSoutput.n304 CSoutput.t11 2.82907
R13569 CSoutput.n302 CSoutput.t42 2.82907
R13570 CSoutput.n302 CSoutput.t44 2.82907
R13571 CSoutput.n301 CSoutput.t26 2.82907
R13572 CSoutput.n301 CSoutput.t16 2.82907
R13573 CSoutput.n336 CSoutput.t12 2.82907
R13574 CSoutput.n336 CSoutput.t24 2.82907
R13575 CSoutput.n337 CSoutput.t41 2.82907
R13576 CSoutput.n337 CSoutput.t4 2.82907
R13577 CSoutput.n339 CSoutput.t8 2.82907
R13578 CSoutput.n339 CSoutput.t18 2.82907
R13579 CSoutput.n341 CSoutput.t23 2.82907
R13580 CSoutput.n341 CSoutput.t10 2.82907
R13581 CSoutput.n343 CSoutput.t15 2.82907
R13582 CSoutput.n343 CSoutput.t27 2.82907
R13583 CSoutput.n345 CSoutput.t32 2.82907
R13584 CSoutput.n345 CSoutput.t45 2.82907
R13585 CSoutput.n325 CSoutput.t5 2.82907
R13586 CSoutput.n325 CSoutput.t13 2.82907
R13587 CSoutput.n326 CSoutput.t34 2.82907
R13588 CSoutput.n326 CSoutput.t46 2.82907
R13589 CSoutput.n328 CSoutput.t49 2.82907
R13590 CSoutput.n328 CSoutput.t9 2.82907
R13591 CSoutput.n330 CSoutput.t14 2.82907
R13592 CSoutput.n330 CSoutput.t3 2.82907
R13593 CSoutput.n332 CSoutput.t7 2.82907
R13594 CSoutput.n332 CSoutput.t17 2.82907
R13595 CSoutput.n334 CSoutput.t22 2.82907
R13596 CSoutput.n334 CSoutput.t38 2.82907
R13597 CSoutput.n348 CSoutput.n324 2.75627
R13598 CSoutput.n75 CSoutput.n1 2.45513
R13599 CSoutput.n205 CSoutput.n203 2.251
R13600 CSoutput.n205 CSoutput.n202 2.251
R13601 CSoutput.n205 CSoutput.n201 2.251
R13602 CSoutput.n205 CSoutput.n200 2.251
R13603 CSoutput.n174 CSoutput.n173 2.251
R13604 CSoutput.n174 CSoutput.n172 2.251
R13605 CSoutput.n174 CSoutput.n171 2.251
R13606 CSoutput.n174 CSoutput.n170 2.251
R13607 CSoutput.n247 CSoutput.n246 2.251
R13608 CSoutput.n212 CSoutput.n210 2.251
R13609 CSoutput.n212 CSoutput.n209 2.251
R13610 CSoutput.n212 CSoutput.n208 2.251
R13611 CSoutput.n230 CSoutput.n212 2.251
R13612 CSoutput.n218 CSoutput.n217 2.251
R13613 CSoutput.n218 CSoutput.n216 2.251
R13614 CSoutput.n218 CSoutput.n215 2.251
R13615 CSoutput.n218 CSoutput.n214 2.251
R13616 CSoutput.n244 CSoutput.n184 2.251
R13617 CSoutput.n239 CSoutput.n237 2.251
R13618 CSoutput.n239 CSoutput.n236 2.251
R13619 CSoutput.n239 CSoutput.n235 2.251
R13620 CSoutput.n239 CSoutput.n234 2.251
R13621 CSoutput.n140 CSoutput.n139 2.251
R13622 CSoutput.n140 CSoutput.n138 2.251
R13623 CSoutput.n140 CSoutput.n137 2.251
R13624 CSoutput.n140 CSoutput.n136 2.251
R13625 CSoutput.n257 CSoutput.n256 2.251
R13626 CSoutput.n174 CSoutput.n154 2.2505
R13627 CSoutput.n169 CSoutput.n154 2.2505
R13628 CSoutput.n167 CSoutput.n154 2.2505
R13629 CSoutput.n166 CSoutput.n154 2.2505
R13630 CSoutput.n251 CSoutput.n154 2.2505
R13631 CSoutput.n249 CSoutput.n154 2.2505
R13632 CSoutput.n247 CSoutput.n154 2.2505
R13633 CSoutput.n177 CSoutput.n154 2.2505
R13634 CSoutput.n176 CSoutput.n154 2.2505
R13635 CSoutput.n180 CSoutput.n154 2.2505
R13636 CSoutput.n179 CSoutput.n154 2.2505
R13637 CSoutput.n162 CSoutput.n154 2.2505
R13638 CSoutput.n254 CSoutput.n154 2.2505
R13639 CSoutput.n254 CSoutput.n253 2.2505
R13640 CSoutput.n218 CSoutput.n189 2.2505
R13641 CSoutput.n199 CSoutput.n189 2.2505
R13642 CSoutput.n220 CSoutput.n189 2.2505
R13643 CSoutput.n198 CSoutput.n189 2.2505
R13644 CSoutput.n222 CSoutput.n189 2.2505
R13645 CSoutput.n189 CSoutput.n183 2.2505
R13646 CSoutput.n244 CSoutput.n189 2.2505
R13647 CSoutput.n242 CSoutput.n189 2.2505
R13648 CSoutput.n224 CSoutput.n189 2.2505
R13649 CSoutput.n196 CSoutput.n189 2.2505
R13650 CSoutput.n226 CSoutput.n189 2.2505
R13651 CSoutput.n195 CSoutput.n189 2.2505
R13652 CSoutput.n240 CSoutput.n189 2.2505
R13653 CSoutput.n240 CSoutput.n193 2.2505
R13654 CSoutput.n140 CSoutput.n120 2.2505
R13655 CSoutput.n135 CSoutput.n120 2.2505
R13656 CSoutput.n133 CSoutput.n120 2.2505
R13657 CSoutput.n132 CSoutput.n120 2.2505
R13658 CSoutput.n261 CSoutput.n120 2.2505
R13659 CSoutput.n259 CSoutput.n120 2.2505
R13660 CSoutput.n257 CSoutput.n120 2.2505
R13661 CSoutput.n143 CSoutput.n120 2.2505
R13662 CSoutput.n142 CSoutput.n120 2.2505
R13663 CSoutput.n146 CSoutput.n120 2.2505
R13664 CSoutput.n145 CSoutput.n120 2.2505
R13665 CSoutput.n128 CSoutput.n120 2.2505
R13666 CSoutput.n264 CSoutput.n120 2.2505
R13667 CSoutput.n264 CSoutput.n263 2.2505
R13668 CSoutput.n182 CSoutput.n175 2.25024
R13669 CSoutput.n182 CSoutput.n168 2.25024
R13670 CSoutput.n250 CSoutput.n182 2.25024
R13671 CSoutput.n182 CSoutput.n178 2.25024
R13672 CSoutput.n182 CSoutput.n181 2.25024
R13673 CSoutput.n182 CSoutput.n149 2.25024
R13674 CSoutput.n232 CSoutput.n229 2.25024
R13675 CSoutput.n232 CSoutput.n228 2.25024
R13676 CSoutput.n232 CSoutput.n227 2.25024
R13677 CSoutput.n232 CSoutput.n194 2.25024
R13678 CSoutput.n232 CSoutput.n231 2.25024
R13679 CSoutput.n233 CSoutput.n232 2.25024
R13680 CSoutput.n148 CSoutput.n141 2.25024
R13681 CSoutput.n148 CSoutput.n134 2.25024
R13682 CSoutput.n260 CSoutput.n148 2.25024
R13683 CSoutput.n148 CSoutput.n144 2.25024
R13684 CSoutput.n148 CSoutput.n147 2.25024
R13685 CSoutput.n148 CSoutput.n115 2.25024
R13686 CSoutput.n300 CSoutput.n114 2.15937
R13687 CSoutput.n249 CSoutput.n159 1.50111
R13688 CSoutput.n197 CSoutput.n183 1.50111
R13689 CSoutput.n259 CSoutput.n125 1.50111
R13690 CSoutput.n205 CSoutput.n204 1.501
R13691 CSoutput.n212 CSoutput.n211 1.501
R13692 CSoutput.n239 CSoutput.n238 1.501
R13693 CSoutput.n253 CSoutput.n164 1.12536
R13694 CSoutput.n253 CSoutput.n165 1.12536
R13695 CSoutput.n253 CSoutput.n252 1.12536
R13696 CSoutput.n213 CSoutput.n193 1.12536
R13697 CSoutput.n219 CSoutput.n193 1.12536
R13698 CSoutput.n221 CSoutput.n193 1.12536
R13699 CSoutput.n263 CSoutput.n130 1.12536
R13700 CSoutput.n263 CSoutput.n131 1.12536
R13701 CSoutput.n263 CSoutput.n262 1.12536
R13702 CSoutput.n253 CSoutput.n160 1.12536
R13703 CSoutput.n253 CSoutput.n161 1.12536
R13704 CSoutput.n253 CSoutput.n163 1.12536
R13705 CSoutput.n243 CSoutput.n193 1.12536
R13706 CSoutput.n223 CSoutput.n193 1.12536
R13707 CSoutput.n225 CSoutput.n193 1.12536
R13708 CSoutput.n263 CSoutput.n126 1.12536
R13709 CSoutput.n263 CSoutput.n127 1.12536
R13710 CSoutput.n263 CSoutput.n129 1.12536
R13711 CSoutput.n31 CSoutput.n30 0.669944
R13712 CSoutput.n62 CSoutput.n61 0.669944
R13713 CSoutput.n316 CSoutput.n314 0.573776
R13714 CSoutput.n318 CSoutput.n316 0.573776
R13715 CSoutput.n320 CSoutput.n318 0.573776
R13716 CSoutput.n322 CSoutput.n320 0.573776
R13717 CSoutput.n305 CSoutput.n303 0.573776
R13718 CSoutput.n307 CSoutput.n305 0.573776
R13719 CSoutput.n309 CSoutput.n307 0.573776
R13720 CSoutput.n311 CSoutput.n309 0.573776
R13721 CSoutput.n346 CSoutput.n344 0.573776
R13722 CSoutput.n344 CSoutput.n342 0.573776
R13723 CSoutput.n342 CSoutput.n340 0.573776
R13724 CSoutput.n340 CSoutput.n338 0.573776
R13725 CSoutput.n335 CSoutput.n333 0.573776
R13726 CSoutput.n333 CSoutput.n331 0.573776
R13727 CSoutput.n331 CSoutput.n329 0.573776
R13728 CSoutput.n329 CSoutput.n327 0.573776
R13729 CSoutput.n349 CSoutput.n264 0.53442
R13730 CSoutput.n292 CSoutput.n290 0.358259
R13731 CSoutput.n294 CSoutput.n292 0.358259
R13732 CSoutput.n296 CSoutput.n294 0.358259
R13733 CSoutput.n298 CSoutput.n296 0.358259
R13734 CSoutput.n280 CSoutput.n278 0.358259
R13735 CSoutput.n282 CSoutput.n280 0.358259
R13736 CSoutput.n284 CSoutput.n282 0.358259
R13737 CSoutput.n286 CSoutput.n284 0.358259
R13738 CSoutput.n269 CSoutput.n267 0.358259
R13739 CSoutput.n271 CSoutput.n269 0.358259
R13740 CSoutput.n273 CSoutput.n271 0.358259
R13741 CSoutput.n275 CSoutput.n273 0.358259
R13742 CSoutput.n112 CSoutput.n110 0.358259
R13743 CSoutput.n110 CSoutput.n108 0.358259
R13744 CSoutput.n108 CSoutput.n106 0.358259
R13745 CSoutput.n106 CSoutput.n104 0.358259
R13746 CSoutput.n100 CSoutput.n98 0.358259
R13747 CSoutput.n98 CSoutput.n96 0.358259
R13748 CSoutput.n96 CSoutput.n94 0.358259
R13749 CSoutput.n94 CSoutput.n92 0.358259
R13750 CSoutput.n89 CSoutput.n87 0.358259
R13751 CSoutput.n87 CSoutput.n85 0.358259
R13752 CSoutput.n85 CSoutput.n83 0.358259
R13753 CSoutput.n83 CSoutput.n81 0.358259
R13754 CSoutput.n21 CSoutput.n20 0.169105
R13755 CSoutput.n21 CSoutput.n16 0.169105
R13756 CSoutput.n26 CSoutput.n16 0.169105
R13757 CSoutput.n27 CSoutput.n26 0.169105
R13758 CSoutput.n27 CSoutput.n14 0.169105
R13759 CSoutput.n32 CSoutput.n14 0.169105
R13760 CSoutput.n33 CSoutput.n32 0.169105
R13761 CSoutput.n34 CSoutput.n33 0.169105
R13762 CSoutput.n34 CSoutput.n12 0.169105
R13763 CSoutput.n39 CSoutput.n12 0.169105
R13764 CSoutput.n40 CSoutput.n39 0.169105
R13765 CSoutput.n40 CSoutput.n10 0.169105
R13766 CSoutput.n45 CSoutput.n10 0.169105
R13767 CSoutput.n46 CSoutput.n45 0.169105
R13768 CSoutput.n47 CSoutput.n46 0.169105
R13769 CSoutput.n47 CSoutput.n8 0.169105
R13770 CSoutput.n52 CSoutput.n8 0.169105
R13771 CSoutput.n53 CSoutput.n52 0.169105
R13772 CSoutput.n53 CSoutput.n6 0.169105
R13773 CSoutput.n58 CSoutput.n6 0.169105
R13774 CSoutput.n59 CSoutput.n58 0.169105
R13775 CSoutput.n60 CSoutput.n59 0.169105
R13776 CSoutput.n60 CSoutput.n4 0.169105
R13777 CSoutput.n66 CSoutput.n4 0.169105
R13778 CSoutput.n67 CSoutput.n66 0.169105
R13779 CSoutput.n68 CSoutput.n67 0.169105
R13780 CSoutput.n68 CSoutput.n2 0.169105
R13781 CSoutput.n73 CSoutput.n2 0.169105
R13782 CSoutput.n74 CSoutput.n73 0.169105
R13783 CSoutput.n74 CSoutput.n0 0.169105
R13784 CSoutput.n78 CSoutput.n0 0.169105
R13785 CSoutput.n207 CSoutput.n206 0.0910737
R13786 CSoutput.n258 CSoutput.n255 0.0723685
R13787 CSoutput.n212 CSoutput.n207 0.0522944
R13788 CSoutput.n255 CSoutput.n254 0.0499135
R13789 CSoutput.n206 CSoutput.n205 0.0499135
R13790 CSoutput.n240 CSoutput.n239 0.0464294
R13791 CSoutput.n248 CSoutput.n245 0.0391444
R13792 CSoutput.n207 CSoutput.t129 0.023435
R13793 CSoutput.n255 CSoutput.t128 0.02262
R13794 CSoutput.n206 CSoutput.t133 0.02262
R13795 CSoutput CSoutput.n349 0.0052
R13796 CSoutput.n177 CSoutput.n160 0.00365111
R13797 CSoutput.n180 CSoutput.n161 0.00365111
R13798 CSoutput.n163 CSoutput.n162 0.00365111
R13799 CSoutput.n205 CSoutput.n164 0.00365111
R13800 CSoutput.n169 CSoutput.n165 0.00365111
R13801 CSoutput.n252 CSoutput.n166 0.00365111
R13802 CSoutput.n243 CSoutput.n242 0.00365111
R13803 CSoutput.n223 CSoutput.n196 0.00365111
R13804 CSoutput.n225 CSoutput.n195 0.00365111
R13805 CSoutput.n213 CSoutput.n212 0.00365111
R13806 CSoutput.n219 CSoutput.n199 0.00365111
R13807 CSoutput.n221 CSoutput.n198 0.00365111
R13808 CSoutput.n143 CSoutput.n126 0.00365111
R13809 CSoutput.n146 CSoutput.n127 0.00365111
R13810 CSoutput.n129 CSoutput.n128 0.00365111
R13811 CSoutput.n239 CSoutput.n130 0.00365111
R13812 CSoutput.n135 CSoutput.n131 0.00365111
R13813 CSoutput.n262 CSoutput.n132 0.00365111
R13814 CSoutput.n174 CSoutput.n164 0.00340054
R13815 CSoutput.n167 CSoutput.n165 0.00340054
R13816 CSoutput.n252 CSoutput.n251 0.00340054
R13817 CSoutput.n247 CSoutput.n160 0.00340054
R13818 CSoutput.n176 CSoutput.n161 0.00340054
R13819 CSoutput.n179 CSoutput.n163 0.00340054
R13820 CSoutput.n218 CSoutput.n213 0.00340054
R13821 CSoutput.n220 CSoutput.n219 0.00340054
R13822 CSoutput.n222 CSoutput.n221 0.00340054
R13823 CSoutput.n244 CSoutput.n243 0.00340054
R13824 CSoutput.n224 CSoutput.n223 0.00340054
R13825 CSoutput.n226 CSoutput.n225 0.00340054
R13826 CSoutput.n140 CSoutput.n130 0.00340054
R13827 CSoutput.n133 CSoutput.n131 0.00340054
R13828 CSoutput.n262 CSoutput.n261 0.00340054
R13829 CSoutput.n257 CSoutput.n126 0.00340054
R13830 CSoutput.n142 CSoutput.n127 0.00340054
R13831 CSoutput.n145 CSoutput.n129 0.00340054
R13832 CSoutput.n175 CSoutput.n169 0.00252698
R13833 CSoutput.n168 CSoutput.n166 0.00252698
R13834 CSoutput.n250 CSoutput.n249 0.00252698
R13835 CSoutput.n178 CSoutput.n176 0.00252698
R13836 CSoutput.n181 CSoutput.n179 0.00252698
R13837 CSoutput.n254 CSoutput.n149 0.00252698
R13838 CSoutput.n175 CSoutput.n174 0.00252698
R13839 CSoutput.n168 CSoutput.n167 0.00252698
R13840 CSoutput.n251 CSoutput.n250 0.00252698
R13841 CSoutput.n178 CSoutput.n177 0.00252698
R13842 CSoutput.n181 CSoutput.n180 0.00252698
R13843 CSoutput.n162 CSoutput.n149 0.00252698
R13844 CSoutput.n229 CSoutput.n199 0.00252698
R13845 CSoutput.n228 CSoutput.n198 0.00252698
R13846 CSoutput.n227 CSoutput.n183 0.00252698
R13847 CSoutput.n224 CSoutput.n194 0.00252698
R13848 CSoutput.n231 CSoutput.n226 0.00252698
R13849 CSoutput.n240 CSoutput.n233 0.00252698
R13850 CSoutput.n229 CSoutput.n218 0.00252698
R13851 CSoutput.n228 CSoutput.n220 0.00252698
R13852 CSoutput.n227 CSoutput.n222 0.00252698
R13853 CSoutput.n242 CSoutput.n194 0.00252698
R13854 CSoutput.n231 CSoutput.n196 0.00252698
R13855 CSoutput.n233 CSoutput.n195 0.00252698
R13856 CSoutput.n141 CSoutput.n135 0.00252698
R13857 CSoutput.n134 CSoutput.n132 0.00252698
R13858 CSoutput.n260 CSoutput.n259 0.00252698
R13859 CSoutput.n144 CSoutput.n142 0.00252698
R13860 CSoutput.n147 CSoutput.n145 0.00252698
R13861 CSoutput.n264 CSoutput.n115 0.00252698
R13862 CSoutput.n141 CSoutput.n140 0.00252698
R13863 CSoutput.n134 CSoutput.n133 0.00252698
R13864 CSoutput.n261 CSoutput.n260 0.00252698
R13865 CSoutput.n144 CSoutput.n143 0.00252698
R13866 CSoutput.n147 CSoutput.n146 0.00252698
R13867 CSoutput.n128 CSoutput.n115 0.00252698
R13868 CSoutput.n249 CSoutput.n248 0.0020275
R13869 CSoutput.n248 CSoutput.n247 0.0020275
R13870 CSoutput.n245 CSoutput.n183 0.0020275
R13871 CSoutput.n245 CSoutput.n244 0.0020275
R13872 CSoutput.n259 CSoutput.n258 0.0020275
R13873 CSoutput.n258 CSoutput.n257 0.0020275
R13874 CSoutput.n159 CSoutput.n158 0.00166668
R13875 CSoutput.n241 CSoutput.n197 0.00166668
R13876 CSoutput.n125 CSoutput.n124 0.00166668
R13877 CSoutput.n263 CSoutput.n125 0.00133328
R13878 CSoutput.n197 CSoutput.n193 0.00133328
R13879 CSoutput.n253 CSoutput.n159 0.00133328
R13880 CSoutput.n256 CSoutput.n148 0.001
R13881 CSoutput.n234 CSoutput.n148 0.001
R13882 CSoutput.n136 CSoutput.n116 0.001
R13883 CSoutput.n235 CSoutput.n116 0.001
R13884 CSoutput.n137 CSoutput.n117 0.001
R13885 CSoutput.n236 CSoutput.n117 0.001
R13886 CSoutput.n138 CSoutput.n118 0.001
R13887 CSoutput.n237 CSoutput.n118 0.001
R13888 CSoutput.n139 CSoutput.n119 0.001
R13889 CSoutput.n238 CSoutput.n119 0.001
R13890 CSoutput.n232 CSoutput.n184 0.001
R13891 CSoutput.n232 CSoutput.n230 0.001
R13892 CSoutput.n214 CSoutput.n185 0.001
R13893 CSoutput.n208 CSoutput.n185 0.001
R13894 CSoutput.n215 CSoutput.n186 0.001
R13895 CSoutput.n209 CSoutput.n186 0.001
R13896 CSoutput.n216 CSoutput.n187 0.001
R13897 CSoutput.n210 CSoutput.n187 0.001
R13898 CSoutput.n217 CSoutput.n188 0.001
R13899 CSoutput.n211 CSoutput.n188 0.001
R13900 CSoutput.n246 CSoutput.n182 0.001
R13901 CSoutput.n200 CSoutput.n182 0.001
R13902 CSoutput.n170 CSoutput.n150 0.001
R13903 CSoutput.n201 CSoutput.n150 0.001
R13904 CSoutput.n171 CSoutput.n151 0.001
R13905 CSoutput.n202 CSoutput.n151 0.001
R13906 CSoutput.n172 CSoutput.n152 0.001
R13907 CSoutput.n203 CSoutput.n152 0.001
R13908 CSoutput.n173 CSoutput.n153 0.001
R13909 CSoutput.n204 CSoutput.n153 0.001
R13910 CSoutput.n204 CSoutput.n154 0.001
R13911 CSoutput.n203 CSoutput.n155 0.001
R13912 CSoutput.n202 CSoutput.n156 0.001
R13913 CSoutput.n201 CSoutput.t126 0.001
R13914 CSoutput.n200 CSoutput.n157 0.001
R13915 CSoutput.n173 CSoutput.n155 0.001
R13916 CSoutput.n172 CSoutput.n156 0.001
R13917 CSoutput.n171 CSoutput.t126 0.001
R13918 CSoutput.n170 CSoutput.n157 0.001
R13919 CSoutput.n246 CSoutput.n158 0.001
R13920 CSoutput.n211 CSoutput.n189 0.001
R13921 CSoutput.n210 CSoutput.n190 0.001
R13922 CSoutput.n209 CSoutput.n191 0.001
R13923 CSoutput.n208 CSoutput.t122 0.001
R13924 CSoutput.n230 CSoutput.n192 0.001
R13925 CSoutput.n217 CSoutput.n190 0.001
R13926 CSoutput.n216 CSoutput.n191 0.001
R13927 CSoutput.n215 CSoutput.t122 0.001
R13928 CSoutput.n214 CSoutput.n192 0.001
R13929 CSoutput.n241 CSoutput.n184 0.001
R13930 CSoutput.n238 CSoutput.n120 0.001
R13931 CSoutput.n237 CSoutput.n121 0.001
R13932 CSoutput.n236 CSoutput.n122 0.001
R13933 CSoutput.n235 CSoutput.t139 0.001
R13934 CSoutput.n234 CSoutput.n123 0.001
R13935 CSoutput.n139 CSoutput.n121 0.001
R13936 CSoutput.n138 CSoutput.n122 0.001
R13937 CSoutput.n137 CSoutput.t139 0.001
R13938 CSoutput.n136 CSoutput.n123 0.001
R13939 CSoutput.n256 CSoutput.n124 0.001
R13940 vdd.n303 vdd.n267 756.745
R13941 vdd.n252 vdd.n216 756.745
R13942 vdd.n209 vdd.n173 756.745
R13943 vdd.n158 vdd.n122 756.745
R13944 vdd.n116 vdd.n80 756.745
R13945 vdd.n65 vdd.n29 756.745
R13946 vdd.n1498 vdd.n1462 756.745
R13947 vdd.n1549 vdd.n1513 756.745
R13948 vdd.n1404 vdd.n1368 756.745
R13949 vdd.n1455 vdd.n1419 756.745
R13950 vdd.n1311 vdd.n1275 756.745
R13951 vdd.n1362 vdd.n1326 756.745
R13952 vdd.n1889 vdd.t129 640.208
R13953 vdd.n793 vdd.t114 640.208
R13954 vdd.n1863 vdd.t156 640.208
R13955 vdd.n785 vdd.t140 640.208
R13956 vdd.n2634 vdd.t101 640.208
R13957 vdd.n2354 vdd.t137 640.208
R13958 vdd.n661 vdd.t118 640.208
R13959 vdd.n2351 vdd.t122 640.208
R13960 vdd.n625 vdd.t126 640.208
R13961 vdd.n855 vdd.t133 640.208
R13962 vdd.n1110 vdd.t150 592.009
R13963 vdd.n1147 vdd.t97 592.009
R13964 vdd.n1021 vdd.t108 592.009
R13965 vdd.n2045 vdd.t93 592.009
R13966 vdd.n1682 vdd.t105 592.009
R13967 vdd.n1642 vdd.t111 592.009
R13968 vdd.n3021 vdd.t153 592.009
R13969 vdd.n427 vdd.t146 592.009
R13970 vdd.n387 vdd.t159 592.009
R13971 vdd.n580 vdd.t86 592.009
R13972 vdd.n543 vdd.t90 592.009
R13973 vdd.n2808 vdd.t143 592.009
R13974 vdd.n304 vdd.n303 585
R13975 vdd.n302 vdd.n269 585
R13976 vdd.n301 vdd.n300 585
R13977 vdd.n272 vdd.n270 585
R13978 vdd.n295 vdd.n294 585
R13979 vdd.n293 vdd.n292 585
R13980 vdd.n276 vdd.n275 585
R13981 vdd.n287 vdd.n286 585
R13982 vdd.n285 vdd.n284 585
R13983 vdd.n280 vdd.n279 585
R13984 vdd.n253 vdd.n252 585
R13985 vdd.n251 vdd.n218 585
R13986 vdd.n250 vdd.n249 585
R13987 vdd.n221 vdd.n219 585
R13988 vdd.n244 vdd.n243 585
R13989 vdd.n242 vdd.n241 585
R13990 vdd.n225 vdd.n224 585
R13991 vdd.n236 vdd.n235 585
R13992 vdd.n234 vdd.n233 585
R13993 vdd.n229 vdd.n228 585
R13994 vdd.n210 vdd.n209 585
R13995 vdd.n208 vdd.n175 585
R13996 vdd.n207 vdd.n206 585
R13997 vdd.n178 vdd.n176 585
R13998 vdd.n201 vdd.n200 585
R13999 vdd.n199 vdd.n198 585
R14000 vdd.n182 vdd.n181 585
R14001 vdd.n193 vdd.n192 585
R14002 vdd.n191 vdd.n190 585
R14003 vdd.n186 vdd.n185 585
R14004 vdd.n159 vdd.n158 585
R14005 vdd.n157 vdd.n124 585
R14006 vdd.n156 vdd.n155 585
R14007 vdd.n127 vdd.n125 585
R14008 vdd.n150 vdd.n149 585
R14009 vdd.n148 vdd.n147 585
R14010 vdd.n131 vdd.n130 585
R14011 vdd.n142 vdd.n141 585
R14012 vdd.n140 vdd.n139 585
R14013 vdd.n135 vdd.n134 585
R14014 vdd.n117 vdd.n116 585
R14015 vdd.n115 vdd.n82 585
R14016 vdd.n114 vdd.n113 585
R14017 vdd.n85 vdd.n83 585
R14018 vdd.n108 vdd.n107 585
R14019 vdd.n106 vdd.n105 585
R14020 vdd.n89 vdd.n88 585
R14021 vdd.n100 vdd.n99 585
R14022 vdd.n98 vdd.n97 585
R14023 vdd.n93 vdd.n92 585
R14024 vdd.n66 vdd.n65 585
R14025 vdd.n64 vdd.n31 585
R14026 vdd.n63 vdd.n62 585
R14027 vdd.n34 vdd.n32 585
R14028 vdd.n57 vdd.n56 585
R14029 vdd.n55 vdd.n54 585
R14030 vdd.n38 vdd.n37 585
R14031 vdd.n49 vdd.n48 585
R14032 vdd.n47 vdd.n46 585
R14033 vdd.n42 vdd.n41 585
R14034 vdd.n1499 vdd.n1498 585
R14035 vdd.n1497 vdd.n1464 585
R14036 vdd.n1496 vdd.n1495 585
R14037 vdd.n1467 vdd.n1465 585
R14038 vdd.n1490 vdd.n1489 585
R14039 vdd.n1488 vdd.n1487 585
R14040 vdd.n1471 vdd.n1470 585
R14041 vdd.n1482 vdd.n1481 585
R14042 vdd.n1480 vdd.n1479 585
R14043 vdd.n1475 vdd.n1474 585
R14044 vdd.n1550 vdd.n1549 585
R14045 vdd.n1548 vdd.n1515 585
R14046 vdd.n1547 vdd.n1546 585
R14047 vdd.n1518 vdd.n1516 585
R14048 vdd.n1541 vdd.n1540 585
R14049 vdd.n1539 vdd.n1538 585
R14050 vdd.n1522 vdd.n1521 585
R14051 vdd.n1533 vdd.n1532 585
R14052 vdd.n1531 vdd.n1530 585
R14053 vdd.n1526 vdd.n1525 585
R14054 vdd.n1405 vdd.n1404 585
R14055 vdd.n1403 vdd.n1370 585
R14056 vdd.n1402 vdd.n1401 585
R14057 vdd.n1373 vdd.n1371 585
R14058 vdd.n1396 vdd.n1395 585
R14059 vdd.n1394 vdd.n1393 585
R14060 vdd.n1377 vdd.n1376 585
R14061 vdd.n1388 vdd.n1387 585
R14062 vdd.n1386 vdd.n1385 585
R14063 vdd.n1381 vdd.n1380 585
R14064 vdd.n1456 vdd.n1455 585
R14065 vdd.n1454 vdd.n1421 585
R14066 vdd.n1453 vdd.n1452 585
R14067 vdd.n1424 vdd.n1422 585
R14068 vdd.n1447 vdd.n1446 585
R14069 vdd.n1445 vdd.n1444 585
R14070 vdd.n1428 vdd.n1427 585
R14071 vdd.n1439 vdd.n1438 585
R14072 vdd.n1437 vdd.n1436 585
R14073 vdd.n1432 vdd.n1431 585
R14074 vdd.n1312 vdd.n1311 585
R14075 vdd.n1310 vdd.n1277 585
R14076 vdd.n1309 vdd.n1308 585
R14077 vdd.n1280 vdd.n1278 585
R14078 vdd.n1303 vdd.n1302 585
R14079 vdd.n1301 vdd.n1300 585
R14080 vdd.n1284 vdd.n1283 585
R14081 vdd.n1295 vdd.n1294 585
R14082 vdd.n1293 vdd.n1292 585
R14083 vdd.n1288 vdd.n1287 585
R14084 vdd.n1363 vdd.n1362 585
R14085 vdd.n1361 vdd.n1328 585
R14086 vdd.n1360 vdd.n1359 585
R14087 vdd.n1331 vdd.n1329 585
R14088 vdd.n1354 vdd.n1353 585
R14089 vdd.n1352 vdd.n1351 585
R14090 vdd.n1335 vdd.n1334 585
R14091 vdd.n1346 vdd.n1345 585
R14092 vdd.n1344 vdd.n1343 585
R14093 vdd.n1339 vdd.n1338 585
R14094 vdd.n3137 vdd.n352 488.781
R14095 vdd.n3019 vdd.n350 488.781
R14096 vdd.n2941 vdd.n515 488.781
R14097 vdd.n2939 vdd.n517 488.781
R14098 vdd.n2040 vdd.n903 488.781
R14099 vdd.n2043 vdd.n2042 488.781
R14100 vdd.n1216 vdd.n981 488.781
R14101 vdd.n1214 vdd.n984 488.781
R14102 vdd.n281 vdd.t198 329.043
R14103 vdd.n230 vdd.t169 329.043
R14104 vdd.n187 vdd.t162 329.043
R14105 vdd.n136 vdd.t224 329.043
R14106 vdd.n94 vdd.t5 329.043
R14107 vdd.n43 vdd.t83 329.043
R14108 vdd.n1476 vdd.t9 329.043
R14109 vdd.n1527 vdd.t187 329.043
R14110 vdd.n1382 vdd.t219 329.043
R14111 vdd.n1433 vdd.t201 329.043
R14112 vdd.n1289 vdd.t84 329.043
R14113 vdd.n1340 vdd.t231 329.043
R14114 vdd.n1110 vdd.t152 319.788
R14115 vdd.n1147 vdd.t100 319.788
R14116 vdd.n1021 vdd.t110 319.788
R14117 vdd.n2045 vdd.t95 319.788
R14118 vdd.n1682 vdd.t106 319.788
R14119 vdd.n1642 vdd.t112 319.788
R14120 vdd.n3021 vdd.t154 319.788
R14121 vdd.n427 vdd.t148 319.788
R14122 vdd.n387 vdd.t160 319.788
R14123 vdd.n580 vdd.t89 319.788
R14124 vdd.n543 vdd.t92 319.788
R14125 vdd.n2808 vdd.t145 319.788
R14126 vdd.n1111 vdd.t151 303.69
R14127 vdd.n1148 vdd.t99 303.69
R14128 vdd.n1022 vdd.t109 303.69
R14129 vdd.n2046 vdd.t96 303.69
R14130 vdd.n1683 vdd.t107 303.69
R14131 vdd.n1643 vdd.t113 303.69
R14132 vdd.n3022 vdd.t155 303.69
R14133 vdd.n428 vdd.t149 303.69
R14134 vdd.n388 vdd.t161 303.69
R14135 vdd.n581 vdd.t88 303.69
R14136 vdd.n544 vdd.t91 303.69
R14137 vdd.n2809 vdd.t144 303.69
R14138 vdd.n2577 vdd.n741 297.074
R14139 vdd.n2770 vdd.n635 297.074
R14140 vdd.n2707 vdd.n632 297.074
R14141 vdd.n2500 vdd.n742 297.074
R14142 vdd.n2315 vdd.n782 297.074
R14143 vdd.n2246 vdd.n2245 297.074
R14144 vdd.n1992 vdd.n878 297.074
R14145 vdd.n2088 vdd.n876 297.074
R14146 vdd.n2686 vdd.n633 297.074
R14147 vdd.n2773 vdd.n2772 297.074
R14148 vdd.n2349 vdd.n743 297.074
R14149 vdd.n2575 vdd.n744 297.074
R14150 vdd.n2243 vdd.n791 297.074
R14151 vdd.n789 vdd.n764 297.074
R14152 vdd.n1929 vdd.n879 297.074
R14153 vdd.n2086 vdd.n880 297.074
R14154 vdd.n2688 vdd.n633 185
R14155 vdd.n2771 vdd.n633 185
R14156 vdd.n2690 vdd.n2689 185
R14157 vdd.n2689 vdd.n631 185
R14158 vdd.n2691 vdd.n667 185
R14159 vdd.n2701 vdd.n667 185
R14160 vdd.n2692 vdd.n676 185
R14161 vdd.n676 vdd.n674 185
R14162 vdd.n2694 vdd.n2693 185
R14163 vdd.n2695 vdd.n2694 185
R14164 vdd.n2647 vdd.n675 185
R14165 vdd.n675 vdd.n671 185
R14166 vdd.n2646 vdd.n2645 185
R14167 vdd.n2645 vdd.n2644 185
R14168 vdd.n678 vdd.n677 185
R14169 vdd.n679 vdd.n678 185
R14170 vdd.n2637 vdd.n2636 185
R14171 vdd.n2638 vdd.n2637 185
R14172 vdd.n2633 vdd.n688 185
R14173 vdd.n688 vdd.n685 185
R14174 vdd.n2632 vdd.n2631 185
R14175 vdd.n2631 vdd.n2630 185
R14176 vdd.n690 vdd.n689 185
R14177 vdd.n698 vdd.n690 185
R14178 vdd.n2623 vdd.n2622 185
R14179 vdd.n2624 vdd.n2623 185
R14180 vdd.n2621 vdd.n699 185
R14181 vdd.n2472 vdd.n699 185
R14182 vdd.n2620 vdd.n2619 185
R14183 vdd.n2619 vdd.n2618 185
R14184 vdd.n701 vdd.n700 185
R14185 vdd.n702 vdd.n701 185
R14186 vdd.n2611 vdd.n2610 185
R14187 vdd.n2612 vdd.n2611 185
R14188 vdd.n2609 vdd.n711 185
R14189 vdd.n711 vdd.n708 185
R14190 vdd.n2608 vdd.n2607 185
R14191 vdd.n2607 vdd.n2606 185
R14192 vdd.n713 vdd.n712 185
R14193 vdd.n721 vdd.n713 185
R14194 vdd.n2599 vdd.n2598 185
R14195 vdd.n2600 vdd.n2599 185
R14196 vdd.n2597 vdd.n722 185
R14197 vdd.n728 vdd.n722 185
R14198 vdd.n2596 vdd.n2595 185
R14199 vdd.n2595 vdd.n2594 185
R14200 vdd.n724 vdd.n723 185
R14201 vdd.n725 vdd.n724 185
R14202 vdd.n2587 vdd.n2586 185
R14203 vdd.n2588 vdd.n2587 185
R14204 vdd.n2585 vdd.n734 185
R14205 vdd.n2493 vdd.n734 185
R14206 vdd.n2584 vdd.n2583 185
R14207 vdd.n2583 vdd.n2582 185
R14208 vdd.n736 vdd.n735 185
R14209 vdd.t209 vdd.n736 185
R14210 vdd.n2575 vdd.n2574 185
R14211 vdd.n2576 vdd.n2575 185
R14212 vdd.n2573 vdd.n744 185
R14213 vdd.n2572 vdd.n2571 185
R14214 vdd.n746 vdd.n745 185
R14215 vdd.n2358 vdd.n2357 185
R14216 vdd.n2360 vdd.n2359 185
R14217 vdd.n2362 vdd.n2361 185
R14218 vdd.n2364 vdd.n2363 185
R14219 vdd.n2366 vdd.n2365 185
R14220 vdd.n2368 vdd.n2367 185
R14221 vdd.n2370 vdd.n2369 185
R14222 vdd.n2372 vdd.n2371 185
R14223 vdd.n2374 vdd.n2373 185
R14224 vdd.n2376 vdd.n2375 185
R14225 vdd.n2378 vdd.n2377 185
R14226 vdd.n2380 vdd.n2379 185
R14227 vdd.n2382 vdd.n2381 185
R14228 vdd.n2384 vdd.n2383 185
R14229 vdd.n2386 vdd.n2385 185
R14230 vdd.n2388 vdd.n2387 185
R14231 vdd.n2390 vdd.n2389 185
R14232 vdd.n2392 vdd.n2391 185
R14233 vdd.n2394 vdd.n2393 185
R14234 vdd.n2396 vdd.n2395 185
R14235 vdd.n2398 vdd.n2397 185
R14236 vdd.n2400 vdd.n2399 185
R14237 vdd.n2402 vdd.n2401 185
R14238 vdd.n2404 vdd.n2403 185
R14239 vdd.n2406 vdd.n2405 185
R14240 vdd.n2408 vdd.n2407 185
R14241 vdd.n2410 vdd.n2409 185
R14242 vdd.n2412 vdd.n2411 185
R14243 vdd.n2414 vdd.n2413 185
R14244 vdd.n2416 vdd.n2415 185
R14245 vdd.n2418 vdd.n2417 185
R14246 vdd.n2419 vdd.n2349 185
R14247 vdd.n2569 vdd.n2349 185
R14248 vdd.n2774 vdd.n2773 185
R14249 vdd.n2775 vdd.n624 185
R14250 vdd.n2777 vdd.n2776 185
R14251 vdd.n2779 vdd.n622 185
R14252 vdd.n2781 vdd.n2780 185
R14253 vdd.n2782 vdd.n621 185
R14254 vdd.n2784 vdd.n2783 185
R14255 vdd.n2786 vdd.n619 185
R14256 vdd.n2788 vdd.n2787 185
R14257 vdd.n2789 vdd.n618 185
R14258 vdd.n2791 vdd.n2790 185
R14259 vdd.n2793 vdd.n616 185
R14260 vdd.n2795 vdd.n2794 185
R14261 vdd.n2796 vdd.n615 185
R14262 vdd.n2798 vdd.n2797 185
R14263 vdd.n2800 vdd.n614 185
R14264 vdd.n2801 vdd.n611 185
R14265 vdd.n2804 vdd.n2803 185
R14266 vdd.n612 vdd.n610 185
R14267 vdd.n2660 vdd.n2659 185
R14268 vdd.n2662 vdd.n2661 185
R14269 vdd.n2664 vdd.n2656 185
R14270 vdd.n2666 vdd.n2665 185
R14271 vdd.n2667 vdd.n2655 185
R14272 vdd.n2669 vdd.n2668 185
R14273 vdd.n2671 vdd.n2653 185
R14274 vdd.n2673 vdd.n2672 185
R14275 vdd.n2674 vdd.n2652 185
R14276 vdd.n2676 vdd.n2675 185
R14277 vdd.n2678 vdd.n2650 185
R14278 vdd.n2680 vdd.n2679 185
R14279 vdd.n2681 vdd.n2649 185
R14280 vdd.n2683 vdd.n2682 185
R14281 vdd.n2685 vdd.n2648 185
R14282 vdd.n2687 vdd.n2686 185
R14283 vdd.n2686 vdd.n613 185
R14284 vdd.n2772 vdd.n628 185
R14285 vdd.n2772 vdd.n2771 185
R14286 vdd.n2424 vdd.n630 185
R14287 vdd.n631 vdd.n630 185
R14288 vdd.n2425 vdd.n666 185
R14289 vdd.n2701 vdd.n666 185
R14290 vdd.n2427 vdd.n2426 185
R14291 vdd.n2426 vdd.n674 185
R14292 vdd.n2428 vdd.n673 185
R14293 vdd.n2695 vdd.n673 185
R14294 vdd.n2430 vdd.n2429 185
R14295 vdd.n2429 vdd.n671 185
R14296 vdd.n2431 vdd.n681 185
R14297 vdd.n2644 vdd.n681 185
R14298 vdd.n2433 vdd.n2432 185
R14299 vdd.n2432 vdd.n679 185
R14300 vdd.n2434 vdd.n687 185
R14301 vdd.n2638 vdd.n687 185
R14302 vdd.n2436 vdd.n2435 185
R14303 vdd.n2435 vdd.n685 185
R14304 vdd.n2437 vdd.n692 185
R14305 vdd.n2630 vdd.n692 185
R14306 vdd.n2439 vdd.n2438 185
R14307 vdd.n2438 vdd.n698 185
R14308 vdd.n2440 vdd.n697 185
R14309 vdd.n2624 vdd.n697 185
R14310 vdd.n2474 vdd.n2473 185
R14311 vdd.n2473 vdd.n2472 185
R14312 vdd.n2475 vdd.n704 185
R14313 vdd.n2618 vdd.n704 185
R14314 vdd.n2477 vdd.n2476 185
R14315 vdd.n2476 vdd.n702 185
R14316 vdd.n2478 vdd.n710 185
R14317 vdd.n2612 vdd.n710 185
R14318 vdd.n2480 vdd.n2479 185
R14319 vdd.n2479 vdd.n708 185
R14320 vdd.n2481 vdd.n715 185
R14321 vdd.n2606 vdd.n715 185
R14322 vdd.n2483 vdd.n2482 185
R14323 vdd.n2482 vdd.n721 185
R14324 vdd.n2484 vdd.n720 185
R14325 vdd.n2600 vdd.n720 185
R14326 vdd.n2486 vdd.n2485 185
R14327 vdd.n2485 vdd.n728 185
R14328 vdd.n2487 vdd.n727 185
R14329 vdd.n2594 vdd.n727 185
R14330 vdd.n2489 vdd.n2488 185
R14331 vdd.n2488 vdd.n725 185
R14332 vdd.n2490 vdd.n733 185
R14333 vdd.n2588 vdd.n733 185
R14334 vdd.n2492 vdd.n2491 185
R14335 vdd.n2493 vdd.n2492 185
R14336 vdd.n2423 vdd.n738 185
R14337 vdd.n2582 vdd.n738 185
R14338 vdd.n2422 vdd.n2421 185
R14339 vdd.n2421 vdd.t209 185
R14340 vdd.n2420 vdd.n743 185
R14341 vdd.n2576 vdd.n743 185
R14342 vdd.n2040 vdd.n2039 185
R14343 vdd.n2041 vdd.n2040 185
R14344 vdd.n904 vdd.n902 185
R14345 vdd.n1606 vdd.n902 185
R14346 vdd.n1609 vdd.n1608 185
R14347 vdd.n1608 vdd.n1607 185
R14348 vdd.n907 vdd.n906 185
R14349 vdd.n908 vdd.n907 185
R14350 vdd.n1595 vdd.n1594 185
R14351 vdd.n1596 vdd.n1595 185
R14352 vdd.n916 vdd.n915 185
R14353 vdd.n1587 vdd.n915 185
R14354 vdd.n1590 vdd.n1589 185
R14355 vdd.n1589 vdd.n1588 185
R14356 vdd.n919 vdd.n918 185
R14357 vdd.n925 vdd.n919 185
R14358 vdd.n1578 vdd.n1577 185
R14359 vdd.n1579 vdd.n1578 185
R14360 vdd.n927 vdd.n926 185
R14361 vdd.n1570 vdd.n926 185
R14362 vdd.n1573 vdd.n1572 185
R14363 vdd.n1572 vdd.n1571 185
R14364 vdd.n930 vdd.n929 185
R14365 vdd.n931 vdd.n930 185
R14366 vdd.n1561 vdd.n1560 185
R14367 vdd.n1562 vdd.n1561 185
R14368 vdd.n939 vdd.n938 185
R14369 vdd.n938 vdd.n937 185
R14370 vdd.n1274 vdd.n1273 185
R14371 vdd.n1273 vdd.n1272 185
R14372 vdd.n942 vdd.n941 185
R14373 vdd.n948 vdd.n942 185
R14374 vdd.n1263 vdd.n1262 185
R14375 vdd.n1264 vdd.n1263 185
R14376 vdd.n950 vdd.n949 185
R14377 vdd.n1255 vdd.n949 185
R14378 vdd.n1258 vdd.n1257 185
R14379 vdd.n1257 vdd.n1256 185
R14380 vdd.n953 vdd.n952 185
R14381 vdd.n960 vdd.n953 185
R14382 vdd.n1246 vdd.n1245 185
R14383 vdd.n1247 vdd.n1246 185
R14384 vdd.n962 vdd.n961 185
R14385 vdd.n961 vdd.n959 185
R14386 vdd.n1241 vdd.n1240 185
R14387 vdd.n1240 vdd.n1239 185
R14388 vdd.n965 vdd.n964 185
R14389 vdd.n966 vdd.n965 185
R14390 vdd.n1230 vdd.n1229 185
R14391 vdd.n1231 vdd.n1230 185
R14392 vdd.n974 vdd.n973 185
R14393 vdd.n973 vdd.n972 185
R14394 vdd.n1225 vdd.n1224 185
R14395 vdd.n1224 vdd.n1223 185
R14396 vdd.n977 vdd.n976 185
R14397 vdd.n983 vdd.n977 185
R14398 vdd.n1214 vdd.n1213 185
R14399 vdd.n1215 vdd.n1214 185
R14400 vdd.n1210 vdd.n984 185
R14401 vdd.n1209 vdd.n987 185
R14402 vdd.n1208 vdd.n988 185
R14403 vdd.n988 vdd.n982 185
R14404 vdd.n991 vdd.n989 185
R14405 vdd.n1204 vdd.n993 185
R14406 vdd.n1203 vdd.n994 185
R14407 vdd.n1202 vdd.n996 185
R14408 vdd.n999 vdd.n997 185
R14409 vdd.n1198 vdd.n1001 185
R14410 vdd.n1197 vdd.n1002 185
R14411 vdd.n1196 vdd.n1004 185
R14412 vdd.n1007 vdd.n1005 185
R14413 vdd.n1192 vdd.n1009 185
R14414 vdd.n1191 vdd.n1010 185
R14415 vdd.n1190 vdd.n1012 185
R14416 vdd.n1015 vdd.n1013 185
R14417 vdd.n1186 vdd.n1017 185
R14418 vdd.n1185 vdd.n1018 185
R14419 vdd.n1184 vdd.n1020 185
R14420 vdd.n1025 vdd.n1023 185
R14421 vdd.n1180 vdd.n1027 185
R14422 vdd.n1179 vdd.n1028 185
R14423 vdd.n1178 vdd.n1030 185
R14424 vdd.n1033 vdd.n1031 185
R14425 vdd.n1174 vdd.n1035 185
R14426 vdd.n1173 vdd.n1036 185
R14427 vdd.n1172 vdd.n1038 185
R14428 vdd.n1041 vdd.n1039 185
R14429 vdd.n1168 vdd.n1043 185
R14430 vdd.n1167 vdd.n1044 185
R14431 vdd.n1166 vdd.n1046 185
R14432 vdd.n1049 vdd.n1047 185
R14433 vdd.n1162 vdd.n1051 185
R14434 vdd.n1161 vdd.n1052 185
R14435 vdd.n1160 vdd.n1054 185
R14436 vdd.n1057 vdd.n1055 185
R14437 vdd.n1156 vdd.n1059 185
R14438 vdd.n1155 vdd.n1060 185
R14439 vdd.n1154 vdd.n1062 185
R14440 vdd.n1065 vdd.n1063 185
R14441 vdd.n1150 vdd.n1067 185
R14442 vdd.n1149 vdd.n1146 185
R14443 vdd.n1144 vdd.n1068 185
R14444 vdd.n1143 vdd.n1142 185
R14445 vdd.n1073 vdd.n1070 185
R14446 vdd.n1138 vdd.n1074 185
R14447 vdd.n1137 vdd.n1076 185
R14448 vdd.n1136 vdd.n1077 185
R14449 vdd.n1081 vdd.n1078 185
R14450 vdd.n1132 vdd.n1082 185
R14451 vdd.n1131 vdd.n1084 185
R14452 vdd.n1130 vdd.n1085 185
R14453 vdd.n1089 vdd.n1086 185
R14454 vdd.n1126 vdd.n1090 185
R14455 vdd.n1125 vdd.n1092 185
R14456 vdd.n1124 vdd.n1093 185
R14457 vdd.n1097 vdd.n1094 185
R14458 vdd.n1120 vdd.n1098 185
R14459 vdd.n1119 vdd.n1100 185
R14460 vdd.n1118 vdd.n1101 185
R14461 vdd.n1105 vdd.n1102 185
R14462 vdd.n1114 vdd.n1106 185
R14463 vdd.n1113 vdd.n1108 185
R14464 vdd.n1109 vdd.n981 185
R14465 vdd.n982 vdd.n981 185
R14466 vdd.n2044 vdd.n2043 185
R14467 vdd.n2048 vdd.n897 185
R14468 vdd.n1711 vdd.n896 185
R14469 vdd.n1714 vdd.n1713 185
R14470 vdd.n1716 vdd.n1715 185
R14471 vdd.n1719 vdd.n1718 185
R14472 vdd.n1721 vdd.n1720 185
R14473 vdd.n1723 vdd.n1709 185
R14474 vdd.n1725 vdd.n1724 185
R14475 vdd.n1726 vdd.n1703 185
R14476 vdd.n1728 vdd.n1727 185
R14477 vdd.n1730 vdd.n1701 185
R14478 vdd.n1732 vdd.n1731 185
R14479 vdd.n1733 vdd.n1696 185
R14480 vdd.n1735 vdd.n1734 185
R14481 vdd.n1737 vdd.n1694 185
R14482 vdd.n1739 vdd.n1738 185
R14483 vdd.n1740 vdd.n1690 185
R14484 vdd.n1742 vdd.n1741 185
R14485 vdd.n1744 vdd.n1687 185
R14486 vdd.n1746 vdd.n1745 185
R14487 vdd.n1688 vdd.n1681 185
R14488 vdd.n1750 vdd.n1685 185
R14489 vdd.n1751 vdd.n1677 185
R14490 vdd.n1753 vdd.n1752 185
R14491 vdd.n1755 vdd.n1675 185
R14492 vdd.n1757 vdd.n1756 185
R14493 vdd.n1758 vdd.n1670 185
R14494 vdd.n1760 vdd.n1759 185
R14495 vdd.n1762 vdd.n1668 185
R14496 vdd.n1764 vdd.n1763 185
R14497 vdd.n1765 vdd.n1663 185
R14498 vdd.n1767 vdd.n1766 185
R14499 vdd.n1769 vdd.n1661 185
R14500 vdd.n1771 vdd.n1770 185
R14501 vdd.n1772 vdd.n1656 185
R14502 vdd.n1774 vdd.n1773 185
R14503 vdd.n1776 vdd.n1654 185
R14504 vdd.n1778 vdd.n1777 185
R14505 vdd.n1779 vdd.n1650 185
R14506 vdd.n1781 vdd.n1780 185
R14507 vdd.n1783 vdd.n1647 185
R14508 vdd.n1785 vdd.n1784 185
R14509 vdd.n1648 vdd.n1641 185
R14510 vdd.n1789 vdd.n1645 185
R14511 vdd.n1790 vdd.n1637 185
R14512 vdd.n1792 vdd.n1791 185
R14513 vdd.n1794 vdd.n1635 185
R14514 vdd.n1796 vdd.n1795 185
R14515 vdd.n1797 vdd.n1630 185
R14516 vdd.n1799 vdd.n1798 185
R14517 vdd.n1801 vdd.n1628 185
R14518 vdd.n1803 vdd.n1802 185
R14519 vdd.n1804 vdd.n1623 185
R14520 vdd.n1806 vdd.n1805 185
R14521 vdd.n1808 vdd.n1622 185
R14522 vdd.n1809 vdd.n1619 185
R14523 vdd.n1812 vdd.n1811 185
R14524 vdd.n1621 vdd.n1617 185
R14525 vdd.n2029 vdd.n1615 185
R14526 vdd.n2031 vdd.n2030 185
R14527 vdd.n2033 vdd.n1613 185
R14528 vdd.n2035 vdd.n2034 185
R14529 vdd.n2036 vdd.n903 185
R14530 vdd.n2042 vdd.n900 185
R14531 vdd.n2042 vdd.n2041 185
R14532 vdd.n911 vdd.n899 185
R14533 vdd.n1606 vdd.n899 185
R14534 vdd.n1605 vdd.n1604 185
R14535 vdd.n1607 vdd.n1605 185
R14536 vdd.n910 vdd.n909 185
R14537 vdd.n909 vdd.n908 185
R14538 vdd.n1598 vdd.n1597 185
R14539 vdd.n1597 vdd.n1596 185
R14540 vdd.n914 vdd.n913 185
R14541 vdd.n1587 vdd.n914 185
R14542 vdd.n1586 vdd.n1585 185
R14543 vdd.n1588 vdd.n1586 185
R14544 vdd.n921 vdd.n920 185
R14545 vdd.n925 vdd.n920 185
R14546 vdd.n1581 vdd.n1580 185
R14547 vdd.n1580 vdd.n1579 185
R14548 vdd.n924 vdd.n923 185
R14549 vdd.n1570 vdd.n924 185
R14550 vdd.n1569 vdd.n1568 185
R14551 vdd.n1571 vdd.n1569 185
R14552 vdd.n933 vdd.n932 185
R14553 vdd.n932 vdd.n931 185
R14554 vdd.n1564 vdd.n1563 185
R14555 vdd.n1563 vdd.n1562 185
R14556 vdd.n936 vdd.n935 185
R14557 vdd.n937 vdd.n936 185
R14558 vdd.n1271 vdd.n1270 185
R14559 vdd.n1272 vdd.n1271 185
R14560 vdd.n944 vdd.n943 185
R14561 vdd.n948 vdd.n943 185
R14562 vdd.n1266 vdd.n1265 185
R14563 vdd.n1265 vdd.n1264 185
R14564 vdd.n947 vdd.n946 185
R14565 vdd.n1255 vdd.n947 185
R14566 vdd.n1254 vdd.n1253 185
R14567 vdd.n1256 vdd.n1254 185
R14568 vdd.n955 vdd.n954 185
R14569 vdd.n960 vdd.n954 185
R14570 vdd.n1249 vdd.n1248 185
R14571 vdd.n1248 vdd.n1247 185
R14572 vdd.n958 vdd.n957 185
R14573 vdd.n959 vdd.n958 185
R14574 vdd.n1238 vdd.n1237 185
R14575 vdd.n1239 vdd.n1238 185
R14576 vdd.n968 vdd.n967 185
R14577 vdd.n967 vdd.n966 185
R14578 vdd.n1233 vdd.n1232 185
R14579 vdd.n1232 vdd.n1231 185
R14580 vdd.n971 vdd.n970 185
R14581 vdd.n972 vdd.n971 185
R14582 vdd.n1222 vdd.n1221 185
R14583 vdd.n1223 vdd.n1222 185
R14584 vdd.n979 vdd.n978 185
R14585 vdd.n983 vdd.n978 185
R14586 vdd.n1217 vdd.n1216 185
R14587 vdd.n1216 vdd.n1215 185
R14588 vdd.n784 vdd.n782 185
R14589 vdd.n2244 vdd.n782 185
R14590 vdd.n2166 vdd.n801 185
R14591 vdd.n801 vdd.t182 185
R14592 vdd.n2168 vdd.n2167 185
R14593 vdd.n2169 vdd.n2168 185
R14594 vdd.n2165 vdd.n800 185
R14595 vdd.n1868 vdd.n800 185
R14596 vdd.n2164 vdd.n2163 185
R14597 vdd.n2163 vdd.n2162 185
R14598 vdd.n803 vdd.n802 185
R14599 vdd.n804 vdd.n803 185
R14600 vdd.n2153 vdd.n2152 185
R14601 vdd.n2154 vdd.n2153 185
R14602 vdd.n2151 vdd.n814 185
R14603 vdd.n814 vdd.n811 185
R14604 vdd.n2150 vdd.n2149 185
R14605 vdd.n2149 vdd.n2148 185
R14606 vdd.n816 vdd.n815 185
R14607 vdd.n817 vdd.n816 185
R14608 vdd.n2141 vdd.n2140 185
R14609 vdd.n2142 vdd.n2141 185
R14610 vdd.n2139 vdd.n825 185
R14611 vdd.n830 vdd.n825 185
R14612 vdd.n2138 vdd.n2137 185
R14613 vdd.n2137 vdd.n2136 185
R14614 vdd.n827 vdd.n826 185
R14615 vdd.n836 vdd.n827 185
R14616 vdd.n2129 vdd.n2128 185
R14617 vdd.n2130 vdd.n2129 185
R14618 vdd.n2127 vdd.n837 185
R14619 vdd.n1969 vdd.n837 185
R14620 vdd.n2126 vdd.n2125 185
R14621 vdd.n2125 vdd.n2124 185
R14622 vdd.n839 vdd.n838 185
R14623 vdd.n840 vdd.n839 185
R14624 vdd.n2117 vdd.n2116 185
R14625 vdd.n2118 vdd.n2117 185
R14626 vdd.n2115 vdd.n849 185
R14627 vdd.n849 vdd.n846 185
R14628 vdd.n2114 vdd.n2113 185
R14629 vdd.n2113 vdd.n2112 185
R14630 vdd.n851 vdd.n850 185
R14631 vdd.n861 vdd.n851 185
R14632 vdd.n2104 vdd.n2103 185
R14633 vdd.n2105 vdd.n2104 185
R14634 vdd.n2102 vdd.n862 185
R14635 vdd.n862 vdd.n858 185
R14636 vdd.n2101 vdd.n2100 185
R14637 vdd.n2100 vdd.n2099 185
R14638 vdd.n864 vdd.n863 185
R14639 vdd.n865 vdd.n864 185
R14640 vdd.n2092 vdd.n2091 185
R14641 vdd.n2093 vdd.n2092 185
R14642 vdd.n2090 vdd.n874 185
R14643 vdd.n874 vdd.n871 185
R14644 vdd.n2089 vdd.n2088 185
R14645 vdd.n2088 vdd.n2087 185
R14646 vdd.n876 vdd.n875 185
R14647 vdd.n1824 vdd.n1823 185
R14648 vdd.n1825 vdd.n1821 185
R14649 vdd.n1821 vdd.n877 185
R14650 vdd.n1827 vdd.n1826 185
R14651 vdd.n1829 vdd.n1820 185
R14652 vdd.n1832 vdd.n1831 185
R14653 vdd.n1833 vdd.n1819 185
R14654 vdd.n1835 vdd.n1834 185
R14655 vdd.n1837 vdd.n1818 185
R14656 vdd.n1840 vdd.n1839 185
R14657 vdd.n1841 vdd.n1817 185
R14658 vdd.n1843 vdd.n1842 185
R14659 vdd.n1845 vdd.n1816 185
R14660 vdd.n1848 vdd.n1847 185
R14661 vdd.n1849 vdd.n1815 185
R14662 vdd.n1851 vdd.n1850 185
R14663 vdd.n1853 vdd.n1814 185
R14664 vdd.n2026 vdd.n1854 185
R14665 vdd.n2025 vdd.n2024 185
R14666 vdd.n2022 vdd.n1855 185
R14667 vdd.n2020 vdd.n2019 185
R14668 vdd.n2018 vdd.n1856 185
R14669 vdd.n2017 vdd.n2016 185
R14670 vdd.n2014 vdd.n1857 185
R14671 vdd.n2012 vdd.n2011 185
R14672 vdd.n2010 vdd.n1858 185
R14673 vdd.n2009 vdd.n2008 185
R14674 vdd.n2006 vdd.n1859 185
R14675 vdd.n2004 vdd.n2003 185
R14676 vdd.n2002 vdd.n1860 185
R14677 vdd.n2001 vdd.n2000 185
R14678 vdd.n1998 vdd.n1861 185
R14679 vdd.n1996 vdd.n1995 185
R14680 vdd.n1994 vdd.n1862 185
R14681 vdd.n1993 vdd.n1992 185
R14682 vdd.n2247 vdd.n2246 185
R14683 vdd.n2249 vdd.n2248 185
R14684 vdd.n2251 vdd.n2250 185
R14685 vdd.n2254 vdd.n2253 185
R14686 vdd.n2256 vdd.n2255 185
R14687 vdd.n2258 vdd.n2257 185
R14688 vdd.n2260 vdd.n2259 185
R14689 vdd.n2262 vdd.n2261 185
R14690 vdd.n2264 vdd.n2263 185
R14691 vdd.n2266 vdd.n2265 185
R14692 vdd.n2268 vdd.n2267 185
R14693 vdd.n2270 vdd.n2269 185
R14694 vdd.n2272 vdd.n2271 185
R14695 vdd.n2274 vdd.n2273 185
R14696 vdd.n2276 vdd.n2275 185
R14697 vdd.n2278 vdd.n2277 185
R14698 vdd.n2280 vdd.n2279 185
R14699 vdd.n2282 vdd.n2281 185
R14700 vdd.n2284 vdd.n2283 185
R14701 vdd.n2286 vdd.n2285 185
R14702 vdd.n2288 vdd.n2287 185
R14703 vdd.n2290 vdd.n2289 185
R14704 vdd.n2292 vdd.n2291 185
R14705 vdd.n2294 vdd.n2293 185
R14706 vdd.n2296 vdd.n2295 185
R14707 vdd.n2298 vdd.n2297 185
R14708 vdd.n2300 vdd.n2299 185
R14709 vdd.n2302 vdd.n2301 185
R14710 vdd.n2304 vdd.n2303 185
R14711 vdd.n2306 vdd.n2305 185
R14712 vdd.n2308 vdd.n2307 185
R14713 vdd.n2310 vdd.n2309 185
R14714 vdd.n2312 vdd.n2311 185
R14715 vdd.n2313 vdd.n783 185
R14716 vdd.n2315 vdd.n2314 185
R14717 vdd.n2316 vdd.n2315 185
R14718 vdd.n2245 vdd.n787 185
R14719 vdd.n2245 vdd.n2244 185
R14720 vdd.n1866 vdd.n788 185
R14721 vdd.t182 vdd.n788 185
R14722 vdd.n1867 vdd.n798 185
R14723 vdd.n2169 vdd.n798 185
R14724 vdd.n1870 vdd.n1869 185
R14725 vdd.n1869 vdd.n1868 185
R14726 vdd.n1871 vdd.n805 185
R14727 vdd.n2162 vdd.n805 185
R14728 vdd.n1873 vdd.n1872 185
R14729 vdd.n1872 vdd.n804 185
R14730 vdd.n1874 vdd.n812 185
R14731 vdd.n2154 vdd.n812 185
R14732 vdd.n1876 vdd.n1875 185
R14733 vdd.n1875 vdd.n811 185
R14734 vdd.n1877 vdd.n818 185
R14735 vdd.n2148 vdd.n818 185
R14736 vdd.n1879 vdd.n1878 185
R14737 vdd.n1878 vdd.n817 185
R14738 vdd.n1880 vdd.n823 185
R14739 vdd.n2142 vdd.n823 185
R14740 vdd.n1882 vdd.n1881 185
R14741 vdd.n1881 vdd.n830 185
R14742 vdd.n1883 vdd.n828 185
R14743 vdd.n2136 vdd.n828 185
R14744 vdd.n1885 vdd.n1884 185
R14745 vdd.n1884 vdd.n836 185
R14746 vdd.n1886 vdd.n834 185
R14747 vdd.n2130 vdd.n834 185
R14748 vdd.n1971 vdd.n1970 185
R14749 vdd.n1970 vdd.n1969 185
R14750 vdd.n1972 vdd.n841 185
R14751 vdd.n2124 vdd.n841 185
R14752 vdd.n1974 vdd.n1973 185
R14753 vdd.n1973 vdd.n840 185
R14754 vdd.n1975 vdd.n847 185
R14755 vdd.n2118 vdd.n847 185
R14756 vdd.n1977 vdd.n1976 185
R14757 vdd.n1976 vdd.n846 185
R14758 vdd.n1978 vdd.n852 185
R14759 vdd.n2112 vdd.n852 185
R14760 vdd.n1980 vdd.n1979 185
R14761 vdd.n1979 vdd.n861 185
R14762 vdd.n1981 vdd.n859 185
R14763 vdd.n2105 vdd.n859 185
R14764 vdd.n1983 vdd.n1982 185
R14765 vdd.n1982 vdd.n858 185
R14766 vdd.n1984 vdd.n866 185
R14767 vdd.n2099 vdd.n866 185
R14768 vdd.n1986 vdd.n1985 185
R14769 vdd.n1985 vdd.n865 185
R14770 vdd.n1987 vdd.n872 185
R14771 vdd.n2093 vdd.n872 185
R14772 vdd.n1989 vdd.n1988 185
R14773 vdd.n1988 vdd.n871 185
R14774 vdd.n1990 vdd.n878 185
R14775 vdd.n2087 vdd.n878 185
R14776 vdd.n3137 vdd.n3136 185
R14777 vdd.n3138 vdd.n3137 185
R14778 vdd.n347 vdd.n346 185
R14779 vdd.n3139 vdd.n347 185
R14780 vdd.n3142 vdd.n3141 185
R14781 vdd.n3141 vdd.n3140 185
R14782 vdd.n3143 vdd.n341 185
R14783 vdd.n341 vdd.n340 185
R14784 vdd.n3145 vdd.n3144 185
R14785 vdd.n3146 vdd.n3145 185
R14786 vdd.n336 vdd.n335 185
R14787 vdd.n3147 vdd.n336 185
R14788 vdd.n3150 vdd.n3149 185
R14789 vdd.n3149 vdd.n3148 185
R14790 vdd.n3151 vdd.n330 185
R14791 vdd.n330 vdd.n329 185
R14792 vdd.n3153 vdd.n3152 185
R14793 vdd.n3154 vdd.n3153 185
R14794 vdd.n324 vdd.n323 185
R14795 vdd.n3155 vdd.n324 185
R14796 vdd.n3158 vdd.n3157 185
R14797 vdd.n3157 vdd.n3156 185
R14798 vdd.n3159 vdd.n319 185
R14799 vdd.n325 vdd.n319 185
R14800 vdd.n3161 vdd.n3160 185
R14801 vdd.n3162 vdd.n3161 185
R14802 vdd.n315 vdd.n313 185
R14803 vdd.n3163 vdd.n315 185
R14804 vdd.n3166 vdd.n3165 185
R14805 vdd.n3165 vdd.n3164 185
R14806 vdd.n314 vdd.n312 185
R14807 vdd.n481 vdd.n314 185
R14808 vdd.n2988 vdd.n2987 185
R14809 vdd.n2989 vdd.n2988 185
R14810 vdd.n483 vdd.n482 185
R14811 vdd.n2980 vdd.n482 185
R14812 vdd.n2983 vdd.n2982 185
R14813 vdd.n2982 vdd.n2981 185
R14814 vdd.n486 vdd.n485 185
R14815 vdd.n493 vdd.n486 185
R14816 vdd.n2971 vdd.n2970 185
R14817 vdd.n2972 vdd.n2971 185
R14818 vdd.n495 vdd.n494 185
R14819 vdd.n494 vdd.n492 185
R14820 vdd.n2966 vdd.n2965 185
R14821 vdd.n2965 vdd.n2964 185
R14822 vdd.n498 vdd.n497 185
R14823 vdd.n499 vdd.n498 185
R14824 vdd.n2955 vdd.n2954 185
R14825 vdd.n2956 vdd.n2955 185
R14826 vdd.n507 vdd.n506 185
R14827 vdd.n506 vdd.n505 185
R14828 vdd.n2950 vdd.n2949 185
R14829 vdd.n2949 vdd.n2948 185
R14830 vdd.n510 vdd.n509 185
R14831 vdd.n511 vdd.n510 185
R14832 vdd.n2939 vdd.n2938 185
R14833 vdd.n2940 vdd.n2939 185
R14834 vdd.n2935 vdd.n517 185
R14835 vdd.n2934 vdd.n2933 185
R14836 vdd.n2931 vdd.n519 185
R14837 vdd.n2931 vdd.n516 185
R14838 vdd.n2930 vdd.n2929 185
R14839 vdd.n2928 vdd.n2927 185
R14840 vdd.n2926 vdd.n2925 185
R14841 vdd.n2924 vdd.n2923 185
R14842 vdd.n2922 vdd.n525 185
R14843 vdd.n2920 vdd.n2919 185
R14844 vdd.n2918 vdd.n526 185
R14845 vdd.n2917 vdd.n2916 185
R14846 vdd.n2914 vdd.n531 185
R14847 vdd.n2912 vdd.n2911 185
R14848 vdd.n2910 vdd.n532 185
R14849 vdd.n2909 vdd.n2908 185
R14850 vdd.n2906 vdd.n537 185
R14851 vdd.n2904 vdd.n2903 185
R14852 vdd.n2902 vdd.n538 185
R14853 vdd.n2901 vdd.n2900 185
R14854 vdd.n2898 vdd.n545 185
R14855 vdd.n2896 vdd.n2895 185
R14856 vdd.n2894 vdd.n546 185
R14857 vdd.n2893 vdd.n2892 185
R14858 vdd.n2890 vdd.n551 185
R14859 vdd.n2888 vdd.n2887 185
R14860 vdd.n2886 vdd.n552 185
R14861 vdd.n2885 vdd.n2884 185
R14862 vdd.n2882 vdd.n557 185
R14863 vdd.n2880 vdd.n2879 185
R14864 vdd.n2878 vdd.n558 185
R14865 vdd.n2877 vdd.n2876 185
R14866 vdd.n2874 vdd.n563 185
R14867 vdd.n2872 vdd.n2871 185
R14868 vdd.n2870 vdd.n564 185
R14869 vdd.n2869 vdd.n2868 185
R14870 vdd.n2866 vdd.n569 185
R14871 vdd.n2864 vdd.n2863 185
R14872 vdd.n2862 vdd.n570 185
R14873 vdd.n2861 vdd.n2860 185
R14874 vdd.n2858 vdd.n575 185
R14875 vdd.n2856 vdd.n2855 185
R14876 vdd.n2854 vdd.n576 185
R14877 vdd.n585 vdd.n579 185
R14878 vdd.n2850 vdd.n2849 185
R14879 vdd.n2847 vdd.n583 185
R14880 vdd.n2846 vdd.n2845 185
R14881 vdd.n2844 vdd.n2843 185
R14882 vdd.n2842 vdd.n589 185
R14883 vdd.n2840 vdd.n2839 185
R14884 vdd.n2838 vdd.n590 185
R14885 vdd.n2837 vdd.n2836 185
R14886 vdd.n2834 vdd.n595 185
R14887 vdd.n2832 vdd.n2831 185
R14888 vdd.n2830 vdd.n596 185
R14889 vdd.n2829 vdd.n2828 185
R14890 vdd.n2826 vdd.n601 185
R14891 vdd.n2824 vdd.n2823 185
R14892 vdd.n2822 vdd.n602 185
R14893 vdd.n2821 vdd.n2820 185
R14894 vdd.n2818 vdd.n2817 185
R14895 vdd.n2816 vdd.n2815 185
R14896 vdd.n2814 vdd.n2813 185
R14897 vdd.n2812 vdd.n2811 185
R14898 vdd.n2807 vdd.n515 185
R14899 vdd.n516 vdd.n515 185
R14900 vdd.n3020 vdd.n3019 185
R14901 vdd.n3024 vdd.n462 185
R14902 vdd.n3026 vdd.n3025 185
R14903 vdd.n3028 vdd.n460 185
R14904 vdd.n3030 vdd.n3029 185
R14905 vdd.n3031 vdd.n455 185
R14906 vdd.n3033 vdd.n3032 185
R14907 vdd.n3035 vdd.n453 185
R14908 vdd.n3037 vdd.n3036 185
R14909 vdd.n3038 vdd.n448 185
R14910 vdd.n3040 vdd.n3039 185
R14911 vdd.n3042 vdd.n446 185
R14912 vdd.n3044 vdd.n3043 185
R14913 vdd.n3045 vdd.n441 185
R14914 vdd.n3047 vdd.n3046 185
R14915 vdd.n3049 vdd.n439 185
R14916 vdd.n3051 vdd.n3050 185
R14917 vdd.n3052 vdd.n435 185
R14918 vdd.n3054 vdd.n3053 185
R14919 vdd.n3056 vdd.n432 185
R14920 vdd.n3058 vdd.n3057 185
R14921 vdd.n433 vdd.n426 185
R14922 vdd.n3062 vdd.n430 185
R14923 vdd.n3063 vdd.n422 185
R14924 vdd.n3065 vdd.n3064 185
R14925 vdd.n3067 vdd.n420 185
R14926 vdd.n3069 vdd.n3068 185
R14927 vdd.n3070 vdd.n415 185
R14928 vdd.n3072 vdd.n3071 185
R14929 vdd.n3074 vdd.n413 185
R14930 vdd.n3076 vdd.n3075 185
R14931 vdd.n3077 vdd.n408 185
R14932 vdd.n3079 vdd.n3078 185
R14933 vdd.n3081 vdd.n406 185
R14934 vdd.n3083 vdd.n3082 185
R14935 vdd.n3084 vdd.n401 185
R14936 vdd.n3086 vdd.n3085 185
R14937 vdd.n3088 vdd.n399 185
R14938 vdd.n3090 vdd.n3089 185
R14939 vdd.n3091 vdd.n395 185
R14940 vdd.n3093 vdd.n3092 185
R14941 vdd.n3095 vdd.n392 185
R14942 vdd.n3097 vdd.n3096 185
R14943 vdd.n393 vdd.n386 185
R14944 vdd.n3101 vdd.n390 185
R14945 vdd.n3102 vdd.n382 185
R14946 vdd.n3104 vdd.n3103 185
R14947 vdd.n3106 vdd.n380 185
R14948 vdd.n3108 vdd.n3107 185
R14949 vdd.n3109 vdd.n375 185
R14950 vdd.n3111 vdd.n3110 185
R14951 vdd.n3113 vdd.n373 185
R14952 vdd.n3115 vdd.n3114 185
R14953 vdd.n3116 vdd.n368 185
R14954 vdd.n3118 vdd.n3117 185
R14955 vdd.n3120 vdd.n366 185
R14956 vdd.n3122 vdd.n3121 185
R14957 vdd.n3123 vdd.n360 185
R14958 vdd.n3125 vdd.n3124 185
R14959 vdd.n3127 vdd.n359 185
R14960 vdd.n3128 vdd.n358 185
R14961 vdd.n3131 vdd.n3130 185
R14962 vdd.n3132 vdd.n356 185
R14963 vdd.n3133 vdd.n352 185
R14964 vdd.n3015 vdd.n350 185
R14965 vdd.n3138 vdd.n350 185
R14966 vdd.n3014 vdd.n349 185
R14967 vdd.n3139 vdd.n349 185
R14968 vdd.n3013 vdd.n348 185
R14969 vdd.n3140 vdd.n348 185
R14970 vdd.n468 vdd.n467 185
R14971 vdd.n467 vdd.n340 185
R14972 vdd.n3009 vdd.n339 185
R14973 vdd.n3146 vdd.n339 185
R14974 vdd.n3008 vdd.n338 185
R14975 vdd.n3147 vdd.n338 185
R14976 vdd.n3007 vdd.n337 185
R14977 vdd.n3148 vdd.n337 185
R14978 vdd.n471 vdd.n470 185
R14979 vdd.n470 vdd.n329 185
R14980 vdd.n3003 vdd.n328 185
R14981 vdd.n3154 vdd.n328 185
R14982 vdd.n3002 vdd.n327 185
R14983 vdd.n3155 vdd.n327 185
R14984 vdd.n3001 vdd.n326 185
R14985 vdd.n3156 vdd.n326 185
R14986 vdd.n474 vdd.n473 185
R14987 vdd.n473 vdd.n325 185
R14988 vdd.n2997 vdd.n318 185
R14989 vdd.n3162 vdd.n318 185
R14990 vdd.n2996 vdd.n317 185
R14991 vdd.n3163 vdd.n317 185
R14992 vdd.n2995 vdd.n316 185
R14993 vdd.n3164 vdd.n316 185
R14994 vdd.n480 vdd.n476 185
R14995 vdd.n481 vdd.n480 185
R14996 vdd.n2991 vdd.n2990 185
R14997 vdd.n2990 vdd.n2989 185
R14998 vdd.n479 vdd.n478 185
R14999 vdd.n2980 vdd.n479 185
R15000 vdd.n2979 vdd.n2978 185
R15001 vdd.n2981 vdd.n2979 185
R15002 vdd.n488 vdd.n487 185
R15003 vdd.n493 vdd.n487 185
R15004 vdd.n2974 vdd.n2973 185
R15005 vdd.n2973 vdd.n2972 185
R15006 vdd.n491 vdd.n490 185
R15007 vdd.n492 vdd.n491 185
R15008 vdd.n2963 vdd.n2962 185
R15009 vdd.n2964 vdd.n2963 185
R15010 vdd.n501 vdd.n500 185
R15011 vdd.n500 vdd.n499 185
R15012 vdd.n2958 vdd.n2957 185
R15013 vdd.n2957 vdd.n2956 185
R15014 vdd.n504 vdd.n503 185
R15015 vdd.n505 vdd.n504 185
R15016 vdd.n2947 vdd.n2946 185
R15017 vdd.n2948 vdd.n2947 185
R15018 vdd.n513 vdd.n512 185
R15019 vdd.n512 vdd.n511 185
R15020 vdd.n2942 vdd.n2941 185
R15021 vdd.n2941 vdd.n2940 185
R15022 vdd.n741 vdd.n740 185
R15023 vdd.n2567 vdd.n2566 185
R15024 vdd.n2565 vdd.n2350 185
R15025 vdd.n2569 vdd.n2350 185
R15026 vdd.n2564 vdd.n2563 185
R15027 vdd.n2562 vdd.n2561 185
R15028 vdd.n2560 vdd.n2559 185
R15029 vdd.n2558 vdd.n2557 185
R15030 vdd.n2556 vdd.n2555 185
R15031 vdd.n2554 vdd.n2553 185
R15032 vdd.n2552 vdd.n2551 185
R15033 vdd.n2550 vdd.n2549 185
R15034 vdd.n2548 vdd.n2547 185
R15035 vdd.n2546 vdd.n2545 185
R15036 vdd.n2544 vdd.n2543 185
R15037 vdd.n2542 vdd.n2541 185
R15038 vdd.n2540 vdd.n2539 185
R15039 vdd.n2538 vdd.n2537 185
R15040 vdd.n2536 vdd.n2535 185
R15041 vdd.n2534 vdd.n2533 185
R15042 vdd.n2532 vdd.n2531 185
R15043 vdd.n2530 vdd.n2529 185
R15044 vdd.n2528 vdd.n2527 185
R15045 vdd.n2526 vdd.n2525 185
R15046 vdd.n2524 vdd.n2523 185
R15047 vdd.n2522 vdd.n2521 185
R15048 vdd.n2520 vdd.n2519 185
R15049 vdd.n2518 vdd.n2517 185
R15050 vdd.n2516 vdd.n2515 185
R15051 vdd.n2514 vdd.n2513 185
R15052 vdd.n2512 vdd.n2511 185
R15053 vdd.n2510 vdd.n2509 185
R15054 vdd.n2508 vdd.n2507 185
R15055 vdd.n2505 vdd.n2504 185
R15056 vdd.n2503 vdd.n2502 185
R15057 vdd.n2501 vdd.n2500 185
R15058 vdd.n2708 vdd.n2707 185
R15059 vdd.n2709 vdd.n660 185
R15060 vdd.n2711 vdd.n2710 185
R15061 vdd.n2713 vdd.n658 185
R15062 vdd.n2715 vdd.n2714 185
R15063 vdd.n2716 vdd.n657 185
R15064 vdd.n2718 vdd.n2717 185
R15065 vdd.n2720 vdd.n655 185
R15066 vdd.n2722 vdd.n2721 185
R15067 vdd.n2723 vdd.n654 185
R15068 vdd.n2725 vdd.n2724 185
R15069 vdd.n2727 vdd.n652 185
R15070 vdd.n2729 vdd.n2728 185
R15071 vdd.n2730 vdd.n651 185
R15072 vdd.n2732 vdd.n2731 185
R15073 vdd.n2734 vdd.n649 185
R15074 vdd.n2736 vdd.n2735 185
R15075 vdd.n2738 vdd.n648 185
R15076 vdd.n2740 vdd.n2739 185
R15077 vdd.n2742 vdd.n646 185
R15078 vdd.n2744 vdd.n2743 185
R15079 vdd.n2745 vdd.n645 185
R15080 vdd.n2747 vdd.n2746 185
R15081 vdd.n2749 vdd.n643 185
R15082 vdd.n2751 vdd.n2750 185
R15083 vdd.n2752 vdd.n642 185
R15084 vdd.n2754 vdd.n2753 185
R15085 vdd.n2756 vdd.n640 185
R15086 vdd.n2758 vdd.n2757 185
R15087 vdd.n2759 vdd.n639 185
R15088 vdd.n2761 vdd.n2760 185
R15089 vdd.n2763 vdd.n638 185
R15090 vdd.n2764 vdd.n637 185
R15091 vdd.n2767 vdd.n2766 185
R15092 vdd.n2768 vdd.n635 185
R15093 vdd.n635 vdd.n613 185
R15094 vdd.n2705 vdd.n632 185
R15095 vdd.n2771 vdd.n632 185
R15096 vdd.n2704 vdd.n2703 185
R15097 vdd.n2703 vdd.n631 185
R15098 vdd.n2702 vdd.n664 185
R15099 vdd.n2702 vdd.n2701 185
R15100 vdd.n2456 vdd.n665 185
R15101 vdd.n674 vdd.n665 185
R15102 vdd.n2457 vdd.n672 185
R15103 vdd.n2695 vdd.n672 185
R15104 vdd.n2459 vdd.n2458 185
R15105 vdd.n2458 vdd.n671 185
R15106 vdd.n2460 vdd.n680 185
R15107 vdd.n2644 vdd.n680 185
R15108 vdd.n2462 vdd.n2461 185
R15109 vdd.n2461 vdd.n679 185
R15110 vdd.n2463 vdd.n686 185
R15111 vdd.n2638 vdd.n686 185
R15112 vdd.n2465 vdd.n2464 185
R15113 vdd.n2464 vdd.n685 185
R15114 vdd.n2466 vdd.n691 185
R15115 vdd.n2630 vdd.n691 185
R15116 vdd.n2468 vdd.n2467 185
R15117 vdd.n2467 vdd.n698 185
R15118 vdd.n2469 vdd.n696 185
R15119 vdd.n2624 vdd.n696 185
R15120 vdd.n2471 vdd.n2470 185
R15121 vdd.n2472 vdd.n2471 185
R15122 vdd.n2455 vdd.n703 185
R15123 vdd.n2618 vdd.n703 185
R15124 vdd.n2454 vdd.n2453 185
R15125 vdd.n2453 vdd.n702 185
R15126 vdd.n2452 vdd.n709 185
R15127 vdd.n2612 vdd.n709 185
R15128 vdd.n2451 vdd.n2450 185
R15129 vdd.n2450 vdd.n708 185
R15130 vdd.n2449 vdd.n714 185
R15131 vdd.n2606 vdd.n714 185
R15132 vdd.n2448 vdd.n2447 185
R15133 vdd.n2447 vdd.n721 185
R15134 vdd.n2446 vdd.n719 185
R15135 vdd.n2600 vdd.n719 185
R15136 vdd.n2445 vdd.n2444 185
R15137 vdd.n2444 vdd.n728 185
R15138 vdd.n2443 vdd.n726 185
R15139 vdd.n2594 vdd.n726 185
R15140 vdd.n2442 vdd.n2441 185
R15141 vdd.n2441 vdd.n725 185
R15142 vdd.n2353 vdd.n732 185
R15143 vdd.n2588 vdd.n732 185
R15144 vdd.n2495 vdd.n2494 185
R15145 vdd.n2494 vdd.n2493 185
R15146 vdd.n2496 vdd.n737 185
R15147 vdd.n2582 vdd.n737 185
R15148 vdd.n2498 vdd.n2497 185
R15149 vdd.n2497 vdd.t209 185
R15150 vdd.n2499 vdd.n742 185
R15151 vdd.n2576 vdd.n742 185
R15152 vdd.n2578 vdd.n2577 185
R15153 vdd.n2577 vdd.n2576 185
R15154 vdd.n2579 vdd.n739 185
R15155 vdd.n739 vdd.t209 185
R15156 vdd.n2581 vdd.n2580 185
R15157 vdd.n2582 vdd.n2581 185
R15158 vdd.n731 vdd.n730 185
R15159 vdd.n2493 vdd.n731 185
R15160 vdd.n2590 vdd.n2589 185
R15161 vdd.n2589 vdd.n2588 185
R15162 vdd.n2591 vdd.n729 185
R15163 vdd.n729 vdd.n725 185
R15164 vdd.n2593 vdd.n2592 185
R15165 vdd.n2594 vdd.n2593 185
R15166 vdd.n718 vdd.n717 185
R15167 vdd.n728 vdd.n718 185
R15168 vdd.n2602 vdd.n2601 185
R15169 vdd.n2601 vdd.n2600 185
R15170 vdd.n2603 vdd.n716 185
R15171 vdd.n721 vdd.n716 185
R15172 vdd.n2605 vdd.n2604 185
R15173 vdd.n2606 vdd.n2605 185
R15174 vdd.n707 vdd.n706 185
R15175 vdd.n708 vdd.n707 185
R15176 vdd.n2614 vdd.n2613 185
R15177 vdd.n2613 vdd.n2612 185
R15178 vdd.n2615 vdd.n705 185
R15179 vdd.n705 vdd.n702 185
R15180 vdd.n2617 vdd.n2616 185
R15181 vdd.n2618 vdd.n2617 185
R15182 vdd.n695 vdd.n694 185
R15183 vdd.n2472 vdd.n695 185
R15184 vdd.n2626 vdd.n2625 185
R15185 vdd.n2625 vdd.n2624 185
R15186 vdd.n2627 vdd.n693 185
R15187 vdd.n698 vdd.n693 185
R15188 vdd.n2629 vdd.n2628 185
R15189 vdd.n2630 vdd.n2629 185
R15190 vdd.n684 vdd.n683 185
R15191 vdd.n685 vdd.n684 185
R15192 vdd.n2640 vdd.n2639 185
R15193 vdd.n2639 vdd.n2638 185
R15194 vdd.n2641 vdd.n682 185
R15195 vdd.n682 vdd.n679 185
R15196 vdd.n2643 vdd.n2642 185
R15197 vdd.n2644 vdd.n2643 185
R15198 vdd.n670 vdd.n669 185
R15199 vdd.n671 vdd.n670 185
R15200 vdd.n2697 vdd.n2696 185
R15201 vdd.n2696 vdd.n2695 185
R15202 vdd.n2698 vdd.n668 185
R15203 vdd.n674 vdd.n668 185
R15204 vdd.n2700 vdd.n2699 185
R15205 vdd.n2701 vdd.n2700 185
R15206 vdd.n636 vdd.n634 185
R15207 vdd.n634 vdd.n631 185
R15208 vdd.n2770 vdd.n2769 185
R15209 vdd.n2771 vdd.n2770 185
R15210 vdd.n2243 vdd.n2242 185
R15211 vdd.n2244 vdd.n2243 185
R15212 vdd.n792 vdd.n790 185
R15213 vdd.n790 vdd.t182 185
R15214 vdd.n2158 vdd.n799 185
R15215 vdd.n2169 vdd.n799 185
R15216 vdd.n2159 vdd.n808 185
R15217 vdd.n1868 vdd.n808 185
R15218 vdd.n2161 vdd.n2160 185
R15219 vdd.n2162 vdd.n2161 185
R15220 vdd.n2157 vdd.n807 185
R15221 vdd.n807 vdd.n804 185
R15222 vdd.n2156 vdd.n2155 185
R15223 vdd.n2155 vdd.n2154 185
R15224 vdd.n810 vdd.n809 185
R15225 vdd.n811 vdd.n810 185
R15226 vdd.n2147 vdd.n2146 185
R15227 vdd.n2148 vdd.n2147 185
R15228 vdd.n2145 vdd.n820 185
R15229 vdd.n820 vdd.n817 185
R15230 vdd.n2144 vdd.n2143 185
R15231 vdd.n2143 vdd.n2142 185
R15232 vdd.n822 vdd.n821 185
R15233 vdd.n830 vdd.n822 185
R15234 vdd.n2135 vdd.n2134 185
R15235 vdd.n2136 vdd.n2135 185
R15236 vdd.n2133 vdd.n831 185
R15237 vdd.n836 vdd.n831 185
R15238 vdd.n2132 vdd.n2131 185
R15239 vdd.n2131 vdd.n2130 185
R15240 vdd.n833 vdd.n832 185
R15241 vdd.n1969 vdd.n833 185
R15242 vdd.n2123 vdd.n2122 185
R15243 vdd.n2124 vdd.n2123 185
R15244 vdd.n2121 vdd.n843 185
R15245 vdd.n843 vdd.n840 185
R15246 vdd.n2120 vdd.n2119 185
R15247 vdd.n2119 vdd.n2118 185
R15248 vdd.n845 vdd.n844 185
R15249 vdd.n846 vdd.n845 185
R15250 vdd.n2111 vdd.n2110 185
R15251 vdd.n2112 vdd.n2111 185
R15252 vdd.n2108 vdd.n854 185
R15253 vdd.n861 vdd.n854 185
R15254 vdd.n2107 vdd.n2106 185
R15255 vdd.n2106 vdd.n2105 185
R15256 vdd.n857 vdd.n856 185
R15257 vdd.n858 vdd.n857 185
R15258 vdd.n2098 vdd.n2097 185
R15259 vdd.n2099 vdd.n2098 185
R15260 vdd.n2096 vdd.n868 185
R15261 vdd.n868 vdd.n865 185
R15262 vdd.n2095 vdd.n2094 185
R15263 vdd.n2094 vdd.n2093 185
R15264 vdd.n870 vdd.n869 185
R15265 vdd.n871 vdd.n870 185
R15266 vdd.n2086 vdd.n2085 185
R15267 vdd.n2087 vdd.n2086 185
R15268 vdd.n2174 vdd.n764 185
R15269 vdd.n2316 vdd.n764 185
R15270 vdd.n2176 vdd.n2175 185
R15271 vdd.n2178 vdd.n2177 185
R15272 vdd.n2180 vdd.n2179 185
R15273 vdd.n2182 vdd.n2181 185
R15274 vdd.n2184 vdd.n2183 185
R15275 vdd.n2186 vdd.n2185 185
R15276 vdd.n2188 vdd.n2187 185
R15277 vdd.n2190 vdd.n2189 185
R15278 vdd.n2192 vdd.n2191 185
R15279 vdd.n2194 vdd.n2193 185
R15280 vdd.n2196 vdd.n2195 185
R15281 vdd.n2198 vdd.n2197 185
R15282 vdd.n2200 vdd.n2199 185
R15283 vdd.n2202 vdd.n2201 185
R15284 vdd.n2204 vdd.n2203 185
R15285 vdd.n2206 vdd.n2205 185
R15286 vdd.n2208 vdd.n2207 185
R15287 vdd.n2210 vdd.n2209 185
R15288 vdd.n2212 vdd.n2211 185
R15289 vdd.n2214 vdd.n2213 185
R15290 vdd.n2216 vdd.n2215 185
R15291 vdd.n2218 vdd.n2217 185
R15292 vdd.n2220 vdd.n2219 185
R15293 vdd.n2222 vdd.n2221 185
R15294 vdd.n2224 vdd.n2223 185
R15295 vdd.n2226 vdd.n2225 185
R15296 vdd.n2228 vdd.n2227 185
R15297 vdd.n2230 vdd.n2229 185
R15298 vdd.n2232 vdd.n2231 185
R15299 vdd.n2234 vdd.n2233 185
R15300 vdd.n2236 vdd.n2235 185
R15301 vdd.n2238 vdd.n2237 185
R15302 vdd.n2240 vdd.n2239 185
R15303 vdd.n2241 vdd.n791 185
R15304 vdd.n2173 vdd.n789 185
R15305 vdd.n2244 vdd.n789 185
R15306 vdd.n2172 vdd.n2171 185
R15307 vdd.n2171 vdd.t182 185
R15308 vdd.n2170 vdd.n796 185
R15309 vdd.n2170 vdd.n2169 185
R15310 vdd.n1950 vdd.n797 185
R15311 vdd.n1868 vdd.n797 185
R15312 vdd.n1951 vdd.n806 185
R15313 vdd.n2162 vdd.n806 185
R15314 vdd.n1953 vdd.n1952 185
R15315 vdd.n1952 vdd.n804 185
R15316 vdd.n1954 vdd.n813 185
R15317 vdd.n2154 vdd.n813 185
R15318 vdd.n1956 vdd.n1955 185
R15319 vdd.n1955 vdd.n811 185
R15320 vdd.n1957 vdd.n819 185
R15321 vdd.n2148 vdd.n819 185
R15322 vdd.n1959 vdd.n1958 185
R15323 vdd.n1958 vdd.n817 185
R15324 vdd.n1960 vdd.n824 185
R15325 vdd.n2142 vdd.n824 185
R15326 vdd.n1962 vdd.n1961 185
R15327 vdd.n1961 vdd.n830 185
R15328 vdd.n1963 vdd.n829 185
R15329 vdd.n2136 vdd.n829 185
R15330 vdd.n1965 vdd.n1964 185
R15331 vdd.n1964 vdd.n836 185
R15332 vdd.n1966 vdd.n835 185
R15333 vdd.n2130 vdd.n835 185
R15334 vdd.n1968 vdd.n1967 185
R15335 vdd.n1969 vdd.n1968 185
R15336 vdd.n1949 vdd.n842 185
R15337 vdd.n2124 vdd.n842 185
R15338 vdd.n1948 vdd.n1947 185
R15339 vdd.n1947 vdd.n840 185
R15340 vdd.n1946 vdd.n848 185
R15341 vdd.n2118 vdd.n848 185
R15342 vdd.n1945 vdd.n1944 185
R15343 vdd.n1944 vdd.n846 185
R15344 vdd.n1943 vdd.n853 185
R15345 vdd.n2112 vdd.n853 185
R15346 vdd.n1942 vdd.n1941 185
R15347 vdd.n1941 vdd.n861 185
R15348 vdd.n1940 vdd.n860 185
R15349 vdd.n2105 vdd.n860 185
R15350 vdd.n1939 vdd.n1938 185
R15351 vdd.n1938 vdd.n858 185
R15352 vdd.n1937 vdd.n867 185
R15353 vdd.n2099 vdd.n867 185
R15354 vdd.n1936 vdd.n1935 185
R15355 vdd.n1935 vdd.n865 185
R15356 vdd.n1934 vdd.n873 185
R15357 vdd.n2093 vdd.n873 185
R15358 vdd.n1933 vdd.n1932 185
R15359 vdd.n1932 vdd.n871 185
R15360 vdd.n1931 vdd.n879 185
R15361 vdd.n2087 vdd.n879 185
R15362 vdd.n2084 vdd.n880 185
R15363 vdd.n2083 vdd.n2082 185
R15364 vdd.n2080 vdd.n881 185
R15365 vdd.n2078 vdd.n2077 185
R15366 vdd.n2076 vdd.n882 185
R15367 vdd.n2075 vdd.n2074 185
R15368 vdd.n2072 vdd.n883 185
R15369 vdd.n2070 vdd.n2069 185
R15370 vdd.n2068 vdd.n884 185
R15371 vdd.n2067 vdd.n2066 185
R15372 vdd.n2064 vdd.n885 185
R15373 vdd.n2062 vdd.n2061 185
R15374 vdd.n2060 vdd.n886 185
R15375 vdd.n2059 vdd.n2058 185
R15376 vdd.n2056 vdd.n887 185
R15377 vdd.n2054 vdd.n2053 185
R15378 vdd.n2052 vdd.n888 185
R15379 vdd.n2051 vdd.n890 185
R15380 vdd.n1896 vdd.n891 185
R15381 vdd.n1899 vdd.n1898 185
R15382 vdd.n1901 vdd.n1900 185
R15383 vdd.n1903 vdd.n1895 185
R15384 vdd.n1906 vdd.n1905 185
R15385 vdd.n1907 vdd.n1894 185
R15386 vdd.n1909 vdd.n1908 185
R15387 vdd.n1911 vdd.n1893 185
R15388 vdd.n1914 vdd.n1913 185
R15389 vdd.n1915 vdd.n1892 185
R15390 vdd.n1917 vdd.n1916 185
R15391 vdd.n1919 vdd.n1891 185
R15392 vdd.n1922 vdd.n1921 185
R15393 vdd.n1923 vdd.n1888 185
R15394 vdd.n1926 vdd.n1925 185
R15395 vdd.n1928 vdd.n1887 185
R15396 vdd.n1930 vdd.n1929 185
R15397 vdd.n1929 vdd.n877 185
R15398 vdd.n303 vdd.n302 171.744
R15399 vdd.n302 vdd.n301 171.744
R15400 vdd.n301 vdd.n270 171.744
R15401 vdd.n294 vdd.n270 171.744
R15402 vdd.n294 vdd.n293 171.744
R15403 vdd.n293 vdd.n275 171.744
R15404 vdd.n286 vdd.n275 171.744
R15405 vdd.n286 vdd.n285 171.744
R15406 vdd.n285 vdd.n279 171.744
R15407 vdd.n252 vdd.n251 171.744
R15408 vdd.n251 vdd.n250 171.744
R15409 vdd.n250 vdd.n219 171.744
R15410 vdd.n243 vdd.n219 171.744
R15411 vdd.n243 vdd.n242 171.744
R15412 vdd.n242 vdd.n224 171.744
R15413 vdd.n235 vdd.n224 171.744
R15414 vdd.n235 vdd.n234 171.744
R15415 vdd.n234 vdd.n228 171.744
R15416 vdd.n209 vdd.n208 171.744
R15417 vdd.n208 vdd.n207 171.744
R15418 vdd.n207 vdd.n176 171.744
R15419 vdd.n200 vdd.n176 171.744
R15420 vdd.n200 vdd.n199 171.744
R15421 vdd.n199 vdd.n181 171.744
R15422 vdd.n192 vdd.n181 171.744
R15423 vdd.n192 vdd.n191 171.744
R15424 vdd.n191 vdd.n185 171.744
R15425 vdd.n158 vdd.n157 171.744
R15426 vdd.n157 vdd.n156 171.744
R15427 vdd.n156 vdd.n125 171.744
R15428 vdd.n149 vdd.n125 171.744
R15429 vdd.n149 vdd.n148 171.744
R15430 vdd.n148 vdd.n130 171.744
R15431 vdd.n141 vdd.n130 171.744
R15432 vdd.n141 vdd.n140 171.744
R15433 vdd.n140 vdd.n134 171.744
R15434 vdd.n116 vdd.n115 171.744
R15435 vdd.n115 vdd.n114 171.744
R15436 vdd.n114 vdd.n83 171.744
R15437 vdd.n107 vdd.n83 171.744
R15438 vdd.n107 vdd.n106 171.744
R15439 vdd.n106 vdd.n88 171.744
R15440 vdd.n99 vdd.n88 171.744
R15441 vdd.n99 vdd.n98 171.744
R15442 vdd.n98 vdd.n92 171.744
R15443 vdd.n65 vdd.n64 171.744
R15444 vdd.n64 vdd.n63 171.744
R15445 vdd.n63 vdd.n32 171.744
R15446 vdd.n56 vdd.n32 171.744
R15447 vdd.n56 vdd.n55 171.744
R15448 vdd.n55 vdd.n37 171.744
R15449 vdd.n48 vdd.n37 171.744
R15450 vdd.n48 vdd.n47 171.744
R15451 vdd.n47 vdd.n41 171.744
R15452 vdd.n1498 vdd.n1497 171.744
R15453 vdd.n1497 vdd.n1496 171.744
R15454 vdd.n1496 vdd.n1465 171.744
R15455 vdd.n1489 vdd.n1465 171.744
R15456 vdd.n1489 vdd.n1488 171.744
R15457 vdd.n1488 vdd.n1470 171.744
R15458 vdd.n1481 vdd.n1470 171.744
R15459 vdd.n1481 vdd.n1480 171.744
R15460 vdd.n1480 vdd.n1474 171.744
R15461 vdd.n1549 vdd.n1548 171.744
R15462 vdd.n1548 vdd.n1547 171.744
R15463 vdd.n1547 vdd.n1516 171.744
R15464 vdd.n1540 vdd.n1516 171.744
R15465 vdd.n1540 vdd.n1539 171.744
R15466 vdd.n1539 vdd.n1521 171.744
R15467 vdd.n1532 vdd.n1521 171.744
R15468 vdd.n1532 vdd.n1531 171.744
R15469 vdd.n1531 vdd.n1525 171.744
R15470 vdd.n1404 vdd.n1403 171.744
R15471 vdd.n1403 vdd.n1402 171.744
R15472 vdd.n1402 vdd.n1371 171.744
R15473 vdd.n1395 vdd.n1371 171.744
R15474 vdd.n1395 vdd.n1394 171.744
R15475 vdd.n1394 vdd.n1376 171.744
R15476 vdd.n1387 vdd.n1376 171.744
R15477 vdd.n1387 vdd.n1386 171.744
R15478 vdd.n1386 vdd.n1380 171.744
R15479 vdd.n1455 vdd.n1454 171.744
R15480 vdd.n1454 vdd.n1453 171.744
R15481 vdd.n1453 vdd.n1422 171.744
R15482 vdd.n1446 vdd.n1422 171.744
R15483 vdd.n1446 vdd.n1445 171.744
R15484 vdd.n1445 vdd.n1427 171.744
R15485 vdd.n1438 vdd.n1427 171.744
R15486 vdd.n1438 vdd.n1437 171.744
R15487 vdd.n1437 vdd.n1431 171.744
R15488 vdd.n1311 vdd.n1310 171.744
R15489 vdd.n1310 vdd.n1309 171.744
R15490 vdd.n1309 vdd.n1278 171.744
R15491 vdd.n1302 vdd.n1278 171.744
R15492 vdd.n1302 vdd.n1301 171.744
R15493 vdd.n1301 vdd.n1283 171.744
R15494 vdd.n1294 vdd.n1283 171.744
R15495 vdd.n1294 vdd.n1293 171.744
R15496 vdd.n1293 vdd.n1287 171.744
R15497 vdd.n1362 vdd.n1361 171.744
R15498 vdd.n1361 vdd.n1360 171.744
R15499 vdd.n1360 vdd.n1329 171.744
R15500 vdd.n1353 vdd.n1329 171.744
R15501 vdd.n1353 vdd.n1352 171.744
R15502 vdd.n1352 vdd.n1334 171.744
R15503 vdd.n1345 vdd.n1334 171.744
R15504 vdd.n1345 vdd.n1344 171.744
R15505 vdd.n1344 vdd.n1338 171.744
R15506 vdd.n3130 vdd.n356 146.341
R15507 vdd.n3128 vdd.n3127 146.341
R15508 vdd.n3125 vdd.n360 146.341
R15509 vdd.n3121 vdd.n3120 146.341
R15510 vdd.n3118 vdd.n368 146.341
R15511 vdd.n3114 vdd.n3113 146.341
R15512 vdd.n3111 vdd.n375 146.341
R15513 vdd.n3107 vdd.n3106 146.341
R15514 vdd.n3104 vdd.n382 146.341
R15515 vdd.n393 vdd.n390 146.341
R15516 vdd.n3096 vdd.n3095 146.341
R15517 vdd.n3093 vdd.n395 146.341
R15518 vdd.n3089 vdd.n3088 146.341
R15519 vdd.n3086 vdd.n401 146.341
R15520 vdd.n3082 vdd.n3081 146.341
R15521 vdd.n3079 vdd.n408 146.341
R15522 vdd.n3075 vdd.n3074 146.341
R15523 vdd.n3072 vdd.n415 146.341
R15524 vdd.n3068 vdd.n3067 146.341
R15525 vdd.n3065 vdd.n422 146.341
R15526 vdd.n433 vdd.n430 146.341
R15527 vdd.n3057 vdd.n3056 146.341
R15528 vdd.n3054 vdd.n435 146.341
R15529 vdd.n3050 vdd.n3049 146.341
R15530 vdd.n3047 vdd.n441 146.341
R15531 vdd.n3043 vdd.n3042 146.341
R15532 vdd.n3040 vdd.n448 146.341
R15533 vdd.n3036 vdd.n3035 146.341
R15534 vdd.n3033 vdd.n455 146.341
R15535 vdd.n3029 vdd.n3028 146.341
R15536 vdd.n3026 vdd.n462 146.341
R15537 vdd.n2941 vdd.n512 146.341
R15538 vdd.n2947 vdd.n512 146.341
R15539 vdd.n2947 vdd.n504 146.341
R15540 vdd.n2957 vdd.n504 146.341
R15541 vdd.n2957 vdd.n500 146.341
R15542 vdd.n2963 vdd.n500 146.341
R15543 vdd.n2963 vdd.n491 146.341
R15544 vdd.n2973 vdd.n491 146.341
R15545 vdd.n2973 vdd.n487 146.341
R15546 vdd.n2979 vdd.n487 146.341
R15547 vdd.n2979 vdd.n479 146.341
R15548 vdd.n2990 vdd.n479 146.341
R15549 vdd.n2990 vdd.n480 146.341
R15550 vdd.n480 vdd.n316 146.341
R15551 vdd.n317 vdd.n316 146.341
R15552 vdd.n318 vdd.n317 146.341
R15553 vdd.n473 vdd.n318 146.341
R15554 vdd.n473 vdd.n326 146.341
R15555 vdd.n327 vdd.n326 146.341
R15556 vdd.n328 vdd.n327 146.341
R15557 vdd.n470 vdd.n328 146.341
R15558 vdd.n470 vdd.n337 146.341
R15559 vdd.n338 vdd.n337 146.341
R15560 vdd.n339 vdd.n338 146.341
R15561 vdd.n467 vdd.n339 146.341
R15562 vdd.n467 vdd.n348 146.341
R15563 vdd.n349 vdd.n348 146.341
R15564 vdd.n350 vdd.n349 146.341
R15565 vdd.n2933 vdd.n2931 146.341
R15566 vdd.n2931 vdd.n2930 146.341
R15567 vdd.n2927 vdd.n2926 146.341
R15568 vdd.n2923 vdd.n2922 146.341
R15569 vdd.n2920 vdd.n526 146.341
R15570 vdd.n2916 vdd.n2914 146.341
R15571 vdd.n2912 vdd.n532 146.341
R15572 vdd.n2908 vdd.n2906 146.341
R15573 vdd.n2904 vdd.n538 146.341
R15574 vdd.n2900 vdd.n2898 146.341
R15575 vdd.n2896 vdd.n546 146.341
R15576 vdd.n2892 vdd.n2890 146.341
R15577 vdd.n2888 vdd.n552 146.341
R15578 vdd.n2884 vdd.n2882 146.341
R15579 vdd.n2880 vdd.n558 146.341
R15580 vdd.n2876 vdd.n2874 146.341
R15581 vdd.n2872 vdd.n564 146.341
R15582 vdd.n2868 vdd.n2866 146.341
R15583 vdd.n2864 vdd.n570 146.341
R15584 vdd.n2860 vdd.n2858 146.341
R15585 vdd.n2856 vdd.n576 146.341
R15586 vdd.n2849 vdd.n585 146.341
R15587 vdd.n2847 vdd.n2846 146.341
R15588 vdd.n2843 vdd.n2842 146.341
R15589 vdd.n2840 vdd.n590 146.341
R15590 vdd.n2836 vdd.n2834 146.341
R15591 vdd.n2832 vdd.n596 146.341
R15592 vdd.n2828 vdd.n2826 146.341
R15593 vdd.n2824 vdd.n602 146.341
R15594 vdd.n2820 vdd.n2818 146.341
R15595 vdd.n2815 vdd.n2814 146.341
R15596 vdd.n2811 vdd.n515 146.341
R15597 vdd.n2939 vdd.n510 146.341
R15598 vdd.n2949 vdd.n510 146.341
R15599 vdd.n2949 vdd.n506 146.341
R15600 vdd.n2955 vdd.n506 146.341
R15601 vdd.n2955 vdd.n498 146.341
R15602 vdd.n2965 vdd.n498 146.341
R15603 vdd.n2965 vdd.n494 146.341
R15604 vdd.n2971 vdd.n494 146.341
R15605 vdd.n2971 vdd.n486 146.341
R15606 vdd.n2982 vdd.n486 146.341
R15607 vdd.n2982 vdd.n482 146.341
R15608 vdd.n2988 vdd.n482 146.341
R15609 vdd.n2988 vdd.n314 146.341
R15610 vdd.n3165 vdd.n314 146.341
R15611 vdd.n3165 vdd.n315 146.341
R15612 vdd.n3161 vdd.n315 146.341
R15613 vdd.n3161 vdd.n319 146.341
R15614 vdd.n3157 vdd.n319 146.341
R15615 vdd.n3157 vdd.n324 146.341
R15616 vdd.n3153 vdd.n324 146.341
R15617 vdd.n3153 vdd.n330 146.341
R15618 vdd.n3149 vdd.n330 146.341
R15619 vdd.n3149 vdd.n336 146.341
R15620 vdd.n3145 vdd.n336 146.341
R15621 vdd.n3145 vdd.n341 146.341
R15622 vdd.n3141 vdd.n341 146.341
R15623 vdd.n3141 vdd.n347 146.341
R15624 vdd.n3137 vdd.n347 146.341
R15625 vdd.n2034 vdd.n2033 146.341
R15626 vdd.n2031 vdd.n1615 146.341
R15627 vdd.n1811 vdd.n1621 146.341
R15628 vdd.n1809 vdd.n1808 146.341
R15629 vdd.n1806 vdd.n1623 146.341
R15630 vdd.n1802 vdd.n1801 146.341
R15631 vdd.n1799 vdd.n1630 146.341
R15632 vdd.n1795 vdd.n1794 146.341
R15633 vdd.n1792 vdd.n1637 146.341
R15634 vdd.n1648 vdd.n1645 146.341
R15635 vdd.n1784 vdd.n1783 146.341
R15636 vdd.n1781 vdd.n1650 146.341
R15637 vdd.n1777 vdd.n1776 146.341
R15638 vdd.n1774 vdd.n1656 146.341
R15639 vdd.n1770 vdd.n1769 146.341
R15640 vdd.n1767 vdd.n1663 146.341
R15641 vdd.n1763 vdd.n1762 146.341
R15642 vdd.n1760 vdd.n1670 146.341
R15643 vdd.n1756 vdd.n1755 146.341
R15644 vdd.n1753 vdd.n1677 146.341
R15645 vdd.n1688 vdd.n1685 146.341
R15646 vdd.n1745 vdd.n1744 146.341
R15647 vdd.n1742 vdd.n1690 146.341
R15648 vdd.n1738 vdd.n1737 146.341
R15649 vdd.n1735 vdd.n1696 146.341
R15650 vdd.n1731 vdd.n1730 146.341
R15651 vdd.n1728 vdd.n1703 146.341
R15652 vdd.n1724 vdd.n1723 146.341
R15653 vdd.n1721 vdd.n1718 146.341
R15654 vdd.n1716 vdd.n1713 146.341
R15655 vdd.n1711 vdd.n897 146.341
R15656 vdd.n1216 vdd.n978 146.341
R15657 vdd.n1222 vdd.n978 146.341
R15658 vdd.n1222 vdd.n971 146.341
R15659 vdd.n1232 vdd.n971 146.341
R15660 vdd.n1232 vdd.n967 146.341
R15661 vdd.n1238 vdd.n967 146.341
R15662 vdd.n1238 vdd.n958 146.341
R15663 vdd.n1248 vdd.n958 146.341
R15664 vdd.n1248 vdd.n954 146.341
R15665 vdd.n1254 vdd.n954 146.341
R15666 vdd.n1254 vdd.n947 146.341
R15667 vdd.n1265 vdd.n947 146.341
R15668 vdd.n1265 vdd.n943 146.341
R15669 vdd.n1271 vdd.n943 146.341
R15670 vdd.n1271 vdd.n936 146.341
R15671 vdd.n1563 vdd.n936 146.341
R15672 vdd.n1563 vdd.n932 146.341
R15673 vdd.n1569 vdd.n932 146.341
R15674 vdd.n1569 vdd.n924 146.341
R15675 vdd.n1580 vdd.n924 146.341
R15676 vdd.n1580 vdd.n920 146.341
R15677 vdd.n1586 vdd.n920 146.341
R15678 vdd.n1586 vdd.n914 146.341
R15679 vdd.n1597 vdd.n914 146.341
R15680 vdd.n1597 vdd.n909 146.341
R15681 vdd.n1605 vdd.n909 146.341
R15682 vdd.n1605 vdd.n899 146.341
R15683 vdd.n2042 vdd.n899 146.341
R15684 vdd.n988 vdd.n987 146.341
R15685 vdd.n991 vdd.n988 146.341
R15686 vdd.n994 vdd.n993 146.341
R15687 vdd.n999 vdd.n996 146.341
R15688 vdd.n1002 vdd.n1001 146.341
R15689 vdd.n1007 vdd.n1004 146.341
R15690 vdd.n1010 vdd.n1009 146.341
R15691 vdd.n1015 vdd.n1012 146.341
R15692 vdd.n1018 vdd.n1017 146.341
R15693 vdd.n1025 vdd.n1020 146.341
R15694 vdd.n1028 vdd.n1027 146.341
R15695 vdd.n1033 vdd.n1030 146.341
R15696 vdd.n1036 vdd.n1035 146.341
R15697 vdd.n1041 vdd.n1038 146.341
R15698 vdd.n1044 vdd.n1043 146.341
R15699 vdd.n1049 vdd.n1046 146.341
R15700 vdd.n1052 vdd.n1051 146.341
R15701 vdd.n1057 vdd.n1054 146.341
R15702 vdd.n1060 vdd.n1059 146.341
R15703 vdd.n1065 vdd.n1062 146.341
R15704 vdd.n1146 vdd.n1067 146.341
R15705 vdd.n1144 vdd.n1143 146.341
R15706 vdd.n1074 vdd.n1073 146.341
R15707 vdd.n1077 vdd.n1076 146.341
R15708 vdd.n1082 vdd.n1081 146.341
R15709 vdd.n1085 vdd.n1084 146.341
R15710 vdd.n1090 vdd.n1089 146.341
R15711 vdd.n1093 vdd.n1092 146.341
R15712 vdd.n1098 vdd.n1097 146.341
R15713 vdd.n1101 vdd.n1100 146.341
R15714 vdd.n1106 vdd.n1105 146.341
R15715 vdd.n1108 vdd.n981 146.341
R15716 vdd.n1214 vdd.n977 146.341
R15717 vdd.n1224 vdd.n977 146.341
R15718 vdd.n1224 vdd.n973 146.341
R15719 vdd.n1230 vdd.n973 146.341
R15720 vdd.n1230 vdd.n965 146.341
R15721 vdd.n1240 vdd.n965 146.341
R15722 vdd.n1240 vdd.n961 146.341
R15723 vdd.n1246 vdd.n961 146.341
R15724 vdd.n1246 vdd.n953 146.341
R15725 vdd.n1257 vdd.n953 146.341
R15726 vdd.n1257 vdd.n949 146.341
R15727 vdd.n1263 vdd.n949 146.341
R15728 vdd.n1263 vdd.n942 146.341
R15729 vdd.n1273 vdd.n942 146.341
R15730 vdd.n1273 vdd.n938 146.341
R15731 vdd.n1561 vdd.n938 146.341
R15732 vdd.n1561 vdd.n930 146.341
R15733 vdd.n1572 vdd.n930 146.341
R15734 vdd.n1572 vdd.n926 146.341
R15735 vdd.n1578 vdd.n926 146.341
R15736 vdd.n1578 vdd.n919 146.341
R15737 vdd.n1589 vdd.n919 146.341
R15738 vdd.n1589 vdd.n915 146.341
R15739 vdd.n1595 vdd.n915 146.341
R15740 vdd.n1595 vdd.n907 146.341
R15741 vdd.n1608 vdd.n907 146.341
R15742 vdd.n1608 vdd.n902 146.341
R15743 vdd.n2040 vdd.n902 146.341
R15744 vdd.n901 vdd.n877 141.707
R15745 vdd.n613 vdd.n516 141.707
R15746 vdd.n1889 vdd.t132 127.284
R15747 vdd.n793 vdd.t116 127.284
R15748 vdd.n1863 vdd.t158 127.284
R15749 vdd.n785 vdd.t141 127.284
R15750 vdd.n2634 vdd.t103 127.284
R15751 vdd.n2634 vdd.t104 127.284
R15752 vdd.n2354 vdd.t139 127.284
R15753 vdd.n661 vdd.t120 127.284
R15754 vdd.n2351 vdd.t125 127.284
R15755 vdd.n625 vdd.t127 127.284
R15756 vdd.n855 vdd.t135 127.284
R15757 vdd.n855 vdd.t136 127.284
R15758 vdd.n22 vdd.n20 117.314
R15759 vdd.n17 vdd.n15 117.314
R15760 vdd.n27 vdd.n26 116.927
R15761 vdd.n24 vdd.n23 116.927
R15762 vdd.n22 vdd.n21 116.927
R15763 vdd.n17 vdd.n16 116.927
R15764 vdd.n19 vdd.n18 116.927
R15765 vdd.n27 vdd.n25 116.927
R15766 vdd.n1890 vdd.t131 111.188
R15767 vdd.n794 vdd.t117 111.188
R15768 vdd.n1864 vdd.t157 111.188
R15769 vdd.n786 vdd.t142 111.188
R15770 vdd.n2355 vdd.t138 111.188
R15771 vdd.n662 vdd.t121 111.188
R15772 vdd.n2352 vdd.t124 111.188
R15773 vdd.n626 vdd.t128 111.188
R15774 vdd.n2577 vdd.n739 99.5127
R15775 vdd.n2581 vdd.n739 99.5127
R15776 vdd.n2581 vdd.n731 99.5127
R15777 vdd.n2589 vdd.n731 99.5127
R15778 vdd.n2589 vdd.n729 99.5127
R15779 vdd.n2593 vdd.n729 99.5127
R15780 vdd.n2593 vdd.n718 99.5127
R15781 vdd.n2601 vdd.n718 99.5127
R15782 vdd.n2601 vdd.n716 99.5127
R15783 vdd.n2605 vdd.n716 99.5127
R15784 vdd.n2605 vdd.n707 99.5127
R15785 vdd.n2613 vdd.n707 99.5127
R15786 vdd.n2613 vdd.n705 99.5127
R15787 vdd.n2617 vdd.n705 99.5127
R15788 vdd.n2617 vdd.n695 99.5127
R15789 vdd.n2625 vdd.n695 99.5127
R15790 vdd.n2625 vdd.n693 99.5127
R15791 vdd.n2629 vdd.n693 99.5127
R15792 vdd.n2629 vdd.n684 99.5127
R15793 vdd.n2639 vdd.n684 99.5127
R15794 vdd.n2639 vdd.n682 99.5127
R15795 vdd.n2643 vdd.n682 99.5127
R15796 vdd.n2643 vdd.n670 99.5127
R15797 vdd.n2696 vdd.n670 99.5127
R15798 vdd.n2696 vdd.n668 99.5127
R15799 vdd.n2700 vdd.n668 99.5127
R15800 vdd.n2700 vdd.n634 99.5127
R15801 vdd.n2770 vdd.n634 99.5127
R15802 vdd.n2766 vdd.n635 99.5127
R15803 vdd.n2764 vdd.n2763 99.5127
R15804 vdd.n2761 vdd.n639 99.5127
R15805 vdd.n2757 vdd.n2756 99.5127
R15806 vdd.n2754 vdd.n642 99.5127
R15807 vdd.n2750 vdd.n2749 99.5127
R15808 vdd.n2747 vdd.n645 99.5127
R15809 vdd.n2743 vdd.n2742 99.5127
R15810 vdd.n2740 vdd.n648 99.5127
R15811 vdd.n2735 vdd.n2734 99.5127
R15812 vdd.n2732 vdd.n651 99.5127
R15813 vdd.n2728 vdd.n2727 99.5127
R15814 vdd.n2725 vdd.n654 99.5127
R15815 vdd.n2721 vdd.n2720 99.5127
R15816 vdd.n2718 vdd.n657 99.5127
R15817 vdd.n2714 vdd.n2713 99.5127
R15818 vdd.n2711 vdd.n660 99.5127
R15819 vdd.n2497 vdd.n742 99.5127
R15820 vdd.n2497 vdd.n737 99.5127
R15821 vdd.n2494 vdd.n737 99.5127
R15822 vdd.n2494 vdd.n732 99.5127
R15823 vdd.n2441 vdd.n732 99.5127
R15824 vdd.n2441 vdd.n726 99.5127
R15825 vdd.n2444 vdd.n726 99.5127
R15826 vdd.n2444 vdd.n719 99.5127
R15827 vdd.n2447 vdd.n719 99.5127
R15828 vdd.n2447 vdd.n714 99.5127
R15829 vdd.n2450 vdd.n714 99.5127
R15830 vdd.n2450 vdd.n709 99.5127
R15831 vdd.n2453 vdd.n709 99.5127
R15832 vdd.n2453 vdd.n703 99.5127
R15833 vdd.n2471 vdd.n703 99.5127
R15834 vdd.n2471 vdd.n696 99.5127
R15835 vdd.n2467 vdd.n696 99.5127
R15836 vdd.n2467 vdd.n691 99.5127
R15837 vdd.n2464 vdd.n691 99.5127
R15838 vdd.n2464 vdd.n686 99.5127
R15839 vdd.n2461 vdd.n686 99.5127
R15840 vdd.n2461 vdd.n680 99.5127
R15841 vdd.n2458 vdd.n680 99.5127
R15842 vdd.n2458 vdd.n672 99.5127
R15843 vdd.n672 vdd.n665 99.5127
R15844 vdd.n2702 vdd.n665 99.5127
R15845 vdd.n2703 vdd.n2702 99.5127
R15846 vdd.n2703 vdd.n632 99.5127
R15847 vdd.n2567 vdd.n2350 99.5127
R15848 vdd.n2563 vdd.n2350 99.5127
R15849 vdd.n2561 vdd.n2560 99.5127
R15850 vdd.n2557 vdd.n2556 99.5127
R15851 vdd.n2553 vdd.n2552 99.5127
R15852 vdd.n2549 vdd.n2548 99.5127
R15853 vdd.n2545 vdd.n2544 99.5127
R15854 vdd.n2541 vdd.n2540 99.5127
R15855 vdd.n2537 vdd.n2536 99.5127
R15856 vdd.n2533 vdd.n2532 99.5127
R15857 vdd.n2529 vdd.n2528 99.5127
R15858 vdd.n2525 vdd.n2524 99.5127
R15859 vdd.n2521 vdd.n2520 99.5127
R15860 vdd.n2517 vdd.n2516 99.5127
R15861 vdd.n2513 vdd.n2512 99.5127
R15862 vdd.n2509 vdd.n2508 99.5127
R15863 vdd.n2504 vdd.n2503 99.5127
R15864 vdd.n2315 vdd.n783 99.5127
R15865 vdd.n2311 vdd.n2310 99.5127
R15866 vdd.n2307 vdd.n2306 99.5127
R15867 vdd.n2303 vdd.n2302 99.5127
R15868 vdd.n2299 vdd.n2298 99.5127
R15869 vdd.n2295 vdd.n2294 99.5127
R15870 vdd.n2291 vdd.n2290 99.5127
R15871 vdd.n2287 vdd.n2286 99.5127
R15872 vdd.n2283 vdd.n2282 99.5127
R15873 vdd.n2279 vdd.n2278 99.5127
R15874 vdd.n2275 vdd.n2274 99.5127
R15875 vdd.n2271 vdd.n2270 99.5127
R15876 vdd.n2267 vdd.n2266 99.5127
R15877 vdd.n2263 vdd.n2262 99.5127
R15878 vdd.n2259 vdd.n2258 99.5127
R15879 vdd.n2255 vdd.n2254 99.5127
R15880 vdd.n2250 vdd.n2249 99.5127
R15881 vdd.n1988 vdd.n878 99.5127
R15882 vdd.n1988 vdd.n872 99.5127
R15883 vdd.n1985 vdd.n872 99.5127
R15884 vdd.n1985 vdd.n866 99.5127
R15885 vdd.n1982 vdd.n866 99.5127
R15886 vdd.n1982 vdd.n859 99.5127
R15887 vdd.n1979 vdd.n859 99.5127
R15888 vdd.n1979 vdd.n852 99.5127
R15889 vdd.n1976 vdd.n852 99.5127
R15890 vdd.n1976 vdd.n847 99.5127
R15891 vdd.n1973 vdd.n847 99.5127
R15892 vdd.n1973 vdd.n841 99.5127
R15893 vdd.n1970 vdd.n841 99.5127
R15894 vdd.n1970 vdd.n834 99.5127
R15895 vdd.n1884 vdd.n834 99.5127
R15896 vdd.n1884 vdd.n828 99.5127
R15897 vdd.n1881 vdd.n828 99.5127
R15898 vdd.n1881 vdd.n823 99.5127
R15899 vdd.n1878 vdd.n823 99.5127
R15900 vdd.n1878 vdd.n818 99.5127
R15901 vdd.n1875 vdd.n818 99.5127
R15902 vdd.n1875 vdd.n812 99.5127
R15903 vdd.n1872 vdd.n812 99.5127
R15904 vdd.n1872 vdd.n805 99.5127
R15905 vdd.n1869 vdd.n805 99.5127
R15906 vdd.n1869 vdd.n798 99.5127
R15907 vdd.n798 vdd.n788 99.5127
R15908 vdd.n2245 vdd.n788 99.5127
R15909 vdd.n1823 vdd.n1821 99.5127
R15910 vdd.n1827 vdd.n1821 99.5127
R15911 vdd.n1831 vdd.n1829 99.5127
R15912 vdd.n1835 vdd.n1819 99.5127
R15913 vdd.n1839 vdd.n1837 99.5127
R15914 vdd.n1843 vdd.n1817 99.5127
R15915 vdd.n1847 vdd.n1845 99.5127
R15916 vdd.n1851 vdd.n1815 99.5127
R15917 vdd.n1854 vdd.n1853 99.5127
R15918 vdd.n2024 vdd.n2022 99.5127
R15919 vdd.n2020 vdd.n1856 99.5127
R15920 vdd.n2016 vdd.n2014 99.5127
R15921 vdd.n2012 vdd.n1858 99.5127
R15922 vdd.n2008 vdd.n2006 99.5127
R15923 vdd.n2004 vdd.n1860 99.5127
R15924 vdd.n2000 vdd.n1998 99.5127
R15925 vdd.n1996 vdd.n1862 99.5127
R15926 vdd.n2088 vdd.n874 99.5127
R15927 vdd.n2092 vdd.n874 99.5127
R15928 vdd.n2092 vdd.n864 99.5127
R15929 vdd.n2100 vdd.n864 99.5127
R15930 vdd.n2100 vdd.n862 99.5127
R15931 vdd.n2104 vdd.n862 99.5127
R15932 vdd.n2104 vdd.n851 99.5127
R15933 vdd.n2113 vdd.n851 99.5127
R15934 vdd.n2113 vdd.n849 99.5127
R15935 vdd.n2117 vdd.n849 99.5127
R15936 vdd.n2117 vdd.n839 99.5127
R15937 vdd.n2125 vdd.n839 99.5127
R15938 vdd.n2125 vdd.n837 99.5127
R15939 vdd.n2129 vdd.n837 99.5127
R15940 vdd.n2129 vdd.n827 99.5127
R15941 vdd.n2137 vdd.n827 99.5127
R15942 vdd.n2137 vdd.n825 99.5127
R15943 vdd.n2141 vdd.n825 99.5127
R15944 vdd.n2141 vdd.n816 99.5127
R15945 vdd.n2149 vdd.n816 99.5127
R15946 vdd.n2149 vdd.n814 99.5127
R15947 vdd.n2153 vdd.n814 99.5127
R15948 vdd.n2153 vdd.n803 99.5127
R15949 vdd.n2163 vdd.n803 99.5127
R15950 vdd.n2163 vdd.n800 99.5127
R15951 vdd.n2168 vdd.n800 99.5127
R15952 vdd.n2168 vdd.n801 99.5127
R15953 vdd.n801 vdd.n782 99.5127
R15954 vdd.n2686 vdd.n2685 99.5127
R15955 vdd.n2683 vdd.n2649 99.5127
R15956 vdd.n2679 vdd.n2678 99.5127
R15957 vdd.n2676 vdd.n2652 99.5127
R15958 vdd.n2672 vdd.n2671 99.5127
R15959 vdd.n2669 vdd.n2655 99.5127
R15960 vdd.n2665 vdd.n2664 99.5127
R15961 vdd.n2662 vdd.n2659 99.5127
R15962 vdd.n2803 vdd.n612 99.5127
R15963 vdd.n2801 vdd.n2800 99.5127
R15964 vdd.n2798 vdd.n615 99.5127
R15965 vdd.n2794 vdd.n2793 99.5127
R15966 vdd.n2791 vdd.n618 99.5127
R15967 vdd.n2787 vdd.n2786 99.5127
R15968 vdd.n2784 vdd.n621 99.5127
R15969 vdd.n2780 vdd.n2779 99.5127
R15970 vdd.n2777 vdd.n624 99.5127
R15971 vdd.n2421 vdd.n743 99.5127
R15972 vdd.n2421 vdd.n738 99.5127
R15973 vdd.n2492 vdd.n738 99.5127
R15974 vdd.n2492 vdd.n733 99.5127
R15975 vdd.n2488 vdd.n733 99.5127
R15976 vdd.n2488 vdd.n727 99.5127
R15977 vdd.n2485 vdd.n727 99.5127
R15978 vdd.n2485 vdd.n720 99.5127
R15979 vdd.n2482 vdd.n720 99.5127
R15980 vdd.n2482 vdd.n715 99.5127
R15981 vdd.n2479 vdd.n715 99.5127
R15982 vdd.n2479 vdd.n710 99.5127
R15983 vdd.n2476 vdd.n710 99.5127
R15984 vdd.n2476 vdd.n704 99.5127
R15985 vdd.n2473 vdd.n704 99.5127
R15986 vdd.n2473 vdd.n697 99.5127
R15987 vdd.n2438 vdd.n697 99.5127
R15988 vdd.n2438 vdd.n692 99.5127
R15989 vdd.n2435 vdd.n692 99.5127
R15990 vdd.n2435 vdd.n687 99.5127
R15991 vdd.n2432 vdd.n687 99.5127
R15992 vdd.n2432 vdd.n681 99.5127
R15993 vdd.n2429 vdd.n681 99.5127
R15994 vdd.n2429 vdd.n673 99.5127
R15995 vdd.n2426 vdd.n673 99.5127
R15996 vdd.n2426 vdd.n666 99.5127
R15997 vdd.n666 vdd.n630 99.5127
R15998 vdd.n2772 vdd.n630 99.5127
R15999 vdd.n2571 vdd.n746 99.5127
R16000 vdd.n2359 vdd.n2358 99.5127
R16001 vdd.n2363 vdd.n2362 99.5127
R16002 vdd.n2367 vdd.n2366 99.5127
R16003 vdd.n2371 vdd.n2370 99.5127
R16004 vdd.n2375 vdd.n2374 99.5127
R16005 vdd.n2379 vdd.n2378 99.5127
R16006 vdd.n2383 vdd.n2382 99.5127
R16007 vdd.n2387 vdd.n2386 99.5127
R16008 vdd.n2391 vdd.n2390 99.5127
R16009 vdd.n2395 vdd.n2394 99.5127
R16010 vdd.n2399 vdd.n2398 99.5127
R16011 vdd.n2403 vdd.n2402 99.5127
R16012 vdd.n2407 vdd.n2406 99.5127
R16013 vdd.n2411 vdd.n2410 99.5127
R16014 vdd.n2415 vdd.n2414 99.5127
R16015 vdd.n2417 vdd.n2349 99.5127
R16016 vdd.n2575 vdd.n736 99.5127
R16017 vdd.n2583 vdd.n736 99.5127
R16018 vdd.n2583 vdd.n734 99.5127
R16019 vdd.n2587 vdd.n734 99.5127
R16020 vdd.n2587 vdd.n724 99.5127
R16021 vdd.n2595 vdd.n724 99.5127
R16022 vdd.n2595 vdd.n722 99.5127
R16023 vdd.n2599 vdd.n722 99.5127
R16024 vdd.n2599 vdd.n713 99.5127
R16025 vdd.n2607 vdd.n713 99.5127
R16026 vdd.n2607 vdd.n711 99.5127
R16027 vdd.n2611 vdd.n711 99.5127
R16028 vdd.n2611 vdd.n701 99.5127
R16029 vdd.n2619 vdd.n701 99.5127
R16030 vdd.n2619 vdd.n699 99.5127
R16031 vdd.n2623 vdd.n699 99.5127
R16032 vdd.n2623 vdd.n690 99.5127
R16033 vdd.n2631 vdd.n690 99.5127
R16034 vdd.n2631 vdd.n688 99.5127
R16035 vdd.n2637 vdd.n688 99.5127
R16036 vdd.n2637 vdd.n678 99.5127
R16037 vdd.n2645 vdd.n678 99.5127
R16038 vdd.n2645 vdd.n675 99.5127
R16039 vdd.n2694 vdd.n675 99.5127
R16040 vdd.n2694 vdd.n676 99.5127
R16041 vdd.n676 vdd.n667 99.5127
R16042 vdd.n2689 vdd.n667 99.5127
R16043 vdd.n2689 vdd.n633 99.5127
R16044 vdd.n2239 vdd.n2238 99.5127
R16045 vdd.n2235 vdd.n2234 99.5127
R16046 vdd.n2231 vdd.n2230 99.5127
R16047 vdd.n2227 vdd.n2226 99.5127
R16048 vdd.n2223 vdd.n2222 99.5127
R16049 vdd.n2219 vdd.n2218 99.5127
R16050 vdd.n2215 vdd.n2214 99.5127
R16051 vdd.n2211 vdd.n2210 99.5127
R16052 vdd.n2207 vdd.n2206 99.5127
R16053 vdd.n2203 vdd.n2202 99.5127
R16054 vdd.n2199 vdd.n2198 99.5127
R16055 vdd.n2195 vdd.n2194 99.5127
R16056 vdd.n2191 vdd.n2190 99.5127
R16057 vdd.n2187 vdd.n2186 99.5127
R16058 vdd.n2183 vdd.n2182 99.5127
R16059 vdd.n2179 vdd.n2178 99.5127
R16060 vdd.n2175 vdd.n764 99.5127
R16061 vdd.n1932 vdd.n879 99.5127
R16062 vdd.n1932 vdd.n873 99.5127
R16063 vdd.n1935 vdd.n873 99.5127
R16064 vdd.n1935 vdd.n867 99.5127
R16065 vdd.n1938 vdd.n867 99.5127
R16066 vdd.n1938 vdd.n860 99.5127
R16067 vdd.n1941 vdd.n860 99.5127
R16068 vdd.n1941 vdd.n853 99.5127
R16069 vdd.n1944 vdd.n853 99.5127
R16070 vdd.n1944 vdd.n848 99.5127
R16071 vdd.n1947 vdd.n848 99.5127
R16072 vdd.n1947 vdd.n842 99.5127
R16073 vdd.n1968 vdd.n842 99.5127
R16074 vdd.n1968 vdd.n835 99.5127
R16075 vdd.n1964 vdd.n835 99.5127
R16076 vdd.n1964 vdd.n829 99.5127
R16077 vdd.n1961 vdd.n829 99.5127
R16078 vdd.n1961 vdd.n824 99.5127
R16079 vdd.n1958 vdd.n824 99.5127
R16080 vdd.n1958 vdd.n819 99.5127
R16081 vdd.n1955 vdd.n819 99.5127
R16082 vdd.n1955 vdd.n813 99.5127
R16083 vdd.n1952 vdd.n813 99.5127
R16084 vdd.n1952 vdd.n806 99.5127
R16085 vdd.n806 vdd.n797 99.5127
R16086 vdd.n2170 vdd.n797 99.5127
R16087 vdd.n2171 vdd.n2170 99.5127
R16088 vdd.n2171 vdd.n789 99.5127
R16089 vdd.n2082 vdd.n2080 99.5127
R16090 vdd.n2078 vdd.n882 99.5127
R16091 vdd.n2074 vdd.n2072 99.5127
R16092 vdd.n2070 vdd.n884 99.5127
R16093 vdd.n2066 vdd.n2064 99.5127
R16094 vdd.n2062 vdd.n886 99.5127
R16095 vdd.n2058 vdd.n2056 99.5127
R16096 vdd.n2054 vdd.n888 99.5127
R16097 vdd.n1896 vdd.n890 99.5127
R16098 vdd.n1901 vdd.n1898 99.5127
R16099 vdd.n1905 vdd.n1903 99.5127
R16100 vdd.n1909 vdd.n1894 99.5127
R16101 vdd.n1913 vdd.n1911 99.5127
R16102 vdd.n1917 vdd.n1892 99.5127
R16103 vdd.n1921 vdd.n1919 99.5127
R16104 vdd.n1926 vdd.n1888 99.5127
R16105 vdd.n1929 vdd.n1928 99.5127
R16106 vdd.n2086 vdd.n870 99.5127
R16107 vdd.n2094 vdd.n870 99.5127
R16108 vdd.n2094 vdd.n868 99.5127
R16109 vdd.n2098 vdd.n868 99.5127
R16110 vdd.n2098 vdd.n857 99.5127
R16111 vdd.n2106 vdd.n857 99.5127
R16112 vdd.n2106 vdd.n854 99.5127
R16113 vdd.n2111 vdd.n854 99.5127
R16114 vdd.n2111 vdd.n845 99.5127
R16115 vdd.n2119 vdd.n845 99.5127
R16116 vdd.n2119 vdd.n843 99.5127
R16117 vdd.n2123 vdd.n843 99.5127
R16118 vdd.n2123 vdd.n833 99.5127
R16119 vdd.n2131 vdd.n833 99.5127
R16120 vdd.n2131 vdd.n831 99.5127
R16121 vdd.n2135 vdd.n831 99.5127
R16122 vdd.n2135 vdd.n822 99.5127
R16123 vdd.n2143 vdd.n822 99.5127
R16124 vdd.n2143 vdd.n820 99.5127
R16125 vdd.n2147 vdd.n820 99.5127
R16126 vdd.n2147 vdd.n810 99.5127
R16127 vdd.n2155 vdd.n810 99.5127
R16128 vdd.n2155 vdd.n807 99.5127
R16129 vdd.n2161 vdd.n807 99.5127
R16130 vdd.n2161 vdd.n808 99.5127
R16131 vdd.n808 vdd.n799 99.5127
R16132 vdd.n799 vdd.n790 99.5127
R16133 vdd.n2243 vdd.n790 99.5127
R16134 vdd.n9 vdd.n7 98.9633
R16135 vdd.n2 vdd.n0 98.9633
R16136 vdd.n9 vdd.n8 98.6055
R16137 vdd.n11 vdd.n10 98.6055
R16138 vdd.n13 vdd.n12 98.6055
R16139 vdd.n6 vdd.n5 98.6055
R16140 vdd.n4 vdd.n3 98.6055
R16141 vdd.n2 vdd.n1 98.6055
R16142 vdd.t198 vdd.n279 85.8723
R16143 vdd.t169 vdd.n228 85.8723
R16144 vdd.t162 vdd.n185 85.8723
R16145 vdd.t224 vdd.n134 85.8723
R16146 vdd.t5 vdd.n92 85.8723
R16147 vdd.t83 vdd.n41 85.8723
R16148 vdd.t9 vdd.n1474 85.8723
R16149 vdd.t187 vdd.n1525 85.8723
R16150 vdd.t219 vdd.n1380 85.8723
R16151 vdd.t201 vdd.n1431 85.8723
R16152 vdd.t84 vdd.n1287 85.8723
R16153 vdd.t231 vdd.n1338 85.8723
R16154 vdd.n2635 vdd.n2634 78.546
R16155 vdd.n2109 vdd.n855 78.546
R16156 vdd.n266 vdd.n265 75.1835
R16157 vdd.n264 vdd.n263 75.1835
R16158 vdd.n262 vdd.n261 75.1835
R16159 vdd.n260 vdd.n259 75.1835
R16160 vdd.n258 vdd.n257 75.1835
R16161 vdd.n172 vdd.n171 75.1835
R16162 vdd.n170 vdd.n169 75.1835
R16163 vdd.n168 vdd.n167 75.1835
R16164 vdd.n166 vdd.n165 75.1835
R16165 vdd.n164 vdd.n163 75.1835
R16166 vdd.n79 vdd.n78 75.1835
R16167 vdd.n77 vdd.n76 75.1835
R16168 vdd.n75 vdd.n74 75.1835
R16169 vdd.n73 vdd.n72 75.1835
R16170 vdd.n71 vdd.n70 75.1835
R16171 vdd.n1504 vdd.n1503 75.1835
R16172 vdd.n1506 vdd.n1505 75.1835
R16173 vdd.n1508 vdd.n1507 75.1835
R16174 vdd.n1510 vdd.n1509 75.1835
R16175 vdd.n1512 vdd.n1511 75.1835
R16176 vdd.n1410 vdd.n1409 75.1835
R16177 vdd.n1412 vdd.n1411 75.1835
R16178 vdd.n1414 vdd.n1413 75.1835
R16179 vdd.n1416 vdd.n1415 75.1835
R16180 vdd.n1418 vdd.n1417 75.1835
R16181 vdd.n1317 vdd.n1316 75.1835
R16182 vdd.n1319 vdd.n1318 75.1835
R16183 vdd.n1321 vdd.n1320 75.1835
R16184 vdd.n1323 vdd.n1322 75.1835
R16185 vdd.n1325 vdd.n1324 75.1835
R16186 vdd.n2570 vdd.n2569 72.8958
R16187 vdd.n2569 vdd.n2333 72.8958
R16188 vdd.n2569 vdd.n2334 72.8958
R16189 vdd.n2569 vdd.n2335 72.8958
R16190 vdd.n2569 vdd.n2336 72.8958
R16191 vdd.n2569 vdd.n2337 72.8958
R16192 vdd.n2569 vdd.n2338 72.8958
R16193 vdd.n2569 vdd.n2339 72.8958
R16194 vdd.n2569 vdd.n2340 72.8958
R16195 vdd.n2569 vdd.n2341 72.8958
R16196 vdd.n2569 vdd.n2342 72.8958
R16197 vdd.n2569 vdd.n2343 72.8958
R16198 vdd.n2569 vdd.n2344 72.8958
R16199 vdd.n2569 vdd.n2345 72.8958
R16200 vdd.n2569 vdd.n2346 72.8958
R16201 vdd.n2569 vdd.n2347 72.8958
R16202 vdd.n2569 vdd.n2348 72.8958
R16203 vdd.n629 vdd.n613 72.8958
R16204 vdd.n2778 vdd.n613 72.8958
R16205 vdd.n623 vdd.n613 72.8958
R16206 vdd.n2785 vdd.n613 72.8958
R16207 vdd.n620 vdd.n613 72.8958
R16208 vdd.n2792 vdd.n613 72.8958
R16209 vdd.n617 vdd.n613 72.8958
R16210 vdd.n2799 vdd.n613 72.8958
R16211 vdd.n2802 vdd.n613 72.8958
R16212 vdd.n2658 vdd.n613 72.8958
R16213 vdd.n2663 vdd.n613 72.8958
R16214 vdd.n2657 vdd.n613 72.8958
R16215 vdd.n2670 vdd.n613 72.8958
R16216 vdd.n2654 vdd.n613 72.8958
R16217 vdd.n2677 vdd.n613 72.8958
R16218 vdd.n2651 vdd.n613 72.8958
R16219 vdd.n2684 vdd.n613 72.8958
R16220 vdd.n1822 vdd.n877 72.8958
R16221 vdd.n1828 vdd.n877 72.8958
R16222 vdd.n1830 vdd.n877 72.8958
R16223 vdd.n1836 vdd.n877 72.8958
R16224 vdd.n1838 vdd.n877 72.8958
R16225 vdd.n1844 vdd.n877 72.8958
R16226 vdd.n1846 vdd.n877 72.8958
R16227 vdd.n1852 vdd.n877 72.8958
R16228 vdd.n2023 vdd.n877 72.8958
R16229 vdd.n2021 vdd.n877 72.8958
R16230 vdd.n2015 vdd.n877 72.8958
R16231 vdd.n2013 vdd.n877 72.8958
R16232 vdd.n2007 vdd.n877 72.8958
R16233 vdd.n2005 vdd.n877 72.8958
R16234 vdd.n1999 vdd.n877 72.8958
R16235 vdd.n1997 vdd.n877 72.8958
R16236 vdd.n1991 vdd.n877 72.8958
R16237 vdd.n2316 vdd.n765 72.8958
R16238 vdd.n2316 vdd.n766 72.8958
R16239 vdd.n2316 vdd.n767 72.8958
R16240 vdd.n2316 vdd.n768 72.8958
R16241 vdd.n2316 vdd.n769 72.8958
R16242 vdd.n2316 vdd.n770 72.8958
R16243 vdd.n2316 vdd.n771 72.8958
R16244 vdd.n2316 vdd.n772 72.8958
R16245 vdd.n2316 vdd.n773 72.8958
R16246 vdd.n2316 vdd.n774 72.8958
R16247 vdd.n2316 vdd.n775 72.8958
R16248 vdd.n2316 vdd.n776 72.8958
R16249 vdd.n2316 vdd.n777 72.8958
R16250 vdd.n2316 vdd.n778 72.8958
R16251 vdd.n2316 vdd.n779 72.8958
R16252 vdd.n2316 vdd.n780 72.8958
R16253 vdd.n2316 vdd.n781 72.8958
R16254 vdd.n2569 vdd.n2568 72.8958
R16255 vdd.n2569 vdd.n2317 72.8958
R16256 vdd.n2569 vdd.n2318 72.8958
R16257 vdd.n2569 vdd.n2319 72.8958
R16258 vdd.n2569 vdd.n2320 72.8958
R16259 vdd.n2569 vdd.n2321 72.8958
R16260 vdd.n2569 vdd.n2322 72.8958
R16261 vdd.n2569 vdd.n2323 72.8958
R16262 vdd.n2569 vdd.n2324 72.8958
R16263 vdd.n2569 vdd.n2325 72.8958
R16264 vdd.n2569 vdd.n2326 72.8958
R16265 vdd.n2569 vdd.n2327 72.8958
R16266 vdd.n2569 vdd.n2328 72.8958
R16267 vdd.n2569 vdd.n2329 72.8958
R16268 vdd.n2569 vdd.n2330 72.8958
R16269 vdd.n2569 vdd.n2331 72.8958
R16270 vdd.n2569 vdd.n2332 72.8958
R16271 vdd.n2706 vdd.n613 72.8958
R16272 vdd.n2712 vdd.n613 72.8958
R16273 vdd.n659 vdd.n613 72.8958
R16274 vdd.n2719 vdd.n613 72.8958
R16275 vdd.n656 vdd.n613 72.8958
R16276 vdd.n2726 vdd.n613 72.8958
R16277 vdd.n653 vdd.n613 72.8958
R16278 vdd.n2733 vdd.n613 72.8958
R16279 vdd.n650 vdd.n613 72.8958
R16280 vdd.n2741 vdd.n613 72.8958
R16281 vdd.n647 vdd.n613 72.8958
R16282 vdd.n2748 vdd.n613 72.8958
R16283 vdd.n644 vdd.n613 72.8958
R16284 vdd.n2755 vdd.n613 72.8958
R16285 vdd.n641 vdd.n613 72.8958
R16286 vdd.n2762 vdd.n613 72.8958
R16287 vdd.n2765 vdd.n613 72.8958
R16288 vdd.n2316 vdd.n763 72.8958
R16289 vdd.n2316 vdd.n762 72.8958
R16290 vdd.n2316 vdd.n761 72.8958
R16291 vdd.n2316 vdd.n760 72.8958
R16292 vdd.n2316 vdd.n759 72.8958
R16293 vdd.n2316 vdd.n758 72.8958
R16294 vdd.n2316 vdd.n757 72.8958
R16295 vdd.n2316 vdd.n756 72.8958
R16296 vdd.n2316 vdd.n755 72.8958
R16297 vdd.n2316 vdd.n754 72.8958
R16298 vdd.n2316 vdd.n753 72.8958
R16299 vdd.n2316 vdd.n752 72.8958
R16300 vdd.n2316 vdd.n751 72.8958
R16301 vdd.n2316 vdd.n750 72.8958
R16302 vdd.n2316 vdd.n749 72.8958
R16303 vdd.n2316 vdd.n748 72.8958
R16304 vdd.n2316 vdd.n747 72.8958
R16305 vdd.n2081 vdd.n877 72.8958
R16306 vdd.n2079 vdd.n877 72.8958
R16307 vdd.n2073 vdd.n877 72.8958
R16308 vdd.n2071 vdd.n877 72.8958
R16309 vdd.n2065 vdd.n877 72.8958
R16310 vdd.n2063 vdd.n877 72.8958
R16311 vdd.n2057 vdd.n877 72.8958
R16312 vdd.n2055 vdd.n877 72.8958
R16313 vdd.n889 vdd.n877 72.8958
R16314 vdd.n1897 vdd.n877 72.8958
R16315 vdd.n1902 vdd.n877 72.8958
R16316 vdd.n1904 vdd.n877 72.8958
R16317 vdd.n1910 vdd.n877 72.8958
R16318 vdd.n1912 vdd.n877 72.8958
R16319 vdd.n1918 vdd.n877 72.8958
R16320 vdd.n1920 vdd.n877 72.8958
R16321 vdd.n1927 vdd.n877 72.8958
R16322 vdd.n986 vdd.n982 66.2847
R16323 vdd.n992 vdd.n982 66.2847
R16324 vdd.n995 vdd.n982 66.2847
R16325 vdd.n1000 vdd.n982 66.2847
R16326 vdd.n1003 vdd.n982 66.2847
R16327 vdd.n1008 vdd.n982 66.2847
R16328 vdd.n1011 vdd.n982 66.2847
R16329 vdd.n1016 vdd.n982 66.2847
R16330 vdd.n1019 vdd.n982 66.2847
R16331 vdd.n1026 vdd.n982 66.2847
R16332 vdd.n1029 vdd.n982 66.2847
R16333 vdd.n1034 vdd.n982 66.2847
R16334 vdd.n1037 vdd.n982 66.2847
R16335 vdd.n1042 vdd.n982 66.2847
R16336 vdd.n1045 vdd.n982 66.2847
R16337 vdd.n1050 vdd.n982 66.2847
R16338 vdd.n1053 vdd.n982 66.2847
R16339 vdd.n1058 vdd.n982 66.2847
R16340 vdd.n1061 vdd.n982 66.2847
R16341 vdd.n1066 vdd.n982 66.2847
R16342 vdd.n1145 vdd.n982 66.2847
R16343 vdd.n1069 vdd.n982 66.2847
R16344 vdd.n1075 vdd.n982 66.2847
R16345 vdd.n1080 vdd.n982 66.2847
R16346 vdd.n1083 vdd.n982 66.2847
R16347 vdd.n1088 vdd.n982 66.2847
R16348 vdd.n1091 vdd.n982 66.2847
R16349 vdd.n1096 vdd.n982 66.2847
R16350 vdd.n1099 vdd.n982 66.2847
R16351 vdd.n1104 vdd.n982 66.2847
R16352 vdd.n1107 vdd.n982 66.2847
R16353 vdd.n901 vdd.n898 66.2847
R16354 vdd.n1712 vdd.n901 66.2847
R16355 vdd.n1717 vdd.n901 66.2847
R16356 vdd.n1722 vdd.n901 66.2847
R16357 vdd.n1710 vdd.n901 66.2847
R16358 vdd.n1729 vdd.n901 66.2847
R16359 vdd.n1702 vdd.n901 66.2847
R16360 vdd.n1736 vdd.n901 66.2847
R16361 vdd.n1695 vdd.n901 66.2847
R16362 vdd.n1743 vdd.n901 66.2847
R16363 vdd.n1689 vdd.n901 66.2847
R16364 vdd.n1684 vdd.n901 66.2847
R16365 vdd.n1754 vdd.n901 66.2847
R16366 vdd.n1676 vdd.n901 66.2847
R16367 vdd.n1761 vdd.n901 66.2847
R16368 vdd.n1669 vdd.n901 66.2847
R16369 vdd.n1768 vdd.n901 66.2847
R16370 vdd.n1662 vdd.n901 66.2847
R16371 vdd.n1775 vdd.n901 66.2847
R16372 vdd.n1655 vdd.n901 66.2847
R16373 vdd.n1782 vdd.n901 66.2847
R16374 vdd.n1649 vdd.n901 66.2847
R16375 vdd.n1644 vdd.n901 66.2847
R16376 vdd.n1793 vdd.n901 66.2847
R16377 vdd.n1636 vdd.n901 66.2847
R16378 vdd.n1800 vdd.n901 66.2847
R16379 vdd.n1629 vdd.n901 66.2847
R16380 vdd.n1807 vdd.n901 66.2847
R16381 vdd.n1810 vdd.n901 66.2847
R16382 vdd.n1620 vdd.n901 66.2847
R16383 vdd.n2032 vdd.n901 66.2847
R16384 vdd.n1614 vdd.n901 66.2847
R16385 vdd.n2932 vdd.n516 66.2847
R16386 vdd.n520 vdd.n516 66.2847
R16387 vdd.n523 vdd.n516 66.2847
R16388 vdd.n2921 vdd.n516 66.2847
R16389 vdd.n2915 vdd.n516 66.2847
R16390 vdd.n2913 vdd.n516 66.2847
R16391 vdd.n2907 vdd.n516 66.2847
R16392 vdd.n2905 vdd.n516 66.2847
R16393 vdd.n2899 vdd.n516 66.2847
R16394 vdd.n2897 vdd.n516 66.2847
R16395 vdd.n2891 vdd.n516 66.2847
R16396 vdd.n2889 vdd.n516 66.2847
R16397 vdd.n2883 vdd.n516 66.2847
R16398 vdd.n2881 vdd.n516 66.2847
R16399 vdd.n2875 vdd.n516 66.2847
R16400 vdd.n2873 vdd.n516 66.2847
R16401 vdd.n2867 vdd.n516 66.2847
R16402 vdd.n2865 vdd.n516 66.2847
R16403 vdd.n2859 vdd.n516 66.2847
R16404 vdd.n2857 vdd.n516 66.2847
R16405 vdd.n584 vdd.n516 66.2847
R16406 vdd.n2848 vdd.n516 66.2847
R16407 vdd.n586 vdd.n516 66.2847
R16408 vdd.n2841 vdd.n516 66.2847
R16409 vdd.n2835 vdd.n516 66.2847
R16410 vdd.n2833 vdd.n516 66.2847
R16411 vdd.n2827 vdd.n516 66.2847
R16412 vdd.n2825 vdd.n516 66.2847
R16413 vdd.n2819 vdd.n516 66.2847
R16414 vdd.n607 vdd.n516 66.2847
R16415 vdd.n609 vdd.n516 66.2847
R16416 vdd.n3018 vdd.n351 66.2847
R16417 vdd.n3027 vdd.n351 66.2847
R16418 vdd.n461 vdd.n351 66.2847
R16419 vdd.n3034 vdd.n351 66.2847
R16420 vdd.n454 vdd.n351 66.2847
R16421 vdd.n3041 vdd.n351 66.2847
R16422 vdd.n447 vdd.n351 66.2847
R16423 vdd.n3048 vdd.n351 66.2847
R16424 vdd.n440 vdd.n351 66.2847
R16425 vdd.n3055 vdd.n351 66.2847
R16426 vdd.n434 vdd.n351 66.2847
R16427 vdd.n429 vdd.n351 66.2847
R16428 vdd.n3066 vdd.n351 66.2847
R16429 vdd.n421 vdd.n351 66.2847
R16430 vdd.n3073 vdd.n351 66.2847
R16431 vdd.n414 vdd.n351 66.2847
R16432 vdd.n3080 vdd.n351 66.2847
R16433 vdd.n407 vdd.n351 66.2847
R16434 vdd.n3087 vdd.n351 66.2847
R16435 vdd.n400 vdd.n351 66.2847
R16436 vdd.n3094 vdd.n351 66.2847
R16437 vdd.n394 vdd.n351 66.2847
R16438 vdd.n389 vdd.n351 66.2847
R16439 vdd.n3105 vdd.n351 66.2847
R16440 vdd.n381 vdd.n351 66.2847
R16441 vdd.n3112 vdd.n351 66.2847
R16442 vdd.n374 vdd.n351 66.2847
R16443 vdd.n3119 vdd.n351 66.2847
R16444 vdd.n367 vdd.n351 66.2847
R16445 vdd.n3126 vdd.n351 66.2847
R16446 vdd.n3129 vdd.n351 66.2847
R16447 vdd.n355 vdd.n351 66.2847
R16448 vdd.n356 vdd.n355 52.4337
R16449 vdd.n3129 vdd.n3128 52.4337
R16450 vdd.n3126 vdd.n3125 52.4337
R16451 vdd.n3121 vdd.n367 52.4337
R16452 vdd.n3119 vdd.n3118 52.4337
R16453 vdd.n3114 vdd.n374 52.4337
R16454 vdd.n3112 vdd.n3111 52.4337
R16455 vdd.n3107 vdd.n381 52.4337
R16456 vdd.n3105 vdd.n3104 52.4337
R16457 vdd.n390 vdd.n389 52.4337
R16458 vdd.n3096 vdd.n394 52.4337
R16459 vdd.n3094 vdd.n3093 52.4337
R16460 vdd.n3089 vdd.n400 52.4337
R16461 vdd.n3087 vdd.n3086 52.4337
R16462 vdd.n3082 vdd.n407 52.4337
R16463 vdd.n3080 vdd.n3079 52.4337
R16464 vdd.n3075 vdd.n414 52.4337
R16465 vdd.n3073 vdd.n3072 52.4337
R16466 vdd.n3068 vdd.n421 52.4337
R16467 vdd.n3066 vdd.n3065 52.4337
R16468 vdd.n430 vdd.n429 52.4337
R16469 vdd.n3057 vdd.n434 52.4337
R16470 vdd.n3055 vdd.n3054 52.4337
R16471 vdd.n3050 vdd.n440 52.4337
R16472 vdd.n3048 vdd.n3047 52.4337
R16473 vdd.n3043 vdd.n447 52.4337
R16474 vdd.n3041 vdd.n3040 52.4337
R16475 vdd.n3036 vdd.n454 52.4337
R16476 vdd.n3034 vdd.n3033 52.4337
R16477 vdd.n3029 vdd.n461 52.4337
R16478 vdd.n3027 vdd.n3026 52.4337
R16479 vdd.n3019 vdd.n3018 52.4337
R16480 vdd.n2932 vdd.n517 52.4337
R16481 vdd.n2930 vdd.n520 52.4337
R16482 vdd.n2926 vdd.n523 52.4337
R16483 vdd.n2922 vdd.n2921 52.4337
R16484 vdd.n2915 vdd.n526 52.4337
R16485 vdd.n2914 vdd.n2913 52.4337
R16486 vdd.n2907 vdd.n532 52.4337
R16487 vdd.n2906 vdd.n2905 52.4337
R16488 vdd.n2899 vdd.n538 52.4337
R16489 vdd.n2898 vdd.n2897 52.4337
R16490 vdd.n2891 vdd.n546 52.4337
R16491 vdd.n2890 vdd.n2889 52.4337
R16492 vdd.n2883 vdd.n552 52.4337
R16493 vdd.n2882 vdd.n2881 52.4337
R16494 vdd.n2875 vdd.n558 52.4337
R16495 vdd.n2874 vdd.n2873 52.4337
R16496 vdd.n2867 vdd.n564 52.4337
R16497 vdd.n2866 vdd.n2865 52.4337
R16498 vdd.n2859 vdd.n570 52.4337
R16499 vdd.n2858 vdd.n2857 52.4337
R16500 vdd.n584 vdd.n576 52.4337
R16501 vdd.n2849 vdd.n2848 52.4337
R16502 vdd.n2846 vdd.n586 52.4337
R16503 vdd.n2842 vdd.n2841 52.4337
R16504 vdd.n2835 vdd.n590 52.4337
R16505 vdd.n2834 vdd.n2833 52.4337
R16506 vdd.n2827 vdd.n596 52.4337
R16507 vdd.n2826 vdd.n2825 52.4337
R16508 vdd.n2819 vdd.n602 52.4337
R16509 vdd.n2818 vdd.n607 52.4337
R16510 vdd.n2814 vdd.n609 52.4337
R16511 vdd.n2034 vdd.n1614 52.4337
R16512 vdd.n2032 vdd.n2031 52.4337
R16513 vdd.n1621 vdd.n1620 52.4337
R16514 vdd.n1810 vdd.n1809 52.4337
R16515 vdd.n1807 vdd.n1806 52.4337
R16516 vdd.n1802 vdd.n1629 52.4337
R16517 vdd.n1800 vdd.n1799 52.4337
R16518 vdd.n1795 vdd.n1636 52.4337
R16519 vdd.n1793 vdd.n1792 52.4337
R16520 vdd.n1645 vdd.n1644 52.4337
R16521 vdd.n1784 vdd.n1649 52.4337
R16522 vdd.n1782 vdd.n1781 52.4337
R16523 vdd.n1777 vdd.n1655 52.4337
R16524 vdd.n1775 vdd.n1774 52.4337
R16525 vdd.n1770 vdd.n1662 52.4337
R16526 vdd.n1768 vdd.n1767 52.4337
R16527 vdd.n1763 vdd.n1669 52.4337
R16528 vdd.n1761 vdd.n1760 52.4337
R16529 vdd.n1756 vdd.n1676 52.4337
R16530 vdd.n1754 vdd.n1753 52.4337
R16531 vdd.n1685 vdd.n1684 52.4337
R16532 vdd.n1745 vdd.n1689 52.4337
R16533 vdd.n1743 vdd.n1742 52.4337
R16534 vdd.n1738 vdd.n1695 52.4337
R16535 vdd.n1736 vdd.n1735 52.4337
R16536 vdd.n1731 vdd.n1702 52.4337
R16537 vdd.n1729 vdd.n1728 52.4337
R16538 vdd.n1724 vdd.n1710 52.4337
R16539 vdd.n1722 vdd.n1721 52.4337
R16540 vdd.n1717 vdd.n1716 52.4337
R16541 vdd.n1712 vdd.n1711 52.4337
R16542 vdd.n2043 vdd.n898 52.4337
R16543 vdd.n986 vdd.n984 52.4337
R16544 vdd.n992 vdd.n991 52.4337
R16545 vdd.n995 vdd.n994 52.4337
R16546 vdd.n1000 vdd.n999 52.4337
R16547 vdd.n1003 vdd.n1002 52.4337
R16548 vdd.n1008 vdd.n1007 52.4337
R16549 vdd.n1011 vdd.n1010 52.4337
R16550 vdd.n1016 vdd.n1015 52.4337
R16551 vdd.n1019 vdd.n1018 52.4337
R16552 vdd.n1026 vdd.n1025 52.4337
R16553 vdd.n1029 vdd.n1028 52.4337
R16554 vdd.n1034 vdd.n1033 52.4337
R16555 vdd.n1037 vdd.n1036 52.4337
R16556 vdd.n1042 vdd.n1041 52.4337
R16557 vdd.n1045 vdd.n1044 52.4337
R16558 vdd.n1050 vdd.n1049 52.4337
R16559 vdd.n1053 vdd.n1052 52.4337
R16560 vdd.n1058 vdd.n1057 52.4337
R16561 vdd.n1061 vdd.n1060 52.4337
R16562 vdd.n1066 vdd.n1065 52.4337
R16563 vdd.n1146 vdd.n1145 52.4337
R16564 vdd.n1143 vdd.n1069 52.4337
R16565 vdd.n1075 vdd.n1074 52.4337
R16566 vdd.n1080 vdd.n1077 52.4337
R16567 vdd.n1083 vdd.n1082 52.4337
R16568 vdd.n1088 vdd.n1085 52.4337
R16569 vdd.n1091 vdd.n1090 52.4337
R16570 vdd.n1096 vdd.n1093 52.4337
R16571 vdd.n1099 vdd.n1098 52.4337
R16572 vdd.n1104 vdd.n1101 52.4337
R16573 vdd.n1107 vdd.n1106 52.4337
R16574 vdd.n987 vdd.n986 52.4337
R16575 vdd.n993 vdd.n992 52.4337
R16576 vdd.n996 vdd.n995 52.4337
R16577 vdd.n1001 vdd.n1000 52.4337
R16578 vdd.n1004 vdd.n1003 52.4337
R16579 vdd.n1009 vdd.n1008 52.4337
R16580 vdd.n1012 vdd.n1011 52.4337
R16581 vdd.n1017 vdd.n1016 52.4337
R16582 vdd.n1020 vdd.n1019 52.4337
R16583 vdd.n1027 vdd.n1026 52.4337
R16584 vdd.n1030 vdd.n1029 52.4337
R16585 vdd.n1035 vdd.n1034 52.4337
R16586 vdd.n1038 vdd.n1037 52.4337
R16587 vdd.n1043 vdd.n1042 52.4337
R16588 vdd.n1046 vdd.n1045 52.4337
R16589 vdd.n1051 vdd.n1050 52.4337
R16590 vdd.n1054 vdd.n1053 52.4337
R16591 vdd.n1059 vdd.n1058 52.4337
R16592 vdd.n1062 vdd.n1061 52.4337
R16593 vdd.n1067 vdd.n1066 52.4337
R16594 vdd.n1145 vdd.n1144 52.4337
R16595 vdd.n1073 vdd.n1069 52.4337
R16596 vdd.n1076 vdd.n1075 52.4337
R16597 vdd.n1081 vdd.n1080 52.4337
R16598 vdd.n1084 vdd.n1083 52.4337
R16599 vdd.n1089 vdd.n1088 52.4337
R16600 vdd.n1092 vdd.n1091 52.4337
R16601 vdd.n1097 vdd.n1096 52.4337
R16602 vdd.n1100 vdd.n1099 52.4337
R16603 vdd.n1105 vdd.n1104 52.4337
R16604 vdd.n1108 vdd.n1107 52.4337
R16605 vdd.n898 vdd.n897 52.4337
R16606 vdd.n1713 vdd.n1712 52.4337
R16607 vdd.n1718 vdd.n1717 52.4337
R16608 vdd.n1723 vdd.n1722 52.4337
R16609 vdd.n1710 vdd.n1703 52.4337
R16610 vdd.n1730 vdd.n1729 52.4337
R16611 vdd.n1702 vdd.n1696 52.4337
R16612 vdd.n1737 vdd.n1736 52.4337
R16613 vdd.n1695 vdd.n1690 52.4337
R16614 vdd.n1744 vdd.n1743 52.4337
R16615 vdd.n1689 vdd.n1688 52.4337
R16616 vdd.n1684 vdd.n1677 52.4337
R16617 vdd.n1755 vdd.n1754 52.4337
R16618 vdd.n1676 vdd.n1670 52.4337
R16619 vdd.n1762 vdd.n1761 52.4337
R16620 vdd.n1669 vdd.n1663 52.4337
R16621 vdd.n1769 vdd.n1768 52.4337
R16622 vdd.n1662 vdd.n1656 52.4337
R16623 vdd.n1776 vdd.n1775 52.4337
R16624 vdd.n1655 vdd.n1650 52.4337
R16625 vdd.n1783 vdd.n1782 52.4337
R16626 vdd.n1649 vdd.n1648 52.4337
R16627 vdd.n1644 vdd.n1637 52.4337
R16628 vdd.n1794 vdd.n1793 52.4337
R16629 vdd.n1636 vdd.n1630 52.4337
R16630 vdd.n1801 vdd.n1800 52.4337
R16631 vdd.n1629 vdd.n1623 52.4337
R16632 vdd.n1808 vdd.n1807 52.4337
R16633 vdd.n1811 vdd.n1810 52.4337
R16634 vdd.n1620 vdd.n1615 52.4337
R16635 vdd.n2033 vdd.n2032 52.4337
R16636 vdd.n1614 vdd.n903 52.4337
R16637 vdd.n2933 vdd.n2932 52.4337
R16638 vdd.n2927 vdd.n520 52.4337
R16639 vdd.n2923 vdd.n523 52.4337
R16640 vdd.n2921 vdd.n2920 52.4337
R16641 vdd.n2916 vdd.n2915 52.4337
R16642 vdd.n2913 vdd.n2912 52.4337
R16643 vdd.n2908 vdd.n2907 52.4337
R16644 vdd.n2905 vdd.n2904 52.4337
R16645 vdd.n2900 vdd.n2899 52.4337
R16646 vdd.n2897 vdd.n2896 52.4337
R16647 vdd.n2892 vdd.n2891 52.4337
R16648 vdd.n2889 vdd.n2888 52.4337
R16649 vdd.n2884 vdd.n2883 52.4337
R16650 vdd.n2881 vdd.n2880 52.4337
R16651 vdd.n2876 vdd.n2875 52.4337
R16652 vdd.n2873 vdd.n2872 52.4337
R16653 vdd.n2868 vdd.n2867 52.4337
R16654 vdd.n2865 vdd.n2864 52.4337
R16655 vdd.n2860 vdd.n2859 52.4337
R16656 vdd.n2857 vdd.n2856 52.4337
R16657 vdd.n585 vdd.n584 52.4337
R16658 vdd.n2848 vdd.n2847 52.4337
R16659 vdd.n2843 vdd.n586 52.4337
R16660 vdd.n2841 vdd.n2840 52.4337
R16661 vdd.n2836 vdd.n2835 52.4337
R16662 vdd.n2833 vdd.n2832 52.4337
R16663 vdd.n2828 vdd.n2827 52.4337
R16664 vdd.n2825 vdd.n2824 52.4337
R16665 vdd.n2820 vdd.n2819 52.4337
R16666 vdd.n2815 vdd.n607 52.4337
R16667 vdd.n2811 vdd.n609 52.4337
R16668 vdd.n3018 vdd.n462 52.4337
R16669 vdd.n3028 vdd.n3027 52.4337
R16670 vdd.n461 vdd.n455 52.4337
R16671 vdd.n3035 vdd.n3034 52.4337
R16672 vdd.n454 vdd.n448 52.4337
R16673 vdd.n3042 vdd.n3041 52.4337
R16674 vdd.n447 vdd.n441 52.4337
R16675 vdd.n3049 vdd.n3048 52.4337
R16676 vdd.n440 vdd.n435 52.4337
R16677 vdd.n3056 vdd.n3055 52.4337
R16678 vdd.n434 vdd.n433 52.4337
R16679 vdd.n429 vdd.n422 52.4337
R16680 vdd.n3067 vdd.n3066 52.4337
R16681 vdd.n421 vdd.n415 52.4337
R16682 vdd.n3074 vdd.n3073 52.4337
R16683 vdd.n414 vdd.n408 52.4337
R16684 vdd.n3081 vdd.n3080 52.4337
R16685 vdd.n407 vdd.n401 52.4337
R16686 vdd.n3088 vdd.n3087 52.4337
R16687 vdd.n400 vdd.n395 52.4337
R16688 vdd.n3095 vdd.n3094 52.4337
R16689 vdd.n394 vdd.n393 52.4337
R16690 vdd.n389 vdd.n382 52.4337
R16691 vdd.n3106 vdd.n3105 52.4337
R16692 vdd.n381 vdd.n375 52.4337
R16693 vdd.n3113 vdd.n3112 52.4337
R16694 vdd.n374 vdd.n368 52.4337
R16695 vdd.n3120 vdd.n3119 52.4337
R16696 vdd.n367 vdd.n360 52.4337
R16697 vdd.n3127 vdd.n3126 52.4337
R16698 vdd.n3130 vdd.n3129 52.4337
R16699 vdd.n355 vdd.n352 52.4337
R16700 vdd.t77 vdd.t176 51.4683
R16701 vdd.n258 vdd.n256 42.0461
R16702 vdd.n164 vdd.n162 42.0461
R16703 vdd.n71 vdd.n69 42.0461
R16704 vdd.n1504 vdd.n1502 42.0461
R16705 vdd.n1410 vdd.n1408 42.0461
R16706 vdd.n1317 vdd.n1315 42.0461
R16707 vdd.n308 vdd.n307 41.6884
R16708 vdd.n214 vdd.n213 41.6884
R16709 vdd.n121 vdd.n120 41.6884
R16710 vdd.n1554 vdd.n1553 41.6884
R16711 vdd.n1460 vdd.n1459 41.6884
R16712 vdd.n1367 vdd.n1366 41.6884
R16713 vdd.n1112 vdd.n1111 41.1157
R16714 vdd.n1149 vdd.n1148 41.1157
R16715 vdd.n1023 vdd.n1022 41.1157
R16716 vdd.n3023 vdd.n3022 41.1157
R16717 vdd.n3062 vdd.n428 41.1157
R16718 vdd.n3101 vdd.n388 41.1157
R16719 vdd.n2765 vdd.n2764 39.2114
R16720 vdd.n2762 vdd.n2761 39.2114
R16721 vdd.n2757 vdd.n641 39.2114
R16722 vdd.n2755 vdd.n2754 39.2114
R16723 vdd.n2750 vdd.n644 39.2114
R16724 vdd.n2748 vdd.n2747 39.2114
R16725 vdd.n2743 vdd.n647 39.2114
R16726 vdd.n2741 vdd.n2740 39.2114
R16727 vdd.n2735 vdd.n650 39.2114
R16728 vdd.n2733 vdd.n2732 39.2114
R16729 vdd.n2728 vdd.n653 39.2114
R16730 vdd.n2726 vdd.n2725 39.2114
R16731 vdd.n2721 vdd.n656 39.2114
R16732 vdd.n2719 vdd.n2718 39.2114
R16733 vdd.n2714 vdd.n659 39.2114
R16734 vdd.n2712 vdd.n2711 39.2114
R16735 vdd.n2707 vdd.n2706 39.2114
R16736 vdd.n2568 vdd.n741 39.2114
R16737 vdd.n2563 vdd.n2317 39.2114
R16738 vdd.n2560 vdd.n2318 39.2114
R16739 vdd.n2556 vdd.n2319 39.2114
R16740 vdd.n2552 vdd.n2320 39.2114
R16741 vdd.n2548 vdd.n2321 39.2114
R16742 vdd.n2544 vdd.n2322 39.2114
R16743 vdd.n2540 vdd.n2323 39.2114
R16744 vdd.n2536 vdd.n2324 39.2114
R16745 vdd.n2532 vdd.n2325 39.2114
R16746 vdd.n2528 vdd.n2326 39.2114
R16747 vdd.n2524 vdd.n2327 39.2114
R16748 vdd.n2520 vdd.n2328 39.2114
R16749 vdd.n2516 vdd.n2329 39.2114
R16750 vdd.n2512 vdd.n2330 39.2114
R16751 vdd.n2508 vdd.n2331 39.2114
R16752 vdd.n2503 vdd.n2332 39.2114
R16753 vdd.n2311 vdd.n781 39.2114
R16754 vdd.n2307 vdd.n780 39.2114
R16755 vdd.n2303 vdd.n779 39.2114
R16756 vdd.n2299 vdd.n778 39.2114
R16757 vdd.n2295 vdd.n777 39.2114
R16758 vdd.n2291 vdd.n776 39.2114
R16759 vdd.n2287 vdd.n775 39.2114
R16760 vdd.n2283 vdd.n774 39.2114
R16761 vdd.n2279 vdd.n773 39.2114
R16762 vdd.n2275 vdd.n772 39.2114
R16763 vdd.n2271 vdd.n771 39.2114
R16764 vdd.n2267 vdd.n770 39.2114
R16765 vdd.n2263 vdd.n769 39.2114
R16766 vdd.n2259 vdd.n768 39.2114
R16767 vdd.n2255 vdd.n767 39.2114
R16768 vdd.n2250 vdd.n766 39.2114
R16769 vdd.n2246 vdd.n765 39.2114
R16770 vdd.n1822 vdd.n876 39.2114
R16771 vdd.n1828 vdd.n1827 39.2114
R16772 vdd.n1831 vdd.n1830 39.2114
R16773 vdd.n1836 vdd.n1835 39.2114
R16774 vdd.n1839 vdd.n1838 39.2114
R16775 vdd.n1844 vdd.n1843 39.2114
R16776 vdd.n1847 vdd.n1846 39.2114
R16777 vdd.n1852 vdd.n1851 39.2114
R16778 vdd.n2023 vdd.n1854 39.2114
R16779 vdd.n2022 vdd.n2021 39.2114
R16780 vdd.n2015 vdd.n1856 39.2114
R16781 vdd.n2014 vdd.n2013 39.2114
R16782 vdd.n2007 vdd.n1858 39.2114
R16783 vdd.n2006 vdd.n2005 39.2114
R16784 vdd.n1999 vdd.n1860 39.2114
R16785 vdd.n1998 vdd.n1997 39.2114
R16786 vdd.n1991 vdd.n1862 39.2114
R16787 vdd.n2684 vdd.n2683 39.2114
R16788 vdd.n2679 vdd.n2651 39.2114
R16789 vdd.n2677 vdd.n2676 39.2114
R16790 vdd.n2672 vdd.n2654 39.2114
R16791 vdd.n2670 vdd.n2669 39.2114
R16792 vdd.n2665 vdd.n2657 39.2114
R16793 vdd.n2663 vdd.n2662 39.2114
R16794 vdd.n2658 vdd.n612 39.2114
R16795 vdd.n2802 vdd.n2801 39.2114
R16796 vdd.n2799 vdd.n2798 39.2114
R16797 vdd.n2794 vdd.n617 39.2114
R16798 vdd.n2792 vdd.n2791 39.2114
R16799 vdd.n2787 vdd.n620 39.2114
R16800 vdd.n2785 vdd.n2784 39.2114
R16801 vdd.n2780 vdd.n623 39.2114
R16802 vdd.n2778 vdd.n2777 39.2114
R16803 vdd.n2773 vdd.n629 39.2114
R16804 vdd.n2570 vdd.n744 39.2114
R16805 vdd.n2333 vdd.n746 39.2114
R16806 vdd.n2359 vdd.n2334 39.2114
R16807 vdd.n2363 vdd.n2335 39.2114
R16808 vdd.n2367 vdd.n2336 39.2114
R16809 vdd.n2371 vdd.n2337 39.2114
R16810 vdd.n2375 vdd.n2338 39.2114
R16811 vdd.n2379 vdd.n2339 39.2114
R16812 vdd.n2383 vdd.n2340 39.2114
R16813 vdd.n2387 vdd.n2341 39.2114
R16814 vdd.n2391 vdd.n2342 39.2114
R16815 vdd.n2395 vdd.n2343 39.2114
R16816 vdd.n2399 vdd.n2344 39.2114
R16817 vdd.n2403 vdd.n2345 39.2114
R16818 vdd.n2407 vdd.n2346 39.2114
R16819 vdd.n2411 vdd.n2347 39.2114
R16820 vdd.n2415 vdd.n2348 39.2114
R16821 vdd.n2571 vdd.n2570 39.2114
R16822 vdd.n2358 vdd.n2333 39.2114
R16823 vdd.n2362 vdd.n2334 39.2114
R16824 vdd.n2366 vdd.n2335 39.2114
R16825 vdd.n2370 vdd.n2336 39.2114
R16826 vdd.n2374 vdd.n2337 39.2114
R16827 vdd.n2378 vdd.n2338 39.2114
R16828 vdd.n2382 vdd.n2339 39.2114
R16829 vdd.n2386 vdd.n2340 39.2114
R16830 vdd.n2390 vdd.n2341 39.2114
R16831 vdd.n2394 vdd.n2342 39.2114
R16832 vdd.n2398 vdd.n2343 39.2114
R16833 vdd.n2402 vdd.n2344 39.2114
R16834 vdd.n2406 vdd.n2345 39.2114
R16835 vdd.n2410 vdd.n2346 39.2114
R16836 vdd.n2414 vdd.n2347 39.2114
R16837 vdd.n2417 vdd.n2348 39.2114
R16838 vdd.n629 vdd.n624 39.2114
R16839 vdd.n2779 vdd.n2778 39.2114
R16840 vdd.n623 vdd.n621 39.2114
R16841 vdd.n2786 vdd.n2785 39.2114
R16842 vdd.n620 vdd.n618 39.2114
R16843 vdd.n2793 vdd.n2792 39.2114
R16844 vdd.n617 vdd.n615 39.2114
R16845 vdd.n2800 vdd.n2799 39.2114
R16846 vdd.n2803 vdd.n2802 39.2114
R16847 vdd.n2659 vdd.n2658 39.2114
R16848 vdd.n2664 vdd.n2663 39.2114
R16849 vdd.n2657 vdd.n2655 39.2114
R16850 vdd.n2671 vdd.n2670 39.2114
R16851 vdd.n2654 vdd.n2652 39.2114
R16852 vdd.n2678 vdd.n2677 39.2114
R16853 vdd.n2651 vdd.n2649 39.2114
R16854 vdd.n2685 vdd.n2684 39.2114
R16855 vdd.n1823 vdd.n1822 39.2114
R16856 vdd.n1829 vdd.n1828 39.2114
R16857 vdd.n1830 vdd.n1819 39.2114
R16858 vdd.n1837 vdd.n1836 39.2114
R16859 vdd.n1838 vdd.n1817 39.2114
R16860 vdd.n1845 vdd.n1844 39.2114
R16861 vdd.n1846 vdd.n1815 39.2114
R16862 vdd.n1853 vdd.n1852 39.2114
R16863 vdd.n2024 vdd.n2023 39.2114
R16864 vdd.n2021 vdd.n2020 39.2114
R16865 vdd.n2016 vdd.n2015 39.2114
R16866 vdd.n2013 vdd.n2012 39.2114
R16867 vdd.n2008 vdd.n2007 39.2114
R16868 vdd.n2005 vdd.n2004 39.2114
R16869 vdd.n2000 vdd.n1999 39.2114
R16870 vdd.n1997 vdd.n1996 39.2114
R16871 vdd.n1992 vdd.n1991 39.2114
R16872 vdd.n2249 vdd.n765 39.2114
R16873 vdd.n2254 vdd.n766 39.2114
R16874 vdd.n2258 vdd.n767 39.2114
R16875 vdd.n2262 vdd.n768 39.2114
R16876 vdd.n2266 vdd.n769 39.2114
R16877 vdd.n2270 vdd.n770 39.2114
R16878 vdd.n2274 vdd.n771 39.2114
R16879 vdd.n2278 vdd.n772 39.2114
R16880 vdd.n2282 vdd.n773 39.2114
R16881 vdd.n2286 vdd.n774 39.2114
R16882 vdd.n2290 vdd.n775 39.2114
R16883 vdd.n2294 vdd.n776 39.2114
R16884 vdd.n2298 vdd.n777 39.2114
R16885 vdd.n2302 vdd.n778 39.2114
R16886 vdd.n2306 vdd.n779 39.2114
R16887 vdd.n2310 vdd.n780 39.2114
R16888 vdd.n783 vdd.n781 39.2114
R16889 vdd.n2568 vdd.n2567 39.2114
R16890 vdd.n2561 vdd.n2317 39.2114
R16891 vdd.n2557 vdd.n2318 39.2114
R16892 vdd.n2553 vdd.n2319 39.2114
R16893 vdd.n2549 vdd.n2320 39.2114
R16894 vdd.n2545 vdd.n2321 39.2114
R16895 vdd.n2541 vdd.n2322 39.2114
R16896 vdd.n2537 vdd.n2323 39.2114
R16897 vdd.n2533 vdd.n2324 39.2114
R16898 vdd.n2529 vdd.n2325 39.2114
R16899 vdd.n2525 vdd.n2326 39.2114
R16900 vdd.n2521 vdd.n2327 39.2114
R16901 vdd.n2517 vdd.n2328 39.2114
R16902 vdd.n2513 vdd.n2329 39.2114
R16903 vdd.n2509 vdd.n2330 39.2114
R16904 vdd.n2504 vdd.n2331 39.2114
R16905 vdd.n2500 vdd.n2332 39.2114
R16906 vdd.n2706 vdd.n660 39.2114
R16907 vdd.n2713 vdd.n2712 39.2114
R16908 vdd.n659 vdd.n657 39.2114
R16909 vdd.n2720 vdd.n2719 39.2114
R16910 vdd.n656 vdd.n654 39.2114
R16911 vdd.n2727 vdd.n2726 39.2114
R16912 vdd.n653 vdd.n651 39.2114
R16913 vdd.n2734 vdd.n2733 39.2114
R16914 vdd.n650 vdd.n648 39.2114
R16915 vdd.n2742 vdd.n2741 39.2114
R16916 vdd.n647 vdd.n645 39.2114
R16917 vdd.n2749 vdd.n2748 39.2114
R16918 vdd.n644 vdd.n642 39.2114
R16919 vdd.n2756 vdd.n2755 39.2114
R16920 vdd.n641 vdd.n639 39.2114
R16921 vdd.n2763 vdd.n2762 39.2114
R16922 vdd.n2766 vdd.n2765 39.2114
R16923 vdd.n791 vdd.n747 39.2114
R16924 vdd.n2238 vdd.n748 39.2114
R16925 vdd.n2234 vdd.n749 39.2114
R16926 vdd.n2230 vdd.n750 39.2114
R16927 vdd.n2226 vdd.n751 39.2114
R16928 vdd.n2222 vdd.n752 39.2114
R16929 vdd.n2218 vdd.n753 39.2114
R16930 vdd.n2214 vdd.n754 39.2114
R16931 vdd.n2210 vdd.n755 39.2114
R16932 vdd.n2206 vdd.n756 39.2114
R16933 vdd.n2202 vdd.n757 39.2114
R16934 vdd.n2198 vdd.n758 39.2114
R16935 vdd.n2194 vdd.n759 39.2114
R16936 vdd.n2190 vdd.n760 39.2114
R16937 vdd.n2186 vdd.n761 39.2114
R16938 vdd.n2182 vdd.n762 39.2114
R16939 vdd.n2178 vdd.n763 39.2114
R16940 vdd.n2081 vdd.n880 39.2114
R16941 vdd.n2080 vdd.n2079 39.2114
R16942 vdd.n2073 vdd.n882 39.2114
R16943 vdd.n2072 vdd.n2071 39.2114
R16944 vdd.n2065 vdd.n884 39.2114
R16945 vdd.n2064 vdd.n2063 39.2114
R16946 vdd.n2057 vdd.n886 39.2114
R16947 vdd.n2056 vdd.n2055 39.2114
R16948 vdd.n889 vdd.n888 39.2114
R16949 vdd.n1897 vdd.n1896 39.2114
R16950 vdd.n1902 vdd.n1901 39.2114
R16951 vdd.n1905 vdd.n1904 39.2114
R16952 vdd.n1910 vdd.n1909 39.2114
R16953 vdd.n1913 vdd.n1912 39.2114
R16954 vdd.n1918 vdd.n1917 39.2114
R16955 vdd.n1921 vdd.n1920 39.2114
R16956 vdd.n1927 vdd.n1926 39.2114
R16957 vdd.n2175 vdd.n763 39.2114
R16958 vdd.n2179 vdd.n762 39.2114
R16959 vdd.n2183 vdd.n761 39.2114
R16960 vdd.n2187 vdd.n760 39.2114
R16961 vdd.n2191 vdd.n759 39.2114
R16962 vdd.n2195 vdd.n758 39.2114
R16963 vdd.n2199 vdd.n757 39.2114
R16964 vdd.n2203 vdd.n756 39.2114
R16965 vdd.n2207 vdd.n755 39.2114
R16966 vdd.n2211 vdd.n754 39.2114
R16967 vdd.n2215 vdd.n753 39.2114
R16968 vdd.n2219 vdd.n752 39.2114
R16969 vdd.n2223 vdd.n751 39.2114
R16970 vdd.n2227 vdd.n750 39.2114
R16971 vdd.n2231 vdd.n749 39.2114
R16972 vdd.n2235 vdd.n748 39.2114
R16973 vdd.n2239 vdd.n747 39.2114
R16974 vdd.n2082 vdd.n2081 39.2114
R16975 vdd.n2079 vdd.n2078 39.2114
R16976 vdd.n2074 vdd.n2073 39.2114
R16977 vdd.n2071 vdd.n2070 39.2114
R16978 vdd.n2066 vdd.n2065 39.2114
R16979 vdd.n2063 vdd.n2062 39.2114
R16980 vdd.n2058 vdd.n2057 39.2114
R16981 vdd.n2055 vdd.n2054 39.2114
R16982 vdd.n890 vdd.n889 39.2114
R16983 vdd.n1898 vdd.n1897 39.2114
R16984 vdd.n1903 vdd.n1902 39.2114
R16985 vdd.n1904 vdd.n1894 39.2114
R16986 vdd.n1911 vdd.n1910 39.2114
R16987 vdd.n1912 vdd.n1892 39.2114
R16988 vdd.n1919 vdd.n1918 39.2114
R16989 vdd.n1920 vdd.n1888 39.2114
R16990 vdd.n1928 vdd.n1927 39.2114
R16991 vdd.n2047 vdd.n2046 37.2369
R16992 vdd.n1750 vdd.n1683 37.2369
R16993 vdd.n1789 vdd.n1643 37.2369
R16994 vdd.n2854 vdd.n581 37.2369
R16995 vdd.n545 vdd.n544 37.2369
R16996 vdd.n2810 vdd.n2809 37.2369
R16997 vdd.n2089 vdd.n875 31.6883
R16998 vdd.n2314 vdd.n784 31.6883
R16999 vdd.n2247 vdd.n787 31.6883
R17000 vdd.n1993 vdd.n1990 31.6883
R17001 vdd.n2501 vdd.n2499 31.6883
R17002 vdd.n2708 vdd.n2705 31.6883
R17003 vdd.n2578 vdd.n740 31.6883
R17004 vdd.n2769 vdd.n2768 31.6883
R17005 vdd.n2688 vdd.n2687 31.6883
R17006 vdd.n2774 vdd.n628 31.6883
R17007 vdd.n2420 vdd.n2419 31.6883
R17008 vdd.n2574 vdd.n2573 31.6883
R17009 vdd.n2085 vdd.n2084 31.6883
R17010 vdd.n2242 vdd.n2241 31.6883
R17011 vdd.n2174 vdd.n2173 31.6883
R17012 vdd.n1931 vdd.n1930 31.6883
R17013 vdd.n1924 vdd.n1890 30.449
R17014 vdd.n795 vdd.n794 30.449
R17015 vdd.n1865 vdd.n1864 30.449
R17016 vdd.n2252 vdd.n786 30.449
R17017 vdd.n2356 vdd.n2355 30.449
R17018 vdd.n663 vdd.n662 30.449
R17019 vdd.n2506 vdd.n2352 30.449
R17020 vdd.n627 vdd.n626 30.449
R17021 vdd.n1215 vdd.n982 20.633
R17022 vdd.n2041 vdd.n901 20.633
R17023 vdd.n2940 vdd.n516 20.633
R17024 vdd.n3138 vdd.n351 20.633
R17025 vdd.n1217 vdd.n979 19.3944
R17026 vdd.n1221 vdd.n979 19.3944
R17027 vdd.n1221 vdd.n970 19.3944
R17028 vdd.n1233 vdd.n970 19.3944
R17029 vdd.n1233 vdd.n968 19.3944
R17030 vdd.n1237 vdd.n968 19.3944
R17031 vdd.n1237 vdd.n957 19.3944
R17032 vdd.n1249 vdd.n957 19.3944
R17033 vdd.n1249 vdd.n955 19.3944
R17034 vdd.n1253 vdd.n955 19.3944
R17035 vdd.n1253 vdd.n946 19.3944
R17036 vdd.n1266 vdd.n946 19.3944
R17037 vdd.n1266 vdd.n944 19.3944
R17038 vdd.n1270 vdd.n944 19.3944
R17039 vdd.n1270 vdd.n935 19.3944
R17040 vdd.n1564 vdd.n935 19.3944
R17041 vdd.n1564 vdd.n933 19.3944
R17042 vdd.n1568 vdd.n933 19.3944
R17043 vdd.n1568 vdd.n923 19.3944
R17044 vdd.n1581 vdd.n923 19.3944
R17045 vdd.n1581 vdd.n921 19.3944
R17046 vdd.n1585 vdd.n921 19.3944
R17047 vdd.n1585 vdd.n913 19.3944
R17048 vdd.n1598 vdd.n913 19.3944
R17049 vdd.n1598 vdd.n910 19.3944
R17050 vdd.n1604 vdd.n910 19.3944
R17051 vdd.n1604 vdd.n911 19.3944
R17052 vdd.n911 vdd.n900 19.3944
R17053 vdd.n1142 vdd.n1068 19.3944
R17054 vdd.n1142 vdd.n1070 19.3944
R17055 vdd.n1138 vdd.n1070 19.3944
R17056 vdd.n1138 vdd.n1137 19.3944
R17057 vdd.n1137 vdd.n1136 19.3944
R17058 vdd.n1136 vdd.n1078 19.3944
R17059 vdd.n1132 vdd.n1078 19.3944
R17060 vdd.n1132 vdd.n1131 19.3944
R17061 vdd.n1131 vdd.n1130 19.3944
R17062 vdd.n1130 vdd.n1086 19.3944
R17063 vdd.n1126 vdd.n1086 19.3944
R17064 vdd.n1126 vdd.n1125 19.3944
R17065 vdd.n1125 vdd.n1124 19.3944
R17066 vdd.n1124 vdd.n1094 19.3944
R17067 vdd.n1120 vdd.n1094 19.3944
R17068 vdd.n1120 vdd.n1119 19.3944
R17069 vdd.n1119 vdd.n1118 19.3944
R17070 vdd.n1118 vdd.n1102 19.3944
R17071 vdd.n1114 vdd.n1102 19.3944
R17072 vdd.n1114 vdd.n1113 19.3944
R17073 vdd.n1180 vdd.n1179 19.3944
R17074 vdd.n1179 vdd.n1178 19.3944
R17075 vdd.n1178 vdd.n1031 19.3944
R17076 vdd.n1174 vdd.n1031 19.3944
R17077 vdd.n1174 vdd.n1173 19.3944
R17078 vdd.n1173 vdd.n1172 19.3944
R17079 vdd.n1172 vdd.n1039 19.3944
R17080 vdd.n1168 vdd.n1039 19.3944
R17081 vdd.n1168 vdd.n1167 19.3944
R17082 vdd.n1167 vdd.n1166 19.3944
R17083 vdd.n1166 vdd.n1047 19.3944
R17084 vdd.n1162 vdd.n1047 19.3944
R17085 vdd.n1162 vdd.n1161 19.3944
R17086 vdd.n1161 vdd.n1160 19.3944
R17087 vdd.n1160 vdd.n1055 19.3944
R17088 vdd.n1156 vdd.n1055 19.3944
R17089 vdd.n1156 vdd.n1155 19.3944
R17090 vdd.n1155 vdd.n1154 19.3944
R17091 vdd.n1154 vdd.n1063 19.3944
R17092 vdd.n1150 vdd.n1063 19.3944
R17093 vdd.n1210 vdd.n1209 19.3944
R17094 vdd.n1209 vdd.n1208 19.3944
R17095 vdd.n1208 vdd.n989 19.3944
R17096 vdd.n1204 vdd.n989 19.3944
R17097 vdd.n1204 vdd.n1203 19.3944
R17098 vdd.n1203 vdd.n1202 19.3944
R17099 vdd.n1202 vdd.n997 19.3944
R17100 vdd.n1198 vdd.n997 19.3944
R17101 vdd.n1198 vdd.n1197 19.3944
R17102 vdd.n1197 vdd.n1196 19.3944
R17103 vdd.n1196 vdd.n1005 19.3944
R17104 vdd.n1192 vdd.n1005 19.3944
R17105 vdd.n1192 vdd.n1191 19.3944
R17106 vdd.n1191 vdd.n1190 19.3944
R17107 vdd.n1190 vdd.n1013 19.3944
R17108 vdd.n1186 vdd.n1013 19.3944
R17109 vdd.n1186 vdd.n1185 19.3944
R17110 vdd.n1185 vdd.n1184 19.3944
R17111 vdd.n1746 vdd.n1681 19.3944
R17112 vdd.n1746 vdd.n1687 19.3944
R17113 vdd.n1741 vdd.n1687 19.3944
R17114 vdd.n1741 vdd.n1740 19.3944
R17115 vdd.n1740 vdd.n1739 19.3944
R17116 vdd.n1739 vdd.n1694 19.3944
R17117 vdd.n1734 vdd.n1694 19.3944
R17118 vdd.n1734 vdd.n1733 19.3944
R17119 vdd.n1733 vdd.n1732 19.3944
R17120 vdd.n1732 vdd.n1701 19.3944
R17121 vdd.n1727 vdd.n1701 19.3944
R17122 vdd.n1727 vdd.n1726 19.3944
R17123 vdd.n1726 vdd.n1725 19.3944
R17124 vdd.n1725 vdd.n1709 19.3944
R17125 vdd.n1720 vdd.n1709 19.3944
R17126 vdd.n1720 vdd.n1719 19.3944
R17127 vdd.n1715 vdd.n1714 19.3944
R17128 vdd.n2048 vdd.n896 19.3944
R17129 vdd.n1785 vdd.n1641 19.3944
R17130 vdd.n1785 vdd.n1647 19.3944
R17131 vdd.n1780 vdd.n1647 19.3944
R17132 vdd.n1780 vdd.n1779 19.3944
R17133 vdd.n1779 vdd.n1778 19.3944
R17134 vdd.n1778 vdd.n1654 19.3944
R17135 vdd.n1773 vdd.n1654 19.3944
R17136 vdd.n1773 vdd.n1772 19.3944
R17137 vdd.n1772 vdd.n1771 19.3944
R17138 vdd.n1771 vdd.n1661 19.3944
R17139 vdd.n1766 vdd.n1661 19.3944
R17140 vdd.n1766 vdd.n1765 19.3944
R17141 vdd.n1765 vdd.n1764 19.3944
R17142 vdd.n1764 vdd.n1668 19.3944
R17143 vdd.n1759 vdd.n1668 19.3944
R17144 vdd.n1759 vdd.n1758 19.3944
R17145 vdd.n1758 vdd.n1757 19.3944
R17146 vdd.n1757 vdd.n1675 19.3944
R17147 vdd.n1752 vdd.n1675 19.3944
R17148 vdd.n1752 vdd.n1751 19.3944
R17149 vdd.n2036 vdd.n2035 19.3944
R17150 vdd.n2035 vdd.n1613 19.3944
R17151 vdd.n2030 vdd.n2029 19.3944
R17152 vdd.n1812 vdd.n1617 19.3944
R17153 vdd.n1812 vdd.n1619 19.3944
R17154 vdd.n1622 vdd.n1619 19.3944
R17155 vdd.n1805 vdd.n1622 19.3944
R17156 vdd.n1805 vdd.n1804 19.3944
R17157 vdd.n1804 vdd.n1803 19.3944
R17158 vdd.n1803 vdd.n1628 19.3944
R17159 vdd.n1798 vdd.n1628 19.3944
R17160 vdd.n1798 vdd.n1797 19.3944
R17161 vdd.n1797 vdd.n1796 19.3944
R17162 vdd.n1796 vdd.n1635 19.3944
R17163 vdd.n1791 vdd.n1635 19.3944
R17164 vdd.n1791 vdd.n1790 19.3944
R17165 vdd.n1213 vdd.n976 19.3944
R17166 vdd.n1225 vdd.n976 19.3944
R17167 vdd.n1225 vdd.n974 19.3944
R17168 vdd.n1229 vdd.n974 19.3944
R17169 vdd.n1229 vdd.n964 19.3944
R17170 vdd.n1241 vdd.n964 19.3944
R17171 vdd.n1241 vdd.n962 19.3944
R17172 vdd.n1245 vdd.n962 19.3944
R17173 vdd.n1245 vdd.n952 19.3944
R17174 vdd.n1258 vdd.n952 19.3944
R17175 vdd.n1258 vdd.n950 19.3944
R17176 vdd.n1262 vdd.n950 19.3944
R17177 vdd.n1262 vdd.n941 19.3944
R17178 vdd.n1274 vdd.n941 19.3944
R17179 vdd.n1274 vdd.n939 19.3944
R17180 vdd.n1560 vdd.n939 19.3944
R17181 vdd.n1560 vdd.n929 19.3944
R17182 vdd.n1573 vdd.n929 19.3944
R17183 vdd.n1573 vdd.n927 19.3944
R17184 vdd.n1577 vdd.n927 19.3944
R17185 vdd.n1577 vdd.n918 19.3944
R17186 vdd.n1590 vdd.n918 19.3944
R17187 vdd.n1590 vdd.n916 19.3944
R17188 vdd.n1594 vdd.n916 19.3944
R17189 vdd.n1594 vdd.n906 19.3944
R17190 vdd.n1609 vdd.n906 19.3944
R17191 vdd.n1609 vdd.n904 19.3944
R17192 vdd.n2039 vdd.n904 19.3944
R17193 vdd.n2942 vdd.n513 19.3944
R17194 vdd.n2946 vdd.n513 19.3944
R17195 vdd.n2946 vdd.n503 19.3944
R17196 vdd.n2958 vdd.n503 19.3944
R17197 vdd.n2958 vdd.n501 19.3944
R17198 vdd.n2962 vdd.n501 19.3944
R17199 vdd.n2962 vdd.n490 19.3944
R17200 vdd.n2974 vdd.n490 19.3944
R17201 vdd.n2974 vdd.n488 19.3944
R17202 vdd.n2978 vdd.n488 19.3944
R17203 vdd.n2978 vdd.n478 19.3944
R17204 vdd.n2991 vdd.n478 19.3944
R17205 vdd.n2991 vdd.n476 19.3944
R17206 vdd.n2995 vdd.n476 19.3944
R17207 vdd.n2996 vdd.n2995 19.3944
R17208 vdd.n2997 vdd.n2996 19.3944
R17209 vdd.n2997 vdd.n474 19.3944
R17210 vdd.n3001 vdd.n474 19.3944
R17211 vdd.n3002 vdd.n3001 19.3944
R17212 vdd.n3003 vdd.n3002 19.3944
R17213 vdd.n3003 vdd.n471 19.3944
R17214 vdd.n3007 vdd.n471 19.3944
R17215 vdd.n3008 vdd.n3007 19.3944
R17216 vdd.n3009 vdd.n3008 19.3944
R17217 vdd.n3009 vdd.n468 19.3944
R17218 vdd.n3013 vdd.n468 19.3944
R17219 vdd.n3014 vdd.n3013 19.3944
R17220 vdd.n3015 vdd.n3014 19.3944
R17221 vdd.n3058 vdd.n426 19.3944
R17222 vdd.n3058 vdd.n432 19.3944
R17223 vdd.n3053 vdd.n432 19.3944
R17224 vdd.n3053 vdd.n3052 19.3944
R17225 vdd.n3052 vdd.n3051 19.3944
R17226 vdd.n3051 vdd.n439 19.3944
R17227 vdd.n3046 vdd.n439 19.3944
R17228 vdd.n3046 vdd.n3045 19.3944
R17229 vdd.n3045 vdd.n3044 19.3944
R17230 vdd.n3044 vdd.n446 19.3944
R17231 vdd.n3039 vdd.n446 19.3944
R17232 vdd.n3039 vdd.n3038 19.3944
R17233 vdd.n3038 vdd.n3037 19.3944
R17234 vdd.n3037 vdd.n453 19.3944
R17235 vdd.n3032 vdd.n453 19.3944
R17236 vdd.n3032 vdd.n3031 19.3944
R17237 vdd.n3031 vdd.n3030 19.3944
R17238 vdd.n3030 vdd.n460 19.3944
R17239 vdd.n3025 vdd.n460 19.3944
R17240 vdd.n3025 vdd.n3024 19.3944
R17241 vdd.n3097 vdd.n386 19.3944
R17242 vdd.n3097 vdd.n392 19.3944
R17243 vdd.n3092 vdd.n392 19.3944
R17244 vdd.n3092 vdd.n3091 19.3944
R17245 vdd.n3091 vdd.n3090 19.3944
R17246 vdd.n3090 vdd.n399 19.3944
R17247 vdd.n3085 vdd.n399 19.3944
R17248 vdd.n3085 vdd.n3084 19.3944
R17249 vdd.n3084 vdd.n3083 19.3944
R17250 vdd.n3083 vdd.n406 19.3944
R17251 vdd.n3078 vdd.n406 19.3944
R17252 vdd.n3078 vdd.n3077 19.3944
R17253 vdd.n3077 vdd.n3076 19.3944
R17254 vdd.n3076 vdd.n413 19.3944
R17255 vdd.n3071 vdd.n413 19.3944
R17256 vdd.n3071 vdd.n3070 19.3944
R17257 vdd.n3070 vdd.n3069 19.3944
R17258 vdd.n3069 vdd.n420 19.3944
R17259 vdd.n3064 vdd.n420 19.3944
R17260 vdd.n3064 vdd.n3063 19.3944
R17261 vdd.n3133 vdd.n3132 19.3944
R17262 vdd.n3132 vdd.n3131 19.3944
R17263 vdd.n3131 vdd.n358 19.3944
R17264 vdd.n359 vdd.n358 19.3944
R17265 vdd.n3124 vdd.n359 19.3944
R17266 vdd.n3124 vdd.n3123 19.3944
R17267 vdd.n3123 vdd.n3122 19.3944
R17268 vdd.n3122 vdd.n366 19.3944
R17269 vdd.n3117 vdd.n366 19.3944
R17270 vdd.n3117 vdd.n3116 19.3944
R17271 vdd.n3116 vdd.n3115 19.3944
R17272 vdd.n3115 vdd.n373 19.3944
R17273 vdd.n3110 vdd.n373 19.3944
R17274 vdd.n3110 vdd.n3109 19.3944
R17275 vdd.n3109 vdd.n3108 19.3944
R17276 vdd.n3108 vdd.n380 19.3944
R17277 vdd.n3103 vdd.n380 19.3944
R17278 vdd.n3103 vdd.n3102 19.3944
R17279 vdd.n2938 vdd.n509 19.3944
R17280 vdd.n2950 vdd.n509 19.3944
R17281 vdd.n2950 vdd.n507 19.3944
R17282 vdd.n2954 vdd.n507 19.3944
R17283 vdd.n2954 vdd.n497 19.3944
R17284 vdd.n2966 vdd.n497 19.3944
R17285 vdd.n2966 vdd.n495 19.3944
R17286 vdd.n2970 vdd.n495 19.3944
R17287 vdd.n2970 vdd.n485 19.3944
R17288 vdd.n2983 vdd.n485 19.3944
R17289 vdd.n2983 vdd.n483 19.3944
R17290 vdd.n2987 vdd.n483 19.3944
R17291 vdd.n2987 vdd.n312 19.3944
R17292 vdd.n3166 vdd.n312 19.3944
R17293 vdd.n3166 vdd.n313 19.3944
R17294 vdd.n3160 vdd.n313 19.3944
R17295 vdd.n3160 vdd.n3159 19.3944
R17296 vdd.n3159 vdd.n3158 19.3944
R17297 vdd.n3158 vdd.n323 19.3944
R17298 vdd.n3152 vdd.n323 19.3944
R17299 vdd.n3152 vdd.n3151 19.3944
R17300 vdd.n3151 vdd.n3150 19.3944
R17301 vdd.n3150 vdd.n335 19.3944
R17302 vdd.n3144 vdd.n335 19.3944
R17303 vdd.n3144 vdd.n3143 19.3944
R17304 vdd.n3143 vdd.n3142 19.3944
R17305 vdd.n3142 vdd.n346 19.3944
R17306 vdd.n3136 vdd.n346 19.3944
R17307 vdd.n2895 vdd.n2894 19.3944
R17308 vdd.n2894 vdd.n2893 19.3944
R17309 vdd.n2893 vdd.n551 19.3944
R17310 vdd.n2887 vdd.n551 19.3944
R17311 vdd.n2887 vdd.n2886 19.3944
R17312 vdd.n2886 vdd.n2885 19.3944
R17313 vdd.n2885 vdd.n557 19.3944
R17314 vdd.n2879 vdd.n557 19.3944
R17315 vdd.n2879 vdd.n2878 19.3944
R17316 vdd.n2878 vdd.n2877 19.3944
R17317 vdd.n2877 vdd.n563 19.3944
R17318 vdd.n2871 vdd.n563 19.3944
R17319 vdd.n2871 vdd.n2870 19.3944
R17320 vdd.n2870 vdd.n2869 19.3944
R17321 vdd.n2869 vdd.n569 19.3944
R17322 vdd.n2863 vdd.n569 19.3944
R17323 vdd.n2863 vdd.n2862 19.3944
R17324 vdd.n2862 vdd.n2861 19.3944
R17325 vdd.n2861 vdd.n575 19.3944
R17326 vdd.n2855 vdd.n575 19.3944
R17327 vdd.n2935 vdd.n2934 19.3944
R17328 vdd.n2934 vdd.n519 19.3944
R17329 vdd.n2929 vdd.n2928 19.3944
R17330 vdd.n2925 vdd.n2924 19.3944
R17331 vdd.n2924 vdd.n525 19.3944
R17332 vdd.n2919 vdd.n525 19.3944
R17333 vdd.n2919 vdd.n2918 19.3944
R17334 vdd.n2918 vdd.n2917 19.3944
R17335 vdd.n2917 vdd.n531 19.3944
R17336 vdd.n2911 vdd.n531 19.3944
R17337 vdd.n2911 vdd.n2910 19.3944
R17338 vdd.n2910 vdd.n2909 19.3944
R17339 vdd.n2909 vdd.n537 19.3944
R17340 vdd.n2903 vdd.n537 19.3944
R17341 vdd.n2903 vdd.n2902 19.3944
R17342 vdd.n2902 vdd.n2901 19.3944
R17343 vdd.n2850 vdd.n579 19.3944
R17344 vdd.n2850 vdd.n583 19.3944
R17345 vdd.n2845 vdd.n583 19.3944
R17346 vdd.n2845 vdd.n2844 19.3944
R17347 vdd.n2844 vdd.n589 19.3944
R17348 vdd.n2839 vdd.n589 19.3944
R17349 vdd.n2839 vdd.n2838 19.3944
R17350 vdd.n2838 vdd.n2837 19.3944
R17351 vdd.n2837 vdd.n595 19.3944
R17352 vdd.n2831 vdd.n595 19.3944
R17353 vdd.n2831 vdd.n2830 19.3944
R17354 vdd.n2830 vdd.n2829 19.3944
R17355 vdd.n2829 vdd.n601 19.3944
R17356 vdd.n2823 vdd.n601 19.3944
R17357 vdd.n2823 vdd.n2822 19.3944
R17358 vdd.n2822 vdd.n2821 19.3944
R17359 vdd.n2817 vdd.n2816 19.3944
R17360 vdd.n2813 vdd.n2812 19.3944
R17361 vdd.n1149 vdd.n1068 19.0066
R17362 vdd.n1750 vdd.n1681 19.0066
R17363 vdd.n3062 vdd.n426 19.0066
R17364 vdd.n2854 vdd.n579 19.0066
R17365 vdd.n1890 vdd.n1889 16.0975
R17366 vdd.n794 vdd.n793 16.0975
R17367 vdd.n1111 vdd.n1110 16.0975
R17368 vdd.n1148 vdd.n1147 16.0975
R17369 vdd.n1022 vdd.n1021 16.0975
R17370 vdd.n2046 vdd.n2045 16.0975
R17371 vdd.n1683 vdd.n1682 16.0975
R17372 vdd.n1643 vdd.n1642 16.0975
R17373 vdd.n1864 vdd.n1863 16.0975
R17374 vdd.n786 vdd.n785 16.0975
R17375 vdd.n2355 vdd.n2354 16.0975
R17376 vdd.n3022 vdd.n3021 16.0975
R17377 vdd.n428 vdd.n427 16.0975
R17378 vdd.n388 vdd.n387 16.0975
R17379 vdd.n581 vdd.n580 16.0975
R17380 vdd.n544 vdd.n543 16.0975
R17381 vdd.n662 vdd.n661 16.0975
R17382 vdd.n2352 vdd.n2351 16.0975
R17383 vdd.n2809 vdd.n2808 16.0975
R17384 vdd.n626 vdd.n625 16.0975
R17385 vdd.t176 vdd.n2316 15.4182
R17386 vdd.n2569 vdd.t77 15.4182
R17387 vdd.n28 vdd.n27 14.5238
R17388 vdd.n2087 vdd.n877 14.5112
R17389 vdd.n2771 vdd.n613 14.5112
R17390 vdd.n304 vdd.n269 13.1884
R17391 vdd.n253 vdd.n218 13.1884
R17392 vdd.n210 vdd.n175 13.1884
R17393 vdd.n159 vdd.n124 13.1884
R17394 vdd.n117 vdd.n82 13.1884
R17395 vdd.n66 vdd.n31 13.1884
R17396 vdd.n1499 vdd.n1464 13.1884
R17397 vdd.n1550 vdd.n1515 13.1884
R17398 vdd.n1405 vdd.n1370 13.1884
R17399 vdd.n1456 vdd.n1421 13.1884
R17400 vdd.n1312 vdd.n1277 13.1884
R17401 vdd.n1363 vdd.n1328 13.1884
R17402 vdd.n1180 vdd.n1023 12.9944
R17403 vdd.n1184 vdd.n1023 12.9944
R17404 vdd.n1789 vdd.n1641 12.9944
R17405 vdd.n1790 vdd.n1789 12.9944
R17406 vdd.n3101 vdd.n386 12.9944
R17407 vdd.n3102 vdd.n3101 12.9944
R17408 vdd.n2895 vdd.n545 12.9944
R17409 vdd.n2901 vdd.n545 12.9944
R17410 vdd.n305 vdd.n267 12.8005
R17411 vdd.n300 vdd.n271 12.8005
R17412 vdd.n254 vdd.n216 12.8005
R17413 vdd.n249 vdd.n220 12.8005
R17414 vdd.n211 vdd.n173 12.8005
R17415 vdd.n206 vdd.n177 12.8005
R17416 vdd.n160 vdd.n122 12.8005
R17417 vdd.n155 vdd.n126 12.8005
R17418 vdd.n118 vdd.n80 12.8005
R17419 vdd.n113 vdd.n84 12.8005
R17420 vdd.n67 vdd.n29 12.8005
R17421 vdd.n62 vdd.n33 12.8005
R17422 vdd.n1500 vdd.n1462 12.8005
R17423 vdd.n1495 vdd.n1466 12.8005
R17424 vdd.n1551 vdd.n1513 12.8005
R17425 vdd.n1546 vdd.n1517 12.8005
R17426 vdd.n1406 vdd.n1368 12.8005
R17427 vdd.n1401 vdd.n1372 12.8005
R17428 vdd.n1457 vdd.n1419 12.8005
R17429 vdd.n1452 vdd.n1423 12.8005
R17430 vdd.n1313 vdd.n1275 12.8005
R17431 vdd.n1308 vdd.n1279 12.8005
R17432 vdd.n1364 vdd.n1326 12.8005
R17433 vdd.n1359 vdd.n1330 12.8005
R17434 vdd.n299 vdd.n272 12.0247
R17435 vdd.n248 vdd.n221 12.0247
R17436 vdd.n205 vdd.n178 12.0247
R17437 vdd.n154 vdd.n127 12.0247
R17438 vdd.n112 vdd.n85 12.0247
R17439 vdd.n61 vdd.n34 12.0247
R17440 vdd.n1494 vdd.n1467 12.0247
R17441 vdd.n1545 vdd.n1518 12.0247
R17442 vdd.n1400 vdd.n1373 12.0247
R17443 vdd.n1451 vdd.n1424 12.0247
R17444 vdd.n1307 vdd.n1280 12.0247
R17445 vdd.n1358 vdd.n1331 12.0247
R17446 vdd.n1215 vdd.n983 11.337
R17447 vdd.n1223 vdd.n972 11.337
R17448 vdd.n1231 vdd.n972 11.337
R17449 vdd.n1239 vdd.n966 11.337
R17450 vdd.n1247 vdd.n959 11.337
R17451 vdd.n1256 vdd.n1255 11.337
R17452 vdd.n1264 vdd.n948 11.337
R17453 vdd.n1562 vdd.n937 11.337
R17454 vdd.n1571 vdd.n931 11.337
R17455 vdd.n1579 vdd.n925 11.337
R17456 vdd.n1588 vdd.n1587 11.337
R17457 vdd.n1596 vdd.n908 11.337
R17458 vdd.n1607 vdd.n908 11.337
R17459 vdd.n1607 vdd.n1606 11.337
R17460 vdd.n2948 vdd.n511 11.337
R17461 vdd.n2948 vdd.n505 11.337
R17462 vdd.n2956 vdd.n505 11.337
R17463 vdd.n2964 vdd.n499 11.337
R17464 vdd.n2972 vdd.n492 11.337
R17465 vdd.n2981 vdd.n2980 11.337
R17466 vdd.n2989 vdd.n481 11.337
R17467 vdd.n3163 vdd.n3162 11.337
R17468 vdd.n3156 vdd.n325 11.337
R17469 vdd.n3154 vdd.n329 11.337
R17470 vdd.n3148 vdd.n3147 11.337
R17471 vdd.n3146 vdd.n340 11.337
R17472 vdd.n3140 vdd.n340 11.337
R17473 vdd.n3139 vdd.n3138 11.337
R17474 vdd.n296 vdd.n295 11.249
R17475 vdd.n245 vdd.n244 11.249
R17476 vdd.n202 vdd.n201 11.249
R17477 vdd.n151 vdd.n150 11.249
R17478 vdd.n109 vdd.n108 11.249
R17479 vdd.n58 vdd.n57 11.249
R17480 vdd.n1491 vdd.n1490 11.249
R17481 vdd.n1542 vdd.n1541 11.249
R17482 vdd.n1397 vdd.n1396 11.249
R17483 vdd.n1448 vdd.n1447 11.249
R17484 vdd.n1304 vdd.n1303 11.249
R17485 vdd.n1355 vdd.n1354 11.249
R17486 vdd.n2244 vdd.t17 11.1103
R17487 vdd.n2576 vdd.t211 11.1103
R17488 vdd.n1231 vdd.t186 10.9969
R17489 vdd.t4 vdd.n3146 10.9969
R17490 vdd.n960 vdd.t66 10.7702
R17491 vdd.t24 vdd.n3155 10.7702
R17492 vdd.n281 vdd.n280 10.7238
R17493 vdd.n230 vdd.n229 10.7238
R17494 vdd.n187 vdd.n186 10.7238
R17495 vdd.n136 vdd.n135 10.7238
R17496 vdd.n94 vdd.n93 10.7238
R17497 vdd.n43 vdd.n42 10.7238
R17498 vdd.n1476 vdd.n1475 10.7238
R17499 vdd.n1527 vdd.n1526 10.7238
R17500 vdd.n1382 vdd.n1381 10.7238
R17501 vdd.n1433 vdd.n1432 10.7238
R17502 vdd.n1289 vdd.n1288 10.7238
R17503 vdd.n1340 vdd.n1339 10.7238
R17504 vdd.n2090 vdd.n2089 10.6151
R17505 vdd.n2091 vdd.n2090 10.6151
R17506 vdd.n2091 vdd.n863 10.6151
R17507 vdd.n2101 vdd.n863 10.6151
R17508 vdd.n2102 vdd.n2101 10.6151
R17509 vdd.n2103 vdd.n2102 10.6151
R17510 vdd.n2103 vdd.n850 10.6151
R17511 vdd.n2114 vdd.n850 10.6151
R17512 vdd.n2115 vdd.n2114 10.6151
R17513 vdd.n2116 vdd.n2115 10.6151
R17514 vdd.n2116 vdd.n838 10.6151
R17515 vdd.n2126 vdd.n838 10.6151
R17516 vdd.n2127 vdd.n2126 10.6151
R17517 vdd.n2128 vdd.n2127 10.6151
R17518 vdd.n2128 vdd.n826 10.6151
R17519 vdd.n2138 vdd.n826 10.6151
R17520 vdd.n2139 vdd.n2138 10.6151
R17521 vdd.n2140 vdd.n2139 10.6151
R17522 vdd.n2140 vdd.n815 10.6151
R17523 vdd.n2150 vdd.n815 10.6151
R17524 vdd.n2151 vdd.n2150 10.6151
R17525 vdd.n2152 vdd.n2151 10.6151
R17526 vdd.n2152 vdd.n802 10.6151
R17527 vdd.n2164 vdd.n802 10.6151
R17528 vdd.n2165 vdd.n2164 10.6151
R17529 vdd.n2167 vdd.n2165 10.6151
R17530 vdd.n2167 vdd.n2166 10.6151
R17531 vdd.n2166 vdd.n784 10.6151
R17532 vdd.n2314 vdd.n2313 10.6151
R17533 vdd.n2313 vdd.n2312 10.6151
R17534 vdd.n2312 vdd.n2309 10.6151
R17535 vdd.n2309 vdd.n2308 10.6151
R17536 vdd.n2308 vdd.n2305 10.6151
R17537 vdd.n2305 vdd.n2304 10.6151
R17538 vdd.n2304 vdd.n2301 10.6151
R17539 vdd.n2301 vdd.n2300 10.6151
R17540 vdd.n2300 vdd.n2297 10.6151
R17541 vdd.n2297 vdd.n2296 10.6151
R17542 vdd.n2296 vdd.n2293 10.6151
R17543 vdd.n2293 vdd.n2292 10.6151
R17544 vdd.n2292 vdd.n2289 10.6151
R17545 vdd.n2289 vdd.n2288 10.6151
R17546 vdd.n2288 vdd.n2285 10.6151
R17547 vdd.n2285 vdd.n2284 10.6151
R17548 vdd.n2284 vdd.n2281 10.6151
R17549 vdd.n2281 vdd.n2280 10.6151
R17550 vdd.n2280 vdd.n2277 10.6151
R17551 vdd.n2277 vdd.n2276 10.6151
R17552 vdd.n2276 vdd.n2273 10.6151
R17553 vdd.n2273 vdd.n2272 10.6151
R17554 vdd.n2272 vdd.n2269 10.6151
R17555 vdd.n2269 vdd.n2268 10.6151
R17556 vdd.n2268 vdd.n2265 10.6151
R17557 vdd.n2265 vdd.n2264 10.6151
R17558 vdd.n2264 vdd.n2261 10.6151
R17559 vdd.n2261 vdd.n2260 10.6151
R17560 vdd.n2260 vdd.n2257 10.6151
R17561 vdd.n2257 vdd.n2256 10.6151
R17562 vdd.n2256 vdd.n2253 10.6151
R17563 vdd.n2251 vdd.n2248 10.6151
R17564 vdd.n2248 vdd.n2247 10.6151
R17565 vdd.n1990 vdd.n1989 10.6151
R17566 vdd.n1989 vdd.n1987 10.6151
R17567 vdd.n1987 vdd.n1986 10.6151
R17568 vdd.n1986 vdd.n1984 10.6151
R17569 vdd.n1984 vdd.n1983 10.6151
R17570 vdd.n1983 vdd.n1981 10.6151
R17571 vdd.n1981 vdd.n1980 10.6151
R17572 vdd.n1980 vdd.n1978 10.6151
R17573 vdd.n1978 vdd.n1977 10.6151
R17574 vdd.n1977 vdd.n1975 10.6151
R17575 vdd.n1975 vdd.n1974 10.6151
R17576 vdd.n1974 vdd.n1972 10.6151
R17577 vdd.n1972 vdd.n1971 10.6151
R17578 vdd.n1971 vdd.n1886 10.6151
R17579 vdd.n1886 vdd.n1885 10.6151
R17580 vdd.n1885 vdd.n1883 10.6151
R17581 vdd.n1883 vdd.n1882 10.6151
R17582 vdd.n1882 vdd.n1880 10.6151
R17583 vdd.n1880 vdd.n1879 10.6151
R17584 vdd.n1879 vdd.n1877 10.6151
R17585 vdd.n1877 vdd.n1876 10.6151
R17586 vdd.n1876 vdd.n1874 10.6151
R17587 vdd.n1874 vdd.n1873 10.6151
R17588 vdd.n1873 vdd.n1871 10.6151
R17589 vdd.n1871 vdd.n1870 10.6151
R17590 vdd.n1870 vdd.n1867 10.6151
R17591 vdd.n1867 vdd.n1866 10.6151
R17592 vdd.n1866 vdd.n787 10.6151
R17593 vdd.n1824 vdd.n875 10.6151
R17594 vdd.n1825 vdd.n1824 10.6151
R17595 vdd.n1826 vdd.n1825 10.6151
R17596 vdd.n1826 vdd.n1820 10.6151
R17597 vdd.n1832 vdd.n1820 10.6151
R17598 vdd.n1833 vdd.n1832 10.6151
R17599 vdd.n1834 vdd.n1833 10.6151
R17600 vdd.n1834 vdd.n1818 10.6151
R17601 vdd.n1840 vdd.n1818 10.6151
R17602 vdd.n1841 vdd.n1840 10.6151
R17603 vdd.n1842 vdd.n1841 10.6151
R17604 vdd.n1842 vdd.n1816 10.6151
R17605 vdd.n1848 vdd.n1816 10.6151
R17606 vdd.n1849 vdd.n1848 10.6151
R17607 vdd.n1850 vdd.n1849 10.6151
R17608 vdd.n1850 vdd.n1814 10.6151
R17609 vdd.n2026 vdd.n1814 10.6151
R17610 vdd.n2026 vdd.n2025 10.6151
R17611 vdd.n2025 vdd.n1855 10.6151
R17612 vdd.n2019 vdd.n1855 10.6151
R17613 vdd.n2019 vdd.n2018 10.6151
R17614 vdd.n2018 vdd.n2017 10.6151
R17615 vdd.n2017 vdd.n1857 10.6151
R17616 vdd.n2011 vdd.n1857 10.6151
R17617 vdd.n2011 vdd.n2010 10.6151
R17618 vdd.n2010 vdd.n2009 10.6151
R17619 vdd.n2009 vdd.n1859 10.6151
R17620 vdd.n2003 vdd.n1859 10.6151
R17621 vdd.n2003 vdd.n2002 10.6151
R17622 vdd.n2002 vdd.n2001 10.6151
R17623 vdd.n2001 vdd.n1861 10.6151
R17624 vdd.n1995 vdd.n1994 10.6151
R17625 vdd.n1994 vdd.n1993 10.6151
R17626 vdd.n2499 vdd.n2498 10.6151
R17627 vdd.n2498 vdd.n2496 10.6151
R17628 vdd.n2496 vdd.n2495 10.6151
R17629 vdd.n2495 vdd.n2353 10.6151
R17630 vdd.n2442 vdd.n2353 10.6151
R17631 vdd.n2443 vdd.n2442 10.6151
R17632 vdd.n2445 vdd.n2443 10.6151
R17633 vdd.n2446 vdd.n2445 10.6151
R17634 vdd.n2448 vdd.n2446 10.6151
R17635 vdd.n2449 vdd.n2448 10.6151
R17636 vdd.n2451 vdd.n2449 10.6151
R17637 vdd.n2452 vdd.n2451 10.6151
R17638 vdd.n2454 vdd.n2452 10.6151
R17639 vdd.n2455 vdd.n2454 10.6151
R17640 vdd.n2470 vdd.n2455 10.6151
R17641 vdd.n2470 vdd.n2469 10.6151
R17642 vdd.n2469 vdd.n2468 10.6151
R17643 vdd.n2468 vdd.n2466 10.6151
R17644 vdd.n2466 vdd.n2465 10.6151
R17645 vdd.n2465 vdd.n2463 10.6151
R17646 vdd.n2463 vdd.n2462 10.6151
R17647 vdd.n2462 vdd.n2460 10.6151
R17648 vdd.n2460 vdd.n2459 10.6151
R17649 vdd.n2459 vdd.n2457 10.6151
R17650 vdd.n2457 vdd.n2456 10.6151
R17651 vdd.n2456 vdd.n664 10.6151
R17652 vdd.n2704 vdd.n664 10.6151
R17653 vdd.n2705 vdd.n2704 10.6151
R17654 vdd.n2566 vdd.n740 10.6151
R17655 vdd.n2566 vdd.n2565 10.6151
R17656 vdd.n2565 vdd.n2564 10.6151
R17657 vdd.n2564 vdd.n2562 10.6151
R17658 vdd.n2562 vdd.n2559 10.6151
R17659 vdd.n2559 vdd.n2558 10.6151
R17660 vdd.n2558 vdd.n2555 10.6151
R17661 vdd.n2555 vdd.n2554 10.6151
R17662 vdd.n2554 vdd.n2551 10.6151
R17663 vdd.n2551 vdd.n2550 10.6151
R17664 vdd.n2550 vdd.n2547 10.6151
R17665 vdd.n2547 vdd.n2546 10.6151
R17666 vdd.n2546 vdd.n2543 10.6151
R17667 vdd.n2543 vdd.n2542 10.6151
R17668 vdd.n2542 vdd.n2539 10.6151
R17669 vdd.n2539 vdd.n2538 10.6151
R17670 vdd.n2538 vdd.n2535 10.6151
R17671 vdd.n2535 vdd.n2534 10.6151
R17672 vdd.n2534 vdd.n2531 10.6151
R17673 vdd.n2531 vdd.n2530 10.6151
R17674 vdd.n2530 vdd.n2527 10.6151
R17675 vdd.n2527 vdd.n2526 10.6151
R17676 vdd.n2526 vdd.n2523 10.6151
R17677 vdd.n2523 vdd.n2522 10.6151
R17678 vdd.n2522 vdd.n2519 10.6151
R17679 vdd.n2519 vdd.n2518 10.6151
R17680 vdd.n2518 vdd.n2515 10.6151
R17681 vdd.n2515 vdd.n2514 10.6151
R17682 vdd.n2514 vdd.n2511 10.6151
R17683 vdd.n2511 vdd.n2510 10.6151
R17684 vdd.n2510 vdd.n2507 10.6151
R17685 vdd.n2505 vdd.n2502 10.6151
R17686 vdd.n2502 vdd.n2501 10.6151
R17687 vdd.n2579 vdd.n2578 10.6151
R17688 vdd.n2580 vdd.n2579 10.6151
R17689 vdd.n2580 vdd.n730 10.6151
R17690 vdd.n2590 vdd.n730 10.6151
R17691 vdd.n2591 vdd.n2590 10.6151
R17692 vdd.n2592 vdd.n2591 10.6151
R17693 vdd.n2592 vdd.n717 10.6151
R17694 vdd.n2602 vdd.n717 10.6151
R17695 vdd.n2603 vdd.n2602 10.6151
R17696 vdd.n2604 vdd.n2603 10.6151
R17697 vdd.n2604 vdd.n706 10.6151
R17698 vdd.n2614 vdd.n706 10.6151
R17699 vdd.n2615 vdd.n2614 10.6151
R17700 vdd.n2616 vdd.n2615 10.6151
R17701 vdd.n2616 vdd.n694 10.6151
R17702 vdd.n2626 vdd.n694 10.6151
R17703 vdd.n2627 vdd.n2626 10.6151
R17704 vdd.n2628 vdd.n2627 10.6151
R17705 vdd.n2628 vdd.n683 10.6151
R17706 vdd.n2640 vdd.n683 10.6151
R17707 vdd.n2641 vdd.n2640 10.6151
R17708 vdd.n2642 vdd.n2641 10.6151
R17709 vdd.n2642 vdd.n669 10.6151
R17710 vdd.n2697 vdd.n669 10.6151
R17711 vdd.n2698 vdd.n2697 10.6151
R17712 vdd.n2699 vdd.n2698 10.6151
R17713 vdd.n2699 vdd.n636 10.6151
R17714 vdd.n2769 vdd.n636 10.6151
R17715 vdd.n2768 vdd.n2767 10.6151
R17716 vdd.n2767 vdd.n637 10.6151
R17717 vdd.n638 vdd.n637 10.6151
R17718 vdd.n2760 vdd.n638 10.6151
R17719 vdd.n2760 vdd.n2759 10.6151
R17720 vdd.n2759 vdd.n2758 10.6151
R17721 vdd.n2758 vdd.n640 10.6151
R17722 vdd.n2753 vdd.n640 10.6151
R17723 vdd.n2753 vdd.n2752 10.6151
R17724 vdd.n2752 vdd.n2751 10.6151
R17725 vdd.n2751 vdd.n643 10.6151
R17726 vdd.n2746 vdd.n643 10.6151
R17727 vdd.n2746 vdd.n2745 10.6151
R17728 vdd.n2745 vdd.n2744 10.6151
R17729 vdd.n2744 vdd.n646 10.6151
R17730 vdd.n2739 vdd.n646 10.6151
R17731 vdd.n2739 vdd.n2738 10.6151
R17732 vdd.n2738 vdd.n2736 10.6151
R17733 vdd.n2736 vdd.n649 10.6151
R17734 vdd.n2731 vdd.n649 10.6151
R17735 vdd.n2731 vdd.n2730 10.6151
R17736 vdd.n2730 vdd.n2729 10.6151
R17737 vdd.n2729 vdd.n652 10.6151
R17738 vdd.n2724 vdd.n652 10.6151
R17739 vdd.n2724 vdd.n2723 10.6151
R17740 vdd.n2723 vdd.n2722 10.6151
R17741 vdd.n2722 vdd.n655 10.6151
R17742 vdd.n2717 vdd.n655 10.6151
R17743 vdd.n2717 vdd.n2716 10.6151
R17744 vdd.n2716 vdd.n2715 10.6151
R17745 vdd.n2715 vdd.n658 10.6151
R17746 vdd.n2710 vdd.n2709 10.6151
R17747 vdd.n2709 vdd.n2708 10.6151
R17748 vdd.n2687 vdd.n2648 10.6151
R17749 vdd.n2682 vdd.n2648 10.6151
R17750 vdd.n2682 vdd.n2681 10.6151
R17751 vdd.n2681 vdd.n2680 10.6151
R17752 vdd.n2680 vdd.n2650 10.6151
R17753 vdd.n2675 vdd.n2650 10.6151
R17754 vdd.n2675 vdd.n2674 10.6151
R17755 vdd.n2674 vdd.n2673 10.6151
R17756 vdd.n2673 vdd.n2653 10.6151
R17757 vdd.n2668 vdd.n2653 10.6151
R17758 vdd.n2668 vdd.n2667 10.6151
R17759 vdd.n2667 vdd.n2666 10.6151
R17760 vdd.n2666 vdd.n2656 10.6151
R17761 vdd.n2661 vdd.n2656 10.6151
R17762 vdd.n2661 vdd.n2660 10.6151
R17763 vdd.n2660 vdd.n610 10.6151
R17764 vdd.n2804 vdd.n610 10.6151
R17765 vdd.n2804 vdd.n611 10.6151
R17766 vdd.n614 vdd.n611 10.6151
R17767 vdd.n2797 vdd.n614 10.6151
R17768 vdd.n2797 vdd.n2796 10.6151
R17769 vdd.n2796 vdd.n2795 10.6151
R17770 vdd.n2795 vdd.n616 10.6151
R17771 vdd.n2790 vdd.n616 10.6151
R17772 vdd.n2790 vdd.n2789 10.6151
R17773 vdd.n2789 vdd.n2788 10.6151
R17774 vdd.n2788 vdd.n619 10.6151
R17775 vdd.n2783 vdd.n619 10.6151
R17776 vdd.n2783 vdd.n2782 10.6151
R17777 vdd.n2782 vdd.n2781 10.6151
R17778 vdd.n2781 vdd.n622 10.6151
R17779 vdd.n2776 vdd.n2775 10.6151
R17780 vdd.n2775 vdd.n2774 10.6151
R17781 vdd.n2422 vdd.n2420 10.6151
R17782 vdd.n2423 vdd.n2422 10.6151
R17783 vdd.n2491 vdd.n2423 10.6151
R17784 vdd.n2491 vdd.n2490 10.6151
R17785 vdd.n2490 vdd.n2489 10.6151
R17786 vdd.n2489 vdd.n2487 10.6151
R17787 vdd.n2487 vdd.n2486 10.6151
R17788 vdd.n2486 vdd.n2484 10.6151
R17789 vdd.n2484 vdd.n2483 10.6151
R17790 vdd.n2483 vdd.n2481 10.6151
R17791 vdd.n2481 vdd.n2480 10.6151
R17792 vdd.n2480 vdd.n2478 10.6151
R17793 vdd.n2478 vdd.n2477 10.6151
R17794 vdd.n2477 vdd.n2475 10.6151
R17795 vdd.n2475 vdd.n2474 10.6151
R17796 vdd.n2474 vdd.n2440 10.6151
R17797 vdd.n2440 vdd.n2439 10.6151
R17798 vdd.n2439 vdd.n2437 10.6151
R17799 vdd.n2437 vdd.n2436 10.6151
R17800 vdd.n2436 vdd.n2434 10.6151
R17801 vdd.n2434 vdd.n2433 10.6151
R17802 vdd.n2433 vdd.n2431 10.6151
R17803 vdd.n2431 vdd.n2430 10.6151
R17804 vdd.n2430 vdd.n2428 10.6151
R17805 vdd.n2428 vdd.n2427 10.6151
R17806 vdd.n2427 vdd.n2425 10.6151
R17807 vdd.n2425 vdd.n2424 10.6151
R17808 vdd.n2424 vdd.n628 10.6151
R17809 vdd.n2573 vdd.n2572 10.6151
R17810 vdd.n2572 vdd.n745 10.6151
R17811 vdd.n2357 vdd.n745 10.6151
R17812 vdd.n2360 vdd.n2357 10.6151
R17813 vdd.n2361 vdd.n2360 10.6151
R17814 vdd.n2364 vdd.n2361 10.6151
R17815 vdd.n2365 vdd.n2364 10.6151
R17816 vdd.n2368 vdd.n2365 10.6151
R17817 vdd.n2369 vdd.n2368 10.6151
R17818 vdd.n2372 vdd.n2369 10.6151
R17819 vdd.n2373 vdd.n2372 10.6151
R17820 vdd.n2376 vdd.n2373 10.6151
R17821 vdd.n2377 vdd.n2376 10.6151
R17822 vdd.n2380 vdd.n2377 10.6151
R17823 vdd.n2381 vdd.n2380 10.6151
R17824 vdd.n2384 vdd.n2381 10.6151
R17825 vdd.n2385 vdd.n2384 10.6151
R17826 vdd.n2388 vdd.n2385 10.6151
R17827 vdd.n2389 vdd.n2388 10.6151
R17828 vdd.n2392 vdd.n2389 10.6151
R17829 vdd.n2393 vdd.n2392 10.6151
R17830 vdd.n2396 vdd.n2393 10.6151
R17831 vdd.n2397 vdd.n2396 10.6151
R17832 vdd.n2400 vdd.n2397 10.6151
R17833 vdd.n2401 vdd.n2400 10.6151
R17834 vdd.n2404 vdd.n2401 10.6151
R17835 vdd.n2405 vdd.n2404 10.6151
R17836 vdd.n2408 vdd.n2405 10.6151
R17837 vdd.n2409 vdd.n2408 10.6151
R17838 vdd.n2412 vdd.n2409 10.6151
R17839 vdd.n2413 vdd.n2412 10.6151
R17840 vdd.n2418 vdd.n2416 10.6151
R17841 vdd.n2419 vdd.n2418 10.6151
R17842 vdd.n2574 vdd.n735 10.6151
R17843 vdd.n2584 vdd.n735 10.6151
R17844 vdd.n2585 vdd.n2584 10.6151
R17845 vdd.n2586 vdd.n2585 10.6151
R17846 vdd.n2586 vdd.n723 10.6151
R17847 vdd.n2596 vdd.n723 10.6151
R17848 vdd.n2597 vdd.n2596 10.6151
R17849 vdd.n2598 vdd.n2597 10.6151
R17850 vdd.n2598 vdd.n712 10.6151
R17851 vdd.n2608 vdd.n712 10.6151
R17852 vdd.n2609 vdd.n2608 10.6151
R17853 vdd.n2610 vdd.n2609 10.6151
R17854 vdd.n2610 vdd.n700 10.6151
R17855 vdd.n2620 vdd.n700 10.6151
R17856 vdd.n2621 vdd.n2620 10.6151
R17857 vdd.n2622 vdd.n2621 10.6151
R17858 vdd.n2622 vdd.n689 10.6151
R17859 vdd.n2632 vdd.n689 10.6151
R17860 vdd.n2633 vdd.n2632 10.6151
R17861 vdd.n2636 vdd.n2633 10.6151
R17862 vdd.n2646 vdd.n677 10.6151
R17863 vdd.n2647 vdd.n2646 10.6151
R17864 vdd.n2693 vdd.n2647 10.6151
R17865 vdd.n2693 vdd.n2692 10.6151
R17866 vdd.n2692 vdd.n2691 10.6151
R17867 vdd.n2691 vdd.n2690 10.6151
R17868 vdd.n2690 vdd.n2688 10.6151
R17869 vdd.n2085 vdd.n869 10.6151
R17870 vdd.n2095 vdd.n869 10.6151
R17871 vdd.n2096 vdd.n2095 10.6151
R17872 vdd.n2097 vdd.n2096 10.6151
R17873 vdd.n2097 vdd.n856 10.6151
R17874 vdd.n2107 vdd.n856 10.6151
R17875 vdd.n2108 vdd.n2107 10.6151
R17876 vdd.n2110 vdd.n844 10.6151
R17877 vdd.n2120 vdd.n844 10.6151
R17878 vdd.n2121 vdd.n2120 10.6151
R17879 vdd.n2122 vdd.n2121 10.6151
R17880 vdd.n2122 vdd.n832 10.6151
R17881 vdd.n2132 vdd.n832 10.6151
R17882 vdd.n2133 vdd.n2132 10.6151
R17883 vdd.n2134 vdd.n2133 10.6151
R17884 vdd.n2134 vdd.n821 10.6151
R17885 vdd.n2144 vdd.n821 10.6151
R17886 vdd.n2145 vdd.n2144 10.6151
R17887 vdd.n2146 vdd.n2145 10.6151
R17888 vdd.n2146 vdd.n809 10.6151
R17889 vdd.n2156 vdd.n809 10.6151
R17890 vdd.n2157 vdd.n2156 10.6151
R17891 vdd.n2160 vdd.n2157 10.6151
R17892 vdd.n2160 vdd.n2159 10.6151
R17893 vdd.n2159 vdd.n2158 10.6151
R17894 vdd.n2158 vdd.n792 10.6151
R17895 vdd.n2242 vdd.n792 10.6151
R17896 vdd.n2241 vdd.n2240 10.6151
R17897 vdd.n2240 vdd.n2237 10.6151
R17898 vdd.n2237 vdd.n2236 10.6151
R17899 vdd.n2236 vdd.n2233 10.6151
R17900 vdd.n2233 vdd.n2232 10.6151
R17901 vdd.n2232 vdd.n2229 10.6151
R17902 vdd.n2229 vdd.n2228 10.6151
R17903 vdd.n2228 vdd.n2225 10.6151
R17904 vdd.n2225 vdd.n2224 10.6151
R17905 vdd.n2224 vdd.n2221 10.6151
R17906 vdd.n2221 vdd.n2220 10.6151
R17907 vdd.n2220 vdd.n2217 10.6151
R17908 vdd.n2217 vdd.n2216 10.6151
R17909 vdd.n2216 vdd.n2213 10.6151
R17910 vdd.n2213 vdd.n2212 10.6151
R17911 vdd.n2212 vdd.n2209 10.6151
R17912 vdd.n2209 vdd.n2208 10.6151
R17913 vdd.n2208 vdd.n2205 10.6151
R17914 vdd.n2205 vdd.n2204 10.6151
R17915 vdd.n2204 vdd.n2201 10.6151
R17916 vdd.n2201 vdd.n2200 10.6151
R17917 vdd.n2200 vdd.n2197 10.6151
R17918 vdd.n2197 vdd.n2196 10.6151
R17919 vdd.n2196 vdd.n2193 10.6151
R17920 vdd.n2193 vdd.n2192 10.6151
R17921 vdd.n2192 vdd.n2189 10.6151
R17922 vdd.n2189 vdd.n2188 10.6151
R17923 vdd.n2188 vdd.n2185 10.6151
R17924 vdd.n2185 vdd.n2184 10.6151
R17925 vdd.n2184 vdd.n2181 10.6151
R17926 vdd.n2181 vdd.n2180 10.6151
R17927 vdd.n2177 vdd.n2176 10.6151
R17928 vdd.n2176 vdd.n2174 10.6151
R17929 vdd.n1933 vdd.n1931 10.6151
R17930 vdd.n1934 vdd.n1933 10.6151
R17931 vdd.n1936 vdd.n1934 10.6151
R17932 vdd.n1937 vdd.n1936 10.6151
R17933 vdd.n1939 vdd.n1937 10.6151
R17934 vdd.n1940 vdd.n1939 10.6151
R17935 vdd.n1942 vdd.n1940 10.6151
R17936 vdd.n1943 vdd.n1942 10.6151
R17937 vdd.n1945 vdd.n1943 10.6151
R17938 vdd.n1946 vdd.n1945 10.6151
R17939 vdd.n1948 vdd.n1946 10.6151
R17940 vdd.n1949 vdd.n1948 10.6151
R17941 vdd.n1967 vdd.n1949 10.6151
R17942 vdd.n1967 vdd.n1966 10.6151
R17943 vdd.n1966 vdd.n1965 10.6151
R17944 vdd.n1965 vdd.n1963 10.6151
R17945 vdd.n1963 vdd.n1962 10.6151
R17946 vdd.n1962 vdd.n1960 10.6151
R17947 vdd.n1960 vdd.n1959 10.6151
R17948 vdd.n1959 vdd.n1957 10.6151
R17949 vdd.n1957 vdd.n1956 10.6151
R17950 vdd.n1956 vdd.n1954 10.6151
R17951 vdd.n1954 vdd.n1953 10.6151
R17952 vdd.n1953 vdd.n1951 10.6151
R17953 vdd.n1951 vdd.n1950 10.6151
R17954 vdd.n1950 vdd.n796 10.6151
R17955 vdd.n2172 vdd.n796 10.6151
R17956 vdd.n2173 vdd.n2172 10.6151
R17957 vdd.n2084 vdd.n2083 10.6151
R17958 vdd.n2083 vdd.n881 10.6151
R17959 vdd.n2077 vdd.n881 10.6151
R17960 vdd.n2077 vdd.n2076 10.6151
R17961 vdd.n2076 vdd.n2075 10.6151
R17962 vdd.n2075 vdd.n883 10.6151
R17963 vdd.n2069 vdd.n883 10.6151
R17964 vdd.n2069 vdd.n2068 10.6151
R17965 vdd.n2068 vdd.n2067 10.6151
R17966 vdd.n2067 vdd.n885 10.6151
R17967 vdd.n2061 vdd.n885 10.6151
R17968 vdd.n2061 vdd.n2060 10.6151
R17969 vdd.n2060 vdd.n2059 10.6151
R17970 vdd.n2059 vdd.n887 10.6151
R17971 vdd.n2053 vdd.n887 10.6151
R17972 vdd.n2053 vdd.n2052 10.6151
R17973 vdd.n2052 vdd.n2051 10.6151
R17974 vdd.n2051 vdd.n891 10.6151
R17975 vdd.n1899 vdd.n891 10.6151
R17976 vdd.n1900 vdd.n1899 10.6151
R17977 vdd.n1900 vdd.n1895 10.6151
R17978 vdd.n1906 vdd.n1895 10.6151
R17979 vdd.n1907 vdd.n1906 10.6151
R17980 vdd.n1908 vdd.n1907 10.6151
R17981 vdd.n1908 vdd.n1893 10.6151
R17982 vdd.n1914 vdd.n1893 10.6151
R17983 vdd.n1915 vdd.n1914 10.6151
R17984 vdd.n1916 vdd.n1915 10.6151
R17985 vdd.n1916 vdd.n1891 10.6151
R17986 vdd.n1922 vdd.n1891 10.6151
R17987 vdd.n1923 vdd.n1922 10.6151
R17988 vdd.n1925 vdd.n1887 10.6151
R17989 vdd.n1930 vdd.n1887 10.6151
R17990 vdd.n1272 vdd.t2 10.5435
R17991 vdd.n2041 vdd.t94 10.5435
R17992 vdd.n2940 vdd.t87 10.5435
R17993 vdd.n3164 vdd.t189 10.5435
R17994 vdd.n292 vdd.n274 10.4732
R17995 vdd.n241 vdd.n223 10.4732
R17996 vdd.n198 vdd.n180 10.4732
R17997 vdd.n147 vdd.n129 10.4732
R17998 vdd.n105 vdd.n87 10.4732
R17999 vdd.n54 vdd.n36 10.4732
R18000 vdd.n1487 vdd.n1469 10.4732
R18001 vdd.n1538 vdd.n1520 10.4732
R18002 vdd.n1393 vdd.n1375 10.4732
R18003 vdd.n1444 vdd.n1426 10.4732
R18004 vdd.n1300 vdd.n1282 10.4732
R18005 vdd.n1351 vdd.n1333 10.4732
R18006 vdd.n1570 vdd.t6 10.3167
R18007 vdd.t213 vdd.n493 10.3167
R18008 vdd.n1223 vdd.t98 9.86327
R18009 vdd.n3140 vdd.t147 9.86327
R18010 vdd.n291 vdd.n276 9.69747
R18011 vdd.n240 vdd.n225 9.69747
R18012 vdd.n197 vdd.n182 9.69747
R18013 vdd.n146 vdd.n131 9.69747
R18014 vdd.n104 vdd.n89 9.69747
R18015 vdd.n53 vdd.n38 9.69747
R18016 vdd.n1486 vdd.n1471 9.69747
R18017 vdd.n1537 vdd.n1522 9.69747
R18018 vdd.n1392 vdd.n1377 9.69747
R18019 vdd.n1443 vdd.n1428 9.69747
R18020 vdd.n1299 vdd.n1284 9.69747
R18021 vdd.n1350 vdd.n1335 9.69747
R18022 vdd.n2027 vdd.n2026 9.67831
R18023 vdd.n2738 vdd.n2737 9.67831
R18024 vdd.n2805 vdd.n2804 9.67831
R18025 vdd.n2051 vdd.n2050 9.67831
R18026 vdd.n307 vdd.n306 9.45567
R18027 vdd.n256 vdd.n255 9.45567
R18028 vdd.n213 vdd.n212 9.45567
R18029 vdd.n162 vdd.n161 9.45567
R18030 vdd.n120 vdd.n119 9.45567
R18031 vdd.n69 vdd.n68 9.45567
R18032 vdd.n1502 vdd.n1501 9.45567
R18033 vdd.n1553 vdd.n1552 9.45567
R18034 vdd.n1408 vdd.n1407 9.45567
R18035 vdd.n1459 vdd.n1458 9.45567
R18036 vdd.n1315 vdd.n1314 9.45567
R18037 vdd.n1366 vdd.n1365 9.45567
R18038 vdd.n1787 vdd.n1641 9.3005
R18039 vdd.n1786 vdd.n1785 9.3005
R18040 vdd.n1647 vdd.n1646 9.3005
R18041 vdd.n1780 vdd.n1651 9.3005
R18042 vdd.n1779 vdd.n1652 9.3005
R18043 vdd.n1778 vdd.n1653 9.3005
R18044 vdd.n1657 vdd.n1654 9.3005
R18045 vdd.n1773 vdd.n1658 9.3005
R18046 vdd.n1772 vdd.n1659 9.3005
R18047 vdd.n1771 vdd.n1660 9.3005
R18048 vdd.n1664 vdd.n1661 9.3005
R18049 vdd.n1766 vdd.n1665 9.3005
R18050 vdd.n1765 vdd.n1666 9.3005
R18051 vdd.n1764 vdd.n1667 9.3005
R18052 vdd.n1671 vdd.n1668 9.3005
R18053 vdd.n1759 vdd.n1672 9.3005
R18054 vdd.n1758 vdd.n1673 9.3005
R18055 vdd.n1757 vdd.n1674 9.3005
R18056 vdd.n1678 vdd.n1675 9.3005
R18057 vdd.n1752 vdd.n1679 9.3005
R18058 vdd.n1751 vdd.n1680 9.3005
R18059 vdd.n1750 vdd.n1749 9.3005
R18060 vdd.n1748 vdd.n1681 9.3005
R18061 vdd.n1747 vdd.n1746 9.3005
R18062 vdd.n1687 vdd.n1686 9.3005
R18063 vdd.n1741 vdd.n1691 9.3005
R18064 vdd.n1740 vdd.n1692 9.3005
R18065 vdd.n1739 vdd.n1693 9.3005
R18066 vdd.n1697 vdd.n1694 9.3005
R18067 vdd.n1734 vdd.n1698 9.3005
R18068 vdd.n1733 vdd.n1699 9.3005
R18069 vdd.n1732 vdd.n1700 9.3005
R18070 vdd.n1704 vdd.n1701 9.3005
R18071 vdd.n1727 vdd.n1705 9.3005
R18072 vdd.n1726 vdd.n1706 9.3005
R18073 vdd.n1725 vdd.n1707 9.3005
R18074 vdd.n1709 vdd.n1708 9.3005
R18075 vdd.n1720 vdd.n892 9.3005
R18076 vdd.n1789 vdd.n1788 9.3005
R18077 vdd.n1813 vdd.n1812 9.3005
R18078 vdd.n1619 vdd.n1618 9.3005
R18079 vdd.n1624 vdd.n1622 9.3005
R18080 vdd.n1805 vdd.n1625 9.3005
R18081 vdd.n1804 vdd.n1626 9.3005
R18082 vdd.n1803 vdd.n1627 9.3005
R18083 vdd.n1631 vdd.n1628 9.3005
R18084 vdd.n1798 vdd.n1632 9.3005
R18085 vdd.n1797 vdd.n1633 9.3005
R18086 vdd.n1796 vdd.n1634 9.3005
R18087 vdd.n1638 vdd.n1635 9.3005
R18088 vdd.n1791 vdd.n1639 9.3005
R18089 vdd.n1790 vdd.n1640 9.3005
R18090 vdd.n2035 vdd.n1612 9.3005
R18091 vdd.n2037 vdd.n2036 9.3005
R18092 vdd.n1558 vdd.n939 9.3005
R18093 vdd.n1560 vdd.n1559 9.3005
R18094 vdd.n929 vdd.n928 9.3005
R18095 vdd.n1574 vdd.n1573 9.3005
R18096 vdd.n1575 vdd.n927 9.3005
R18097 vdd.n1577 vdd.n1576 9.3005
R18098 vdd.n918 vdd.n917 9.3005
R18099 vdd.n1591 vdd.n1590 9.3005
R18100 vdd.n1592 vdd.n916 9.3005
R18101 vdd.n1594 vdd.n1593 9.3005
R18102 vdd.n906 vdd.n905 9.3005
R18103 vdd.n1610 vdd.n1609 9.3005
R18104 vdd.n1611 vdd.n904 9.3005
R18105 vdd.n2039 vdd.n2038 9.3005
R18106 vdd.n283 vdd.n282 9.3005
R18107 vdd.n278 vdd.n277 9.3005
R18108 vdd.n289 vdd.n288 9.3005
R18109 vdd.n291 vdd.n290 9.3005
R18110 vdd.n274 vdd.n273 9.3005
R18111 vdd.n297 vdd.n296 9.3005
R18112 vdd.n299 vdd.n298 9.3005
R18113 vdd.n271 vdd.n268 9.3005
R18114 vdd.n306 vdd.n305 9.3005
R18115 vdd.n232 vdd.n231 9.3005
R18116 vdd.n227 vdd.n226 9.3005
R18117 vdd.n238 vdd.n237 9.3005
R18118 vdd.n240 vdd.n239 9.3005
R18119 vdd.n223 vdd.n222 9.3005
R18120 vdd.n246 vdd.n245 9.3005
R18121 vdd.n248 vdd.n247 9.3005
R18122 vdd.n220 vdd.n217 9.3005
R18123 vdd.n255 vdd.n254 9.3005
R18124 vdd.n189 vdd.n188 9.3005
R18125 vdd.n184 vdd.n183 9.3005
R18126 vdd.n195 vdd.n194 9.3005
R18127 vdd.n197 vdd.n196 9.3005
R18128 vdd.n180 vdd.n179 9.3005
R18129 vdd.n203 vdd.n202 9.3005
R18130 vdd.n205 vdd.n204 9.3005
R18131 vdd.n177 vdd.n174 9.3005
R18132 vdd.n212 vdd.n211 9.3005
R18133 vdd.n138 vdd.n137 9.3005
R18134 vdd.n133 vdd.n132 9.3005
R18135 vdd.n144 vdd.n143 9.3005
R18136 vdd.n146 vdd.n145 9.3005
R18137 vdd.n129 vdd.n128 9.3005
R18138 vdd.n152 vdd.n151 9.3005
R18139 vdd.n154 vdd.n153 9.3005
R18140 vdd.n126 vdd.n123 9.3005
R18141 vdd.n161 vdd.n160 9.3005
R18142 vdd.n96 vdd.n95 9.3005
R18143 vdd.n91 vdd.n90 9.3005
R18144 vdd.n102 vdd.n101 9.3005
R18145 vdd.n104 vdd.n103 9.3005
R18146 vdd.n87 vdd.n86 9.3005
R18147 vdd.n110 vdd.n109 9.3005
R18148 vdd.n112 vdd.n111 9.3005
R18149 vdd.n84 vdd.n81 9.3005
R18150 vdd.n119 vdd.n118 9.3005
R18151 vdd.n45 vdd.n44 9.3005
R18152 vdd.n40 vdd.n39 9.3005
R18153 vdd.n51 vdd.n50 9.3005
R18154 vdd.n53 vdd.n52 9.3005
R18155 vdd.n36 vdd.n35 9.3005
R18156 vdd.n59 vdd.n58 9.3005
R18157 vdd.n61 vdd.n60 9.3005
R18158 vdd.n33 vdd.n30 9.3005
R18159 vdd.n68 vdd.n67 9.3005
R18160 vdd.n2854 vdd.n2853 9.3005
R18161 vdd.n2855 vdd.n578 9.3005
R18162 vdd.n577 vdd.n575 9.3005
R18163 vdd.n2861 vdd.n574 9.3005
R18164 vdd.n2862 vdd.n573 9.3005
R18165 vdd.n2863 vdd.n572 9.3005
R18166 vdd.n571 vdd.n569 9.3005
R18167 vdd.n2869 vdd.n568 9.3005
R18168 vdd.n2870 vdd.n567 9.3005
R18169 vdd.n2871 vdd.n566 9.3005
R18170 vdd.n565 vdd.n563 9.3005
R18171 vdd.n2877 vdd.n562 9.3005
R18172 vdd.n2878 vdd.n561 9.3005
R18173 vdd.n2879 vdd.n560 9.3005
R18174 vdd.n559 vdd.n557 9.3005
R18175 vdd.n2885 vdd.n556 9.3005
R18176 vdd.n2886 vdd.n555 9.3005
R18177 vdd.n2887 vdd.n554 9.3005
R18178 vdd.n553 vdd.n551 9.3005
R18179 vdd.n2893 vdd.n550 9.3005
R18180 vdd.n2894 vdd.n549 9.3005
R18181 vdd.n2895 vdd.n548 9.3005
R18182 vdd.n547 vdd.n545 9.3005
R18183 vdd.n2901 vdd.n542 9.3005
R18184 vdd.n2902 vdd.n541 9.3005
R18185 vdd.n2903 vdd.n540 9.3005
R18186 vdd.n539 vdd.n537 9.3005
R18187 vdd.n2909 vdd.n536 9.3005
R18188 vdd.n2910 vdd.n535 9.3005
R18189 vdd.n2911 vdd.n534 9.3005
R18190 vdd.n533 vdd.n531 9.3005
R18191 vdd.n2917 vdd.n530 9.3005
R18192 vdd.n2918 vdd.n529 9.3005
R18193 vdd.n2919 vdd.n528 9.3005
R18194 vdd.n527 vdd.n525 9.3005
R18195 vdd.n2924 vdd.n524 9.3005
R18196 vdd.n2934 vdd.n518 9.3005
R18197 vdd.n2936 vdd.n2935 9.3005
R18198 vdd.n509 vdd.n508 9.3005
R18199 vdd.n2951 vdd.n2950 9.3005
R18200 vdd.n2952 vdd.n507 9.3005
R18201 vdd.n2954 vdd.n2953 9.3005
R18202 vdd.n497 vdd.n496 9.3005
R18203 vdd.n2967 vdd.n2966 9.3005
R18204 vdd.n2968 vdd.n495 9.3005
R18205 vdd.n2970 vdd.n2969 9.3005
R18206 vdd.n485 vdd.n484 9.3005
R18207 vdd.n2984 vdd.n2983 9.3005
R18208 vdd.n2985 vdd.n483 9.3005
R18209 vdd.n2987 vdd.n2986 9.3005
R18210 vdd.n312 vdd.n310 9.3005
R18211 vdd.n2938 vdd.n2937 9.3005
R18212 vdd.n3167 vdd.n3166 9.3005
R18213 vdd.n313 vdd.n311 9.3005
R18214 vdd.n3160 vdd.n320 9.3005
R18215 vdd.n3159 vdd.n321 9.3005
R18216 vdd.n3158 vdd.n322 9.3005
R18217 vdd.n331 vdd.n323 9.3005
R18218 vdd.n3152 vdd.n332 9.3005
R18219 vdd.n3151 vdd.n333 9.3005
R18220 vdd.n3150 vdd.n334 9.3005
R18221 vdd.n342 vdd.n335 9.3005
R18222 vdd.n3144 vdd.n343 9.3005
R18223 vdd.n3143 vdd.n344 9.3005
R18224 vdd.n3142 vdd.n345 9.3005
R18225 vdd.n353 vdd.n346 9.3005
R18226 vdd.n3136 vdd.n3135 9.3005
R18227 vdd.n3132 vdd.n354 9.3005
R18228 vdd.n3131 vdd.n357 9.3005
R18229 vdd.n361 vdd.n358 9.3005
R18230 vdd.n362 vdd.n359 9.3005
R18231 vdd.n3124 vdd.n363 9.3005
R18232 vdd.n3123 vdd.n364 9.3005
R18233 vdd.n3122 vdd.n365 9.3005
R18234 vdd.n369 vdd.n366 9.3005
R18235 vdd.n3117 vdd.n370 9.3005
R18236 vdd.n3116 vdd.n371 9.3005
R18237 vdd.n3115 vdd.n372 9.3005
R18238 vdd.n376 vdd.n373 9.3005
R18239 vdd.n3110 vdd.n377 9.3005
R18240 vdd.n3109 vdd.n378 9.3005
R18241 vdd.n3108 vdd.n379 9.3005
R18242 vdd.n383 vdd.n380 9.3005
R18243 vdd.n3103 vdd.n384 9.3005
R18244 vdd.n3102 vdd.n385 9.3005
R18245 vdd.n3101 vdd.n3100 9.3005
R18246 vdd.n3099 vdd.n386 9.3005
R18247 vdd.n3098 vdd.n3097 9.3005
R18248 vdd.n392 vdd.n391 9.3005
R18249 vdd.n3092 vdd.n396 9.3005
R18250 vdd.n3091 vdd.n397 9.3005
R18251 vdd.n3090 vdd.n398 9.3005
R18252 vdd.n402 vdd.n399 9.3005
R18253 vdd.n3085 vdd.n403 9.3005
R18254 vdd.n3084 vdd.n404 9.3005
R18255 vdd.n3083 vdd.n405 9.3005
R18256 vdd.n409 vdd.n406 9.3005
R18257 vdd.n3078 vdd.n410 9.3005
R18258 vdd.n3077 vdd.n411 9.3005
R18259 vdd.n3076 vdd.n412 9.3005
R18260 vdd.n416 vdd.n413 9.3005
R18261 vdd.n3071 vdd.n417 9.3005
R18262 vdd.n3070 vdd.n418 9.3005
R18263 vdd.n3069 vdd.n419 9.3005
R18264 vdd.n423 vdd.n420 9.3005
R18265 vdd.n3064 vdd.n424 9.3005
R18266 vdd.n3063 vdd.n425 9.3005
R18267 vdd.n3062 vdd.n3061 9.3005
R18268 vdd.n3060 vdd.n426 9.3005
R18269 vdd.n3059 vdd.n3058 9.3005
R18270 vdd.n432 vdd.n431 9.3005
R18271 vdd.n3053 vdd.n436 9.3005
R18272 vdd.n3052 vdd.n437 9.3005
R18273 vdd.n3051 vdd.n438 9.3005
R18274 vdd.n442 vdd.n439 9.3005
R18275 vdd.n3046 vdd.n443 9.3005
R18276 vdd.n3045 vdd.n444 9.3005
R18277 vdd.n3044 vdd.n445 9.3005
R18278 vdd.n449 vdd.n446 9.3005
R18279 vdd.n3039 vdd.n450 9.3005
R18280 vdd.n3038 vdd.n451 9.3005
R18281 vdd.n3037 vdd.n452 9.3005
R18282 vdd.n456 vdd.n453 9.3005
R18283 vdd.n3032 vdd.n457 9.3005
R18284 vdd.n3031 vdd.n458 9.3005
R18285 vdd.n3030 vdd.n459 9.3005
R18286 vdd.n463 vdd.n460 9.3005
R18287 vdd.n3025 vdd.n464 9.3005
R18288 vdd.n3024 vdd.n465 9.3005
R18289 vdd.n3020 vdd.n3017 9.3005
R18290 vdd.n3134 vdd.n3133 9.3005
R18291 vdd.n2944 vdd.n513 9.3005
R18292 vdd.n2946 vdd.n2945 9.3005
R18293 vdd.n503 vdd.n502 9.3005
R18294 vdd.n2959 vdd.n2958 9.3005
R18295 vdd.n2960 vdd.n501 9.3005
R18296 vdd.n2962 vdd.n2961 9.3005
R18297 vdd.n490 vdd.n489 9.3005
R18298 vdd.n2975 vdd.n2974 9.3005
R18299 vdd.n2976 vdd.n488 9.3005
R18300 vdd.n2978 vdd.n2977 9.3005
R18301 vdd.n478 vdd.n477 9.3005
R18302 vdd.n2992 vdd.n2991 9.3005
R18303 vdd.n2993 vdd.n476 9.3005
R18304 vdd.n2995 vdd.n2994 9.3005
R18305 vdd.n2996 vdd.n475 9.3005
R18306 vdd.n2998 vdd.n2997 9.3005
R18307 vdd.n2999 vdd.n474 9.3005
R18308 vdd.n3001 vdd.n3000 9.3005
R18309 vdd.n3002 vdd.n472 9.3005
R18310 vdd.n3004 vdd.n3003 9.3005
R18311 vdd.n3005 vdd.n471 9.3005
R18312 vdd.n3007 vdd.n3006 9.3005
R18313 vdd.n3008 vdd.n469 9.3005
R18314 vdd.n3010 vdd.n3009 9.3005
R18315 vdd.n3011 vdd.n468 9.3005
R18316 vdd.n3013 vdd.n3012 9.3005
R18317 vdd.n3014 vdd.n466 9.3005
R18318 vdd.n3016 vdd.n3015 9.3005
R18319 vdd.n2943 vdd.n2942 9.3005
R18320 vdd.n2807 vdd.n514 9.3005
R18321 vdd.n2812 vdd.n2806 9.3005
R18322 vdd.n2822 vdd.n605 9.3005
R18323 vdd.n2823 vdd.n604 9.3005
R18324 vdd.n603 vdd.n601 9.3005
R18325 vdd.n2829 vdd.n600 9.3005
R18326 vdd.n2830 vdd.n599 9.3005
R18327 vdd.n2831 vdd.n598 9.3005
R18328 vdd.n597 vdd.n595 9.3005
R18329 vdd.n2837 vdd.n594 9.3005
R18330 vdd.n2838 vdd.n593 9.3005
R18331 vdd.n2839 vdd.n592 9.3005
R18332 vdd.n591 vdd.n589 9.3005
R18333 vdd.n2844 vdd.n588 9.3005
R18334 vdd.n2845 vdd.n587 9.3005
R18335 vdd.n583 vdd.n582 9.3005
R18336 vdd.n2851 vdd.n2850 9.3005
R18337 vdd.n2852 vdd.n579 9.3005
R18338 vdd.n2049 vdd.n2048 9.3005
R18339 vdd.n2044 vdd.n895 9.3005
R18340 vdd.n1219 vdd.n979 9.3005
R18341 vdd.n1221 vdd.n1220 9.3005
R18342 vdd.n970 vdd.n969 9.3005
R18343 vdd.n1234 vdd.n1233 9.3005
R18344 vdd.n1235 vdd.n968 9.3005
R18345 vdd.n1237 vdd.n1236 9.3005
R18346 vdd.n957 vdd.n956 9.3005
R18347 vdd.n1250 vdd.n1249 9.3005
R18348 vdd.n1251 vdd.n955 9.3005
R18349 vdd.n1253 vdd.n1252 9.3005
R18350 vdd.n946 vdd.n945 9.3005
R18351 vdd.n1267 vdd.n1266 9.3005
R18352 vdd.n1268 vdd.n944 9.3005
R18353 vdd.n1270 vdd.n1269 9.3005
R18354 vdd.n935 vdd.n934 9.3005
R18355 vdd.n1565 vdd.n1564 9.3005
R18356 vdd.n1566 vdd.n933 9.3005
R18357 vdd.n1568 vdd.n1567 9.3005
R18358 vdd.n923 vdd.n922 9.3005
R18359 vdd.n1582 vdd.n1581 9.3005
R18360 vdd.n1583 vdd.n921 9.3005
R18361 vdd.n1585 vdd.n1584 9.3005
R18362 vdd.n913 vdd.n912 9.3005
R18363 vdd.n1599 vdd.n1598 9.3005
R18364 vdd.n1600 vdd.n910 9.3005
R18365 vdd.n1604 vdd.n1603 9.3005
R18366 vdd.n1602 vdd.n911 9.3005
R18367 vdd.n1601 vdd.n900 9.3005
R18368 vdd.n1218 vdd.n1217 9.3005
R18369 vdd.n1113 vdd.n1103 9.3005
R18370 vdd.n1115 vdd.n1114 9.3005
R18371 vdd.n1116 vdd.n1102 9.3005
R18372 vdd.n1118 vdd.n1117 9.3005
R18373 vdd.n1119 vdd.n1095 9.3005
R18374 vdd.n1121 vdd.n1120 9.3005
R18375 vdd.n1122 vdd.n1094 9.3005
R18376 vdd.n1124 vdd.n1123 9.3005
R18377 vdd.n1125 vdd.n1087 9.3005
R18378 vdd.n1127 vdd.n1126 9.3005
R18379 vdd.n1128 vdd.n1086 9.3005
R18380 vdd.n1130 vdd.n1129 9.3005
R18381 vdd.n1131 vdd.n1079 9.3005
R18382 vdd.n1133 vdd.n1132 9.3005
R18383 vdd.n1134 vdd.n1078 9.3005
R18384 vdd.n1136 vdd.n1135 9.3005
R18385 vdd.n1137 vdd.n1072 9.3005
R18386 vdd.n1139 vdd.n1138 9.3005
R18387 vdd.n1140 vdd.n1070 9.3005
R18388 vdd.n1142 vdd.n1141 9.3005
R18389 vdd.n1071 vdd.n1068 9.3005
R18390 vdd.n1149 vdd.n1064 9.3005
R18391 vdd.n1151 vdd.n1150 9.3005
R18392 vdd.n1152 vdd.n1063 9.3005
R18393 vdd.n1154 vdd.n1153 9.3005
R18394 vdd.n1155 vdd.n1056 9.3005
R18395 vdd.n1157 vdd.n1156 9.3005
R18396 vdd.n1158 vdd.n1055 9.3005
R18397 vdd.n1160 vdd.n1159 9.3005
R18398 vdd.n1161 vdd.n1048 9.3005
R18399 vdd.n1163 vdd.n1162 9.3005
R18400 vdd.n1164 vdd.n1047 9.3005
R18401 vdd.n1166 vdd.n1165 9.3005
R18402 vdd.n1167 vdd.n1040 9.3005
R18403 vdd.n1169 vdd.n1168 9.3005
R18404 vdd.n1170 vdd.n1039 9.3005
R18405 vdd.n1172 vdd.n1171 9.3005
R18406 vdd.n1173 vdd.n1032 9.3005
R18407 vdd.n1175 vdd.n1174 9.3005
R18408 vdd.n1176 vdd.n1031 9.3005
R18409 vdd.n1178 vdd.n1177 9.3005
R18410 vdd.n1179 vdd.n1024 9.3005
R18411 vdd.n1181 vdd.n1180 9.3005
R18412 vdd.n1182 vdd.n1023 9.3005
R18413 vdd.n1184 vdd.n1183 9.3005
R18414 vdd.n1185 vdd.n1014 9.3005
R18415 vdd.n1187 vdd.n1186 9.3005
R18416 vdd.n1188 vdd.n1013 9.3005
R18417 vdd.n1190 vdd.n1189 9.3005
R18418 vdd.n1191 vdd.n1006 9.3005
R18419 vdd.n1193 vdd.n1192 9.3005
R18420 vdd.n1194 vdd.n1005 9.3005
R18421 vdd.n1196 vdd.n1195 9.3005
R18422 vdd.n1197 vdd.n998 9.3005
R18423 vdd.n1199 vdd.n1198 9.3005
R18424 vdd.n1200 vdd.n997 9.3005
R18425 vdd.n1202 vdd.n1201 9.3005
R18426 vdd.n1203 vdd.n990 9.3005
R18427 vdd.n1205 vdd.n1204 9.3005
R18428 vdd.n1206 vdd.n989 9.3005
R18429 vdd.n1208 vdd.n1207 9.3005
R18430 vdd.n1209 vdd.n985 9.3005
R18431 vdd.n1211 vdd.n1210 9.3005
R18432 vdd.n1109 vdd.n980 9.3005
R18433 vdd.n976 vdd.n975 9.3005
R18434 vdd.n1226 vdd.n1225 9.3005
R18435 vdd.n1227 vdd.n974 9.3005
R18436 vdd.n1229 vdd.n1228 9.3005
R18437 vdd.n964 vdd.n963 9.3005
R18438 vdd.n1242 vdd.n1241 9.3005
R18439 vdd.n1243 vdd.n962 9.3005
R18440 vdd.n1245 vdd.n1244 9.3005
R18441 vdd.n952 vdd.n951 9.3005
R18442 vdd.n1259 vdd.n1258 9.3005
R18443 vdd.n1260 vdd.n950 9.3005
R18444 vdd.n1262 vdd.n1261 9.3005
R18445 vdd.n941 vdd.n940 9.3005
R18446 vdd.n1213 vdd.n1212 9.3005
R18447 vdd.n1557 vdd.n1274 9.3005
R18448 vdd.n1478 vdd.n1477 9.3005
R18449 vdd.n1473 vdd.n1472 9.3005
R18450 vdd.n1484 vdd.n1483 9.3005
R18451 vdd.n1486 vdd.n1485 9.3005
R18452 vdd.n1469 vdd.n1468 9.3005
R18453 vdd.n1492 vdd.n1491 9.3005
R18454 vdd.n1494 vdd.n1493 9.3005
R18455 vdd.n1466 vdd.n1463 9.3005
R18456 vdd.n1501 vdd.n1500 9.3005
R18457 vdd.n1529 vdd.n1528 9.3005
R18458 vdd.n1524 vdd.n1523 9.3005
R18459 vdd.n1535 vdd.n1534 9.3005
R18460 vdd.n1537 vdd.n1536 9.3005
R18461 vdd.n1520 vdd.n1519 9.3005
R18462 vdd.n1543 vdd.n1542 9.3005
R18463 vdd.n1545 vdd.n1544 9.3005
R18464 vdd.n1517 vdd.n1514 9.3005
R18465 vdd.n1552 vdd.n1551 9.3005
R18466 vdd.n1384 vdd.n1383 9.3005
R18467 vdd.n1379 vdd.n1378 9.3005
R18468 vdd.n1390 vdd.n1389 9.3005
R18469 vdd.n1392 vdd.n1391 9.3005
R18470 vdd.n1375 vdd.n1374 9.3005
R18471 vdd.n1398 vdd.n1397 9.3005
R18472 vdd.n1400 vdd.n1399 9.3005
R18473 vdd.n1372 vdd.n1369 9.3005
R18474 vdd.n1407 vdd.n1406 9.3005
R18475 vdd.n1435 vdd.n1434 9.3005
R18476 vdd.n1430 vdd.n1429 9.3005
R18477 vdd.n1441 vdd.n1440 9.3005
R18478 vdd.n1443 vdd.n1442 9.3005
R18479 vdd.n1426 vdd.n1425 9.3005
R18480 vdd.n1449 vdd.n1448 9.3005
R18481 vdd.n1451 vdd.n1450 9.3005
R18482 vdd.n1423 vdd.n1420 9.3005
R18483 vdd.n1458 vdd.n1457 9.3005
R18484 vdd.n1291 vdd.n1290 9.3005
R18485 vdd.n1286 vdd.n1285 9.3005
R18486 vdd.n1297 vdd.n1296 9.3005
R18487 vdd.n1299 vdd.n1298 9.3005
R18488 vdd.n1282 vdd.n1281 9.3005
R18489 vdd.n1305 vdd.n1304 9.3005
R18490 vdd.n1307 vdd.n1306 9.3005
R18491 vdd.n1279 vdd.n1276 9.3005
R18492 vdd.n1314 vdd.n1313 9.3005
R18493 vdd.n1342 vdd.n1341 9.3005
R18494 vdd.n1337 vdd.n1336 9.3005
R18495 vdd.n1348 vdd.n1347 9.3005
R18496 vdd.n1350 vdd.n1349 9.3005
R18497 vdd.n1333 vdd.n1332 9.3005
R18498 vdd.n1356 vdd.n1355 9.3005
R18499 vdd.n1358 vdd.n1357 9.3005
R18500 vdd.n1330 vdd.n1327 9.3005
R18501 vdd.n1365 vdd.n1364 9.3005
R18502 vdd.n288 vdd.n287 8.92171
R18503 vdd.n237 vdd.n236 8.92171
R18504 vdd.n194 vdd.n193 8.92171
R18505 vdd.n143 vdd.n142 8.92171
R18506 vdd.n101 vdd.n100 8.92171
R18507 vdd.n50 vdd.n49 8.92171
R18508 vdd.n1483 vdd.n1482 8.92171
R18509 vdd.n1534 vdd.n1533 8.92171
R18510 vdd.n1389 vdd.n1388 8.92171
R18511 vdd.n1440 vdd.n1439 8.92171
R18512 vdd.n1296 vdd.n1295 8.92171
R18513 vdd.n1347 vdd.n1346 8.92171
R18514 vdd.n215 vdd.n121 8.81535
R18515 vdd.n1461 vdd.n1367 8.81535
R18516 vdd.n1596 vdd.t8 8.72962
R18517 vdd.n2956 vdd.t82 8.72962
R18518 vdd.t29 vdd.n1570 8.50289
R18519 vdd.n493 vdd.t0 8.50289
R18520 vdd.n28 vdd.n14 8.42249
R18521 vdd.n1272 vdd.t26 8.27616
R18522 vdd.n3164 vdd.t63 8.27616
R18523 vdd.n3168 vdd.n3167 8.16225
R18524 vdd.n1557 vdd.n1556 8.16225
R18525 vdd.n284 vdd.n278 8.14595
R18526 vdd.n233 vdd.n227 8.14595
R18527 vdd.n190 vdd.n184 8.14595
R18528 vdd.n139 vdd.n133 8.14595
R18529 vdd.n97 vdd.n91 8.14595
R18530 vdd.n46 vdd.n40 8.14595
R18531 vdd.n1479 vdd.n1473 8.14595
R18532 vdd.n1530 vdd.n1524 8.14595
R18533 vdd.n1385 vdd.n1379 8.14595
R18534 vdd.n1436 vdd.n1430 8.14595
R18535 vdd.n1292 vdd.n1286 8.14595
R18536 vdd.n1343 vdd.n1337 8.14595
R18537 vdd.n2635 vdd.n677 8.11757
R18538 vdd.n2109 vdd.n2108 8.11757
R18539 vdd.t55 vdd.n960 8.04943
R18540 vdd.n3155 vdd.t72 8.04943
R18541 vdd.n2087 vdd.n871 7.70933
R18542 vdd.n2093 vdd.n871 7.70933
R18543 vdd.n2099 vdd.n865 7.70933
R18544 vdd.n2099 vdd.n858 7.70933
R18545 vdd.n2105 vdd.n858 7.70933
R18546 vdd.n2105 vdd.n861 7.70933
R18547 vdd.n2112 vdd.n846 7.70933
R18548 vdd.n2118 vdd.n846 7.70933
R18549 vdd.n2124 vdd.n840 7.70933
R18550 vdd.n2130 vdd.n836 7.70933
R18551 vdd.n2136 vdd.n830 7.70933
R18552 vdd.n2148 vdd.n817 7.70933
R18553 vdd.n2154 vdd.n811 7.70933
R18554 vdd.n2154 vdd.n804 7.70933
R18555 vdd.n2162 vdd.n804 7.70933
R18556 vdd.n2169 vdd.t182 7.70933
R18557 vdd.n2244 vdd.t182 7.70933
R18558 vdd.n2576 vdd.t209 7.70933
R18559 vdd.n2582 vdd.t209 7.70933
R18560 vdd.n2588 vdd.n725 7.70933
R18561 vdd.n2594 vdd.n725 7.70933
R18562 vdd.n2594 vdd.n728 7.70933
R18563 vdd.n2600 vdd.n721 7.70933
R18564 vdd.n2612 vdd.n708 7.70933
R18565 vdd.n2618 vdd.n702 7.70933
R18566 vdd.n2624 vdd.n698 7.70933
R18567 vdd.n2630 vdd.n685 7.70933
R18568 vdd.n2638 vdd.n685 7.70933
R18569 vdd.n2644 vdd.n679 7.70933
R18570 vdd.n2644 vdd.n671 7.70933
R18571 vdd.n2695 vdd.n671 7.70933
R18572 vdd.n2695 vdd.n674 7.70933
R18573 vdd.n2701 vdd.n631 7.70933
R18574 vdd.n2771 vdd.n631 7.70933
R18575 vdd.n283 vdd.n280 7.3702
R18576 vdd.n232 vdd.n229 7.3702
R18577 vdd.n189 vdd.n186 7.3702
R18578 vdd.n138 vdd.n135 7.3702
R18579 vdd.n96 vdd.n93 7.3702
R18580 vdd.n45 vdd.n42 7.3702
R18581 vdd.n1478 vdd.n1475 7.3702
R18582 vdd.n1529 vdd.n1526 7.3702
R18583 vdd.n1384 vdd.n1381 7.3702
R18584 vdd.n1435 vdd.n1432 7.3702
R18585 vdd.n1291 vdd.n1288 7.3702
R18586 vdd.n1342 vdd.n1339 7.3702
R18587 vdd.n1239 vdd.t166 7.1425
R18588 vdd.n3148 vdd.t163 7.1425
R18589 vdd.n1150 vdd.n1149 6.98232
R18590 vdd.n1751 vdd.n1750 6.98232
R18591 vdd.n3063 vdd.n3062 6.98232
R18592 vdd.n2855 vdd.n2854 6.98232
R18593 vdd.n1255 vdd.t69 6.91577
R18594 vdd.n325 vdd.t60 6.91577
R18595 vdd.n1562 vdd.t32 6.68904
R18596 vdd.n2989 vdd.t57 6.68904
R18597 vdd.n925 vdd.t10 6.46231
R18598 vdd.t34 vdd.n492 6.46231
R18599 vdd.n3168 vdd.n309 6.27748
R18600 vdd.n1556 vdd.n1555 6.27748
R18601 vdd.n2124 vdd.t85 6.00885
R18602 vdd.n2624 vdd.t181 6.00885
R18603 vdd.n861 vdd.t134 5.89549
R18604 vdd.t102 vdd.n679 5.89549
R18605 vdd.n284 vdd.n283 5.81868
R18606 vdd.n233 vdd.n232 5.81868
R18607 vdd.n190 vdd.n189 5.81868
R18608 vdd.n139 vdd.n138 5.81868
R18609 vdd.n97 vdd.n96 5.81868
R18610 vdd.n46 vdd.n45 5.81868
R18611 vdd.n1479 vdd.n1478 5.81868
R18612 vdd.n1530 vdd.n1529 5.81868
R18613 vdd.n1385 vdd.n1384 5.81868
R18614 vdd.n1436 vdd.n1435 5.81868
R18615 vdd.n1292 vdd.n1291 5.81868
R18616 vdd.n1343 vdd.n1342 5.81868
R18617 vdd.t130 vdd.n865 5.78212
R18618 vdd.n1868 vdd.t115 5.78212
R18619 vdd.n2493 vdd.t123 5.78212
R18620 vdd.n674 vdd.t119 5.78212
R18621 vdd.n2252 vdd.n2251 5.77611
R18622 vdd.n1995 vdd.n1865 5.77611
R18623 vdd.n2506 vdd.n2505 5.77611
R18624 vdd.n2710 vdd.n663 5.77611
R18625 vdd.n2776 vdd.n627 5.77611
R18626 vdd.n2416 vdd.n2356 5.77611
R18627 vdd.n2177 vdd.n795 5.77611
R18628 vdd.n1925 vdd.n1924 5.77611
R18629 vdd.n1112 vdd.n1109 5.62474
R18630 vdd.n2047 vdd.n2044 5.62474
R18631 vdd.n3023 vdd.n3020 5.62474
R18632 vdd.n2810 vdd.n2807 5.62474
R18633 vdd.t12 vdd.n817 5.44203
R18634 vdd.n721 vdd.t19 5.44203
R18635 vdd.t16 vdd.n840 5.10193
R18636 vdd.n830 vdd.t38 5.10193
R18637 vdd.t21 vdd.n708 5.10193
R18638 vdd.n698 vdd.t192 5.10193
R18639 vdd.n287 vdd.n278 5.04292
R18640 vdd.n236 vdd.n227 5.04292
R18641 vdd.n193 vdd.n184 5.04292
R18642 vdd.n142 vdd.n133 5.04292
R18643 vdd.n100 vdd.n91 5.04292
R18644 vdd.n49 vdd.n40 5.04292
R18645 vdd.n1482 vdd.n1473 5.04292
R18646 vdd.n1533 vdd.n1524 5.04292
R18647 vdd.n1388 vdd.n1379 5.04292
R18648 vdd.n1439 vdd.n1430 5.04292
R18649 vdd.n1295 vdd.n1286 5.04292
R18650 vdd.n1346 vdd.n1337 5.04292
R18651 vdd.n1588 vdd.t10 4.8752
R18652 vdd.t37 vdd.t207 4.8752
R18653 vdd.t180 vdd.t178 4.8752
R18654 vdd.t80 vdd.t76 4.8752
R18655 vdd.t14 vdd.t175 4.8752
R18656 vdd.n2964 vdd.t34 4.8752
R18657 vdd.n2253 vdd.n2252 4.83952
R18658 vdd.n1865 vdd.n1861 4.83952
R18659 vdd.n2507 vdd.n2506 4.83952
R18660 vdd.n663 vdd.n658 4.83952
R18661 vdd.n627 vdd.n622 4.83952
R18662 vdd.n2413 vdd.n2356 4.83952
R18663 vdd.n2180 vdd.n795 4.83952
R18664 vdd.n1924 vdd.n1923 4.83952
R18665 vdd.n1719 vdd.n893 4.74817
R18666 vdd.n1714 vdd.n894 4.74817
R18667 vdd.n1616 vdd.n1613 4.74817
R18668 vdd.n2028 vdd.n1617 4.74817
R18669 vdd.n2030 vdd.n1616 4.74817
R18670 vdd.n2029 vdd.n2028 4.74817
R18671 vdd.n521 vdd.n519 4.74817
R18672 vdd.n2925 vdd.n522 4.74817
R18673 vdd.n2928 vdd.n522 4.74817
R18674 vdd.n2929 vdd.n521 4.74817
R18675 vdd.n2817 vdd.n606 4.74817
R18676 vdd.n2813 vdd.n608 4.74817
R18677 vdd.n2816 vdd.n608 4.74817
R18678 vdd.n2821 vdd.n606 4.74817
R18679 vdd.n1715 vdd.n893 4.74817
R18680 vdd.n896 vdd.n894 4.74817
R18681 vdd.n309 vdd.n308 4.7074
R18682 vdd.n215 vdd.n214 4.7074
R18683 vdd.n1555 vdd.n1554 4.7074
R18684 vdd.n1461 vdd.n1460 4.7074
R18685 vdd.t32 vdd.n931 4.64847
R18686 vdd.n2980 vdd.t57 4.64847
R18687 vdd.n2130 vdd.t220 4.53511
R18688 vdd.n2618 vdd.t205 4.53511
R18689 vdd.n1264 vdd.t69 4.42174
R18690 vdd.n3162 vdd.t60 4.42174
R18691 vdd.n2162 vdd.t203 4.30838
R18692 vdd.n2588 vdd.t74 4.30838
R18693 vdd.n288 vdd.n276 4.26717
R18694 vdd.n237 vdd.n225 4.26717
R18695 vdd.n194 vdd.n182 4.26717
R18696 vdd.n143 vdd.n131 4.26717
R18697 vdd.n101 vdd.n89 4.26717
R18698 vdd.n50 vdd.n38 4.26717
R18699 vdd.n1483 vdd.n1471 4.26717
R18700 vdd.n1534 vdd.n1522 4.26717
R18701 vdd.n1389 vdd.n1377 4.26717
R18702 vdd.n1440 vdd.n1428 4.26717
R18703 vdd.n1296 vdd.n1284 4.26717
R18704 vdd.n1347 vdd.n1335 4.26717
R18705 vdd.t166 vdd.n959 4.19501
R18706 vdd.t163 vdd.n329 4.19501
R18707 vdd.n309 vdd.n215 4.10845
R18708 vdd.n1555 vdd.n1461 4.10845
R18709 vdd.n265 vdd.t73 4.06363
R18710 vdd.n265 vdd.t195 4.06363
R18711 vdd.n263 vdd.t62 4.06363
R18712 vdd.n263 vdd.t25 4.06363
R18713 vdd.n261 vdd.t191 4.06363
R18714 vdd.n261 vdd.t230 4.06363
R18715 vdd.n259 vdd.t22 4.06363
R18716 vdd.n259 vdd.t65 4.06363
R18717 vdd.n257 vdd.t168 4.06363
R18718 vdd.n257 vdd.t218 4.06363
R18719 vdd.n171 vdd.t226 4.06363
R18720 vdd.n171 vdd.t164 4.06363
R18721 vdd.n169 vdd.t61 4.06363
R18722 vdd.n169 vdd.t59 4.06363
R18723 vdd.n167 vdd.t215 4.06363
R18724 vdd.n167 vdd.t172 4.06363
R18725 vdd.n165 vdd.t1 4.06363
R18726 vdd.n165 vdd.t229 4.06363
R18727 vdd.n163 vdd.t200 4.06363
R18728 vdd.n163 vdd.t214 4.06363
R18729 vdd.n78 vdd.t184 4.06363
R18730 vdd.n78 vdd.t165 4.06363
R18731 vdd.n76 vdd.t68 4.06363
R18732 vdd.n76 vdd.t28 4.06363
R18733 vdd.n74 vdd.t190 4.06363
R18734 vdd.n74 vdd.t64 4.06363
R18735 vdd.n72 vdd.t71 4.06363
R18736 vdd.n72 vdd.t58 4.06363
R18737 vdd.n70 vdd.t35 4.06363
R18738 vdd.n70 vdd.t225 4.06363
R18739 vdd.n1503 vdd.t194 4.06363
R18740 vdd.n1503 vdd.t11 4.06363
R18741 vdd.n1505 vdd.t222 4.06363
R18742 vdd.n1505 vdd.t216 4.06363
R18743 vdd.n1507 vdd.t199 4.06363
R18744 vdd.n1507 vdd.t23 4.06363
R18745 vdd.n1509 vdd.t173 4.06363
R18746 vdd.n1509 vdd.t217 4.06363
R18747 vdd.n1511 vdd.t188 4.06363
R18748 vdd.n1511 vdd.t196 4.06363
R18749 vdd.n1409 vdd.t7 4.06363
R18750 vdd.n1409 vdd.t36 4.06363
R18751 vdd.n1411 vdd.t33 4.06363
R18752 vdd.n1411 vdd.t170 4.06363
R18753 vdd.n1413 vdd.t27 4.06363
R18754 vdd.n1413 vdd.t3 4.06363
R18755 vdd.n1415 vdd.t223 4.06363
R18756 vdd.n1415 vdd.t171 4.06363
R18757 vdd.n1417 vdd.t202 4.06363
R18758 vdd.n1417 vdd.t56 4.06363
R18759 vdd.n1316 vdd.t228 4.06363
R18760 vdd.n1316 vdd.t227 4.06363
R18761 vdd.n1318 vdd.t193 4.06363
R18762 vdd.n1318 vdd.t30 4.06363
R18763 vdd.n1320 vdd.t197 4.06363
R18764 vdd.n1320 vdd.t31 4.06363
R18765 vdd.n1322 vdd.t67 4.06363
R18766 vdd.n1322 vdd.t70 4.06363
R18767 vdd.n1324 vdd.t167 4.06363
R18768 vdd.n1324 vdd.t185 4.06363
R18769 vdd.n26 vdd.t48 3.9605
R18770 vdd.n26 vdd.t47 3.9605
R18771 vdd.n23 vdd.t40 3.9605
R18772 vdd.n23 vdd.t42 3.9605
R18773 vdd.n21 vdd.t54 3.9605
R18774 vdd.n21 vdd.t44 3.9605
R18775 vdd.n20 vdd.t52 3.9605
R18776 vdd.n20 vdd.t39 3.9605
R18777 vdd.n15 vdd.t41 3.9605
R18778 vdd.n15 vdd.t45 3.9605
R18779 vdd.n16 vdd.t51 3.9605
R18780 vdd.n16 vdd.t53 3.9605
R18781 vdd.n18 vdd.t49 3.9605
R18782 vdd.n18 vdd.t50 3.9605
R18783 vdd.n25 vdd.t46 3.9605
R18784 vdd.n25 vdd.t43 3.9605
R18785 vdd.n7 vdd.t15 3.61217
R18786 vdd.n7 vdd.t206 3.61217
R18787 vdd.n8 vdd.t81 3.61217
R18788 vdd.n8 vdd.t20 3.61217
R18789 vdd.n10 vdd.t210 3.61217
R18790 vdd.n10 vdd.t75 3.61217
R18791 vdd.n12 vdd.t78 3.61217
R18792 vdd.n12 vdd.t212 3.61217
R18793 vdd.n5 vdd.t18 3.61217
R18794 vdd.n5 vdd.t177 3.61217
R18795 vdd.n3 vdd.t204 3.61217
R18796 vdd.n3 vdd.t183 3.61217
R18797 vdd.n1 vdd.t13 3.61217
R18798 vdd.n1 vdd.t179 3.61217
R18799 vdd.n0 vdd.t221 3.61217
R18800 vdd.n0 vdd.t208 3.61217
R18801 vdd.n292 vdd.n291 3.49141
R18802 vdd.n241 vdd.n240 3.49141
R18803 vdd.n198 vdd.n197 3.49141
R18804 vdd.n147 vdd.n146 3.49141
R18805 vdd.n105 vdd.n104 3.49141
R18806 vdd.n54 vdd.n53 3.49141
R18807 vdd.n1487 vdd.n1486 3.49141
R18808 vdd.n1538 vdd.n1537 3.49141
R18809 vdd.n1393 vdd.n1392 3.49141
R18810 vdd.n1444 vdd.n1443 3.49141
R18811 vdd.n1300 vdd.n1299 3.49141
R18812 vdd.n1351 vdd.n1350 3.49141
R18813 vdd.n1868 vdd.t203 3.40145
R18814 vdd.n2316 vdd.t17 3.40145
R18815 vdd.n2569 vdd.t211 3.40145
R18816 vdd.n2493 vdd.t74 3.40145
R18817 vdd.n1247 vdd.t55 3.28809
R18818 vdd.t72 vdd.n3154 3.28809
R18819 vdd.n1969 vdd.t220 3.17472
R18820 vdd.n2472 vdd.t205 3.17472
R18821 vdd.n948 vdd.t26 3.06136
R18822 vdd.t63 vdd.n3163 3.06136
R18823 vdd.n1571 vdd.t29 2.83463
R18824 vdd.n2981 vdd.t0 2.83463
R18825 vdd.n295 vdd.n274 2.71565
R18826 vdd.n244 vdd.n223 2.71565
R18827 vdd.n201 vdd.n180 2.71565
R18828 vdd.n150 vdd.n129 2.71565
R18829 vdd.n108 vdd.n87 2.71565
R18830 vdd.n57 vdd.n36 2.71565
R18831 vdd.n1490 vdd.n1469 2.71565
R18832 vdd.n1541 vdd.n1520 2.71565
R18833 vdd.n1396 vdd.n1375 2.71565
R18834 vdd.n1447 vdd.n1426 2.71565
R18835 vdd.n1303 vdd.n1282 2.71565
R18836 vdd.n1354 vdd.n1333 2.71565
R18837 vdd.n1587 vdd.t8 2.6079
R18838 vdd.n2118 vdd.t16 2.6079
R18839 vdd.n2142 vdd.t38 2.6079
R18840 vdd.n2606 vdd.t21 2.6079
R18841 vdd.n2630 vdd.t192 2.6079
R18842 vdd.t82 vdd.n499 2.6079
R18843 vdd.n2636 vdd.n2635 2.49806
R18844 vdd.n2110 vdd.n2109 2.49806
R18845 vdd.n282 vdd.n281 2.4129
R18846 vdd.n231 vdd.n230 2.4129
R18847 vdd.n188 vdd.n187 2.4129
R18848 vdd.n137 vdd.n136 2.4129
R18849 vdd.n95 vdd.n94 2.4129
R18850 vdd.n44 vdd.n43 2.4129
R18851 vdd.n1477 vdd.n1476 2.4129
R18852 vdd.n1528 vdd.n1527 2.4129
R18853 vdd.n1383 vdd.n1382 2.4129
R18854 vdd.n1434 vdd.n1433 2.4129
R18855 vdd.n1290 vdd.n1289 2.4129
R18856 vdd.n1341 vdd.n1340 2.4129
R18857 vdd.n2027 vdd.n1616 2.27742
R18858 vdd.n2028 vdd.n2027 2.27742
R18859 vdd.n2737 vdd.n522 2.27742
R18860 vdd.n2737 vdd.n521 2.27742
R18861 vdd.n2805 vdd.n608 2.27742
R18862 vdd.n2805 vdd.n606 2.27742
R18863 vdd.n2050 vdd.n893 2.27742
R18864 vdd.n2050 vdd.n894 2.27742
R18865 vdd.n2142 vdd.t12 2.2678
R18866 vdd.n2606 vdd.t19 2.2678
R18867 vdd.t178 vdd.n811 2.04107
R18868 vdd.n728 vdd.t80 2.04107
R18869 vdd.n296 vdd.n272 1.93989
R18870 vdd.n245 vdd.n221 1.93989
R18871 vdd.n202 vdd.n178 1.93989
R18872 vdd.n151 vdd.n127 1.93989
R18873 vdd.n109 vdd.n85 1.93989
R18874 vdd.n58 vdd.n34 1.93989
R18875 vdd.n1491 vdd.n1467 1.93989
R18876 vdd.n1542 vdd.n1518 1.93989
R18877 vdd.n1397 vdd.n1373 1.93989
R18878 vdd.n1448 vdd.n1424 1.93989
R18879 vdd.n1304 vdd.n1280 1.93989
R18880 vdd.n1355 vdd.n1331 1.93989
R18881 vdd.n2093 vdd.t130 1.92771
R18882 vdd.n2169 vdd.t115 1.92771
R18883 vdd.n2582 vdd.t123 1.92771
R18884 vdd.n2701 vdd.t119 1.92771
R18885 vdd.n1969 vdd.t85 1.70098
R18886 vdd.n836 vdd.t37 1.70098
R18887 vdd.t175 vdd.n702 1.70098
R18888 vdd.n2472 vdd.t181 1.70098
R18889 vdd.n983 vdd.t98 1.47425
R18890 vdd.t147 vdd.n3139 1.47425
R18891 vdd.n307 vdd.n267 1.16414
R18892 vdd.n300 vdd.n299 1.16414
R18893 vdd.n256 vdd.n216 1.16414
R18894 vdd.n249 vdd.n248 1.16414
R18895 vdd.n213 vdd.n173 1.16414
R18896 vdd.n206 vdd.n205 1.16414
R18897 vdd.n162 vdd.n122 1.16414
R18898 vdd.n155 vdd.n154 1.16414
R18899 vdd.n120 vdd.n80 1.16414
R18900 vdd.n113 vdd.n112 1.16414
R18901 vdd.n69 vdd.n29 1.16414
R18902 vdd.n62 vdd.n61 1.16414
R18903 vdd.n1502 vdd.n1462 1.16414
R18904 vdd.n1495 vdd.n1494 1.16414
R18905 vdd.n1553 vdd.n1513 1.16414
R18906 vdd.n1546 vdd.n1545 1.16414
R18907 vdd.n1408 vdd.n1368 1.16414
R18908 vdd.n1401 vdd.n1400 1.16414
R18909 vdd.n1459 vdd.n1419 1.16414
R18910 vdd.n1452 vdd.n1451 1.16414
R18911 vdd.n1315 vdd.n1275 1.16414
R18912 vdd.n1308 vdd.n1307 1.16414
R18913 vdd.n1366 vdd.n1326 1.16414
R18914 vdd.n1359 vdd.n1358 1.16414
R18915 vdd.n2136 vdd.t207 1.13415
R18916 vdd.n2612 vdd.t14 1.13415
R18917 vdd.n1579 vdd.t6 1.02079
R18918 vdd.t134 vdd.t174 1.02079
R18919 vdd.t79 vdd.t102 1.02079
R18920 vdd.n2972 vdd.t213 1.02079
R18921 vdd.n1113 vdd.n1112 0.970197
R18922 vdd.n2048 vdd.n2047 0.970197
R18923 vdd.n3024 vdd.n3023 0.970197
R18924 vdd.n2812 vdd.n2810 0.970197
R18925 vdd.n1556 vdd.n28 0.800283
R18926 vdd.t2 vdd.n937 0.794056
R18927 vdd.n1606 vdd.t94 0.794056
R18928 vdd.n2112 vdd.t174 0.794056
R18929 vdd.n2148 vdd.t180 0.794056
R18930 vdd.n2600 vdd.t76 0.794056
R18931 vdd.n2638 vdd.t79 0.794056
R18932 vdd.t87 vdd.n511 0.794056
R18933 vdd.n481 vdd.t189 0.794056
R18934 vdd vdd.n3168 0.79245
R18935 vdd.n1256 vdd.t66 0.567326
R18936 vdd.n3156 vdd.t24 0.567326
R18937 vdd.n2038 vdd.n2037 0.509646
R18938 vdd.n2937 vdd.n2936 0.509646
R18939 vdd.n3135 vdd.n3134 0.509646
R18940 vdd.n3017 vdd.n3016 0.509646
R18941 vdd.n2943 vdd.n514 0.509646
R18942 vdd.n1601 vdd.n895 0.509646
R18943 vdd.n1218 vdd.n980 0.509646
R18944 vdd.n1212 vdd.n1211 0.509646
R18945 vdd.n4 vdd.n2 0.459552
R18946 vdd.n11 vdd.n9 0.459552
R18947 vdd.n305 vdd.n304 0.388379
R18948 vdd.n271 vdd.n269 0.388379
R18949 vdd.n254 vdd.n253 0.388379
R18950 vdd.n220 vdd.n218 0.388379
R18951 vdd.n211 vdd.n210 0.388379
R18952 vdd.n177 vdd.n175 0.388379
R18953 vdd.n160 vdd.n159 0.388379
R18954 vdd.n126 vdd.n124 0.388379
R18955 vdd.n118 vdd.n117 0.388379
R18956 vdd.n84 vdd.n82 0.388379
R18957 vdd.n67 vdd.n66 0.388379
R18958 vdd.n33 vdd.n31 0.388379
R18959 vdd.n1500 vdd.n1499 0.388379
R18960 vdd.n1466 vdd.n1464 0.388379
R18961 vdd.n1551 vdd.n1550 0.388379
R18962 vdd.n1517 vdd.n1515 0.388379
R18963 vdd.n1406 vdd.n1405 0.388379
R18964 vdd.n1372 vdd.n1370 0.388379
R18965 vdd.n1457 vdd.n1456 0.388379
R18966 vdd.n1423 vdd.n1421 0.388379
R18967 vdd.n1313 vdd.n1312 0.388379
R18968 vdd.n1279 vdd.n1277 0.388379
R18969 vdd.n1364 vdd.n1363 0.388379
R18970 vdd.n1330 vdd.n1328 0.388379
R18971 vdd.n19 vdd.n17 0.387128
R18972 vdd.n24 vdd.n22 0.387128
R18973 vdd.n6 vdd.n4 0.358259
R18974 vdd.n13 vdd.n11 0.358259
R18975 vdd.n260 vdd.n258 0.358259
R18976 vdd.n262 vdd.n260 0.358259
R18977 vdd.n264 vdd.n262 0.358259
R18978 vdd.n266 vdd.n264 0.358259
R18979 vdd.n308 vdd.n266 0.358259
R18980 vdd.n166 vdd.n164 0.358259
R18981 vdd.n168 vdd.n166 0.358259
R18982 vdd.n170 vdd.n168 0.358259
R18983 vdd.n172 vdd.n170 0.358259
R18984 vdd.n214 vdd.n172 0.358259
R18985 vdd.n73 vdd.n71 0.358259
R18986 vdd.n75 vdd.n73 0.358259
R18987 vdd.n77 vdd.n75 0.358259
R18988 vdd.n79 vdd.n77 0.358259
R18989 vdd.n121 vdd.n79 0.358259
R18990 vdd.n1554 vdd.n1512 0.358259
R18991 vdd.n1512 vdd.n1510 0.358259
R18992 vdd.n1510 vdd.n1508 0.358259
R18993 vdd.n1508 vdd.n1506 0.358259
R18994 vdd.n1506 vdd.n1504 0.358259
R18995 vdd.n1460 vdd.n1418 0.358259
R18996 vdd.n1418 vdd.n1416 0.358259
R18997 vdd.n1416 vdd.n1414 0.358259
R18998 vdd.n1414 vdd.n1412 0.358259
R18999 vdd.n1412 vdd.n1410 0.358259
R19000 vdd.n1367 vdd.n1325 0.358259
R19001 vdd.n1325 vdd.n1323 0.358259
R19002 vdd.n1323 vdd.n1321 0.358259
R19003 vdd.n1321 vdd.n1319 0.358259
R19004 vdd.n1319 vdd.n1317 0.358259
R19005 vdd.t186 vdd.n966 0.340595
R19006 vdd.n3147 vdd.t4 0.340595
R19007 vdd.n14 vdd.n6 0.334552
R19008 vdd.n14 vdd.n13 0.334552
R19009 vdd.n27 vdd.n19 0.21707
R19010 vdd.n27 vdd.n24 0.21707
R19011 vdd.n306 vdd.n268 0.155672
R19012 vdd.n298 vdd.n268 0.155672
R19013 vdd.n298 vdd.n297 0.155672
R19014 vdd.n297 vdd.n273 0.155672
R19015 vdd.n290 vdd.n273 0.155672
R19016 vdd.n290 vdd.n289 0.155672
R19017 vdd.n289 vdd.n277 0.155672
R19018 vdd.n282 vdd.n277 0.155672
R19019 vdd.n255 vdd.n217 0.155672
R19020 vdd.n247 vdd.n217 0.155672
R19021 vdd.n247 vdd.n246 0.155672
R19022 vdd.n246 vdd.n222 0.155672
R19023 vdd.n239 vdd.n222 0.155672
R19024 vdd.n239 vdd.n238 0.155672
R19025 vdd.n238 vdd.n226 0.155672
R19026 vdd.n231 vdd.n226 0.155672
R19027 vdd.n212 vdd.n174 0.155672
R19028 vdd.n204 vdd.n174 0.155672
R19029 vdd.n204 vdd.n203 0.155672
R19030 vdd.n203 vdd.n179 0.155672
R19031 vdd.n196 vdd.n179 0.155672
R19032 vdd.n196 vdd.n195 0.155672
R19033 vdd.n195 vdd.n183 0.155672
R19034 vdd.n188 vdd.n183 0.155672
R19035 vdd.n161 vdd.n123 0.155672
R19036 vdd.n153 vdd.n123 0.155672
R19037 vdd.n153 vdd.n152 0.155672
R19038 vdd.n152 vdd.n128 0.155672
R19039 vdd.n145 vdd.n128 0.155672
R19040 vdd.n145 vdd.n144 0.155672
R19041 vdd.n144 vdd.n132 0.155672
R19042 vdd.n137 vdd.n132 0.155672
R19043 vdd.n119 vdd.n81 0.155672
R19044 vdd.n111 vdd.n81 0.155672
R19045 vdd.n111 vdd.n110 0.155672
R19046 vdd.n110 vdd.n86 0.155672
R19047 vdd.n103 vdd.n86 0.155672
R19048 vdd.n103 vdd.n102 0.155672
R19049 vdd.n102 vdd.n90 0.155672
R19050 vdd.n95 vdd.n90 0.155672
R19051 vdd.n68 vdd.n30 0.155672
R19052 vdd.n60 vdd.n30 0.155672
R19053 vdd.n60 vdd.n59 0.155672
R19054 vdd.n59 vdd.n35 0.155672
R19055 vdd.n52 vdd.n35 0.155672
R19056 vdd.n52 vdd.n51 0.155672
R19057 vdd.n51 vdd.n39 0.155672
R19058 vdd.n44 vdd.n39 0.155672
R19059 vdd.n1501 vdd.n1463 0.155672
R19060 vdd.n1493 vdd.n1463 0.155672
R19061 vdd.n1493 vdd.n1492 0.155672
R19062 vdd.n1492 vdd.n1468 0.155672
R19063 vdd.n1485 vdd.n1468 0.155672
R19064 vdd.n1485 vdd.n1484 0.155672
R19065 vdd.n1484 vdd.n1472 0.155672
R19066 vdd.n1477 vdd.n1472 0.155672
R19067 vdd.n1552 vdd.n1514 0.155672
R19068 vdd.n1544 vdd.n1514 0.155672
R19069 vdd.n1544 vdd.n1543 0.155672
R19070 vdd.n1543 vdd.n1519 0.155672
R19071 vdd.n1536 vdd.n1519 0.155672
R19072 vdd.n1536 vdd.n1535 0.155672
R19073 vdd.n1535 vdd.n1523 0.155672
R19074 vdd.n1528 vdd.n1523 0.155672
R19075 vdd.n1407 vdd.n1369 0.155672
R19076 vdd.n1399 vdd.n1369 0.155672
R19077 vdd.n1399 vdd.n1398 0.155672
R19078 vdd.n1398 vdd.n1374 0.155672
R19079 vdd.n1391 vdd.n1374 0.155672
R19080 vdd.n1391 vdd.n1390 0.155672
R19081 vdd.n1390 vdd.n1378 0.155672
R19082 vdd.n1383 vdd.n1378 0.155672
R19083 vdd.n1458 vdd.n1420 0.155672
R19084 vdd.n1450 vdd.n1420 0.155672
R19085 vdd.n1450 vdd.n1449 0.155672
R19086 vdd.n1449 vdd.n1425 0.155672
R19087 vdd.n1442 vdd.n1425 0.155672
R19088 vdd.n1442 vdd.n1441 0.155672
R19089 vdd.n1441 vdd.n1429 0.155672
R19090 vdd.n1434 vdd.n1429 0.155672
R19091 vdd.n1314 vdd.n1276 0.155672
R19092 vdd.n1306 vdd.n1276 0.155672
R19093 vdd.n1306 vdd.n1305 0.155672
R19094 vdd.n1305 vdd.n1281 0.155672
R19095 vdd.n1298 vdd.n1281 0.155672
R19096 vdd.n1298 vdd.n1297 0.155672
R19097 vdd.n1297 vdd.n1285 0.155672
R19098 vdd.n1290 vdd.n1285 0.155672
R19099 vdd.n1365 vdd.n1327 0.155672
R19100 vdd.n1357 vdd.n1327 0.155672
R19101 vdd.n1357 vdd.n1356 0.155672
R19102 vdd.n1356 vdd.n1332 0.155672
R19103 vdd.n1349 vdd.n1332 0.155672
R19104 vdd.n1349 vdd.n1348 0.155672
R19105 vdd.n1348 vdd.n1336 0.155672
R19106 vdd.n1341 vdd.n1336 0.155672
R19107 vdd.n1813 vdd.n1618 0.152939
R19108 vdd.n1624 vdd.n1618 0.152939
R19109 vdd.n1625 vdd.n1624 0.152939
R19110 vdd.n1626 vdd.n1625 0.152939
R19111 vdd.n1627 vdd.n1626 0.152939
R19112 vdd.n1631 vdd.n1627 0.152939
R19113 vdd.n1632 vdd.n1631 0.152939
R19114 vdd.n1633 vdd.n1632 0.152939
R19115 vdd.n1634 vdd.n1633 0.152939
R19116 vdd.n1638 vdd.n1634 0.152939
R19117 vdd.n1639 vdd.n1638 0.152939
R19118 vdd.n1640 vdd.n1639 0.152939
R19119 vdd.n1788 vdd.n1640 0.152939
R19120 vdd.n1788 vdd.n1787 0.152939
R19121 vdd.n1787 vdd.n1786 0.152939
R19122 vdd.n1786 vdd.n1646 0.152939
R19123 vdd.n1651 vdd.n1646 0.152939
R19124 vdd.n1652 vdd.n1651 0.152939
R19125 vdd.n1653 vdd.n1652 0.152939
R19126 vdd.n1657 vdd.n1653 0.152939
R19127 vdd.n1658 vdd.n1657 0.152939
R19128 vdd.n1659 vdd.n1658 0.152939
R19129 vdd.n1660 vdd.n1659 0.152939
R19130 vdd.n1664 vdd.n1660 0.152939
R19131 vdd.n1665 vdd.n1664 0.152939
R19132 vdd.n1666 vdd.n1665 0.152939
R19133 vdd.n1667 vdd.n1666 0.152939
R19134 vdd.n1671 vdd.n1667 0.152939
R19135 vdd.n1672 vdd.n1671 0.152939
R19136 vdd.n1673 vdd.n1672 0.152939
R19137 vdd.n1674 vdd.n1673 0.152939
R19138 vdd.n1678 vdd.n1674 0.152939
R19139 vdd.n1679 vdd.n1678 0.152939
R19140 vdd.n1680 vdd.n1679 0.152939
R19141 vdd.n1749 vdd.n1680 0.152939
R19142 vdd.n1749 vdd.n1748 0.152939
R19143 vdd.n1748 vdd.n1747 0.152939
R19144 vdd.n1747 vdd.n1686 0.152939
R19145 vdd.n1691 vdd.n1686 0.152939
R19146 vdd.n1692 vdd.n1691 0.152939
R19147 vdd.n1693 vdd.n1692 0.152939
R19148 vdd.n1697 vdd.n1693 0.152939
R19149 vdd.n1698 vdd.n1697 0.152939
R19150 vdd.n1699 vdd.n1698 0.152939
R19151 vdd.n1700 vdd.n1699 0.152939
R19152 vdd.n1704 vdd.n1700 0.152939
R19153 vdd.n1705 vdd.n1704 0.152939
R19154 vdd.n1706 vdd.n1705 0.152939
R19155 vdd.n1707 vdd.n1706 0.152939
R19156 vdd.n1708 vdd.n1707 0.152939
R19157 vdd.n1708 vdd.n892 0.152939
R19158 vdd.n2037 vdd.n1612 0.152939
R19159 vdd.n1559 vdd.n1558 0.152939
R19160 vdd.n1559 vdd.n928 0.152939
R19161 vdd.n1574 vdd.n928 0.152939
R19162 vdd.n1575 vdd.n1574 0.152939
R19163 vdd.n1576 vdd.n1575 0.152939
R19164 vdd.n1576 vdd.n917 0.152939
R19165 vdd.n1591 vdd.n917 0.152939
R19166 vdd.n1592 vdd.n1591 0.152939
R19167 vdd.n1593 vdd.n1592 0.152939
R19168 vdd.n1593 vdd.n905 0.152939
R19169 vdd.n1610 vdd.n905 0.152939
R19170 vdd.n1611 vdd.n1610 0.152939
R19171 vdd.n2038 vdd.n1611 0.152939
R19172 vdd.n527 vdd.n524 0.152939
R19173 vdd.n528 vdd.n527 0.152939
R19174 vdd.n529 vdd.n528 0.152939
R19175 vdd.n530 vdd.n529 0.152939
R19176 vdd.n533 vdd.n530 0.152939
R19177 vdd.n534 vdd.n533 0.152939
R19178 vdd.n535 vdd.n534 0.152939
R19179 vdd.n536 vdd.n535 0.152939
R19180 vdd.n539 vdd.n536 0.152939
R19181 vdd.n540 vdd.n539 0.152939
R19182 vdd.n541 vdd.n540 0.152939
R19183 vdd.n542 vdd.n541 0.152939
R19184 vdd.n547 vdd.n542 0.152939
R19185 vdd.n548 vdd.n547 0.152939
R19186 vdd.n549 vdd.n548 0.152939
R19187 vdd.n550 vdd.n549 0.152939
R19188 vdd.n553 vdd.n550 0.152939
R19189 vdd.n554 vdd.n553 0.152939
R19190 vdd.n555 vdd.n554 0.152939
R19191 vdd.n556 vdd.n555 0.152939
R19192 vdd.n559 vdd.n556 0.152939
R19193 vdd.n560 vdd.n559 0.152939
R19194 vdd.n561 vdd.n560 0.152939
R19195 vdd.n562 vdd.n561 0.152939
R19196 vdd.n565 vdd.n562 0.152939
R19197 vdd.n566 vdd.n565 0.152939
R19198 vdd.n567 vdd.n566 0.152939
R19199 vdd.n568 vdd.n567 0.152939
R19200 vdd.n571 vdd.n568 0.152939
R19201 vdd.n572 vdd.n571 0.152939
R19202 vdd.n573 vdd.n572 0.152939
R19203 vdd.n574 vdd.n573 0.152939
R19204 vdd.n577 vdd.n574 0.152939
R19205 vdd.n578 vdd.n577 0.152939
R19206 vdd.n2853 vdd.n578 0.152939
R19207 vdd.n2853 vdd.n2852 0.152939
R19208 vdd.n2852 vdd.n2851 0.152939
R19209 vdd.n2851 vdd.n582 0.152939
R19210 vdd.n587 vdd.n582 0.152939
R19211 vdd.n588 vdd.n587 0.152939
R19212 vdd.n591 vdd.n588 0.152939
R19213 vdd.n592 vdd.n591 0.152939
R19214 vdd.n593 vdd.n592 0.152939
R19215 vdd.n594 vdd.n593 0.152939
R19216 vdd.n597 vdd.n594 0.152939
R19217 vdd.n598 vdd.n597 0.152939
R19218 vdd.n599 vdd.n598 0.152939
R19219 vdd.n600 vdd.n599 0.152939
R19220 vdd.n603 vdd.n600 0.152939
R19221 vdd.n604 vdd.n603 0.152939
R19222 vdd.n605 vdd.n604 0.152939
R19223 vdd.n2936 vdd.n518 0.152939
R19224 vdd.n2937 vdd.n508 0.152939
R19225 vdd.n2951 vdd.n508 0.152939
R19226 vdd.n2952 vdd.n2951 0.152939
R19227 vdd.n2953 vdd.n2952 0.152939
R19228 vdd.n2953 vdd.n496 0.152939
R19229 vdd.n2967 vdd.n496 0.152939
R19230 vdd.n2968 vdd.n2967 0.152939
R19231 vdd.n2969 vdd.n2968 0.152939
R19232 vdd.n2969 vdd.n484 0.152939
R19233 vdd.n2984 vdd.n484 0.152939
R19234 vdd.n2985 vdd.n2984 0.152939
R19235 vdd.n2986 vdd.n2985 0.152939
R19236 vdd.n2986 vdd.n310 0.152939
R19237 vdd.n320 vdd.n311 0.152939
R19238 vdd.n321 vdd.n320 0.152939
R19239 vdd.n322 vdd.n321 0.152939
R19240 vdd.n331 vdd.n322 0.152939
R19241 vdd.n332 vdd.n331 0.152939
R19242 vdd.n333 vdd.n332 0.152939
R19243 vdd.n334 vdd.n333 0.152939
R19244 vdd.n342 vdd.n334 0.152939
R19245 vdd.n343 vdd.n342 0.152939
R19246 vdd.n344 vdd.n343 0.152939
R19247 vdd.n345 vdd.n344 0.152939
R19248 vdd.n353 vdd.n345 0.152939
R19249 vdd.n3135 vdd.n353 0.152939
R19250 vdd.n3134 vdd.n354 0.152939
R19251 vdd.n357 vdd.n354 0.152939
R19252 vdd.n361 vdd.n357 0.152939
R19253 vdd.n362 vdd.n361 0.152939
R19254 vdd.n363 vdd.n362 0.152939
R19255 vdd.n364 vdd.n363 0.152939
R19256 vdd.n365 vdd.n364 0.152939
R19257 vdd.n369 vdd.n365 0.152939
R19258 vdd.n370 vdd.n369 0.152939
R19259 vdd.n371 vdd.n370 0.152939
R19260 vdd.n372 vdd.n371 0.152939
R19261 vdd.n376 vdd.n372 0.152939
R19262 vdd.n377 vdd.n376 0.152939
R19263 vdd.n378 vdd.n377 0.152939
R19264 vdd.n379 vdd.n378 0.152939
R19265 vdd.n383 vdd.n379 0.152939
R19266 vdd.n384 vdd.n383 0.152939
R19267 vdd.n385 vdd.n384 0.152939
R19268 vdd.n3100 vdd.n385 0.152939
R19269 vdd.n3100 vdd.n3099 0.152939
R19270 vdd.n3099 vdd.n3098 0.152939
R19271 vdd.n3098 vdd.n391 0.152939
R19272 vdd.n396 vdd.n391 0.152939
R19273 vdd.n397 vdd.n396 0.152939
R19274 vdd.n398 vdd.n397 0.152939
R19275 vdd.n402 vdd.n398 0.152939
R19276 vdd.n403 vdd.n402 0.152939
R19277 vdd.n404 vdd.n403 0.152939
R19278 vdd.n405 vdd.n404 0.152939
R19279 vdd.n409 vdd.n405 0.152939
R19280 vdd.n410 vdd.n409 0.152939
R19281 vdd.n411 vdd.n410 0.152939
R19282 vdd.n412 vdd.n411 0.152939
R19283 vdd.n416 vdd.n412 0.152939
R19284 vdd.n417 vdd.n416 0.152939
R19285 vdd.n418 vdd.n417 0.152939
R19286 vdd.n419 vdd.n418 0.152939
R19287 vdd.n423 vdd.n419 0.152939
R19288 vdd.n424 vdd.n423 0.152939
R19289 vdd.n425 vdd.n424 0.152939
R19290 vdd.n3061 vdd.n425 0.152939
R19291 vdd.n3061 vdd.n3060 0.152939
R19292 vdd.n3060 vdd.n3059 0.152939
R19293 vdd.n3059 vdd.n431 0.152939
R19294 vdd.n436 vdd.n431 0.152939
R19295 vdd.n437 vdd.n436 0.152939
R19296 vdd.n438 vdd.n437 0.152939
R19297 vdd.n442 vdd.n438 0.152939
R19298 vdd.n443 vdd.n442 0.152939
R19299 vdd.n444 vdd.n443 0.152939
R19300 vdd.n445 vdd.n444 0.152939
R19301 vdd.n449 vdd.n445 0.152939
R19302 vdd.n450 vdd.n449 0.152939
R19303 vdd.n451 vdd.n450 0.152939
R19304 vdd.n452 vdd.n451 0.152939
R19305 vdd.n456 vdd.n452 0.152939
R19306 vdd.n457 vdd.n456 0.152939
R19307 vdd.n458 vdd.n457 0.152939
R19308 vdd.n459 vdd.n458 0.152939
R19309 vdd.n463 vdd.n459 0.152939
R19310 vdd.n464 vdd.n463 0.152939
R19311 vdd.n465 vdd.n464 0.152939
R19312 vdd.n3017 vdd.n465 0.152939
R19313 vdd.n2944 vdd.n2943 0.152939
R19314 vdd.n2945 vdd.n2944 0.152939
R19315 vdd.n2945 vdd.n502 0.152939
R19316 vdd.n2959 vdd.n502 0.152939
R19317 vdd.n2960 vdd.n2959 0.152939
R19318 vdd.n2961 vdd.n2960 0.152939
R19319 vdd.n2961 vdd.n489 0.152939
R19320 vdd.n2975 vdd.n489 0.152939
R19321 vdd.n2976 vdd.n2975 0.152939
R19322 vdd.n2977 vdd.n2976 0.152939
R19323 vdd.n2977 vdd.n477 0.152939
R19324 vdd.n2992 vdd.n477 0.152939
R19325 vdd.n2993 vdd.n2992 0.152939
R19326 vdd.n2994 vdd.n2993 0.152939
R19327 vdd.n2994 vdd.n475 0.152939
R19328 vdd.n2998 vdd.n475 0.152939
R19329 vdd.n2999 vdd.n2998 0.152939
R19330 vdd.n3000 vdd.n2999 0.152939
R19331 vdd.n3000 vdd.n472 0.152939
R19332 vdd.n3004 vdd.n472 0.152939
R19333 vdd.n3005 vdd.n3004 0.152939
R19334 vdd.n3006 vdd.n3005 0.152939
R19335 vdd.n3006 vdd.n469 0.152939
R19336 vdd.n3010 vdd.n469 0.152939
R19337 vdd.n3011 vdd.n3010 0.152939
R19338 vdd.n3012 vdd.n3011 0.152939
R19339 vdd.n3012 vdd.n466 0.152939
R19340 vdd.n3016 vdd.n466 0.152939
R19341 vdd.n2806 vdd.n514 0.152939
R19342 vdd.n2049 vdd.n895 0.152939
R19343 vdd.n1219 vdd.n1218 0.152939
R19344 vdd.n1220 vdd.n1219 0.152939
R19345 vdd.n1220 vdd.n969 0.152939
R19346 vdd.n1234 vdd.n969 0.152939
R19347 vdd.n1235 vdd.n1234 0.152939
R19348 vdd.n1236 vdd.n1235 0.152939
R19349 vdd.n1236 vdd.n956 0.152939
R19350 vdd.n1250 vdd.n956 0.152939
R19351 vdd.n1251 vdd.n1250 0.152939
R19352 vdd.n1252 vdd.n1251 0.152939
R19353 vdd.n1252 vdd.n945 0.152939
R19354 vdd.n1267 vdd.n945 0.152939
R19355 vdd.n1268 vdd.n1267 0.152939
R19356 vdd.n1269 vdd.n1268 0.152939
R19357 vdd.n1269 vdd.n934 0.152939
R19358 vdd.n1565 vdd.n934 0.152939
R19359 vdd.n1566 vdd.n1565 0.152939
R19360 vdd.n1567 vdd.n1566 0.152939
R19361 vdd.n1567 vdd.n922 0.152939
R19362 vdd.n1582 vdd.n922 0.152939
R19363 vdd.n1583 vdd.n1582 0.152939
R19364 vdd.n1584 vdd.n1583 0.152939
R19365 vdd.n1584 vdd.n912 0.152939
R19366 vdd.n1599 vdd.n912 0.152939
R19367 vdd.n1600 vdd.n1599 0.152939
R19368 vdd.n1603 vdd.n1600 0.152939
R19369 vdd.n1603 vdd.n1602 0.152939
R19370 vdd.n1602 vdd.n1601 0.152939
R19371 vdd.n1211 vdd.n985 0.152939
R19372 vdd.n1207 vdd.n985 0.152939
R19373 vdd.n1207 vdd.n1206 0.152939
R19374 vdd.n1206 vdd.n1205 0.152939
R19375 vdd.n1205 vdd.n990 0.152939
R19376 vdd.n1201 vdd.n990 0.152939
R19377 vdd.n1201 vdd.n1200 0.152939
R19378 vdd.n1200 vdd.n1199 0.152939
R19379 vdd.n1199 vdd.n998 0.152939
R19380 vdd.n1195 vdd.n998 0.152939
R19381 vdd.n1195 vdd.n1194 0.152939
R19382 vdd.n1194 vdd.n1193 0.152939
R19383 vdd.n1193 vdd.n1006 0.152939
R19384 vdd.n1189 vdd.n1006 0.152939
R19385 vdd.n1189 vdd.n1188 0.152939
R19386 vdd.n1188 vdd.n1187 0.152939
R19387 vdd.n1187 vdd.n1014 0.152939
R19388 vdd.n1183 vdd.n1014 0.152939
R19389 vdd.n1183 vdd.n1182 0.152939
R19390 vdd.n1182 vdd.n1181 0.152939
R19391 vdd.n1181 vdd.n1024 0.152939
R19392 vdd.n1177 vdd.n1024 0.152939
R19393 vdd.n1177 vdd.n1176 0.152939
R19394 vdd.n1176 vdd.n1175 0.152939
R19395 vdd.n1175 vdd.n1032 0.152939
R19396 vdd.n1171 vdd.n1032 0.152939
R19397 vdd.n1171 vdd.n1170 0.152939
R19398 vdd.n1170 vdd.n1169 0.152939
R19399 vdd.n1169 vdd.n1040 0.152939
R19400 vdd.n1165 vdd.n1040 0.152939
R19401 vdd.n1165 vdd.n1164 0.152939
R19402 vdd.n1164 vdd.n1163 0.152939
R19403 vdd.n1163 vdd.n1048 0.152939
R19404 vdd.n1159 vdd.n1048 0.152939
R19405 vdd.n1159 vdd.n1158 0.152939
R19406 vdd.n1158 vdd.n1157 0.152939
R19407 vdd.n1157 vdd.n1056 0.152939
R19408 vdd.n1153 vdd.n1056 0.152939
R19409 vdd.n1153 vdd.n1152 0.152939
R19410 vdd.n1152 vdd.n1151 0.152939
R19411 vdd.n1151 vdd.n1064 0.152939
R19412 vdd.n1071 vdd.n1064 0.152939
R19413 vdd.n1141 vdd.n1071 0.152939
R19414 vdd.n1141 vdd.n1140 0.152939
R19415 vdd.n1140 vdd.n1139 0.152939
R19416 vdd.n1139 vdd.n1072 0.152939
R19417 vdd.n1135 vdd.n1072 0.152939
R19418 vdd.n1135 vdd.n1134 0.152939
R19419 vdd.n1134 vdd.n1133 0.152939
R19420 vdd.n1133 vdd.n1079 0.152939
R19421 vdd.n1129 vdd.n1079 0.152939
R19422 vdd.n1129 vdd.n1128 0.152939
R19423 vdd.n1128 vdd.n1127 0.152939
R19424 vdd.n1127 vdd.n1087 0.152939
R19425 vdd.n1123 vdd.n1087 0.152939
R19426 vdd.n1123 vdd.n1122 0.152939
R19427 vdd.n1122 vdd.n1121 0.152939
R19428 vdd.n1121 vdd.n1095 0.152939
R19429 vdd.n1117 vdd.n1095 0.152939
R19430 vdd.n1117 vdd.n1116 0.152939
R19431 vdd.n1116 vdd.n1115 0.152939
R19432 vdd.n1115 vdd.n1103 0.152939
R19433 vdd.n1103 vdd.n980 0.152939
R19434 vdd.n1212 vdd.n975 0.152939
R19435 vdd.n1226 vdd.n975 0.152939
R19436 vdd.n1227 vdd.n1226 0.152939
R19437 vdd.n1228 vdd.n1227 0.152939
R19438 vdd.n1228 vdd.n963 0.152939
R19439 vdd.n1242 vdd.n963 0.152939
R19440 vdd.n1243 vdd.n1242 0.152939
R19441 vdd.n1244 vdd.n1243 0.152939
R19442 vdd.n1244 vdd.n951 0.152939
R19443 vdd.n1259 vdd.n951 0.152939
R19444 vdd.n1260 vdd.n1259 0.152939
R19445 vdd.n1261 vdd.n1260 0.152939
R19446 vdd.n1261 vdd.n940 0.152939
R19447 vdd.n1558 vdd.n1557 0.145814
R19448 vdd.n3167 vdd.n310 0.145814
R19449 vdd.n3167 vdd.n311 0.145814
R19450 vdd.n1557 vdd.n940 0.145814
R19451 vdd.n2027 vdd.n1612 0.110256
R19452 vdd.n2737 vdd.n518 0.110256
R19453 vdd.n2806 vdd.n2805 0.110256
R19454 vdd.n2050 vdd.n2049 0.110256
R19455 vdd.n2027 vdd.n1813 0.0431829
R19456 vdd.n2050 vdd.n892 0.0431829
R19457 vdd.n2737 vdd.n524 0.0431829
R19458 vdd.n2805 vdd.n605 0.0431829
R19459 vdd vdd.n28 0.00833333
R19460 a_n6308_8799.n138 a_n6308_8799.t83 490.524
R19461 a_n6308_8799.n149 a_n6308_8799.t90 490.524
R19462 a_n6308_8799.n161 a_n6308_8799.t100 490.524
R19463 a_n6308_8799.n104 a_n6308_8799.t60 490.524
R19464 a_n6308_8799.n115 a_n6308_8799.t66 490.524
R19465 a_n6308_8799.n127 a_n6308_8799.t99 490.524
R19466 a_n6308_8799.n30 a_n6308_8799.t69 484.3
R19467 a_n6308_8799.n144 a_n6308_8799.t68 464.166
R19468 a_n6308_8799.n143 a_n6308_8799.t50 464.166
R19469 a_n6308_8799.n134 a_n6308_8799.t96 464.166
R19470 a_n6308_8799.n142 a_n6308_8799.t70 464.166
R19471 a_n6308_8799.n141 a_n6308_8799.t55 464.166
R19472 a_n6308_8799.n135 a_n6308_8799.t98 464.166
R19473 a_n6308_8799.n140 a_n6308_8799.t80 464.166
R19474 a_n6308_8799.n139 a_n6308_8799.t78 464.166
R19475 a_n6308_8799.n136 a_n6308_8799.t39 464.166
R19476 a_n6308_8799.n137 a_n6308_8799.t84 464.166
R19477 a_n6308_8799.n39 a_n6308_8799.t74 484.3
R19478 a_n6308_8799.n155 a_n6308_8799.t73 464.166
R19479 a_n6308_8799.n154 a_n6308_8799.t62 464.166
R19480 a_n6308_8799.n145 a_n6308_8799.t104 464.166
R19481 a_n6308_8799.n153 a_n6308_8799.t77 464.166
R19482 a_n6308_8799.n152 a_n6308_8799.t63 464.166
R19483 a_n6308_8799.n146 a_n6308_8799.t36 464.166
R19484 a_n6308_8799.n151 a_n6308_8799.t89 464.166
R19485 a_n6308_8799.n150 a_n6308_8799.t88 464.166
R19486 a_n6308_8799.n147 a_n6308_8799.t46 464.166
R19487 a_n6308_8799.n148 a_n6308_8799.t91 464.166
R19488 a_n6308_8799.n48 a_n6308_8799.t106 484.3
R19489 a_n6308_8799.n167 a_n6308_8799.t48 464.166
R19490 a_n6308_8799.n166 a_n6308_8799.t75 464.166
R19491 a_n6308_8799.n157 a_n6308_8799.t38 464.166
R19492 a_n6308_8799.n165 a_n6308_8799.t93 464.166
R19493 a_n6308_8799.n164 a_n6308_8799.t54 464.166
R19494 a_n6308_8799.n158 a_n6308_8799.t81 464.166
R19495 a_n6308_8799.n163 a_n6308_8799.t40 464.166
R19496 a_n6308_8799.n162 a_n6308_8799.t58 464.166
R19497 a_n6308_8799.n159 a_n6308_8799.t102 464.166
R19498 a_n6308_8799.n160 a_n6308_8799.t86 464.166
R19499 a_n6308_8799.n103 a_n6308_8799.t61 464.166
R19500 a_n6308_8799.n102 a_n6308_8799.t85 464.166
R19501 a_n6308_8799.n105 a_n6308_8799.t37 464.166
R19502 a_n6308_8799.n101 a_n6308_8799.t57 464.166
R19503 a_n6308_8799.n106 a_n6308_8799.t72 464.166
R19504 a_n6308_8799.n107 a_n6308_8799.t97 464.166
R19505 a_n6308_8799.n100 a_n6308_8799.t44 464.166
R19506 a_n6308_8799.n108 a_n6308_8799.t56 464.166
R19507 a_n6308_8799.n99 a_n6308_8799.t95 464.166
R19508 a_n6308_8799.n109 a_n6308_8799.t43 464.166
R19509 a_n6308_8799.n114 a_n6308_8799.t67 464.166
R19510 a_n6308_8799.n113 a_n6308_8799.t92 464.166
R19511 a_n6308_8799.n116 a_n6308_8799.t45 464.166
R19512 a_n6308_8799.n112 a_n6308_8799.t65 464.166
R19513 a_n6308_8799.n117 a_n6308_8799.t79 464.166
R19514 a_n6308_8799.n118 a_n6308_8799.t105 464.166
R19515 a_n6308_8799.n111 a_n6308_8799.t53 464.166
R19516 a_n6308_8799.n119 a_n6308_8799.t64 464.166
R19517 a_n6308_8799.n110 a_n6308_8799.t101 464.166
R19518 a_n6308_8799.n120 a_n6308_8799.t49 464.166
R19519 a_n6308_8799.n126 a_n6308_8799.t87 464.166
R19520 a_n6308_8799.n125 a_n6308_8799.t103 464.166
R19521 a_n6308_8799.n128 a_n6308_8799.t71 464.166
R19522 a_n6308_8799.n124 a_n6308_8799.t41 464.166
R19523 a_n6308_8799.n129 a_n6308_8799.t82 464.166
R19524 a_n6308_8799.n130 a_n6308_8799.t52 464.166
R19525 a_n6308_8799.n123 a_n6308_8799.t94 464.166
R19526 a_n6308_8799.n131 a_n6308_8799.t59 464.166
R19527 a_n6308_8799.n122 a_n6308_8799.t76 464.166
R19528 a_n6308_8799.n132 a_n6308_8799.t47 464.166
R19529 a_n6308_8799.n38 a_n6308_8799.n37 75.3623
R19530 a_n6308_8799.n36 a_n6308_8799.n20 70.3058
R19531 a_n6308_8799.n20 a_n6308_8799.n35 70.1674
R19532 a_n6308_8799.n35 a_n6308_8799.n135 20.9683
R19533 a_n6308_8799.n34 a_n6308_8799.n21 75.0448
R19534 a_n6308_8799.n141 a_n6308_8799.n34 11.2134
R19535 a_n6308_8799.n33 a_n6308_8799.n21 80.4688
R19536 a_n6308_8799.n23 a_n6308_8799.n32 74.73
R19537 a_n6308_8799.n31 a_n6308_8799.n23 70.1674
R19538 a_n6308_8799.n144 a_n6308_8799.n31 20.9683
R19539 a_n6308_8799.n22 a_n6308_8799.n30 70.5844
R19540 a_n6308_8799.n47 a_n6308_8799.n46 75.3623
R19541 a_n6308_8799.n45 a_n6308_8799.n16 70.3058
R19542 a_n6308_8799.n16 a_n6308_8799.n44 70.1674
R19543 a_n6308_8799.n44 a_n6308_8799.n146 20.9683
R19544 a_n6308_8799.n43 a_n6308_8799.n17 75.0448
R19545 a_n6308_8799.n152 a_n6308_8799.n43 11.2134
R19546 a_n6308_8799.n42 a_n6308_8799.n17 80.4688
R19547 a_n6308_8799.n19 a_n6308_8799.n41 74.73
R19548 a_n6308_8799.n40 a_n6308_8799.n19 70.1674
R19549 a_n6308_8799.n155 a_n6308_8799.n40 20.9683
R19550 a_n6308_8799.n18 a_n6308_8799.n39 70.5844
R19551 a_n6308_8799.n56 a_n6308_8799.n55 75.3623
R19552 a_n6308_8799.n54 a_n6308_8799.n12 70.3058
R19553 a_n6308_8799.n12 a_n6308_8799.n53 70.1674
R19554 a_n6308_8799.n53 a_n6308_8799.n158 20.9683
R19555 a_n6308_8799.n52 a_n6308_8799.n13 75.0448
R19556 a_n6308_8799.n164 a_n6308_8799.n52 11.2134
R19557 a_n6308_8799.n51 a_n6308_8799.n13 80.4688
R19558 a_n6308_8799.n15 a_n6308_8799.n50 74.73
R19559 a_n6308_8799.n49 a_n6308_8799.n15 70.1674
R19560 a_n6308_8799.n167 a_n6308_8799.n49 20.9683
R19561 a_n6308_8799.n14 a_n6308_8799.n48 70.5844
R19562 a_n6308_8799.n8 a_n6308_8799.n65 70.5844
R19563 a_n6308_8799.n64 a_n6308_8799.n9 70.1674
R19564 a_n6308_8799.n64 a_n6308_8799.n99 20.9683
R19565 a_n6308_8799.n9 a_n6308_8799.n63 74.73
R19566 a_n6308_8799.n108 a_n6308_8799.n63 11.843
R19567 a_n6308_8799.n62 a_n6308_8799.n10 80.4688
R19568 a_n6308_8799.n62 a_n6308_8799.n100 0.365327
R19569 a_n6308_8799.n10 a_n6308_8799.n61 75.0448
R19570 a_n6308_8799.n60 a_n6308_8799.n11 70.1674
R19571 a_n6308_8799.n60 a_n6308_8799.n101 20.9683
R19572 a_n6308_8799.n11 a_n6308_8799.n59 70.3058
R19573 a_n6308_8799.n105 a_n6308_8799.n59 20.6913
R19574 a_n6308_8799.n58 a_n6308_8799.n57 75.3623
R19575 a_n6308_8799.n4 a_n6308_8799.n74 70.5844
R19576 a_n6308_8799.n73 a_n6308_8799.n5 70.1674
R19577 a_n6308_8799.n73 a_n6308_8799.n110 20.9683
R19578 a_n6308_8799.n5 a_n6308_8799.n72 74.73
R19579 a_n6308_8799.n119 a_n6308_8799.n72 11.843
R19580 a_n6308_8799.n71 a_n6308_8799.n6 80.4688
R19581 a_n6308_8799.n71 a_n6308_8799.n111 0.365327
R19582 a_n6308_8799.n6 a_n6308_8799.n70 75.0448
R19583 a_n6308_8799.n69 a_n6308_8799.n7 70.1674
R19584 a_n6308_8799.n69 a_n6308_8799.n112 20.9683
R19585 a_n6308_8799.n7 a_n6308_8799.n68 70.3058
R19586 a_n6308_8799.n116 a_n6308_8799.n68 20.6913
R19587 a_n6308_8799.n67 a_n6308_8799.n66 75.3623
R19588 a_n6308_8799.n0 a_n6308_8799.n83 70.5844
R19589 a_n6308_8799.n82 a_n6308_8799.n1 70.1674
R19590 a_n6308_8799.n82 a_n6308_8799.n122 20.9683
R19591 a_n6308_8799.n1 a_n6308_8799.n81 74.73
R19592 a_n6308_8799.n131 a_n6308_8799.n81 11.843
R19593 a_n6308_8799.n80 a_n6308_8799.n2 80.4688
R19594 a_n6308_8799.n80 a_n6308_8799.n123 0.365327
R19595 a_n6308_8799.n2 a_n6308_8799.n79 75.0448
R19596 a_n6308_8799.n78 a_n6308_8799.n3 70.1674
R19597 a_n6308_8799.n78 a_n6308_8799.n124 20.9683
R19598 a_n6308_8799.n3 a_n6308_8799.n77 70.3058
R19599 a_n6308_8799.n128 a_n6308_8799.n77 20.6913
R19600 a_n6308_8799.n76 a_n6308_8799.n75 75.3623
R19601 a_n6308_8799.n174 a_n6308_8799.n28 98.9632
R19602 a_n6308_8799.n27 a_n6308_8799.n84 98.9631
R19603 a_n6308_8799.n28 a_n6308_8799.n172 98.6055
R19604 a_n6308_8799.n28 a_n6308_8799.n173 98.6055
R19605 a_n6308_8799.n27 a_n6308_8799.n85 98.6055
R19606 a_n6308_8799.n27 a_n6308_8799.n86 98.6055
R19607 a_n6308_8799.n25 a_n6308_8799.n87 81.2902
R19608 a_n6308_8799.n29 a_n6308_8799.n93 81.2902
R19609 a_n6308_8799.n24 a_n6308_8799.n90 81.2902
R19610 a_n6308_8799.n26 a_n6308_8799.n96 80.9324
R19611 a_n6308_8799.n26 a_n6308_8799.n97 80.9324
R19612 a_n6308_8799.n25 a_n6308_8799.n98 80.9324
R19613 a_n6308_8799.n25 a_n6308_8799.n89 80.9324
R19614 a_n6308_8799.n25 a_n6308_8799.n88 80.9324
R19615 a_n6308_8799.n29 a_n6308_8799.n94 80.9324
R19616 a_n6308_8799.n24 a_n6308_8799.n95 80.9324
R19617 a_n6308_8799.n24 a_n6308_8799.n92 80.9324
R19618 a_n6308_8799.n24 a_n6308_8799.n91 80.9324
R19619 a_n6308_8799.n31 a_n6308_8799.n143 20.9683
R19620 a_n6308_8799.n142 a_n6308_8799.n141 48.2005
R19621 a_n6308_8799.n140 a_n6308_8799.n35 20.9683
R19622 a_n6308_8799.n137 a_n6308_8799.n136 48.2005
R19623 a_n6308_8799.n40 a_n6308_8799.n154 20.9683
R19624 a_n6308_8799.n153 a_n6308_8799.n152 48.2005
R19625 a_n6308_8799.n151 a_n6308_8799.n44 20.9683
R19626 a_n6308_8799.n148 a_n6308_8799.n147 48.2005
R19627 a_n6308_8799.n49 a_n6308_8799.n166 20.9683
R19628 a_n6308_8799.n165 a_n6308_8799.n164 48.2005
R19629 a_n6308_8799.n163 a_n6308_8799.n53 20.9683
R19630 a_n6308_8799.n160 a_n6308_8799.n159 48.2005
R19631 a_n6308_8799.n103 a_n6308_8799.n102 48.2005
R19632 a_n6308_8799.n106 a_n6308_8799.n60 20.9683
R19633 a_n6308_8799.n107 a_n6308_8799.n100 48.2005
R19634 a_n6308_8799.n109 a_n6308_8799.n64 20.9683
R19635 a_n6308_8799.n114 a_n6308_8799.n113 48.2005
R19636 a_n6308_8799.n117 a_n6308_8799.n69 20.9683
R19637 a_n6308_8799.n118 a_n6308_8799.n111 48.2005
R19638 a_n6308_8799.n120 a_n6308_8799.n73 20.9683
R19639 a_n6308_8799.n126 a_n6308_8799.n125 48.2005
R19640 a_n6308_8799.n129 a_n6308_8799.n78 20.9683
R19641 a_n6308_8799.n130 a_n6308_8799.n123 48.2005
R19642 a_n6308_8799.n132 a_n6308_8799.n82 20.9683
R19643 a_n6308_8799.n33 a_n6308_8799.n134 47.835
R19644 a_n6308_8799.n36 a_n6308_8799.n139 20.6913
R19645 a_n6308_8799.n42 a_n6308_8799.n145 47.835
R19646 a_n6308_8799.n45 a_n6308_8799.n150 20.6913
R19647 a_n6308_8799.n51 a_n6308_8799.n157 47.835
R19648 a_n6308_8799.n54 a_n6308_8799.n162 20.6913
R19649 a_n6308_8799.n101 a_n6308_8799.n59 21.4216
R19650 a_n6308_8799.n112 a_n6308_8799.n68 21.4216
R19651 a_n6308_8799.n124 a_n6308_8799.n77 21.4216
R19652 a_n6308_8799.t42 a_n6308_8799.n65 484.3
R19653 a_n6308_8799.t51 a_n6308_8799.n74 484.3
R19654 a_n6308_8799.t107 a_n6308_8799.n83 484.3
R19655 a_n6308_8799.n58 a_n6308_8799.n104 45.0871
R19656 a_n6308_8799.n67 a_n6308_8799.n115 45.0871
R19657 a_n6308_8799.n76 a_n6308_8799.n127 45.0871
R19658 a_n6308_8799.n38 a_n6308_8799.n138 45.0871
R19659 a_n6308_8799.n47 a_n6308_8799.n149 45.0871
R19660 a_n6308_8799.n56 a_n6308_8799.n161 45.0871
R19661 a_n6308_8799.n26 a_n6308_8799.n24 32.5134
R19662 a_n6308_8799.n32 a_n6308_8799.n134 11.843
R19663 a_n6308_8799.n139 a_n6308_8799.n37 36.139
R19664 a_n6308_8799.n41 a_n6308_8799.n145 11.843
R19665 a_n6308_8799.n150 a_n6308_8799.n46 36.139
R19666 a_n6308_8799.n50 a_n6308_8799.n157 11.843
R19667 a_n6308_8799.n162 a_n6308_8799.n55 36.139
R19668 a_n6308_8799.n105 a_n6308_8799.n57 36.139
R19669 a_n6308_8799.n99 a_n6308_8799.n63 34.4824
R19670 a_n6308_8799.n116 a_n6308_8799.n66 36.139
R19671 a_n6308_8799.n110 a_n6308_8799.n72 34.4824
R19672 a_n6308_8799.n128 a_n6308_8799.n75 36.139
R19673 a_n6308_8799.n122 a_n6308_8799.n81 34.4824
R19674 a_n6308_8799.n34 a_n6308_8799.n135 35.3134
R19675 a_n6308_8799.n43 a_n6308_8799.n146 35.3134
R19676 a_n6308_8799.n52 a_n6308_8799.n158 35.3134
R19677 a_n6308_8799.n61 a_n6308_8799.n106 35.3134
R19678 a_n6308_8799.n107 a_n6308_8799.n61 11.2134
R19679 a_n6308_8799.n70 a_n6308_8799.n117 35.3134
R19680 a_n6308_8799.n118 a_n6308_8799.n70 11.2134
R19681 a_n6308_8799.n79 a_n6308_8799.n129 35.3134
R19682 a_n6308_8799.n130 a_n6308_8799.n79 11.2134
R19683 a_n6308_8799.n143 a_n6308_8799.n32 34.4824
R19684 a_n6308_8799.n37 a_n6308_8799.n136 10.5784
R19685 a_n6308_8799.n154 a_n6308_8799.n41 34.4824
R19686 a_n6308_8799.n46 a_n6308_8799.n147 10.5784
R19687 a_n6308_8799.n166 a_n6308_8799.n50 34.4824
R19688 a_n6308_8799.n55 a_n6308_8799.n159 10.5784
R19689 a_n6308_8799.n57 a_n6308_8799.n102 10.5784
R19690 a_n6308_8799.n66 a_n6308_8799.n113 10.5784
R19691 a_n6308_8799.n75 a_n6308_8799.n125 10.5784
R19692 a_n6308_8799.n138 a_n6308_8799.n137 14.1472
R19693 a_n6308_8799.n149 a_n6308_8799.n148 14.1472
R19694 a_n6308_8799.n161 a_n6308_8799.n160 14.1472
R19695 a_n6308_8799.n104 a_n6308_8799.n103 14.1472
R19696 a_n6308_8799.n115 a_n6308_8799.n114 14.1472
R19697 a_n6308_8799.n127 a_n6308_8799.n126 14.1472
R19698 a_n6308_8799.n170 a_n6308_8799.n25 12.3339
R19699 a_n6308_8799.n171 a_n6308_8799.n170 11.4887
R19700 a_n6308_8799.n156 a_n6308_8799.n22 9.01755
R19701 a_n6308_8799.n121 a_n6308_8799.n8 9.01755
R19702 a_n6308_8799.n169 a_n6308_8799.n133 6.86452
R19703 a_n6308_8799.n169 a_n6308_8799.n168 6.51829
R19704 a_n6308_8799.n156 a_n6308_8799.n18 4.90959
R19705 a_n6308_8799.n168 a_n6308_8799.n14 4.90959
R19706 a_n6308_8799.n121 a_n6308_8799.n4 4.90959
R19707 a_n6308_8799.n133 a_n6308_8799.n0 4.90959
R19708 a_n6308_8799.n168 a_n6308_8799.n156 4.10845
R19709 a_n6308_8799.n133 a_n6308_8799.n121 4.10845
R19710 a_n6308_8799.n172 a_n6308_8799.t25 3.61217
R19711 a_n6308_8799.n172 a_n6308_8799.t8 3.61217
R19712 a_n6308_8799.n173 a_n6308_8799.t15 3.61217
R19713 a_n6308_8799.n173 a_n6308_8799.t22 3.61217
R19714 a_n6308_8799.n84 a_n6308_8799.t9 3.61217
R19715 a_n6308_8799.n84 a_n6308_8799.t21 3.61217
R19716 a_n6308_8799.n85 a_n6308_8799.t20 3.61217
R19717 a_n6308_8799.n85 a_n6308_8799.t28 3.61217
R19718 a_n6308_8799.n86 a_n6308_8799.t13 3.61217
R19719 a_n6308_8799.n86 a_n6308_8799.t14 3.61217
R19720 a_n6308_8799.t7 a_n6308_8799.n174 3.61217
R19721 a_n6308_8799.n174 a_n6308_8799.t16 3.61217
R19722 a_n6308_8799.n170 a_n6308_8799.n169 3.4105
R19723 a_n6308_8799.n96 a_n6308_8799.t27 2.82907
R19724 a_n6308_8799.n96 a_n6308_8799.t1 2.82907
R19725 a_n6308_8799.n97 a_n6308_8799.t23 2.82907
R19726 a_n6308_8799.n97 a_n6308_8799.t33 2.82907
R19727 a_n6308_8799.n98 a_n6308_8799.t24 2.82907
R19728 a_n6308_8799.n98 a_n6308_8799.t18 2.82907
R19729 a_n6308_8799.n89 a_n6308_8799.t4 2.82907
R19730 a_n6308_8799.n89 a_n6308_8799.t12 2.82907
R19731 a_n6308_8799.n88 a_n6308_8799.t30 2.82907
R19732 a_n6308_8799.n88 a_n6308_8799.t11 2.82907
R19733 a_n6308_8799.n87 a_n6308_8799.t6 2.82907
R19734 a_n6308_8799.n87 a_n6308_8799.t29 2.82907
R19735 a_n6308_8799.n93 a_n6308_8799.t32 2.82907
R19736 a_n6308_8799.n93 a_n6308_8799.t2 2.82907
R19737 a_n6308_8799.n94 a_n6308_8799.t34 2.82907
R19738 a_n6308_8799.n94 a_n6308_8799.t26 2.82907
R19739 a_n6308_8799.n95 a_n6308_8799.t3 2.82907
R19740 a_n6308_8799.n95 a_n6308_8799.t31 2.82907
R19741 a_n6308_8799.n92 a_n6308_8799.t5 2.82907
R19742 a_n6308_8799.n92 a_n6308_8799.t17 2.82907
R19743 a_n6308_8799.n91 a_n6308_8799.t10 2.82907
R19744 a_n6308_8799.n91 a_n6308_8799.t35 2.82907
R19745 a_n6308_8799.n90 a_n6308_8799.t19 2.82907
R19746 a_n6308_8799.n90 a_n6308_8799.t0 2.82907
R19747 a_n6308_8799.n30 a_n6308_8799.n144 22.3251
R19748 a_n6308_8799.n39 a_n6308_8799.n155 22.3251
R19749 a_n6308_8799.n48 a_n6308_8799.n167 22.3251
R19750 a_n6308_8799.n65 a_n6308_8799.n109 22.3251
R19751 a_n6308_8799.n74 a_n6308_8799.n120 22.3251
R19752 a_n6308_8799.n83 a_n6308_8799.n132 22.3251
R19753 a_n6308_8799.n33 a_n6308_8799.n142 0.365327
R19754 a_n6308_8799.n140 a_n6308_8799.n36 21.4216
R19755 a_n6308_8799.n42 a_n6308_8799.n153 0.365327
R19756 a_n6308_8799.n151 a_n6308_8799.n45 21.4216
R19757 a_n6308_8799.n51 a_n6308_8799.n165 0.365327
R19758 a_n6308_8799.n163 a_n6308_8799.n54 21.4216
R19759 a_n6308_8799.n108 a_n6308_8799.n62 47.835
R19760 a_n6308_8799.n119 a_n6308_8799.n71 47.835
R19761 a_n6308_8799.n131 a_n6308_8799.n80 47.835
R19762 a_n6308_8799.n171 a_n6308_8799.n27 31.0347
R19763 a_n6308_8799.n28 a_n6308_8799.n171 18.1305
R19764 a_n6308_8799.n25 a_n6308_8799.n26 1.43153
R19765 a_n6308_8799.n24 a_n6308_8799.n29 1.07378
R19766 a_n6308_8799.n23 a_n6308_8799.n21 0.758076
R19767 a_n6308_8799.n21 a_n6308_8799.n20 0.758076
R19768 a_n6308_8799.n38 a_n6308_8799.n20 0.758076
R19769 a_n6308_8799.n19 a_n6308_8799.n17 0.758076
R19770 a_n6308_8799.n17 a_n6308_8799.n16 0.758076
R19771 a_n6308_8799.n47 a_n6308_8799.n16 0.758076
R19772 a_n6308_8799.n15 a_n6308_8799.n13 0.758076
R19773 a_n6308_8799.n13 a_n6308_8799.n12 0.758076
R19774 a_n6308_8799.n56 a_n6308_8799.n12 0.758076
R19775 a_n6308_8799.n11 a_n6308_8799.n10 0.758076
R19776 a_n6308_8799.n10 a_n6308_8799.n9 0.758076
R19777 a_n6308_8799.n9 a_n6308_8799.n8 0.758076
R19778 a_n6308_8799.n7 a_n6308_8799.n6 0.758076
R19779 a_n6308_8799.n6 a_n6308_8799.n5 0.758076
R19780 a_n6308_8799.n5 a_n6308_8799.n4 0.758076
R19781 a_n6308_8799.n3 a_n6308_8799.n2 0.758076
R19782 a_n6308_8799.n2 a_n6308_8799.n1 0.758076
R19783 a_n6308_8799.n1 a_n6308_8799.n0 0.758076
R19784 a_n6308_8799.n76 a_n6308_8799.n3 0.568682
R19785 a_n6308_8799.n67 a_n6308_8799.n7 0.568682
R19786 a_n6308_8799.n58 a_n6308_8799.n11 0.568682
R19787 a_n6308_8799.n15 a_n6308_8799.n14 0.568682
R19788 a_n6308_8799.n19 a_n6308_8799.n18 0.568682
R19789 a_n6308_8799.n23 a_n6308_8799.n22 0.568682
R19790 a_n1986_13878.n88 a_n1986_13878.t64 512.366
R19791 a_n1986_13878.n78 a_n1986_13878.t55 512.366
R19792 a_n1986_13878.n89 a_n1986_13878.t49 512.366
R19793 a_n1986_13878.n86 a_n1986_13878.t72 512.366
R19794 a_n1986_13878.n79 a_n1986_13878.t61 512.366
R19795 a_n1986_13878.n87 a_n1986_13878.t60 512.366
R19796 a_n1986_13878.n84 a_n1986_13878.t68 512.366
R19797 a_n1986_13878.n80 a_n1986_13878.t53 512.366
R19798 a_n1986_13878.n85 a_n1986_13878.t54 512.366
R19799 a_n1986_13878.n82 a_n1986_13878.t57 512.366
R19800 a_n1986_13878.n81 a_n1986_13878.t66 512.366
R19801 a_n1986_13878.n83 a_n1986_13878.t48 512.366
R19802 a_n1986_13878.n20 a_n1986_13878.t75 539.01
R19803 a_n1986_13878.n93 a_n1986_13878.t58 512.366
R19804 a_n1986_13878.n92 a_n1986_13878.t62 512.366
R19805 a_n1986_13878.n66 a_n1986_13878.t52 512.366
R19806 a_n1986_13878.n91 a_n1986_13878.t67 512.366
R19807 a_n1986_13878.n52 a_n1986_13878.t16 533.058
R19808 a_n1986_13878.n22 a_n1986_13878.t0 539.01
R19809 a_n1986_13878.n96 a_n1986_13878.t2 512.366
R19810 a_n1986_13878.n95 a_n1986_13878.t6 512.366
R19811 a_n1986_13878.n53 a_n1986_13878.t20 512.366
R19812 a_n1986_13878.n94 a_n1986_13878.t12 512.366
R19813 a_n1986_13878.n12 a_n1986_13878.t18 539.01
R19814 a_n1986_13878.n74 a_n1986_13878.t8 512.366
R19815 a_n1986_13878.n75 a_n1986_13878.t4 512.366
R19816 a_n1986_13878.n69 a_n1986_13878.t10 512.366
R19817 a_n1986_13878.n76 a_n1986_13878.t14 512.366
R19818 a_n1986_13878.n16 a_n1986_13878.t70 539.01
R19819 a_n1986_13878.n71 a_n1986_13878.t71 512.366
R19820 a_n1986_13878.n72 a_n1986_13878.t50 512.366
R19821 a_n1986_13878.n70 a_n1986_13878.t56 512.366
R19822 a_n1986_13878.n73 a_n1986_13878.t65 512.366
R19823 a_n1986_13878.n0 a_n1986_13878.n51 70.1674
R19824 a_n1986_13878.n2 a_n1986_13878.n49 70.1674
R19825 a_n1986_13878.n4 a_n1986_13878.n47 70.1674
R19826 a_n1986_13878.n7 a_n1986_13878.n45 70.1674
R19827 a_n1986_13878.n37 a_n1986_13878.n18 70.3058
R19828 a_n1986_13878.n31 a_n1986_13878.n34 70.1674
R19829 a_n1986_13878.n34 a_n1986_13878.n53 20.9683
R19830 a_n1986_13878.n33 a_n1986_13878.n32 75.0448
R19831 a_n1986_13878.n95 a_n1986_13878.n33 11.2134
R19832 a_n1986_13878.n21 a_n1986_13878.n22 44.8194
R19833 a_n1986_13878.n52 a_n1986_13878.n31 70.3058
R19834 a_n1986_13878.n19 a_n1986_13878.n36 70.1674
R19835 a_n1986_13878.n36 a_n1986_13878.n66 20.9683
R19836 a_n1986_13878.n35 a_n1986_13878.n19 75.0448
R19837 a_n1986_13878.n92 a_n1986_13878.n35 11.2134
R19838 a_n1986_13878.n17 a_n1986_13878.n20 44.8194
R19839 a_n1986_13878.n9 a_n1986_13878.n43 70.3058
R19840 a_n1986_13878.n13 a_n1986_13878.n40 70.3058
R19841 a_n1986_13878.n39 a_n1986_13878.n14 70.1674
R19842 a_n1986_13878.n39 a_n1986_13878.n70 20.9683
R19843 a_n1986_13878.n14 a_n1986_13878.n38 75.0448
R19844 a_n1986_13878.n72 a_n1986_13878.n38 11.2134
R19845 a_n1986_13878.n15 a_n1986_13878.n16 44.8194
R19846 a_n1986_13878.n42 a_n1986_13878.n10 70.1674
R19847 a_n1986_13878.n42 a_n1986_13878.n69 20.9683
R19848 a_n1986_13878.n10 a_n1986_13878.n41 75.0448
R19849 a_n1986_13878.n75 a_n1986_13878.n41 11.2134
R19850 a_n1986_13878.n11 a_n1986_13878.n12 44.8194
R19851 a_n1986_13878.n83 a_n1986_13878.n45 20.9683
R19852 a_n1986_13878.n44 a_n1986_13878.n8 75.0448
R19853 a_n1986_13878.n44 a_n1986_13878.n81 11.2134
R19854 a_n1986_13878.n8 a_n1986_13878.n82 161.3
R19855 a_n1986_13878.n85 a_n1986_13878.n47 20.9683
R19856 a_n1986_13878.n46 a_n1986_13878.n5 75.0448
R19857 a_n1986_13878.n46 a_n1986_13878.n80 11.2134
R19858 a_n1986_13878.n5 a_n1986_13878.n84 161.3
R19859 a_n1986_13878.n87 a_n1986_13878.n49 20.9683
R19860 a_n1986_13878.n48 a_n1986_13878.n3 75.0448
R19861 a_n1986_13878.n48 a_n1986_13878.n79 11.2134
R19862 a_n1986_13878.n3 a_n1986_13878.n86 161.3
R19863 a_n1986_13878.n89 a_n1986_13878.n51 20.9683
R19864 a_n1986_13878.n50 a_n1986_13878.n1 75.0448
R19865 a_n1986_13878.n50 a_n1986_13878.n78 11.2134
R19866 a_n1986_13878.n1 a_n1986_13878.n88 161.3
R19867 a_n1986_13878.n29 a_n1986_13878.n63 81.2902
R19868 a_n1986_13878.n30 a_n1986_13878.n57 81.2902
R19869 a_n1986_13878.n23 a_n1986_13878.n54 81.2902
R19870 a_n1986_13878.n29 a_n1986_13878.n64 80.9324
R19871 a_n1986_13878.n25 a_n1986_13878.n65 80.9324
R19872 a_n1986_13878.n25 a_n1986_13878.n62 80.9324
R19873 a_n1986_13878.n25 a_n1986_13878.n61 80.9324
R19874 a_n1986_13878.n24 a_n1986_13878.n60 80.9324
R19875 a_n1986_13878.n30 a_n1986_13878.n58 80.9324
R19876 a_n1986_13878.n23 a_n1986_13878.n59 80.9324
R19877 a_n1986_13878.n23 a_n1986_13878.n56 80.9324
R19878 a_n1986_13878.n23 a_n1986_13878.n55 80.9324
R19879 a_n1986_13878.n28 a_n1986_13878.t17 74.6477
R19880 a_n1986_13878.n26 a_n1986_13878.t19 74.6477
R19881 a_n1986_13878.t1 a_n1986_13878.n100 74.2899
R19882 a_n1986_13878.n27 a_n1986_13878.t23 74.2897
R19883 a_n1986_13878.n28 a_n1986_13878.n98 70.6783
R19884 a_n1986_13878.n28 a_n1986_13878.n99 70.6783
R19885 a_n1986_13878.n27 a_n1986_13878.n68 70.6783
R19886 a_n1986_13878.n26 a_n1986_13878.n67 70.6783
R19887 a_n1986_13878.n88 a_n1986_13878.n78 48.2005
R19888 a_n1986_13878.t69 a_n1986_13878.n51 533.335
R19889 a_n1986_13878.n86 a_n1986_13878.n79 48.2005
R19890 a_n1986_13878.t74 a_n1986_13878.n49 533.335
R19891 a_n1986_13878.n84 a_n1986_13878.n80 48.2005
R19892 a_n1986_13878.t63 a_n1986_13878.n47 533.335
R19893 a_n1986_13878.n82 a_n1986_13878.n81 48.2005
R19894 a_n1986_13878.t59 a_n1986_13878.n45 533.335
R19895 a_n1986_13878.n93 a_n1986_13878.n92 48.2005
R19896 a_n1986_13878.n91 a_n1986_13878.n36 20.9683
R19897 a_n1986_13878.n96 a_n1986_13878.n95 48.2005
R19898 a_n1986_13878.n94 a_n1986_13878.n34 20.9683
R19899 a_n1986_13878.n75 a_n1986_13878.n74 48.2005
R19900 a_n1986_13878.n76 a_n1986_13878.n42 20.9683
R19901 a_n1986_13878.n72 a_n1986_13878.n71 48.2005
R19902 a_n1986_13878.n73 a_n1986_13878.n39 20.9683
R19903 a_n1986_13878.n37 a_n1986_13878.t73 533.058
R19904 a_n1986_13878.t22 a_n1986_13878.n43 533.058
R19905 a_n1986_13878.t51 a_n1986_13878.n40 533.058
R19906 a_n1986_13878.n24 a_n1986_13878.n23 31.7747
R19907 a_n1986_13878.n89 a_n1986_13878.n50 35.3134
R19908 a_n1986_13878.n87 a_n1986_13878.n48 35.3134
R19909 a_n1986_13878.n85 a_n1986_13878.n46 35.3134
R19910 a_n1986_13878.n83 a_n1986_13878.n44 35.3134
R19911 a_n1986_13878.n35 a_n1986_13878.n66 35.3134
R19912 a_n1986_13878.n33 a_n1986_13878.n53 35.3134
R19913 a_n1986_13878.n69 a_n1986_13878.n41 35.3134
R19914 a_n1986_13878.n70 a_n1986_13878.n38 35.3134
R19915 a_n1986_13878.n31 a_n1986_13878.n25 23.891
R19916 a_n1986_13878.n15 a_n1986_13878.n6 12.046
R19917 a_n1986_13878.n18 a_n1986_13878.n90 11.8414
R19918 a_n1986_13878.n97 a_n1986_13878.n21 10.5365
R19919 a_n1986_13878.n77 a_n1986_13878.n27 9.50122
R19920 a_n1986_13878.n90 a_n1986_13878.n0 7.47588
R19921 a_n1986_13878.n8 a_n1986_13878.n6 7.47588
R19922 a_n1986_13878.n77 a_n1986_13878.n9 6.70126
R19923 a_n1986_13878.n100 a_n1986_13878.n97 5.65783
R19924 a_n1986_13878.n90 a_n1986_13878.n77 5.3452
R19925 a_n1986_13878.n31 a_n1986_13878.n17 3.95126
R19926 a_n1986_13878.n11 a_n1986_13878.n13 3.95126
R19927 a_n1986_13878.n98 a_n1986_13878.t21 3.61217
R19928 a_n1986_13878.n98 a_n1986_13878.t13 3.61217
R19929 a_n1986_13878.n99 a_n1986_13878.t3 3.61217
R19930 a_n1986_13878.n99 a_n1986_13878.t7 3.61217
R19931 a_n1986_13878.n68 a_n1986_13878.t11 3.61217
R19932 a_n1986_13878.n68 a_n1986_13878.t15 3.61217
R19933 a_n1986_13878.n67 a_n1986_13878.t9 3.61217
R19934 a_n1986_13878.n67 a_n1986_13878.t5 3.61217
R19935 a_n1986_13878.n63 a_n1986_13878.t39 2.82907
R19936 a_n1986_13878.n63 a_n1986_13878.t24 2.82907
R19937 a_n1986_13878.n64 a_n1986_13878.t36 2.82907
R19938 a_n1986_13878.n64 a_n1986_13878.t25 2.82907
R19939 a_n1986_13878.n65 a_n1986_13878.t47 2.82907
R19940 a_n1986_13878.n65 a_n1986_13878.t32 2.82907
R19941 a_n1986_13878.n62 a_n1986_13878.t27 2.82907
R19942 a_n1986_13878.n62 a_n1986_13878.t43 2.82907
R19943 a_n1986_13878.n61 a_n1986_13878.t41 2.82907
R19944 a_n1986_13878.n61 a_n1986_13878.t40 2.82907
R19945 a_n1986_13878.n60 a_n1986_13878.t30 2.82907
R19946 a_n1986_13878.n60 a_n1986_13878.t31 2.82907
R19947 a_n1986_13878.n57 a_n1986_13878.t33 2.82907
R19948 a_n1986_13878.n57 a_n1986_13878.t37 2.82907
R19949 a_n1986_13878.n58 a_n1986_13878.t42 2.82907
R19950 a_n1986_13878.n58 a_n1986_13878.t28 2.82907
R19951 a_n1986_13878.n59 a_n1986_13878.t34 2.82907
R19952 a_n1986_13878.n59 a_n1986_13878.t44 2.82907
R19953 a_n1986_13878.n56 a_n1986_13878.t26 2.82907
R19954 a_n1986_13878.n56 a_n1986_13878.t35 2.82907
R19955 a_n1986_13878.n55 a_n1986_13878.t38 2.82907
R19956 a_n1986_13878.n55 a_n1986_13878.t46 2.82907
R19957 a_n1986_13878.n54 a_n1986_13878.t45 2.82907
R19958 a_n1986_13878.n54 a_n1986_13878.t29 2.82907
R19959 a_n1986_13878.n97 a_n1986_13878.n6 1.30542
R19960 a_n1986_13878.n3 a_n1986_13878.n4 1.04595
R19961 a_n1986_13878.n20 a_n1986_13878.n93 13.657
R19962 a_n1986_13878.n91 a_n1986_13878.n37 21.4216
R19963 a_n1986_13878.n22 a_n1986_13878.n96 13.657
R19964 a_n1986_13878.n94 a_n1986_13878.n52 21.4216
R19965 a_n1986_13878.n74 a_n1986_13878.n12 13.657
R19966 a_n1986_13878.n43 a_n1986_13878.n76 21.4216
R19967 a_n1986_13878.n71 a_n1986_13878.n16 13.657
R19968 a_n1986_13878.n40 a_n1986_13878.n73 21.4216
R19969 a_n1986_13878.n23 a_n1986_13878.n30 1.07378
R19970 a_n1986_13878.n32 a_n1986_13878.n21 0.758076
R19971 a_n1986_13878.n19 a_n1986_13878.n17 0.758076
R19972 a_n1986_13878.n19 a_n1986_13878.n18 0.758076
R19973 a_n1986_13878.n15 a_n1986_13878.n14 0.758076
R19974 a_n1986_13878.n14 a_n1986_13878.n13 0.758076
R19975 a_n1986_13878.n11 a_n1986_13878.n10 0.758076
R19976 a_n1986_13878.n10 a_n1986_13878.n9 0.758076
R19977 a_n1986_13878.n8 a_n1986_13878.n7 0.758076
R19978 a_n1986_13878.n5 a_n1986_13878.n4 0.758076
R19979 a_n1986_13878.n3 a_n1986_13878.n2 0.758076
R19980 a_n1986_13878.n1 a_n1986_13878.n0 0.758076
R19981 a_n1986_13878.n32 a_n1986_13878.n31 0.720197
R19982 a_n1986_13878.n25 a_n1986_13878.n29 0.716017
R19983 a_n1986_13878.n100 a_n1986_13878.n28 0.716017
R19984 a_n1986_13878.n27 a_n1986_13878.n26 0.716017
R19985 a_n1986_13878.n25 a_n1986_13878.n24 0.716017
R19986 a_n1986_13878.n5 a_n1986_13878.n7 0.67853
R19987 a_n1986_13878.n1 a_n1986_13878.n2 0.67853
R19988 a_n1986_8322.n6 a_n1986_8322.t18 74.6477
R19989 a_n1986_8322.n1 a_n1986_8322.t5 74.6477
R19990 a_n1986_8322.n16 a_n1986_8322.t14 74.6474
R19991 a_n1986_8322.n14 a_n1986_8322.t7 74.2899
R19992 a_n1986_8322.n7 a_n1986_8322.t16 74.2899
R19993 a_n1986_8322.n8 a_n1986_8322.t19 74.2899
R19994 a_n1986_8322.n11 a_n1986_8322.t20 74.2899
R19995 a_n1986_8322.n4 a_n1986_8322.t4 74.2899
R19996 a_n1986_8322.n16 a_n1986_8322.n15 70.6783
R19997 a_n1986_8322.n6 a_n1986_8322.n5 70.6783
R19998 a_n1986_8322.n10 a_n1986_8322.n9 70.6783
R19999 a_n1986_8322.n1 a_n1986_8322.n0 70.6783
R20000 a_n1986_8322.n3 a_n1986_8322.n2 70.6783
R20001 a_n1986_8322.n18 a_n1986_8322.n17 70.6782
R20002 a_n1986_8322.n12 a_n1986_8322.n4 22.7556
R20003 a_n1986_8322.n13 a_n1986_8322.t2 9.7972
R20004 a_n1986_8322.n12 a_n1986_8322.n11 6.2408
R20005 a_n1986_8322.n14 a_n1986_8322.n13 5.83671
R20006 a_n1986_8322.n13 a_n1986_8322.n12 5.3452
R20007 a_n1986_8322.n15 a_n1986_8322.t12 3.61217
R20008 a_n1986_8322.n15 a_n1986_8322.t9 3.61217
R20009 a_n1986_8322.n5 a_n1986_8322.t22 3.61217
R20010 a_n1986_8322.n5 a_n1986_8322.t21 3.61217
R20011 a_n1986_8322.n9 a_n1986_8322.t17 3.61217
R20012 a_n1986_8322.n9 a_n1986_8322.t23 3.61217
R20013 a_n1986_8322.n0 a_n1986_8322.t13 3.61217
R20014 a_n1986_8322.n0 a_n1986_8322.t8 3.61217
R20015 a_n1986_8322.n2 a_n1986_8322.t11 3.61217
R20016 a_n1986_8322.n2 a_n1986_8322.t10 3.61217
R20017 a_n1986_8322.n18 a_n1986_8322.t6 3.61217
R20018 a_n1986_8322.t15 a_n1986_8322.n18 3.61217
R20019 a_n1986_8322.n11 a_n1986_8322.n10 0.358259
R20020 a_n1986_8322.n10 a_n1986_8322.n8 0.358259
R20021 a_n1986_8322.n7 a_n1986_8322.n6 0.358259
R20022 a_n1986_8322.n4 a_n1986_8322.n3 0.358259
R20023 a_n1986_8322.n3 a_n1986_8322.n1 0.358259
R20024 a_n1986_8322.n17 a_n1986_8322.n14 0.358259
R20025 a_n1986_8322.n17 a_n1986_8322.n16 0.358259
R20026 a_n1986_8322.n8 a_n1986_8322.n7 0.101793
R20027 a_n1986_8322.t3 a_n1986_8322.t0 0.0788333
R20028 a_n1986_8322.t1 a_n1986_8322.t3 0.0631667
R20029 a_n1986_8322.t2 a_n1986_8322.t1 0.0471944
R20030 a_n1986_8322.t2 a_n1986_8322.t0 0.0453889
R20031 a_n1808_13878.n16 a_n1808_13878.n0 98.9633
R20032 a_n1808_13878.n3 a_n1808_13878.n1 98.7517
R20033 a_n1808_13878.n5 a_n1808_13878.n4 98.6055
R20034 a_n1808_13878.n3 a_n1808_13878.n2 98.6055
R20035 a_n1808_13878.n17 a_n1808_13878.n16 98.6054
R20036 a_n1808_13878.n15 a_n1808_13878.n14 98.6054
R20037 a_n1808_13878.n7 a_n1808_13878.t1 74.6477
R20038 a_n1808_13878.n12 a_n1808_13878.t2 74.2899
R20039 a_n1808_13878.n9 a_n1808_13878.t3 74.2899
R20040 a_n1808_13878.n8 a_n1808_13878.t0 74.2899
R20041 a_n1808_13878.n11 a_n1808_13878.n10 70.6783
R20042 a_n1808_13878.n7 a_n1808_13878.n6 70.6783
R20043 a_n1808_13878.n13 a_n1808_13878.n5 13.5694
R20044 a_n1808_13878.n15 a_n1808_13878.n13 11.5762
R20045 a_n1808_13878.n13 a_n1808_13878.n12 6.2408
R20046 a_n1808_13878.n14 a_n1808_13878.t15 3.61217
R20047 a_n1808_13878.n14 a_n1808_13878.t16 3.61217
R20048 a_n1808_13878.n0 a_n1808_13878.t13 3.61217
R20049 a_n1808_13878.n0 a_n1808_13878.t17 3.61217
R20050 a_n1808_13878.n10 a_n1808_13878.t6 3.61217
R20051 a_n1808_13878.n10 a_n1808_13878.t7 3.61217
R20052 a_n1808_13878.n6 a_n1808_13878.t4 3.61217
R20053 a_n1808_13878.n6 a_n1808_13878.t5 3.61217
R20054 a_n1808_13878.n4 a_n1808_13878.t12 3.61217
R20055 a_n1808_13878.n4 a_n1808_13878.t19 3.61217
R20056 a_n1808_13878.n2 a_n1808_13878.t14 3.61217
R20057 a_n1808_13878.n2 a_n1808_13878.t9 3.61217
R20058 a_n1808_13878.n1 a_n1808_13878.t8 3.61217
R20059 a_n1808_13878.n1 a_n1808_13878.t10 3.61217
R20060 a_n1808_13878.t18 a_n1808_13878.n17 3.61217
R20061 a_n1808_13878.n17 a_n1808_13878.t11 3.61217
R20062 a_n1808_13878.n8 a_n1808_13878.n7 0.358259
R20063 a_n1808_13878.n11 a_n1808_13878.n9 0.358259
R20064 a_n1808_13878.n12 a_n1808_13878.n11 0.358259
R20065 a_n1808_13878.n16 a_n1808_13878.n15 0.358259
R20066 a_n1808_13878.n5 a_n1808_13878.n3 0.146627
R20067 a_n1808_13878.n9 a_n1808_13878.n8 0.101793
R20068 outputibias.n27 outputibias.n1 289.615
R20069 outputibias.n58 outputibias.n32 289.615
R20070 outputibias.n90 outputibias.n64 289.615
R20071 outputibias.n122 outputibias.n96 289.615
R20072 outputibias.n28 outputibias.n27 185
R20073 outputibias.n26 outputibias.n25 185
R20074 outputibias.n5 outputibias.n4 185
R20075 outputibias.n20 outputibias.n19 185
R20076 outputibias.n18 outputibias.n17 185
R20077 outputibias.n9 outputibias.n8 185
R20078 outputibias.n12 outputibias.n11 185
R20079 outputibias.n59 outputibias.n58 185
R20080 outputibias.n57 outputibias.n56 185
R20081 outputibias.n36 outputibias.n35 185
R20082 outputibias.n51 outputibias.n50 185
R20083 outputibias.n49 outputibias.n48 185
R20084 outputibias.n40 outputibias.n39 185
R20085 outputibias.n43 outputibias.n42 185
R20086 outputibias.n91 outputibias.n90 185
R20087 outputibias.n89 outputibias.n88 185
R20088 outputibias.n68 outputibias.n67 185
R20089 outputibias.n83 outputibias.n82 185
R20090 outputibias.n81 outputibias.n80 185
R20091 outputibias.n72 outputibias.n71 185
R20092 outputibias.n75 outputibias.n74 185
R20093 outputibias.n123 outputibias.n122 185
R20094 outputibias.n121 outputibias.n120 185
R20095 outputibias.n100 outputibias.n99 185
R20096 outputibias.n115 outputibias.n114 185
R20097 outputibias.n113 outputibias.n112 185
R20098 outputibias.n104 outputibias.n103 185
R20099 outputibias.n107 outputibias.n106 185
R20100 outputibias.n0 outputibias.t8 178.945
R20101 outputibias.n133 outputibias.t10 177.018
R20102 outputibias.n132 outputibias.t11 177.018
R20103 outputibias.n0 outputibias.t9 177.018
R20104 outputibias.t5 outputibias.n10 147.661
R20105 outputibias.t7 outputibias.n41 147.661
R20106 outputibias.t1 outputibias.n73 147.661
R20107 outputibias.t3 outputibias.n105 147.661
R20108 outputibias.n128 outputibias.t4 132.363
R20109 outputibias.n128 outputibias.t6 130.436
R20110 outputibias.n129 outputibias.t0 130.436
R20111 outputibias.n130 outputibias.t2 130.436
R20112 outputibias.n27 outputibias.n26 104.615
R20113 outputibias.n26 outputibias.n4 104.615
R20114 outputibias.n19 outputibias.n4 104.615
R20115 outputibias.n19 outputibias.n18 104.615
R20116 outputibias.n18 outputibias.n8 104.615
R20117 outputibias.n11 outputibias.n8 104.615
R20118 outputibias.n58 outputibias.n57 104.615
R20119 outputibias.n57 outputibias.n35 104.615
R20120 outputibias.n50 outputibias.n35 104.615
R20121 outputibias.n50 outputibias.n49 104.615
R20122 outputibias.n49 outputibias.n39 104.615
R20123 outputibias.n42 outputibias.n39 104.615
R20124 outputibias.n90 outputibias.n89 104.615
R20125 outputibias.n89 outputibias.n67 104.615
R20126 outputibias.n82 outputibias.n67 104.615
R20127 outputibias.n82 outputibias.n81 104.615
R20128 outputibias.n81 outputibias.n71 104.615
R20129 outputibias.n74 outputibias.n71 104.615
R20130 outputibias.n122 outputibias.n121 104.615
R20131 outputibias.n121 outputibias.n99 104.615
R20132 outputibias.n114 outputibias.n99 104.615
R20133 outputibias.n114 outputibias.n113 104.615
R20134 outputibias.n113 outputibias.n103 104.615
R20135 outputibias.n106 outputibias.n103 104.615
R20136 outputibias.n63 outputibias.n31 95.6354
R20137 outputibias.n63 outputibias.n62 94.6732
R20138 outputibias.n95 outputibias.n94 94.6732
R20139 outputibias.n127 outputibias.n126 94.6732
R20140 outputibias.n11 outputibias.t5 52.3082
R20141 outputibias.n42 outputibias.t7 52.3082
R20142 outputibias.n74 outputibias.t1 52.3082
R20143 outputibias.n106 outputibias.t3 52.3082
R20144 outputibias.n12 outputibias.n10 15.6674
R20145 outputibias.n43 outputibias.n41 15.6674
R20146 outputibias.n75 outputibias.n73 15.6674
R20147 outputibias.n107 outputibias.n105 15.6674
R20148 outputibias.n13 outputibias.n9 12.8005
R20149 outputibias.n44 outputibias.n40 12.8005
R20150 outputibias.n76 outputibias.n72 12.8005
R20151 outputibias.n108 outputibias.n104 12.8005
R20152 outputibias.n17 outputibias.n16 12.0247
R20153 outputibias.n48 outputibias.n47 12.0247
R20154 outputibias.n80 outputibias.n79 12.0247
R20155 outputibias.n112 outputibias.n111 12.0247
R20156 outputibias.n20 outputibias.n7 11.249
R20157 outputibias.n51 outputibias.n38 11.249
R20158 outputibias.n83 outputibias.n70 11.249
R20159 outputibias.n115 outputibias.n102 11.249
R20160 outputibias.n21 outputibias.n5 10.4732
R20161 outputibias.n52 outputibias.n36 10.4732
R20162 outputibias.n84 outputibias.n68 10.4732
R20163 outputibias.n116 outputibias.n100 10.4732
R20164 outputibias.n25 outputibias.n24 9.69747
R20165 outputibias.n56 outputibias.n55 9.69747
R20166 outputibias.n88 outputibias.n87 9.69747
R20167 outputibias.n120 outputibias.n119 9.69747
R20168 outputibias.n31 outputibias.n30 9.45567
R20169 outputibias.n62 outputibias.n61 9.45567
R20170 outputibias.n94 outputibias.n93 9.45567
R20171 outputibias.n126 outputibias.n125 9.45567
R20172 outputibias.n30 outputibias.n29 9.3005
R20173 outputibias.n3 outputibias.n2 9.3005
R20174 outputibias.n24 outputibias.n23 9.3005
R20175 outputibias.n22 outputibias.n21 9.3005
R20176 outputibias.n7 outputibias.n6 9.3005
R20177 outputibias.n16 outputibias.n15 9.3005
R20178 outputibias.n14 outputibias.n13 9.3005
R20179 outputibias.n61 outputibias.n60 9.3005
R20180 outputibias.n34 outputibias.n33 9.3005
R20181 outputibias.n55 outputibias.n54 9.3005
R20182 outputibias.n53 outputibias.n52 9.3005
R20183 outputibias.n38 outputibias.n37 9.3005
R20184 outputibias.n47 outputibias.n46 9.3005
R20185 outputibias.n45 outputibias.n44 9.3005
R20186 outputibias.n93 outputibias.n92 9.3005
R20187 outputibias.n66 outputibias.n65 9.3005
R20188 outputibias.n87 outputibias.n86 9.3005
R20189 outputibias.n85 outputibias.n84 9.3005
R20190 outputibias.n70 outputibias.n69 9.3005
R20191 outputibias.n79 outputibias.n78 9.3005
R20192 outputibias.n77 outputibias.n76 9.3005
R20193 outputibias.n125 outputibias.n124 9.3005
R20194 outputibias.n98 outputibias.n97 9.3005
R20195 outputibias.n119 outputibias.n118 9.3005
R20196 outputibias.n117 outputibias.n116 9.3005
R20197 outputibias.n102 outputibias.n101 9.3005
R20198 outputibias.n111 outputibias.n110 9.3005
R20199 outputibias.n109 outputibias.n108 9.3005
R20200 outputibias.n28 outputibias.n3 8.92171
R20201 outputibias.n59 outputibias.n34 8.92171
R20202 outputibias.n91 outputibias.n66 8.92171
R20203 outputibias.n123 outputibias.n98 8.92171
R20204 outputibias.n29 outputibias.n1 8.14595
R20205 outputibias.n60 outputibias.n32 8.14595
R20206 outputibias.n92 outputibias.n64 8.14595
R20207 outputibias.n124 outputibias.n96 8.14595
R20208 outputibias.n31 outputibias.n1 5.81868
R20209 outputibias.n62 outputibias.n32 5.81868
R20210 outputibias.n94 outputibias.n64 5.81868
R20211 outputibias.n126 outputibias.n96 5.81868
R20212 outputibias.n131 outputibias.n130 5.20947
R20213 outputibias.n29 outputibias.n28 5.04292
R20214 outputibias.n60 outputibias.n59 5.04292
R20215 outputibias.n92 outputibias.n91 5.04292
R20216 outputibias.n124 outputibias.n123 5.04292
R20217 outputibias.n131 outputibias.n127 4.42209
R20218 outputibias.n14 outputibias.n10 4.38594
R20219 outputibias.n45 outputibias.n41 4.38594
R20220 outputibias.n77 outputibias.n73 4.38594
R20221 outputibias.n109 outputibias.n105 4.38594
R20222 outputibias.n132 outputibias.n131 4.28454
R20223 outputibias.n25 outputibias.n3 4.26717
R20224 outputibias.n56 outputibias.n34 4.26717
R20225 outputibias.n88 outputibias.n66 4.26717
R20226 outputibias.n120 outputibias.n98 4.26717
R20227 outputibias.n24 outputibias.n5 3.49141
R20228 outputibias.n55 outputibias.n36 3.49141
R20229 outputibias.n87 outputibias.n68 3.49141
R20230 outputibias.n119 outputibias.n100 3.49141
R20231 outputibias.n21 outputibias.n20 2.71565
R20232 outputibias.n52 outputibias.n51 2.71565
R20233 outputibias.n84 outputibias.n83 2.71565
R20234 outputibias.n116 outputibias.n115 2.71565
R20235 outputibias.n17 outputibias.n7 1.93989
R20236 outputibias.n48 outputibias.n38 1.93989
R20237 outputibias.n80 outputibias.n70 1.93989
R20238 outputibias.n112 outputibias.n102 1.93989
R20239 outputibias.n130 outputibias.n129 1.9266
R20240 outputibias.n129 outputibias.n128 1.9266
R20241 outputibias.n133 outputibias.n132 1.92658
R20242 outputibias.n134 outputibias.n133 1.29913
R20243 outputibias.n16 outputibias.n9 1.16414
R20244 outputibias.n47 outputibias.n40 1.16414
R20245 outputibias.n79 outputibias.n72 1.16414
R20246 outputibias.n111 outputibias.n104 1.16414
R20247 outputibias.n127 outputibias.n95 0.962709
R20248 outputibias.n95 outputibias.n63 0.962709
R20249 outputibias.n13 outputibias.n12 0.388379
R20250 outputibias.n44 outputibias.n43 0.388379
R20251 outputibias.n76 outputibias.n75 0.388379
R20252 outputibias.n108 outputibias.n107 0.388379
R20253 outputibias.n134 outputibias.n0 0.337251
R20254 outputibias outputibias.n134 0.302375
R20255 outputibias.n30 outputibias.n2 0.155672
R20256 outputibias.n23 outputibias.n2 0.155672
R20257 outputibias.n23 outputibias.n22 0.155672
R20258 outputibias.n22 outputibias.n6 0.155672
R20259 outputibias.n15 outputibias.n6 0.155672
R20260 outputibias.n15 outputibias.n14 0.155672
R20261 outputibias.n61 outputibias.n33 0.155672
R20262 outputibias.n54 outputibias.n33 0.155672
R20263 outputibias.n54 outputibias.n53 0.155672
R20264 outputibias.n53 outputibias.n37 0.155672
R20265 outputibias.n46 outputibias.n37 0.155672
R20266 outputibias.n46 outputibias.n45 0.155672
R20267 outputibias.n93 outputibias.n65 0.155672
R20268 outputibias.n86 outputibias.n65 0.155672
R20269 outputibias.n86 outputibias.n85 0.155672
R20270 outputibias.n85 outputibias.n69 0.155672
R20271 outputibias.n78 outputibias.n69 0.155672
R20272 outputibias.n78 outputibias.n77 0.155672
R20273 outputibias.n125 outputibias.n97 0.155672
R20274 outputibias.n118 outputibias.n97 0.155672
R20275 outputibias.n118 outputibias.n117 0.155672
R20276 outputibias.n117 outputibias.n101 0.155672
R20277 outputibias.n110 outputibias.n101 0.155672
R20278 outputibias.n110 outputibias.n109 0.155672
R20279 output.n41 output.n15 289.615
R20280 output.n72 output.n46 289.615
R20281 output.n104 output.n78 289.615
R20282 output.n136 output.n110 289.615
R20283 output.n77 output.n45 197.26
R20284 output.n77 output.n76 196.298
R20285 output.n109 output.n108 196.298
R20286 output.n141 output.n140 196.298
R20287 output.n42 output.n41 185
R20288 output.n40 output.n39 185
R20289 output.n19 output.n18 185
R20290 output.n34 output.n33 185
R20291 output.n32 output.n31 185
R20292 output.n23 output.n22 185
R20293 output.n26 output.n25 185
R20294 output.n73 output.n72 185
R20295 output.n71 output.n70 185
R20296 output.n50 output.n49 185
R20297 output.n65 output.n64 185
R20298 output.n63 output.n62 185
R20299 output.n54 output.n53 185
R20300 output.n57 output.n56 185
R20301 output.n105 output.n104 185
R20302 output.n103 output.n102 185
R20303 output.n82 output.n81 185
R20304 output.n97 output.n96 185
R20305 output.n95 output.n94 185
R20306 output.n86 output.n85 185
R20307 output.n89 output.n88 185
R20308 output.n137 output.n136 185
R20309 output.n135 output.n134 185
R20310 output.n114 output.n113 185
R20311 output.n129 output.n128 185
R20312 output.n127 output.n126 185
R20313 output.n118 output.n117 185
R20314 output.n121 output.n120 185
R20315 output.t19 output.n24 147.661
R20316 output.t18 output.n55 147.661
R20317 output.t17 output.n87 147.661
R20318 output.t16 output.n119 147.661
R20319 output.n41 output.n40 104.615
R20320 output.n40 output.n18 104.615
R20321 output.n33 output.n18 104.615
R20322 output.n33 output.n32 104.615
R20323 output.n32 output.n22 104.615
R20324 output.n25 output.n22 104.615
R20325 output.n72 output.n71 104.615
R20326 output.n71 output.n49 104.615
R20327 output.n64 output.n49 104.615
R20328 output.n64 output.n63 104.615
R20329 output.n63 output.n53 104.615
R20330 output.n56 output.n53 104.615
R20331 output.n104 output.n103 104.615
R20332 output.n103 output.n81 104.615
R20333 output.n96 output.n81 104.615
R20334 output.n96 output.n95 104.615
R20335 output.n95 output.n85 104.615
R20336 output.n88 output.n85 104.615
R20337 output.n136 output.n135 104.615
R20338 output.n135 output.n113 104.615
R20339 output.n128 output.n113 104.615
R20340 output.n128 output.n127 104.615
R20341 output.n127 output.n117 104.615
R20342 output.n120 output.n117 104.615
R20343 output.n1 output.t15 77.056
R20344 output.n14 output.t0 76.6694
R20345 output.n1 output.n0 72.7095
R20346 output.n3 output.n2 72.7095
R20347 output.n5 output.n4 72.7095
R20348 output.n7 output.n6 72.7095
R20349 output.n9 output.n8 72.7095
R20350 output.n11 output.n10 72.7095
R20351 output.n13 output.n12 72.7095
R20352 output.n25 output.t19 52.3082
R20353 output.n56 output.t18 52.3082
R20354 output.n88 output.t17 52.3082
R20355 output.n120 output.t16 52.3082
R20356 output.n26 output.n24 15.6674
R20357 output.n57 output.n55 15.6674
R20358 output.n89 output.n87 15.6674
R20359 output.n121 output.n119 15.6674
R20360 output.n27 output.n23 12.8005
R20361 output.n58 output.n54 12.8005
R20362 output.n90 output.n86 12.8005
R20363 output.n122 output.n118 12.8005
R20364 output.n31 output.n30 12.0247
R20365 output.n62 output.n61 12.0247
R20366 output.n94 output.n93 12.0247
R20367 output.n126 output.n125 12.0247
R20368 output.n34 output.n21 11.249
R20369 output.n65 output.n52 11.249
R20370 output.n97 output.n84 11.249
R20371 output.n129 output.n116 11.249
R20372 output.n35 output.n19 10.4732
R20373 output.n66 output.n50 10.4732
R20374 output.n98 output.n82 10.4732
R20375 output.n130 output.n114 10.4732
R20376 output.n39 output.n38 9.69747
R20377 output.n70 output.n69 9.69747
R20378 output.n102 output.n101 9.69747
R20379 output.n134 output.n133 9.69747
R20380 output.n45 output.n44 9.45567
R20381 output.n76 output.n75 9.45567
R20382 output.n108 output.n107 9.45567
R20383 output.n140 output.n139 9.45567
R20384 output.n44 output.n43 9.3005
R20385 output.n17 output.n16 9.3005
R20386 output.n38 output.n37 9.3005
R20387 output.n36 output.n35 9.3005
R20388 output.n21 output.n20 9.3005
R20389 output.n30 output.n29 9.3005
R20390 output.n28 output.n27 9.3005
R20391 output.n75 output.n74 9.3005
R20392 output.n48 output.n47 9.3005
R20393 output.n69 output.n68 9.3005
R20394 output.n67 output.n66 9.3005
R20395 output.n52 output.n51 9.3005
R20396 output.n61 output.n60 9.3005
R20397 output.n59 output.n58 9.3005
R20398 output.n107 output.n106 9.3005
R20399 output.n80 output.n79 9.3005
R20400 output.n101 output.n100 9.3005
R20401 output.n99 output.n98 9.3005
R20402 output.n84 output.n83 9.3005
R20403 output.n93 output.n92 9.3005
R20404 output.n91 output.n90 9.3005
R20405 output.n139 output.n138 9.3005
R20406 output.n112 output.n111 9.3005
R20407 output.n133 output.n132 9.3005
R20408 output.n131 output.n130 9.3005
R20409 output.n116 output.n115 9.3005
R20410 output.n125 output.n124 9.3005
R20411 output.n123 output.n122 9.3005
R20412 output.n42 output.n17 8.92171
R20413 output.n73 output.n48 8.92171
R20414 output.n105 output.n80 8.92171
R20415 output.n137 output.n112 8.92171
R20416 output output.n141 8.15037
R20417 output.n43 output.n15 8.14595
R20418 output.n74 output.n46 8.14595
R20419 output.n106 output.n78 8.14595
R20420 output.n138 output.n110 8.14595
R20421 output.n45 output.n15 5.81868
R20422 output.n76 output.n46 5.81868
R20423 output.n108 output.n78 5.81868
R20424 output.n140 output.n110 5.81868
R20425 output.n43 output.n42 5.04292
R20426 output.n74 output.n73 5.04292
R20427 output.n106 output.n105 5.04292
R20428 output.n138 output.n137 5.04292
R20429 output.n28 output.n24 4.38594
R20430 output.n59 output.n55 4.38594
R20431 output.n91 output.n87 4.38594
R20432 output.n123 output.n119 4.38594
R20433 output.n39 output.n17 4.26717
R20434 output.n70 output.n48 4.26717
R20435 output.n102 output.n80 4.26717
R20436 output.n134 output.n112 4.26717
R20437 output.n0 output.t5 3.9605
R20438 output.n0 output.t9 3.9605
R20439 output.n2 output.t12 3.9605
R20440 output.n2 output.t1 3.9605
R20441 output.n4 output.t2 3.9605
R20442 output.n4 output.t7 3.9605
R20443 output.n6 output.t11 3.9605
R20444 output.n6 output.t3 3.9605
R20445 output.n8 output.t6 3.9605
R20446 output.n8 output.t4 3.9605
R20447 output.n10 output.t10 3.9605
R20448 output.n10 output.t13 3.9605
R20449 output.n12 output.t14 3.9605
R20450 output.n12 output.t8 3.9605
R20451 output.n38 output.n19 3.49141
R20452 output.n69 output.n50 3.49141
R20453 output.n101 output.n82 3.49141
R20454 output.n133 output.n114 3.49141
R20455 output.n35 output.n34 2.71565
R20456 output.n66 output.n65 2.71565
R20457 output.n98 output.n97 2.71565
R20458 output.n130 output.n129 2.71565
R20459 output.n31 output.n21 1.93989
R20460 output.n62 output.n52 1.93989
R20461 output.n94 output.n84 1.93989
R20462 output.n126 output.n116 1.93989
R20463 output.n30 output.n23 1.16414
R20464 output.n61 output.n54 1.16414
R20465 output.n93 output.n86 1.16414
R20466 output.n125 output.n118 1.16414
R20467 output.n141 output.n109 0.962709
R20468 output.n109 output.n77 0.962709
R20469 output.n27 output.n26 0.388379
R20470 output.n58 output.n57 0.388379
R20471 output.n90 output.n89 0.388379
R20472 output.n122 output.n121 0.388379
R20473 output.n14 output.n13 0.387128
R20474 output.n13 output.n11 0.387128
R20475 output.n11 output.n9 0.387128
R20476 output.n9 output.n7 0.387128
R20477 output.n7 output.n5 0.387128
R20478 output.n5 output.n3 0.387128
R20479 output.n3 output.n1 0.387128
R20480 output.n44 output.n16 0.155672
R20481 output.n37 output.n16 0.155672
R20482 output.n37 output.n36 0.155672
R20483 output.n36 output.n20 0.155672
R20484 output.n29 output.n20 0.155672
R20485 output.n29 output.n28 0.155672
R20486 output.n75 output.n47 0.155672
R20487 output.n68 output.n47 0.155672
R20488 output.n68 output.n67 0.155672
R20489 output.n67 output.n51 0.155672
R20490 output.n60 output.n51 0.155672
R20491 output.n60 output.n59 0.155672
R20492 output.n107 output.n79 0.155672
R20493 output.n100 output.n79 0.155672
R20494 output.n100 output.n99 0.155672
R20495 output.n99 output.n83 0.155672
R20496 output.n92 output.n83 0.155672
R20497 output.n92 output.n91 0.155672
R20498 output.n139 output.n111 0.155672
R20499 output.n132 output.n111 0.155672
R20500 output.n132 output.n131 0.155672
R20501 output.n131 output.n115 0.155672
R20502 output.n124 output.n115 0.155672
R20503 output.n124 output.n123 0.155672
R20504 output output.n14 0.126227
R20505 minus.n45 minus.t26 442.325
R20506 minus.n9 minus.t12 442.325
R20507 minus.n66 minus.t15 415.966
R20508 minus.n64 minus.t28 415.966
R20509 minus.n63 minus.t21 415.966
R20510 minus.n37 minus.t14 415.966
R20511 minus.n57 minus.t23 415.966
R20512 minus.n56 minus.t11 415.966
R20513 minus.n40 minus.t5 415.966
R20514 minus.n51 minus.t17 415.966
R20515 minus.n49 minus.t10 415.966
R20516 minus.n43 minus.t25 415.966
R20517 minus.n44 minus.t7 415.966
R20518 minus.n8 minus.t18 415.966
R20519 minus.n7 minus.t8 415.966
R20520 minus.n13 minus.t13 415.966
R20521 minus.n5 minus.t24 415.966
R20522 minus.n18 minus.t19 415.966
R20523 minus.n20 minus.t22 415.966
R20524 minus.n3 minus.t6 415.966
R20525 minus.n25 minus.t20 415.966
R20526 minus.n1 minus.t27 415.966
R20527 minus.n30 minus.t16 415.966
R20528 minus.n32 minus.t9 415.966
R20529 minus.n72 minus.t3 243.255
R20530 minus.n71 minus.n69 224.169
R20531 minus.n71 minus.n70 223.454
R20532 minus.n46 minus.n43 161.3
R20533 minus.n48 minus.n47 161.3
R20534 minus.n49 minus.n42 161.3
R20535 minus.n50 minus.n41 161.3
R20536 minus.n52 minus.n51 161.3
R20537 minus.n53 minus.n40 161.3
R20538 minus.n55 minus.n54 161.3
R20539 minus.n56 minus.n39 161.3
R20540 minus.n57 minus.n38 161.3
R20541 minus.n59 minus.n58 161.3
R20542 minus.n60 minus.n37 161.3
R20543 minus.n62 minus.n61 161.3
R20544 minus.n63 minus.n36 161.3
R20545 minus.n64 minus.n35 161.3
R20546 minus.n65 minus.n34 161.3
R20547 minus.n67 minus.n66 161.3
R20548 minus.n33 minus.n32 161.3
R20549 minus.n31 minus.n0 161.3
R20550 minus.n30 minus.n29 161.3
R20551 minus.n28 minus.n1 161.3
R20552 minus.n27 minus.n26 161.3
R20553 minus.n25 minus.n2 161.3
R20554 minus.n24 minus.n23 161.3
R20555 minus.n22 minus.n3 161.3
R20556 minus.n21 minus.n20 161.3
R20557 minus.n19 minus.n4 161.3
R20558 minus.n18 minus.n17 161.3
R20559 minus.n16 minus.n5 161.3
R20560 minus.n15 minus.n14 161.3
R20561 minus.n13 minus.n6 161.3
R20562 minus.n12 minus.n11 161.3
R20563 minus.n10 minus.n7 161.3
R20564 minus.n64 minus.n63 48.2005
R20565 minus.n57 minus.n56 48.2005
R20566 minus.n51 minus.n40 48.2005
R20567 minus.n44 minus.n43 48.2005
R20568 minus.n8 minus.n7 48.2005
R20569 minus.n18 minus.n5 48.2005
R20570 minus.n20 minus.n3 48.2005
R20571 minus.n30 minus.n1 48.2005
R20572 minus.n58 minus.n37 47.4702
R20573 minus.n50 minus.n49 47.4702
R20574 minus.n14 minus.n13 47.4702
R20575 minus.n25 minus.n24 47.4702
R20576 minus.n66 minus.n65 46.0096
R20577 minus.n32 minus.n31 46.0096
R20578 minus.n10 minus.n9 45.0871
R20579 minus.n46 minus.n45 45.0871
R20580 minus.n68 minus.n67 31.2713
R20581 minus.n62 minus.n37 25.5611
R20582 minus.n49 minus.n48 25.5611
R20583 minus.n13 minus.n12 25.5611
R20584 minus.n26 minus.n25 25.5611
R20585 minus.n56 minus.n55 24.1005
R20586 minus.n55 minus.n40 24.1005
R20587 minus.n19 minus.n18 24.1005
R20588 minus.n20 minus.n19 24.1005
R20589 minus.n63 minus.n62 22.6399
R20590 minus.n48 minus.n43 22.6399
R20591 minus.n12 minus.n7 22.6399
R20592 minus.n26 minus.n1 22.6399
R20593 minus.n70 minus.t2 19.8005
R20594 minus.n70 minus.t0 19.8005
R20595 minus.n69 minus.t1 19.8005
R20596 minus.n69 minus.t4 19.8005
R20597 minus.n45 minus.n44 14.1472
R20598 minus.n9 minus.n8 14.1472
R20599 minus.n68 minus.n33 11.9418
R20600 minus minus.n73 11.2412
R20601 minus.n73 minus.n72 4.80222
R20602 minus.n65 minus.n64 2.19141
R20603 minus.n31 minus.n30 2.19141
R20604 minus.n73 minus.n68 0.972091
R20605 minus.n58 minus.n57 0.730803
R20606 minus.n51 minus.n50 0.730803
R20607 minus.n14 minus.n5 0.730803
R20608 minus.n24 minus.n3 0.730803
R20609 minus.n72 minus.n71 0.716017
R20610 minus.n67 minus.n34 0.189894
R20611 minus.n35 minus.n34 0.189894
R20612 minus.n36 minus.n35 0.189894
R20613 minus.n61 minus.n36 0.189894
R20614 minus.n61 minus.n60 0.189894
R20615 minus.n60 minus.n59 0.189894
R20616 minus.n59 minus.n38 0.189894
R20617 minus.n39 minus.n38 0.189894
R20618 minus.n54 minus.n39 0.189894
R20619 minus.n54 minus.n53 0.189894
R20620 minus.n53 minus.n52 0.189894
R20621 minus.n52 minus.n41 0.189894
R20622 minus.n42 minus.n41 0.189894
R20623 minus.n47 minus.n42 0.189894
R20624 minus.n47 minus.n46 0.189894
R20625 minus.n11 minus.n10 0.189894
R20626 minus.n11 minus.n6 0.189894
R20627 minus.n15 minus.n6 0.189894
R20628 minus.n16 minus.n15 0.189894
R20629 minus.n17 minus.n16 0.189894
R20630 minus.n17 minus.n4 0.189894
R20631 minus.n21 minus.n4 0.189894
R20632 minus.n22 minus.n21 0.189894
R20633 minus.n23 minus.n22 0.189894
R20634 minus.n23 minus.n2 0.189894
R20635 minus.n27 minus.n2 0.189894
R20636 minus.n28 minus.n27 0.189894
R20637 minus.n29 minus.n28 0.189894
R20638 minus.n29 minus.n0 0.189894
R20639 minus.n33 minus.n0 0.189894
R20640 plus.n43 plus.t25 442.325
R20641 plus.n11 plus.t12 442.325
R20642 plus.n42 plus.t5 415.966
R20643 plus.n41 plus.t20 415.966
R20644 plus.n47 plus.t26 415.966
R20645 plus.n39 plus.t11 415.966
R20646 plus.n52 plus.t6 415.966
R20647 plus.n54 plus.t10 415.966
R20648 plus.n37 plus.t19 415.966
R20649 plus.n59 plus.t8 415.966
R20650 plus.n35 plus.t16 415.966
R20651 plus.n64 plus.t28 415.966
R20652 plus.n66 plus.t21 415.966
R20653 plus.n32 plus.t23 415.966
R20654 plus.n30 plus.t13 415.966
R20655 plus.n29 plus.t27 415.966
R20656 plus.n3 plus.t22 415.966
R20657 plus.n23 plus.t7 415.966
R20658 plus.n22 plus.t18 415.966
R20659 plus.n6 plus.t14 415.966
R20660 plus.n17 plus.t24 415.966
R20661 plus.n15 plus.t17 415.966
R20662 plus.n9 plus.t9 415.966
R20663 plus.n10 plus.t15 415.966
R20664 plus.n70 plus.t3 243.97
R20665 plus.n70 plus.n69 223.454
R20666 plus.n72 plus.n71 223.454
R20667 plus.n67 plus.n66 161.3
R20668 plus.n65 plus.n34 161.3
R20669 plus.n64 plus.n63 161.3
R20670 plus.n62 plus.n35 161.3
R20671 plus.n61 plus.n60 161.3
R20672 plus.n59 plus.n36 161.3
R20673 plus.n58 plus.n57 161.3
R20674 plus.n56 plus.n37 161.3
R20675 plus.n55 plus.n54 161.3
R20676 plus.n53 plus.n38 161.3
R20677 plus.n52 plus.n51 161.3
R20678 plus.n50 plus.n39 161.3
R20679 plus.n49 plus.n48 161.3
R20680 plus.n47 plus.n40 161.3
R20681 plus.n46 plus.n45 161.3
R20682 plus.n44 plus.n41 161.3
R20683 plus.n12 plus.n9 161.3
R20684 plus.n14 plus.n13 161.3
R20685 plus.n15 plus.n8 161.3
R20686 plus.n16 plus.n7 161.3
R20687 plus.n18 plus.n17 161.3
R20688 plus.n19 plus.n6 161.3
R20689 plus.n21 plus.n20 161.3
R20690 plus.n22 plus.n5 161.3
R20691 plus.n23 plus.n4 161.3
R20692 plus.n25 plus.n24 161.3
R20693 plus.n26 plus.n3 161.3
R20694 plus.n28 plus.n27 161.3
R20695 plus.n29 plus.n2 161.3
R20696 plus.n30 plus.n1 161.3
R20697 plus.n31 plus.n0 161.3
R20698 plus.n33 plus.n32 161.3
R20699 plus.n42 plus.n41 48.2005
R20700 plus.n52 plus.n39 48.2005
R20701 plus.n54 plus.n37 48.2005
R20702 plus.n64 plus.n35 48.2005
R20703 plus.n30 plus.n29 48.2005
R20704 plus.n23 plus.n22 48.2005
R20705 plus.n17 plus.n6 48.2005
R20706 plus.n10 plus.n9 48.2005
R20707 plus.n48 plus.n47 47.4702
R20708 plus.n59 plus.n58 47.4702
R20709 plus.n24 plus.n3 47.4702
R20710 plus.n16 plus.n15 47.4702
R20711 plus.n66 plus.n65 46.0096
R20712 plus.n32 plus.n31 46.0096
R20713 plus.n44 plus.n43 45.0871
R20714 plus.n12 plus.n11 45.0871
R20715 plus.n68 plus.n67 31.0554
R20716 plus.n47 plus.n46 25.5611
R20717 plus.n60 plus.n59 25.5611
R20718 plus.n28 plus.n3 25.5611
R20719 plus.n15 plus.n14 25.5611
R20720 plus.n53 plus.n52 24.1005
R20721 plus.n54 plus.n53 24.1005
R20722 plus.n22 plus.n21 24.1005
R20723 plus.n21 plus.n6 24.1005
R20724 plus.n46 plus.n41 22.6399
R20725 plus.n60 plus.n35 22.6399
R20726 plus.n29 plus.n28 22.6399
R20727 plus.n14 plus.n9 22.6399
R20728 plus.n69 plus.t4 19.8005
R20729 plus.n69 plus.t1 19.8005
R20730 plus.n71 plus.t0 19.8005
R20731 plus.n71 plus.t2 19.8005
R20732 plus.n43 plus.n42 14.1472
R20733 plus.n11 plus.n10 14.1472
R20734 plus plus.n73 14.0784
R20735 plus.n68 plus.n33 11.7259
R20736 plus.n73 plus.n72 5.40567
R20737 plus.n65 plus.n64 2.19141
R20738 plus.n31 plus.n30 2.19141
R20739 plus.n73 plus.n68 1.188
R20740 plus.n48 plus.n39 0.730803
R20741 plus.n58 plus.n37 0.730803
R20742 plus.n24 plus.n23 0.730803
R20743 plus.n17 plus.n16 0.730803
R20744 plus.n72 plus.n70 0.716017
R20745 plus.n45 plus.n44 0.189894
R20746 plus.n45 plus.n40 0.189894
R20747 plus.n49 plus.n40 0.189894
R20748 plus.n50 plus.n49 0.189894
R20749 plus.n51 plus.n50 0.189894
R20750 plus.n51 plus.n38 0.189894
R20751 plus.n55 plus.n38 0.189894
R20752 plus.n56 plus.n55 0.189894
R20753 plus.n57 plus.n56 0.189894
R20754 plus.n57 plus.n36 0.189894
R20755 plus.n61 plus.n36 0.189894
R20756 plus.n62 plus.n61 0.189894
R20757 plus.n63 plus.n62 0.189894
R20758 plus.n63 plus.n34 0.189894
R20759 plus.n67 plus.n34 0.189894
R20760 plus.n33 plus.n0 0.189894
R20761 plus.n1 plus.n0 0.189894
R20762 plus.n2 plus.n1 0.189894
R20763 plus.n27 plus.n2 0.189894
R20764 plus.n27 plus.n26 0.189894
R20765 plus.n26 plus.n25 0.189894
R20766 plus.n25 plus.n4 0.189894
R20767 plus.n5 plus.n4 0.189894
R20768 plus.n20 plus.n5 0.189894
R20769 plus.n20 plus.n19 0.189894
R20770 plus.n19 plus.n18 0.189894
R20771 plus.n18 plus.n7 0.189894
R20772 plus.n8 plus.n7 0.189894
R20773 plus.n13 plus.n8 0.189894
R20774 plus.n13 plus.n12 0.189894
R20775 a_n2903_n3924.n14 a_n2903_n3924.t27 214.994
R20776 a_n2903_n3924.n1 a_n2903_n3924.t30 214.493
R20777 a_n2903_n3924.n15 a_n2903_n3924.t55 214.321
R20778 a_n2903_n3924.n16 a_n2903_n3924.t29 214.321
R20779 a_n2903_n3924.n17 a_n2903_n3924.t28 214.321
R20780 a_n2903_n3924.n18 a_n2903_n3924.t0 214.321
R20781 a_n2903_n3924.n19 a_n2903_n3924.t1 214.321
R20782 a_n2903_n3924.n14 a_n2903_n3924.t26 214.321
R20783 a_n2903_n3924.n0 a_n2903_n3924.t5 55.8337
R20784 a_n2903_n3924.n2 a_n2903_n3924.t33 55.8337
R20785 a_n2903_n3924.n13 a_n2903_n3924.t44 55.8337
R20786 a_n2903_n3924.n47 a_n2903_n3924.t9 55.8335
R20787 a_n2903_n3924.n45 a_n2903_n3924.t50 55.8335
R20788 a_n2903_n3924.n34 a_n2903_n3924.t47 55.8335
R20789 a_n2903_n3924.n33 a_n2903_n3924.t18 55.8335
R20790 a_n2903_n3924.n22 a_n2903_n3924.t7 55.8335
R20791 a_n2903_n3924.n49 a_n2903_n3924.n48 53.0052
R20792 a_n2903_n3924.n51 a_n2903_n3924.n50 53.0052
R20793 a_n2903_n3924.n53 a_n2903_n3924.n52 53.0052
R20794 a_n2903_n3924.n55 a_n2903_n3924.n54 53.0052
R20795 a_n2903_n3924.n4 a_n2903_n3924.n3 53.0052
R20796 a_n2903_n3924.n6 a_n2903_n3924.n5 53.0052
R20797 a_n2903_n3924.n8 a_n2903_n3924.n7 53.0052
R20798 a_n2903_n3924.n10 a_n2903_n3924.n9 53.0052
R20799 a_n2903_n3924.n12 a_n2903_n3924.n11 53.0052
R20800 a_n2903_n3924.n44 a_n2903_n3924.n43 53.0051
R20801 a_n2903_n3924.n42 a_n2903_n3924.n41 53.0051
R20802 a_n2903_n3924.n40 a_n2903_n3924.n39 53.0051
R20803 a_n2903_n3924.n38 a_n2903_n3924.n37 53.0051
R20804 a_n2903_n3924.n36 a_n2903_n3924.n35 53.0051
R20805 a_n2903_n3924.n32 a_n2903_n3924.n31 53.0051
R20806 a_n2903_n3924.n30 a_n2903_n3924.n29 53.0051
R20807 a_n2903_n3924.n28 a_n2903_n3924.n27 53.0051
R20808 a_n2903_n3924.n26 a_n2903_n3924.n25 53.0051
R20809 a_n2903_n3924.n24 a_n2903_n3924.n23 53.0051
R20810 a_n2903_n3924.n57 a_n2903_n3924.n56 53.0051
R20811 a_n2903_n3924.n21 a_n2903_n3924.n13 12.1555
R20812 a_n2903_n3924.n47 a_n2903_n3924.n46 12.1555
R20813 a_n2903_n3924.n22 a_n2903_n3924.n21 5.07593
R20814 a_n2903_n3924.n46 a_n2903_n3924.n45 5.07593
R20815 a_n2903_n3924.n48 a_n2903_n3924.t14 2.82907
R20816 a_n2903_n3924.n48 a_n2903_n3924.t2 2.82907
R20817 a_n2903_n3924.n50 a_n2903_n3924.t11 2.82907
R20818 a_n2903_n3924.n50 a_n2903_n3924.t22 2.82907
R20819 a_n2903_n3924.n52 a_n2903_n3924.t24 2.82907
R20820 a_n2903_n3924.n52 a_n2903_n3924.t20 2.82907
R20821 a_n2903_n3924.n54 a_n2903_n3924.t4 2.82907
R20822 a_n2903_n3924.n54 a_n2903_n3924.t19 2.82907
R20823 a_n2903_n3924.n3 a_n2903_n3924.t34 2.82907
R20824 a_n2903_n3924.n3 a_n2903_n3924.t52 2.82907
R20825 a_n2903_n3924.n5 a_n2903_n3924.t42 2.82907
R20826 a_n2903_n3924.n5 a_n2903_n3924.t49 2.82907
R20827 a_n2903_n3924.n7 a_n2903_n3924.t48 2.82907
R20828 a_n2903_n3924.n7 a_n2903_n3924.t54 2.82907
R20829 a_n2903_n3924.n9 a_n2903_n3924.t45 2.82907
R20830 a_n2903_n3924.n9 a_n2903_n3924.t36 2.82907
R20831 a_n2903_n3924.n11 a_n2903_n3924.t31 2.82907
R20832 a_n2903_n3924.n11 a_n2903_n3924.t38 2.82907
R20833 a_n2903_n3924.n43 a_n2903_n3924.t32 2.82907
R20834 a_n2903_n3924.n43 a_n2903_n3924.t43 2.82907
R20835 a_n2903_n3924.n41 a_n2903_n3924.t53 2.82907
R20836 a_n2903_n3924.n41 a_n2903_n3924.t39 2.82907
R20837 a_n2903_n3924.n39 a_n2903_n3924.t40 2.82907
R20838 a_n2903_n3924.n39 a_n2903_n3924.t37 2.82907
R20839 a_n2903_n3924.n37 a_n2903_n3924.t46 2.82907
R20840 a_n2903_n3924.n37 a_n2903_n3924.t35 2.82907
R20841 a_n2903_n3924.n35 a_n2903_n3924.t41 2.82907
R20842 a_n2903_n3924.n35 a_n2903_n3924.t51 2.82907
R20843 a_n2903_n3924.n31 a_n2903_n3924.t21 2.82907
R20844 a_n2903_n3924.n31 a_n2903_n3924.t15 2.82907
R20845 a_n2903_n3924.n29 a_n2903_n3924.t6 2.82907
R20846 a_n2903_n3924.n29 a_n2903_n3924.t13 2.82907
R20847 a_n2903_n3924.n27 a_n2903_n3924.t12 2.82907
R20848 a_n2903_n3924.n27 a_n2903_n3924.t16 2.82907
R20849 a_n2903_n3924.n25 a_n2903_n3924.t8 2.82907
R20850 a_n2903_n3924.n25 a_n2903_n3924.t23 2.82907
R20851 a_n2903_n3924.n23 a_n2903_n3924.t17 2.82907
R20852 a_n2903_n3924.n23 a_n2903_n3924.t3 2.82907
R20853 a_n2903_n3924.t25 a_n2903_n3924.n57 2.82907
R20854 a_n2903_n3924.n57 a_n2903_n3924.t10 2.82907
R20855 a_n2903_n3924.n46 a_n2903_n3924.n1 1.95694
R20856 a_n2903_n3924.n21 a_n2903_n3924.n20 1.95694
R20857 a_n2903_n3924.n19 a_n2903_n3924.n18 0.672012
R20858 a_n2903_n3924.n18 a_n2903_n3924.n17 0.672012
R20859 a_n2903_n3924.n17 a_n2903_n3924.n16 0.672012
R20860 a_n2903_n3924.n16 a_n2903_n3924.n15 0.672012
R20861 a_n2903_n3924.n20 a_n2903_n3924.n19 0.643669
R20862 a_n2903_n3924.n15 a_n2903_n3924.n1 0.501227
R20863 a_n2903_n3924.n24 a_n2903_n3924.n22 0.358259
R20864 a_n2903_n3924.n26 a_n2903_n3924.n24 0.358259
R20865 a_n2903_n3924.n28 a_n2903_n3924.n26 0.358259
R20866 a_n2903_n3924.n30 a_n2903_n3924.n28 0.358259
R20867 a_n2903_n3924.n32 a_n2903_n3924.n30 0.358259
R20868 a_n2903_n3924.n33 a_n2903_n3924.n32 0.358259
R20869 a_n2903_n3924.n36 a_n2903_n3924.n34 0.358259
R20870 a_n2903_n3924.n38 a_n2903_n3924.n36 0.358259
R20871 a_n2903_n3924.n40 a_n2903_n3924.n38 0.358259
R20872 a_n2903_n3924.n42 a_n2903_n3924.n40 0.358259
R20873 a_n2903_n3924.n44 a_n2903_n3924.n42 0.358259
R20874 a_n2903_n3924.n45 a_n2903_n3924.n44 0.358259
R20875 a_n2903_n3924.n13 a_n2903_n3924.n12 0.358259
R20876 a_n2903_n3924.n12 a_n2903_n3924.n10 0.358259
R20877 a_n2903_n3924.n10 a_n2903_n3924.n8 0.358259
R20878 a_n2903_n3924.n8 a_n2903_n3924.n6 0.358259
R20879 a_n2903_n3924.n6 a_n2903_n3924.n4 0.358259
R20880 a_n2903_n3924.n4 a_n2903_n3924.n2 0.358259
R20881 a_n2903_n3924.n56 a_n2903_n3924.n0 0.358259
R20882 a_n2903_n3924.n56 a_n2903_n3924.n55 0.358259
R20883 a_n2903_n3924.n55 a_n2903_n3924.n53 0.358259
R20884 a_n2903_n3924.n53 a_n2903_n3924.n51 0.358259
R20885 a_n2903_n3924.n51 a_n2903_n3924.n49 0.358259
R20886 a_n2903_n3924.n49 a_n2903_n3924.n47 0.358259
R20887 a_n2903_n3924.n34 a_n2903_n3924.n33 0.235414
R20888 a_n2903_n3924.n2 a_n2903_n3924.n0 0.235414
R20889 a_n2903_n3924.n20 a_n2903_n3924.n14 0.028843
R20890 diffpairibias.n0 diffpairibias.t18 436.822
R20891 diffpairibias.n21 diffpairibias.t19 435.479
R20892 diffpairibias.n20 diffpairibias.t16 435.479
R20893 diffpairibias.n19 diffpairibias.t17 435.479
R20894 diffpairibias.n18 diffpairibias.t21 435.479
R20895 diffpairibias.n0 diffpairibias.t22 435.479
R20896 diffpairibias.n1 diffpairibias.t20 435.479
R20897 diffpairibias.n2 diffpairibias.t23 435.479
R20898 diffpairibias.n10 diffpairibias.t0 377.536
R20899 diffpairibias.n10 diffpairibias.t8 376.193
R20900 diffpairibias.n11 diffpairibias.t10 376.193
R20901 diffpairibias.n12 diffpairibias.t6 376.193
R20902 diffpairibias.n13 diffpairibias.t2 376.193
R20903 diffpairibias.n14 diffpairibias.t12 376.193
R20904 diffpairibias.n15 diffpairibias.t4 376.193
R20905 diffpairibias.n16 diffpairibias.t14 376.193
R20906 diffpairibias.n3 diffpairibias.t1 113.368
R20907 diffpairibias.n3 diffpairibias.t9 112.698
R20908 diffpairibias.n4 diffpairibias.t11 112.698
R20909 diffpairibias.n5 diffpairibias.t7 112.698
R20910 diffpairibias.n6 diffpairibias.t3 112.698
R20911 diffpairibias.n7 diffpairibias.t13 112.698
R20912 diffpairibias.n8 diffpairibias.t5 112.698
R20913 diffpairibias.n9 diffpairibias.t15 112.698
R20914 diffpairibias.n17 diffpairibias.n16 4.77242
R20915 diffpairibias.n17 diffpairibias.n9 4.30807
R20916 diffpairibias.n18 diffpairibias.n17 4.13945
R20917 diffpairibias.n16 diffpairibias.n15 1.34352
R20918 diffpairibias.n15 diffpairibias.n14 1.34352
R20919 diffpairibias.n14 diffpairibias.n13 1.34352
R20920 diffpairibias.n13 diffpairibias.n12 1.34352
R20921 diffpairibias.n12 diffpairibias.n11 1.34352
R20922 diffpairibias.n11 diffpairibias.n10 1.34352
R20923 diffpairibias.n2 diffpairibias.n1 1.34352
R20924 diffpairibias.n1 diffpairibias.n0 1.34352
R20925 diffpairibias.n19 diffpairibias.n18 1.34352
R20926 diffpairibias.n20 diffpairibias.n19 1.34352
R20927 diffpairibias.n21 diffpairibias.n20 1.34352
R20928 diffpairibias.n22 diffpairibias.n21 0.862419
R20929 diffpairibias diffpairibias.n22 0.684875
R20930 diffpairibias.n9 diffpairibias.n8 0.672012
R20931 diffpairibias.n8 diffpairibias.n7 0.672012
R20932 diffpairibias.n7 diffpairibias.n6 0.672012
R20933 diffpairibias.n6 diffpairibias.n5 0.672012
R20934 diffpairibias.n5 diffpairibias.n4 0.672012
R20935 diffpairibias.n4 diffpairibias.n3 0.672012
R20936 diffpairibias.n22 diffpairibias.n2 0.190907
C0 minus diffpairibias 2.98e-19
C1 commonsourceibias output 0.006808f
C2 CSoutput minus 2.51572f
C3 vdd plus 0.073313f
C4 commonsourceibias outputibias 0.003832f
C5 plus diffpairibias 2.75e-19
C6 vdd commonsourceibias 0.004218f
C7 CSoutput plus 0.834874f
C8 commonsourceibias diffpairibias 0.052851f
C9 CSoutput commonsourceibias 29.0223f
C10 minus plus 8.7598f
C11 minus commonsourceibias 0.322616f
C12 plus commonsourceibias 0.276969f
C13 output outputibias 2.34152f
C14 vdd output 7.23429f
C15 CSoutput output 6.13571f
C16 CSoutput outputibias 0.032386f
C17 vdd CSoutput 91.981f
C18 diffpairibias gnd 48.968437f
C19 outputibias gnd 32.465668f
C20 output gnd 15.47879f
C21 commonsourceibias gnd 0.118808p
C22 plus gnd 32.3879f
C23 minus gnd 26.34968f
C24 CSoutput gnd 88.49096f
C25 vdd gnd 0.376956p
C26 diffpairibias.t18 gnd 0.087401f
C27 diffpairibias.t22 gnd 0.087239f
C28 diffpairibias.n0 gnd 0.102784f
C29 diffpairibias.t20 gnd 0.087239f
C30 diffpairibias.n1 gnd 0.050171f
C31 diffpairibias.t23 gnd 0.087239f
C32 diffpairibias.n2 gnd 0.039841f
C33 diffpairibias.t1 gnd 0.083757f
C34 diffpairibias.t9 gnd 0.083392f
C35 diffpairibias.n3 gnd 0.131682f
C36 diffpairibias.t11 gnd 0.083392f
C37 diffpairibias.n4 gnd 0.07027f
C38 diffpairibias.t7 gnd 0.083392f
C39 diffpairibias.n5 gnd 0.07027f
C40 diffpairibias.t3 gnd 0.083392f
C41 diffpairibias.n6 gnd 0.07027f
C42 diffpairibias.t13 gnd 0.083392f
C43 diffpairibias.n7 gnd 0.07027f
C44 diffpairibias.t5 gnd 0.083392f
C45 diffpairibias.n8 gnd 0.07027f
C46 diffpairibias.t15 gnd 0.083392f
C47 diffpairibias.n9 gnd 0.099771f
C48 diffpairibias.t0 gnd 0.08427f
C49 diffpairibias.t8 gnd 0.084123f
C50 diffpairibias.n10 gnd 0.091784f
C51 diffpairibias.t10 gnd 0.084123f
C52 diffpairibias.n11 gnd 0.050681f
C53 diffpairibias.t6 gnd 0.084123f
C54 diffpairibias.n12 gnd 0.050681f
C55 diffpairibias.t2 gnd 0.084123f
C56 diffpairibias.n13 gnd 0.050681f
C57 diffpairibias.t12 gnd 0.084123f
C58 diffpairibias.n14 gnd 0.050681f
C59 diffpairibias.t4 gnd 0.084123f
C60 diffpairibias.n15 gnd 0.050681f
C61 diffpairibias.t14 gnd 0.084123f
C62 diffpairibias.n16 gnd 0.059977f
C63 diffpairibias.n17 gnd 0.226448f
C64 diffpairibias.t21 gnd 0.087239f
C65 diffpairibias.n18 gnd 0.050181f
C66 diffpairibias.t17 gnd 0.087239f
C67 diffpairibias.n19 gnd 0.050171f
C68 diffpairibias.t16 gnd 0.087239f
C69 diffpairibias.n20 gnd 0.050171f
C70 diffpairibias.t19 gnd 0.087239f
C71 diffpairibias.n21 gnd 0.045859f
C72 diffpairibias.n22 gnd 0.046268f
C73 a_n2903_n3924.t10 gnd 0.108618f
C74 a_n2903_n3924.t5 gnd 1.12888f
C75 a_n2903_n3924.n0 gnd 0.383133f
C76 a_n2903_n3924.t30 gnd 1.40337f
C77 a_n2903_n3924.n1 gnd 1.48426f
C78 a_n2903_n3924.t33 gnd 1.12888f
C79 a_n2903_n3924.n2 gnd 0.383133f
C80 a_n2903_n3924.t34 gnd 0.108618f
C81 a_n2903_n3924.t52 gnd 0.108618f
C82 a_n2903_n3924.n3 gnd 0.887099f
C83 a_n2903_n3924.n4 gnd 0.359777f
C84 a_n2903_n3924.t42 gnd 0.108618f
C85 a_n2903_n3924.t49 gnd 0.108618f
C86 a_n2903_n3924.n5 gnd 0.887099f
C87 a_n2903_n3924.n6 gnd 0.359777f
C88 a_n2903_n3924.t48 gnd 0.108618f
C89 a_n2903_n3924.t54 gnd 0.108618f
C90 a_n2903_n3924.n7 gnd 0.887099f
C91 a_n2903_n3924.n8 gnd 0.359777f
C92 a_n2903_n3924.t45 gnd 0.108618f
C93 a_n2903_n3924.t36 gnd 0.108618f
C94 a_n2903_n3924.n9 gnd 0.887099f
C95 a_n2903_n3924.n10 gnd 0.359777f
C96 a_n2903_n3924.t31 gnd 0.108618f
C97 a_n2903_n3924.t38 gnd 0.108618f
C98 a_n2903_n3924.n11 gnd 0.887099f
C99 a_n2903_n3924.n12 gnd 0.359777f
C100 a_n2903_n3924.t44 gnd 1.12888f
C101 a_n2903_n3924.n13 gnd 0.974186f
C102 a_n2903_n3924.t27 gnd 1.40461f
C103 a_n2903_n3924.t26 gnd 1.40261f
C104 a_n2903_n3924.n14 gnd 1.26893f
C105 a_n2903_n3924.t55 gnd 1.40261f
C106 a_n2903_n3924.n15 gnd 0.892855f
C107 a_n2903_n3924.t29 gnd 1.40261f
C108 a_n2903_n3924.n16 gnd 0.987884f
C109 a_n2903_n3924.t28 gnd 1.40261f
C110 a_n2903_n3924.n17 gnd 0.987884f
C111 a_n2903_n3924.t0 gnd 1.40261f
C112 a_n2903_n3924.n18 gnd 0.987884f
C113 a_n2903_n3924.t1 gnd 1.40261f
C114 a_n2903_n3924.n19 gnd 0.972113f
C115 a_n2903_n3924.n20 gnd 0.533935f
C116 a_n2903_n3924.n21 gnd 1.01395f
C117 a_n2903_n3924.t7 gnd 1.12888f
C118 a_n2903_n3924.n22 gnd 0.619233f
C119 a_n2903_n3924.t17 gnd 0.108618f
C120 a_n2903_n3924.t3 gnd 0.108618f
C121 a_n2903_n3924.n23 gnd 0.887098f
C122 a_n2903_n3924.n24 gnd 0.359779f
C123 a_n2903_n3924.t8 gnd 0.108618f
C124 a_n2903_n3924.t23 gnd 0.108618f
C125 a_n2903_n3924.n25 gnd 0.887098f
C126 a_n2903_n3924.n26 gnd 0.359779f
C127 a_n2903_n3924.t12 gnd 0.108618f
C128 a_n2903_n3924.t16 gnd 0.108618f
C129 a_n2903_n3924.n27 gnd 0.887098f
C130 a_n2903_n3924.n28 gnd 0.359779f
C131 a_n2903_n3924.t6 gnd 0.108618f
C132 a_n2903_n3924.t13 gnd 0.108618f
C133 a_n2903_n3924.n29 gnd 0.887098f
C134 a_n2903_n3924.n30 gnd 0.359779f
C135 a_n2903_n3924.t21 gnd 0.108618f
C136 a_n2903_n3924.t15 gnd 0.108618f
C137 a_n2903_n3924.n31 gnd 0.887098f
C138 a_n2903_n3924.n32 gnd 0.359779f
C139 a_n2903_n3924.t18 gnd 1.12888f
C140 a_n2903_n3924.n33 gnd 0.383138f
C141 a_n2903_n3924.t47 gnd 1.12888f
C142 a_n2903_n3924.n34 gnd 0.383138f
C143 a_n2903_n3924.t41 gnd 0.108618f
C144 a_n2903_n3924.t51 gnd 0.108618f
C145 a_n2903_n3924.n35 gnd 0.887098f
C146 a_n2903_n3924.n36 gnd 0.359779f
C147 a_n2903_n3924.t46 gnd 0.108618f
C148 a_n2903_n3924.t35 gnd 0.108618f
C149 a_n2903_n3924.n37 gnd 0.887098f
C150 a_n2903_n3924.n38 gnd 0.359779f
C151 a_n2903_n3924.t40 gnd 0.108618f
C152 a_n2903_n3924.t37 gnd 0.108618f
C153 a_n2903_n3924.n39 gnd 0.887098f
C154 a_n2903_n3924.n40 gnd 0.359779f
C155 a_n2903_n3924.t53 gnd 0.108618f
C156 a_n2903_n3924.t39 gnd 0.108618f
C157 a_n2903_n3924.n41 gnd 0.887098f
C158 a_n2903_n3924.n42 gnd 0.359779f
C159 a_n2903_n3924.t32 gnd 0.108618f
C160 a_n2903_n3924.t43 gnd 0.108618f
C161 a_n2903_n3924.n43 gnd 0.887098f
C162 a_n2903_n3924.n44 gnd 0.359779f
C163 a_n2903_n3924.t50 gnd 1.12888f
C164 a_n2903_n3924.n45 gnd 0.619233f
C165 a_n2903_n3924.n46 gnd 1.01395f
C166 a_n2903_n3924.t9 gnd 1.12888f
C167 a_n2903_n3924.n47 gnd 0.97419f
C168 a_n2903_n3924.t14 gnd 0.108618f
C169 a_n2903_n3924.t2 gnd 0.108618f
C170 a_n2903_n3924.n48 gnd 0.887099f
C171 a_n2903_n3924.n49 gnd 0.359777f
C172 a_n2903_n3924.t11 gnd 0.108618f
C173 a_n2903_n3924.t22 gnd 0.108618f
C174 a_n2903_n3924.n50 gnd 0.887099f
C175 a_n2903_n3924.n51 gnd 0.359777f
C176 a_n2903_n3924.t24 gnd 0.108618f
C177 a_n2903_n3924.t20 gnd 0.108618f
C178 a_n2903_n3924.n52 gnd 0.887099f
C179 a_n2903_n3924.n53 gnd 0.359777f
C180 a_n2903_n3924.t4 gnd 0.108618f
C181 a_n2903_n3924.t19 gnd 0.108618f
C182 a_n2903_n3924.n54 gnd 0.887099f
C183 a_n2903_n3924.n55 gnd 0.359777f
C184 a_n2903_n3924.n56 gnd 0.359776f
C185 a_n2903_n3924.n57 gnd 0.887101f
C186 a_n2903_n3924.t25 gnd 0.108618f
C187 plus.n0 gnd 0.024493f
C188 plus.t23 gnd 0.247447f
C189 plus.n1 gnd 0.024493f
C190 plus.t13 gnd 0.247447f
C191 plus.n2 gnd 0.024493f
C192 plus.t27 gnd 0.247447f
C193 plus.t22 gnd 0.247447f
C194 plus.n3 gnd 0.114403f
C195 plus.n4 gnd 0.024493f
C196 plus.t7 gnd 0.247447f
C197 plus.n5 gnd 0.024493f
C198 plus.t18 gnd 0.247447f
C199 plus.t14 gnd 0.247447f
C200 plus.n6 gnd 0.114327f
C201 plus.n7 gnd 0.024493f
C202 plus.t24 gnd 0.247447f
C203 plus.n8 gnd 0.024493f
C204 plus.t17 gnd 0.247447f
C205 plus.t9 gnd 0.247447f
C206 plus.n9 gnd 0.114176f
C207 plus.t12 gnd 0.254109f
C208 plus.t15 gnd 0.247447f
C209 plus.n10 gnd 0.117074f
C210 plus.n11 gnd 0.105976f
C211 plus.n12 gnd 0.09945f
C212 plus.n13 gnd 0.024493f
C213 plus.n14 gnd 0.005558f
C214 plus.n15 gnd 0.114403f
C215 plus.n16 gnd 0.005558f
C216 plus.n17 gnd 0.111911f
C217 plus.n18 gnd 0.024493f
C218 plus.n19 gnd 0.024493f
C219 plus.n20 gnd 0.024493f
C220 plus.n21 gnd 0.005558f
C221 plus.n22 gnd 0.114327f
C222 plus.n23 gnd 0.111911f
C223 plus.n24 gnd 0.005558f
C224 plus.n25 gnd 0.024493f
C225 plus.n26 gnd 0.024493f
C226 plus.n27 gnd 0.024493f
C227 plus.n28 gnd 0.005558f
C228 plus.n29 gnd 0.114176f
C229 plus.n30 gnd 0.112062f
C230 plus.n31 gnd 0.005558f
C231 plus.n32 gnd 0.111609f
C232 plus.n33 gnd 0.268547f
C233 plus.n34 gnd 0.024493f
C234 plus.t16 gnd 0.247447f
C235 plus.n35 gnd 0.114176f
C236 plus.t28 gnd 0.247447f
C237 plus.n36 gnd 0.024493f
C238 plus.t19 gnd 0.247447f
C239 plus.n37 gnd 0.111911f
C240 plus.n38 gnd 0.024493f
C241 plus.t11 gnd 0.247447f
C242 plus.n39 gnd 0.111911f
C243 plus.t6 gnd 0.247447f
C244 plus.n40 gnd 0.024493f
C245 plus.t20 gnd 0.247447f
C246 plus.n41 gnd 0.114176f
C247 plus.t25 gnd 0.254109f
C248 plus.t5 gnd 0.247447f
C249 plus.n42 gnd 0.117074f
C250 plus.n43 gnd 0.105976f
C251 plus.n44 gnd 0.09945f
C252 plus.n45 gnd 0.024493f
C253 plus.n46 gnd 0.005558f
C254 plus.t26 gnd 0.247447f
C255 plus.n47 gnd 0.114403f
C256 plus.n48 gnd 0.005558f
C257 plus.n49 gnd 0.024493f
C258 plus.n50 gnd 0.024493f
C259 plus.n51 gnd 0.024493f
C260 plus.n52 gnd 0.114327f
C261 plus.n53 gnd 0.005558f
C262 plus.t10 gnd 0.247447f
C263 plus.n54 gnd 0.114327f
C264 plus.n55 gnd 0.024493f
C265 plus.n56 gnd 0.024493f
C266 plus.n57 gnd 0.024493f
C267 plus.n58 gnd 0.005558f
C268 plus.t8 gnd 0.247447f
C269 plus.n59 gnd 0.114403f
C270 plus.n60 gnd 0.005558f
C271 plus.n61 gnd 0.024493f
C272 plus.n62 gnd 0.024493f
C273 plus.n63 gnd 0.024493f
C274 plus.n64 gnd 0.112062f
C275 plus.n65 gnd 0.005558f
C276 plus.t21 gnd 0.247447f
C277 plus.n66 gnd 0.111609f
C278 plus.n67 gnd 0.733391f
C279 plus.n68 gnd 1.11778f
C280 plus.t3 gnd 0.042281f
C281 plus.t4 gnd 0.00755f
C282 plus.t1 gnd 0.00755f
C283 plus.n69 gnd 0.024487f
C284 plus.n70 gnd 0.190096f
C285 plus.t0 gnd 0.00755f
C286 plus.t2 gnd 0.00755f
C287 plus.n71 gnd 0.024487f
C288 plus.n72 gnd 0.14269f
C289 plus.n73 gnd 2.50198f
C290 minus.n0 gnd 0.033787f
C291 minus.t27 gnd 0.341345f
C292 minus.n1 gnd 0.157502f
C293 minus.n2 gnd 0.033787f
C294 minus.t6 gnd 0.341345f
C295 minus.n3 gnd 0.154377f
C296 minus.n4 gnd 0.033787f
C297 minus.t24 gnd 0.341345f
C298 minus.n5 gnd 0.154377f
C299 minus.n6 gnd 0.033787f
C300 minus.t8 gnd 0.341345f
C301 minus.n7 gnd 0.157502f
C302 minus.t12 gnd 0.350535f
C303 minus.t18 gnd 0.341345f
C304 minus.n8 gnd 0.1615f
C305 minus.n9 gnd 0.14619f
C306 minus.n10 gnd 0.137189f
C307 minus.n11 gnd 0.033787f
C308 minus.n12 gnd 0.007667f
C309 minus.t13 gnd 0.341345f
C310 minus.n13 gnd 0.157815f
C311 minus.n14 gnd 0.007667f
C312 minus.n15 gnd 0.033787f
C313 minus.n16 gnd 0.033787f
C314 minus.n17 gnd 0.033787f
C315 minus.t19 gnd 0.341345f
C316 minus.n18 gnd 0.15771f
C317 minus.n19 gnd 0.007667f
C318 minus.t22 gnd 0.341345f
C319 minus.n20 gnd 0.15771f
C320 minus.n21 gnd 0.033787f
C321 minus.n22 gnd 0.033787f
C322 minus.n23 gnd 0.033787f
C323 minus.n24 gnd 0.007667f
C324 minus.t20 gnd 0.341345f
C325 minus.n25 gnd 0.157815f
C326 minus.n26 gnd 0.007667f
C327 minus.n27 gnd 0.033787f
C328 minus.n28 gnd 0.033787f
C329 minus.n29 gnd 0.033787f
C330 minus.t16 gnd 0.341345f
C331 minus.n30 gnd 0.154586f
C332 minus.n31 gnd 0.007667f
C333 minus.t9 gnd 0.341345f
C334 minus.n32 gnd 0.153961f
C335 minus.n33 gnd 0.379182f
C336 minus.n34 gnd 0.033787f
C337 minus.t15 gnd 0.341345f
C338 minus.t28 gnd 0.341345f
C339 minus.n35 gnd 0.033787f
C340 minus.t21 gnd 0.341345f
C341 minus.n36 gnd 0.033787f
C342 minus.t14 gnd 0.341345f
C343 minus.n37 gnd 0.157815f
C344 minus.n38 gnd 0.033787f
C345 minus.t23 gnd 0.341345f
C346 minus.t11 gnd 0.341345f
C347 minus.n39 gnd 0.033787f
C348 minus.t5 gnd 0.341345f
C349 minus.n40 gnd 0.15771f
C350 minus.n41 gnd 0.033787f
C351 minus.t17 gnd 0.341345f
C352 minus.t10 gnd 0.341345f
C353 minus.n42 gnd 0.033787f
C354 minus.t25 gnd 0.341345f
C355 minus.n43 gnd 0.157502f
C356 minus.t26 gnd 0.350535f
C357 minus.t7 gnd 0.341345f
C358 minus.n44 gnd 0.1615f
C359 minus.n45 gnd 0.14619f
C360 minus.n46 gnd 0.137189f
C361 minus.n47 gnd 0.033787f
C362 minus.n48 gnd 0.007667f
C363 minus.n49 gnd 0.157815f
C364 minus.n50 gnd 0.007667f
C365 minus.n51 gnd 0.154377f
C366 minus.n52 gnd 0.033787f
C367 minus.n53 gnd 0.033787f
C368 minus.n54 gnd 0.033787f
C369 minus.n55 gnd 0.007667f
C370 minus.n56 gnd 0.15771f
C371 minus.n57 gnd 0.154377f
C372 minus.n58 gnd 0.007667f
C373 minus.n59 gnd 0.033787f
C374 minus.n60 gnd 0.033787f
C375 minus.n61 gnd 0.033787f
C376 minus.n62 gnd 0.007667f
C377 minus.n63 gnd 0.157502f
C378 minus.n64 gnd 0.154586f
C379 minus.n65 gnd 0.007667f
C380 minus.n66 gnd 0.153961f
C381 minus.n67 gnd 1.02527f
C382 minus.n68 gnd 1.55525f
C383 minus.t1 gnd 0.010415f
C384 minus.t4 gnd 0.010415f
C385 minus.n69 gnd 0.034249f
C386 minus.t2 gnd 0.010415f
C387 minus.t0 gnd 0.010415f
C388 minus.n70 gnd 0.033779f
C389 minus.n71 gnd 0.28829f
C390 minus.t3 gnd 0.057971f
C391 minus.n72 gnd 0.157317f
C392 minus.n73 gnd 1.91669f
C393 output.t15 gnd 0.464308f
C394 output.t5 gnd 0.044422f
C395 output.t9 gnd 0.044422f
C396 output.n0 gnd 0.364624f
C397 output.n1 gnd 0.614102f
C398 output.t12 gnd 0.044422f
C399 output.t1 gnd 0.044422f
C400 output.n2 gnd 0.364624f
C401 output.n3 gnd 0.350265f
C402 output.t2 gnd 0.044422f
C403 output.t7 gnd 0.044422f
C404 output.n4 gnd 0.364624f
C405 output.n5 gnd 0.350265f
C406 output.t11 gnd 0.044422f
C407 output.t3 gnd 0.044422f
C408 output.n6 gnd 0.364624f
C409 output.n7 gnd 0.350265f
C410 output.t6 gnd 0.044422f
C411 output.t4 gnd 0.044422f
C412 output.n8 gnd 0.364624f
C413 output.n9 gnd 0.350265f
C414 output.t10 gnd 0.044422f
C415 output.t13 gnd 0.044422f
C416 output.n10 gnd 0.364624f
C417 output.n11 gnd 0.350265f
C418 output.t14 gnd 0.044422f
C419 output.t8 gnd 0.044422f
C420 output.n12 gnd 0.364624f
C421 output.n13 gnd 0.350265f
C422 output.t0 gnd 0.462979f
C423 output.n14 gnd 0.28994f
C424 output.n15 gnd 0.015803f
C425 output.n16 gnd 0.011243f
C426 output.n17 gnd 0.006041f
C427 output.n18 gnd 0.01428f
C428 output.n19 gnd 0.006397f
C429 output.n20 gnd 0.011243f
C430 output.n21 gnd 0.006041f
C431 output.n22 gnd 0.01428f
C432 output.n23 gnd 0.006397f
C433 output.n24 gnd 0.048111f
C434 output.t19 gnd 0.023274f
C435 output.n25 gnd 0.01071f
C436 output.n26 gnd 0.008435f
C437 output.n27 gnd 0.006041f
C438 output.n28 gnd 0.267512f
C439 output.n29 gnd 0.011243f
C440 output.n30 gnd 0.006041f
C441 output.n31 gnd 0.006397f
C442 output.n32 gnd 0.01428f
C443 output.n33 gnd 0.01428f
C444 output.n34 gnd 0.006397f
C445 output.n35 gnd 0.006041f
C446 output.n36 gnd 0.011243f
C447 output.n37 gnd 0.011243f
C448 output.n38 gnd 0.006041f
C449 output.n39 gnd 0.006397f
C450 output.n40 gnd 0.01428f
C451 output.n41 gnd 0.030913f
C452 output.n42 gnd 0.006397f
C453 output.n43 gnd 0.006041f
C454 output.n44 gnd 0.025987f
C455 output.n45 gnd 0.097665f
C456 output.n46 gnd 0.015803f
C457 output.n47 gnd 0.011243f
C458 output.n48 gnd 0.006041f
C459 output.n49 gnd 0.01428f
C460 output.n50 gnd 0.006397f
C461 output.n51 gnd 0.011243f
C462 output.n52 gnd 0.006041f
C463 output.n53 gnd 0.01428f
C464 output.n54 gnd 0.006397f
C465 output.n55 gnd 0.048111f
C466 output.t18 gnd 0.023274f
C467 output.n56 gnd 0.01071f
C468 output.n57 gnd 0.008435f
C469 output.n58 gnd 0.006041f
C470 output.n59 gnd 0.267512f
C471 output.n60 gnd 0.011243f
C472 output.n61 gnd 0.006041f
C473 output.n62 gnd 0.006397f
C474 output.n63 gnd 0.01428f
C475 output.n64 gnd 0.01428f
C476 output.n65 gnd 0.006397f
C477 output.n66 gnd 0.006041f
C478 output.n67 gnd 0.011243f
C479 output.n68 gnd 0.011243f
C480 output.n69 gnd 0.006041f
C481 output.n70 gnd 0.006397f
C482 output.n71 gnd 0.01428f
C483 output.n72 gnd 0.030913f
C484 output.n73 gnd 0.006397f
C485 output.n74 gnd 0.006041f
C486 output.n75 gnd 0.025987f
C487 output.n76 gnd 0.09306f
C488 output.n77 gnd 1.65264f
C489 output.n78 gnd 0.015803f
C490 output.n79 gnd 0.011243f
C491 output.n80 gnd 0.006041f
C492 output.n81 gnd 0.01428f
C493 output.n82 gnd 0.006397f
C494 output.n83 gnd 0.011243f
C495 output.n84 gnd 0.006041f
C496 output.n85 gnd 0.01428f
C497 output.n86 gnd 0.006397f
C498 output.n87 gnd 0.048111f
C499 output.t17 gnd 0.023274f
C500 output.n88 gnd 0.01071f
C501 output.n89 gnd 0.008435f
C502 output.n90 gnd 0.006041f
C503 output.n91 gnd 0.267512f
C504 output.n92 gnd 0.011243f
C505 output.n93 gnd 0.006041f
C506 output.n94 gnd 0.006397f
C507 output.n95 gnd 0.01428f
C508 output.n96 gnd 0.01428f
C509 output.n97 gnd 0.006397f
C510 output.n98 gnd 0.006041f
C511 output.n99 gnd 0.011243f
C512 output.n100 gnd 0.011243f
C513 output.n101 gnd 0.006041f
C514 output.n102 gnd 0.006397f
C515 output.n103 gnd 0.01428f
C516 output.n104 gnd 0.030913f
C517 output.n105 gnd 0.006397f
C518 output.n106 gnd 0.006041f
C519 output.n107 gnd 0.025987f
C520 output.n108 gnd 0.09306f
C521 output.n109 gnd 0.713089f
C522 output.n110 gnd 0.015803f
C523 output.n111 gnd 0.011243f
C524 output.n112 gnd 0.006041f
C525 output.n113 gnd 0.01428f
C526 output.n114 gnd 0.006397f
C527 output.n115 gnd 0.011243f
C528 output.n116 gnd 0.006041f
C529 output.n117 gnd 0.01428f
C530 output.n118 gnd 0.006397f
C531 output.n119 gnd 0.048111f
C532 output.t16 gnd 0.023274f
C533 output.n120 gnd 0.01071f
C534 output.n121 gnd 0.008435f
C535 output.n122 gnd 0.006041f
C536 output.n123 gnd 0.267512f
C537 output.n124 gnd 0.011243f
C538 output.n125 gnd 0.006041f
C539 output.n126 gnd 0.006397f
C540 output.n127 gnd 0.01428f
C541 output.n128 gnd 0.01428f
C542 output.n129 gnd 0.006397f
C543 output.n130 gnd 0.006041f
C544 output.n131 gnd 0.011243f
C545 output.n132 gnd 0.011243f
C546 output.n133 gnd 0.006041f
C547 output.n134 gnd 0.006397f
C548 output.n135 gnd 0.01428f
C549 output.n136 gnd 0.030913f
C550 output.n137 gnd 0.006397f
C551 output.n138 gnd 0.006041f
C552 output.n139 gnd 0.025987f
C553 output.n140 gnd 0.09306f
C554 output.n141 gnd 1.67353f
C555 outputibias.t9 gnd 0.11477f
C556 outputibias.t8 gnd 0.115567f
C557 outputibias.n0 gnd 0.130108f
C558 outputibias.n1 gnd 0.001372f
C559 outputibias.n2 gnd 9.76e-19
C560 outputibias.n3 gnd 5.24e-19
C561 outputibias.n4 gnd 0.001239f
C562 outputibias.n5 gnd 5.55e-19
C563 outputibias.n6 gnd 9.76e-19
C564 outputibias.n7 gnd 5.24e-19
C565 outputibias.n8 gnd 0.001239f
C566 outputibias.n9 gnd 5.55e-19
C567 outputibias.n10 gnd 0.004176f
C568 outputibias.t5 gnd 0.00202f
C569 outputibias.n11 gnd 9.3e-19
C570 outputibias.n12 gnd 7.32e-19
C571 outputibias.n13 gnd 5.24e-19
C572 outputibias.n14 gnd 0.02322f
C573 outputibias.n15 gnd 9.76e-19
C574 outputibias.n16 gnd 5.24e-19
C575 outputibias.n17 gnd 5.55e-19
C576 outputibias.n18 gnd 0.001239f
C577 outputibias.n19 gnd 0.001239f
C578 outputibias.n20 gnd 5.55e-19
C579 outputibias.n21 gnd 5.24e-19
C580 outputibias.n22 gnd 9.76e-19
C581 outputibias.n23 gnd 9.76e-19
C582 outputibias.n24 gnd 5.24e-19
C583 outputibias.n25 gnd 5.55e-19
C584 outputibias.n26 gnd 0.001239f
C585 outputibias.n27 gnd 0.002683f
C586 outputibias.n28 gnd 5.55e-19
C587 outputibias.n29 gnd 5.24e-19
C588 outputibias.n30 gnd 0.002256f
C589 outputibias.n31 gnd 0.005781f
C590 outputibias.n32 gnd 0.001372f
C591 outputibias.n33 gnd 9.76e-19
C592 outputibias.n34 gnd 5.24e-19
C593 outputibias.n35 gnd 0.001239f
C594 outputibias.n36 gnd 5.55e-19
C595 outputibias.n37 gnd 9.76e-19
C596 outputibias.n38 gnd 5.24e-19
C597 outputibias.n39 gnd 0.001239f
C598 outputibias.n40 gnd 5.55e-19
C599 outputibias.n41 gnd 0.004176f
C600 outputibias.t7 gnd 0.00202f
C601 outputibias.n42 gnd 9.3e-19
C602 outputibias.n43 gnd 7.32e-19
C603 outputibias.n44 gnd 5.24e-19
C604 outputibias.n45 gnd 0.02322f
C605 outputibias.n46 gnd 9.76e-19
C606 outputibias.n47 gnd 5.24e-19
C607 outputibias.n48 gnd 5.55e-19
C608 outputibias.n49 gnd 0.001239f
C609 outputibias.n50 gnd 0.001239f
C610 outputibias.n51 gnd 5.55e-19
C611 outputibias.n52 gnd 5.24e-19
C612 outputibias.n53 gnd 9.76e-19
C613 outputibias.n54 gnd 9.76e-19
C614 outputibias.n55 gnd 5.24e-19
C615 outputibias.n56 gnd 5.55e-19
C616 outputibias.n57 gnd 0.001239f
C617 outputibias.n58 gnd 0.002683f
C618 outputibias.n59 gnd 5.55e-19
C619 outputibias.n60 gnd 5.24e-19
C620 outputibias.n61 gnd 0.002256f
C621 outputibias.n62 gnd 0.005197f
C622 outputibias.n63 gnd 0.121892f
C623 outputibias.n64 gnd 0.001372f
C624 outputibias.n65 gnd 9.76e-19
C625 outputibias.n66 gnd 5.24e-19
C626 outputibias.n67 gnd 0.001239f
C627 outputibias.n68 gnd 5.55e-19
C628 outputibias.n69 gnd 9.76e-19
C629 outputibias.n70 gnd 5.24e-19
C630 outputibias.n71 gnd 0.001239f
C631 outputibias.n72 gnd 5.55e-19
C632 outputibias.n73 gnd 0.004176f
C633 outputibias.t1 gnd 0.00202f
C634 outputibias.n74 gnd 9.3e-19
C635 outputibias.n75 gnd 7.32e-19
C636 outputibias.n76 gnd 5.24e-19
C637 outputibias.n77 gnd 0.02322f
C638 outputibias.n78 gnd 9.76e-19
C639 outputibias.n79 gnd 5.24e-19
C640 outputibias.n80 gnd 5.55e-19
C641 outputibias.n81 gnd 0.001239f
C642 outputibias.n82 gnd 0.001239f
C643 outputibias.n83 gnd 5.55e-19
C644 outputibias.n84 gnd 5.24e-19
C645 outputibias.n85 gnd 9.76e-19
C646 outputibias.n86 gnd 9.76e-19
C647 outputibias.n87 gnd 5.24e-19
C648 outputibias.n88 gnd 5.55e-19
C649 outputibias.n89 gnd 0.001239f
C650 outputibias.n90 gnd 0.002683f
C651 outputibias.n91 gnd 5.55e-19
C652 outputibias.n92 gnd 5.24e-19
C653 outputibias.n93 gnd 0.002256f
C654 outputibias.n94 gnd 0.005197f
C655 outputibias.n95 gnd 0.064513f
C656 outputibias.n96 gnd 0.001372f
C657 outputibias.n97 gnd 9.76e-19
C658 outputibias.n98 gnd 5.24e-19
C659 outputibias.n99 gnd 0.001239f
C660 outputibias.n100 gnd 5.55e-19
C661 outputibias.n101 gnd 9.76e-19
C662 outputibias.n102 gnd 5.24e-19
C663 outputibias.n103 gnd 0.001239f
C664 outputibias.n104 gnd 5.55e-19
C665 outputibias.n105 gnd 0.004176f
C666 outputibias.t3 gnd 0.00202f
C667 outputibias.n106 gnd 9.3e-19
C668 outputibias.n107 gnd 7.32e-19
C669 outputibias.n108 gnd 5.24e-19
C670 outputibias.n109 gnd 0.02322f
C671 outputibias.n110 gnd 9.76e-19
C672 outputibias.n111 gnd 5.24e-19
C673 outputibias.n112 gnd 5.55e-19
C674 outputibias.n113 gnd 0.001239f
C675 outputibias.n114 gnd 0.001239f
C676 outputibias.n115 gnd 5.55e-19
C677 outputibias.n116 gnd 5.24e-19
C678 outputibias.n117 gnd 9.76e-19
C679 outputibias.n118 gnd 9.76e-19
C680 outputibias.n119 gnd 5.24e-19
C681 outputibias.n120 gnd 5.55e-19
C682 outputibias.n121 gnd 0.001239f
C683 outputibias.n122 gnd 0.002683f
C684 outputibias.n123 gnd 5.55e-19
C685 outputibias.n124 gnd 5.24e-19
C686 outputibias.n125 gnd 0.002256f
C687 outputibias.n126 gnd 0.005197f
C688 outputibias.n127 gnd 0.084814f
C689 outputibias.t2 gnd 0.108319f
C690 outputibias.t0 gnd 0.108319f
C691 outputibias.t6 gnd 0.108319f
C692 outputibias.t4 gnd 0.109238f
C693 outputibias.n128 gnd 0.134674f
C694 outputibias.n129 gnd 0.07244f
C695 outputibias.n130 gnd 0.079818f
C696 outputibias.n131 gnd 0.164901f
C697 outputibias.t11 gnd 0.11477f
C698 outputibias.n132 gnd 0.067481f
C699 outputibias.t10 gnd 0.11477f
C700 outputibias.n133 gnd 0.065115f
C701 outputibias.n134 gnd 0.029159f
C702 a_n1808_13878.t11 gnd 0.185195f
C703 a_n1808_13878.t13 gnd 0.185195f
C704 a_n1808_13878.t17 gnd 0.185195f
C705 a_n1808_13878.n0 gnd 1.46067f
C706 a_n1808_13878.t8 gnd 0.185195f
C707 a_n1808_13878.t10 gnd 0.185195f
C708 a_n1808_13878.n1 gnd 1.4598f
C709 a_n1808_13878.t14 gnd 0.185195f
C710 a_n1808_13878.t9 gnd 0.185195f
C711 a_n1808_13878.n2 gnd 1.45825f
C712 a_n1808_13878.n3 gnd 2.03762f
C713 a_n1808_13878.t12 gnd 0.185195f
C714 a_n1808_13878.t19 gnd 0.185195f
C715 a_n1808_13878.n4 gnd 1.45825f
C716 a_n1808_13878.n5 gnd 3.69301f
C717 a_n1808_13878.t1 gnd 1.73408f
C718 a_n1808_13878.t4 gnd 0.185195f
C719 a_n1808_13878.t5 gnd 0.185195f
C720 a_n1808_13878.n6 gnd 1.30452f
C721 a_n1808_13878.n7 gnd 1.4576f
C722 a_n1808_13878.t0 gnd 1.73062f
C723 a_n1808_13878.n8 gnd 0.733487f
C724 a_n1808_13878.t3 gnd 1.73062f
C725 a_n1808_13878.n9 gnd 0.733487f
C726 a_n1808_13878.t6 gnd 0.185195f
C727 a_n1808_13878.t7 gnd 0.185195f
C728 a_n1808_13878.n10 gnd 1.30452f
C729 a_n1808_13878.n11 gnd 0.74059f
C730 a_n1808_13878.t2 gnd 1.73062f
C731 a_n1808_13878.n12 gnd 1.7272f
C732 a_n1808_13878.n13 gnd 2.51438f
C733 a_n1808_13878.t15 gnd 0.185195f
C734 a_n1808_13878.t16 gnd 0.185195f
C735 a_n1808_13878.n14 gnd 1.45825f
C736 a_n1808_13878.n15 gnd 1.80025f
C737 a_n1808_13878.n16 gnd 1.31079f
C738 a_n1808_13878.n17 gnd 1.45826f
C739 a_n1808_13878.t18 gnd 0.185195f
C740 a_n1986_8322.t0 gnd 38.672398f
C741 a_n1986_8322.t2 gnd 27.512402f
C742 a_n1986_8322.t3 gnd 19.268198f
C743 a_n1986_8322.t1 gnd 38.672398f
C744 a_n1986_8322.t6 gnd 0.093533f
C745 a_n1986_8322.t5 gnd 0.875792f
C746 a_n1986_8322.t13 gnd 0.093533f
C747 a_n1986_8322.t8 gnd 0.093533f
C748 a_n1986_8322.n0 gnd 0.658844f
C749 a_n1986_8322.n1 gnd 0.736161f
C750 a_n1986_8322.t11 gnd 0.093533f
C751 a_n1986_8322.t10 gnd 0.093533f
C752 a_n1986_8322.n2 gnd 0.658844f
C753 a_n1986_8322.n3 gnd 0.374034f
C754 a_n1986_8322.t4 gnd 0.874048f
C755 a_n1986_8322.n4 gnd 1.39896f
C756 a_n1986_8322.t18 gnd 0.875792f
C757 a_n1986_8322.t22 gnd 0.093533f
C758 a_n1986_8322.t21 gnd 0.093533f
C759 a_n1986_8322.n5 gnd 0.658844f
C760 a_n1986_8322.n6 gnd 0.736161f
C761 a_n1986_8322.t16 gnd 0.874048f
C762 a_n1986_8322.n7 gnd 0.370446f
C763 a_n1986_8322.t19 gnd 0.874048f
C764 a_n1986_8322.n8 gnd 0.370446f
C765 a_n1986_8322.t17 gnd 0.093533f
C766 a_n1986_8322.t23 gnd 0.093533f
C767 a_n1986_8322.n9 gnd 0.658844f
C768 a_n1986_8322.n10 gnd 0.374034f
C769 a_n1986_8322.t20 gnd 0.874048f
C770 a_n1986_8322.n11 gnd 0.872317f
C771 a_n1986_8322.n12 gnd 1.59071f
C772 a_n1986_8322.n13 gnd 3.20172f
C773 a_n1986_8322.t7 gnd 0.874048f
C774 a_n1986_8322.n14 gnd 0.76652f
C775 a_n1986_8322.t14 gnd 0.875789f
C776 a_n1986_8322.t12 gnd 0.093533f
C777 a_n1986_8322.t9 gnd 0.093533f
C778 a_n1986_8322.n15 gnd 0.658844f
C779 a_n1986_8322.n16 gnd 0.736163f
C780 a_n1986_8322.n17 gnd 0.374032f
C781 a_n1986_8322.n18 gnd 0.658845f
C782 a_n1986_8322.t15 gnd 0.093533f
C783 a_n1986_13878.n0 gnd 0.543543f
C784 a_n1986_13878.n1 gnd 0.211712f
C785 a_n1986_13878.n2 gnd 0.15593f
C786 a_n1986_13878.n3 gnd 0.245072f
C787 a_n1986_13878.n4 gnd 0.18929f
C788 a_n1986_13878.n5 gnd 0.211712f
C789 a_n1986_13878.n6 gnd 1.03979f
C790 a_n1986_13878.n7 gnd 0.15593f
C791 a_n1986_13878.n8 gnd 0.599325f
C792 a_n1986_13878.n9 gnd 0.446674f
C793 a_n1986_13878.n10 gnd 0.223128f
C794 a_n1986_13878.n11 gnd 0.508859f
C795 a_n1986_13878.n12 gnd 0.291913f
C796 a_n1986_13878.n13 gnd 0.453077f
C797 a_n1986_13878.n14 gnd 0.223128f
C798 a_n1986_13878.n15 gnd 0.755878f
C799 a_n1986_13878.n16 gnd 0.291913f
C800 a_n1986_13878.n17 gnd 0.508859f
C801 a_n1986_13878.n18 gnd 0.686545f
C802 a_n1986_13878.n19 gnd 0.223128f
C803 a_n1986_13878.n20 gnd 0.291913f
C804 a_n1986_13878.n21 gnd 0.66047f
C805 a_n1986_13878.n22 gnd 0.291913f
C806 a_n1986_13878.n23 gnd 3.60937f
C807 a_n1986_13878.n24 gnd 2.74915f
C808 a_n1986_13878.n25 gnd 3.87242f
C809 a_n1986_13878.n26 gnd 1.21809f
C810 a_n1986_13878.n27 gnd 1.97943f
C811 a_n1986_13878.n28 gnd 1.83699f
C812 a_n1986_13878.n29 gnd 0.751202f
C813 a_n1986_13878.n30 gnd 0.751204f
C814 a_n1986_13878.n31 gnd 3.32125f
C815 a_n1986_13878.n32 gnd 0.111564f
C816 a_n1986_13878.n33 gnd 0.008639f
C817 a_n1986_13878.n35 gnd 0.008639f
C818 a_n1986_13878.n37 gnd 0.295172f
C819 a_n1986_13878.n38 gnd 0.008639f
C820 a_n1986_13878.n40 gnd 0.295172f
C821 a_n1986_13878.n41 gnd 0.008639f
C822 a_n1986_13878.n43 gnd 0.295172f
C823 a_n1986_13878.n44 gnd 0.008639f
C824 a_n1986_13878.n45 gnd 0.294752f
C825 a_n1986_13878.n46 gnd 0.008639f
C826 a_n1986_13878.n47 gnd 0.294752f
C827 a_n1986_13878.n48 gnd 0.008639f
C828 a_n1986_13878.n49 gnd 0.294752f
C829 a_n1986_13878.n50 gnd 0.008639f
C830 a_n1986_13878.n51 gnd 0.294752f
C831 a_n1986_13878.n52 gnd 0.295172f
C832 a_n1986_13878.t0 gnd 0.73505f
C833 a_n1986_13878.t2 gnd 0.719888f
C834 a_n1986_13878.t6 gnd 0.719888f
C835 a_n1986_13878.t20 gnd 0.719888f
C836 a_n1986_13878.n53 gnd 0.316508f
C837 a_n1986_13878.t16 gnd 0.731791f
C838 a_n1986_13878.t45 gnd 0.120372f
C839 a_n1986_13878.t29 gnd 0.120372f
C840 a_n1986_13878.n54 gnd 1.06535f
C841 a_n1986_13878.t38 gnd 0.120372f
C842 a_n1986_13878.t46 gnd 0.120372f
C843 a_n1986_13878.n55 gnd 1.06365f
C844 a_n1986_13878.t26 gnd 0.120372f
C845 a_n1986_13878.t35 gnd 0.120372f
C846 a_n1986_13878.n56 gnd 1.06365f
C847 a_n1986_13878.t33 gnd 0.120372f
C848 a_n1986_13878.t37 gnd 0.120372f
C849 a_n1986_13878.n57 gnd 1.06535f
C850 a_n1986_13878.t42 gnd 0.120372f
C851 a_n1986_13878.t28 gnd 0.120372f
C852 a_n1986_13878.n58 gnd 1.06365f
C853 a_n1986_13878.t34 gnd 0.120372f
C854 a_n1986_13878.t44 gnd 0.120372f
C855 a_n1986_13878.n59 gnd 1.06365f
C856 a_n1986_13878.t30 gnd 0.120372f
C857 a_n1986_13878.t31 gnd 0.120372f
C858 a_n1986_13878.n60 gnd 1.06365f
C859 a_n1986_13878.t41 gnd 0.120372f
C860 a_n1986_13878.t40 gnd 0.120372f
C861 a_n1986_13878.n61 gnd 1.06365f
C862 a_n1986_13878.t27 gnd 0.120372f
C863 a_n1986_13878.t43 gnd 0.120372f
C864 a_n1986_13878.n62 gnd 1.06365f
C865 a_n1986_13878.t39 gnd 0.120372f
C866 a_n1986_13878.t24 gnd 0.120372f
C867 a_n1986_13878.n63 gnd 1.06535f
C868 a_n1986_13878.t36 gnd 0.120372f
C869 a_n1986_13878.t25 gnd 0.120372f
C870 a_n1986_13878.n64 gnd 1.06365f
C871 a_n1986_13878.t47 gnd 0.120372f
C872 a_n1986_13878.t32 gnd 0.120372f
C873 a_n1986_13878.n65 gnd 1.06365f
C874 a_n1986_13878.t75 gnd 0.73505f
C875 a_n1986_13878.t58 gnd 0.719888f
C876 a_n1986_13878.t62 gnd 0.719888f
C877 a_n1986_13878.t52 gnd 0.719888f
C878 a_n1986_13878.n66 gnd 0.316508f
C879 a_n1986_13878.t67 gnd 0.719888f
C880 a_n1986_13878.t73 gnd 0.731791f
C881 a_n1986_13878.t19 gnd 1.44913f
C882 a_n1986_13878.t9 gnd 0.154764f
C883 a_n1986_13878.t5 gnd 0.154764f
C884 a_n1986_13878.n67 gnd 1.09016f
C885 a_n1986_13878.t11 gnd 0.154764f
C886 a_n1986_13878.t15 gnd 0.154764f
C887 a_n1986_13878.n68 gnd 1.09016f
C888 a_n1986_13878.t23 gnd 1.44624f
C889 a_n1986_13878.t10 gnd 0.719888f
C890 a_n1986_13878.n69 gnd 0.316508f
C891 a_n1986_13878.t14 gnd 0.719888f
C892 a_n1986_13878.t8 gnd 0.719888f
C893 a_n1986_13878.t56 gnd 0.719888f
C894 a_n1986_13878.n70 gnd 0.316508f
C895 a_n1986_13878.t65 gnd 0.719888f
C896 a_n1986_13878.t71 gnd 0.719888f
C897 a_n1986_13878.t70 gnd 0.73505f
C898 a_n1986_13878.n71 gnd 0.319212f
C899 a_n1986_13878.t50 gnd 0.719888f
C900 a_n1986_13878.n72 gnd 0.312489f
C901 a_n1986_13878.n73 gnd 0.319213f
C902 a_n1986_13878.t51 gnd 0.731791f
C903 a_n1986_13878.t18 gnd 0.73505f
C904 a_n1986_13878.n74 gnd 0.319212f
C905 a_n1986_13878.t4 gnd 0.719888f
C906 a_n1986_13878.n75 gnd 0.312489f
C907 a_n1986_13878.n76 gnd 0.319213f
C908 a_n1986_13878.t22 gnd 0.731791f
C909 a_n1986_13878.n77 gnd 1.16971f
C910 a_n1986_13878.t55 gnd 0.719888f
C911 a_n1986_13878.n78 gnd 0.312489f
C912 a_n1986_13878.t61 gnd 0.719888f
C913 a_n1986_13878.n79 gnd 0.312489f
C914 a_n1986_13878.t53 gnd 0.719888f
C915 a_n1986_13878.n80 gnd 0.312489f
C916 a_n1986_13878.t66 gnd 0.719888f
C917 a_n1986_13878.n81 gnd 0.312489f
C918 a_n1986_13878.t57 gnd 0.719888f
C919 a_n1986_13878.n82 gnd 0.306814f
C920 a_n1986_13878.t48 gnd 0.719888f
C921 a_n1986_13878.n83 gnd 0.316508f
C922 a_n1986_13878.t59 gnd 0.731951f
C923 a_n1986_13878.t68 gnd 0.719888f
C924 a_n1986_13878.n84 gnd 0.306814f
C925 a_n1986_13878.t54 gnd 0.719888f
C926 a_n1986_13878.n85 gnd 0.316508f
C927 a_n1986_13878.t63 gnd 0.731951f
C928 a_n1986_13878.t72 gnd 0.719888f
C929 a_n1986_13878.n86 gnd 0.306814f
C930 a_n1986_13878.t60 gnd 0.719888f
C931 a_n1986_13878.n87 gnd 0.316508f
C932 a_n1986_13878.t74 gnd 0.731951f
C933 a_n1986_13878.t64 gnd 0.719888f
C934 a_n1986_13878.n88 gnd 0.306814f
C935 a_n1986_13878.t49 gnd 0.719888f
C936 a_n1986_13878.n89 gnd 0.316508f
C937 a_n1986_13878.t69 gnd 0.731951f
C938 a_n1986_13878.n90 gnd 1.38299f
C939 a_n1986_13878.n91 gnd 0.319213f
C940 a_n1986_13878.n92 gnd 0.312489f
C941 a_n1986_13878.n93 gnd 0.319212f
C942 a_n1986_13878.t12 gnd 0.719888f
C943 a_n1986_13878.n94 gnd 0.319213f
C944 a_n1986_13878.n95 gnd 0.312489f
C945 a_n1986_13878.n96 gnd 0.319212f
C946 a_n1986_13878.n97 gnd 0.813122f
C947 a_n1986_13878.t17 gnd 1.44913f
C948 a_n1986_13878.t21 gnd 0.154764f
C949 a_n1986_13878.t13 gnd 0.154764f
C950 a_n1986_13878.n98 gnd 1.09016f
C951 a_n1986_13878.t3 gnd 0.154764f
C952 a_n1986_13878.t7 gnd 0.154764f
C953 a_n1986_13878.n99 gnd 1.09016f
C954 a_n1986_13878.n100 gnd 1.18267f
C955 a_n1986_13878.t1 gnd 1.44625f
C956 a_n6308_8799.n0 gnd 0.181284f
C957 a_n6308_8799.n1 gnd 0.212295f
C958 a_n6308_8799.n2 gnd 0.212295f
C959 a_n6308_8799.n3 gnd 0.212295f
C960 a_n6308_8799.n4 gnd 0.181284f
C961 a_n6308_8799.n5 gnd 0.212295f
C962 a_n6308_8799.n6 gnd 0.212295f
C963 a_n6308_8799.n7 gnd 0.212295f
C964 a_n6308_8799.n8 gnd 0.350177f
C965 a_n6308_8799.n9 gnd 0.212295f
C966 a_n6308_8799.n10 gnd 0.212295f
C967 a_n6308_8799.n11 gnd 0.212295f
C968 a_n6308_8799.n12 gnd 0.212295f
C969 a_n6308_8799.n13 gnd 0.212295f
C970 a_n6308_8799.n14 gnd 0.181284f
C971 a_n6308_8799.n15 gnd 0.212295f
C972 a_n6308_8799.n16 gnd 0.212295f
C973 a_n6308_8799.n17 gnd 0.212295f
C974 a_n6308_8799.n18 gnd 0.181284f
C975 a_n6308_8799.n19 gnd 0.212295f
C976 a_n6308_8799.n20 gnd 0.212295f
C977 a_n6308_8799.n21 gnd 0.212295f
C978 a_n6308_8799.n22 gnd 0.350177f
C979 a_n6308_8799.n23 gnd 0.212295f
C980 a_n6308_8799.n24 gnd 3.48405f
C981 a_n6308_8799.n25 gnd 1.77648f
C982 a_n6308_8799.n26 gnd 3.02258f
C983 a_n6308_8799.n27 gnd 4.05465f
C984 a_n6308_8799.n28 gnd 2.89712f
C985 a_n6308_8799.n29 gnd 0.714731f
C986 a_n6308_8799.n30 gnd 0.256734f
C987 a_n6308_8799.n32 gnd 0.007907f
C988 a_n6308_8799.n33 gnd 0.011952f
C989 a_n6308_8799.n34 gnd 0.008219f
C990 a_n6308_8799.n36 gnd 4.11e-19
C991 a_n6308_8799.n37 gnd 0.008518f
C992 a_n6308_8799.n38 gnd 0.268575f
C993 a_n6308_8799.n39 gnd 0.256734f
C994 a_n6308_8799.n41 gnd 0.007907f
C995 a_n6308_8799.n42 gnd 0.011952f
C996 a_n6308_8799.n43 gnd 0.008219f
C997 a_n6308_8799.n45 gnd 4.11e-19
C998 a_n6308_8799.n46 gnd 0.008518f
C999 a_n6308_8799.n47 gnd 0.268575f
C1000 a_n6308_8799.n48 gnd 0.256734f
C1001 a_n6308_8799.n50 gnd 0.007907f
C1002 a_n6308_8799.n51 gnd 0.011952f
C1003 a_n6308_8799.n52 gnd 0.008219f
C1004 a_n6308_8799.n54 gnd 4.11e-19
C1005 a_n6308_8799.n55 gnd 0.008518f
C1006 a_n6308_8799.n56 gnd 0.268575f
C1007 a_n6308_8799.n57 gnd 0.008518f
C1008 a_n6308_8799.n58 gnd 0.268575f
C1009 a_n6308_8799.n59 gnd 4.11e-19
C1010 a_n6308_8799.n61 gnd 0.008219f
C1011 a_n6308_8799.n62 gnd 0.011952f
C1012 a_n6308_8799.n63 gnd 0.007907f
C1013 a_n6308_8799.n65 gnd 0.256734f
C1014 a_n6308_8799.n66 gnd 0.008518f
C1015 a_n6308_8799.n67 gnd 0.268575f
C1016 a_n6308_8799.n68 gnd 4.11e-19
C1017 a_n6308_8799.n70 gnd 0.008219f
C1018 a_n6308_8799.n71 gnd 0.011952f
C1019 a_n6308_8799.n72 gnd 0.007907f
C1020 a_n6308_8799.n74 gnd 0.256734f
C1021 a_n6308_8799.n75 gnd 0.008518f
C1022 a_n6308_8799.n76 gnd 0.268575f
C1023 a_n6308_8799.n77 gnd 4.11e-19
C1024 a_n6308_8799.n79 gnd 0.008219f
C1025 a_n6308_8799.n80 gnd 0.011952f
C1026 a_n6308_8799.n81 gnd 0.007907f
C1027 a_n6308_8799.n83 gnd 0.256734f
C1028 a_n6308_8799.t16 gnd 0.14725f
C1029 a_n6308_8799.t9 gnd 0.14725f
C1030 a_n6308_8799.t21 gnd 0.14725f
C1031 a_n6308_8799.n84 gnd 1.16138f
C1032 a_n6308_8799.t20 gnd 0.14725f
C1033 a_n6308_8799.t28 gnd 0.14725f
C1034 a_n6308_8799.n85 gnd 1.15947f
C1035 a_n6308_8799.t13 gnd 0.14725f
C1036 a_n6308_8799.t14 gnd 0.14725f
C1037 a_n6308_8799.n86 gnd 1.15947f
C1038 a_n6308_8799.t6 gnd 0.114528f
C1039 a_n6308_8799.t29 gnd 0.114528f
C1040 a_n6308_8799.n87 gnd 1.01362f
C1041 a_n6308_8799.t30 gnd 0.114528f
C1042 a_n6308_8799.t11 gnd 0.114528f
C1043 a_n6308_8799.n88 gnd 1.01201f
C1044 a_n6308_8799.t4 gnd 0.114528f
C1045 a_n6308_8799.t12 gnd 0.114528f
C1046 a_n6308_8799.n89 gnd 1.01201f
C1047 a_n6308_8799.t19 gnd 0.114528f
C1048 a_n6308_8799.t0 gnd 0.114528f
C1049 a_n6308_8799.n90 gnd 1.01362f
C1050 a_n6308_8799.t10 gnd 0.114528f
C1051 a_n6308_8799.t35 gnd 0.114528f
C1052 a_n6308_8799.n91 gnd 1.01201f
C1053 a_n6308_8799.t5 gnd 0.114528f
C1054 a_n6308_8799.t17 gnd 0.114528f
C1055 a_n6308_8799.n92 gnd 1.01201f
C1056 a_n6308_8799.t32 gnd 0.114528f
C1057 a_n6308_8799.t2 gnd 0.114528f
C1058 a_n6308_8799.n93 gnd 1.01362f
C1059 a_n6308_8799.t34 gnd 0.114528f
C1060 a_n6308_8799.t26 gnd 0.114528f
C1061 a_n6308_8799.n94 gnd 1.01201f
C1062 a_n6308_8799.t3 gnd 0.114528f
C1063 a_n6308_8799.t31 gnd 0.114528f
C1064 a_n6308_8799.n95 gnd 1.01201f
C1065 a_n6308_8799.t27 gnd 0.114528f
C1066 a_n6308_8799.t1 gnd 0.114528f
C1067 a_n6308_8799.n96 gnd 1.01201f
C1068 a_n6308_8799.t23 gnd 0.114528f
C1069 a_n6308_8799.t33 gnd 0.114528f
C1070 a_n6308_8799.n97 gnd 1.01201f
C1071 a_n6308_8799.t24 gnd 0.114528f
C1072 a_n6308_8799.t18 gnd 0.114528f
C1073 a_n6308_8799.n98 gnd 1.01201f
C1074 a_n6308_8799.t95 gnd 0.610567f
C1075 a_n6308_8799.n99 gnd 0.276336f
C1076 a_n6308_8799.t43 gnd 0.610567f
C1077 a_n6308_8799.t44 gnd 0.610567f
C1078 a_n6308_8799.n100 gnd 0.267292f
C1079 a_n6308_8799.t57 gnd 0.610567f
C1080 a_n6308_8799.n101 gnd 0.278925f
C1081 a_n6308_8799.t72 gnd 0.610567f
C1082 a_n6308_8799.t85 gnd 0.610567f
C1083 a_n6308_8799.n102 gnd 0.2722f
C1084 a_n6308_8799.t60 gnd 0.624917f
C1085 a_n6308_8799.t61 gnd 0.610567f
C1086 a_n6308_8799.n103 gnd 0.27848f
C1087 a_n6308_8799.n104 gnd 0.254517f
C1088 a_n6308_8799.t37 gnd 0.610567f
C1089 a_n6308_8799.n105 gnd 0.276216f
C1090 a_n6308_8799.n106 gnd 0.276351f
C1091 a_n6308_8799.t97 gnd 0.610567f
C1092 a_n6308_8799.n107 gnd 0.272527f
C1093 a_n6308_8799.t56 gnd 0.610567f
C1094 a_n6308_8799.n108 gnd 0.272783f
C1095 a_n6308_8799.n109 gnd 0.27848f
C1096 a_n6308_8799.t42 gnd 0.621652f
C1097 a_n6308_8799.t101 gnd 0.610567f
C1098 a_n6308_8799.n110 gnd 0.276336f
C1099 a_n6308_8799.t49 gnd 0.610567f
C1100 a_n6308_8799.t53 gnd 0.610567f
C1101 a_n6308_8799.n111 gnd 0.267292f
C1102 a_n6308_8799.t65 gnd 0.610567f
C1103 a_n6308_8799.n112 gnd 0.278925f
C1104 a_n6308_8799.t79 gnd 0.610567f
C1105 a_n6308_8799.t92 gnd 0.610567f
C1106 a_n6308_8799.n113 gnd 0.2722f
C1107 a_n6308_8799.t66 gnd 0.624917f
C1108 a_n6308_8799.t67 gnd 0.610567f
C1109 a_n6308_8799.n114 gnd 0.27848f
C1110 a_n6308_8799.n115 gnd 0.254517f
C1111 a_n6308_8799.t45 gnd 0.610567f
C1112 a_n6308_8799.n116 gnd 0.276216f
C1113 a_n6308_8799.n117 gnd 0.276351f
C1114 a_n6308_8799.t105 gnd 0.610567f
C1115 a_n6308_8799.n118 gnd 0.272527f
C1116 a_n6308_8799.t64 gnd 0.610567f
C1117 a_n6308_8799.n119 gnd 0.272783f
C1118 a_n6308_8799.n120 gnd 0.27848f
C1119 a_n6308_8799.t51 gnd 0.621652f
C1120 a_n6308_8799.n121 gnd 0.916628f
C1121 a_n6308_8799.t76 gnd 0.610567f
C1122 a_n6308_8799.n122 gnd 0.276336f
C1123 a_n6308_8799.t47 gnd 0.610567f
C1124 a_n6308_8799.t94 gnd 0.610567f
C1125 a_n6308_8799.n123 gnd 0.267292f
C1126 a_n6308_8799.t41 gnd 0.610567f
C1127 a_n6308_8799.n124 gnd 0.278925f
C1128 a_n6308_8799.t82 gnd 0.610567f
C1129 a_n6308_8799.t103 gnd 0.610567f
C1130 a_n6308_8799.n125 gnd 0.2722f
C1131 a_n6308_8799.t99 gnd 0.624917f
C1132 a_n6308_8799.t87 gnd 0.610567f
C1133 a_n6308_8799.n126 gnd 0.27848f
C1134 a_n6308_8799.n127 gnd 0.254517f
C1135 a_n6308_8799.t71 gnd 0.610567f
C1136 a_n6308_8799.n128 gnd 0.276216f
C1137 a_n6308_8799.n129 gnd 0.276351f
C1138 a_n6308_8799.t52 gnd 0.610567f
C1139 a_n6308_8799.n130 gnd 0.272527f
C1140 a_n6308_8799.t59 gnd 0.610567f
C1141 a_n6308_8799.n131 gnd 0.272783f
C1142 a_n6308_8799.n132 gnd 0.27848f
C1143 a_n6308_8799.t107 gnd 0.621652f
C1144 a_n6308_8799.n133 gnd 1.4839f
C1145 a_n6308_8799.t69 gnd 0.621652f
C1146 a_n6308_8799.t68 gnd 0.610567f
C1147 a_n6308_8799.t50 gnd 0.610567f
C1148 a_n6308_8799.t96 gnd 0.610567f
C1149 a_n6308_8799.n134 gnd 0.272783f
C1150 a_n6308_8799.t70 gnd 0.610567f
C1151 a_n6308_8799.t55 gnd 0.610567f
C1152 a_n6308_8799.t98 gnd 0.610567f
C1153 a_n6308_8799.n135 gnd 0.276351f
C1154 a_n6308_8799.t80 gnd 0.610567f
C1155 a_n6308_8799.t78 gnd 0.610567f
C1156 a_n6308_8799.t39 gnd 0.610567f
C1157 a_n6308_8799.n136 gnd 0.2722f
C1158 a_n6308_8799.t83 gnd 0.624917f
C1159 a_n6308_8799.t84 gnd 0.610567f
C1160 a_n6308_8799.n137 gnd 0.27848f
C1161 a_n6308_8799.n138 gnd 0.254517f
C1162 a_n6308_8799.n139 gnd 0.276216f
C1163 a_n6308_8799.n140 gnd 0.278925f
C1164 a_n6308_8799.n141 gnd 0.272527f
C1165 a_n6308_8799.n142 gnd 0.267292f
C1166 a_n6308_8799.n143 gnd 0.276336f
C1167 a_n6308_8799.n144 gnd 0.27848f
C1168 a_n6308_8799.t74 gnd 0.621652f
C1169 a_n6308_8799.t73 gnd 0.610567f
C1170 a_n6308_8799.t62 gnd 0.610567f
C1171 a_n6308_8799.t104 gnd 0.610567f
C1172 a_n6308_8799.n145 gnd 0.272783f
C1173 a_n6308_8799.t77 gnd 0.610567f
C1174 a_n6308_8799.t63 gnd 0.610567f
C1175 a_n6308_8799.t36 gnd 0.610567f
C1176 a_n6308_8799.n146 gnd 0.276351f
C1177 a_n6308_8799.t89 gnd 0.610567f
C1178 a_n6308_8799.t88 gnd 0.610567f
C1179 a_n6308_8799.t46 gnd 0.610567f
C1180 a_n6308_8799.n147 gnd 0.2722f
C1181 a_n6308_8799.t90 gnd 0.624917f
C1182 a_n6308_8799.t91 gnd 0.610567f
C1183 a_n6308_8799.n148 gnd 0.27848f
C1184 a_n6308_8799.n149 gnd 0.254517f
C1185 a_n6308_8799.n150 gnd 0.276216f
C1186 a_n6308_8799.n151 gnd 0.278925f
C1187 a_n6308_8799.n152 gnd 0.272527f
C1188 a_n6308_8799.n153 gnd 0.267292f
C1189 a_n6308_8799.n154 gnd 0.276336f
C1190 a_n6308_8799.n155 gnd 0.27848f
C1191 a_n6308_8799.n156 gnd 0.916628f
C1192 a_n6308_8799.t106 gnd 0.621652f
C1193 a_n6308_8799.t48 gnd 0.610567f
C1194 a_n6308_8799.t75 gnd 0.610567f
C1195 a_n6308_8799.t38 gnd 0.610567f
C1196 a_n6308_8799.n157 gnd 0.272783f
C1197 a_n6308_8799.t93 gnd 0.610567f
C1198 a_n6308_8799.t54 gnd 0.610567f
C1199 a_n6308_8799.t81 gnd 0.610567f
C1200 a_n6308_8799.n158 gnd 0.276351f
C1201 a_n6308_8799.t40 gnd 0.610567f
C1202 a_n6308_8799.t58 gnd 0.610567f
C1203 a_n6308_8799.t102 gnd 0.610567f
C1204 a_n6308_8799.n159 gnd 0.2722f
C1205 a_n6308_8799.t100 gnd 0.624917f
C1206 a_n6308_8799.t86 gnd 0.610567f
C1207 a_n6308_8799.n160 gnd 0.27848f
C1208 a_n6308_8799.n161 gnd 0.254517f
C1209 a_n6308_8799.n162 gnd 0.276216f
C1210 a_n6308_8799.n163 gnd 0.278925f
C1211 a_n6308_8799.n164 gnd 0.272527f
C1212 a_n6308_8799.n165 gnd 0.267292f
C1213 a_n6308_8799.n166 gnd 0.276336f
C1214 a_n6308_8799.n167 gnd 0.27848f
C1215 a_n6308_8799.n168 gnd 1.16031f
C1216 a_n6308_8799.n169 gnd 12.5067f
C1217 a_n6308_8799.n170 gnd 4.46846f
C1218 a_n6308_8799.n171 gnd 5.81379f
C1219 a_n6308_8799.t25 gnd 0.14725f
C1220 a_n6308_8799.t8 gnd 0.14725f
C1221 a_n6308_8799.n172 gnd 1.15947f
C1222 a_n6308_8799.t15 gnd 0.14725f
C1223 a_n6308_8799.t22 gnd 0.14725f
C1224 a_n6308_8799.n173 gnd 1.15947f
C1225 a_n6308_8799.n174 gnd 1.16139f
C1226 a_n6308_8799.t7 gnd 0.14725f
C1227 vdd.t221 gnd 0.035753f
C1228 vdd.t208 gnd 0.035753f
C1229 vdd.n0 gnd 0.281991f
C1230 vdd.t13 gnd 0.035753f
C1231 vdd.t179 gnd 0.035753f
C1232 vdd.n1 gnd 0.281525f
C1233 vdd.n2 gnd 0.25962f
C1234 vdd.t204 gnd 0.035753f
C1235 vdd.t183 gnd 0.035753f
C1236 vdd.n3 gnd 0.281525f
C1237 vdd.n4 gnd 0.1313f
C1238 vdd.t18 gnd 0.035753f
C1239 vdd.t177 gnd 0.035753f
C1240 vdd.n5 gnd 0.281525f
C1241 vdd.n6 gnd 0.1232f
C1242 vdd.t15 gnd 0.035753f
C1243 vdd.t206 gnd 0.035753f
C1244 vdd.n7 gnd 0.281991f
C1245 vdd.t81 gnd 0.035753f
C1246 vdd.t20 gnd 0.035753f
C1247 vdd.n8 gnd 0.281525f
C1248 vdd.n9 gnd 0.25962f
C1249 vdd.t210 gnd 0.035753f
C1250 vdd.t75 gnd 0.035753f
C1251 vdd.n10 gnd 0.281525f
C1252 vdd.n11 gnd 0.1313f
C1253 vdd.t78 gnd 0.035753f
C1254 vdd.t212 gnd 0.035753f
C1255 vdd.n12 gnd 0.281525f
C1256 vdd.n13 gnd 0.1232f
C1257 vdd.n14 gnd 0.0871f
C1258 vdd.t41 gnd 0.019863f
C1259 vdd.t45 gnd 0.019863f
C1260 vdd.n15 gnd 0.182829f
C1261 vdd.t51 gnd 0.019863f
C1262 vdd.t53 gnd 0.019863f
C1263 vdd.n16 gnd 0.182294f
C1264 vdd.n17 gnd 0.317249f
C1265 vdd.t49 gnd 0.019863f
C1266 vdd.t50 gnd 0.019863f
C1267 vdd.n18 gnd 0.182294f
C1268 vdd.n19 gnd 0.13125f
C1269 vdd.t52 gnd 0.019863f
C1270 vdd.t39 gnd 0.019863f
C1271 vdd.n20 gnd 0.182829f
C1272 vdd.t54 gnd 0.019863f
C1273 vdd.t44 gnd 0.019863f
C1274 vdd.n21 gnd 0.182294f
C1275 vdd.n22 gnd 0.317249f
C1276 vdd.t40 gnd 0.019863f
C1277 vdd.t42 gnd 0.019863f
C1278 vdd.n23 gnd 0.182294f
C1279 vdd.n24 gnd 0.13125f
C1280 vdd.t46 gnd 0.019863f
C1281 vdd.t43 gnd 0.019863f
C1282 vdd.n25 gnd 0.182294f
C1283 vdd.t48 gnd 0.019863f
C1284 vdd.t47 gnd 0.019863f
C1285 vdd.n26 gnd 0.182294f
C1286 vdd.n27 gnd 20.783f
C1287 vdd.n28 gnd 7.52955f
C1288 vdd.n29 gnd 0.005417f
C1289 vdd.n30 gnd 0.005027f
C1290 vdd.n31 gnd 0.002781f
C1291 vdd.n32 gnd 0.006385f
C1292 vdd.n33 gnd 0.002701f
C1293 vdd.n34 gnd 0.00286f
C1294 vdd.n35 gnd 0.005027f
C1295 vdd.n36 gnd 0.002701f
C1296 vdd.n37 gnd 0.006385f
C1297 vdd.n38 gnd 0.00286f
C1298 vdd.n39 gnd 0.005027f
C1299 vdd.n40 gnd 0.002701f
C1300 vdd.n41 gnd 0.004789f
C1301 vdd.n42 gnd 0.004803f
C1302 vdd.t83 gnd 0.013718f
C1303 vdd.n43 gnd 0.030521f
C1304 vdd.n44 gnd 0.158841f
C1305 vdd.n45 gnd 0.002701f
C1306 vdd.n46 gnd 0.00286f
C1307 vdd.n47 gnd 0.006385f
C1308 vdd.n48 gnd 0.006385f
C1309 vdd.n49 gnd 0.00286f
C1310 vdd.n50 gnd 0.002701f
C1311 vdd.n51 gnd 0.005027f
C1312 vdd.n52 gnd 0.005027f
C1313 vdd.n53 gnd 0.002701f
C1314 vdd.n54 gnd 0.00286f
C1315 vdd.n55 gnd 0.006385f
C1316 vdd.n56 gnd 0.006385f
C1317 vdd.n57 gnd 0.00286f
C1318 vdd.n58 gnd 0.002701f
C1319 vdd.n59 gnd 0.005027f
C1320 vdd.n60 gnd 0.005027f
C1321 vdd.n61 gnd 0.002701f
C1322 vdd.n62 gnd 0.00286f
C1323 vdd.n63 gnd 0.006385f
C1324 vdd.n64 gnd 0.006385f
C1325 vdd.n65 gnd 0.015096f
C1326 vdd.n66 gnd 0.002781f
C1327 vdd.n67 gnd 0.002701f
C1328 vdd.n68 gnd 0.012993f
C1329 vdd.n69 gnd 0.009071f
C1330 vdd.t35 gnd 0.031781f
C1331 vdd.t225 gnd 0.031781f
C1332 vdd.n70 gnd 0.218418f
C1333 vdd.n71 gnd 0.171752f
C1334 vdd.t71 gnd 0.031781f
C1335 vdd.t58 gnd 0.031781f
C1336 vdd.n72 gnd 0.218418f
C1337 vdd.n73 gnd 0.138603f
C1338 vdd.t190 gnd 0.031781f
C1339 vdd.t64 gnd 0.031781f
C1340 vdd.n74 gnd 0.218418f
C1341 vdd.n75 gnd 0.138603f
C1342 vdd.t68 gnd 0.031781f
C1343 vdd.t28 gnd 0.031781f
C1344 vdd.n76 gnd 0.218418f
C1345 vdd.n77 gnd 0.138603f
C1346 vdd.t184 gnd 0.031781f
C1347 vdd.t165 gnd 0.031781f
C1348 vdd.n78 gnd 0.218418f
C1349 vdd.n79 gnd 0.138603f
C1350 vdd.n80 gnd 0.005417f
C1351 vdd.n81 gnd 0.005027f
C1352 vdd.n82 gnd 0.002781f
C1353 vdd.n83 gnd 0.006385f
C1354 vdd.n84 gnd 0.002701f
C1355 vdd.n85 gnd 0.00286f
C1356 vdd.n86 gnd 0.005027f
C1357 vdd.n87 gnd 0.002701f
C1358 vdd.n88 gnd 0.006385f
C1359 vdd.n89 gnd 0.00286f
C1360 vdd.n90 gnd 0.005027f
C1361 vdd.n91 gnd 0.002701f
C1362 vdd.n92 gnd 0.004789f
C1363 vdd.n93 gnd 0.004803f
C1364 vdd.t5 gnd 0.013718f
C1365 vdd.n94 gnd 0.030521f
C1366 vdd.n95 gnd 0.158841f
C1367 vdd.n96 gnd 0.002701f
C1368 vdd.n97 gnd 0.00286f
C1369 vdd.n98 gnd 0.006385f
C1370 vdd.n99 gnd 0.006385f
C1371 vdd.n100 gnd 0.00286f
C1372 vdd.n101 gnd 0.002701f
C1373 vdd.n102 gnd 0.005027f
C1374 vdd.n103 gnd 0.005027f
C1375 vdd.n104 gnd 0.002701f
C1376 vdd.n105 gnd 0.00286f
C1377 vdd.n106 gnd 0.006385f
C1378 vdd.n107 gnd 0.006385f
C1379 vdd.n108 gnd 0.00286f
C1380 vdd.n109 gnd 0.002701f
C1381 vdd.n110 gnd 0.005027f
C1382 vdd.n111 gnd 0.005027f
C1383 vdd.n112 gnd 0.002701f
C1384 vdd.n113 gnd 0.00286f
C1385 vdd.n114 gnd 0.006385f
C1386 vdd.n115 gnd 0.006385f
C1387 vdd.n116 gnd 0.015096f
C1388 vdd.n117 gnd 0.002781f
C1389 vdd.n118 gnd 0.002701f
C1390 vdd.n119 gnd 0.012993f
C1391 vdd.n120 gnd 0.008787f
C1392 vdd.n121 gnd 0.103122f
C1393 vdd.n122 gnd 0.005417f
C1394 vdd.n123 gnd 0.005027f
C1395 vdd.n124 gnd 0.002781f
C1396 vdd.n125 gnd 0.006385f
C1397 vdd.n126 gnd 0.002701f
C1398 vdd.n127 gnd 0.00286f
C1399 vdd.n128 gnd 0.005027f
C1400 vdd.n129 gnd 0.002701f
C1401 vdd.n130 gnd 0.006385f
C1402 vdd.n131 gnd 0.00286f
C1403 vdd.n132 gnd 0.005027f
C1404 vdd.n133 gnd 0.002701f
C1405 vdd.n134 gnd 0.004789f
C1406 vdd.n135 gnd 0.004803f
C1407 vdd.t224 gnd 0.013718f
C1408 vdd.n136 gnd 0.030521f
C1409 vdd.n137 gnd 0.158841f
C1410 vdd.n138 gnd 0.002701f
C1411 vdd.n139 gnd 0.00286f
C1412 vdd.n140 gnd 0.006385f
C1413 vdd.n141 gnd 0.006385f
C1414 vdd.n142 gnd 0.00286f
C1415 vdd.n143 gnd 0.002701f
C1416 vdd.n144 gnd 0.005027f
C1417 vdd.n145 gnd 0.005027f
C1418 vdd.n146 gnd 0.002701f
C1419 vdd.n147 gnd 0.00286f
C1420 vdd.n148 gnd 0.006385f
C1421 vdd.n149 gnd 0.006385f
C1422 vdd.n150 gnd 0.00286f
C1423 vdd.n151 gnd 0.002701f
C1424 vdd.n152 gnd 0.005027f
C1425 vdd.n153 gnd 0.005027f
C1426 vdd.n154 gnd 0.002701f
C1427 vdd.n155 gnd 0.00286f
C1428 vdd.n156 gnd 0.006385f
C1429 vdd.n157 gnd 0.006385f
C1430 vdd.n158 gnd 0.015096f
C1431 vdd.n159 gnd 0.002781f
C1432 vdd.n160 gnd 0.002701f
C1433 vdd.n161 gnd 0.012993f
C1434 vdd.n162 gnd 0.009071f
C1435 vdd.t200 gnd 0.031781f
C1436 vdd.t214 gnd 0.031781f
C1437 vdd.n163 gnd 0.218418f
C1438 vdd.n164 gnd 0.171752f
C1439 vdd.t1 gnd 0.031781f
C1440 vdd.t229 gnd 0.031781f
C1441 vdd.n165 gnd 0.218418f
C1442 vdd.n166 gnd 0.138603f
C1443 vdd.t215 gnd 0.031781f
C1444 vdd.t172 gnd 0.031781f
C1445 vdd.n167 gnd 0.218418f
C1446 vdd.n168 gnd 0.138603f
C1447 vdd.t61 gnd 0.031781f
C1448 vdd.t59 gnd 0.031781f
C1449 vdd.n169 gnd 0.218418f
C1450 vdd.n170 gnd 0.138603f
C1451 vdd.t226 gnd 0.031781f
C1452 vdd.t164 gnd 0.031781f
C1453 vdd.n171 gnd 0.218418f
C1454 vdd.n172 gnd 0.138603f
C1455 vdd.n173 gnd 0.005417f
C1456 vdd.n174 gnd 0.005027f
C1457 vdd.n175 gnd 0.002781f
C1458 vdd.n176 gnd 0.006385f
C1459 vdd.n177 gnd 0.002701f
C1460 vdd.n178 gnd 0.00286f
C1461 vdd.n179 gnd 0.005027f
C1462 vdd.n180 gnd 0.002701f
C1463 vdd.n181 gnd 0.006385f
C1464 vdd.n182 gnd 0.00286f
C1465 vdd.n183 gnd 0.005027f
C1466 vdd.n184 gnd 0.002701f
C1467 vdd.n185 gnd 0.004789f
C1468 vdd.n186 gnd 0.004803f
C1469 vdd.t162 gnd 0.013718f
C1470 vdd.n187 gnd 0.030521f
C1471 vdd.n188 gnd 0.158841f
C1472 vdd.n189 gnd 0.002701f
C1473 vdd.n190 gnd 0.00286f
C1474 vdd.n191 gnd 0.006385f
C1475 vdd.n192 gnd 0.006385f
C1476 vdd.n193 gnd 0.00286f
C1477 vdd.n194 gnd 0.002701f
C1478 vdd.n195 gnd 0.005027f
C1479 vdd.n196 gnd 0.005027f
C1480 vdd.n197 gnd 0.002701f
C1481 vdd.n198 gnd 0.00286f
C1482 vdd.n199 gnd 0.006385f
C1483 vdd.n200 gnd 0.006385f
C1484 vdd.n201 gnd 0.00286f
C1485 vdd.n202 gnd 0.002701f
C1486 vdd.n203 gnd 0.005027f
C1487 vdd.n204 gnd 0.005027f
C1488 vdd.n205 gnd 0.002701f
C1489 vdd.n206 gnd 0.00286f
C1490 vdd.n207 gnd 0.006385f
C1491 vdd.n208 gnd 0.006385f
C1492 vdd.n209 gnd 0.015096f
C1493 vdd.n210 gnd 0.002781f
C1494 vdd.n211 gnd 0.002701f
C1495 vdd.n212 gnd 0.012993f
C1496 vdd.n213 gnd 0.008787f
C1497 vdd.n214 gnd 0.061347f
C1498 vdd.n215 gnd 0.221049f
C1499 vdd.n216 gnd 0.005417f
C1500 vdd.n217 gnd 0.005027f
C1501 vdd.n218 gnd 0.002781f
C1502 vdd.n219 gnd 0.006385f
C1503 vdd.n220 gnd 0.002701f
C1504 vdd.n221 gnd 0.00286f
C1505 vdd.n222 gnd 0.005027f
C1506 vdd.n223 gnd 0.002701f
C1507 vdd.n224 gnd 0.006385f
C1508 vdd.n225 gnd 0.00286f
C1509 vdd.n226 gnd 0.005027f
C1510 vdd.n227 gnd 0.002701f
C1511 vdd.n228 gnd 0.004789f
C1512 vdd.n229 gnd 0.004803f
C1513 vdd.t169 gnd 0.013718f
C1514 vdd.n230 gnd 0.030521f
C1515 vdd.n231 gnd 0.158841f
C1516 vdd.n232 gnd 0.002701f
C1517 vdd.n233 gnd 0.00286f
C1518 vdd.n234 gnd 0.006385f
C1519 vdd.n235 gnd 0.006385f
C1520 vdd.n236 gnd 0.00286f
C1521 vdd.n237 gnd 0.002701f
C1522 vdd.n238 gnd 0.005027f
C1523 vdd.n239 gnd 0.005027f
C1524 vdd.n240 gnd 0.002701f
C1525 vdd.n241 gnd 0.00286f
C1526 vdd.n242 gnd 0.006385f
C1527 vdd.n243 gnd 0.006385f
C1528 vdd.n244 gnd 0.00286f
C1529 vdd.n245 gnd 0.002701f
C1530 vdd.n246 gnd 0.005027f
C1531 vdd.n247 gnd 0.005027f
C1532 vdd.n248 gnd 0.002701f
C1533 vdd.n249 gnd 0.00286f
C1534 vdd.n250 gnd 0.006385f
C1535 vdd.n251 gnd 0.006385f
C1536 vdd.n252 gnd 0.015096f
C1537 vdd.n253 gnd 0.002781f
C1538 vdd.n254 gnd 0.002701f
C1539 vdd.n255 gnd 0.012993f
C1540 vdd.n256 gnd 0.009071f
C1541 vdd.t168 gnd 0.031781f
C1542 vdd.t218 gnd 0.031781f
C1543 vdd.n257 gnd 0.218418f
C1544 vdd.n258 gnd 0.171752f
C1545 vdd.t22 gnd 0.031781f
C1546 vdd.t65 gnd 0.031781f
C1547 vdd.n259 gnd 0.218418f
C1548 vdd.n260 gnd 0.138603f
C1549 vdd.t191 gnd 0.031781f
C1550 vdd.t230 gnd 0.031781f
C1551 vdd.n261 gnd 0.218418f
C1552 vdd.n262 gnd 0.138603f
C1553 vdd.t62 gnd 0.031781f
C1554 vdd.t25 gnd 0.031781f
C1555 vdd.n263 gnd 0.218418f
C1556 vdd.n264 gnd 0.138603f
C1557 vdd.t73 gnd 0.031781f
C1558 vdd.t195 gnd 0.031781f
C1559 vdd.n265 gnd 0.218418f
C1560 vdd.n266 gnd 0.138603f
C1561 vdd.n267 gnd 0.005417f
C1562 vdd.n268 gnd 0.005027f
C1563 vdd.n269 gnd 0.002781f
C1564 vdd.n270 gnd 0.006385f
C1565 vdd.n271 gnd 0.002701f
C1566 vdd.n272 gnd 0.00286f
C1567 vdd.n273 gnd 0.005027f
C1568 vdd.n274 gnd 0.002701f
C1569 vdd.n275 gnd 0.006385f
C1570 vdd.n276 gnd 0.00286f
C1571 vdd.n277 gnd 0.005027f
C1572 vdd.n278 gnd 0.002701f
C1573 vdd.n279 gnd 0.004789f
C1574 vdd.n280 gnd 0.004803f
C1575 vdd.t198 gnd 0.013718f
C1576 vdd.n281 gnd 0.030521f
C1577 vdd.n282 gnd 0.158841f
C1578 vdd.n283 gnd 0.002701f
C1579 vdd.n284 gnd 0.00286f
C1580 vdd.n285 gnd 0.006385f
C1581 vdd.n286 gnd 0.006385f
C1582 vdd.n287 gnd 0.00286f
C1583 vdd.n288 gnd 0.002701f
C1584 vdd.n289 gnd 0.005027f
C1585 vdd.n290 gnd 0.005027f
C1586 vdd.n291 gnd 0.002701f
C1587 vdd.n292 gnd 0.00286f
C1588 vdd.n293 gnd 0.006385f
C1589 vdd.n294 gnd 0.006385f
C1590 vdd.n295 gnd 0.00286f
C1591 vdd.n296 gnd 0.002701f
C1592 vdd.n297 gnd 0.005027f
C1593 vdd.n298 gnd 0.005027f
C1594 vdd.n299 gnd 0.002701f
C1595 vdd.n300 gnd 0.00286f
C1596 vdd.n301 gnd 0.006385f
C1597 vdd.n302 gnd 0.006385f
C1598 vdd.n303 gnd 0.015096f
C1599 vdd.n304 gnd 0.002781f
C1600 vdd.n305 gnd 0.002701f
C1601 vdd.n306 gnd 0.012993f
C1602 vdd.n307 gnd 0.008787f
C1603 vdd.n308 gnd 0.061347f
C1604 vdd.n309 gnd 0.24294f
C1605 vdd.n310 gnd 0.009837f
C1606 vdd.n311 gnd 0.009837f
C1607 vdd.n312 gnd 0.007945f
C1608 vdd.n313 gnd 0.007945f
C1609 vdd.n314 gnd 0.009871f
C1610 vdd.n315 gnd 0.009871f
C1611 vdd.t189 gnd 0.504397f
C1612 vdd.n316 gnd 0.009871f
C1613 vdd.n317 gnd 0.009871f
C1614 vdd.n318 gnd 0.009871f
C1615 vdd.t60 gnd 0.504397f
C1616 vdd.n319 gnd 0.009871f
C1617 vdd.n320 gnd 0.009871f
C1618 vdd.n321 gnd 0.009871f
C1619 vdd.n322 gnd 0.009871f
C1620 vdd.n323 gnd 0.007945f
C1621 vdd.n324 gnd 0.009871f
C1622 vdd.n325 gnd 0.812078f
C1623 vdd.n326 gnd 0.009871f
C1624 vdd.n327 gnd 0.009871f
C1625 vdd.n328 gnd 0.009871f
C1626 vdd.n329 gnd 0.691023f
C1627 vdd.n330 gnd 0.009871f
C1628 vdd.n331 gnd 0.009871f
C1629 vdd.n332 gnd 0.009871f
C1630 vdd.n333 gnd 0.009871f
C1631 vdd.n334 gnd 0.009871f
C1632 vdd.n335 gnd 0.007945f
C1633 vdd.n336 gnd 0.009871f
C1634 vdd.t163 gnd 0.504397f
C1635 vdd.n337 gnd 0.009871f
C1636 vdd.n338 gnd 0.009871f
C1637 vdd.n339 gnd 0.009871f
C1638 vdd.n340 gnd 1.00879f
C1639 vdd.n341 gnd 0.009871f
C1640 vdd.n342 gnd 0.009871f
C1641 vdd.n343 gnd 0.009871f
C1642 vdd.n344 gnd 0.009871f
C1643 vdd.n345 gnd 0.009871f
C1644 vdd.n346 gnd 0.007945f
C1645 vdd.n347 gnd 0.009871f
C1646 vdd.n348 gnd 0.009871f
C1647 vdd.n349 gnd 0.009871f
C1648 vdd.n350 gnd 0.023262f
C1649 vdd.n351 gnd 2.32022f
C1650 vdd.n352 gnd 0.023626f
C1651 vdd.n353 gnd 0.009871f
C1652 vdd.n354 gnd 0.009871f
C1653 vdd.n356 gnd 0.009871f
C1654 vdd.n357 gnd 0.009871f
C1655 vdd.n358 gnd 0.007945f
C1656 vdd.n359 gnd 0.007945f
C1657 vdd.n360 gnd 0.009871f
C1658 vdd.n361 gnd 0.009871f
C1659 vdd.n362 gnd 0.009871f
C1660 vdd.n363 gnd 0.009871f
C1661 vdd.n364 gnd 0.009871f
C1662 vdd.n365 gnd 0.009871f
C1663 vdd.n366 gnd 0.007945f
C1664 vdd.n368 gnd 0.009871f
C1665 vdd.n369 gnd 0.009871f
C1666 vdd.n370 gnd 0.009871f
C1667 vdd.n371 gnd 0.009871f
C1668 vdd.n372 gnd 0.009871f
C1669 vdd.n373 gnd 0.007945f
C1670 vdd.n375 gnd 0.009871f
C1671 vdd.n376 gnd 0.009871f
C1672 vdd.n377 gnd 0.009871f
C1673 vdd.n378 gnd 0.009871f
C1674 vdd.n379 gnd 0.009871f
C1675 vdd.n380 gnd 0.007945f
C1676 vdd.n382 gnd 0.009871f
C1677 vdd.n383 gnd 0.009871f
C1678 vdd.n384 gnd 0.009871f
C1679 vdd.n385 gnd 0.009871f
C1680 vdd.n386 gnd 0.006634f
C1681 vdd.t161 gnd 0.121442f
C1682 vdd.t160 gnd 0.129788f
C1683 vdd.t159 gnd 0.158602f
C1684 vdd.n387 gnd 0.203305f
C1685 vdd.n388 gnd 0.171608f
C1686 vdd.n390 gnd 0.009871f
C1687 vdd.n391 gnd 0.009871f
C1688 vdd.n392 gnd 0.007945f
C1689 vdd.n393 gnd 0.009871f
C1690 vdd.n395 gnd 0.009871f
C1691 vdd.n396 gnd 0.009871f
C1692 vdd.n397 gnd 0.009871f
C1693 vdd.n398 gnd 0.009871f
C1694 vdd.n399 gnd 0.007945f
C1695 vdd.n401 gnd 0.009871f
C1696 vdd.n402 gnd 0.009871f
C1697 vdd.n403 gnd 0.009871f
C1698 vdd.n404 gnd 0.009871f
C1699 vdd.n405 gnd 0.009871f
C1700 vdd.n406 gnd 0.007945f
C1701 vdd.n408 gnd 0.009871f
C1702 vdd.n409 gnd 0.009871f
C1703 vdd.n410 gnd 0.009871f
C1704 vdd.n411 gnd 0.009871f
C1705 vdd.n412 gnd 0.009871f
C1706 vdd.n413 gnd 0.007945f
C1707 vdd.n415 gnd 0.009871f
C1708 vdd.n416 gnd 0.009871f
C1709 vdd.n417 gnd 0.009871f
C1710 vdd.n418 gnd 0.009871f
C1711 vdd.n419 gnd 0.009871f
C1712 vdd.n420 gnd 0.007945f
C1713 vdd.n422 gnd 0.009871f
C1714 vdd.n423 gnd 0.009871f
C1715 vdd.n424 gnd 0.009871f
C1716 vdd.n425 gnd 0.009871f
C1717 vdd.n426 gnd 0.007866f
C1718 vdd.t149 gnd 0.121442f
C1719 vdd.t148 gnd 0.129788f
C1720 vdd.t146 gnd 0.158602f
C1721 vdd.n427 gnd 0.203305f
C1722 vdd.n428 gnd 0.171608f
C1723 vdd.n430 gnd 0.009871f
C1724 vdd.n431 gnd 0.009871f
C1725 vdd.n432 gnd 0.007945f
C1726 vdd.n433 gnd 0.009871f
C1727 vdd.n435 gnd 0.009871f
C1728 vdd.n436 gnd 0.009871f
C1729 vdd.n437 gnd 0.009871f
C1730 vdd.n438 gnd 0.009871f
C1731 vdd.n439 gnd 0.007945f
C1732 vdd.n441 gnd 0.009871f
C1733 vdd.n442 gnd 0.009871f
C1734 vdd.n443 gnd 0.009871f
C1735 vdd.n444 gnd 0.009871f
C1736 vdd.n445 gnd 0.009871f
C1737 vdd.n446 gnd 0.007945f
C1738 vdd.n448 gnd 0.009871f
C1739 vdd.n449 gnd 0.009871f
C1740 vdd.n450 gnd 0.009871f
C1741 vdd.n451 gnd 0.009871f
C1742 vdd.n452 gnd 0.009871f
C1743 vdd.n453 gnd 0.007945f
C1744 vdd.n455 gnd 0.009871f
C1745 vdd.n456 gnd 0.009871f
C1746 vdd.n457 gnd 0.009871f
C1747 vdd.n458 gnd 0.009871f
C1748 vdd.n459 gnd 0.009871f
C1749 vdd.n460 gnd 0.007945f
C1750 vdd.n462 gnd 0.009871f
C1751 vdd.n463 gnd 0.009871f
C1752 vdd.n464 gnd 0.009871f
C1753 vdd.n465 gnd 0.009871f
C1754 vdd.n466 gnd 0.009871f
C1755 vdd.n467 gnd 0.009871f
C1756 vdd.n468 gnd 0.007945f
C1757 vdd.n469 gnd 0.009871f
C1758 vdd.n470 gnd 0.009871f
C1759 vdd.n471 gnd 0.007945f
C1760 vdd.n472 gnd 0.009871f
C1761 vdd.n473 gnd 0.009871f
C1762 vdd.n474 gnd 0.007945f
C1763 vdd.n475 gnd 0.009871f
C1764 vdd.n476 gnd 0.007945f
C1765 vdd.n477 gnd 0.009871f
C1766 vdd.n478 gnd 0.007945f
C1767 vdd.n479 gnd 0.009871f
C1768 vdd.n480 gnd 0.009871f
C1769 vdd.t57 gnd 0.504397f
C1770 vdd.n481 gnd 0.539704f
C1771 vdd.n482 gnd 0.009871f
C1772 vdd.n483 gnd 0.007945f
C1773 vdd.n484 gnd 0.009871f
C1774 vdd.n485 gnd 0.007945f
C1775 vdd.n486 gnd 0.009871f
C1776 vdd.t0 gnd 0.504397f
C1777 vdd.n487 gnd 0.009871f
C1778 vdd.n488 gnd 0.007945f
C1779 vdd.n489 gnd 0.009871f
C1780 vdd.n490 gnd 0.007945f
C1781 vdd.n491 gnd 0.009871f
C1782 vdd.n492 gnd 0.791903f
C1783 vdd.n493 gnd 0.837298f
C1784 vdd.t213 gnd 0.504397f
C1785 vdd.n494 gnd 0.009871f
C1786 vdd.n495 gnd 0.007945f
C1787 vdd.n496 gnd 0.009871f
C1788 vdd.n497 gnd 0.007945f
C1789 vdd.n498 gnd 0.009871f
C1790 vdd.n499 gnd 0.620408f
C1791 vdd.n500 gnd 0.009871f
C1792 vdd.n501 gnd 0.007945f
C1793 vdd.n502 gnd 0.009871f
C1794 vdd.n503 gnd 0.007945f
C1795 vdd.n504 gnd 0.009871f
C1796 vdd.n505 gnd 1.00879f
C1797 vdd.t82 gnd 0.504397f
C1798 vdd.n506 gnd 0.009871f
C1799 vdd.n507 gnd 0.007945f
C1800 vdd.n508 gnd 0.009871f
C1801 vdd.n509 gnd 0.007945f
C1802 vdd.n510 gnd 0.009871f
C1803 vdd.n511 gnd 0.539704f
C1804 vdd.n512 gnd 0.009871f
C1805 vdd.n513 gnd 0.007945f
C1806 vdd.n514 gnd 0.023626f
C1807 vdd.n515 gnd 0.023626f
C1808 vdd.n516 gnd 7.22296f
C1809 vdd.t87 gnd 0.504397f
C1810 vdd.n517 gnd 0.023626f
C1811 vdd.n518 gnd 0.008489f
C1812 vdd.n519 gnd 0.007945f
C1813 vdd.n524 gnd 0.006318f
C1814 vdd.n525 gnd 0.007945f
C1815 vdd.n526 gnd 0.009871f
C1816 vdd.n527 gnd 0.009871f
C1817 vdd.n528 gnd 0.009871f
C1818 vdd.n529 gnd 0.009871f
C1819 vdd.n530 gnd 0.009871f
C1820 vdd.n531 gnd 0.007945f
C1821 vdd.n532 gnd 0.009871f
C1822 vdd.n533 gnd 0.009871f
C1823 vdd.n534 gnd 0.009871f
C1824 vdd.n535 gnd 0.009871f
C1825 vdd.n536 gnd 0.009871f
C1826 vdd.n537 gnd 0.007945f
C1827 vdd.n538 gnd 0.009871f
C1828 vdd.n539 gnd 0.009871f
C1829 vdd.n540 gnd 0.009871f
C1830 vdd.n541 gnd 0.009871f
C1831 vdd.n542 gnd 0.009871f
C1832 vdd.t91 gnd 0.121442f
C1833 vdd.t92 gnd 0.129788f
C1834 vdd.t90 gnd 0.158602f
C1835 vdd.n543 gnd 0.203305f
C1836 vdd.n544 gnd 0.170813f
C1837 vdd.n545 gnd 0.016208f
C1838 vdd.n546 gnd 0.009871f
C1839 vdd.n547 gnd 0.009871f
C1840 vdd.n548 gnd 0.009871f
C1841 vdd.n549 gnd 0.009871f
C1842 vdd.n550 gnd 0.009871f
C1843 vdd.n551 gnd 0.007945f
C1844 vdd.n552 gnd 0.009871f
C1845 vdd.n553 gnd 0.009871f
C1846 vdd.n554 gnd 0.009871f
C1847 vdd.n555 gnd 0.009871f
C1848 vdd.n556 gnd 0.009871f
C1849 vdd.n557 gnd 0.007945f
C1850 vdd.n558 gnd 0.009871f
C1851 vdd.n559 gnd 0.009871f
C1852 vdd.n560 gnd 0.009871f
C1853 vdd.n561 gnd 0.009871f
C1854 vdd.n562 gnd 0.009871f
C1855 vdd.n563 gnd 0.007945f
C1856 vdd.n564 gnd 0.009871f
C1857 vdd.n565 gnd 0.009871f
C1858 vdd.n566 gnd 0.009871f
C1859 vdd.n567 gnd 0.009871f
C1860 vdd.n568 gnd 0.009871f
C1861 vdd.n569 gnd 0.007945f
C1862 vdd.n570 gnd 0.009871f
C1863 vdd.n571 gnd 0.009871f
C1864 vdd.n572 gnd 0.009871f
C1865 vdd.n573 gnd 0.009871f
C1866 vdd.n574 gnd 0.009871f
C1867 vdd.n575 gnd 0.007945f
C1868 vdd.n576 gnd 0.009871f
C1869 vdd.n577 gnd 0.009871f
C1870 vdd.n578 gnd 0.009871f
C1871 vdd.n579 gnd 0.007866f
C1872 vdd.t88 gnd 0.121442f
C1873 vdd.t89 gnd 0.129788f
C1874 vdd.t86 gnd 0.158602f
C1875 vdd.n580 gnd 0.203305f
C1876 vdd.n581 gnd 0.170813f
C1877 vdd.n582 gnd 0.009871f
C1878 vdd.n583 gnd 0.007945f
C1879 vdd.n585 gnd 0.009871f
C1880 vdd.n587 gnd 0.009871f
C1881 vdd.n588 gnd 0.009871f
C1882 vdd.n589 gnd 0.007945f
C1883 vdd.n590 gnd 0.009871f
C1884 vdd.n591 gnd 0.009871f
C1885 vdd.n592 gnd 0.009871f
C1886 vdd.n593 gnd 0.009871f
C1887 vdd.n594 gnd 0.009871f
C1888 vdd.n595 gnd 0.007945f
C1889 vdd.n596 gnd 0.009871f
C1890 vdd.n597 gnd 0.009871f
C1891 vdd.n598 gnd 0.009871f
C1892 vdd.n599 gnd 0.009871f
C1893 vdd.n600 gnd 0.009871f
C1894 vdd.n601 gnd 0.007945f
C1895 vdd.n602 gnd 0.009871f
C1896 vdd.n603 gnd 0.009871f
C1897 vdd.n604 gnd 0.009871f
C1898 vdd.n605 gnd 0.006318f
C1899 vdd.n610 gnd 0.006712f
C1900 vdd.n611 gnd 0.006712f
C1901 vdd.n612 gnd 0.006712f
C1902 vdd.n613 gnd 6.95058f
C1903 vdd.n614 gnd 0.006712f
C1904 vdd.n615 gnd 0.006712f
C1905 vdd.n616 gnd 0.006712f
C1906 vdd.n618 gnd 0.006712f
C1907 vdd.n619 gnd 0.006712f
C1908 vdd.n621 gnd 0.006712f
C1909 vdd.n622 gnd 0.004886f
C1910 vdd.n624 gnd 0.006712f
C1911 vdd.t128 gnd 0.271249f
C1912 vdd.t127 gnd 0.277657f
C1913 vdd.t126 gnd 0.177082f
C1914 vdd.n625 gnd 0.095703f
C1915 vdd.n626 gnd 0.054286f
C1916 vdd.n627 gnd 0.009593f
C1917 vdd.n628 gnd 0.015688f
C1918 vdd.n630 gnd 0.006712f
C1919 vdd.n631 gnd 0.685979f
C1920 vdd.n632 gnd 0.014871f
C1921 vdd.n633 gnd 0.014871f
C1922 vdd.n634 gnd 0.006712f
C1923 vdd.n635 gnd 0.015927f
C1924 vdd.n636 gnd 0.006712f
C1925 vdd.n637 gnd 0.006712f
C1926 vdd.n638 gnd 0.006712f
C1927 vdd.n639 gnd 0.006712f
C1928 vdd.n640 gnd 0.006712f
C1929 vdd.n642 gnd 0.006712f
C1930 vdd.n643 gnd 0.006712f
C1931 vdd.n645 gnd 0.006712f
C1932 vdd.n646 gnd 0.006712f
C1933 vdd.n648 gnd 0.006712f
C1934 vdd.n649 gnd 0.006712f
C1935 vdd.n651 gnd 0.006712f
C1936 vdd.n652 gnd 0.006712f
C1937 vdd.n654 gnd 0.006712f
C1938 vdd.n655 gnd 0.006712f
C1939 vdd.n657 gnd 0.006712f
C1940 vdd.n658 gnd 0.004886f
C1941 vdd.n660 gnd 0.006712f
C1942 vdd.t121 gnd 0.271249f
C1943 vdd.t120 gnd 0.277657f
C1944 vdd.t118 gnd 0.177082f
C1945 vdd.n661 gnd 0.095703f
C1946 vdd.n662 gnd 0.054286f
C1947 vdd.n663 gnd 0.009593f
C1948 vdd.n664 gnd 0.006712f
C1949 vdd.n665 gnd 0.006712f
C1950 vdd.t119 gnd 0.34299f
C1951 vdd.n666 gnd 0.006712f
C1952 vdd.n667 gnd 0.006712f
C1953 vdd.n668 gnd 0.006712f
C1954 vdd.n669 gnd 0.006712f
C1955 vdd.n670 gnd 0.006712f
C1956 vdd.n671 gnd 0.685979f
C1957 vdd.n672 gnd 0.006712f
C1958 vdd.n673 gnd 0.006712f
C1959 vdd.n674 gnd 0.600232f
C1960 vdd.n675 gnd 0.006712f
C1961 vdd.n676 gnd 0.006712f
C1962 vdd.n677 gnd 0.005923f
C1963 vdd.n678 gnd 0.006712f
C1964 vdd.n679 gnd 0.605276f
C1965 vdd.n680 gnd 0.006712f
C1966 vdd.n681 gnd 0.006712f
C1967 vdd.n682 gnd 0.006712f
C1968 vdd.n683 gnd 0.006712f
C1969 vdd.n684 gnd 0.006712f
C1970 vdd.n685 gnd 0.685979f
C1971 vdd.n686 gnd 0.006712f
C1972 vdd.n687 gnd 0.006712f
C1973 vdd.t102 gnd 0.307682f
C1974 vdd.t79 gnd 0.080703f
C1975 vdd.n688 gnd 0.006712f
C1976 vdd.n689 gnd 0.006712f
C1977 vdd.n690 gnd 0.006712f
C1978 vdd.t192 gnd 0.34299f
C1979 vdd.n691 gnd 0.006712f
C1980 vdd.n692 gnd 0.006712f
C1981 vdd.n693 gnd 0.006712f
C1982 vdd.n694 gnd 0.006712f
C1983 vdd.n695 gnd 0.006712f
C1984 vdd.t181 gnd 0.34299f
C1985 vdd.n696 gnd 0.006712f
C1986 vdd.n697 gnd 0.006712f
C1987 vdd.n698 gnd 0.569968f
C1988 vdd.n699 gnd 0.006712f
C1989 vdd.n700 gnd 0.006712f
C1990 vdd.n701 gnd 0.006712f
C1991 vdd.n702 gnd 0.418649f
C1992 vdd.n703 gnd 0.006712f
C1993 vdd.n704 gnd 0.006712f
C1994 vdd.t205 gnd 0.34299f
C1995 vdd.n705 gnd 0.006712f
C1996 vdd.n706 gnd 0.006712f
C1997 vdd.n707 gnd 0.006712f
C1998 vdd.n708 gnd 0.569968f
C1999 vdd.n709 gnd 0.006712f
C2000 vdd.n710 gnd 0.006712f
C2001 vdd.t175 gnd 0.29255f
C2002 vdd.t14 gnd 0.26733f
C2003 vdd.n711 gnd 0.006712f
C2004 vdd.n712 gnd 0.006712f
C2005 vdd.n713 gnd 0.006712f
C2006 vdd.t19 gnd 0.34299f
C2007 vdd.n714 gnd 0.006712f
C2008 vdd.n715 gnd 0.006712f
C2009 vdd.t21 gnd 0.34299f
C2010 vdd.n716 gnd 0.006712f
C2011 vdd.n717 gnd 0.006712f
C2012 vdd.n718 gnd 0.006712f
C2013 vdd.t76 gnd 0.252198f
C2014 vdd.n719 gnd 0.006712f
C2015 vdd.n720 gnd 0.006712f
C2016 vdd.n721 gnd 0.5851f
C2017 vdd.n722 gnd 0.006712f
C2018 vdd.n723 gnd 0.006712f
C2019 vdd.n724 gnd 0.006712f
C2020 vdd.n725 gnd 0.685979f
C2021 vdd.n726 gnd 0.006712f
C2022 vdd.n727 gnd 0.006712f
C2023 vdd.t80 gnd 0.307682f
C2024 vdd.n728 gnd 0.433781f
C2025 vdd.n729 gnd 0.006712f
C2026 vdd.n730 gnd 0.006712f
C2027 vdd.n731 gnd 0.006712f
C2028 vdd.t74 gnd 0.34299f
C2029 vdd.n732 gnd 0.006712f
C2030 vdd.n733 gnd 0.006712f
C2031 vdd.n734 gnd 0.006712f
C2032 vdd.n735 gnd 0.006712f
C2033 vdd.n736 gnd 0.006712f
C2034 vdd.t209 gnd 0.685979f
C2035 vdd.n737 gnd 0.006712f
C2036 vdd.n738 gnd 0.006712f
C2037 vdd.t123 gnd 0.34299f
C2038 vdd.n739 gnd 0.006712f
C2039 vdd.n740 gnd 0.015927f
C2040 vdd.n741 gnd 0.015927f
C2041 vdd.t211 gnd 0.645628f
C2042 vdd.n742 gnd 0.014871f
C2043 vdd.n743 gnd 0.014871f
C2044 vdd.n744 gnd 0.015927f
C2045 vdd.n745 gnd 0.006712f
C2046 vdd.n746 gnd 0.006712f
C2047 vdd.t17 gnd 0.645628f
C2048 vdd.n764 gnd 0.015927f
C2049 vdd.n782 gnd 0.014871f
C2050 vdd.n783 gnd 0.006712f
C2051 vdd.n784 gnd 0.014871f
C2052 vdd.t142 gnd 0.271249f
C2053 vdd.t141 gnd 0.277657f
C2054 vdd.t140 gnd 0.177082f
C2055 vdd.n785 gnd 0.095703f
C2056 vdd.n786 gnd 0.054286f
C2057 vdd.n787 gnd 0.015688f
C2058 vdd.n788 gnd 0.006712f
C2059 vdd.t182 gnd 0.685979f
C2060 vdd.n789 gnd 0.014871f
C2061 vdd.n790 gnd 0.006712f
C2062 vdd.n791 gnd 0.015927f
C2063 vdd.n792 gnd 0.006712f
C2064 vdd.t117 gnd 0.271249f
C2065 vdd.t116 gnd 0.277657f
C2066 vdd.t114 gnd 0.177082f
C2067 vdd.n793 gnd 0.095703f
C2068 vdd.n794 gnd 0.054286f
C2069 vdd.n795 gnd 0.009593f
C2070 vdd.n796 gnd 0.006712f
C2071 vdd.n797 gnd 0.006712f
C2072 vdd.t115 gnd 0.34299f
C2073 vdd.n798 gnd 0.006712f
C2074 vdd.n799 gnd 0.006712f
C2075 vdd.n800 gnd 0.006712f
C2076 vdd.n801 gnd 0.006712f
C2077 vdd.n802 gnd 0.006712f
C2078 vdd.n803 gnd 0.006712f
C2079 vdd.n804 gnd 0.685979f
C2080 vdd.n805 gnd 0.006712f
C2081 vdd.n806 gnd 0.006712f
C2082 vdd.t203 gnd 0.34299f
C2083 vdd.n807 gnd 0.006712f
C2084 vdd.n808 gnd 0.006712f
C2085 vdd.n809 gnd 0.006712f
C2086 vdd.n810 gnd 0.006712f
C2087 vdd.n811 gnd 0.433781f
C2088 vdd.n812 gnd 0.006712f
C2089 vdd.n813 gnd 0.006712f
C2090 vdd.n814 gnd 0.006712f
C2091 vdd.n815 gnd 0.006712f
C2092 vdd.n816 gnd 0.006712f
C2093 vdd.n817 gnd 0.5851f
C2094 vdd.n818 gnd 0.006712f
C2095 vdd.n819 gnd 0.006712f
C2096 vdd.t178 gnd 0.307682f
C2097 vdd.t180 gnd 0.252198f
C2098 vdd.n820 gnd 0.006712f
C2099 vdd.n821 gnd 0.006712f
C2100 vdd.n822 gnd 0.006712f
C2101 vdd.t38 gnd 0.34299f
C2102 vdd.n823 gnd 0.006712f
C2103 vdd.n824 gnd 0.006712f
C2104 vdd.t12 gnd 0.34299f
C2105 vdd.n825 gnd 0.006712f
C2106 vdd.n826 gnd 0.006712f
C2107 vdd.n827 gnd 0.006712f
C2108 vdd.t207 gnd 0.26733f
C2109 vdd.n828 gnd 0.006712f
C2110 vdd.n829 gnd 0.006712f
C2111 vdd.n830 gnd 0.569968f
C2112 vdd.n831 gnd 0.006712f
C2113 vdd.n832 gnd 0.006712f
C2114 vdd.n833 gnd 0.006712f
C2115 vdd.t220 gnd 0.34299f
C2116 vdd.n834 gnd 0.006712f
C2117 vdd.n835 gnd 0.006712f
C2118 vdd.t37 gnd 0.29255f
C2119 vdd.n836 gnd 0.418649f
C2120 vdd.n837 gnd 0.006712f
C2121 vdd.n838 gnd 0.006712f
C2122 vdd.n839 gnd 0.006712f
C2123 vdd.n840 gnd 0.569968f
C2124 vdd.n841 gnd 0.006712f
C2125 vdd.n842 gnd 0.006712f
C2126 vdd.t85 gnd 0.34299f
C2127 vdd.n843 gnd 0.006712f
C2128 vdd.n844 gnd 0.006712f
C2129 vdd.n845 gnd 0.006712f
C2130 vdd.n846 gnd 0.685979f
C2131 vdd.n847 gnd 0.006712f
C2132 vdd.n848 gnd 0.006712f
C2133 vdd.t16 gnd 0.34299f
C2134 vdd.n849 gnd 0.006712f
C2135 vdd.n850 gnd 0.006712f
C2136 vdd.n851 gnd 0.006712f
C2137 vdd.t174 gnd 0.080703f
C2138 vdd.n852 gnd 0.006712f
C2139 vdd.n853 gnd 0.006712f
C2140 vdd.n854 gnd 0.006712f
C2141 vdd.t135 gnd 0.277657f
C2142 vdd.t133 gnd 0.177082f
C2143 vdd.t136 gnd 0.277657f
C2144 vdd.n855 gnd 0.156054f
C2145 vdd.n856 gnd 0.006712f
C2146 vdd.n857 gnd 0.006712f
C2147 vdd.n858 gnd 0.685979f
C2148 vdd.n859 gnd 0.006712f
C2149 vdd.n860 gnd 0.006712f
C2150 vdd.t134 gnd 0.307682f
C2151 vdd.n861 gnd 0.605276f
C2152 vdd.n862 gnd 0.006712f
C2153 vdd.n863 gnd 0.006712f
C2154 vdd.n864 gnd 0.006712f
C2155 vdd.n865 gnd 0.600232f
C2156 vdd.n866 gnd 0.006712f
C2157 vdd.n867 gnd 0.006712f
C2158 vdd.n868 gnd 0.006712f
C2159 vdd.n869 gnd 0.006712f
C2160 vdd.n870 gnd 0.006712f
C2161 vdd.n871 gnd 0.685979f
C2162 vdd.n872 gnd 0.006712f
C2163 vdd.n873 gnd 0.006712f
C2164 vdd.t130 gnd 0.34299f
C2165 vdd.n874 gnd 0.006712f
C2166 vdd.n875 gnd 0.015927f
C2167 vdd.n876 gnd 0.015927f
C2168 vdd.n877 gnd 6.95058f
C2169 vdd.n878 gnd 0.014871f
C2170 vdd.n879 gnd 0.014871f
C2171 vdd.n880 gnd 0.015927f
C2172 vdd.n881 gnd 0.006712f
C2173 vdd.n882 gnd 0.006712f
C2174 vdd.n883 gnd 0.006712f
C2175 vdd.n884 gnd 0.006712f
C2176 vdd.n885 gnd 0.006712f
C2177 vdd.n886 gnd 0.006712f
C2178 vdd.n887 gnd 0.006712f
C2179 vdd.n888 gnd 0.006712f
C2180 vdd.n890 gnd 0.006712f
C2181 vdd.n891 gnd 0.006712f
C2182 vdd.n892 gnd 0.006318f
C2183 vdd.n895 gnd 0.023626f
C2184 vdd.n896 gnd 0.007945f
C2185 vdd.n897 gnd 0.009871f
C2186 vdd.n899 gnd 0.009871f
C2187 vdd.n900 gnd 0.006594f
C2188 vdd.t94 gnd 0.504397f
C2189 vdd.n901 gnd 7.22296f
C2190 vdd.n902 gnd 0.009871f
C2191 vdd.n903 gnd 0.023626f
C2192 vdd.n904 gnd 0.007945f
C2193 vdd.n905 gnd 0.009871f
C2194 vdd.n906 gnd 0.007945f
C2195 vdd.n907 gnd 0.009871f
C2196 vdd.n908 gnd 1.00879f
C2197 vdd.n909 gnd 0.009871f
C2198 vdd.n910 gnd 0.007945f
C2199 vdd.n911 gnd 0.007945f
C2200 vdd.n912 gnd 0.009871f
C2201 vdd.n913 gnd 0.007945f
C2202 vdd.n914 gnd 0.009871f
C2203 vdd.t8 gnd 0.504397f
C2204 vdd.n915 gnd 0.009871f
C2205 vdd.n916 gnd 0.007945f
C2206 vdd.n917 gnd 0.009871f
C2207 vdd.n918 gnd 0.007945f
C2208 vdd.n919 gnd 0.009871f
C2209 vdd.t10 gnd 0.504397f
C2210 vdd.n920 gnd 0.009871f
C2211 vdd.n921 gnd 0.007945f
C2212 vdd.n922 gnd 0.009871f
C2213 vdd.n923 gnd 0.007945f
C2214 vdd.n924 gnd 0.009871f
C2215 vdd.t6 gnd 0.504397f
C2216 vdd.n925 gnd 0.791903f
C2217 vdd.n926 gnd 0.009871f
C2218 vdd.n927 gnd 0.007945f
C2219 vdd.n928 gnd 0.009871f
C2220 vdd.n929 gnd 0.007945f
C2221 vdd.n930 gnd 0.009871f
C2222 vdd.n931 gnd 0.711199f
C2223 vdd.n932 gnd 0.009871f
C2224 vdd.n933 gnd 0.007945f
C2225 vdd.n934 gnd 0.009871f
C2226 vdd.n935 gnd 0.007945f
C2227 vdd.n936 gnd 0.009871f
C2228 vdd.n937 gnd 0.539704f
C2229 vdd.t32 gnd 0.504397f
C2230 vdd.n938 gnd 0.009871f
C2231 vdd.n939 gnd 0.007945f
C2232 vdd.n940 gnd 0.009837f
C2233 vdd.n941 gnd 0.007945f
C2234 vdd.n942 gnd 0.009871f
C2235 vdd.t26 gnd 0.504397f
C2236 vdd.n943 gnd 0.009871f
C2237 vdd.n944 gnd 0.007945f
C2238 vdd.n945 gnd 0.009871f
C2239 vdd.n946 gnd 0.007945f
C2240 vdd.n947 gnd 0.009871f
C2241 vdd.t69 gnd 0.504397f
C2242 vdd.n948 gnd 0.640584f
C2243 vdd.n949 gnd 0.009871f
C2244 vdd.n950 gnd 0.007945f
C2245 vdd.n951 gnd 0.009871f
C2246 vdd.n952 gnd 0.007945f
C2247 vdd.n953 gnd 0.009871f
C2248 vdd.t66 gnd 0.504397f
C2249 vdd.n954 gnd 0.009871f
C2250 vdd.n955 gnd 0.007945f
C2251 vdd.n956 gnd 0.009871f
C2252 vdd.n957 gnd 0.007945f
C2253 vdd.n958 gnd 0.009871f
C2254 vdd.n959 gnd 0.691023f
C2255 vdd.n960 gnd 0.837298f
C2256 vdd.t55 gnd 0.504397f
C2257 vdd.n961 gnd 0.009871f
C2258 vdd.n962 gnd 0.007945f
C2259 vdd.n963 gnd 0.009871f
C2260 vdd.n964 gnd 0.007945f
C2261 vdd.n965 gnd 0.009871f
C2262 vdd.n966 gnd 0.519529f
C2263 vdd.n967 gnd 0.009871f
C2264 vdd.n968 gnd 0.007945f
C2265 vdd.n969 gnd 0.009871f
C2266 vdd.n970 gnd 0.007945f
C2267 vdd.n971 gnd 0.009871f
C2268 vdd.n972 gnd 1.00879f
C2269 vdd.t186 gnd 0.504397f
C2270 vdd.n973 gnd 0.009871f
C2271 vdd.n974 gnd 0.007945f
C2272 vdd.n975 gnd 0.009871f
C2273 vdd.n976 gnd 0.007945f
C2274 vdd.n977 gnd 0.009871f
C2275 vdd.t98 gnd 0.504397f
C2276 vdd.n978 gnd 0.009871f
C2277 vdd.n979 gnd 0.007945f
C2278 vdd.n980 gnd 0.023626f
C2279 vdd.n981 gnd 0.023626f
C2280 vdd.n982 gnd 2.32022f
C2281 vdd.n983 gnd 0.569968f
C2282 vdd.n984 gnd 0.023626f
C2283 vdd.n985 gnd 0.009871f
C2284 vdd.n987 gnd 0.009871f
C2285 vdd.n988 gnd 0.009871f
C2286 vdd.n989 gnd 0.007945f
C2287 vdd.n990 gnd 0.009871f
C2288 vdd.n991 gnd 0.009871f
C2289 vdd.n993 gnd 0.009871f
C2290 vdd.n994 gnd 0.009871f
C2291 vdd.n996 gnd 0.009871f
C2292 vdd.n997 gnd 0.007945f
C2293 vdd.n998 gnd 0.009871f
C2294 vdd.n999 gnd 0.009871f
C2295 vdd.n1001 gnd 0.009871f
C2296 vdd.n1002 gnd 0.009871f
C2297 vdd.n1004 gnd 0.009871f
C2298 vdd.n1005 gnd 0.007945f
C2299 vdd.n1006 gnd 0.009871f
C2300 vdd.n1007 gnd 0.009871f
C2301 vdd.n1009 gnd 0.009871f
C2302 vdd.n1010 gnd 0.009871f
C2303 vdd.n1012 gnd 0.009871f
C2304 vdd.n1013 gnd 0.007945f
C2305 vdd.n1014 gnd 0.009871f
C2306 vdd.n1015 gnd 0.009871f
C2307 vdd.n1017 gnd 0.009871f
C2308 vdd.n1018 gnd 0.009871f
C2309 vdd.n1020 gnd 0.009871f
C2310 vdd.t109 gnd 0.121442f
C2311 vdd.t110 gnd 0.129788f
C2312 vdd.t108 gnd 0.158602f
C2313 vdd.n1021 gnd 0.203305f
C2314 vdd.n1022 gnd 0.171608f
C2315 vdd.n1023 gnd 0.017003f
C2316 vdd.n1024 gnd 0.009871f
C2317 vdd.n1025 gnd 0.009871f
C2318 vdd.n1027 gnd 0.009871f
C2319 vdd.n1028 gnd 0.009871f
C2320 vdd.n1030 gnd 0.009871f
C2321 vdd.n1031 gnd 0.007945f
C2322 vdd.n1032 gnd 0.009871f
C2323 vdd.n1033 gnd 0.009871f
C2324 vdd.n1035 gnd 0.009871f
C2325 vdd.n1036 gnd 0.009871f
C2326 vdd.n1038 gnd 0.009871f
C2327 vdd.n1039 gnd 0.007945f
C2328 vdd.n1040 gnd 0.009871f
C2329 vdd.n1041 gnd 0.009871f
C2330 vdd.n1043 gnd 0.009871f
C2331 vdd.n1044 gnd 0.009871f
C2332 vdd.n1046 gnd 0.009871f
C2333 vdd.n1047 gnd 0.007945f
C2334 vdd.n1048 gnd 0.009871f
C2335 vdd.n1049 gnd 0.009871f
C2336 vdd.n1051 gnd 0.009871f
C2337 vdd.n1052 gnd 0.009871f
C2338 vdd.n1054 gnd 0.009871f
C2339 vdd.n1055 gnd 0.007945f
C2340 vdd.n1056 gnd 0.009871f
C2341 vdd.n1057 gnd 0.009871f
C2342 vdd.n1059 gnd 0.009871f
C2343 vdd.n1060 gnd 0.009871f
C2344 vdd.n1062 gnd 0.009871f
C2345 vdd.n1063 gnd 0.007945f
C2346 vdd.n1064 gnd 0.009871f
C2347 vdd.n1065 gnd 0.009871f
C2348 vdd.n1067 gnd 0.009871f
C2349 vdd.n1068 gnd 0.007866f
C2350 vdd.n1070 gnd 0.007945f
C2351 vdd.n1071 gnd 0.009871f
C2352 vdd.n1072 gnd 0.009871f
C2353 vdd.n1073 gnd 0.009871f
C2354 vdd.n1074 gnd 0.009871f
C2355 vdd.n1076 gnd 0.009871f
C2356 vdd.n1077 gnd 0.009871f
C2357 vdd.n1078 gnd 0.007945f
C2358 vdd.n1079 gnd 0.009871f
C2359 vdd.n1081 gnd 0.009871f
C2360 vdd.n1082 gnd 0.009871f
C2361 vdd.n1084 gnd 0.009871f
C2362 vdd.n1085 gnd 0.009871f
C2363 vdd.n1086 gnd 0.007945f
C2364 vdd.n1087 gnd 0.009871f
C2365 vdd.n1089 gnd 0.009871f
C2366 vdd.n1090 gnd 0.009871f
C2367 vdd.n1092 gnd 0.009871f
C2368 vdd.n1093 gnd 0.009871f
C2369 vdd.n1094 gnd 0.007945f
C2370 vdd.n1095 gnd 0.009871f
C2371 vdd.n1097 gnd 0.009871f
C2372 vdd.n1098 gnd 0.009871f
C2373 vdd.n1100 gnd 0.009871f
C2374 vdd.n1101 gnd 0.009871f
C2375 vdd.n1102 gnd 0.007945f
C2376 vdd.n1103 gnd 0.009871f
C2377 vdd.n1105 gnd 0.009871f
C2378 vdd.n1106 gnd 0.009871f
C2379 vdd.n1108 gnd 0.009871f
C2380 vdd.n1109 gnd 0.003774f
C2381 vdd.t151 gnd 0.121442f
C2382 vdd.t152 gnd 0.129788f
C2383 vdd.t150 gnd 0.158602f
C2384 vdd.n1110 gnd 0.203305f
C2385 vdd.n1111 gnd 0.171608f
C2386 vdd.n1112 gnd 0.01303f
C2387 vdd.n1113 gnd 0.004171f
C2388 vdd.n1114 gnd 0.007945f
C2389 vdd.n1115 gnd 0.009871f
C2390 vdd.n1116 gnd 0.009871f
C2391 vdd.n1117 gnd 0.009871f
C2392 vdd.n1118 gnd 0.007945f
C2393 vdd.n1119 gnd 0.007945f
C2394 vdd.n1120 gnd 0.007945f
C2395 vdd.n1121 gnd 0.009871f
C2396 vdd.n1122 gnd 0.009871f
C2397 vdd.n1123 gnd 0.009871f
C2398 vdd.n1124 gnd 0.007945f
C2399 vdd.n1125 gnd 0.007945f
C2400 vdd.n1126 gnd 0.007945f
C2401 vdd.n1127 gnd 0.009871f
C2402 vdd.n1128 gnd 0.009871f
C2403 vdd.n1129 gnd 0.009871f
C2404 vdd.n1130 gnd 0.007945f
C2405 vdd.n1131 gnd 0.007945f
C2406 vdd.n1132 gnd 0.007945f
C2407 vdd.n1133 gnd 0.009871f
C2408 vdd.n1134 gnd 0.009871f
C2409 vdd.n1135 gnd 0.009871f
C2410 vdd.n1136 gnd 0.007945f
C2411 vdd.n1137 gnd 0.007945f
C2412 vdd.n1138 gnd 0.007945f
C2413 vdd.n1139 gnd 0.009871f
C2414 vdd.n1140 gnd 0.009871f
C2415 vdd.n1141 gnd 0.009871f
C2416 vdd.n1142 gnd 0.007945f
C2417 vdd.n1143 gnd 0.009871f
C2418 vdd.n1144 gnd 0.009871f
C2419 vdd.n1146 gnd 0.009871f
C2420 vdd.t99 gnd 0.121442f
C2421 vdd.t100 gnd 0.129788f
C2422 vdd.t97 gnd 0.158602f
C2423 vdd.n1147 gnd 0.203305f
C2424 vdd.n1148 gnd 0.171608f
C2425 vdd.n1149 gnd 0.017003f
C2426 vdd.n1150 gnd 0.005403f
C2427 vdd.n1151 gnd 0.009871f
C2428 vdd.n1152 gnd 0.009871f
C2429 vdd.n1153 gnd 0.009871f
C2430 vdd.n1154 gnd 0.007945f
C2431 vdd.n1155 gnd 0.007945f
C2432 vdd.n1156 gnd 0.007945f
C2433 vdd.n1157 gnd 0.009871f
C2434 vdd.n1158 gnd 0.009871f
C2435 vdd.n1159 gnd 0.009871f
C2436 vdd.n1160 gnd 0.007945f
C2437 vdd.n1161 gnd 0.007945f
C2438 vdd.n1162 gnd 0.007945f
C2439 vdd.n1163 gnd 0.009871f
C2440 vdd.n1164 gnd 0.009871f
C2441 vdd.n1165 gnd 0.009871f
C2442 vdd.n1166 gnd 0.007945f
C2443 vdd.n1167 gnd 0.007945f
C2444 vdd.n1168 gnd 0.007945f
C2445 vdd.n1169 gnd 0.009871f
C2446 vdd.n1170 gnd 0.009871f
C2447 vdd.n1171 gnd 0.009871f
C2448 vdd.n1172 gnd 0.007945f
C2449 vdd.n1173 gnd 0.007945f
C2450 vdd.n1174 gnd 0.007945f
C2451 vdd.n1175 gnd 0.009871f
C2452 vdd.n1176 gnd 0.009871f
C2453 vdd.n1177 gnd 0.009871f
C2454 vdd.n1178 gnd 0.007945f
C2455 vdd.n1179 gnd 0.007945f
C2456 vdd.n1180 gnd 0.006634f
C2457 vdd.n1181 gnd 0.009871f
C2458 vdd.n1182 gnd 0.009871f
C2459 vdd.n1183 gnd 0.009871f
C2460 vdd.n1184 gnd 0.006634f
C2461 vdd.n1185 gnd 0.007945f
C2462 vdd.n1186 gnd 0.007945f
C2463 vdd.n1187 gnd 0.009871f
C2464 vdd.n1188 gnd 0.009871f
C2465 vdd.n1189 gnd 0.009871f
C2466 vdd.n1190 gnd 0.007945f
C2467 vdd.n1191 gnd 0.007945f
C2468 vdd.n1192 gnd 0.007945f
C2469 vdd.n1193 gnd 0.009871f
C2470 vdd.n1194 gnd 0.009871f
C2471 vdd.n1195 gnd 0.009871f
C2472 vdd.n1196 gnd 0.007945f
C2473 vdd.n1197 gnd 0.007945f
C2474 vdd.n1198 gnd 0.007945f
C2475 vdd.n1199 gnd 0.009871f
C2476 vdd.n1200 gnd 0.009871f
C2477 vdd.n1201 gnd 0.009871f
C2478 vdd.n1202 gnd 0.007945f
C2479 vdd.n1203 gnd 0.007945f
C2480 vdd.n1204 gnd 0.007945f
C2481 vdd.n1205 gnd 0.009871f
C2482 vdd.n1206 gnd 0.009871f
C2483 vdd.n1207 gnd 0.009871f
C2484 vdd.n1208 gnd 0.007945f
C2485 vdd.n1209 gnd 0.007945f
C2486 vdd.n1210 gnd 0.006594f
C2487 vdd.n1211 gnd 0.023626f
C2488 vdd.n1212 gnd 0.023262f
C2489 vdd.n1213 gnd 0.006594f
C2490 vdd.n1214 gnd 0.023262f
C2491 vdd.n1215 gnd 1.4224f
C2492 vdd.n1216 gnd 0.023262f
C2493 vdd.n1217 gnd 0.006594f
C2494 vdd.n1218 gnd 0.023262f
C2495 vdd.n1219 gnd 0.009871f
C2496 vdd.n1220 gnd 0.009871f
C2497 vdd.n1221 gnd 0.007945f
C2498 vdd.n1222 gnd 0.009871f
C2499 vdd.n1223 gnd 0.943222f
C2500 vdd.n1224 gnd 0.009871f
C2501 vdd.n1225 gnd 0.007945f
C2502 vdd.n1226 gnd 0.009871f
C2503 vdd.n1227 gnd 0.009871f
C2504 vdd.n1228 gnd 0.009871f
C2505 vdd.n1229 gnd 0.007945f
C2506 vdd.n1230 gnd 0.009871f
C2507 vdd.n1231 gnd 0.993661f
C2508 vdd.n1232 gnd 0.009871f
C2509 vdd.n1233 gnd 0.007945f
C2510 vdd.n1234 gnd 0.009871f
C2511 vdd.n1235 gnd 0.009871f
C2512 vdd.n1236 gnd 0.009871f
C2513 vdd.n1237 gnd 0.007945f
C2514 vdd.n1238 gnd 0.009871f
C2515 vdd.t166 gnd 0.504397f
C2516 vdd.n1239 gnd 0.822166f
C2517 vdd.n1240 gnd 0.009871f
C2518 vdd.n1241 gnd 0.007945f
C2519 vdd.n1242 gnd 0.009871f
C2520 vdd.n1243 gnd 0.009871f
C2521 vdd.n1244 gnd 0.009871f
C2522 vdd.n1245 gnd 0.007945f
C2523 vdd.n1246 gnd 0.009871f
C2524 vdd.n1247 gnd 0.650672f
C2525 vdd.n1248 gnd 0.009871f
C2526 vdd.n1249 gnd 0.007945f
C2527 vdd.n1250 gnd 0.009871f
C2528 vdd.n1251 gnd 0.009871f
C2529 vdd.n1252 gnd 0.009871f
C2530 vdd.n1253 gnd 0.007945f
C2531 vdd.n1254 gnd 0.009871f
C2532 vdd.n1255 gnd 0.812078f
C2533 vdd.n1256 gnd 0.529616f
C2534 vdd.n1257 gnd 0.009871f
C2535 vdd.n1258 gnd 0.007945f
C2536 vdd.n1259 gnd 0.009871f
C2537 vdd.n1260 gnd 0.009871f
C2538 vdd.n1261 gnd 0.009871f
C2539 vdd.n1262 gnd 0.007945f
C2540 vdd.n1263 gnd 0.009871f
C2541 vdd.n1264 gnd 0.701111f
C2542 vdd.n1265 gnd 0.009871f
C2543 vdd.n1266 gnd 0.007945f
C2544 vdd.n1267 gnd 0.009871f
C2545 vdd.n1268 gnd 0.009871f
C2546 vdd.n1269 gnd 0.009871f
C2547 vdd.n1270 gnd 0.007945f
C2548 vdd.n1271 gnd 0.009871f
C2549 vdd.t2 gnd 0.504397f
C2550 vdd.n1272 gnd 0.837298f
C2551 vdd.n1273 gnd 0.009871f
C2552 vdd.n1274 gnd 0.007945f
C2553 vdd.n1275 gnd 0.005417f
C2554 vdd.n1276 gnd 0.005027f
C2555 vdd.n1277 gnd 0.002781f
C2556 vdd.n1278 gnd 0.006385f
C2557 vdd.n1279 gnd 0.002701f
C2558 vdd.n1280 gnd 0.00286f
C2559 vdd.n1281 gnd 0.005027f
C2560 vdd.n1282 gnd 0.002701f
C2561 vdd.n1283 gnd 0.006385f
C2562 vdd.n1284 gnd 0.00286f
C2563 vdd.n1285 gnd 0.005027f
C2564 vdd.n1286 gnd 0.002701f
C2565 vdd.n1287 gnd 0.004789f
C2566 vdd.n1288 gnd 0.004803f
C2567 vdd.t84 gnd 0.013718f
C2568 vdd.n1289 gnd 0.030521f
C2569 vdd.n1290 gnd 0.158841f
C2570 vdd.n1291 gnd 0.002701f
C2571 vdd.n1292 gnd 0.00286f
C2572 vdd.n1293 gnd 0.006385f
C2573 vdd.n1294 gnd 0.006385f
C2574 vdd.n1295 gnd 0.00286f
C2575 vdd.n1296 gnd 0.002701f
C2576 vdd.n1297 gnd 0.005027f
C2577 vdd.n1298 gnd 0.005027f
C2578 vdd.n1299 gnd 0.002701f
C2579 vdd.n1300 gnd 0.00286f
C2580 vdd.n1301 gnd 0.006385f
C2581 vdd.n1302 gnd 0.006385f
C2582 vdd.n1303 gnd 0.00286f
C2583 vdd.n1304 gnd 0.002701f
C2584 vdd.n1305 gnd 0.005027f
C2585 vdd.n1306 gnd 0.005027f
C2586 vdd.n1307 gnd 0.002701f
C2587 vdd.n1308 gnd 0.00286f
C2588 vdd.n1309 gnd 0.006385f
C2589 vdd.n1310 gnd 0.006385f
C2590 vdd.n1311 gnd 0.015096f
C2591 vdd.n1312 gnd 0.002781f
C2592 vdd.n1313 gnd 0.002701f
C2593 vdd.n1314 gnd 0.012993f
C2594 vdd.n1315 gnd 0.009071f
C2595 vdd.t228 gnd 0.031781f
C2596 vdd.t227 gnd 0.031781f
C2597 vdd.n1316 gnd 0.218418f
C2598 vdd.n1317 gnd 0.171752f
C2599 vdd.t193 gnd 0.031781f
C2600 vdd.t30 gnd 0.031781f
C2601 vdd.n1318 gnd 0.218418f
C2602 vdd.n1319 gnd 0.138603f
C2603 vdd.t197 gnd 0.031781f
C2604 vdd.t31 gnd 0.031781f
C2605 vdd.n1320 gnd 0.218418f
C2606 vdd.n1321 gnd 0.138603f
C2607 vdd.t67 gnd 0.031781f
C2608 vdd.t70 gnd 0.031781f
C2609 vdd.n1322 gnd 0.218418f
C2610 vdd.n1323 gnd 0.138603f
C2611 vdd.t167 gnd 0.031781f
C2612 vdd.t185 gnd 0.031781f
C2613 vdd.n1324 gnd 0.218418f
C2614 vdd.n1325 gnd 0.138603f
C2615 vdd.n1326 gnd 0.005417f
C2616 vdd.n1327 gnd 0.005027f
C2617 vdd.n1328 gnd 0.002781f
C2618 vdd.n1329 gnd 0.006385f
C2619 vdd.n1330 gnd 0.002701f
C2620 vdd.n1331 gnd 0.00286f
C2621 vdd.n1332 gnd 0.005027f
C2622 vdd.n1333 gnd 0.002701f
C2623 vdd.n1334 gnd 0.006385f
C2624 vdd.n1335 gnd 0.00286f
C2625 vdd.n1336 gnd 0.005027f
C2626 vdd.n1337 gnd 0.002701f
C2627 vdd.n1338 gnd 0.004789f
C2628 vdd.n1339 gnd 0.004803f
C2629 vdd.t231 gnd 0.013718f
C2630 vdd.n1340 gnd 0.030521f
C2631 vdd.n1341 gnd 0.158841f
C2632 vdd.n1342 gnd 0.002701f
C2633 vdd.n1343 gnd 0.00286f
C2634 vdd.n1344 gnd 0.006385f
C2635 vdd.n1345 gnd 0.006385f
C2636 vdd.n1346 gnd 0.00286f
C2637 vdd.n1347 gnd 0.002701f
C2638 vdd.n1348 gnd 0.005027f
C2639 vdd.n1349 gnd 0.005027f
C2640 vdd.n1350 gnd 0.002701f
C2641 vdd.n1351 gnd 0.00286f
C2642 vdd.n1352 gnd 0.006385f
C2643 vdd.n1353 gnd 0.006385f
C2644 vdd.n1354 gnd 0.00286f
C2645 vdd.n1355 gnd 0.002701f
C2646 vdd.n1356 gnd 0.005027f
C2647 vdd.n1357 gnd 0.005027f
C2648 vdd.n1358 gnd 0.002701f
C2649 vdd.n1359 gnd 0.00286f
C2650 vdd.n1360 gnd 0.006385f
C2651 vdd.n1361 gnd 0.006385f
C2652 vdd.n1362 gnd 0.015096f
C2653 vdd.n1363 gnd 0.002781f
C2654 vdd.n1364 gnd 0.002701f
C2655 vdd.n1365 gnd 0.012993f
C2656 vdd.n1366 gnd 0.008787f
C2657 vdd.n1367 gnd 0.103122f
C2658 vdd.n1368 gnd 0.005417f
C2659 vdd.n1369 gnd 0.005027f
C2660 vdd.n1370 gnd 0.002781f
C2661 vdd.n1371 gnd 0.006385f
C2662 vdd.n1372 gnd 0.002701f
C2663 vdd.n1373 gnd 0.00286f
C2664 vdd.n1374 gnd 0.005027f
C2665 vdd.n1375 gnd 0.002701f
C2666 vdd.n1376 gnd 0.006385f
C2667 vdd.n1377 gnd 0.00286f
C2668 vdd.n1378 gnd 0.005027f
C2669 vdd.n1379 gnd 0.002701f
C2670 vdd.n1380 gnd 0.004789f
C2671 vdd.n1381 gnd 0.004803f
C2672 vdd.t219 gnd 0.013718f
C2673 vdd.n1382 gnd 0.030521f
C2674 vdd.n1383 gnd 0.158841f
C2675 vdd.n1384 gnd 0.002701f
C2676 vdd.n1385 gnd 0.00286f
C2677 vdd.n1386 gnd 0.006385f
C2678 vdd.n1387 gnd 0.006385f
C2679 vdd.n1388 gnd 0.00286f
C2680 vdd.n1389 gnd 0.002701f
C2681 vdd.n1390 gnd 0.005027f
C2682 vdd.n1391 gnd 0.005027f
C2683 vdd.n1392 gnd 0.002701f
C2684 vdd.n1393 gnd 0.00286f
C2685 vdd.n1394 gnd 0.006385f
C2686 vdd.n1395 gnd 0.006385f
C2687 vdd.n1396 gnd 0.00286f
C2688 vdd.n1397 gnd 0.002701f
C2689 vdd.n1398 gnd 0.005027f
C2690 vdd.n1399 gnd 0.005027f
C2691 vdd.n1400 gnd 0.002701f
C2692 vdd.n1401 gnd 0.00286f
C2693 vdd.n1402 gnd 0.006385f
C2694 vdd.n1403 gnd 0.006385f
C2695 vdd.n1404 gnd 0.015096f
C2696 vdd.n1405 gnd 0.002781f
C2697 vdd.n1406 gnd 0.002701f
C2698 vdd.n1407 gnd 0.012993f
C2699 vdd.n1408 gnd 0.009071f
C2700 vdd.t7 gnd 0.031781f
C2701 vdd.t36 gnd 0.031781f
C2702 vdd.n1409 gnd 0.218418f
C2703 vdd.n1410 gnd 0.171752f
C2704 vdd.t33 gnd 0.031781f
C2705 vdd.t170 gnd 0.031781f
C2706 vdd.n1411 gnd 0.218418f
C2707 vdd.n1412 gnd 0.138603f
C2708 vdd.t27 gnd 0.031781f
C2709 vdd.t3 gnd 0.031781f
C2710 vdd.n1413 gnd 0.218418f
C2711 vdd.n1414 gnd 0.138603f
C2712 vdd.t223 gnd 0.031781f
C2713 vdd.t171 gnd 0.031781f
C2714 vdd.n1415 gnd 0.218418f
C2715 vdd.n1416 gnd 0.138603f
C2716 vdd.t202 gnd 0.031781f
C2717 vdd.t56 gnd 0.031781f
C2718 vdd.n1417 gnd 0.218418f
C2719 vdd.n1418 gnd 0.138603f
C2720 vdd.n1419 gnd 0.005417f
C2721 vdd.n1420 gnd 0.005027f
C2722 vdd.n1421 gnd 0.002781f
C2723 vdd.n1422 gnd 0.006385f
C2724 vdd.n1423 gnd 0.002701f
C2725 vdd.n1424 gnd 0.00286f
C2726 vdd.n1425 gnd 0.005027f
C2727 vdd.n1426 gnd 0.002701f
C2728 vdd.n1427 gnd 0.006385f
C2729 vdd.n1428 gnd 0.00286f
C2730 vdd.n1429 gnd 0.005027f
C2731 vdd.n1430 gnd 0.002701f
C2732 vdd.n1431 gnd 0.004789f
C2733 vdd.n1432 gnd 0.004803f
C2734 vdd.t201 gnd 0.013718f
C2735 vdd.n1433 gnd 0.030521f
C2736 vdd.n1434 gnd 0.158841f
C2737 vdd.n1435 gnd 0.002701f
C2738 vdd.n1436 gnd 0.00286f
C2739 vdd.n1437 gnd 0.006385f
C2740 vdd.n1438 gnd 0.006385f
C2741 vdd.n1439 gnd 0.00286f
C2742 vdd.n1440 gnd 0.002701f
C2743 vdd.n1441 gnd 0.005027f
C2744 vdd.n1442 gnd 0.005027f
C2745 vdd.n1443 gnd 0.002701f
C2746 vdd.n1444 gnd 0.00286f
C2747 vdd.n1445 gnd 0.006385f
C2748 vdd.n1446 gnd 0.006385f
C2749 vdd.n1447 gnd 0.00286f
C2750 vdd.n1448 gnd 0.002701f
C2751 vdd.n1449 gnd 0.005027f
C2752 vdd.n1450 gnd 0.005027f
C2753 vdd.n1451 gnd 0.002701f
C2754 vdd.n1452 gnd 0.00286f
C2755 vdd.n1453 gnd 0.006385f
C2756 vdd.n1454 gnd 0.006385f
C2757 vdd.n1455 gnd 0.015096f
C2758 vdd.n1456 gnd 0.002781f
C2759 vdd.n1457 gnd 0.002701f
C2760 vdd.n1458 gnd 0.012993f
C2761 vdd.n1459 gnd 0.008787f
C2762 vdd.n1460 gnd 0.061347f
C2763 vdd.n1461 gnd 0.221049f
C2764 vdd.n1462 gnd 0.005417f
C2765 vdd.n1463 gnd 0.005027f
C2766 vdd.n1464 gnd 0.002781f
C2767 vdd.n1465 gnd 0.006385f
C2768 vdd.n1466 gnd 0.002701f
C2769 vdd.n1467 gnd 0.00286f
C2770 vdd.n1468 gnd 0.005027f
C2771 vdd.n1469 gnd 0.002701f
C2772 vdd.n1470 gnd 0.006385f
C2773 vdd.n1471 gnd 0.00286f
C2774 vdd.n1472 gnd 0.005027f
C2775 vdd.n1473 gnd 0.002701f
C2776 vdd.n1474 gnd 0.004789f
C2777 vdd.n1475 gnd 0.004803f
C2778 vdd.t9 gnd 0.013718f
C2779 vdd.n1476 gnd 0.030521f
C2780 vdd.n1477 gnd 0.158841f
C2781 vdd.n1478 gnd 0.002701f
C2782 vdd.n1479 gnd 0.00286f
C2783 vdd.n1480 gnd 0.006385f
C2784 vdd.n1481 gnd 0.006385f
C2785 vdd.n1482 gnd 0.00286f
C2786 vdd.n1483 gnd 0.002701f
C2787 vdd.n1484 gnd 0.005027f
C2788 vdd.n1485 gnd 0.005027f
C2789 vdd.n1486 gnd 0.002701f
C2790 vdd.n1487 gnd 0.00286f
C2791 vdd.n1488 gnd 0.006385f
C2792 vdd.n1489 gnd 0.006385f
C2793 vdd.n1490 gnd 0.00286f
C2794 vdd.n1491 gnd 0.002701f
C2795 vdd.n1492 gnd 0.005027f
C2796 vdd.n1493 gnd 0.005027f
C2797 vdd.n1494 gnd 0.002701f
C2798 vdd.n1495 gnd 0.00286f
C2799 vdd.n1496 gnd 0.006385f
C2800 vdd.n1497 gnd 0.006385f
C2801 vdd.n1498 gnd 0.015096f
C2802 vdd.n1499 gnd 0.002781f
C2803 vdd.n1500 gnd 0.002701f
C2804 vdd.n1501 gnd 0.012993f
C2805 vdd.n1502 gnd 0.009071f
C2806 vdd.t194 gnd 0.031781f
C2807 vdd.t11 gnd 0.031781f
C2808 vdd.n1503 gnd 0.218418f
C2809 vdd.n1504 gnd 0.171752f
C2810 vdd.t222 gnd 0.031781f
C2811 vdd.t216 gnd 0.031781f
C2812 vdd.n1505 gnd 0.218418f
C2813 vdd.n1506 gnd 0.138603f
C2814 vdd.t199 gnd 0.031781f
C2815 vdd.t23 gnd 0.031781f
C2816 vdd.n1507 gnd 0.218418f
C2817 vdd.n1508 gnd 0.138603f
C2818 vdd.t173 gnd 0.031781f
C2819 vdd.t217 gnd 0.031781f
C2820 vdd.n1509 gnd 0.218418f
C2821 vdd.n1510 gnd 0.138603f
C2822 vdd.t188 gnd 0.031781f
C2823 vdd.t196 gnd 0.031781f
C2824 vdd.n1511 gnd 0.218418f
C2825 vdd.n1512 gnd 0.138603f
C2826 vdd.n1513 gnd 0.005417f
C2827 vdd.n1514 gnd 0.005027f
C2828 vdd.n1515 gnd 0.002781f
C2829 vdd.n1516 gnd 0.006385f
C2830 vdd.n1517 gnd 0.002701f
C2831 vdd.n1518 gnd 0.00286f
C2832 vdd.n1519 gnd 0.005027f
C2833 vdd.n1520 gnd 0.002701f
C2834 vdd.n1521 gnd 0.006385f
C2835 vdd.n1522 gnd 0.00286f
C2836 vdd.n1523 gnd 0.005027f
C2837 vdd.n1524 gnd 0.002701f
C2838 vdd.n1525 gnd 0.004789f
C2839 vdd.n1526 gnd 0.004803f
C2840 vdd.t187 gnd 0.013718f
C2841 vdd.n1527 gnd 0.030521f
C2842 vdd.n1528 gnd 0.158841f
C2843 vdd.n1529 gnd 0.002701f
C2844 vdd.n1530 gnd 0.00286f
C2845 vdd.n1531 gnd 0.006385f
C2846 vdd.n1532 gnd 0.006385f
C2847 vdd.n1533 gnd 0.00286f
C2848 vdd.n1534 gnd 0.002701f
C2849 vdd.n1535 gnd 0.005027f
C2850 vdd.n1536 gnd 0.005027f
C2851 vdd.n1537 gnd 0.002701f
C2852 vdd.n1538 gnd 0.00286f
C2853 vdd.n1539 gnd 0.006385f
C2854 vdd.n1540 gnd 0.006385f
C2855 vdd.n1541 gnd 0.00286f
C2856 vdd.n1542 gnd 0.002701f
C2857 vdd.n1543 gnd 0.005027f
C2858 vdd.n1544 gnd 0.005027f
C2859 vdd.n1545 gnd 0.002701f
C2860 vdd.n1546 gnd 0.00286f
C2861 vdd.n1547 gnd 0.006385f
C2862 vdd.n1548 gnd 0.006385f
C2863 vdd.n1549 gnd 0.015096f
C2864 vdd.n1550 gnd 0.002781f
C2865 vdd.n1551 gnd 0.002701f
C2866 vdd.n1552 gnd 0.012993f
C2867 vdd.n1553 gnd 0.008787f
C2868 vdd.n1554 gnd 0.061347f
C2869 vdd.n1555 gnd 0.24294f
C2870 vdd.n1556 gnd 2.1865f
C2871 vdd.n1557 gnd 0.587613f
C2872 vdd.n1558 gnd 0.009837f
C2873 vdd.n1559 gnd 0.009871f
C2874 vdd.n1560 gnd 0.007945f
C2875 vdd.n1561 gnd 0.009871f
C2876 vdd.n1562 gnd 0.801991f
C2877 vdd.n1563 gnd 0.009871f
C2878 vdd.n1564 gnd 0.007945f
C2879 vdd.n1565 gnd 0.009871f
C2880 vdd.n1566 gnd 0.009871f
C2881 vdd.n1567 gnd 0.009871f
C2882 vdd.n1568 gnd 0.007945f
C2883 vdd.n1569 gnd 0.009871f
C2884 vdd.n1570 gnd 0.837298f
C2885 vdd.t29 gnd 0.504397f
C2886 vdd.n1571 gnd 0.630496f
C2887 vdd.n1572 gnd 0.009871f
C2888 vdd.n1573 gnd 0.007945f
C2889 vdd.n1574 gnd 0.009871f
C2890 vdd.n1575 gnd 0.009871f
C2891 vdd.n1576 gnd 0.009871f
C2892 vdd.n1577 gnd 0.007945f
C2893 vdd.n1578 gnd 0.009871f
C2894 vdd.n1579 gnd 0.549792f
C2895 vdd.n1580 gnd 0.009871f
C2896 vdd.n1581 gnd 0.007945f
C2897 vdd.n1582 gnd 0.009871f
C2898 vdd.n1583 gnd 0.009871f
C2899 vdd.n1584 gnd 0.009871f
C2900 vdd.n1585 gnd 0.007945f
C2901 vdd.n1586 gnd 0.009871f
C2902 vdd.n1587 gnd 0.620408f
C2903 vdd.n1588 gnd 0.721287f
C2904 vdd.n1589 gnd 0.009871f
C2905 vdd.n1590 gnd 0.007945f
C2906 vdd.n1591 gnd 0.009871f
C2907 vdd.n1592 gnd 0.009871f
C2908 vdd.n1593 gnd 0.009871f
C2909 vdd.n1594 gnd 0.007945f
C2910 vdd.n1595 gnd 0.009871f
C2911 vdd.n1596 gnd 0.892782f
C2912 vdd.n1597 gnd 0.009871f
C2913 vdd.n1598 gnd 0.007945f
C2914 vdd.n1599 gnd 0.009871f
C2915 vdd.n1600 gnd 0.009871f
C2916 vdd.n1601 gnd 0.023262f
C2917 vdd.n1602 gnd 0.009871f
C2918 vdd.n1603 gnd 0.009871f
C2919 vdd.n1604 gnd 0.007945f
C2920 vdd.n1605 gnd 0.009871f
C2921 vdd.n1606 gnd 0.539704f
C2922 vdd.n1607 gnd 1.00879f
C2923 vdd.n1608 gnd 0.009871f
C2924 vdd.n1609 gnd 0.007945f
C2925 vdd.n1610 gnd 0.009871f
C2926 vdd.n1611 gnd 0.009871f
C2927 vdd.n1612 gnd 0.008489f
C2928 vdd.n1613 gnd 0.007945f
C2929 vdd.n1615 gnd 0.009871f
C2930 vdd.n1617 gnd 0.007945f
C2931 vdd.n1618 gnd 0.009871f
C2932 vdd.n1619 gnd 0.007945f
C2933 vdd.n1621 gnd 0.009871f
C2934 vdd.n1622 gnd 0.007945f
C2935 vdd.n1623 gnd 0.009871f
C2936 vdd.n1624 gnd 0.009871f
C2937 vdd.n1625 gnd 0.009871f
C2938 vdd.n1626 gnd 0.009871f
C2939 vdd.n1627 gnd 0.009871f
C2940 vdd.n1628 gnd 0.007945f
C2941 vdd.n1630 gnd 0.009871f
C2942 vdd.n1631 gnd 0.009871f
C2943 vdd.n1632 gnd 0.009871f
C2944 vdd.n1633 gnd 0.009871f
C2945 vdd.n1634 gnd 0.009871f
C2946 vdd.n1635 gnd 0.007945f
C2947 vdd.n1637 gnd 0.009871f
C2948 vdd.n1638 gnd 0.009871f
C2949 vdd.n1639 gnd 0.009871f
C2950 vdd.n1640 gnd 0.009871f
C2951 vdd.n1641 gnd 0.006634f
C2952 vdd.t113 gnd 0.121442f
C2953 vdd.t112 gnd 0.129788f
C2954 vdd.t111 gnd 0.158602f
C2955 vdd.n1642 gnd 0.203305f
C2956 vdd.n1643 gnd 0.170813f
C2957 vdd.n1645 gnd 0.009871f
C2958 vdd.n1646 gnd 0.009871f
C2959 vdd.n1647 gnd 0.007945f
C2960 vdd.n1648 gnd 0.009871f
C2961 vdd.n1650 gnd 0.009871f
C2962 vdd.n1651 gnd 0.009871f
C2963 vdd.n1652 gnd 0.009871f
C2964 vdd.n1653 gnd 0.009871f
C2965 vdd.n1654 gnd 0.007945f
C2966 vdd.n1656 gnd 0.009871f
C2967 vdd.n1657 gnd 0.009871f
C2968 vdd.n1658 gnd 0.009871f
C2969 vdd.n1659 gnd 0.009871f
C2970 vdd.n1660 gnd 0.009871f
C2971 vdd.n1661 gnd 0.007945f
C2972 vdd.n1663 gnd 0.009871f
C2973 vdd.n1664 gnd 0.009871f
C2974 vdd.n1665 gnd 0.009871f
C2975 vdd.n1666 gnd 0.009871f
C2976 vdd.n1667 gnd 0.009871f
C2977 vdd.n1668 gnd 0.007945f
C2978 vdd.n1670 gnd 0.009871f
C2979 vdd.n1671 gnd 0.009871f
C2980 vdd.n1672 gnd 0.009871f
C2981 vdd.n1673 gnd 0.009871f
C2982 vdd.n1674 gnd 0.009871f
C2983 vdd.n1675 gnd 0.007945f
C2984 vdd.n1677 gnd 0.009871f
C2985 vdd.n1678 gnd 0.009871f
C2986 vdd.n1679 gnd 0.009871f
C2987 vdd.n1680 gnd 0.009871f
C2988 vdd.n1681 gnd 0.007866f
C2989 vdd.t107 gnd 0.121442f
C2990 vdd.t106 gnd 0.129788f
C2991 vdd.t105 gnd 0.158602f
C2992 vdd.n1682 gnd 0.203305f
C2993 vdd.n1683 gnd 0.170813f
C2994 vdd.n1685 gnd 0.009871f
C2995 vdd.n1686 gnd 0.009871f
C2996 vdd.n1687 gnd 0.007945f
C2997 vdd.n1688 gnd 0.009871f
C2998 vdd.n1690 gnd 0.009871f
C2999 vdd.n1691 gnd 0.009871f
C3000 vdd.n1692 gnd 0.009871f
C3001 vdd.n1693 gnd 0.009871f
C3002 vdd.n1694 gnd 0.007945f
C3003 vdd.n1696 gnd 0.009871f
C3004 vdd.n1697 gnd 0.009871f
C3005 vdd.n1698 gnd 0.009871f
C3006 vdd.n1699 gnd 0.009871f
C3007 vdd.n1700 gnd 0.009871f
C3008 vdd.n1701 gnd 0.007945f
C3009 vdd.n1703 gnd 0.009871f
C3010 vdd.n1704 gnd 0.009871f
C3011 vdd.n1705 gnd 0.009871f
C3012 vdd.n1706 gnd 0.009871f
C3013 vdd.n1707 gnd 0.009871f
C3014 vdd.n1708 gnd 0.009871f
C3015 vdd.n1709 gnd 0.007945f
C3016 vdd.n1711 gnd 0.009871f
C3017 vdd.n1713 gnd 0.009871f
C3018 vdd.n1714 gnd 0.007945f
C3019 vdd.n1715 gnd 0.007945f
C3020 vdd.n1716 gnd 0.009871f
C3021 vdd.n1718 gnd 0.009871f
C3022 vdd.n1719 gnd 0.007945f
C3023 vdd.n1720 gnd 0.007945f
C3024 vdd.n1721 gnd 0.009871f
C3025 vdd.n1723 gnd 0.009871f
C3026 vdd.n1724 gnd 0.009871f
C3027 vdd.n1725 gnd 0.007945f
C3028 vdd.n1726 gnd 0.007945f
C3029 vdd.n1727 gnd 0.007945f
C3030 vdd.n1728 gnd 0.009871f
C3031 vdd.n1730 gnd 0.009871f
C3032 vdd.n1731 gnd 0.009871f
C3033 vdd.n1732 gnd 0.007945f
C3034 vdd.n1733 gnd 0.007945f
C3035 vdd.n1734 gnd 0.007945f
C3036 vdd.n1735 gnd 0.009871f
C3037 vdd.n1737 gnd 0.009871f
C3038 vdd.n1738 gnd 0.009871f
C3039 vdd.n1739 gnd 0.007945f
C3040 vdd.n1740 gnd 0.007945f
C3041 vdd.n1741 gnd 0.007945f
C3042 vdd.n1742 gnd 0.009871f
C3043 vdd.n1744 gnd 0.009871f
C3044 vdd.n1745 gnd 0.009871f
C3045 vdd.n1746 gnd 0.007945f
C3046 vdd.n1747 gnd 0.009871f
C3047 vdd.n1748 gnd 0.009871f
C3048 vdd.n1749 gnd 0.009871f
C3049 vdd.n1750 gnd 0.016208f
C3050 vdd.n1751 gnd 0.005403f
C3051 vdd.n1752 gnd 0.007945f
C3052 vdd.n1753 gnd 0.009871f
C3053 vdd.n1755 gnd 0.009871f
C3054 vdd.n1756 gnd 0.009871f
C3055 vdd.n1757 gnd 0.007945f
C3056 vdd.n1758 gnd 0.007945f
C3057 vdd.n1759 gnd 0.007945f
C3058 vdd.n1760 gnd 0.009871f
C3059 vdd.n1762 gnd 0.009871f
C3060 vdd.n1763 gnd 0.009871f
C3061 vdd.n1764 gnd 0.007945f
C3062 vdd.n1765 gnd 0.007945f
C3063 vdd.n1766 gnd 0.007945f
C3064 vdd.n1767 gnd 0.009871f
C3065 vdd.n1769 gnd 0.009871f
C3066 vdd.n1770 gnd 0.009871f
C3067 vdd.n1771 gnd 0.007945f
C3068 vdd.n1772 gnd 0.007945f
C3069 vdd.n1773 gnd 0.007945f
C3070 vdd.n1774 gnd 0.009871f
C3071 vdd.n1776 gnd 0.009871f
C3072 vdd.n1777 gnd 0.009871f
C3073 vdd.n1778 gnd 0.007945f
C3074 vdd.n1779 gnd 0.007945f
C3075 vdd.n1780 gnd 0.007945f
C3076 vdd.n1781 gnd 0.009871f
C3077 vdd.n1783 gnd 0.009871f
C3078 vdd.n1784 gnd 0.009871f
C3079 vdd.n1785 gnd 0.007945f
C3080 vdd.n1786 gnd 0.009871f
C3081 vdd.n1787 gnd 0.009871f
C3082 vdd.n1788 gnd 0.009871f
C3083 vdd.n1789 gnd 0.016208f
C3084 vdd.n1790 gnd 0.006634f
C3085 vdd.n1791 gnd 0.007945f
C3086 vdd.n1792 gnd 0.009871f
C3087 vdd.n1794 gnd 0.009871f
C3088 vdd.n1795 gnd 0.009871f
C3089 vdd.n1796 gnd 0.007945f
C3090 vdd.n1797 gnd 0.007945f
C3091 vdd.n1798 gnd 0.007945f
C3092 vdd.n1799 gnd 0.009871f
C3093 vdd.n1801 gnd 0.009871f
C3094 vdd.n1802 gnd 0.009871f
C3095 vdd.n1803 gnd 0.007945f
C3096 vdd.n1804 gnd 0.007945f
C3097 vdd.n1805 gnd 0.007945f
C3098 vdd.n1806 gnd 0.009871f
C3099 vdd.n1808 gnd 0.009871f
C3100 vdd.n1809 gnd 0.009871f
C3101 vdd.n1811 gnd 0.009871f
C3102 vdd.n1812 gnd 0.007945f
C3103 vdd.n1813 gnd 0.006318f
C3104 vdd.n1814 gnd 0.006712f
C3105 vdd.n1815 gnd 0.006712f
C3106 vdd.n1816 gnd 0.006712f
C3107 vdd.n1817 gnd 0.006712f
C3108 vdd.n1818 gnd 0.006712f
C3109 vdd.n1819 gnd 0.006712f
C3110 vdd.n1820 gnd 0.006712f
C3111 vdd.n1821 gnd 0.006712f
C3112 vdd.n1823 gnd 0.006712f
C3113 vdd.n1824 gnd 0.006712f
C3114 vdd.n1825 gnd 0.006712f
C3115 vdd.n1826 gnd 0.006712f
C3116 vdd.n1827 gnd 0.006712f
C3117 vdd.n1829 gnd 0.006712f
C3118 vdd.n1831 gnd 0.006712f
C3119 vdd.n1832 gnd 0.006712f
C3120 vdd.n1833 gnd 0.006712f
C3121 vdd.n1834 gnd 0.006712f
C3122 vdd.n1835 gnd 0.006712f
C3123 vdd.n1837 gnd 0.006712f
C3124 vdd.n1839 gnd 0.006712f
C3125 vdd.n1840 gnd 0.006712f
C3126 vdd.n1841 gnd 0.006712f
C3127 vdd.n1842 gnd 0.006712f
C3128 vdd.n1843 gnd 0.006712f
C3129 vdd.n1845 gnd 0.006712f
C3130 vdd.n1847 gnd 0.006712f
C3131 vdd.n1848 gnd 0.006712f
C3132 vdd.n1849 gnd 0.006712f
C3133 vdd.n1850 gnd 0.006712f
C3134 vdd.n1851 gnd 0.006712f
C3135 vdd.n1853 gnd 0.006712f
C3136 vdd.n1854 gnd 0.006712f
C3137 vdd.n1855 gnd 0.006712f
C3138 vdd.n1856 gnd 0.006712f
C3139 vdd.n1857 gnd 0.006712f
C3140 vdd.n1858 gnd 0.006712f
C3141 vdd.n1859 gnd 0.006712f
C3142 vdd.n1860 gnd 0.006712f
C3143 vdd.n1861 gnd 0.004886f
C3144 vdd.n1862 gnd 0.006712f
C3145 vdd.t157 gnd 0.271249f
C3146 vdd.t158 gnd 0.277657f
C3147 vdd.t156 gnd 0.177082f
C3148 vdd.n1863 gnd 0.095703f
C3149 vdd.n1864 gnd 0.054286f
C3150 vdd.n1865 gnd 0.009593f
C3151 vdd.n1866 gnd 0.006712f
C3152 vdd.n1867 gnd 0.006712f
C3153 vdd.n1868 gnd 0.408561f
C3154 vdd.n1869 gnd 0.006712f
C3155 vdd.n1870 gnd 0.006712f
C3156 vdd.n1871 gnd 0.006712f
C3157 vdd.n1872 gnd 0.006712f
C3158 vdd.n1873 gnd 0.006712f
C3159 vdd.n1874 gnd 0.006712f
C3160 vdd.n1875 gnd 0.006712f
C3161 vdd.n1876 gnd 0.006712f
C3162 vdd.n1877 gnd 0.006712f
C3163 vdd.n1878 gnd 0.006712f
C3164 vdd.n1879 gnd 0.006712f
C3165 vdd.n1880 gnd 0.006712f
C3166 vdd.n1881 gnd 0.006712f
C3167 vdd.n1882 gnd 0.006712f
C3168 vdd.n1883 gnd 0.006712f
C3169 vdd.n1884 gnd 0.006712f
C3170 vdd.n1885 gnd 0.006712f
C3171 vdd.n1886 gnd 0.006712f
C3172 vdd.n1887 gnd 0.006712f
C3173 vdd.n1888 gnd 0.006712f
C3174 vdd.t131 gnd 0.271249f
C3175 vdd.t132 gnd 0.277657f
C3176 vdd.t129 gnd 0.177082f
C3177 vdd.n1889 gnd 0.095703f
C3178 vdd.n1890 gnd 0.054286f
C3179 vdd.n1891 gnd 0.006712f
C3180 vdd.n1892 gnd 0.006712f
C3181 vdd.n1893 gnd 0.006712f
C3182 vdd.n1894 gnd 0.006712f
C3183 vdd.n1895 gnd 0.006712f
C3184 vdd.n1896 gnd 0.006712f
C3185 vdd.n1898 gnd 0.006712f
C3186 vdd.n1899 gnd 0.006712f
C3187 vdd.n1900 gnd 0.006712f
C3188 vdd.n1901 gnd 0.006712f
C3189 vdd.n1903 gnd 0.006712f
C3190 vdd.n1905 gnd 0.006712f
C3191 vdd.n1906 gnd 0.006712f
C3192 vdd.n1907 gnd 0.006712f
C3193 vdd.n1908 gnd 0.006712f
C3194 vdd.n1909 gnd 0.006712f
C3195 vdd.n1911 gnd 0.006712f
C3196 vdd.n1913 gnd 0.006712f
C3197 vdd.n1914 gnd 0.006712f
C3198 vdd.n1915 gnd 0.006712f
C3199 vdd.n1916 gnd 0.006712f
C3200 vdd.n1917 gnd 0.006712f
C3201 vdd.n1919 gnd 0.006712f
C3202 vdd.n1921 gnd 0.006712f
C3203 vdd.n1922 gnd 0.006712f
C3204 vdd.n1923 gnd 0.004886f
C3205 vdd.n1924 gnd 0.009593f
C3206 vdd.n1925 gnd 0.005182f
C3207 vdd.n1926 gnd 0.006712f
C3208 vdd.n1928 gnd 0.006712f
C3209 vdd.n1929 gnd 0.015927f
C3210 vdd.n1930 gnd 0.015927f
C3211 vdd.n1931 gnd 0.014871f
C3212 vdd.n1932 gnd 0.006712f
C3213 vdd.n1933 gnd 0.006712f
C3214 vdd.n1934 gnd 0.006712f
C3215 vdd.n1935 gnd 0.006712f
C3216 vdd.n1936 gnd 0.006712f
C3217 vdd.n1937 gnd 0.006712f
C3218 vdd.n1938 gnd 0.006712f
C3219 vdd.n1939 gnd 0.006712f
C3220 vdd.n1940 gnd 0.006712f
C3221 vdd.n1941 gnd 0.006712f
C3222 vdd.n1942 gnd 0.006712f
C3223 vdd.n1943 gnd 0.006712f
C3224 vdd.n1944 gnd 0.006712f
C3225 vdd.n1945 gnd 0.006712f
C3226 vdd.n1946 gnd 0.006712f
C3227 vdd.n1947 gnd 0.006712f
C3228 vdd.n1948 gnd 0.006712f
C3229 vdd.n1949 gnd 0.006712f
C3230 vdd.n1950 gnd 0.006712f
C3231 vdd.n1951 gnd 0.006712f
C3232 vdd.n1952 gnd 0.006712f
C3233 vdd.n1953 gnd 0.006712f
C3234 vdd.n1954 gnd 0.006712f
C3235 vdd.n1955 gnd 0.006712f
C3236 vdd.n1956 gnd 0.006712f
C3237 vdd.n1957 gnd 0.006712f
C3238 vdd.n1958 gnd 0.006712f
C3239 vdd.n1959 gnd 0.006712f
C3240 vdd.n1960 gnd 0.006712f
C3241 vdd.n1961 gnd 0.006712f
C3242 vdd.n1962 gnd 0.006712f
C3243 vdd.n1963 gnd 0.006712f
C3244 vdd.n1964 gnd 0.006712f
C3245 vdd.n1965 gnd 0.006712f
C3246 vdd.n1966 gnd 0.006712f
C3247 vdd.n1967 gnd 0.006712f
C3248 vdd.n1968 gnd 0.006712f
C3249 vdd.n1969 gnd 0.216891f
C3250 vdd.n1970 gnd 0.006712f
C3251 vdd.n1971 gnd 0.006712f
C3252 vdd.n1972 gnd 0.006712f
C3253 vdd.n1973 gnd 0.006712f
C3254 vdd.n1974 gnd 0.006712f
C3255 vdd.n1975 gnd 0.006712f
C3256 vdd.n1976 gnd 0.006712f
C3257 vdd.n1977 gnd 0.006712f
C3258 vdd.n1978 gnd 0.006712f
C3259 vdd.n1979 gnd 0.006712f
C3260 vdd.n1980 gnd 0.006712f
C3261 vdd.n1981 gnd 0.006712f
C3262 vdd.n1982 gnd 0.006712f
C3263 vdd.n1983 gnd 0.006712f
C3264 vdd.n1984 gnd 0.006712f
C3265 vdd.n1985 gnd 0.006712f
C3266 vdd.n1986 gnd 0.006712f
C3267 vdd.n1987 gnd 0.006712f
C3268 vdd.n1988 gnd 0.006712f
C3269 vdd.n1989 gnd 0.006712f
C3270 vdd.n1990 gnd 0.014871f
C3271 vdd.n1992 gnd 0.015927f
C3272 vdd.n1993 gnd 0.015927f
C3273 vdd.n1994 gnd 0.006712f
C3274 vdd.n1995 gnd 0.005182f
C3275 vdd.n1996 gnd 0.006712f
C3276 vdd.n1998 gnd 0.006712f
C3277 vdd.n2000 gnd 0.006712f
C3278 vdd.n2001 gnd 0.006712f
C3279 vdd.n2002 gnd 0.006712f
C3280 vdd.n2003 gnd 0.006712f
C3281 vdd.n2004 gnd 0.006712f
C3282 vdd.n2006 gnd 0.006712f
C3283 vdd.n2008 gnd 0.006712f
C3284 vdd.n2009 gnd 0.006712f
C3285 vdd.n2010 gnd 0.006712f
C3286 vdd.n2011 gnd 0.006712f
C3287 vdd.n2012 gnd 0.006712f
C3288 vdd.n2014 gnd 0.006712f
C3289 vdd.n2016 gnd 0.006712f
C3290 vdd.n2017 gnd 0.006712f
C3291 vdd.n2018 gnd 0.006712f
C3292 vdd.n2019 gnd 0.006712f
C3293 vdd.n2020 gnd 0.006712f
C3294 vdd.n2022 gnd 0.006712f
C3295 vdd.n2024 gnd 0.006712f
C3296 vdd.n2025 gnd 0.006712f
C3297 vdd.n2026 gnd 0.020022f
C3298 vdd.n2027 gnd 0.593532f
C3299 vdd.n2029 gnd 0.007945f
C3300 vdd.n2030 gnd 0.007945f
C3301 vdd.n2031 gnd 0.009871f
C3302 vdd.n2033 gnd 0.009871f
C3303 vdd.n2034 gnd 0.009871f
C3304 vdd.n2035 gnd 0.007945f
C3305 vdd.n2036 gnd 0.006594f
C3306 vdd.n2037 gnd 0.023626f
C3307 vdd.n2038 gnd 0.023262f
C3308 vdd.n2039 gnd 0.006594f
C3309 vdd.n2040 gnd 0.023262f
C3310 vdd.n2041 gnd 1.38709f
C3311 vdd.n2042 gnd 0.023262f
C3312 vdd.n2043 gnd 0.023626f
C3313 vdd.n2044 gnd 0.003774f
C3314 vdd.t96 gnd 0.121442f
C3315 vdd.t95 gnd 0.129788f
C3316 vdd.t93 gnd 0.158602f
C3317 vdd.n2045 gnd 0.203305f
C3318 vdd.n2046 gnd 0.170813f
C3319 vdd.n2047 gnd 0.012235f
C3320 vdd.n2048 gnd 0.004171f
C3321 vdd.n2049 gnd 0.008489f
C3322 vdd.n2050 gnd 0.593532f
C3323 vdd.n2051 gnd 0.020022f
C3324 vdd.n2052 gnd 0.006712f
C3325 vdd.n2053 gnd 0.006712f
C3326 vdd.n2054 gnd 0.006712f
C3327 vdd.n2056 gnd 0.006712f
C3328 vdd.n2058 gnd 0.006712f
C3329 vdd.n2059 gnd 0.006712f
C3330 vdd.n2060 gnd 0.006712f
C3331 vdd.n2061 gnd 0.006712f
C3332 vdd.n2062 gnd 0.006712f
C3333 vdd.n2064 gnd 0.006712f
C3334 vdd.n2066 gnd 0.006712f
C3335 vdd.n2067 gnd 0.006712f
C3336 vdd.n2068 gnd 0.006712f
C3337 vdd.n2069 gnd 0.006712f
C3338 vdd.n2070 gnd 0.006712f
C3339 vdd.n2072 gnd 0.006712f
C3340 vdd.n2074 gnd 0.006712f
C3341 vdd.n2075 gnd 0.006712f
C3342 vdd.n2076 gnd 0.006712f
C3343 vdd.n2077 gnd 0.006712f
C3344 vdd.n2078 gnd 0.006712f
C3345 vdd.n2080 gnd 0.006712f
C3346 vdd.n2082 gnd 0.006712f
C3347 vdd.n2083 gnd 0.006712f
C3348 vdd.n2084 gnd 0.015927f
C3349 vdd.n2085 gnd 0.014871f
C3350 vdd.n2086 gnd 0.014871f
C3351 vdd.n2087 gnd 0.988617f
C3352 vdd.n2088 gnd 0.014871f
C3353 vdd.n2089 gnd 0.014871f
C3354 vdd.n2090 gnd 0.006712f
C3355 vdd.n2091 gnd 0.006712f
C3356 vdd.n2092 gnd 0.006712f
C3357 vdd.n2093 gnd 0.428737f
C3358 vdd.n2094 gnd 0.006712f
C3359 vdd.n2095 gnd 0.006712f
C3360 vdd.n2096 gnd 0.006712f
C3361 vdd.n2097 gnd 0.006712f
C3362 vdd.n2098 gnd 0.006712f
C3363 vdd.n2099 gnd 0.685979f
C3364 vdd.n2100 gnd 0.006712f
C3365 vdd.n2101 gnd 0.006712f
C3366 vdd.n2102 gnd 0.006712f
C3367 vdd.n2103 gnd 0.006712f
C3368 vdd.n2104 gnd 0.006712f
C3369 vdd.n2105 gnd 0.685979f
C3370 vdd.n2106 gnd 0.006712f
C3371 vdd.n2107 gnd 0.006712f
C3372 vdd.n2108 gnd 0.005923f
C3373 vdd.n2109 gnd 0.019445f
C3374 vdd.n2110 gnd 0.004146f
C3375 vdd.n2111 gnd 0.006712f
C3376 vdd.n2112 gnd 0.378297f
C3377 vdd.n2113 gnd 0.006712f
C3378 vdd.n2114 gnd 0.006712f
C3379 vdd.n2115 gnd 0.006712f
C3380 vdd.n2116 gnd 0.006712f
C3381 vdd.n2117 gnd 0.006712f
C3382 vdd.n2118 gnd 0.459001f
C3383 vdd.n2119 gnd 0.006712f
C3384 vdd.n2120 gnd 0.006712f
C3385 vdd.n2121 gnd 0.006712f
C3386 vdd.n2122 gnd 0.006712f
C3387 vdd.n2123 gnd 0.006712f
C3388 vdd.n2124 gnd 0.61032f
C3389 vdd.n2125 gnd 0.006712f
C3390 vdd.n2126 gnd 0.006712f
C3391 vdd.n2127 gnd 0.006712f
C3392 vdd.n2128 gnd 0.006712f
C3393 vdd.n2129 gnd 0.006712f
C3394 vdd.n2130 gnd 0.544748f
C3395 vdd.n2131 gnd 0.006712f
C3396 vdd.n2132 gnd 0.006712f
C3397 vdd.n2133 gnd 0.006712f
C3398 vdd.n2134 gnd 0.006712f
C3399 vdd.n2135 gnd 0.006712f
C3400 vdd.n2136 gnd 0.393429f
C3401 vdd.n2137 gnd 0.006712f
C3402 vdd.n2138 gnd 0.006712f
C3403 vdd.n2139 gnd 0.006712f
C3404 vdd.n2140 gnd 0.006712f
C3405 vdd.n2141 gnd 0.006712f
C3406 vdd.n2142 gnd 0.216891f
C3407 vdd.n2143 gnd 0.006712f
C3408 vdd.n2144 gnd 0.006712f
C3409 vdd.n2145 gnd 0.006712f
C3410 vdd.n2146 gnd 0.006712f
C3411 vdd.n2147 gnd 0.006712f
C3412 vdd.n2148 gnd 0.378297f
C3413 vdd.n2149 gnd 0.006712f
C3414 vdd.n2150 gnd 0.006712f
C3415 vdd.n2151 gnd 0.006712f
C3416 vdd.n2152 gnd 0.006712f
C3417 vdd.n2153 gnd 0.006712f
C3418 vdd.n2154 gnd 0.685979f
C3419 vdd.n2155 gnd 0.006712f
C3420 vdd.n2156 gnd 0.006712f
C3421 vdd.n2157 gnd 0.006712f
C3422 vdd.n2158 gnd 0.006712f
C3423 vdd.n2159 gnd 0.006712f
C3424 vdd.n2160 gnd 0.006712f
C3425 vdd.n2161 gnd 0.006712f
C3426 vdd.n2162 gnd 0.53466f
C3427 vdd.n2163 gnd 0.006712f
C3428 vdd.n2164 gnd 0.006712f
C3429 vdd.n2165 gnd 0.006712f
C3430 vdd.n2166 gnd 0.006712f
C3431 vdd.n2167 gnd 0.006712f
C3432 vdd.n2168 gnd 0.006712f
C3433 vdd.n2169 gnd 0.428737f
C3434 vdd.n2170 gnd 0.006712f
C3435 vdd.n2171 gnd 0.006712f
C3436 vdd.n2172 gnd 0.006712f
C3437 vdd.n2173 gnd 0.015688f
C3438 vdd.n2174 gnd 0.01511f
C3439 vdd.n2175 gnd 0.006712f
C3440 vdd.n2176 gnd 0.006712f
C3441 vdd.n2177 gnd 0.005182f
C3442 vdd.n2178 gnd 0.006712f
C3443 vdd.n2179 gnd 0.006712f
C3444 vdd.n2180 gnd 0.004886f
C3445 vdd.n2181 gnd 0.006712f
C3446 vdd.n2182 gnd 0.006712f
C3447 vdd.n2183 gnd 0.006712f
C3448 vdd.n2184 gnd 0.006712f
C3449 vdd.n2185 gnd 0.006712f
C3450 vdd.n2186 gnd 0.006712f
C3451 vdd.n2187 gnd 0.006712f
C3452 vdd.n2188 gnd 0.006712f
C3453 vdd.n2189 gnd 0.006712f
C3454 vdd.n2190 gnd 0.006712f
C3455 vdd.n2191 gnd 0.006712f
C3456 vdd.n2192 gnd 0.006712f
C3457 vdd.n2193 gnd 0.006712f
C3458 vdd.n2194 gnd 0.006712f
C3459 vdd.n2195 gnd 0.006712f
C3460 vdd.n2196 gnd 0.006712f
C3461 vdd.n2197 gnd 0.006712f
C3462 vdd.n2198 gnd 0.006712f
C3463 vdd.n2199 gnd 0.006712f
C3464 vdd.n2200 gnd 0.006712f
C3465 vdd.n2201 gnd 0.006712f
C3466 vdd.n2202 gnd 0.006712f
C3467 vdd.n2203 gnd 0.006712f
C3468 vdd.n2204 gnd 0.006712f
C3469 vdd.n2205 gnd 0.006712f
C3470 vdd.n2206 gnd 0.006712f
C3471 vdd.n2207 gnd 0.006712f
C3472 vdd.n2208 gnd 0.006712f
C3473 vdd.n2209 gnd 0.006712f
C3474 vdd.n2210 gnd 0.006712f
C3475 vdd.n2211 gnd 0.006712f
C3476 vdd.n2212 gnd 0.006712f
C3477 vdd.n2213 gnd 0.006712f
C3478 vdd.n2214 gnd 0.006712f
C3479 vdd.n2215 gnd 0.006712f
C3480 vdd.n2216 gnd 0.006712f
C3481 vdd.n2217 gnd 0.006712f
C3482 vdd.n2218 gnd 0.006712f
C3483 vdd.n2219 gnd 0.006712f
C3484 vdd.n2220 gnd 0.006712f
C3485 vdd.n2221 gnd 0.006712f
C3486 vdd.n2222 gnd 0.006712f
C3487 vdd.n2223 gnd 0.006712f
C3488 vdd.n2224 gnd 0.006712f
C3489 vdd.n2225 gnd 0.006712f
C3490 vdd.n2226 gnd 0.006712f
C3491 vdd.n2227 gnd 0.006712f
C3492 vdd.n2228 gnd 0.006712f
C3493 vdd.n2229 gnd 0.006712f
C3494 vdd.n2230 gnd 0.006712f
C3495 vdd.n2231 gnd 0.006712f
C3496 vdd.n2232 gnd 0.006712f
C3497 vdd.n2233 gnd 0.006712f
C3498 vdd.n2234 gnd 0.006712f
C3499 vdd.n2235 gnd 0.006712f
C3500 vdd.n2236 gnd 0.006712f
C3501 vdd.n2237 gnd 0.006712f
C3502 vdd.n2238 gnd 0.006712f
C3503 vdd.n2239 gnd 0.006712f
C3504 vdd.n2240 gnd 0.006712f
C3505 vdd.n2241 gnd 0.015927f
C3506 vdd.n2242 gnd 0.014871f
C3507 vdd.n2243 gnd 0.014871f
C3508 vdd.n2244 gnd 0.837298f
C3509 vdd.n2245 gnd 0.014871f
C3510 vdd.n2246 gnd 0.015927f
C3511 vdd.n2247 gnd 0.01511f
C3512 vdd.n2248 gnd 0.006712f
C3513 vdd.n2249 gnd 0.006712f
C3514 vdd.n2250 gnd 0.006712f
C3515 vdd.n2251 gnd 0.005182f
C3516 vdd.n2252 gnd 0.009593f
C3517 vdd.n2253 gnd 0.004886f
C3518 vdd.n2254 gnd 0.006712f
C3519 vdd.n2255 gnd 0.006712f
C3520 vdd.n2256 gnd 0.006712f
C3521 vdd.n2257 gnd 0.006712f
C3522 vdd.n2258 gnd 0.006712f
C3523 vdd.n2259 gnd 0.006712f
C3524 vdd.n2260 gnd 0.006712f
C3525 vdd.n2261 gnd 0.006712f
C3526 vdd.n2262 gnd 0.006712f
C3527 vdd.n2263 gnd 0.006712f
C3528 vdd.n2264 gnd 0.006712f
C3529 vdd.n2265 gnd 0.006712f
C3530 vdd.n2266 gnd 0.006712f
C3531 vdd.n2267 gnd 0.006712f
C3532 vdd.n2268 gnd 0.006712f
C3533 vdd.n2269 gnd 0.006712f
C3534 vdd.n2270 gnd 0.006712f
C3535 vdd.n2271 gnd 0.006712f
C3536 vdd.n2272 gnd 0.006712f
C3537 vdd.n2273 gnd 0.006712f
C3538 vdd.n2274 gnd 0.006712f
C3539 vdd.n2275 gnd 0.006712f
C3540 vdd.n2276 gnd 0.006712f
C3541 vdd.n2277 gnd 0.006712f
C3542 vdd.n2278 gnd 0.006712f
C3543 vdd.n2279 gnd 0.006712f
C3544 vdd.n2280 gnd 0.006712f
C3545 vdd.n2281 gnd 0.006712f
C3546 vdd.n2282 gnd 0.006712f
C3547 vdd.n2283 gnd 0.006712f
C3548 vdd.n2284 gnd 0.006712f
C3549 vdd.n2285 gnd 0.006712f
C3550 vdd.n2286 gnd 0.006712f
C3551 vdd.n2287 gnd 0.006712f
C3552 vdd.n2288 gnd 0.006712f
C3553 vdd.n2289 gnd 0.006712f
C3554 vdd.n2290 gnd 0.006712f
C3555 vdd.n2291 gnd 0.006712f
C3556 vdd.n2292 gnd 0.006712f
C3557 vdd.n2293 gnd 0.006712f
C3558 vdd.n2294 gnd 0.006712f
C3559 vdd.n2295 gnd 0.006712f
C3560 vdd.n2296 gnd 0.006712f
C3561 vdd.n2297 gnd 0.006712f
C3562 vdd.n2298 gnd 0.006712f
C3563 vdd.n2299 gnd 0.006712f
C3564 vdd.n2300 gnd 0.006712f
C3565 vdd.n2301 gnd 0.006712f
C3566 vdd.n2302 gnd 0.006712f
C3567 vdd.n2303 gnd 0.006712f
C3568 vdd.n2304 gnd 0.006712f
C3569 vdd.n2305 gnd 0.006712f
C3570 vdd.n2306 gnd 0.006712f
C3571 vdd.n2307 gnd 0.006712f
C3572 vdd.n2308 gnd 0.006712f
C3573 vdd.n2309 gnd 0.006712f
C3574 vdd.n2310 gnd 0.006712f
C3575 vdd.n2311 gnd 0.006712f
C3576 vdd.n2312 gnd 0.006712f
C3577 vdd.n2313 gnd 0.006712f
C3578 vdd.n2314 gnd 0.015927f
C3579 vdd.n2315 gnd 0.015927f
C3580 vdd.n2316 gnd 0.837298f
C3581 vdd.t176 gnd 2.97594f
C3582 vdd.t77 gnd 2.97594f
C3583 vdd.n2349 gnd 0.015927f
C3584 vdd.n2350 gnd 0.006712f
C3585 vdd.t124 gnd 0.271249f
C3586 vdd.t125 gnd 0.277657f
C3587 vdd.t122 gnd 0.177082f
C3588 vdd.n2351 gnd 0.095703f
C3589 vdd.n2352 gnd 0.054286f
C3590 vdd.n2353 gnd 0.006712f
C3591 vdd.t138 gnd 0.271249f
C3592 vdd.t139 gnd 0.277657f
C3593 vdd.t137 gnd 0.177082f
C3594 vdd.n2354 gnd 0.095703f
C3595 vdd.n2355 gnd 0.054286f
C3596 vdd.n2356 gnd 0.009593f
C3597 vdd.n2357 gnd 0.006712f
C3598 vdd.n2358 gnd 0.006712f
C3599 vdd.n2359 gnd 0.006712f
C3600 vdd.n2360 gnd 0.006712f
C3601 vdd.n2361 gnd 0.006712f
C3602 vdd.n2362 gnd 0.006712f
C3603 vdd.n2363 gnd 0.006712f
C3604 vdd.n2364 gnd 0.006712f
C3605 vdd.n2365 gnd 0.006712f
C3606 vdd.n2366 gnd 0.006712f
C3607 vdd.n2367 gnd 0.006712f
C3608 vdd.n2368 gnd 0.006712f
C3609 vdd.n2369 gnd 0.006712f
C3610 vdd.n2370 gnd 0.006712f
C3611 vdd.n2371 gnd 0.006712f
C3612 vdd.n2372 gnd 0.006712f
C3613 vdd.n2373 gnd 0.006712f
C3614 vdd.n2374 gnd 0.006712f
C3615 vdd.n2375 gnd 0.006712f
C3616 vdd.n2376 gnd 0.006712f
C3617 vdd.n2377 gnd 0.006712f
C3618 vdd.n2378 gnd 0.006712f
C3619 vdd.n2379 gnd 0.006712f
C3620 vdd.n2380 gnd 0.006712f
C3621 vdd.n2381 gnd 0.006712f
C3622 vdd.n2382 gnd 0.006712f
C3623 vdd.n2383 gnd 0.006712f
C3624 vdd.n2384 gnd 0.006712f
C3625 vdd.n2385 gnd 0.006712f
C3626 vdd.n2386 gnd 0.006712f
C3627 vdd.n2387 gnd 0.006712f
C3628 vdd.n2388 gnd 0.006712f
C3629 vdd.n2389 gnd 0.006712f
C3630 vdd.n2390 gnd 0.006712f
C3631 vdd.n2391 gnd 0.006712f
C3632 vdd.n2392 gnd 0.006712f
C3633 vdd.n2393 gnd 0.006712f
C3634 vdd.n2394 gnd 0.006712f
C3635 vdd.n2395 gnd 0.006712f
C3636 vdd.n2396 gnd 0.006712f
C3637 vdd.n2397 gnd 0.006712f
C3638 vdd.n2398 gnd 0.006712f
C3639 vdd.n2399 gnd 0.006712f
C3640 vdd.n2400 gnd 0.006712f
C3641 vdd.n2401 gnd 0.006712f
C3642 vdd.n2402 gnd 0.006712f
C3643 vdd.n2403 gnd 0.006712f
C3644 vdd.n2404 gnd 0.006712f
C3645 vdd.n2405 gnd 0.006712f
C3646 vdd.n2406 gnd 0.006712f
C3647 vdd.n2407 gnd 0.006712f
C3648 vdd.n2408 gnd 0.006712f
C3649 vdd.n2409 gnd 0.006712f
C3650 vdd.n2410 gnd 0.006712f
C3651 vdd.n2411 gnd 0.006712f
C3652 vdd.n2412 gnd 0.006712f
C3653 vdd.n2413 gnd 0.004886f
C3654 vdd.n2414 gnd 0.006712f
C3655 vdd.n2415 gnd 0.006712f
C3656 vdd.n2416 gnd 0.005182f
C3657 vdd.n2417 gnd 0.006712f
C3658 vdd.n2418 gnd 0.006712f
C3659 vdd.n2419 gnd 0.015927f
C3660 vdd.n2420 gnd 0.014871f
C3661 vdd.n2421 gnd 0.006712f
C3662 vdd.n2422 gnd 0.006712f
C3663 vdd.n2423 gnd 0.006712f
C3664 vdd.n2424 gnd 0.006712f
C3665 vdd.n2425 gnd 0.006712f
C3666 vdd.n2426 gnd 0.006712f
C3667 vdd.n2427 gnd 0.006712f
C3668 vdd.n2428 gnd 0.006712f
C3669 vdd.n2429 gnd 0.006712f
C3670 vdd.n2430 gnd 0.006712f
C3671 vdd.n2431 gnd 0.006712f
C3672 vdd.n2432 gnd 0.006712f
C3673 vdd.n2433 gnd 0.006712f
C3674 vdd.n2434 gnd 0.006712f
C3675 vdd.n2435 gnd 0.006712f
C3676 vdd.n2436 gnd 0.006712f
C3677 vdd.n2437 gnd 0.006712f
C3678 vdd.n2438 gnd 0.006712f
C3679 vdd.n2439 gnd 0.006712f
C3680 vdd.n2440 gnd 0.006712f
C3681 vdd.n2441 gnd 0.006712f
C3682 vdd.n2442 gnd 0.006712f
C3683 vdd.n2443 gnd 0.006712f
C3684 vdd.n2444 gnd 0.006712f
C3685 vdd.n2445 gnd 0.006712f
C3686 vdd.n2446 gnd 0.006712f
C3687 vdd.n2447 gnd 0.006712f
C3688 vdd.n2448 gnd 0.006712f
C3689 vdd.n2449 gnd 0.006712f
C3690 vdd.n2450 gnd 0.006712f
C3691 vdd.n2451 gnd 0.006712f
C3692 vdd.n2452 gnd 0.006712f
C3693 vdd.n2453 gnd 0.006712f
C3694 vdd.n2454 gnd 0.006712f
C3695 vdd.n2455 gnd 0.006712f
C3696 vdd.n2456 gnd 0.006712f
C3697 vdd.n2457 gnd 0.006712f
C3698 vdd.n2458 gnd 0.006712f
C3699 vdd.n2459 gnd 0.006712f
C3700 vdd.n2460 gnd 0.006712f
C3701 vdd.n2461 gnd 0.006712f
C3702 vdd.n2462 gnd 0.006712f
C3703 vdd.n2463 gnd 0.006712f
C3704 vdd.n2464 gnd 0.006712f
C3705 vdd.n2465 gnd 0.006712f
C3706 vdd.n2466 gnd 0.006712f
C3707 vdd.n2467 gnd 0.006712f
C3708 vdd.n2468 gnd 0.006712f
C3709 vdd.n2469 gnd 0.006712f
C3710 vdd.n2470 gnd 0.006712f
C3711 vdd.n2471 gnd 0.006712f
C3712 vdd.n2472 gnd 0.216891f
C3713 vdd.n2473 gnd 0.006712f
C3714 vdd.n2474 gnd 0.006712f
C3715 vdd.n2475 gnd 0.006712f
C3716 vdd.n2476 gnd 0.006712f
C3717 vdd.n2477 gnd 0.006712f
C3718 vdd.n2478 gnd 0.006712f
C3719 vdd.n2479 gnd 0.006712f
C3720 vdd.n2480 gnd 0.006712f
C3721 vdd.n2481 gnd 0.006712f
C3722 vdd.n2482 gnd 0.006712f
C3723 vdd.n2483 gnd 0.006712f
C3724 vdd.n2484 gnd 0.006712f
C3725 vdd.n2485 gnd 0.006712f
C3726 vdd.n2486 gnd 0.006712f
C3727 vdd.n2487 gnd 0.006712f
C3728 vdd.n2488 gnd 0.006712f
C3729 vdd.n2489 gnd 0.006712f
C3730 vdd.n2490 gnd 0.006712f
C3731 vdd.n2491 gnd 0.006712f
C3732 vdd.n2492 gnd 0.006712f
C3733 vdd.n2493 gnd 0.408561f
C3734 vdd.n2494 gnd 0.006712f
C3735 vdd.n2495 gnd 0.006712f
C3736 vdd.n2496 gnd 0.006712f
C3737 vdd.n2497 gnd 0.006712f
C3738 vdd.n2498 gnd 0.006712f
C3739 vdd.n2499 gnd 0.014871f
C3740 vdd.n2500 gnd 0.015927f
C3741 vdd.n2501 gnd 0.015927f
C3742 vdd.n2502 gnd 0.006712f
C3743 vdd.n2503 gnd 0.006712f
C3744 vdd.n2504 gnd 0.006712f
C3745 vdd.n2505 gnd 0.005182f
C3746 vdd.n2506 gnd 0.009593f
C3747 vdd.n2507 gnd 0.004886f
C3748 vdd.n2508 gnd 0.006712f
C3749 vdd.n2509 gnd 0.006712f
C3750 vdd.n2510 gnd 0.006712f
C3751 vdd.n2511 gnd 0.006712f
C3752 vdd.n2512 gnd 0.006712f
C3753 vdd.n2513 gnd 0.006712f
C3754 vdd.n2514 gnd 0.006712f
C3755 vdd.n2515 gnd 0.006712f
C3756 vdd.n2516 gnd 0.006712f
C3757 vdd.n2517 gnd 0.006712f
C3758 vdd.n2518 gnd 0.006712f
C3759 vdd.n2519 gnd 0.006712f
C3760 vdd.n2520 gnd 0.006712f
C3761 vdd.n2521 gnd 0.006712f
C3762 vdd.n2522 gnd 0.006712f
C3763 vdd.n2523 gnd 0.006712f
C3764 vdd.n2524 gnd 0.006712f
C3765 vdd.n2525 gnd 0.006712f
C3766 vdd.n2526 gnd 0.006712f
C3767 vdd.n2527 gnd 0.006712f
C3768 vdd.n2528 gnd 0.006712f
C3769 vdd.n2529 gnd 0.006712f
C3770 vdd.n2530 gnd 0.006712f
C3771 vdd.n2531 gnd 0.006712f
C3772 vdd.n2532 gnd 0.006712f
C3773 vdd.n2533 gnd 0.006712f
C3774 vdd.n2534 gnd 0.006712f
C3775 vdd.n2535 gnd 0.006712f
C3776 vdd.n2536 gnd 0.006712f
C3777 vdd.n2537 gnd 0.006712f
C3778 vdd.n2538 gnd 0.006712f
C3779 vdd.n2539 gnd 0.006712f
C3780 vdd.n2540 gnd 0.006712f
C3781 vdd.n2541 gnd 0.006712f
C3782 vdd.n2542 gnd 0.006712f
C3783 vdd.n2543 gnd 0.006712f
C3784 vdd.n2544 gnd 0.006712f
C3785 vdd.n2545 gnd 0.006712f
C3786 vdd.n2546 gnd 0.006712f
C3787 vdd.n2547 gnd 0.006712f
C3788 vdd.n2548 gnd 0.006712f
C3789 vdd.n2549 gnd 0.006712f
C3790 vdd.n2550 gnd 0.006712f
C3791 vdd.n2551 gnd 0.006712f
C3792 vdd.n2552 gnd 0.006712f
C3793 vdd.n2553 gnd 0.006712f
C3794 vdd.n2554 gnd 0.006712f
C3795 vdd.n2555 gnd 0.006712f
C3796 vdd.n2556 gnd 0.006712f
C3797 vdd.n2557 gnd 0.006712f
C3798 vdd.n2558 gnd 0.006712f
C3799 vdd.n2559 gnd 0.006712f
C3800 vdd.n2560 gnd 0.006712f
C3801 vdd.n2561 gnd 0.006712f
C3802 vdd.n2562 gnd 0.006712f
C3803 vdd.n2563 gnd 0.006712f
C3804 vdd.n2564 gnd 0.006712f
C3805 vdd.n2565 gnd 0.006712f
C3806 vdd.n2566 gnd 0.006712f
C3807 vdd.n2567 gnd 0.006712f
C3808 vdd.n2569 gnd 0.837298f
C3809 vdd.n2571 gnd 0.006712f
C3810 vdd.n2572 gnd 0.006712f
C3811 vdd.n2573 gnd 0.015927f
C3812 vdd.n2574 gnd 0.014871f
C3813 vdd.n2575 gnd 0.014871f
C3814 vdd.n2576 gnd 0.837298f
C3815 vdd.n2577 gnd 0.014871f
C3816 vdd.n2578 gnd 0.014871f
C3817 vdd.n2579 gnd 0.006712f
C3818 vdd.n2580 gnd 0.006712f
C3819 vdd.n2581 gnd 0.006712f
C3820 vdd.n2582 gnd 0.428737f
C3821 vdd.n2583 gnd 0.006712f
C3822 vdd.n2584 gnd 0.006712f
C3823 vdd.n2585 gnd 0.006712f
C3824 vdd.n2586 gnd 0.006712f
C3825 vdd.n2587 gnd 0.006712f
C3826 vdd.n2588 gnd 0.53466f
C3827 vdd.n2589 gnd 0.006712f
C3828 vdd.n2590 gnd 0.006712f
C3829 vdd.n2591 gnd 0.006712f
C3830 vdd.n2592 gnd 0.006712f
C3831 vdd.n2593 gnd 0.006712f
C3832 vdd.n2594 gnd 0.685979f
C3833 vdd.n2595 gnd 0.006712f
C3834 vdd.n2596 gnd 0.006712f
C3835 vdd.n2597 gnd 0.006712f
C3836 vdd.n2598 gnd 0.006712f
C3837 vdd.n2599 gnd 0.006712f
C3838 vdd.n2600 gnd 0.378297f
C3839 vdd.n2601 gnd 0.006712f
C3840 vdd.n2602 gnd 0.006712f
C3841 vdd.n2603 gnd 0.006712f
C3842 vdd.n2604 gnd 0.006712f
C3843 vdd.n2605 gnd 0.006712f
C3844 vdd.n2606 gnd 0.216891f
C3845 vdd.n2607 gnd 0.006712f
C3846 vdd.n2608 gnd 0.006712f
C3847 vdd.n2609 gnd 0.006712f
C3848 vdd.n2610 gnd 0.006712f
C3849 vdd.n2611 gnd 0.006712f
C3850 vdd.n2612 gnd 0.393429f
C3851 vdd.n2613 gnd 0.006712f
C3852 vdd.n2614 gnd 0.006712f
C3853 vdd.n2615 gnd 0.006712f
C3854 vdd.n2616 gnd 0.006712f
C3855 vdd.n2617 gnd 0.006712f
C3856 vdd.n2618 gnd 0.544748f
C3857 vdd.n2619 gnd 0.006712f
C3858 vdd.n2620 gnd 0.006712f
C3859 vdd.n2621 gnd 0.006712f
C3860 vdd.n2622 gnd 0.006712f
C3861 vdd.n2623 gnd 0.006712f
C3862 vdd.n2624 gnd 0.61032f
C3863 vdd.n2625 gnd 0.006712f
C3864 vdd.n2626 gnd 0.006712f
C3865 vdd.n2627 gnd 0.006712f
C3866 vdd.n2628 gnd 0.006712f
C3867 vdd.n2629 gnd 0.006712f
C3868 vdd.n2630 gnd 0.459001f
C3869 vdd.n2631 gnd 0.006712f
C3870 vdd.n2632 gnd 0.006712f
C3871 vdd.n2633 gnd 0.006712f
C3872 vdd.t103 gnd 0.277657f
C3873 vdd.t101 gnd 0.177082f
C3874 vdd.t104 gnd 0.277657f
C3875 vdd.n2634 gnd 0.156054f
C3876 vdd.n2635 gnd 0.019445f
C3877 vdd.n2636 gnd 0.004146f
C3878 vdd.n2637 gnd 0.006712f
C3879 vdd.n2638 gnd 0.378297f
C3880 vdd.n2639 gnd 0.006712f
C3881 vdd.n2640 gnd 0.006712f
C3882 vdd.n2641 gnd 0.006712f
C3883 vdd.n2642 gnd 0.006712f
C3884 vdd.n2643 gnd 0.006712f
C3885 vdd.n2644 gnd 0.685979f
C3886 vdd.n2645 gnd 0.006712f
C3887 vdd.n2646 gnd 0.006712f
C3888 vdd.n2647 gnd 0.006712f
C3889 vdd.n2648 gnd 0.006712f
C3890 vdd.n2649 gnd 0.006712f
C3891 vdd.n2650 gnd 0.006712f
C3892 vdd.n2652 gnd 0.006712f
C3893 vdd.n2653 gnd 0.006712f
C3894 vdd.n2655 gnd 0.006712f
C3895 vdd.n2656 gnd 0.006712f
C3896 vdd.n2659 gnd 0.006712f
C3897 vdd.n2660 gnd 0.006712f
C3898 vdd.n2661 gnd 0.006712f
C3899 vdd.n2662 gnd 0.006712f
C3900 vdd.n2664 gnd 0.006712f
C3901 vdd.n2665 gnd 0.006712f
C3902 vdd.n2666 gnd 0.006712f
C3903 vdd.n2667 gnd 0.006712f
C3904 vdd.n2668 gnd 0.006712f
C3905 vdd.n2669 gnd 0.006712f
C3906 vdd.n2671 gnd 0.006712f
C3907 vdd.n2672 gnd 0.006712f
C3908 vdd.n2673 gnd 0.006712f
C3909 vdd.n2674 gnd 0.006712f
C3910 vdd.n2675 gnd 0.006712f
C3911 vdd.n2676 gnd 0.006712f
C3912 vdd.n2678 gnd 0.006712f
C3913 vdd.n2679 gnd 0.006712f
C3914 vdd.n2680 gnd 0.006712f
C3915 vdd.n2681 gnd 0.006712f
C3916 vdd.n2682 gnd 0.006712f
C3917 vdd.n2683 gnd 0.006712f
C3918 vdd.n2685 gnd 0.006712f
C3919 vdd.n2686 gnd 0.015927f
C3920 vdd.n2687 gnd 0.015927f
C3921 vdd.n2688 gnd 0.014871f
C3922 vdd.n2689 gnd 0.006712f
C3923 vdd.n2690 gnd 0.006712f
C3924 vdd.n2691 gnd 0.006712f
C3925 vdd.n2692 gnd 0.006712f
C3926 vdd.n2693 gnd 0.006712f
C3927 vdd.n2694 gnd 0.006712f
C3928 vdd.n2695 gnd 0.685979f
C3929 vdd.n2696 gnd 0.006712f
C3930 vdd.n2697 gnd 0.006712f
C3931 vdd.n2698 gnd 0.006712f
C3932 vdd.n2699 gnd 0.006712f
C3933 vdd.n2700 gnd 0.006712f
C3934 vdd.n2701 gnd 0.428737f
C3935 vdd.n2702 gnd 0.006712f
C3936 vdd.n2703 gnd 0.006712f
C3937 vdd.n2704 gnd 0.006712f
C3938 vdd.n2705 gnd 0.015688f
C3939 vdd.n2707 gnd 0.015927f
C3940 vdd.n2708 gnd 0.01511f
C3941 vdd.n2709 gnd 0.006712f
C3942 vdd.n2710 gnd 0.005182f
C3943 vdd.n2711 gnd 0.006712f
C3944 vdd.n2713 gnd 0.006712f
C3945 vdd.n2714 gnd 0.006712f
C3946 vdd.n2715 gnd 0.006712f
C3947 vdd.n2716 gnd 0.006712f
C3948 vdd.n2717 gnd 0.006712f
C3949 vdd.n2718 gnd 0.006712f
C3950 vdd.n2720 gnd 0.006712f
C3951 vdd.n2721 gnd 0.006712f
C3952 vdd.n2722 gnd 0.006712f
C3953 vdd.n2723 gnd 0.006712f
C3954 vdd.n2724 gnd 0.006712f
C3955 vdd.n2725 gnd 0.006712f
C3956 vdd.n2727 gnd 0.006712f
C3957 vdd.n2728 gnd 0.006712f
C3958 vdd.n2729 gnd 0.006712f
C3959 vdd.n2730 gnd 0.006712f
C3960 vdd.n2731 gnd 0.006712f
C3961 vdd.n2732 gnd 0.006712f
C3962 vdd.n2734 gnd 0.006712f
C3963 vdd.n2735 gnd 0.006712f
C3964 vdd.n2736 gnd 0.006712f
C3965 vdd.n2737 gnd 0.597423f
C3966 vdd.n2738 gnd 0.01613f
C3967 vdd.n2739 gnd 0.006712f
C3968 vdd.n2740 gnd 0.006712f
C3969 vdd.n2742 gnd 0.006712f
C3970 vdd.n2743 gnd 0.006712f
C3971 vdd.n2744 gnd 0.006712f
C3972 vdd.n2745 gnd 0.006712f
C3973 vdd.n2746 gnd 0.006712f
C3974 vdd.n2747 gnd 0.006712f
C3975 vdd.n2749 gnd 0.006712f
C3976 vdd.n2750 gnd 0.006712f
C3977 vdd.n2751 gnd 0.006712f
C3978 vdd.n2752 gnd 0.006712f
C3979 vdd.n2753 gnd 0.006712f
C3980 vdd.n2754 gnd 0.006712f
C3981 vdd.n2756 gnd 0.006712f
C3982 vdd.n2757 gnd 0.006712f
C3983 vdd.n2758 gnd 0.006712f
C3984 vdd.n2759 gnd 0.006712f
C3985 vdd.n2760 gnd 0.006712f
C3986 vdd.n2761 gnd 0.006712f
C3987 vdd.n2763 gnd 0.006712f
C3988 vdd.n2764 gnd 0.006712f
C3989 vdd.n2766 gnd 0.006712f
C3990 vdd.n2767 gnd 0.006712f
C3991 vdd.n2768 gnd 0.015927f
C3992 vdd.n2769 gnd 0.014871f
C3993 vdd.n2770 gnd 0.014871f
C3994 vdd.n2771 gnd 0.988617f
C3995 vdd.n2772 gnd 0.014871f
C3996 vdd.n2773 gnd 0.015927f
C3997 vdd.n2774 gnd 0.01511f
C3998 vdd.n2775 gnd 0.006712f
C3999 vdd.n2776 gnd 0.005182f
C4000 vdd.n2777 gnd 0.006712f
C4001 vdd.n2779 gnd 0.006712f
C4002 vdd.n2780 gnd 0.006712f
C4003 vdd.n2781 gnd 0.006712f
C4004 vdd.n2782 gnd 0.006712f
C4005 vdd.n2783 gnd 0.006712f
C4006 vdd.n2784 gnd 0.006712f
C4007 vdd.n2786 gnd 0.006712f
C4008 vdd.n2787 gnd 0.006712f
C4009 vdd.n2788 gnd 0.006712f
C4010 vdd.n2789 gnd 0.006712f
C4011 vdd.n2790 gnd 0.006712f
C4012 vdd.n2791 gnd 0.006712f
C4013 vdd.n2793 gnd 0.006712f
C4014 vdd.n2794 gnd 0.006712f
C4015 vdd.n2795 gnd 0.006712f
C4016 vdd.n2796 gnd 0.006712f
C4017 vdd.n2797 gnd 0.006712f
C4018 vdd.n2798 gnd 0.006712f
C4019 vdd.n2800 gnd 0.006712f
C4020 vdd.n2801 gnd 0.006712f
C4021 vdd.n2803 gnd 0.006712f
C4022 vdd.n2804 gnd 0.01613f
C4023 vdd.n2805 gnd 0.597423f
C4024 vdd.n2806 gnd 0.008489f
C4025 vdd.n2807 gnd 0.003774f
C4026 vdd.t144 gnd 0.121442f
C4027 vdd.t145 gnd 0.129788f
C4028 vdd.t143 gnd 0.158602f
C4029 vdd.n2808 gnd 0.203305f
C4030 vdd.n2809 gnd 0.170813f
C4031 vdd.n2810 gnd 0.012235f
C4032 vdd.n2811 gnd 0.009871f
C4033 vdd.n2812 gnd 0.004171f
C4034 vdd.n2813 gnd 0.007945f
C4035 vdd.n2814 gnd 0.009871f
C4036 vdd.n2815 gnd 0.009871f
C4037 vdd.n2816 gnd 0.007945f
C4038 vdd.n2817 gnd 0.007945f
C4039 vdd.n2818 gnd 0.009871f
C4040 vdd.n2820 gnd 0.009871f
C4041 vdd.n2821 gnd 0.007945f
C4042 vdd.n2822 gnd 0.007945f
C4043 vdd.n2823 gnd 0.007945f
C4044 vdd.n2824 gnd 0.009871f
C4045 vdd.n2826 gnd 0.009871f
C4046 vdd.n2828 gnd 0.009871f
C4047 vdd.n2829 gnd 0.007945f
C4048 vdd.n2830 gnd 0.007945f
C4049 vdd.n2831 gnd 0.007945f
C4050 vdd.n2832 gnd 0.009871f
C4051 vdd.n2834 gnd 0.009871f
C4052 vdd.n2836 gnd 0.009871f
C4053 vdd.n2837 gnd 0.007945f
C4054 vdd.n2838 gnd 0.007945f
C4055 vdd.n2839 gnd 0.007945f
C4056 vdd.n2840 gnd 0.009871f
C4057 vdd.n2842 gnd 0.009871f
C4058 vdd.n2843 gnd 0.009871f
C4059 vdd.n2844 gnd 0.007945f
C4060 vdd.n2845 gnd 0.007945f
C4061 vdd.n2846 gnd 0.009871f
C4062 vdd.n2847 gnd 0.009871f
C4063 vdd.n2849 gnd 0.009871f
C4064 vdd.n2850 gnd 0.007945f
C4065 vdd.n2851 gnd 0.009871f
C4066 vdd.n2852 gnd 0.009871f
C4067 vdd.n2853 gnd 0.009871f
C4068 vdd.n2854 gnd 0.016208f
C4069 vdd.n2855 gnd 0.005403f
C4070 vdd.n2856 gnd 0.009871f
C4071 vdd.n2858 gnd 0.009871f
C4072 vdd.n2860 gnd 0.009871f
C4073 vdd.n2861 gnd 0.007945f
C4074 vdd.n2862 gnd 0.007945f
C4075 vdd.n2863 gnd 0.007945f
C4076 vdd.n2864 gnd 0.009871f
C4077 vdd.n2866 gnd 0.009871f
C4078 vdd.n2868 gnd 0.009871f
C4079 vdd.n2869 gnd 0.007945f
C4080 vdd.n2870 gnd 0.007945f
C4081 vdd.n2871 gnd 0.007945f
C4082 vdd.n2872 gnd 0.009871f
C4083 vdd.n2874 gnd 0.009871f
C4084 vdd.n2876 gnd 0.009871f
C4085 vdd.n2877 gnd 0.007945f
C4086 vdd.n2878 gnd 0.007945f
C4087 vdd.n2879 gnd 0.007945f
C4088 vdd.n2880 gnd 0.009871f
C4089 vdd.n2882 gnd 0.009871f
C4090 vdd.n2884 gnd 0.009871f
C4091 vdd.n2885 gnd 0.007945f
C4092 vdd.n2886 gnd 0.007945f
C4093 vdd.n2887 gnd 0.007945f
C4094 vdd.n2888 gnd 0.009871f
C4095 vdd.n2890 gnd 0.009871f
C4096 vdd.n2892 gnd 0.009871f
C4097 vdd.n2893 gnd 0.007945f
C4098 vdd.n2894 gnd 0.007945f
C4099 vdd.n2895 gnd 0.006634f
C4100 vdd.n2896 gnd 0.009871f
C4101 vdd.n2898 gnd 0.009871f
C4102 vdd.n2900 gnd 0.009871f
C4103 vdd.n2901 gnd 0.006634f
C4104 vdd.n2902 gnd 0.007945f
C4105 vdd.n2903 gnd 0.007945f
C4106 vdd.n2904 gnd 0.009871f
C4107 vdd.n2906 gnd 0.009871f
C4108 vdd.n2908 gnd 0.009871f
C4109 vdd.n2909 gnd 0.007945f
C4110 vdd.n2910 gnd 0.007945f
C4111 vdd.n2911 gnd 0.007945f
C4112 vdd.n2912 gnd 0.009871f
C4113 vdd.n2914 gnd 0.009871f
C4114 vdd.n2916 gnd 0.009871f
C4115 vdd.n2917 gnd 0.007945f
C4116 vdd.n2918 gnd 0.007945f
C4117 vdd.n2919 gnd 0.007945f
C4118 vdd.n2920 gnd 0.009871f
C4119 vdd.n2922 gnd 0.009871f
C4120 vdd.n2923 gnd 0.009871f
C4121 vdd.n2924 gnd 0.007945f
C4122 vdd.n2925 gnd 0.007945f
C4123 vdd.n2926 gnd 0.009871f
C4124 vdd.n2927 gnd 0.009871f
C4125 vdd.n2928 gnd 0.007945f
C4126 vdd.n2929 gnd 0.007945f
C4127 vdd.n2930 gnd 0.009871f
C4128 vdd.n2931 gnd 0.009871f
C4129 vdd.n2933 gnd 0.009871f
C4130 vdd.n2934 gnd 0.007945f
C4131 vdd.n2935 gnd 0.006594f
C4132 vdd.n2936 gnd 0.023626f
C4133 vdd.n2937 gnd 0.023262f
C4134 vdd.n2938 gnd 0.006594f
C4135 vdd.n2939 gnd 0.023262f
C4136 vdd.n2940 gnd 1.38709f
C4137 vdd.n2941 gnd 0.023262f
C4138 vdd.n2942 gnd 0.006594f
C4139 vdd.n2943 gnd 0.023262f
C4140 vdd.n2944 gnd 0.009871f
C4141 vdd.n2945 gnd 0.009871f
C4142 vdd.n2946 gnd 0.007945f
C4143 vdd.n2947 gnd 0.009871f
C4144 vdd.n2948 gnd 1.00879f
C4145 vdd.n2949 gnd 0.009871f
C4146 vdd.n2950 gnd 0.007945f
C4147 vdd.n2951 gnd 0.009871f
C4148 vdd.n2952 gnd 0.009871f
C4149 vdd.n2953 gnd 0.009871f
C4150 vdd.n2954 gnd 0.007945f
C4151 vdd.n2955 gnd 0.009871f
C4152 vdd.n2956 gnd 0.892782f
C4153 vdd.n2957 gnd 0.009871f
C4154 vdd.n2958 gnd 0.007945f
C4155 vdd.n2959 gnd 0.009871f
C4156 vdd.n2960 gnd 0.009871f
C4157 vdd.n2961 gnd 0.009871f
C4158 vdd.n2962 gnd 0.007945f
C4159 vdd.n2963 gnd 0.009871f
C4160 vdd.t34 gnd 0.504397f
C4161 vdd.n2964 gnd 0.721287f
C4162 vdd.n2965 gnd 0.009871f
C4163 vdd.n2966 gnd 0.007945f
C4164 vdd.n2967 gnd 0.009871f
C4165 vdd.n2968 gnd 0.009871f
C4166 vdd.n2969 gnd 0.009871f
C4167 vdd.n2970 gnd 0.007945f
C4168 vdd.n2971 gnd 0.009871f
C4169 vdd.n2972 gnd 0.549792f
C4170 vdd.n2973 gnd 0.009871f
C4171 vdd.n2974 gnd 0.007945f
C4172 vdd.n2975 gnd 0.009871f
C4173 vdd.n2976 gnd 0.009871f
C4174 vdd.n2977 gnd 0.009871f
C4175 vdd.n2978 gnd 0.007945f
C4176 vdd.n2979 gnd 0.009871f
C4177 vdd.n2980 gnd 0.711199f
C4178 vdd.n2981 gnd 0.630496f
C4179 vdd.n2982 gnd 0.009871f
C4180 vdd.n2983 gnd 0.007945f
C4181 vdd.n2984 gnd 0.009871f
C4182 vdd.n2985 gnd 0.009871f
C4183 vdd.n2986 gnd 0.009871f
C4184 vdd.n2987 gnd 0.007945f
C4185 vdd.n2988 gnd 0.009871f
C4186 vdd.n2989 gnd 0.801991f
C4187 vdd.n2990 gnd 0.009871f
C4188 vdd.n2991 gnd 0.007945f
C4189 vdd.n2992 gnd 0.009871f
C4190 vdd.n2993 gnd 0.009871f
C4191 vdd.n2994 gnd 0.009871f
C4192 vdd.n2995 gnd 0.007945f
C4193 vdd.n2996 gnd 0.007945f
C4194 vdd.n2997 gnd 0.007945f
C4195 vdd.n2998 gnd 0.009871f
C4196 vdd.n2999 gnd 0.009871f
C4197 vdd.n3000 gnd 0.009871f
C4198 vdd.n3001 gnd 0.007945f
C4199 vdd.n3002 gnd 0.007945f
C4200 vdd.n3003 gnd 0.007945f
C4201 vdd.n3004 gnd 0.009871f
C4202 vdd.n3005 gnd 0.009871f
C4203 vdd.n3006 gnd 0.009871f
C4204 vdd.n3007 gnd 0.007945f
C4205 vdd.n3008 gnd 0.007945f
C4206 vdd.n3009 gnd 0.007945f
C4207 vdd.n3010 gnd 0.009871f
C4208 vdd.n3011 gnd 0.009871f
C4209 vdd.n3012 gnd 0.009871f
C4210 vdd.n3013 gnd 0.007945f
C4211 vdd.n3014 gnd 0.007945f
C4212 vdd.n3015 gnd 0.006594f
C4213 vdd.n3016 gnd 0.023262f
C4214 vdd.n3017 gnd 0.023626f
C4215 vdd.n3019 gnd 0.023626f
C4216 vdd.n3020 gnd 0.003774f
C4217 vdd.t155 gnd 0.121442f
C4218 vdd.t154 gnd 0.129788f
C4219 vdd.t153 gnd 0.158602f
C4220 vdd.n3021 gnd 0.203305f
C4221 vdd.n3022 gnd 0.171608f
C4222 vdd.n3023 gnd 0.01303f
C4223 vdd.n3024 gnd 0.004171f
C4224 vdd.n3025 gnd 0.007945f
C4225 vdd.n3026 gnd 0.009871f
C4226 vdd.n3028 gnd 0.009871f
C4227 vdd.n3029 gnd 0.009871f
C4228 vdd.n3030 gnd 0.007945f
C4229 vdd.n3031 gnd 0.007945f
C4230 vdd.n3032 gnd 0.007945f
C4231 vdd.n3033 gnd 0.009871f
C4232 vdd.n3035 gnd 0.009871f
C4233 vdd.n3036 gnd 0.009871f
C4234 vdd.n3037 gnd 0.007945f
C4235 vdd.n3038 gnd 0.007945f
C4236 vdd.n3039 gnd 0.007945f
C4237 vdd.n3040 gnd 0.009871f
C4238 vdd.n3042 gnd 0.009871f
C4239 vdd.n3043 gnd 0.009871f
C4240 vdd.n3044 gnd 0.007945f
C4241 vdd.n3045 gnd 0.007945f
C4242 vdd.n3046 gnd 0.007945f
C4243 vdd.n3047 gnd 0.009871f
C4244 vdd.n3049 gnd 0.009871f
C4245 vdd.n3050 gnd 0.009871f
C4246 vdd.n3051 gnd 0.007945f
C4247 vdd.n3052 gnd 0.007945f
C4248 vdd.n3053 gnd 0.007945f
C4249 vdd.n3054 gnd 0.009871f
C4250 vdd.n3056 gnd 0.009871f
C4251 vdd.n3057 gnd 0.009871f
C4252 vdd.n3058 gnd 0.007945f
C4253 vdd.n3059 gnd 0.009871f
C4254 vdd.n3060 gnd 0.009871f
C4255 vdd.n3061 gnd 0.009871f
C4256 vdd.n3062 gnd 0.017003f
C4257 vdd.n3063 gnd 0.005403f
C4258 vdd.n3064 gnd 0.007945f
C4259 vdd.n3065 gnd 0.009871f
C4260 vdd.n3067 gnd 0.009871f
C4261 vdd.n3068 gnd 0.009871f
C4262 vdd.n3069 gnd 0.007945f
C4263 vdd.n3070 gnd 0.007945f
C4264 vdd.n3071 gnd 0.007945f
C4265 vdd.n3072 gnd 0.009871f
C4266 vdd.n3074 gnd 0.009871f
C4267 vdd.n3075 gnd 0.009871f
C4268 vdd.n3076 gnd 0.007945f
C4269 vdd.n3077 gnd 0.007945f
C4270 vdd.n3078 gnd 0.007945f
C4271 vdd.n3079 gnd 0.009871f
C4272 vdd.n3081 gnd 0.009871f
C4273 vdd.n3082 gnd 0.009871f
C4274 vdd.n3083 gnd 0.007945f
C4275 vdd.n3084 gnd 0.007945f
C4276 vdd.n3085 gnd 0.007945f
C4277 vdd.n3086 gnd 0.009871f
C4278 vdd.n3088 gnd 0.009871f
C4279 vdd.n3089 gnd 0.009871f
C4280 vdd.n3090 gnd 0.007945f
C4281 vdd.n3091 gnd 0.007945f
C4282 vdd.n3092 gnd 0.007945f
C4283 vdd.n3093 gnd 0.009871f
C4284 vdd.n3095 gnd 0.009871f
C4285 vdd.n3096 gnd 0.009871f
C4286 vdd.n3097 gnd 0.007945f
C4287 vdd.n3098 gnd 0.009871f
C4288 vdd.n3099 gnd 0.009871f
C4289 vdd.n3100 gnd 0.009871f
C4290 vdd.n3101 gnd 0.017003f
C4291 vdd.n3102 gnd 0.006634f
C4292 vdd.n3103 gnd 0.007945f
C4293 vdd.n3104 gnd 0.009871f
C4294 vdd.n3106 gnd 0.009871f
C4295 vdd.n3107 gnd 0.009871f
C4296 vdd.n3108 gnd 0.007945f
C4297 vdd.n3109 gnd 0.007945f
C4298 vdd.n3110 gnd 0.007945f
C4299 vdd.n3111 gnd 0.009871f
C4300 vdd.n3113 gnd 0.009871f
C4301 vdd.n3114 gnd 0.009871f
C4302 vdd.n3115 gnd 0.007945f
C4303 vdd.n3116 gnd 0.007945f
C4304 vdd.n3117 gnd 0.007945f
C4305 vdd.n3118 gnd 0.009871f
C4306 vdd.n3120 gnd 0.009871f
C4307 vdd.n3121 gnd 0.009871f
C4308 vdd.n3122 gnd 0.007945f
C4309 vdd.n3123 gnd 0.007945f
C4310 vdd.n3124 gnd 0.007945f
C4311 vdd.n3125 gnd 0.009871f
C4312 vdd.n3127 gnd 0.009871f
C4313 vdd.n3128 gnd 0.009871f
C4314 vdd.n3130 gnd 0.009871f
C4315 vdd.n3131 gnd 0.007945f
C4316 vdd.n3132 gnd 0.007945f
C4317 vdd.n3133 gnd 0.006594f
C4318 vdd.n3134 gnd 0.023626f
C4319 vdd.n3135 gnd 0.023262f
C4320 vdd.n3136 gnd 0.006594f
C4321 vdd.n3137 gnd 0.023262f
C4322 vdd.n3138 gnd 1.4224f
C4323 vdd.n3139 gnd 0.569968f
C4324 vdd.t147 gnd 0.504397f
C4325 vdd.n3140 gnd 0.943222f
C4326 vdd.n3141 gnd 0.009871f
C4327 vdd.n3142 gnd 0.007945f
C4328 vdd.n3143 gnd 0.007945f
C4329 vdd.n3144 gnd 0.007945f
C4330 vdd.n3145 gnd 0.009871f
C4331 vdd.n3146 gnd 0.993661f
C4332 vdd.t4 gnd 0.504397f
C4333 vdd.n3147 gnd 0.519529f
C4334 vdd.n3148 gnd 0.822166f
C4335 vdd.n3149 gnd 0.009871f
C4336 vdd.n3150 gnd 0.007945f
C4337 vdd.n3151 gnd 0.007945f
C4338 vdd.n3152 gnd 0.007945f
C4339 vdd.n3153 gnd 0.009871f
C4340 vdd.n3154 gnd 0.650672f
C4341 vdd.t72 gnd 0.504397f
C4342 vdd.n3155 gnd 0.837298f
C4343 vdd.t24 gnd 0.504397f
C4344 vdd.n3156 gnd 0.529616f
C4345 vdd.n3157 gnd 0.009871f
C4346 vdd.n3158 gnd 0.007945f
C4347 vdd.n3159 gnd 0.007945f
C4348 vdd.n3160 gnd 0.007945f
C4349 vdd.n3161 gnd 0.009871f
C4350 vdd.n3162 gnd 0.701111f
C4351 vdd.n3163 gnd 0.640584f
C4352 vdd.t63 gnd 0.504397f
C4353 vdd.n3164 gnd 0.837298f
C4354 vdd.n3165 gnd 0.009871f
C4355 vdd.n3166 gnd 0.007945f
C4356 vdd.n3167 gnd 0.587612f
C4357 vdd.n3168 gnd 2.17513f
C4358 CSoutput.n0 gnd 0.040642f
C4359 CSoutput.t130 gnd 0.268837f
C4360 CSoutput.n1 gnd 0.121393f
C4361 CSoutput.n2 gnd 0.040642f
C4362 CSoutput.t135 gnd 0.268837f
C4363 CSoutput.n3 gnd 0.032212f
C4364 CSoutput.n4 gnd 0.040642f
C4365 CSoutput.t124 gnd 0.268837f
C4366 CSoutput.n5 gnd 0.027777f
C4367 CSoutput.n6 gnd 0.040642f
C4368 CSoutput.t132 gnd 0.268837f
C4369 CSoutput.t138 gnd 0.268837f
C4370 CSoutput.n7 gnd 0.12007f
C4371 CSoutput.n8 gnd 0.040642f
C4372 CSoutput.t137 gnd 0.268837f
C4373 CSoutput.n9 gnd 0.026483f
C4374 CSoutput.n10 gnd 0.040642f
C4375 CSoutput.t125 gnd 0.268837f
C4376 CSoutput.t136 gnd 0.268837f
C4377 CSoutput.n11 gnd 0.12007f
C4378 CSoutput.n12 gnd 0.040642f
C4379 CSoutput.t134 gnd 0.268837f
C4380 CSoutput.n13 gnd 0.027777f
C4381 CSoutput.n14 gnd 0.040642f
C4382 CSoutput.t123 gnd 0.268837f
C4383 CSoutput.t127 gnd 0.268837f
C4384 CSoutput.n15 gnd 0.12007f
C4385 CSoutput.n16 gnd 0.040642f
C4386 CSoutput.t131 gnd 0.268837f
C4387 CSoutput.n17 gnd 0.029667f
C4388 CSoutput.t141 gnd 0.321268f
C4389 CSoutput.t121 gnd 0.268837f
C4390 CSoutput.n18 gnd 0.153283f
C4391 CSoutput.n19 gnd 0.148738f
C4392 CSoutput.n20 gnd 0.172554f
C4393 CSoutput.n21 gnd 0.040642f
C4394 CSoutput.n22 gnd 0.03392f
C4395 CSoutput.n23 gnd 0.12007f
C4396 CSoutput.n24 gnd 0.032698f
C4397 CSoutput.n25 gnd 0.032212f
C4398 CSoutput.n26 gnd 0.040642f
C4399 CSoutput.n27 gnd 0.040642f
C4400 CSoutput.n28 gnd 0.033659f
C4401 CSoutput.n29 gnd 0.028578f
C4402 CSoutput.n30 gnd 0.122743f
C4403 CSoutput.n31 gnd 0.028971f
C4404 CSoutput.n32 gnd 0.040642f
C4405 CSoutput.n33 gnd 0.040642f
C4406 CSoutput.n34 gnd 0.040642f
C4407 CSoutput.n35 gnd 0.033301f
C4408 CSoutput.n36 gnd 0.12007f
C4409 CSoutput.n37 gnd 0.031847f
C4410 CSoutput.n38 gnd 0.033063f
C4411 CSoutput.n39 gnd 0.040642f
C4412 CSoutput.n40 gnd 0.040642f
C4413 CSoutput.n41 gnd 0.033913f
C4414 CSoutput.n42 gnd 0.030997f
C4415 CSoutput.n43 gnd 0.12007f
C4416 CSoutput.n44 gnd 0.031783f
C4417 CSoutput.n45 gnd 0.040642f
C4418 CSoutput.n46 gnd 0.040642f
C4419 CSoutput.n47 gnd 0.040642f
C4420 CSoutput.n48 gnd 0.031783f
C4421 CSoutput.n49 gnd 0.12007f
C4422 CSoutput.n50 gnd 0.030997f
C4423 CSoutput.n51 gnd 0.033913f
C4424 CSoutput.n52 gnd 0.040642f
C4425 CSoutput.n53 gnd 0.040642f
C4426 CSoutput.n54 gnd 0.033063f
C4427 CSoutput.n55 gnd 0.031847f
C4428 CSoutput.n56 gnd 0.12007f
C4429 CSoutput.n57 gnd 0.033301f
C4430 CSoutput.n58 gnd 0.040642f
C4431 CSoutput.n59 gnd 0.040642f
C4432 CSoutput.n60 gnd 0.040642f
C4433 CSoutput.n61 gnd 0.028971f
C4434 CSoutput.n62 gnd 0.122743f
C4435 CSoutput.n63 gnd 0.028578f
C4436 CSoutput.t140 gnd 0.268837f
C4437 CSoutput.n64 gnd 0.12007f
C4438 CSoutput.n65 gnd 0.033659f
C4439 CSoutput.n66 gnd 0.040642f
C4440 CSoutput.n67 gnd 0.040642f
C4441 CSoutput.n68 gnd 0.040642f
C4442 CSoutput.n69 gnd 0.032698f
C4443 CSoutput.n70 gnd 0.12007f
C4444 CSoutput.n71 gnd 0.03392f
C4445 CSoutput.n72 gnd 0.029667f
C4446 CSoutput.n73 gnd 0.040642f
C4447 CSoutput.n74 gnd 0.040642f
C4448 CSoutput.n75 gnd 0.030767f
C4449 CSoutput.n76 gnd 0.018272f
C4450 CSoutput.t120 gnd 0.302058f
C4451 CSoutput.n77 gnd 0.15005f
C4452 CSoutput.n78 gnd 0.642051f
C4453 CSoutput.t115 gnd 0.050695f
C4454 CSoutput.t77 gnd 0.050695f
C4455 CSoutput.n79 gnd 0.392498f
C4456 CSoutput.t59 gnd 0.050695f
C4457 CSoutput.t116 gnd 0.050695f
C4458 CSoutput.n80 gnd 0.391798f
C4459 CSoutput.n81 gnd 0.397674f
C4460 CSoutput.t60 gnd 0.050695f
C4461 CSoutput.t94 gnd 0.050695f
C4462 CSoutput.n82 gnd 0.391798f
C4463 CSoutput.n83 gnd 0.195957f
C4464 CSoutput.t73 gnd 0.050695f
C4465 CSoutput.t98 gnd 0.050695f
C4466 CSoutput.n84 gnd 0.391798f
C4467 CSoutput.n85 gnd 0.195957f
C4468 CSoutput.t89 gnd 0.050695f
C4469 CSoutput.t71 gnd 0.050695f
C4470 CSoutput.n86 gnd 0.391798f
C4471 CSoutput.n87 gnd 0.195957f
C4472 CSoutput.t119 gnd 0.050695f
C4473 CSoutput.t81 gnd 0.050695f
C4474 CSoutput.n88 gnd 0.391798f
C4475 CSoutput.n89 gnd 0.35934f
C4476 CSoutput.t63 gnd 0.050695f
C4477 CSoutput.t109 gnd 0.050695f
C4478 CSoutput.n90 gnd 0.392498f
C4479 CSoutput.t84 gnd 0.050695f
C4480 CSoutput.t51 gnd 0.050695f
C4481 CSoutput.n91 gnd 0.391798f
C4482 CSoutput.n92 gnd 0.397674f
C4483 CSoutput.t1 gnd 0.050695f
C4484 CSoutput.t61 gnd 0.050695f
C4485 CSoutput.n93 gnd 0.391798f
C4486 CSoutput.n94 gnd 0.195957f
C4487 CSoutput.t85 gnd 0.050695f
C4488 CSoutput.t57 gnd 0.050695f
C4489 CSoutput.n95 gnd 0.391798f
C4490 CSoutput.n96 gnd 0.195957f
C4491 CSoutput.t64 gnd 0.050695f
C4492 CSoutput.t111 gnd 0.050695f
C4493 CSoutput.n97 gnd 0.391798f
C4494 CSoutput.n98 gnd 0.195957f
C4495 CSoutput.t102 gnd 0.050695f
C4496 CSoutput.t103 gnd 0.050695f
C4497 CSoutput.n99 gnd 0.391798f
C4498 CSoutput.n100 gnd 0.292221f
C4499 CSoutput.n101 gnd 0.368489f
C4500 CSoutput.t53 gnd 0.050695f
C4501 CSoutput.t52 gnd 0.050695f
C4502 CSoutput.n102 gnd 0.392498f
C4503 CSoutput.t106 gnd 0.050695f
C4504 CSoutput.t95 gnd 0.050695f
C4505 CSoutput.n103 gnd 0.391798f
C4506 CSoutput.n104 gnd 0.397674f
C4507 CSoutput.t55 gnd 0.050695f
C4508 CSoutput.t110 gnd 0.050695f
C4509 CSoutput.n105 gnd 0.391798f
C4510 CSoutput.n106 gnd 0.195957f
C4511 CSoutput.t107 gnd 0.050695f
C4512 CSoutput.t100 gnd 0.050695f
C4513 CSoutput.n107 gnd 0.391798f
C4514 CSoutput.n108 gnd 0.195957f
C4515 CSoutput.t97 gnd 0.050695f
C4516 CSoutput.t87 gnd 0.050695f
C4517 CSoutput.n109 gnd 0.391798f
C4518 CSoutput.n110 gnd 0.195957f
C4519 CSoutput.t90 gnd 0.050695f
C4520 CSoutput.t91 gnd 0.050695f
C4521 CSoutput.n111 gnd 0.391798f
C4522 CSoutput.n112 gnd 0.292221f
C4523 CSoutput.n113 gnd 0.411877f
C4524 CSoutput.n114 gnd 6.98446f
C4525 CSoutput.n116 gnd 0.718948f
C4526 CSoutput.n117 gnd 0.539211f
C4527 CSoutput.n118 gnd 0.718948f
C4528 CSoutput.n119 gnd 0.718948f
C4529 CSoutput.n120 gnd 1.93563f
C4530 CSoutput.n121 gnd 0.718948f
C4531 CSoutput.n122 gnd 0.718948f
C4532 CSoutput.t139 gnd 0.898685f
C4533 CSoutput.n123 gnd 0.718948f
C4534 CSoutput.n124 gnd 0.718948f
C4535 CSoutput.n128 gnd 0.718948f
C4536 CSoutput.n132 gnd 0.718948f
C4537 CSoutput.n133 gnd 0.718948f
C4538 CSoutput.n135 gnd 0.718948f
C4539 CSoutput.n140 gnd 0.718948f
C4540 CSoutput.n142 gnd 0.718948f
C4541 CSoutput.n143 gnd 0.718948f
C4542 CSoutput.n145 gnd 0.718948f
C4543 CSoutput.n146 gnd 0.718948f
C4544 CSoutput.n148 gnd 0.718948f
C4545 CSoutput.t128 gnd 12.013499f
C4546 CSoutput.n150 gnd 0.718948f
C4547 CSoutput.n151 gnd 0.539211f
C4548 CSoutput.n152 gnd 0.718948f
C4549 CSoutput.n153 gnd 0.718948f
C4550 CSoutput.n154 gnd 1.93563f
C4551 CSoutput.n155 gnd 0.718948f
C4552 CSoutput.n156 gnd 0.718948f
C4553 CSoutput.t126 gnd 0.898685f
C4554 CSoutput.n157 gnd 0.718948f
C4555 CSoutput.n158 gnd 0.718948f
C4556 CSoutput.n162 gnd 0.718948f
C4557 CSoutput.n166 gnd 0.718948f
C4558 CSoutput.n167 gnd 0.718948f
C4559 CSoutput.n169 gnd 0.718948f
C4560 CSoutput.n174 gnd 0.718948f
C4561 CSoutput.n176 gnd 0.718948f
C4562 CSoutput.n177 gnd 0.718948f
C4563 CSoutput.n179 gnd 0.718948f
C4564 CSoutput.n180 gnd 0.718948f
C4565 CSoutput.n182 gnd 0.718948f
C4566 CSoutput.n183 gnd 0.539211f
C4567 CSoutput.n185 gnd 0.718948f
C4568 CSoutput.n186 gnd 0.539211f
C4569 CSoutput.n187 gnd 0.718948f
C4570 CSoutput.n188 gnd 0.718948f
C4571 CSoutput.n189 gnd 1.93563f
C4572 CSoutput.n190 gnd 0.718948f
C4573 CSoutput.n191 gnd 0.718948f
C4574 CSoutput.t122 gnd 0.898685f
C4575 CSoutput.n192 gnd 0.718948f
C4576 CSoutput.n193 gnd 1.93563f
C4577 CSoutput.n195 gnd 0.718948f
C4578 CSoutput.n196 gnd 0.718948f
C4579 CSoutput.n198 gnd 0.718948f
C4580 CSoutput.n199 gnd 0.718948f
C4581 CSoutput.t129 gnd 11.8178f
C4582 CSoutput.t133 gnd 12.013499f
C4583 CSoutput.n205 gnd 2.25544f
C4584 CSoutput.n206 gnd 9.18786f
C4585 CSoutput.n207 gnd 9.57232f
C4586 CSoutput.n212 gnd 2.44325f
C4587 CSoutput.n218 gnd 0.718948f
C4588 CSoutput.n220 gnd 0.718948f
C4589 CSoutput.n222 gnd 0.718948f
C4590 CSoutput.n224 gnd 0.718948f
C4591 CSoutput.n226 gnd 0.718948f
C4592 CSoutput.n232 gnd 0.718948f
C4593 CSoutput.n239 gnd 1.31899f
C4594 CSoutput.n240 gnd 1.31899f
C4595 CSoutput.n241 gnd 0.718948f
C4596 CSoutput.n242 gnd 0.718948f
C4597 CSoutput.n244 gnd 0.539211f
C4598 CSoutput.n245 gnd 0.461786f
C4599 CSoutput.n247 gnd 0.539211f
C4600 CSoutput.n248 gnd 0.461786f
C4601 CSoutput.n249 gnd 0.539211f
C4602 CSoutput.n251 gnd 0.718948f
C4603 CSoutput.n253 gnd 1.93563f
C4604 CSoutput.n254 gnd 2.25544f
C4605 CSoutput.n255 gnd 8.45047f
C4606 CSoutput.n257 gnd 0.539211f
C4607 CSoutput.n258 gnd 1.38742f
C4608 CSoutput.n259 gnd 0.539211f
C4609 CSoutput.n261 gnd 0.718948f
C4610 CSoutput.n263 gnd 1.93563f
C4611 CSoutput.n264 gnd 4.21611f
C4612 CSoutput.t76 gnd 0.050695f
C4613 CSoutput.t62 gnd 0.050695f
C4614 CSoutput.n265 gnd 0.392498f
C4615 CSoutput.t113 gnd 0.050695f
C4616 CSoutput.t74 gnd 0.050695f
C4617 CSoutput.n266 gnd 0.391798f
C4618 CSoutput.n267 gnd 0.397674f
C4619 CSoutput.t65 gnd 0.050695f
C4620 CSoutput.t92 gnd 0.050695f
C4621 CSoutput.n268 gnd 0.391798f
C4622 CSoutput.n269 gnd 0.195957f
C4623 CSoutput.t69 gnd 0.050695f
C4624 CSoutput.t72 gnd 0.050695f
C4625 CSoutput.n270 gnd 0.391798f
C4626 CSoutput.n271 gnd 0.195957f
C4627 CSoutput.t58 gnd 0.050695f
C4628 CSoutput.t88 gnd 0.050695f
C4629 CSoutput.n272 gnd 0.391798f
C4630 CSoutput.n273 gnd 0.195957f
C4631 CSoutput.t80 gnd 0.050695f
C4632 CSoutput.t50 gnd 0.050695f
C4633 CSoutput.n274 gnd 0.391798f
C4634 CSoutput.n275 gnd 0.35934f
C4635 CSoutput.t112 gnd 0.050695f
C4636 CSoutput.t101 gnd 0.050695f
C4637 CSoutput.n276 gnd 0.392498f
C4638 CSoutput.t104 gnd 0.050695f
C4639 CSoutput.t0 gnd 0.050695f
C4640 CSoutput.n277 gnd 0.391798f
C4641 CSoutput.n278 gnd 0.397674f
C4642 CSoutput.t117 gnd 0.050695f
C4643 CSoutput.t105 gnd 0.050695f
C4644 CSoutput.n279 gnd 0.391798f
C4645 CSoutput.n280 gnd 0.195957f
C4646 CSoutput.t86 gnd 0.050695f
C4647 CSoutput.t67 gnd 0.050695f
C4648 CSoutput.n281 gnd 0.391798f
C4649 CSoutput.n282 gnd 0.195957f
C4650 CSoutput.t66 gnd 0.050695f
C4651 CSoutput.t114 gnd 0.050695f
C4652 CSoutput.n283 gnd 0.391798f
C4653 CSoutput.n284 gnd 0.195957f
C4654 CSoutput.t79 gnd 0.050695f
C4655 CSoutput.t78 gnd 0.050695f
C4656 CSoutput.n285 gnd 0.391798f
C4657 CSoutput.n286 gnd 0.292221f
C4658 CSoutput.n287 gnd 0.368489f
C4659 CSoutput.t83 gnd 0.050695f
C4660 CSoutput.t82 gnd 0.050695f
C4661 CSoutput.n288 gnd 0.392498f
C4662 CSoutput.t108 gnd 0.050695f
C4663 CSoutput.t54 gnd 0.050695f
C4664 CSoutput.n289 gnd 0.391798f
C4665 CSoutput.n290 gnd 0.397674f
C4666 CSoutput.t70 gnd 0.050695f
C4667 CSoutput.t93 gnd 0.050695f
C4668 CSoutput.n291 gnd 0.391798f
C4669 CSoutput.n292 gnd 0.195957f
C4670 CSoutput.t118 gnd 0.050695f
C4671 CSoutput.t68 gnd 0.050695f
C4672 CSoutput.n293 gnd 0.391798f
C4673 CSoutput.n294 gnd 0.195957f
C4674 CSoutput.t56 gnd 0.050695f
C4675 CSoutput.t75 gnd 0.050695f
C4676 CSoutput.n295 gnd 0.391798f
C4677 CSoutput.n296 gnd 0.195957f
C4678 CSoutput.t96 gnd 0.050695f
C4679 CSoutput.t99 gnd 0.050695f
C4680 CSoutput.n297 gnd 0.391797f
C4681 CSoutput.n298 gnd 0.292223f
C4682 CSoutput.n299 gnd 0.411877f
C4683 CSoutput.n300 gnd 10.2443f
C4684 CSoutput.t26 gnd 0.044358f
C4685 CSoutput.t16 gnd 0.044358f
C4686 CSoutput.n301 gnd 0.393276f
C4687 CSoutput.t42 gnd 0.044358f
C4688 CSoutput.t44 gnd 0.044358f
C4689 CSoutput.n302 gnd 0.391964f
C4690 CSoutput.n303 gnd 0.365237f
C4691 CSoutput.t21 gnd 0.044358f
C4692 CSoutput.t11 gnd 0.044358f
C4693 CSoutput.n304 gnd 0.391964f
C4694 CSoutput.n305 gnd 0.180045f
C4695 CSoutput.t47 gnd 0.044358f
C4696 CSoutput.t28 gnd 0.044358f
C4697 CSoutput.n306 gnd 0.391964f
C4698 CSoutput.n307 gnd 0.180045f
C4699 CSoutput.t30 gnd 0.044358f
C4700 CSoutput.t19 gnd 0.044358f
C4701 CSoutput.n308 gnd 0.391964f
C4702 CSoutput.n309 gnd 0.180045f
C4703 CSoutput.t33 gnd 0.044358f
C4704 CSoutput.t35 gnd 0.044358f
C4705 CSoutput.n310 gnd 0.391964f
C4706 CSoutput.n311 gnd 0.332039f
C4707 CSoutput.t36 gnd 0.044358f
C4708 CSoutput.t25 gnd 0.044358f
C4709 CSoutput.n312 gnd 0.393276f
C4710 CSoutput.t48 gnd 0.044358f
C4711 CSoutput.t2 gnd 0.044358f
C4712 CSoutput.n313 gnd 0.391964f
C4713 CSoutput.n314 gnd 0.365237f
C4714 CSoutput.t31 gnd 0.044358f
C4715 CSoutput.t20 gnd 0.044358f
C4716 CSoutput.n315 gnd 0.391964f
C4717 CSoutput.n316 gnd 0.180045f
C4718 CSoutput.t6 gnd 0.044358f
C4719 CSoutput.t37 gnd 0.044358f
C4720 CSoutput.n317 gnd 0.391964f
C4721 CSoutput.n318 gnd 0.180045f
C4722 CSoutput.t39 gnd 0.044358f
C4723 CSoutput.t29 gnd 0.044358f
C4724 CSoutput.n319 gnd 0.391964f
C4725 CSoutput.n320 gnd 0.180045f
C4726 CSoutput.t40 gnd 0.044358f
C4727 CSoutput.t43 gnd 0.044358f
C4728 CSoutput.n321 gnd 0.391964f
C4729 CSoutput.n322 gnd 0.273347f
C4730 CSoutput.n323 gnd 0.507899f
C4731 CSoutput.n324 gnd 10.6628f
C4732 CSoutput.t5 gnd 0.044358f
C4733 CSoutput.t13 gnd 0.044358f
C4734 CSoutput.n325 gnd 0.393276f
C4735 CSoutput.t34 gnd 0.044358f
C4736 CSoutput.t46 gnd 0.044358f
C4737 CSoutput.n326 gnd 0.391964f
C4738 CSoutput.n327 gnd 0.365237f
C4739 CSoutput.t49 gnd 0.044358f
C4740 CSoutput.t9 gnd 0.044358f
C4741 CSoutput.n328 gnd 0.391964f
C4742 CSoutput.n329 gnd 0.180045f
C4743 CSoutput.t14 gnd 0.044358f
C4744 CSoutput.t3 gnd 0.044358f
C4745 CSoutput.n330 gnd 0.391964f
C4746 CSoutput.n331 gnd 0.180045f
C4747 CSoutput.t7 gnd 0.044358f
C4748 CSoutput.t17 gnd 0.044358f
C4749 CSoutput.n332 gnd 0.391964f
C4750 CSoutput.n333 gnd 0.180045f
C4751 CSoutput.t22 gnd 0.044358f
C4752 CSoutput.t38 gnd 0.044358f
C4753 CSoutput.n334 gnd 0.391964f
C4754 CSoutput.n335 gnd 0.332039f
C4755 CSoutput.t12 gnd 0.044358f
C4756 CSoutput.t24 gnd 0.044358f
C4757 CSoutput.n336 gnd 0.393276f
C4758 CSoutput.t41 gnd 0.044358f
C4759 CSoutput.t4 gnd 0.044358f
C4760 CSoutput.n337 gnd 0.391964f
C4761 CSoutput.n338 gnd 0.365237f
C4762 CSoutput.t8 gnd 0.044358f
C4763 CSoutput.t18 gnd 0.044358f
C4764 CSoutput.n339 gnd 0.391964f
C4765 CSoutput.n340 gnd 0.180045f
C4766 CSoutput.t23 gnd 0.044358f
C4767 CSoutput.t10 gnd 0.044358f
C4768 CSoutput.n341 gnd 0.391964f
C4769 CSoutput.n342 gnd 0.180045f
C4770 CSoutput.t15 gnd 0.044358f
C4771 CSoutput.t27 gnd 0.044358f
C4772 CSoutput.n343 gnd 0.391964f
C4773 CSoutput.n344 gnd 0.180045f
C4774 CSoutput.t32 gnd 0.044358f
C4775 CSoutput.t45 gnd 0.044358f
C4776 CSoutput.n345 gnd 0.391964f
C4777 CSoutput.n346 gnd 0.273347f
C4778 CSoutput.n347 gnd 0.507899f
C4779 CSoutput.n348 gnd 5.91521f
C4780 CSoutput.n349 gnd 13.0833f
C4781 commonsourceibias.n0 gnd 0.010301f
C4782 commonsourceibias.t71 gnd 0.155981f
C4783 commonsourceibias.t81 gnd 0.144227f
C4784 commonsourceibias.n1 gnd 0.057546f
C4785 commonsourceibias.n2 gnd 0.00772f
C4786 commonsourceibias.t55 gnd 0.144227f
C4787 commonsourceibias.n3 gnd 0.006245f
C4788 commonsourceibias.n4 gnd 0.00772f
C4789 commonsourceibias.t53 gnd 0.144227f
C4790 commonsourceibias.n5 gnd 0.007453f
C4791 commonsourceibias.n6 gnd 0.00772f
C4792 commonsourceibias.t76 gnd 0.144227f
C4793 commonsourceibias.n7 gnd 0.057546f
C4794 commonsourceibias.t86 gnd 0.144227f
C4795 commonsourceibias.n8 gnd 0.006235f
C4796 commonsourceibias.n9 gnd 0.010301f
C4797 commonsourceibias.t32 gnd 0.155981f
C4798 commonsourceibias.t14 gnd 0.144227f
C4799 commonsourceibias.n10 gnd 0.057546f
C4800 commonsourceibias.n11 gnd 0.00772f
C4801 commonsourceibias.t24 gnd 0.144227f
C4802 commonsourceibias.n12 gnd 0.006245f
C4803 commonsourceibias.n13 gnd 0.00772f
C4804 commonsourceibias.t30 gnd 0.144227f
C4805 commonsourceibias.n14 gnd 0.007453f
C4806 commonsourceibias.n15 gnd 0.00772f
C4807 commonsourceibias.t20 gnd 0.144227f
C4808 commonsourceibias.n16 gnd 0.057546f
C4809 commonsourceibias.t36 gnd 0.144227f
C4810 commonsourceibias.n17 gnd 0.006235f
C4811 commonsourceibias.n18 gnd 0.00772f
C4812 commonsourceibias.t44 gnd 0.144227f
C4813 commonsourceibias.t26 gnd 0.144227f
C4814 commonsourceibias.n19 gnd 0.057546f
C4815 commonsourceibias.n20 gnd 0.00772f
C4816 commonsourceibias.t34 gnd 0.144227f
C4817 commonsourceibias.n21 gnd 0.057546f
C4818 commonsourceibias.n22 gnd 0.00772f
C4819 commonsourceibias.t10 gnd 0.144227f
C4820 commonsourceibias.n23 gnd 0.057546f
C4821 commonsourceibias.n24 gnd 0.038863f
C4822 commonsourceibias.t40 gnd 0.144227f
C4823 commonsourceibias.t46 gnd 0.162743f
C4824 commonsourceibias.n25 gnd 0.066782f
C4825 commonsourceibias.n26 gnd 0.069137f
C4826 commonsourceibias.n27 gnd 0.009515f
C4827 commonsourceibias.n28 gnd 0.010526f
C4828 commonsourceibias.n29 gnd 0.00772f
C4829 commonsourceibias.n30 gnd 0.00772f
C4830 commonsourceibias.n31 gnd 0.010457f
C4831 commonsourceibias.n32 gnd 0.006245f
C4832 commonsourceibias.n33 gnd 0.010587f
C4833 commonsourceibias.n34 gnd 0.00772f
C4834 commonsourceibias.n35 gnd 0.00772f
C4835 commonsourceibias.n36 gnd 0.010651f
C4836 commonsourceibias.n37 gnd 0.009185f
C4837 commonsourceibias.n38 gnd 0.007453f
C4838 commonsourceibias.n39 gnd 0.00772f
C4839 commonsourceibias.n40 gnd 0.00772f
C4840 commonsourceibias.n41 gnd 0.009442f
C4841 commonsourceibias.n42 gnd 0.010598f
C4842 commonsourceibias.n43 gnd 0.057546f
C4843 commonsourceibias.n44 gnd 0.010527f
C4844 commonsourceibias.n45 gnd 0.00772f
C4845 commonsourceibias.n46 gnd 0.00772f
C4846 commonsourceibias.n47 gnd 0.00772f
C4847 commonsourceibias.n48 gnd 0.010527f
C4848 commonsourceibias.n49 gnd 0.057546f
C4849 commonsourceibias.n50 gnd 0.010598f
C4850 commonsourceibias.n51 gnd 0.009442f
C4851 commonsourceibias.n52 gnd 0.00772f
C4852 commonsourceibias.n53 gnd 0.00772f
C4853 commonsourceibias.n54 gnd 0.00772f
C4854 commonsourceibias.n55 gnd 0.009185f
C4855 commonsourceibias.n56 gnd 0.010651f
C4856 commonsourceibias.n57 gnd 0.057546f
C4857 commonsourceibias.n58 gnd 0.010587f
C4858 commonsourceibias.n59 gnd 0.00772f
C4859 commonsourceibias.n60 gnd 0.00772f
C4860 commonsourceibias.n61 gnd 0.00772f
C4861 commonsourceibias.n62 gnd 0.010457f
C4862 commonsourceibias.n63 gnd 0.057546f
C4863 commonsourceibias.n64 gnd 0.010526f
C4864 commonsourceibias.n65 gnd 0.009515f
C4865 commonsourceibias.n66 gnd 0.00772f
C4866 commonsourceibias.n67 gnd 0.00772f
C4867 commonsourceibias.n68 gnd 0.007831f
C4868 commonsourceibias.n69 gnd 0.008096f
C4869 commonsourceibias.n70 gnd 0.068855f
C4870 commonsourceibias.n71 gnd 0.076384f
C4871 commonsourceibias.t33 gnd 0.016658f
C4872 commonsourceibias.t15 gnd 0.016658f
C4873 commonsourceibias.n72 gnd 0.147197f
C4874 commonsourceibias.n73 gnd 0.12719f
C4875 commonsourceibias.t25 gnd 0.016658f
C4876 commonsourceibias.t31 gnd 0.016658f
C4877 commonsourceibias.n74 gnd 0.147197f
C4878 commonsourceibias.n75 gnd 0.067614f
C4879 commonsourceibias.t21 gnd 0.016658f
C4880 commonsourceibias.t37 gnd 0.016658f
C4881 commonsourceibias.n76 gnd 0.147197f
C4882 commonsourceibias.n77 gnd 0.056488f
C4883 commonsourceibias.t41 gnd 0.016658f
C4884 commonsourceibias.t47 gnd 0.016658f
C4885 commonsourceibias.n78 gnd 0.14769f
C4886 commonsourceibias.t35 gnd 0.016658f
C4887 commonsourceibias.t11 gnd 0.016658f
C4888 commonsourceibias.n79 gnd 0.147197f
C4889 commonsourceibias.n80 gnd 0.13716f
C4890 commonsourceibias.t45 gnd 0.016658f
C4891 commonsourceibias.t27 gnd 0.016658f
C4892 commonsourceibias.n81 gnd 0.147197f
C4893 commonsourceibias.n82 gnd 0.056488f
C4894 commonsourceibias.n83 gnd 0.068401f
C4895 commonsourceibias.n84 gnd 0.00772f
C4896 commonsourceibias.t50 gnd 0.144227f
C4897 commonsourceibias.t69 gnd 0.144227f
C4898 commonsourceibias.n85 gnd 0.057546f
C4899 commonsourceibias.n86 gnd 0.00772f
C4900 commonsourceibias.t67 gnd 0.144227f
C4901 commonsourceibias.n87 gnd 0.057546f
C4902 commonsourceibias.n88 gnd 0.00772f
C4903 commonsourceibias.t78 gnd 0.144227f
C4904 commonsourceibias.n89 gnd 0.057546f
C4905 commonsourceibias.n90 gnd 0.038863f
C4906 commonsourceibias.t64 gnd 0.144227f
C4907 commonsourceibias.t62 gnd 0.162743f
C4908 commonsourceibias.n91 gnd 0.066782f
C4909 commonsourceibias.n92 gnd 0.069137f
C4910 commonsourceibias.n93 gnd 0.009515f
C4911 commonsourceibias.n94 gnd 0.010526f
C4912 commonsourceibias.n95 gnd 0.00772f
C4913 commonsourceibias.n96 gnd 0.00772f
C4914 commonsourceibias.n97 gnd 0.010457f
C4915 commonsourceibias.n98 gnd 0.006245f
C4916 commonsourceibias.n99 gnd 0.010587f
C4917 commonsourceibias.n100 gnd 0.00772f
C4918 commonsourceibias.n101 gnd 0.00772f
C4919 commonsourceibias.n102 gnd 0.010651f
C4920 commonsourceibias.n103 gnd 0.009185f
C4921 commonsourceibias.n104 gnd 0.007453f
C4922 commonsourceibias.n105 gnd 0.00772f
C4923 commonsourceibias.n106 gnd 0.00772f
C4924 commonsourceibias.n107 gnd 0.009442f
C4925 commonsourceibias.n108 gnd 0.010598f
C4926 commonsourceibias.n109 gnd 0.057546f
C4927 commonsourceibias.n110 gnd 0.010527f
C4928 commonsourceibias.n111 gnd 0.007683f
C4929 commonsourceibias.n112 gnd 0.055804f
C4930 commonsourceibias.n113 gnd 0.007683f
C4931 commonsourceibias.n114 gnd 0.010527f
C4932 commonsourceibias.n115 gnd 0.057546f
C4933 commonsourceibias.n116 gnd 0.010598f
C4934 commonsourceibias.n117 gnd 0.009442f
C4935 commonsourceibias.n118 gnd 0.00772f
C4936 commonsourceibias.n119 gnd 0.00772f
C4937 commonsourceibias.n120 gnd 0.00772f
C4938 commonsourceibias.n121 gnd 0.009185f
C4939 commonsourceibias.n122 gnd 0.010651f
C4940 commonsourceibias.n123 gnd 0.057546f
C4941 commonsourceibias.n124 gnd 0.010587f
C4942 commonsourceibias.n125 gnd 0.00772f
C4943 commonsourceibias.n126 gnd 0.00772f
C4944 commonsourceibias.n127 gnd 0.00772f
C4945 commonsourceibias.n128 gnd 0.010457f
C4946 commonsourceibias.n129 gnd 0.057546f
C4947 commonsourceibias.n130 gnd 0.010526f
C4948 commonsourceibias.n131 gnd 0.009515f
C4949 commonsourceibias.n132 gnd 0.00772f
C4950 commonsourceibias.n133 gnd 0.00772f
C4951 commonsourceibias.n134 gnd 0.007831f
C4952 commonsourceibias.n135 gnd 0.008096f
C4953 commonsourceibias.n136 gnd 0.068855f
C4954 commonsourceibias.n137 gnd 0.04456f
C4955 commonsourceibias.n138 gnd 0.010301f
C4956 commonsourceibias.t72 gnd 0.144227f
C4957 commonsourceibias.n139 gnd 0.057546f
C4958 commonsourceibias.n140 gnd 0.00772f
C4959 commonsourceibias.t49 gnd 0.144227f
C4960 commonsourceibias.n141 gnd 0.006245f
C4961 commonsourceibias.n142 gnd 0.00772f
C4962 commonsourceibias.t95 gnd 0.144227f
C4963 commonsourceibias.n143 gnd 0.007453f
C4964 commonsourceibias.n144 gnd 0.00772f
C4965 commonsourceibias.t66 gnd 0.144227f
C4966 commonsourceibias.n145 gnd 0.057546f
C4967 commonsourceibias.t77 gnd 0.144227f
C4968 commonsourceibias.n146 gnd 0.006235f
C4969 commonsourceibias.n147 gnd 0.00772f
C4970 commonsourceibias.t91 gnd 0.144227f
C4971 commonsourceibias.t60 gnd 0.144227f
C4972 commonsourceibias.n148 gnd 0.057546f
C4973 commonsourceibias.n149 gnd 0.00772f
C4974 commonsourceibias.t58 gnd 0.144227f
C4975 commonsourceibias.n150 gnd 0.057546f
C4976 commonsourceibias.n151 gnd 0.00772f
C4977 commonsourceibias.t68 gnd 0.144227f
C4978 commonsourceibias.n152 gnd 0.057546f
C4979 commonsourceibias.n153 gnd 0.038863f
C4980 commonsourceibias.t57 gnd 0.144227f
C4981 commonsourceibias.t54 gnd 0.162743f
C4982 commonsourceibias.n154 gnd 0.066782f
C4983 commonsourceibias.n155 gnd 0.069137f
C4984 commonsourceibias.n156 gnd 0.009515f
C4985 commonsourceibias.n157 gnd 0.010526f
C4986 commonsourceibias.n158 gnd 0.00772f
C4987 commonsourceibias.n159 gnd 0.00772f
C4988 commonsourceibias.n160 gnd 0.010457f
C4989 commonsourceibias.n161 gnd 0.006245f
C4990 commonsourceibias.n162 gnd 0.010587f
C4991 commonsourceibias.n163 gnd 0.00772f
C4992 commonsourceibias.n164 gnd 0.00772f
C4993 commonsourceibias.n165 gnd 0.010651f
C4994 commonsourceibias.n166 gnd 0.009185f
C4995 commonsourceibias.n167 gnd 0.007453f
C4996 commonsourceibias.n168 gnd 0.00772f
C4997 commonsourceibias.n169 gnd 0.00772f
C4998 commonsourceibias.n170 gnd 0.009442f
C4999 commonsourceibias.n171 gnd 0.010598f
C5000 commonsourceibias.n172 gnd 0.057546f
C5001 commonsourceibias.n173 gnd 0.010527f
C5002 commonsourceibias.n174 gnd 0.00772f
C5003 commonsourceibias.n175 gnd 0.00772f
C5004 commonsourceibias.n176 gnd 0.00772f
C5005 commonsourceibias.n177 gnd 0.010527f
C5006 commonsourceibias.n178 gnd 0.057546f
C5007 commonsourceibias.n179 gnd 0.010598f
C5008 commonsourceibias.n180 gnd 0.009442f
C5009 commonsourceibias.n181 gnd 0.00772f
C5010 commonsourceibias.n182 gnd 0.00772f
C5011 commonsourceibias.n183 gnd 0.00772f
C5012 commonsourceibias.n184 gnd 0.009185f
C5013 commonsourceibias.n185 gnd 0.010651f
C5014 commonsourceibias.n186 gnd 0.057546f
C5015 commonsourceibias.n187 gnd 0.010587f
C5016 commonsourceibias.n188 gnd 0.00772f
C5017 commonsourceibias.n189 gnd 0.00772f
C5018 commonsourceibias.n190 gnd 0.00772f
C5019 commonsourceibias.n191 gnd 0.010457f
C5020 commonsourceibias.n192 gnd 0.057546f
C5021 commonsourceibias.n193 gnd 0.010526f
C5022 commonsourceibias.n194 gnd 0.009515f
C5023 commonsourceibias.n195 gnd 0.00772f
C5024 commonsourceibias.n196 gnd 0.00772f
C5025 commonsourceibias.n197 gnd 0.007831f
C5026 commonsourceibias.n198 gnd 0.008096f
C5027 commonsourceibias.t61 gnd 0.155981f
C5028 commonsourceibias.n199 gnd 0.068855f
C5029 commonsourceibias.n200 gnd 0.023432f
C5030 commonsourceibias.n201 gnd 0.388694f
C5031 commonsourceibias.n202 gnd 0.010301f
C5032 commonsourceibias.t84 gnd 0.155981f
C5033 commonsourceibias.t92 gnd 0.144227f
C5034 commonsourceibias.n203 gnd 0.057546f
C5035 commonsourceibias.n204 gnd 0.00772f
C5036 commonsourceibias.t51 gnd 0.144227f
C5037 commonsourceibias.n205 gnd 0.006245f
C5038 commonsourceibias.n206 gnd 0.00772f
C5039 commonsourceibias.t63 gnd 0.144227f
C5040 commonsourceibias.n207 gnd 0.007453f
C5041 commonsourceibias.n208 gnd 0.00772f
C5042 commonsourceibias.t48 gnd 0.144227f
C5043 commonsourceibias.n209 gnd 0.006235f
C5044 commonsourceibias.n210 gnd 0.00772f
C5045 commonsourceibias.t94 gnd 0.144227f
C5046 commonsourceibias.t83 gnd 0.144227f
C5047 commonsourceibias.n211 gnd 0.057546f
C5048 commonsourceibias.n212 gnd 0.00772f
C5049 commonsourceibias.t80 gnd 0.144227f
C5050 commonsourceibias.n213 gnd 0.057546f
C5051 commonsourceibias.n214 gnd 0.00772f
C5052 commonsourceibias.t90 gnd 0.144227f
C5053 commonsourceibias.n215 gnd 0.057546f
C5054 commonsourceibias.n216 gnd 0.038863f
C5055 commonsourceibias.t59 gnd 0.144227f
C5056 commonsourceibias.t75 gnd 0.162743f
C5057 commonsourceibias.n217 gnd 0.066782f
C5058 commonsourceibias.n218 gnd 0.069137f
C5059 commonsourceibias.n219 gnd 0.009515f
C5060 commonsourceibias.n220 gnd 0.010526f
C5061 commonsourceibias.n221 gnd 0.00772f
C5062 commonsourceibias.n222 gnd 0.00772f
C5063 commonsourceibias.n223 gnd 0.010457f
C5064 commonsourceibias.n224 gnd 0.006245f
C5065 commonsourceibias.n225 gnd 0.010587f
C5066 commonsourceibias.n226 gnd 0.00772f
C5067 commonsourceibias.n227 gnd 0.00772f
C5068 commonsourceibias.n228 gnd 0.010651f
C5069 commonsourceibias.n229 gnd 0.009185f
C5070 commonsourceibias.n230 gnd 0.007453f
C5071 commonsourceibias.n231 gnd 0.00772f
C5072 commonsourceibias.n232 gnd 0.00772f
C5073 commonsourceibias.n233 gnd 0.009442f
C5074 commonsourceibias.n234 gnd 0.010598f
C5075 commonsourceibias.n235 gnd 0.057546f
C5076 commonsourceibias.n236 gnd 0.010527f
C5077 commonsourceibias.n237 gnd 0.007683f
C5078 commonsourceibias.t17 gnd 0.016658f
C5079 commonsourceibias.t9 gnd 0.016658f
C5080 commonsourceibias.n238 gnd 0.14769f
C5081 commonsourceibias.t19 gnd 0.016658f
C5082 commonsourceibias.t5 gnd 0.016658f
C5083 commonsourceibias.n239 gnd 0.147197f
C5084 commonsourceibias.n240 gnd 0.13716f
C5085 commonsourceibias.t43 gnd 0.016658f
C5086 commonsourceibias.t13 gnd 0.016658f
C5087 commonsourceibias.n241 gnd 0.147197f
C5088 commonsourceibias.n242 gnd 0.056488f
C5089 commonsourceibias.n243 gnd 0.010301f
C5090 commonsourceibias.t22 gnd 0.144227f
C5091 commonsourceibias.n244 gnd 0.057546f
C5092 commonsourceibias.n245 gnd 0.00772f
C5093 commonsourceibias.t38 gnd 0.144227f
C5094 commonsourceibias.n246 gnd 0.006245f
C5095 commonsourceibias.n247 gnd 0.00772f
C5096 commonsourceibias.t0 gnd 0.144227f
C5097 commonsourceibias.n248 gnd 0.007453f
C5098 commonsourceibias.n249 gnd 0.00772f
C5099 commonsourceibias.t6 gnd 0.144227f
C5100 commonsourceibias.n250 gnd 0.006235f
C5101 commonsourceibias.n251 gnd 0.00772f
C5102 commonsourceibias.t12 gnd 0.144227f
C5103 commonsourceibias.t42 gnd 0.144227f
C5104 commonsourceibias.n252 gnd 0.057546f
C5105 commonsourceibias.n253 gnd 0.00772f
C5106 commonsourceibias.t4 gnd 0.144227f
C5107 commonsourceibias.n254 gnd 0.057546f
C5108 commonsourceibias.n255 gnd 0.00772f
C5109 commonsourceibias.t18 gnd 0.144227f
C5110 commonsourceibias.n256 gnd 0.057546f
C5111 commonsourceibias.n257 gnd 0.038863f
C5112 commonsourceibias.t8 gnd 0.144227f
C5113 commonsourceibias.t16 gnd 0.162743f
C5114 commonsourceibias.n258 gnd 0.066782f
C5115 commonsourceibias.n259 gnd 0.069137f
C5116 commonsourceibias.n260 gnd 0.009515f
C5117 commonsourceibias.n261 gnd 0.010526f
C5118 commonsourceibias.n262 gnd 0.00772f
C5119 commonsourceibias.n263 gnd 0.00772f
C5120 commonsourceibias.n264 gnd 0.010457f
C5121 commonsourceibias.n265 gnd 0.006245f
C5122 commonsourceibias.n266 gnd 0.010587f
C5123 commonsourceibias.n267 gnd 0.00772f
C5124 commonsourceibias.n268 gnd 0.00772f
C5125 commonsourceibias.n269 gnd 0.010651f
C5126 commonsourceibias.n270 gnd 0.009185f
C5127 commonsourceibias.n271 gnd 0.007453f
C5128 commonsourceibias.n272 gnd 0.00772f
C5129 commonsourceibias.n273 gnd 0.00772f
C5130 commonsourceibias.n274 gnd 0.009442f
C5131 commonsourceibias.n275 gnd 0.010598f
C5132 commonsourceibias.n276 gnd 0.057546f
C5133 commonsourceibias.n277 gnd 0.010527f
C5134 commonsourceibias.n278 gnd 0.00772f
C5135 commonsourceibias.n279 gnd 0.00772f
C5136 commonsourceibias.n280 gnd 0.00772f
C5137 commonsourceibias.n281 gnd 0.010527f
C5138 commonsourceibias.n282 gnd 0.057546f
C5139 commonsourceibias.n283 gnd 0.010598f
C5140 commonsourceibias.t28 gnd 0.144227f
C5141 commonsourceibias.n284 gnd 0.057546f
C5142 commonsourceibias.n285 gnd 0.009442f
C5143 commonsourceibias.n286 gnd 0.00772f
C5144 commonsourceibias.n287 gnd 0.00772f
C5145 commonsourceibias.n288 gnd 0.00772f
C5146 commonsourceibias.n289 gnd 0.009185f
C5147 commonsourceibias.n290 gnd 0.010651f
C5148 commonsourceibias.n291 gnd 0.057546f
C5149 commonsourceibias.n292 gnd 0.010587f
C5150 commonsourceibias.n293 gnd 0.00772f
C5151 commonsourceibias.n294 gnd 0.00772f
C5152 commonsourceibias.n295 gnd 0.00772f
C5153 commonsourceibias.n296 gnd 0.010457f
C5154 commonsourceibias.n297 gnd 0.057546f
C5155 commonsourceibias.n298 gnd 0.010526f
C5156 commonsourceibias.n299 gnd 0.009515f
C5157 commonsourceibias.n300 gnd 0.00772f
C5158 commonsourceibias.n301 gnd 0.00772f
C5159 commonsourceibias.n302 gnd 0.007831f
C5160 commonsourceibias.n303 gnd 0.008096f
C5161 commonsourceibias.t2 gnd 0.155981f
C5162 commonsourceibias.n304 gnd 0.068855f
C5163 commonsourceibias.n305 gnd 0.076384f
C5164 commonsourceibias.t23 gnd 0.016658f
C5165 commonsourceibias.t3 gnd 0.016658f
C5166 commonsourceibias.n306 gnd 0.147197f
C5167 commonsourceibias.n307 gnd 0.12719f
C5168 commonsourceibias.t1 gnd 0.016658f
C5169 commonsourceibias.t39 gnd 0.016658f
C5170 commonsourceibias.n308 gnd 0.147197f
C5171 commonsourceibias.n309 gnd 0.067614f
C5172 commonsourceibias.t7 gnd 0.016658f
C5173 commonsourceibias.t29 gnd 0.016658f
C5174 commonsourceibias.n310 gnd 0.147197f
C5175 commonsourceibias.n311 gnd 0.056488f
C5176 commonsourceibias.n312 gnd 0.068401f
C5177 commonsourceibias.n313 gnd 0.055804f
C5178 commonsourceibias.n314 gnd 0.007683f
C5179 commonsourceibias.n315 gnd 0.010527f
C5180 commonsourceibias.n316 gnd 0.057546f
C5181 commonsourceibias.n317 gnd 0.010598f
C5182 commonsourceibias.t88 gnd 0.144227f
C5183 commonsourceibias.n318 gnd 0.057546f
C5184 commonsourceibias.n319 gnd 0.009442f
C5185 commonsourceibias.n320 gnd 0.00772f
C5186 commonsourceibias.n321 gnd 0.00772f
C5187 commonsourceibias.n322 gnd 0.00772f
C5188 commonsourceibias.n323 gnd 0.009185f
C5189 commonsourceibias.n324 gnd 0.010651f
C5190 commonsourceibias.n325 gnd 0.057546f
C5191 commonsourceibias.n326 gnd 0.010587f
C5192 commonsourceibias.n327 gnd 0.00772f
C5193 commonsourceibias.n328 gnd 0.00772f
C5194 commonsourceibias.n329 gnd 0.00772f
C5195 commonsourceibias.n330 gnd 0.010457f
C5196 commonsourceibias.n331 gnd 0.057546f
C5197 commonsourceibias.n332 gnd 0.010526f
C5198 commonsourceibias.n333 gnd 0.009515f
C5199 commonsourceibias.n334 gnd 0.00772f
C5200 commonsourceibias.n335 gnd 0.00772f
C5201 commonsourceibias.n336 gnd 0.007831f
C5202 commonsourceibias.n337 gnd 0.008096f
C5203 commonsourceibias.n338 gnd 0.068855f
C5204 commonsourceibias.n339 gnd 0.04456f
C5205 commonsourceibias.n340 gnd 0.010301f
C5206 commonsourceibias.t85 gnd 0.144227f
C5207 commonsourceibias.n341 gnd 0.057546f
C5208 commonsourceibias.n342 gnd 0.00772f
C5209 commonsourceibias.t93 gnd 0.144227f
C5210 commonsourceibias.n343 gnd 0.006245f
C5211 commonsourceibias.n344 gnd 0.00772f
C5212 commonsourceibias.t56 gnd 0.144227f
C5213 commonsourceibias.n345 gnd 0.007453f
C5214 commonsourceibias.n346 gnd 0.00772f
C5215 commonsourceibias.t89 gnd 0.144227f
C5216 commonsourceibias.n347 gnd 0.006235f
C5217 commonsourceibias.n348 gnd 0.00772f
C5218 commonsourceibias.t87 gnd 0.144227f
C5219 commonsourceibias.t74 gnd 0.144227f
C5220 commonsourceibias.n349 gnd 0.057546f
C5221 commonsourceibias.n350 gnd 0.00772f
C5222 commonsourceibias.t70 gnd 0.144227f
C5223 commonsourceibias.n351 gnd 0.057546f
C5224 commonsourceibias.n352 gnd 0.00772f
C5225 commonsourceibias.t82 gnd 0.144227f
C5226 commonsourceibias.n353 gnd 0.057546f
C5227 commonsourceibias.n354 gnd 0.038863f
C5228 commonsourceibias.t52 gnd 0.144227f
C5229 commonsourceibias.t65 gnd 0.162743f
C5230 commonsourceibias.n355 gnd 0.066782f
C5231 commonsourceibias.n356 gnd 0.069137f
C5232 commonsourceibias.n357 gnd 0.009515f
C5233 commonsourceibias.n358 gnd 0.010526f
C5234 commonsourceibias.n359 gnd 0.00772f
C5235 commonsourceibias.n360 gnd 0.00772f
C5236 commonsourceibias.n361 gnd 0.010457f
C5237 commonsourceibias.n362 gnd 0.006245f
C5238 commonsourceibias.n363 gnd 0.010587f
C5239 commonsourceibias.n364 gnd 0.00772f
C5240 commonsourceibias.n365 gnd 0.00772f
C5241 commonsourceibias.n366 gnd 0.010651f
C5242 commonsourceibias.n367 gnd 0.009185f
C5243 commonsourceibias.n368 gnd 0.007453f
C5244 commonsourceibias.n369 gnd 0.00772f
C5245 commonsourceibias.n370 gnd 0.00772f
C5246 commonsourceibias.n371 gnd 0.009442f
C5247 commonsourceibias.n372 gnd 0.010598f
C5248 commonsourceibias.n373 gnd 0.057546f
C5249 commonsourceibias.n374 gnd 0.010527f
C5250 commonsourceibias.n375 gnd 0.00772f
C5251 commonsourceibias.n376 gnd 0.00772f
C5252 commonsourceibias.n377 gnd 0.00772f
C5253 commonsourceibias.n378 gnd 0.010527f
C5254 commonsourceibias.n379 gnd 0.057546f
C5255 commonsourceibias.n380 gnd 0.010598f
C5256 commonsourceibias.t79 gnd 0.144227f
C5257 commonsourceibias.n381 gnd 0.057546f
C5258 commonsourceibias.n382 gnd 0.009442f
C5259 commonsourceibias.n383 gnd 0.00772f
C5260 commonsourceibias.n384 gnd 0.00772f
C5261 commonsourceibias.n385 gnd 0.00772f
C5262 commonsourceibias.n386 gnd 0.009185f
C5263 commonsourceibias.n387 gnd 0.010651f
C5264 commonsourceibias.n388 gnd 0.057546f
C5265 commonsourceibias.n389 gnd 0.010587f
C5266 commonsourceibias.n390 gnd 0.00772f
C5267 commonsourceibias.n391 gnd 0.00772f
C5268 commonsourceibias.n392 gnd 0.00772f
C5269 commonsourceibias.n393 gnd 0.010457f
C5270 commonsourceibias.n394 gnd 0.057546f
C5271 commonsourceibias.n395 gnd 0.010526f
C5272 commonsourceibias.n396 gnd 0.009515f
C5273 commonsourceibias.n397 gnd 0.00772f
C5274 commonsourceibias.n398 gnd 0.00772f
C5275 commonsourceibias.n399 gnd 0.007831f
C5276 commonsourceibias.n400 gnd 0.008096f
C5277 commonsourceibias.t73 gnd 0.155981f
C5278 commonsourceibias.n401 gnd 0.068855f
C5279 commonsourceibias.n402 gnd 0.023432f
C5280 commonsourceibias.n403 gnd 0.212991f
C5281 commonsourceibias.n404 gnd 4.01312f
.ends

