* NGSPICE file created from opamp61.ext - technology: sky130A

.subckt opamp61 gnd CSoutput output vdd plus minus commonsourceibias outputibias diffpairibias
X0 a_n8300_8799.t37 plus.t5 a_n2903_n3924.t28 gnd.t316 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.7
X1 CSoutput.t95 commonsourceibias.t64 gnd.t30 gnd.t29 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X2 a_n2804_13878.t7 a_n2982_13878.t64 vdd.t131 vdd.t130 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X3 a_n2804_13878.t31 a_n2982_13878.t55 a_n2982_13878.t56 vdd.t118 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X4 CSoutput.t168 a_n2982_8322.t37 sky130_fd_pr__cap_mim_m3_1 l=12 w=12
X5 vdd.t243 a_n8300_8799.t40 CSoutput.t134 vdd.t207 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X6 gnd.t199 commonsourceibias.t65 CSoutput.t94 gnd.t12 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X7 CSoutput.t93 commonsourceibias.t66 gnd.t70 gnd.t69 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X8 CSoutput.t92 commonsourceibias.t67 gnd.t282 gnd.t44 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X9 CSoutput.t133 a_n8300_8799.t41 vdd.t242 vdd.t160 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=3.12 ps=16.78 w=8 l=0.5
X10 a_n2903_n3924.t36 plus.t6 a_n8300_8799.t36 gnd.t315 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.7
X11 plus.t3 gnd.t194 gnd.t196 gnd.t195 sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.5
X12 a_n2982_8322.t31 a_n2982_13878.t65 a_n8300_8799.t7 vdd.t128 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X13 vdd.t135 CSoutput.t169 output.t18 gnd.t318 sky130_fd_pr__nfet_01v8 ad=0.825 pd=5.33 as=0.825 ps=5.33 w=5 l=1
X14 CSoutput.t162 a_n8300_8799.t42 vdd.t241 vdd.t180 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X15 CSoutput.t91 commonsourceibias.t68 gnd.t251 gnd.t18 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X16 gnd.t284 commonsourceibias.t69 CSoutput.t90 gnd.t6 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X17 CSoutput.t89 commonsourceibias.t70 gnd.t275 gnd.t233 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X18 gnd.t220 commonsourceibias.t71 CSoutput.t88 gnd.t16 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=1.155 ps=7.33 w=7 l=1
X19 vdd.t240 a_n8300_8799.t43 CSoutput.t161 vdd.t200 sky130_fd_pr__pfet_01v8 ad=3.12 pd=16.78 as=1.32 ps=8.33 w=8 l=0.5
X20 CSoutput.t87 commonsourceibias.t72 gnd.t240 gnd.t233 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X21 CSoutput.t86 commonsourceibias.t73 gnd.t64 gnd.t63 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X22 gnd.t261 commonsourceibias.t74 CSoutput.t85 gnd.t53 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=1.155 ps=7.33 w=7 l=1
X23 commonsourceibias.t63 commonsourceibias.t62 gnd.t198 gnd.t18 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X24 CSoutput.t84 commonsourceibias.t75 gnd.t202 gnd.t44 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X25 a_n8300_8799.t38 a_n2982_13878.t66 a_n2982_8322.t30 vdd.t114 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X26 vdd.t239 a_n8300_8799.t44 CSoutput.t160 vdd.t152 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X27 a_n2982_13878.t4 minus.t5 a_n2903_n3924.t6 gnd.t37 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.7
X28 vdd.t238 a_n8300_8799.t45 CSoutput.t122 vdd.t216 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X29 CSoutput.t170 a_n2982_8322.t36 sky130_fd_pr__cap_mim_m3_1 l=12 w=12
X30 a_n8300_8799.t12 a_n2982_13878.t67 a_n2982_8322.t29 vdd.t77 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=3.51 ps=18.78 w=9 l=0.5
X31 CSoutput.t83 commonsourceibias.t76 gnd.t254 gnd.t29 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X32 gnd.t204 commonsourceibias.t77 CSoutput.t82 gnd.t0 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X33 gnd.t193 gnd.t191 gnd.t192 gnd.t111 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=0 ps=0 w=7 l=1
X34 CSoutput.t81 commonsourceibias.t78 gnd.t72 gnd.t71 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X35 CSoutput.t80 commonsourceibias.t79 gnd.t304 gnd.t241 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X36 a_n2903_n3924.t11 minus.t6 a_n2982_13878.t7 gnd.t223 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=1.155 ps=7.33 w=7 l=0.7
X37 gnd.t190 gnd.t188 gnd.t189 gnd.t103 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=0 ps=0 w=7 l=1
X38 gnd.t187 gnd.t185 minus.t4 gnd.t186 sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.39 ps=2.78 w=1 l=0.5
X39 CSoutput.t79 commonsourceibias.t80 gnd.t279 gnd.t4 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X40 a_n2903_n3924.t7 diffpairibias.t16 gnd.t41 gnd.t40 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=2.73 ps=14.78 w=7 l=1
X41 CSoutput.t121 a_n8300_8799.t46 vdd.t237 vdd.t189 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X42 gnd.t73 commonsourceibias.t81 CSoutput.t78 gnd.t24 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X43 gnd.t184 gnd.t182 gnd.t183 gnd.t131 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=0 ps=0 w=7 l=0.7
X44 vdd.t236 a_n8300_8799.t47 CSoutput.t120 vdd.t152 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X45 CSoutput.t77 commonsourceibias.t82 gnd.t205 gnd.t2 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=2.73 ps=14.78 w=7 l=1
X46 gnd.t267 commonsourceibias.t60 commonsourceibias.t61 gnd.t61 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X47 CSoutput.t76 commonsourceibias.t83 gnd.t27 gnd.t4 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X48 output.t2 outputibias.t8 gnd.t271 gnd.t270 sky130_fd_pr__nfet_01v8 ad=2.34 pd=12.78 as=2.34 ps=12.78 w=6 l=2
X49 gnd.t246 commonsourceibias.t84 CSoutput.t75 gnd.t200 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X50 a_n2903_n3924.t32 plus.t7 a_n8300_8799.t35 gnd.t66 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.7
X51 CSoutput.t74 commonsourceibias.t85 gnd.t347 gnd.t42 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X52 a_n2804_13878.t30 a_n2982_13878.t59 a_n2982_13878.t60 vdd.t85 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X53 gnd.t289 commonsourceibias.t86 CSoutput.t73 gnd.t200 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X54 vdd.t137 CSoutput.t171 output.t17 gnd.t319 sky130_fd_pr__nfet_01v8 ad=0.825 pd=5.33 as=0.825 ps=5.33 w=5 l=1
X55 CSoutput.t72 commonsourceibias.t87 gnd.t203 gnd.t56 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X56 a_n2982_13878.t14 a_n2982_13878.t13 a_n2804_13878.t29 vdd.t98 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X57 gnd.t212 commonsourceibias.t88 CSoutput.t71 gnd.t12 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X58 a_n8300_8799.t34 plus.t8 a_n2903_n3924.t23 gnd.t35 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.7
X59 CSoutput.t145 a_n8300_8799.t48 vdd.t235 vdd.t180 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X60 gnd.t350 commonsourceibias.t58 commonsourceibias.t59 gnd.t20 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X61 vdd.t75 vdd.t73 vdd.t74 vdd.t50 sky130_fd_pr__pfet_01v8 ad=3.51 pd=18.78 as=0 ps=0 w=9 l=0.5
X62 CSoutput.t70 commonsourceibias.t89 gnd.t234 gnd.t233 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X63 gnd.t181 gnd.t178 gnd.t180 gnd.t179 sky130_fd_pr__nfet_01v8 ad=1.95 pd=10.78 as=0 ps=0 w=5 l=1
X64 vdd.t234 a_n8300_8799.t49 CSoutput.t144 vdd.t200 sky130_fd_pr__pfet_01v8 ad=3.12 pd=16.78 as=1.32 ps=8.33 w=8 l=0.5
X65 gnd.t177 gnd.t175 gnd.t176 gnd.t111 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=0 ps=0 w=7 l=1
X66 CSoutput.t69 commonsourceibias.t90 gnd.t43 gnd.t42 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X67 diffpairibias.t15 diffpairibias.t14 gnd.t256 gnd.t255 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=2.73 ps=14.78 w=7 l=1
X68 a_n2982_13878.t12 minus.t7 a_n2903_n3924.t19 gnd.t288 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.7
X69 a_n2982_13878.t42 a_n2982_13878.t41 a_n2804_13878.t28 vdd.t113 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X70 CSoutput.t68 commonsourceibias.t91 gnd.t3 gnd.t2 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=2.73 ps=14.78 w=7 l=1
X71 CSoutput.t67 commonsourceibias.t92 gnd.t274 gnd.t259 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X72 gnd.t230 commonsourceibias.t93 CSoutput.t66 gnd.t38 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X73 gnd.t239 commonsourceibias.t94 CSoutput.t65 gnd.t22 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X74 a_n8300_8799.t4 a_n2982_13878.t68 a_n2982_8322.t28 vdd.t108 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X75 CSoutput.t143 a_n8300_8799.t50 vdd.t233 vdd.t209 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X76 gnd.t217 commonsourceibias.t95 CSoutput.t64 gnd.t206 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X77 a_n2982_13878.t34 a_n2982_13878.t33 a_n2804_13878.t27 vdd.t129 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X78 vdd.t232 a_n8300_8799.t51 CSoutput.t98 vdd.t162 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X79 vdd.t231 a_n8300_8799.t52 CSoutput.t97 vdd.t216 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X80 a_n8300_8799.t3 a_n2982_13878.t69 a_n2982_8322.t27 vdd.t106 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X81 CSoutput.t63 commonsourceibias.t96 gnd.t273 gnd.t259 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X82 diffpairibias.t13 diffpairibias.t12 gnd.t355 gnd.t354 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=2.73 ps=14.78 w=7 l=1
X83 CSoutput.t96 a_n8300_8799.t53 vdd.t230 vdd.t165 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X84 gnd.t323 commonsourceibias.t56 commonsourceibias.t57 gnd.t248 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X85 gnd.t215 commonsourceibias.t97 CSoutput.t62 gnd.t53 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=1.155 ps=7.33 w=7 l=1
X86 CSoutput.t61 commonsourceibias.t98 gnd.t216 gnd.t56 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X87 a_n8300_8799.t16 a_n2982_13878.t70 a_n2982_8322.t26 vdd.t121 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X88 gnd.t283 commonsourceibias.t99 CSoutput.t60 gnd.t248 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X89 gnd.t174 gnd.t172 gnd.t173 gnd.t93 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=0 ps=0 w=7 l=1
X90 CSoutput.t59 commonsourceibias.t100 gnd.t278 gnd.t63 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X91 CSoutput.t58 commonsourceibias.t101 gnd.t339 gnd.t48 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X92 a_n2982_8322.t25 a_n2982_13878.t71 a_n8300_8799.t1 vdd.t129 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X93 gnd.t340 commonsourceibias.t102 CSoutput.t57 gnd.t0 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X94 vdd.t72 vdd.t70 vdd.t71 vdd.t37 sky130_fd_pr__pfet_01v8 ad=3.12 pd=16.78 as=0 ps=0 w=8 l=0.5
X95 CSoutput.t148 a_n8300_8799.t54 vdd.t229 vdd.t192 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X96 CSoutput.t172 a_n2982_8322.t35 sky130_fd_pr__cap_mim_m3_1 l=12 w=12
X97 gnd.t329 commonsourceibias.t54 commonsourceibias.t55 gnd.t58 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X98 output.t16 CSoutput.t173 vdd.t133 gnd.t321 sky130_fd_pr__nfet_01v8 ad=0.825 pd=5.33 as=0.825 ps=5.33 w=5 l=1
X99 a_n2903_n3924.t21 plus.t9 a_n8300_8799.t33 gnd.t33 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=1.155 ps=7.33 w=7 l=0.7
X100 gnd.t171 gnd.t169 minus.t3 gnd.t170 sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.5
X101 gnd.t342 commonsourceibias.t103 CSoutput.t56 gnd.t248 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X102 a_n2903_n3924.t0 diffpairibias.t17 gnd.t11 gnd.t10 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=2.73 ps=14.78 w=7 l=1
X103 vdd.t228 a_n8300_8799.t55 CSoutput.t147 vdd.t198 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X104 gnd.t168 gnd.t166 gnd.t167 gnd.t89 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=0 ps=0 w=7 l=1
X105 vdd.t227 a_n8300_8799.t56 CSoutput.t146 vdd.t220 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X106 a_n2982_13878.t54 a_n2982_13878.t53 a_n2804_13878.t26 vdd.t128 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X107 vdd.t226 a_n8300_8799.t57 CSoutput.t110 vdd.t205 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X108 gnd.t52 commonsourceibias.t104 CSoutput.t55 gnd.t24 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X109 a_n8300_8799.t10 a_n2982_13878.t72 a_n2982_8322.t24 vdd.t117 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X110 a_n2982_13878.t40 a_n2982_13878.t39 a_n2804_13878.t25 vdd.t80 sky130_fd_pr__pfet_01v8 ad=3.51 pd=18.78 as=1.485 ps=9.33 w=9 l=0.5
X111 gnd.t165 gnd.t163 gnd.t164 gnd.t89 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=0 ps=0 w=7 l=1
X112 CSoutput.t54 commonsourceibias.t105 gnd.t343 gnd.t241 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X113 gnd.t312 commonsourceibias.t106 CSoutput.t53 gnd.t46 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X114 a_n2982_13878.t1 minus.t8 a_n2903_n3924.t3 gnd.t34 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.7
X115 output.t15 CSoutput.t174 vdd.t145 gnd.t322 sky130_fd_pr__nfet_01v8 ad=0.825 pd=5.33 as=0.825 ps=5.33 w=5 l=1
X116 vdd.t69 vdd.t67 vdd.t68 vdd.t57 sky130_fd_pr__pfet_01v8 ad=3.51 pd=18.78 as=0 ps=0 w=9 l=0.5
X117 gnd.t7 commonsourceibias.t52 commonsourceibias.t53 gnd.t6 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X118 gnd.t308 commonsourceibias.t107 CSoutput.t52 gnd.t61 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X119 CSoutput.t109 a_n8300_8799.t58 vdd.t225 vdd.t165 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X120 vdd.t66 vdd.t63 vdd.t65 vdd.t64 sky130_fd_pr__pfet_01v8 ad=3.51 pd=18.78 as=0 ps=0 w=9 l=0.5
X121 output.t1 outputibias.t9 gnd.t236 gnd.t235 sky130_fd_pr__nfet_01v8 ad=2.34 pd=12.78 as=2.34 ps=12.78 w=6 l=2
X122 gnd.t162 gnd.t160 gnd.t161 gnd.t107 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=0 ps=0 w=7 l=0.7
X123 a_n2804_13878.t24 a_n2982_13878.t31 a_n2982_13878.t32 vdd.t90 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=3.51 ps=18.78 w=9 l=0.5
X124 a_n2903_n3924.t16 minus.t9 a_n2982_13878.t10 gnd.t272 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.7
X125 CSoutput.t108 a_n8300_8799.t59 vdd.t224 vdd.t148 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X126 CSoutput.t175 a_n2982_8322.t34 sky130_fd_pr__cap_mim_m3_1 l=12 w=12
X127 vdd.t223 a_n8300_8799.t60 CSoutput.t115 vdd.t220 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X128 vdd.t127 a_n2982_13878.t73 a_n2982_8322.t7 vdd.t126 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X129 a_n2982_13878.t38 a_n2982_13878.t37 a_n2804_13878.t23 vdd.t88 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X130 vdd.t62 vdd.t60 vdd.t61 vdd.t37 sky130_fd_pr__pfet_01v8 ad=3.12 pd=16.78 as=0 ps=0 w=8 l=0.5
X131 a_n2982_8322.t6 a_n2982_13878.t74 vdd.t125 vdd.t124 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X132 gnd.t54 commonsourceibias.t108 CSoutput.t51 gnd.t53 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=1.155 ps=7.33 w=7 l=1
X133 a_n2903_n3924.t1 diffpairibias.t18 gnd.t32 gnd.t31 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=2.73 ps=14.78 w=7 l=1
X134 output.t14 CSoutput.t176 vdd.t141 gnd.t344 sky130_fd_pr__nfet_01v8 ad=0.825 pd=5.33 as=0.825 ps=5.33 w=5 l=1
X135 CSoutput.t114 a_n8300_8799.t61 vdd.t222 vdd.t192 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X136 vdd.t140 CSoutput.t177 output.t13 gnd.t345 sky130_fd_pr__nfet_01v8 ad=0.825 pd=5.33 as=0.825 ps=5.33 w=5 l=1
X137 gnd.t331 commonsourceibias.t109 CSoutput.t50 gnd.t200 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X138 gnd.t225 commonsourceibias.t50 commonsourceibias.t51 gnd.t38 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X139 CSoutput.t49 commonsourceibias.t110 gnd.t333 gnd.t63 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X140 gnd.t334 commonsourceibias.t111 CSoutput.t48 gnd.t58 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X141 CSoutput.t47 commonsourceibias.t112 gnd.t309 gnd.t297 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=2.73 ps=14.78 w=7 l=1
X142 CSoutput.t46 commonsourceibias.t113 gnd.t338 gnd.t29 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X143 a_n2903_n3924.t37 minus.t10 a_n2982_13878.t61 gnd.t314 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.7
X144 CSoutput.t178 a_n2982_8322.t33 sky130_fd_pr__cap_mim_m3_1 l=12 w=12
X145 gnd.t159 gnd.t157 plus.t0 gnd.t158 sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.39 ps=2.78 w=1 l=0.5
X146 vdd.t123 a_n2982_13878.t75 a_n2804_13878.t6 vdd.t122 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X147 a_n2903_n3924.t22 plus.t10 a_n8300_8799.t32 gnd.t243 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.7
X148 vdd.t59 vdd.t56 vdd.t58 vdd.t57 sky130_fd_pr__pfet_01v8 ad=3.51 pd=18.78 as=0 ps=0 w=9 l=0.5
X149 gnd.t156 gnd.t154 gnd.t155 gnd.t89 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=0 ps=0 w=7 l=1
X150 a_n2804_13878.t22 a_n2982_13878.t15 a_n2982_13878.t16 vdd.t121 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X151 vdd.t221 a_n8300_8799.t62 CSoutput.t113 vdd.t220 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X152 vdd.t219 a_n8300_8799.t63 CSoutput.t159 vdd.t205 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X153 a_n2982_8322.t23 a_n2982_13878.t76 a_n8300_8799.t0 vdd.t107 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X154 a_n8300_8799.t31 plus.t11 a_n2903_n3924.t24 gnd.t65 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=2.73 ps=14.78 w=7 l=0.7
X155 a_n8300_8799.t30 plus.t12 a_n2903_n3924.t25 gnd.t287 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=2.73 ps=14.78 w=7 l=0.7
X156 vdd.t55 vdd.t53 vdd.t54 vdd.t19 sky130_fd_pr__pfet_01v8 ad=3.12 pd=16.78 as=0 ps=0 w=8 l=0.5
X157 vdd.t52 vdd.t49 vdd.t51 vdd.t50 sky130_fd_pr__pfet_01v8 ad=3.51 pd=18.78 as=0 ps=0 w=9 l=0.5
X158 a_n2982_8322.t5 a_n2982_13878.t77 vdd.t120 vdd.t119 sky130_fd_pr__pfet_01v8 ad=3.51 pd=18.78 as=1.485 ps=9.33 w=9 l=0.5
X159 a_n8300_8799.t21 a_n2982_13878.t78 a_n2982_8322.t22 vdd.t87 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X160 CSoutput.t158 a_n8300_8799.t64 vdd.t218 vdd.t173 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X161 diffpairibias.t11 diffpairibias.t10 gnd.t349 gnd.t348 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=2.73 ps=14.78 w=7 l=1
X162 vdd.t217 a_n8300_8799.t65 CSoutput.t136 vdd.t216 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X163 a_n2982_13878.t9 minus.t11 a_n2903_n3924.t15 gnd.t266 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.7
X164 a_n2982_13878.t36 a_n2982_13878.t35 a_n2804_13878.t21 vdd.t99 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X165 CSoutput.t45 commonsourceibias.t114 gnd.t310 gnd.t69 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X166 a_n8300_8799.t20 a_n2982_13878.t79 a_n2982_8322.t21 vdd.t118 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X167 commonsourceibias.t49 commonsourceibias.t48 gnd.t45 gnd.t44 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X168 output.t12 CSoutput.t179 vdd.t139 gnd.t293 sky130_fd_pr__nfet_01v8 ad=0.825 pd=5.33 as=0.825 ps=5.33 w=5 l=1
X169 gnd.t237 commonsourceibias.t115 CSoutput.t44 gnd.t12 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X170 a_n2804_13878.t20 a_n2982_13878.t43 a_n2982_13878.t44 vdd.t117 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X171 a_n2903_n3924.t5 minus.t12 a_n2982_13878.t3 gnd.t36 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.7
X172 gnd.t153 gnd.t150 gnd.t152 gnd.t151 sky130_fd_pr__nfet_01v8 ad=1.95 pd=10.78 as=0 ps=0 w=5 l=1
X173 CSoutput.t43 commonsourceibias.t116 gnd.t242 gnd.t241 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X174 minus.t2 gnd.t147 gnd.t149 gnd.t148 sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.5
X175 vdd.t48 vdd.t46 vdd.t47 vdd.t5 sky130_fd_pr__pfet_01v8 ad=3.51 pd=18.78 as=0 ps=0 w=9 l=0.5
X176 output.t11 CSoutput.t180 vdd.t146 gnd.t294 sky130_fd_pr__nfet_01v8 ad=0.825 pd=5.33 as=0.825 ps=5.33 w=5 l=1
X177 CSoutput.t135 a_n8300_8799.t66 vdd.t215 vdd.t209 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X178 CSoutput.t42 commonsourceibias.t117 gnd.t353 gnd.t42 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X179 gnd.t146 gnd.t144 gnd.t145 gnd.t103 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=0 ps=0 w=7 l=1
X180 vdd.t116 a_n2982_13878.t80 a_n2982_8322.t4 vdd.t115 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=3.51 ps=18.78 w=9 l=0.5
X181 a_n2804_13878.t19 a_n2982_13878.t19 a_n2982_13878.t20 vdd.t114 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X182 outputibias.t7 outputibias.t6 gnd.t258 gnd.t257 sky130_fd_pr__nfet_01v8 ad=2.34 pd=12.78 as=2.34 ps=12.78 w=6 l=2
X183 vdd.t214 a_n8300_8799.t67 CSoutput.t125 vdd.t207 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X184 gnd.t341 commonsourceibias.t118 CSoutput.t41 gnd.t22 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X185 gnd.t346 commonsourceibias.t119 CSoutput.t40 gnd.t0 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X186 a_n2982_13878.t28 a_n2982_13878.t27 a_n2804_13878.t18 vdd.t84 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X187 commonsourceibias.t47 commonsourceibias.t46 gnd.t291 gnd.t63 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X188 gnd.t224 commonsourceibias.t120 CSoutput.t39 gnd.t16 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=1.155 ps=7.33 w=7 l=1
X189 outputibias.t5 outputibias.t4 gnd.t253 gnd.t252 sky130_fd_pr__nfet_01v8 ad=2.34 pd=12.78 as=2.34 ps=12.78 w=6 l=2
X190 vdd.t213 a_n8300_8799.t68 CSoutput.t124 vdd.t175 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X191 CSoutput.t38 commonsourceibias.t121 gnd.t197 gnd.t71 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X192 a_n2903_n3924.t10 diffpairibias.t19 gnd.t209 gnd.t208 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=2.73 ps=14.78 w=7 l=1
X193 gnd.t143 gnd.t140 gnd.t142 gnd.t141 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=0 ps=0 w=7 l=1
X194 a_n2903_n3924.t14 diffpairibias.t20 gnd.t265 gnd.t264 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=2.73 ps=14.78 w=7 l=1
X195 commonsourceibias.t45 commonsourceibias.t44 gnd.t238 gnd.t29 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X196 vdd.t212 a_n8300_8799.t69 CSoutput.t123 vdd.t198 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X197 gnd.t139 gnd.t137 gnd.t138 gnd.t111 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=0 ps=0 w=7 l=1
X198 gnd.t136 gnd.t134 gnd.t135 gnd.t103 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=0 ps=0 w=7 l=1
X199 vdd.t45 vdd.t43 vdd.t44 vdd.t19 sky130_fd_pr__pfet_01v8 ad=3.12 pd=16.78 as=0 ps=0 w=8 l=0.5
X200 vdd.t132 CSoutput.t181 output.t10 gnd.t295 sky130_fd_pr__nfet_01v8 ad=0.825 pd=5.33 as=0.825 ps=5.33 w=5 l=1
X201 CSoutput.t37 commonsourceibias.t122 gnd.t250 gnd.t69 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X202 CSoutput.t36 commonsourceibias.t123 gnd.t281 gnd.t48 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X203 a_n2804_13878.t17 a_n2982_13878.t45 a_n2982_13878.t46 vdd.t89 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X204 a_n2982_8322.t20 a_n2982_13878.t81 a_n8300_8799.t18 vdd.t113 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X205 CSoutput.t164 a_n8300_8799.t70 vdd.t211 vdd.t150 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X206 commonsourceibias.t43 commonsourceibias.t42 gnd.t5 gnd.t4 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X207 gnd.t201 commonsourceibias.t40 commonsourceibias.t41 gnd.t200 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X208 vdd.t134 CSoutput.t182 output.t9 gnd.t324 sky130_fd_pr__nfet_01v8 ad=0.825 pd=5.33 as=0.825 ps=5.33 w=5 l=1
X209 diffpairibias.t9 diffpairibias.t8 gnd.t357 gnd.t356 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=2.73 ps=14.78 w=7 l=1
X210 a_n2804_13878.t5 a_n2982_13878.t82 vdd.t112 vdd.t111 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X211 vdd.t110 a_n2982_13878.t83 a_n2804_13878.t4 vdd.t109 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X212 CSoutput.t35 commonsourceibias.t124 gnd.t245 gnd.t71 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X213 CSoutput.t34 commonsourceibias.t125 gnd.t9 gnd.t8 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X214 CSoutput.t163 a_n8300_8799.t71 vdd.t210 vdd.t209 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X215 gnd.t13 commonsourceibias.t38 commonsourceibias.t39 gnd.t12 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X216 vdd.t208 a_n8300_8799.t72 CSoutput.t119 vdd.t207 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X217 gnd.t133 gnd.t130 gnd.t132 gnd.t131 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=0 ps=0 w=7 l=0.7
X218 gnd.t129 gnd.t127 plus.t4 gnd.t128 sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.5
X219 vdd.t206 a_n8300_8799.t73 CSoutput.t118 vdd.t205 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X220 commonsourceibias.t37 commonsourceibias.t36 gnd.t313 gnd.t233 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X221 outputibias.t3 outputibias.t2 gnd.t352 gnd.t351 sky130_fd_pr__nfet_01v8 ad=2.34 pd=12.78 as=2.34 ps=12.78 w=6 l=2
X222 CSoutput.t107 a_n8300_8799.t74 vdd.t204 vdd.t186 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X223 a_n2804_13878.t16 a_n2982_13878.t51 a_n2982_13878.t52 vdd.t108 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X224 a_n2903_n3924.t9 minus.t13 a_n2982_13878.t6 gnd.t66 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.7
X225 gnd.t296 commonsourceibias.t126 CSoutput.t33 gnd.t14 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X226 commonsourceibias.t35 commonsourceibias.t34 gnd.t26 gnd.t2 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=2.73 ps=14.78 w=7 l=1
X227 vdd.t203 a_n8300_8799.t75 CSoutput.t106 vdd.t175 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X228 gnd.t218 commonsourceibias.t32 commonsourceibias.t33 gnd.t206 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X229 a_n2982_8322.t19 a_n2982_13878.t84 a_n8300_8799.t17 vdd.t76 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X230 CSoutput.t32 commonsourceibias.t127 gnd.t226 gnd.t56 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X231 CSoutput.t105 a_n8300_8799.t76 vdd.t202 vdd.t177 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=3.12 ps=16.78 w=8 l=0.5
X232 a_n2982_13878.t18 a_n2982_13878.t17 a_n2804_13878.t15 vdd.t107 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X233 diffpairibias.t7 diffpairibias.t6 gnd.t232 gnd.t231 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=2.73 ps=14.78 w=7 l=1
X234 vdd.t201 a_n8300_8799.t77 CSoutput.t138 vdd.t200 sky130_fd_pr__pfet_01v8 ad=3.12 pd=16.78 as=1.32 ps=8.33 w=8 l=0.5
X235 commonsourceibias.t31 commonsourceibias.t30 gnd.t260 gnd.t259 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X236 a_n2982_13878.t2 minus.t14 a_n2903_n3924.t4 gnd.t35 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.7
X237 a_n2804_13878.t14 a_n2982_13878.t57 a_n2982_13878.t58 vdd.t106 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X238 a_n2982_13878.t62 minus.t15 a_n2903_n3924.t38 gnd.t316 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.7
X239 vdd.t42 vdd.t40 vdd.t41 vdd.t23 sky130_fd_pr__pfet_01v8 ad=3.12 pd=16.78 as=0 ps=0 w=8 l=0.5
X240 vdd.t105 a_n2982_13878.t85 a_n2982_8322.t3 vdd.t104 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=3.51 ps=18.78 w=9 l=0.5
X241 vdd.t199 a_n8300_8799.t78 CSoutput.t137 vdd.t198 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X242 a_n8300_8799.t29 plus.t13 a_n2903_n3924.t31 gnd.t288 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.7
X243 gnd.t15 commonsourceibias.t128 CSoutput.t31 gnd.t14 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X244 a_n2903_n3924.t39 minus.t16 a_n2982_13878.t63 gnd.t315 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.7
X245 CSoutput.t166 a_n8300_8799.t79 vdd.t197 vdd.t189 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X246 gnd.t1 commonsourceibias.t28 commonsourceibias.t29 gnd.t0 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X247 CSoutput.t30 commonsourceibias.t129 gnd.t298 gnd.t297 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=2.73 ps=14.78 w=7 l=1
X248 a_n2804_13878.t3 a_n2982_13878.t86 vdd.t103 vdd.t102 sky130_fd_pr__pfet_01v8 ad=3.51 pd=18.78 as=1.485 ps=9.33 w=9 l=0.5
X249 vdd.t39 vdd.t36 vdd.t38 vdd.t37 sky130_fd_pr__pfet_01v8 ad=3.12 pd=16.78 as=0 ps=0 w=8 l=0.5
X250 vdd.t35 vdd.t33 vdd.t34 vdd.t23 sky130_fd_pr__pfet_01v8 ad=3.12 pd=16.78 as=0 ps=0 w=8 l=0.5
X251 output.t8 CSoutput.t183 vdd.t142 gnd.t325 sky130_fd_pr__nfet_01v8 ad=0.825 pd=5.33 as=0.825 ps=5.33 w=5 l=1
X252 CSoutput.t165 a_n8300_8799.t80 vdd.t196 vdd.t186 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X253 gnd.t39 commonsourceibias.t130 CSoutput.t29 gnd.t38 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X254 gnd.t126 gnd.t123 gnd.t125 gnd.t124 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=0 ps=0 w=7 l=1
X255 vdd.t32 vdd.t30 vdd.t31 vdd.t9 sky130_fd_pr__pfet_01v8 ad=3.12 pd=16.78 as=0 ps=0 w=8 l=0.5
X256 vdd.t195 a_n8300_8799.t81 CSoutput.t128 vdd.t182 sky130_fd_pr__pfet_01v8 ad=3.12 pd=16.78 as=1.32 ps=8.33 w=8 l=0.5
X257 a_n2903_n3924.t13 diffpairibias.t21 gnd.t263 gnd.t262 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=2.73 ps=14.78 w=7 l=1
X258 vdd.t101 a_n2982_13878.t87 a_n2982_8322.t2 vdd.t100 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X259 a_n2982_8322.t18 a_n2982_13878.t88 a_n8300_8799.t19 vdd.t99 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X260 gnd.t292 commonsourceibias.t26 commonsourceibias.t27 gnd.t24 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X261 a_n8300_8799.t28 plus.t14 a_n2903_n3924.t34 gnd.t37 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.7
X262 gnd.t122 gnd.t120 plus.t1 gnd.t121 sky130_fd_pr__nfet_01v8 ad=0.39 pd=2.78 as=0.165 ps=1.33 w=1 l=0.5
X263 output.t19 outputibias.t10 gnd.t359 gnd.t358 sky130_fd_pr__nfet_01v8 ad=2.34 pd=12.78 as=2.34 ps=12.78 w=6 l=2
X264 gnd.t119 gnd.t117 gnd.t118 gnd.t93 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=0 ps=0 w=7 l=1
X265 gnd.t60 commonsourceibias.t24 commonsourceibias.t25 gnd.t46 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X266 vdd.t29 vdd.t26 vdd.t28 vdd.t27 sky130_fd_pr__pfet_01v8 ad=3.51 pd=18.78 as=0 ps=0 w=9 l=0.5
X267 gnd.t116 gnd.t114 gnd.t115 gnd.t93 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=0 ps=0 w=7 l=1
X268 CSoutput.t28 commonsourceibias.t131 gnd.t19 gnd.t18 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X269 a_n2903_n3924.t27 plus.t15 a_n8300_8799.t27 gnd.t223 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=1.155 ps=7.33 w=7 l=0.7
X270 vdd.t194 a_n8300_8799.t82 CSoutput.t127 vdd.t154 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X271 vdd.t138 CSoutput.t184 output.t7 gnd.t326 sky130_fd_pr__nfet_01v8 ad=0.825 pd=5.33 as=0.825 ps=5.33 w=5 l=1
X272 CSoutput.t126 a_n8300_8799.t83 vdd.t193 vdd.t192 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X273 CSoutput.t27 commonsourceibias.t132 gnd.t311 gnd.t4 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X274 output.t0 outputibias.t11 gnd.t222 gnd.t221 sky130_fd_pr__nfet_01v8 ad=2.34 pd=12.78 as=2.34 ps=12.78 w=6 l=2
X275 a_n2804_13878.t13 a_n2982_13878.t23 a_n2982_13878.t24 vdd.t93 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X276 CSoutput.t142 a_n8300_8799.t84 vdd.t191 vdd.t177 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=3.12 ps=16.78 w=8 l=0.5
X277 a_n2982_8322.t17 a_n2982_13878.t89 a_n8300_8799.t2 vdd.t98 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X278 vdd.t25 vdd.t22 vdd.t24 vdd.t23 sky130_fd_pr__pfet_01v8 ad=3.12 pd=16.78 as=0 ps=0 w=8 l=0.5
X279 diffpairibias.t5 diffpairibias.t4 gnd.t211 gnd.t210 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=2.73 ps=14.78 w=7 l=1
X280 gnd.t113 gnd.t110 gnd.t112 gnd.t111 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=0 ps=0 w=7 l=1
X281 CSoutput.t141 a_n8300_8799.t85 vdd.t190 vdd.t189 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X282 CSoutput.t100 a_n8300_8799.t86 vdd.t188 vdd.t173 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X283 gnd.t229 commonsourceibias.t22 commonsourceibias.t23 gnd.t53 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=1.155 ps=7.33 w=7 l=1
X284 output.t6 CSoutput.t185 vdd.t143 gnd.t305 sky130_fd_pr__nfet_01v8 ad=1.95 pd=10.78 as=0.825 ps=5.33 w=5 l=1
X285 vdd.t21 vdd.t18 vdd.t20 vdd.t19 sky130_fd_pr__pfet_01v8 ad=3.12 pd=16.78 as=0 ps=0 w=8 l=0.5
X286 CSoutput.t26 commonsourceibias.t133 gnd.t299 gnd.t259 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X287 a_n2982_8322.t1 a_n2982_13878.t90 vdd.t97 vdd.t96 sky130_fd_pr__pfet_01v8 ad=3.51 pd=18.78 as=1.485 ps=9.33 w=9 l=0.5
X288 CSoutput.t99 a_n8300_8799.t87 vdd.t187 vdd.t186 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X289 gnd.t109 gnd.t106 gnd.t108 gnd.t107 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=0 ps=0 w=7 l=0.7
X290 vdd.t185 a_n8300_8799.t88 CSoutput.t154 vdd.t182 sky130_fd_pr__pfet_01v8 ad=3.12 pd=16.78 as=1.32 ps=8.33 w=8 l=0.5
X291 gnd.t227 commonsourceibias.t134 CSoutput.t25 gnd.t61 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X292 CSoutput.t153 a_n8300_8799.t89 vdd.t184 vdd.t160 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=3.12 ps=16.78 w=8 l=0.5
X293 vdd.t95 a_n2982_13878.t91 a_n2804_13878.t2 vdd.t94 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=3.51 ps=18.78 w=9 l=0.5
X294 vdd.t183 a_n8300_8799.t90 CSoutput.t104 vdd.t182 sky130_fd_pr__pfet_01v8 ad=3.12 pd=16.78 as=1.32 ps=8.33 w=8 l=0.5
X295 CSoutput.t103 a_n8300_8799.t91 vdd.t181 vdd.t180 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X296 gnd.t247 commonsourceibias.t135 CSoutput.t24 gnd.t206 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X297 gnd.t21 commonsourceibias.t136 CSoutput.t23 gnd.t20 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X298 output.t5 CSoutput.t186 vdd.t147 gnd.t306 sky130_fd_pr__nfet_01v8 ad=0.825 pd=5.33 as=0.825 ps=5.33 w=5 l=1
X299 a_n2982_8322.t16 a_n2982_13878.t92 a_n8300_8799.t9 vdd.t86 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X300 commonsourceibias.t21 commonsourceibias.t20 gnd.t76 gnd.t69 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X301 vdd.t144 CSoutput.t187 output.t4 gnd.t307 sky130_fd_pr__nfet_01v8 ad=0.825 pd=5.33 as=1.95 ps=10.78 w=5 l=1
X302 gnd.t101 gnd.t99 minus.t1 gnd.t100 sky130_fd_pr__nfet_01v8 ad=0.39 pd=2.78 as=0.165 ps=1.33 w=1 l=0.5
X303 a_n8300_8799.t11 a_n2982_13878.t93 a_n2982_8322.t15 vdd.t93 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X304 a_n2804_13878.t1 a_n2982_13878.t94 vdd.t92 vdd.t91 sky130_fd_pr__pfet_01v8 ad=3.51 pd=18.78 as=1.485 ps=9.33 w=9 l=0.5
X305 gnd.t47 commonsourceibias.t137 CSoutput.t22 gnd.t46 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X306 vdd.t17 vdd.t15 vdd.t16 vdd.t1 sky130_fd_pr__pfet_01v8 ad=3.51 pd=18.78 as=0 ps=0 w=9 l=0.5
X307 vdd.t179 a_n8300_8799.t92 CSoutput.t150 vdd.t162 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X308 a_n2982_13878.t5 minus.t17 a_n2903_n3924.t8 gnd.t65 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=2.73 ps=14.78 w=7 l=0.7
X309 CSoutput.t149 a_n8300_8799.t93 vdd.t178 vdd.t177 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=3.12 ps=16.78 w=8 l=0.5
X310 commonsourceibias.t19 commonsourceibias.t18 gnd.t336 gnd.t241 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X311 a_n2982_13878.t50 a_n2982_13878.t49 a_n2804_13878.t12 vdd.t81 sky130_fd_pr__pfet_01v8 ad=3.51 pd=18.78 as=1.485 ps=9.33 w=9 l=0.5
X312 a_n8300_8799.t14 a_n2982_13878.t95 a_n2982_8322.t14 vdd.t90 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=3.51 ps=18.78 w=9 l=0.5
X313 gnd.t105 gnd.t102 gnd.t104 gnd.t103 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=0 ps=0 w=7 l=1
X314 minus.t0 gnd.t96 gnd.t98 gnd.t97 sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.5
X315 a_n8300_8799.t8 a_n2982_13878.t96 a_n2982_8322.t13 vdd.t89 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X316 gnd.t23 commonsourceibias.t138 CSoutput.t21 gnd.t22 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X317 commonsourceibias.t17 commonsourceibias.t16 gnd.t67 gnd.t42 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X318 a_n8300_8799.t26 plus.t16 a_n2903_n3924.t26 gnd.t266 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.7
X319 a_n2982_8322.t12 a_n2982_13878.t97 a_n8300_8799.t5 vdd.t88 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X320 gnd.t249 commonsourceibias.t139 CSoutput.t20 gnd.t248 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X321 CSoutput.t19 commonsourceibias.t140 gnd.t302 gnd.t297 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=2.73 ps=14.78 w=7 l=1
X322 a_n2903_n3924.t2 minus.t18 a_n2982_13878.t0 gnd.t33 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=1.155 ps=7.33 w=7 l=0.7
X323 vdd.t176 a_n8300_8799.t94 CSoutput.t152 vdd.t175 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X324 gnd.t290 commonsourceibias.t14 commonsourceibias.t15 gnd.t22 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X325 CSoutput.t151 a_n8300_8799.t95 vdd.t174 vdd.t173 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X326 CSoutput.t102 a_n8300_8799.t96 vdd.t172 vdd.t158 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X327 CSoutput.t101 a_n8300_8799.t97 vdd.t171 vdd.t158 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X328 gnd.t95 gnd.t92 gnd.t94 gnd.t93 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=0 ps=0 w=7 l=1
X329 a_n2804_13878.t11 a_n2982_13878.t25 a_n2982_13878.t26 vdd.t87 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X330 a_n2903_n3924.t35 plus.t17 a_n8300_8799.t25 gnd.t36 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.7
X331 vdd.t170 a_n8300_8799.t98 CSoutput.t157 vdd.t156 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X332 gnd.t17 commonsourceibias.t12 commonsourceibias.t13 gnd.t16 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=1.155 ps=7.33 w=7 l=1
X333 commonsourceibias.t11 commonsourceibias.t10 gnd.t280 gnd.t71 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X334 gnd.t228 commonsourceibias.t141 CSoutput.t18 gnd.t58 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X335 a_n2903_n3924.t17 diffpairibias.t22 gnd.t286 gnd.t285 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=2.73 ps=14.78 w=7 l=1
X336 gnd.t25 commonsourceibias.t142 CSoutput.t17 gnd.t24 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X337 CSoutput.t16 commonsourceibias.t143 gnd.t49 gnd.t48 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X338 vdd.t169 a_n8300_8799.t99 CSoutput.t156 vdd.t154 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X339 gnd.t62 commonsourceibias.t144 CSoutput.t15 gnd.t61 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X340 CSoutput.t155 a_n8300_8799.t100 vdd.t168 vdd.t150 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X341 CSoutput.t14 commonsourceibias.t145 gnd.t68 gnd.t18 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X342 a_n2982_13878.t30 a_n2982_13878.t29 a_n2804_13878.t10 vdd.t86 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X343 gnd.t91 gnd.t88 gnd.t90 gnd.t89 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=0 ps=0 w=7 l=1
X344 a_n8300_8799.t13 a_n2982_13878.t98 a_n2982_8322.t11 vdd.t85 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X345 vdd.t136 CSoutput.t188 output.t3 gnd.t328 sky130_fd_pr__nfet_01v8 ad=0.825 pd=5.33 as=0.825 ps=5.33 w=5 l=1
X346 vdd.t167 a_n8300_8799.t101 CSoutput.t112 vdd.t156 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X347 CSoutput.t111 a_n8300_8799.t102 vdd.t166 vdd.t165 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X348 a_n8300_8799.t24 plus.t18 a_n2903_n3924.t30 gnd.t34 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.7
X349 vdd.t14 vdd.t12 vdd.t13 vdd.t9 sky130_fd_pr__pfet_01v8 ad=3.12 pd=16.78 as=0 ps=0 w=8 l=0.5
X350 CSoutput.t13 commonsourceibias.t146 gnd.t75 gnd.t8 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X351 gnd.t214 commonsourceibias.t147 CSoutput.t12 gnd.t16 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=1.155 ps=7.33 w=7 l=1
X352 commonsourceibias.t9 commonsourceibias.t8 gnd.t55 gnd.t48 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X353 diffpairibias.t3 diffpairibias.t2 gnd.t269 gnd.t268 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=2.73 ps=14.78 w=7 l=1
X354 CSoutput.t117 a_n8300_8799.t103 vdd.t164 vdd.t148 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X355 CSoutput.t189 a_n2982_8322.t32 sky130_fd_pr__cap_mim_m3_1 l=12 w=12
X356 a_n2982_8322.t10 a_n2982_13878.t99 a_n8300_8799.t15 vdd.t84 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X357 gnd.t244 commonsourceibias.t148 CSoutput.t11 gnd.t14 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X358 a_n2903_n3924.t33 plus.t19 a_n8300_8799.t23 gnd.t272 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.7
X359 vdd.t163 a_n8300_8799.t104 CSoutput.t116 vdd.t162 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X360 gnd.t87 gnd.t84 gnd.t86 gnd.t85 sky130_fd_pr__nfet_01v8 ad=2.34 pd=12.78 as=0 ps=0 w=6 l=2
X361 CSoutput.t140 a_n8300_8799.t105 vdd.t161 vdd.t160 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=3.12 ps=16.78 w=8 l=0.5
X362 diffpairibias.t1 diffpairibias.t0 gnd.t51 gnd.t50 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=2.73 ps=14.78 w=7 l=1
X363 gnd.t59 commonsourceibias.t149 CSoutput.t10 gnd.t58 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X364 commonsourceibias.t7 commonsourceibias.t6 gnd.t28 gnd.t8 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X365 gnd.t327 commonsourceibias.t150 CSoutput.t9 gnd.t6 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X366 a_n2903_n3924.t29 plus.t20 a_n8300_8799.t22 gnd.t314 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.7
X367 CSoutput.t8 commonsourceibias.t151 gnd.t213 gnd.t2 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=2.73 ps=14.78 w=7 l=1
X368 vdd.t83 a_n2982_13878.t100 a_n2804_13878.t0 vdd.t82 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=3.51 ps=18.78 w=9 l=0.5
X369 CSoutput.t139 a_n8300_8799.t106 vdd.t159 vdd.t158 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X370 a_n2903_n3924.t12 minus.t19 a_n2982_13878.t8 gnd.t243 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.7
X371 vdd.t157 a_n8300_8799.t107 CSoutput.t132 vdd.t156 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X372 gnd.t219 commonsourceibias.t4 commonsourceibias.t5 gnd.t14 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X373 gnd.t320 commonsourceibias.t152 CSoutput.t7 gnd.t38 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X374 a_n2982_8322.t9 a_n2982_13878.t101 a_n8300_8799.t39 vdd.t81 sky130_fd_pr__pfet_01v8 ad=3.51 pd=18.78 as=1.485 ps=9.33 w=9 l=0.5
X375 a_n2982_13878.t11 minus.t20 a_n2903_n3924.t18 gnd.t287 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=2.73 ps=14.78 w=7 l=0.7
X376 commonsourceibias.t3 commonsourceibias.t2 gnd.t57 gnd.t56 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X377 gnd.t317 commonsourceibias.t153 CSoutput.t6 gnd.t6 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X378 gnd.t83 gnd.t80 gnd.t82 gnd.t81 sky130_fd_pr__nfet_01v8 ad=2.34 pd=12.78 as=0 ps=0 w=6 l=2
X379 gnd.t207 commonsourceibias.t154 CSoutput.t5 gnd.t206 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X380 a_n2982_8322.t8 a_n2982_13878.t102 a_n8300_8799.t6 vdd.t80 sky130_fd_pr__pfet_01v8 ad=3.51 pd=18.78 as=1.485 ps=9.33 w=9 l=0.5
X381 vdd.t155 a_n8300_8799.t108 CSoutput.t131 vdd.t154 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X382 vdd.t153 a_n8300_8799.t109 CSoutput.t130 vdd.t152 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X383 CSoutput.t129 a_n8300_8799.t110 vdd.t151 vdd.t150 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X384 gnd.t337 commonsourceibias.t155 CSoutput.t4 gnd.t20 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X385 plus.t2 gnd.t77 gnd.t79 gnd.t78 sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.5
X386 vdd.t11 vdd.t8 vdd.t10 vdd.t9 sky130_fd_pr__pfet_01v8 ad=3.12 pd=16.78 as=0 ps=0 w=8 l=0.5
X387 a_n2982_8322.t0 a_n2982_13878.t103 vdd.t79 vdd.t78 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X388 gnd.t335 commonsourceibias.t156 CSoutput.t3 gnd.t46 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X389 a_n2804_13878.t9 a_n2982_13878.t21 a_n2982_13878.t22 vdd.t77 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=3.51 ps=18.78 w=9 l=0.5
X390 gnd.t74 commonsourceibias.t157 CSoutput.t2 gnd.t20 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X391 CSoutput.t1 commonsourceibias.t158 gnd.t332 gnd.t8 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X392 commonsourceibias.t1 commonsourceibias.t0 gnd.t303 gnd.t297 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=2.73 ps=14.78 w=7 l=1
X393 CSoutput.t0 commonsourceibias.t159 gnd.t330 gnd.t44 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X394 outputibias.t1 outputibias.t0 gnd.t277 gnd.t276 sky130_fd_pr__nfet_01v8 ad=2.34 pd=12.78 as=2.34 ps=12.78 w=6 l=2
X395 vdd.t7 vdd.t4 vdd.t6 vdd.t5 sky130_fd_pr__pfet_01v8 ad=3.51 pd=18.78 as=0 ps=0 w=9 l=0.5
X396 a_n2903_n3924.t20 diffpairibias.t23 gnd.t301 gnd.t300 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=2.73 ps=14.78 w=7 l=1
X397 vdd.t3 vdd.t0 vdd.t2 vdd.t1 sky130_fd_pr__pfet_01v8 ad=3.51 pd=18.78 as=0 ps=0 w=9 l=0.5
X398 CSoutput.t167 a_n8300_8799.t111 vdd.t149 vdd.t148 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X399 a_n2982_13878.t48 a_n2982_13878.t47 a_n2804_13878.t8 vdd.t76 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
R0 plus.n33 plus.t15 321.495
R1 plus.n7 plus.t12 321.495
R2 plus.n32 plus.t14 297.12
R3 plus.n36 plus.t19 297.12
R4 plus.n38 plus.t18 297.12
R5 plus.n42 plus.t20 297.12
R6 plus.n44 plus.t8 297.12
R7 plus.n48 plus.t7 297.12
R8 plus.n50 plus.t11 297.12
R9 plus.n24 plus.t9 297.12
R10 plus.n22 plus.t5 297.12
R11 plus.n2 plus.t6 297.12
R12 plus.n16 plus.t16 297.12
R13 plus.n4 plus.t17 297.12
R14 plus.n10 plus.t13 297.12
R15 plus.n6 plus.t10 297.12
R16 plus.n54 plus.t0 243.97
R17 plus.n54 plus.n53 223.454
R18 plus.n56 plus.n55 223.454
R19 plus.n51 plus.n50 161.3
R20 plus.n49 plus.n26 161.3
R21 plus.n48 plus.n47 161.3
R22 plus.n46 plus.n27 161.3
R23 plus.n45 plus.n44 161.3
R24 plus.n43 plus.n28 161.3
R25 plus.n42 plus.n41 161.3
R26 plus.n40 plus.n29 161.3
R27 plus.n39 plus.n38 161.3
R28 plus.n37 plus.n30 161.3
R29 plus.n36 plus.n35 161.3
R30 plus.n34 plus.n31 161.3
R31 plus.n9 plus.n8 161.3
R32 plus.n10 plus.n5 161.3
R33 plus.n12 plus.n11 161.3
R34 plus.n13 plus.n4 161.3
R35 plus.n15 plus.n14 161.3
R36 plus.n16 plus.n3 161.3
R37 plus.n18 plus.n17 161.3
R38 plus.n19 plus.n2 161.3
R39 plus.n21 plus.n20 161.3
R40 plus.n22 plus.n1 161.3
R41 plus.n23 plus.n0 161.3
R42 plus.n25 plus.n24 161.3
R43 plus.n34 plus.n33 44.9377
R44 plus.n8 plus.n7 44.9377
R45 plus.n50 plus.n49 37.246
R46 plus.n24 plus.n23 37.246
R47 plus.n32 plus.n31 32.8641
R48 plus.n48 plus.n27 32.8641
R49 plus.n22 plus.n21 32.8641
R50 plus.n9 plus.n6 32.8641
R51 plus.n52 plus.n51 30.0327
R52 plus.n37 plus.n36 28.4823
R53 plus.n44 plus.n43 28.4823
R54 plus.n17 plus.n2 28.4823
R55 plus.n11 plus.n10 28.4823
R56 plus.n38 plus.n29 24.1005
R57 plus.n42 plus.n29 24.1005
R58 plus.n16 plus.n15 24.1005
R59 plus.n15 plus.n4 24.1005
R60 plus.n53 plus.t4 19.8005
R61 plus.n53 plus.t3 19.8005
R62 plus.n55 plus.t1 19.8005
R63 plus.n55 plus.t2 19.8005
R64 plus.n38 plus.n37 19.7187
R65 plus.n43 plus.n42 19.7187
R66 plus.n17 plus.n16 19.7187
R67 plus.n11 plus.n4 19.7187
R68 plus.n33 plus.n32 17.0522
R69 plus.n7 plus.n6 17.0522
R70 plus.n36 plus.n31 15.3369
R71 plus.n44 plus.n27 15.3369
R72 plus.n21 plus.n2 15.3369
R73 plus.n10 plus.n9 15.3369
R74 plus plus.n57 14.3159
R75 plus.n52 plus.n25 11.8547
R76 plus.n49 plus.n48 10.955
R77 plus.n23 plus.n22 10.955
R78 plus.n57 plus.n56 5.40567
R79 plus.n57 plus.n52 1.188
R80 plus.n56 plus.n54 0.716017
R81 plus.n35 plus.n34 0.189894
R82 plus.n35 plus.n30 0.189894
R83 plus.n39 plus.n30 0.189894
R84 plus.n40 plus.n39 0.189894
R85 plus.n41 plus.n40 0.189894
R86 plus.n41 plus.n28 0.189894
R87 plus.n45 plus.n28 0.189894
R88 plus.n46 plus.n45 0.189894
R89 plus.n47 plus.n46 0.189894
R90 plus.n47 plus.n26 0.189894
R91 plus.n51 plus.n26 0.189894
R92 plus.n25 plus.n0 0.189894
R93 plus.n1 plus.n0 0.189894
R94 plus.n20 plus.n1 0.189894
R95 plus.n20 plus.n19 0.189894
R96 plus.n19 plus.n18 0.189894
R97 plus.n18 plus.n3 0.189894
R98 plus.n14 plus.n3 0.189894
R99 plus.n14 plus.n13 0.189894
R100 plus.n13 plus.n12 0.189894
R101 plus.n12 plus.n5 0.189894
R102 plus.n8 plus.n5 0.189894
R103 a_n2903_n3924.n7 a_n2903_n3924.t13 214.994
R104 a_n2903_n3924.n10 a_n2903_n3924.t1 214.714
R105 a_n2903_n3924.n10 a_n2903_n3924.t17 214.321
R106 a_n2903_n3924.n6 a_n2903_n3924.t14 214.321
R107 a_n2903_n3924.n6 a_n2903_n3924.t20 214.321
R108 a_n2903_n3924.n5 a_n2903_n3924.t10 214.321
R109 a_n2903_n3924.n7 a_n2903_n3924.t7 214.321
R110 a_n2903_n3924.n7 a_n2903_n3924.t0 214.321
R111 a_n2903_n3924.n4 a_n2903_n3924.t27 55.8337
R112 a_n2903_n3924.n4 a_n2903_n3924.t18 55.8337
R113 a_n2903_n3924.t2 a_n2903_n3924.n9 55.8337
R114 a_n2903_n3924.n0 a_n2903_n3924.t24 55.8335
R115 a_n2903_n3924.n1 a_n2903_n3924.t8 55.8335
R116 a_n2903_n3924.n8 a_n2903_n3924.t11 55.8335
R117 a_n2903_n3924.n8 a_n2903_n3924.t25 55.8335
R118 a_n2903_n3924.n3 a_n2903_n3924.t21 55.8335
R119 a_n2903_n3924.n0 a_n2903_n3924.n18 53.0052
R120 a_n2903_n3924.n0 a_n2903_n3924.n19 53.0052
R121 a_n2903_n3924.n0 a_n2903_n3924.n20 53.0052
R122 a_n2903_n3924.n4 a_n2903_n3924.n21 53.0052
R123 a_n2903_n3924.n4 a_n2903_n3924.n22 53.0052
R124 a_n2903_n3924.n9 a_n2903_n3924.n23 53.0052
R125 a_n2903_n3924.n1 a_n2903_n3924.n16 53.0051
R126 a_n2903_n3924.n1 a_n2903_n3924.n15 53.0051
R127 a_n2903_n3924.n1 a_n2903_n3924.n14 53.0051
R128 a_n2903_n3924.n8 a_n2903_n3924.n13 53.0051
R129 a_n2903_n3924.n3 a_n2903_n3924.n12 53.0051
R130 a_n2903_n3924.n3 a_n2903_n3924.n11 53.0051
R131 a_n2903_n3924.n9 a_n2903_n3924.n2 12.1986
R132 a_n2903_n3924.n0 a_n2903_n3924.n17 12.1986
R133 a_n2903_n3924.n3 a_n2903_n3924.n2 5.11903
R134 a_n2903_n3924.n17 a_n2903_n3924.n1 5.11903
R135 a_n2903_n3924.n18 a_n2903_n3924.t23 2.82907
R136 a_n2903_n3924.n18 a_n2903_n3924.t32 2.82907
R137 a_n2903_n3924.n19 a_n2903_n3924.t30 2.82907
R138 a_n2903_n3924.n19 a_n2903_n3924.t29 2.82907
R139 a_n2903_n3924.n20 a_n2903_n3924.t34 2.82907
R140 a_n2903_n3924.n20 a_n2903_n3924.t33 2.82907
R141 a_n2903_n3924.n21 a_n2903_n3924.t19 2.82907
R142 a_n2903_n3924.n21 a_n2903_n3924.t12 2.82907
R143 a_n2903_n3924.n22 a_n2903_n3924.t15 2.82907
R144 a_n2903_n3924.n22 a_n2903_n3924.t5 2.82907
R145 a_n2903_n3924.n23 a_n2903_n3924.t38 2.82907
R146 a_n2903_n3924.n23 a_n2903_n3924.t39 2.82907
R147 a_n2903_n3924.n16 a_n2903_n3924.t4 2.82907
R148 a_n2903_n3924.n16 a_n2903_n3924.t9 2.82907
R149 a_n2903_n3924.n15 a_n2903_n3924.t3 2.82907
R150 a_n2903_n3924.n15 a_n2903_n3924.t37 2.82907
R151 a_n2903_n3924.n14 a_n2903_n3924.t6 2.82907
R152 a_n2903_n3924.n14 a_n2903_n3924.t16 2.82907
R153 a_n2903_n3924.n13 a_n2903_n3924.t31 2.82907
R154 a_n2903_n3924.n13 a_n2903_n3924.t22 2.82907
R155 a_n2903_n3924.n12 a_n2903_n3924.t26 2.82907
R156 a_n2903_n3924.n12 a_n2903_n3924.t35 2.82907
R157 a_n2903_n3924.n11 a_n2903_n3924.t28 2.82907
R158 a_n2903_n3924.n11 a_n2903_n3924.t36 2.82907
R159 a_n2903_n3924.n4 a_n2903_n3924.n0 2.45524
R160 a_n2903_n3924.n1 a_n2903_n3924.n8 2.01128
R161 a_n2903_n3924.n17 a_n2903_n3924.n10 1.95694
R162 a_n2903_n3924.n7 a_n2903_n3924.n2 1.95694
R163 a_n2903_n3924.n8 a_n2903_n3924.n3 1.77636
R164 a_n2903_n3924.n6 a_n2903_n3924.n5 1.34352
R165 a_n2903_n3924.n5 a_n2903_n3924.n7 1.34352
R166 a_n2903_n3924.n9 a_n2903_n3924.n4 1.3324
R167 a_n2903_n3924.n10 a_n2903_n3924.n6 0.951808
R168 a_n8300_8799.n138 a_n8300_8799.t105 490.524
R169 a_n8300_8799.n172 a_n8300_8799.t41 490.524
R170 a_n8300_8799.n207 a_n8300_8799.t89 490.524
R171 a_n8300_8799.n32 a_n8300_8799.t81 490.524
R172 a_n8300_8799.n66 a_n8300_8799.t88 490.524
R173 a_n8300_8799.n101 a_n8300_8799.t90 490.524
R174 a_n8300_8799.n159 a_n8300_8799.t43 464.166
R175 a_n8300_8799.n157 a_n8300_8799.t42 464.166
R176 a_n8300_8799.n156 a_n8300_8799.t92 464.166
R177 a_n8300_8799.n130 a_n8300_8799.t53 464.166
R178 a_n8300_8799.n150 a_n8300_8799.t45 464.166
R179 a_n8300_8799.n149 a_n8300_8799.t96 464.166
R180 a_n8300_8799.n133 a_n8300_8799.t69 464.166
R181 a_n8300_8799.n144 a_n8300_8799.t54 464.166
R182 a_n8300_8799.n142 a_n8300_8799.t109 464.166
R183 a_n8300_8799.n136 a_n8300_8799.t80 464.166
R184 a_n8300_8799.n137 a_n8300_8799.t56 464.166
R185 a_n8300_8799.n193 a_n8300_8799.t49 464.166
R186 a_n8300_8799.n191 a_n8300_8799.t48 464.166
R187 a_n8300_8799.n190 a_n8300_8799.t104 464.166
R188 a_n8300_8799.n164 a_n8300_8799.t58 464.166
R189 a_n8300_8799.n184 a_n8300_8799.t52 464.166
R190 a_n8300_8799.n183 a_n8300_8799.t106 464.166
R191 a_n8300_8799.n167 a_n8300_8799.t78 464.166
R192 a_n8300_8799.n178 a_n8300_8799.t61 464.166
R193 a_n8300_8799.n176 a_n8300_8799.t44 464.166
R194 a_n8300_8799.n170 a_n8300_8799.t87 464.166
R195 a_n8300_8799.n171 a_n8300_8799.t62 464.166
R196 a_n8300_8799.n228 a_n8300_8799.t77 464.166
R197 a_n8300_8799.n226 a_n8300_8799.t91 464.166
R198 a_n8300_8799.n225 a_n8300_8799.t51 464.166
R199 a_n8300_8799.n199 a_n8300_8799.t102 464.166
R200 a_n8300_8799.n219 a_n8300_8799.t65 464.166
R201 a_n8300_8799.n218 a_n8300_8799.t97 464.166
R202 a_n8300_8799.n202 a_n8300_8799.t55 464.166
R203 a_n8300_8799.n213 a_n8300_8799.t83 464.166
R204 a_n8300_8799.n211 a_n8300_8799.t47 464.166
R205 a_n8300_8799.n205 a_n8300_8799.t74 464.166
R206 a_n8300_8799.n206 a_n8300_8799.t60 464.166
R207 a_n8300_8799.n31 a_n8300_8799.t103 464.166
R208 a_n8300_8799.n30 a_n8300_8799.t57 464.166
R209 a_n8300_8799.n36 a_n8300_8799.t79 464.166
R210 a_n8300_8799.n28 a_n8300_8799.t99 464.166
R211 a_n8300_8799.n41 a_n8300_8799.t100 464.166
R212 a_n8300_8799.n43 a_n8300_8799.t68 464.166
R213 a_n8300_8799.n26 a_n8300_8799.t86 464.166
R214 a_n8300_8799.n48 a_n8300_8799.t98 464.166
R215 a_n8300_8799.n24 a_n8300_8799.t66 464.166
R216 a_n8300_8799.n53 a_n8300_8799.t67 464.166
R217 a_n8300_8799.n55 a_n8300_8799.t84 464.166
R218 a_n8300_8799.n65 a_n8300_8799.t111 464.166
R219 a_n8300_8799.n64 a_n8300_8799.t63 464.166
R220 a_n8300_8799.n70 a_n8300_8799.t85 464.166
R221 a_n8300_8799.n62 a_n8300_8799.t108 464.166
R222 a_n8300_8799.n75 a_n8300_8799.t110 464.166
R223 a_n8300_8799.n77 a_n8300_8799.t75 464.166
R224 a_n8300_8799.n60 a_n8300_8799.t95 464.166
R225 a_n8300_8799.n82 a_n8300_8799.t107 464.166
R226 a_n8300_8799.n58 a_n8300_8799.t71 464.166
R227 a_n8300_8799.n87 a_n8300_8799.t72 464.166
R228 a_n8300_8799.n89 a_n8300_8799.t93 464.166
R229 a_n8300_8799.n100 a_n8300_8799.t59 464.166
R230 a_n8300_8799.n99 a_n8300_8799.t73 464.166
R231 a_n8300_8799.n105 a_n8300_8799.t46 464.166
R232 a_n8300_8799.n97 a_n8300_8799.t82 464.166
R233 a_n8300_8799.n110 a_n8300_8799.t70 464.166
R234 a_n8300_8799.n112 a_n8300_8799.t94 464.166
R235 a_n8300_8799.n95 a_n8300_8799.t64 464.166
R236 a_n8300_8799.n117 a_n8300_8799.t101 464.166
R237 a_n8300_8799.n93 a_n8300_8799.t50 464.166
R238 a_n8300_8799.n122 a_n8300_8799.t40 464.166
R239 a_n8300_8799.n124 a_n8300_8799.t76 464.166
R240 a_n8300_8799.n139 a_n8300_8799.n136 161.3
R241 a_n8300_8799.n141 a_n8300_8799.n140 161.3
R242 a_n8300_8799.n142 a_n8300_8799.n135 161.3
R243 a_n8300_8799.n143 a_n8300_8799.n134 161.3
R244 a_n8300_8799.n145 a_n8300_8799.n144 161.3
R245 a_n8300_8799.n146 a_n8300_8799.n133 161.3
R246 a_n8300_8799.n148 a_n8300_8799.n147 161.3
R247 a_n8300_8799.n149 a_n8300_8799.n132 161.3
R248 a_n8300_8799.n150 a_n8300_8799.n131 161.3
R249 a_n8300_8799.n152 a_n8300_8799.n151 161.3
R250 a_n8300_8799.n153 a_n8300_8799.n130 161.3
R251 a_n8300_8799.n155 a_n8300_8799.n154 161.3
R252 a_n8300_8799.n156 a_n8300_8799.n129 161.3
R253 a_n8300_8799.n157 a_n8300_8799.n128 161.3
R254 a_n8300_8799.n158 a_n8300_8799.n127 161.3
R255 a_n8300_8799.n160 a_n8300_8799.n159 161.3
R256 a_n8300_8799.n173 a_n8300_8799.n170 161.3
R257 a_n8300_8799.n175 a_n8300_8799.n174 161.3
R258 a_n8300_8799.n176 a_n8300_8799.n169 161.3
R259 a_n8300_8799.n177 a_n8300_8799.n168 161.3
R260 a_n8300_8799.n179 a_n8300_8799.n178 161.3
R261 a_n8300_8799.n180 a_n8300_8799.n167 161.3
R262 a_n8300_8799.n182 a_n8300_8799.n181 161.3
R263 a_n8300_8799.n183 a_n8300_8799.n166 161.3
R264 a_n8300_8799.n184 a_n8300_8799.n165 161.3
R265 a_n8300_8799.n186 a_n8300_8799.n185 161.3
R266 a_n8300_8799.n187 a_n8300_8799.n164 161.3
R267 a_n8300_8799.n189 a_n8300_8799.n188 161.3
R268 a_n8300_8799.n190 a_n8300_8799.n163 161.3
R269 a_n8300_8799.n191 a_n8300_8799.n162 161.3
R270 a_n8300_8799.n192 a_n8300_8799.n161 161.3
R271 a_n8300_8799.n194 a_n8300_8799.n193 161.3
R272 a_n8300_8799.n208 a_n8300_8799.n205 161.3
R273 a_n8300_8799.n210 a_n8300_8799.n209 161.3
R274 a_n8300_8799.n211 a_n8300_8799.n204 161.3
R275 a_n8300_8799.n212 a_n8300_8799.n203 161.3
R276 a_n8300_8799.n214 a_n8300_8799.n213 161.3
R277 a_n8300_8799.n215 a_n8300_8799.n202 161.3
R278 a_n8300_8799.n217 a_n8300_8799.n216 161.3
R279 a_n8300_8799.n218 a_n8300_8799.n201 161.3
R280 a_n8300_8799.n219 a_n8300_8799.n200 161.3
R281 a_n8300_8799.n221 a_n8300_8799.n220 161.3
R282 a_n8300_8799.n222 a_n8300_8799.n199 161.3
R283 a_n8300_8799.n224 a_n8300_8799.n223 161.3
R284 a_n8300_8799.n225 a_n8300_8799.n198 161.3
R285 a_n8300_8799.n226 a_n8300_8799.n197 161.3
R286 a_n8300_8799.n227 a_n8300_8799.n196 161.3
R287 a_n8300_8799.n229 a_n8300_8799.n228 161.3
R288 a_n8300_8799.n56 a_n8300_8799.n55 161.3
R289 a_n8300_8799.n54 a_n8300_8799.n23 161.3
R290 a_n8300_8799.n53 a_n8300_8799.n52 161.3
R291 a_n8300_8799.n51 a_n8300_8799.n24 161.3
R292 a_n8300_8799.n50 a_n8300_8799.n49 161.3
R293 a_n8300_8799.n48 a_n8300_8799.n25 161.3
R294 a_n8300_8799.n47 a_n8300_8799.n46 161.3
R295 a_n8300_8799.n45 a_n8300_8799.n26 161.3
R296 a_n8300_8799.n44 a_n8300_8799.n43 161.3
R297 a_n8300_8799.n42 a_n8300_8799.n27 161.3
R298 a_n8300_8799.n41 a_n8300_8799.n40 161.3
R299 a_n8300_8799.n39 a_n8300_8799.n28 161.3
R300 a_n8300_8799.n38 a_n8300_8799.n37 161.3
R301 a_n8300_8799.n36 a_n8300_8799.n29 161.3
R302 a_n8300_8799.n35 a_n8300_8799.n34 161.3
R303 a_n8300_8799.n33 a_n8300_8799.n30 161.3
R304 a_n8300_8799.n90 a_n8300_8799.n89 161.3
R305 a_n8300_8799.n88 a_n8300_8799.n57 161.3
R306 a_n8300_8799.n87 a_n8300_8799.n86 161.3
R307 a_n8300_8799.n85 a_n8300_8799.n58 161.3
R308 a_n8300_8799.n84 a_n8300_8799.n83 161.3
R309 a_n8300_8799.n82 a_n8300_8799.n59 161.3
R310 a_n8300_8799.n81 a_n8300_8799.n80 161.3
R311 a_n8300_8799.n79 a_n8300_8799.n60 161.3
R312 a_n8300_8799.n78 a_n8300_8799.n77 161.3
R313 a_n8300_8799.n76 a_n8300_8799.n61 161.3
R314 a_n8300_8799.n75 a_n8300_8799.n74 161.3
R315 a_n8300_8799.n73 a_n8300_8799.n62 161.3
R316 a_n8300_8799.n72 a_n8300_8799.n71 161.3
R317 a_n8300_8799.n70 a_n8300_8799.n63 161.3
R318 a_n8300_8799.n69 a_n8300_8799.n68 161.3
R319 a_n8300_8799.n67 a_n8300_8799.n64 161.3
R320 a_n8300_8799.n125 a_n8300_8799.n124 161.3
R321 a_n8300_8799.n123 a_n8300_8799.n92 161.3
R322 a_n8300_8799.n122 a_n8300_8799.n121 161.3
R323 a_n8300_8799.n120 a_n8300_8799.n93 161.3
R324 a_n8300_8799.n119 a_n8300_8799.n118 161.3
R325 a_n8300_8799.n117 a_n8300_8799.n94 161.3
R326 a_n8300_8799.n116 a_n8300_8799.n115 161.3
R327 a_n8300_8799.n114 a_n8300_8799.n95 161.3
R328 a_n8300_8799.n113 a_n8300_8799.n112 161.3
R329 a_n8300_8799.n111 a_n8300_8799.n96 161.3
R330 a_n8300_8799.n110 a_n8300_8799.n109 161.3
R331 a_n8300_8799.n108 a_n8300_8799.n97 161.3
R332 a_n8300_8799.n107 a_n8300_8799.n106 161.3
R333 a_n8300_8799.n105 a_n8300_8799.n98 161.3
R334 a_n8300_8799.n104 a_n8300_8799.n103 161.3
R335 a_n8300_8799.n102 a_n8300_8799.n99 161.3
R336 a_n8300_8799.n13 a_n8300_8799.n11 98.9633
R337 a_n8300_8799.n2 a_n8300_8799.n0 98.9631
R338 a_n8300_8799.n21 a_n8300_8799.n20 98.6055
R339 a_n8300_8799.n19 a_n8300_8799.n18 98.6055
R340 a_n8300_8799.n17 a_n8300_8799.n16 98.6055
R341 a_n8300_8799.n15 a_n8300_8799.n14 98.6055
R342 a_n8300_8799.n13 a_n8300_8799.n12 98.6055
R343 a_n8300_8799.n2 a_n8300_8799.n1 98.6055
R344 a_n8300_8799.n4 a_n8300_8799.n3 98.6055
R345 a_n8300_8799.n6 a_n8300_8799.n5 98.6055
R346 a_n8300_8799.n8 a_n8300_8799.n7 98.6055
R347 a_n8300_8799.n10 a_n8300_8799.n9 98.6055
R348 a_n8300_8799.n247 a_n8300_8799.n246 81.3766
R349 a_n8300_8799.n235 a_n8300_8799.n233 81.3764
R350 a_n8300_8799.n243 a_n8300_8799.n241 81.3764
R351 a_n8300_8799.n240 a_n8300_8799.n239 80.9324
R352 a_n8300_8799.n238 a_n8300_8799.n237 80.9324
R353 a_n8300_8799.n235 a_n8300_8799.n234 80.9324
R354 a_n8300_8799.n243 a_n8300_8799.n242 80.9324
R355 a_n8300_8799.n246 a_n8300_8799.n245 80.9324
R356 a_n8300_8799.n157 a_n8300_8799.n156 48.2005
R357 a_n8300_8799.n150 a_n8300_8799.n149 48.2005
R358 a_n8300_8799.n144 a_n8300_8799.n133 48.2005
R359 a_n8300_8799.n137 a_n8300_8799.n136 48.2005
R360 a_n8300_8799.n191 a_n8300_8799.n190 48.2005
R361 a_n8300_8799.n184 a_n8300_8799.n183 48.2005
R362 a_n8300_8799.n178 a_n8300_8799.n167 48.2005
R363 a_n8300_8799.n171 a_n8300_8799.n170 48.2005
R364 a_n8300_8799.n226 a_n8300_8799.n225 48.2005
R365 a_n8300_8799.n219 a_n8300_8799.n218 48.2005
R366 a_n8300_8799.n213 a_n8300_8799.n202 48.2005
R367 a_n8300_8799.n206 a_n8300_8799.n205 48.2005
R368 a_n8300_8799.n31 a_n8300_8799.n30 48.2005
R369 a_n8300_8799.n41 a_n8300_8799.n28 48.2005
R370 a_n8300_8799.n43 a_n8300_8799.n26 48.2005
R371 a_n8300_8799.n53 a_n8300_8799.n24 48.2005
R372 a_n8300_8799.n65 a_n8300_8799.n64 48.2005
R373 a_n8300_8799.n75 a_n8300_8799.n62 48.2005
R374 a_n8300_8799.n77 a_n8300_8799.n60 48.2005
R375 a_n8300_8799.n87 a_n8300_8799.n58 48.2005
R376 a_n8300_8799.n100 a_n8300_8799.n99 48.2005
R377 a_n8300_8799.n110 a_n8300_8799.n97 48.2005
R378 a_n8300_8799.n112 a_n8300_8799.n95 48.2005
R379 a_n8300_8799.n122 a_n8300_8799.n93 48.2005
R380 a_n8300_8799.n151 a_n8300_8799.n130 47.4702
R381 a_n8300_8799.n143 a_n8300_8799.n142 47.4702
R382 a_n8300_8799.n185 a_n8300_8799.n164 47.4702
R383 a_n8300_8799.n177 a_n8300_8799.n176 47.4702
R384 a_n8300_8799.n220 a_n8300_8799.n199 47.4702
R385 a_n8300_8799.n212 a_n8300_8799.n211 47.4702
R386 a_n8300_8799.n37 a_n8300_8799.n36 47.4702
R387 a_n8300_8799.n48 a_n8300_8799.n47 47.4702
R388 a_n8300_8799.n71 a_n8300_8799.n70 47.4702
R389 a_n8300_8799.n82 a_n8300_8799.n81 47.4702
R390 a_n8300_8799.n106 a_n8300_8799.n105 47.4702
R391 a_n8300_8799.n117 a_n8300_8799.n116 47.4702
R392 a_n8300_8799.n159 a_n8300_8799.n158 46.0096
R393 a_n8300_8799.n193 a_n8300_8799.n192 46.0096
R394 a_n8300_8799.n228 a_n8300_8799.n227 46.0096
R395 a_n8300_8799.n55 a_n8300_8799.n54 46.0096
R396 a_n8300_8799.n89 a_n8300_8799.n88 46.0096
R397 a_n8300_8799.n124 a_n8300_8799.n123 46.0096
R398 a_n8300_8799.n33 a_n8300_8799.n32 45.0871
R399 a_n8300_8799.n67 a_n8300_8799.n66 45.0871
R400 a_n8300_8799.n102 a_n8300_8799.n101 45.0871
R401 a_n8300_8799.n139 a_n8300_8799.n138 45.0871
R402 a_n8300_8799.n173 a_n8300_8799.n172 45.0871
R403 a_n8300_8799.n208 a_n8300_8799.n207 45.0871
R404 a_n8300_8799.n22 a_n8300_8799.n10 33.7114
R405 a_n8300_8799.n244 a_n8300_8799.n240 32.0866
R406 a_n8300_8799.n155 a_n8300_8799.n130 25.5611
R407 a_n8300_8799.n142 a_n8300_8799.n141 25.5611
R408 a_n8300_8799.n189 a_n8300_8799.n164 25.5611
R409 a_n8300_8799.n176 a_n8300_8799.n175 25.5611
R410 a_n8300_8799.n224 a_n8300_8799.n199 25.5611
R411 a_n8300_8799.n211 a_n8300_8799.n210 25.5611
R412 a_n8300_8799.n36 a_n8300_8799.n35 25.5611
R413 a_n8300_8799.n49 a_n8300_8799.n48 25.5611
R414 a_n8300_8799.n70 a_n8300_8799.n69 25.5611
R415 a_n8300_8799.n83 a_n8300_8799.n82 25.5611
R416 a_n8300_8799.n105 a_n8300_8799.n104 25.5611
R417 a_n8300_8799.n118 a_n8300_8799.n117 25.5611
R418 a_n8300_8799.n149 a_n8300_8799.n148 24.1005
R419 a_n8300_8799.n148 a_n8300_8799.n133 24.1005
R420 a_n8300_8799.n183 a_n8300_8799.n182 24.1005
R421 a_n8300_8799.n182 a_n8300_8799.n167 24.1005
R422 a_n8300_8799.n218 a_n8300_8799.n217 24.1005
R423 a_n8300_8799.n217 a_n8300_8799.n202 24.1005
R424 a_n8300_8799.n42 a_n8300_8799.n41 24.1005
R425 a_n8300_8799.n43 a_n8300_8799.n42 24.1005
R426 a_n8300_8799.n76 a_n8300_8799.n75 24.1005
R427 a_n8300_8799.n77 a_n8300_8799.n76 24.1005
R428 a_n8300_8799.n111 a_n8300_8799.n110 24.1005
R429 a_n8300_8799.n112 a_n8300_8799.n111 24.1005
R430 a_n8300_8799.n156 a_n8300_8799.n155 22.6399
R431 a_n8300_8799.n141 a_n8300_8799.n136 22.6399
R432 a_n8300_8799.n190 a_n8300_8799.n189 22.6399
R433 a_n8300_8799.n175 a_n8300_8799.n170 22.6399
R434 a_n8300_8799.n225 a_n8300_8799.n224 22.6399
R435 a_n8300_8799.n210 a_n8300_8799.n205 22.6399
R436 a_n8300_8799.n35 a_n8300_8799.n30 22.6399
R437 a_n8300_8799.n49 a_n8300_8799.n24 22.6399
R438 a_n8300_8799.n69 a_n8300_8799.n64 22.6399
R439 a_n8300_8799.n83 a_n8300_8799.n58 22.6399
R440 a_n8300_8799.n104 a_n8300_8799.n99 22.6399
R441 a_n8300_8799.n118 a_n8300_8799.n93 22.6399
R442 a_n8300_8799.n22 a_n8300_8799.n21 21.1779
R443 a_n8300_8799.n138 a_n8300_8799.n137 14.1472
R444 a_n8300_8799.n172 a_n8300_8799.n171 14.1472
R445 a_n8300_8799.n207 a_n8300_8799.n206 14.1472
R446 a_n8300_8799.n32 a_n8300_8799.n31 14.1472
R447 a_n8300_8799.n66 a_n8300_8799.n65 14.1472
R448 a_n8300_8799.n101 a_n8300_8799.n100 14.1472
R449 a_n8300_8799.n236 a_n8300_8799.n232 12.3339
R450 a_n8300_8799.n232 a_n8300_8799.n22 11.4887
R451 a_n8300_8799.n195 a_n8300_8799.n160 9.01755
R452 a_n8300_8799.n91 a_n8300_8799.n56 9.01755
R453 a_n8300_8799.n231 a_n8300_8799.n126 7.14965
R454 a_n8300_8799.n231 a_n8300_8799.n230 6.85731
R455 a_n8300_8799.n195 a_n8300_8799.n194 4.90959
R456 a_n8300_8799.n230 a_n8300_8799.n229 4.90959
R457 a_n8300_8799.n91 a_n8300_8799.n90 4.90959
R458 a_n8300_8799.n126 a_n8300_8799.n125 4.90959
R459 a_n8300_8799.n230 a_n8300_8799.n195 4.10845
R460 a_n8300_8799.n126 a_n8300_8799.n91 4.10845
R461 a_n8300_8799.n20 a_n8300_8799.t0 3.61217
R462 a_n8300_8799.n20 a_n8300_8799.t14 3.61217
R463 a_n8300_8799.n18 a_n8300_8799.t18 3.61217
R464 a_n8300_8799.n18 a_n8300_8799.t3 3.61217
R465 a_n8300_8799.n16 a_n8300_8799.t15 3.61217
R466 a_n8300_8799.n16 a_n8300_8799.t38 3.61217
R467 a_n8300_8799.n14 a_n8300_8799.t2 3.61217
R468 a_n8300_8799.n14 a_n8300_8799.t13 3.61217
R469 a_n8300_8799.n12 a_n8300_8799.t17 3.61217
R470 a_n8300_8799.n12 a_n8300_8799.t10 3.61217
R471 a_n8300_8799.n11 a_n8300_8799.t6 3.61217
R472 a_n8300_8799.n11 a_n8300_8799.t20 3.61217
R473 a_n8300_8799.n0 a_n8300_8799.t19 3.61217
R474 a_n8300_8799.n0 a_n8300_8799.t12 3.61217
R475 a_n8300_8799.n1 a_n8300_8799.t7 3.61217
R476 a_n8300_8799.n1 a_n8300_8799.t21 3.61217
R477 a_n8300_8799.n3 a_n8300_8799.t9 3.61217
R478 a_n8300_8799.n3 a_n8300_8799.t11 3.61217
R479 a_n8300_8799.n5 a_n8300_8799.t5 3.61217
R480 a_n8300_8799.n5 a_n8300_8799.t4 3.61217
R481 a_n8300_8799.n7 a_n8300_8799.t1 3.61217
R482 a_n8300_8799.n7 a_n8300_8799.t8 3.61217
R483 a_n8300_8799.n9 a_n8300_8799.t39 3.61217
R484 a_n8300_8799.n9 a_n8300_8799.t16 3.61217
R485 a_n8300_8799.n232 a_n8300_8799.n231 3.4105
R486 a_n8300_8799.n241 a_n8300_8799.t32 2.82907
R487 a_n8300_8799.n241 a_n8300_8799.t30 2.82907
R488 a_n8300_8799.n242 a_n8300_8799.t25 2.82907
R489 a_n8300_8799.n242 a_n8300_8799.t29 2.82907
R490 a_n8300_8799.n245 a_n8300_8799.t36 2.82907
R491 a_n8300_8799.n245 a_n8300_8799.t26 2.82907
R492 a_n8300_8799.n239 a_n8300_8799.t35 2.82907
R493 a_n8300_8799.n239 a_n8300_8799.t31 2.82907
R494 a_n8300_8799.n237 a_n8300_8799.t22 2.82907
R495 a_n8300_8799.n237 a_n8300_8799.t34 2.82907
R496 a_n8300_8799.n234 a_n8300_8799.t23 2.82907
R497 a_n8300_8799.n234 a_n8300_8799.t24 2.82907
R498 a_n8300_8799.n233 a_n8300_8799.t27 2.82907
R499 a_n8300_8799.n233 a_n8300_8799.t28 2.82907
R500 a_n8300_8799.n247 a_n8300_8799.t33 2.82907
R501 a_n8300_8799.t37 a_n8300_8799.n247 2.82907
R502 a_n8300_8799.n158 a_n8300_8799.n157 2.19141
R503 a_n8300_8799.n192 a_n8300_8799.n191 2.19141
R504 a_n8300_8799.n227 a_n8300_8799.n226 2.19141
R505 a_n8300_8799.n54 a_n8300_8799.n53 2.19141
R506 a_n8300_8799.n88 a_n8300_8799.n87 2.19141
R507 a_n8300_8799.n123 a_n8300_8799.n122 2.19141
R508 a_n8300_8799.n151 a_n8300_8799.n150 0.730803
R509 a_n8300_8799.n144 a_n8300_8799.n143 0.730803
R510 a_n8300_8799.n185 a_n8300_8799.n184 0.730803
R511 a_n8300_8799.n178 a_n8300_8799.n177 0.730803
R512 a_n8300_8799.n220 a_n8300_8799.n219 0.730803
R513 a_n8300_8799.n213 a_n8300_8799.n212 0.730803
R514 a_n8300_8799.n37 a_n8300_8799.n28 0.730803
R515 a_n8300_8799.n47 a_n8300_8799.n26 0.730803
R516 a_n8300_8799.n71 a_n8300_8799.n62 0.730803
R517 a_n8300_8799.n81 a_n8300_8799.n60 0.730803
R518 a_n8300_8799.n106 a_n8300_8799.n97 0.730803
R519 a_n8300_8799.n116 a_n8300_8799.n95 0.730803
R520 a_n8300_8799.n240 a_n8300_8799.n238 0.444466
R521 a_n8300_8799.n15 a_n8300_8799.n13 0.358259
R522 a_n8300_8799.n17 a_n8300_8799.n15 0.358259
R523 a_n8300_8799.n19 a_n8300_8799.n17 0.358259
R524 a_n8300_8799.n21 a_n8300_8799.n19 0.358259
R525 a_n8300_8799.n10 a_n8300_8799.n8 0.358259
R526 a_n8300_8799.n8 a_n8300_8799.n6 0.358259
R527 a_n8300_8799.n6 a_n8300_8799.n4 0.358259
R528 a_n8300_8799.n4 a_n8300_8799.n2 0.358259
R529 a_n8300_8799.n236 a_n8300_8799.n235 0.222483
R530 a_n8300_8799.n238 a_n8300_8799.n236 0.222483
R531 a_n8300_8799.n246 a_n8300_8799.n244 0.222483
R532 a_n8300_8799.n244 a_n8300_8799.n243 0.222483
R533 a_n8300_8799.n160 a_n8300_8799.n127 0.189894
R534 a_n8300_8799.n128 a_n8300_8799.n127 0.189894
R535 a_n8300_8799.n129 a_n8300_8799.n128 0.189894
R536 a_n8300_8799.n154 a_n8300_8799.n129 0.189894
R537 a_n8300_8799.n154 a_n8300_8799.n153 0.189894
R538 a_n8300_8799.n153 a_n8300_8799.n152 0.189894
R539 a_n8300_8799.n152 a_n8300_8799.n131 0.189894
R540 a_n8300_8799.n132 a_n8300_8799.n131 0.189894
R541 a_n8300_8799.n147 a_n8300_8799.n132 0.189894
R542 a_n8300_8799.n147 a_n8300_8799.n146 0.189894
R543 a_n8300_8799.n146 a_n8300_8799.n145 0.189894
R544 a_n8300_8799.n145 a_n8300_8799.n134 0.189894
R545 a_n8300_8799.n135 a_n8300_8799.n134 0.189894
R546 a_n8300_8799.n140 a_n8300_8799.n135 0.189894
R547 a_n8300_8799.n140 a_n8300_8799.n139 0.189894
R548 a_n8300_8799.n194 a_n8300_8799.n161 0.189894
R549 a_n8300_8799.n162 a_n8300_8799.n161 0.189894
R550 a_n8300_8799.n163 a_n8300_8799.n162 0.189894
R551 a_n8300_8799.n188 a_n8300_8799.n163 0.189894
R552 a_n8300_8799.n188 a_n8300_8799.n187 0.189894
R553 a_n8300_8799.n187 a_n8300_8799.n186 0.189894
R554 a_n8300_8799.n186 a_n8300_8799.n165 0.189894
R555 a_n8300_8799.n166 a_n8300_8799.n165 0.189894
R556 a_n8300_8799.n181 a_n8300_8799.n166 0.189894
R557 a_n8300_8799.n181 a_n8300_8799.n180 0.189894
R558 a_n8300_8799.n180 a_n8300_8799.n179 0.189894
R559 a_n8300_8799.n179 a_n8300_8799.n168 0.189894
R560 a_n8300_8799.n169 a_n8300_8799.n168 0.189894
R561 a_n8300_8799.n174 a_n8300_8799.n169 0.189894
R562 a_n8300_8799.n174 a_n8300_8799.n173 0.189894
R563 a_n8300_8799.n229 a_n8300_8799.n196 0.189894
R564 a_n8300_8799.n197 a_n8300_8799.n196 0.189894
R565 a_n8300_8799.n198 a_n8300_8799.n197 0.189894
R566 a_n8300_8799.n223 a_n8300_8799.n198 0.189894
R567 a_n8300_8799.n223 a_n8300_8799.n222 0.189894
R568 a_n8300_8799.n222 a_n8300_8799.n221 0.189894
R569 a_n8300_8799.n221 a_n8300_8799.n200 0.189894
R570 a_n8300_8799.n201 a_n8300_8799.n200 0.189894
R571 a_n8300_8799.n216 a_n8300_8799.n201 0.189894
R572 a_n8300_8799.n216 a_n8300_8799.n215 0.189894
R573 a_n8300_8799.n215 a_n8300_8799.n214 0.189894
R574 a_n8300_8799.n214 a_n8300_8799.n203 0.189894
R575 a_n8300_8799.n204 a_n8300_8799.n203 0.189894
R576 a_n8300_8799.n209 a_n8300_8799.n204 0.189894
R577 a_n8300_8799.n209 a_n8300_8799.n208 0.189894
R578 a_n8300_8799.n34 a_n8300_8799.n33 0.189894
R579 a_n8300_8799.n34 a_n8300_8799.n29 0.189894
R580 a_n8300_8799.n38 a_n8300_8799.n29 0.189894
R581 a_n8300_8799.n39 a_n8300_8799.n38 0.189894
R582 a_n8300_8799.n40 a_n8300_8799.n39 0.189894
R583 a_n8300_8799.n40 a_n8300_8799.n27 0.189894
R584 a_n8300_8799.n44 a_n8300_8799.n27 0.189894
R585 a_n8300_8799.n45 a_n8300_8799.n44 0.189894
R586 a_n8300_8799.n46 a_n8300_8799.n45 0.189894
R587 a_n8300_8799.n46 a_n8300_8799.n25 0.189894
R588 a_n8300_8799.n50 a_n8300_8799.n25 0.189894
R589 a_n8300_8799.n51 a_n8300_8799.n50 0.189894
R590 a_n8300_8799.n52 a_n8300_8799.n51 0.189894
R591 a_n8300_8799.n52 a_n8300_8799.n23 0.189894
R592 a_n8300_8799.n56 a_n8300_8799.n23 0.189894
R593 a_n8300_8799.n68 a_n8300_8799.n67 0.189894
R594 a_n8300_8799.n68 a_n8300_8799.n63 0.189894
R595 a_n8300_8799.n72 a_n8300_8799.n63 0.189894
R596 a_n8300_8799.n73 a_n8300_8799.n72 0.189894
R597 a_n8300_8799.n74 a_n8300_8799.n73 0.189894
R598 a_n8300_8799.n74 a_n8300_8799.n61 0.189894
R599 a_n8300_8799.n78 a_n8300_8799.n61 0.189894
R600 a_n8300_8799.n79 a_n8300_8799.n78 0.189894
R601 a_n8300_8799.n80 a_n8300_8799.n79 0.189894
R602 a_n8300_8799.n80 a_n8300_8799.n59 0.189894
R603 a_n8300_8799.n84 a_n8300_8799.n59 0.189894
R604 a_n8300_8799.n85 a_n8300_8799.n84 0.189894
R605 a_n8300_8799.n86 a_n8300_8799.n85 0.189894
R606 a_n8300_8799.n86 a_n8300_8799.n57 0.189894
R607 a_n8300_8799.n90 a_n8300_8799.n57 0.189894
R608 a_n8300_8799.n103 a_n8300_8799.n102 0.189894
R609 a_n8300_8799.n103 a_n8300_8799.n98 0.189894
R610 a_n8300_8799.n107 a_n8300_8799.n98 0.189894
R611 a_n8300_8799.n108 a_n8300_8799.n107 0.189894
R612 a_n8300_8799.n109 a_n8300_8799.n108 0.189894
R613 a_n8300_8799.n109 a_n8300_8799.n96 0.189894
R614 a_n8300_8799.n113 a_n8300_8799.n96 0.189894
R615 a_n8300_8799.n114 a_n8300_8799.n113 0.189894
R616 a_n8300_8799.n115 a_n8300_8799.n114 0.189894
R617 a_n8300_8799.n115 a_n8300_8799.n94 0.189894
R618 a_n8300_8799.n119 a_n8300_8799.n94 0.189894
R619 a_n8300_8799.n120 a_n8300_8799.n119 0.189894
R620 a_n8300_8799.n121 a_n8300_8799.n120 0.189894
R621 a_n8300_8799.n121 a_n8300_8799.n92 0.189894
R622 a_n8300_8799.n125 a_n8300_8799.n92 0.189894
R623 gnd.n7083 gnd.n525 1768.67
R624 gnd.n5047 gnd.n5046 939.716
R625 gnd.n7558 gnd.n208 795.207
R626 gnd.n348 gnd.n211 795.207
R627 gnd.n3771 gnd.n1601 795.207
R628 gnd.n3840 gnd.n1603 795.207
R629 gnd.n4789 gnd.n1372 795.207
R630 gnd.n3078 gnd.n1375 795.207
R631 gnd.n2743 gnd.n1067 795.207
R632 gnd.n2700 gnd.n2699 795.207
R633 gnd.n3143 gnd.n2335 771.183
R634 gnd.n4563 gnd.n1578 771.183
R635 gnd.n3145 gnd.n2332 771.183
R636 gnd.n3928 gnd.n1580 771.183
R637 gnd.n6429 gnd.n1026 766.379
R638 gnd.n6345 gnd.n1028 766.379
R639 gnd.n5557 gnd.n5456 766.379
R640 gnd.n5555 gnd.n5458 766.379
R641 gnd.n6426 gnd.n5049 756.769
R642 gnd.n6395 gnd.n1029 756.769
R643 gnd.n5689 gnd.n5418 756.769
R644 gnd.n5675 gnd.n5407 756.769
R645 gnd.n7556 gnd.n213 739.952
R646 gnd.n7447 gnd.n210 739.952
R647 gnd.n4322 gnd.n1600 739.952
R648 gnd.n4545 gnd.n1604 739.952
R649 gnd.n4787 gnd.n1377 739.952
R650 gnd.n2456 gnd.n1374 739.952
R651 gnd.n4924 gnd.n1140 739.952
R652 gnd.n5044 gnd.n1071 739.952
R653 gnd.n6630 gnd.n800 670.282
R654 gnd.n7084 gnd.n526 670.282
R655 gnd.n7297 gnd.n399 670.282
R656 gnd.n2791 gnd.n2785 670.282
R657 gnd.n6630 gnd.n6629 585
R658 gnd.n6631 gnd.n6630 585
R659 gnd.n6628 gnd.n802 585
R660 gnd.n802 gnd.n801 585
R661 gnd.n6627 gnd.n6626 585
R662 gnd.n6626 gnd.n6625 585
R663 gnd.n807 gnd.n806 585
R664 gnd.n6624 gnd.n807 585
R665 gnd.n6622 gnd.n6621 585
R666 gnd.n6623 gnd.n6622 585
R667 gnd.n6620 gnd.n809 585
R668 gnd.n809 gnd.n808 585
R669 gnd.n6619 gnd.n6618 585
R670 gnd.n6618 gnd.n6617 585
R671 gnd.n815 gnd.n814 585
R672 gnd.n6616 gnd.n815 585
R673 gnd.n6614 gnd.n6613 585
R674 gnd.n6615 gnd.n6614 585
R675 gnd.n6612 gnd.n817 585
R676 gnd.n817 gnd.n816 585
R677 gnd.n6611 gnd.n6610 585
R678 gnd.n6610 gnd.n6609 585
R679 gnd.n823 gnd.n822 585
R680 gnd.n6608 gnd.n823 585
R681 gnd.n6606 gnd.n6605 585
R682 gnd.n6607 gnd.n6606 585
R683 gnd.n6604 gnd.n825 585
R684 gnd.n825 gnd.n824 585
R685 gnd.n6603 gnd.n6602 585
R686 gnd.n6602 gnd.n6601 585
R687 gnd.n831 gnd.n830 585
R688 gnd.n6600 gnd.n831 585
R689 gnd.n6598 gnd.n6597 585
R690 gnd.n6599 gnd.n6598 585
R691 gnd.n6596 gnd.n833 585
R692 gnd.n833 gnd.n832 585
R693 gnd.n6595 gnd.n6594 585
R694 gnd.n6594 gnd.n6593 585
R695 gnd.n839 gnd.n838 585
R696 gnd.n6592 gnd.n839 585
R697 gnd.n6590 gnd.n6589 585
R698 gnd.n6591 gnd.n6590 585
R699 gnd.n6588 gnd.n841 585
R700 gnd.n841 gnd.n840 585
R701 gnd.n6587 gnd.n6586 585
R702 gnd.n6586 gnd.n6585 585
R703 gnd.n847 gnd.n846 585
R704 gnd.n6584 gnd.n847 585
R705 gnd.n6582 gnd.n6581 585
R706 gnd.n6583 gnd.n6582 585
R707 gnd.n6580 gnd.n849 585
R708 gnd.n849 gnd.n848 585
R709 gnd.n6579 gnd.n6578 585
R710 gnd.n6578 gnd.n6577 585
R711 gnd.n855 gnd.n854 585
R712 gnd.n6576 gnd.n855 585
R713 gnd.n6574 gnd.n6573 585
R714 gnd.n6575 gnd.n6574 585
R715 gnd.n6572 gnd.n857 585
R716 gnd.n857 gnd.n856 585
R717 gnd.n6571 gnd.n6570 585
R718 gnd.n6570 gnd.n6569 585
R719 gnd.n863 gnd.n862 585
R720 gnd.n6568 gnd.n863 585
R721 gnd.n6566 gnd.n6565 585
R722 gnd.n6567 gnd.n6566 585
R723 gnd.n6564 gnd.n865 585
R724 gnd.n865 gnd.n864 585
R725 gnd.n6563 gnd.n6562 585
R726 gnd.n6562 gnd.n6561 585
R727 gnd.n871 gnd.n870 585
R728 gnd.n6560 gnd.n871 585
R729 gnd.n6558 gnd.n6557 585
R730 gnd.n6559 gnd.n6558 585
R731 gnd.n6556 gnd.n873 585
R732 gnd.n873 gnd.n872 585
R733 gnd.n6555 gnd.n6554 585
R734 gnd.n6554 gnd.n6553 585
R735 gnd.n879 gnd.n878 585
R736 gnd.n6552 gnd.n879 585
R737 gnd.n6550 gnd.n6549 585
R738 gnd.n6551 gnd.n6550 585
R739 gnd.n6548 gnd.n881 585
R740 gnd.n881 gnd.n880 585
R741 gnd.n6547 gnd.n6546 585
R742 gnd.n6546 gnd.n6545 585
R743 gnd.n887 gnd.n886 585
R744 gnd.n6544 gnd.n887 585
R745 gnd.n6542 gnd.n6541 585
R746 gnd.n6543 gnd.n6542 585
R747 gnd.n6540 gnd.n889 585
R748 gnd.n889 gnd.n888 585
R749 gnd.n6539 gnd.n6538 585
R750 gnd.n6538 gnd.n6537 585
R751 gnd.n895 gnd.n894 585
R752 gnd.n6536 gnd.n895 585
R753 gnd.n6534 gnd.n6533 585
R754 gnd.n6535 gnd.n6534 585
R755 gnd.n6532 gnd.n897 585
R756 gnd.n897 gnd.n896 585
R757 gnd.n6531 gnd.n6530 585
R758 gnd.n6530 gnd.n6529 585
R759 gnd.n903 gnd.n902 585
R760 gnd.n6528 gnd.n903 585
R761 gnd.n6526 gnd.n6525 585
R762 gnd.n6527 gnd.n6526 585
R763 gnd.n6524 gnd.n905 585
R764 gnd.n905 gnd.n904 585
R765 gnd.n6523 gnd.n6522 585
R766 gnd.n6522 gnd.n6521 585
R767 gnd.n911 gnd.n910 585
R768 gnd.n6520 gnd.n911 585
R769 gnd.n6518 gnd.n6517 585
R770 gnd.n6519 gnd.n6518 585
R771 gnd.n6516 gnd.n913 585
R772 gnd.n913 gnd.n912 585
R773 gnd.n6515 gnd.n6514 585
R774 gnd.n6514 gnd.n6513 585
R775 gnd.n919 gnd.n918 585
R776 gnd.n6512 gnd.n919 585
R777 gnd.n6510 gnd.n6509 585
R778 gnd.n6511 gnd.n6510 585
R779 gnd.n6508 gnd.n921 585
R780 gnd.n921 gnd.n920 585
R781 gnd.n6507 gnd.n6506 585
R782 gnd.n6506 gnd.n6505 585
R783 gnd.n927 gnd.n926 585
R784 gnd.n6504 gnd.n927 585
R785 gnd.n6502 gnd.n6501 585
R786 gnd.n6503 gnd.n6502 585
R787 gnd.n6500 gnd.n929 585
R788 gnd.n929 gnd.n928 585
R789 gnd.n6499 gnd.n6498 585
R790 gnd.n6498 gnd.n6497 585
R791 gnd.n935 gnd.n934 585
R792 gnd.n6496 gnd.n935 585
R793 gnd.n6494 gnd.n6493 585
R794 gnd.n6495 gnd.n6494 585
R795 gnd.n6492 gnd.n937 585
R796 gnd.n937 gnd.n936 585
R797 gnd.n6491 gnd.n6490 585
R798 gnd.n6490 gnd.n6489 585
R799 gnd.n943 gnd.n942 585
R800 gnd.n6488 gnd.n943 585
R801 gnd.n6486 gnd.n6485 585
R802 gnd.n6487 gnd.n6486 585
R803 gnd.n6484 gnd.n945 585
R804 gnd.n945 gnd.n944 585
R805 gnd.n6483 gnd.n6482 585
R806 gnd.n6482 gnd.n6481 585
R807 gnd.n951 gnd.n950 585
R808 gnd.n6480 gnd.n951 585
R809 gnd.n6478 gnd.n6477 585
R810 gnd.n6479 gnd.n6478 585
R811 gnd.n6476 gnd.n953 585
R812 gnd.n953 gnd.n952 585
R813 gnd.n6475 gnd.n6474 585
R814 gnd.n6474 gnd.n6473 585
R815 gnd.n959 gnd.n958 585
R816 gnd.n6472 gnd.n959 585
R817 gnd.n6470 gnd.n6469 585
R818 gnd.n6471 gnd.n6470 585
R819 gnd.n6468 gnd.n961 585
R820 gnd.n961 gnd.n960 585
R821 gnd.n6467 gnd.n6466 585
R822 gnd.n6466 gnd.n6465 585
R823 gnd.n967 gnd.n966 585
R824 gnd.n6464 gnd.n967 585
R825 gnd.n800 gnd.n799 585
R826 gnd.n6632 gnd.n800 585
R827 gnd.n6635 gnd.n6634 585
R828 gnd.n6634 gnd.n6633 585
R829 gnd.n797 gnd.n796 585
R830 gnd.n796 gnd.n795 585
R831 gnd.n6640 gnd.n6639 585
R832 gnd.n6641 gnd.n6640 585
R833 gnd.n794 gnd.n793 585
R834 gnd.n6642 gnd.n794 585
R835 gnd.n6645 gnd.n6644 585
R836 gnd.n6644 gnd.n6643 585
R837 gnd.n791 gnd.n790 585
R838 gnd.n790 gnd.n789 585
R839 gnd.n6650 gnd.n6649 585
R840 gnd.n6651 gnd.n6650 585
R841 gnd.n788 gnd.n787 585
R842 gnd.n6652 gnd.n788 585
R843 gnd.n6655 gnd.n6654 585
R844 gnd.n6654 gnd.n6653 585
R845 gnd.n785 gnd.n784 585
R846 gnd.n784 gnd.n783 585
R847 gnd.n6660 gnd.n6659 585
R848 gnd.n6661 gnd.n6660 585
R849 gnd.n782 gnd.n781 585
R850 gnd.n6662 gnd.n782 585
R851 gnd.n6665 gnd.n6664 585
R852 gnd.n6664 gnd.n6663 585
R853 gnd.n779 gnd.n778 585
R854 gnd.n778 gnd.n777 585
R855 gnd.n6670 gnd.n6669 585
R856 gnd.n6671 gnd.n6670 585
R857 gnd.n776 gnd.n775 585
R858 gnd.n6672 gnd.n776 585
R859 gnd.n6675 gnd.n6674 585
R860 gnd.n6674 gnd.n6673 585
R861 gnd.n773 gnd.n772 585
R862 gnd.n772 gnd.n771 585
R863 gnd.n6680 gnd.n6679 585
R864 gnd.n6681 gnd.n6680 585
R865 gnd.n770 gnd.n769 585
R866 gnd.n6682 gnd.n770 585
R867 gnd.n6685 gnd.n6684 585
R868 gnd.n6684 gnd.n6683 585
R869 gnd.n767 gnd.n766 585
R870 gnd.n766 gnd.n765 585
R871 gnd.n6690 gnd.n6689 585
R872 gnd.n6691 gnd.n6690 585
R873 gnd.n764 gnd.n763 585
R874 gnd.n6692 gnd.n764 585
R875 gnd.n6695 gnd.n6694 585
R876 gnd.n6694 gnd.n6693 585
R877 gnd.n761 gnd.n760 585
R878 gnd.n760 gnd.n759 585
R879 gnd.n6700 gnd.n6699 585
R880 gnd.n6701 gnd.n6700 585
R881 gnd.n758 gnd.n757 585
R882 gnd.n6702 gnd.n758 585
R883 gnd.n6705 gnd.n6704 585
R884 gnd.n6704 gnd.n6703 585
R885 gnd.n755 gnd.n754 585
R886 gnd.n754 gnd.n753 585
R887 gnd.n6710 gnd.n6709 585
R888 gnd.n6711 gnd.n6710 585
R889 gnd.n752 gnd.n751 585
R890 gnd.n6712 gnd.n752 585
R891 gnd.n6715 gnd.n6714 585
R892 gnd.n6714 gnd.n6713 585
R893 gnd.n749 gnd.n748 585
R894 gnd.n748 gnd.n747 585
R895 gnd.n6720 gnd.n6719 585
R896 gnd.n6721 gnd.n6720 585
R897 gnd.n746 gnd.n745 585
R898 gnd.n6722 gnd.n746 585
R899 gnd.n6725 gnd.n6724 585
R900 gnd.n6724 gnd.n6723 585
R901 gnd.n743 gnd.n742 585
R902 gnd.n742 gnd.n741 585
R903 gnd.n6730 gnd.n6729 585
R904 gnd.n6731 gnd.n6730 585
R905 gnd.n740 gnd.n739 585
R906 gnd.n6732 gnd.n740 585
R907 gnd.n6735 gnd.n6734 585
R908 gnd.n6734 gnd.n6733 585
R909 gnd.n737 gnd.n736 585
R910 gnd.n736 gnd.n735 585
R911 gnd.n6740 gnd.n6739 585
R912 gnd.n6741 gnd.n6740 585
R913 gnd.n734 gnd.n733 585
R914 gnd.n6742 gnd.n734 585
R915 gnd.n6745 gnd.n6744 585
R916 gnd.n6744 gnd.n6743 585
R917 gnd.n731 gnd.n730 585
R918 gnd.n730 gnd.n729 585
R919 gnd.n6750 gnd.n6749 585
R920 gnd.n6751 gnd.n6750 585
R921 gnd.n728 gnd.n727 585
R922 gnd.n6752 gnd.n728 585
R923 gnd.n6755 gnd.n6754 585
R924 gnd.n6754 gnd.n6753 585
R925 gnd.n725 gnd.n724 585
R926 gnd.n724 gnd.n723 585
R927 gnd.n6760 gnd.n6759 585
R928 gnd.n6761 gnd.n6760 585
R929 gnd.n722 gnd.n721 585
R930 gnd.n6762 gnd.n722 585
R931 gnd.n6765 gnd.n6764 585
R932 gnd.n6764 gnd.n6763 585
R933 gnd.n719 gnd.n718 585
R934 gnd.n718 gnd.n717 585
R935 gnd.n6770 gnd.n6769 585
R936 gnd.n6771 gnd.n6770 585
R937 gnd.n716 gnd.n715 585
R938 gnd.n6772 gnd.n716 585
R939 gnd.n6775 gnd.n6774 585
R940 gnd.n6774 gnd.n6773 585
R941 gnd.n713 gnd.n712 585
R942 gnd.n712 gnd.n711 585
R943 gnd.n6780 gnd.n6779 585
R944 gnd.n6781 gnd.n6780 585
R945 gnd.n710 gnd.n709 585
R946 gnd.n6782 gnd.n710 585
R947 gnd.n6785 gnd.n6784 585
R948 gnd.n6784 gnd.n6783 585
R949 gnd.n707 gnd.n706 585
R950 gnd.n706 gnd.n705 585
R951 gnd.n6790 gnd.n6789 585
R952 gnd.n6791 gnd.n6790 585
R953 gnd.n704 gnd.n703 585
R954 gnd.n6792 gnd.n704 585
R955 gnd.n6795 gnd.n6794 585
R956 gnd.n6794 gnd.n6793 585
R957 gnd.n701 gnd.n700 585
R958 gnd.n700 gnd.n699 585
R959 gnd.n6800 gnd.n6799 585
R960 gnd.n6801 gnd.n6800 585
R961 gnd.n698 gnd.n697 585
R962 gnd.n6802 gnd.n698 585
R963 gnd.n6805 gnd.n6804 585
R964 gnd.n6804 gnd.n6803 585
R965 gnd.n695 gnd.n694 585
R966 gnd.n694 gnd.n693 585
R967 gnd.n6810 gnd.n6809 585
R968 gnd.n6811 gnd.n6810 585
R969 gnd.n692 gnd.n691 585
R970 gnd.n6812 gnd.n692 585
R971 gnd.n6815 gnd.n6814 585
R972 gnd.n6814 gnd.n6813 585
R973 gnd.n689 gnd.n688 585
R974 gnd.n688 gnd.n687 585
R975 gnd.n6820 gnd.n6819 585
R976 gnd.n6821 gnd.n6820 585
R977 gnd.n686 gnd.n685 585
R978 gnd.n6822 gnd.n686 585
R979 gnd.n6825 gnd.n6824 585
R980 gnd.n6824 gnd.n6823 585
R981 gnd.n683 gnd.n682 585
R982 gnd.n682 gnd.n681 585
R983 gnd.n6830 gnd.n6829 585
R984 gnd.n6831 gnd.n6830 585
R985 gnd.n680 gnd.n679 585
R986 gnd.n6832 gnd.n680 585
R987 gnd.n6835 gnd.n6834 585
R988 gnd.n6834 gnd.n6833 585
R989 gnd.n677 gnd.n676 585
R990 gnd.n676 gnd.n675 585
R991 gnd.n6840 gnd.n6839 585
R992 gnd.n6841 gnd.n6840 585
R993 gnd.n674 gnd.n673 585
R994 gnd.n6842 gnd.n674 585
R995 gnd.n6845 gnd.n6844 585
R996 gnd.n6844 gnd.n6843 585
R997 gnd.n671 gnd.n670 585
R998 gnd.n670 gnd.n669 585
R999 gnd.n6850 gnd.n6849 585
R1000 gnd.n6851 gnd.n6850 585
R1001 gnd.n668 gnd.n667 585
R1002 gnd.n6852 gnd.n668 585
R1003 gnd.n6855 gnd.n6854 585
R1004 gnd.n6854 gnd.n6853 585
R1005 gnd.n665 gnd.n664 585
R1006 gnd.n664 gnd.n663 585
R1007 gnd.n6860 gnd.n6859 585
R1008 gnd.n6861 gnd.n6860 585
R1009 gnd.n662 gnd.n661 585
R1010 gnd.n6862 gnd.n662 585
R1011 gnd.n6865 gnd.n6864 585
R1012 gnd.n6864 gnd.n6863 585
R1013 gnd.n659 gnd.n658 585
R1014 gnd.n658 gnd.n657 585
R1015 gnd.n6870 gnd.n6869 585
R1016 gnd.n6871 gnd.n6870 585
R1017 gnd.n656 gnd.n655 585
R1018 gnd.n6872 gnd.n656 585
R1019 gnd.n6875 gnd.n6874 585
R1020 gnd.n6874 gnd.n6873 585
R1021 gnd.n653 gnd.n652 585
R1022 gnd.n652 gnd.n651 585
R1023 gnd.n6880 gnd.n6879 585
R1024 gnd.n6881 gnd.n6880 585
R1025 gnd.n650 gnd.n649 585
R1026 gnd.n6882 gnd.n650 585
R1027 gnd.n6885 gnd.n6884 585
R1028 gnd.n6884 gnd.n6883 585
R1029 gnd.n647 gnd.n646 585
R1030 gnd.n646 gnd.n645 585
R1031 gnd.n6890 gnd.n6889 585
R1032 gnd.n6891 gnd.n6890 585
R1033 gnd.n644 gnd.n643 585
R1034 gnd.n6892 gnd.n644 585
R1035 gnd.n6895 gnd.n6894 585
R1036 gnd.n6894 gnd.n6893 585
R1037 gnd.n641 gnd.n640 585
R1038 gnd.n640 gnd.n639 585
R1039 gnd.n6900 gnd.n6899 585
R1040 gnd.n6901 gnd.n6900 585
R1041 gnd.n638 gnd.n637 585
R1042 gnd.n6902 gnd.n638 585
R1043 gnd.n6905 gnd.n6904 585
R1044 gnd.n6904 gnd.n6903 585
R1045 gnd.n635 gnd.n634 585
R1046 gnd.n634 gnd.n633 585
R1047 gnd.n6910 gnd.n6909 585
R1048 gnd.n6911 gnd.n6910 585
R1049 gnd.n632 gnd.n631 585
R1050 gnd.n6912 gnd.n632 585
R1051 gnd.n6915 gnd.n6914 585
R1052 gnd.n6914 gnd.n6913 585
R1053 gnd.n629 gnd.n628 585
R1054 gnd.n628 gnd.n627 585
R1055 gnd.n6920 gnd.n6919 585
R1056 gnd.n6921 gnd.n6920 585
R1057 gnd.n626 gnd.n625 585
R1058 gnd.n6922 gnd.n626 585
R1059 gnd.n6925 gnd.n6924 585
R1060 gnd.n6924 gnd.n6923 585
R1061 gnd.n623 gnd.n622 585
R1062 gnd.n622 gnd.n621 585
R1063 gnd.n6930 gnd.n6929 585
R1064 gnd.n6931 gnd.n6930 585
R1065 gnd.n620 gnd.n619 585
R1066 gnd.n6932 gnd.n620 585
R1067 gnd.n6935 gnd.n6934 585
R1068 gnd.n6934 gnd.n6933 585
R1069 gnd.n617 gnd.n616 585
R1070 gnd.n616 gnd.n615 585
R1071 gnd.n6940 gnd.n6939 585
R1072 gnd.n6941 gnd.n6940 585
R1073 gnd.n614 gnd.n613 585
R1074 gnd.n6942 gnd.n614 585
R1075 gnd.n6945 gnd.n6944 585
R1076 gnd.n6944 gnd.n6943 585
R1077 gnd.n611 gnd.n610 585
R1078 gnd.n610 gnd.n609 585
R1079 gnd.n6950 gnd.n6949 585
R1080 gnd.n6951 gnd.n6950 585
R1081 gnd.n608 gnd.n607 585
R1082 gnd.n6952 gnd.n608 585
R1083 gnd.n6955 gnd.n6954 585
R1084 gnd.n6954 gnd.n6953 585
R1085 gnd.n605 gnd.n604 585
R1086 gnd.n604 gnd.n603 585
R1087 gnd.n6960 gnd.n6959 585
R1088 gnd.n6961 gnd.n6960 585
R1089 gnd.n602 gnd.n601 585
R1090 gnd.n6962 gnd.n602 585
R1091 gnd.n6965 gnd.n6964 585
R1092 gnd.n6964 gnd.n6963 585
R1093 gnd.n599 gnd.n598 585
R1094 gnd.n598 gnd.n597 585
R1095 gnd.n6970 gnd.n6969 585
R1096 gnd.n6971 gnd.n6970 585
R1097 gnd.n596 gnd.n595 585
R1098 gnd.n6972 gnd.n596 585
R1099 gnd.n6975 gnd.n6974 585
R1100 gnd.n6974 gnd.n6973 585
R1101 gnd.n593 gnd.n592 585
R1102 gnd.n592 gnd.n591 585
R1103 gnd.n6980 gnd.n6979 585
R1104 gnd.n6981 gnd.n6980 585
R1105 gnd.n590 gnd.n589 585
R1106 gnd.n6982 gnd.n590 585
R1107 gnd.n6985 gnd.n6984 585
R1108 gnd.n6984 gnd.n6983 585
R1109 gnd.n587 gnd.n586 585
R1110 gnd.n586 gnd.n585 585
R1111 gnd.n6990 gnd.n6989 585
R1112 gnd.n6991 gnd.n6990 585
R1113 gnd.n584 gnd.n583 585
R1114 gnd.n6992 gnd.n584 585
R1115 gnd.n6995 gnd.n6994 585
R1116 gnd.n6994 gnd.n6993 585
R1117 gnd.n581 gnd.n580 585
R1118 gnd.n580 gnd.n579 585
R1119 gnd.n7000 gnd.n6999 585
R1120 gnd.n7001 gnd.n7000 585
R1121 gnd.n578 gnd.n577 585
R1122 gnd.n7002 gnd.n578 585
R1123 gnd.n7005 gnd.n7004 585
R1124 gnd.n7004 gnd.n7003 585
R1125 gnd.n575 gnd.n574 585
R1126 gnd.n574 gnd.n573 585
R1127 gnd.n7010 gnd.n7009 585
R1128 gnd.n7011 gnd.n7010 585
R1129 gnd.n572 gnd.n571 585
R1130 gnd.n7012 gnd.n572 585
R1131 gnd.n7015 gnd.n7014 585
R1132 gnd.n7014 gnd.n7013 585
R1133 gnd.n569 gnd.n568 585
R1134 gnd.n568 gnd.n567 585
R1135 gnd.n7020 gnd.n7019 585
R1136 gnd.n7021 gnd.n7020 585
R1137 gnd.n566 gnd.n565 585
R1138 gnd.n7022 gnd.n566 585
R1139 gnd.n7025 gnd.n7024 585
R1140 gnd.n7024 gnd.n7023 585
R1141 gnd.n563 gnd.n562 585
R1142 gnd.n562 gnd.n561 585
R1143 gnd.n7030 gnd.n7029 585
R1144 gnd.n7031 gnd.n7030 585
R1145 gnd.n560 gnd.n559 585
R1146 gnd.n7032 gnd.n560 585
R1147 gnd.n7035 gnd.n7034 585
R1148 gnd.n7034 gnd.n7033 585
R1149 gnd.n557 gnd.n556 585
R1150 gnd.n556 gnd.n555 585
R1151 gnd.n7040 gnd.n7039 585
R1152 gnd.n7041 gnd.n7040 585
R1153 gnd.n554 gnd.n553 585
R1154 gnd.n7042 gnd.n554 585
R1155 gnd.n7045 gnd.n7044 585
R1156 gnd.n7044 gnd.n7043 585
R1157 gnd.n551 gnd.n550 585
R1158 gnd.n550 gnd.n549 585
R1159 gnd.n7050 gnd.n7049 585
R1160 gnd.n7051 gnd.n7050 585
R1161 gnd.n548 gnd.n547 585
R1162 gnd.n7052 gnd.n548 585
R1163 gnd.n7055 gnd.n7054 585
R1164 gnd.n7054 gnd.n7053 585
R1165 gnd.n545 gnd.n544 585
R1166 gnd.n544 gnd.n543 585
R1167 gnd.n7060 gnd.n7059 585
R1168 gnd.n7061 gnd.n7060 585
R1169 gnd.n542 gnd.n541 585
R1170 gnd.n7062 gnd.n542 585
R1171 gnd.n7065 gnd.n7064 585
R1172 gnd.n7064 gnd.n7063 585
R1173 gnd.n539 gnd.n538 585
R1174 gnd.n538 gnd.n537 585
R1175 gnd.n7070 gnd.n7069 585
R1176 gnd.n7071 gnd.n7070 585
R1177 gnd.n536 gnd.n535 585
R1178 gnd.n7072 gnd.n536 585
R1179 gnd.n7075 gnd.n7074 585
R1180 gnd.n7074 gnd.n7073 585
R1181 gnd.n533 gnd.n532 585
R1182 gnd.n532 gnd.n531 585
R1183 gnd.n7080 gnd.n7079 585
R1184 gnd.n7081 gnd.n7080 585
R1185 gnd.n530 gnd.n529 585
R1186 gnd.n7082 gnd.n530 585
R1187 gnd.n7085 gnd.n7084 585
R1188 gnd.n7084 gnd.n7083 585
R1189 gnd.n7296 gnd.n403 585
R1190 gnd.n7296 gnd.n7295 585
R1191 gnd.n7290 gnd.n404 585
R1192 gnd.n7294 gnd.n404 585
R1193 gnd.n7292 gnd.n7291 585
R1194 gnd.n7293 gnd.n7292 585
R1195 gnd.n407 gnd.n406 585
R1196 gnd.n406 gnd.n405 585
R1197 gnd.n7285 gnd.n7284 585
R1198 gnd.n7284 gnd.n7283 585
R1199 gnd.n410 gnd.n409 585
R1200 gnd.n7282 gnd.n410 585
R1201 gnd.n7280 gnd.n7279 585
R1202 gnd.n7281 gnd.n7280 585
R1203 gnd.n413 gnd.n412 585
R1204 gnd.n412 gnd.n411 585
R1205 gnd.n7275 gnd.n7274 585
R1206 gnd.n7274 gnd.n7273 585
R1207 gnd.n416 gnd.n415 585
R1208 gnd.n7272 gnd.n416 585
R1209 gnd.n7270 gnd.n7269 585
R1210 gnd.n7271 gnd.n7270 585
R1211 gnd.n419 gnd.n418 585
R1212 gnd.n418 gnd.n417 585
R1213 gnd.n7265 gnd.n7264 585
R1214 gnd.n7264 gnd.n7263 585
R1215 gnd.n422 gnd.n421 585
R1216 gnd.n7262 gnd.n422 585
R1217 gnd.n7260 gnd.n7259 585
R1218 gnd.n7261 gnd.n7260 585
R1219 gnd.n425 gnd.n424 585
R1220 gnd.n424 gnd.n423 585
R1221 gnd.n7255 gnd.n7254 585
R1222 gnd.n7254 gnd.n7253 585
R1223 gnd.n428 gnd.n427 585
R1224 gnd.n7252 gnd.n428 585
R1225 gnd.n7250 gnd.n7249 585
R1226 gnd.n7251 gnd.n7250 585
R1227 gnd.n431 gnd.n430 585
R1228 gnd.n430 gnd.n429 585
R1229 gnd.n7245 gnd.n7244 585
R1230 gnd.n7244 gnd.n7243 585
R1231 gnd.n434 gnd.n433 585
R1232 gnd.n7242 gnd.n434 585
R1233 gnd.n7240 gnd.n7239 585
R1234 gnd.n7241 gnd.n7240 585
R1235 gnd.n437 gnd.n436 585
R1236 gnd.n436 gnd.n435 585
R1237 gnd.n7235 gnd.n7234 585
R1238 gnd.n7234 gnd.n7233 585
R1239 gnd.n440 gnd.n439 585
R1240 gnd.n7232 gnd.n440 585
R1241 gnd.n7230 gnd.n7229 585
R1242 gnd.n7231 gnd.n7230 585
R1243 gnd.n443 gnd.n442 585
R1244 gnd.n442 gnd.n441 585
R1245 gnd.n7225 gnd.n7224 585
R1246 gnd.n7224 gnd.n7223 585
R1247 gnd.n446 gnd.n445 585
R1248 gnd.n7222 gnd.n446 585
R1249 gnd.n7220 gnd.n7219 585
R1250 gnd.n7221 gnd.n7220 585
R1251 gnd.n449 gnd.n448 585
R1252 gnd.n448 gnd.n447 585
R1253 gnd.n7215 gnd.n7214 585
R1254 gnd.n7214 gnd.n7213 585
R1255 gnd.n452 gnd.n451 585
R1256 gnd.n7212 gnd.n452 585
R1257 gnd.n7210 gnd.n7209 585
R1258 gnd.n7211 gnd.n7210 585
R1259 gnd.n455 gnd.n454 585
R1260 gnd.n454 gnd.n453 585
R1261 gnd.n7205 gnd.n7204 585
R1262 gnd.n7204 gnd.n7203 585
R1263 gnd.n458 gnd.n457 585
R1264 gnd.n7202 gnd.n458 585
R1265 gnd.n7200 gnd.n7199 585
R1266 gnd.n7201 gnd.n7200 585
R1267 gnd.n461 gnd.n460 585
R1268 gnd.n460 gnd.n459 585
R1269 gnd.n7195 gnd.n7194 585
R1270 gnd.n7194 gnd.n7193 585
R1271 gnd.n464 gnd.n463 585
R1272 gnd.n7192 gnd.n464 585
R1273 gnd.n7190 gnd.n7189 585
R1274 gnd.n7191 gnd.n7190 585
R1275 gnd.n467 gnd.n466 585
R1276 gnd.n466 gnd.n465 585
R1277 gnd.n7185 gnd.n7184 585
R1278 gnd.n7184 gnd.n7183 585
R1279 gnd.n470 gnd.n469 585
R1280 gnd.n7182 gnd.n470 585
R1281 gnd.n7180 gnd.n7179 585
R1282 gnd.n7181 gnd.n7180 585
R1283 gnd.n473 gnd.n472 585
R1284 gnd.n472 gnd.n471 585
R1285 gnd.n7175 gnd.n7174 585
R1286 gnd.n7174 gnd.n7173 585
R1287 gnd.n476 gnd.n475 585
R1288 gnd.n7172 gnd.n476 585
R1289 gnd.n7170 gnd.n7169 585
R1290 gnd.n7171 gnd.n7170 585
R1291 gnd.n479 gnd.n478 585
R1292 gnd.n478 gnd.n477 585
R1293 gnd.n7165 gnd.n7164 585
R1294 gnd.n7164 gnd.n7163 585
R1295 gnd.n482 gnd.n481 585
R1296 gnd.n7162 gnd.n482 585
R1297 gnd.n7160 gnd.n7159 585
R1298 gnd.n7161 gnd.n7160 585
R1299 gnd.n485 gnd.n484 585
R1300 gnd.n484 gnd.n483 585
R1301 gnd.n7155 gnd.n7154 585
R1302 gnd.n7154 gnd.n7153 585
R1303 gnd.n488 gnd.n487 585
R1304 gnd.n7152 gnd.n488 585
R1305 gnd.n7150 gnd.n7149 585
R1306 gnd.n7151 gnd.n7150 585
R1307 gnd.n491 gnd.n490 585
R1308 gnd.n490 gnd.n489 585
R1309 gnd.n7145 gnd.n7144 585
R1310 gnd.n7144 gnd.n7143 585
R1311 gnd.n494 gnd.n493 585
R1312 gnd.n7142 gnd.n494 585
R1313 gnd.n7140 gnd.n7139 585
R1314 gnd.n7141 gnd.n7140 585
R1315 gnd.n497 gnd.n496 585
R1316 gnd.n496 gnd.n495 585
R1317 gnd.n7135 gnd.n7134 585
R1318 gnd.n7134 gnd.n7133 585
R1319 gnd.n500 gnd.n499 585
R1320 gnd.n7132 gnd.n500 585
R1321 gnd.n7130 gnd.n7129 585
R1322 gnd.n7131 gnd.n7130 585
R1323 gnd.n503 gnd.n502 585
R1324 gnd.n502 gnd.n501 585
R1325 gnd.n7125 gnd.n7124 585
R1326 gnd.n7124 gnd.n7123 585
R1327 gnd.n506 gnd.n505 585
R1328 gnd.n7122 gnd.n506 585
R1329 gnd.n7120 gnd.n7119 585
R1330 gnd.n7121 gnd.n7120 585
R1331 gnd.n509 gnd.n508 585
R1332 gnd.n508 gnd.n507 585
R1333 gnd.n7115 gnd.n7114 585
R1334 gnd.n7114 gnd.n7113 585
R1335 gnd.n512 gnd.n511 585
R1336 gnd.n7112 gnd.n512 585
R1337 gnd.n7110 gnd.n7109 585
R1338 gnd.n7111 gnd.n7110 585
R1339 gnd.n515 gnd.n514 585
R1340 gnd.n514 gnd.n513 585
R1341 gnd.n7105 gnd.n7104 585
R1342 gnd.n7104 gnd.n7103 585
R1343 gnd.n518 gnd.n517 585
R1344 gnd.n7102 gnd.n518 585
R1345 gnd.n7100 gnd.n7099 585
R1346 gnd.n7101 gnd.n7100 585
R1347 gnd.n521 gnd.n520 585
R1348 gnd.n520 gnd.n519 585
R1349 gnd.n7095 gnd.n7094 585
R1350 gnd.n7094 gnd.n7093 585
R1351 gnd.n524 gnd.n523 585
R1352 gnd.n7092 gnd.n524 585
R1353 gnd.n7090 gnd.n7089 585
R1354 gnd.n7091 gnd.n7090 585
R1355 gnd.n527 gnd.n526 585
R1356 gnd.n526 gnd.n525 585
R1357 gnd.n4790 gnd.n4789 585
R1358 gnd.n4789 gnd.n4788 585
R1359 gnd.n4791 gnd.n1368 585
R1360 gnd.n3021 gnd.n1368 585
R1361 gnd.n4793 gnd.n4792 585
R1362 gnd.n4794 gnd.n4793 585
R1363 gnd.n1352 gnd.n1351 585
R1364 gnd.n3014 gnd.n1352 585
R1365 gnd.n4802 gnd.n4801 585
R1366 gnd.n4801 gnd.n4800 585
R1367 gnd.n4803 gnd.n1347 585
R1368 gnd.n3009 gnd.n1347 585
R1369 gnd.n4805 gnd.n4804 585
R1370 gnd.n4806 gnd.n4805 585
R1371 gnd.n1332 gnd.n1331 585
R1372 gnd.n3036 gnd.n1332 585
R1373 gnd.n4814 gnd.n4813 585
R1374 gnd.n4813 gnd.n4812 585
R1375 gnd.n4815 gnd.n1327 585
R1376 gnd.n3002 gnd.n1327 585
R1377 gnd.n4817 gnd.n4816 585
R1378 gnd.n4818 gnd.n4817 585
R1379 gnd.n1312 gnd.n1311 585
R1380 gnd.n2994 gnd.n1312 585
R1381 gnd.n4826 gnd.n4825 585
R1382 gnd.n4825 gnd.n4824 585
R1383 gnd.n4827 gnd.n1307 585
R1384 gnd.n2987 gnd.n1307 585
R1385 gnd.n4829 gnd.n4828 585
R1386 gnd.n4830 gnd.n4829 585
R1387 gnd.n1292 gnd.n1291 585
R1388 gnd.n2979 gnd.n1292 585
R1389 gnd.n4838 gnd.n4837 585
R1390 gnd.n4837 gnd.n4836 585
R1391 gnd.n4839 gnd.n1287 585
R1392 gnd.n2925 gnd.n1287 585
R1393 gnd.n4841 gnd.n4840 585
R1394 gnd.n4842 gnd.n4841 585
R1395 gnd.n1273 gnd.n1272 585
R1396 gnd.n2916 gnd.n1273 585
R1397 gnd.n4850 gnd.n4849 585
R1398 gnd.n4849 gnd.n4848 585
R1399 gnd.n4851 gnd.n1267 585
R1400 gnd.n2910 gnd.n1267 585
R1401 gnd.n4853 gnd.n4852 585
R1402 gnd.n4854 gnd.n4853 585
R1403 gnd.n1268 gnd.n1266 585
R1404 gnd.n2939 gnd.n1266 585
R1405 gnd.n2905 gnd.n2904 585
R1406 gnd.n2904 gnd.n2903 585
R1407 gnd.n2610 gnd.n2609 585
R1408 gnd.n2898 gnd.n2610 585
R1409 gnd.n2880 gnd.n2879 585
R1410 gnd.n2879 gnd.n2878 585
R1411 gnd.n2881 gnd.n2622 585
R1412 gnd.n2889 gnd.n2622 585
R1413 gnd.n2883 gnd.n2882 585
R1414 gnd.n2884 gnd.n2883 585
R1415 gnd.n2629 gnd.n2628 585
R1416 gnd.n2852 gnd.n2628 585
R1417 gnd.n2858 gnd.n2857 585
R1418 gnd.n2860 gnd.n2858 585
R1419 gnd.n1244 gnd.n1243 585
R1420 gnd.n2640 gnd.n1244 585
R1421 gnd.n4864 gnd.n4863 585
R1422 gnd.n4863 gnd.n4862 585
R1423 gnd.n4865 gnd.n1239 585
R1424 gnd.n2841 gnd.n1239 585
R1425 gnd.n4867 gnd.n4866 585
R1426 gnd.n4868 gnd.n4867 585
R1427 gnd.n1223 gnd.n1222 585
R1428 gnd.n2834 gnd.n1223 585
R1429 gnd.n4876 gnd.n4875 585
R1430 gnd.n4875 gnd.n4874 585
R1431 gnd.n4877 gnd.n1218 585
R1432 gnd.n2825 gnd.n1218 585
R1433 gnd.n4879 gnd.n4878 585
R1434 gnd.n4880 gnd.n4879 585
R1435 gnd.n1203 gnd.n1202 585
R1436 gnd.n2819 gnd.n1203 585
R1437 gnd.n4888 gnd.n4887 585
R1438 gnd.n4887 gnd.n4886 585
R1439 gnd.n4889 gnd.n1198 585
R1440 gnd.n2772 gnd.n1198 585
R1441 gnd.n4891 gnd.n4890 585
R1442 gnd.n4892 gnd.n4891 585
R1443 gnd.n1183 gnd.n1182 585
R1444 gnd.n2766 gnd.n1183 585
R1445 gnd.n4900 gnd.n4899 585
R1446 gnd.n4899 gnd.n4898 585
R1447 gnd.n4901 gnd.n1178 585
R1448 gnd.n1178 gnd.n1177 585
R1449 gnd.n4903 gnd.n4902 585
R1450 gnd.n4904 gnd.n4903 585
R1451 gnd.n1164 gnd.n1163 585
R1452 gnd.n1167 gnd.n1164 585
R1453 gnd.n4912 gnd.n4911 585
R1454 gnd.n4911 gnd.n4910 585
R1455 gnd.n4913 gnd.n1157 585
R1456 gnd.n1157 gnd.n1155 585
R1457 gnd.n4915 gnd.n4914 585
R1458 gnd.n4916 gnd.n4915 585
R1459 gnd.n1159 gnd.n1156 585
R1460 gnd.n1156 gnd.n1152 585
R1461 gnd.n1158 gnd.n1143 585
R1462 gnd.n4922 gnd.n1143 585
R1463 gnd.n2699 gnd.n1137 585
R1464 gnd.n2699 gnd.n1068 585
R1465 gnd.n2701 gnd.n2700 585
R1466 gnd.n2703 gnd.n2702 585
R1467 gnd.n2705 gnd.n2704 585
R1468 gnd.n2709 gnd.n2697 585
R1469 gnd.n2711 gnd.n2710 585
R1470 gnd.n2713 gnd.n2712 585
R1471 gnd.n2715 gnd.n2714 585
R1472 gnd.n2719 gnd.n2695 585
R1473 gnd.n2721 gnd.n2720 585
R1474 gnd.n2723 gnd.n2722 585
R1475 gnd.n2725 gnd.n2724 585
R1476 gnd.n2729 gnd.n2693 585
R1477 gnd.n2731 gnd.n2730 585
R1478 gnd.n2733 gnd.n2732 585
R1479 gnd.n2735 gnd.n2734 585
R1480 gnd.n2690 gnd.n2689 585
R1481 gnd.n2739 gnd.n2691 585
R1482 gnd.n2740 gnd.n2686 585
R1483 gnd.n2741 gnd.n1067 585
R1484 gnd.n5046 gnd.n1067 585
R1485 gnd.n3079 gnd.n3078 585
R1486 gnd.n3080 gnd.n2525 585
R1487 gnd.n3081 gnd.n2521 585
R1488 gnd.n2519 gnd.n2511 585
R1489 gnd.n3088 gnd.n2510 585
R1490 gnd.n3089 gnd.n2508 585
R1491 gnd.n2507 gnd.n2500 585
R1492 gnd.n3096 gnd.n2499 585
R1493 gnd.n3097 gnd.n2498 585
R1494 gnd.n2496 gnd.n2490 585
R1495 gnd.n3104 gnd.n2489 585
R1496 gnd.n3105 gnd.n2487 585
R1497 gnd.n2486 gnd.n2479 585
R1498 gnd.n3112 gnd.n2478 585
R1499 gnd.n3113 gnd.n2477 585
R1500 gnd.n2475 gnd.n2469 585
R1501 gnd.n3120 gnd.n2468 585
R1502 gnd.n3121 gnd.n2466 585
R1503 gnd.n2465 gnd.n1372 585
R1504 gnd.n1381 gnd.n1372 585
R1505 gnd.n3023 gnd.n1375 585
R1506 gnd.n4788 gnd.n1375 585
R1507 gnd.n3024 gnd.n3022 585
R1508 gnd.n3022 gnd.n3021 585
R1509 gnd.n2574 gnd.n1366 585
R1510 gnd.n4794 gnd.n1366 585
R1511 gnd.n3028 gnd.n2573 585
R1512 gnd.n3014 gnd.n2573 585
R1513 gnd.n3029 gnd.n1355 585
R1514 gnd.n4800 gnd.n1355 585
R1515 gnd.n3030 gnd.n2572 585
R1516 gnd.n3009 gnd.n2572 585
R1517 gnd.n2569 gnd.n1345 585
R1518 gnd.n4806 gnd.n1345 585
R1519 gnd.n3035 gnd.n3034 585
R1520 gnd.n3036 gnd.n3035 585
R1521 gnd.n2568 gnd.n1335 585
R1522 gnd.n4812 gnd.n1335 585
R1523 gnd.n3001 gnd.n3000 585
R1524 gnd.n3002 gnd.n3001 585
R1525 gnd.n2577 gnd.n1325 585
R1526 gnd.n4818 gnd.n1325 585
R1527 gnd.n2996 gnd.n2995 585
R1528 gnd.n2995 gnd.n2994 585
R1529 gnd.n2579 gnd.n1315 585
R1530 gnd.n4824 gnd.n1315 585
R1531 gnd.n2986 gnd.n2985 585
R1532 gnd.n2987 gnd.n2986 585
R1533 gnd.n2582 gnd.n1305 585
R1534 gnd.n4830 gnd.n1305 585
R1535 gnd.n2981 gnd.n2980 585
R1536 gnd.n2980 gnd.n2979 585
R1537 gnd.n2584 gnd.n1295 585
R1538 gnd.n4836 gnd.n1295 585
R1539 gnd.n2927 gnd.n2926 585
R1540 gnd.n2926 gnd.n2925 585
R1541 gnd.n2606 gnd.n1285 585
R1542 gnd.n4842 gnd.n1285 585
R1543 gnd.n2931 gnd.n2605 585
R1544 gnd.n2916 gnd.n2605 585
R1545 gnd.n2932 gnd.n1276 585
R1546 gnd.n4848 gnd.n1276 585
R1547 gnd.n2933 gnd.n2604 585
R1548 gnd.n2910 gnd.n2604 585
R1549 gnd.n2601 gnd.n1264 585
R1550 gnd.n4854 gnd.n1264 585
R1551 gnd.n2938 gnd.n2937 585
R1552 gnd.n2939 gnd.n2938 585
R1553 gnd.n2600 gnd.n2599 585
R1554 gnd.n2903 gnd.n2599 585
R1555 gnd.n2897 gnd.n2896 585
R1556 gnd.n2898 gnd.n2897 585
R1557 gnd.n2616 gnd.n2615 585
R1558 gnd.n2878 gnd.n2615 585
R1559 gnd.n2891 gnd.n2890 585
R1560 gnd.n2890 gnd.n2889 585
R1561 gnd.n2619 gnd.n2618 585
R1562 gnd.n2884 gnd.n2619 585
R1563 gnd.n2851 gnd.n2850 585
R1564 gnd.n2852 gnd.n2851 585
R1565 gnd.n2652 gnd.n2642 585
R1566 gnd.n2860 gnd.n2642 585
R1567 gnd.n2846 gnd.n2845 585
R1568 gnd.n2845 gnd.n2640 585
R1569 gnd.n2844 gnd.n1247 585
R1570 gnd.n4862 gnd.n1247 585
R1571 gnd.n2843 gnd.n2842 585
R1572 gnd.n2842 gnd.n2841 585
R1573 gnd.n2654 gnd.n1237 585
R1574 gnd.n4868 gnd.n1237 585
R1575 gnd.n2833 gnd.n2832 585
R1576 gnd.n2834 gnd.n2833 585
R1577 gnd.n2658 gnd.n1226 585
R1578 gnd.n4874 gnd.n1226 585
R1579 gnd.n2827 gnd.n2826 585
R1580 gnd.n2826 gnd.n2825 585
R1581 gnd.n2660 gnd.n1216 585
R1582 gnd.n4880 gnd.n1216 585
R1583 gnd.n2779 gnd.n2778 585
R1584 gnd.n2819 gnd.n2779 585
R1585 gnd.n2663 gnd.n1206 585
R1586 gnd.n4886 gnd.n1206 585
R1587 gnd.n2774 gnd.n2773 585
R1588 gnd.n2773 gnd.n2772 585
R1589 gnd.n2665 gnd.n1196 585
R1590 gnd.n4892 gnd.n1196 585
R1591 gnd.n2765 gnd.n2764 585
R1592 gnd.n2766 gnd.n2765 585
R1593 gnd.n2680 gnd.n1186 585
R1594 gnd.n4898 gnd.n1186 585
R1595 gnd.n2760 gnd.n2759 585
R1596 gnd.n2759 gnd.n1177 585
R1597 gnd.n2758 gnd.n1176 585
R1598 gnd.n4904 gnd.n1176 585
R1599 gnd.n2757 gnd.n2756 585
R1600 gnd.n2756 gnd.n1167 585
R1601 gnd.n2682 gnd.n1166 585
R1602 gnd.n4910 gnd.n1166 585
R1603 gnd.n2752 gnd.n2751 585
R1604 gnd.n2751 gnd.n1155 585
R1605 gnd.n2750 gnd.n1154 585
R1606 gnd.n4916 gnd.n1154 585
R1607 gnd.n2749 gnd.n2748 585
R1608 gnd.n2748 gnd.n1152 585
R1609 gnd.n2684 gnd.n1142 585
R1610 gnd.n4922 gnd.n1142 585
R1611 gnd.n2744 gnd.n2743 585
R1612 gnd.n2743 gnd.n1068 585
R1613 gnd.n6430 gnd.n6429 585
R1614 gnd.n6429 gnd.n6428 585
R1615 gnd.n6431 gnd.n1021 585
R1616 gnd.n6338 gnd.n1021 585
R1617 gnd.n6433 gnd.n6432 585
R1618 gnd.n6434 gnd.n6433 585
R1619 gnd.n1022 gnd.n1020 585
R1620 gnd.n1020 gnd.n1016 585
R1621 gnd.n1001 gnd.n1000 585
R1622 gnd.n1005 gnd.n1001 585
R1623 gnd.n6444 gnd.n6443 585
R1624 gnd.n6443 gnd.n6442 585
R1625 gnd.n6445 gnd.n995 585
R1626 gnd.n6327 gnd.n995 585
R1627 gnd.n6447 gnd.n6446 585
R1628 gnd.n6448 gnd.n6447 585
R1629 gnd.n996 gnd.n994 585
R1630 gnd.n994 gnd.n990 585
R1631 gnd.n978 gnd.n977 585
R1632 gnd.n6320 gnd.n978 585
R1633 gnd.n6458 gnd.n6457 585
R1634 gnd.n6457 gnd.n6456 585
R1635 gnd.n6459 gnd.n972 585
R1636 gnd.n5983 gnd.n972 585
R1637 gnd.n6461 gnd.n6460 585
R1638 gnd.n6462 gnd.n6461 585
R1639 gnd.n973 gnd.n971 585
R1640 gnd.n5145 gnd.n971 585
R1641 gnd.n6021 gnd.n6020 585
R1642 gnd.n6020 gnd.n6019 585
R1643 gnd.n5143 gnd.n5142 585
R1644 gnd.n6003 gnd.n5143 585
R1645 gnd.n5995 gnd.n5994 585
R1646 gnd.n5994 gnd.n5993 585
R1647 gnd.n5157 gnd.n5156 585
R1648 gnd.n5165 gnd.n5157 585
R1649 gnd.n5969 gnd.n5968 585
R1650 gnd.n5970 gnd.n5969 585
R1651 gnd.n5168 gnd.n5167 585
R1652 gnd.n5175 gnd.n5167 585
R1653 gnd.n5943 gnd.n5187 585
R1654 gnd.n5187 gnd.n5174 585
R1655 gnd.n5945 gnd.n5944 585
R1656 gnd.n5946 gnd.n5945 585
R1657 gnd.n5188 gnd.n5186 585
R1658 gnd.n5186 gnd.n5182 585
R1659 gnd.n5932 gnd.n5931 585
R1660 gnd.n5931 gnd.n5930 585
R1661 gnd.n5193 gnd.n5192 585
R1662 gnd.n5203 gnd.n5193 585
R1663 gnd.n5921 gnd.n5920 585
R1664 gnd.n5920 gnd.n5919 585
R1665 gnd.n5200 gnd.n5199 585
R1666 gnd.n5907 gnd.n5200 585
R1667 gnd.n5881 gnd.n5285 585
R1668 gnd.n5285 gnd.n5210 585
R1669 gnd.n5883 gnd.n5882 585
R1670 gnd.n5884 gnd.n5883 585
R1671 gnd.n5286 gnd.n5284 585
R1672 gnd.n5294 gnd.n5284 585
R1673 gnd.n5859 gnd.n5306 585
R1674 gnd.n5306 gnd.n5293 585
R1675 gnd.n5861 gnd.n5860 585
R1676 gnd.n5862 gnd.n5861 585
R1677 gnd.n5307 gnd.n5305 585
R1678 gnd.n5305 gnd.n5301 585
R1679 gnd.n5847 gnd.n5846 585
R1680 gnd.n5846 gnd.n5845 585
R1681 gnd.n5312 gnd.n5311 585
R1682 gnd.n5321 gnd.n5312 585
R1683 gnd.n5836 gnd.n5835 585
R1684 gnd.n5835 gnd.n5834 585
R1685 gnd.n5319 gnd.n5318 585
R1686 gnd.n5822 gnd.n5319 585
R1687 gnd.n5794 gnd.n5793 585
R1688 gnd.n5793 gnd.n5328 585
R1689 gnd.n5795 gnd.n5339 585
R1690 gnd.n5786 gnd.n5339 585
R1691 gnd.n5797 gnd.n5796 585
R1692 gnd.n5798 gnd.n5797 585
R1693 gnd.n5340 gnd.n5338 585
R1694 gnd.n5354 gnd.n5338 585
R1695 gnd.n5778 gnd.n5777 585
R1696 gnd.n5777 gnd.n5776 585
R1697 gnd.n5351 gnd.n5350 585
R1698 gnd.n5761 gnd.n5351 585
R1699 gnd.n5748 gnd.n5371 585
R1700 gnd.n5371 gnd.n5361 585
R1701 gnd.n5750 gnd.n5749 585
R1702 gnd.n5751 gnd.n5750 585
R1703 gnd.n5372 gnd.n5370 585
R1704 gnd.n5380 gnd.n5370 585
R1705 gnd.n5724 gnd.n5392 585
R1706 gnd.n5392 gnd.n5379 585
R1707 gnd.n5726 gnd.n5725 585
R1708 gnd.n5727 gnd.n5726 585
R1709 gnd.n5393 gnd.n5391 585
R1710 gnd.n5391 gnd.n5387 585
R1711 gnd.n5712 gnd.n5711 585
R1712 gnd.n5711 gnd.n5710 585
R1713 gnd.n5398 gnd.n5397 585
R1714 gnd.n5402 gnd.n5398 585
R1715 gnd.n5696 gnd.n5695 585
R1716 gnd.n5697 gnd.n5696 585
R1717 gnd.n5413 gnd.n5412 585
R1718 gnd.n5412 gnd.n5408 585
R1719 gnd.n5686 gnd.n5685 585
R1720 gnd.n5687 gnd.n5686 585
R1721 gnd.n5422 gnd.n5421 585
R1722 gnd.n5421 gnd.n5419 585
R1723 gnd.n5680 gnd.n5679 585
R1724 gnd.n5679 gnd.n5678 585
R1725 gnd.n5426 gnd.n5425 585
R1726 gnd.n5434 gnd.n5426 585
R1727 gnd.n5587 gnd.n5586 585
R1728 gnd.n5588 gnd.n5587 585
R1729 gnd.n5436 gnd.n5435 585
R1730 gnd.n5435 gnd.n5433 585
R1731 gnd.n5582 gnd.n5581 585
R1732 gnd.n5581 gnd.n5580 585
R1733 gnd.n5439 gnd.n5438 585
R1734 gnd.n5440 gnd.n5439 585
R1735 gnd.n5571 gnd.n5570 585
R1736 gnd.n5572 gnd.n5571 585
R1737 gnd.n5448 gnd.n5447 585
R1738 gnd.n5447 gnd.n5446 585
R1739 gnd.n5566 gnd.n5565 585
R1740 gnd.n5565 gnd.n5564 585
R1741 gnd.n5451 gnd.n5450 585
R1742 gnd.n5452 gnd.n5451 585
R1743 gnd.n5555 gnd.n5554 585
R1744 gnd.n5556 gnd.n5555 585
R1745 gnd.n5551 gnd.n5458 585
R1746 gnd.n5550 gnd.n5549 585
R1747 gnd.n5547 gnd.n5460 585
R1748 gnd.n5547 gnd.n5457 585
R1749 gnd.n5546 gnd.n5545 585
R1750 gnd.n5544 gnd.n5543 585
R1751 gnd.n5542 gnd.n5465 585
R1752 gnd.n5540 gnd.n5539 585
R1753 gnd.n5538 gnd.n5466 585
R1754 gnd.n5537 gnd.n5536 585
R1755 gnd.n5534 gnd.n5471 585
R1756 gnd.n5532 gnd.n5531 585
R1757 gnd.n5530 gnd.n5472 585
R1758 gnd.n5529 gnd.n5528 585
R1759 gnd.n5526 gnd.n5477 585
R1760 gnd.n5524 gnd.n5523 585
R1761 gnd.n5522 gnd.n5478 585
R1762 gnd.n5521 gnd.n5520 585
R1763 gnd.n5518 gnd.n5483 585
R1764 gnd.n5516 gnd.n5515 585
R1765 gnd.n5514 gnd.n5484 585
R1766 gnd.n5513 gnd.n5512 585
R1767 gnd.n5510 gnd.n5489 585
R1768 gnd.n5508 gnd.n5507 585
R1769 gnd.n5505 gnd.n5490 585
R1770 gnd.n5504 gnd.n5503 585
R1771 gnd.n5501 gnd.n5499 585
R1772 gnd.n5497 gnd.n5456 585
R1773 gnd.n6346 gnd.n6345 585
R1774 gnd.n6347 gnd.n5126 585
R1775 gnd.n6349 gnd.n6348 585
R1776 gnd.n6351 gnd.n5125 585
R1777 gnd.n6353 gnd.n6352 585
R1778 gnd.n6354 gnd.n5116 585
R1779 gnd.n6356 gnd.n6355 585
R1780 gnd.n6358 gnd.n5114 585
R1781 gnd.n6360 gnd.n6359 585
R1782 gnd.n6361 gnd.n5109 585
R1783 gnd.n6363 gnd.n6362 585
R1784 gnd.n6365 gnd.n5107 585
R1785 gnd.n6367 gnd.n6366 585
R1786 gnd.n6368 gnd.n5102 585
R1787 gnd.n6370 gnd.n6369 585
R1788 gnd.n6372 gnd.n5100 585
R1789 gnd.n6374 gnd.n6373 585
R1790 gnd.n6375 gnd.n5095 585
R1791 gnd.n6377 gnd.n6376 585
R1792 gnd.n6379 gnd.n5093 585
R1793 gnd.n6381 gnd.n6380 585
R1794 gnd.n6382 gnd.n5088 585
R1795 gnd.n6384 gnd.n6383 585
R1796 gnd.n6386 gnd.n5086 585
R1797 gnd.n6388 gnd.n6387 585
R1798 gnd.n6389 gnd.n5084 585
R1799 gnd.n6390 gnd.n1026 585
R1800 gnd.n5047 gnd.n1026 585
R1801 gnd.n6341 gnd.n1028 585
R1802 gnd.n6428 gnd.n1028 585
R1803 gnd.n6340 gnd.n6339 585
R1804 gnd.n6339 gnd.n6338 585
R1805 gnd.n6337 gnd.n1018 585
R1806 gnd.n6434 gnd.n1018 585
R1807 gnd.n6331 gnd.n5131 585
R1808 gnd.n6331 gnd.n1016 585
R1809 gnd.n6333 gnd.n6332 585
R1810 gnd.n6332 gnd.n1005 585
R1811 gnd.n6330 gnd.n1003 585
R1812 gnd.n6442 gnd.n1003 585
R1813 gnd.n6329 gnd.n6328 585
R1814 gnd.n6328 gnd.n6327 585
R1815 gnd.n5133 gnd.n992 585
R1816 gnd.n6448 gnd.n992 585
R1817 gnd.n6323 gnd.n6322 585
R1818 gnd.n6322 gnd.n990 585
R1819 gnd.n6321 gnd.n5135 585
R1820 gnd.n6321 gnd.n6320 585
R1821 gnd.n5982 gnd.n980 585
R1822 gnd.n6456 gnd.n980 585
R1823 gnd.n5985 gnd.n5984 585
R1824 gnd.n5984 gnd.n5983 585
R1825 gnd.n5986 gnd.n969 585
R1826 gnd.n6462 gnd.n969 585
R1827 gnd.n5988 gnd.n5987 585
R1828 gnd.n5987 gnd.n5145 585
R1829 gnd.n5989 gnd.n5144 585
R1830 gnd.n6019 gnd.n5144 585
R1831 gnd.n5990 gnd.n5153 585
R1832 gnd.n6003 gnd.n5153 585
R1833 gnd.n5992 gnd.n5991 585
R1834 gnd.n5993 gnd.n5992 585
R1835 gnd.n5160 gnd.n5159 585
R1836 gnd.n5165 gnd.n5159 585
R1837 gnd.n5972 gnd.n5971 585
R1838 gnd.n5971 gnd.n5970 585
R1839 gnd.n5163 gnd.n5162 585
R1840 gnd.n5175 gnd.n5163 585
R1841 gnd.n5897 gnd.n5896 585
R1842 gnd.n5896 gnd.n5174 585
R1843 gnd.n5898 gnd.n5184 585
R1844 gnd.n5946 gnd.n5184 585
R1845 gnd.n5900 gnd.n5899 585
R1846 gnd.n5899 gnd.n5182 585
R1847 gnd.n5901 gnd.n5195 585
R1848 gnd.n5930 gnd.n5195 585
R1849 gnd.n5903 gnd.n5902 585
R1850 gnd.n5902 gnd.n5203 585
R1851 gnd.n5904 gnd.n5202 585
R1852 gnd.n5919 gnd.n5202 585
R1853 gnd.n5906 gnd.n5905 585
R1854 gnd.n5907 gnd.n5906 585
R1855 gnd.n5214 gnd.n5213 585
R1856 gnd.n5213 gnd.n5210 585
R1857 gnd.n5886 gnd.n5885 585
R1858 gnd.n5885 gnd.n5884 585
R1859 gnd.n5281 gnd.n5280 585
R1860 gnd.n5294 gnd.n5281 585
R1861 gnd.n5807 gnd.n5806 585
R1862 gnd.n5806 gnd.n5293 585
R1863 gnd.n5808 gnd.n5303 585
R1864 gnd.n5862 gnd.n5303 585
R1865 gnd.n5811 gnd.n5810 585
R1866 gnd.n5810 gnd.n5301 585
R1867 gnd.n5812 gnd.n5314 585
R1868 gnd.n5845 gnd.n5314 585
R1869 gnd.n5815 gnd.n5814 585
R1870 gnd.n5814 gnd.n5321 585
R1871 gnd.n5816 gnd.n5320 585
R1872 gnd.n5834 gnd.n5320 585
R1873 gnd.n5819 gnd.n5818 585
R1874 gnd.n5822 gnd.n5819 585
R1875 gnd.n5804 gnd.n5330 585
R1876 gnd.n5330 gnd.n5328 585
R1877 gnd.n5335 gnd.n5331 585
R1878 gnd.n5786 gnd.n5335 585
R1879 gnd.n5800 gnd.n5799 585
R1880 gnd.n5799 gnd.n5798 585
R1881 gnd.n5334 gnd.n5333 585
R1882 gnd.n5354 gnd.n5334 585
R1883 gnd.n5758 gnd.n5353 585
R1884 gnd.n5776 gnd.n5353 585
R1885 gnd.n5760 gnd.n5759 585
R1886 gnd.n5761 gnd.n5760 585
R1887 gnd.n5364 gnd.n5363 585
R1888 gnd.n5363 gnd.n5361 585
R1889 gnd.n5753 gnd.n5752 585
R1890 gnd.n5752 gnd.n5751 585
R1891 gnd.n5367 gnd.n5366 585
R1892 gnd.n5380 gnd.n5367 585
R1893 gnd.n5604 gnd.n5603 585
R1894 gnd.n5603 gnd.n5379 585
R1895 gnd.n5605 gnd.n5389 585
R1896 gnd.n5727 gnd.n5389 585
R1897 gnd.n5607 gnd.n5606 585
R1898 gnd.n5606 gnd.n5387 585
R1899 gnd.n5608 gnd.n5399 585
R1900 gnd.n5710 gnd.n5399 585
R1901 gnd.n5610 gnd.n5609 585
R1902 gnd.n5609 gnd.n5402 585
R1903 gnd.n5611 gnd.n5410 585
R1904 gnd.n5697 gnd.n5410 585
R1905 gnd.n5613 gnd.n5612 585
R1906 gnd.n5612 gnd.n5408 585
R1907 gnd.n5614 gnd.n5420 585
R1908 gnd.n5687 gnd.n5420 585
R1909 gnd.n5615 gnd.n5428 585
R1910 gnd.n5428 gnd.n5419 585
R1911 gnd.n5617 gnd.n5616 585
R1912 gnd.n5678 gnd.n5617 585
R1913 gnd.n5429 gnd.n5427 585
R1914 gnd.n5434 gnd.n5427 585
R1915 gnd.n5590 gnd.n5589 585
R1916 gnd.n5589 gnd.n5588 585
R1917 gnd.n5432 gnd.n5431 585
R1918 gnd.n5433 gnd.n5432 585
R1919 gnd.n5579 gnd.n5578 585
R1920 gnd.n5580 gnd.n5579 585
R1921 gnd.n5442 gnd.n5441 585
R1922 gnd.n5441 gnd.n5440 585
R1923 gnd.n5574 gnd.n5573 585
R1924 gnd.n5573 gnd.n5572 585
R1925 gnd.n5445 gnd.n5444 585
R1926 gnd.n5446 gnd.n5445 585
R1927 gnd.n5563 gnd.n5562 585
R1928 gnd.n5564 gnd.n5563 585
R1929 gnd.n5454 gnd.n5453 585
R1930 gnd.n5453 gnd.n5452 585
R1931 gnd.n5558 gnd.n5557 585
R1932 gnd.n5557 gnd.n5556 585
R1933 gnd.n7559 gnd.n7558 585
R1934 gnd.n7558 gnd.n7557 585
R1935 gnd.n7560 gnd.n204 585
R1936 gnd.n209 gnd.n204 585
R1937 gnd.n7562 gnd.n7561 585
R1938 gnd.n7563 gnd.n7562 585
R1939 gnd.n191 gnd.n190 585
R1940 gnd.n194 gnd.n191 585
R1941 gnd.n7571 gnd.n7570 585
R1942 gnd.n7570 gnd.n7569 585
R1943 gnd.n7572 gnd.n186 585
R1944 gnd.n186 gnd.n185 585
R1945 gnd.n7574 gnd.n7573 585
R1946 gnd.n7575 gnd.n7574 585
R1947 gnd.n171 gnd.n170 585
R1948 gnd.n175 gnd.n171 585
R1949 gnd.n7583 gnd.n7582 585
R1950 gnd.n7582 gnd.n7581 585
R1951 gnd.n7584 gnd.n166 585
R1952 gnd.n7392 gnd.n166 585
R1953 gnd.n7586 gnd.n7585 585
R1954 gnd.n7587 gnd.n7586 585
R1955 gnd.n152 gnd.n151 585
R1956 gnd.n7371 gnd.n152 585
R1957 gnd.n7595 gnd.n7594 585
R1958 gnd.n7594 gnd.n7593 585
R1959 gnd.n7596 gnd.n147 585
R1960 gnd.n7362 gnd.n147 585
R1961 gnd.n7598 gnd.n7597 585
R1962 gnd.n7599 gnd.n7598 585
R1963 gnd.n131 gnd.n130 585
R1964 gnd.n7356 gnd.n131 585
R1965 gnd.n7607 gnd.n7606 585
R1966 gnd.n7606 gnd.n7605 585
R1967 gnd.n7608 gnd.n126 585
R1968 gnd.n7348 gnd.n126 585
R1969 gnd.n7610 gnd.n7609 585
R1970 gnd.n7611 gnd.n7610 585
R1971 gnd.n113 gnd.n112 585
R1972 gnd.n7342 gnd.n113 585
R1973 gnd.n7619 gnd.n7618 585
R1974 gnd.n7618 gnd.n7617 585
R1975 gnd.n7620 gnd.n107 585
R1976 gnd.n7334 gnd.n107 585
R1977 gnd.n7622 gnd.n7621 585
R1978 gnd.n7623 gnd.n7622 585
R1979 gnd.n108 gnd.n106 585
R1980 gnd.n7328 gnd.n106 585
R1981 gnd.n4431 gnd.n4430 585
R1982 gnd.n4430 gnd.n381 585
R1983 gnd.n4432 gnd.n88 585
R1984 gnd.n7631 gnd.n88 585
R1985 gnd.n4434 gnd.n4433 585
R1986 gnd.n4435 gnd.n4434 585
R1987 gnd.n4425 gnd.n4424 585
R1988 gnd.n4424 gnd.n1732 585
R1989 gnd.n1720 gnd.n1719 585
R1990 gnd.n4471 gnd.n1720 585
R1991 gnd.n4476 gnd.n4475 585
R1992 gnd.n4475 gnd.n4474 585
R1993 gnd.n4477 gnd.n1715 585
R1994 gnd.n4456 gnd.n1715 585
R1995 gnd.n4479 gnd.n4478 585
R1996 gnd.n4480 gnd.n4479 585
R1997 gnd.n1703 gnd.n1702 585
R1998 gnd.n4445 gnd.n1703 585
R1999 gnd.n4488 gnd.n4487 585
R2000 gnd.n4487 gnd.n4486 585
R2001 gnd.n4489 gnd.n1698 585
R2002 gnd.n4415 gnd.n1698 585
R2003 gnd.n4491 gnd.n4490 585
R2004 gnd.n4492 gnd.n4491 585
R2005 gnd.n1682 gnd.n1681 585
R2006 gnd.n4374 gnd.n1682 585
R2007 gnd.n4500 gnd.n4499 585
R2008 gnd.n4499 gnd.n4498 585
R2009 gnd.n4501 gnd.n1677 585
R2010 gnd.n4367 gnd.n1677 585
R2011 gnd.n4503 gnd.n4502 585
R2012 gnd.n4504 gnd.n4503 585
R2013 gnd.n1663 gnd.n1662 585
R2014 gnd.n4362 gnd.n1663 585
R2015 gnd.n4512 gnd.n4511 585
R2016 gnd.n4511 gnd.n4510 585
R2017 gnd.n4513 gnd.n1658 585
R2018 gnd.n4391 gnd.n1658 585
R2019 gnd.n4515 gnd.n4514 585
R2020 gnd.n4516 gnd.n4515 585
R2021 gnd.n1642 gnd.n1641 585
R2022 gnd.n4355 gnd.n1642 585
R2023 gnd.n4524 gnd.n4523 585
R2024 gnd.n4523 gnd.n4522 585
R2025 gnd.n4525 gnd.n1637 585
R2026 gnd.n4347 gnd.n1637 585
R2027 gnd.n4527 gnd.n4526 585
R2028 gnd.n4528 gnd.n4527 585
R2029 gnd.n1622 gnd.n1621 585
R2030 gnd.n4341 gnd.n1622 585
R2031 gnd.n4536 gnd.n4535 585
R2032 gnd.n4535 gnd.n4534 585
R2033 gnd.n4537 gnd.n1616 585
R2034 gnd.n4333 gnd.n1616 585
R2035 gnd.n4539 gnd.n4538 585
R2036 gnd.n4540 gnd.n4539 585
R2037 gnd.n1617 gnd.n1615 585
R2038 gnd.n3754 gnd.n1615 585
R2039 gnd.n4326 gnd.n1603 585
R2040 gnd.n4546 gnd.n1603 585
R2041 gnd.n3841 gnd.n3840 585
R2042 gnd.n3804 gnd.n3803 585
R2043 gnd.n3855 gnd.n3854 585
R2044 gnd.n3857 gnd.n3802 585
R2045 gnd.n3860 gnd.n3859 585
R2046 gnd.n3795 gnd.n3794 585
R2047 gnd.n3874 gnd.n3873 585
R2048 gnd.n3876 gnd.n3793 585
R2049 gnd.n3879 gnd.n3878 585
R2050 gnd.n3786 gnd.n3785 585
R2051 gnd.n3893 gnd.n3892 585
R2052 gnd.n3895 gnd.n3784 585
R2053 gnd.n3898 gnd.n3897 585
R2054 gnd.n3777 gnd.n3776 585
R2055 gnd.n3913 gnd.n3912 585
R2056 gnd.n3915 gnd.n3775 585
R2057 gnd.n3918 gnd.n3917 585
R2058 gnd.n3919 gnd.n3772 585
R2059 gnd.n3771 gnd.n3770 585
R2060 gnd.n3771 gnd.n1591 585
R2061 gnd.n349 gnd.n348 585
R2062 gnd.n7413 gnd.n344 585
R2063 gnd.n7415 gnd.n7414 585
R2064 gnd.n7417 gnd.n342 585
R2065 gnd.n7419 gnd.n7418 585
R2066 gnd.n7420 gnd.n337 585
R2067 gnd.n7422 gnd.n7421 585
R2068 gnd.n7424 gnd.n335 585
R2069 gnd.n7426 gnd.n7425 585
R2070 gnd.n7427 gnd.n330 585
R2071 gnd.n7429 gnd.n7428 585
R2072 gnd.n7431 gnd.n328 585
R2073 gnd.n7433 gnd.n7432 585
R2074 gnd.n7434 gnd.n323 585
R2075 gnd.n7436 gnd.n7435 585
R2076 gnd.n7438 gnd.n321 585
R2077 gnd.n7440 gnd.n7439 585
R2078 gnd.n7441 gnd.n319 585
R2079 gnd.n7442 gnd.n208 585
R2080 gnd.n212 gnd.n208 585
R2081 gnd.n7409 gnd.n211 585
R2082 gnd.n7557 gnd.n211 585
R2083 gnd.n7408 gnd.n7407 585
R2084 gnd.n7407 gnd.n209 585
R2085 gnd.n7406 gnd.n203 585
R2086 gnd.n7563 gnd.n203 585
R2087 gnd.n354 gnd.n353 585
R2088 gnd.n353 gnd.n194 585
R2089 gnd.n7402 gnd.n193 585
R2090 gnd.n7569 gnd.n193 585
R2091 gnd.n7401 gnd.n7400 585
R2092 gnd.n7400 gnd.n185 585
R2093 gnd.n7399 gnd.n184 585
R2094 gnd.n7575 gnd.n184 585
R2095 gnd.n357 gnd.n356 585
R2096 gnd.n356 gnd.n175 585
R2097 gnd.n7395 gnd.n174 585
R2098 gnd.n7581 gnd.n174 585
R2099 gnd.n7394 gnd.n7393 585
R2100 gnd.n7393 gnd.n7392 585
R2101 gnd.n359 gnd.n165 585
R2102 gnd.n7587 gnd.n165 585
R2103 gnd.n7370 gnd.n7369 585
R2104 gnd.n7371 gnd.n7370 585
R2105 gnd.n363 gnd.n155 585
R2106 gnd.n7593 gnd.n155 585
R2107 gnd.n7364 gnd.n7363 585
R2108 gnd.n7363 gnd.n7362 585
R2109 gnd.n365 gnd.n145 585
R2110 gnd.n7599 gnd.n145 585
R2111 gnd.n7355 gnd.n7354 585
R2112 gnd.n7356 gnd.n7355 585
R2113 gnd.n368 gnd.n134 585
R2114 gnd.n7605 gnd.n134 585
R2115 gnd.n7350 gnd.n7349 585
R2116 gnd.n7349 gnd.n7348 585
R2117 gnd.n370 gnd.n125 585
R2118 gnd.n7611 gnd.n125 585
R2119 gnd.n7341 gnd.n7340 585
R2120 gnd.n7342 gnd.n7341 585
R2121 gnd.n375 gnd.n116 585
R2122 gnd.n7617 gnd.n116 585
R2123 gnd.n7336 gnd.n7335 585
R2124 gnd.n7335 gnd.n7334 585
R2125 gnd.n377 gnd.n104 585
R2126 gnd.n7623 gnd.n104 585
R2127 gnd.n7327 gnd.n7326 585
R2128 gnd.n7328 gnd.n7327 585
R2129 gnd.n84 gnd.n83 585
R2130 gnd.n381 gnd.n84 585
R2131 gnd.n7633 gnd.n7632 585
R2132 gnd.n7632 gnd.n7631 585
R2133 gnd.n7634 gnd.n82 585
R2134 gnd.n4435 gnd.n82 585
R2135 gnd.n1731 gnd.n81 585
R2136 gnd.n1732 gnd.n1731 585
R2137 gnd.n4450 gnd.n1730 585
R2138 gnd.n4471 gnd.n1730 585
R2139 gnd.n1739 gnd.n1723 585
R2140 gnd.n4474 gnd.n1723 585
R2141 gnd.n4455 gnd.n4454 585
R2142 gnd.n4456 gnd.n4455 585
R2143 gnd.n1738 gnd.n1714 585
R2144 gnd.n4480 gnd.n1714 585
R2145 gnd.n4447 gnd.n4446 585
R2146 gnd.n4446 gnd.n4445 585
R2147 gnd.n1741 gnd.n1705 585
R2148 gnd.n4486 gnd.n1705 585
R2149 gnd.n4377 gnd.n1743 585
R2150 gnd.n4415 gnd.n1743 585
R2151 gnd.n4378 gnd.n1696 585
R2152 gnd.n4492 gnd.n1696 585
R2153 gnd.n4379 gnd.n4375 585
R2154 gnd.n4375 gnd.n4374 585
R2155 gnd.n1762 gnd.n1685 585
R2156 gnd.n4498 gnd.n1685 585
R2157 gnd.n4383 gnd.n1761 585
R2158 gnd.n4367 gnd.n1761 585
R2159 gnd.n4384 gnd.n1676 585
R2160 gnd.n4504 gnd.n1676 585
R2161 gnd.n4385 gnd.n1760 585
R2162 gnd.n4362 gnd.n1760 585
R2163 gnd.n1757 gnd.n1665 585
R2164 gnd.n4510 gnd.n1665 585
R2165 gnd.n4390 gnd.n4389 585
R2166 gnd.n4391 gnd.n4390 585
R2167 gnd.n1756 gnd.n1656 585
R2168 gnd.n4516 gnd.n1656 585
R2169 gnd.n4354 gnd.n4353 585
R2170 gnd.n4355 gnd.n4354 585
R2171 gnd.n1766 gnd.n1645 585
R2172 gnd.n4522 gnd.n1645 585
R2173 gnd.n4349 gnd.n4348 585
R2174 gnd.n4348 gnd.n4347 585
R2175 gnd.n1768 gnd.n1636 585
R2176 gnd.n4528 gnd.n1636 585
R2177 gnd.n4340 gnd.n4339 585
R2178 gnd.n4341 gnd.n4340 585
R2179 gnd.n1803 gnd.n1625 585
R2180 gnd.n4534 gnd.n1625 585
R2181 gnd.n4335 gnd.n4334 585
R2182 gnd.n4334 gnd.n4333 585
R2183 gnd.n1805 gnd.n1613 585
R2184 gnd.n4540 gnd.n1613 585
R2185 gnd.n3756 gnd.n3755 585
R2186 gnd.n3755 gnd.n3754 585
R2187 gnd.n3757 gnd.n1601 585
R2188 gnd.n4546 gnd.n1601 585
R2189 gnd.n6426 gnd.n6425 585
R2190 gnd.n6427 gnd.n6426 585
R2191 gnd.n5050 gnd.n5048 585
R2192 gnd.n5048 gnd.n1027 585
R2193 gnd.n1015 gnd.n1014 585
R2194 gnd.n1019 gnd.n1015 585
R2195 gnd.n6437 gnd.n6436 585
R2196 gnd.n6436 gnd.n6435 585
R2197 gnd.n6438 gnd.n1007 585
R2198 gnd.n6308 gnd.n1007 585
R2199 gnd.n6440 gnd.n6439 585
R2200 gnd.n6441 gnd.n6440 585
R2201 gnd.n1008 gnd.n1006 585
R2202 gnd.n1006 gnd.n1002 585
R2203 gnd.n989 gnd.n988 585
R2204 gnd.n993 gnd.n989 585
R2205 gnd.n6451 gnd.n6450 585
R2206 gnd.n6450 gnd.n6449 585
R2207 gnd.n6452 gnd.n983 585
R2208 gnd.n6319 gnd.n983 585
R2209 gnd.n6454 gnd.n6453 585
R2210 gnd.n6455 gnd.n6454 585
R2211 gnd.n984 gnd.n982 585
R2212 gnd.n982 gnd.n979 585
R2213 gnd.n6014 gnd.n6013 585
R2214 gnd.n6013 gnd.n970 585
R2215 gnd.n6015 gnd.n5147 585
R2216 gnd.n5147 gnd.n968 585
R2217 gnd.n6017 gnd.n6016 585
R2218 gnd.n6018 gnd.n6017 585
R2219 gnd.n5148 gnd.n5146 585
R2220 gnd.n6002 gnd.n5146 585
R2221 gnd.n6006 gnd.n6005 585
R2222 gnd.n6005 gnd.n6004 585
R2223 gnd.n5151 gnd.n5150 585
R2224 gnd.n5158 gnd.n5151 585
R2225 gnd.n5956 gnd.n5955 585
R2226 gnd.n5955 gnd.n5166 585
R2227 gnd.n5957 gnd.n5177 585
R2228 gnd.n5177 gnd.n5164 585
R2229 gnd.n5959 gnd.n5958 585
R2230 gnd.n5960 gnd.n5959 585
R2231 gnd.n5178 gnd.n5176 585
R2232 gnd.n5185 gnd.n5176 585
R2233 gnd.n5949 gnd.n5948 585
R2234 gnd.n5948 gnd.n5947 585
R2235 gnd.n5181 gnd.n5180 585
R2236 gnd.n5929 gnd.n5181 585
R2237 gnd.n5915 gnd.n5205 585
R2238 gnd.n5205 gnd.n5194 585
R2239 gnd.n5917 gnd.n5916 585
R2240 gnd.n5918 gnd.n5917 585
R2241 gnd.n5206 gnd.n5204 585
R2242 gnd.n5204 gnd.n5201 585
R2243 gnd.n5910 gnd.n5909 585
R2244 gnd.n5909 gnd.n5908 585
R2245 gnd.n5209 gnd.n5208 585
R2246 gnd.n5283 gnd.n5209 585
R2247 gnd.n5870 gnd.n5296 585
R2248 gnd.n5296 gnd.n5282 585
R2249 gnd.n5872 gnd.n5871 585
R2250 gnd.n5873 gnd.n5872 585
R2251 gnd.n5297 gnd.n5295 585
R2252 gnd.n5304 gnd.n5295 585
R2253 gnd.n5865 gnd.n5864 585
R2254 gnd.n5864 gnd.n5863 585
R2255 gnd.n5300 gnd.n5299 585
R2256 gnd.n5844 gnd.n5300 585
R2257 gnd.n5830 gnd.n5323 585
R2258 gnd.n5323 gnd.n5313 585
R2259 gnd.n5832 gnd.n5831 585
R2260 gnd.n5833 gnd.n5832 585
R2261 gnd.n5324 gnd.n5322 585
R2262 gnd.n5821 gnd.n5322 585
R2263 gnd.n5825 gnd.n5824 585
R2264 gnd.n5824 gnd.n5823 585
R2265 gnd.n5327 gnd.n5326 585
R2266 gnd.n5787 gnd.n5327 585
R2267 gnd.n5771 gnd.n5770 585
R2268 gnd.n5770 gnd.n5337 585
R2269 gnd.n5772 gnd.n5356 585
R2270 gnd.n5356 gnd.n5336 585
R2271 gnd.n5774 gnd.n5773 585
R2272 gnd.n5775 gnd.n5774 585
R2273 gnd.n5357 gnd.n5355 585
R2274 gnd.n5355 gnd.n5352 585
R2275 gnd.n5764 gnd.n5763 585
R2276 gnd.n5763 gnd.n5762 585
R2277 gnd.n5360 gnd.n5359 585
R2278 gnd.n5369 gnd.n5360 585
R2279 gnd.n5735 gnd.n5382 585
R2280 gnd.n5382 gnd.n5368 585
R2281 gnd.n5737 gnd.n5736 585
R2282 gnd.n5738 gnd.n5737 585
R2283 gnd.n5383 gnd.n5381 585
R2284 gnd.n5390 gnd.n5381 585
R2285 gnd.n5730 gnd.n5729 585
R2286 gnd.n5729 gnd.n5728 585
R2287 gnd.n5386 gnd.n5385 585
R2288 gnd.n5709 gnd.n5386 585
R2289 gnd.n5705 gnd.n5704 585
R2290 gnd.n5706 gnd.n5705 585
R2291 gnd.n5404 gnd.n5403 585
R2292 gnd.n5411 gnd.n5403 585
R2293 gnd.n5700 gnd.n5699 585
R2294 gnd.n5699 gnd.n5698 585
R2295 gnd.n5407 gnd.n5406 585
R2296 gnd.n5688 gnd.n5407 585
R2297 gnd.n5675 gnd.n5674 585
R2298 gnd.n5673 gnd.n5626 585
R2299 gnd.n5672 gnd.n5625 585
R2300 gnd.n5677 gnd.n5625 585
R2301 gnd.n5671 gnd.n5670 585
R2302 gnd.n5669 gnd.n5668 585
R2303 gnd.n5667 gnd.n5666 585
R2304 gnd.n5665 gnd.n5664 585
R2305 gnd.n5663 gnd.n5662 585
R2306 gnd.n5661 gnd.n5660 585
R2307 gnd.n5659 gnd.n5658 585
R2308 gnd.n5657 gnd.n5656 585
R2309 gnd.n5655 gnd.n5654 585
R2310 gnd.n5653 gnd.n5652 585
R2311 gnd.n5651 gnd.n5650 585
R2312 gnd.n5649 gnd.n5648 585
R2313 gnd.n5647 gnd.n5646 585
R2314 gnd.n5642 gnd.n5418 585
R2315 gnd.n6395 gnd.n6394 585
R2316 gnd.n6397 gnd.n5079 585
R2317 gnd.n6399 gnd.n6398 585
R2318 gnd.n6400 gnd.n5072 585
R2319 gnd.n6402 gnd.n6401 585
R2320 gnd.n6404 gnd.n5070 585
R2321 gnd.n6406 gnd.n6405 585
R2322 gnd.n6407 gnd.n5065 585
R2323 gnd.n6409 gnd.n6408 585
R2324 gnd.n6411 gnd.n5063 585
R2325 gnd.n6413 gnd.n6412 585
R2326 gnd.n6414 gnd.n5058 585
R2327 gnd.n6416 gnd.n6415 585
R2328 gnd.n6418 gnd.n5056 585
R2329 gnd.n6420 gnd.n6419 585
R2330 gnd.n6421 gnd.n5054 585
R2331 gnd.n6422 gnd.n5049 585
R2332 gnd.n5049 gnd.n5047 585
R2333 gnd.n6302 gnd.n1029 585
R2334 gnd.n6427 gnd.n1029 585
R2335 gnd.n6304 gnd.n6303 585
R2336 gnd.n6304 gnd.n1027 585
R2337 gnd.n6306 gnd.n6305 585
R2338 gnd.n6305 gnd.n1019 585
R2339 gnd.n6307 gnd.n1017 585
R2340 gnd.n6435 gnd.n1017 585
R2341 gnd.n6310 gnd.n6309 585
R2342 gnd.n6309 gnd.n6308 585
R2343 gnd.n6311 gnd.n1004 585
R2344 gnd.n6441 gnd.n1004 585
R2345 gnd.n6313 gnd.n6312 585
R2346 gnd.n6313 gnd.n1002 585
R2347 gnd.n6315 gnd.n6314 585
R2348 gnd.n6314 gnd.n993 585
R2349 gnd.n6316 gnd.n991 585
R2350 gnd.n6449 gnd.n991 585
R2351 gnd.n6318 gnd.n6317 585
R2352 gnd.n6319 gnd.n6318 585
R2353 gnd.n6031 gnd.n981 585
R2354 gnd.n6455 gnd.n981 585
R2355 gnd.n6030 gnd.n6029 585
R2356 gnd.n6029 gnd.n979 585
R2357 gnd.n6028 gnd.n5137 585
R2358 gnd.n6028 gnd.n970 585
R2359 gnd.n6027 gnd.n6026 585
R2360 gnd.n6027 gnd.n968 585
R2361 gnd.n5140 gnd.n5139 585
R2362 gnd.n6018 gnd.n5139 585
R2363 gnd.n6001 gnd.n6000 585
R2364 gnd.n6002 gnd.n6001 585
R2365 gnd.n5999 gnd.n5152 585
R2366 gnd.n6004 gnd.n5152 585
R2367 gnd.n5963 gnd.n5154 585
R2368 gnd.n5963 gnd.n5158 585
R2369 gnd.n5965 gnd.n5964 585
R2370 gnd.n5964 gnd.n5166 585
R2371 gnd.n5962 gnd.n5171 585
R2372 gnd.n5962 gnd.n5164 585
R2373 gnd.n5961 gnd.n5173 585
R2374 gnd.n5961 gnd.n5960 585
R2375 gnd.n5938 gnd.n5172 585
R2376 gnd.n5185 gnd.n5172 585
R2377 gnd.n5937 gnd.n5183 585
R2378 gnd.n5947 gnd.n5183 585
R2379 gnd.n5928 gnd.n5190 585
R2380 gnd.n5929 gnd.n5928 585
R2381 gnd.n5927 gnd.n5926 585
R2382 gnd.n5927 gnd.n5194 585
R2383 gnd.n5925 gnd.n5196 585
R2384 gnd.n5918 gnd.n5196 585
R2385 gnd.n5211 gnd.n5197 585
R2386 gnd.n5211 gnd.n5201 585
R2387 gnd.n5878 gnd.n5212 585
R2388 gnd.n5908 gnd.n5212 585
R2389 gnd.n5877 gnd.n5876 585
R2390 gnd.n5876 gnd.n5283 585
R2391 gnd.n5875 gnd.n5290 585
R2392 gnd.n5875 gnd.n5282 585
R2393 gnd.n5874 gnd.n5292 585
R2394 gnd.n5874 gnd.n5873 585
R2395 gnd.n5853 gnd.n5291 585
R2396 gnd.n5304 gnd.n5291 585
R2397 gnd.n5852 gnd.n5302 585
R2398 gnd.n5863 gnd.n5302 585
R2399 gnd.n5843 gnd.n5309 585
R2400 gnd.n5844 gnd.n5843 585
R2401 gnd.n5842 gnd.n5841 585
R2402 gnd.n5842 gnd.n5313 585
R2403 gnd.n5840 gnd.n5315 585
R2404 gnd.n5833 gnd.n5315 585
R2405 gnd.n5820 gnd.n5316 585
R2406 gnd.n5821 gnd.n5820 585
R2407 gnd.n5790 gnd.n5329 585
R2408 gnd.n5823 gnd.n5329 585
R2409 gnd.n5789 gnd.n5788 585
R2410 gnd.n5788 gnd.n5787 585
R2411 gnd.n5785 gnd.n5346 585
R2412 gnd.n5785 gnd.n5337 585
R2413 gnd.n5784 gnd.n5783 585
R2414 gnd.n5784 gnd.n5336 585
R2415 gnd.n5348 gnd.n5347 585
R2416 gnd.n5775 gnd.n5347 585
R2417 gnd.n5744 gnd.n5743 585
R2418 gnd.n5743 gnd.n5352 585
R2419 gnd.n5745 gnd.n5362 585
R2420 gnd.n5762 gnd.n5362 585
R2421 gnd.n5742 gnd.n5741 585
R2422 gnd.n5741 gnd.n5369 585
R2423 gnd.n5740 gnd.n5376 585
R2424 gnd.n5740 gnd.n5368 585
R2425 gnd.n5739 gnd.n5378 585
R2426 gnd.n5739 gnd.n5738 585
R2427 gnd.n5718 gnd.n5377 585
R2428 gnd.n5390 gnd.n5377 585
R2429 gnd.n5717 gnd.n5388 585
R2430 gnd.n5728 gnd.n5388 585
R2431 gnd.n5708 gnd.n5395 585
R2432 gnd.n5709 gnd.n5708 585
R2433 gnd.n5707 gnd.n5401 585
R2434 gnd.n5707 gnd.n5706 585
R2435 gnd.n5692 gnd.n5400 585
R2436 gnd.n5411 gnd.n5400 585
R2437 gnd.n5691 gnd.n5409 585
R2438 gnd.n5698 gnd.n5409 585
R2439 gnd.n5690 gnd.n5689 585
R2440 gnd.n5689 gnd.n5688 585
R2441 gnd.n4077 gnd.n4076 585
R2442 gnd.n4078 gnd.n4077 585
R2443 gnd.n3991 gnd.n1885 585
R2444 gnd.n3986 gnd.n1885 585
R2445 gnd.n3990 gnd.n3989 585
R2446 gnd.n3989 gnd.n3988 585
R2447 gnd.n1888 gnd.n1887 585
R2448 gnd.n3714 gnd.n1888 585
R2449 gnd.n3703 gnd.n1959 585
R2450 gnd.n1959 gnd.n1958 585
R2451 gnd.n3705 gnd.n3704 585
R2452 gnd.n3706 gnd.n3705 585
R2453 gnd.n3702 gnd.n1956 585
R2454 gnd.n1964 gnd.n1956 585
R2455 gnd.n3701 gnd.n3700 585
R2456 gnd.n3700 gnd.n3699 585
R2457 gnd.n1961 gnd.n1960 585
R2458 gnd.n3581 gnd.n1961 585
R2459 gnd.n3680 gnd.n3679 585
R2460 gnd.n3681 gnd.n3680 585
R2461 gnd.n3678 gnd.n1976 585
R2462 gnd.n1976 gnd.n1972 585
R2463 gnd.n3677 gnd.n3676 585
R2464 gnd.n3676 gnd.n3675 585
R2465 gnd.n1978 gnd.n1977 585
R2466 gnd.n3590 gnd.n1978 585
R2467 gnd.n3657 gnd.n3656 585
R2468 gnd.n3658 gnd.n3657 585
R2469 gnd.n3655 gnd.n1989 585
R2470 gnd.n1989 gnd.n1986 585
R2471 gnd.n3654 gnd.n3653 585
R2472 gnd.n3653 gnd.n3652 585
R2473 gnd.n1991 gnd.n1990 585
R2474 gnd.n3597 gnd.n1991 585
R2475 gnd.n3637 gnd.n3636 585
R2476 gnd.n3638 gnd.n3637 585
R2477 gnd.n3635 gnd.n2002 585
R2478 gnd.n3630 gnd.n2002 585
R2479 gnd.n3634 gnd.n3633 585
R2480 gnd.n3633 gnd.n3632 585
R2481 gnd.n2004 gnd.n2003 585
R2482 gnd.n2016 gnd.n2004 585
R2483 gnd.n3567 gnd.n3566 585
R2484 gnd.n3567 gnd.n2015 585
R2485 gnd.n3571 gnd.n3570 585
R2486 gnd.n3570 gnd.n3569 585
R2487 gnd.n3572 gnd.n2022 585
R2488 gnd.n3610 gnd.n2022 585
R2489 gnd.n3573 gnd.n2031 585
R2490 gnd.n3498 gnd.n2031 585
R2491 gnd.n3575 gnd.n3574 585
R2492 gnd.n3576 gnd.n3575 585
R2493 gnd.n3565 gnd.n2030 585
R2494 gnd.n3559 gnd.n2030 585
R2495 gnd.n3564 gnd.n3563 585
R2496 gnd.n3563 gnd.n3562 585
R2497 gnd.n2033 gnd.n2032 585
R2498 gnd.n3548 gnd.n2033 585
R2499 gnd.n3538 gnd.n2050 585
R2500 gnd.n2050 gnd.n2042 585
R2501 gnd.n3540 gnd.n3539 585
R2502 gnd.n3541 gnd.n3540 585
R2503 gnd.n3537 gnd.n2049 585
R2504 gnd.n2054 gnd.n2049 585
R2505 gnd.n3536 gnd.n3535 585
R2506 gnd.n3535 gnd.n3534 585
R2507 gnd.n2052 gnd.n2051 585
R2508 gnd.n3489 gnd.n2052 585
R2509 gnd.n3522 gnd.n3521 585
R2510 gnd.n3523 gnd.n3522 585
R2511 gnd.n3520 gnd.n2065 585
R2512 gnd.n2065 gnd.n2061 585
R2513 gnd.n3519 gnd.n3518 585
R2514 gnd.n3518 gnd.n3517 585
R2515 gnd.n2067 gnd.n2066 585
R2516 gnd.n3479 gnd.n2067 585
R2517 gnd.n3464 gnd.n3463 585
R2518 gnd.n3463 gnd.n2077 585
R2519 gnd.n3465 gnd.n2087 585
R2520 gnd.n3448 gnd.n2087 585
R2521 gnd.n3467 gnd.n3466 585
R2522 gnd.n3468 gnd.n3467 585
R2523 gnd.n3462 gnd.n2086 585
R2524 gnd.n2086 gnd.n2083 585
R2525 gnd.n3461 gnd.n3460 585
R2526 gnd.n3460 gnd.n3459 585
R2527 gnd.n2089 gnd.n2088 585
R2528 gnd.n3439 gnd.n2089 585
R2529 gnd.n3424 gnd.n3423 585
R2530 gnd.n3423 gnd.n2100 585
R2531 gnd.n3425 gnd.n2110 585
R2532 gnd.n3412 gnd.n2110 585
R2533 gnd.n3427 gnd.n3426 585
R2534 gnd.n3428 gnd.n3427 585
R2535 gnd.n3422 gnd.n2109 585
R2536 gnd.n2109 gnd.n2106 585
R2537 gnd.n3421 gnd.n3420 585
R2538 gnd.n3420 gnd.n3419 585
R2539 gnd.n2112 gnd.n2111 585
R2540 gnd.n2125 gnd.n2112 585
R2541 gnd.n3396 gnd.n3395 585
R2542 gnd.n3397 gnd.n3396 585
R2543 gnd.n3394 gnd.n2127 585
R2544 gnd.n3389 gnd.n2127 585
R2545 gnd.n3393 gnd.n3392 585
R2546 gnd.n3392 gnd.n3391 585
R2547 gnd.n2129 gnd.n2128 585
R2548 gnd.n3376 gnd.n2129 585
R2549 gnd.n3364 gnd.n2147 585
R2550 gnd.n2147 gnd.n2139 585
R2551 gnd.n3366 gnd.n3365 585
R2552 gnd.n3367 gnd.n3366 585
R2553 gnd.n3363 gnd.n2146 585
R2554 gnd.n3307 gnd.n2146 585
R2555 gnd.n3362 gnd.n3361 585
R2556 gnd.n3361 gnd.n3360 585
R2557 gnd.n2149 gnd.n2148 585
R2558 gnd.n3335 gnd.n2149 585
R2559 gnd.n3348 gnd.n3347 585
R2560 gnd.n3349 gnd.n3348 585
R2561 gnd.n3346 gnd.n2160 585
R2562 gnd.n3341 gnd.n2160 585
R2563 gnd.n3345 gnd.n3344 585
R2564 gnd.n3344 gnd.n3343 585
R2565 gnd.n2162 gnd.n2161 585
R2566 gnd.n3330 gnd.n2162 585
R2567 gnd.n3281 gnd.n3278 585
R2568 gnd.n3281 gnd.n3280 585
R2569 gnd.n3282 gnd.n3277 585
R2570 gnd.n3282 gnd.n2176 585
R2571 gnd.n3284 gnd.n3283 585
R2572 gnd.n3283 gnd.n2175 585
R2573 gnd.n3285 gnd.n3275 585
R2574 gnd.n3275 gnd.n3274 585
R2575 gnd.n3287 gnd.n3286 585
R2576 gnd.n3288 gnd.n3287 585
R2577 gnd.n3276 gnd.n2186 585
R2578 gnd.n3264 gnd.n2186 585
R2579 gnd.n1489 gnd.n1488 585
R2580 gnd.n1493 gnd.n1489 585
R2581 gnd.n4665 gnd.n4664 585
R2582 gnd.n4664 gnd.n4663 585
R2583 gnd.n4666 gnd.n1467 585
R2584 gnd.n3257 gnd.n1467 585
R2585 gnd.n4731 gnd.n4730 585
R2586 gnd.n4729 gnd.n1466 585
R2587 gnd.n4728 gnd.n1465 585
R2588 gnd.n4733 gnd.n1465 585
R2589 gnd.n4727 gnd.n4726 585
R2590 gnd.n4725 gnd.n4724 585
R2591 gnd.n4723 gnd.n4722 585
R2592 gnd.n4721 gnd.n4720 585
R2593 gnd.n4719 gnd.n4718 585
R2594 gnd.n4717 gnd.n4716 585
R2595 gnd.n4715 gnd.n4714 585
R2596 gnd.n4713 gnd.n4712 585
R2597 gnd.n4711 gnd.n4710 585
R2598 gnd.n4709 gnd.n4708 585
R2599 gnd.n4707 gnd.n4706 585
R2600 gnd.n4705 gnd.n4704 585
R2601 gnd.n4703 gnd.n4702 585
R2602 gnd.n4701 gnd.n4700 585
R2603 gnd.n4699 gnd.n4698 585
R2604 gnd.n4697 gnd.n4696 585
R2605 gnd.n4695 gnd.n4694 585
R2606 gnd.n4693 gnd.n4692 585
R2607 gnd.n4691 gnd.n4690 585
R2608 gnd.n4689 gnd.n4688 585
R2609 gnd.n4687 gnd.n4686 585
R2610 gnd.n4685 gnd.n4684 585
R2611 gnd.n4683 gnd.n4682 585
R2612 gnd.n4681 gnd.n4680 585
R2613 gnd.n4679 gnd.n4678 585
R2614 gnd.n4677 gnd.n4676 585
R2615 gnd.n4675 gnd.n4674 585
R2616 gnd.n4673 gnd.n4672 585
R2617 gnd.n4671 gnd.n1430 585
R2618 gnd.n4736 gnd.n4735 585
R2619 gnd.n1432 gnd.n1429 585
R2620 gnd.n2191 gnd.n2190 585
R2621 gnd.n2193 gnd.n2192 585
R2622 gnd.n2196 gnd.n2195 585
R2623 gnd.n2198 gnd.n2197 585
R2624 gnd.n2200 gnd.n2199 585
R2625 gnd.n2202 gnd.n2201 585
R2626 gnd.n2204 gnd.n2203 585
R2627 gnd.n2206 gnd.n2205 585
R2628 gnd.n2208 gnd.n2207 585
R2629 gnd.n2210 gnd.n2209 585
R2630 gnd.n2212 gnd.n2211 585
R2631 gnd.n2214 gnd.n2213 585
R2632 gnd.n2216 gnd.n2215 585
R2633 gnd.n2218 gnd.n2217 585
R2634 gnd.n2220 gnd.n2219 585
R2635 gnd.n2222 gnd.n2221 585
R2636 gnd.n2224 gnd.n2223 585
R2637 gnd.n2226 gnd.n2225 585
R2638 gnd.n2228 gnd.n2227 585
R2639 gnd.n2230 gnd.n2229 585
R2640 gnd.n2232 gnd.n2231 585
R2641 gnd.n2234 gnd.n2233 585
R2642 gnd.n2236 gnd.n2235 585
R2643 gnd.n2238 gnd.n2237 585
R2644 gnd.n2240 gnd.n2239 585
R2645 gnd.n2242 gnd.n2241 585
R2646 gnd.n2244 gnd.n2243 585
R2647 gnd.n2246 gnd.n2245 585
R2648 gnd.n2248 gnd.n2247 585
R2649 gnd.n2250 gnd.n2249 585
R2650 gnd.n2252 gnd.n2251 585
R2651 gnd.n4081 gnd.n4080 585
R2652 gnd.n4083 gnd.n4082 585
R2653 gnd.n4085 gnd.n4084 585
R2654 gnd.n4087 gnd.n4086 585
R2655 gnd.n4089 gnd.n4088 585
R2656 gnd.n4091 gnd.n4090 585
R2657 gnd.n4093 gnd.n4092 585
R2658 gnd.n4095 gnd.n4094 585
R2659 gnd.n4097 gnd.n4096 585
R2660 gnd.n4099 gnd.n4098 585
R2661 gnd.n4101 gnd.n4100 585
R2662 gnd.n4103 gnd.n4102 585
R2663 gnd.n4105 gnd.n4104 585
R2664 gnd.n4107 gnd.n4106 585
R2665 gnd.n4109 gnd.n4108 585
R2666 gnd.n4111 gnd.n4110 585
R2667 gnd.n4113 gnd.n4112 585
R2668 gnd.n4115 gnd.n4114 585
R2669 gnd.n4117 gnd.n4116 585
R2670 gnd.n4119 gnd.n4118 585
R2671 gnd.n4121 gnd.n4120 585
R2672 gnd.n4123 gnd.n4122 585
R2673 gnd.n4125 gnd.n4124 585
R2674 gnd.n4127 gnd.n4126 585
R2675 gnd.n4129 gnd.n4128 585
R2676 gnd.n4131 gnd.n4130 585
R2677 gnd.n4133 gnd.n4132 585
R2678 gnd.n4135 gnd.n4134 585
R2679 gnd.n4137 gnd.n4136 585
R2680 gnd.n4139 gnd.n1878 585
R2681 gnd.n4141 gnd.n4140 585
R2682 gnd.n4143 gnd.n1842 585
R2683 gnd.n4145 gnd.n4144 585
R2684 gnd.n4148 gnd.n4147 585
R2685 gnd.n1845 gnd.n1843 585
R2686 gnd.n4014 gnd.n4013 585
R2687 gnd.n4016 gnd.n4015 585
R2688 gnd.n4019 gnd.n4018 585
R2689 gnd.n4021 gnd.n4020 585
R2690 gnd.n4023 gnd.n4022 585
R2691 gnd.n4025 gnd.n4024 585
R2692 gnd.n4027 gnd.n4026 585
R2693 gnd.n4029 gnd.n4028 585
R2694 gnd.n4031 gnd.n4030 585
R2695 gnd.n4033 gnd.n4032 585
R2696 gnd.n4035 gnd.n4034 585
R2697 gnd.n4037 gnd.n4036 585
R2698 gnd.n4039 gnd.n4038 585
R2699 gnd.n4041 gnd.n4040 585
R2700 gnd.n4043 gnd.n4042 585
R2701 gnd.n4045 gnd.n4044 585
R2702 gnd.n4047 gnd.n4046 585
R2703 gnd.n4049 gnd.n4048 585
R2704 gnd.n4051 gnd.n4050 585
R2705 gnd.n4053 gnd.n4052 585
R2706 gnd.n4055 gnd.n4054 585
R2707 gnd.n4057 gnd.n4056 585
R2708 gnd.n4059 gnd.n4058 585
R2709 gnd.n4061 gnd.n4060 585
R2710 gnd.n4063 gnd.n4062 585
R2711 gnd.n4065 gnd.n4064 585
R2712 gnd.n4067 gnd.n4066 585
R2713 gnd.n4069 gnd.n4068 585
R2714 gnd.n4071 gnd.n4070 585
R2715 gnd.n4073 gnd.n4072 585
R2716 gnd.n4074 gnd.n1886 585
R2717 gnd.n4079 gnd.n1881 585
R2718 gnd.n4079 gnd.n4078 585
R2719 gnd.n3710 gnd.n1882 585
R2720 gnd.n3986 gnd.n1882 585
R2721 gnd.n3711 gnd.n1890 585
R2722 gnd.n3988 gnd.n1890 585
R2723 gnd.n3713 gnd.n3712 585
R2724 gnd.n3714 gnd.n3713 585
R2725 gnd.n3709 gnd.n1952 585
R2726 gnd.n1958 gnd.n1952 585
R2727 gnd.n3708 gnd.n3707 585
R2728 gnd.n3707 gnd.n3706 585
R2729 gnd.n1954 gnd.n1953 585
R2730 gnd.n1964 gnd.n1954 585
R2731 gnd.n3580 gnd.n1963 585
R2732 gnd.n3699 gnd.n1963 585
R2733 gnd.n3583 gnd.n3582 585
R2734 gnd.n3582 gnd.n3581 585
R2735 gnd.n3584 gnd.n1974 585
R2736 gnd.n3681 gnd.n1974 585
R2737 gnd.n3586 gnd.n3585 585
R2738 gnd.n3585 gnd.n1972 585
R2739 gnd.n3587 gnd.n1979 585
R2740 gnd.n3675 gnd.n1979 585
R2741 gnd.n3592 gnd.n3591 585
R2742 gnd.n3591 gnd.n3590 585
R2743 gnd.n3593 gnd.n1987 585
R2744 gnd.n3658 gnd.n1987 585
R2745 gnd.n3595 gnd.n3594 585
R2746 gnd.n3594 gnd.n1986 585
R2747 gnd.n3596 gnd.n1993 585
R2748 gnd.n3652 gnd.n1993 585
R2749 gnd.n3599 gnd.n3598 585
R2750 gnd.n3598 gnd.n3597 585
R2751 gnd.n3600 gnd.n2000 585
R2752 gnd.n3638 gnd.n2000 585
R2753 gnd.n3601 gnd.n2007 585
R2754 gnd.n3630 gnd.n2007 585
R2755 gnd.n3602 gnd.n2006 585
R2756 gnd.n3632 gnd.n2006 585
R2757 gnd.n3604 gnd.n3603 585
R2758 gnd.n3604 gnd.n2016 585
R2759 gnd.n3606 gnd.n3605 585
R2760 gnd.n3605 gnd.n2015 585
R2761 gnd.n3607 gnd.n2025 585
R2762 gnd.n3569 gnd.n2025 585
R2763 gnd.n3609 gnd.n3608 585
R2764 gnd.n3610 gnd.n3609 585
R2765 gnd.n3579 gnd.n2024 585
R2766 gnd.n3498 gnd.n2024 585
R2767 gnd.n3578 gnd.n3577 585
R2768 gnd.n3577 gnd.n3576 585
R2769 gnd.n2027 gnd.n2026 585
R2770 gnd.n3559 gnd.n2027 585
R2771 gnd.n3545 gnd.n2035 585
R2772 gnd.n3562 gnd.n2035 585
R2773 gnd.n3547 gnd.n3546 585
R2774 gnd.n3548 gnd.n3547 585
R2775 gnd.n3544 gnd.n2044 585
R2776 gnd.n2044 gnd.n2042 585
R2777 gnd.n3543 gnd.n3542 585
R2778 gnd.n3542 gnd.n3541 585
R2779 gnd.n2046 gnd.n2045 585
R2780 gnd.n2054 gnd.n2046 585
R2781 gnd.n3486 gnd.n2053 585
R2782 gnd.n3534 gnd.n2053 585
R2783 gnd.n3488 gnd.n3487 585
R2784 gnd.n3489 gnd.n3488 585
R2785 gnd.n3485 gnd.n2063 585
R2786 gnd.n3523 gnd.n2063 585
R2787 gnd.n3484 gnd.n3483 585
R2788 gnd.n3483 gnd.n2061 585
R2789 gnd.n3482 gnd.n2069 585
R2790 gnd.n3517 gnd.n2069 585
R2791 gnd.n3481 gnd.n3480 585
R2792 gnd.n3480 gnd.n3479 585
R2793 gnd.n2076 gnd.n2075 585
R2794 gnd.n2077 gnd.n2076 585
R2795 gnd.n3447 gnd.n3446 585
R2796 gnd.n3448 gnd.n3447 585
R2797 gnd.n3445 gnd.n2084 585
R2798 gnd.n3468 gnd.n2084 585
R2799 gnd.n3444 gnd.n3443 585
R2800 gnd.n3443 gnd.n2083 585
R2801 gnd.n3442 gnd.n2091 585
R2802 gnd.n3459 gnd.n2091 585
R2803 gnd.n3441 gnd.n3440 585
R2804 gnd.n3440 gnd.n3439 585
R2805 gnd.n2099 gnd.n2098 585
R2806 gnd.n2100 gnd.n2099 585
R2807 gnd.n3414 gnd.n3413 585
R2808 gnd.n3413 gnd.n3412 585
R2809 gnd.n3415 gnd.n2107 585
R2810 gnd.n3428 gnd.n2107 585
R2811 gnd.n3416 gnd.n2115 585
R2812 gnd.n2115 gnd.n2106 585
R2813 gnd.n3418 gnd.n3417 585
R2814 gnd.n3419 gnd.n3418 585
R2815 gnd.n2116 gnd.n2114 585
R2816 gnd.n2125 gnd.n2114 585
R2817 gnd.n3371 gnd.n2124 585
R2818 gnd.n3397 gnd.n2124 585
R2819 gnd.n3372 gnd.n2132 585
R2820 gnd.n3389 gnd.n2132 585
R2821 gnd.n3373 gnd.n2131 585
R2822 gnd.n3391 gnd.n2131 585
R2823 gnd.n3375 gnd.n3374 585
R2824 gnd.n3376 gnd.n3375 585
R2825 gnd.n3370 gnd.n2141 585
R2826 gnd.n2141 gnd.n2139 585
R2827 gnd.n3369 gnd.n3368 585
R2828 gnd.n3368 gnd.n3367 585
R2829 gnd.n2143 gnd.n2142 585
R2830 gnd.n3307 gnd.n2143 585
R2831 gnd.n3334 gnd.n2151 585
R2832 gnd.n3360 gnd.n2151 585
R2833 gnd.n3337 gnd.n3336 585
R2834 gnd.n3336 gnd.n3335 585
R2835 gnd.n3338 gnd.n2158 585
R2836 gnd.n3349 gnd.n2158 585
R2837 gnd.n3340 gnd.n3339 585
R2838 gnd.n3341 gnd.n3340 585
R2839 gnd.n3333 gnd.n2164 585
R2840 gnd.n3343 gnd.n2164 585
R2841 gnd.n3332 gnd.n3331 585
R2842 gnd.n3331 gnd.n3330 585
R2843 gnd.n2167 gnd.n2166 585
R2844 gnd.n3280 gnd.n2167 585
R2845 gnd.n3269 gnd.n3268 585
R2846 gnd.n3268 gnd.n2176 585
R2847 gnd.n3270 gnd.n2187 585
R2848 gnd.n2187 gnd.n2175 585
R2849 gnd.n3272 gnd.n3271 585
R2850 gnd.n3274 gnd.n3272 585
R2851 gnd.n3267 gnd.n2184 585
R2852 gnd.n3288 gnd.n2184 585
R2853 gnd.n3266 gnd.n3265 585
R2854 gnd.n3265 gnd.n3264 585
R2855 gnd.n3262 gnd.n3261 585
R2856 gnd.n3262 gnd.n1493 585
R2857 gnd.n3260 gnd.n1491 585
R2858 gnd.n4663 gnd.n1491 585
R2859 gnd.n3259 gnd.n3258 585
R2860 gnd.n3258 gnd.n3257 585
R2861 gnd.n4787 gnd.n4786 585
R2862 gnd.n4788 gnd.n4787 585
R2863 gnd.n1363 gnd.n1362 585
R2864 gnd.n3021 gnd.n1363 585
R2865 gnd.n4796 gnd.n4795 585
R2866 gnd.n4795 gnd.n4794 585
R2867 gnd.n4797 gnd.n1357 585
R2868 gnd.n3014 gnd.n1357 585
R2869 gnd.n4799 gnd.n4798 585
R2870 gnd.n4800 gnd.n4799 585
R2871 gnd.n1343 gnd.n1342 585
R2872 gnd.n3009 gnd.n1343 585
R2873 gnd.n4808 gnd.n4807 585
R2874 gnd.n4807 gnd.n4806 585
R2875 gnd.n4809 gnd.n1337 585
R2876 gnd.n3036 gnd.n1337 585
R2877 gnd.n4811 gnd.n4810 585
R2878 gnd.n4812 gnd.n4811 585
R2879 gnd.n1322 gnd.n1321 585
R2880 gnd.n3002 gnd.n1322 585
R2881 gnd.n4820 gnd.n4819 585
R2882 gnd.n4819 gnd.n4818 585
R2883 gnd.n4821 gnd.n1316 585
R2884 gnd.n2994 gnd.n1316 585
R2885 gnd.n4823 gnd.n4822 585
R2886 gnd.n4824 gnd.n4823 585
R2887 gnd.n1303 gnd.n1302 585
R2888 gnd.n2987 gnd.n1303 585
R2889 gnd.n4832 gnd.n4831 585
R2890 gnd.n4831 gnd.n4830 585
R2891 gnd.n4833 gnd.n1297 585
R2892 gnd.n2979 gnd.n1297 585
R2893 gnd.n4835 gnd.n4834 585
R2894 gnd.n4836 gnd.n4835 585
R2895 gnd.n1282 gnd.n1281 585
R2896 gnd.n2925 gnd.n1282 585
R2897 gnd.n4844 gnd.n4843 585
R2898 gnd.n4843 gnd.n4842 585
R2899 gnd.n4845 gnd.n1277 585
R2900 gnd.n2916 gnd.n1277 585
R2901 gnd.n4847 gnd.n4846 585
R2902 gnd.n4848 gnd.n4847 585
R2903 gnd.n1262 gnd.n1260 585
R2904 gnd.n2910 gnd.n1262 585
R2905 gnd.n4856 gnd.n4855 585
R2906 gnd.n4855 gnd.n4854 585
R2907 gnd.n1261 gnd.n1259 585
R2908 gnd.n2939 gnd.n1261 585
R2909 gnd.n2902 gnd.n2901 585
R2910 gnd.n2903 gnd.n2902 585
R2911 gnd.n2900 gnd.n2899 585
R2912 gnd.n2899 gnd.n2898 585
R2913 gnd.n2886 gnd.n2613 585
R2914 gnd.n2878 gnd.n2613 585
R2915 gnd.n2888 gnd.n2887 585
R2916 gnd.n2889 gnd.n2888 585
R2917 gnd.n2885 gnd.n2624 585
R2918 gnd.n2885 gnd.n2884 585
R2919 gnd.n2623 gnd.n1258 585
R2920 gnd.n2852 gnd.n2623 585
R2921 gnd.n2859 gnd.n1252 585
R2922 gnd.n2860 gnd.n2859 585
R2923 gnd.n4859 gnd.n1249 585
R2924 gnd.n2640 gnd.n1249 585
R2925 gnd.n4861 gnd.n4860 585
R2926 gnd.n4862 gnd.n4861 585
R2927 gnd.n1234 gnd.n1233 585
R2928 gnd.n2841 gnd.n1234 585
R2929 gnd.n4870 gnd.n4869 585
R2930 gnd.n4869 gnd.n4868 585
R2931 gnd.n4871 gnd.n1228 585
R2932 gnd.n2834 gnd.n1228 585
R2933 gnd.n4873 gnd.n4872 585
R2934 gnd.n4874 gnd.n4873 585
R2935 gnd.n1214 gnd.n1213 585
R2936 gnd.n2825 gnd.n1214 585
R2937 gnd.n4882 gnd.n4881 585
R2938 gnd.n4881 gnd.n4880 585
R2939 gnd.n4883 gnd.n1208 585
R2940 gnd.n2819 gnd.n1208 585
R2941 gnd.n4885 gnd.n4884 585
R2942 gnd.n4886 gnd.n4885 585
R2943 gnd.n1193 gnd.n1192 585
R2944 gnd.n2772 gnd.n1193 585
R2945 gnd.n4894 gnd.n4893 585
R2946 gnd.n4893 gnd.n4892 585
R2947 gnd.n4895 gnd.n1187 585
R2948 gnd.n2766 gnd.n1187 585
R2949 gnd.n4897 gnd.n4896 585
R2950 gnd.n4898 gnd.n4897 585
R2951 gnd.n1174 gnd.n1173 585
R2952 gnd.n1177 gnd.n1174 585
R2953 gnd.n4906 gnd.n4905 585
R2954 gnd.n4905 gnd.n4904 585
R2955 gnd.n4907 gnd.n1168 585
R2956 gnd.n1168 gnd.n1167 585
R2957 gnd.n4909 gnd.n4908 585
R2958 gnd.n4910 gnd.n4909 585
R2959 gnd.n1151 gnd.n1150 585
R2960 gnd.n1155 gnd.n1151 585
R2961 gnd.n4918 gnd.n4917 585
R2962 gnd.n4917 gnd.n4916 585
R2963 gnd.n4919 gnd.n1144 585
R2964 gnd.n1152 gnd.n1144 585
R2965 gnd.n4921 gnd.n4920 585
R2966 gnd.n4922 gnd.n4921 585
R2967 gnd.n1145 gnd.n1071 585
R2968 gnd.n1071 gnd.n1068 585
R2969 gnd.n5044 gnd.n5043 585
R2970 gnd.n5042 gnd.n1070 585
R2971 gnd.n5041 gnd.n1069 585
R2972 gnd.n5046 gnd.n1069 585
R2973 gnd.n5040 gnd.n5039 585
R2974 gnd.n5038 gnd.n5037 585
R2975 gnd.n5036 gnd.n5035 585
R2976 gnd.n5034 gnd.n5033 585
R2977 gnd.n5032 gnd.n5031 585
R2978 gnd.n5030 gnd.n5029 585
R2979 gnd.n5028 gnd.n5027 585
R2980 gnd.n5026 gnd.n5025 585
R2981 gnd.n5024 gnd.n5023 585
R2982 gnd.n5022 gnd.n5021 585
R2983 gnd.n5020 gnd.n5019 585
R2984 gnd.n5018 gnd.n5017 585
R2985 gnd.n5016 gnd.n5015 585
R2986 gnd.n5014 gnd.n5013 585
R2987 gnd.n5012 gnd.n5011 585
R2988 gnd.n5009 gnd.n5008 585
R2989 gnd.n5007 gnd.n5006 585
R2990 gnd.n5005 gnd.n5004 585
R2991 gnd.n5003 gnd.n5002 585
R2992 gnd.n5001 gnd.n5000 585
R2993 gnd.n4999 gnd.n4998 585
R2994 gnd.n4997 gnd.n4996 585
R2995 gnd.n4995 gnd.n4994 585
R2996 gnd.n4993 gnd.n4992 585
R2997 gnd.n4991 gnd.n4990 585
R2998 gnd.n4989 gnd.n4988 585
R2999 gnd.n4987 gnd.n4986 585
R3000 gnd.n4985 gnd.n4984 585
R3001 gnd.n4983 gnd.n4982 585
R3002 gnd.n4981 gnd.n4980 585
R3003 gnd.n4979 gnd.n4978 585
R3004 gnd.n4977 gnd.n4976 585
R3005 gnd.n4975 gnd.n4974 585
R3006 gnd.n4973 gnd.n4972 585
R3007 gnd.n4971 gnd.n4970 585
R3008 gnd.n4969 gnd.n4968 585
R3009 gnd.n4967 gnd.n4966 585
R3010 gnd.n4965 gnd.n4964 585
R3011 gnd.n4963 gnd.n4962 585
R3012 gnd.n4961 gnd.n4960 585
R3013 gnd.n4959 gnd.n4958 585
R3014 gnd.n4957 gnd.n4956 585
R3015 gnd.n4955 gnd.n4954 585
R3016 gnd.n4953 gnd.n4952 585
R3017 gnd.n4951 gnd.n4950 585
R3018 gnd.n4949 gnd.n4948 585
R3019 gnd.n4947 gnd.n4946 585
R3020 gnd.n4945 gnd.n4944 585
R3021 gnd.n4943 gnd.n4942 585
R3022 gnd.n4941 gnd.n4940 585
R3023 gnd.n4939 gnd.n4938 585
R3024 gnd.n4937 gnd.n4936 585
R3025 gnd.n4935 gnd.n4934 585
R3026 gnd.n4933 gnd.n4932 585
R3027 gnd.n4931 gnd.n4930 585
R3028 gnd.n1140 gnd.n1133 585
R3029 gnd.n2457 gnd.n2456 585
R3030 gnd.n2454 gnd.n2350 585
R3031 gnd.n2453 gnd.n2452 585
R3032 gnd.n2446 gnd.n2352 585
R3033 gnd.n2448 gnd.n2447 585
R3034 gnd.n2444 gnd.n2354 585
R3035 gnd.n2443 gnd.n2442 585
R3036 gnd.n2436 gnd.n2356 585
R3037 gnd.n2438 gnd.n2437 585
R3038 gnd.n2434 gnd.n2358 585
R3039 gnd.n2433 gnd.n2432 585
R3040 gnd.n2426 gnd.n2360 585
R3041 gnd.n2428 gnd.n2427 585
R3042 gnd.n2424 gnd.n2362 585
R3043 gnd.n2423 gnd.n2422 585
R3044 gnd.n2416 gnd.n2364 585
R3045 gnd.n2418 gnd.n2417 585
R3046 gnd.n2414 gnd.n2366 585
R3047 gnd.n2413 gnd.n2412 585
R3048 gnd.n2406 gnd.n2368 585
R3049 gnd.n2408 gnd.n2407 585
R3050 gnd.n2404 gnd.n2372 585
R3051 gnd.n2403 gnd.n2402 585
R3052 gnd.n2396 gnd.n2374 585
R3053 gnd.n2398 gnd.n2397 585
R3054 gnd.n2394 gnd.n2376 585
R3055 gnd.n2393 gnd.n2392 585
R3056 gnd.n2386 gnd.n2378 585
R3057 gnd.n2388 gnd.n2387 585
R3058 gnd.n2384 gnd.n2381 585
R3059 gnd.n2383 gnd.n1425 585
R3060 gnd.n4738 gnd.n1421 585
R3061 gnd.n4740 gnd.n4739 585
R3062 gnd.n4742 gnd.n1419 585
R3063 gnd.n4744 gnd.n4743 585
R3064 gnd.n4745 gnd.n1414 585
R3065 gnd.n4747 gnd.n4746 585
R3066 gnd.n4749 gnd.n1412 585
R3067 gnd.n4751 gnd.n4750 585
R3068 gnd.n4753 gnd.n1405 585
R3069 gnd.n4755 gnd.n4754 585
R3070 gnd.n4757 gnd.n1403 585
R3071 gnd.n4759 gnd.n4758 585
R3072 gnd.n4760 gnd.n1398 585
R3073 gnd.n4762 gnd.n4761 585
R3074 gnd.n4764 gnd.n1396 585
R3075 gnd.n4766 gnd.n4765 585
R3076 gnd.n4767 gnd.n1391 585
R3077 gnd.n4769 gnd.n4768 585
R3078 gnd.n4771 gnd.n1389 585
R3079 gnd.n4773 gnd.n4772 585
R3080 gnd.n4774 gnd.n1383 585
R3081 gnd.n4776 gnd.n4775 585
R3082 gnd.n4778 gnd.n1382 585
R3083 gnd.n4779 gnd.n1380 585
R3084 gnd.n4782 gnd.n4781 585
R3085 gnd.n4783 gnd.n1377 585
R3086 gnd.n1381 gnd.n1377 585
R3087 gnd.n3018 gnd.n1374 585
R3088 gnd.n4788 gnd.n1374 585
R3089 gnd.n3020 gnd.n3019 585
R3090 gnd.n3021 gnd.n3020 585
R3091 gnd.n3017 gnd.n1365 585
R3092 gnd.n4794 gnd.n1365 585
R3093 gnd.n3016 gnd.n3015 585
R3094 gnd.n3015 gnd.n3014 585
R3095 gnd.n3012 gnd.n1354 585
R3096 gnd.n4800 gnd.n1354 585
R3097 gnd.n3011 gnd.n3010 585
R3098 gnd.n3010 gnd.n3009 585
R3099 gnd.n3008 gnd.n1344 585
R3100 gnd.n4806 gnd.n1344 585
R3101 gnd.n3007 gnd.n2567 585
R3102 gnd.n3036 gnd.n2567 585
R3103 gnd.n3005 gnd.n1334 585
R3104 gnd.n4812 gnd.n1334 585
R3105 gnd.n3004 gnd.n3003 585
R3106 gnd.n3003 gnd.n3002 585
R3107 gnd.n2576 gnd.n1324 585
R3108 gnd.n4818 gnd.n1324 585
R3109 gnd.n2993 gnd.n2992 585
R3110 gnd.n2994 gnd.n2993 585
R3111 gnd.n2990 gnd.n1314 585
R3112 gnd.n4824 gnd.n1314 585
R3113 gnd.n2989 gnd.n2988 585
R3114 gnd.n2988 gnd.n2987 585
R3115 gnd.n2581 gnd.n1304 585
R3116 gnd.n4830 gnd.n1304 585
R3117 gnd.n2921 gnd.n2585 585
R3118 gnd.n2979 gnd.n2585 585
R3119 gnd.n2922 gnd.n1294 585
R3120 gnd.n4836 gnd.n1294 585
R3121 gnd.n2924 gnd.n2923 585
R3122 gnd.n2925 gnd.n2924 585
R3123 gnd.n2919 gnd.n1284 585
R3124 gnd.n4842 gnd.n1284 585
R3125 gnd.n2918 gnd.n2917 585
R3126 gnd.n2917 gnd.n2916 585
R3127 gnd.n2913 gnd.n1275 585
R3128 gnd.n4848 gnd.n1275 585
R3129 gnd.n2912 gnd.n2911 585
R3130 gnd.n2911 gnd.n2910 585
R3131 gnd.n2909 gnd.n1263 585
R3132 gnd.n4854 gnd.n1263 585
R3133 gnd.n2908 gnd.n2598 585
R3134 gnd.n2939 gnd.n2598 585
R3135 gnd.n2612 gnd.n2607 585
R3136 gnd.n2903 gnd.n2612 585
R3137 gnd.n2648 gnd.n2614 585
R3138 gnd.n2898 gnd.n2614 585
R3139 gnd.n2649 gnd.n2633 585
R3140 gnd.n2878 gnd.n2633 585
R3141 gnd.n2650 gnd.n2620 585
R3142 gnd.n2889 gnd.n2620 585
R3143 gnd.n2651 gnd.n2626 585
R3144 gnd.n2884 gnd.n2626 585
R3145 gnd.n2854 gnd.n2853 585
R3146 gnd.n2853 gnd.n2852 585
R3147 gnd.n2855 gnd.n2641 585
R3148 gnd.n2860 gnd.n2641 585
R3149 gnd.n2647 gnd.n2646 585
R3150 gnd.n2646 gnd.n2640 585
R3151 gnd.n2838 gnd.n1246 585
R3152 gnd.n4862 gnd.n1246 585
R3153 gnd.n2840 gnd.n2839 585
R3154 gnd.n2841 gnd.n2840 585
R3155 gnd.n2837 gnd.n1236 585
R3156 gnd.n4868 gnd.n1236 585
R3157 gnd.n2836 gnd.n2835 585
R3158 gnd.n2835 gnd.n2834 585
R3159 gnd.n2656 gnd.n1225 585
R3160 gnd.n4874 gnd.n1225 585
R3161 gnd.n2824 gnd.n2823 585
R3162 gnd.n2825 gnd.n2824 585
R3163 gnd.n2822 gnd.n1215 585
R3164 gnd.n4880 gnd.n1215 585
R3165 gnd.n2821 gnd.n2820 585
R3166 gnd.n2820 gnd.n2819 585
R3167 gnd.n2661 gnd.n1205 585
R3168 gnd.n4886 gnd.n1205 585
R3169 gnd.n2771 gnd.n2770 585
R3170 gnd.n2772 gnd.n2771 585
R3171 gnd.n2769 gnd.n1195 585
R3172 gnd.n4892 gnd.n1195 585
R3173 gnd.n2768 gnd.n2767 585
R3174 gnd.n2767 gnd.n2766 585
R3175 gnd.n2678 gnd.n1185 585
R3176 gnd.n4898 gnd.n1185 585
R3177 gnd.n2677 gnd.n2676 585
R3178 gnd.n2676 gnd.n1177 585
R3179 gnd.n2675 gnd.n1175 585
R3180 gnd.n4904 gnd.n1175 585
R3181 gnd.n2674 gnd.n2673 585
R3182 gnd.n2673 gnd.n1167 585
R3183 gnd.n2671 gnd.n1165 585
R3184 gnd.n4910 gnd.n1165 585
R3185 gnd.n2670 gnd.n2669 585
R3186 gnd.n2669 gnd.n1155 585
R3187 gnd.n2668 gnd.n1153 585
R3188 gnd.n4916 gnd.n1153 585
R3189 gnd.n2667 gnd.n1141 585
R3190 gnd.n1152 gnd.n1141 585
R3191 gnd.n4923 gnd.n1139 585
R3192 gnd.n4923 gnd.n4922 585
R3193 gnd.n4925 gnd.n4924 585
R3194 gnd.n4924 gnd.n1068 585
R3195 gnd.n7556 gnd.n7555 585
R3196 gnd.n7557 gnd.n7556 585
R3197 gnd.n201 gnd.n200 585
R3198 gnd.n209 gnd.n201 585
R3199 gnd.n7565 gnd.n7564 585
R3200 gnd.n7564 gnd.n7563 585
R3201 gnd.n7566 gnd.n195 585
R3202 gnd.n195 gnd.n194 585
R3203 gnd.n7568 gnd.n7567 585
R3204 gnd.n7569 gnd.n7568 585
R3205 gnd.n182 gnd.n181 585
R3206 gnd.n185 gnd.n182 585
R3207 gnd.n7577 gnd.n7576 585
R3208 gnd.n7576 gnd.n7575 585
R3209 gnd.n7578 gnd.n176 585
R3210 gnd.n176 gnd.n175 585
R3211 gnd.n7580 gnd.n7579 585
R3212 gnd.n7581 gnd.n7580 585
R3213 gnd.n162 gnd.n161 585
R3214 gnd.n7392 gnd.n162 585
R3215 gnd.n7589 gnd.n7588 585
R3216 gnd.n7588 gnd.n7587 585
R3217 gnd.n7590 gnd.n156 585
R3218 gnd.n7371 gnd.n156 585
R3219 gnd.n7592 gnd.n7591 585
R3220 gnd.n7593 gnd.n7592 585
R3221 gnd.n142 gnd.n141 585
R3222 gnd.n7362 gnd.n142 585
R3223 gnd.n7601 gnd.n7600 585
R3224 gnd.n7600 gnd.n7599 585
R3225 gnd.n7602 gnd.n136 585
R3226 gnd.n7356 gnd.n136 585
R3227 gnd.n7604 gnd.n7603 585
R3228 gnd.n7605 gnd.n7604 585
R3229 gnd.n122 gnd.n121 585
R3230 gnd.n7348 gnd.n122 585
R3231 gnd.n7613 gnd.n7612 585
R3232 gnd.n7612 gnd.n7611 585
R3233 gnd.n7614 gnd.n117 585
R3234 gnd.n7342 gnd.n117 585
R3235 gnd.n7616 gnd.n7615 585
R3236 gnd.n7617 gnd.n7616 585
R3237 gnd.n101 gnd.n99 585
R3238 gnd.n7334 gnd.n101 585
R3239 gnd.n7625 gnd.n7624 585
R3240 gnd.n7624 gnd.n7623 585
R3241 gnd.n100 gnd.n92 585
R3242 gnd.n7328 gnd.n100 585
R3243 gnd.n7628 gnd.n90 585
R3244 gnd.n381 gnd.n90 585
R3245 gnd.n7630 gnd.n7629 585
R3246 gnd.n7631 gnd.n7630 585
R3247 gnd.n1725 gnd.n89 585
R3248 gnd.n4435 gnd.n89 585
R3249 gnd.n1727 gnd.n1726 585
R3250 gnd.n1732 gnd.n1727 585
R3251 gnd.n4472 gnd.n1728 585
R3252 gnd.n4472 gnd.n4471 585
R3253 gnd.n4473 gnd.n97 585
R3254 gnd.n4474 gnd.n4473 585
R3255 gnd.n1711 gnd.n1710 585
R3256 gnd.n4456 gnd.n1711 585
R3257 gnd.n4482 gnd.n4481 585
R3258 gnd.n4481 gnd.n4480 585
R3259 gnd.n4483 gnd.n1707 585
R3260 gnd.n4445 gnd.n1707 585
R3261 gnd.n4485 gnd.n4484 585
R3262 gnd.n4486 gnd.n4485 585
R3263 gnd.n1693 gnd.n1692 585
R3264 gnd.n4415 gnd.n1693 585
R3265 gnd.n4494 gnd.n4493 585
R3266 gnd.n4493 gnd.n4492 585
R3267 gnd.n4495 gnd.n1687 585
R3268 gnd.n4374 gnd.n1687 585
R3269 gnd.n4497 gnd.n4496 585
R3270 gnd.n4498 gnd.n4497 585
R3271 gnd.n1673 gnd.n1672 585
R3272 gnd.n4367 gnd.n1673 585
R3273 gnd.n4506 gnd.n4505 585
R3274 gnd.n4505 gnd.n4504 585
R3275 gnd.n4507 gnd.n1667 585
R3276 gnd.n4362 gnd.n1667 585
R3277 gnd.n4509 gnd.n4508 585
R3278 gnd.n4510 gnd.n4509 585
R3279 gnd.n1653 gnd.n1652 585
R3280 gnd.n4391 gnd.n1653 585
R3281 gnd.n4518 gnd.n4517 585
R3282 gnd.n4517 gnd.n4516 585
R3283 gnd.n4519 gnd.n1647 585
R3284 gnd.n4355 gnd.n1647 585
R3285 gnd.n4521 gnd.n4520 585
R3286 gnd.n4522 gnd.n4521 585
R3287 gnd.n1633 gnd.n1632 585
R3288 gnd.n4347 gnd.n1633 585
R3289 gnd.n4530 gnd.n4529 585
R3290 gnd.n4529 gnd.n4528 585
R3291 gnd.n4531 gnd.n1627 585
R3292 gnd.n4341 gnd.n1627 585
R3293 gnd.n4533 gnd.n4532 585
R3294 gnd.n4534 gnd.n4533 585
R3295 gnd.n1610 gnd.n1609 585
R3296 gnd.n4333 gnd.n1610 585
R3297 gnd.n4542 gnd.n4541 585
R3298 gnd.n4541 gnd.n4540 585
R3299 gnd.n4543 gnd.n1605 585
R3300 gnd.n3754 gnd.n1605 585
R3301 gnd.n4545 gnd.n4544 585
R3302 gnd.n4546 gnd.n4545 585
R3303 gnd.n4174 gnd.n1604 585
R3304 gnd.n4179 gnd.n4177 585
R3305 gnd.n4180 gnd.n4173 585
R3306 gnd.n4180 gnd.n1591 585
R3307 gnd.n4183 gnd.n4182 585
R3308 gnd.n4171 gnd.n4170 585
R3309 gnd.n4188 gnd.n4187 585
R3310 gnd.n4190 gnd.n4169 585
R3311 gnd.n4193 gnd.n4192 585
R3312 gnd.n4167 gnd.n4166 585
R3313 gnd.n4198 gnd.n4197 585
R3314 gnd.n4200 gnd.n4165 585
R3315 gnd.n4203 gnd.n4202 585
R3316 gnd.n4163 gnd.n4162 585
R3317 gnd.n4208 gnd.n4207 585
R3318 gnd.n4210 gnd.n4161 585
R3319 gnd.n4213 gnd.n4212 585
R3320 gnd.n4159 gnd.n4158 585
R3321 gnd.n4221 gnd.n4220 585
R3322 gnd.n4223 gnd.n4157 585
R3323 gnd.n4226 gnd.n4225 585
R3324 gnd.n4155 gnd.n4154 585
R3325 gnd.n4231 gnd.n4230 585
R3326 gnd.n4233 gnd.n4153 585
R3327 gnd.n4236 gnd.n4235 585
R3328 gnd.n4151 gnd.n4150 585
R3329 gnd.n4242 gnd.n4241 585
R3330 gnd.n4246 gnd.n1841 585
R3331 gnd.n4249 gnd.n4248 585
R3332 gnd.n1839 gnd.n1838 585
R3333 gnd.n4254 gnd.n4253 585
R3334 gnd.n4256 gnd.n1837 585
R3335 gnd.n4259 gnd.n4258 585
R3336 gnd.n1835 gnd.n1834 585
R3337 gnd.n4264 gnd.n4263 585
R3338 gnd.n4266 gnd.n1833 585
R3339 gnd.n4271 gnd.n4268 585
R3340 gnd.n1831 gnd.n1830 585
R3341 gnd.n4276 gnd.n4275 585
R3342 gnd.n4278 gnd.n1829 585
R3343 gnd.n4281 gnd.n4280 585
R3344 gnd.n1827 gnd.n1826 585
R3345 gnd.n4286 gnd.n4285 585
R3346 gnd.n4288 gnd.n1825 585
R3347 gnd.n4291 gnd.n4290 585
R3348 gnd.n1823 gnd.n1822 585
R3349 gnd.n4296 gnd.n4295 585
R3350 gnd.n4298 gnd.n1821 585
R3351 gnd.n4301 gnd.n4300 585
R3352 gnd.n1819 gnd.n1818 585
R3353 gnd.n4306 gnd.n4305 585
R3354 gnd.n4308 gnd.n1817 585
R3355 gnd.n4311 gnd.n4310 585
R3356 gnd.n1815 gnd.n1814 585
R3357 gnd.n4317 gnd.n4316 585
R3358 gnd.n4319 gnd.n1813 585
R3359 gnd.n4320 gnd.n1812 585
R3360 gnd.n4323 gnd.n4322 585
R3361 gnd.n7447 gnd.n7446 585
R3362 gnd.n7449 gnd.n315 585
R3363 gnd.n7451 gnd.n7450 585
R3364 gnd.n7452 gnd.n308 585
R3365 gnd.n7454 gnd.n7453 585
R3366 gnd.n7456 gnd.n306 585
R3367 gnd.n7458 gnd.n7457 585
R3368 gnd.n7459 gnd.n301 585
R3369 gnd.n7461 gnd.n7460 585
R3370 gnd.n7463 gnd.n299 585
R3371 gnd.n7465 gnd.n7464 585
R3372 gnd.n7466 gnd.n294 585
R3373 gnd.n7468 gnd.n7467 585
R3374 gnd.n7470 gnd.n292 585
R3375 gnd.n7472 gnd.n7471 585
R3376 gnd.n7473 gnd.n287 585
R3377 gnd.n7475 gnd.n7474 585
R3378 gnd.n7477 gnd.n286 585
R3379 gnd.n7478 gnd.n283 585
R3380 gnd.n7481 gnd.n7480 585
R3381 gnd.n285 gnd.n279 585
R3382 gnd.n7485 gnd.n276 585
R3383 gnd.n7487 gnd.n7486 585
R3384 gnd.n7489 gnd.n274 585
R3385 gnd.n7491 gnd.n7490 585
R3386 gnd.n7492 gnd.n269 585
R3387 gnd.n7494 gnd.n7493 585
R3388 gnd.n7496 gnd.n267 585
R3389 gnd.n7498 gnd.n7497 585
R3390 gnd.n7499 gnd.n262 585
R3391 gnd.n7501 gnd.n7500 585
R3392 gnd.n7503 gnd.n260 585
R3393 gnd.n7505 gnd.n7504 585
R3394 gnd.n7506 gnd.n255 585
R3395 gnd.n7508 gnd.n7507 585
R3396 gnd.n7510 gnd.n253 585
R3397 gnd.n7512 gnd.n7511 585
R3398 gnd.n7513 gnd.n248 585
R3399 gnd.n7515 gnd.n7514 585
R3400 gnd.n7517 gnd.n246 585
R3401 gnd.n7519 gnd.n7518 585
R3402 gnd.n7523 gnd.n241 585
R3403 gnd.n7525 gnd.n7524 585
R3404 gnd.n7527 gnd.n239 585
R3405 gnd.n7529 gnd.n7528 585
R3406 gnd.n7530 gnd.n234 585
R3407 gnd.n7532 gnd.n7531 585
R3408 gnd.n7534 gnd.n232 585
R3409 gnd.n7536 gnd.n7535 585
R3410 gnd.n7537 gnd.n227 585
R3411 gnd.n7539 gnd.n7538 585
R3412 gnd.n7541 gnd.n225 585
R3413 gnd.n7543 gnd.n7542 585
R3414 gnd.n7544 gnd.n220 585
R3415 gnd.n7546 gnd.n7545 585
R3416 gnd.n7548 gnd.n218 585
R3417 gnd.n7550 gnd.n7549 585
R3418 gnd.n7551 gnd.n216 585
R3419 gnd.n7552 gnd.n213 585
R3420 gnd.n213 gnd.n212 585
R3421 gnd.n7377 gnd.n210 585
R3422 gnd.n7557 gnd.n210 585
R3423 gnd.n7379 gnd.n7378 585
R3424 gnd.n7378 gnd.n209 585
R3425 gnd.n7380 gnd.n202 585
R3426 gnd.n7563 gnd.n202 585
R3427 gnd.n7382 gnd.n7381 585
R3428 gnd.n7381 gnd.n194 585
R3429 gnd.n7383 gnd.n192 585
R3430 gnd.n7569 gnd.n192 585
R3431 gnd.n7385 gnd.n7384 585
R3432 gnd.n7384 gnd.n185 585
R3433 gnd.n7386 gnd.n183 585
R3434 gnd.n7575 gnd.n183 585
R3435 gnd.n7388 gnd.n7387 585
R3436 gnd.n7387 gnd.n175 585
R3437 gnd.n7389 gnd.n173 585
R3438 gnd.n7581 gnd.n173 585
R3439 gnd.n7391 gnd.n7390 585
R3440 gnd.n7392 gnd.n7391 585
R3441 gnd.n7374 gnd.n164 585
R3442 gnd.n7587 gnd.n164 585
R3443 gnd.n7373 gnd.n7372 585
R3444 gnd.n7372 gnd.n7371 585
R3445 gnd.n360 gnd.n154 585
R3446 gnd.n7593 gnd.n154 585
R3447 gnd.n7361 gnd.n7360 585
R3448 gnd.n7362 gnd.n7361 585
R3449 gnd.n7359 gnd.n144 585
R3450 gnd.n7599 gnd.n144 585
R3451 gnd.n7358 gnd.n7357 585
R3452 gnd.n7357 gnd.n7356 585
R3453 gnd.n366 gnd.n133 585
R3454 gnd.n7605 gnd.n133 585
R3455 gnd.n7347 gnd.n7346 585
R3456 gnd.n7348 gnd.n7347 585
R3457 gnd.n7345 gnd.n124 585
R3458 gnd.n7611 gnd.n124 585
R3459 gnd.n7344 gnd.n7343 585
R3460 gnd.n7343 gnd.n7342 585
R3461 gnd.n372 gnd.n115 585
R3462 gnd.n7617 gnd.n115 585
R3463 gnd.n7333 gnd.n7332 585
R3464 gnd.n7334 gnd.n7333 585
R3465 gnd.n7331 gnd.n103 585
R3466 gnd.n7623 gnd.n103 585
R3467 gnd.n7330 gnd.n7329 585
R3468 gnd.n7329 gnd.n7328 585
R3469 gnd.n380 gnd.n378 585
R3470 gnd.n381 gnd.n380 585
R3471 gnd.n4427 gnd.n86 585
R3472 gnd.n7631 gnd.n86 585
R3473 gnd.n4436 gnd.n4422 585
R3474 gnd.n4436 gnd.n4435 585
R3475 gnd.n4438 gnd.n4437 585
R3476 gnd.n4437 gnd.n1732 585
R3477 gnd.n4439 gnd.n1729 585
R3478 gnd.n4471 gnd.n1729 585
R3479 gnd.n4440 gnd.n1722 585
R3480 gnd.n4474 gnd.n1722 585
R3481 gnd.n4441 gnd.n1737 585
R3482 gnd.n4456 gnd.n1737 585
R3483 gnd.n4442 gnd.n1713 585
R3484 gnd.n4480 gnd.n1713 585
R3485 gnd.n4444 gnd.n4443 585
R3486 gnd.n4445 gnd.n4444 585
R3487 gnd.n4418 gnd.n1704 585
R3488 gnd.n4486 gnd.n1704 585
R3489 gnd.n4417 gnd.n4416 585
R3490 gnd.n4416 gnd.n4415 585
R3491 gnd.n1742 gnd.n1695 585
R3492 gnd.n4492 gnd.n1695 585
R3493 gnd.n4373 gnd.n4372 585
R3494 gnd.n4374 gnd.n4373 585
R3495 gnd.n4370 gnd.n1684 585
R3496 gnd.n4498 gnd.n1684 585
R3497 gnd.n4369 gnd.n4368 585
R3498 gnd.n4368 gnd.n4367 585
R3499 gnd.n4365 gnd.n1675 585
R3500 gnd.n4504 gnd.n1675 585
R3501 gnd.n4364 gnd.n4363 585
R3502 gnd.n4363 gnd.n4362 585
R3503 gnd.n4360 gnd.n1664 585
R3504 gnd.n4510 gnd.n1664 585
R3505 gnd.n4359 gnd.n1755 585
R3506 gnd.n4391 gnd.n1755 585
R3507 gnd.n4358 gnd.n1655 585
R3508 gnd.n4516 gnd.n1655 585
R3509 gnd.n4357 gnd.n4356 585
R3510 gnd.n4356 gnd.n4355 585
R3511 gnd.n1764 gnd.n1644 585
R3512 gnd.n4522 gnd.n1644 585
R3513 gnd.n4346 gnd.n4345 585
R3514 gnd.n4347 gnd.n4346 585
R3515 gnd.n4344 gnd.n1635 585
R3516 gnd.n4528 gnd.n1635 585
R3517 gnd.n4343 gnd.n4342 585
R3518 gnd.n4342 gnd.n4341 585
R3519 gnd.n1801 gnd.n1624 585
R3520 gnd.n4534 gnd.n1624 585
R3521 gnd.n4332 gnd.n4331 585
R3522 gnd.n4333 gnd.n4332 585
R3523 gnd.n4330 gnd.n1612 585
R3524 gnd.n4540 gnd.n1612 585
R3525 gnd.n4329 gnd.n1807 585
R3526 gnd.n3754 gnd.n1807 585
R3527 gnd.n1806 gnd.n1600 585
R3528 gnd.n4546 gnd.n1600 585
R3529 gnd.n2787 gnd.n2785 585
R3530 gnd.n2785 gnd.n1184 585
R3531 gnd.n7298 gnd.n7297 585
R3532 gnd.n7297 gnd.n172 585
R3533 gnd.n7301 gnd.n399 585
R3534 gnd.n399 gnd.n163 585
R3535 gnd.n7303 gnd.n7302 585
R3536 gnd.n7303 gnd.n362 585
R3537 gnd.n7304 gnd.n398 585
R3538 gnd.n7304 gnd.n153 585
R3539 gnd.n7306 gnd.n7305 585
R3540 gnd.n7305 gnd.n146 585
R3541 gnd.n7307 gnd.n393 585
R3542 gnd.n393 gnd.n143 585
R3543 gnd.n7309 gnd.n7308 585
R3544 gnd.n7309 gnd.n135 585
R3545 gnd.n7310 gnd.n392 585
R3546 gnd.n7310 gnd.n132 585
R3547 gnd.n7312 gnd.n7311 585
R3548 gnd.n7311 gnd.n371 585
R3549 gnd.n7313 gnd.n387 585
R3550 gnd.n387 gnd.n123 585
R3551 gnd.n7315 gnd.n7314 585
R3552 gnd.n7315 gnd.n374 585
R3553 gnd.n7316 gnd.n386 585
R3554 gnd.n7316 gnd.n114 585
R3555 gnd.n7318 gnd.n7317 585
R3556 gnd.n7317 gnd.n105 585
R3557 gnd.n7319 gnd.n383 585
R3558 gnd.n383 gnd.n102 585
R3559 gnd.n7322 gnd.n7321 585
R3560 gnd.n7323 gnd.n7322 585
R3561 gnd.n384 gnd.n382 585
R3562 gnd.n382 gnd.n87 585
R3563 gnd.n4465 gnd.n4464 585
R3564 gnd.n4464 gnd.n85 585
R3565 gnd.n4466 gnd.n1734 585
R3566 gnd.n4423 gnd.n1734 585
R3567 gnd.n4469 gnd.n4468 585
R3568 gnd.n4470 gnd.n4469 585
R3569 gnd.n4462 gnd.n1733 585
R3570 gnd.n1733 gnd.n1724 585
R3571 gnd.n4460 gnd.n4459 585
R3572 gnd.n4459 gnd.n1721 585
R3573 gnd.n4458 gnd.n1735 585
R3574 gnd.n4458 gnd.n4457 585
R3575 gnd.n4410 gnd.n1736 585
R3576 gnd.n1736 gnd.n1712 585
R3577 gnd.n4411 gnd.n1745 585
R3578 gnd.n1745 gnd.n1706 585
R3579 gnd.n4413 gnd.n4412 585
R3580 gnd.n4414 gnd.n4413 585
R3581 gnd.n1746 gnd.n1744 585
R3582 gnd.n1744 gnd.n1697 585
R3583 gnd.n4404 gnd.n4403 585
R3584 gnd.n4403 gnd.n1694 585
R3585 gnd.n4402 gnd.n1748 585
R3586 gnd.n4402 gnd.n1686 585
R3587 gnd.n4401 gnd.n4400 585
R3588 gnd.n4401 gnd.n1683 585
R3589 gnd.n1750 gnd.n1749 585
R3590 gnd.n4366 gnd.n1749 585
R3591 gnd.n4396 gnd.n4395 585
R3592 gnd.n4395 gnd.n1674 585
R3593 gnd.n4394 gnd.n1752 585
R3594 gnd.n4394 gnd.n1666 585
R3595 gnd.n4393 gnd.n1754 585
R3596 gnd.n4393 gnd.n4392 585
R3597 gnd.n1792 gnd.n1753 585
R3598 gnd.n1753 gnd.n1657 585
R3599 gnd.n1794 gnd.n1793 585
R3600 gnd.n1794 gnd.n1654 585
R3601 gnd.n1796 gnd.n1795 585
R3602 gnd.n1795 gnd.n1646 585
R3603 gnd.n1797 gnd.n1770 585
R3604 gnd.n1770 gnd.n1643 585
R3605 gnd.n1799 gnd.n1798 585
R3606 gnd.n1800 gnd.n1799 585
R3607 gnd.n1771 gnd.n1769 585
R3608 gnd.n1769 gnd.n1634 585
R3609 gnd.n1783 gnd.n1782 585
R3610 gnd.n1782 gnd.n1626 585
R3611 gnd.n1781 gnd.n1773 585
R3612 gnd.n1781 gnd.n1623 585
R3613 gnd.n1780 gnd.n1779 585
R3614 gnd.n1780 gnd.n1614 585
R3615 gnd.n1775 gnd.n1774 585
R3616 gnd.n1774 gnd.n1611 585
R3617 gnd.n1598 gnd.n1597 585
R3618 gnd.n1602 gnd.n1598 585
R3619 gnd.n4549 gnd.n4548 585
R3620 gnd.n4548 gnd.n4547 585
R3621 gnd.n4550 gnd.n1592 585
R3622 gnd.n1599 gnd.n1592 585
R3623 gnd.n4552 gnd.n4551 585
R3624 gnd.n4553 gnd.n4552 585
R3625 gnd.n1589 gnd.n1588 585
R3626 gnd.n4554 gnd.n1589 585
R3627 gnd.n4557 gnd.n4556 585
R3628 gnd.n4556 gnd.n4555 585
R3629 gnd.n4558 gnd.n1583 585
R3630 gnd.n1583 gnd.n1581 585
R3631 gnd.n4560 gnd.n4559 585
R3632 gnd.n4561 gnd.n4560 585
R3633 gnd.n1584 gnd.n1582 585
R3634 gnd.n1582 gnd.n1579 585
R3635 gnd.n3940 gnd.n3939 585
R3636 gnd.n3941 gnd.n3940 585
R3637 gnd.n1933 gnd.n1932 585
R3638 gnd.n3943 gnd.n1933 585
R3639 gnd.n3948 gnd.n3947 585
R3640 gnd.n3947 gnd.n3946 585
R3641 gnd.n3949 gnd.n1927 585
R3642 gnd.n1934 gnd.n1927 585
R3643 gnd.n3951 gnd.n3950 585
R3644 gnd.n3952 gnd.n3951 585
R3645 gnd.n1921 gnd.n1920 585
R3646 gnd.n3954 gnd.n1921 585
R3647 gnd.n3959 gnd.n3958 585
R3648 gnd.n3958 gnd.n3957 585
R3649 gnd.n3960 gnd.n1915 585
R3650 gnd.n1922 gnd.n1915 585
R3651 gnd.n3962 gnd.n3961 585
R3652 gnd.n3963 gnd.n3962 585
R3653 gnd.n1909 gnd.n1908 585
R3654 gnd.n3965 gnd.n1909 585
R3655 gnd.n3970 gnd.n3969 585
R3656 gnd.n3969 gnd.n3968 585
R3657 gnd.n3971 gnd.n1903 585
R3658 gnd.n1910 gnd.n1903 585
R3659 gnd.n3973 gnd.n3972 585
R3660 gnd.n3974 gnd.n3973 585
R3661 gnd.n1899 gnd.n1898 585
R3662 gnd.n3976 gnd.n1899 585
R3663 gnd.n3981 gnd.n3980 585
R3664 gnd.n3980 gnd.n3979 585
R3665 gnd.n3982 gnd.n1893 585
R3666 gnd.n1893 gnd.n1884 585
R3667 gnd.n3984 gnd.n3983 585
R3668 gnd.n3985 gnd.n3984 585
R3669 gnd.n1894 gnd.n1892 585
R3670 gnd.n1892 gnd.n1889 585
R3671 gnd.n3694 gnd.n3693 585
R3672 gnd.n3693 gnd.n1951 585
R3673 gnd.n3695 gnd.n1967 585
R3674 gnd.n1967 gnd.n1955 585
R3675 gnd.n3697 gnd.n3696 585
R3676 gnd.n3698 gnd.n3697 585
R3677 gnd.n1968 gnd.n1966 585
R3678 gnd.n1975 gnd.n1966 585
R3679 gnd.n3686 gnd.n3685 585
R3680 gnd.n3685 gnd.n3684 585
R3681 gnd.n1971 gnd.n1970 585
R3682 gnd.n3588 gnd.n1971 585
R3683 gnd.n3646 gnd.n1995 585
R3684 gnd.n1995 gnd.n1988 585
R3685 gnd.n3648 gnd.n3647 585
R3686 gnd.n3649 gnd.n3648 585
R3687 gnd.n1996 gnd.n1994 585
R3688 gnd.n1994 gnd.n1992 585
R3689 gnd.n3641 gnd.n3640 585
R3690 gnd.n3640 gnd.n3639 585
R3691 gnd.n1999 gnd.n1998 585
R3692 gnd.n3631 gnd.n1999 585
R3693 gnd.n3617 gnd.n3616 585
R3694 gnd.n3618 gnd.n3617 585
R3695 gnd.n2018 gnd.n2017 585
R3696 gnd.n3568 gnd.n2017 585
R3697 gnd.n3612 gnd.n3611 585
R3698 gnd.n3611 gnd.n3610 585
R3699 gnd.n2021 gnd.n2020 585
R3700 gnd.n2029 gnd.n2021 585
R3701 gnd.n3557 gnd.n3556 585
R3702 gnd.n3558 gnd.n3557 585
R3703 gnd.n2038 gnd.n2037 585
R3704 gnd.n2037 gnd.n2034 585
R3705 gnd.n3552 gnd.n3551 585
R3706 gnd.n3551 gnd.n3550 585
R3707 gnd.n2041 gnd.n2040 585
R3708 gnd.n2047 gnd.n2041 585
R3709 gnd.n3532 gnd.n3531 585
R3710 gnd.n3533 gnd.n3532 585
R3711 gnd.n2057 gnd.n2056 585
R3712 gnd.n2064 gnd.n2056 585
R3713 gnd.n3527 gnd.n3526 585
R3714 gnd.n3526 gnd.n3525 585
R3715 gnd.n2060 gnd.n2059 585
R3716 gnd.n2068 gnd.n2060 585
R3717 gnd.n3476 gnd.n3475 585
R3718 gnd.n3477 gnd.n3476 585
R3719 gnd.n2079 gnd.n2078 585
R3720 gnd.n2097 gnd.n2078 585
R3721 gnd.n3471 gnd.n3470 585
R3722 gnd.n3470 gnd.n3469 585
R3723 gnd.n2082 gnd.n2081 585
R3724 gnd.n2090 gnd.n2082 585
R3725 gnd.n3436 gnd.n3435 585
R3726 gnd.n3437 gnd.n3436 585
R3727 gnd.n2102 gnd.n2101 585
R3728 gnd.n2117 gnd.n2101 585
R3729 gnd.n3431 gnd.n3430 585
R3730 gnd.n3430 gnd.n3429 585
R3731 gnd.n2105 gnd.n2104 585
R3732 gnd.n3419 gnd.n2105 585
R3733 gnd.n3385 gnd.n2134 585
R3734 gnd.n2134 gnd.n2126 585
R3735 gnd.n3387 gnd.n3386 585
R3736 gnd.n3388 gnd.n3387 585
R3737 gnd.n2135 gnd.n2133 585
R3738 gnd.n2133 gnd.n2130 585
R3739 gnd.n3380 gnd.n3379 585
R3740 gnd.n3379 gnd.n3378 585
R3741 gnd.n2138 gnd.n2137 585
R3742 gnd.n2144 gnd.n2138 585
R3743 gnd.n3358 gnd.n3357 585
R3744 gnd.n3359 gnd.n3358 585
R3745 gnd.n2153 gnd.n2152 585
R3746 gnd.n2159 gnd.n2152 585
R3747 gnd.n3353 gnd.n3352 585
R3748 gnd.n3352 gnd.n3351 585
R3749 gnd.n2156 gnd.n2155 585
R3750 gnd.n2163 gnd.n2156 585
R3751 gnd.n3296 gnd.n2178 585
R3752 gnd.n2178 gnd.n2168 585
R3753 gnd.n3298 gnd.n3297 585
R3754 gnd.n3299 gnd.n3298 585
R3755 gnd.n2179 gnd.n2177 585
R3756 gnd.n3273 gnd.n2177 585
R3757 gnd.n3291 gnd.n3290 585
R3758 gnd.n3290 gnd.n3289 585
R3759 gnd.n2182 gnd.n2181 585
R3760 gnd.n3263 gnd.n2182 585
R3761 gnd.n3226 gnd.n3225 585
R3762 gnd.n3226 gnd.n1490 585
R3763 gnd.n3228 gnd.n3222 585
R3764 gnd.n3228 gnd.n3227 585
R3765 gnd.n3230 gnd.n3229 585
R3766 gnd.n3229 gnd.n2260 585
R3767 gnd.n3231 gnd.n2272 585
R3768 gnd.n2272 gnd.n2259 585
R3769 gnd.n3233 gnd.n3232 585
R3770 gnd.n3234 gnd.n3233 585
R3771 gnd.n2273 gnd.n2271 585
R3772 gnd.n2271 gnd.n2268 585
R3773 gnd.n3216 gnd.n3215 585
R3774 gnd.n3215 gnd.n3214 585
R3775 gnd.n2276 gnd.n2275 585
R3776 gnd.n2285 gnd.n2276 585
R3777 gnd.n3191 gnd.n2297 585
R3778 gnd.n2297 gnd.n2284 585
R3779 gnd.n3193 gnd.n3192 585
R3780 gnd.n3194 gnd.n3193 585
R3781 gnd.n2298 gnd.n2296 585
R3782 gnd.n2296 gnd.n2293 585
R3783 gnd.n3186 gnd.n3185 585
R3784 gnd.n3185 gnd.n3184 585
R3785 gnd.n2301 gnd.n2300 585
R3786 gnd.n2309 gnd.n2301 585
R3787 gnd.n3161 gnd.n2322 585
R3788 gnd.n2322 gnd.n2308 585
R3789 gnd.n3163 gnd.n3162 585
R3790 gnd.n3164 gnd.n3163 585
R3791 gnd.n2323 gnd.n2321 585
R3792 gnd.n2321 gnd.n2318 585
R3793 gnd.n3156 gnd.n3155 585
R3794 gnd.n3155 gnd.n3154 585
R3795 gnd.n2326 gnd.n2325 585
R3796 gnd.n2334 gnd.n2326 585
R3797 gnd.n3065 gnd.n2553 585
R3798 gnd.n2553 gnd.n2333 585
R3799 gnd.n3067 gnd.n3066 585
R3800 gnd.n3068 gnd.n3067 585
R3801 gnd.n2554 gnd.n2552 585
R3802 gnd.n2552 gnd.n2530 585
R3803 gnd.n3060 gnd.n3059 585
R3804 gnd.n3059 gnd.n3058 585
R3805 gnd.n3056 gnd.n2556 585
R3806 gnd.n3057 gnd.n3056 585
R3807 gnd.n3055 gnd.n3053 585
R3808 gnd.n3055 gnd.n3054 585
R3809 gnd.n2558 gnd.n2557 585
R3810 gnd.n2557 gnd.n1376 585
R3811 gnd.n3049 gnd.n3048 585
R3812 gnd.n3048 gnd.n1373 585
R3813 gnd.n3047 gnd.n2560 585
R3814 gnd.n3047 gnd.n1367 585
R3815 gnd.n3046 gnd.n3045 585
R3816 gnd.n3046 gnd.n1364 585
R3817 gnd.n2562 gnd.n2561 585
R3818 gnd.n2561 gnd.n1356 585
R3819 gnd.n3041 gnd.n3040 585
R3820 gnd.n3040 gnd.n1353 585
R3821 gnd.n3039 gnd.n2564 585
R3822 gnd.n3039 gnd.n1346 585
R3823 gnd.n3038 gnd.n2566 585
R3824 gnd.n3038 gnd.n3037 585
R3825 gnd.n2966 gnd.n2565 585
R3826 gnd.n2565 gnd.n1336 585
R3827 gnd.n2968 gnd.n2967 585
R3828 gnd.n2967 gnd.n1333 585
R3829 gnd.n2969 gnd.n2959 585
R3830 gnd.n2959 gnd.n1326 585
R3831 gnd.n2971 gnd.n2970 585
R3832 gnd.n2971 gnd.n1323 585
R3833 gnd.n2972 gnd.n2958 585
R3834 gnd.n2972 gnd.n2580 585
R3835 gnd.n2974 gnd.n2973 585
R3836 gnd.n2973 gnd.n1313 585
R3837 gnd.n2975 gnd.n2587 585
R3838 gnd.n2587 gnd.n1306 585
R3839 gnd.n2977 gnd.n2976 585
R3840 gnd.n2978 gnd.n2977 585
R3841 gnd.n2588 gnd.n2586 585
R3842 gnd.n2586 gnd.n1296 585
R3843 gnd.n2952 gnd.n2951 585
R3844 gnd.n2951 gnd.n1293 585
R3845 gnd.n2950 gnd.n2590 585
R3846 gnd.n2950 gnd.n1286 585
R3847 gnd.n2949 gnd.n2948 585
R3848 gnd.n2949 gnd.n1283 585
R3849 gnd.n2592 gnd.n2591 585
R3850 gnd.n2915 gnd.n2591 585
R3851 gnd.n2944 gnd.n2943 585
R3852 gnd.n2943 gnd.n1274 585
R3853 gnd.n2942 gnd.n2593 585
R3854 gnd.n2942 gnd.n1265 585
R3855 gnd.n2941 gnd.n2596 585
R3856 gnd.n2941 gnd.n2940 585
R3857 gnd.n2872 gnd.n2594 585
R3858 gnd.n2597 gnd.n2594 585
R3859 gnd.n2874 gnd.n2635 585
R3860 gnd.n2635 gnd.n2611 585
R3861 gnd.n2876 gnd.n2875 585
R3862 gnd.n2877 gnd.n2876 585
R3863 gnd.n2870 gnd.n2634 585
R3864 gnd.n2634 gnd.n2621 585
R3865 gnd.n2869 gnd.n2868 585
R3866 gnd.n2868 gnd.n2627 585
R3867 gnd.n2867 gnd.n2866 585
R3868 gnd.n2867 gnd.n2625 585
R3869 gnd.n2865 gnd.n2637 585
R3870 gnd.n2643 gnd.n2637 585
R3871 gnd.n2863 gnd.n2862 585
R3872 gnd.n2862 gnd.n2861 585
R3873 gnd.n2639 gnd.n2638 585
R3874 gnd.n2639 gnd.n1248 585
R3875 gnd.n2808 gnd.n2807 585
R3876 gnd.n2807 gnd.n1245 585
R3877 gnd.n2809 gnd.n2801 585
R3878 gnd.n2801 gnd.n1238 585
R3879 gnd.n2811 gnd.n2810 585
R3880 gnd.n2811 gnd.n1235 585
R3881 gnd.n2812 gnd.n2800 585
R3882 gnd.n2812 gnd.n1227 585
R3883 gnd.n2814 gnd.n2813 585
R3884 gnd.n2813 gnd.n1224 585
R3885 gnd.n2815 gnd.n2781 585
R3886 gnd.n2781 gnd.n1217 585
R3887 gnd.n2817 gnd.n2816 585
R3888 gnd.n2818 gnd.n2817 585
R3889 gnd.n2782 gnd.n2780 585
R3890 gnd.n2780 gnd.n1207 585
R3891 gnd.n2794 gnd.n2793 585
R3892 gnd.n2793 gnd.n1204 585
R3893 gnd.n2792 gnd.n2784 585
R3894 gnd.n2792 gnd.n1197 585
R3895 gnd.n2791 gnd.n2790 585
R3896 gnd.n2791 gnd.n1194 585
R3897 gnd.n4564 gnd.n4563 585
R3898 gnd.n4563 gnd.n4562 585
R3899 gnd.n4565 gnd.n1576 585
R3900 gnd.n3935 gnd.n1576 585
R3901 gnd.n4566 gnd.n1575 585
R3902 gnd.n3942 gnd.n1575 585
R3903 gnd.n3944 gnd.n1573 585
R3904 gnd.n3945 gnd.n3944 585
R3905 gnd.n4570 gnd.n1572 585
R3906 gnd.n1935 gnd.n1572 585
R3907 gnd.n4571 gnd.n1571 585
R3908 gnd.n1926 gnd.n1571 585
R3909 gnd.n4572 gnd.n1570 585
R3910 gnd.n3953 gnd.n1570 585
R3911 gnd.n3955 gnd.n1568 585
R3912 gnd.n3956 gnd.n3955 585
R3913 gnd.n4576 gnd.n1567 585
R3914 gnd.n1923 gnd.n1567 585
R3915 gnd.n4577 gnd.n1566 585
R3916 gnd.n1914 gnd.n1566 585
R3917 gnd.n4578 gnd.n1565 585
R3918 gnd.n3964 gnd.n1565 585
R3919 gnd.n3966 gnd.n1563 585
R3920 gnd.n3967 gnd.n3966 585
R3921 gnd.n4582 gnd.n1562 585
R3922 gnd.n1911 gnd.n1562 585
R3923 gnd.n4583 gnd.n1561 585
R3924 gnd.n1902 gnd.n1561 585
R3925 gnd.n4584 gnd.n1560 585
R3926 gnd.n3975 gnd.n1560 585
R3927 gnd.n3977 gnd.n1558 585
R3928 gnd.n3978 gnd.n3977 585
R3929 gnd.n4588 gnd.n1557 585
R3930 gnd.n1846 gnd.n1557 585
R3931 gnd.n4589 gnd.n1556 585
R3932 gnd.n1883 gnd.n1556 585
R3933 gnd.n4590 gnd.n1555 585
R3934 gnd.n3987 gnd.n1555 585
R3935 gnd.n3715 gnd.n1553 585
R3936 gnd.n3716 gnd.n3715 585
R3937 gnd.n4594 gnd.n1552 585
R3938 gnd.n1957 gnd.n1552 585
R3939 gnd.n4595 gnd.n1551 585
R3940 gnd.n1965 gnd.n1551 585
R3941 gnd.n4596 gnd.n1550 585
R3942 gnd.n1962 gnd.n1550 585
R3943 gnd.n3682 gnd.n1548 585
R3944 gnd.n3683 gnd.n3682 585
R3945 gnd.n4600 gnd.n1547 585
R3946 gnd.n3674 gnd.n1547 585
R3947 gnd.n4601 gnd.n1546 585
R3948 gnd.n3589 gnd.n1546 585
R3949 gnd.n4602 gnd.n1545 585
R3950 gnd.n3659 gnd.n1545 585
R3951 gnd.n3650 gnd.n1543 585
R3952 gnd.n3651 gnd.n3650 585
R3953 gnd.n4606 gnd.n1542 585
R3954 gnd.n2001 gnd.n1542 585
R3955 gnd.n4607 gnd.n1541 585
R3956 gnd.n3629 gnd.n1541 585
R3957 gnd.n4608 gnd.n1540 585
R3958 gnd.n2005 gnd.n1540 585
R3959 gnd.n3619 gnd.n1538 585
R3960 gnd.n3620 gnd.n3619 585
R3961 gnd.n4612 gnd.n1537 585
R3962 gnd.n2023 gnd.n1537 585
R3963 gnd.n4613 gnd.n1536 585
R3964 gnd.n3499 gnd.n1536 585
R3965 gnd.n4614 gnd.n1535 585
R3966 gnd.n2028 gnd.n1535 585
R3967 gnd.n3560 gnd.n1533 585
R3968 gnd.n3561 gnd.n3560 585
R3969 gnd.n4618 gnd.n1532 585
R3970 gnd.n3549 gnd.n1532 585
R3971 gnd.n4619 gnd.n1531 585
R3972 gnd.n2048 gnd.n1531 585
R3973 gnd.n4620 gnd.n1530 585
R3974 gnd.n2055 gnd.n1530 585
R3975 gnd.n3490 gnd.n1528 585
R3976 gnd.n3491 gnd.n3490 585
R3977 gnd.n4624 gnd.n1527 585
R3978 gnd.n3524 gnd.n1527 585
R3979 gnd.n4625 gnd.n1526 585
R3980 gnd.n3516 gnd.n1526 585
R3981 gnd.n4626 gnd.n1525 585
R3982 gnd.n3478 gnd.n1525 585
R3983 gnd.n3449 gnd.n1523 585
R3984 gnd.n3450 gnd.n3449 585
R3985 gnd.n4630 gnd.n1522 585
R3986 gnd.n2085 gnd.n1522 585
R3987 gnd.n4631 gnd.n1521 585
R3988 gnd.n3458 gnd.n1521 585
R3989 gnd.n4632 gnd.n1520 585
R3990 gnd.n3438 gnd.n1520 585
R3991 gnd.n3410 gnd.n1518 585
R3992 gnd.n3411 gnd.n3410 585
R3993 gnd.n4636 gnd.n1517 585
R3994 gnd.n2108 gnd.n1517 585
R3995 gnd.n4637 gnd.n1516 585
R3996 gnd.n3402 gnd.n1516 585
R3997 gnd.n4638 gnd.n1515 585
R3998 gnd.n2113 gnd.n1515 585
R3999 gnd.n3398 gnd.n1513 585
R4000 gnd.n3399 gnd.n3398 585
R4001 gnd.n4642 gnd.n1512 585
R4002 gnd.n3390 gnd.n1512 585
R4003 gnd.n4643 gnd.n1511 585
R4004 gnd.n3377 gnd.n1511 585
R4005 gnd.n4644 gnd.n1510 585
R4006 gnd.n2145 gnd.n1510 585
R4007 gnd.n3308 gnd.n1508 585
R4008 gnd.n3309 gnd.n3308 585
R4009 gnd.n4648 gnd.n1507 585
R4010 gnd.n2150 gnd.n1507 585
R4011 gnd.n4649 gnd.n1506 585
R4012 gnd.n3350 gnd.n1506 585
R4013 gnd.n4650 gnd.n1505 585
R4014 gnd.n3342 gnd.n1505 585
R4015 gnd.n3328 gnd.n1503 585
R4016 gnd.n3329 gnd.n3328 585
R4017 gnd.n4654 gnd.n1502 585
R4018 gnd.n3279 gnd.n1502 585
R4019 gnd.n4655 gnd.n1501 585
R4020 gnd.n3300 gnd.n1501 585
R4021 gnd.n4656 gnd.n1500 585
R4022 gnd.n2185 gnd.n1500 585
R4023 gnd.n1497 gnd.n1495 585
R4024 gnd.n2183 gnd.n1495 585
R4025 gnd.n4661 gnd.n4660 585
R4026 gnd.n4662 gnd.n4661 585
R4027 gnd.n1496 gnd.n1494 585
R4028 gnd.n3256 gnd.n1494 585
R4029 gnd.n2264 gnd.n2262 585
R4030 gnd.n2262 gnd.n1464 585
R4031 gnd.n3243 gnd.n3242 585
R4032 gnd.n3244 gnd.n3243 585
R4033 gnd.n2263 gnd.n2261 585
R4034 gnd.n2270 gnd.n2261 585
R4035 gnd.n3237 gnd.n3236 585
R4036 gnd.n3236 gnd.n3235 585
R4037 gnd.n2267 gnd.n2266 585
R4038 gnd.n3213 gnd.n2267 585
R4039 gnd.n2289 gnd.n2287 585
R4040 gnd.n2287 gnd.n2277 585
R4041 gnd.n3203 gnd.n3202 585
R4042 gnd.n3204 gnd.n3203 585
R4043 gnd.n2288 gnd.n2286 585
R4044 gnd.n2295 gnd.n2286 585
R4045 gnd.n3197 gnd.n3196 585
R4046 gnd.n3196 gnd.n3195 585
R4047 gnd.n2292 gnd.n2291 585
R4048 gnd.n3183 gnd.n2292 585
R4049 gnd.n2314 gnd.n2312 585
R4050 gnd.n2312 gnd.n2311 585
R4051 gnd.n3173 gnd.n3172 585
R4052 gnd.n3174 gnd.n3173 585
R4053 gnd.n2313 gnd.n2310 585
R4054 gnd.n2320 gnd.n2310 585
R4055 gnd.n3167 gnd.n3166 585
R4056 gnd.n3166 gnd.n3165 585
R4057 gnd.n2317 gnd.n2316 585
R4058 gnd.n3153 gnd.n2317 585
R4059 gnd.n2337 gnd.n2336 585
R4060 gnd.n2336 gnd.n2327 585
R4061 gnd.n3143 gnd.n3142 585
R4062 gnd.n3144 gnd.n3143 585
R4063 gnd.n3138 gnd.n2335 585
R4064 gnd.n3137 gnd.n2339 585
R4065 gnd.n3136 gnd.n2340 585
R4066 gnd.n3070 gnd.n2340 585
R4067 gnd.n2531 gnd.n2341 585
R4068 gnd.n3132 gnd.n2343 585
R4069 gnd.n3131 gnd.n2344 585
R4070 gnd.n3130 gnd.n2345 585
R4071 gnd.n2534 gnd.n2346 585
R4072 gnd.n3125 gnd.n2461 585
R4073 gnd.n3124 gnd.n2462 585
R4074 gnd.n2536 gnd.n2463 585
R4075 gnd.n3117 gnd.n2471 585
R4076 gnd.n3116 gnd.n2472 585
R4077 gnd.n2539 gnd.n2473 585
R4078 gnd.n3109 gnd.n2481 585
R4079 gnd.n3108 gnd.n2482 585
R4080 gnd.n2541 gnd.n2483 585
R4081 gnd.n3101 gnd.n2492 585
R4082 gnd.n3100 gnd.n2493 585
R4083 gnd.n2544 gnd.n2494 585
R4084 gnd.n3093 gnd.n2502 585
R4085 gnd.n3092 gnd.n2503 585
R4086 gnd.n2546 gnd.n2504 585
R4087 gnd.n3085 gnd.n2513 585
R4088 gnd.n3084 gnd.n2514 585
R4089 gnd.n2550 gnd.n2549 585
R4090 gnd.n2529 gnd.n2528 585
R4091 gnd.n3074 gnd.n3072 585
R4092 gnd.n3073 gnd.n2332 585
R4093 gnd.n1939 gnd.n1580 585
R4094 gnd.n4562 gnd.n1580 585
R4095 gnd.n3934 gnd.n3933 585
R4096 gnd.n3935 gnd.n3934 585
R4097 gnd.n1938 gnd.n1937 585
R4098 gnd.n3942 gnd.n1937 585
R4099 gnd.n3750 gnd.n1936 585
R4100 gnd.n3945 gnd.n1936 585
R4101 gnd.n3749 gnd.n3748 585
R4102 gnd.n3748 gnd.n1935 585
R4103 gnd.n3747 gnd.n3746 585
R4104 gnd.n3747 gnd.n1926 585
R4105 gnd.n1941 gnd.n1925 585
R4106 gnd.n3953 gnd.n1925 585
R4107 gnd.n3742 gnd.n1924 585
R4108 gnd.n3956 gnd.n1924 585
R4109 gnd.n3741 gnd.n3740 585
R4110 gnd.n3740 gnd.n1923 585
R4111 gnd.n3739 gnd.n3738 585
R4112 gnd.n3739 gnd.n1914 585
R4113 gnd.n1943 gnd.n1913 585
R4114 gnd.n3964 gnd.n1913 585
R4115 gnd.n3734 gnd.n1912 585
R4116 gnd.n3967 gnd.n1912 585
R4117 gnd.n3733 gnd.n3732 585
R4118 gnd.n3732 gnd.n1911 585
R4119 gnd.n3731 gnd.n3730 585
R4120 gnd.n3731 gnd.n1902 585
R4121 gnd.n1945 gnd.n1901 585
R4122 gnd.n3975 gnd.n1901 585
R4123 gnd.n3726 gnd.n1900 585
R4124 gnd.n3978 gnd.n1900 585
R4125 gnd.n3725 gnd.n3724 585
R4126 gnd.n3724 gnd.n1846 585
R4127 gnd.n3723 gnd.n3722 585
R4128 gnd.n3723 gnd.n1883 585
R4129 gnd.n1947 gnd.n1891 585
R4130 gnd.n3987 gnd.n1891 585
R4131 gnd.n3718 gnd.n3717 585
R4132 gnd.n3717 gnd.n3716 585
R4133 gnd.n1950 gnd.n1949 585
R4134 gnd.n1957 gnd.n1950 585
R4135 gnd.n3667 gnd.n3666 585
R4136 gnd.n3666 gnd.n1965 585
R4137 gnd.n3668 gnd.n3665 585
R4138 gnd.n3665 gnd.n1962 585
R4139 gnd.n1982 gnd.n1973 585
R4140 gnd.n3683 gnd.n1973 585
R4141 gnd.n3673 gnd.n3672 585
R4142 gnd.n3674 gnd.n3673 585
R4143 gnd.n1981 gnd.n1980 585
R4144 gnd.n3589 gnd.n1980 585
R4145 gnd.n3661 gnd.n3660 585
R4146 gnd.n3660 gnd.n3659 585
R4147 gnd.n1985 gnd.n1984 585
R4148 gnd.n3651 gnd.n1985 585
R4149 gnd.n2011 gnd.n2009 585
R4150 gnd.n2009 gnd.n2001 585
R4151 gnd.n3628 gnd.n3627 585
R4152 gnd.n3629 gnd.n3628 585
R4153 gnd.n2010 gnd.n2008 585
R4154 gnd.n2008 gnd.n2005 585
R4155 gnd.n3622 gnd.n3621 585
R4156 gnd.n3621 gnd.n3620 585
R4157 gnd.n2014 gnd.n2013 585
R4158 gnd.n2023 gnd.n2014 585
R4159 gnd.n3502 gnd.n3500 585
R4160 gnd.n3500 gnd.n3499 585
R4161 gnd.n3503 gnd.n3497 585
R4162 gnd.n3497 gnd.n2028 585
R4163 gnd.n3504 gnd.n2036 585
R4164 gnd.n3561 gnd.n2036 585
R4165 gnd.n3495 gnd.n2043 585
R4166 gnd.n3549 gnd.n2043 585
R4167 gnd.n3508 gnd.n3494 585
R4168 gnd.n3494 gnd.n2048 585
R4169 gnd.n3509 gnd.n3493 585
R4170 gnd.n3493 gnd.n2055 585
R4171 gnd.n3510 gnd.n3492 585
R4172 gnd.n3492 gnd.n3491 585
R4173 gnd.n2072 gnd.n2062 585
R4174 gnd.n3524 gnd.n2062 585
R4175 gnd.n3515 gnd.n3514 585
R4176 gnd.n3516 gnd.n3515 585
R4177 gnd.n2071 gnd.n2070 585
R4178 gnd.n3478 gnd.n2070 585
R4179 gnd.n3452 gnd.n3451 585
R4180 gnd.n3451 gnd.n3450 585
R4181 gnd.n2095 gnd.n2093 585
R4182 gnd.n2093 gnd.n2085 585
R4183 gnd.n3457 gnd.n3456 585
R4184 gnd.n3458 gnd.n3457 585
R4185 gnd.n2094 gnd.n2092 585
R4186 gnd.n3438 gnd.n2092 585
R4187 gnd.n3409 gnd.n3408 585
R4188 gnd.n3411 gnd.n3409 585
R4189 gnd.n2119 gnd.n2118 585
R4190 gnd.n2118 gnd.n2108 585
R4191 gnd.n3404 gnd.n3403 585
R4192 gnd.n3403 gnd.n3402 585
R4193 gnd.n3401 gnd.n2121 585
R4194 gnd.n3401 gnd.n2113 585
R4195 gnd.n3400 gnd.n2123 585
R4196 gnd.n3400 gnd.n3399 585
R4197 gnd.n3315 gnd.n2122 585
R4198 gnd.n3390 gnd.n2122 585
R4199 gnd.n3316 gnd.n2140 585
R4200 gnd.n3377 gnd.n2140 585
R4201 gnd.n3312 gnd.n3311 585
R4202 gnd.n3311 gnd.n2145 585
R4203 gnd.n3320 gnd.n3310 585
R4204 gnd.n3310 gnd.n3309 585
R4205 gnd.n3321 gnd.n3306 585
R4206 gnd.n3306 gnd.n2150 585
R4207 gnd.n3322 gnd.n2157 585
R4208 gnd.n3350 gnd.n2157 585
R4209 gnd.n2171 gnd.n2165 585
R4210 gnd.n3342 gnd.n2165 585
R4211 gnd.n3327 gnd.n3326 585
R4212 gnd.n3329 gnd.n3327 585
R4213 gnd.n2170 gnd.n2169 585
R4214 gnd.n3279 gnd.n2169 585
R4215 gnd.n3302 gnd.n3301 585
R4216 gnd.n3301 gnd.n3300 585
R4217 gnd.n2174 gnd.n2173 585
R4218 gnd.n2185 gnd.n2174 585
R4219 gnd.n3250 gnd.n3249 585
R4220 gnd.n3249 gnd.n2183 585
R4221 gnd.n2255 gnd.n1492 585
R4222 gnd.n4662 gnd.n1492 585
R4223 gnd.n3255 gnd.n3254 585
R4224 gnd.n3256 gnd.n3255 585
R4225 gnd.n2254 gnd.n2253 585
R4226 gnd.n2253 gnd.n1464 585
R4227 gnd.n3246 gnd.n3245 585
R4228 gnd.n3245 gnd.n3244 585
R4229 gnd.n2258 gnd.n2257 585
R4230 gnd.n2270 gnd.n2258 585
R4231 gnd.n2280 gnd.n2269 585
R4232 gnd.n3235 gnd.n2269 585
R4233 gnd.n3212 gnd.n3211 585
R4234 gnd.n3213 gnd.n3212 585
R4235 gnd.n2279 gnd.n2278 585
R4236 gnd.n2278 gnd.n2277 585
R4237 gnd.n3206 gnd.n3205 585
R4238 gnd.n3205 gnd.n3204 585
R4239 gnd.n2283 gnd.n2282 585
R4240 gnd.n2295 gnd.n2283 585
R4241 gnd.n2304 gnd.n2294 585
R4242 gnd.n3195 gnd.n2294 585
R4243 gnd.n3182 gnd.n3181 585
R4244 gnd.n3183 gnd.n3182 585
R4245 gnd.n2303 gnd.n2302 585
R4246 gnd.n2311 gnd.n2302 585
R4247 gnd.n3176 gnd.n3175 585
R4248 gnd.n3175 gnd.n3174 585
R4249 gnd.n2307 gnd.n2306 585
R4250 gnd.n2320 gnd.n2307 585
R4251 gnd.n2330 gnd.n2319 585
R4252 gnd.n3165 gnd.n2319 585
R4253 gnd.n3152 gnd.n3151 585
R4254 gnd.n3153 gnd.n3152 585
R4255 gnd.n2329 gnd.n2328 585
R4256 gnd.n2328 gnd.n2327 585
R4257 gnd.n3146 gnd.n3145 585
R4258 gnd.n3145 gnd.n3144 585
R4259 gnd.n3908 gnd.n3762 585
R4260 gnd.n3762 gnd.n1590 585
R4261 gnd.n3909 gnd.n3906 585
R4262 gnd.n3904 gnd.n3780 585
R4263 gnd.n3903 gnd.n3902 585
R4264 gnd.n3887 gnd.n3782 585
R4265 gnd.n3889 gnd.n3888 585
R4266 gnd.n3885 gnd.n3789 585
R4267 gnd.n3884 gnd.n3883 585
R4268 gnd.n3868 gnd.n3791 585
R4269 gnd.n3870 gnd.n3869 585
R4270 gnd.n3866 gnd.n3798 585
R4271 gnd.n3865 gnd.n3864 585
R4272 gnd.n3849 gnd.n3800 585
R4273 gnd.n3851 gnd.n3850 585
R4274 gnd.n3847 gnd.n3807 585
R4275 gnd.n3846 gnd.n3845 585
R4276 gnd.n3834 gnd.n3809 585
R4277 gnd.n3836 gnd.n3835 585
R4278 gnd.n3832 gnd.n3810 585
R4279 gnd.n3831 gnd.n3830 585
R4280 gnd.n3823 gnd.n3812 585
R4281 gnd.n3825 gnd.n3824 585
R4282 gnd.n3821 gnd.n3814 585
R4283 gnd.n3820 gnd.n3819 585
R4284 gnd.n3816 gnd.n1578 585
R4285 gnd.n3929 gnd.n3928 585
R4286 gnd.n3926 gnd.n3760 585
R4287 gnd.n3925 gnd.n3761 585
R4288 gnd.n3923 gnd.n3922 585
R4289 gnd.n4077 gnd.n1886 463.671
R4290 gnd.n4080 gnd.n4079 463.671
R4291 gnd.n3258 gnd.n2252 463.671
R4292 gnd.n4731 gnd.n1467 463.671
R4293 gnd.n2188 gnd.t106 443.966
R4294 gnd.n1879 gnd.t130 443.966
R4295 gnd.n4668 gnd.t160 443.966
R4296 gnd.n4011 gnd.t182 443.966
R4297 gnd.n6632 gnd.n6631 434.747
R4298 gnd.n2515 gnd.t140 371.625
R4299 gnd.n3773 gnd.t166 371.625
R4300 gnd.n2522 gnd.t191 371.625
R4301 gnd.n4217 gnd.t163 371.625
R4302 gnd.n4269 gnd.t154 371.625
R4303 gnd.n1810 gnd.t88 371.625
R4304 gnd.n313 gnd.t188 371.625
R4305 gnd.n280 gnd.t102 371.625
R4306 gnd.n7520 gnd.t144 371.625
R4307 gnd.n350 gnd.t134 371.625
R4308 gnd.n1090 gnd.t117 371.625
R4309 gnd.n1112 gnd.t114 371.625
R4310 gnd.n1134 gnd.t92 371.625
R4311 gnd.n2687 gnd.t172 371.625
R4312 gnd.n1409 gnd.t175 371.625
R4313 gnd.n2348 gnd.t110 371.625
R4314 gnd.n2370 gnd.t137 371.625
R4315 gnd.n3763 gnd.t123 371.625
R4316 gnd.n5643 gnd.t150 323.425
R4317 gnd.n5077 gnd.t178 323.425
R4318 gnd.n6288 gnd.n6262 289.615
R4319 gnd.n6256 gnd.n6230 289.615
R4320 gnd.n6224 gnd.n6198 289.615
R4321 gnd.n6193 gnd.n6167 289.615
R4322 gnd.n6161 gnd.n6135 289.615
R4323 gnd.n6129 gnd.n6103 289.615
R4324 gnd.n6097 gnd.n6071 289.615
R4325 gnd.n6066 gnd.n6040 289.615
R4326 gnd.n5493 gnd.t84 279.217
R4327 gnd.n5121 gnd.t80 279.217
R4328 gnd.n1474 gnd.t122 260.649
R4329 gnd.n4003 gnd.t101 260.649
R4330 gnd.n4733 gnd.n4732 256.663
R4331 gnd.n4733 gnd.n1433 256.663
R4332 gnd.n4733 gnd.n1434 256.663
R4333 gnd.n4733 gnd.n1435 256.663
R4334 gnd.n4733 gnd.n1436 256.663
R4335 gnd.n4733 gnd.n1437 256.663
R4336 gnd.n4733 gnd.n1438 256.663
R4337 gnd.n4733 gnd.n1439 256.663
R4338 gnd.n4733 gnd.n1440 256.663
R4339 gnd.n4733 gnd.n1441 256.663
R4340 gnd.n4733 gnd.n1442 256.663
R4341 gnd.n4733 gnd.n1443 256.663
R4342 gnd.n4733 gnd.n1444 256.663
R4343 gnd.n4733 gnd.n1445 256.663
R4344 gnd.n4733 gnd.n1446 256.663
R4345 gnd.n4733 gnd.n1447 256.663
R4346 gnd.n4736 gnd.n1431 256.663
R4347 gnd.n4734 gnd.n4733 256.663
R4348 gnd.n4733 gnd.n1448 256.663
R4349 gnd.n4733 gnd.n1449 256.663
R4350 gnd.n4733 gnd.n1450 256.663
R4351 gnd.n4733 gnd.n1451 256.663
R4352 gnd.n4733 gnd.n1452 256.663
R4353 gnd.n4733 gnd.n1453 256.663
R4354 gnd.n4733 gnd.n1454 256.663
R4355 gnd.n4733 gnd.n1455 256.663
R4356 gnd.n4733 gnd.n1456 256.663
R4357 gnd.n4733 gnd.n1457 256.663
R4358 gnd.n4733 gnd.n1458 256.663
R4359 gnd.n4733 gnd.n1459 256.663
R4360 gnd.n4733 gnd.n1460 256.663
R4361 gnd.n4733 gnd.n1461 256.663
R4362 gnd.n4733 gnd.n1462 256.663
R4363 gnd.n4733 gnd.n1463 256.663
R4364 gnd.n4145 gnd.n1863 256.663
R4365 gnd.n4145 gnd.n1864 256.663
R4366 gnd.n4145 gnd.n1865 256.663
R4367 gnd.n4145 gnd.n1866 256.663
R4368 gnd.n4145 gnd.n1867 256.663
R4369 gnd.n4145 gnd.n1868 256.663
R4370 gnd.n4145 gnd.n1869 256.663
R4371 gnd.n4145 gnd.n1870 256.663
R4372 gnd.n4145 gnd.n1871 256.663
R4373 gnd.n4145 gnd.n1872 256.663
R4374 gnd.n4145 gnd.n1873 256.663
R4375 gnd.n4145 gnd.n1874 256.663
R4376 gnd.n4145 gnd.n1875 256.663
R4377 gnd.n4145 gnd.n1876 256.663
R4378 gnd.n4145 gnd.n1877 256.663
R4379 gnd.n4145 gnd.n4142 256.663
R4380 gnd.n4148 gnd.n1844 256.663
R4381 gnd.n4146 gnd.n4145 256.663
R4382 gnd.n4145 gnd.n1862 256.663
R4383 gnd.n4145 gnd.n1861 256.663
R4384 gnd.n4145 gnd.n1860 256.663
R4385 gnd.n4145 gnd.n1859 256.663
R4386 gnd.n4145 gnd.n1858 256.663
R4387 gnd.n4145 gnd.n1857 256.663
R4388 gnd.n4145 gnd.n1856 256.663
R4389 gnd.n4145 gnd.n1855 256.663
R4390 gnd.n4145 gnd.n1854 256.663
R4391 gnd.n4145 gnd.n1853 256.663
R4392 gnd.n4145 gnd.n1852 256.663
R4393 gnd.n4145 gnd.n1851 256.663
R4394 gnd.n4145 gnd.n1850 256.663
R4395 gnd.n4145 gnd.n1849 256.663
R4396 gnd.n4145 gnd.n1848 256.663
R4397 gnd.n4145 gnd.n1847 256.663
R4398 gnd.n5046 gnd.n1058 242.672
R4399 gnd.n5046 gnd.n1059 242.672
R4400 gnd.n5046 gnd.n1060 242.672
R4401 gnd.n5046 gnd.n1061 242.672
R4402 gnd.n5046 gnd.n1062 242.672
R4403 gnd.n5046 gnd.n1063 242.672
R4404 gnd.n5046 gnd.n1064 242.672
R4405 gnd.n5046 gnd.n1065 242.672
R4406 gnd.n5046 gnd.n1066 242.672
R4407 gnd.n3077 gnd.n1381 242.672
R4408 gnd.n2520 gnd.n1381 242.672
R4409 gnd.n2509 gnd.n1381 242.672
R4410 gnd.n2506 gnd.n1381 242.672
R4411 gnd.n2497 gnd.n1381 242.672
R4412 gnd.n2488 gnd.n1381 242.672
R4413 gnd.n2485 gnd.n1381 242.672
R4414 gnd.n2476 gnd.n1381 242.672
R4415 gnd.n2467 gnd.n1381 242.672
R4416 gnd.n5548 gnd.n5457 242.672
R4417 gnd.n5461 gnd.n5457 242.672
R4418 gnd.n5541 gnd.n5457 242.672
R4419 gnd.n5535 gnd.n5457 242.672
R4420 gnd.n5533 gnd.n5457 242.672
R4421 gnd.n5527 gnd.n5457 242.672
R4422 gnd.n5525 gnd.n5457 242.672
R4423 gnd.n5519 gnd.n5457 242.672
R4424 gnd.n5517 gnd.n5457 242.672
R4425 gnd.n5511 gnd.n5457 242.672
R4426 gnd.n5509 gnd.n5457 242.672
R4427 gnd.n5502 gnd.n5457 242.672
R4428 gnd.n5500 gnd.n5457 242.672
R4429 gnd.n6344 gnd.n5047 242.672
R4430 gnd.n6350 gnd.n5047 242.672
R4431 gnd.n5124 gnd.n5047 242.672
R4432 gnd.n6357 gnd.n5047 242.672
R4433 gnd.n5115 gnd.n5047 242.672
R4434 gnd.n6364 gnd.n5047 242.672
R4435 gnd.n5108 gnd.n5047 242.672
R4436 gnd.n6371 gnd.n5047 242.672
R4437 gnd.n5101 gnd.n5047 242.672
R4438 gnd.n6378 gnd.n5047 242.672
R4439 gnd.n5094 gnd.n5047 242.672
R4440 gnd.n6385 gnd.n5047 242.672
R4441 gnd.n5087 gnd.n5047 242.672
R4442 gnd.n3839 gnd.n1591 242.672
R4443 gnd.n3856 gnd.n1591 242.672
R4444 gnd.n3858 gnd.n1591 242.672
R4445 gnd.n3875 gnd.n1591 242.672
R4446 gnd.n3877 gnd.n1591 242.672
R4447 gnd.n3894 gnd.n1591 242.672
R4448 gnd.n3896 gnd.n1591 242.672
R4449 gnd.n3914 gnd.n1591 242.672
R4450 gnd.n3916 gnd.n1591 242.672
R4451 gnd.n347 gnd.n212 242.672
R4452 gnd.n7416 gnd.n212 242.672
R4453 gnd.n343 gnd.n212 242.672
R4454 gnd.n7423 gnd.n212 242.672
R4455 gnd.n336 gnd.n212 242.672
R4456 gnd.n7430 gnd.n212 242.672
R4457 gnd.n329 gnd.n212 242.672
R4458 gnd.n7437 gnd.n212 242.672
R4459 gnd.n322 gnd.n212 242.672
R4460 gnd.n5677 gnd.n5676 242.672
R4461 gnd.n5677 gnd.n5618 242.672
R4462 gnd.n5677 gnd.n5619 242.672
R4463 gnd.n5677 gnd.n5620 242.672
R4464 gnd.n5677 gnd.n5621 242.672
R4465 gnd.n5677 gnd.n5622 242.672
R4466 gnd.n5677 gnd.n5623 242.672
R4467 gnd.n5677 gnd.n5624 242.672
R4468 gnd.n6396 gnd.n5047 242.672
R4469 gnd.n5080 gnd.n5047 242.672
R4470 gnd.n6403 gnd.n5047 242.672
R4471 gnd.n5071 gnd.n5047 242.672
R4472 gnd.n6410 gnd.n5047 242.672
R4473 gnd.n5064 gnd.n5047 242.672
R4474 gnd.n6417 gnd.n5047 242.672
R4475 gnd.n5057 gnd.n5047 242.672
R4476 gnd.n5046 gnd.n5045 242.672
R4477 gnd.n5046 gnd.n1030 242.672
R4478 gnd.n5046 gnd.n1031 242.672
R4479 gnd.n5046 gnd.n1032 242.672
R4480 gnd.n5046 gnd.n1033 242.672
R4481 gnd.n5046 gnd.n1034 242.672
R4482 gnd.n5046 gnd.n1035 242.672
R4483 gnd.n5046 gnd.n1036 242.672
R4484 gnd.n5046 gnd.n1037 242.672
R4485 gnd.n5046 gnd.n1038 242.672
R4486 gnd.n5046 gnd.n1039 242.672
R4487 gnd.n5046 gnd.n1040 242.672
R4488 gnd.n5046 gnd.n1041 242.672
R4489 gnd.n5046 gnd.n1042 242.672
R4490 gnd.n5046 gnd.n1043 242.672
R4491 gnd.n5046 gnd.n1044 242.672
R4492 gnd.n5046 gnd.n1045 242.672
R4493 gnd.n5046 gnd.n1046 242.672
R4494 gnd.n5046 gnd.n1047 242.672
R4495 gnd.n5046 gnd.n1048 242.672
R4496 gnd.n5046 gnd.n1049 242.672
R4497 gnd.n5046 gnd.n1050 242.672
R4498 gnd.n5046 gnd.n1051 242.672
R4499 gnd.n5046 gnd.n1052 242.672
R4500 gnd.n5046 gnd.n1053 242.672
R4501 gnd.n5046 gnd.n1054 242.672
R4502 gnd.n5046 gnd.n1055 242.672
R4503 gnd.n5046 gnd.n1056 242.672
R4504 gnd.n5046 gnd.n1057 242.672
R4505 gnd.n2455 gnd.n1381 242.672
R4506 gnd.n2351 gnd.n1381 242.672
R4507 gnd.n2445 gnd.n1381 242.672
R4508 gnd.n2355 gnd.n1381 242.672
R4509 gnd.n2435 gnd.n1381 242.672
R4510 gnd.n2359 gnd.n1381 242.672
R4511 gnd.n2425 gnd.n1381 242.672
R4512 gnd.n2363 gnd.n1381 242.672
R4513 gnd.n2415 gnd.n1381 242.672
R4514 gnd.n2367 gnd.n1381 242.672
R4515 gnd.n2405 gnd.n1381 242.672
R4516 gnd.n2373 gnd.n1381 242.672
R4517 gnd.n2395 gnd.n1381 242.672
R4518 gnd.n2377 gnd.n1381 242.672
R4519 gnd.n2385 gnd.n1381 242.672
R4520 gnd.n2382 gnd.n1381 242.672
R4521 gnd.n4737 gnd.n1427 242.672
R4522 gnd.n1426 gnd.n1381 242.672
R4523 gnd.n4741 gnd.n1381 242.672
R4524 gnd.n1420 gnd.n1381 242.672
R4525 gnd.n4748 gnd.n1381 242.672
R4526 gnd.n1413 gnd.n1381 242.672
R4527 gnd.n4756 gnd.n1381 242.672
R4528 gnd.n1404 gnd.n1381 242.672
R4529 gnd.n4763 gnd.n1381 242.672
R4530 gnd.n1397 gnd.n1381 242.672
R4531 gnd.n4770 gnd.n1381 242.672
R4532 gnd.n1390 gnd.n1381 242.672
R4533 gnd.n4777 gnd.n1381 242.672
R4534 gnd.n4780 gnd.n1381 242.672
R4535 gnd.n4178 gnd.n1591 242.672
R4536 gnd.n4181 gnd.n1591 242.672
R4537 gnd.n4189 gnd.n1591 242.672
R4538 gnd.n4191 gnd.n1591 242.672
R4539 gnd.n4199 gnd.n1591 242.672
R4540 gnd.n4201 gnd.n1591 242.672
R4541 gnd.n4209 gnd.n1591 242.672
R4542 gnd.n4211 gnd.n1591 242.672
R4543 gnd.n4222 gnd.n1591 242.672
R4544 gnd.n4224 gnd.n1591 242.672
R4545 gnd.n4232 gnd.n1591 242.672
R4546 gnd.n4234 gnd.n1591 242.672
R4547 gnd.n4243 gnd.n1591 242.672
R4548 gnd.n4244 gnd.n4149 242.672
R4549 gnd.n4245 gnd.n1591 242.672
R4550 gnd.n4247 gnd.n1591 242.672
R4551 gnd.n4255 gnd.n1591 242.672
R4552 gnd.n4257 gnd.n1591 242.672
R4553 gnd.n4265 gnd.n1591 242.672
R4554 gnd.n4267 gnd.n1591 242.672
R4555 gnd.n4277 gnd.n1591 242.672
R4556 gnd.n4279 gnd.n1591 242.672
R4557 gnd.n4287 gnd.n1591 242.672
R4558 gnd.n4289 gnd.n1591 242.672
R4559 gnd.n4297 gnd.n1591 242.672
R4560 gnd.n4299 gnd.n1591 242.672
R4561 gnd.n4307 gnd.n1591 242.672
R4562 gnd.n4309 gnd.n1591 242.672
R4563 gnd.n4318 gnd.n1591 242.672
R4564 gnd.n4321 gnd.n1591 242.672
R4565 gnd.n7448 gnd.n212 242.672
R4566 gnd.n316 gnd.n212 242.672
R4567 gnd.n7455 gnd.n212 242.672
R4568 gnd.n307 gnd.n212 242.672
R4569 gnd.n7462 gnd.n212 242.672
R4570 gnd.n300 gnd.n212 242.672
R4571 gnd.n7469 gnd.n212 242.672
R4572 gnd.n293 gnd.n212 242.672
R4573 gnd.n7476 gnd.n212 242.672
R4574 gnd.n7479 gnd.n212 242.672
R4575 gnd.n284 gnd.n212 242.672
R4576 gnd.n7488 gnd.n212 242.672
R4577 gnd.n275 gnd.n212 242.672
R4578 gnd.n7495 gnd.n212 242.672
R4579 gnd.n268 gnd.n212 242.672
R4580 gnd.n7502 gnd.n212 242.672
R4581 gnd.n261 gnd.n212 242.672
R4582 gnd.n7509 gnd.n212 242.672
R4583 gnd.n254 gnd.n212 242.672
R4584 gnd.n7516 gnd.n212 242.672
R4585 gnd.n247 gnd.n212 242.672
R4586 gnd.n7526 gnd.n212 242.672
R4587 gnd.n240 gnd.n212 242.672
R4588 gnd.n7533 gnd.n212 242.672
R4589 gnd.n233 gnd.n212 242.672
R4590 gnd.n7540 gnd.n212 242.672
R4591 gnd.n226 gnd.n212 242.672
R4592 gnd.n7547 gnd.n212 242.672
R4593 gnd.n219 gnd.n212 242.672
R4594 gnd.n3070 gnd.n3069 242.672
R4595 gnd.n3070 gnd.n2532 242.672
R4596 gnd.n3070 gnd.n2533 242.672
R4597 gnd.n3070 gnd.n2535 242.672
R4598 gnd.n3070 gnd.n2537 242.672
R4599 gnd.n3070 gnd.n2538 242.672
R4600 gnd.n3070 gnd.n2540 242.672
R4601 gnd.n3070 gnd.n2542 242.672
R4602 gnd.n3070 gnd.n2543 242.672
R4603 gnd.n3070 gnd.n2545 242.672
R4604 gnd.n3070 gnd.n2547 242.672
R4605 gnd.n3070 gnd.n2548 242.672
R4606 gnd.n3070 gnd.n2551 242.672
R4607 gnd.n3071 gnd.n3070 242.672
R4608 gnd.n3905 gnd.n1590 242.672
R4609 gnd.n3781 gnd.n1590 242.672
R4610 gnd.n3886 gnd.n1590 242.672
R4611 gnd.n3790 gnd.n1590 242.672
R4612 gnd.n3867 gnd.n1590 242.672
R4613 gnd.n3799 gnd.n1590 242.672
R4614 gnd.n3848 gnd.n1590 242.672
R4615 gnd.n3808 gnd.n1590 242.672
R4616 gnd.n3833 gnd.n1590 242.672
R4617 gnd.n3811 gnd.n1590 242.672
R4618 gnd.n3822 gnd.n1590 242.672
R4619 gnd.n3815 gnd.n1590 242.672
R4620 gnd.n3927 gnd.n1590 242.672
R4621 gnd.n3924 gnd.n1590 242.672
R4622 gnd.n216 gnd.n213 240.244
R4623 gnd.n7549 gnd.n7548 240.244
R4624 gnd.n7546 gnd.n220 240.244
R4625 gnd.n7542 gnd.n7541 240.244
R4626 gnd.n7539 gnd.n227 240.244
R4627 gnd.n7535 gnd.n7534 240.244
R4628 gnd.n7532 gnd.n234 240.244
R4629 gnd.n7528 gnd.n7527 240.244
R4630 gnd.n7525 gnd.n241 240.244
R4631 gnd.n7518 gnd.n7517 240.244
R4632 gnd.n7515 gnd.n248 240.244
R4633 gnd.n7511 gnd.n7510 240.244
R4634 gnd.n7508 gnd.n255 240.244
R4635 gnd.n7504 gnd.n7503 240.244
R4636 gnd.n7501 gnd.n262 240.244
R4637 gnd.n7497 gnd.n7496 240.244
R4638 gnd.n7494 gnd.n269 240.244
R4639 gnd.n7490 gnd.n7489 240.244
R4640 gnd.n7487 gnd.n276 240.244
R4641 gnd.n7480 gnd.n285 240.244
R4642 gnd.n7478 gnd.n7477 240.244
R4643 gnd.n7475 gnd.n287 240.244
R4644 gnd.n7471 gnd.n7470 240.244
R4645 gnd.n7468 gnd.n294 240.244
R4646 gnd.n7464 gnd.n7463 240.244
R4647 gnd.n7461 gnd.n301 240.244
R4648 gnd.n7457 gnd.n7456 240.244
R4649 gnd.n7454 gnd.n308 240.244
R4650 gnd.n7450 gnd.n7449 240.244
R4651 gnd.n1807 gnd.n1600 240.244
R4652 gnd.n1807 gnd.n1612 240.244
R4653 gnd.n4332 gnd.n1612 240.244
R4654 gnd.n4332 gnd.n1624 240.244
R4655 gnd.n4342 gnd.n1624 240.244
R4656 gnd.n4342 gnd.n1635 240.244
R4657 gnd.n4346 gnd.n1635 240.244
R4658 gnd.n4346 gnd.n1644 240.244
R4659 gnd.n4356 gnd.n1644 240.244
R4660 gnd.n4356 gnd.n1655 240.244
R4661 gnd.n1755 gnd.n1655 240.244
R4662 gnd.n1755 gnd.n1664 240.244
R4663 gnd.n4363 gnd.n1664 240.244
R4664 gnd.n4363 gnd.n1675 240.244
R4665 gnd.n4368 gnd.n1675 240.244
R4666 gnd.n4368 gnd.n1684 240.244
R4667 gnd.n4373 gnd.n1684 240.244
R4668 gnd.n4373 gnd.n1695 240.244
R4669 gnd.n4416 gnd.n1695 240.244
R4670 gnd.n4416 gnd.n1704 240.244
R4671 gnd.n4444 gnd.n1704 240.244
R4672 gnd.n4444 gnd.n1713 240.244
R4673 gnd.n1737 gnd.n1713 240.244
R4674 gnd.n1737 gnd.n1722 240.244
R4675 gnd.n1729 gnd.n1722 240.244
R4676 gnd.n4437 gnd.n1729 240.244
R4677 gnd.n4437 gnd.n4436 240.244
R4678 gnd.n4436 gnd.n86 240.244
R4679 gnd.n380 gnd.n86 240.244
R4680 gnd.n7329 gnd.n380 240.244
R4681 gnd.n7329 gnd.n103 240.244
R4682 gnd.n7333 gnd.n103 240.244
R4683 gnd.n7333 gnd.n115 240.244
R4684 gnd.n7343 gnd.n115 240.244
R4685 gnd.n7343 gnd.n124 240.244
R4686 gnd.n7347 gnd.n124 240.244
R4687 gnd.n7347 gnd.n133 240.244
R4688 gnd.n7357 gnd.n133 240.244
R4689 gnd.n7357 gnd.n144 240.244
R4690 gnd.n7361 gnd.n144 240.244
R4691 gnd.n7361 gnd.n154 240.244
R4692 gnd.n7372 gnd.n154 240.244
R4693 gnd.n7372 gnd.n164 240.244
R4694 gnd.n7391 gnd.n164 240.244
R4695 gnd.n7391 gnd.n173 240.244
R4696 gnd.n7387 gnd.n173 240.244
R4697 gnd.n7387 gnd.n183 240.244
R4698 gnd.n7384 gnd.n183 240.244
R4699 gnd.n7384 gnd.n192 240.244
R4700 gnd.n7381 gnd.n192 240.244
R4701 gnd.n7381 gnd.n202 240.244
R4702 gnd.n7378 gnd.n202 240.244
R4703 gnd.n7378 gnd.n210 240.244
R4704 gnd.n4180 gnd.n4179 240.244
R4705 gnd.n4182 gnd.n4180 240.244
R4706 gnd.n4188 gnd.n4170 240.244
R4707 gnd.n4192 gnd.n4190 240.244
R4708 gnd.n4198 gnd.n4166 240.244
R4709 gnd.n4202 gnd.n4200 240.244
R4710 gnd.n4208 gnd.n4162 240.244
R4711 gnd.n4212 gnd.n4210 240.244
R4712 gnd.n4221 gnd.n4158 240.244
R4713 gnd.n4225 gnd.n4223 240.244
R4714 gnd.n4231 gnd.n4154 240.244
R4715 gnd.n4235 gnd.n4233 240.244
R4716 gnd.n4242 gnd.n4150 240.244
R4717 gnd.n4248 gnd.n4246 240.244
R4718 gnd.n4254 gnd.n1838 240.244
R4719 gnd.n4258 gnd.n4256 240.244
R4720 gnd.n4264 gnd.n1834 240.244
R4721 gnd.n4268 gnd.n4266 240.244
R4722 gnd.n4276 gnd.n1830 240.244
R4723 gnd.n4280 gnd.n4278 240.244
R4724 gnd.n4286 gnd.n1826 240.244
R4725 gnd.n4290 gnd.n4288 240.244
R4726 gnd.n4296 gnd.n1822 240.244
R4727 gnd.n4300 gnd.n4298 240.244
R4728 gnd.n4306 gnd.n1818 240.244
R4729 gnd.n4310 gnd.n4308 240.244
R4730 gnd.n4317 gnd.n1814 240.244
R4731 gnd.n4320 gnd.n4319 240.244
R4732 gnd.n4545 gnd.n1605 240.244
R4733 gnd.n4541 gnd.n1605 240.244
R4734 gnd.n4541 gnd.n1610 240.244
R4735 gnd.n4533 gnd.n1610 240.244
R4736 gnd.n4533 gnd.n1627 240.244
R4737 gnd.n4529 gnd.n1627 240.244
R4738 gnd.n4529 gnd.n1633 240.244
R4739 gnd.n4521 gnd.n1633 240.244
R4740 gnd.n4521 gnd.n1647 240.244
R4741 gnd.n4517 gnd.n1647 240.244
R4742 gnd.n4517 gnd.n1653 240.244
R4743 gnd.n4509 gnd.n1653 240.244
R4744 gnd.n4509 gnd.n1667 240.244
R4745 gnd.n4505 gnd.n1667 240.244
R4746 gnd.n4505 gnd.n1673 240.244
R4747 gnd.n4497 gnd.n1673 240.244
R4748 gnd.n4497 gnd.n1687 240.244
R4749 gnd.n4493 gnd.n1687 240.244
R4750 gnd.n4493 gnd.n1693 240.244
R4751 gnd.n4485 gnd.n1693 240.244
R4752 gnd.n4485 gnd.n1707 240.244
R4753 gnd.n4481 gnd.n1707 240.244
R4754 gnd.n4481 gnd.n1711 240.244
R4755 gnd.n4473 gnd.n1711 240.244
R4756 gnd.n4473 gnd.n4472 240.244
R4757 gnd.n4472 gnd.n1727 240.244
R4758 gnd.n1727 gnd.n89 240.244
R4759 gnd.n7630 gnd.n89 240.244
R4760 gnd.n7630 gnd.n90 240.244
R4761 gnd.n100 gnd.n90 240.244
R4762 gnd.n7624 gnd.n100 240.244
R4763 gnd.n7624 gnd.n101 240.244
R4764 gnd.n7616 gnd.n101 240.244
R4765 gnd.n7616 gnd.n117 240.244
R4766 gnd.n7612 gnd.n117 240.244
R4767 gnd.n7612 gnd.n122 240.244
R4768 gnd.n7604 gnd.n122 240.244
R4769 gnd.n7604 gnd.n136 240.244
R4770 gnd.n7600 gnd.n136 240.244
R4771 gnd.n7600 gnd.n142 240.244
R4772 gnd.n7592 gnd.n142 240.244
R4773 gnd.n7592 gnd.n156 240.244
R4774 gnd.n7588 gnd.n156 240.244
R4775 gnd.n7588 gnd.n162 240.244
R4776 gnd.n7580 gnd.n162 240.244
R4777 gnd.n7580 gnd.n176 240.244
R4778 gnd.n7576 gnd.n176 240.244
R4779 gnd.n7576 gnd.n182 240.244
R4780 gnd.n7568 gnd.n182 240.244
R4781 gnd.n7568 gnd.n195 240.244
R4782 gnd.n7564 gnd.n195 240.244
R4783 gnd.n7564 gnd.n201 240.244
R4784 gnd.n7556 gnd.n201 240.244
R4785 gnd.n4781 gnd.n1377 240.244
R4786 gnd.n4779 gnd.n4778 240.244
R4787 gnd.n4776 gnd.n1383 240.244
R4788 gnd.n4772 gnd.n4771 240.244
R4789 gnd.n4769 gnd.n1391 240.244
R4790 gnd.n4765 gnd.n4764 240.244
R4791 gnd.n4762 gnd.n1398 240.244
R4792 gnd.n4758 gnd.n4757 240.244
R4793 gnd.n4755 gnd.n1405 240.244
R4794 gnd.n4750 gnd.n4749 240.244
R4795 gnd.n4747 gnd.n1414 240.244
R4796 gnd.n4743 gnd.n4742 240.244
R4797 gnd.n4740 gnd.n1421 240.244
R4798 gnd.n2384 gnd.n2383 240.244
R4799 gnd.n2387 gnd.n2386 240.244
R4800 gnd.n2394 gnd.n2393 240.244
R4801 gnd.n2397 gnd.n2396 240.244
R4802 gnd.n2404 gnd.n2403 240.244
R4803 gnd.n2407 gnd.n2406 240.244
R4804 gnd.n2414 gnd.n2413 240.244
R4805 gnd.n2417 gnd.n2416 240.244
R4806 gnd.n2424 gnd.n2423 240.244
R4807 gnd.n2427 gnd.n2426 240.244
R4808 gnd.n2434 gnd.n2433 240.244
R4809 gnd.n2437 gnd.n2436 240.244
R4810 gnd.n2444 gnd.n2443 240.244
R4811 gnd.n2447 gnd.n2446 240.244
R4812 gnd.n2454 gnd.n2453 240.244
R4813 gnd.n4924 gnd.n4923 240.244
R4814 gnd.n4923 gnd.n1141 240.244
R4815 gnd.n1153 gnd.n1141 240.244
R4816 gnd.n2669 gnd.n1153 240.244
R4817 gnd.n2669 gnd.n1165 240.244
R4818 gnd.n2673 gnd.n1165 240.244
R4819 gnd.n2673 gnd.n1175 240.244
R4820 gnd.n2676 gnd.n1175 240.244
R4821 gnd.n2676 gnd.n1185 240.244
R4822 gnd.n2767 gnd.n1185 240.244
R4823 gnd.n2767 gnd.n1195 240.244
R4824 gnd.n2771 gnd.n1195 240.244
R4825 gnd.n2771 gnd.n1205 240.244
R4826 gnd.n2820 gnd.n1205 240.244
R4827 gnd.n2820 gnd.n1215 240.244
R4828 gnd.n2824 gnd.n1215 240.244
R4829 gnd.n2824 gnd.n1225 240.244
R4830 gnd.n2835 gnd.n1225 240.244
R4831 gnd.n2835 gnd.n1236 240.244
R4832 gnd.n2840 gnd.n1236 240.244
R4833 gnd.n2840 gnd.n1246 240.244
R4834 gnd.n2646 gnd.n1246 240.244
R4835 gnd.n2646 gnd.n2641 240.244
R4836 gnd.n2853 gnd.n2641 240.244
R4837 gnd.n2853 gnd.n2626 240.244
R4838 gnd.n2626 gnd.n2620 240.244
R4839 gnd.n2633 gnd.n2620 240.244
R4840 gnd.n2633 gnd.n2614 240.244
R4841 gnd.n2614 gnd.n2612 240.244
R4842 gnd.n2612 gnd.n2598 240.244
R4843 gnd.n2598 gnd.n1263 240.244
R4844 gnd.n2911 gnd.n1263 240.244
R4845 gnd.n2911 gnd.n1275 240.244
R4846 gnd.n2917 gnd.n1275 240.244
R4847 gnd.n2917 gnd.n1284 240.244
R4848 gnd.n2924 gnd.n1284 240.244
R4849 gnd.n2924 gnd.n1294 240.244
R4850 gnd.n2585 gnd.n1294 240.244
R4851 gnd.n2585 gnd.n1304 240.244
R4852 gnd.n2988 gnd.n1304 240.244
R4853 gnd.n2988 gnd.n1314 240.244
R4854 gnd.n2993 gnd.n1314 240.244
R4855 gnd.n2993 gnd.n1324 240.244
R4856 gnd.n3003 gnd.n1324 240.244
R4857 gnd.n3003 gnd.n1334 240.244
R4858 gnd.n2567 gnd.n1334 240.244
R4859 gnd.n2567 gnd.n1344 240.244
R4860 gnd.n3010 gnd.n1344 240.244
R4861 gnd.n3010 gnd.n1354 240.244
R4862 gnd.n3015 gnd.n1354 240.244
R4863 gnd.n3015 gnd.n1365 240.244
R4864 gnd.n3020 gnd.n1365 240.244
R4865 gnd.n3020 gnd.n1374 240.244
R4866 gnd.n1070 gnd.n1069 240.244
R4867 gnd.n5039 gnd.n1069 240.244
R4868 gnd.n5037 gnd.n5036 240.244
R4869 gnd.n5033 gnd.n5032 240.244
R4870 gnd.n5029 gnd.n5028 240.244
R4871 gnd.n5025 gnd.n5024 240.244
R4872 gnd.n5021 gnd.n5020 240.244
R4873 gnd.n5017 gnd.n5016 240.244
R4874 gnd.n5013 gnd.n5012 240.244
R4875 gnd.n5008 gnd.n5007 240.244
R4876 gnd.n5004 gnd.n5003 240.244
R4877 gnd.n5000 gnd.n4999 240.244
R4878 gnd.n4996 gnd.n4995 240.244
R4879 gnd.n4992 gnd.n4991 240.244
R4880 gnd.n4988 gnd.n4987 240.244
R4881 gnd.n4984 gnd.n4983 240.244
R4882 gnd.n4980 gnd.n4979 240.244
R4883 gnd.n4976 gnd.n4975 240.244
R4884 gnd.n4972 gnd.n4971 240.244
R4885 gnd.n4968 gnd.n4967 240.244
R4886 gnd.n4964 gnd.n4963 240.244
R4887 gnd.n4960 gnd.n4959 240.244
R4888 gnd.n4956 gnd.n4955 240.244
R4889 gnd.n4952 gnd.n4951 240.244
R4890 gnd.n4948 gnd.n4947 240.244
R4891 gnd.n4944 gnd.n4943 240.244
R4892 gnd.n4940 gnd.n4939 240.244
R4893 gnd.n4936 gnd.n4935 240.244
R4894 gnd.n4932 gnd.n4931 240.244
R4895 gnd.n4921 gnd.n1071 240.244
R4896 gnd.n4921 gnd.n1144 240.244
R4897 gnd.n4917 gnd.n1144 240.244
R4898 gnd.n4917 gnd.n1151 240.244
R4899 gnd.n4909 gnd.n1151 240.244
R4900 gnd.n4909 gnd.n1168 240.244
R4901 gnd.n4905 gnd.n1168 240.244
R4902 gnd.n4905 gnd.n1174 240.244
R4903 gnd.n4897 gnd.n1174 240.244
R4904 gnd.n4897 gnd.n1187 240.244
R4905 gnd.n4893 gnd.n1187 240.244
R4906 gnd.n4893 gnd.n1193 240.244
R4907 gnd.n4885 gnd.n1193 240.244
R4908 gnd.n4885 gnd.n1208 240.244
R4909 gnd.n4881 gnd.n1208 240.244
R4910 gnd.n4881 gnd.n1214 240.244
R4911 gnd.n4873 gnd.n1214 240.244
R4912 gnd.n4873 gnd.n1228 240.244
R4913 gnd.n4869 gnd.n1228 240.244
R4914 gnd.n4869 gnd.n1234 240.244
R4915 gnd.n4861 gnd.n1234 240.244
R4916 gnd.n4861 gnd.n1249 240.244
R4917 gnd.n2859 gnd.n1249 240.244
R4918 gnd.n2859 gnd.n2623 240.244
R4919 gnd.n2885 gnd.n2623 240.244
R4920 gnd.n2888 gnd.n2885 240.244
R4921 gnd.n2888 gnd.n2613 240.244
R4922 gnd.n2899 gnd.n2613 240.244
R4923 gnd.n2902 gnd.n2899 240.244
R4924 gnd.n2902 gnd.n1261 240.244
R4925 gnd.n4855 gnd.n1261 240.244
R4926 gnd.n4855 gnd.n1262 240.244
R4927 gnd.n4847 gnd.n1262 240.244
R4928 gnd.n4847 gnd.n1277 240.244
R4929 gnd.n4843 gnd.n1277 240.244
R4930 gnd.n4843 gnd.n1282 240.244
R4931 gnd.n4835 gnd.n1282 240.244
R4932 gnd.n4835 gnd.n1297 240.244
R4933 gnd.n4831 gnd.n1297 240.244
R4934 gnd.n4831 gnd.n1303 240.244
R4935 gnd.n4823 gnd.n1303 240.244
R4936 gnd.n4823 gnd.n1316 240.244
R4937 gnd.n4819 gnd.n1316 240.244
R4938 gnd.n4819 gnd.n1322 240.244
R4939 gnd.n4811 gnd.n1322 240.244
R4940 gnd.n4811 gnd.n1337 240.244
R4941 gnd.n4807 gnd.n1337 240.244
R4942 gnd.n4807 gnd.n1343 240.244
R4943 gnd.n4799 gnd.n1343 240.244
R4944 gnd.n4799 gnd.n1357 240.244
R4945 gnd.n4795 gnd.n1357 240.244
R4946 gnd.n4795 gnd.n1363 240.244
R4947 gnd.n4787 gnd.n1363 240.244
R4948 gnd.n5054 gnd.n5049 240.244
R4949 gnd.n6419 gnd.n6418 240.244
R4950 gnd.n6416 gnd.n5058 240.244
R4951 gnd.n6412 gnd.n6411 240.244
R4952 gnd.n6409 gnd.n5065 240.244
R4953 gnd.n6405 gnd.n6404 240.244
R4954 gnd.n6402 gnd.n5072 240.244
R4955 gnd.n6398 gnd.n6397 240.244
R4956 gnd.n5689 gnd.n5409 240.244
R4957 gnd.n5409 gnd.n5400 240.244
R4958 gnd.n5707 gnd.n5400 240.244
R4959 gnd.n5708 gnd.n5707 240.244
R4960 gnd.n5708 gnd.n5388 240.244
R4961 gnd.n5388 gnd.n5377 240.244
R4962 gnd.n5739 gnd.n5377 240.244
R4963 gnd.n5740 gnd.n5739 240.244
R4964 gnd.n5741 gnd.n5740 240.244
R4965 gnd.n5741 gnd.n5362 240.244
R4966 gnd.n5743 gnd.n5362 240.244
R4967 gnd.n5743 gnd.n5347 240.244
R4968 gnd.n5784 gnd.n5347 240.244
R4969 gnd.n5785 gnd.n5784 240.244
R4970 gnd.n5788 gnd.n5785 240.244
R4971 gnd.n5788 gnd.n5329 240.244
R4972 gnd.n5820 gnd.n5329 240.244
R4973 gnd.n5820 gnd.n5315 240.244
R4974 gnd.n5842 gnd.n5315 240.244
R4975 gnd.n5843 gnd.n5842 240.244
R4976 gnd.n5843 gnd.n5302 240.244
R4977 gnd.n5302 gnd.n5291 240.244
R4978 gnd.n5874 gnd.n5291 240.244
R4979 gnd.n5875 gnd.n5874 240.244
R4980 gnd.n5876 gnd.n5875 240.244
R4981 gnd.n5876 gnd.n5212 240.244
R4982 gnd.n5212 gnd.n5211 240.244
R4983 gnd.n5211 gnd.n5196 240.244
R4984 gnd.n5927 gnd.n5196 240.244
R4985 gnd.n5928 gnd.n5927 240.244
R4986 gnd.n5928 gnd.n5183 240.244
R4987 gnd.n5183 gnd.n5172 240.244
R4988 gnd.n5961 gnd.n5172 240.244
R4989 gnd.n5962 gnd.n5961 240.244
R4990 gnd.n5964 gnd.n5962 240.244
R4991 gnd.n5964 gnd.n5963 240.244
R4992 gnd.n5963 gnd.n5152 240.244
R4993 gnd.n6001 gnd.n5152 240.244
R4994 gnd.n6001 gnd.n5139 240.244
R4995 gnd.n6027 gnd.n5139 240.244
R4996 gnd.n6028 gnd.n6027 240.244
R4997 gnd.n6029 gnd.n6028 240.244
R4998 gnd.n6029 gnd.n981 240.244
R4999 gnd.n6318 gnd.n981 240.244
R5000 gnd.n6318 gnd.n991 240.244
R5001 gnd.n6314 gnd.n991 240.244
R5002 gnd.n6314 gnd.n6313 240.244
R5003 gnd.n6313 gnd.n1004 240.244
R5004 gnd.n6309 gnd.n1004 240.244
R5005 gnd.n6309 gnd.n1017 240.244
R5006 gnd.n6305 gnd.n1017 240.244
R5007 gnd.n6305 gnd.n6304 240.244
R5008 gnd.n6304 gnd.n1029 240.244
R5009 gnd.n5626 gnd.n5625 240.244
R5010 gnd.n5670 gnd.n5625 240.244
R5011 gnd.n5668 gnd.n5667 240.244
R5012 gnd.n5664 gnd.n5663 240.244
R5013 gnd.n5660 gnd.n5659 240.244
R5014 gnd.n5656 gnd.n5655 240.244
R5015 gnd.n5652 gnd.n5651 240.244
R5016 gnd.n5648 gnd.n5647 240.244
R5017 gnd.n5699 gnd.n5407 240.244
R5018 gnd.n5699 gnd.n5403 240.244
R5019 gnd.n5705 gnd.n5403 240.244
R5020 gnd.n5705 gnd.n5386 240.244
R5021 gnd.n5729 gnd.n5386 240.244
R5022 gnd.n5729 gnd.n5381 240.244
R5023 gnd.n5737 gnd.n5381 240.244
R5024 gnd.n5737 gnd.n5382 240.244
R5025 gnd.n5382 gnd.n5360 240.244
R5026 gnd.n5763 gnd.n5360 240.244
R5027 gnd.n5763 gnd.n5355 240.244
R5028 gnd.n5774 gnd.n5355 240.244
R5029 gnd.n5774 gnd.n5356 240.244
R5030 gnd.n5770 gnd.n5356 240.244
R5031 gnd.n5770 gnd.n5327 240.244
R5032 gnd.n5824 gnd.n5327 240.244
R5033 gnd.n5824 gnd.n5322 240.244
R5034 gnd.n5832 gnd.n5322 240.244
R5035 gnd.n5832 gnd.n5323 240.244
R5036 gnd.n5323 gnd.n5300 240.244
R5037 gnd.n5864 gnd.n5300 240.244
R5038 gnd.n5864 gnd.n5295 240.244
R5039 gnd.n5872 gnd.n5295 240.244
R5040 gnd.n5872 gnd.n5296 240.244
R5041 gnd.n5296 gnd.n5209 240.244
R5042 gnd.n5909 gnd.n5209 240.244
R5043 gnd.n5909 gnd.n5204 240.244
R5044 gnd.n5917 gnd.n5204 240.244
R5045 gnd.n5917 gnd.n5205 240.244
R5046 gnd.n5205 gnd.n5181 240.244
R5047 gnd.n5948 gnd.n5181 240.244
R5048 gnd.n5948 gnd.n5176 240.244
R5049 gnd.n5959 gnd.n5176 240.244
R5050 gnd.n5959 gnd.n5177 240.244
R5051 gnd.n5955 gnd.n5177 240.244
R5052 gnd.n5955 gnd.n5151 240.244
R5053 gnd.n6005 gnd.n5151 240.244
R5054 gnd.n6005 gnd.n5146 240.244
R5055 gnd.n6017 gnd.n5146 240.244
R5056 gnd.n6017 gnd.n5147 240.244
R5057 gnd.n6013 gnd.n5147 240.244
R5058 gnd.n6013 gnd.n982 240.244
R5059 gnd.n6454 gnd.n982 240.244
R5060 gnd.n6454 gnd.n983 240.244
R5061 gnd.n6450 gnd.n983 240.244
R5062 gnd.n6450 gnd.n989 240.244
R5063 gnd.n1006 gnd.n989 240.244
R5064 gnd.n6440 gnd.n1006 240.244
R5065 gnd.n6440 gnd.n1007 240.244
R5066 gnd.n6436 gnd.n1007 240.244
R5067 gnd.n6436 gnd.n1015 240.244
R5068 gnd.n5048 gnd.n1015 240.244
R5069 gnd.n6426 gnd.n5048 240.244
R5070 gnd.n319 gnd.n208 240.244
R5071 gnd.n7439 gnd.n7438 240.244
R5072 gnd.n7436 gnd.n323 240.244
R5073 gnd.n7432 gnd.n7431 240.244
R5074 gnd.n7429 gnd.n330 240.244
R5075 gnd.n7425 gnd.n7424 240.244
R5076 gnd.n7422 gnd.n337 240.244
R5077 gnd.n7418 gnd.n7417 240.244
R5078 gnd.n7415 gnd.n344 240.244
R5079 gnd.n3755 gnd.n1601 240.244
R5080 gnd.n3755 gnd.n1613 240.244
R5081 gnd.n4334 gnd.n1613 240.244
R5082 gnd.n4334 gnd.n1625 240.244
R5083 gnd.n4340 gnd.n1625 240.244
R5084 gnd.n4340 gnd.n1636 240.244
R5085 gnd.n4348 gnd.n1636 240.244
R5086 gnd.n4348 gnd.n1645 240.244
R5087 gnd.n4354 gnd.n1645 240.244
R5088 gnd.n4354 gnd.n1656 240.244
R5089 gnd.n4390 gnd.n1656 240.244
R5090 gnd.n4390 gnd.n1665 240.244
R5091 gnd.n1760 gnd.n1665 240.244
R5092 gnd.n1760 gnd.n1676 240.244
R5093 gnd.n1761 gnd.n1676 240.244
R5094 gnd.n1761 gnd.n1685 240.244
R5095 gnd.n4375 gnd.n1685 240.244
R5096 gnd.n4375 gnd.n1696 240.244
R5097 gnd.n1743 gnd.n1696 240.244
R5098 gnd.n1743 gnd.n1705 240.244
R5099 gnd.n4446 gnd.n1705 240.244
R5100 gnd.n4446 gnd.n1714 240.244
R5101 gnd.n4455 gnd.n1714 240.244
R5102 gnd.n4455 gnd.n1723 240.244
R5103 gnd.n1730 gnd.n1723 240.244
R5104 gnd.n1731 gnd.n1730 240.244
R5105 gnd.n1731 gnd.n82 240.244
R5106 gnd.n7632 gnd.n82 240.244
R5107 gnd.n7632 gnd.n84 240.244
R5108 gnd.n7327 gnd.n84 240.244
R5109 gnd.n7327 gnd.n104 240.244
R5110 gnd.n7335 gnd.n104 240.244
R5111 gnd.n7335 gnd.n116 240.244
R5112 gnd.n7341 gnd.n116 240.244
R5113 gnd.n7341 gnd.n125 240.244
R5114 gnd.n7349 gnd.n125 240.244
R5115 gnd.n7349 gnd.n134 240.244
R5116 gnd.n7355 gnd.n134 240.244
R5117 gnd.n7355 gnd.n145 240.244
R5118 gnd.n7363 gnd.n145 240.244
R5119 gnd.n7363 gnd.n155 240.244
R5120 gnd.n7370 gnd.n155 240.244
R5121 gnd.n7370 gnd.n165 240.244
R5122 gnd.n7393 gnd.n165 240.244
R5123 gnd.n7393 gnd.n174 240.244
R5124 gnd.n356 gnd.n174 240.244
R5125 gnd.n356 gnd.n184 240.244
R5126 gnd.n7400 gnd.n184 240.244
R5127 gnd.n7400 gnd.n193 240.244
R5128 gnd.n353 gnd.n193 240.244
R5129 gnd.n353 gnd.n203 240.244
R5130 gnd.n7407 gnd.n203 240.244
R5131 gnd.n7407 gnd.n211 240.244
R5132 gnd.n3855 gnd.n3803 240.244
R5133 gnd.n3859 gnd.n3857 240.244
R5134 gnd.n3874 gnd.n3794 240.244
R5135 gnd.n3878 gnd.n3876 240.244
R5136 gnd.n3893 gnd.n3785 240.244
R5137 gnd.n3897 gnd.n3895 240.244
R5138 gnd.n3913 gnd.n3776 240.244
R5139 gnd.n3917 gnd.n3915 240.244
R5140 gnd.n3772 gnd.n3771 240.244
R5141 gnd.n1615 gnd.n1603 240.244
R5142 gnd.n4539 gnd.n1615 240.244
R5143 gnd.n4539 gnd.n1616 240.244
R5144 gnd.n4535 gnd.n1616 240.244
R5145 gnd.n4535 gnd.n1622 240.244
R5146 gnd.n4527 gnd.n1622 240.244
R5147 gnd.n4527 gnd.n1637 240.244
R5148 gnd.n4523 gnd.n1637 240.244
R5149 gnd.n4523 gnd.n1642 240.244
R5150 gnd.n4515 gnd.n1642 240.244
R5151 gnd.n4515 gnd.n1658 240.244
R5152 gnd.n4511 gnd.n1658 240.244
R5153 gnd.n4511 gnd.n1663 240.244
R5154 gnd.n4503 gnd.n1663 240.244
R5155 gnd.n4503 gnd.n1677 240.244
R5156 gnd.n4499 gnd.n1677 240.244
R5157 gnd.n4499 gnd.n1682 240.244
R5158 gnd.n4491 gnd.n1682 240.244
R5159 gnd.n4491 gnd.n1698 240.244
R5160 gnd.n4487 gnd.n1698 240.244
R5161 gnd.n4487 gnd.n1703 240.244
R5162 gnd.n4479 gnd.n1703 240.244
R5163 gnd.n4479 gnd.n1715 240.244
R5164 gnd.n4475 gnd.n1715 240.244
R5165 gnd.n4475 gnd.n1720 240.244
R5166 gnd.n4424 gnd.n1720 240.244
R5167 gnd.n4434 gnd.n4424 240.244
R5168 gnd.n4434 gnd.n88 240.244
R5169 gnd.n4430 gnd.n88 240.244
R5170 gnd.n4430 gnd.n106 240.244
R5171 gnd.n7622 gnd.n106 240.244
R5172 gnd.n7622 gnd.n107 240.244
R5173 gnd.n7618 gnd.n107 240.244
R5174 gnd.n7618 gnd.n113 240.244
R5175 gnd.n7610 gnd.n113 240.244
R5176 gnd.n7610 gnd.n126 240.244
R5177 gnd.n7606 gnd.n126 240.244
R5178 gnd.n7606 gnd.n131 240.244
R5179 gnd.n7598 gnd.n131 240.244
R5180 gnd.n7598 gnd.n147 240.244
R5181 gnd.n7594 gnd.n147 240.244
R5182 gnd.n7594 gnd.n152 240.244
R5183 gnd.n7586 gnd.n152 240.244
R5184 gnd.n7586 gnd.n166 240.244
R5185 gnd.n7582 gnd.n166 240.244
R5186 gnd.n7582 gnd.n171 240.244
R5187 gnd.n7574 gnd.n171 240.244
R5188 gnd.n7574 gnd.n186 240.244
R5189 gnd.n7570 gnd.n186 240.244
R5190 gnd.n7570 gnd.n191 240.244
R5191 gnd.n7562 gnd.n191 240.244
R5192 gnd.n7562 gnd.n204 240.244
R5193 gnd.n7558 gnd.n204 240.244
R5194 gnd.n5084 gnd.n1026 240.244
R5195 gnd.n6387 gnd.n6386 240.244
R5196 gnd.n6384 gnd.n5088 240.244
R5197 gnd.n6380 gnd.n6379 240.244
R5198 gnd.n6377 gnd.n5095 240.244
R5199 gnd.n6373 gnd.n6372 240.244
R5200 gnd.n6370 gnd.n5102 240.244
R5201 gnd.n6366 gnd.n6365 240.244
R5202 gnd.n6363 gnd.n5109 240.244
R5203 gnd.n6359 gnd.n6358 240.244
R5204 gnd.n6356 gnd.n5116 240.244
R5205 gnd.n6352 gnd.n6351 240.244
R5206 gnd.n6349 gnd.n5126 240.244
R5207 gnd.n5557 gnd.n5453 240.244
R5208 gnd.n5563 gnd.n5453 240.244
R5209 gnd.n5563 gnd.n5445 240.244
R5210 gnd.n5573 gnd.n5445 240.244
R5211 gnd.n5573 gnd.n5441 240.244
R5212 gnd.n5579 gnd.n5441 240.244
R5213 gnd.n5579 gnd.n5432 240.244
R5214 gnd.n5589 gnd.n5432 240.244
R5215 gnd.n5589 gnd.n5427 240.244
R5216 gnd.n5617 gnd.n5427 240.244
R5217 gnd.n5617 gnd.n5428 240.244
R5218 gnd.n5428 gnd.n5420 240.244
R5219 gnd.n5612 gnd.n5420 240.244
R5220 gnd.n5612 gnd.n5410 240.244
R5221 gnd.n5609 gnd.n5410 240.244
R5222 gnd.n5609 gnd.n5399 240.244
R5223 gnd.n5606 gnd.n5399 240.244
R5224 gnd.n5606 gnd.n5389 240.244
R5225 gnd.n5603 gnd.n5389 240.244
R5226 gnd.n5603 gnd.n5367 240.244
R5227 gnd.n5752 gnd.n5367 240.244
R5228 gnd.n5752 gnd.n5363 240.244
R5229 gnd.n5760 gnd.n5363 240.244
R5230 gnd.n5760 gnd.n5353 240.244
R5231 gnd.n5353 gnd.n5334 240.244
R5232 gnd.n5799 gnd.n5334 240.244
R5233 gnd.n5799 gnd.n5335 240.244
R5234 gnd.n5335 gnd.n5330 240.244
R5235 gnd.n5819 gnd.n5330 240.244
R5236 gnd.n5819 gnd.n5320 240.244
R5237 gnd.n5814 gnd.n5320 240.244
R5238 gnd.n5814 gnd.n5314 240.244
R5239 gnd.n5810 gnd.n5314 240.244
R5240 gnd.n5810 gnd.n5303 240.244
R5241 gnd.n5806 gnd.n5303 240.244
R5242 gnd.n5806 gnd.n5281 240.244
R5243 gnd.n5885 gnd.n5281 240.244
R5244 gnd.n5885 gnd.n5213 240.244
R5245 gnd.n5906 gnd.n5213 240.244
R5246 gnd.n5906 gnd.n5202 240.244
R5247 gnd.n5902 gnd.n5202 240.244
R5248 gnd.n5902 gnd.n5195 240.244
R5249 gnd.n5899 gnd.n5195 240.244
R5250 gnd.n5899 gnd.n5184 240.244
R5251 gnd.n5896 gnd.n5184 240.244
R5252 gnd.n5896 gnd.n5163 240.244
R5253 gnd.n5971 gnd.n5163 240.244
R5254 gnd.n5971 gnd.n5159 240.244
R5255 gnd.n5992 gnd.n5159 240.244
R5256 gnd.n5992 gnd.n5153 240.244
R5257 gnd.n5153 gnd.n5144 240.244
R5258 gnd.n5987 gnd.n5144 240.244
R5259 gnd.n5987 gnd.n969 240.244
R5260 gnd.n5984 gnd.n969 240.244
R5261 gnd.n5984 gnd.n980 240.244
R5262 gnd.n6321 gnd.n980 240.244
R5263 gnd.n6322 gnd.n6321 240.244
R5264 gnd.n6322 gnd.n992 240.244
R5265 gnd.n6328 gnd.n992 240.244
R5266 gnd.n6328 gnd.n1003 240.244
R5267 gnd.n6332 gnd.n1003 240.244
R5268 gnd.n6332 gnd.n6331 240.244
R5269 gnd.n6331 gnd.n1018 240.244
R5270 gnd.n6339 gnd.n1018 240.244
R5271 gnd.n6339 gnd.n1028 240.244
R5272 gnd.n5549 gnd.n5547 240.244
R5273 gnd.n5547 gnd.n5546 240.244
R5274 gnd.n5543 gnd.n5542 240.244
R5275 gnd.n5540 gnd.n5466 240.244
R5276 gnd.n5536 gnd.n5534 240.244
R5277 gnd.n5532 gnd.n5472 240.244
R5278 gnd.n5528 gnd.n5526 240.244
R5279 gnd.n5524 gnd.n5478 240.244
R5280 gnd.n5520 gnd.n5518 240.244
R5281 gnd.n5516 gnd.n5484 240.244
R5282 gnd.n5512 gnd.n5510 240.244
R5283 gnd.n5508 gnd.n5490 240.244
R5284 gnd.n5503 gnd.n5501 240.244
R5285 gnd.n5555 gnd.n5451 240.244
R5286 gnd.n5565 gnd.n5451 240.244
R5287 gnd.n5565 gnd.n5447 240.244
R5288 gnd.n5571 gnd.n5447 240.244
R5289 gnd.n5571 gnd.n5439 240.244
R5290 gnd.n5581 gnd.n5439 240.244
R5291 gnd.n5581 gnd.n5435 240.244
R5292 gnd.n5587 gnd.n5435 240.244
R5293 gnd.n5587 gnd.n5426 240.244
R5294 gnd.n5679 gnd.n5426 240.244
R5295 gnd.n5679 gnd.n5421 240.244
R5296 gnd.n5686 gnd.n5421 240.244
R5297 gnd.n5686 gnd.n5412 240.244
R5298 gnd.n5696 gnd.n5412 240.244
R5299 gnd.n5696 gnd.n5398 240.244
R5300 gnd.n5711 gnd.n5398 240.244
R5301 gnd.n5711 gnd.n5391 240.244
R5302 gnd.n5726 gnd.n5391 240.244
R5303 gnd.n5726 gnd.n5392 240.244
R5304 gnd.n5392 gnd.n5370 240.244
R5305 gnd.n5750 gnd.n5370 240.244
R5306 gnd.n5750 gnd.n5371 240.244
R5307 gnd.n5371 gnd.n5351 240.244
R5308 gnd.n5777 gnd.n5351 240.244
R5309 gnd.n5777 gnd.n5338 240.244
R5310 gnd.n5797 gnd.n5338 240.244
R5311 gnd.n5797 gnd.n5339 240.244
R5312 gnd.n5793 gnd.n5339 240.244
R5313 gnd.n5793 gnd.n5319 240.244
R5314 gnd.n5835 gnd.n5319 240.244
R5315 gnd.n5835 gnd.n5312 240.244
R5316 gnd.n5846 gnd.n5312 240.244
R5317 gnd.n5846 gnd.n5305 240.244
R5318 gnd.n5861 gnd.n5305 240.244
R5319 gnd.n5861 gnd.n5306 240.244
R5320 gnd.n5306 gnd.n5284 240.244
R5321 gnd.n5883 gnd.n5284 240.244
R5322 gnd.n5883 gnd.n5285 240.244
R5323 gnd.n5285 gnd.n5200 240.244
R5324 gnd.n5920 gnd.n5200 240.244
R5325 gnd.n5920 gnd.n5193 240.244
R5326 gnd.n5931 gnd.n5193 240.244
R5327 gnd.n5931 gnd.n5186 240.244
R5328 gnd.n5945 gnd.n5186 240.244
R5329 gnd.n5945 gnd.n5187 240.244
R5330 gnd.n5187 gnd.n5167 240.244
R5331 gnd.n5969 gnd.n5167 240.244
R5332 gnd.n5969 gnd.n5157 240.244
R5333 gnd.n5994 gnd.n5157 240.244
R5334 gnd.n5994 gnd.n5143 240.244
R5335 gnd.n6020 gnd.n5143 240.244
R5336 gnd.n6020 gnd.n971 240.244
R5337 gnd.n6461 gnd.n971 240.244
R5338 gnd.n6461 gnd.n972 240.244
R5339 gnd.n6457 gnd.n972 240.244
R5340 gnd.n6457 gnd.n978 240.244
R5341 gnd.n994 gnd.n978 240.244
R5342 gnd.n6447 gnd.n994 240.244
R5343 gnd.n6447 gnd.n995 240.244
R5344 gnd.n6443 gnd.n995 240.244
R5345 gnd.n6443 gnd.n1001 240.244
R5346 gnd.n1020 gnd.n1001 240.244
R5347 gnd.n6433 gnd.n1020 240.244
R5348 gnd.n6433 gnd.n1021 240.244
R5349 gnd.n6429 gnd.n1021 240.244
R5350 gnd.n2466 gnd.n1372 240.244
R5351 gnd.n2475 gnd.n2468 240.244
R5352 gnd.n2478 gnd.n2477 240.244
R5353 gnd.n2487 gnd.n2486 240.244
R5354 gnd.n2496 gnd.n2489 240.244
R5355 gnd.n2499 gnd.n2498 240.244
R5356 gnd.n2508 gnd.n2507 240.244
R5357 gnd.n2519 gnd.n2510 240.244
R5358 gnd.n2525 gnd.n2521 240.244
R5359 gnd.n2743 gnd.n1142 240.244
R5360 gnd.n2748 gnd.n1142 240.244
R5361 gnd.n2748 gnd.n1154 240.244
R5362 gnd.n2751 gnd.n1154 240.244
R5363 gnd.n2751 gnd.n1166 240.244
R5364 gnd.n2756 gnd.n1166 240.244
R5365 gnd.n2756 gnd.n1176 240.244
R5366 gnd.n2759 gnd.n1176 240.244
R5367 gnd.n2759 gnd.n1186 240.244
R5368 gnd.n2765 gnd.n1186 240.244
R5369 gnd.n2765 gnd.n1196 240.244
R5370 gnd.n2773 gnd.n1196 240.244
R5371 gnd.n2773 gnd.n1206 240.244
R5372 gnd.n2779 gnd.n1206 240.244
R5373 gnd.n2779 gnd.n1216 240.244
R5374 gnd.n2826 gnd.n1216 240.244
R5375 gnd.n2826 gnd.n1226 240.244
R5376 gnd.n2833 gnd.n1226 240.244
R5377 gnd.n2833 gnd.n1237 240.244
R5378 gnd.n2842 gnd.n1237 240.244
R5379 gnd.n2842 gnd.n1247 240.244
R5380 gnd.n2845 gnd.n1247 240.244
R5381 gnd.n2845 gnd.n2642 240.244
R5382 gnd.n2851 gnd.n2642 240.244
R5383 gnd.n2851 gnd.n2619 240.244
R5384 gnd.n2890 gnd.n2619 240.244
R5385 gnd.n2890 gnd.n2615 240.244
R5386 gnd.n2897 gnd.n2615 240.244
R5387 gnd.n2897 gnd.n2599 240.244
R5388 gnd.n2938 gnd.n2599 240.244
R5389 gnd.n2938 gnd.n1264 240.244
R5390 gnd.n2604 gnd.n1264 240.244
R5391 gnd.n2604 gnd.n1276 240.244
R5392 gnd.n2605 gnd.n1276 240.244
R5393 gnd.n2605 gnd.n1285 240.244
R5394 gnd.n2926 gnd.n1285 240.244
R5395 gnd.n2926 gnd.n1295 240.244
R5396 gnd.n2980 gnd.n1295 240.244
R5397 gnd.n2980 gnd.n1305 240.244
R5398 gnd.n2986 gnd.n1305 240.244
R5399 gnd.n2986 gnd.n1315 240.244
R5400 gnd.n2995 gnd.n1315 240.244
R5401 gnd.n2995 gnd.n1325 240.244
R5402 gnd.n3001 gnd.n1325 240.244
R5403 gnd.n3001 gnd.n1335 240.244
R5404 gnd.n3035 gnd.n1335 240.244
R5405 gnd.n3035 gnd.n1345 240.244
R5406 gnd.n2572 gnd.n1345 240.244
R5407 gnd.n2572 gnd.n1355 240.244
R5408 gnd.n2573 gnd.n1355 240.244
R5409 gnd.n2573 gnd.n1366 240.244
R5410 gnd.n3022 gnd.n1366 240.244
R5411 gnd.n3022 gnd.n1375 240.244
R5412 gnd.n2704 gnd.n2703 240.244
R5413 gnd.n2710 gnd.n2709 240.244
R5414 gnd.n2714 gnd.n2713 240.244
R5415 gnd.n2720 gnd.n2719 240.244
R5416 gnd.n2724 gnd.n2723 240.244
R5417 gnd.n2730 gnd.n2729 240.244
R5418 gnd.n2734 gnd.n2733 240.244
R5419 gnd.n2691 gnd.n2690 240.244
R5420 gnd.n2686 gnd.n1067 240.244
R5421 gnd.n2699 gnd.n1143 240.244
R5422 gnd.n1156 gnd.n1143 240.244
R5423 gnd.n4915 gnd.n1156 240.244
R5424 gnd.n4915 gnd.n1157 240.244
R5425 gnd.n4911 gnd.n1157 240.244
R5426 gnd.n4911 gnd.n1164 240.244
R5427 gnd.n4903 gnd.n1164 240.244
R5428 gnd.n4903 gnd.n1178 240.244
R5429 gnd.n4899 gnd.n1178 240.244
R5430 gnd.n4899 gnd.n1183 240.244
R5431 gnd.n4891 gnd.n1183 240.244
R5432 gnd.n4891 gnd.n1198 240.244
R5433 gnd.n4887 gnd.n1198 240.244
R5434 gnd.n4887 gnd.n1203 240.244
R5435 gnd.n4879 gnd.n1203 240.244
R5436 gnd.n4879 gnd.n1218 240.244
R5437 gnd.n4875 gnd.n1218 240.244
R5438 gnd.n4875 gnd.n1223 240.244
R5439 gnd.n4867 gnd.n1223 240.244
R5440 gnd.n4867 gnd.n1239 240.244
R5441 gnd.n4863 gnd.n1239 240.244
R5442 gnd.n4863 gnd.n1244 240.244
R5443 gnd.n2858 gnd.n1244 240.244
R5444 gnd.n2858 gnd.n2628 240.244
R5445 gnd.n2883 gnd.n2628 240.244
R5446 gnd.n2883 gnd.n2622 240.244
R5447 gnd.n2879 gnd.n2622 240.244
R5448 gnd.n2879 gnd.n2610 240.244
R5449 gnd.n2904 gnd.n2610 240.244
R5450 gnd.n2904 gnd.n1266 240.244
R5451 gnd.n4853 gnd.n1266 240.244
R5452 gnd.n4853 gnd.n1267 240.244
R5453 gnd.n4849 gnd.n1267 240.244
R5454 gnd.n4849 gnd.n1273 240.244
R5455 gnd.n4841 gnd.n1273 240.244
R5456 gnd.n4841 gnd.n1287 240.244
R5457 gnd.n4837 gnd.n1287 240.244
R5458 gnd.n4837 gnd.n1292 240.244
R5459 gnd.n4829 gnd.n1292 240.244
R5460 gnd.n4829 gnd.n1307 240.244
R5461 gnd.n4825 gnd.n1307 240.244
R5462 gnd.n4825 gnd.n1312 240.244
R5463 gnd.n4817 gnd.n1312 240.244
R5464 gnd.n4817 gnd.n1327 240.244
R5465 gnd.n4813 gnd.n1327 240.244
R5466 gnd.n4813 gnd.n1332 240.244
R5467 gnd.n4805 gnd.n1332 240.244
R5468 gnd.n4805 gnd.n1347 240.244
R5469 gnd.n4801 gnd.n1347 240.244
R5470 gnd.n4801 gnd.n1352 240.244
R5471 gnd.n4793 gnd.n1352 240.244
R5472 gnd.n4793 gnd.n1368 240.244
R5473 gnd.n4789 gnd.n1368 240.244
R5474 gnd.n6634 gnd.n800 240.244
R5475 gnd.n6634 gnd.n796 240.244
R5476 gnd.n6640 gnd.n796 240.244
R5477 gnd.n6640 gnd.n794 240.244
R5478 gnd.n6644 gnd.n794 240.244
R5479 gnd.n6644 gnd.n790 240.244
R5480 gnd.n6650 gnd.n790 240.244
R5481 gnd.n6650 gnd.n788 240.244
R5482 gnd.n6654 gnd.n788 240.244
R5483 gnd.n6654 gnd.n784 240.244
R5484 gnd.n6660 gnd.n784 240.244
R5485 gnd.n6660 gnd.n782 240.244
R5486 gnd.n6664 gnd.n782 240.244
R5487 gnd.n6664 gnd.n778 240.244
R5488 gnd.n6670 gnd.n778 240.244
R5489 gnd.n6670 gnd.n776 240.244
R5490 gnd.n6674 gnd.n776 240.244
R5491 gnd.n6674 gnd.n772 240.244
R5492 gnd.n6680 gnd.n772 240.244
R5493 gnd.n6680 gnd.n770 240.244
R5494 gnd.n6684 gnd.n770 240.244
R5495 gnd.n6684 gnd.n766 240.244
R5496 gnd.n6690 gnd.n766 240.244
R5497 gnd.n6690 gnd.n764 240.244
R5498 gnd.n6694 gnd.n764 240.244
R5499 gnd.n6694 gnd.n760 240.244
R5500 gnd.n6700 gnd.n760 240.244
R5501 gnd.n6700 gnd.n758 240.244
R5502 gnd.n6704 gnd.n758 240.244
R5503 gnd.n6704 gnd.n754 240.244
R5504 gnd.n6710 gnd.n754 240.244
R5505 gnd.n6710 gnd.n752 240.244
R5506 gnd.n6714 gnd.n752 240.244
R5507 gnd.n6714 gnd.n748 240.244
R5508 gnd.n6720 gnd.n748 240.244
R5509 gnd.n6720 gnd.n746 240.244
R5510 gnd.n6724 gnd.n746 240.244
R5511 gnd.n6724 gnd.n742 240.244
R5512 gnd.n6730 gnd.n742 240.244
R5513 gnd.n6730 gnd.n740 240.244
R5514 gnd.n6734 gnd.n740 240.244
R5515 gnd.n6734 gnd.n736 240.244
R5516 gnd.n6740 gnd.n736 240.244
R5517 gnd.n6740 gnd.n734 240.244
R5518 gnd.n6744 gnd.n734 240.244
R5519 gnd.n6744 gnd.n730 240.244
R5520 gnd.n6750 gnd.n730 240.244
R5521 gnd.n6750 gnd.n728 240.244
R5522 gnd.n6754 gnd.n728 240.244
R5523 gnd.n6754 gnd.n724 240.244
R5524 gnd.n6760 gnd.n724 240.244
R5525 gnd.n6760 gnd.n722 240.244
R5526 gnd.n6764 gnd.n722 240.244
R5527 gnd.n6764 gnd.n718 240.244
R5528 gnd.n6770 gnd.n718 240.244
R5529 gnd.n6770 gnd.n716 240.244
R5530 gnd.n6774 gnd.n716 240.244
R5531 gnd.n6774 gnd.n712 240.244
R5532 gnd.n6780 gnd.n712 240.244
R5533 gnd.n6780 gnd.n710 240.244
R5534 gnd.n6784 gnd.n710 240.244
R5535 gnd.n6784 gnd.n706 240.244
R5536 gnd.n6790 gnd.n706 240.244
R5537 gnd.n6790 gnd.n704 240.244
R5538 gnd.n6794 gnd.n704 240.244
R5539 gnd.n6794 gnd.n700 240.244
R5540 gnd.n6800 gnd.n700 240.244
R5541 gnd.n6800 gnd.n698 240.244
R5542 gnd.n6804 gnd.n698 240.244
R5543 gnd.n6804 gnd.n694 240.244
R5544 gnd.n6810 gnd.n694 240.244
R5545 gnd.n6810 gnd.n692 240.244
R5546 gnd.n6814 gnd.n692 240.244
R5547 gnd.n6814 gnd.n688 240.244
R5548 gnd.n6820 gnd.n688 240.244
R5549 gnd.n6820 gnd.n686 240.244
R5550 gnd.n6824 gnd.n686 240.244
R5551 gnd.n6824 gnd.n682 240.244
R5552 gnd.n6830 gnd.n682 240.244
R5553 gnd.n6830 gnd.n680 240.244
R5554 gnd.n6834 gnd.n680 240.244
R5555 gnd.n6834 gnd.n676 240.244
R5556 gnd.n6840 gnd.n676 240.244
R5557 gnd.n6840 gnd.n674 240.244
R5558 gnd.n6844 gnd.n674 240.244
R5559 gnd.n6844 gnd.n670 240.244
R5560 gnd.n6850 gnd.n670 240.244
R5561 gnd.n6850 gnd.n668 240.244
R5562 gnd.n6854 gnd.n668 240.244
R5563 gnd.n6854 gnd.n664 240.244
R5564 gnd.n6860 gnd.n664 240.244
R5565 gnd.n6860 gnd.n662 240.244
R5566 gnd.n6864 gnd.n662 240.244
R5567 gnd.n6864 gnd.n658 240.244
R5568 gnd.n6870 gnd.n658 240.244
R5569 gnd.n6870 gnd.n656 240.244
R5570 gnd.n6874 gnd.n656 240.244
R5571 gnd.n6874 gnd.n652 240.244
R5572 gnd.n6880 gnd.n652 240.244
R5573 gnd.n6880 gnd.n650 240.244
R5574 gnd.n6884 gnd.n650 240.244
R5575 gnd.n6884 gnd.n646 240.244
R5576 gnd.n6890 gnd.n646 240.244
R5577 gnd.n6890 gnd.n644 240.244
R5578 gnd.n6894 gnd.n644 240.244
R5579 gnd.n6894 gnd.n640 240.244
R5580 gnd.n6900 gnd.n640 240.244
R5581 gnd.n6900 gnd.n638 240.244
R5582 gnd.n6904 gnd.n638 240.244
R5583 gnd.n6904 gnd.n634 240.244
R5584 gnd.n6910 gnd.n634 240.244
R5585 gnd.n6910 gnd.n632 240.244
R5586 gnd.n6914 gnd.n632 240.244
R5587 gnd.n6914 gnd.n628 240.244
R5588 gnd.n6920 gnd.n628 240.244
R5589 gnd.n6920 gnd.n626 240.244
R5590 gnd.n6924 gnd.n626 240.244
R5591 gnd.n6924 gnd.n622 240.244
R5592 gnd.n6930 gnd.n622 240.244
R5593 gnd.n6930 gnd.n620 240.244
R5594 gnd.n6934 gnd.n620 240.244
R5595 gnd.n6934 gnd.n616 240.244
R5596 gnd.n6940 gnd.n616 240.244
R5597 gnd.n6940 gnd.n614 240.244
R5598 gnd.n6944 gnd.n614 240.244
R5599 gnd.n6944 gnd.n610 240.244
R5600 gnd.n6950 gnd.n610 240.244
R5601 gnd.n6950 gnd.n608 240.244
R5602 gnd.n6954 gnd.n608 240.244
R5603 gnd.n6954 gnd.n604 240.244
R5604 gnd.n6960 gnd.n604 240.244
R5605 gnd.n6960 gnd.n602 240.244
R5606 gnd.n6964 gnd.n602 240.244
R5607 gnd.n6964 gnd.n598 240.244
R5608 gnd.n6970 gnd.n598 240.244
R5609 gnd.n6970 gnd.n596 240.244
R5610 gnd.n6974 gnd.n596 240.244
R5611 gnd.n6974 gnd.n592 240.244
R5612 gnd.n6980 gnd.n592 240.244
R5613 gnd.n6980 gnd.n590 240.244
R5614 gnd.n6984 gnd.n590 240.244
R5615 gnd.n6984 gnd.n586 240.244
R5616 gnd.n6990 gnd.n586 240.244
R5617 gnd.n6990 gnd.n584 240.244
R5618 gnd.n6994 gnd.n584 240.244
R5619 gnd.n6994 gnd.n580 240.244
R5620 gnd.n7000 gnd.n580 240.244
R5621 gnd.n7000 gnd.n578 240.244
R5622 gnd.n7004 gnd.n578 240.244
R5623 gnd.n7004 gnd.n574 240.244
R5624 gnd.n7010 gnd.n574 240.244
R5625 gnd.n7010 gnd.n572 240.244
R5626 gnd.n7014 gnd.n572 240.244
R5627 gnd.n7014 gnd.n568 240.244
R5628 gnd.n7020 gnd.n568 240.244
R5629 gnd.n7020 gnd.n566 240.244
R5630 gnd.n7024 gnd.n566 240.244
R5631 gnd.n7024 gnd.n562 240.244
R5632 gnd.n7030 gnd.n562 240.244
R5633 gnd.n7030 gnd.n560 240.244
R5634 gnd.n7034 gnd.n560 240.244
R5635 gnd.n7034 gnd.n556 240.244
R5636 gnd.n7040 gnd.n556 240.244
R5637 gnd.n7040 gnd.n554 240.244
R5638 gnd.n7044 gnd.n554 240.244
R5639 gnd.n7044 gnd.n550 240.244
R5640 gnd.n7050 gnd.n550 240.244
R5641 gnd.n7050 gnd.n548 240.244
R5642 gnd.n7054 gnd.n548 240.244
R5643 gnd.n7054 gnd.n544 240.244
R5644 gnd.n7060 gnd.n544 240.244
R5645 gnd.n7060 gnd.n542 240.244
R5646 gnd.n7064 gnd.n542 240.244
R5647 gnd.n7064 gnd.n538 240.244
R5648 gnd.n7070 gnd.n538 240.244
R5649 gnd.n7070 gnd.n536 240.244
R5650 gnd.n7074 gnd.n536 240.244
R5651 gnd.n7074 gnd.n532 240.244
R5652 gnd.n7080 gnd.n532 240.244
R5653 gnd.n7080 gnd.n530 240.244
R5654 gnd.n7084 gnd.n530 240.244
R5655 gnd.n7090 gnd.n526 240.244
R5656 gnd.n7090 gnd.n524 240.244
R5657 gnd.n7094 gnd.n524 240.244
R5658 gnd.n7094 gnd.n520 240.244
R5659 gnd.n7100 gnd.n520 240.244
R5660 gnd.n7100 gnd.n518 240.244
R5661 gnd.n7104 gnd.n518 240.244
R5662 gnd.n7104 gnd.n514 240.244
R5663 gnd.n7110 gnd.n514 240.244
R5664 gnd.n7110 gnd.n512 240.244
R5665 gnd.n7114 gnd.n512 240.244
R5666 gnd.n7114 gnd.n508 240.244
R5667 gnd.n7120 gnd.n508 240.244
R5668 gnd.n7120 gnd.n506 240.244
R5669 gnd.n7124 gnd.n506 240.244
R5670 gnd.n7124 gnd.n502 240.244
R5671 gnd.n7130 gnd.n502 240.244
R5672 gnd.n7130 gnd.n500 240.244
R5673 gnd.n7134 gnd.n500 240.244
R5674 gnd.n7134 gnd.n496 240.244
R5675 gnd.n7140 gnd.n496 240.244
R5676 gnd.n7140 gnd.n494 240.244
R5677 gnd.n7144 gnd.n494 240.244
R5678 gnd.n7144 gnd.n490 240.244
R5679 gnd.n7150 gnd.n490 240.244
R5680 gnd.n7150 gnd.n488 240.244
R5681 gnd.n7154 gnd.n488 240.244
R5682 gnd.n7154 gnd.n484 240.244
R5683 gnd.n7160 gnd.n484 240.244
R5684 gnd.n7160 gnd.n482 240.244
R5685 gnd.n7164 gnd.n482 240.244
R5686 gnd.n7164 gnd.n478 240.244
R5687 gnd.n7170 gnd.n478 240.244
R5688 gnd.n7170 gnd.n476 240.244
R5689 gnd.n7174 gnd.n476 240.244
R5690 gnd.n7174 gnd.n472 240.244
R5691 gnd.n7180 gnd.n472 240.244
R5692 gnd.n7180 gnd.n470 240.244
R5693 gnd.n7184 gnd.n470 240.244
R5694 gnd.n7184 gnd.n466 240.244
R5695 gnd.n7190 gnd.n466 240.244
R5696 gnd.n7190 gnd.n464 240.244
R5697 gnd.n7194 gnd.n464 240.244
R5698 gnd.n7194 gnd.n460 240.244
R5699 gnd.n7200 gnd.n460 240.244
R5700 gnd.n7200 gnd.n458 240.244
R5701 gnd.n7204 gnd.n458 240.244
R5702 gnd.n7204 gnd.n454 240.244
R5703 gnd.n7210 gnd.n454 240.244
R5704 gnd.n7210 gnd.n452 240.244
R5705 gnd.n7214 gnd.n452 240.244
R5706 gnd.n7214 gnd.n448 240.244
R5707 gnd.n7220 gnd.n448 240.244
R5708 gnd.n7220 gnd.n446 240.244
R5709 gnd.n7224 gnd.n446 240.244
R5710 gnd.n7224 gnd.n442 240.244
R5711 gnd.n7230 gnd.n442 240.244
R5712 gnd.n7230 gnd.n440 240.244
R5713 gnd.n7234 gnd.n440 240.244
R5714 gnd.n7234 gnd.n436 240.244
R5715 gnd.n7240 gnd.n436 240.244
R5716 gnd.n7240 gnd.n434 240.244
R5717 gnd.n7244 gnd.n434 240.244
R5718 gnd.n7244 gnd.n430 240.244
R5719 gnd.n7250 gnd.n430 240.244
R5720 gnd.n7250 gnd.n428 240.244
R5721 gnd.n7254 gnd.n428 240.244
R5722 gnd.n7254 gnd.n424 240.244
R5723 gnd.n7260 gnd.n424 240.244
R5724 gnd.n7260 gnd.n422 240.244
R5725 gnd.n7264 gnd.n422 240.244
R5726 gnd.n7264 gnd.n418 240.244
R5727 gnd.n7270 gnd.n418 240.244
R5728 gnd.n7270 gnd.n416 240.244
R5729 gnd.n7274 gnd.n416 240.244
R5730 gnd.n7274 gnd.n412 240.244
R5731 gnd.n7280 gnd.n412 240.244
R5732 gnd.n7280 gnd.n410 240.244
R5733 gnd.n7284 gnd.n410 240.244
R5734 gnd.n7284 gnd.n406 240.244
R5735 gnd.n7292 gnd.n406 240.244
R5736 gnd.n7292 gnd.n404 240.244
R5737 gnd.n7296 gnd.n404 240.244
R5738 gnd.n7297 gnd.n7296 240.244
R5739 gnd.n2792 gnd.n2791 240.244
R5740 gnd.n2793 gnd.n2792 240.244
R5741 gnd.n2793 gnd.n2780 240.244
R5742 gnd.n2817 gnd.n2780 240.244
R5743 gnd.n2817 gnd.n2781 240.244
R5744 gnd.n2813 gnd.n2781 240.244
R5745 gnd.n2813 gnd.n2812 240.244
R5746 gnd.n2812 gnd.n2811 240.244
R5747 gnd.n2811 gnd.n2801 240.244
R5748 gnd.n2807 gnd.n2801 240.244
R5749 gnd.n2807 gnd.n2639 240.244
R5750 gnd.n2862 gnd.n2639 240.244
R5751 gnd.n2862 gnd.n2637 240.244
R5752 gnd.n2867 gnd.n2637 240.244
R5753 gnd.n2868 gnd.n2867 240.244
R5754 gnd.n2868 gnd.n2634 240.244
R5755 gnd.n2876 gnd.n2634 240.244
R5756 gnd.n2876 gnd.n2635 240.244
R5757 gnd.n2635 gnd.n2594 240.244
R5758 gnd.n2941 gnd.n2594 240.244
R5759 gnd.n2942 gnd.n2941 240.244
R5760 gnd.n2943 gnd.n2942 240.244
R5761 gnd.n2943 gnd.n2591 240.244
R5762 gnd.n2949 gnd.n2591 240.244
R5763 gnd.n2950 gnd.n2949 240.244
R5764 gnd.n2951 gnd.n2950 240.244
R5765 gnd.n2951 gnd.n2586 240.244
R5766 gnd.n2977 gnd.n2586 240.244
R5767 gnd.n2977 gnd.n2587 240.244
R5768 gnd.n2973 gnd.n2587 240.244
R5769 gnd.n2973 gnd.n2972 240.244
R5770 gnd.n2972 gnd.n2971 240.244
R5771 gnd.n2971 gnd.n2959 240.244
R5772 gnd.n2967 gnd.n2959 240.244
R5773 gnd.n2967 gnd.n2565 240.244
R5774 gnd.n3038 gnd.n2565 240.244
R5775 gnd.n3039 gnd.n3038 240.244
R5776 gnd.n3040 gnd.n3039 240.244
R5777 gnd.n3040 gnd.n2561 240.244
R5778 gnd.n3046 gnd.n2561 240.244
R5779 gnd.n3047 gnd.n3046 240.244
R5780 gnd.n3048 gnd.n3047 240.244
R5781 gnd.n3048 gnd.n2557 240.244
R5782 gnd.n3055 gnd.n2557 240.244
R5783 gnd.n3056 gnd.n3055 240.244
R5784 gnd.n3059 gnd.n3056 240.244
R5785 gnd.n3059 gnd.n2552 240.244
R5786 gnd.n3067 gnd.n2552 240.244
R5787 gnd.n3067 gnd.n2553 240.244
R5788 gnd.n2553 gnd.n2326 240.244
R5789 gnd.n3155 gnd.n2326 240.244
R5790 gnd.n3155 gnd.n2321 240.244
R5791 gnd.n3163 gnd.n2321 240.244
R5792 gnd.n3163 gnd.n2322 240.244
R5793 gnd.n2322 gnd.n2301 240.244
R5794 gnd.n3185 gnd.n2301 240.244
R5795 gnd.n3185 gnd.n2296 240.244
R5796 gnd.n3193 gnd.n2296 240.244
R5797 gnd.n3193 gnd.n2297 240.244
R5798 gnd.n2297 gnd.n2276 240.244
R5799 gnd.n3215 gnd.n2276 240.244
R5800 gnd.n3215 gnd.n2271 240.244
R5801 gnd.n3233 gnd.n2271 240.244
R5802 gnd.n3233 gnd.n2272 240.244
R5803 gnd.n3229 gnd.n2272 240.244
R5804 gnd.n3229 gnd.n3228 240.244
R5805 gnd.n3228 gnd.n3226 240.244
R5806 gnd.n3226 gnd.n2182 240.244
R5807 gnd.n3290 gnd.n2182 240.244
R5808 gnd.n3290 gnd.n2177 240.244
R5809 gnd.n3298 gnd.n2177 240.244
R5810 gnd.n3298 gnd.n2178 240.244
R5811 gnd.n2178 gnd.n2156 240.244
R5812 gnd.n3352 gnd.n2156 240.244
R5813 gnd.n3352 gnd.n2152 240.244
R5814 gnd.n3358 gnd.n2152 240.244
R5815 gnd.n3358 gnd.n2138 240.244
R5816 gnd.n3379 gnd.n2138 240.244
R5817 gnd.n3379 gnd.n2133 240.244
R5818 gnd.n3387 gnd.n2133 240.244
R5819 gnd.n3387 gnd.n2134 240.244
R5820 gnd.n2134 gnd.n2105 240.244
R5821 gnd.n3430 gnd.n2105 240.244
R5822 gnd.n3430 gnd.n2101 240.244
R5823 gnd.n3436 gnd.n2101 240.244
R5824 gnd.n3436 gnd.n2082 240.244
R5825 gnd.n3470 gnd.n2082 240.244
R5826 gnd.n3470 gnd.n2078 240.244
R5827 gnd.n3476 gnd.n2078 240.244
R5828 gnd.n3476 gnd.n2060 240.244
R5829 gnd.n3526 gnd.n2060 240.244
R5830 gnd.n3526 gnd.n2056 240.244
R5831 gnd.n3532 gnd.n2056 240.244
R5832 gnd.n3532 gnd.n2041 240.244
R5833 gnd.n3551 gnd.n2041 240.244
R5834 gnd.n3551 gnd.n2037 240.244
R5835 gnd.n3557 gnd.n2037 240.244
R5836 gnd.n3557 gnd.n2021 240.244
R5837 gnd.n3611 gnd.n2021 240.244
R5838 gnd.n3611 gnd.n2017 240.244
R5839 gnd.n3617 gnd.n2017 240.244
R5840 gnd.n3617 gnd.n1999 240.244
R5841 gnd.n3640 gnd.n1999 240.244
R5842 gnd.n3640 gnd.n1994 240.244
R5843 gnd.n3648 gnd.n1994 240.244
R5844 gnd.n3648 gnd.n1995 240.244
R5845 gnd.n1995 gnd.n1971 240.244
R5846 gnd.n3685 gnd.n1971 240.244
R5847 gnd.n3685 gnd.n1966 240.244
R5848 gnd.n3697 gnd.n1966 240.244
R5849 gnd.n3697 gnd.n1967 240.244
R5850 gnd.n3693 gnd.n1967 240.244
R5851 gnd.n3693 gnd.n1892 240.244
R5852 gnd.n3984 gnd.n1892 240.244
R5853 gnd.n3984 gnd.n1893 240.244
R5854 gnd.n3980 gnd.n1893 240.244
R5855 gnd.n3980 gnd.n1899 240.244
R5856 gnd.n3973 gnd.n1899 240.244
R5857 gnd.n3973 gnd.n1903 240.244
R5858 gnd.n3969 gnd.n1903 240.244
R5859 gnd.n3969 gnd.n1909 240.244
R5860 gnd.n3962 gnd.n1909 240.244
R5861 gnd.n3962 gnd.n1915 240.244
R5862 gnd.n3958 gnd.n1915 240.244
R5863 gnd.n3958 gnd.n1921 240.244
R5864 gnd.n3951 gnd.n1921 240.244
R5865 gnd.n3951 gnd.n1927 240.244
R5866 gnd.n3947 gnd.n1927 240.244
R5867 gnd.n3947 gnd.n1933 240.244
R5868 gnd.n3940 gnd.n1933 240.244
R5869 gnd.n3940 gnd.n1582 240.244
R5870 gnd.n4560 gnd.n1582 240.244
R5871 gnd.n4560 gnd.n1583 240.244
R5872 gnd.n4556 gnd.n1583 240.244
R5873 gnd.n4556 gnd.n1589 240.244
R5874 gnd.n4552 gnd.n1589 240.244
R5875 gnd.n4552 gnd.n1592 240.244
R5876 gnd.n4548 gnd.n1592 240.244
R5877 gnd.n4548 gnd.n1598 240.244
R5878 gnd.n1774 gnd.n1598 240.244
R5879 gnd.n1780 gnd.n1774 240.244
R5880 gnd.n1781 gnd.n1780 240.244
R5881 gnd.n1782 gnd.n1781 240.244
R5882 gnd.n1782 gnd.n1769 240.244
R5883 gnd.n1799 gnd.n1769 240.244
R5884 gnd.n1799 gnd.n1770 240.244
R5885 gnd.n1795 gnd.n1770 240.244
R5886 gnd.n1795 gnd.n1794 240.244
R5887 gnd.n1794 gnd.n1753 240.244
R5888 gnd.n4393 gnd.n1753 240.244
R5889 gnd.n4394 gnd.n4393 240.244
R5890 gnd.n4395 gnd.n4394 240.244
R5891 gnd.n4395 gnd.n1749 240.244
R5892 gnd.n4401 gnd.n1749 240.244
R5893 gnd.n4402 gnd.n4401 240.244
R5894 gnd.n4403 gnd.n4402 240.244
R5895 gnd.n4403 gnd.n1744 240.244
R5896 gnd.n4413 gnd.n1744 240.244
R5897 gnd.n4413 gnd.n1745 240.244
R5898 gnd.n1745 gnd.n1736 240.244
R5899 gnd.n4458 gnd.n1736 240.244
R5900 gnd.n4459 gnd.n4458 240.244
R5901 gnd.n4459 gnd.n1733 240.244
R5902 gnd.n4469 gnd.n1733 240.244
R5903 gnd.n4469 gnd.n1734 240.244
R5904 gnd.n4464 gnd.n1734 240.244
R5905 gnd.n4464 gnd.n382 240.244
R5906 gnd.n7322 gnd.n382 240.244
R5907 gnd.n7322 gnd.n383 240.244
R5908 gnd.n7317 gnd.n383 240.244
R5909 gnd.n7317 gnd.n7316 240.244
R5910 gnd.n7316 gnd.n7315 240.244
R5911 gnd.n7315 gnd.n387 240.244
R5912 gnd.n7311 gnd.n387 240.244
R5913 gnd.n7311 gnd.n7310 240.244
R5914 gnd.n7310 gnd.n7309 240.244
R5915 gnd.n7309 gnd.n393 240.244
R5916 gnd.n7305 gnd.n393 240.244
R5917 gnd.n7305 gnd.n7304 240.244
R5918 gnd.n7304 gnd.n7303 240.244
R5919 gnd.n7303 gnd.n399 240.244
R5920 gnd.n6630 gnd.n802 240.244
R5921 gnd.n6626 gnd.n802 240.244
R5922 gnd.n6626 gnd.n807 240.244
R5923 gnd.n6622 gnd.n807 240.244
R5924 gnd.n6622 gnd.n809 240.244
R5925 gnd.n6618 gnd.n809 240.244
R5926 gnd.n6618 gnd.n815 240.244
R5927 gnd.n6614 gnd.n815 240.244
R5928 gnd.n6614 gnd.n817 240.244
R5929 gnd.n6610 gnd.n817 240.244
R5930 gnd.n6610 gnd.n823 240.244
R5931 gnd.n6606 gnd.n823 240.244
R5932 gnd.n6606 gnd.n825 240.244
R5933 gnd.n6602 gnd.n825 240.244
R5934 gnd.n6602 gnd.n831 240.244
R5935 gnd.n6598 gnd.n831 240.244
R5936 gnd.n6598 gnd.n833 240.244
R5937 gnd.n6594 gnd.n833 240.244
R5938 gnd.n6594 gnd.n839 240.244
R5939 gnd.n6590 gnd.n839 240.244
R5940 gnd.n6590 gnd.n841 240.244
R5941 gnd.n6586 gnd.n841 240.244
R5942 gnd.n6586 gnd.n847 240.244
R5943 gnd.n6582 gnd.n847 240.244
R5944 gnd.n6582 gnd.n849 240.244
R5945 gnd.n6578 gnd.n849 240.244
R5946 gnd.n6578 gnd.n855 240.244
R5947 gnd.n6574 gnd.n855 240.244
R5948 gnd.n6574 gnd.n857 240.244
R5949 gnd.n6570 gnd.n857 240.244
R5950 gnd.n6570 gnd.n863 240.244
R5951 gnd.n6566 gnd.n863 240.244
R5952 gnd.n6566 gnd.n865 240.244
R5953 gnd.n6562 gnd.n865 240.244
R5954 gnd.n6562 gnd.n871 240.244
R5955 gnd.n6558 gnd.n871 240.244
R5956 gnd.n6558 gnd.n873 240.244
R5957 gnd.n6554 gnd.n873 240.244
R5958 gnd.n6554 gnd.n879 240.244
R5959 gnd.n6550 gnd.n879 240.244
R5960 gnd.n6550 gnd.n881 240.244
R5961 gnd.n6546 gnd.n881 240.244
R5962 gnd.n6546 gnd.n887 240.244
R5963 gnd.n6542 gnd.n887 240.244
R5964 gnd.n6542 gnd.n889 240.244
R5965 gnd.n6538 gnd.n889 240.244
R5966 gnd.n6538 gnd.n895 240.244
R5967 gnd.n6534 gnd.n895 240.244
R5968 gnd.n6534 gnd.n897 240.244
R5969 gnd.n6530 gnd.n897 240.244
R5970 gnd.n6530 gnd.n903 240.244
R5971 gnd.n6526 gnd.n903 240.244
R5972 gnd.n6526 gnd.n905 240.244
R5973 gnd.n6522 gnd.n905 240.244
R5974 gnd.n6522 gnd.n911 240.244
R5975 gnd.n6518 gnd.n911 240.244
R5976 gnd.n6518 gnd.n913 240.244
R5977 gnd.n6514 gnd.n913 240.244
R5978 gnd.n6514 gnd.n919 240.244
R5979 gnd.n6510 gnd.n919 240.244
R5980 gnd.n6510 gnd.n921 240.244
R5981 gnd.n6506 gnd.n921 240.244
R5982 gnd.n6506 gnd.n927 240.244
R5983 gnd.n6502 gnd.n927 240.244
R5984 gnd.n6502 gnd.n929 240.244
R5985 gnd.n6498 gnd.n929 240.244
R5986 gnd.n6498 gnd.n935 240.244
R5987 gnd.n6494 gnd.n935 240.244
R5988 gnd.n6494 gnd.n937 240.244
R5989 gnd.n6490 gnd.n937 240.244
R5990 gnd.n6490 gnd.n943 240.244
R5991 gnd.n6486 gnd.n943 240.244
R5992 gnd.n6486 gnd.n945 240.244
R5993 gnd.n6482 gnd.n945 240.244
R5994 gnd.n6482 gnd.n951 240.244
R5995 gnd.n6478 gnd.n951 240.244
R5996 gnd.n6478 gnd.n953 240.244
R5997 gnd.n6474 gnd.n953 240.244
R5998 gnd.n6474 gnd.n959 240.244
R5999 gnd.n6470 gnd.n959 240.244
R6000 gnd.n6470 gnd.n961 240.244
R6001 gnd.n6466 gnd.n961 240.244
R6002 gnd.n6466 gnd.n967 240.244
R6003 gnd.n2785 gnd.n967 240.244
R6004 gnd.n3143 gnd.n2336 240.244
R6005 gnd.n2336 gnd.n2317 240.244
R6006 gnd.n3166 gnd.n2317 240.244
R6007 gnd.n3166 gnd.n2310 240.244
R6008 gnd.n3173 gnd.n2310 240.244
R6009 gnd.n3173 gnd.n2312 240.244
R6010 gnd.n2312 gnd.n2292 240.244
R6011 gnd.n3196 gnd.n2292 240.244
R6012 gnd.n3196 gnd.n2286 240.244
R6013 gnd.n3203 gnd.n2286 240.244
R6014 gnd.n3203 gnd.n2287 240.244
R6015 gnd.n2287 gnd.n2267 240.244
R6016 gnd.n3236 gnd.n2267 240.244
R6017 gnd.n3236 gnd.n2261 240.244
R6018 gnd.n3243 gnd.n2261 240.244
R6019 gnd.n3243 gnd.n2262 240.244
R6020 gnd.n2262 gnd.n1494 240.244
R6021 gnd.n4661 gnd.n1494 240.244
R6022 gnd.n4661 gnd.n1495 240.244
R6023 gnd.n1500 gnd.n1495 240.244
R6024 gnd.n1501 gnd.n1500 240.244
R6025 gnd.n1502 gnd.n1501 240.244
R6026 gnd.n3328 gnd.n1502 240.244
R6027 gnd.n3328 gnd.n1505 240.244
R6028 gnd.n1506 gnd.n1505 240.244
R6029 gnd.n1507 gnd.n1506 240.244
R6030 gnd.n3308 gnd.n1507 240.244
R6031 gnd.n3308 gnd.n1510 240.244
R6032 gnd.n1511 gnd.n1510 240.244
R6033 gnd.n1512 gnd.n1511 240.244
R6034 gnd.n3398 gnd.n1512 240.244
R6035 gnd.n3398 gnd.n1515 240.244
R6036 gnd.n1516 gnd.n1515 240.244
R6037 gnd.n1517 gnd.n1516 240.244
R6038 gnd.n3410 gnd.n1517 240.244
R6039 gnd.n3410 gnd.n1520 240.244
R6040 gnd.n1521 gnd.n1520 240.244
R6041 gnd.n1522 gnd.n1521 240.244
R6042 gnd.n3449 gnd.n1522 240.244
R6043 gnd.n3449 gnd.n1525 240.244
R6044 gnd.n1526 gnd.n1525 240.244
R6045 gnd.n1527 gnd.n1526 240.244
R6046 gnd.n3490 gnd.n1527 240.244
R6047 gnd.n3490 gnd.n1530 240.244
R6048 gnd.n1531 gnd.n1530 240.244
R6049 gnd.n1532 gnd.n1531 240.244
R6050 gnd.n3560 gnd.n1532 240.244
R6051 gnd.n3560 gnd.n1535 240.244
R6052 gnd.n1536 gnd.n1535 240.244
R6053 gnd.n1537 gnd.n1536 240.244
R6054 gnd.n3619 gnd.n1537 240.244
R6055 gnd.n3619 gnd.n1540 240.244
R6056 gnd.n1541 gnd.n1540 240.244
R6057 gnd.n1542 gnd.n1541 240.244
R6058 gnd.n3650 gnd.n1542 240.244
R6059 gnd.n3650 gnd.n1545 240.244
R6060 gnd.n1546 gnd.n1545 240.244
R6061 gnd.n1547 gnd.n1546 240.244
R6062 gnd.n3682 gnd.n1547 240.244
R6063 gnd.n3682 gnd.n1550 240.244
R6064 gnd.n1551 gnd.n1550 240.244
R6065 gnd.n1552 gnd.n1551 240.244
R6066 gnd.n3715 gnd.n1552 240.244
R6067 gnd.n3715 gnd.n1555 240.244
R6068 gnd.n1556 gnd.n1555 240.244
R6069 gnd.n1557 gnd.n1556 240.244
R6070 gnd.n3977 gnd.n1557 240.244
R6071 gnd.n3977 gnd.n1560 240.244
R6072 gnd.n1561 gnd.n1560 240.244
R6073 gnd.n1562 gnd.n1561 240.244
R6074 gnd.n3966 gnd.n1562 240.244
R6075 gnd.n3966 gnd.n1565 240.244
R6076 gnd.n1566 gnd.n1565 240.244
R6077 gnd.n1567 gnd.n1566 240.244
R6078 gnd.n3955 gnd.n1567 240.244
R6079 gnd.n3955 gnd.n1570 240.244
R6080 gnd.n1571 gnd.n1570 240.244
R6081 gnd.n1572 gnd.n1571 240.244
R6082 gnd.n3944 gnd.n1572 240.244
R6083 gnd.n3944 gnd.n1575 240.244
R6084 gnd.n1576 gnd.n1575 240.244
R6085 gnd.n4563 gnd.n1576 240.244
R6086 gnd.n2340 gnd.n2339 240.244
R6087 gnd.n2531 gnd.n2340 240.244
R6088 gnd.n2344 gnd.n2343 240.244
R6089 gnd.n2534 gnd.n2345 240.244
R6090 gnd.n2462 gnd.n2461 240.244
R6091 gnd.n2536 gnd.n2471 240.244
R6092 gnd.n2539 gnd.n2472 240.244
R6093 gnd.n2482 gnd.n2481 240.244
R6094 gnd.n2541 gnd.n2492 240.244
R6095 gnd.n2544 gnd.n2493 240.244
R6096 gnd.n2503 gnd.n2502 240.244
R6097 gnd.n2546 gnd.n2513 240.244
R6098 gnd.n2550 gnd.n2514 240.244
R6099 gnd.n3072 gnd.n2529 240.244
R6100 gnd.n3145 gnd.n2328 240.244
R6101 gnd.n3152 gnd.n2328 240.244
R6102 gnd.n3152 gnd.n2319 240.244
R6103 gnd.n2319 gnd.n2307 240.244
R6104 gnd.n3175 gnd.n2307 240.244
R6105 gnd.n3175 gnd.n2302 240.244
R6106 gnd.n3182 gnd.n2302 240.244
R6107 gnd.n3182 gnd.n2294 240.244
R6108 gnd.n2294 gnd.n2283 240.244
R6109 gnd.n3205 gnd.n2283 240.244
R6110 gnd.n3205 gnd.n2278 240.244
R6111 gnd.n3212 gnd.n2278 240.244
R6112 gnd.n3212 gnd.n2269 240.244
R6113 gnd.n2269 gnd.n2258 240.244
R6114 gnd.n3245 gnd.n2258 240.244
R6115 gnd.n3245 gnd.n2253 240.244
R6116 gnd.n3255 gnd.n2253 240.244
R6117 gnd.n3255 gnd.n1492 240.244
R6118 gnd.n3249 gnd.n1492 240.244
R6119 gnd.n3249 gnd.n2174 240.244
R6120 gnd.n3301 gnd.n2174 240.244
R6121 gnd.n3301 gnd.n2169 240.244
R6122 gnd.n3327 gnd.n2169 240.244
R6123 gnd.n3327 gnd.n2165 240.244
R6124 gnd.n2165 gnd.n2157 240.244
R6125 gnd.n3306 gnd.n2157 240.244
R6126 gnd.n3310 gnd.n3306 240.244
R6127 gnd.n3311 gnd.n3310 240.244
R6128 gnd.n3311 gnd.n2140 240.244
R6129 gnd.n2140 gnd.n2122 240.244
R6130 gnd.n3400 gnd.n2122 240.244
R6131 gnd.n3401 gnd.n3400 240.244
R6132 gnd.n3403 gnd.n3401 240.244
R6133 gnd.n3403 gnd.n2118 240.244
R6134 gnd.n3409 gnd.n2118 240.244
R6135 gnd.n3409 gnd.n2092 240.244
R6136 gnd.n3457 gnd.n2092 240.244
R6137 gnd.n3457 gnd.n2093 240.244
R6138 gnd.n3451 gnd.n2093 240.244
R6139 gnd.n3451 gnd.n2070 240.244
R6140 gnd.n3515 gnd.n2070 240.244
R6141 gnd.n3515 gnd.n2062 240.244
R6142 gnd.n3492 gnd.n2062 240.244
R6143 gnd.n3493 gnd.n3492 240.244
R6144 gnd.n3494 gnd.n3493 240.244
R6145 gnd.n3494 gnd.n2043 240.244
R6146 gnd.n2043 gnd.n2036 240.244
R6147 gnd.n3497 gnd.n2036 240.244
R6148 gnd.n3500 gnd.n3497 240.244
R6149 gnd.n3500 gnd.n2014 240.244
R6150 gnd.n3621 gnd.n2014 240.244
R6151 gnd.n3621 gnd.n2008 240.244
R6152 gnd.n3628 gnd.n2008 240.244
R6153 gnd.n3628 gnd.n2009 240.244
R6154 gnd.n2009 gnd.n1985 240.244
R6155 gnd.n3660 gnd.n1985 240.244
R6156 gnd.n3660 gnd.n1980 240.244
R6157 gnd.n3673 gnd.n1980 240.244
R6158 gnd.n3673 gnd.n1973 240.244
R6159 gnd.n3665 gnd.n1973 240.244
R6160 gnd.n3666 gnd.n3665 240.244
R6161 gnd.n3666 gnd.n1950 240.244
R6162 gnd.n3717 gnd.n1950 240.244
R6163 gnd.n3717 gnd.n1891 240.244
R6164 gnd.n3723 gnd.n1891 240.244
R6165 gnd.n3724 gnd.n3723 240.244
R6166 gnd.n3724 gnd.n1900 240.244
R6167 gnd.n1901 gnd.n1900 240.244
R6168 gnd.n3731 gnd.n1901 240.244
R6169 gnd.n3732 gnd.n3731 240.244
R6170 gnd.n3732 gnd.n1912 240.244
R6171 gnd.n1913 gnd.n1912 240.244
R6172 gnd.n3739 gnd.n1913 240.244
R6173 gnd.n3740 gnd.n3739 240.244
R6174 gnd.n3740 gnd.n1924 240.244
R6175 gnd.n1925 gnd.n1924 240.244
R6176 gnd.n3747 gnd.n1925 240.244
R6177 gnd.n3748 gnd.n3747 240.244
R6178 gnd.n3748 gnd.n1936 240.244
R6179 gnd.n1937 gnd.n1936 240.244
R6180 gnd.n3934 gnd.n1937 240.244
R6181 gnd.n3934 gnd.n1580 240.244
R6182 gnd.n3821 gnd.n3820 240.244
R6183 gnd.n3824 gnd.n3823 240.244
R6184 gnd.n3832 gnd.n3831 240.244
R6185 gnd.n3835 gnd.n3834 240.244
R6186 gnd.n3847 gnd.n3846 240.244
R6187 gnd.n3850 gnd.n3849 240.244
R6188 gnd.n3866 gnd.n3865 240.244
R6189 gnd.n3869 gnd.n3868 240.244
R6190 gnd.n3885 gnd.n3884 240.244
R6191 gnd.n3888 gnd.n3887 240.244
R6192 gnd.n3904 gnd.n3903 240.244
R6193 gnd.n3906 gnd.n3762 240.244
R6194 gnd.n3923 gnd.n3762 240.244
R6195 gnd.n3926 gnd.n3925 240.244
R6196 gnd.n1474 gnd.n1473 240.132
R6197 gnd.n4003 gnd.n4002 240.132
R6198 gnd.n6633 gnd.n6632 225.874
R6199 gnd.n6633 gnd.n795 225.874
R6200 gnd.n6641 gnd.n795 225.874
R6201 gnd.n6642 gnd.n6641 225.874
R6202 gnd.n6643 gnd.n6642 225.874
R6203 gnd.n6643 gnd.n789 225.874
R6204 gnd.n6651 gnd.n789 225.874
R6205 gnd.n6652 gnd.n6651 225.874
R6206 gnd.n6653 gnd.n6652 225.874
R6207 gnd.n6653 gnd.n783 225.874
R6208 gnd.n6661 gnd.n783 225.874
R6209 gnd.n6662 gnd.n6661 225.874
R6210 gnd.n6663 gnd.n6662 225.874
R6211 gnd.n6663 gnd.n777 225.874
R6212 gnd.n6671 gnd.n777 225.874
R6213 gnd.n6672 gnd.n6671 225.874
R6214 gnd.n6673 gnd.n6672 225.874
R6215 gnd.n6673 gnd.n771 225.874
R6216 gnd.n6681 gnd.n771 225.874
R6217 gnd.n6682 gnd.n6681 225.874
R6218 gnd.n6683 gnd.n6682 225.874
R6219 gnd.n6683 gnd.n765 225.874
R6220 gnd.n6691 gnd.n765 225.874
R6221 gnd.n6692 gnd.n6691 225.874
R6222 gnd.n6693 gnd.n6692 225.874
R6223 gnd.n6693 gnd.n759 225.874
R6224 gnd.n6701 gnd.n759 225.874
R6225 gnd.n6702 gnd.n6701 225.874
R6226 gnd.n6703 gnd.n6702 225.874
R6227 gnd.n6703 gnd.n753 225.874
R6228 gnd.n6711 gnd.n753 225.874
R6229 gnd.n6712 gnd.n6711 225.874
R6230 gnd.n6713 gnd.n6712 225.874
R6231 gnd.n6713 gnd.n747 225.874
R6232 gnd.n6721 gnd.n747 225.874
R6233 gnd.n6722 gnd.n6721 225.874
R6234 gnd.n6723 gnd.n6722 225.874
R6235 gnd.n6723 gnd.n741 225.874
R6236 gnd.n6731 gnd.n741 225.874
R6237 gnd.n6732 gnd.n6731 225.874
R6238 gnd.n6733 gnd.n6732 225.874
R6239 gnd.n6733 gnd.n735 225.874
R6240 gnd.n6741 gnd.n735 225.874
R6241 gnd.n6742 gnd.n6741 225.874
R6242 gnd.n6743 gnd.n6742 225.874
R6243 gnd.n6743 gnd.n729 225.874
R6244 gnd.n6751 gnd.n729 225.874
R6245 gnd.n6752 gnd.n6751 225.874
R6246 gnd.n6753 gnd.n6752 225.874
R6247 gnd.n6753 gnd.n723 225.874
R6248 gnd.n6761 gnd.n723 225.874
R6249 gnd.n6762 gnd.n6761 225.874
R6250 gnd.n6763 gnd.n6762 225.874
R6251 gnd.n6763 gnd.n717 225.874
R6252 gnd.n6771 gnd.n717 225.874
R6253 gnd.n6772 gnd.n6771 225.874
R6254 gnd.n6773 gnd.n6772 225.874
R6255 gnd.n6773 gnd.n711 225.874
R6256 gnd.n6781 gnd.n711 225.874
R6257 gnd.n6782 gnd.n6781 225.874
R6258 gnd.n6783 gnd.n6782 225.874
R6259 gnd.n6783 gnd.n705 225.874
R6260 gnd.n6791 gnd.n705 225.874
R6261 gnd.n6792 gnd.n6791 225.874
R6262 gnd.n6793 gnd.n6792 225.874
R6263 gnd.n6793 gnd.n699 225.874
R6264 gnd.n6801 gnd.n699 225.874
R6265 gnd.n6802 gnd.n6801 225.874
R6266 gnd.n6803 gnd.n6802 225.874
R6267 gnd.n6803 gnd.n693 225.874
R6268 gnd.n6811 gnd.n693 225.874
R6269 gnd.n6812 gnd.n6811 225.874
R6270 gnd.n6813 gnd.n6812 225.874
R6271 gnd.n6813 gnd.n687 225.874
R6272 gnd.n6821 gnd.n687 225.874
R6273 gnd.n6822 gnd.n6821 225.874
R6274 gnd.n6823 gnd.n6822 225.874
R6275 gnd.n6823 gnd.n681 225.874
R6276 gnd.n6831 gnd.n681 225.874
R6277 gnd.n6832 gnd.n6831 225.874
R6278 gnd.n6833 gnd.n6832 225.874
R6279 gnd.n6833 gnd.n675 225.874
R6280 gnd.n6841 gnd.n675 225.874
R6281 gnd.n6842 gnd.n6841 225.874
R6282 gnd.n6843 gnd.n6842 225.874
R6283 gnd.n6843 gnd.n669 225.874
R6284 gnd.n6851 gnd.n669 225.874
R6285 gnd.n6852 gnd.n6851 225.874
R6286 gnd.n6853 gnd.n6852 225.874
R6287 gnd.n6853 gnd.n663 225.874
R6288 gnd.n6861 gnd.n663 225.874
R6289 gnd.n6862 gnd.n6861 225.874
R6290 gnd.n6863 gnd.n6862 225.874
R6291 gnd.n6863 gnd.n657 225.874
R6292 gnd.n6871 gnd.n657 225.874
R6293 gnd.n6872 gnd.n6871 225.874
R6294 gnd.n6873 gnd.n6872 225.874
R6295 gnd.n6873 gnd.n651 225.874
R6296 gnd.n6881 gnd.n651 225.874
R6297 gnd.n6882 gnd.n6881 225.874
R6298 gnd.n6883 gnd.n6882 225.874
R6299 gnd.n6883 gnd.n645 225.874
R6300 gnd.n6891 gnd.n645 225.874
R6301 gnd.n6892 gnd.n6891 225.874
R6302 gnd.n6893 gnd.n6892 225.874
R6303 gnd.n6893 gnd.n639 225.874
R6304 gnd.n6901 gnd.n639 225.874
R6305 gnd.n6902 gnd.n6901 225.874
R6306 gnd.n6903 gnd.n6902 225.874
R6307 gnd.n6903 gnd.n633 225.874
R6308 gnd.n6911 gnd.n633 225.874
R6309 gnd.n6912 gnd.n6911 225.874
R6310 gnd.n6913 gnd.n6912 225.874
R6311 gnd.n6913 gnd.n627 225.874
R6312 gnd.n6921 gnd.n627 225.874
R6313 gnd.n6922 gnd.n6921 225.874
R6314 gnd.n6923 gnd.n6922 225.874
R6315 gnd.n6923 gnd.n621 225.874
R6316 gnd.n6931 gnd.n621 225.874
R6317 gnd.n6932 gnd.n6931 225.874
R6318 gnd.n6933 gnd.n6932 225.874
R6319 gnd.n6933 gnd.n615 225.874
R6320 gnd.n6941 gnd.n615 225.874
R6321 gnd.n6942 gnd.n6941 225.874
R6322 gnd.n6943 gnd.n6942 225.874
R6323 gnd.n6943 gnd.n609 225.874
R6324 gnd.n6951 gnd.n609 225.874
R6325 gnd.n6952 gnd.n6951 225.874
R6326 gnd.n6953 gnd.n6952 225.874
R6327 gnd.n6953 gnd.n603 225.874
R6328 gnd.n6961 gnd.n603 225.874
R6329 gnd.n6962 gnd.n6961 225.874
R6330 gnd.n6963 gnd.n6962 225.874
R6331 gnd.n6963 gnd.n597 225.874
R6332 gnd.n6971 gnd.n597 225.874
R6333 gnd.n6972 gnd.n6971 225.874
R6334 gnd.n6973 gnd.n6972 225.874
R6335 gnd.n6973 gnd.n591 225.874
R6336 gnd.n6981 gnd.n591 225.874
R6337 gnd.n6982 gnd.n6981 225.874
R6338 gnd.n6983 gnd.n6982 225.874
R6339 gnd.n6983 gnd.n585 225.874
R6340 gnd.n6991 gnd.n585 225.874
R6341 gnd.n6992 gnd.n6991 225.874
R6342 gnd.n6993 gnd.n6992 225.874
R6343 gnd.n6993 gnd.n579 225.874
R6344 gnd.n7001 gnd.n579 225.874
R6345 gnd.n7002 gnd.n7001 225.874
R6346 gnd.n7003 gnd.n7002 225.874
R6347 gnd.n7003 gnd.n573 225.874
R6348 gnd.n7011 gnd.n573 225.874
R6349 gnd.n7012 gnd.n7011 225.874
R6350 gnd.n7013 gnd.n7012 225.874
R6351 gnd.n7013 gnd.n567 225.874
R6352 gnd.n7021 gnd.n567 225.874
R6353 gnd.n7022 gnd.n7021 225.874
R6354 gnd.n7023 gnd.n7022 225.874
R6355 gnd.n7023 gnd.n561 225.874
R6356 gnd.n7031 gnd.n561 225.874
R6357 gnd.n7032 gnd.n7031 225.874
R6358 gnd.n7033 gnd.n7032 225.874
R6359 gnd.n7033 gnd.n555 225.874
R6360 gnd.n7041 gnd.n555 225.874
R6361 gnd.n7042 gnd.n7041 225.874
R6362 gnd.n7043 gnd.n7042 225.874
R6363 gnd.n7043 gnd.n549 225.874
R6364 gnd.n7051 gnd.n549 225.874
R6365 gnd.n7052 gnd.n7051 225.874
R6366 gnd.n7053 gnd.n7052 225.874
R6367 gnd.n7053 gnd.n543 225.874
R6368 gnd.n7061 gnd.n543 225.874
R6369 gnd.n7062 gnd.n7061 225.874
R6370 gnd.n7063 gnd.n7062 225.874
R6371 gnd.n7063 gnd.n537 225.874
R6372 gnd.n7071 gnd.n537 225.874
R6373 gnd.n7072 gnd.n7071 225.874
R6374 gnd.n7073 gnd.n7072 225.874
R6375 gnd.n7073 gnd.n531 225.874
R6376 gnd.n7081 gnd.n531 225.874
R6377 gnd.n7082 gnd.n7081 225.874
R6378 gnd.n7083 gnd.n7082 225.874
R6379 gnd.n5493 gnd.t87 224.174
R6380 gnd.n5121 gnd.t82 224.174
R6381 gnd.n4244 gnd.n4243 199.319
R6382 gnd.n4245 gnd.n4244 199.319
R6383 gnd.n1427 gnd.n1426 199.319
R6384 gnd.n2382 gnd.n1427 199.319
R6385 gnd.n1475 gnd.n1472 186.49
R6386 gnd.n4004 gnd.n4001 186.49
R6387 gnd.n6289 gnd.n6288 185
R6388 gnd.n6287 gnd.n6286 185
R6389 gnd.n6266 gnd.n6265 185
R6390 gnd.n6281 gnd.n6280 185
R6391 gnd.n6279 gnd.n6278 185
R6392 gnd.n6270 gnd.n6269 185
R6393 gnd.n6273 gnd.n6272 185
R6394 gnd.n6257 gnd.n6256 185
R6395 gnd.n6255 gnd.n6254 185
R6396 gnd.n6234 gnd.n6233 185
R6397 gnd.n6249 gnd.n6248 185
R6398 gnd.n6247 gnd.n6246 185
R6399 gnd.n6238 gnd.n6237 185
R6400 gnd.n6241 gnd.n6240 185
R6401 gnd.n6225 gnd.n6224 185
R6402 gnd.n6223 gnd.n6222 185
R6403 gnd.n6202 gnd.n6201 185
R6404 gnd.n6217 gnd.n6216 185
R6405 gnd.n6215 gnd.n6214 185
R6406 gnd.n6206 gnd.n6205 185
R6407 gnd.n6209 gnd.n6208 185
R6408 gnd.n6194 gnd.n6193 185
R6409 gnd.n6192 gnd.n6191 185
R6410 gnd.n6171 gnd.n6170 185
R6411 gnd.n6186 gnd.n6185 185
R6412 gnd.n6184 gnd.n6183 185
R6413 gnd.n6175 gnd.n6174 185
R6414 gnd.n6178 gnd.n6177 185
R6415 gnd.n6162 gnd.n6161 185
R6416 gnd.n6160 gnd.n6159 185
R6417 gnd.n6139 gnd.n6138 185
R6418 gnd.n6154 gnd.n6153 185
R6419 gnd.n6152 gnd.n6151 185
R6420 gnd.n6143 gnd.n6142 185
R6421 gnd.n6146 gnd.n6145 185
R6422 gnd.n6130 gnd.n6129 185
R6423 gnd.n6128 gnd.n6127 185
R6424 gnd.n6107 gnd.n6106 185
R6425 gnd.n6122 gnd.n6121 185
R6426 gnd.n6120 gnd.n6119 185
R6427 gnd.n6111 gnd.n6110 185
R6428 gnd.n6114 gnd.n6113 185
R6429 gnd.n6098 gnd.n6097 185
R6430 gnd.n6096 gnd.n6095 185
R6431 gnd.n6075 gnd.n6074 185
R6432 gnd.n6090 gnd.n6089 185
R6433 gnd.n6088 gnd.n6087 185
R6434 gnd.n6079 gnd.n6078 185
R6435 gnd.n6082 gnd.n6081 185
R6436 gnd.n6067 gnd.n6066 185
R6437 gnd.n6065 gnd.n6064 185
R6438 gnd.n6044 gnd.n6043 185
R6439 gnd.n6059 gnd.n6058 185
R6440 gnd.n6057 gnd.n6056 185
R6441 gnd.n6048 gnd.n6047 185
R6442 gnd.n6051 gnd.n6050 185
R6443 gnd.n5494 gnd.t86 178.987
R6444 gnd.n5122 gnd.t83 178.987
R6445 gnd.n7091 gnd.n525 173.845
R6446 gnd.n7092 gnd.n7091 173.845
R6447 gnd.n7093 gnd.n7092 173.845
R6448 gnd.n7093 gnd.n519 173.845
R6449 gnd.n7101 gnd.n519 173.845
R6450 gnd.n7102 gnd.n7101 173.845
R6451 gnd.n7103 gnd.n7102 173.845
R6452 gnd.n7103 gnd.n513 173.845
R6453 gnd.n7111 gnd.n513 173.845
R6454 gnd.n7112 gnd.n7111 173.845
R6455 gnd.n7113 gnd.n7112 173.845
R6456 gnd.n7113 gnd.n507 173.845
R6457 gnd.n7121 gnd.n507 173.845
R6458 gnd.n7122 gnd.n7121 173.845
R6459 gnd.n7123 gnd.n7122 173.845
R6460 gnd.n7123 gnd.n501 173.845
R6461 gnd.n7131 gnd.n501 173.845
R6462 gnd.n7132 gnd.n7131 173.845
R6463 gnd.n7133 gnd.n7132 173.845
R6464 gnd.n7133 gnd.n495 173.845
R6465 gnd.n7141 gnd.n495 173.845
R6466 gnd.n7142 gnd.n7141 173.845
R6467 gnd.n7143 gnd.n7142 173.845
R6468 gnd.n7143 gnd.n489 173.845
R6469 gnd.n7151 gnd.n489 173.845
R6470 gnd.n7152 gnd.n7151 173.845
R6471 gnd.n7153 gnd.n7152 173.845
R6472 gnd.n7153 gnd.n483 173.845
R6473 gnd.n7161 gnd.n483 173.845
R6474 gnd.n7162 gnd.n7161 173.845
R6475 gnd.n7163 gnd.n7162 173.845
R6476 gnd.n7163 gnd.n477 173.845
R6477 gnd.n7171 gnd.n477 173.845
R6478 gnd.n7172 gnd.n7171 173.845
R6479 gnd.n7173 gnd.n7172 173.845
R6480 gnd.n7173 gnd.n471 173.845
R6481 gnd.n7181 gnd.n471 173.845
R6482 gnd.n7182 gnd.n7181 173.845
R6483 gnd.n7183 gnd.n7182 173.845
R6484 gnd.n7183 gnd.n465 173.845
R6485 gnd.n7191 gnd.n465 173.845
R6486 gnd.n7192 gnd.n7191 173.845
R6487 gnd.n7193 gnd.n7192 173.845
R6488 gnd.n7193 gnd.n459 173.845
R6489 gnd.n7201 gnd.n459 173.845
R6490 gnd.n7202 gnd.n7201 173.845
R6491 gnd.n7203 gnd.n7202 173.845
R6492 gnd.n7203 gnd.n453 173.845
R6493 gnd.n7211 gnd.n453 173.845
R6494 gnd.n7212 gnd.n7211 173.845
R6495 gnd.n7213 gnd.n7212 173.845
R6496 gnd.n7213 gnd.n447 173.845
R6497 gnd.n7221 gnd.n447 173.845
R6498 gnd.n7222 gnd.n7221 173.845
R6499 gnd.n7223 gnd.n7222 173.845
R6500 gnd.n7223 gnd.n441 173.845
R6501 gnd.n7231 gnd.n441 173.845
R6502 gnd.n7232 gnd.n7231 173.845
R6503 gnd.n7233 gnd.n7232 173.845
R6504 gnd.n7233 gnd.n435 173.845
R6505 gnd.n7241 gnd.n435 173.845
R6506 gnd.n7242 gnd.n7241 173.845
R6507 gnd.n7243 gnd.n7242 173.845
R6508 gnd.n7243 gnd.n429 173.845
R6509 gnd.n7251 gnd.n429 173.845
R6510 gnd.n7252 gnd.n7251 173.845
R6511 gnd.n7253 gnd.n7252 173.845
R6512 gnd.n7253 gnd.n423 173.845
R6513 gnd.n7261 gnd.n423 173.845
R6514 gnd.n7262 gnd.n7261 173.845
R6515 gnd.n7263 gnd.n7262 173.845
R6516 gnd.n7263 gnd.n417 173.845
R6517 gnd.n7271 gnd.n417 173.845
R6518 gnd.n7272 gnd.n7271 173.845
R6519 gnd.n7273 gnd.n7272 173.845
R6520 gnd.n7273 gnd.n411 173.845
R6521 gnd.n7281 gnd.n411 173.845
R6522 gnd.n7282 gnd.n7281 173.845
R6523 gnd.n7283 gnd.n7282 173.845
R6524 gnd.n7283 gnd.n405 173.845
R6525 gnd.n7293 gnd.n405 173.845
R6526 gnd.n7294 gnd.n7293 173.845
R6527 gnd.n7295 gnd.n7294 173.845
R6528 gnd.n1 gnd.t263 170.774
R6529 gnd.n7 gnd.t32 170.103
R6530 gnd.n6 gnd.t286 170.103
R6531 gnd.n5 gnd.t265 170.103
R6532 gnd.n4 gnd.t301 170.103
R6533 gnd.n3 gnd.t209 170.103
R6534 gnd.n2 gnd.t41 170.103
R6535 gnd.n1 gnd.t11 170.103
R6536 gnd.n4072 gnd.n4071 163.367
R6537 gnd.n4068 gnd.n4067 163.367
R6538 gnd.n4064 gnd.n4063 163.367
R6539 gnd.n4060 gnd.n4059 163.367
R6540 gnd.n4056 gnd.n4055 163.367
R6541 gnd.n4052 gnd.n4051 163.367
R6542 gnd.n4048 gnd.n4047 163.367
R6543 gnd.n4044 gnd.n4043 163.367
R6544 gnd.n4040 gnd.n4039 163.367
R6545 gnd.n4036 gnd.n4035 163.367
R6546 gnd.n4032 gnd.n4031 163.367
R6547 gnd.n4028 gnd.n4027 163.367
R6548 gnd.n4024 gnd.n4023 163.367
R6549 gnd.n4020 gnd.n4019 163.367
R6550 gnd.n4015 gnd.n4014 163.367
R6551 gnd.n4147 gnd.n1845 163.367
R6552 gnd.n4144 gnd.n4143 163.367
R6553 gnd.n4141 gnd.n1878 163.367
R6554 gnd.n4136 gnd.n4135 163.367
R6555 gnd.n4132 gnd.n4131 163.367
R6556 gnd.n4128 gnd.n4127 163.367
R6557 gnd.n4124 gnd.n4123 163.367
R6558 gnd.n4120 gnd.n4119 163.367
R6559 gnd.n4116 gnd.n4115 163.367
R6560 gnd.n4112 gnd.n4111 163.367
R6561 gnd.n4108 gnd.n4107 163.367
R6562 gnd.n4104 gnd.n4103 163.367
R6563 gnd.n4100 gnd.n4099 163.367
R6564 gnd.n4096 gnd.n4095 163.367
R6565 gnd.n4092 gnd.n4091 163.367
R6566 gnd.n4088 gnd.n4087 163.367
R6567 gnd.n4084 gnd.n4083 163.367
R6568 gnd.n3258 gnd.n1491 163.367
R6569 gnd.n3262 gnd.n1491 163.367
R6570 gnd.n3265 gnd.n3262 163.367
R6571 gnd.n3265 gnd.n2184 163.367
R6572 gnd.n3272 gnd.n2184 163.367
R6573 gnd.n3272 gnd.n2187 163.367
R6574 gnd.n3268 gnd.n2187 163.367
R6575 gnd.n3268 gnd.n2167 163.367
R6576 gnd.n3331 gnd.n2167 163.367
R6577 gnd.n3331 gnd.n2164 163.367
R6578 gnd.n3340 gnd.n2164 163.367
R6579 gnd.n3340 gnd.n2158 163.367
R6580 gnd.n3336 gnd.n2158 163.367
R6581 gnd.n3336 gnd.n2151 163.367
R6582 gnd.n2151 gnd.n2143 163.367
R6583 gnd.n3368 gnd.n2143 163.367
R6584 gnd.n3368 gnd.n2141 163.367
R6585 gnd.n3375 gnd.n2141 163.367
R6586 gnd.n3375 gnd.n2131 163.367
R6587 gnd.n2132 gnd.n2131 163.367
R6588 gnd.n2132 gnd.n2124 163.367
R6589 gnd.n2124 gnd.n2114 163.367
R6590 gnd.n3418 gnd.n2114 163.367
R6591 gnd.n3418 gnd.n2115 163.367
R6592 gnd.n2115 gnd.n2107 163.367
R6593 gnd.n3413 gnd.n2107 163.367
R6594 gnd.n3413 gnd.n2099 163.367
R6595 gnd.n3440 gnd.n2099 163.367
R6596 gnd.n3440 gnd.n2091 163.367
R6597 gnd.n3443 gnd.n2091 163.367
R6598 gnd.n3443 gnd.n2084 163.367
R6599 gnd.n3447 gnd.n2084 163.367
R6600 gnd.n3447 gnd.n2076 163.367
R6601 gnd.n3480 gnd.n2076 163.367
R6602 gnd.n3480 gnd.n2069 163.367
R6603 gnd.n3483 gnd.n2069 163.367
R6604 gnd.n3483 gnd.n2063 163.367
R6605 gnd.n3488 gnd.n2063 163.367
R6606 gnd.n3488 gnd.n2053 163.367
R6607 gnd.n2053 gnd.n2046 163.367
R6608 gnd.n3542 gnd.n2046 163.367
R6609 gnd.n3542 gnd.n2044 163.367
R6610 gnd.n3547 gnd.n2044 163.367
R6611 gnd.n3547 gnd.n2035 163.367
R6612 gnd.n2035 gnd.n2027 163.367
R6613 gnd.n3577 gnd.n2027 163.367
R6614 gnd.n3577 gnd.n2024 163.367
R6615 gnd.n3609 gnd.n2024 163.367
R6616 gnd.n3609 gnd.n2025 163.367
R6617 gnd.n3605 gnd.n2025 163.367
R6618 gnd.n3605 gnd.n3604 163.367
R6619 gnd.n3604 gnd.n2006 163.367
R6620 gnd.n2007 gnd.n2006 163.367
R6621 gnd.n2007 gnd.n2000 163.367
R6622 gnd.n3598 gnd.n2000 163.367
R6623 gnd.n3598 gnd.n1993 163.367
R6624 gnd.n3594 gnd.n1993 163.367
R6625 gnd.n3594 gnd.n1987 163.367
R6626 gnd.n3591 gnd.n1987 163.367
R6627 gnd.n3591 gnd.n1979 163.367
R6628 gnd.n3585 gnd.n1979 163.367
R6629 gnd.n3585 gnd.n1974 163.367
R6630 gnd.n3582 gnd.n1974 163.367
R6631 gnd.n3582 gnd.n1963 163.367
R6632 gnd.n1963 gnd.n1954 163.367
R6633 gnd.n3707 gnd.n1954 163.367
R6634 gnd.n3707 gnd.n1952 163.367
R6635 gnd.n3713 gnd.n1952 163.367
R6636 gnd.n3713 gnd.n1890 163.367
R6637 gnd.n1890 gnd.n1882 163.367
R6638 gnd.n4079 gnd.n1882 163.367
R6639 gnd.n1466 gnd.n1465 163.367
R6640 gnd.n4726 gnd.n1465 163.367
R6641 gnd.n4724 gnd.n4723 163.367
R6642 gnd.n4720 gnd.n4719 163.367
R6643 gnd.n4716 gnd.n4715 163.367
R6644 gnd.n4712 gnd.n4711 163.367
R6645 gnd.n4708 gnd.n4707 163.367
R6646 gnd.n4704 gnd.n4703 163.367
R6647 gnd.n4700 gnd.n4699 163.367
R6648 gnd.n4696 gnd.n4695 163.367
R6649 gnd.n4692 gnd.n4691 163.367
R6650 gnd.n4688 gnd.n4687 163.367
R6651 gnd.n4684 gnd.n4683 163.367
R6652 gnd.n4680 gnd.n4679 163.367
R6653 gnd.n4676 gnd.n4675 163.367
R6654 gnd.n4672 gnd.n4671 163.367
R6655 gnd.n4735 gnd.n1432 163.367
R6656 gnd.n2192 gnd.n2191 163.367
R6657 gnd.n2197 gnd.n2196 163.367
R6658 gnd.n2201 gnd.n2200 163.367
R6659 gnd.n2205 gnd.n2204 163.367
R6660 gnd.n2209 gnd.n2208 163.367
R6661 gnd.n2213 gnd.n2212 163.367
R6662 gnd.n2217 gnd.n2216 163.367
R6663 gnd.n2221 gnd.n2220 163.367
R6664 gnd.n2225 gnd.n2224 163.367
R6665 gnd.n2229 gnd.n2228 163.367
R6666 gnd.n2233 gnd.n2232 163.367
R6667 gnd.n2237 gnd.n2236 163.367
R6668 gnd.n2241 gnd.n2240 163.367
R6669 gnd.n2245 gnd.n2244 163.367
R6670 gnd.n2249 gnd.n2248 163.367
R6671 gnd.n4664 gnd.n1467 163.367
R6672 gnd.n4664 gnd.n1489 163.367
R6673 gnd.n2186 gnd.n1489 163.367
R6674 gnd.n3287 gnd.n2186 163.367
R6675 gnd.n3287 gnd.n3275 163.367
R6676 gnd.n3283 gnd.n3275 163.367
R6677 gnd.n3283 gnd.n3282 163.367
R6678 gnd.n3282 gnd.n3281 163.367
R6679 gnd.n3281 gnd.n2162 163.367
R6680 gnd.n3344 gnd.n2162 163.367
R6681 gnd.n3344 gnd.n2160 163.367
R6682 gnd.n3348 gnd.n2160 163.367
R6683 gnd.n3348 gnd.n2149 163.367
R6684 gnd.n3361 gnd.n2149 163.367
R6685 gnd.n3361 gnd.n2146 163.367
R6686 gnd.n3366 gnd.n2146 163.367
R6687 gnd.n3366 gnd.n2147 163.367
R6688 gnd.n2147 gnd.n2129 163.367
R6689 gnd.n3392 gnd.n2129 163.367
R6690 gnd.n3392 gnd.n2127 163.367
R6691 gnd.n3396 gnd.n2127 163.367
R6692 gnd.n3396 gnd.n2112 163.367
R6693 gnd.n3420 gnd.n2112 163.367
R6694 gnd.n3420 gnd.n2109 163.367
R6695 gnd.n3427 gnd.n2109 163.367
R6696 gnd.n3427 gnd.n2110 163.367
R6697 gnd.n3423 gnd.n2110 163.367
R6698 gnd.n3423 gnd.n2089 163.367
R6699 gnd.n3460 gnd.n2089 163.367
R6700 gnd.n3460 gnd.n2086 163.367
R6701 gnd.n3467 gnd.n2086 163.367
R6702 gnd.n3467 gnd.n2087 163.367
R6703 gnd.n3463 gnd.n2087 163.367
R6704 gnd.n3463 gnd.n2067 163.367
R6705 gnd.n3518 gnd.n2067 163.367
R6706 gnd.n3518 gnd.n2065 163.367
R6707 gnd.n3522 gnd.n2065 163.367
R6708 gnd.n3522 gnd.n2052 163.367
R6709 gnd.n3535 gnd.n2052 163.367
R6710 gnd.n3535 gnd.n2049 163.367
R6711 gnd.n3540 gnd.n2049 163.367
R6712 gnd.n3540 gnd.n2050 163.367
R6713 gnd.n2050 gnd.n2033 163.367
R6714 gnd.n3563 gnd.n2033 163.367
R6715 gnd.n3563 gnd.n2030 163.367
R6716 gnd.n3575 gnd.n2030 163.367
R6717 gnd.n3575 gnd.n2031 163.367
R6718 gnd.n2031 gnd.n2022 163.367
R6719 gnd.n3570 gnd.n2022 163.367
R6720 gnd.n3570 gnd.n3567 163.367
R6721 gnd.n3567 gnd.n2004 163.367
R6722 gnd.n3633 gnd.n2004 163.367
R6723 gnd.n3633 gnd.n2002 163.367
R6724 gnd.n3637 gnd.n2002 163.367
R6725 gnd.n3637 gnd.n1991 163.367
R6726 gnd.n3653 gnd.n1991 163.367
R6727 gnd.n3653 gnd.n1989 163.367
R6728 gnd.n3657 gnd.n1989 163.367
R6729 gnd.n3657 gnd.n1978 163.367
R6730 gnd.n3676 gnd.n1978 163.367
R6731 gnd.n3676 gnd.n1976 163.367
R6732 gnd.n3680 gnd.n1976 163.367
R6733 gnd.n3680 gnd.n1961 163.367
R6734 gnd.n3700 gnd.n1961 163.367
R6735 gnd.n3700 gnd.n1956 163.367
R6736 gnd.n3705 gnd.n1956 163.367
R6737 gnd.n3705 gnd.n1959 163.367
R6738 gnd.n1959 gnd.n1888 163.367
R6739 gnd.n3989 gnd.n1888 163.367
R6740 gnd.n3989 gnd.n1885 163.367
R6741 gnd.n4077 gnd.n1885 163.367
R6742 gnd.n4010 gnd.n4009 156.462
R6743 gnd.n6229 gnd.n6197 153.042
R6744 gnd.n6293 gnd.n6292 152.079
R6745 gnd.n6261 gnd.n6260 152.079
R6746 gnd.n6229 gnd.n6228 152.079
R6747 gnd.n1480 gnd.n1479 152
R6748 gnd.n1481 gnd.n1470 152
R6749 gnd.n1483 gnd.n1482 152
R6750 gnd.n1485 gnd.n1468 152
R6751 gnd.n1487 gnd.n1486 152
R6752 gnd.n4008 gnd.n3992 152
R6753 gnd.n4000 gnd.n3993 152
R6754 gnd.n3999 gnd.n3998 152
R6755 gnd.n3997 gnd.n3994 152
R6756 gnd.n3995 gnd.t99 150.546
R6757 gnd.t359 gnd.n6271 147.661
R6758 gnd.t236 gnd.n6239 147.661
R6759 gnd.t271 gnd.n6207 147.661
R6760 gnd.t222 gnd.n6176 147.661
R6761 gnd.t258 gnd.n6144 147.661
R6762 gnd.t277 gnd.n6112 147.661
R6763 gnd.t352 gnd.n6080 147.661
R6764 gnd.t253 gnd.n6049 147.661
R6765 gnd.n4146 gnd.n1844 143.351
R6766 gnd.n1447 gnd.n1431 143.351
R6767 gnd.n4734 gnd.n1431 143.351
R6768 gnd.n7295 gnd.n212 132.349
R6769 gnd.n4149 gnd.n4148 131.649
R6770 gnd.n4737 gnd.n4736 131.649
R6771 gnd.n1477 gnd.t157 130.484
R6772 gnd.n1486 gnd.t120 126.766
R6773 gnd.n1484 gnd.t77 126.766
R6774 gnd.n1470 gnd.t127 126.766
R6775 gnd.n1478 gnd.t194 126.766
R6776 gnd.n3996 gnd.t96 126.766
R6777 gnd.n3998 gnd.t169 126.766
R6778 gnd.n4007 gnd.t147 126.766
R6779 gnd.n4009 gnd.t185 126.766
R6780 gnd.n6288 gnd.n6287 104.615
R6781 gnd.n6287 gnd.n6265 104.615
R6782 gnd.n6280 gnd.n6265 104.615
R6783 gnd.n6280 gnd.n6279 104.615
R6784 gnd.n6279 gnd.n6269 104.615
R6785 gnd.n6272 gnd.n6269 104.615
R6786 gnd.n6256 gnd.n6255 104.615
R6787 gnd.n6255 gnd.n6233 104.615
R6788 gnd.n6248 gnd.n6233 104.615
R6789 gnd.n6248 gnd.n6247 104.615
R6790 gnd.n6247 gnd.n6237 104.615
R6791 gnd.n6240 gnd.n6237 104.615
R6792 gnd.n6224 gnd.n6223 104.615
R6793 gnd.n6223 gnd.n6201 104.615
R6794 gnd.n6216 gnd.n6201 104.615
R6795 gnd.n6216 gnd.n6215 104.615
R6796 gnd.n6215 gnd.n6205 104.615
R6797 gnd.n6208 gnd.n6205 104.615
R6798 gnd.n6193 gnd.n6192 104.615
R6799 gnd.n6192 gnd.n6170 104.615
R6800 gnd.n6185 gnd.n6170 104.615
R6801 gnd.n6185 gnd.n6184 104.615
R6802 gnd.n6184 gnd.n6174 104.615
R6803 gnd.n6177 gnd.n6174 104.615
R6804 gnd.n6161 gnd.n6160 104.615
R6805 gnd.n6160 gnd.n6138 104.615
R6806 gnd.n6153 gnd.n6138 104.615
R6807 gnd.n6153 gnd.n6152 104.615
R6808 gnd.n6152 gnd.n6142 104.615
R6809 gnd.n6145 gnd.n6142 104.615
R6810 gnd.n6129 gnd.n6128 104.615
R6811 gnd.n6128 gnd.n6106 104.615
R6812 gnd.n6121 gnd.n6106 104.615
R6813 gnd.n6121 gnd.n6120 104.615
R6814 gnd.n6120 gnd.n6110 104.615
R6815 gnd.n6113 gnd.n6110 104.615
R6816 gnd.n6097 gnd.n6096 104.615
R6817 gnd.n6096 gnd.n6074 104.615
R6818 gnd.n6089 gnd.n6074 104.615
R6819 gnd.n6089 gnd.n6088 104.615
R6820 gnd.n6088 gnd.n6078 104.615
R6821 gnd.n6081 gnd.n6078 104.615
R6822 gnd.n6066 gnd.n6065 104.615
R6823 gnd.n6065 gnd.n6043 104.615
R6824 gnd.n6058 gnd.n6043 104.615
R6825 gnd.n6058 gnd.n6057 104.615
R6826 gnd.n6057 gnd.n6047 104.615
R6827 gnd.n6050 gnd.n6047 104.615
R6828 gnd.n5643 gnd.t153 100.632
R6829 gnd.n5077 gnd.t180 100.632
R6830 gnd.n7549 gnd.n219 99.6594
R6831 gnd.n7547 gnd.n7546 99.6594
R6832 gnd.n7542 gnd.n226 99.6594
R6833 gnd.n7540 gnd.n7539 99.6594
R6834 gnd.n7535 gnd.n233 99.6594
R6835 gnd.n7533 gnd.n7532 99.6594
R6836 gnd.n7528 gnd.n240 99.6594
R6837 gnd.n7526 gnd.n7525 99.6594
R6838 gnd.n7518 gnd.n247 99.6594
R6839 gnd.n7516 gnd.n7515 99.6594
R6840 gnd.n7511 gnd.n254 99.6594
R6841 gnd.n7509 gnd.n7508 99.6594
R6842 gnd.n7504 gnd.n261 99.6594
R6843 gnd.n7502 gnd.n7501 99.6594
R6844 gnd.n7497 gnd.n268 99.6594
R6845 gnd.n7495 gnd.n7494 99.6594
R6846 gnd.n7490 gnd.n275 99.6594
R6847 gnd.n7488 gnd.n7487 99.6594
R6848 gnd.n285 gnd.n284 99.6594
R6849 gnd.n7479 gnd.n7478 99.6594
R6850 gnd.n7476 gnd.n7475 99.6594
R6851 gnd.n7471 gnd.n293 99.6594
R6852 gnd.n7469 gnd.n7468 99.6594
R6853 gnd.n7464 gnd.n300 99.6594
R6854 gnd.n7462 gnd.n7461 99.6594
R6855 gnd.n7457 gnd.n307 99.6594
R6856 gnd.n7455 gnd.n7454 99.6594
R6857 gnd.n7450 gnd.n316 99.6594
R6858 gnd.n7448 gnd.n7447 99.6594
R6859 gnd.n4178 gnd.n1604 99.6594
R6860 gnd.n4182 gnd.n4181 99.6594
R6861 gnd.n4189 gnd.n4188 99.6594
R6862 gnd.n4192 gnd.n4191 99.6594
R6863 gnd.n4199 gnd.n4198 99.6594
R6864 gnd.n4202 gnd.n4201 99.6594
R6865 gnd.n4209 gnd.n4208 99.6594
R6866 gnd.n4212 gnd.n4211 99.6594
R6867 gnd.n4222 gnd.n4221 99.6594
R6868 gnd.n4225 gnd.n4224 99.6594
R6869 gnd.n4232 gnd.n4231 99.6594
R6870 gnd.n4235 gnd.n4234 99.6594
R6871 gnd.n4243 gnd.n4242 99.6594
R6872 gnd.n4248 gnd.n4247 99.6594
R6873 gnd.n4255 gnd.n4254 99.6594
R6874 gnd.n4258 gnd.n4257 99.6594
R6875 gnd.n4265 gnd.n4264 99.6594
R6876 gnd.n4268 gnd.n4267 99.6594
R6877 gnd.n4277 gnd.n4276 99.6594
R6878 gnd.n4280 gnd.n4279 99.6594
R6879 gnd.n4287 gnd.n4286 99.6594
R6880 gnd.n4290 gnd.n4289 99.6594
R6881 gnd.n4297 gnd.n4296 99.6594
R6882 gnd.n4300 gnd.n4299 99.6594
R6883 gnd.n4307 gnd.n4306 99.6594
R6884 gnd.n4310 gnd.n4309 99.6594
R6885 gnd.n4318 gnd.n4317 99.6594
R6886 gnd.n4321 gnd.n4320 99.6594
R6887 gnd.n4780 gnd.n4779 99.6594
R6888 gnd.n4777 gnd.n4776 99.6594
R6889 gnd.n4772 gnd.n1390 99.6594
R6890 gnd.n4770 gnd.n4769 99.6594
R6891 gnd.n4765 gnd.n1397 99.6594
R6892 gnd.n4763 gnd.n4762 99.6594
R6893 gnd.n4758 gnd.n1404 99.6594
R6894 gnd.n4756 gnd.n4755 99.6594
R6895 gnd.n4750 gnd.n1413 99.6594
R6896 gnd.n4748 gnd.n4747 99.6594
R6897 gnd.n4743 gnd.n1420 99.6594
R6898 gnd.n4741 gnd.n4740 99.6594
R6899 gnd.n2383 gnd.n2382 99.6594
R6900 gnd.n2387 gnd.n2385 99.6594
R6901 gnd.n2393 gnd.n2377 99.6594
R6902 gnd.n2397 gnd.n2395 99.6594
R6903 gnd.n2403 gnd.n2373 99.6594
R6904 gnd.n2407 gnd.n2405 99.6594
R6905 gnd.n2413 gnd.n2367 99.6594
R6906 gnd.n2417 gnd.n2415 99.6594
R6907 gnd.n2423 gnd.n2363 99.6594
R6908 gnd.n2427 gnd.n2425 99.6594
R6909 gnd.n2433 gnd.n2359 99.6594
R6910 gnd.n2437 gnd.n2435 99.6594
R6911 gnd.n2443 gnd.n2355 99.6594
R6912 gnd.n2447 gnd.n2445 99.6594
R6913 gnd.n2453 gnd.n2351 99.6594
R6914 gnd.n2456 gnd.n2455 99.6594
R6915 gnd.n5045 gnd.n5044 99.6594
R6916 gnd.n5039 gnd.n1030 99.6594
R6917 gnd.n5036 gnd.n1031 99.6594
R6918 gnd.n5032 gnd.n1032 99.6594
R6919 gnd.n5028 gnd.n1033 99.6594
R6920 gnd.n5024 gnd.n1034 99.6594
R6921 gnd.n5020 gnd.n1035 99.6594
R6922 gnd.n5016 gnd.n1036 99.6594
R6923 gnd.n5012 gnd.n1037 99.6594
R6924 gnd.n5007 gnd.n1038 99.6594
R6925 gnd.n5003 gnd.n1039 99.6594
R6926 gnd.n4999 gnd.n1040 99.6594
R6927 gnd.n4995 gnd.n1041 99.6594
R6928 gnd.n4991 gnd.n1042 99.6594
R6929 gnd.n4987 gnd.n1043 99.6594
R6930 gnd.n4983 gnd.n1044 99.6594
R6931 gnd.n4979 gnd.n1045 99.6594
R6932 gnd.n4975 gnd.n1046 99.6594
R6933 gnd.n4971 gnd.n1047 99.6594
R6934 gnd.n4967 gnd.n1048 99.6594
R6935 gnd.n4963 gnd.n1049 99.6594
R6936 gnd.n4959 gnd.n1050 99.6594
R6937 gnd.n4955 gnd.n1051 99.6594
R6938 gnd.n4951 gnd.n1052 99.6594
R6939 gnd.n4947 gnd.n1053 99.6594
R6940 gnd.n4943 gnd.n1054 99.6594
R6941 gnd.n4939 gnd.n1055 99.6594
R6942 gnd.n4935 gnd.n1056 99.6594
R6943 gnd.n4931 gnd.n1057 99.6594
R6944 gnd.n6419 gnd.n5057 99.6594
R6945 gnd.n6417 gnd.n6416 99.6594
R6946 gnd.n6412 gnd.n5064 99.6594
R6947 gnd.n6410 gnd.n6409 99.6594
R6948 gnd.n6405 gnd.n5071 99.6594
R6949 gnd.n6403 gnd.n6402 99.6594
R6950 gnd.n6398 gnd.n5080 99.6594
R6951 gnd.n6396 gnd.n6395 99.6594
R6952 gnd.n5676 gnd.n5675 99.6594
R6953 gnd.n5670 gnd.n5618 99.6594
R6954 gnd.n5667 gnd.n5619 99.6594
R6955 gnd.n5663 gnd.n5620 99.6594
R6956 gnd.n5659 gnd.n5621 99.6594
R6957 gnd.n5655 gnd.n5622 99.6594
R6958 gnd.n5651 gnd.n5623 99.6594
R6959 gnd.n5647 gnd.n5624 99.6594
R6960 gnd.n7439 gnd.n322 99.6594
R6961 gnd.n7437 gnd.n7436 99.6594
R6962 gnd.n7432 gnd.n329 99.6594
R6963 gnd.n7430 gnd.n7429 99.6594
R6964 gnd.n7425 gnd.n336 99.6594
R6965 gnd.n7423 gnd.n7422 99.6594
R6966 gnd.n7418 gnd.n343 99.6594
R6967 gnd.n7416 gnd.n7415 99.6594
R6968 gnd.n348 gnd.n347 99.6594
R6969 gnd.n3840 gnd.n3839 99.6594
R6970 gnd.n3856 gnd.n3855 99.6594
R6971 gnd.n3859 gnd.n3858 99.6594
R6972 gnd.n3875 gnd.n3874 99.6594
R6973 gnd.n3878 gnd.n3877 99.6594
R6974 gnd.n3894 gnd.n3893 99.6594
R6975 gnd.n3897 gnd.n3896 99.6594
R6976 gnd.n3914 gnd.n3913 99.6594
R6977 gnd.n3917 gnd.n3916 99.6594
R6978 gnd.n6387 gnd.n5087 99.6594
R6979 gnd.n6385 gnd.n6384 99.6594
R6980 gnd.n6380 gnd.n5094 99.6594
R6981 gnd.n6378 gnd.n6377 99.6594
R6982 gnd.n6373 gnd.n5101 99.6594
R6983 gnd.n6371 gnd.n6370 99.6594
R6984 gnd.n6366 gnd.n5108 99.6594
R6985 gnd.n6364 gnd.n6363 99.6594
R6986 gnd.n6359 gnd.n5115 99.6594
R6987 gnd.n6357 gnd.n6356 99.6594
R6988 gnd.n6352 gnd.n5124 99.6594
R6989 gnd.n6350 gnd.n6349 99.6594
R6990 gnd.n6345 gnd.n6344 99.6594
R6991 gnd.n5548 gnd.n5458 99.6594
R6992 gnd.n5546 gnd.n5461 99.6594
R6993 gnd.n5542 gnd.n5541 99.6594
R6994 gnd.n5535 gnd.n5466 99.6594
R6995 gnd.n5534 gnd.n5533 99.6594
R6996 gnd.n5527 gnd.n5472 99.6594
R6997 gnd.n5526 gnd.n5525 99.6594
R6998 gnd.n5519 gnd.n5478 99.6594
R6999 gnd.n5518 gnd.n5517 99.6594
R7000 gnd.n5511 gnd.n5484 99.6594
R7001 gnd.n5510 gnd.n5509 99.6594
R7002 gnd.n5502 gnd.n5490 99.6594
R7003 gnd.n5501 gnd.n5500 99.6594
R7004 gnd.n2468 gnd.n2467 99.6594
R7005 gnd.n2477 gnd.n2476 99.6594
R7006 gnd.n2486 gnd.n2485 99.6594
R7007 gnd.n2489 gnd.n2488 99.6594
R7008 gnd.n2498 gnd.n2497 99.6594
R7009 gnd.n2507 gnd.n2506 99.6594
R7010 gnd.n2510 gnd.n2509 99.6594
R7011 gnd.n2521 gnd.n2520 99.6594
R7012 gnd.n3078 gnd.n3077 99.6594
R7013 gnd.n2700 gnd.n1058 99.6594
R7014 gnd.n2704 gnd.n1059 99.6594
R7015 gnd.n2710 gnd.n1060 99.6594
R7016 gnd.n2714 gnd.n1061 99.6594
R7017 gnd.n2720 gnd.n1062 99.6594
R7018 gnd.n2724 gnd.n1063 99.6594
R7019 gnd.n2730 gnd.n1064 99.6594
R7020 gnd.n2734 gnd.n1065 99.6594
R7021 gnd.n2691 gnd.n1066 99.6594
R7022 gnd.n2703 gnd.n1058 99.6594
R7023 gnd.n2709 gnd.n1059 99.6594
R7024 gnd.n2713 gnd.n1060 99.6594
R7025 gnd.n2719 gnd.n1061 99.6594
R7026 gnd.n2723 gnd.n1062 99.6594
R7027 gnd.n2729 gnd.n1063 99.6594
R7028 gnd.n2733 gnd.n1064 99.6594
R7029 gnd.n2690 gnd.n1065 99.6594
R7030 gnd.n2686 gnd.n1066 99.6594
R7031 gnd.n3077 gnd.n2525 99.6594
R7032 gnd.n2520 gnd.n2519 99.6594
R7033 gnd.n2509 gnd.n2508 99.6594
R7034 gnd.n2506 gnd.n2499 99.6594
R7035 gnd.n2497 gnd.n2496 99.6594
R7036 gnd.n2488 gnd.n2487 99.6594
R7037 gnd.n2485 gnd.n2478 99.6594
R7038 gnd.n2476 gnd.n2475 99.6594
R7039 gnd.n2467 gnd.n2466 99.6594
R7040 gnd.n5549 gnd.n5548 99.6594
R7041 gnd.n5543 gnd.n5461 99.6594
R7042 gnd.n5541 gnd.n5540 99.6594
R7043 gnd.n5536 gnd.n5535 99.6594
R7044 gnd.n5533 gnd.n5532 99.6594
R7045 gnd.n5528 gnd.n5527 99.6594
R7046 gnd.n5525 gnd.n5524 99.6594
R7047 gnd.n5520 gnd.n5519 99.6594
R7048 gnd.n5517 gnd.n5516 99.6594
R7049 gnd.n5512 gnd.n5511 99.6594
R7050 gnd.n5509 gnd.n5508 99.6594
R7051 gnd.n5503 gnd.n5502 99.6594
R7052 gnd.n5500 gnd.n5456 99.6594
R7053 gnd.n6344 gnd.n5126 99.6594
R7054 gnd.n6351 gnd.n6350 99.6594
R7055 gnd.n5124 gnd.n5116 99.6594
R7056 gnd.n6358 gnd.n6357 99.6594
R7057 gnd.n5115 gnd.n5109 99.6594
R7058 gnd.n6365 gnd.n6364 99.6594
R7059 gnd.n5108 gnd.n5102 99.6594
R7060 gnd.n6372 gnd.n6371 99.6594
R7061 gnd.n5101 gnd.n5095 99.6594
R7062 gnd.n6379 gnd.n6378 99.6594
R7063 gnd.n5094 gnd.n5088 99.6594
R7064 gnd.n6386 gnd.n6385 99.6594
R7065 gnd.n5087 gnd.n5084 99.6594
R7066 gnd.n3839 gnd.n3803 99.6594
R7067 gnd.n3857 gnd.n3856 99.6594
R7068 gnd.n3858 gnd.n3794 99.6594
R7069 gnd.n3876 gnd.n3875 99.6594
R7070 gnd.n3877 gnd.n3785 99.6594
R7071 gnd.n3895 gnd.n3894 99.6594
R7072 gnd.n3896 gnd.n3776 99.6594
R7073 gnd.n3915 gnd.n3914 99.6594
R7074 gnd.n3916 gnd.n3772 99.6594
R7075 gnd.n347 gnd.n344 99.6594
R7076 gnd.n7417 gnd.n7416 99.6594
R7077 gnd.n343 gnd.n337 99.6594
R7078 gnd.n7424 gnd.n7423 99.6594
R7079 gnd.n336 gnd.n330 99.6594
R7080 gnd.n7431 gnd.n7430 99.6594
R7081 gnd.n329 gnd.n323 99.6594
R7082 gnd.n7438 gnd.n7437 99.6594
R7083 gnd.n322 gnd.n319 99.6594
R7084 gnd.n5676 gnd.n5626 99.6594
R7085 gnd.n5668 gnd.n5618 99.6594
R7086 gnd.n5664 gnd.n5619 99.6594
R7087 gnd.n5660 gnd.n5620 99.6594
R7088 gnd.n5656 gnd.n5621 99.6594
R7089 gnd.n5652 gnd.n5622 99.6594
R7090 gnd.n5648 gnd.n5623 99.6594
R7091 gnd.n5624 gnd.n5418 99.6594
R7092 gnd.n6397 gnd.n6396 99.6594
R7093 gnd.n5080 gnd.n5072 99.6594
R7094 gnd.n6404 gnd.n6403 99.6594
R7095 gnd.n5071 gnd.n5065 99.6594
R7096 gnd.n6411 gnd.n6410 99.6594
R7097 gnd.n5064 gnd.n5058 99.6594
R7098 gnd.n6418 gnd.n6417 99.6594
R7099 gnd.n5057 gnd.n5054 99.6594
R7100 gnd.n5045 gnd.n1070 99.6594
R7101 gnd.n5037 gnd.n1030 99.6594
R7102 gnd.n5033 gnd.n1031 99.6594
R7103 gnd.n5029 gnd.n1032 99.6594
R7104 gnd.n5025 gnd.n1033 99.6594
R7105 gnd.n5021 gnd.n1034 99.6594
R7106 gnd.n5017 gnd.n1035 99.6594
R7107 gnd.n5013 gnd.n1036 99.6594
R7108 gnd.n5008 gnd.n1037 99.6594
R7109 gnd.n5004 gnd.n1038 99.6594
R7110 gnd.n5000 gnd.n1039 99.6594
R7111 gnd.n4996 gnd.n1040 99.6594
R7112 gnd.n4992 gnd.n1041 99.6594
R7113 gnd.n4988 gnd.n1042 99.6594
R7114 gnd.n4984 gnd.n1043 99.6594
R7115 gnd.n4980 gnd.n1044 99.6594
R7116 gnd.n4976 gnd.n1045 99.6594
R7117 gnd.n4972 gnd.n1046 99.6594
R7118 gnd.n4968 gnd.n1047 99.6594
R7119 gnd.n4964 gnd.n1048 99.6594
R7120 gnd.n4960 gnd.n1049 99.6594
R7121 gnd.n4956 gnd.n1050 99.6594
R7122 gnd.n4952 gnd.n1051 99.6594
R7123 gnd.n4948 gnd.n1052 99.6594
R7124 gnd.n4944 gnd.n1053 99.6594
R7125 gnd.n4940 gnd.n1054 99.6594
R7126 gnd.n4936 gnd.n1055 99.6594
R7127 gnd.n4932 gnd.n1056 99.6594
R7128 gnd.n1140 gnd.n1057 99.6594
R7129 gnd.n2455 gnd.n2454 99.6594
R7130 gnd.n2446 gnd.n2351 99.6594
R7131 gnd.n2445 gnd.n2444 99.6594
R7132 gnd.n2436 gnd.n2355 99.6594
R7133 gnd.n2435 gnd.n2434 99.6594
R7134 gnd.n2426 gnd.n2359 99.6594
R7135 gnd.n2425 gnd.n2424 99.6594
R7136 gnd.n2416 gnd.n2363 99.6594
R7137 gnd.n2415 gnd.n2414 99.6594
R7138 gnd.n2406 gnd.n2367 99.6594
R7139 gnd.n2405 gnd.n2404 99.6594
R7140 gnd.n2396 gnd.n2373 99.6594
R7141 gnd.n2395 gnd.n2394 99.6594
R7142 gnd.n2386 gnd.n2377 99.6594
R7143 gnd.n2385 gnd.n2384 99.6594
R7144 gnd.n1426 gnd.n1421 99.6594
R7145 gnd.n4742 gnd.n4741 99.6594
R7146 gnd.n1420 gnd.n1414 99.6594
R7147 gnd.n4749 gnd.n4748 99.6594
R7148 gnd.n1413 gnd.n1405 99.6594
R7149 gnd.n4757 gnd.n4756 99.6594
R7150 gnd.n1404 gnd.n1398 99.6594
R7151 gnd.n4764 gnd.n4763 99.6594
R7152 gnd.n1397 gnd.n1391 99.6594
R7153 gnd.n4771 gnd.n4770 99.6594
R7154 gnd.n1390 gnd.n1383 99.6594
R7155 gnd.n4778 gnd.n4777 99.6594
R7156 gnd.n4781 gnd.n4780 99.6594
R7157 gnd.n4179 gnd.n4178 99.6594
R7158 gnd.n4181 gnd.n4170 99.6594
R7159 gnd.n4190 gnd.n4189 99.6594
R7160 gnd.n4191 gnd.n4166 99.6594
R7161 gnd.n4200 gnd.n4199 99.6594
R7162 gnd.n4201 gnd.n4162 99.6594
R7163 gnd.n4210 gnd.n4209 99.6594
R7164 gnd.n4211 gnd.n4158 99.6594
R7165 gnd.n4223 gnd.n4222 99.6594
R7166 gnd.n4224 gnd.n4154 99.6594
R7167 gnd.n4233 gnd.n4232 99.6594
R7168 gnd.n4234 gnd.n4150 99.6594
R7169 gnd.n4246 gnd.n4245 99.6594
R7170 gnd.n4247 gnd.n1838 99.6594
R7171 gnd.n4256 gnd.n4255 99.6594
R7172 gnd.n4257 gnd.n1834 99.6594
R7173 gnd.n4266 gnd.n4265 99.6594
R7174 gnd.n4267 gnd.n1830 99.6594
R7175 gnd.n4278 gnd.n4277 99.6594
R7176 gnd.n4279 gnd.n1826 99.6594
R7177 gnd.n4288 gnd.n4287 99.6594
R7178 gnd.n4289 gnd.n1822 99.6594
R7179 gnd.n4298 gnd.n4297 99.6594
R7180 gnd.n4299 gnd.n1818 99.6594
R7181 gnd.n4308 gnd.n4307 99.6594
R7182 gnd.n4309 gnd.n1814 99.6594
R7183 gnd.n4319 gnd.n4318 99.6594
R7184 gnd.n4322 gnd.n4321 99.6594
R7185 gnd.n7449 gnd.n7448 99.6594
R7186 gnd.n316 gnd.n308 99.6594
R7187 gnd.n7456 gnd.n7455 99.6594
R7188 gnd.n307 gnd.n301 99.6594
R7189 gnd.n7463 gnd.n7462 99.6594
R7190 gnd.n300 gnd.n294 99.6594
R7191 gnd.n7470 gnd.n7469 99.6594
R7192 gnd.n293 gnd.n287 99.6594
R7193 gnd.n7477 gnd.n7476 99.6594
R7194 gnd.n7480 gnd.n7479 99.6594
R7195 gnd.n284 gnd.n276 99.6594
R7196 gnd.n7489 gnd.n7488 99.6594
R7197 gnd.n275 gnd.n269 99.6594
R7198 gnd.n7496 gnd.n7495 99.6594
R7199 gnd.n268 gnd.n262 99.6594
R7200 gnd.n7503 gnd.n7502 99.6594
R7201 gnd.n261 gnd.n255 99.6594
R7202 gnd.n7510 gnd.n7509 99.6594
R7203 gnd.n254 gnd.n248 99.6594
R7204 gnd.n7517 gnd.n7516 99.6594
R7205 gnd.n247 gnd.n241 99.6594
R7206 gnd.n7527 gnd.n7526 99.6594
R7207 gnd.n240 gnd.n234 99.6594
R7208 gnd.n7534 gnd.n7533 99.6594
R7209 gnd.n233 gnd.n227 99.6594
R7210 gnd.n7541 gnd.n7540 99.6594
R7211 gnd.n226 gnd.n220 99.6594
R7212 gnd.n7548 gnd.n7547 99.6594
R7213 gnd.n219 gnd.n216 99.6594
R7214 gnd.n3069 gnd.n2335 99.6594
R7215 gnd.n2532 gnd.n2531 99.6594
R7216 gnd.n2533 gnd.n2344 99.6594
R7217 gnd.n2535 gnd.n2534 99.6594
R7218 gnd.n2537 gnd.n2462 99.6594
R7219 gnd.n2538 gnd.n2471 99.6594
R7220 gnd.n2540 gnd.n2539 99.6594
R7221 gnd.n2542 gnd.n2482 99.6594
R7222 gnd.n2543 gnd.n2492 99.6594
R7223 gnd.n2545 gnd.n2544 99.6594
R7224 gnd.n2547 gnd.n2503 99.6594
R7225 gnd.n2548 gnd.n2513 99.6594
R7226 gnd.n2551 gnd.n2550 99.6594
R7227 gnd.n3072 gnd.n3071 99.6594
R7228 gnd.n3069 gnd.n2339 99.6594
R7229 gnd.n2532 gnd.n2343 99.6594
R7230 gnd.n2533 gnd.n2345 99.6594
R7231 gnd.n2535 gnd.n2461 99.6594
R7232 gnd.n2537 gnd.n2536 99.6594
R7233 gnd.n2538 gnd.n2472 99.6594
R7234 gnd.n2540 gnd.n2481 99.6594
R7235 gnd.n2542 gnd.n2541 99.6594
R7236 gnd.n2543 gnd.n2493 99.6594
R7237 gnd.n2545 gnd.n2502 99.6594
R7238 gnd.n2547 gnd.n2546 99.6594
R7239 gnd.n2548 gnd.n2514 99.6594
R7240 gnd.n2551 gnd.n2529 99.6594
R7241 gnd.n3071 gnd.n2332 99.6594
R7242 gnd.n3820 gnd.n3815 99.6594
R7243 gnd.n3824 gnd.n3822 99.6594
R7244 gnd.n3831 gnd.n3811 99.6594
R7245 gnd.n3835 gnd.n3833 99.6594
R7246 gnd.n3846 gnd.n3808 99.6594
R7247 gnd.n3850 gnd.n3848 99.6594
R7248 gnd.n3865 gnd.n3799 99.6594
R7249 gnd.n3869 gnd.n3867 99.6594
R7250 gnd.n3884 gnd.n3790 99.6594
R7251 gnd.n3888 gnd.n3886 99.6594
R7252 gnd.n3903 gnd.n3781 99.6594
R7253 gnd.n3906 gnd.n3905 99.6594
R7254 gnd.n3924 gnd.n3923 99.6594
R7255 gnd.n3927 gnd.n3926 99.6594
R7256 gnd.n3905 gnd.n3904 99.6594
R7257 gnd.n3887 gnd.n3781 99.6594
R7258 gnd.n3886 gnd.n3885 99.6594
R7259 gnd.n3868 gnd.n3790 99.6594
R7260 gnd.n3867 gnd.n3866 99.6594
R7261 gnd.n3849 gnd.n3799 99.6594
R7262 gnd.n3848 gnd.n3847 99.6594
R7263 gnd.n3834 gnd.n3808 99.6594
R7264 gnd.n3833 gnd.n3832 99.6594
R7265 gnd.n3823 gnd.n3811 99.6594
R7266 gnd.n3822 gnd.n3821 99.6594
R7267 gnd.n3815 gnd.n1578 99.6594
R7268 gnd.n3928 gnd.n3927 99.6594
R7269 gnd.n3925 gnd.n3924 99.6594
R7270 gnd.n2515 gnd.t143 98.63
R7271 gnd.n3773 gnd.t168 98.63
R7272 gnd.n2522 gnd.t192 98.63
R7273 gnd.n4217 gnd.t165 98.63
R7274 gnd.n4269 gnd.t156 98.63
R7275 gnd.n1810 gnd.t91 98.63
R7276 gnd.n313 gnd.t189 98.63
R7277 gnd.n280 gnd.t104 98.63
R7278 gnd.n7520 gnd.t145 98.63
R7279 gnd.n350 gnd.t135 98.63
R7280 gnd.n1090 gnd.t119 98.63
R7281 gnd.n1112 gnd.t116 98.63
R7282 gnd.n1134 gnd.t95 98.63
R7283 gnd.n2687 gnd.t174 98.63
R7284 gnd.n1409 gnd.t176 98.63
R7285 gnd.n2348 gnd.t112 98.63
R7286 gnd.n2370 gnd.t138 98.63
R7287 gnd.n3763 gnd.t125 98.63
R7288 gnd.n2188 gnd.t109 92.8196
R7289 gnd.n1879 gnd.t132 92.8196
R7290 gnd.n4668 gnd.t162 92.8118
R7291 gnd.n4011 gnd.t183 92.8118
R7292 gnd.n1477 gnd.n1476 81.8399
R7293 gnd.n5644 gnd.t152 74.8376
R7294 gnd.n5078 gnd.t181 74.8376
R7295 gnd.n2189 gnd.t108 72.8438
R7296 gnd.n1880 gnd.t133 72.8438
R7297 gnd.n1478 gnd.n1471 72.8411
R7298 gnd.n1484 gnd.n1469 72.8411
R7299 gnd.n4007 gnd.n4006 72.8411
R7300 gnd.n2516 gnd.t142 72.836
R7301 gnd.n4669 gnd.t161 72.836
R7302 gnd.n4012 gnd.t184 72.836
R7303 gnd.n3774 gnd.t167 72.836
R7304 gnd.n2523 gnd.t193 72.836
R7305 gnd.n4218 gnd.t164 72.836
R7306 gnd.n4270 gnd.t155 72.836
R7307 gnd.n1811 gnd.t90 72.836
R7308 gnd.n314 gnd.t190 72.836
R7309 gnd.n281 gnd.t105 72.836
R7310 gnd.n7521 gnd.t146 72.836
R7311 gnd.n351 gnd.t136 72.836
R7312 gnd.n1091 gnd.t118 72.836
R7313 gnd.n1113 gnd.t115 72.836
R7314 gnd.n1135 gnd.t94 72.836
R7315 gnd.n2688 gnd.t173 72.836
R7316 gnd.n1410 gnd.t177 72.836
R7317 gnd.n2349 gnd.t113 72.836
R7318 gnd.n2371 gnd.t139 72.836
R7319 gnd.n3764 gnd.t126 72.836
R7320 gnd.n4072 gnd.n1847 71.676
R7321 gnd.n4068 gnd.n1848 71.676
R7322 gnd.n4064 gnd.n1849 71.676
R7323 gnd.n4060 gnd.n1850 71.676
R7324 gnd.n4056 gnd.n1851 71.676
R7325 gnd.n4052 gnd.n1852 71.676
R7326 gnd.n4048 gnd.n1853 71.676
R7327 gnd.n4044 gnd.n1854 71.676
R7328 gnd.n4040 gnd.n1855 71.676
R7329 gnd.n4036 gnd.n1856 71.676
R7330 gnd.n4032 gnd.n1857 71.676
R7331 gnd.n4028 gnd.n1858 71.676
R7332 gnd.n4024 gnd.n1859 71.676
R7333 gnd.n4020 gnd.n1860 71.676
R7334 gnd.n4015 gnd.n1861 71.676
R7335 gnd.n1862 gnd.n1845 71.676
R7336 gnd.n4144 gnd.n1844 71.676
R7337 gnd.n4142 gnd.n4141 71.676
R7338 gnd.n4136 gnd.n1877 71.676
R7339 gnd.n4132 gnd.n1876 71.676
R7340 gnd.n4128 gnd.n1875 71.676
R7341 gnd.n4124 gnd.n1874 71.676
R7342 gnd.n4120 gnd.n1873 71.676
R7343 gnd.n4116 gnd.n1872 71.676
R7344 gnd.n4112 gnd.n1871 71.676
R7345 gnd.n4108 gnd.n1870 71.676
R7346 gnd.n4104 gnd.n1869 71.676
R7347 gnd.n4100 gnd.n1868 71.676
R7348 gnd.n4096 gnd.n1867 71.676
R7349 gnd.n4092 gnd.n1866 71.676
R7350 gnd.n4088 gnd.n1865 71.676
R7351 gnd.n4084 gnd.n1864 71.676
R7352 gnd.n4080 gnd.n1863 71.676
R7353 gnd.n4732 gnd.n4731 71.676
R7354 gnd.n4726 gnd.n1433 71.676
R7355 gnd.n4723 gnd.n1434 71.676
R7356 gnd.n4719 gnd.n1435 71.676
R7357 gnd.n4715 gnd.n1436 71.676
R7358 gnd.n4711 gnd.n1437 71.676
R7359 gnd.n4707 gnd.n1438 71.676
R7360 gnd.n4703 gnd.n1439 71.676
R7361 gnd.n4699 gnd.n1440 71.676
R7362 gnd.n4695 gnd.n1441 71.676
R7363 gnd.n4691 gnd.n1442 71.676
R7364 gnd.n4687 gnd.n1443 71.676
R7365 gnd.n4683 gnd.n1444 71.676
R7366 gnd.n4679 gnd.n1445 71.676
R7367 gnd.n4675 gnd.n1446 71.676
R7368 gnd.n4671 gnd.n1447 71.676
R7369 gnd.n1448 gnd.n1432 71.676
R7370 gnd.n2192 gnd.n1449 71.676
R7371 gnd.n2197 gnd.n1450 71.676
R7372 gnd.n2201 gnd.n1451 71.676
R7373 gnd.n2205 gnd.n1452 71.676
R7374 gnd.n2209 gnd.n1453 71.676
R7375 gnd.n2213 gnd.n1454 71.676
R7376 gnd.n2217 gnd.n1455 71.676
R7377 gnd.n2221 gnd.n1456 71.676
R7378 gnd.n2225 gnd.n1457 71.676
R7379 gnd.n2229 gnd.n1458 71.676
R7380 gnd.n2233 gnd.n1459 71.676
R7381 gnd.n2237 gnd.n1460 71.676
R7382 gnd.n2241 gnd.n1461 71.676
R7383 gnd.n2245 gnd.n1462 71.676
R7384 gnd.n2249 gnd.n1463 71.676
R7385 gnd.n4732 gnd.n1466 71.676
R7386 gnd.n4724 gnd.n1433 71.676
R7387 gnd.n4720 gnd.n1434 71.676
R7388 gnd.n4716 gnd.n1435 71.676
R7389 gnd.n4712 gnd.n1436 71.676
R7390 gnd.n4708 gnd.n1437 71.676
R7391 gnd.n4704 gnd.n1438 71.676
R7392 gnd.n4700 gnd.n1439 71.676
R7393 gnd.n4696 gnd.n1440 71.676
R7394 gnd.n4692 gnd.n1441 71.676
R7395 gnd.n4688 gnd.n1442 71.676
R7396 gnd.n4684 gnd.n1443 71.676
R7397 gnd.n4680 gnd.n1444 71.676
R7398 gnd.n4676 gnd.n1445 71.676
R7399 gnd.n4672 gnd.n1446 71.676
R7400 gnd.n4735 gnd.n4734 71.676
R7401 gnd.n2191 gnd.n1448 71.676
R7402 gnd.n2196 gnd.n1449 71.676
R7403 gnd.n2200 gnd.n1450 71.676
R7404 gnd.n2204 gnd.n1451 71.676
R7405 gnd.n2208 gnd.n1452 71.676
R7406 gnd.n2212 gnd.n1453 71.676
R7407 gnd.n2216 gnd.n1454 71.676
R7408 gnd.n2220 gnd.n1455 71.676
R7409 gnd.n2224 gnd.n1456 71.676
R7410 gnd.n2228 gnd.n1457 71.676
R7411 gnd.n2232 gnd.n1458 71.676
R7412 gnd.n2236 gnd.n1459 71.676
R7413 gnd.n2240 gnd.n1460 71.676
R7414 gnd.n2244 gnd.n1461 71.676
R7415 gnd.n2248 gnd.n1462 71.676
R7416 gnd.n2252 gnd.n1463 71.676
R7417 gnd.n4083 gnd.n1863 71.676
R7418 gnd.n4087 gnd.n1864 71.676
R7419 gnd.n4091 gnd.n1865 71.676
R7420 gnd.n4095 gnd.n1866 71.676
R7421 gnd.n4099 gnd.n1867 71.676
R7422 gnd.n4103 gnd.n1868 71.676
R7423 gnd.n4107 gnd.n1869 71.676
R7424 gnd.n4111 gnd.n1870 71.676
R7425 gnd.n4115 gnd.n1871 71.676
R7426 gnd.n4119 gnd.n1872 71.676
R7427 gnd.n4123 gnd.n1873 71.676
R7428 gnd.n4127 gnd.n1874 71.676
R7429 gnd.n4131 gnd.n1875 71.676
R7430 gnd.n4135 gnd.n1876 71.676
R7431 gnd.n1878 gnd.n1877 71.676
R7432 gnd.n4143 gnd.n4142 71.676
R7433 gnd.n4147 gnd.n4146 71.676
R7434 gnd.n4014 gnd.n1862 71.676
R7435 gnd.n4019 gnd.n1861 71.676
R7436 gnd.n4023 gnd.n1860 71.676
R7437 gnd.n4027 gnd.n1859 71.676
R7438 gnd.n4031 gnd.n1858 71.676
R7439 gnd.n4035 gnd.n1857 71.676
R7440 gnd.n4039 gnd.n1856 71.676
R7441 gnd.n4043 gnd.n1855 71.676
R7442 gnd.n4047 gnd.n1854 71.676
R7443 gnd.n4051 gnd.n1853 71.676
R7444 gnd.n4055 gnd.n1852 71.676
R7445 gnd.n4059 gnd.n1851 71.676
R7446 gnd.n4063 gnd.n1850 71.676
R7447 gnd.n4067 gnd.n1849 71.676
R7448 gnd.n4071 gnd.n1848 71.676
R7449 gnd.n1886 gnd.n1847 71.676
R7450 gnd.n8 gnd.t256 69.1507
R7451 gnd.n14 gnd.t51 68.4792
R7452 gnd.n13 gnd.t357 68.4792
R7453 gnd.n12 gnd.t349 68.4792
R7454 gnd.n11 gnd.t232 68.4792
R7455 gnd.n10 gnd.t269 68.4792
R7456 gnd.n9 gnd.t355 68.4792
R7457 gnd.n8 gnd.t211 68.4792
R7458 gnd.n5556 gnd.n5457 64.369
R7459 gnd.n2194 gnd.n2189 59.5399
R7460 gnd.n4138 gnd.n1880 59.5399
R7461 gnd.n4670 gnd.n4669 59.5399
R7462 gnd.n4017 gnd.n4012 59.5399
R7463 gnd.n4667 gnd.n1487 59.1804
R7464 gnd.n6427 gnd.n5047 57.3586
R7465 gnd.n5046 gnd.n1068 57.3586
R7466 gnd.n7557 gnd.n212 57.3586
R7467 gnd.n5263 gnd.t26 56.407
R7468 gnd.n5216 gnd.t205 56.407
R7469 gnd.n5231 gnd.t213 56.407
R7470 gnd.n5247 gnd.t3 56.407
R7471 gnd.n64 gnd.t17 56.407
R7472 gnd.n17 gnd.t214 56.407
R7473 gnd.n32 gnd.t220 56.407
R7474 gnd.n48 gnd.t224 56.407
R7475 gnd.n5276 gnd.t229 55.8337
R7476 gnd.n5229 gnd.t261 55.8337
R7477 gnd.n5244 gnd.t215 55.8337
R7478 gnd.n5260 gnd.t54 55.8337
R7479 gnd.n77 gnd.t303 55.8337
R7480 gnd.n30 gnd.t302 55.8337
R7481 gnd.n45 gnd.t309 55.8337
R7482 gnd.n61 gnd.t298 55.8337
R7483 gnd.n1475 gnd.n1474 54.358
R7484 gnd.n4004 gnd.n4003 54.358
R7485 gnd.n5263 gnd.n5262 53.0052
R7486 gnd.n5265 gnd.n5264 53.0052
R7487 gnd.n5267 gnd.n5266 53.0052
R7488 gnd.n5269 gnd.n5268 53.0052
R7489 gnd.n5271 gnd.n5270 53.0052
R7490 gnd.n5273 gnd.n5272 53.0052
R7491 gnd.n5275 gnd.n5274 53.0052
R7492 gnd.n5216 gnd.n5215 53.0052
R7493 gnd.n5218 gnd.n5217 53.0052
R7494 gnd.n5220 gnd.n5219 53.0052
R7495 gnd.n5222 gnd.n5221 53.0052
R7496 gnd.n5224 gnd.n5223 53.0052
R7497 gnd.n5226 gnd.n5225 53.0052
R7498 gnd.n5228 gnd.n5227 53.0052
R7499 gnd.n5231 gnd.n5230 53.0052
R7500 gnd.n5233 gnd.n5232 53.0052
R7501 gnd.n5235 gnd.n5234 53.0052
R7502 gnd.n5237 gnd.n5236 53.0052
R7503 gnd.n5239 gnd.n5238 53.0052
R7504 gnd.n5241 gnd.n5240 53.0052
R7505 gnd.n5243 gnd.n5242 53.0052
R7506 gnd.n5247 gnd.n5246 53.0052
R7507 gnd.n5249 gnd.n5248 53.0052
R7508 gnd.n5251 gnd.n5250 53.0052
R7509 gnd.n5253 gnd.n5252 53.0052
R7510 gnd.n5255 gnd.n5254 53.0052
R7511 gnd.n5257 gnd.n5256 53.0052
R7512 gnd.n5259 gnd.n5258 53.0052
R7513 gnd.n76 gnd.n75 53.0052
R7514 gnd.n74 gnd.n73 53.0052
R7515 gnd.n72 gnd.n71 53.0052
R7516 gnd.n70 gnd.n69 53.0052
R7517 gnd.n68 gnd.n67 53.0052
R7518 gnd.n66 gnd.n65 53.0052
R7519 gnd.n64 gnd.n63 53.0052
R7520 gnd.n29 gnd.n28 53.0052
R7521 gnd.n27 gnd.n26 53.0052
R7522 gnd.n25 gnd.n24 53.0052
R7523 gnd.n23 gnd.n22 53.0052
R7524 gnd.n21 gnd.n20 53.0052
R7525 gnd.n19 gnd.n18 53.0052
R7526 gnd.n17 gnd.n16 53.0052
R7527 gnd.n44 gnd.n43 53.0052
R7528 gnd.n42 gnd.n41 53.0052
R7529 gnd.n40 gnd.n39 53.0052
R7530 gnd.n38 gnd.n37 53.0052
R7531 gnd.n36 gnd.n35 53.0052
R7532 gnd.n34 gnd.n33 53.0052
R7533 gnd.n32 gnd.n31 53.0052
R7534 gnd.n60 gnd.n59 53.0052
R7535 gnd.n58 gnd.n57 53.0052
R7536 gnd.n56 gnd.n55 53.0052
R7537 gnd.n54 gnd.n53 53.0052
R7538 gnd.n52 gnd.n51 53.0052
R7539 gnd.n50 gnd.n49 53.0052
R7540 gnd.n48 gnd.n47 53.0052
R7541 gnd.n3995 gnd.n3994 52.4801
R7542 gnd.n6272 gnd.t359 52.3082
R7543 gnd.n6240 gnd.t236 52.3082
R7544 gnd.n6208 gnd.t271 52.3082
R7545 gnd.n6177 gnd.t222 52.3082
R7546 gnd.n6145 gnd.t258 52.3082
R7547 gnd.n6113 gnd.t277 52.3082
R7548 gnd.n6081 gnd.t352 52.3082
R7549 gnd.n6050 gnd.t253 52.3082
R7550 gnd.n6102 gnd.n6070 51.4173
R7551 gnd.n6166 gnd.n6165 50.455
R7552 gnd.n6134 gnd.n6133 50.455
R7553 gnd.n6102 gnd.n6101 50.455
R7554 gnd.n5494 gnd.n5493 45.1884
R7555 gnd.n5122 gnd.n5121 45.1884
R7556 gnd.n4075 gnd.n4010 44.3322
R7557 gnd.n1478 gnd.n1477 44.3189
R7558 gnd.n2517 gnd.n2516 42.2793
R7559 gnd.n3919 gnd.n3774 42.2793
R7560 gnd.n5506 gnd.n5494 42.2793
R7561 gnd.n5123 gnd.n5122 42.2793
R7562 gnd.n5646 gnd.n5644 42.2793
R7563 gnd.n5079 gnd.n5078 42.2793
R7564 gnd.n3080 gnd.n2523 42.2793
R7565 gnd.n4219 gnd.n4218 42.2793
R7566 gnd.n4271 gnd.n4270 42.2793
R7567 gnd.n1812 gnd.n1811 42.2793
R7568 gnd.n315 gnd.n314 42.2793
R7569 gnd.n7485 gnd.n281 42.2793
R7570 gnd.n7522 gnd.n7521 42.2793
R7571 gnd.n7413 gnd.n351 42.2793
R7572 gnd.n5010 gnd.n1091 42.2793
R7573 gnd.n4970 gnd.n1113 42.2793
R7574 gnd.n4930 gnd.n1135 42.2793
R7575 gnd.n2740 gnd.n2688 42.2793
R7576 gnd.n4752 gnd.n1410 42.2793
R7577 gnd.n2350 gnd.n2349 42.2793
R7578 gnd.n2372 gnd.n2371 42.2793
R7579 gnd.n3765 gnd.n3764 42.2793
R7580 gnd.n1476 gnd.n1475 41.6274
R7581 gnd.n4005 gnd.n4004 41.6274
R7582 gnd.n1485 gnd.n1484 40.8975
R7583 gnd.n4008 gnd.n4007 40.8975
R7584 gnd.n6631 gnd.n801 39.6473
R7585 gnd.n6625 gnd.n801 39.6473
R7586 gnd.n6625 gnd.n6624 39.6473
R7587 gnd.n6624 gnd.n6623 39.6473
R7588 gnd.n6623 gnd.n808 39.6473
R7589 gnd.n6617 gnd.n808 39.6473
R7590 gnd.n6617 gnd.n6616 39.6473
R7591 gnd.n6616 gnd.n6615 39.6473
R7592 gnd.n6615 gnd.n816 39.6473
R7593 gnd.n6609 gnd.n816 39.6473
R7594 gnd.n6609 gnd.n6608 39.6473
R7595 gnd.n6608 gnd.n6607 39.6473
R7596 gnd.n6607 gnd.n824 39.6473
R7597 gnd.n6601 gnd.n824 39.6473
R7598 gnd.n6601 gnd.n6600 39.6473
R7599 gnd.n6600 gnd.n6599 39.6473
R7600 gnd.n6599 gnd.n832 39.6473
R7601 gnd.n6593 gnd.n832 39.6473
R7602 gnd.n6593 gnd.n6592 39.6473
R7603 gnd.n6592 gnd.n6591 39.6473
R7604 gnd.n6591 gnd.n840 39.6473
R7605 gnd.n6585 gnd.n840 39.6473
R7606 gnd.n6585 gnd.n6584 39.6473
R7607 gnd.n6584 gnd.n6583 39.6473
R7608 gnd.n6583 gnd.n848 39.6473
R7609 gnd.n6577 gnd.n848 39.6473
R7610 gnd.n6577 gnd.n6576 39.6473
R7611 gnd.n6576 gnd.n6575 39.6473
R7612 gnd.n6575 gnd.n856 39.6473
R7613 gnd.n6569 gnd.n856 39.6473
R7614 gnd.n6569 gnd.n6568 39.6473
R7615 gnd.n6568 gnd.n6567 39.6473
R7616 gnd.n6567 gnd.n864 39.6473
R7617 gnd.n6561 gnd.n864 39.6473
R7618 gnd.n6561 gnd.n6560 39.6473
R7619 gnd.n6560 gnd.n6559 39.6473
R7620 gnd.n6559 gnd.n872 39.6473
R7621 gnd.n6553 gnd.n872 39.6473
R7622 gnd.n6553 gnd.n6552 39.6473
R7623 gnd.n6552 gnd.n6551 39.6473
R7624 gnd.n6551 gnd.n880 39.6473
R7625 gnd.n6545 gnd.n880 39.6473
R7626 gnd.n6545 gnd.n6544 39.6473
R7627 gnd.n6544 gnd.n6543 39.6473
R7628 gnd.n6543 gnd.n888 39.6473
R7629 gnd.n6537 gnd.n888 39.6473
R7630 gnd.n6537 gnd.n6536 39.6473
R7631 gnd.n6536 gnd.n6535 39.6473
R7632 gnd.n6535 gnd.n896 39.6473
R7633 gnd.n6529 gnd.n896 39.6473
R7634 gnd.n6529 gnd.n6528 39.6473
R7635 gnd.n6528 gnd.n6527 39.6473
R7636 gnd.n6527 gnd.n904 39.6473
R7637 gnd.n6521 gnd.n904 39.6473
R7638 gnd.n6521 gnd.n6520 39.6473
R7639 gnd.n6520 gnd.n6519 39.6473
R7640 gnd.n6519 gnd.n912 39.6473
R7641 gnd.n6513 gnd.n912 39.6473
R7642 gnd.n6513 gnd.n6512 39.6473
R7643 gnd.n6512 gnd.n6511 39.6473
R7644 gnd.n6511 gnd.n920 39.6473
R7645 gnd.n6505 gnd.n920 39.6473
R7646 gnd.n6505 gnd.n6504 39.6473
R7647 gnd.n6504 gnd.n6503 39.6473
R7648 gnd.n6503 gnd.n928 39.6473
R7649 gnd.n6497 gnd.n928 39.6473
R7650 gnd.n6497 gnd.n6496 39.6473
R7651 gnd.n6496 gnd.n6495 39.6473
R7652 gnd.n6495 gnd.n936 39.6473
R7653 gnd.n6489 gnd.n936 39.6473
R7654 gnd.n6489 gnd.n6488 39.6473
R7655 gnd.n6488 gnd.n6487 39.6473
R7656 gnd.n6487 gnd.n944 39.6473
R7657 gnd.n6481 gnd.n944 39.6473
R7658 gnd.n6481 gnd.n6480 39.6473
R7659 gnd.n6480 gnd.n6479 39.6473
R7660 gnd.n6479 gnd.n952 39.6473
R7661 gnd.n6473 gnd.n952 39.6473
R7662 gnd.n6473 gnd.n6472 39.6473
R7663 gnd.n6472 gnd.n6471 39.6473
R7664 gnd.n6471 gnd.n960 39.6473
R7665 gnd.n6465 gnd.n960 39.6473
R7666 gnd.n6465 gnd.n6464 39.6473
R7667 gnd.n1484 gnd.n1483 35.055
R7668 gnd.n1479 gnd.n1478 35.055
R7669 gnd.n3997 gnd.n3996 35.055
R7670 gnd.n4007 gnd.n3993 35.055
R7671 gnd.n5556 gnd.n5452 31.8661
R7672 gnd.n5564 gnd.n5452 31.8661
R7673 gnd.n5572 gnd.n5446 31.8661
R7674 gnd.n5572 gnd.n5440 31.8661
R7675 gnd.n5580 gnd.n5440 31.8661
R7676 gnd.n5580 gnd.n5433 31.8661
R7677 gnd.n5588 gnd.n5433 31.8661
R7678 gnd.n5588 gnd.n5434 31.8661
R7679 gnd.n5687 gnd.n5419 31.8661
R7680 gnd.n4922 gnd.n1068 31.8661
R7681 gnd.n4916 gnd.n1152 31.8661
R7682 gnd.n4916 gnd.n1155 31.8661
R7683 gnd.n4910 gnd.n1155 31.8661
R7684 gnd.n4910 gnd.n1167 31.8661
R7685 gnd.n4904 gnd.n1177 31.8661
R7686 gnd.n3054 gnd.n1376 31.8661
R7687 gnd.n3058 gnd.n3057 31.8661
R7688 gnd.n3058 gnd.n2530 31.8661
R7689 gnd.n3068 gnd.n2333 31.8661
R7690 gnd.n4561 gnd.n1581 31.8661
R7691 gnd.n4555 gnd.n4554 31.8661
R7692 gnd.n4554 gnd.n4553 31.8661
R7693 gnd.n4547 gnd.n1599 31.8661
R7694 gnd.n7581 gnd.n175 31.8661
R7695 gnd.n7575 gnd.n185 31.8661
R7696 gnd.n7569 gnd.n185 31.8661
R7697 gnd.n7569 gnd.n194 31.8661
R7698 gnd.n7563 gnd.n194 31.8661
R7699 gnd.n7557 gnd.n209 31.8661
R7700 gnd.n4081 gnd.n1881 30.1273
R7701 gnd.n3259 gnd.n2251 30.1273
R7702 gnd.n4892 gnd.n1194 26.7676
R7703 gnd.n4886 gnd.n1204 26.7676
R7704 gnd.n2819 gnd.n1207 26.7676
R7705 gnd.n2825 gnd.n1217 26.7676
R7706 gnd.n4874 gnd.n1224 26.7676
R7707 gnd.n4868 gnd.n1235 26.7676
R7708 gnd.n4862 gnd.n1245 26.7676
R7709 gnd.n2640 gnd.n1248 26.7676
R7710 gnd.n2852 gnd.n2643 26.7676
R7711 gnd.n2884 gnd.n2625 26.7676
R7712 gnd.n2878 gnd.n2621 26.7676
R7713 gnd.n2903 gnd.n2611 26.7676
R7714 gnd.n2939 gnd.n2597 26.7676
R7715 gnd.n2910 gnd.n1265 26.7676
R7716 gnd.n4848 gnd.n1274 26.7676
R7717 gnd.n2916 gnd.n2915 26.7676
R7718 gnd.n4842 gnd.n1283 26.7676
R7719 gnd.n4836 gnd.n1293 26.7676
R7720 gnd.n2979 gnd.n1296 26.7676
R7721 gnd.n2987 gnd.n1306 26.7676
R7722 gnd.n4824 gnd.n1313 26.7676
R7723 gnd.n2994 gnd.n2580 26.7676
R7724 gnd.n4818 gnd.n1323 26.7676
R7725 gnd.n4812 gnd.n1333 26.7676
R7726 gnd.n3036 gnd.n1336 26.7676
R7727 gnd.n3009 gnd.n1346 26.7676
R7728 gnd.n4800 gnd.n1353 26.7676
R7729 gnd.n3014 gnd.n1356 26.7676
R7730 gnd.n4794 gnd.n1364 26.7676
R7731 gnd.n4788 gnd.n1373 26.7676
R7732 gnd.n4546 gnd.n1602 26.7676
R7733 gnd.n4540 gnd.n1614 26.7676
R7734 gnd.n4333 gnd.n1623 26.7676
R7735 gnd.n4534 gnd.n1626 26.7676
R7736 gnd.n4341 gnd.n1634 26.7676
R7737 gnd.n4347 gnd.n1643 26.7676
R7738 gnd.n4522 gnd.n1646 26.7676
R7739 gnd.n4516 gnd.n1657 26.7676
R7740 gnd.n4392 gnd.n4391 26.7676
R7741 gnd.n4510 gnd.n1666 26.7676
R7742 gnd.n4362 gnd.n1674 26.7676
R7743 gnd.n4367 gnd.n1683 26.7676
R7744 gnd.n4498 gnd.n1686 26.7676
R7745 gnd.n4492 gnd.n1697 26.7676
R7746 gnd.n4415 gnd.n4414 26.7676
R7747 gnd.n4486 gnd.n1706 26.7676
R7748 gnd.n4445 gnd.n1712 26.7676
R7749 gnd.n4456 gnd.n1721 26.7676
R7750 gnd.n4474 gnd.n1724 26.7676
R7751 gnd.n4423 gnd.n1732 26.7676
R7752 gnd.n7631 gnd.n87 26.7676
R7753 gnd.n7323 gnd.n381 26.7676
R7754 gnd.n7623 gnd.n105 26.7676
R7755 gnd.n7334 gnd.n114 26.7676
R7756 gnd.n7342 gnd.n123 26.7676
R7757 gnd.n7348 gnd.n132 26.7676
R7758 gnd.n7605 gnd.n135 26.7676
R7759 gnd.n7599 gnd.n146 26.7676
R7760 gnd.n7362 gnd.n153 26.7676
R7761 gnd.n7371 gnd.n163 26.7676
R7762 gnd.n2889 gnd.t233 26.4489
R7763 gnd.n4435 gnd.t22 26.4489
R7764 gnd.n2834 gnd.t6 25.8116
R7765 gnd.n7611 gnd.t259 25.8116
R7766 gnd.n2516 gnd.n2515 25.7944
R7767 gnd.n3774 gnd.n3773 25.7944
R7768 gnd.n5644 gnd.n5643 25.7944
R7769 gnd.n5078 gnd.n5077 25.7944
R7770 gnd.n2523 gnd.n2522 25.7944
R7771 gnd.n4218 gnd.n4217 25.7944
R7772 gnd.n4270 gnd.n4269 25.7944
R7773 gnd.n1811 gnd.n1810 25.7944
R7774 gnd.n314 gnd.n313 25.7944
R7775 gnd.n281 gnd.n280 25.7944
R7776 gnd.n7521 gnd.n7520 25.7944
R7777 gnd.n351 gnd.n350 25.7944
R7778 gnd.n1091 gnd.n1090 25.7944
R7779 gnd.n1113 gnd.n1112 25.7944
R7780 gnd.n1135 gnd.n1134 25.7944
R7781 gnd.n2688 gnd.n2687 25.7944
R7782 gnd.n1410 gnd.n1409 25.7944
R7783 gnd.n2349 gnd.n2348 25.7944
R7784 gnd.n2371 gnd.n2370 25.7944
R7785 gnd.n3764 gnd.n3763 25.7944
R7786 gnd.n2766 gnd.t18 25.1743
R7787 gnd.n7587 gnd.t38 25.1743
R7788 gnd.n5688 gnd.n5408 24.8557
R7789 gnd.n5411 gnd.n5402 24.8557
R7790 gnd.n5709 gnd.n5387 24.8557
R7791 gnd.n5728 gnd.n5727 24.8557
R7792 gnd.n5738 gnd.n5380 24.8557
R7793 gnd.n5751 gnd.n5368 24.8557
R7794 gnd.n5776 gnd.n5352 24.8557
R7795 gnd.n5775 gnd.n5354 24.8557
R7796 gnd.n5798 gnd.n5336 24.8557
R7797 gnd.n5787 gnd.n5328 24.8557
R7798 gnd.n5823 gnd.n5822 24.8557
R7799 gnd.n5833 gnd.n5321 24.8557
R7800 gnd.n5845 gnd.n5313 24.8557
R7801 gnd.n5844 gnd.n5301 24.8557
R7802 gnd.n5863 gnd.n5862 24.8557
R7803 gnd.n5884 gnd.n5282 24.8557
R7804 gnd.n5908 gnd.n5907 24.8557
R7805 gnd.n5919 gnd.n5201 24.8557
R7806 gnd.n5918 gnd.n5203 24.8557
R7807 gnd.n5930 gnd.n5194 24.8557
R7808 gnd.n5947 gnd.n5946 24.8557
R7809 gnd.n5185 gnd.n5174 24.8557
R7810 gnd.n5970 gnd.n5164 24.8557
R7811 gnd.n5166 gnd.n5165 24.8557
R7812 gnd.n5993 gnd.n5158 24.8557
R7813 gnd.n6004 gnd.n6003 24.8557
R7814 gnd.n6018 gnd.n5145 24.8557
R7815 gnd.n6456 gnd.n979 24.8557
R7816 gnd.n6319 gnd.n990 24.8557
R7817 gnd.n6449 gnd.n6448 24.8557
R7818 gnd.n6442 gnd.n1002 24.8557
R7819 gnd.n6441 gnd.n1005 24.8557
R7820 gnd.n6308 gnd.n1016 24.8557
R7821 gnd.n6428 gnd.n1027 24.8557
R7822 gnd.n6464 gnd.n6463 23.7886
R7823 gnd.n5706 gnd.t252 23.2624
R7824 gnd.n5698 gnd.t151 22.6251
R7825 gnd.n4922 gnd.t93 22.6251
R7826 gnd.t200 gnd.n1197 22.6251
R7827 gnd.n3021 gnd.t111 22.6251
R7828 gnd.n3754 gnd.t89 22.6251
R7829 gnd.n362 gnd.t241 22.6251
R7830 gnd.n209 gnd.t103 22.6251
R7831 gnd.t4 gnd.n1238 21.9878
R7832 gnd.n374 gnd.t46 21.9878
R7833 gnd.n5678 gnd.t221 21.3504
R7834 gnd.n2877 gnd.t24 21.3504
R7835 gnd.t8 gnd.n4470 21.3504
R7836 gnd.n5983 gnd.t295 20.7131
R7837 gnd.t48 gnd.n1286 20.7131
R7838 gnd.t20 gnd.n1694 20.7131
R7839 gnd.n3054 gnd.n1381 20.3945
R7840 gnd.n1599 gnd.n1591 20.3945
R7841 gnd.t293 gnd.n5175 20.0758
R7842 gnd.t61 gnd.n1326 20.0758
R7843 gnd.t44 gnd.n1654 20.0758
R7844 gnd.n2189 gnd.n2188 19.9763
R7845 gnd.n1880 gnd.n1879 19.9763
R7846 gnd.n4669 gnd.n4668 19.9763
R7847 gnd.n4012 gnd.n4011 19.9763
R7848 gnd.n1473 gnd.t79 19.8005
R7849 gnd.n1473 gnd.t129 19.8005
R7850 gnd.n1472 gnd.t196 19.8005
R7851 gnd.n1472 gnd.t159 19.8005
R7852 gnd.n4002 gnd.t98 19.8005
R7853 gnd.n4002 gnd.t171 19.8005
R7854 gnd.n4001 gnd.t149 19.8005
R7855 gnd.n4001 gnd.t187 19.8005
R7856 gnd.n1469 gnd.n1468 19.5087
R7857 gnd.n1482 gnd.n1469 19.5087
R7858 gnd.n1480 gnd.n1471 19.5087
R7859 gnd.n4006 gnd.n4000 19.5087
R7860 gnd.t318 gnd.n5210 19.4385
R7861 gnd.n3146 gnd.n2329 19.3944
R7862 gnd.n3151 gnd.n2329 19.3944
R7863 gnd.n3151 gnd.n2330 19.3944
R7864 gnd.n2330 gnd.n2306 19.3944
R7865 gnd.n3176 gnd.n2306 19.3944
R7866 gnd.n3176 gnd.n2303 19.3944
R7867 gnd.n3181 gnd.n2303 19.3944
R7868 gnd.n3181 gnd.n2304 19.3944
R7869 gnd.n2304 gnd.n2282 19.3944
R7870 gnd.n3206 gnd.n2282 19.3944
R7871 gnd.n3206 gnd.n2279 19.3944
R7872 gnd.n3211 gnd.n2279 19.3944
R7873 gnd.n3211 gnd.n2280 19.3944
R7874 gnd.n2280 gnd.n2257 19.3944
R7875 gnd.n3246 gnd.n2257 19.3944
R7876 gnd.n3246 gnd.n2254 19.3944
R7877 gnd.n3254 gnd.n2254 19.3944
R7878 gnd.n3254 gnd.n2255 19.3944
R7879 gnd.n3250 gnd.n2255 19.3944
R7880 gnd.n3250 gnd.n2173 19.3944
R7881 gnd.n3302 gnd.n2173 19.3944
R7882 gnd.n3302 gnd.n2170 19.3944
R7883 gnd.n3326 gnd.n2170 19.3944
R7884 gnd.n3326 gnd.n2171 19.3944
R7885 gnd.n3322 gnd.n2171 19.3944
R7886 gnd.n3322 gnd.n3321 19.3944
R7887 gnd.n3321 gnd.n3320 19.3944
R7888 gnd.n3320 gnd.n3312 19.3944
R7889 gnd.n3316 gnd.n3312 19.3944
R7890 gnd.n3316 gnd.n3315 19.3944
R7891 gnd.n3315 gnd.n2123 19.3944
R7892 gnd.n2123 gnd.n2121 19.3944
R7893 gnd.n3404 gnd.n2121 19.3944
R7894 gnd.n3404 gnd.n2119 19.3944
R7895 gnd.n3408 gnd.n2119 19.3944
R7896 gnd.n3408 gnd.n2094 19.3944
R7897 gnd.n3456 gnd.n2094 19.3944
R7898 gnd.n3456 gnd.n2095 19.3944
R7899 gnd.n3452 gnd.n2095 19.3944
R7900 gnd.n3452 gnd.n2071 19.3944
R7901 gnd.n3514 gnd.n2071 19.3944
R7902 gnd.n3514 gnd.n2072 19.3944
R7903 gnd.n3510 gnd.n2072 19.3944
R7904 gnd.n3510 gnd.n3509 19.3944
R7905 gnd.n3509 gnd.n3508 19.3944
R7906 gnd.n3508 gnd.n3495 19.3944
R7907 gnd.n3504 gnd.n3495 19.3944
R7908 gnd.n3504 gnd.n3503 19.3944
R7909 gnd.n3503 gnd.n3502 19.3944
R7910 gnd.n3502 gnd.n2013 19.3944
R7911 gnd.n3622 gnd.n2013 19.3944
R7912 gnd.n3622 gnd.n2010 19.3944
R7913 gnd.n3627 gnd.n2010 19.3944
R7914 gnd.n3627 gnd.n2011 19.3944
R7915 gnd.n2011 gnd.n1984 19.3944
R7916 gnd.n3661 gnd.n1984 19.3944
R7917 gnd.n3661 gnd.n1981 19.3944
R7918 gnd.n3672 gnd.n1981 19.3944
R7919 gnd.n3672 gnd.n1982 19.3944
R7920 gnd.n3668 gnd.n1982 19.3944
R7921 gnd.n3668 gnd.n3667 19.3944
R7922 gnd.n3667 gnd.n1949 19.3944
R7923 gnd.n3718 gnd.n1949 19.3944
R7924 gnd.n3718 gnd.n1947 19.3944
R7925 gnd.n3722 gnd.n1947 19.3944
R7926 gnd.n3725 gnd.n3722 19.3944
R7927 gnd.n3726 gnd.n3725 19.3944
R7928 gnd.n3726 gnd.n1945 19.3944
R7929 gnd.n3730 gnd.n1945 19.3944
R7930 gnd.n3733 gnd.n3730 19.3944
R7931 gnd.n3734 gnd.n3733 19.3944
R7932 gnd.n3734 gnd.n1943 19.3944
R7933 gnd.n3738 gnd.n1943 19.3944
R7934 gnd.n3741 gnd.n3738 19.3944
R7935 gnd.n3742 gnd.n3741 19.3944
R7936 gnd.n3742 gnd.n1941 19.3944
R7937 gnd.n3746 gnd.n1941 19.3944
R7938 gnd.n3749 gnd.n3746 19.3944
R7939 gnd.n3750 gnd.n3749 19.3944
R7940 gnd.n3750 gnd.n1938 19.3944
R7941 gnd.n3933 gnd.n1938 19.3944
R7942 gnd.n3933 gnd.n1939 19.3944
R7943 gnd.n2549 gnd.n2528 19.3944
R7944 gnd.n3074 gnd.n2528 19.3944
R7945 gnd.n3074 gnd.n3073 19.3944
R7946 gnd.n3138 gnd.n3137 19.3944
R7947 gnd.n3137 gnd.n3136 19.3944
R7948 gnd.n3136 gnd.n2341 19.3944
R7949 gnd.n3132 gnd.n2341 19.3944
R7950 gnd.n3132 gnd.n3131 19.3944
R7951 gnd.n3131 gnd.n3130 19.3944
R7952 gnd.n3130 gnd.n2346 19.3944
R7953 gnd.n3125 gnd.n2346 19.3944
R7954 gnd.n3125 gnd.n3124 19.3944
R7955 gnd.n3124 gnd.n2463 19.3944
R7956 gnd.n3117 gnd.n2463 19.3944
R7957 gnd.n3117 gnd.n3116 19.3944
R7958 gnd.n3116 gnd.n2473 19.3944
R7959 gnd.n3109 gnd.n2473 19.3944
R7960 gnd.n3109 gnd.n3108 19.3944
R7961 gnd.n3108 gnd.n2483 19.3944
R7962 gnd.n3101 gnd.n2483 19.3944
R7963 gnd.n3101 gnd.n3100 19.3944
R7964 gnd.n3100 gnd.n2494 19.3944
R7965 gnd.n3093 gnd.n2494 19.3944
R7966 gnd.n3093 gnd.n3092 19.3944
R7967 gnd.n3092 gnd.n2504 19.3944
R7968 gnd.n3085 gnd.n2504 19.3944
R7969 gnd.n3085 gnd.n3084 19.3944
R7970 gnd.n3841 gnd.n3804 19.3944
R7971 gnd.n3854 gnd.n3804 19.3944
R7972 gnd.n3854 gnd.n3802 19.3944
R7973 gnd.n3860 gnd.n3802 19.3944
R7974 gnd.n3860 gnd.n3795 19.3944
R7975 gnd.n3873 gnd.n3795 19.3944
R7976 gnd.n3873 gnd.n3793 19.3944
R7977 gnd.n3879 gnd.n3793 19.3944
R7978 gnd.n3879 gnd.n3786 19.3944
R7979 gnd.n3892 gnd.n3786 19.3944
R7980 gnd.n3892 gnd.n3784 19.3944
R7981 gnd.n3898 gnd.n3784 19.3944
R7982 gnd.n3898 gnd.n3777 19.3944
R7983 gnd.n3912 gnd.n3777 19.3944
R7984 gnd.n3912 gnd.n3775 19.3944
R7985 gnd.n3918 gnd.n3775 19.3944
R7986 gnd.n5551 gnd.n5550 19.3944
R7987 gnd.n5550 gnd.n5460 19.3944
R7988 gnd.n5545 gnd.n5460 19.3944
R7989 gnd.n5545 gnd.n5544 19.3944
R7990 gnd.n5544 gnd.n5465 19.3944
R7991 gnd.n5539 gnd.n5465 19.3944
R7992 gnd.n5539 gnd.n5538 19.3944
R7993 gnd.n5538 gnd.n5537 19.3944
R7994 gnd.n5537 gnd.n5471 19.3944
R7995 gnd.n5531 gnd.n5471 19.3944
R7996 gnd.n5531 gnd.n5530 19.3944
R7997 gnd.n5530 gnd.n5529 19.3944
R7998 gnd.n5529 gnd.n5477 19.3944
R7999 gnd.n5523 gnd.n5477 19.3944
R8000 gnd.n5523 gnd.n5522 19.3944
R8001 gnd.n5522 gnd.n5521 19.3944
R8002 gnd.n5521 gnd.n5483 19.3944
R8003 gnd.n5515 gnd.n5483 19.3944
R8004 gnd.n5515 gnd.n5514 19.3944
R8005 gnd.n5514 gnd.n5513 19.3944
R8006 gnd.n5513 gnd.n5489 19.3944
R8007 gnd.n5507 gnd.n5489 19.3944
R8008 gnd.n5505 gnd.n5504 19.3944
R8009 gnd.n5504 gnd.n5499 19.3944
R8010 gnd.n5499 gnd.n5497 19.3944
R8011 gnd.n6348 gnd.n5125 19.3944
R8012 gnd.n6348 gnd.n6347 19.3944
R8013 gnd.n6347 gnd.n6346 19.3944
R8014 gnd.n6390 gnd.n6389 19.3944
R8015 gnd.n6389 gnd.n6388 19.3944
R8016 gnd.n6388 gnd.n5086 19.3944
R8017 gnd.n6383 gnd.n5086 19.3944
R8018 gnd.n6383 gnd.n6382 19.3944
R8019 gnd.n6382 gnd.n6381 19.3944
R8020 gnd.n6381 gnd.n5093 19.3944
R8021 gnd.n6376 gnd.n5093 19.3944
R8022 gnd.n6376 gnd.n6375 19.3944
R8023 gnd.n6375 gnd.n6374 19.3944
R8024 gnd.n6374 gnd.n5100 19.3944
R8025 gnd.n6369 gnd.n5100 19.3944
R8026 gnd.n6369 gnd.n6368 19.3944
R8027 gnd.n6368 gnd.n6367 19.3944
R8028 gnd.n6367 gnd.n5107 19.3944
R8029 gnd.n6362 gnd.n5107 19.3944
R8030 gnd.n6362 gnd.n6361 19.3944
R8031 gnd.n6361 gnd.n6360 19.3944
R8032 gnd.n6360 gnd.n5114 19.3944
R8033 gnd.n6355 gnd.n5114 19.3944
R8034 gnd.n6355 gnd.n6354 19.3944
R8035 gnd.n6354 gnd.n6353 19.3944
R8036 gnd.n5691 gnd.n5690 19.3944
R8037 gnd.n5692 gnd.n5691 19.3944
R8038 gnd.n5692 gnd.n5401 19.3944
R8039 gnd.n5401 gnd.n5395 19.3944
R8040 gnd.n5717 gnd.n5395 19.3944
R8041 gnd.n5718 gnd.n5717 19.3944
R8042 gnd.n5718 gnd.n5378 19.3944
R8043 gnd.n5378 gnd.n5376 19.3944
R8044 gnd.n5742 gnd.n5376 19.3944
R8045 gnd.n5745 gnd.n5742 19.3944
R8046 gnd.n5745 gnd.n5744 19.3944
R8047 gnd.n5744 gnd.n5348 19.3944
R8048 gnd.n5783 gnd.n5348 19.3944
R8049 gnd.n5783 gnd.n5346 19.3944
R8050 gnd.n5789 gnd.n5346 19.3944
R8051 gnd.n5790 gnd.n5789 19.3944
R8052 gnd.n5790 gnd.n5316 19.3944
R8053 gnd.n5840 gnd.n5316 19.3944
R8054 gnd.n5841 gnd.n5840 19.3944
R8055 gnd.n5841 gnd.n5309 19.3944
R8056 gnd.n5852 gnd.n5309 19.3944
R8057 gnd.n5853 gnd.n5852 19.3944
R8058 gnd.n5853 gnd.n5292 19.3944
R8059 gnd.n5292 gnd.n5290 19.3944
R8060 gnd.n5877 gnd.n5290 19.3944
R8061 gnd.n5878 gnd.n5877 19.3944
R8062 gnd.n5878 gnd.n5197 19.3944
R8063 gnd.n5925 gnd.n5197 19.3944
R8064 gnd.n5926 gnd.n5925 19.3944
R8065 gnd.n5926 gnd.n5190 19.3944
R8066 gnd.n5937 gnd.n5190 19.3944
R8067 gnd.n5938 gnd.n5937 19.3944
R8068 gnd.n5938 gnd.n5173 19.3944
R8069 gnd.n5173 gnd.n5171 19.3944
R8070 gnd.n5965 gnd.n5171 19.3944
R8071 gnd.n5965 gnd.n5154 19.3944
R8072 gnd.n5999 gnd.n5154 19.3944
R8073 gnd.n6000 gnd.n5999 19.3944
R8074 gnd.n6000 gnd.n5140 19.3944
R8075 gnd.n6026 gnd.n5140 19.3944
R8076 gnd.n6026 gnd.n5137 19.3944
R8077 gnd.n6030 gnd.n5137 19.3944
R8078 gnd.n6031 gnd.n6030 19.3944
R8079 gnd.n6317 gnd.n6031 19.3944
R8080 gnd.n6317 gnd.n6316 19.3944
R8081 gnd.n6316 gnd.n6315 19.3944
R8082 gnd.n6315 gnd.n6312 19.3944
R8083 gnd.n6312 gnd.n6311 19.3944
R8084 gnd.n6311 gnd.n6310 19.3944
R8085 gnd.n6310 gnd.n6307 19.3944
R8086 gnd.n6307 gnd.n6306 19.3944
R8087 gnd.n6306 gnd.n6303 19.3944
R8088 gnd.n6303 gnd.n6302 19.3944
R8089 gnd.n5674 gnd.n5673 19.3944
R8090 gnd.n5673 gnd.n5672 19.3944
R8091 gnd.n5672 gnd.n5671 19.3944
R8092 gnd.n5671 gnd.n5669 19.3944
R8093 gnd.n5669 gnd.n5666 19.3944
R8094 gnd.n5666 gnd.n5665 19.3944
R8095 gnd.n5665 gnd.n5662 19.3944
R8096 gnd.n5662 gnd.n5661 19.3944
R8097 gnd.n5661 gnd.n5658 19.3944
R8098 gnd.n5658 gnd.n5657 19.3944
R8099 gnd.n5657 gnd.n5654 19.3944
R8100 gnd.n5654 gnd.n5653 19.3944
R8101 gnd.n5653 gnd.n5650 19.3944
R8102 gnd.n5650 gnd.n5649 19.3944
R8103 gnd.n5700 gnd.n5406 19.3944
R8104 gnd.n5700 gnd.n5404 19.3944
R8105 gnd.n5704 gnd.n5404 19.3944
R8106 gnd.n5704 gnd.n5385 19.3944
R8107 gnd.n5730 gnd.n5385 19.3944
R8108 gnd.n5730 gnd.n5383 19.3944
R8109 gnd.n5736 gnd.n5383 19.3944
R8110 gnd.n5736 gnd.n5735 19.3944
R8111 gnd.n5735 gnd.n5359 19.3944
R8112 gnd.n5764 gnd.n5359 19.3944
R8113 gnd.n5764 gnd.n5357 19.3944
R8114 gnd.n5773 gnd.n5357 19.3944
R8115 gnd.n5773 gnd.n5772 19.3944
R8116 gnd.n5772 gnd.n5771 19.3944
R8117 gnd.n5771 gnd.n5326 19.3944
R8118 gnd.n5825 gnd.n5326 19.3944
R8119 gnd.n5825 gnd.n5324 19.3944
R8120 gnd.n5831 gnd.n5324 19.3944
R8121 gnd.n5831 gnd.n5830 19.3944
R8122 gnd.n5830 gnd.n5299 19.3944
R8123 gnd.n5865 gnd.n5299 19.3944
R8124 gnd.n5865 gnd.n5297 19.3944
R8125 gnd.n5871 gnd.n5297 19.3944
R8126 gnd.n5871 gnd.n5870 19.3944
R8127 gnd.n5870 gnd.n5208 19.3944
R8128 gnd.n5910 gnd.n5208 19.3944
R8129 gnd.n5910 gnd.n5206 19.3944
R8130 gnd.n5916 gnd.n5206 19.3944
R8131 gnd.n5916 gnd.n5915 19.3944
R8132 gnd.n5915 gnd.n5180 19.3944
R8133 gnd.n5949 gnd.n5180 19.3944
R8134 gnd.n5949 gnd.n5178 19.3944
R8135 gnd.n5958 gnd.n5178 19.3944
R8136 gnd.n5958 gnd.n5957 19.3944
R8137 gnd.n5957 gnd.n5956 19.3944
R8138 gnd.n5956 gnd.n5150 19.3944
R8139 gnd.n6006 gnd.n5150 19.3944
R8140 gnd.n6006 gnd.n5148 19.3944
R8141 gnd.n6016 gnd.n5148 19.3944
R8142 gnd.n6016 gnd.n6015 19.3944
R8143 gnd.n6015 gnd.n6014 19.3944
R8144 gnd.n6014 gnd.n984 19.3944
R8145 gnd.n6453 gnd.n984 19.3944
R8146 gnd.n6453 gnd.n6452 19.3944
R8147 gnd.n6452 gnd.n6451 19.3944
R8148 gnd.n6451 gnd.n988 19.3944
R8149 gnd.n1008 gnd.n988 19.3944
R8150 gnd.n6439 gnd.n1008 19.3944
R8151 gnd.n6439 gnd.n6438 19.3944
R8152 gnd.n6438 gnd.n6437 19.3944
R8153 gnd.n6437 gnd.n1014 19.3944
R8154 gnd.n5050 gnd.n1014 19.3944
R8155 gnd.n6425 gnd.n5050 19.3944
R8156 gnd.n6422 gnd.n6421 19.3944
R8157 gnd.n6421 gnd.n6420 19.3944
R8158 gnd.n6420 gnd.n5056 19.3944
R8159 gnd.n6415 gnd.n5056 19.3944
R8160 gnd.n6415 gnd.n6414 19.3944
R8161 gnd.n6414 gnd.n6413 19.3944
R8162 gnd.n6413 gnd.n5063 19.3944
R8163 gnd.n6408 gnd.n5063 19.3944
R8164 gnd.n6408 gnd.n6407 19.3944
R8165 gnd.n6407 gnd.n6406 19.3944
R8166 gnd.n6406 gnd.n5070 19.3944
R8167 gnd.n6401 gnd.n5070 19.3944
R8168 gnd.n6401 gnd.n6400 19.3944
R8169 gnd.n6400 gnd.n6399 19.3944
R8170 gnd.n5558 gnd.n5454 19.3944
R8171 gnd.n5562 gnd.n5454 19.3944
R8172 gnd.n5562 gnd.n5444 19.3944
R8173 gnd.n5574 gnd.n5444 19.3944
R8174 gnd.n5574 gnd.n5442 19.3944
R8175 gnd.n5578 gnd.n5442 19.3944
R8176 gnd.n5578 gnd.n5431 19.3944
R8177 gnd.n5590 gnd.n5431 19.3944
R8178 gnd.n5590 gnd.n5429 19.3944
R8179 gnd.n5616 gnd.n5429 19.3944
R8180 gnd.n5616 gnd.n5615 19.3944
R8181 gnd.n5615 gnd.n5614 19.3944
R8182 gnd.n5614 gnd.n5613 19.3944
R8183 gnd.n5613 gnd.n5611 19.3944
R8184 gnd.n5611 gnd.n5610 19.3944
R8185 gnd.n5610 gnd.n5608 19.3944
R8186 gnd.n5608 gnd.n5607 19.3944
R8187 gnd.n5607 gnd.n5605 19.3944
R8188 gnd.n5605 gnd.n5604 19.3944
R8189 gnd.n5604 gnd.n5366 19.3944
R8190 gnd.n5753 gnd.n5366 19.3944
R8191 gnd.n5753 gnd.n5364 19.3944
R8192 gnd.n5759 gnd.n5364 19.3944
R8193 gnd.n5759 gnd.n5758 19.3944
R8194 gnd.n5758 gnd.n5333 19.3944
R8195 gnd.n5800 gnd.n5333 19.3944
R8196 gnd.n5800 gnd.n5331 19.3944
R8197 gnd.n5804 gnd.n5331 19.3944
R8198 gnd.n5818 gnd.n5804 19.3944
R8199 gnd.n5816 gnd.n5815 19.3944
R8200 gnd.n5812 gnd.n5811 19.3944
R8201 gnd.n5808 gnd.n5807 19.3944
R8202 gnd.n5886 gnd.n5280 19.3944
R8203 gnd.n5886 gnd.n5214 19.3944
R8204 gnd.n5905 gnd.n5214 19.3944
R8205 gnd.n5905 gnd.n5904 19.3944
R8206 gnd.n5904 gnd.n5903 19.3944
R8207 gnd.n5903 gnd.n5901 19.3944
R8208 gnd.n5901 gnd.n5900 19.3944
R8209 gnd.n5900 gnd.n5898 19.3944
R8210 gnd.n5898 gnd.n5897 19.3944
R8211 gnd.n5897 gnd.n5162 19.3944
R8212 gnd.n5972 gnd.n5162 19.3944
R8213 gnd.n5972 gnd.n5160 19.3944
R8214 gnd.n5991 gnd.n5160 19.3944
R8215 gnd.n5991 gnd.n5990 19.3944
R8216 gnd.n5990 gnd.n5989 19.3944
R8217 gnd.n5989 gnd.n5988 19.3944
R8218 gnd.n5988 gnd.n5986 19.3944
R8219 gnd.n5986 gnd.n5985 19.3944
R8220 gnd.n5985 gnd.n5982 19.3944
R8221 gnd.n5982 gnd.n5135 19.3944
R8222 gnd.n6323 gnd.n5135 19.3944
R8223 gnd.n6323 gnd.n5133 19.3944
R8224 gnd.n6329 gnd.n5133 19.3944
R8225 gnd.n6330 gnd.n6329 19.3944
R8226 gnd.n6333 gnd.n6330 19.3944
R8227 gnd.n6333 gnd.n5131 19.3944
R8228 gnd.n6337 gnd.n5131 19.3944
R8229 gnd.n6340 gnd.n6337 19.3944
R8230 gnd.n6341 gnd.n6340 19.3944
R8231 gnd.n5554 gnd.n5450 19.3944
R8232 gnd.n5566 gnd.n5450 19.3944
R8233 gnd.n5566 gnd.n5448 19.3944
R8234 gnd.n5570 gnd.n5448 19.3944
R8235 gnd.n5570 gnd.n5438 19.3944
R8236 gnd.n5582 gnd.n5438 19.3944
R8237 gnd.n5582 gnd.n5436 19.3944
R8238 gnd.n5586 gnd.n5436 19.3944
R8239 gnd.n5586 gnd.n5425 19.3944
R8240 gnd.n5680 gnd.n5425 19.3944
R8241 gnd.n5680 gnd.n5422 19.3944
R8242 gnd.n5685 gnd.n5422 19.3944
R8243 gnd.n5685 gnd.n5413 19.3944
R8244 gnd.n5695 gnd.n5413 19.3944
R8245 gnd.n5695 gnd.n5397 19.3944
R8246 gnd.n5712 gnd.n5397 19.3944
R8247 gnd.n5712 gnd.n5393 19.3944
R8248 gnd.n5725 gnd.n5393 19.3944
R8249 gnd.n5725 gnd.n5724 19.3944
R8250 gnd.n5724 gnd.n5372 19.3944
R8251 gnd.n5749 gnd.n5372 19.3944
R8252 gnd.n5749 gnd.n5748 19.3944
R8253 gnd.n5748 gnd.n5350 19.3944
R8254 gnd.n5778 gnd.n5350 19.3944
R8255 gnd.n5778 gnd.n5340 19.3944
R8256 gnd.n5796 gnd.n5340 19.3944
R8257 gnd.n5796 gnd.n5795 19.3944
R8258 gnd.n5795 gnd.n5794 19.3944
R8259 gnd.n5794 gnd.n5318 19.3944
R8260 gnd.n5836 gnd.n5318 19.3944
R8261 gnd.n5836 gnd.n5311 19.3944
R8262 gnd.n5847 gnd.n5311 19.3944
R8263 gnd.n5847 gnd.n5307 19.3944
R8264 gnd.n5860 gnd.n5307 19.3944
R8265 gnd.n5860 gnd.n5859 19.3944
R8266 gnd.n5859 gnd.n5286 19.3944
R8267 gnd.n5882 gnd.n5286 19.3944
R8268 gnd.n5882 gnd.n5881 19.3944
R8269 gnd.n5881 gnd.n5199 19.3944
R8270 gnd.n5921 gnd.n5199 19.3944
R8271 gnd.n5921 gnd.n5192 19.3944
R8272 gnd.n5932 gnd.n5192 19.3944
R8273 gnd.n5932 gnd.n5188 19.3944
R8274 gnd.n5944 gnd.n5188 19.3944
R8275 gnd.n5944 gnd.n5943 19.3944
R8276 gnd.n5943 gnd.n5168 19.3944
R8277 gnd.n5968 gnd.n5168 19.3944
R8278 gnd.n5968 gnd.n5156 19.3944
R8279 gnd.n5995 gnd.n5156 19.3944
R8280 gnd.n5995 gnd.n5142 19.3944
R8281 gnd.n6021 gnd.n5142 19.3944
R8282 gnd.n6021 gnd.n973 19.3944
R8283 gnd.n6460 gnd.n973 19.3944
R8284 gnd.n6460 gnd.n6459 19.3944
R8285 gnd.n6459 gnd.n6458 19.3944
R8286 gnd.n6458 gnd.n977 19.3944
R8287 gnd.n996 gnd.n977 19.3944
R8288 gnd.n6446 gnd.n996 19.3944
R8289 gnd.n6446 gnd.n6445 19.3944
R8290 gnd.n6445 gnd.n6444 19.3944
R8291 gnd.n6444 gnd.n1000 19.3944
R8292 gnd.n1022 gnd.n1000 19.3944
R8293 gnd.n6432 gnd.n1022 19.3944
R8294 gnd.n6432 gnd.n6431 19.3944
R8295 gnd.n6431 gnd.n6430 19.3944
R8296 gnd.n3121 gnd.n2465 19.3944
R8297 gnd.n3121 gnd.n3120 19.3944
R8298 gnd.n3120 gnd.n2469 19.3944
R8299 gnd.n3113 gnd.n2469 19.3944
R8300 gnd.n3113 gnd.n3112 19.3944
R8301 gnd.n3112 gnd.n2479 19.3944
R8302 gnd.n3105 gnd.n2479 19.3944
R8303 gnd.n3105 gnd.n3104 19.3944
R8304 gnd.n3104 gnd.n2490 19.3944
R8305 gnd.n3097 gnd.n2490 19.3944
R8306 gnd.n3097 gnd.n3096 19.3944
R8307 gnd.n3096 gnd.n2500 19.3944
R8308 gnd.n3089 gnd.n2500 19.3944
R8309 gnd.n3089 gnd.n3088 19.3944
R8310 gnd.n3088 gnd.n2511 19.3944
R8311 gnd.n3081 gnd.n2511 19.3944
R8312 gnd.n7089 gnd.n527 19.3944
R8313 gnd.n7089 gnd.n523 19.3944
R8314 gnd.n7095 gnd.n523 19.3944
R8315 gnd.n7095 gnd.n521 19.3944
R8316 gnd.n7099 gnd.n521 19.3944
R8317 gnd.n7099 gnd.n517 19.3944
R8318 gnd.n7105 gnd.n517 19.3944
R8319 gnd.n7105 gnd.n515 19.3944
R8320 gnd.n7109 gnd.n515 19.3944
R8321 gnd.n7109 gnd.n511 19.3944
R8322 gnd.n7115 gnd.n511 19.3944
R8323 gnd.n7115 gnd.n509 19.3944
R8324 gnd.n7119 gnd.n509 19.3944
R8325 gnd.n7119 gnd.n505 19.3944
R8326 gnd.n7125 gnd.n505 19.3944
R8327 gnd.n7125 gnd.n503 19.3944
R8328 gnd.n7129 gnd.n503 19.3944
R8329 gnd.n7129 gnd.n499 19.3944
R8330 gnd.n7135 gnd.n499 19.3944
R8331 gnd.n7135 gnd.n497 19.3944
R8332 gnd.n7139 gnd.n497 19.3944
R8333 gnd.n7139 gnd.n493 19.3944
R8334 gnd.n7145 gnd.n493 19.3944
R8335 gnd.n7145 gnd.n491 19.3944
R8336 gnd.n7149 gnd.n491 19.3944
R8337 gnd.n7149 gnd.n487 19.3944
R8338 gnd.n7155 gnd.n487 19.3944
R8339 gnd.n7155 gnd.n485 19.3944
R8340 gnd.n7159 gnd.n485 19.3944
R8341 gnd.n7159 gnd.n481 19.3944
R8342 gnd.n7165 gnd.n481 19.3944
R8343 gnd.n7165 gnd.n479 19.3944
R8344 gnd.n7169 gnd.n479 19.3944
R8345 gnd.n7169 gnd.n475 19.3944
R8346 gnd.n7175 gnd.n475 19.3944
R8347 gnd.n7175 gnd.n473 19.3944
R8348 gnd.n7179 gnd.n473 19.3944
R8349 gnd.n7179 gnd.n469 19.3944
R8350 gnd.n7185 gnd.n469 19.3944
R8351 gnd.n7185 gnd.n467 19.3944
R8352 gnd.n7189 gnd.n467 19.3944
R8353 gnd.n7189 gnd.n463 19.3944
R8354 gnd.n7195 gnd.n463 19.3944
R8355 gnd.n7195 gnd.n461 19.3944
R8356 gnd.n7199 gnd.n461 19.3944
R8357 gnd.n7199 gnd.n457 19.3944
R8358 gnd.n7205 gnd.n457 19.3944
R8359 gnd.n7205 gnd.n455 19.3944
R8360 gnd.n7209 gnd.n455 19.3944
R8361 gnd.n7209 gnd.n451 19.3944
R8362 gnd.n7215 gnd.n451 19.3944
R8363 gnd.n7215 gnd.n449 19.3944
R8364 gnd.n7219 gnd.n449 19.3944
R8365 gnd.n7219 gnd.n445 19.3944
R8366 gnd.n7225 gnd.n445 19.3944
R8367 gnd.n7225 gnd.n443 19.3944
R8368 gnd.n7229 gnd.n443 19.3944
R8369 gnd.n7229 gnd.n439 19.3944
R8370 gnd.n7235 gnd.n439 19.3944
R8371 gnd.n7235 gnd.n437 19.3944
R8372 gnd.n7239 gnd.n437 19.3944
R8373 gnd.n7239 gnd.n433 19.3944
R8374 gnd.n7245 gnd.n433 19.3944
R8375 gnd.n7245 gnd.n431 19.3944
R8376 gnd.n7249 gnd.n431 19.3944
R8377 gnd.n7249 gnd.n427 19.3944
R8378 gnd.n7255 gnd.n427 19.3944
R8379 gnd.n7255 gnd.n425 19.3944
R8380 gnd.n7259 gnd.n425 19.3944
R8381 gnd.n7259 gnd.n421 19.3944
R8382 gnd.n7265 gnd.n421 19.3944
R8383 gnd.n7265 gnd.n419 19.3944
R8384 gnd.n7269 gnd.n419 19.3944
R8385 gnd.n7269 gnd.n415 19.3944
R8386 gnd.n7275 gnd.n415 19.3944
R8387 gnd.n7275 gnd.n413 19.3944
R8388 gnd.n7279 gnd.n413 19.3944
R8389 gnd.n7279 gnd.n409 19.3944
R8390 gnd.n7285 gnd.n409 19.3944
R8391 gnd.n7285 gnd.n407 19.3944
R8392 gnd.n7291 gnd.n407 19.3944
R8393 gnd.n7291 gnd.n7290 19.3944
R8394 gnd.n7290 gnd.n403 19.3944
R8395 gnd.n7298 gnd.n403 19.3944
R8396 gnd.n6635 gnd.n799 19.3944
R8397 gnd.n6635 gnd.n797 19.3944
R8398 gnd.n6639 gnd.n797 19.3944
R8399 gnd.n6639 gnd.n793 19.3944
R8400 gnd.n6645 gnd.n793 19.3944
R8401 gnd.n6645 gnd.n791 19.3944
R8402 gnd.n6649 gnd.n791 19.3944
R8403 gnd.n6649 gnd.n787 19.3944
R8404 gnd.n6655 gnd.n787 19.3944
R8405 gnd.n6655 gnd.n785 19.3944
R8406 gnd.n6659 gnd.n785 19.3944
R8407 gnd.n6659 gnd.n781 19.3944
R8408 gnd.n6665 gnd.n781 19.3944
R8409 gnd.n6665 gnd.n779 19.3944
R8410 gnd.n6669 gnd.n779 19.3944
R8411 gnd.n6669 gnd.n775 19.3944
R8412 gnd.n6675 gnd.n775 19.3944
R8413 gnd.n6675 gnd.n773 19.3944
R8414 gnd.n6679 gnd.n773 19.3944
R8415 gnd.n6679 gnd.n769 19.3944
R8416 gnd.n6685 gnd.n769 19.3944
R8417 gnd.n6685 gnd.n767 19.3944
R8418 gnd.n6689 gnd.n767 19.3944
R8419 gnd.n6689 gnd.n763 19.3944
R8420 gnd.n6695 gnd.n763 19.3944
R8421 gnd.n6695 gnd.n761 19.3944
R8422 gnd.n6699 gnd.n761 19.3944
R8423 gnd.n6699 gnd.n757 19.3944
R8424 gnd.n6705 gnd.n757 19.3944
R8425 gnd.n6705 gnd.n755 19.3944
R8426 gnd.n6709 gnd.n755 19.3944
R8427 gnd.n6709 gnd.n751 19.3944
R8428 gnd.n6715 gnd.n751 19.3944
R8429 gnd.n6715 gnd.n749 19.3944
R8430 gnd.n6719 gnd.n749 19.3944
R8431 gnd.n6719 gnd.n745 19.3944
R8432 gnd.n6725 gnd.n745 19.3944
R8433 gnd.n6725 gnd.n743 19.3944
R8434 gnd.n6729 gnd.n743 19.3944
R8435 gnd.n6729 gnd.n739 19.3944
R8436 gnd.n6735 gnd.n739 19.3944
R8437 gnd.n6735 gnd.n737 19.3944
R8438 gnd.n6739 gnd.n737 19.3944
R8439 gnd.n6739 gnd.n733 19.3944
R8440 gnd.n6745 gnd.n733 19.3944
R8441 gnd.n6745 gnd.n731 19.3944
R8442 gnd.n6749 gnd.n731 19.3944
R8443 gnd.n6749 gnd.n727 19.3944
R8444 gnd.n6755 gnd.n727 19.3944
R8445 gnd.n6755 gnd.n725 19.3944
R8446 gnd.n6759 gnd.n725 19.3944
R8447 gnd.n6759 gnd.n721 19.3944
R8448 gnd.n6765 gnd.n721 19.3944
R8449 gnd.n6765 gnd.n719 19.3944
R8450 gnd.n6769 gnd.n719 19.3944
R8451 gnd.n6769 gnd.n715 19.3944
R8452 gnd.n6775 gnd.n715 19.3944
R8453 gnd.n6775 gnd.n713 19.3944
R8454 gnd.n6779 gnd.n713 19.3944
R8455 gnd.n6779 gnd.n709 19.3944
R8456 gnd.n6785 gnd.n709 19.3944
R8457 gnd.n6785 gnd.n707 19.3944
R8458 gnd.n6789 gnd.n707 19.3944
R8459 gnd.n6789 gnd.n703 19.3944
R8460 gnd.n6795 gnd.n703 19.3944
R8461 gnd.n6795 gnd.n701 19.3944
R8462 gnd.n6799 gnd.n701 19.3944
R8463 gnd.n6799 gnd.n697 19.3944
R8464 gnd.n6805 gnd.n697 19.3944
R8465 gnd.n6805 gnd.n695 19.3944
R8466 gnd.n6809 gnd.n695 19.3944
R8467 gnd.n6809 gnd.n691 19.3944
R8468 gnd.n6815 gnd.n691 19.3944
R8469 gnd.n6815 gnd.n689 19.3944
R8470 gnd.n6819 gnd.n689 19.3944
R8471 gnd.n6819 gnd.n685 19.3944
R8472 gnd.n6825 gnd.n685 19.3944
R8473 gnd.n6825 gnd.n683 19.3944
R8474 gnd.n6829 gnd.n683 19.3944
R8475 gnd.n6829 gnd.n679 19.3944
R8476 gnd.n6835 gnd.n679 19.3944
R8477 gnd.n6835 gnd.n677 19.3944
R8478 gnd.n6839 gnd.n677 19.3944
R8479 gnd.n6839 gnd.n673 19.3944
R8480 gnd.n6845 gnd.n673 19.3944
R8481 gnd.n6845 gnd.n671 19.3944
R8482 gnd.n6849 gnd.n671 19.3944
R8483 gnd.n6849 gnd.n667 19.3944
R8484 gnd.n6855 gnd.n667 19.3944
R8485 gnd.n6855 gnd.n665 19.3944
R8486 gnd.n6859 gnd.n665 19.3944
R8487 gnd.n6859 gnd.n661 19.3944
R8488 gnd.n6865 gnd.n661 19.3944
R8489 gnd.n6865 gnd.n659 19.3944
R8490 gnd.n6869 gnd.n659 19.3944
R8491 gnd.n6869 gnd.n655 19.3944
R8492 gnd.n6875 gnd.n655 19.3944
R8493 gnd.n6875 gnd.n653 19.3944
R8494 gnd.n6879 gnd.n653 19.3944
R8495 gnd.n6879 gnd.n649 19.3944
R8496 gnd.n6885 gnd.n649 19.3944
R8497 gnd.n6885 gnd.n647 19.3944
R8498 gnd.n6889 gnd.n647 19.3944
R8499 gnd.n6889 gnd.n643 19.3944
R8500 gnd.n6895 gnd.n643 19.3944
R8501 gnd.n6895 gnd.n641 19.3944
R8502 gnd.n6899 gnd.n641 19.3944
R8503 gnd.n6899 gnd.n637 19.3944
R8504 gnd.n6905 gnd.n637 19.3944
R8505 gnd.n6905 gnd.n635 19.3944
R8506 gnd.n6909 gnd.n635 19.3944
R8507 gnd.n6909 gnd.n631 19.3944
R8508 gnd.n6915 gnd.n631 19.3944
R8509 gnd.n6915 gnd.n629 19.3944
R8510 gnd.n6919 gnd.n629 19.3944
R8511 gnd.n6919 gnd.n625 19.3944
R8512 gnd.n6925 gnd.n625 19.3944
R8513 gnd.n6925 gnd.n623 19.3944
R8514 gnd.n6929 gnd.n623 19.3944
R8515 gnd.n6929 gnd.n619 19.3944
R8516 gnd.n6935 gnd.n619 19.3944
R8517 gnd.n6935 gnd.n617 19.3944
R8518 gnd.n6939 gnd.n617 19.3944
R8519 gnd.n6939 gnd.n613 19.3944
R8520 gnd.n6945 gnd.n613 19.3944
R8521 gnd.n6945 gnd.n611 19.3944
R8522 gnd.n6949 gnd.n611 19.3944
R8523 gnd.n6949 gnd.n607 19.3944
R8524 gnd.n6955 gnd.n607 19.3944
R8525 gnd.n6955 gnd.n605 19.3944
R8526 gnd.n6959 gnd.n605 19.3944
R8527 gnd.n6959 gnd.n601 19.3944
R8528 gnd.n6965 gnd.n601 19.3944
R8529 gnd.n6965 gnd.n599 19.3944
R8530 gnd.n6969 gnd.n599 19.3944
R8531 gnd.n6969 gnd.n595 19.3944
R8532 gnd.n6975 gnd.n595 19.3944
R8533 gnd.n6975 gnd.n593 19.3944
R8534 gnd.n6979 gnd.n593 19.3944
R8535 gnd.n6979 gnd.n589 19.3944
R8536 gnd.n6985 gnd.n589 19.3944
R8537 gnd.n6985 gnd.n587 19.3944
R8538 gnd.n6989 gnd.n587 19.3944
R8539 gnd.n6989 gnd.n583 19.3944
R8540 gnd.n6995 gnd.n583 19.3944
R8541 gnd.n6995 gnd.n581 19.3944
R8542 gnd.n6999 gnd.n581 19.3944
R8543 gnd.n6999 gnd.n577 19.3944
R8544 gnd.n7005 gnd.n577 19.3944
R8545 gnd.n7005 gnd.n575 19.3944
R8546 gnd.n7009 gnd.n575 19.3944
R8547 gnd.n7009 gnd.n571 19.3944
R8548 gnd.n7015 gnd.n571 19.3944
R8549 gnd.n7015 gnd.n569 19.3944
R8550 gnd.n7019 gnd.n569 19.3944
R8551 gnd.n7019 gnd.n565 19.3944
R8552 gnd.n7025 gnd.n565 19.3944
R8553 gnd.n7025 gnd.n563 19.3944
R8554 gnd.n7029 gnd.n563 19.3944
R8555 gnd.n7029 gnd.n559 19.3944
R8556 gnd.n7035 gnd.n559 19.3944
R8557 gnd.n7035 gnd.n557 19.3944
R8558 gnd.n7039 gnd.n557 19.3944
R8559 gnd.n7039 gnd.n553 19.3944
R8560 gnd.n7045 gnd.n553 19.3944
R8561 gnd.n7045 gnd.n551 19.3944
R8562 gnd.n7049 gnd.n551 19.3944
R8563 gnd.n7049 gnd.n547 19.3944
R8564 gnd.n7055 gnd.n547 19.3944
R8565 gnd.n7055 gnd.n545 19.3944
R8566 gnd.n7059 gnd.n545 19.3944
R8567 gnd.n7059 gnd.n541 19.3944
R8568 gnd.n7065 gnd.n541 19.3944
R8569 gnd.n7065 gnd.n539 19.3944
R8570 gnd.n7069 gnd.n539 19.3944
R8571 gnd.n7069 gnd.n535 19.3944
R8572 gnd.n7075 gnd.n535 19.3944
R8573 gnd.n7075 gnd.n533 19.3944
R8574 gnd.n7079 gnd.n533 19.3944
R8575 gnd.n7079 gnd.n529 19.3944
R8576 gnd.n7085 gnd.n529 19.3944
R8577 gnd.n4177 gnd.n4174 19.3944
R8578 gnd.n4177 gnd.n4173 19.3944
R8579 gnd.n4183 gnd.n4173 19.3944
R8580 gnd.n4183 gnd.n4171 19.3944
R8581 gnd.n4187 gnd.n4171 19.3944
R8582 gnd.n4187 gnd.n4169 19.3944
R8583 gnd.n4193 gnd.n4169 19.3944
R8584 gnd.n4193 gnd.n4167 19.3944
R8585 gnd.n4197 gnd.n4167 19.3944
R8586 gnd.n4197 gnd.n4165 19.3944
R8587 gnd.n4203 gnd.n4165 19.3944
R8588 gnd.n4203 gnd.n4163 19.3944
R8589 gnd.n4207 gnd.n4163 19.3944
R8590 gnd.n4207 gnd.n4161 19.3944
R8591 gnd.n4213 gnd.n4161 19.3944
R8592 gnd.n4213 gnd.n4159 19.3944
R8593 gnd.n4220 gnd.n4159 19.3944
R8594 gnd.n4226 gnd.n4157 19.3944
R8595 gnd.n4226 gnd.n4155 19.3944
R8596 gnd.n4230 gnd.n4155 19.3944
R8597 gnd.n4230 gnd.n4153 19.3944
R8598 gnd.n4236 gnd.n4153 19.3944
R8599 gnd.n4236 gnd.n4151 19.3944
R8600 gnd.n4241 gnd.n4151 19.3944
R8601 gnd.n4249 gnd.n1841 19.3944
R8602 gnd.n4249 gnd.n1839 19.3944
R8603 gnd.n4253 gnd.n1839 19.3944
R8604 gnd.n4253 gnd.n1837 19.3944
R8605 gnd.n4259 gnd.n1837 19.3944
R8606 gnd.n4259 gnd.n1835 19.3944
R8607 gnd.n4263 gnd.n1835 19.3944
R8608 gnd.n4263 gnd.n1833 19.3944
R8609 gnd.n4275 gnd.n1831 19.3944
R8610 gnd.n4275 gnd.n1829 19.3944
R8611 gnd.n4281 gnd.n1829 19.3944
R8612 gnd.n4281 gnd.n1827 19.3944
R8613 gnd.n4285 gnd.n1827 19.3944
R8614 gnd.n4285 gnd.n1825 19.3944
R8615 gnd.n4291 gnd.n1825 19.3944
R8616 gnd.n4291 gnd.n1823 19.3944
R8617 gnd.n4295 gnd.n1823 19.3944
R8618 gnd.n4295 gnd.n1821 19.3944
R8619 gnd.n4301 gnd.n1821 19.3944
R8620 gnd.n4301 gnd.n1819 19.3944
R8621 gnd.n4305 gnd.n1819 19.3944
R8622 gnd.n4305 gnd.n1817 19.3944
R8623 gnd.n4311 gnd.n1817 19.3944
R8624 gnd.n4311 gnd.n1815 19.3944
R8625 gnd.n4316 gnd.n1815 19.3944
R8626 gnd.n4316 gnd.n1813 19.3944
R8627 gnd.n4329 gnd.n1806 19.3944
R8628 gnd.n4330 gnd.n4329 19.3944
R8629 gnd.n4331 gnd.n4330 19.3944
R8630 gnd.n4331 gnd.n1801 19.3944
R8631 gnd.n4343 gnd.n1801 19.3944
R8632 gnd.n4344 gnd.n4343 19.3944
R8633 gnd.n4345 gnd.n4344 19.3944
R8634 gnd.n4345 gnd.n1764 19.3944
R8635 gnd.n4357 gnd.n1764 19.3944
R8636 gnd.n4358 gnd.n4357 19.3944
R8637 gnd.n4359 gnd.n4358 19.3944
R8638 gnd.n4360 gnd.n4359 19.3944
R8639 gnd.n4364 gnd.n4360 19.3944
R8640 gnd.n4365 gnd.n4364 19.3944
R8641 gnd.n4369 gnd.n4365 19.3944
R8642 gnd.n4370 gnd.n4369 19.3944
R8643 gnd.n4372 gnd.n4370 19.3944
R8644 gnd.n4372 gnd.n1742 19.3944
R8645 gnd.n4417 gnd.n1742 19.3944
R8646 gnd.n4418 gnd.n4417 19.3944
R8647 gnd.n4443 gnd.n4418 19.3944
R8648 gnd.n4443 gnd.n4442 19.3944
R8649 gnd.n4442 gnd.n4441 19.3944
R8650 gnd.n4441 gnd.n4440 19.3944
R8651 gnd.n4440 gnd.n4439 19.3944
R8652 gnd.n4439 gnd.n4438 19.3944
R8653 gnd.n4438 gnd.n4422 19.3944
R8654 gnd.n4427 gnd.n4422 19.3944
R8655 gnd.n4427 gnd.n378 19.3944
R8656 gnd.n7330 gnd.n378 19.3944
R8657 gnd.n7331 gnd.n7330 19.3944
R8658 gnd.n7332 gnd.n7331 19.3944
R8659 gnd.n7332 gnd.n372 19.3944
R8660 gnd.n7344 gnd.n372 19.3944
R8661 gnd.n7345 gnd.n7344 19.3944
R8662 gnd.n7346 gnd.n7345 19.3944
R8663 gnd.n7346 gnd.n366 19.3944
R8664 gnd.n7358 gnd.n366 19.3944
R8665 gnd.n7359 gnd.n7358 19.3944
R8666 gnd.n7360 gnd.n7359 19.3944
R8667 gnd.n7360 gnd.n360 19.3944
R8668 gnd.n7373 gnd.n360 19.3944
R8669 gnd.n7374 gnd.n7373 19.3944
R8670 gnd.n7390 gnd.n7374 19.3944
R8671 gnd.n7390 gnd.n7389 19.3944
R8672 gnd.n7389 gnd.n7388 19.3944
R8673 gnd.n7388 gnd.n7386 19.3944
R8674 gnd.n7386 gnd.n7385 19.3944
R8675 gnd.n7385 gnd.n7383 19.3944
R8676 gnd.n7383 gnd.n7382 19.3944
R8677 gnd.n7382 gnd.n7380 19.3944
R8678 gnd.n7380 gnd.n7379 19.3944
R8679 gnd.n7379 gnd.n7377 19.3944
R8680 gnd.n4326 gnd.n1617 19.3944
R8681 gnd.n4538 gnd.n1617 19.3944
R8682 gnd.n4538 gnd.n4537 19.3944
R8683 gnd.n4537 gnd.n4536 19.3944
R8684 gnd.n4536 gnd.n1621 19.3944
R8685 gnd.n4526 gnd.n1621 19.3944
R8686 gnd.n4526 gnd.n4525 19.3944
R8687 gnd.n4525 gnd.n4524 19.3944
R8688 gnd.n4524 gnd.n1641 19.3944
R8689 gnd.n4514 gnd.n1641 19.3944
R8690 gnd.n4514 gnd.n4513 19.3944
R8691 gnd.n4513 gnd.n4512 19.3944
R8692 gnd.n4512 gnd.n1662 19.3944
R8693 gnd.n4502 gnd.n1662 19.3944
R8694 gnd.n4502 gnd.n4501 19.3944
R8695 gnd.n4501 gnd.n4500 19.3944
R8696 gnd.n4500 gnd.n1681 19.3944
R8697 gnd.n4490 gnd.n1681 19.3944
R8698 gnd.n4490 gnd.n4489 19.3944
R8699 gnd.n4489 gnd.n4488 19.3944
R8700 gnd.n4488 gnd.n1702 19.3944
R8701 gnd.n4478 gnd.n1702 19.3944
R8702 gnd.n4478 gnd.n4477 19.3944
R8703 gnd.n4477 gnd.n4476 19.3944
R8704 gnd.n4476 gnd.n1719 19.3944
R8705 gnd.n4425 gnd.n1719 19.3944
R8706 gnd.n4433 gnd.n4425 19.3944
R8707 gnd.n4433 gnd.n4432 19.3944
R8708 gnd.n4432 gnd.n4431 19.3944
R8709 gnd.n4431 gnd.n108 19.3944
R8710 gnd.n7621 gnd.n108 19.3944
R8711 gnd.n7621 gnd.n7620 19.3944
R8712 gnd.n7620 gnd.n7619 19.3944
R8713 gnd.n7619 gnd.n112 19.3944
R8714 gnd.n7609 gnd.n112 19.3944
R8715 gnd.n7609 gnd.n7608 19.3944
R8716 gnd.n7608 gnd.n7607 19.3944
R8717 gnd.n7607 gnd.n130 19.3944
R8718 gnd.n7597 gnd.n130 19.3944
R8719 gnd.n7597 gnd.n7596 19.3944
R8720 gnd.n7596 gnd.n7595 19.3944
R8721 gnd.n7595 gnd.n151 19.3944
R8722 gnd.n7585 gnd.n151 19.3944
R8723 gnd.n7585 gnd.n7584 19.3944
R8724 gnd.n7584 gnd.n7583 19.3944
R8725 gnd.n7583 gnd.n170 19.3944
R8726 gnd.n7573 gnd.n170 19.3944
R8727 gnd.n7573 gnd.n7572 19.3944
R8728 gnd.n7572 gnd.n7571 19.3944
R8729 gnd.n7571 gnd.n190 19.3944
R8730 gnd.n7561 gnd.n190 19.3944
R8731 gnd.n7561 gnd.n7560 19.3944
R8732 gnd.n7560 gnd.n7559 19.3944
R8733 gnd.n7481 gnd.n279 19.3944
R8734 gnd.n7481 gnd.n283 19.3944
R8735 gnd.n286 gnd.n283 19.3944
R8736 gnd.n7474 gnd.n286 19.3944
R8737 gnd.n7474 gnd.n7473 19.3944
R8738 gnd.n7473 gnd.n7472 19.3944
R8739 gnd.n7472 gnd.n292 19.3944
R8740 gnd.n7467 gnd.n292 19.3944
R8741 gnd.n7467 gnd.n7466 19.3944
R8742 gnd.n7466 gnd.n7465 19.3944
R8743 gnd.n7465 gnd.n299 19.3944
R8744 gnd.n7460 gnd.n299 19.3944
R8745 gnd.n7460 gnd.n7459 19.3944
R8746 gnd.n7459 gnd.n7458 19.3944
R8747 gnd.n7458 gnd.n306 19.3944
R8748 gnd.n7453 gnd.n306 19.3944
R8749 gnd.n7453 gnd.n7452 19.3944
R8750 gnd.n7452 gnd.n7451 19.3944
R8751 gnd.n7519 gnd.n246 19.3944
R8752 gnd.n7514 gnd.n246 19.3944
R8753 gnd.n7514 gnd.n7513 19.3944
R8754 gnd.n7513 gnd.n7512 19.3944
R8755 gnd.n7512 gnd.n253 19.3944
R8756 gnd.n7507 gnd.n253 19.3944
R8757 gnd.n7507 gnd.n7506 19.3944
R8758 gnd.n7506 gnd.n7505 19.3944
R8759 gnd.n7505 gnd.n260 19.3944
R8760 gnd.n7500 gnd.n260 19.3944
R8761 gnd.n7500 gnd.n7499 19.3944
R8762 gnd.n7499 gnd.n7498 19.3944
R8763 gnd.n7498 gnd.n267 19.3944
R8764 gnd.n7493 gnd.n267 19.3944
R8765 gnd.n7493 gnd.n7492 19.3944
R8766 gnd.n7492 gnd.n7491 19.3944
R8767 gnd.n7491 gnd.n274 19.3944
R8768 gnd.n7486 gnd.n274 19.3944
R8769 gnd.n7552 gnd.n7551 19.3944
R8770 gnd.n7551 gnd.n7550 19.3944
R8771 gnd.n7550 gnd.n218 19.3944
R8772 gnd.n7545 gnd.n218 19.3944
R8773 gnd.n7545 gnd.n7544 19.3944
R8774 gnd.n7544 gnd.n7543 19.3944
R8775 gnd.n7543 gnd.n225 19.3944
R8776 gnd.n7538 gnd.n225 19.3944
R8777 gnd.n7538 gnd.n7537 19.3944
R8778 gnd.n7537 gnd.n7536 19.3944
R8779 gnd.n7536 gnd.n232 19.3944
R8780 gnd.n7531 gnd.n232 19.3944
R8781 gnd.n7531 gnd.n7530 19.3944
R8782 gnd.n7530 gnd.n7529 19.3944
R8783 gnd.n7529 gnd.n239 19.3944
R8784 gnd.n7524 gnd.n239 19.3944
R8785 gnd.n7524 gnd.n7523 19.3944
R8786 gnd.n7442 gnd.n7441 19.3944
R8787 gnd.n7441 gnd.n7440 19.3944
R8788 gnd.n7440 gnd.n321 19.3944
R8789 gnd.n7435 gnd.n321 19.3944
R8790 gnd.n7435 gnd.n7434 19.3944
R8791 gnd.n7434 gnd.n7433 19.3944
R8792 gnd.n7433 gnd.n328 19.3944
R8793 gnd.n7428 gnd.n328 19.3944
R8794 gnd.n7428 gnd.n7427 19.3944
R8795 gnd.n7427 gnd.n7426 19.3944
R8796 gnd.n7426 gnd.n335 19.3944
R8797 gnd.n7421 gnd.n335 19.3944
R8798 gnd.n7421 gnd.n7420 19.3944
R8799 gnd.n7420 gnd.n7419 19.3944
R8800 gnd.n7419 gnd.n342 19.3944
R8801 gnd.n7414 gnd.n342 19.3944
R8802 gnd.n3757 gnd.n3756 19.3944
R8803 gnd.n3756 gnd.n1805 19.3944
R8804 gnd.n4335 gnd.n1805 19.3944
R8805 gnd.n4335 gnd.n1803 19.3944
R8806 gnd.n4339 gnd.n1803 19.3944
R8807 gnd.n4339 gnd.n1768 19.3944
R8808 gnd.n4349 gnd.n1768 19.3944
R8809 gnd.n4349 gnd.n1766 19.3944
R8810 gnd.n4353 gnd.n1766 19.3944
R8811 gnd.n4353 gnd.n1756 19.3944
R8812 gnd.n4389 gnd.n1756 19.3944
R8813 gnd.n4389 gnd.n1757 19.3944
R8814 gnd.n4385 gnd.n1757 19.3944
R8815 gnd.n4385 gnd.n4384 19.3944
R8816 gnd.n4384 gnd.n4383 19.3944
R8817 gnd.n4383 gnd.n1762 19.3944
R8818 gnd.n4379 gnd.n1762 19.3944
R8819 gnd.n4379 gnd.n4378 19.3944
R8820 gnd.n4378 gnd.n4377 19.3944
R8821 gnd.n4377 gnd.n1741 19.3944
R8822 gnd.n4447 gnd.n1741 19.3944
R8823 gnd.n4447 gnd.n1738 19.3944
R8824 gnd.n4454 gnd.n1738 19.3944
R8825 gnd.n4454 gnd.n1739 19.3944
R8826 gnd.n4450 gnd.n1739 19.3944
R8827 gnd.n4450 gnd.n81 19.3944
R8828 gnd.n7634 gnd.n81 19.3944
R8829 gnd.n7634 gnd.n7633 19.3944
R8830 gnd.n7633 gnd.n83 19.3944
R8831 gnd.n7326 gnd.n83 19.3944
R8832 gnd.n7326 gnd.n377 19.3944
R8833 gnd.n7336 gnd.n377 19.3944
R8834 gnd.n7336 gnd.n375 19.3944
R8835 gnd.n7340 gnd.n375 19.3944
R8836 gnd.n7340 gnd.n370 19.3944
R8837 gnd.n7350 gnd.n370 19.3944
R8838 gnd.n7350 gnd.n368 19.3944
R8839 gnd.n7354 gnd.n368 19.3944
R8840 gnd.n7354 gnd.n365 19.3944
R8841 gnd.n7364 gnd.n365 19.3944
R8842 gnd.n7364 gnd.n363 19.3944
R8843 gnd.n7369 gnd.n363 19.3944
R8844 gnd.n7369 gnd.n359 19.3944
R8845 gnd.n7394 gnd.n359 19.3944
R8846 gnd.n7395 gnd.n7394 19.3944
R8847 gnd.n7395 gnd.n357 19.3944
R8848 gnd.n7399 gnd.n357 19.3944
R8849 gnd.n7401 gnd.n7399 19.3944
R8850 gnd.n7402 gnd.n7401 19.3944
R8851 gnd.n7402 gnd.n354 19.3944
R8852 gnd.n7406 gnd.n354 19.3944
R8853 gnd.n7408 gnd.n7406 19.3944
R8854 gnd.n7409 gnd.n7408 19.3944
R8855 gnd.n4544 gnd.n4543 19.3944
R8856 gnd.n4543 gnd.n4542 19.3944
R8857 gnd.n4542 gnd.n1609 19.3944
R8858 gnd.n4532 gnd.n1609 19.3944
R8859 gnd.n4532 gnd.n4531 19.3944
R8860 gnd.n4531 gnd.n4530 19.3944
R8861 gnd.n4530 gnd.n1632 19.3944
R8862 gnd.n4520 gnd.n1632 19.3944
R8863 gnd.n4520 gnd.n4519 19.3944
R8864 gnd.n4519 gnd.n4518 19.3944
R8865 gnd.n4518 gnd.n1652 19.3944
R8866 gnd.n4508 gnd.n1652 19.3944
R8867 gnd.n4508 gnd.n4507 19.3944
R8868 gnd.n4507 gnd.n4506 19.3944
R8869 gnd.n4506 gnd.n1672 19.3944
R8870 gnd.n4496 gnd.n1672 19.3944
R8871 gnd.n4496 gnd.n4495 19.3944
R8872 gnd.n4495 gnd.n4494 19.3944
R8873 gnd.n4494 gnd.n1692 19.3944
R8874 gnd.n4484 gnd.n1692 19.3944
R8875 gnd.n4484 gnd.n4483 19.3944
R8876 gnd.n4483 gnd.n4482 19.3944
R8877 gnd.n1710 gnd.n97 19.3944
R8878 gnd.n1728 gnd.n97 19.3944
R8879 gnd.n1726 gnd.n1725 19.3944
R8880 gnd.n7629 gnd.n7628 19.3944
R8881 gnd.n7625 gnd.n92 19.3944
R8882 gnd.n7625 gnd.n99 19.3944
R8883 gnd.n7615 gnd.n99 19.3944
R8884 gnd.n7615 gnd.n7614 19.3944
R8885 gnd.n7614 gnd.n7613 19.3944
R8886 gnd.n7613 gnd.n121 19.3944
R8887 gnd.n7603 gnd.n121 19.3944
R8888 gnd.n7603 gnd.n7602 19.3944
R8889 gnd.n7602 gnd.n7601 19.3944
R8890 gnd.n7601 gnd.n141 19.3944
R8891 gnd.n7591 gnd.n141 19.3944
R8892 gnd.n7591 gnd.n7590 19.3944
R8893 gnd.n7590 gnd.n7589 19.3944
R8894 gnd.n7589 gnd.n161 19.3944
R8895 gnd.n7579 gnd.n161 19.3944
R8896 gnd.n7579 gnd.n7578 19.3944
R8897 gnd.n7578 gnd.n7577 19.3944
R8898 gnd.n7577 gnd.n181 19.3944
R8899 gnd.n7567 gnd.n181 19.3944
R8900 gnd.n7567 gnd.n7566 19.3944
R8901 gnd.n7566 gnd.n7565 19.3944
R8902 gnd.n7565 gnd.n200 19.3944
R8903 gnd.n7555 gnd.n200 19.3944
R8904 gnd.n2790 gnd.n2784 19.3944
R8905 gnd.n2794 gnd.n2784 19.3944
R8906 gnd.n2794 gnd.n2782 19.3944
R8907 gnd.n2816 gnd.n2782 19.3944
R8908 gnd.n2816 gnd.n2815 19.3944
R8909 gnd.n2815 gnd.n2814 19.3944
R8910 gnd.n2814 gnd.n2800 19.3944
R8911 gnd.n2810 gnd.n2800 19.3944
R8912 gnd.n2810 gnd.n2809 19.3944
R8913 gnd.n2809 gnd.n2808 19.3944
R8914 gnd.n2808 gnd.n2638 19.3944
R8915 gnd.n2863 gnd.n2638 19.3944
R8916 gnd.n2866 gnd.n2865 19.3944
R8917 gnd.n2870 gnd.n2869 19.3944
R8918 gnd.n2875 gnd.n2874 19.3944
R8919 gnd.n2872 gnd.n2596 19.3944
R8920 gnd.n2944 gnd.n2593 19.3944
R8921 gnd.n2944 gnd.n2592 19.3944
R8922 gnd.n2948 gnd.n2592 19.3944
R8923 gnd.n2948 gnd.n2590 19.3944
R8924 gnd.n2952 gnd.n2590 19.3944
R8925 gnd.n2952 gnd.n2588 19.3944
R8926 gnd.n2976 gnd.n2588 19.3944
R8927 gnd.n2976 gnd.n2975 19.3944
R8928 gnd.n2975 gnd.n2974 19.3944
R8929 gnd.n2974 gnd.n2958 19.3944
R8930 gnd.n2970 gnd.n2958 19.3944
R8931 gnd.n2970 gnd.n2969 19.3944
R8932 gnd.n2969 gnd.n2968 19.3944
R8933 gnd.n2968 gnd.n2966 19.3944
R8934 gnd.n2966 gnd.n2566 19.3944
R8935 gnd.n2566 gnd.n2564 19.3944
R8936 gnd.n3041 gnd.n2564 19.3944
R8937 gnd.n3041 gnd.n2562 19.3944
R8938 gnd.n3045 gnd.n2562 19.3944
R8939 gnd.n3045 gnd.n2560 19.3944
R8940 gnd.n3049 gnd.n2560 19.3944
R8941 gnd.n3049 gnd.n2558 19.3944
R8942 gnd.n3053 gnd.n2558 19.3944
R8943 gnd.n3053 gnd.n2556 19.3944
R8944 gnd.n3060 gnd.n2556 19.3944
R8945 gnd.n3060 gnd.n2554 19.3944
R8946 gnd.n3066 gnd.n2554 19.3944
R8947 gnd.n3066 gnd.n3065 19.3944
R8948 gnd.n3065 gnd.n2325 19.3944
R8949 gnd.n3156 gnd.n2325 19.3944
R8950 gnd.n3156 gnd.n2323 19.3944
R8951 gnd.n3162 gnd.n2323 19.3944
R8952 gnd.n3162 gnd.n3161 19.3944
R8953 gnd.n3161 gnd.n2300 19.3944
R8954 gnd.n3186 gnd.n2300 19.3944
R8955 gnd.n3186 gnd.n2298 19.3944
R8956 gnd.n3192 gnd.n2298 19.3944
R8957 gnd.n3192 gnd.n3191 19.3944
R8958 gnd.n3191 gnd.n2275 19.3944
R8959 gnd.n3216 gnd.n2275 19.3944
R8960 gnd.n3216 gnd.n2273 19.3944
R8961 gnd.n3232 gnd.n2273 19.3944
R8962 gnd.n3232 gnd.n3231 19.3944
R8963 gnd.n3231 gnd.n3230 19.3944
R8964 gnd.n3230 gnd.n3222 19.3944
R8965 gnd.n3225 gnd.n3222 19.3944
R8966 gnd.n3225 gnd.n2181 19.3944
R8967 gnd.n3291 gnd.n2181 19.3944
R8968 gnd.n3291 gnd.n2179 19.3944
R8969 gnd.n3297 gnd.n2179 19.3944
R8970 gnd.n3297 gnd.n3296 19.3944
R8971 gnd.n3296 gnd.n2155 19.3944
R8972 gnd.n3353 gnd.n2155 19.3944
R8973 gnd.n3353 gnd.n2153 19.3944
R8974 gnd.n3357 gnd.n2153 19.3944
R8975 gnd.n3357 gnd.n2137 19.3944
R8976 gnd.n3380 gnd.n2137 19.3944
R8977 gnd.n3380 gnd.n2135 19.3944
R8978 gnd.n3386 gnd.n2135 19.3944
R8979 gnd.n3386 gnd.n3385 19.3944
R8980 gnd.n3385 gnd.n2104 19.3944
R8981 gnd.n3431 gnd.n2104 19.3944
R8982 gnd.n3431 gnd.n2102 19.3944
R8983 gnd.n3435 gnd.n2102 19.3944
R8984 gnd.n3435 gnd.n2081 19.3944
R8985 gnd.n3471 gnd.n2081 19.3944
R8986 gnd.n3471 gnd.n2079 19.3944
R8987 gnd.n3475 gnd.n2079 19.3944
R8988 gnd.n3475 gnd.n2059 19.3944
R8989 gnd.n3527 gnd.n2059 19.3944
R8990 gnd.n3527 gnd.n2057 19.3944
R8991 gnd.n3531 gnd.n2057 19.3944
R8992 gnd.n3531 gnd.n2040 19.3944
R8993 gnd.n3552 gnd.n2040 19.3944
R8994 gnd.n3552 gnd.n2038 19.3944
R8995 gnd.n3556 gnd.n2038 19.3944
R8996 gnd.n3556 gnd.n2020 19.3944
R8997 gnd.n3612 gnd.n2020 19.3944
R8998 gnd.n3612 gnd.n2018 19.3944
R8999 gnd.n3616 gnd.n2018 19.3944
R9000 gnd.n3616 gnd.n1998 19.3944
R9001 gnd.n3641 gnd.n1998 19.3944
R9002 gnd.n3641 gnd.n1996 19.3944
R9003 gnd.n3647 gnd.n1996 19.3944
R9004 gnd.n3647 gnd.n3646 19.3944
R9005 gnd.n3646 gnd.n1970 19.3944
R9006 gnd.n3686 gnd.n1970 19.3944
R9007 gnd.n3686 gnd.n1968 19.3944
R9008 gnd.n3696 gnd.n1968 19.3944
R9009 gnd.n3696 gnd.n3695 19.3944
R9010 gnd.n3695 gnd.n3694 19.3944
R9011 gnd.n3694 gnd.n1894 19.3944
R9012 gnd.n3983 gnd.n1894 19.3944
R9013 gnd.n3983 gnd.n3982 19.3944
R9014 gnd.n3982 gnd.n3981 19.3944
R9015 gnd.n3981 gnd.n1898 19.3944
R9016 gnd.n3972 gnd.n1898 19.3944
R9017 gnd.n3972 gnd.n3971 19.3944
R9018 gnd.n3971 gnd.n3970 19.3944
R9019 gnd.n3970 gnd.n1908 19.3944
R9020 gnd.n3961 gnd.n1908 19.3944
R9021 gnd.n3961 gnd.n3960 19.3944
R9022 gnd.n3960 gnd.n3959 19.3944
R9023 gnd.n3959 gnd.n1920 19.3944
R9024 gnd.n3950 gnd.n1920 19.3944
R9025 gnd.n3950 gnd.n3949 19.3944
R9026 gnd.n3949 gnd.n3948 19.3944
R9027 gnd.n3948 gnd.n1932 19.3944
R9028 gnd.n3939 gnd.n1932 19.3944
R9029 gnd.n3939 gnd.n1584 19.3944
R9030 gnd.n4559 gnd.n1584 19.3944
R9031 gnd.n4559 gnd.n4558 19.3944
R9032 gnd.n4558 gnd.n4557 19.3944
R9033 gnd.n4557 gnd.n1588 19.3944
R9034 gnd.n4551 gnd.n1588 19.3944
R9035 gnd.n4551 gnd.n4550 19.3944
R9036 gnd.n4550 gnd.n4549 19.3944
R9037 gnd.n4549 gnd.n1597 19.3944
R9038 gnd.n1775 gnd.n1597 19.3944
R9039 gnd.n1779 gnd.n1775 19.3944
R9040 gnd.n1779 gnd.n1773 19.3944
R9041 gnd.n1783 gnd.n1773 19.3944
R9042 gnd.n1783 gnd.n1771 19.3944
R9043 gnd.n1798 gnd.n1771 19.3944
R9044 gnd.n1798 gnd.n1797 19.3944
R9045 gnd.n1797 gnd.n1796 19.3944
R9046 gnd.n1796 gnd.n1793 19.3944
R9047 gnd.n1793 gnd.n1792 19.3944
R9048 gnd.n1792 gnd.n1754 19.3944
R9049 gnd.n1754 gnd.n1752 19.3944
R9050 gnd.n4396 gnd.n1752 19.3944
R9051 gnd.n4396 gnd.n1750 19.3944
R9052 gnd.n4400 gnd.n1750 19.3944
R9053 gnd.n4400 gnd.n1748 19.3944
R9054 gnd.n4404 gnd.n1748 19.3944
R9055 gnd.n4404 gnd.n1746 19.3944
R9056 gnd.n4412 gnd.n1746 19.3944
R9057 gnd.n4412 gnd.n4411 19.3944
R9058 gnd.n4411 gnd.n4410 19.3944
R9059 gnd.n4460 gnd.n1735 19.3944
R9060 gnd.n4468 gnd.n4462 19.3944
R9061 gnd.n4466 gnd.n4465 19.3944
R9062 gnd.n7321 gnd.n384 19.3944
R9063 gnd.n7319 gnd.n7318 19.3944
R9064 gnd.n7318 gnd.n386 19.3944
R9065 gnd.n7314 gnd.n386 19.3944
R9066 gnd.n7314 gnd.n7313 19.3944
R9067 gnd.n7313 gnd.n7312 19.3944
R9068 gnd.n7312 gnd.n392 19.3944
R9069 gnd.n7308 gnd.n392 19.3944
R9070 gnd.n7308 gnd.n7307 19.3944
R9071 gnd.n7307 gnd.n7306 19.3944
R9072 gnd.n7306 gnd.n398 19.3944
R9073 gnd.n7302 gnd.n398 19.3944
R9074 gnd.n7302 gnd.n7301 19.3944
R9075 gnd.n5043 gnd.n5042 19.3944
R9076 gnd.n5042 gnd.n5041 19.3944
R9077 gnd.n5041 gnd.n5040 19.3944
R9078 gnd.n5040 gnd.n5038 19.3944
R9079 gnd.n5038 gnd.n5035 19.3944
R9080 gnd.n5035 gnd.n5034 19.3944
R9081 gnd.n5034 gnd.n5031 19.3944
R9082 gnd.n5031 gnd.n5030 19.3944
R9083 gnd.n5030 gnd.n5027 19.3944
R9084 gnd.n5027 gnd.n5026 19.3944
R9085 gnd.n5026 gnd.n5023 19.3944
R9086 gnd.n5023 gnd.n5022 19.3944
R9087 gnd.n5022 gnd.n5019 19.3944
R9088 gnd.n5019 gnd.n5018 19.3944
R9089 gnd.n5018 gnd.n5015 19.3944
R9090 gnd.n5015 gnd.n5014 19.3944
R9091 gnd.n5014 gnd.n5011 19.3944
R9092 gnd.n5009 gnd.n5006 19.3944
R9093 gnd.n5006 gnd.n5005 19.3944
R9094 gnd.n5005 gnd.n5002 19.3944
R9095 gnd.n5002 gnd.n5001 19.3944
R9096 gnd.n5001 gnd.n4998 19.3944
R9097 gnd.n4998 gnd.n4997 19.3944
R9098 gnd.n4997 gnd.n4994 19.3944
R9099 gnd.n4994 gnd.n4993 19.3944
R9100 gnd.n4993 gnd.n4990 19.3944
R9101 gnd.n4990 gnd.n4989 19.3944
R9102 gnd.n4989 gnd.n4986 19.3944
R9103 gnd.n4986 gnd.n4985 19.3944
R9104 gnd.n4985 gnd.n4982 19.3944
R9105 gnd.n4982 gnd.n4981 19.3944
R9106 gnd.n4981 gnd.n4978 19.3944
R9107 gnd.n4978 gnd.n4977 19.3944
R9108 gnd.n4977 gnd.n4974 19.3944
R9109 gnd.n4974 gnd.n4973 19.3944
R9110 gnd.n4969 gnd.n4966 19.3944
R9111 gnd.n4966 gnd.n4965 19.3944
R9112 gnd.n4965 gnd.n4962 19.3944
R9113 gnd.n4962 gnd.n4961 19.3944
R9114 gnd.n4961 gnd.n4958 19.3944
R9115 gnd.n4958 gnd.n4957 19.3944
R9116 gnd.n4957 gnd.n4954 19.3944
R9117 gnd.n4954 gnd.n4953 19.3944
R9118 gnd.n4953 gnd.n4950 19.3944
R9119 gnd.n4950 gnd.n4949 19.3944
R9120 gnd.n4949 gnd.n4946 19.3944
R9121 gnd.n4946 gnd.n4945 19.3944
R9122 gnd.n4945 gnd.n4942 19.3944
R9123 gnd.n4942 gnd.n4941 19.3944
R9124 gnd.n4941 gnd.n4938 19.3944
R9125 gnd.n4938 gnd.n4937 19.3944
R9126 gnd.n4937 gnd.n4934 19.3944
R9127 gnd.n4934 gnd.n4933 19.3944
R9128 gnd.n2702 gnd.n2701 19.3944
R9129 gnd.n2705 gnd.n2702 19.3944
R9130 gnd.n2705 gnd.n2697 19.3944
R9131 gnd.n2711 gnd.n2697 19.3944
R9132 gnd.n2712 gnd.n2711 19.3944
R9133 gnd.n2715 gnd.n2712 19.3944
R9134 gnd.n2715 gnd.n2695 19.3944
R9135 gnd.n2721 gnd.n2695 19.3944
R9136 gnd.n2722 gnd.n2721 19.3944
R9137 gnd.n2725 gnd.n2722 19.3944
R9138 gnd.n2725 gnd.n2693 19.3944
R9139 gnd.n2731 gnd.n2693 19.3944
R9140 gnd.n2732 gnd.n2731 19.3944
R9141 gnd.n2735 gnd.n2732 19.3944
R9142 gnd.n2735 gnd.n2689 19.3944
R9143 gnd.n2739 gnd.n2689 19.3944
R9144 gnd.n2744 gnd.n2684 19.3944
R9145 gnd.n2749 gnd.n2684 19.3944
R9146 gnd.n2750 gnd.n2749 19.3944
R9147 gnd.n2752 gnd.n2750 19.3944
R9148 gnd.n2752 gnd.n2682 19.3944
R9149 gnd.n2757 gnd.n2682 19.3944
R9150 gnd.n2758 gnd.n2757 19.3944
R9151 gnd.n2760 gnd.n2758 19.3944
R9152 gnd.n2760 gnd.n2680 19.3944
R9153 gnd.n2764 gnd.n2680 19.3944
R9154 gnd.n2764 gnd.n2665 19.3944
R9155 gnd.n2774 gnd.n2665 19.3944
R9156 gnd.n2774 gnd.n2663 19.3944
R9157 gnd.n2778 gnd.n2663 19.3944
R9158 gnd.n2778 gnd.n2660 19.3944
R9159 gnd.n2827 gnd.n2660 19.3944
R9160 gnd.n2827 gnd.n2658 19.3944
R9161 gnd.n2832 gnd.n2658 19.3944
R9162 gnd.n2832 gnd.n2654 19.3944
R9163 gnd.n2843 gnd.n2654 19.3944
R9164 gnd.n2844 gnd.n2843 19.3944
R9165 gnd.n2846 gnd.n2844 19.3944
R9166 gnd.n2846 gnd.n2652 19.3944
R9167 gnd.n2850 gnd.n2652 19.3944
R9168 gnd.n2850 gnd.n2618 19.3944
R9169 gnd.n2891 gnd.n2618 19.3944
R9170 gnd.n2891 gnd.n2616 19.3944
R9171 gnd.n2896 gnd.n2616 19.3944
R9172 gnd.n2896 gnd.n2600 19.3944
R9173 gnd.n2937 gnd.n2600 19.3944
R9174 gnd.n2937 gnd.n2601 19.3944
R9175 gnd.n2933 gnd.n2601 19.3944
R9176 gnd.n2933 gnd.n2932 19.3944
R9177 gnd.n2932 gnd.n2931 19.3944
R9178 gnd.n2931 gnd.n2606 19.3944
R9179 gnd.n2927 gnd.n2606 19.3944
R9180 gnd.n2927 gnd.n2584 19.3944
R9181 gnd.n2981 gnd.n2584 19.3944
R9182 gnd.n2981 gnd.n2582 19.3944
R9183 gnd.n2985 gnd.n2582 19.3944
R9184 gnd.n2985 gnd.n2579 19.3944
R9185 gnd.n2996 gnd.n2579 19.3944
R9186 gnd.n2996 gnd.n2577 19.3944
R9187 gnd.n3000 gnd.n2577 19.3944
R9188 gnd.n3000 gnd.n2568 19.3944
R9189 gnd.n3034 gnd.n2568 19.3944
R9190 gnd.n3034 gnd.n2569 19.3944
R9191 gnd.n3030 gnd.n2569 19.3944
R9192 gnd.n3030 gnd.n3029 19.3944
R9193 gnd.n3029 gnd.n3028 19.3944
R9194 gnd.n3028 gnd.n2574 19.3944
R9195 gnd.n3024 gnd.n2574 19.3944
R9196 gnd.n3024 gnd.n3023 19.3944
R9197 gnd.n4925 gnd.n1139 19.3944
R9198 gnd.n2667 gnd.n1139 19.3944
R9199 gnd.n2668 gnd.n2667 19.3944
R9200 gnd.n2670 gnd.n2668 19.3944
R9201 gnd.n2671 gnd.n2670 19.3944
R9202 gnd.n2674 gnd.n2671 19.3944
R9203 gnd.n2675 gnd.n2674 19.3944
R9204 gnd.n2677 gnd.n2675 19.3944
R9205 gnd.n2678 gnd.n2677 19.3944
R9206 gnd.n2768 gnd.n2678 19.3944
R9207 gnd.n2769 gnd.n2768 19.3944
R9208 gnd.n2770 gnd.n2769 19.3944
R9209 gnd.n2770 gnd.n2661 19.3944
R9210 gnd.n2821 gnd.n2661 19.3944
R9211 gnd.n2822 gnd.n2821 19.3944
R9212 gnd.n2823 gnd.n2822 19.3944
R9213 gnd.n2823 gnd.n2656 19.3944
R9214 gnd.n2836 gnd.n2656 19.3944
R9215 gnd.n2837 gnd.n2836 19.3944
R9216 gnd.n2839 gnd.n2837 19.3944
R9217 gnd.n2839 gnd.n2838 19.3944
R9218 gnd.n2838 gnd.n2647 19.3944
R9219 gnd.n2855 gnd.n2647 19.3944
R9220 gnd.n2855 gnd.n2854 19.3944
R9221 gnd.n2854 gnd.n2651 19.3944
R9222 gnd.n2651 gnd.n2650 19.3944
R9223 gnd.n2650 gnd.n2649 19.3944
R9224 gnd.n2649 gnd.n2648 19.3944
R9225 gnd.n2648 gnd.n2607 19.3944
R9226 gnd.n2908 gnd.n2607 19.3944
R9227 gnd.n2909 gnd.n2908 19.3944
R9228 gnd.n2912 gnd.n2909 19.3944
R9229 gnd.n2913 gnd.n2912 19.3944
R9230 gnd.n2918 gnd.n2913 19.3944
R9231 gnd.n2919 gnd.n2918 19.3944
R9232 gnd.n2923 gnd.n2919 19.3944
R9233 gnd.n2923 gnd.n2922 19.3944
R9234 gnd.n2922 gnd.n2921 19.3944
R9235 gnd.n2921 gnd.n2581 19.3944
R9236 gnd.n2989 gnd.n2581 19.3944
R9237 gnd.n2990 gnd.n2989 19.3944
R9238 gnd.n2992 gnd.n2990 19.3944
R9239 gnd.n2992 gnd.n2576 19.3944
R9240 gnd.n3004 gnd.n2576 19.3944
R9241 gnd.n3005 gnd.n3004 19.3944
R9242 gnd.n3007 gnd.n3005 19.3944
R9243 gnd.n3008 gnd.n3007 19.3944
R9244 gnd.n3011 gnd.n3008 19.3944
R9245 gnd.n3012 gnd.n3011 19.3944
R9246 gnd.n3016 gnd.n3012 19.3944
R9247 gnd.n3017 gnd.n3016 19.3944
R9248 gnd.n3019 gnd.n3017 19.3944
R9249 gnd.n3019 gnd.n3018 19.3944
R9250 gnd.n1158 gnd.n1137 19.3944
R9251 gnd.n1159 gnd.n1158 19.3944
R9252 gnd.n4914 gnd.n1159 19.3944
R9253 gnd.n4914 gnd.n4913 19.3944
R9254 gnd.n4913 gnd.n4912 19.3944
R9255 gnd.n4912 gnd.n1163 19.3944
R9256 gnd.n4902 gnd.n1163 19.3944
R9257 gnd.n4902 gnd.n4901 19.3944
R9258 gnd.n4901 gnd.n4900 19.3944
R9259 gnd.n4900 gnd.n1182 19.3944
R9260 gnd.n4890 gnd.n1182 19.3944
R9261 gnd.n4890 gnd.n4889 19.3944
R9262 gnd.n4889 gnd.n4888 19.3944
R9263 gnd.n4888 gnd.n1202 19.3944
R9264 gnd.n4878 gnd.n1202 19.3944
R9265 gnd.n4878 gnd.n4877 19.3944
R9266 gnd.n4877 gnd.n4876 19.3944
R9267 gnd.n4876 gnd.n1222 19.3944
R9268 gnd.n4866 gnd.n1222 19.3944
R9269 gnd.n4866 gnd.n4865 19.3944
R9270 gnd.n4865 gnd.n4864 19.3944
R9271 gnd.n4864 gnd.n1243 19.3944
R9272 gnd.n2857 gnd.n1243 19.3944
R9273 gnd.n2857 gnd.n2629 19.3944
R9274 gnd.n2882 gnd.n2629 19.3944
R9275 gnd.n2882 gnd.n2881 19.3944
R9276 gnd.n2881 gnd.n2880 19.3944
R9277 gnd.n2880 gnd.n2609 19.3944
R9278 gnd.n2905 gnd.n2609 19.3944
R9279 gnd.n2905 gnd.n1268 19.3944
R9280 gnd.n4852 gnd.n1268 19.3944
R9281 gnd.n4852 gnd.n4851 19.3944
R9282 gnd.n4851 gnd.n4850 19.3944
R9283 gnd.n4850 gnd.n1272 19.3944
R9284 gnd.n4840 gnd.n1272 19.3944
R9285 gnd.n4840 gnd.n4839 19.3944
R9286 gnd.n4839 gnd.n4838 19.3944
R9287 gnd.n4838 gnd.n1291 19.3944
R9288 gnd.n4828 gnd.n1291 19.3944
R9289 gnd.n4828 gnd.n4827 19.3944
R9290 gnd.n4827 gnd.n4826 19.3944
R9291 gnd.n4826 gnd.n1311 19.3944
R9292 gnd.n4816 gnd.n1311 19.3944
R9293 gnd.n4816 gnd.n4815 19.3944
R9294 gnd.n4815 gnd.n4814 19.3944
R9295 gnd.n4814 gnd.n1331 19.3944
R9296 gnd.n4804 gnd.n1331 19.3944
R9297 gnd.n4804 gnd.n4803 19.3944
R9298 gnd.n4803 gnd.n4802 19.3944
R9299 gnd.n4802 gnd.n1351 19.3944
R9300 gnd.n4792 gnd.n1351 19.3944
R9301 gnd.n4792 gnd.n4791 19.3944
R9302 gnd.n4791 gnd.n4790 19.3944
R9303 gnd.n4783 gnd.n4782 19.3944
R9304 gnd.n4782 gnd.n1380 19.3944
R9305 gnd.n1382 gnd.n1380 19.3944
R9306 gnd.n4775 gnd.n1382 19.3944
R9307 gnd.n4775 gnd.n4774 19.3944
R9308 gnd.n4774 gnd.n4773 19.3944
R9309 gnd.n4773 gnd.n1389 19.3944
R9310 gnd.n4768 gnd.n1389 19.3944
R9311 gnd.n4768 gnd.n4767 19.3944
R9312 gnd.n4767 gnd.n4766 19.3944
R9313 gnd.n4766 gnd.n1396 19.3944
R9314 gnd.n4761 gnd.n1396 19.3944
R9315 gnd.n4761 gnd.n4760 19.3944
R9316 gnd.n4760 gnd.n4759 19.3944
R9317 gnd.n4759 gnd.n1403 19.3944
R9318 gnd.n4754 gnd.n1403 19.3944
R9319 gnd.n4754 gnd.n4753 19.3944
R9320 gnd.n2408 gnd.n2368 19.3944
R9321 gnd.n2412 gnd.n2368 19.3944
R9322 gnd.n2412 gnd.n2366 19.3944
R9323 gnd.n2418 gnd.n2366 19.3944
R9324 gnd.n2418 gnd.n2364 19.3944
R9325 gnd.n2422 gnd.n2364 19.3944
R9326 gnd.n2422 gnd.n2362 19.3944
R9327 gnd.n2428 gnd.n2362 19.3944
R9328 gnd.n2428 gnd.n2360 19.3944
R9329 gnd.n2432 gnd.n2360 19.3944
R9330 gnd.n2432 gnd.n2358 19.3944
R9331 gnd.n2438 gnd.n2358 19.3944
R9332 gnd.n2438 gnd.n2356 19.3944
R9333 gnd.n2442 gnd.n2356 19.3944
R9334 gnd.n2442 gnd.n2354 19.3944
R9335 gnd.n2448 gnd.n2354 19.3944
R9336 gnd.n2448 gnd.n2352 19.3944
R9337 gnd.n2452 gnd.n2352 19.3944
R9338 gnd.n2381 gnd.n1425 19.3944
R9339 gnd.n2388 gnd.n2381 19.3944
R9340 gnd.n2388 gnd.n2378 19.3944
R9341 gnd.n2392 gnd.n2378 19.3944
R9342 gnd.n2392 gnd.n2376 19.3944
R9343 gnd.n2398 gnd.n2376 19.3944
R9344 gnd.n2398 gnd.n2374 19.3944
R9345 gnd.n2402 gnd.n2374 19.3944
R9346 gnd.n4751 gnd.n1412 19.3944
R9347 gnd.n4746 gnd.n1412 19.3944
R9348 gnd.n4746 gnd.n4745 19.3944
R9349 gnd.n4745 gnd.n4744 19.3944
R9350 gnd.n4744 gnd.n1419 19.3944
R9351 gnd.n4739 gnd.n1419 19.3944
R9352 gnd.n4739 gnd.n4738 19.3944
R9353 gnd.n4920 gnd.n1145 19.3944
R9354 gnd.n4920 gnd.n4919 19.3944
R9355 gnd.n4919 gnd.n4918 19.3944
R9356 gnd.n4918 gnd.n1150 19.3944
R9357 gnd.n4908 gnd.n1150 19.3944
R9358 gnd.n4908 gnd.n4907 19.3944
R9359 gnd.n4907 gnd.n4906 19.3944
R9360 gnd.n4906 gnd.n1173 19.3944
R9361 gnd.n4896 gnd.n1173 19.3944
R9362 gnd.n4896 gnd.n4895 19.3944
R9363 gnd.n4895 gnd.n4894 19.3944
R9364 gnd.n4894 gnd.n1192 19.3944
R9365 gnd.n4884 gnd.n1192 19.3944
R9366 gnd.n4884 gnd.n4883 19.3944
R9367 gnd.n4883 gnd.n4882 19.3944
R9368 gnd.n4882 gnd.n1213 19.3944
R9369 gnd.n4872 gnd.n1213 19.3944
R9370 gnd.n4872 gnd.n4871 19.3944
R9371 gnd.n4871 gnd.n4870 19.3944
R9372 gnd.n4870 gnd.n1233 19.3944
R9373 gnd.n4860 gnd.n1233 19.3944
R9374 gnd.n4860 gnd.n4859 19.3944
R9375 gnd.n1258 gnd.n1252 19.3944
R9376 gnd.n2624 gnd.n1258 19.3944
R9377 gnd.n2887 gnd.n2886 19.3944
R9378 gnd.n2901 gnd.n2900 19.3944
R9379 gnd.n4856 gnd.n1259 19.3944
R9380 gnd.n4856 gnd.n1260 19.3944
R9381 gnd.n4846 gnd.n1260 19.3944
R9382 gnd.n4846 gnd.n4845 19.3944
R9383 gnd.n4845 gnd.n4844 19.3944
R9384 gnd.n4844 gnd.n1281 19.3944
R9385 gnd.n4834 gnd.n1281 19.3944
R9386 gnd.n4834 gnd.n4833 19.3944
R9387 gnd.n4833 gnd.n4832 19.3944
R9388 gnd.n4832 gnd.n1302 19.3944
R9389 gnd.n4822 gnd.n1302 19.3944
R9390 gnd.n4822 gnd.n4821 19.3944
R9391 gnd.n4821 gnd.n4820 19.3944
R9392 gnd.n4820 gnd.n1321 19.3944
R9393 gnd.n4810 gnd.n1321 19.3944
R9394 gnd.n4810 gnd.n4809 19.3944
R9395 gnd.n4809 gnd.n4808 19.3944
R9396 gnd.n4808 gnd.n1342 19.3944
R9397 gnd.n4798 gnd.n1342 19.3944
R9398 gnd.n4798 gnd.n4797 19.3944
R9399 gnd.n4797 gnd.n4796 19.3944
R9400 gnd.n4796 gnd.n1362 19.3944
R9401 gnd.n4786 gnd.n1362 19.3944
R9402 gnd.n6629 gnd.n6628 19.3944
R9403 gnd.n6628 gnd.n6627 19.3944
R9404 gnd.n6627 gnd.n806 19.3944
R9405 gnd.n6621 gnd.n806 19.3944
R9406 gnd.n6621 gnd.n6620 19.3944
R9407 gnd.n6620 gnd.n6619 19.3944
R9408 gnd.n6619 gnd.n814 19.3944
R9409 gnd.n6613 gnd.n814 19.3944
R9410 gnd.n6613 gnd.n6612 19.3944
R9411 gnd.n6612 gnd.n6611 19.3944
R9412 gnd.n6611 gnd.n822 19.3944
R9413 gnd.n6605 gnd.n822 19.3944
R9414 gnd.n6605 gnd.n6604 19.3944
R9415 gnd.n6604 gnd.n6603 19.3944
R9416 gnd.n6603 gnd.n830 19.3944
R9417 gnd.n6597 gnd.n830 19.3944
R9418 gnd.n6597 gnd.n6596 19.3944
R9419 gnd.n6596 gnd.n6595 19.3944
R9420 gnd.n6595 gnd.n838 19.3944
R9421 gnd.n6589 gnd.n838 19.3944
R9422 gnd.n6589 gnd.n6588 19.3944
R9423 gnd.n6588 gnd.n6587 19.3944
R9424 gnd.n6587 gnd.n846 19.3944
R9425 gnd.n6581 gnd.n846 19.3944
R9426 gnd.n6581 gnd.n6580 19.3944
R9427 gnd.n6580 gnd.n6579 19.3944
R9428 gnd.n6579 gnd.n854 19.3944
R9429 gnd.n6573 gnd.n854 19.3944
R9430 gnd.n6573 gnd.n6572 19.3944
R9431 gnd.n6572 gnd.n6571 19.3944
R9432 gnd.n6571 gnd.n862 19.3944
R9433 gnd.n6565 gnd.n862 19.3944
R9434 gnd.n6565 gnd.n6564 19.3944
R9435 gnd.n6564 gnd.n6563 19.3944
R9436 gnd.n6563 gnd.n870 19.3944
R9437 gnd.n6557 gnd.n870 19.3944
R9438 gnd.n6557 gnd.n6556 19.3944
R9439 gnd.n6556 gnd.n6555 19.3944
R9440 gnd.n6555 gnd.n878 19.3944
R9441 gnd.n6549 gnd.n878 19.3944
R9442 gnd.n6549 gnd.n6548 19.3944
R9443 gnd.n6548 gnd.n6547 19.3944
R9444 gnd.n6547 gnd.n886 19.3944
R9445 gnd.n6541 gnd.n886 19.3944
R9446 gnd.n6541 gnd.n6540 19.3944
R9447 gnd.n6540 gnd.n6539 19.3944
R9448 gnd.n6539 gnd.n894 19.3944
R9449 gnd.n6533 gnd.n894 19.3944
R9450 gnd.n6533 gnd.n6532 19.3944
R9451 gnd.n6532 gnd.n6531 19.3944
R9452 gnd.n6531 gnd.n902 19.3944
R9453 gnd.n6525 gnd.n902 19.3944
R9454 gnd.n6525 gnd.n6524 19.3944
R9455 gnd.n6524 gnd.n6523 19.3944
R9456 gnd.n6523 gnd.n910 19.3944
R9457 gnd.n6517 gnd.n910 19.3944
R9458 gnd.n6517 gnd.n6516 19.3944
R9459 gnd.n6516 gnd.n6515 19.3944
R9460 gnd.n6515 gnd.n918 19.3944
R9461 gnd.n6509 gnd.n918 19.3944
R9462 gnd.n6509 gnd.n6508 19.3944
R9463 gnd.n6508 gnd.n6507 19.3944
R9464 gnd.n6507 gnd.n926 19.3944
R9465 gnd.n6501 gnd.n926 19.3944
R9466 gnd.n6501 gnd.n6500 19.3944
R9467 gnd.n6500 gnd.n6499 19.3944
R9468 gnd.n6499 gnd.n934 19.3944
R9469 gnd.n6493 gnd.n934 19.3944
R9470 gnd.n6493 gnd.n6492 19.3944
R9471 gnd.n6492 gnd.n6491 19.3944
R9472 gnd.n6491 gnd.n942 19.3944
R9473 gnd.n6485 gnd.n942 19.3944
R9474 gnd.n6485 gnd.n6484 19.3944
R9475 gnd.n6484 gnd.n6483 19.3944
R9476 gnd.n6483 gnd.n950 19.3944
R9477 gnd.n6477 gnd.n950 19.3944
R9478 gnd.n6477 gnd.n6476 19.3944
R9479 gnd.n6476 gnd.n6475 19.3944
R9480 gnd.n6475 gnd.n958 19.3944
R9481 gnd.n6469 gnd.n958 19.3944
R9482 gnd.n6469 gnd.n6468 19.3944
R9483 gnd.n6468 gnd.n6467 19.3944
R9484 gnd.n6467 gnd.n966 19.3944
R9485 gnd.n2787 gnd.n966 19.3944
R9486 gnd.n3142 gnd.n2337 19.3944
R9487 gnd.n2337 gnd.n2316 19.3944
R9488 gnd.n3167 gnd.n2316 19.3944
R9489 gnd.n3167 gnd.n2313 19.3944
R9490 gnd.n3172 gnd.n2313 19.3944
R9491 gnd.n3172 gnd.n2314 19.3944
R9492 gnd.n2314 gnd.n2291 19.3944
R9493 gnd.n3197 gnd.n2291 19.3944
R9494 gnd.n3197 gnd.n2288 19.3944
R9495 gnd.n3202 gnd.n2288 19.3944
R9496 gnd.n3202 gnd.n2289 19.3944
R9497 gnd.n2289 gnd.n2266 19.3944
R9498 gnd.n3237 gnd.n2266 19.3944
R9499 gnd.n3237 gnd.n2263 19.3944
R9500 gnd.n3242 gnd.n2263 19.3944
R9501 gnd.n3242 gnd.n2264 19.3944
R9502 gnd.n2264 gnd.n1496 19.3944
R9503 gnd.n4660 gnd.n1496 19.3944
R9504 gnd.n4660 gnd.n1497 19.3944
R9505 gnd.n4656 gnd.n1497 19.3944
R9506 gnd.n4656 gnd.n4655 19.3944
R9507 gnd.n4655 gnd.n4654 19.3944
R9508 gnd.n4654 gnd.n1503 19.3944
R9509 gnd.n4650 gnd.n1503 19.3944
R9510 gnd.n4650 gnd.n4649 19.3944
R9511 gnd.n4649 gnd.n4648 19.3944
R9512 gnd.n4648 gnd.n1508 19.3944
R9513 gnd.n4644 gnd.n1508 19.3944
R9514 gnd.n4644 gnd.n4643 19.3944
R9515 gnd.n4643 gnd.n4642 19.3944
R9516 gnd.n4642 gnd.n1513 19.3944
R9517 gnd.n4638 gnd.n1513 19.3944
R9518 gnd.n4638 gnd.n4637 19.3944
R9519 gnd.n4637 gnd.n4636 19.3944
R9520 gnd.n4636 gnd.n1518 19.3944
R9521 gnd.n4632 gnd.n1518 19.3944
R9522 gnd.n4632 gnd.n4631 19.3944
R9523 gnd.n4631 gnd.n4630 19.3944
R9524 gnd.n4630 gnd.n1523 19.3944
R9525 gnd.n4626 gnd.n1523 19.3944
R9526 gnd.n4626 gnd.n4625 19.3944
R9527 gnd.n4625 gnd.n4624 19.3944
R9528 gnd.n4624 gnd.n1528 19.3944
R9529 gnd.n4620 gnd.n1528 19.3944
R9530 gnd.n4620 gnd.n4619 19.3944
R9531 gnd.n4619 gnd.n4618 19.3944
R9532 gnd.n4618 gnd.n1533 19.3944
R9533 gnd.n4614 gnd.n1533 19.3944
R9534 gnd.n4614 gnd.n4613 19.3944
R9535 gnd.n4613 gnd.n4612 19.3944
R9536 gnd.n4612 gnd.n1538 19.3944
R9537 gnd.n4608 gnd.n1538 19.3944
R9538 gnd.n4608 gnd.n4607 19.3944
R9539 gnd.n4607 gnd.n4606 19.3944
R9540 gnd.n4606 gnd.n1543 19.3944
R9541 gnd.n4602 gnd.n1543 19.3944
R9542 gnd.n4602 gnd.n4601 19.3944
R9543 gnd.n4601 gnd.n4600 19.3944
R9544 gnd.n4600 gnd.n1548 19.3944
R9545 gnd.n4596 gnd.n1548 19.3944
R9546 gnd.n4596 gnd.n4595 19.3944
R9547 gnd.n4595 gnd.n4594 19.3944
R9548 gnd.n4594 gnd.n1553 19.3944
R9549 gnd.n4590 gnd.n1553 19.3944
R9550 gnd.n4590 gnd.n4589 19.3944
R9551 gnd.n4589 gnd.n4588 19.3944
R9552 gnd.n4588 gnd.n1558 19.3944
R9553 gnd.n4584 gnd.n1558 19.3944
R9554 gnd.n4584 gnd.n4583 19.3944
R9555 gnd.n4583 gnd.n4582 19.3944
R9556 gnd.n4582 gnd.n1563 19.3944
R9557 gnd.n4578 gnd.n1563 19.3944
R9558 gnd.n4578 gnd.n4577 19.3944
R9559 gnd.n4577 gnd.n4576 19.3944
R9560 gnd.n4576 gnd.n1568 19.3944
R9561 gnd.n4572 gnd.n1568 19.3944
R9562 gnd.n4572 gnd.n4571 19.3944
R9563 gnd.n4571 gnd.n4570 19.3944
R9564 gnd.n4570 gnd.n1573 19.3944
R9565 gnd.n4566 gnd.n1573 19.3944
R9566 gnd.n4566 gnd.n4565 19.3944
R9567 gnd.n4565 gnd.n4564 19.3944
R9568 gnd.n3819 gnd.n3816 19.3944
R9569 gnd.n3819 gnd.n3814 19.3944
R9570 gnd.n3825 gnd.n3814 19.3944
R9571 gnd.n3825 gnd.n3812 19.3944
R9572 gnd.n3830 gnd.n3812 19.3944
R9573 gnd.n3830 gnd.n3810 19.3944
R9574 gnd.n3836 gnd.n3810 19.3944
R9575 gnd.n3836 gnd.n3809 19.3944
R9576 gnd.n3845 gnd.n3809 19.3944
R9577 gnd.n3845 gnd.n3807 19.3944
R9578 gnd.n3851 gnd.n3807 19.3944
R9579 gnd.n3851 gnd.n3800 19.3944
R9580 gnd.n3864 gnd.n3800 19.3944
R9581 gnd.n3864 gnd.n3798 19.3944
R9582 gnd.n3870 gnd.n3798 19.3944
R9583 gnd.n3870 gnd.n3791 19.3944
R9584 gnd.n3883 gnd.n3791 19.3944
R9585 gnd.n3883 gnd.n3789 19.3944
R9586 gnd.n3889 gnd.n3789 19.3944
R9587 gnd.n3889 gnd.n3782 19.3944
R9588 gnd.n3902 gnd.n3782 19.3944
R9589 gnd.n3902 gnd.n3780 19.3944
R9590 gnd.n3909 gnd.n3780 19.3944
R9591 gnd.n3909 gnd.n3908 19.3944
R9592 gnd.n3922 gnd.n3761 19.3944
R9593 gnd.n3761 gnd.n3760 19.3944
R9594 gnd.n3929 gnd.n3760 19.3944
R9595 gnd.n5834 gnd.t325 18.8012
R9596 gnd.n5873 gnd.t235 18.8012
R9597 gnd.n5677 gnd.n5419 18.4825
R9598 gnd.n6463 gnd.n968 18.4825
R9599 gnd.n4241 gnd.n4149 18.4247
R9600 gnd.n4738 gnd.n4737 18.4247
R9601 gnd.n3919 gnd.n3918 18.2308
R9602 gnd.n3081 gnd.n3080 18.2308
R9603 gnd.n7414 gnd.n7413 18.2308
R9604 gnd.n2740 gnd.n2739 18.2308
R9605 gnd.t324 gnd.n5361 18.1639
R9606 gnd.n1184 gnd.n1177 18.1639
R9607 gnd.n7581 gnd.n172 18.1639
R9608 gnd.n4667 gnd.n4666 17.9517
R9609 gnd.n4076 gnd.n4075 17.9517
R9610 gnd.n5390 gnd.t305 17.5266
R9611 gnd.t53 gnd.n1167 17.5266
R9612 gnd.n4806 gnd.t2 17.5266
R9613 gnd.n4528 gnd.t16 17.5266
R9614 gnd.n7575 gnd.t297 17.5266
R9615 gnd.t319 gnd.n5337 16.8893
R9616 gnd.n4830 gnd.t206 16.8893
R9617 gnd.n4504 gnd.t71 16.8893
R9618 gnd.n4271 gnd.n1833 16.6793
R9619 gnd.n7486 gnd.n7485 16.6793
R9620 gnd.n4973 gnd.n4970 16.6793
R9621 gnd.n2402 gnd.n2372 16.6793
R9622 gnd.t85 gnd.n5446 16.2519
R9623 gnd.n5304 gnd.t321 16.2519
R9624 gnd.n4854 gnd.t63 16.2519
R9625 gnd.n4480 gnd.t0 16.2519
R9626 gnd.n3070 gnd.n2530 15.9333
R9627 gnd.n3070 gnd.n3068 15.9333
R9628 gnd.n3144 gnd.n2333 15.9333
R9629 gnd.n3144 gnd.n2334 15.9333
R9630 gnd.n2334 gnd.n2327 15.9333
R9631 gnd.n3154 gnd.n2327 15.9333
R9632 gnd.n3153 gnd.n2318 15.9333
R9633 gnd.n3165 gnd.n2318 15.9333
R9634 gnd.n3165 gnd.n3164 15.9333
R9635 gnd.n3164 gnd.n2320 15.9333
R9636 gnd.n2320 gnd.n2308 15.9333
R9637 gnd.n3174 gnd.n2308 15.9333
R9638 gnd.n3174 gnd.n2309 15.9333
R9639 gnd.n2311 gnd.n2309 15.9333
R9640 gnd.n3184 gnd.n3183 15.9333
R9641 gnd.n3183 gnd.n2293 15.9333
R9642 gnd.n3195 gnd.n2293 15.9333
R9643 gnd.n3195 gnd.n3194 15.9333
R9644 gnd.n3194 gnd.n2295 15.9333
R9645 gnd.n2295 gnd.n2284 15.9333
R9646 gnd.n3204 gnd.n2284 15.9333
R9647 gnd.n3204 gnd.n2285 15.9333
R9648 gnd.n3214 gnd.n2277 15.9333
R9649 gnd.n3214 gnd.n3213 15.9333
R9650 gnd.n3213 gnd.n2268 15.9333
R9651 gnd.n3235 gnd.n2268 15.9333
R9652 gnd.n3235 gnd.n3234 15.9333
R9653 gnd.n3234 gnd.n2270 15.9333
R9654 gnd.n2270 gnd.n2259 15.9333
R9655 gnd.n3244 gnd.n2259 15.9333
R9656 gnd.n3244 gnd.n2260 15.9333
R9657 gnd.n3227 gnd.n1464 15.9333
R9658 gnd.n3256 gnd.n1490 15.9333
R9659 gnd.n3289 gnd.n2183 15.9333
R9660 gnd.n3300 gnd.n3299 15.9333
R9661 gnd.n3419 gnd.n2113 15.9333
R9662 gnd.n3438 gnd.n2090 15.9333
R9663 gnd.n2097 gnd.n2085 15.9333
R9664 gnd.n3478 gnd.n2068 15.9333
R9665 gnd.n3525 gnd.n3524 15.9333
R9666 gnd.n3533 gnd.n2055 15.9333
R9667 gnd.n3550 gnd.n3549 15.9333
R9668 gnd.n3610 gnd.n2023 15.9333
R9669 gnd.n3684 gnd.n3683 15.9333
R9670 gnd.n3698 gnd.n1965 15.9333
R9671 gnd.n3716 gnd.n1951 15.9333
R9672 gnd.n1884 gnd.n1846 15.9333
R9673 gnd.n3979 gnd.n3978 15.9333
R9674 gnd.n3978 gnd.n3976 15.9333
R9675 gnd.n3976 gnd.n3975 15.9333
R9676 gnd.n3975 gnd.n3974 15.9333
R9677 gnd.n3974 gnd.n1902 15.9333
R9678 gnd.n1910 gnd.n1902 15.9333
R9679 gnd.n1911 gnd.n1910 15.9333
R9680 gnd.n3968 gnd.n1911 15.9333
R9681 gnd.n3968 gnd.n3967 15.9333
R9682 gnd.n3965 gnd.n3964 15.9333
R9683 gnd.n3964 gnd.n3963 15.9333
R9684 gnd.n3963 gnd.n1914 15.9333
R9685 gnd.n1922 gnd.n1914 15.9333
R9686 gnd.n1923 gnd.n1922 15.9333
R9687 gnd.n3957 gnd.n1923 15.9333
R9688 gnd.n3957 gnd.n3956 15.9333
R9689 gnd.n3956 gnd.n3954 15.9333
R9690 gnd.n3953 gnd.n3952 15.9333
R9691 gnd.n3952 gnd.n1926 15.9333
R9692 gnd.n1934 gnd.n1926 15.9333
R9693 gnd.n1935 gnd.n1934 15.9333
R9694 gnd.n3946 gnd.n1935 15.9333
R9695 gnd.n3946 gnd.n3945 15.9333
R9696 gnd.n3945 gnd.n3943 15.9333
R9697 gnd.n3943 gnd.n3942 15.9333
R9698 gnd.n3941 gnd.n3935 15.9333
R9699 gnd.n3935 gnd.n1579 15.9333
R9700 gnd.n4562 gnd.n1579 15.9333
R9701 gnd.n4562 gnd.n4561 15.9333
R9702 gnd.n1590 gnd.n1581 15.9333
R9703 gnd.n4555 gnd.n1590 15.9333
R9704 gnd.n6273 gnd.n6271 15.6674
R9705 gnd.n6241 gnd.n6239 15.6674
R9706 gnd.n6209 gnd.n6207 15.6674
R9707 gnd.n6178 gnd.n6176 15.6674
R9708 gnd.n6146 gnd.n6144 15.6674
R9709 gnd.n6114 gnd.n6112 15.6674
R9710 gnd.n6082 gnd.n6080 15.6674
R9711 gnd.n6051 gnd.n6049 15.6674
R9712 gnd.n5564 gnd.t85 15.6146
R9713 gnd.t81 gnd.n6434 15.6146
R9714 gnd.n6338 gnd.t179 15.6146
R9715 gnd.t248 gnd.n2860 15.6146
R9716 gnd.t141 gnd.n3153 15.6146
R9717 gnd.n3942 gnd.t124 15.6146
R9718 gnd.n7328 gnd.t29 15.6146
R9719 gnd.n4323 gnd.n1812 15.3217
R9720 gnd.n7446 gnd.n315 15.3217
R9721 gnd.n4930 gnd.n1133 15.3217
R9722 gnd.n2457 gnd.n2350 15.3217
R9723 gnd.n3330 gnd.n2168 15.296
R9724 gnd.n3349 gnd.n2159 15.296
R9725 gnd.n3309 gnd.t316 15.296
R9726 gnd.n3479 gnd.n3477 15.296
R9727 gnd.n3523 gnd.n2064 15.296
R9728 gnd.n3651 gnd.t66 15.296
R9729 gnd.n3590 gnd.n1988 15.296
R9730 gnd.n3681 gnd.n1975 15.296
R9731 gnd.n3996 gnd.n3995 15.0827
R9732 gnd.n1476 gnd.n1471 15.0481
R9733 gnd.n4006 gnd.n4005 15.0481
R9734 gnd.n6002 gnd.t294 14.9773
R9735 gnd.n4880 gnd.t56 14.9773
R9736 gnd.n2285 gnd.t255 14.9773
R9737 gnd.t31 gnd.n3965 14.9773
R9738 gnd.n7356 gnd.t58 14.9773
R9739 gnd.n4663 gnd.n4662 14.6587
R9740 gnd.n3390 gnd.n3389 14.6587
R9741 gnd.n2016 gnd.n2005 14.6587
R9742 gnd.n3987 gnd.n3986 14.6587
R9743 gnd.n6455 gnd.t257 14.34
R9744 gnd.t307 gnd.n993 14.34
R9745 gnd.n4904 gnd.t53 14.34
R9746 gnd.t297 gnd.n175 14.34
R9747 gnd.n3273 gnd.n2175 14.0214
R9748 gnd.n3307 gnd.n2144 14.0214
R9749 gnd.n3469 gnd.n3468 14.0214
R9750 gnd.n2054 gnd.n2047 14.0214
R9751 gnd.n3652 gnd.n1992 14.0214
R9752 gnd.t270 gnd.n5761 13.7027
R9753 gnd.n4898 gnd.n1184 13.7027
R9754 gnd.n2117 gnd.t208 13.7027
R9755 gnd.n3558 gnd.t231 13.7027
R9756 gnd.n7392 gnd.n172 13.7027
R9757 gnd.n5646 gnd.n5642 13.5763
R9758 gnd.n6394 gnd.n5079 13.5763
R9759 gnd.n5678 gnd.n5677 13.384
R9760 gnd.n3288 gnd.n2185 13.384
R9761 gnd.n2145 gnd.n2139 13.384
R9762 gnd.t315 gnd.n3377 13.384
R9763 gnd.n3629 gnd.t35 13.384
R9764 gnd.n3638 gnd.n2001 13.384
R9765 gnd.n1958 gnd.n1957 13.384
R9766 gnd.n1487 gnd.n1468 13.1884
R9767 gnd.n1482 gnd.n1481 13.1884
R9768 gnd.n1481 gnd.n1480 13.1884
R9769 gnd.n3999 gnd.n3994 13.1884
R9770 gnd.n4000 gnd.n3999 13.1884
R9771 gnd.n1483 gnd.n1470 13.146
R9772 gnd.n1479 gnd.n1470 13.146
R9773 gnd.n3998 gnd.n3997 13.146
R9774 gnd.n3998 gnd.n3993 13.146
R9775 gnd.n6274 gnd.n6270 12.8005
R9776 gnd.n6242 gnd.n6238 12.8005
R9777 gnd.n6210 gnd.n6206 12.8005
R9778 gnd.n6179 gnd.n6175 12.8005
R9779 gnd.n6147 gnd.n6143 12.8005
R9780 gnd.n6115 gnd.n6111 12.8005
R9781 gnd.n6083 gnd.n6079 12.8005
R9782 gnd.n6052 gnd.n6048 12.8005
R9783 gnd.n3264 gnd.n3263 12.7467
R9784 gnd.n3439 gnd.n3437 12.7467
R9785 gnd.n3548 gnd.n2034 12.7467
R9786 gnd.n1964 gnd.t97 12.7467
R9787 gnd.n5649 gnd.n5646 12.4126
R9788 gnd.n6399 gnd.n5079 12.4126
R9789 gnd.n4730 gnd.n4667 12.1761
R9790 gnd.n4075 gnd.n4074 12.1761
R9791 gnd.n3360 gnd.n2150 12.1094
R9792 gnd.n3659 gnd.n1986 12.1094
R9793 gnd.n3699 gnd.n1962 12.1094
R9794 gnd.t170 gnd.n1889 12.1094
R9795 gnd.n6278 gnd.n6277 12.0247
R9796 gnd.n6246 gnd.n6245 12.0247
R9797 gnd.n6214 gnd.n6213 12.0247
R9798 gnd.n6183 gnd.n6182 12.0247
R9799 gnd.n6151 gnd.n6150 12.0247
R9800 gnd.n6119 gnd.n6118 12.0247
R9801 gnd.n6087 gnd.n6086 12.0247
R9802 gnd.n6056 gnd.n6055 12.0247
R9803 gnd.n2818 gnd.t56 11.7908
R9804 gnd.t58 gnd.n143 11.7908
R9805 gnd.n3057 gnd.n1381 11.4721
R9806 gnd.n3399 gnd.t266 11.4721
R9807 gnd.n3397 gnd.n2126 11.4721
R9808 gnd.n3429 gnd.n3428 11.4721
R9809 gnd.n3576 gnd.n2029 11.4721
R9810 gnd.n3568 gnd.n2015 11.4721
R9811 gnd.n3620 gnd.t314 11.4721
R9812 gnd.n4078 gnd.n1884 11.4721
R9813 gnd.n4553 gnd.n1591 11.4721
R9814 gnd.n6281 gnd.n6268 11.249
R9815 gnd.n6249 gnd.n6236 11.249
R9816 gnd.n6217 gnd.n6204 11.249
R9817 gnd.n6186 gnd.n6173 11.249
R9818 gnd.n6154 gnd.n6141 11.249
R9819 gnd.n6122 gnd.n6109 11.249
R9820 gnd.n6090 gnd.n6077 11.249
R9821 gnd.n6059 gnd.n6046 11.249
R9822 gnd.n5762 gnd.t270 11.1535
R9823 gnd.n2861 gnd.t248 11.1535
R9824 gnd.n2311 gnd.t262 11.1535
R9825 gnd.n3376 gnd.t354 11.1535
R9826 gnd.t264 gnd.n3630 11.1535
R9827 gnd.t50 gnd.n3953 11.1535
R9828 gnd.t29 gnd.n102 11.1535
R9829 gnd.n3329 gnd.t158 10.8348
R9830 gnd.n3343 gnd.n3342 10.8348
R9831 gnd.n3342 gnd.n3341 10.8348
R9832 gnd.n3517 gnd.n3516 10.8348
R9833 gnd.n3516 gnd.n2061 10.8348
R9834 gnd.n3675 gnd.n3674 10.8348
R9835 gnd.n3674 gnd.n1972 10.8348
R9836 gnd.n1813 gnd.n1812 10.6672
R9837 gnd.n7451 gnd.n315 10.6672
R9838 gnd.n4933 gnd.n4930 10.6672
R9839 gnd.n2452 gnd.n2350 10.6672
R9840 gnd.n4140 gnd.n1842 10.6151
R9841 gnd.n4140 gnd.n4139 10.6151
R9842 gnd.n4137 gnd.n4134 10.6151
R9843 gnd.n4134 gnd.n4133 10.6151
R9844 gnd.n4133 gnd.n4130 10.6151
R9845 gnd.n4130 gnd.n4129 10.6151
R9846 gnd.n4129 gnd.n4126 10.6151
R9847 gnd.n4126 gnd.n4125 10.6151
R9848 gnd.n4125 gnd.n4122 10.6151
R9849 gnd.n4122 gnd.n4121 10.6151
R9850 gnd.n4121 gnd.n4118 10.6151
R9851 gnd.n4118 gnd.n4117 10.6151
R9852 gnd.n4117 gnd.n4114 10.6151
R9853 gnd.n4114 gnd.n4113 10.6151
R9854 gnd.n4113 gnd.n4110 10.6151
R9855 gnd.n4110 gnd.n4109 10.6151
R9856 gnd.n4109 gnd.n4106 10.6151
R9857 gnd.n4106 gnd.n4105 10.6151
R9858 gnd.n4105 gnd.n4102 10.6151
R9859 gnd.n4102 gnd.n4101 10.6151
R9860 gnd.n4101 gnd.n4098 10.6151
R9861 gnd.n4098 gnd.n4097 10.6151
R9862 gnd.n4097 gnd.n4094 10.6151
R9863 gnd.n4094 gnd.n4093 10.6151
R9864 gnd.n4093 gnd.n4090 10.6151
R9865 gnd.n4090 gnd.n4089 10.6151
R9866 gnd.n4089 gnd.n4086 10.6151
R9867 gnd.n4086 gnd.n4085 10.6151
R9868 gnd.n4085 gnd.n4082 10.6151
R9869 gnd.n4082 gnd.n4081 10.6151
R9870 gnd.n3260 gnd.n3259 10.6151
R9871 gnd.n3261 gnd.n3260 10.6151
R9872 gnd.n3266 gnd.n3261 10.6151
R9873 gnd.n3267 gnd.n3266 10.6151
R9874 gnd.n3271 gnd.n3267 10.6151
R9875 gnd.n3271 gnd.n3270 10.6151
R9876 gnd.n3270 gnd.n3269 10.6151
R9877 gnd.n3269 gnd.n2166 10.6151
R9878 gnd.n3332 gnd.n2166 10.6151
R9879 gnd.n3333 gnd.n3332 10.6151
R9880 gnd.n3339 gnd.n3333 10.6151
R9881 gnd.n3339 gnd.n3338 10.6151
R9882 gnd.n3338 gnd.n3337 10.6151
R9883 gnd.n3337 gnd.n3334 10.6151
R9884 gnd.n3334 gnd.n2142 10.6151
R9885 gnd.n3369 gnd.n2142 10.6151
R9886 gnd.n3370 gnd.n3369 10.6151
R9887 gnd.n3374 gnd.n3370 10.6151
R9888 gnd.n3374 gnd.n3373 10.6151
R9889 gnd.n3373 gnd.n3372 10.6151
R9890 gnd.n3372 gnd.n3371 10.6151
R9891 gnd.n3371 gnd.n2116 10.6151
R9892 gnd.n3417 gnd.n2116 10.6151
R9893 gnd.n3417 gnd.n3416 10.6151
R9894 gnd.n3416 gnd.n3415 10.6151
R9895 gnd.n3415 gnd.n3414 10.6151
R9896 gnd.n3414 gnd.n2098 10.6151
R9897 gnd.n3441 gnd.n2098 10.6151
R9898 gnd.n3442 gnd.n3441 10.6151
R9899 gnd.n3444 gnd.n3442 10.6151
R9900 gnd.n3445 gnd.n3444 10.6151
R9901 gnd.n3446 gnd.n3445 10.6151
R9902 gnd.n3446 gnd.n2075 10.6151
R9903 gnd.n3481 gnd.n2075 10.6151
R9904 gnd.n3482 gnd.n3481 10.6151
R9905 gnd.n3484 gnd.n3482 10.6151
R9906 gnd.n3485 gnd.n3484 10.6151
R9907 gnd.n3487 gnd.n3485 10.6151
R9908 gnd.n3487 gnd.n3486 10.6151
R9909 gnd.n3486 gnd.n2045 10.6151
R9910 gnd.n3543 gnd.n2045 10.6151
R9911 gnd.n3544 gnd.n3543 10.6151
R9912 gnd.n3546 gnd.n3544 10.6151
R9913 gnd.n3546 gnd.n3545 10.6151
R9914 gnd.n3545 gnd.n2026 10.6151
R9915 gnd.n3578 gnd.n2026 10.6151
R9916 gnd.n3579 gnd.n3578 10.6151
R9917 gnd.n3608 gnd.n3579 10.6151
R9918 gnd.n3608 gnd.n3607 10.6151
R9919 gnd.n3607 gnd.n3606 10.6151
R9920 gnd.n3606 gnd.n3603 10.6151
R9921 gnd.n3603 gnd.n3602 10.6151
R9922 gnd.n3602 gnd.n3601 10.6151
R9923 gnd.n3601 gnd.n3600 10.6151
R9924 gnd.n3600 gnd.n3599 10.6151
R9925 gnd.n3599 gnd.n3596 10.6151
R9926 gnd.n3596 gnd.n3595 10.6151
R9927 gnd.n3595 gnd.n3593 10.6151
R9928 gnd.n3593 gnd.n3592 10.6151
R9929 gnd.n3592 gnd.n3587 10.6151
R9930 gnd.n3587 gnd.n3586 10.6151
R9931 gnd.n3586 gnd.n3584 10.6151
R9932 gnd.n3584 gnd.n3583 10.6151
R9933 gnd.n3583 gnd.n3580 10.6151
R9934 gnd.n3580 gnd.n1953 10.6151
R9935 gnd.n3708 gnd.n1953 10.6151
R9936 gnd.n3709 gnd.n3708 10.6151
R9937 gnd.n3712 gnd.n3709 10.6151
R9938 gnd.n3712 gnd.n3711 10.6151
R9939 gnd.n3711 gnd.n3710 10.6151
R9940 gnd.n3710 gnd.n1881 10.6151
R9941 gnd.n2190 gnd.n1429 10.6151
R9942 gnd.n2193 gnd.n2190 10.6151
R9943 gnd.n2198 gnd.n2195 10.6151
R9944 gnd.n2199 gnd.n2198 10.6151
R9945 gnd.n2202 gnd.n2199 10.6151
R9946 gnd.n2203 gnd.n2202 10.6151
R9947 gnd.n2206 gnd.n2203 10.6151
R9948 gnd.n2207 gnd.n2206 10.6151
R9949 gnd.n2210 gnd.n2207 10.6151
R9950 gnd.n2211 gnd.n2210 10.6151
R9951 gnd.n2214 gnd.n2211 10.6151
R9952 gnd.n2215 gnd.n2214 10.6151
R9953 gnd.n2218 gnd.n2215 10.6151
R9954 gnd.n2219 gnd.n2218 10.6151
R9955 gnd.n2222 gnd.n2219 10.6151
R9956 gnd.n2223 gnd.n2222 10.6151
R9957 gnd.n2226 gnd.n2223 10.6151
R9958 gnd.n2227 gnd.n2226 10.6151
R9959 gnd.n2230 gnd.n2227 10.6151
R9960 gnd.n2231 gnd.n2230 10.6151
R9961 gnd.n2234 gnd.n2231 10.6151
R9962 gnd.n2235 gnd.n2234 10.6151
R9963 gnd.n2238 gnd.n2235 10.6151
R9964 gnd.n2239 gnd.n2238 10.6151
R9965 gnd.n2242 gnd.n2239 10.6151
R9966 gnd.n2243 gnd.n2242 10.6151
R9967 gnd.n2246 gnd.n2243 10.6151
R9968 gnd.n2247 gnd.n2246 10.6151
R9969 gnd.n2250 gnd.n2247 10.6151
R9970 gnd.n2251 gnd.n2250 10.6151
R9971 gnd.n4730 gnd.n4729 10.6151
R9972 gnd.n4729 gnd.n4728 10.6151
R9973 gnd.n4728 gnd.n4727 10.6151
R9974 gnd.n4727 gnd.n4725 10.6151
R9975 gnd.n4725 gnd.n4722 10.6151
R9976 gnd.n4722 gnd.n4721 10.6151
R9977 gnd.n4721 gnd.n4718 10.6151
R9978 gnd.n4718 gnd.n4717 10.6151
R9979 gnd.n4717 gnd.n4714 10.6151
R9980 gnd.n4714 gnd.n4713 10.6151
R9981 gnd.n4713 gnd.n4710 10.6151
R9982 gnd.n4710 gnd.n4709 10.6151
R9983 gnd.n4709 gnd.n4706 10.6151
R9984 gnd.n4706 gnd.n4705 10.6151
R9985 gnd.n4705 gnd.n4702 10.6151
R9986 gnd.n4702 gnd.n4701 10.6151
R9987 gnd.n4701 gnd.n4698 10.6151
R9988 gnd.n4698 gnd.n4697 10.6151
R9989 gnd.n4697 gnd.n4694 10.6151
R9990 gnd.n4694 gnd.n4693 10.6151
R9991 gnd.n4693 gnd.n4690 10.6151
R9992 gnd.n4690 gnd.n4689 10.6151
R9993 gnd.n4689 gnd.n4686 10.6151
R9994 gnd.n4686 gnd.n4685 10.6151
R9995 gnd.n4685 gnd.n4682 10.6151
R9996 gnd.n4682 gnd.n4681 10.6151
R9997 gnd.n4681 gnd.n4678 10.6151
R9998 gnd.n4678 gnd.n4677 10.6151
R9999 gnd.n4674 gnd.n4673 10.6151
R10000 gnd.n4673 gnd.n1430 10.6151
R10001 gnd.n4074 gnd.n4073 10.6151
R10002 gnd.n4073 gnd.n4070 10.6151
R10003 gnd.n4070 gnd.n4069 10.6151
R10004 gnd.n4069 gnd.n4066 10.6151
R10005 gnd.n4066 gnd.n4065 10.6151
R10006 gnd.n4065 gnd.n4062 10.6151
R10007 gnd.n4062 gnd.n4061 10.6151
R10008 gnd.n4061 gnd.n4058 10.6151
R10009 gnd.n4058 gnd.n4057 10.6151
R10010 gnd.n4057 gnd.n4054 10.6151
R10011 gnd.n4054 gnd.n4053 10.6151
R10012 gnd.n4053 gnd.n4050 10.6151
R10013 gnd.n4050 gnd.n4049 10.6151
R10014 gnd.n4049 gnd.n4046 10.6151
R10015 gnd.n4046 gnd.n4045 10.6151
R10016 gnd.n4045 gnd.n4042 10.6151
R10017 gnd.n4042 gnd.n4041 10.6151
R10018 gnd.n4041 gnd.n4038 10.6151
R10019 gnd.n4038 gnd.n4037 10.6151
R10020 gnd.n4037 gnd.n4034 10.6151
R10021 gnd.n4034 gnd.n4033 10.6151
R10022 gnd.n4033 gnd.n4030 10.6151
R10023 gnd.n4030 gnd.n4029 10.6151
R10024 gnd.n4029 gnd.n4026 10.6151
R10025 gnd.n4026 gnd.n4025 10.6151
R10026 gnd.n4025 gnd.n4022 10.6151
R10027 gnd.n4022 gnd.n4021 10.6151
R10028 gnd.n4021 gnd.n4018 10.6151
R10029 gnd.n4016 gnd.n4013 10.6151
R10030 gnd.n4013 gnd.n1843 10.6151
R10031 gnd.n4666 gnd.n4665 10.6151
R10032 gnd.n4665 gnd.n1488 10.6151
R10033 gnd.n3276 gnd.n1488 10.6151
R10034 gnd.n3286 gnd.n3276 10.6151
R10035 gnd.n3286 gnd.n3285 10.6151
R10036 gnd.n3285 gnd.n3284 10.6151
R10037 gnd.n3284 gnd.n3277 10.6151
R10038 gnd.n3278 gnd.n3277 10.6151
R10039 gnd.n3278 gnd.n2161 10.6151
R10040 gnd.n3345 gnd.n2161 10.6151
R10041 gnd.n3346 gnd.n3345 10.6151
R10042 gnd.n3347 gnd.n3346 10.6151
R10043 gnd.n3347 gnd.n2148 10.6151
R10044 gnd.n3362 gnd.n2148 10.6151
R10045 gnd.n3363 gnd.n3362 10.6151
R10046 gnd.n3365 gnd.n3363 10.6151
R10047 gnd.n3365 gnd.n3364 10.6151
R10048 gnd.n3364 gnd.n2128 10.6151
R10049 gnd.n3393 gnd.n2128 10.6151
R10050 gnd.n3394 gnd.n3393 10.6151
R10051 gnd.n3395 gnd.n3394 10.6151
R10052 gnd.n3395 gnd.n2111 10.6151
R10053 gnd.n3421 gnd.n2111 10.6151
R10054 gnd.n3422 gnd.n3421 10.6151
R10055 gnd.n3426 gnd.n3422 10.6151
R10056 gnd.n3426 gnd.n3425 10.6151
R10057 gnd.n3425 gnd.n3424 10.6151
R10058 gnd.n3424 gnd.n2088 10.6151
R10059 gnd.n3461 gnd.n2088 10.6151
R10060 gnd.n3462 gnd.n3461 10.6151
R10061 gnd.n3466 gnd.n3462 10.6151
R10062 gnd.n3466 gnd.n3465 10.6151
R10063 gnd.n3465 gnd.n3464 10.6151
R10064 gnd.n3464 gnd.n2066 10.6151
R10065 gnd.n3519 gnd.n2066 10.6151
R10066 gnd.n3520 gnd.n3519 10.6151
R10067 gnd.n3521 gnd.n3520 10.6151
R10068 gnd.n3521 gnd.n2051 10.6151
R10069 gnd.n3536 gnd.n2051 10.6151
R10070 gnd.n3537 gnd.n3536 10.6151
R10071 gnd.n3539 gnd.n3537 10.6151
R10072 gnd.n3539 gnd.n3538 10.6151
R10073 gnd.n3538 gnd.n2032 10.6151
R10074 gnd.n3564 gnd.n2032 10.6151
R10075 gnd.n3565 gnd.n3564 10.6151
R10076 gnd.n3574 gnd.n3565 10.6151
R10077 gnd.n3574 gnd.n3573 10.6151
R10078 gnd.n3573 gnd.n3572 10.6151
R10079 gnd.n3572 gnd.n3571 10.6151
R10080 gnd.n3571 gnd.n3566 10.6151
R10081 gnd.n3566 gnd.n2003 10.6151
R10082 gnd.n3634 gnd.n2003 10.6151
R10083 gnd.n3635 gnd.n3634 10.6151
R10084 gnd.n3636 gnd.n3635 10.6151
R10085 gnd.n3636 gnd.n1990 10.6151
R10086 gnd.n3654 gnd.n1990 10.6151
R10087 gnd.n3655 gnd.n3654 10.6151
R10088 gnd.n3656 gnd.n3655 10.6151
R10089 gnd.n3656 gnd.n1977 10.6151
R10090 gnd.n3677 gnd.n1977 10.6151
R10091 gnd.n3678 gnd.n3677 10.6151
R10092 gnd.n3679 gnd.n3678 10.6151
R10093 gnd.n3679 gnd.n1960 10.6151
R10094 gnd.n3701 gnd.n1960 10.6151
R10095 gnd.n3702 gnd.n3701 10.6151
R10096 gnd.n3704 gnd.n3702 10.6151
R10097 gnd.n3704 gnd.n3703 10.6151
R10098 gnd.n3703 gnd.n1887 10.6151
R10099 gnd.n3990 gnd.n1887 10.6151
R10100 gnd.n3991 gnd.n3990 10.6151
R10101 gnd.n4076 gnd.n3991 10.6151
R10102 gnd.n5434 gnd.t221 10.5161
R10103 gnd.n6320 gnd.t257 10.5161
R10104 gnd.n6327 gnd.t307 10.5161
R10105 gnd.n2940 gnd.t63 10.5161
R10106 gnd.n3351 gnd.t40 10.5161
R10107 gnd.t348 gnd.n3588 10.5161
R10108 gnd.n4457 gnd.t0 10.5161
R10109 gnd.n6282 gnd.n6266 10.4732
R10110 gnd.n6250 gnd.n6234 10.4732
R10111 gnd.n6218 gnd.n6202 10.4732
R10112 gnd.n6187 gnd.n6171 10.4732
R10113 gnd.n6155 gnd.n6139 10.4732
R10114 gnd.n6123 gnd.n6107 10.4732
R10115 gnd.n6091 gnd.n6075 10.4732
R10116 gnd.n6060 gnd.n6044 10.4732
R10117 gnd.n3279 gnd.t195 10.1975
R10118 gnd.n2126 gnd.n2125 10.1975
R10119 gnd.n3429 gnd.n2106 10.1975
R10120 gnd.n3498 gnd.n2029 10.1975
R10121 gnd.n3569 gnd.n3568 10.1975
R10122 gnd.n6019 gnd.t294 9.87883
R10123 gnd.n2978 gnd.t206 9.87883
R10124 gnd.n4366 gnd.t71 9.87883
R10125 gnd.n6286 gnd.n6285 9.69747
R10126 gnd.n6254 gnd.n6253 9.69747
R10127 gnd.n6222 gnd.n6221 9.69747
R10128 gnd.n6191 gnd.n6190 9.69747
R10129 gnd.n6159 gnd.n6158 9.69747
R10130 gnd.n6127 gnd.n6126 9.69747
R10131 gnd.n6095 gnd.n6094 9.69747
R10132 gnd.n6064 gnd.n6063 9.69747
R10133 gnd.n3280 gnd.n3279 9.56018
R10134 gnd.n3335 gnd.n2150 9.56018
R10135 gnd.n3402 gnd.t36 9.56018
R10136 gnd.n3450 gnd.n2077 9.56018
R10137 gnd.n3491 gnd.n3489 9.56018
R10138 gnd.n3499 gnd.t34 9.56018
R10139 gnd.n3659 gnd.n3658 9.56018
R10140 gnd.n6292 gnd.n6291 9.45567
R10141 gnd.n6260 gnd.n6259 9.45567
R10142 gnd.n6228 gnd.n6227 9.45567
R10143 gnd.n6197 gnd.n6196 9.45567
R10144 gnd.n6165 gnd.n6164 9.45567
R10145 gnd.n6133 gnd.n6132 9.45567
R10146 gnd.n6101 gnd.n6100 9.45567
R10147 gnd.n6070 gnd.n6069 9.45567
R10148 gnd.n4271 gnd.n1831 9.30959
R10149 gnd.n7485 gnd.n279 9.30959
R10150 gnd.n4970 gnd.n4969 9.30959
R10151 gnd.n2408 gnd.n2372 9.30959
R10152 gnd.n6291 gnd.n6290 9.3005
R10153 gnd.n6264 gnd.n6263 9.3005
R10154 gnd.n6285 gnd.n6284 9.3005
R10155 gnd.n6283 gnd.n6282 9.3005
R10156 gnd.n6268 gnd.n6267 9.3005
R10157 gnd.n6277 gnd.n6276 9.3005
R10158 gnd.n6275 gnd.n6274 9.3005
R10159 gnd.n6259 gnd.n6258 9.3005
R10160 gnd.n6232 gnd.n6231 9.3005
R10161 gnd.n6253 gnd.n6252 9.3005
R10162 gnd.n6251 gnd.n6250 9.3005
R10163 gnd.n6236 gnd.n6235 9.3005
R10164 gnd.n6245 gnd.n6244 9.3005
R10165 gnd.n6243 gnd.n6242 9.3005
R10166 gnd.n6227 gnd.n6226 9.3005
R10167 gnd.n6200 gnd.n6199 9.3005
R10168 gnd.n6221 gnd.n6220 9.3005
R10169 gnd.n6219 gnd.n6218 9.3005
R10170 gnd.n6204 gnd.n6203 9.3005
R10171 gnd.n6213 gnd.n6212 9.3005
R10172 gnd.n6211 gnd.n6210 9.3005
R10173 gnd.n6196 gnd.n6195 9.3005
R10174 gnd.n6169 gnd.n6168 9.3005
R10175 gnd.n6190 gnd.n6189 9.3005
R10176 gnd.n6188 gnd.n6187 9.3005
R10177 gnd.n6173 gnd.n6172 9.3005
R10178 gnd.n6182 gnd.n6181 9.3005
R10179 gnd.n6180 gnd.n6179 9.3005
R10180 gnd.n6164 gnd.n6163 9.3005
R10181 gnd.n6137 gnd.n6136 9.3005
R10182 gnd.n6158 gnd.n6157 9.3005
R10183 gnd.n6156 gnd.n6155 9.3005
R10184 gnd.n6141 gnd.n6140 9.3005
R10185 gnd.n6150 gnd.n6149 9.3005
R10186 gnd.n6148 gnd.n6147 9.3005
R10187 gnd.n6132 gnd.n6131 9.3005
R10188 gnd.n6105 gnd.n6104 9.3005
R10189 gnd.n6126 gnd.n6125 9.3005
R10190 gnd.n6124 gnd.n6123 9.3005
R10191 gnd.n6109 gnd.n6108 9.3005
R10192 gnd.n6118 gnd.n6117 9.3005
R10193 gnd.n6116 gnd.n6115 9.3005
R10194 gnd.n6100 gnd.n6099 9.3005
R10195 gnd.n6073 gnd.n6072 9.3005
R10196 gnd.n6094 gnd.n6093 9.3005
R10197 gnd.n6092 gnd.n6091 9.3005
R10198 gnd.n6077 gnd.n6076 9.3005
R10199 gnd.n6086 gnd.n6085 9.3005
R10200 gnd.n6084 gnd.n6083 9.3005
R10201 gnd.n6069 gnd.n6068 9.3005
R10202 gnd.n6042 gnd.n6041 9.3005
R10203 gnd.n6063 gnd.n6062 9.3005
R10204 gnd.n6061 gnd.n6060 9.3005
R10205 gnd.n6046 gnd.n6045 9.3005
R10206 gnd.n6055 gnd.n6054 9.3005
R10207 gnd.n6053 gnd.n6052 9.3005
R10208 gnd.n6421 gnd.n5053 9.3005
R10209 gnd.n6420 gnd.n5055 9.3005
R10210 gnd.n5059 gnd.n5056 9.3005
R10211 gnd.n6415 gnd.n5060 9.3005
R10212 gnd.n6414 gnd.n5061 9.3005
R10213 gnd.n6413 gnd.n5062 9.3005
R10214 gnd.n5066 gnd.n5063 9.3005
R10215 gnd.n6408 gnd.n5067 9.3005
R10216 gnd.n6407 gnd.n5068 9.3005
R10217 gnd.n6406 gnd.n5069 9.3005
R10218 gnd.n5073 gnd.n5070 9.3005
R10219 gnd.n6401 gnd.n5074 9.3005
R10220 gnd.n6400 gnd.n5075 9.3005
R10221 gnd.n6399 gnd.n5076 9.3005
R10222 gnd.n5081 gnd.n5079 9.3005
R10223 gnd.n6394 gnd.n6393 9.3005
R10224 gnd.n6423 gnd.n6422 9.3005
R10225 gnd.n5701 gnd.n5700 9.3005
R10226 gnd.n5702 gnd.n5404 9.3005
R10227 gnd.n5704 gnd.n5703 9.3005
R10228 gnd.n5385 gnd.n5384 9.3005
R10229 gnd.n5731 gnd.n5730 9.3005
R10230 gnd.n5732 gnd.n5383 9.3005
R10231 gnd.n5736 gnd.n5733 9.3005
R10232 gnd.n5735 gnd.n5734 9.3005
R10233 gnd.n5359 gnd.n5358 9.3005
R10234 gnd.n5765 gnd.n5764 9.3005
R10235 gnd.n5766 gnd.n5357 9.3005
R10236 gnd.n5773 gnd.n5767 9.3005
R10237 gnd.n5772 gnd.n5768 9.3005
R10238 gnd.n5771 gnd.n5769 9.3005
R10239 gnd.n5326 gnd.n5325 9.3005
R10240 gnd.n5826 gnd.n5825 9.3005
R10241 gnd.n5827 gnd.n5324 9.3005
R10242 gnd.n5831 gnd.n5828 9.3005
R10243 gnd.n5830 gnd.n5829 9.3005
R10244 gnd.n5299 gnd.n5298 9.3005
R10245 gnd.n5866 gnd.n5865 9.3005
R10246 gnd.n5867 gnd.n5297 9.3005
R10247 gnd.n5871 gnd.n5868 9.3005
R10248 gnd.n5870 gnd.n5869 9.3005
R10249 gnd.n5208 gnd.n5207 9.3005
R10250 gnd.n5911 gnd.n5910 9.3005
R10251 gnd.n5912 gnd.n5206 9.3005
R10252 gnd.n5916 gnd.n5913 9.3005
R10253 gnd.n5915 gnd.n5914 9.3005
R10254 gnd.n5180 gnd.n5179 9.3005
R10255 gnd.n5950 gnd.n5949 9.3005
R10256 gnd.n5951 gnd.n5178 9.3005
R10257 gnd.n5958 gnd.n5952 9.3005
R10258 gnd.n5957 gnd.n5953 9.3005
R10259 gnd.n5956 gnd.n5954 9.3005
R10260 gnd.n5150 gnd.n5149 9.3005
R10261 gnd.n6007 gnd.n6006 9.3005
R10262 gnd.n6008 gnd.n5148 9.3005
R10263 gnd.n6016 gnd.n6009 9.3005
R10264 gnd.n6015 gnd.n6010 9.3005
R10265 gnd.n6014 gnd.n6012 9.3005
R10266 gnd.n6011 gnd.n984 9.3005
R10267 gnd.n6453 gnd.n985 9.3005
R10268 gnd.n6452 gnd.n986 9.3005
R10269 gnd.n6451 gnd.n987 9.3005
R10270 gnd.n1009 gnd.n988 9.3005
R10271 gnd.n1010 gnd.n1008 9.3005
R10272 gnd.n6439 gnd.n1011 9.3005
R10273 gnd.n6438 gnd.n1012 9.3005
R10274 gnd.n6437 gnd.n1013 9.3005
R10275 gnd.n5051 gnd.n1014 9.3005
R10276 gnd.n5052 gnd.n5050 9.3005
R10277 gnd.n6425 gnd.n6424 9.3005
R10278 gnd.n5406 gnd.n5405 9.3005
R10279 gnd.n5646 gnd.n5645 9.3005
R10280 gnd.n5649 gnd.n5641 9.3005
R10281 gnd.n5650 gnd.n5640 9.3005
R10282 gnd.n5653 gnd.n5639 9.3005
R10283 gnd.n5654 gnd.n5638 9.3005
R10284 gnd.n5657 gnd.n5637 9.3005
R10285 gnd.n5658 gnd.n5636 9.3005
R10286 gnd.n5661 gnd.n5635 9.3005
R10287 gnd.n5662 gnd.n5634 9.3005
R10288 gnd.n5665 gnd.n5633 9.3005
R10289 gnd.n5666 gnd.n5632 9.3005
R10290 gnd.n5669 gnd.n5631 9.3005
R10291 gnd.n5671 gnd.n5630 9.3005
R10292 gnd.n5672 gnd.n5629 9.3005
R10293 gnd.n5673 gnd.n5628 9.3005
R10294 gnd.n5674 gnd.n5627 9.3005
R10295 gnd.n5642 gnd.n5423 9.3005
R10296 gnd.n5691 gnd.n5414 9.3005
R10297 gnd.n5693 gnd.n5692 9.3005
R10298 gnd.n5401 gnd.n5396 9.3005
R10299 gnd.n5714 gnd.n5395 9.3005
R10300 gnd.n5717 gnd.n5716 9.3005
R10301 gnd.n5719 gnd.n5718 9.3005
R10302 gnd.n5722 gnd.n5378 9.3005
R10303 gnd.n5720 gnd.n5376 9.3005
R10304 gnd.n5742 gnd.n5374 9.3005
R10305 gnd.n5746 gnd.n5745 9.3005
R10306 gnd.n5744 gnd.n5349 9.3005
R10307 gnd.n5780 gnd.n5348 9.3005
R10308 gnd.n5783 gnd.n5782 9.3005
R10309 gnd.n5346 gnd.n5345 9.3005
R10310 gnd.n5789 gnd.n5343 9.3005
R10311 gnd.n5791 gnd.n5790 9.3005
R10312 gnd.n5317 gnd.n5316 9.3005
R10313 gnd.n5840 gnd.n5839 9.3005
R10314 gnd.n5841 gnd.n5310 9.3005
R10315 gnd.n5849 gnd.n5309 9.3005
R10316 gnd.n5852 gnd.n5851 9.3005
R10317 gnd.n5854 gnd.n5853 9.3005
R10318 gnd.n5857 gnd.n5292 9.3005
R10319 gnd.n5855 gnd.n5290 9.3005
R10320 gnd.n5877 gnd.n5288 9.3005
R10321 gnd.n5879 gnd.n5878 9.3005
R10322 gnd.n5198 gnd.n5197 9.3005
R10323 gnd.n5925 gnd.n5924 9.3005
R10324 gnd.n5926 gnd.n5191 9.3005
R10325 gnd.n5934 gnd.n5190 9.3005
R10326 gnd.n5937 gnd.n5936 9.3005
R10327 gnd.n5939 gnd.n5938 9.3005
R10328 gnd.n5941 gnd.n5173 9.3005
R10329 gnd.n5171 gnd.n5169 9.3005
R10330 gnd.n5966 gnd.n5965 9.3005
R10331 gnd.n5155 gnd.n5154 9.3005
R10332 gnd.n5999 gnd.n5998 9.3005
R10333 gnd.n6000 gnd.n5141 9.3005
R10334 gnd.n6023 gnd.n5140 9.3005
R10335 gnd.n6026 gnd.n6025 9.3005
R10336 gnd.n5137 gnd.n5136 9.3005
R10337 gnd.n6030 gnd.n5138 9.3005
R10338 gnd.n6032 gnd.n6031 9.3005
R10339 gnd.n6317 gnd.n6034 9.3005
R10340 gnd.n6316 gnd.n6036 9.3005
R10341 gnd.n6315 gnd.n6037 9.3005
R10342 gnd.n6312 gnd.n6038 9.3005
R10343 gnd.n6311 gnd.n6039 9.3005
R10344 gnd.n6310 gnd.n6297 9.3005
R10345 gnd.n6307 gnd.n6299 9.3005
R10346 gnd.n6306 gnd.n6300 9.3005
R10347 gnd.n6303 gnd.n6301 9.3005
R10348 gnd.n6302 gnd.n5082 9.3005
R10349 gnd.n5690 gnd.n5417 9.3005
R10350 gnd.n6389 gnd.n5083 9.3005
R10351 gnd.n6388 gnd.n5085 9.3005
R10352 gnd.n5089 gnd.n5086 9.3005
R10353 gnd.n6383 gnd.n5090 9.3005
R10354 gnd.n6382 gnd.n5091 9.3005
R10355 gnd.n6381 gnd.n5092 9.3005
R10356 gnd.n5096 gnd.n5093 9.3005
R10357 gnd.n6376 gnd.n5097 9.3005
R10358 gnd.n6375 gnd.n5098 9.3005
R10359 gnd.n6374 gnd.n5099 9.3005
R10360 gnd.n5103 gnd.n5100 9.3005
R10361 gnd.n6369 gnd.n5104 9.3005
R10362 gnd.n6368 gnd.n5105 9.3005
R10363 gnd.n6367 gnd.n5106 9.3005
R10364 gnd.n5110 gnd.n5107 9.3005
R10365 gnd.n6362 gnd.n5111 9.3005
R10366 gnd.n6361 gnd.n5112 9.3005
R10367 gnd.n6360 gnd.n5113 9.3005
R10368 gnd.n5117 gnd.n5114 9.3005
R10369 gnd.n6355 gnd.n5118 9.3005
R10370 gnd.n6354 gnd.n5119 9.3005
R10371 gnd.n6353 gnd.n5120 9.3005
R10372 gnd.n5127 gnd.n5125 9.3005
R10373 gnd.n6348 gnd.n5128 9.3005
R10374 gnd.n6347 gnd.n5129 9.3005
R10375 gnd.n6346 gnd.n6343 9.3005
R10376 gnd.n6391 gnd.n6390 9.3005
R10377 gnd.n5887 gnd.n5886 9.3005
R10378 gnd.n5888 gnd.n5214 9.3005
R10379 gnd.n5905 gnd.n5889 9.3005
R10380 gnd.n5904 gnd.n5890 9.3005
R10381 gnd.n5903 gnd.n5891 9.3005
R10382 gnd.n5901 gnd.n5892 9.3005
R10383 gnd.n5900 gnd.n5893 9.3005
R10384 gnd.n5898 gnd.n5894 9.3005
R10385 gnd.n5897 gnd.n5895 9.3005
R10386 gnd.n5162 gnd.n5161 9.3005
R10387 gnd.n5973 gnd.n5972 9.3005
R10388 gnd.n5974 gnd.n5160 9.3005
R10389 gnd.n5991 gnd.n5975 9.3005
R10390 gnd.n5990 gnd.n5976 9.3005
R10391 gnd.n5989 gnd.n5977 9.3005
R10392 gnd.n5988 gnd.n5978 9.3005
R10393 gnd.n5986 gnd.n5979 9.3005
R10394 gnd.n5985 gnd.n5980 9.3005
R10395 gnd.n5982 gnd.n5981 9.3005
R10396 gnd.n5135 gnd.n5134 9.3005
R10397 gnd.n6324 gnd.n6323 9.3005
R10398 gnd.n6325 gnd.n5133 9.3005
R10399 gnd.n6329 gnd.n6326 9.3005
R10400 gnd.n6330 gnd.n5132 9.3005
R10401 gnd.n6334 gnd.n6333 9.3005
R10402 gnd.n6335 gnd.n5131 9.3005
R10403 gnd.n6337 gnd.n6336 9.3005
R10404 gnd.n6340 gnd.n5130 9.3005
R10405 gnd.n6342 gnd.n6341 9.3005
R10406 gnd.n5560 gnd.n5454 9.3005
R10407 gnd.n5562 gnd.n5561 9.3005
R10408 gnd.n5444 gnd.n5443 9.3005
R10409 gnd.n5575 gnd.n5574 9.3005
R10410 gnd.n5576 gnd.n5442 9.3005
R10411 gnd.n5578 gnd.n5577 9.3005
R10412 gnd.n5431 gnd.n5430 9.3005
R10413 gnd.n5591 gnd.n5590 9.3005
R10414 gnd.n5592 gnd.n5429 9.3005
R10415 gnd.n5616 gnd.n5593 9.3005
R10416 gnd.n5615 gnd.n5594 9.3005
R10417 gnd.n5614 gnd.n5595 9.3005
R10418 gnd.n5613 gnd.n5596 9.3005
R10419 gnd.n5611 gnd.n5597 9.3005
R10420 gnd.n5610 gnd.n5598 9.3005
R10421 gnd.n5608 gnd.n5599 9.3005
R10422 gnd.n5607 gnd.n5600 9.3005
R10423 gnd.n5605 gnd.n5601 9.3005
R10424 gnd.n5604 gnd.n5602 9.3005
R10425 gnd.n5366 gnd.n5365 9.3005
R10426 gnd.n5754 gnd.n5753 9.3005
R10427 gnd.n5755 gnd.n5364 9.3005
R10428 gnd.n5759 gnd.n5756 9.3005
R10429 gnd.n5758 gnd.n5757 9.3005
R10430 gnd.n5333 gnd.n5332 9.3005
R10431 gnd.n5801 gnd.n5800 9.3005
R10432 gnd.n5802 gnd.n5331 9.3005
R10433 gnd.n5804 gnd.n5803 9.3005
R10434 gnd.n5559 gnd.n5558 9.3005
R10435 gnd.n5499 gnd.n5498 9.3005
R10436 gnd.n5504 gnd.n5496 9.3005
R10437 gnd.n5505 gnd.n5495 9.3005
R10438 gnd.n5507 gnd.n5492 9.3005
R10439 gnd.n5491 gnd.n5489 9.3005
R10440 gnd.n5513 gnd.n5488 9.3005
R10441 gnd.n5514 gnd.n5487 9.3005
R10442 gnd.n5515 gnd.n5486 9.3005
R10443 gnd.n5485 gnd.n5483 9.3005
R10444 gnd.n5521 gnd.n5482 9.3005
R10445 gnd.n5522 gnd.n5481 9.3005
R10446 gnd.n5523 gnd.n5480 9.3005
R10447 gnd.n5479 gnd.n5477 9.3005
R10448 gnd.n5529 gnd.n5476 9.3005
R10449 gnd.n5530 gnd.n5475 9.3005
R10450 gnd.n5531 gnd.n5474 9.3005
R10451 gnd.n5473 gnd.n5471 9.3005
R10452 gnd.n5537 gnd.n5470 9.3005
R10453 gnd.n5538 gnd.n5469 9.3005
R10454 gnd.n5539 gnd.n5468 9.3005
R10455 gnd.n5467 gnd.n5465 9.3005
R10456 gnd.n5544 gnd.n5464 9.3005
R10457 gnd.n5545 gnd.n5463 9.3005
R10458 gnd.n5462 gnd.n5460 9.3005
R10459 gnd.n5550 gnd.n5459 9.3005
R10460 gnd.n5552 gnd.n5551 9.3005
R10461 gnd.n5497 gnd.n5455 9.3005
R10462 gnd.n5450 gnd.n5449 9.3005
R10463 gnd.n5567 gnd.n5566 9.3005
R10464 gnd.n5568 gnd.n5448 9.3005
R10465 gnd.n5570 gnd.n5569 9.3005
R10466 gnd.n5438 gnd.n5437 9.3005
R10467 gnd.n5583 gnd.n5582 9.3005
R10468 gnd.n5584 gnd.n5436 9.3005
R10469 gnd.n5586 gnd.n5585 9.3005
R10470 gnd.n5425 gnd.n5424 9.3005
R10471 gnd.n5681 gnd.n5680 9.3005
R10472 gnd.n5683 gnd.n5422 9.3005
R10473 gnd.n5685 gnd.n5684 9.3005
R10474 gnd.n5416 gnd.n5413 9.3005
R10475 gnd.n5695 gnd.n5694 9.3005
R10476 gnd.n5415 gnd.n5397 9.3005
R10477 gnd.n5713 gnd.n5712 9.3005
R10478 gnd.n5715 gnd.n5393 9.3005
R10479 gnd.n5725 gnd.n5394 9.3005
R10480 gnd.n5724 gnd.n5723 9.3005
R10481 gnd.n5721 gnd.n5372 9.3005
R10482 gnd.n5749 gnd.n5373 9.3005
R10483 gnd.n5748 gnd.n5747 9.3005
R10484 gnd.n5375 gnd.n5350 9.3005
R10485 gnd.n5779 gnd.n5778 9.3005
R10486 gnd.n5781 gnd.n5340 9.3005
R10487 gnd.n5796 gnd.n5341 9.3005
R10488 gnd.n5795 gnd.n5342 9.3005
R10489 gnd.n5794 gnd.n5792 9.3005
R10490 gnd.n5344 gnd.n5318 9.3005
R10491 gnd.n5837 gnd.n5836 9.3005
R10492 gnd.n5838 gnd.n5311 9.3005
R10493 gnd.n5848 gnd.n5847 9.3005
R10494 gnd.n5850 gnd.n5307 9.3005
R10495 gnd.n5860 gnd.n5308 9.3005
R10496 gnd.n5859 gnd.n5858 9.3005
R10497 gnd.n5856 gnd.n5286 9.3005
R10498 gnd.n5882 gnd.n5287 9.3005
R10499 gnd.n5881 gnd.n5880 9.3005
R10500 gnd.n5289 gnd.n5199 9.3005
R10501 gnd.n5922 gnd.n5921 9.3005
R10502 gnd.n5923 gnd.n5192 9.3005
R10503 gnd.n5933 gnd.n5932 9.3005
R10504 gnd.n5935 gnd.n5188 9.3005
R10505 gnd.n5944 gnd.n5189 9.3005
R10506 gnd.n5943 gnd.n5942 9.3005
R10507 gnd.n5940 gnd.n5168 9.3005
R10508 gnd.n5968 gnd.n5967 9.3005
R10509 gnd.n5170 gnd.n5156 9.3005
R10510 gnd.n5996 gnd.n5995 9.3005
R10511 gnd.n5997 gnd.n5142 9.3005
R10512 gnd.n6022 gnd.n6021 9.3005
R10513 gnd.n6024 gnd.n973 9.3005
R10514 gnd.n6460 gnd.n974 9.3005
R10515 gnd.n6459 gnd.n975 9.3005
R10516 gnd.n6458 gnd.n976 9.3005
R10517 gnd.n6033 gnd.n977 9.3005
R10518 gnd.n6035 gnd.n996 9.3005
R10519 gnd.n6446 gnd.n997 9.3005
R10520 gnd.n6445 gnd.n998 9.3005
R10521 gnd.n6444 gnd.n999 9.3005
R10522 gnd.n6296 gnd.n1000 9.3005
R10523 gnd.n6298 gnd.n1022 9.3005
R10524 gnd.n6432 gnd.n1023 9.3005
R10525 gnd.n6431 gnd.n1024 9.3005
R10526 gnd.n6430 gnd.n1025 9.3005
R10527 gnd.n5554 gnd.n5553 9.3005
R10528 gnd.n799 gnd.n798 9.3005
R10529 gnd.n6636 gnd.n6635 9.3005
R10530 gnd.n6637 gnd.n797 9.3005
R10531 gnd.n6639 gnd.n6638 9.3005
R10532 gnd.n793 gnd.n792 9.3005
R10533 gnd.n6646 gnd.n6645 9.3005
R10534 gnd.n6647 gnd.n791 9.3005
R10535 gnd.n6649 gnd.n6648 9.3005
R10536 gnd.n787 gnd.n786 9.3005
R10537 gnd.n6656 gnd.n6655 9.3005
R10538 gnd.n6657 gnd.n785 9.3005
R10539 gnd.n6659 gnd.n6658 9.3005
R10540 gnd.n781 gnd.n780 9.3005
R10541 gnd.n6666 gnd.n6665 9.3005
R10542 gnd.n6667 gnd.n779 9.3005
R10543 gnd.n6669 gnd.n6668 9.3005
R10544 gnd.n775 gnd.n774 9.3005
R10545 gnd.n6676 gnd.n6675 9.3005
R10546 gnd.n6677 gnd.n773 9.3005
R10547 gnd.n6679 gnd.n6678 9.3005
R10548 gnd.n769 gnd.n768 9.3005
R10549 gnd.n6686 gnd.n6685 9.3005
R10550 gnd.n6687 gnd.n767 9.3005
R10551 gnd.n6689 gnd.n6688 9.3005
R10552 gnd.n763 gnd.n762 9.3005
R10553 gnd.n6696 gnd.n6695 9.3005
R10554 gnd.n6697 gnd.n761 9.3005
R10555 gnd.n6699 gnd.n6698 9.3005
R10556 gnd.n757 gnd.n756 9.3005
R10557 gnd.n6706 gnd.n6705 9.3005
R10558 gnd.n6707 gnd.n755 9.3005
R10559 gnd.n6709 gnd.n6708 9.3005
R10560 gnd.n751 gnd.n750 9.3005
R10561 gnd.n6716 gnd.n6715 9.3005
R10562 gnd.n6717 gnd.n749 9.3005
R10563 gnd.n6719 gnd.n6718 9.3005
R10564 gnd.n745 gnd.n744 9.3005
R10565 gnd.n6726 gnd.n6725 9.3005
R10566 gnd.n6727 gnd.n743 9.3005
R10567 gnd.n6729 gnd.n6728 9.3005
R10568 gnd.n739 gnd.n738 9.3005
R10569 gnd.n6736 gnd.n6735 9.3005
R10570 gnd.n6737 gnd.n737 9.3005
R10571 gnd.n6739 gnd.n6738 9.3005
R10572 gnd.n733 gnd.n732 9.3005
R10573 gnd.n6746 gnd.n6745 9.3005
R10574 gnd.n6747 gnd.n731 9.3005
R10575 gnd.n6749 gnd.n6748 9.3005
R10576 gnd.n727 gnd.n726 9.3005
R10577 gnd.n6756 gnd.n6755 9.3005
R10578 gnd.n6757 gnd.n725 9.3005
R10579 gnd.n6759 gnd.n6758 9.3005
R10580 gnd.n721 gnd.n720 9.3005
R10581 gnd.n6766 gnd.n6765 9.3005
R10582 gnd.n6767 gnd.n719 9.3005
R10583 gnd.n6769 gnd.n6768 9.3005
R10584 gnd.n715 gnd.n714 9.3005
R10585 gnd.n6776 gnd.n6775 9.3005
R10586 gnd.n6777 gnd.n713 9.3005
R10587 gnd.n6779 gnd.n6778 9.3005
R10588 gnd.n709 gnd.n708 9.3005
R10589 gnd.n6786 gnd.n6785 9.3005
R10590 gnd.n6787 gnd.n707 9.3005
R10591 gnd.n6789 gnd.n6788 9.3005
R10592 gnd.n703 gnd.n702 9.3005
R10593 gnd.n6796 gnd.n6795 9.3005
R10594 gnd.n6797 gnd.n701 9.3005
R10595 gnd.n6799 gnd.n6798 9.3005
R10596 gnd.n697 gnd.n696 9.3005
R10597 gnd.n6806 gnd.n6805 9.3005
R10598 gnd.n6807 gnd.n695 9.3005
R10599 gnd.n6809 gnd.n6808 9.3005
R10600 gnd.n691 gnd.n690 9.3005
R10601 gnd.n6816 gnd.n6815 9.3005
R10602 gnd.n6817 gnd.n689 9.3005
R10603 gnd.n6819 gnd.n6818 9.3005
R10604 gnd.n685 gnd.n684 9.3005
R10605 gnd.n6826 gnd.n6825 9.3005
R10606 gnd.n6827 gnd.n683 9.3005
R10607 gnd.n6829 gnd.n6828 9.3005
R10608 gnd.n679 gnd.n678 9.3005
R10609 gnd.n6836 gnd.n6835 9.3005
R10610 gnd.n6837 gnd.n677 9.3005
R10611 gnd.n6839 gnd.n6838 9.3005
R10612 gnd.n673 gnd.n672 9.3005
R10613 gnd.n6846 gnd.n6845 9.3005
R10614 gnd.n6847 gnd.n671 9.3005
R10615 gnd.n6849 gnd.n6848 9.3005
R10616 gnd.n667 gnd.n666 9.3005
R10617 gnd.n6856 gnd.n6855 9.3005
R10618 gnd.n6857 gnd.n665 9.3005
R10619 gnd.n6859 gnd.n6858 9.3005
R10620 gnd.n661 gnd.n660 9.3005
R10621 gnd.n6866 gnd.n6865 9.3005
R10622 gnd.n6867 gnd.n659 9.3005
R10623 gnd.n6869 gnd.n6868 9.3005
R10624 gnd.n655 gnd.n654 9.3005
R10625 gnd.n6876 gnd.n6875 9.3005
R10626 gnd.n6877 gnd.n653 9.3005
R10627 gnd.n6879 gnd.n6878 9.3005
R10628 gnd.n649 gnd.n648 9.3005
R10629 gnd.n6886 gnd.n6885 9.3005
R10630 gnd.n6887 gnd.n647 9.3005
R10631 gnd.n6889 gnd.n6888 9.3005
R10632 gnd.n643 gnd.n642 9.3005
R10633 gnd.n6896 gnd.n6895 9.3005
R10634 gnd.n6897 gnd.n641 9.3005
R10635 gnd.n6899 gnd.n6898 9.3005
R10636 gnd.n637 gnd.n636 9.3005
R10637 gnd.n6906 gnd.n6905 9.3005
R10638 gnd.n6907 gnd.n635 9.3005
R10639 gnd.n6909 gnd.n6908 9.3005
R10640 gnd.n631 gnd.n630 9.3005
R10641 gnd.n6916 gnd.n6915 9.3005
R10642 gnd.n6917 gnd.n629 9.3005
R10643 gnd.n6919 gnd.n6918 9.3005
R10644 gnd.n625 gnd.n624 9.3005
R10645 gnd.n6926 gnd.n6925 9.3005
R10646 gnd.n6927 gnd.n623 9.3005
R10647 gnd.n6929 gnd.n6928 9.3005
R10648 gnd.n619 gnd.n618 9.3005
R10649 gnd.n6936 gnd.n6935 9.3005
R10650 gnd.n6937 gnd.n617 9.3005
R10651 gnd.n6939 gnd.n6938 9.3005
R10652 gnd.n613 gnd.n612 9.3005
R10653 gnd.n6946 gnd.n6945 9.3005
R10654 gnd.n6947 gnd.n611 9.3005
R10655 gnd.n6949 gnd.n6948 9.3005
R10656 gnd.n607 gnd.n606 9.3005
R10657 gnd.n6956 gnd.n6955 9.3005
R10658 gnd.n6957 gnd.n605 9.3005
R10659 gnd.n6959 gnd.n6958 9.3005
R10660 gnd.n601 gnd.n600 9.3005
R10661 gnd.n6966 gnd.n6965 9.3005
R10662 gnd.n6967 gnd.n599 9.3005
R10663 gnd.n6969 gnd.n6968 9.3005
R10664 gnd.n595 gnd.n594 9.3005
R10665 gnd.n6976 gnd.n6975 9.3005
R10666 gnd.n6977 gnd.n593 9.3005
R10667 gnd.n6979 gnd.n6978 9.3005
R10668 gnd.n589 gnd.n588 9.3005
R10669 gnd.n6986 gnd.n6985 9.3005
R10670 gnd.n6987 gnd.n587 9.3005
R10671 gnd.n6989 gnd.n6988 9.3005
R10672 gnd.n583 gnd.n582 9.3005
R10673 gnd.n6996 gnd.n6995 9.3005
R10674 gnd.n6997 gnd.n581 9.3005
R10675 gnd.n6999 gnd.n6998 9.3005
R10676 gnd.n577 gnd.n576 9.3005
R10677 gnd.n7006 gnd.n7005 9.3005
R10678 gnd.n7007 gnd.n575 9.3005
R10679 gnd.n7009 gnd.n7008 9.3005
R10680 gnd.n571 gnd.n570 9.3005
R10681 gnd.n7016 gnd.n7015 9.3005
R10682 gnd.n7017 gnd.n569 9.3005
R10683 gnd.n7019 gnd.n7018 9.3005
R10684 gnd.n565 gnd.n564 9.3005
R10685 gnd.n7026 gnd.n7025 9.3005
R10686 gnd.n7027 gnd.n563 9.3005
R10687 gnd.n7029 gnd.n7028 9.3005
R10688 gnd.n559 gnd.n558 9.3005
R10689 gnd.n7036 gnd.n7035 9.3005
R10690 gnd.n7037 gnd.n557 9.3005
R10691 gnd.n7039 gnd.n7038 9.3005
R10692 gnd.n553 gnd.n552 9.3005
R10693 gnd.n7046 gnd.n7045 9.3005
R10694 gnd.n7047 gnd.n551 9.3005
R10695 gnd.n7049 gnd.n7048 9.3005
R10696 gnd.n547 gnd.n546 9.3005
R10697 gnd.n7056 gnd.n7055 9.3005
R10698 gnd.n7057 gnd.n545 9.3005
R10699 gnd.n7059 gnd.n7058 9.3005
R10700 gnd.n541 gnd.n540 9.3005
R10701 gnd.n7066 gnd.n7065 9.3005
R10702 gnd.n7067 gnd.n539 9.3005
R10703 gnd.n7069 gnd.n7068 9.3005
R10704 gnd.n535 gnd.n534 9.3005
R10705 gnd.n7076 gnd.n7075 9.3005
R10706 gnd.n7077 gnd.n533 9.3005
R10707 gnd.n7079 gnd.n7078 9.3005
R10708 gnd.n529 gnd.n528 9.3005
R10709 gnd.n7086 gnd.n7085 9.3005
R10710 gnd.n7089 gnd.n7088 9.3005
R10711 gnd.n523 gnd.n522 9.3005
R10712 gnd.n7096 gnd.n7095 9.3005
R10713 gnd.n7097 gnd.n521 9.3005
R10714 gnd.n7099 gnd.n7098 9.3005
R10715 gnd.n517 gnd.n516 9.3005
R10716 gnd.n7106 gnd.n7105 9.3005
R10717 gnd.n7107 gnd.n515 9.3005
R10718 gnd.n7109 gnd.n7108 9.3005
R10719 gnd.n511 gnd.n510 9.3005
R10720 gnd.n7116 gnd.n7115 9.3005
R10721 gnd.n7117 gnd.n509 9.3005
R10722 gnd.n7119 gnd.n7118 9.3005
R10723 gnd.n505 gnd.n504 9.3005
R10724 gnd.n7126 gnd.n7125 9.3005
R10725 gnd.n7127 gnd.n503 9.3005
R10726 gnd.n7129 gnd.n7128 9.3005
R10727 gnd.n499 gnd.n498 9.3005
R10728 gnd.n7136 gnd.n7135 9.3005
R10729 gnd.n7137 gnd.n497 9.3005
R10730 gnd.n7139 gnd.n7138 9.3005
R10731 gnd.n493 gnd.n492 9.3005
R10732 gnd.n7146 gnd.n7145 9.3005
R10733 gnd.n7147 gnd.n491 9.3005
R10734 gnd.n7149 gnd.n7148 9.3005
R10735 gnd.n487 gnd.n486 9.3005
R10736 gnd.n7156 gnd.n7155 9.3005
R10737 gnd.n7157 gnd.n485 9.3005
R10738 gnd.n7159 gnd.n7158 9.3005
R10739 gnd.n481 gnd.n480 9.3005
R10740 gnd.n7166 gnd.n7165 9.3005
R10741 gnd.n7167 gnd.n479 9.3005
R10742 gnd.n7169 gnd.n7168 9.3005
R10743 gnd.n475 gnd.n474 9.3005
R10744 gnd.n7176 gnd.n7175 9.3005
R10745 gnd.n7177 gnd.n473 9.3005
R10746 gnd.n7179 gnd.n7178 9.3005
R10747 gnd.n469 gnd.n468 9.3005
R10748 gnd.n7186 gnd.n7185 9.3005
R10749 gnd.n7187 gnd.n467 9.3005
R10750 gnd.n7189 gnd.n7188 9.3005
R10751 gnd.n463 gnd.n462 9.3005
R10752 gnd.n7196 gnd.n7195 9.3005
R10753 gnd.n7197 gnd.n461 9.3005
R10754 gnd.n7199 gnd.n7198 9.3005
R10755 gnd.n457 gnd.n456 9.3005
R10756 gnd.n7206 gnd.n7205 9.3005
R10757 gnd.n7207 gnd.n455 9.3005
R10758 gnd.n7209 gnd.n7208 9.3005
R10759 gnd.n451 gnd.n450 9.3005
R10760 gnd.n7216 gnd.n7215 9.3005
R10761 gnd.n7217 gnd.n449 9.3005
R10762 gnd.n7219 gnd.n7218 9.3005
R10763 gnd.n445 gnd.n444 9.3005
R10764 gnd.n7226 gnd.n7225 9.3005
R10765 gnd.n7227 gnd.n443 9.3005
R10766 gnd.n7229 gnd.n7228 9.3005
R10767 gnd.n439 gnd.n438 9.3005
R10768 gnd.n7236 gnd.n7235 9.3005
R10769 gnd.n7237 gnd.n437 9.3005
R10770 gnd.n7239 gnd.n7238 9.3005
R10771 gnd.n433 gnd.n432 9.3005
R10772 gnd.n7246 gnd.n7245 9.3005
R10773 gnd.n7247 gnd.n431 9.3005
R10774 gnd.n7249 gnd.n7248 9.3005
R10775 gnd.n427 gnd.n426 9.3005
R10776 gnd.n7256 gnd.n7255 9.3005
R10777 gnd.n7257 gnd.n425 9.3005
R10778 gnd.n7259 gnd.n7258 9.3005
R10779 gnd.n421 gnd.n420 9.3005
R10780 gnd.n7266 gnd.n7265 9.3005
R10781 gnd.n7267 gnd.n419 9.3005
R10782 gnd.n7269 gnd.n7268 9.3005
R10783 gnd.n415 gnd.n414 9.3005
R10784 gnd.n7276 gnd.n7275 9.3005
R10785 gnd.n7277 gnd.n413 9.3005
R10786 gnd.n7279 gnd.n7278 9.3005
R10787 gnd.n409 gnd.n408 9.3005
R10788 gnd.n7286 gnd.n7285 9.3005
R10789 gnd.n7287 gnd.n407 9.3005
R10790 gnd.n7291 gnd.n7288 9.3005
R10791 gnd.n7290 gnd.n7289 9.3005
R10792 gnd.n403 gnd.n402 9.3005
R10793 gnd.n7299 gnd.n7298 9.3005
R10794 gnd.n7087 gnd.n527 9.3005
R10795 gnd.n7635 gnd.n7634 9.3005
R10796 gnd.n7633 gnd.n80 9.3005
R10797 gnd.n7324 gnd.n83 9.3005
R10798 gnd.n7326 gnd.n7325 9.3005
R10799 gnd.n377 gnd.n376 9.3005
R10800 gnd.n7337 gnd.n7336 9.3005
R10801 gnd.n7338 gnd.n375 9.3005
R10802 gnd.n7340 gnd.n7339 9.3005
R10803 gnd.n370 gnd.n369 9.3005
R10804 gnd.n7351 gnd.n7350 9.3005
R10805 gnd.n7352 gnd.n368 9.3005
R10806 gnd.n7354 gnd.n7353 9.3005
R10807 gnd.n365 gnd.n364 9.3005
R10808 gnd.n7365 gnd.n7364 9.3005
R10809 gnd.n7366 gnd.n363 9.3005
R10810 gnd.n7369 gnd.n7368 9.3005
R10811 gnd.n7367 gnd.n359 9.3005
R10812 gnd.n7394 gnd.n358 9.3005
R10813 gnd.n7396 gnd.n7395 9.3005
R10814 gnd.n7397 gnd.n357 9.3005
R10815 gnd.n7399 gnd.n7398 9.3005
R10816 gnd.n7401 gnd.n355 9.3005
R10817 gnd.n7403 gnd.n7402 9.3005
R10818 gnd.n7404 gnd.n354 9.3005
R10819 gnd.n7406 gnd.n7405 9.3005
R10820 gnd.n7408 gnd.n352 9.3005
R10821 gnd.n7410 gnd.n7409 9.3005
R10822 gnd.n7441 gnd.n318 9.3005
R10823 gnd.n7440 gnd.n320 9.3005
R10824 gnd.n324 gnd.n321 9.3005
R10825 gnd.n7435 gnd.n325 9.3005
R10826 gnd.n7434 gnd.n326 9.3005
R10827 gnd.n7433 gnd.n327 9.3005
R10828 gnd.n331 gnd.n328 9.3005
R10829 gnd.n7428 gnd.n332 9.3005
R10830 gnd.n7427 gnd.n333 9.3005
R10831 gnd.n7426 gnd.n334 9.3005
R10832 gnd.n338 gnd.n335 9.3005
R10833 gnd.n7421 gnd.n339 9.3005
R10834 gnd.n7420 gnd.n340 9.3005
R10835 gnd.n7419 gnd.n341 9.3005
R10836 gnd.n345 gnd.n342 9.3005
R10837 gnd.n7414 gnd.n346 9.3005
R10838 gnd.n7413 gnd.n7412 9.3005
R10839 gnd.n7411 gnd.n349 9.3005
R10840 gnd.n7443 gnd.n7442 9.3005
R10841 gnd.n7551 gnd.n215 9.3005
R10842 gnd.n7550 gnd.n217 9.3005
R10843 gnd.n221 gnd.n218 9.3005
R10844 gnd.n7545 gnd.n222 9.3005
R10845 gnd.n7544 gnd.n223 9.3005
R10846 gnd.n7543 gnd.n224 9.3005
R10847 gnd.n228 gnd.n225 9.3005
R10848 gnd.n7538 gnd.n229 9.3005
R10849 gnd.n7537 gnd.n230 9.3005
R10850 gnd.n7536 gnd.n231 9.3005
R10851 gnd.n235 gnd.n232 9.3005
R10852 gnd.n7531 gnd.n236 9.3005
R10853 gnd.n7530 gnd.n237 9.3005
R10854 gnd.n7529 gnd.n238 9.3005
R10855 gnd.n242 gnd.n239 9.3005
R10856 gnd.n7524 gnd.n243 9.3005
R10857 gnd.n7523 gnd.n244 9.3005
R10858 gnd.n7519 gnd.n245 9.3005
R10859 gnd.n249 gnd.n246 9.3005
R10860 gnd.n7514 gnd.n250 9.3005
R10861 gnd.n7513 gnd.n251 9.3005
R10862 gnd.n7512 gnd.n252 9.3005
R10863 gnd.n256 gnd.n253 9.3005
R10864 gnd.n7507 gnd.n257 9.3005
R10865 gnd.n7506 gnd.n258 9.3005
R10866 gnd.n7505 gnd.n259 9.3005
R10867 gnd.n263 gnd.n260 9.3005
R10868 gnd.n7500 gnd.n264 9.3005
R10869 gnd.n7499 gnd.n265 9.3005
R10870 gnd.n7498 gnd.n266 9.3005
R10871 gnd.n270 gnd.n267 9.3005
R10872 gnd.n7493 gnd.n271 9.3005
R10873 gnd.n7492 gnd.n272 9.3005
R10874 gnd.n7491 gnd.n273 9.3005
R10875 gnd.n277 gnd.n274 9.3005
R10876 gnd.n7486 gnd.n278 9.3005
R10877 gnd.n7485 gnd.n7484 9.3005
R10878 gnd.n7483 gnd.n279 9.3005
R10879 gnd.n7482 gnd.n7481 9.3005
R10880 gnd.n283 gnd.n282 9.3005
R10881 gnd.n288 gnd.n286 9.3005
R10882 gnd.n7474 gnd.n289 9.3005
R10883 gnd.n7473 gnd.n290 9.3005
R10884 gnd.n7472 gnd.n291 9.3005
R10885 gnd.n295 gnd.n292 9.3005
R10886 gnd.n7467 gnd.n296 9.3005
R10887 gnd.n7466 gnd.n297 9.3005
R10888 gnd.n7465 gnd.n298 9.3005
R10889 gnd.n302 gnd.n299 9.3005
R10890 gnd.n7460 gnd.n303 9.3005
R10891 gnd.n7459 gnd.n304 9.3005
R10892 gnd.n7458 gnd.n305 9.3005
R10893 gnd.n309 gnd.n306 9.3005
R10894 gnd.n7453 gnd.n310 9.3005
R10895 gnd.n7452 gnd.n311 9.3005
R10896 gnd.n7451 gnd.n312 9.3005
R10897 gnd.n317 gnd.n315 9.3005
R10898 gnd.n7446 gnd.n7445 9.3005
R10899 gnd.n7553 gnd.n7552 9.3005
R10900 gnd.n4328 gnd.n1617 9.3005
R10901 gnd.n4538 gnd.n1618 9.3005
R10902 gnd.n4537 gnd.n1619 9.3005
R10903 gnd.n4536 gnd.n1620 9.3005
R10904 gnd.n1802 gnd.n1621 9.3005
R10905 gnd.n4526 gnd.n1638 9.3005
R10906 gnd.n4525 gnd.n1639 9.3005
R10907 gnd.n4524 gnd.n1640 9.3005
R10908 gnd.n1765 gnd.n1641 9.3005
R10909 gnd.n4514 gnd.n1659 9.3005
R10910 gnd.n4513 gnd.n1660 9.3005
R10911 gnd.n4512 gnd.n1661 9.3005
R10912 gnd.n4361 gnd.n1662 9.3005
R10913 gnd.n4502 gnd.n1678 9.3005
R10914 gnd.n4501 gnd.n1679 9.3005
R10915 gnd.n4500 gnd.n1680 9.3005
R10916 gnd.n4371 gnd.n1681 9.3005
R10917 gnd.n4490 gnd.n1699 9.3005
R10918 gnd.n4489 gnd.n1700 9.3005
R10919 gnd.n4488 gnd.n1701 9.3005
R10920 gnd.n4419 gnd.n1702 9.3005
R10921 gnd.n4478 gnd.n1716 9.3005
R10922 gnd.n4477 gnd.n1717 9.3005
R10923 gnd.n4476 gnd.n1718 9.3005
R10924 gnd.n4420 gnd.n1719 9.3005
R10925 gnd.n4425 gnd.n4421 9.3005
R10926 gnd.n4433 gnd.n4426 9.3005
R10927 gnd.n4432 gnd.n4428 9.3005
R10928 gnd.n4431 gnd.n4429 9.3005
R10929 gnd.n379 gnd.n108 9.3005
R10930 gnd.n7621 gnd.n109 9.3005
R10931 gnd.n7620 gnd.n110 9.3005
R10932 gnd.n7619 gnd.n111 9.3005
R10933 gnd.n373 gnd.n112 9.3005
R10934 gnd.n7609 gnd.n127 9.3005
R10935 gnd.n7608 gnd.n128 9.3005
R10936 gnd.n7607 gnd.n129 9.3005
R10937 gnd.n367 gnd.n130 9.3005
R10938 gnd.n7597 gnd.n148 9.3005
R10939 gnd.n7596 gnd.n149 9.3005
R10940 gnd.n7595 gnd.n150 9.3005
R10941 gnd.n361 gnd.n151 9.3005
R10942 gnd.n7585 gnd.n167 9.3005
R10943 gnd.n7584 gnd.n168 9.3005
R10944 gnd.n7583 gnd.n169 9.3005
R10945 gnd.n7375 gnd.n170 9.3005
R10946 gnd.n7573 gnd.n187 9.3005
R10947 gnd.n7572 gnd.n188 9.3005
R10948 gnd.n7571 gnd.n189 9.3005
R10949 gnd.n7376 gnd.n190 9.3005
R10950 gnd.n7561 gnd.n205 9.3005
R10951 gnd.n7560 gnd.n206 9.3005
R10952 gnd.n7559 gnd.n207 9.3005
R10953 gnd.n4327 gnd.n4326 9.3005
R10954 gnd.n4329 gnd.n4328 9.3005
R10955 gnd.n4330 gnd.n1618 9.3005
R10956 gnd.n4331 gnd.n1619 9.3005
R10957 gnd.n1801 gnd.n1620 9.3005
R10958 gnd.n4343 gnd.n1802 9.3005
R10959 gnd.n4344 gnd.n1638 9.3005
R10960 gnd.n4345 gnd.n1639 9.3005
R10961 gnd.n1764 gnd.n1640 9.3005
R10962 gnd.n4357 gnd.n1765 9.3005
R10963 gnd.n4358 gnd.n1659 9.3005
R10964 gnd.n4359 gnd.n1660 9.3005
R10965 gnd.n4360 gnd.n1661 9.3005
R10966 gnd.n4364 gnd.n4361 9.3005
R10967 gnd.n4365 gnd.n1678 9.3005
R10968 gnd.n4369 gnd.n1679 9.3005
R10969 gnd.n4370 gnd.n1680 9.3005
R10970 gnd.n4372 gnd.n4371 9.3005
R10971 gnd.n1742 gnd.n1699 9.3005
R10972 gnd.n4417 gnd.n1700 9.3005
R10973 gnd.n4418 gnd.n1701 9.3005
R10974 gnd.n4443 gnd.n4419 9.3005
R10975 gnd.n4442 gnd.n1716 9.3005
R10976 gnd.n4441 gnd.n1717 9.3005
R10977 gnd.n4440 gnd.n1718 9.3005
R10978 gnd.n4439 gnd.n4420 9.3005
R10979 gnd.n4438 gnd.n4421 9.3005
R10980 gnd.n4426 gnd.n4422 9.3005
R10981 gnd.n4428 gnd.n4427 9.3005
R10982 gnd.n4429 gnd.n378 9.3005
R10983 gnd.n7330 gnd.n379 9.3005
R10984 gnd.n7331 gnd.n109 9.3005
R10985 gnd.n7332 gnd.n110 9.3005
R10986 gnd.n372 gnd.n111 9.3005
R10987 gnd.n7344 gnd.n373 9.3005
R10988 gnd.n7345 gnd.n127 9.3005
R10989 gnd.n7346 gnd.n128 9.3005
R10990 gnd.n366 gnd.n129 9.3005
R10991 gnd.n7358 gnd.n367 9.3005
R10992 gnd.n7359 gnd.n148 9.3005
R10993 gnd.n7360 gnd.n149 9.3005
R10994 gnd.n360 gnd.n150 9.3005
R10995 gnd.n7373 gnd.n361 9.3005
R10996 gnd.n7374 gnd.n167 9.3005
R10997 gnd.n7390 gnd.n168 9.3005
R10998 gnd.n7389 gnd.n169 9.3005
R10999 gnd.n7388 gnd.n7375 9.3005
R11000 gnd.n7386 gnd.n187 9.3005
R11001 gnd.n7385 gnd.n188 9.3005
R11002 gnd.n7383 gnd.n189 9.3005
R11003 gnd.n7382 gnd.n7376 9.3005
R11004 gnd.n7380 gnd.n205 9.3005
R11005 gnd.n7379 gnd.n206 9.3005
R11006 gnd.n7377 gnd.n207 9.3005
R11007 gnd.n4327 gnd.n1806 9.3005
R11008 gnd.n1812 gnd.n1809 9.3005
R11009 gnd.n4314 gnd.n1813 9.3005
R11010 gnd.n4316 gnd.n4315 9.3005
R11011 gnd.n4313 gnd.n1815 9.3005
R11012 gnd.n4312 gnd.n4311 9.3005
R11013 gnd.n1817 gnd.n1816 9.3005
R11014 gnd.n4305 gnd.n4304 9.3005
R11015 gnd.n4303 gnd.n1819 9.3005
R11016 gnd.n4302 gnd.n4301 9.3005
R11017 gnd.n1821 gnd.n1820 9.3005
R11018 gnd.n4295 gnd.n4294 9.3005
R11019 gnd.n4293 gnd.n1823 9.3005
R11020 gnd.n4292 gnd.n4291 9.3005
R11021 gnd.n1825 gnd.n1824 9.3005
R11022 gnd.n4285 gnd.n4284 9.3005
R11023 gnd.n4283 gnd.n1827 9.3005
R11024 gnd.n4282 gnd.n4281 9.3005
R11025 gnd.n1829 gnd.n1828 9.3005
R11026 gnd.n4275 gnd.n4274 9.3005
R11027 gnd.n4273 gnd.n1831 9.3005
R11028 gnd.n1833 gnd.n1832 9.3005
R11029 gnd.n4263 gnd.n4262 9.3005
R11030 gnd.n4261 gnd.n1835 9.3005
R11031 gnd.n4260 gnd.n4259 9.3005
R11032 gnd.n1837 gnd.n1836 9.3005
R11033 gnd.n4253 gnd.n4252 9.3005
R11034 gnd.n4251 gnd.n1839 9.3005
R11035 gnd.n4250 gnd.n4249 9.3005
R11036 gnd.n1841 gnd.n1840 9.3005
R11037 gnd.n4241 gnd.n4240 9.3005
R11038 gnd.n4238 gnd.n4151 9.3005
R11039 gnd.n4237 gnd.n4236 9.3005
R11040 gnd.n4153 gnd.n4152 9.3005
R11041 gnd.n4230 gnd.n4229 9.3005
R11042 gnd.n4228 gnd.n4155 9.3005
R11043 gnd.n4227 gnd.n4226 9.3005
R11044 gnd.n4157 gnd.n4156 9.3005
R11045 gnd.n4220 gnd.n4216 9.3005
R11046 gnd.n4215 gnd.n4159 9.3005
R11047 gnd.n4214 gnd.n4213 9.3005
R11048 gnd.n4161 gnd.n4160 9.3005
R11049 gnd.n4207 gnd.n4206 9.3005
R11050 gnd.n4205 gnd.n4163 9.3005
R11051 gnd.n4204 gnd.n4203 9.3005
R11052 gnd.n4165 gnd.n4164 9.3005
R11053 gnd.n4197 gnd.n4196 9.3005
R11054 gnd.n4195 gnd.n4167 9.3005
R11055 gnd.n4194 gnd.n4193 9.3005
R11056 gnd.n4169 gnd.n4168 9.3005
R11057 gnd.n4187 gnd.n4186 9.3005
R11058 gnd.n4185 gnd.n4171 9.3005
R11059 gnd.n4184 gnd.n4183 9.3005
R11060 gnd.n4173 gnd.n4172 9.3005
R11061 gnd.n4177 gnd.n4176 9.3005
R11062 gnd.n4175 gnd.n4174 9.3005
R11063 gnd.n4272 gnd.n4271 9.3005
R11064 gnd.n4324 gnd.n4323 9.3005
R11065 gnd.n4543 gnd.n1607 9.3005
R11066 gnd.n4542 gnd.n1608 9.3005
R11067 gnd.n1628 gnd.n1609 9.3005
R11068 gnd.n4532 gnd.n1629 9.3005
R11069 gnd.n4531 gnd.n1630 9.3005
R11070 gnd.n4530 gnd.n1631 9.3005
R11071 gnd.n1648 gnd.n1632 9.3005
R11072 gnd.n4520 gnd.n1649 9.3005
R11073 gnd.n4519 gnd.n1650 9.3005
R11074 gnd.n4518 gnd.n1651 9.3005
R11075 gnd.n1668 gnd.n1652 9.3005
R11076 gnd.n4508 gnd.n1669 9.3005
R11077 gnd.n4507 gnd.n1670 9.3005
R11078 gnd.n4506 gnd.n1671 9.3005
R11079 gnd.n1688 gnd.n1672 9.3005
R11080 gnd.n4496 gnd.n1689 9.3005
R11081 gnd.n4495 gnd.n1690 9.3005
R11082 gnd.n4494 gnd.n1691 9.3005
R11083 gnd.n1708 gnd.n1692 9.3005
R11084 gnd.n4484 gnd.n1709 9.3005
R11085 gnd.n4483 gnd.n94 9.3005
R11086 gnd.n99 gnd.n93 9.3005
R11087 gnd.n7615 gnd.n118 9.3005
R11088 gnd.n7614 gnd.n119 9.3005
R11089 gnd.n7613 gnd.n120 9.3005
R11090 gnd.n137 gnd.n121 9.3005
R11091 gnd.n7603 gnd.n138 9.3005
R11092 gnd.n7602 gnd.n139 9.3005
R11093 gnd.n7601 gnd.n140 9.3005
R11094 gnd.n157 gnd.n141 9.3005
R11095 gnd.n7591 gnd.n158 9.3005
R11096 gnd.n7590 gnd.n159 9.3005
R11097 gnd.n7589 gnd.n160 9.3005
R11098 gnd.n177 gnd.n161 9.3005
R11099 gnd.n7579 gnd.n178 9.3005
R11100 gnd.n7578 gnd.n179 9.3005
R11101 gnd.n7577 gnd.n180 9.3005
R11102 gnd.n196 gnd.n181 9.3005
R11103 gnd.n7567 gnd.n197 9.3005
R11104 gnd.n7566 gnd.n198 9.3005
R11105 gnd.n7565 gnd.n199 9.3005
R11106 gnd.n214 gnd.n200 9.3005
R11107 gnd.n7555 gnd.n7554 9.3005
R11108 gnd.n4544 gnd.n1606 9.3005
R11109 gnd.n7626 gnd.n97 9.3005
R11110 gnd.n7626 gnd.n7625 9.3005
R11111 gnd.n2945 gnd.n2944 9.3005
R11112 gnd.n2946 gnd.n2592 9.3005
R11113 gnd.n2948 gnd.n2947 9.3005
R11114 gnd.n2590 gnd.n2589 9.3005
R11115 gnd.n2953 gnd.n2952 9.3005
R11116 gnd.n2954 gnd.n2588 9.3005
R11117 gnd.n2976 gnd.n2955 9.3005
R11118 gnd.n2975 gnd.n2956 9.3005
R11119 gnd.n2974 gnd.n2957 9.3005
R11120 gnd.n2960 gnd.n2958 9.3005
R11121 gnd.n2970 gnd.n2961 9.3005
R11122 gnd.n2969 gnd.n2962 9.3005
R11123 gnd.n2968 gnd.n2963 9.3005
R11124 gnd.n2966 gnd.n2965 9.3005
R11125 gnd.n2964 gnd.n2566 9.3005
R11126 gnd.n2564 gnd.n2563 9.3005
R11127 gnd.n3042 gnd.n3041 9.3005
R11128 gnd.n3043 gnd.n2562 9.3005
R11129 gnd.n3045 gnd.n3044 9.3005
R11130 gnd.n2560 gnd.n2559 9.3005
R11131 gnd.n3050 gnd.n3049 9.3005
R11132 gnd.n3051 gnd.n2558 9.3005
R11133 gnd.n3053 gnd.n3052 9.3005
R11134 gnd.n2556 gnd.n2555 9.3005
R11135 gnd.n3061 gnd.n3060 9.3005
R11136 gnd.n3062 gnd.n2554 9.3005
R11137 gnd.n3066 gnd.n3063 9.3005
R11138 gnd.n3065 gnd.n3064 9.3005
R11139 gnd.n2325 gnd.n2324 9.3005
R11140 gnd.n3157 gnd.n3156 9.3005
R11141 gnd.n3158 gnd.n2323 9.3005
R11142 gnd.n3162 gnd.n3159 9.3005
R11143 gnd.n3161 gnd.n3160 9.3005
R11144 gnd.n2300 gnd.n2299 9.3005
R11145 gnd.n3187 gnd.n3186 9.3005
R11146 gnd.n3188 gnd.n2298 9.3005
R11147 gnd.n3192 gnd.n3189 9.3005
R11148 gnd.n3191 gnd.n3190 9.3005
R11149 gnd.n2275 gnd.n2274 9.3005
R11150 gnd.n3217 gnd.n3216 9.3005
R11151 gnd.n3218 gnd.n2273 9.3005
R11152 gnd.n3232 gnd.n3219 9.3005
R11153 gnd.n3231 gnd.n3220 9.3005
R11154 gnd.n3230 gnd.n3221 9.3005
R11155 gnd.n3223 gnd.n3222 9.3005
R11156 gnd.n3225 gnd.n3224 9.3005
R11157 gnd.n2181 gnd.n2180 9.3005
R11158 gnd.n3292 gnd.n3291 9.3005
R11159 gnd.n3293 gnd.n2179 9.3005
R11160 gnd.n3297 gnd.n3294 9.3005
R11161 gnd.n3296 gnd.n3295 9.3005
R11162 gnd.n2155 gnd.n2154 9.3005
R11163 gnd.n3354 gnd.n3353 9.3005
R11164 gnd.n3355 gnd.n2153 9.3005
R11165 gnd.n3357 gnd.n3356 9.3005
R11166 gnd.n2137 gnd.n2136 9.3005
R11167 gnd.n3381 gnd.n3380 9.3005
R11168 gnd.n3382 gnd.n2135 9.3005
R11169 gnd.n3386 gnd.n3383 9.3005
R11170 gnd.n3385 gnd.n3384 9.3005
R11171 gnd.n2104 gnd.n2103 9.3005
R11172 gnd.n3432 gnd.n3431 9.3005
R11173 gnd.n3433 gnd.n2102 9.3005
R11174 gnd.n3435 gnd.n3434 9.3005
R11175 gnd.n2081 gnd.n2080 9.3005
R11176 gnd.n3472 gnd.n3471 9.3005
R11177 gnd.n3473 gnd.n2079 9.3005
R11178 gnd.n3475 gnd.n3474 9.3005
R11179 gnd.n2059 gnd.n2058 9.3005
R11180 gnd.n3528 gnd.n3527 9.3005
R11181 gnd.n3529 gnd.n2057 9.3005
R11182 gnd.n3531 gnd.n3530 9.3005
R11183 gnd.n2040 gnd.n2039 9.3005
R11184 gnd.n3553 gnd.n3552 9.3005
R11185 gnd.n3554 gnd.n2038 9.3005
R11186 gnd.n3556 gnd.n3555 9.3005
R11187 gnd.n2020 gnd.n2019 9.3005
R11188 gnd.n3613 gnd.n3612 9.3005
R11189 gnd.n3614 gnd.n2018 9.3005
R11190 gnd.n3616 gnd.n3615 9.3005
R11191 gnd.n1998 gnd.n1997 9.3005
R11192 gnd.n3642 gnd.n3641 9.3005
R11193 gnd.n3643 gnd.n1996 9.3005
R11194 gnd.n3647 gnd.n3644 9.3005
R11195 gnd.n3646 gnd.n3645 9.3005
R11196 gnd.n1970 gnd.n1969 9.3005
R11197 gnd.n3687 gnd.n3686 9.3005
R11198 gnd.n3688 gnd.n1968 9.3005
R11199 gnd.n3696 gnd.n3689 9.3005
R11200 gnd.n3695 gnd.n3690 9.3005
R11201 gnd.n3694 gnd.n3692 9.3005
R11202 gnd.n3691 gnd.n1894 9.3005
R11203 gnd.n3983 gnd.n1895 9.3005
R11204 gnd.n3982 gnd.n1896 9.3005
R11205 gnd.n3981 gnd.n1897 9.3005
R11206 gnd.n1904 gnd.n1898 9.3005
R11207 gnd.n3972 gnd.n1905 9.3005
R11208 gnd.n3971 gnd.n1906 9.3005
R11209 gnd.n3970 gnd.n1907 9.3005
R11210 gnd.n1916 gnd.n1908 9.3005
R11211 gnd.n3961 gnd.n1917 9.3005
R11212 gnd.n3960 gnd.n1918 9.3005
R11213 gnd.n3959 gnd.n1919 9.3005
R11214 gnd.n1928 gnd.n1920 9.3005
R11215 gnd.n3950 gnd.n1929 9.3005
R11216 gnd.n3949 gnd.n1930 9.3005
R11217 gnd.n3948 gnd.n1931 9.3005
R11218 gnd.n3936 gnd.n1932 9.3005
R11219 gnd.n3939 gnd.n3938 9.3005
R11220 gnd.n3937 gnd.n1584 9.3005
R11221 gnd.n4559 gnd.n1585 9.3005
R11222 gnd.n4558 gnd.n1586 9.3005
R11223 gnd.n4557 gnd.n1587 9.3005
R11224 gnd.n1593 gnd.n1588 9.3005
R11225 gnd.n4551 gnd.n1594 9.3005
R11226 gnd.n4550 gnd.n1595 9.3005
R11227 gnd.n4549 gnd.n1596 9.3005
R11228 gnd.n1776 gnd.n1597 9.3005
R11229 gnd.n1777 gnd.n1775 9.3005
R11230 gnd.n1779 gnd.n1778 9.3005
R11231 gnd.n1773 gnd.n1772 9.3005
R11232 gnd.n1784 gnd.n1783 9.3005
R11233 gnd.n1785 gnd.n1771 9.3005
R11234 gnd.n1798 gnd.n1786 9.3005
R11235 gnd.n1797 gnd.n1787 9.3005
R11236 gnd.n1796 gnd.n1788 9.3005
R11237 gnd.n1793 gnd.n1789 9.3005
R11238 gnd.n1792 gnd.n1791 9.3005
R11239 gnd.n1790 gnd.n1754 9.3005
R11240 gnd.n1752 gnd.n1751 9.3005
R11241 gnd.n4397 gnd.n4396 9.3005
R11242 gnd.n4398 gnd.n1750 9.3005
R11243 gnd.n4400 gnd.n4399 9.3005
R11244 gnd.n1748 gnd.n1747 9.3005
R11245 gnd.n4405 gnd.n4404 9.3005
R11246 gnd.n4406 gnd.n1746 9.3005
R11247 gnd.n4412 gnd.n4407 9.3005
R11248 gnd.n4411 gnd.n4408 9.3005
R11249 gnd.n7318 gnd.n385 9.3005
R11250 gnd.n388 gnd.n386 9.3005
R11251 gnd.n7314 gnd.n389 9.3005
R11252 gnd.n7313 gnd.n390 9.3005
R11253 gnd.n7312 gnd.n391 9.3005
R11254 gnd.n394 gnd.n392 9.3005
R11255 gnd.n7308 gnd.n395 9.3005
R11256 gnd.n7307 gnd.n396 9.3005
R11257 gnd.n7306 gnd.n397 9.3005
R11258 gnd.n400 gnd.n398 9.3005
R11259 gnd.n7302 gnd.n401 9.3005
R11260 gnd.n7301 gnd.n7300 9.3005
R11261 gnd.n2746 gnd.n2684 9.3005
R11262 gnd.n2749 gnd.n2747 9.3005
R11263 gnd.n2750 gnd.n2683 9.3005
R11264 gnd.n2753 gnd.n2752 9.3005
R11265 gnd.n2754 gnd.n2682 9.3005
R11266 gnd.n2757 gnd.n2755 9.3005
R11267 gnd.n2758 gnd.n2681 9.3005
R11268 gnd.n2761 gnd.n2760 9.3005
R11269 gnd.n2762 gnd.n2680 9.3005
R11270 gnd.n2764 gnd.n2763 9.3005
R11271 gnd.n2665 gnd.n2664 9.3005
R11272 gnd.n2775 gnd.n2774 9.3005
R11273 gnd.n2776 gnd.n2663 9.3005
R11274 gnd.n2778 gnd.n2777 9.3005
R11275 gnd.n2660 gnd.n2659 9.3005
R11276 gnd.n2828 gnd.n2827 9.3005
R11277 gnd.n2829 gnd.n2658 9.3005
R11278 gnd.n2832 gnd.n2831 9.3005
R11279 gnd.n2830 gnd.n2654 9.3005
R11280 gnd.n2843 gnd.n2655 9.3005
R11281 gnd.n2844 gnd.n2653 9.3005
R11282 gnd.n2847 gnd.n2846 9.3005
R11283 gnd.n2848 gnd.n2652 9.3005
R11284 gnd.n2850 gnd.n2849 9.3005
R11285 gnd.n2618 gnd.n2617 9.3005
R11286 gnd.n2892 gnd.n2891 9.3005
R11287 gnd.n2745 gnd.n2744 9.3005
R11288 gnd.n2739 gnd.n2738 9.3005
R11289 gnd.n2737 gnd.n2689 9.3005
R11290 gnd.n2736 gnd.n2735 9.3005
R11291 gnd.n2732 gnd.n2692 9.3005
R11292 gnd.n2731 gnd.n2728 9.3005
R11293 gnd.n2727 gnd.n2693 9.3005
R11294 gnd.n2726 gnd.n2725 9.3005
R11295 gnd.n2722 gnd.n2694 9.3005
R11296 gnd.n2721 gnd.n2718 9.3005
R11297 gnd.n2717 gnd.n2695 9.3005
R11298 gnd.n2716 gnd.n2715 9.3005
R11299 gnd.n2712 gnd.n2696 9.3005
R11300 gnd.n2711 gnd.n2708 9.3005
R11301 gnd.n2707 gnd.n2697 9.3005
R11302 gnd.n2706 gnd.n2705 9.3005
R11303 gnd.n2702 gnd.n2698 9.3005
R11304 gnd.n2701 gnd.n1136 9.3005
R11305 gnd.n2740 gnd.n2685 9.3005
R11306 gnd.n2742 gnd.n2741 9.3005
R11307 gnd.n4738 gnd.n1424 9.3005
R11308 gnd.n4739 gnd.n1423 9.3005
R11309 gnd.n1422 gnd.n1419 9.3005
R11310 gnd.n4744 gnd.n1418 9.3005
R11311 gnd.n4745 gnd.n1417 9.3005
R11312 gnd.n4746 gnd.n1416 9.3005
R11313 gnd.n1415 gnd.n1412 9.3005
R11314 gnd.n4751 gnd.n1411 9.3005
R11315 gnd.n4753 gnd.n1408 9.3005
R11316 gnd.n4754 gnd.n1407 9.3005
R11317 gnd.n1406 gnd.n1403 9.3005
R11318 gnd.n4759 gnd.n1402 9.3005
R11319 gnd.n4760 gnd.n1401 9.3005
R11320 gnd.n4761 gnd.n1400 9.3005
R11321 gnd.n1399 gnd.n1396 9.3005
R11322 gnd.n4766 gnd.n1395 9.3005
R11323 gnd.n4767 gnd.n1394 9.3005
R11324 gnd.n4768 gnd.n1393 9.3005
R11325 gnd.n1392 gnd.n1389 9.3005
R11326 gnd.n4773 gnd.n1388 9.3005
R11327 gnd.n4774 gnd.n1387 9.3005
R11328 gnd.n4775 gnd.n1386 9.3005
R11329 gnd.n1385 gnd.n1382 9.3005
R11330 gnd.n1384 gnd.n1380 9.3005
R11331 gnd.n4782 gnd.n1379 9.3005
R11332 gnd.n4784 gnd.n4783 9.3005
R11333 gnd.n2381 gnd.n2380 9.3005
R11334 gnd.n2389 gnd.n2388 9.3005
R11335 gnd.n2390 gnd.n2378 9.3005
R11336 gnd.n2392 gnd.n2391 9.3005
R11337 gnd.n2376 gnd.n2375 9.3005
R11338 gnd.n2399 gnd.n2398 9.3005
R11339 gnd.n2400 gnd.n2374 9.3005
R11340 gnd.n2402 gnd.n2401 9.3005
R11341 gnd.n2372 gnd.n2369 9.3005
R11342 gnd.n2409 gnd.n2408 9.3005
R11343 gnd.n2410 gnd.n2368 9.3005
R11344 gnd.n2412 gnd.n2411 9.3005
R11345 gnd.n2366 gnd.n2365 9.3005
R11346 gnd.n2419 gnd.n2418 9.3005
R11347 gnd.n2420 gnd.n2364 9.3005
R11348 gnd.n2422 gnd.n2421 9.3005
R11349 gnd.n2362 gnd.n2361 9.3005
R11350 gnd.n2429 gnd.n2428 9.3005
R11351 gnd.n2430 gnd.n2360 9.3005
R11352 gnd.n2432 gnd.n2431 9.3005
R11353 gnd.n2358 gnd.n2357 9.3005
R11354 gnd.n2439 gnd.n2438 9.3005
R11355 gnd.n2440 gnd.n2356 9.3005
R11356 gnd.n2442 gnd.n2441 9.3005
R11357 gnd.n2354 gnd.n2353 9.3005
R11358 gnd.n2449 gnd.n2448 9.3005
R11359 gnd.n2450 gnd.n2352 9.3005
R11360 gnd.n2452 gnd.n2451 9.3005
R11361 gnd.n2350 gnd.n2347 9.3005
R11362 gnd.n2458 gnd.n2457 9.3005
R11363 gnd.n2379 gnd.n1425 9.3005
R11364 gnd.n1158 gnd.n1138 9.3005
R11365 gnd.n2666 gnd.n1159 9.3005
R11366 gnd.n4914 gnd.n1160 9.3005
R11367 gnd.n4913 gnd.n1161 9.3005
R11368 gnd.n4912 gnd.n1162 9.3005
R11369 gnd.n2672 gnd.n1163 9.3005
R11370 gnd.n4902 gnd.n1179 9.3005
R11371 gnd.n4901 gnd.n1180 9.3005
R11372 gnd.n4900 gnd.n1181 9.3005
R11373 gnd.n2679 gnd.n1182 9.3005
R11374 gnd.n4890 gnd.n1199 9.3005
R11375 gnd.n4889 gnd.n1200 9.3005
R11376 gnd.n4888 gnd.n1201 9.3005
R11377 gnd.n2662 gnd.n1202 9.3005
R11378 gnd.n4878 gnd.n1219 9.3005
R11379 gnd.n4877 gnd.n1220 9.3005
R11380 gnd.n4876 gnd.n1221 9.3005
R11381 gnd.n2657 gnd.n1222 9.3005
R11382 gnd.n4866 gnd.n1240 9.3005
R11383 gnd.n4865 gnd.n1241 9.3005
R11384 gnd.n4864 gnd.n1242 9.3005
R11385 gnd.n2644 gnd.n1243 9.3005
R11386 gnd.n2857 gnd.n2856 9.3005
R11387 gnd.n2645 gnd.n2629 9.3005
R11388 gnd.n2882 gnd.n2630 9.3005
R11389 gnd.n2881 gnd.n2631 9.3005
R11390 gnd.n2880 gnd.n2632 9.3005
R11391 gnd.n2609 gnd.n2608 9.3005
R11392 gnd.n2906 gnd.n2905 9.3005
R11393 gnd.n2907 gnd.n1268 9.3005
R11394 gnd.n4852 gnd.n1269 9.3005
R11395 gnd.n4851 gnd.n1270 9.3005
R11396 gnd.n4850 gnd.n1271 9.3005
R11397 gnd.n2914 gnd.n1272 9.3005
R11398 gnd.n4840 gnd.n1288 9.3005
R11399 gnd.n4839 gnd.n1289 9.3005
R11400 gnd.n4838 gnd.n1290 9.3005
R11401 gnd.n2920 gnd.n1291 9.3005
R11402 gnd.n4828 gnd.n1308 9.3005
R11403 gnd.n4827 gnd.n1309 9.3005
R11404 gnd.n4826 gnd.n1310 9.3005
R11405 gnd.n2991 gnd.n1311 9.3005
R11406 gnd.n4816 gnd.n1328 9.3005
R11407 gnd.n4815 gnd.n1329 9.3005
R11408 gnd.n4814 gnd.n1330 9.3005
R11409 gnd.n3006 gnd.n1331 9.3005
R11410 gnd.n4804 gnd.n1348 9.3005
R11411 gnd.n4803 gnd.n1349 9.3005
R11412 gnd.n4802 gnd.n1350 9.3005
R11413 gnd.n3013 gnd.n1351 9.3005
R11414 gnd.n4792 gnd.n1369 9.3005
R11415 gnd.n4791 gnd.n1370 9.3005
R11416 gnd.n4790 gnd.n1371 9.3005
R11417 gnd.n4926 gnd.n1137 9.3005
R11418 gnd.n1139 gnd.n1138 9.3005
R11419 gnd.n2667 gnd.n2666 9.3005
R11420 gnd.n2668 gnd.n1160 9.3005
R11421 gnd.n2670 gnd.n1161 9.3005
R11422 gnd.n2671 gnd.n1162 9.3005
R11423 gnd.n2674 gnd.n2672 9.3005
R11424 gnd.n2675 gnd.n1179 9.3005
R11425 gnd.n2677 gnd.n1180 9.3005
R11426 gnd.n2678 gnd.n1181 9.3005
R11427 gnd.n2768 gnd.n2679 9.3005
R11428 gnd.n2769 gnd.n1199 9.3005
R11429 gnd.n2770 gnd.n1200 9.3005
R11430 gnd.n2661 gnd.n1201 9.3005
R11431 gnd.n2821 gnd.n2662 9.3005
R11432 gnd.n2822 gnd.n1219 9.3005
R11433 gnd.n2823 gnd.n1220 9.3005
R11434 gnd.n2656 gnd.n1221 9.3005
R11435 gnd.n2836 gnd.n2657 9.3005
R11436 gnd.n2837 gnd.n1240 9.3005
R11437 gnd.n2839 gnd.n1241 9.3005
R11438 gnd.n2838 gnd.n1242 9.3005
R11439 gnd.n2647 gnd.n2644 9.3005
R11440 gnd.n2856 gnd.n2855 9.3005
R11441 gnd.n2854 gnd.n2645 9.3005
R11442 gnd.n2651 gnd.n2630 9.3005
R11443 gnd.n2650 gnd.n2631 9.3005
R11444 gnd.n2649 gnd.n2632 9.3005
R11445 gnd.n2648 gnd.n2608 9.3005
R11446 gnd.n2906 gnd.n2607 9.3005
R11447 gnd.n2908 gnd.n2907 9.3005
R11448 gnd.n2909 gnd.n1269 9.3005
R11449 gnd.n2912 gnd.n1270 9.3005
R11450 gnd.n2913 gnd.n1271 9.3005
R11451 gnd.n2918 gnd.n2914 9.3005
R11452 gnd.n2919 gnd.n1288 9.3005
R11453 gnd.n2923 gnd.n1289 9.3005
R11454 gnd.n2922 gnd.n1290 9.3005
R11455 gnd.n2921 gnd.n2920 9.3005
R11456 gnd.n2581 gnd.n1308 9.3005
R11457 gnd.n2989 gnd.n1309 9.3005
R11458 gnd.n2990 gnd.n1310 9.3005
R11459 gnd.n2992 gnd.n2991 9.3005
R11460 gnd.n2576 gnd.n1328 9.3005
R11461 gnd.n3004 gnd.n1329 9.3005
R11462 gnd.n3005 gnd.n1330 9.3005
R11463 gnd.n3007 gnd.n3006 9.3005
R11464 gnd.n3008 gnd.n1348 9.3005
R11465 gnd.n3011 gnd.n1349 9.3005
R11466 gnd.n3012 gnd.n1350 9.3005
R11467 gnd.n3016 gnd.n3013 9.3005
R11468 gnd.n3017 gnd.n1369 9.3005
R11469 gnd.n3019 gnd.n1370 9.3005
R11470 gnd.n3018 gnd.n1371 9.3005
R11471 gnd.n4926 gnd.n4925 9.3005
R11472 gnd.n4930 gnd.n4929 9.3005
R11473 gnd.n4933 gnd.n1132 9.3005
R11474 gnd.n4934 gnd.n1131 9.3005
R11475 gnd.n4937 gnd.n1130 9.3005
R11476 gnd.n4938 gnd.n1129 9.3005
R11477 gnd.n4941 gnd.n1128 9.3005
R11478 gnd.n4942 gnd.n1127 9.3005
R11479 gnd.n4945 gnd.n1126 9.3005
R11480 gnd.n4946 gnd.n1125 9.3005
R11481 gnd.n4949 gnd.n1124 9.3005
R11482 gnd.n4950 gnd.n1123 9.3005
R11483 gnd.n4953 gnd.n1122 9.3005
R11484 gnd.n4954 gnd.n1121 9.3005
R11485 gnd.n4957 gnd.n1120 9.3005
R11486 gnd.n4958 gnd.n1119 9.3005
R11487 gnd.n4961 gnd.n1118 9.3005
R11488 gnd.n4962 gnd.n1117 9.3005
R11489 gnd.n4965 gnd.n1116 9.3005
R11490 gnd.n4966 gnd.n1115 9.3005
R11491 gnd.n4969 gnd.n1114 9.3005
R11492 gnd.n4973 gnd.n1110 9.3005
R11493 gnd.n4974 gnd.n1109 9.3005
R11494 gnd.n4977 gnd.n1108 9.3005
R11495 gnd.n4978 gnd.n1107 9.3005
R11496 gnd.n4981 gnd.n1106 9.3005
R11497 gnd.n4982 gnd.n1105 9.3005
R11498 gnd.n4985 gnd.n1104 9.3005
R11499 gnd.n4986 gnd.n1103 9.3005
R11500 gnd.n4989 gnd.n1102 9.3005
R11501 gnd.n4990 gnd.n1101 9.3005
R11502 gnd.n4993 gnd.n1100 9.3005
R11503 gnd.n4994 gnd.n1099 9.3005
R11504 gnd.n4997 gnd.n1098 9.3005
R11505 gnd.n4998 gnd.n1097 9.3005
R11506 gnd.n5001 gnd.n1096 9.3005
R11507 gnd.n5002 gnd.n1095 9.3005
R11508 gnd.n5005 gnd.n1094 9.3005
R11509 gnd.n5006 gnd.n1093 9.3005
R11510 gnd.n5009 gnd.n1092 9.3005
R11511 gnd.n5011 gnd.n1089 9.3005
R11512 gnd.n5014 gnd.n1088 9.3005
R11513 gnd.n5015 gnd.n1087 9.3005
R11514 gnd.n5018 gnd.n1086 9.3005
R11515 gnd.n5019 gnd.n1085 9.3005
R11516 gnd.n5022 gnd.n1084 9.3005
R11517 gnd.n5023 gnd.n1083 9.3005
R11518 gnd.n5026 gnd.n1082 9.3005
R11519 gnd.n5027 gnd.n1081 9.3005
R11520 gnd.n5030 gnd.n1080 9.3005
R11521 gnd.n5031 gnd.n1079 9.3005
R11522 gnd.n5034 gnd.n1078 9.3005
R11523 gnd.n5035 gnd.n1077 9.3005
R11524 gnd.n5038 gnd.n1076 9.3005
R11525 gnd.n5040 gnd.n1075 9.3005
R11526 gnd.n5041 gnd.n1074 9.3005
R11527 gnd.n5042 gnd.n1073 9.3005
R11528 gnd.n5043 gnd.n1072 9.3005
R11529 gnd.n4970 gnd.n1111 9.3005
R11530 gnd.n4928 gnd.n1133 9.3005
R11531 gnd.n4920 gnd.n1147 9.3005
R11532 gnd.n4919 gnd.n1148 9.3005
R11533 gnd.n4918 gnd.n1149 9.3005
R11534 gnd.n1169 gnd.n1150 9.3005
R11535 gnd.n4908 gnd.n1170 9.3005
R11536 gnd.n4907 gnd.n1171 9.3005
R11537 gnd.n4906 gnd.n1172 9.3005
R11538 gnd.n1188 gnd.n1173 9.3005
R11539 gnd.n4896 gnd.n1189 9.3005
R11540 gnd.n4895 gnd.n1190 9.3005
R11541 gnd.n4894 gnd.n1191 9.3005
R11542 gnd.n1209 gnd.n1192 9.3005
R11543 gnd.n4884 gnd.n1210 9.3005
R11544 gnd.n4883 gnd.n1211 9.3005
R11545 gnd.n4882 gnd.n1212 9.3005
R11546 gnd.n1229 gnd.n1213 9.3005
R11547 gnd.n4872 gnd.n1230 9.3005
R11548 gnd.n4871 gnd.n1231 9.3005
R11549 gnd.n4870 gnd.n1232 9.3005
R11550 gnd.n1250 gnd.n1233 9.3005
R11551 gnd.n4860 gnd.n1251 9.3005
R11552 gnd.n1260 gnd.n1253 9.3005
R11553 gnd.n4846 gnd.n1278 9.3005
R11554 gnd.n4845 gnd.n1279 9.3005
R11555 gnd.n4844 gnd.n1280 9.3005
R11556 gnd.n1298 gnd.n1281 9.3005
R11557 gnd.n4834 gnd.n1299 9.3005
R11558 gnd.n4833 gnd.n1300 9.3005
R11559 gnd.n4832 gnd.n1301 9.3005
R11560 gnd.n1317 gnd.n1302 9.3005
R11561 gnd.n4822 gnd.n1318 9.3005
R11562 gnd.n4821 gnd.n1319 9.3005
R11563 gnd.n4820 gnd.n1320 9.3005
R11564 gnd.n1338 gnd.n1321 9.3005
R11565 gnd.n4810 gnd.n1339 9.3005
R11566 gnd.n4809 gnd.n1340 9.3005
R11567 gnd.n4808 gnd.n1341 9.3005
R11568 gnd.n1358 gnd.n1342 9.3005
R11569 gnd.n4798 gnd.n1359 9.3005
R11570 gnd.n4797 gnd.n1360 9.3005
R11571 gnd.n4796 gnd.n1361 9.3005
R11572 gnd.n1378 gnd.n1362 9.3005
R11573 gnd.n4786 gnd.n4785 9.3005
R11574 gnd.n1146 gnd.n1145 9.3005
R11575 gnd.n4857 gnd.n1258 9.3005
R11576 gnd.n4857 gnd.n4856 9.3005
R11577 gnd.n2784 gnd.n2783 9.3005
R11578 gnd.n2795 gnd.n2794 9.3005
R11579 gnd.n2796 gnd.n2782 9.3005
R11580 gnd.n2816 gnd.n2797 9.3005
R11581 gnd.n2815 gnd.n2798 9.3005
R11582 gnd.n2814 gnd.n2799 9.3005
R11583 gnd.n2802 gnd.n2800 9.3005
R11584 gnd.n2810 gnd.n2803 9.3005
R11585 gnd.n2809 gnd.n2804 9.3005
R11586 gnd.n2808 gnd.n2806 9.3005
R11587 gnd.n2805 gnd.n2638 9.3005
R11588 gnd.n2790 gnd.n2789 9.3005
R11589 gnd.n2786 gnd.n966 9.3005
R11590 gnd.n6467 gnd.n965 9.3005
R11591 gnd.n6468 gnd.n964 9.3005
R11592 gnd.n6469 gnd.n963 9.3005
R11593 gnd.n962 gnd.n958 9.3005
R11594 gnd.n6475 gnd.n957 9.3005
R11595 gnd.n6476 gnd.n956 9.3005
R11596 gnd.n6477 gnd.n955 9.3005
R11597 gnd.n954 gnd.n950 9.3005
R11598 gnd.n6483 gnd.n949 9.3005
R11599 gnd.n6484 gnd.n948 9.3005
R11600 gnd.n6485 gnd.n947 9.3005
R11601 gnd.n946 gnd.n942 9.3005
R11602 gnd.n6491 gnd.n941 9.3005
R11603 gnd.n6492 gnd.n940 9.3005
R11604 gnd.n6493 gnd.n939 9.3005
R11605 gnd.n938 gnd.n934 9.3005
R11606 gnd.n6499 gnd.n933 9.3005
R11607 gnd.n6500 gnd.n932 9.3005
R11608 gnd.n6501 gnd.n931 9.3005
R11609 gnd.n930 gnd.n926 9.3005
R11610 gnd.n6507 gnd.n925 9.3005
R11611 gnd.n6508 gnd.n924 9.3005
R11612 gnd.n6509 gnd.n923 9.3005
R11613 gnd.n922 gnd.n918 9.3005
R11614 gnd.n6515 gnd.n917 9.3005
R11615 gnd.n6516 gnd.n916 9.3005
R11616 gnd.n6517 gnd.n915 9.3005
R11617 gnd.n914 gnd.n910 9.3005
R11618 gnd.n6523 gnd.n909 9.3005
R11619 gnd.n6524 gnd.n908 9.3005
R11620 gnd.n6525 gnd.n907 9.3005
R11621 gnd.n906 gnd.n902 9.3005
R11622 gnd.n6531 gnd.n901 9.3005
R11623 gnd.n6532 gnd.n900 9.3005
R11624 gnd.n6533 gnd.n899 9.3005
R11625 gnd.n898 gnd.n894 9.3005
R11626 gnd.n6539 gnd.n893 9.3005
R11627 gnd.n6540 gnd.n892 9.3005
R11628 gnd.n6541 gnd.n891 9.3005
R11629 gnd.n890 gnd.n886 9.3005
R11630 gnd.n6547 gnd.n885 9.3005
R11631 gnd.n6548 gnd.n884 9.3005
R11632 gnd.n6549 gnd.n883 9.3005
R11633 gnd.n882 gnd.n878 9.3005
R11634 gnd.n6555 gnd.n877 9.3005
R11635 gnd.n6556 gnd.n876 9.3005
R11636 gnd.n6557 gnd.n875 9.3005
R11637 gnd.n874 gnd.n870 9.3005
R11638 gnd.n6563 gnd.n869 9.3005
R11639 gnd.n6564 gnd.n868 9.3005
R11640 gnd.n6565 gnd.n867 9.3005
R11641 gnd.n866 gnd.n862 9.3005
R11642 gnd.n6571 gnd.n861 9.3005
R11643 gnd.n6572 gnd.n860 9.3005
R11644 gnd.n6573 gnd.n859 9.3005
R11645 gnd.n858 gnd.n854 9.3005
R11646 gnd.n6579 gnd.n853 9.3005
R11647 gnd.n6580 gnd.n852 9.3005
R11648 gnd.n6581 gnd.n851 9.3005
R11649 gnd.n850 gnd.n846 9.3005
R11650 gnd.n6587 gnd.n845 9.3005
R11651 gnd.n6588 gnd.n844 9.3005
R11652 gnd.n6589 gnd.n843 9.3005
R11653 gnd.n842 gnd.n838 9.3005
R11654 gnd.n6595 gnd.n837 9.3005
R11655 gnd.n6596 gnd.n836 9.3005
R11656 gnd.n6597 gnd.n835 9.3005
R11657 gnd.n834 gnd.n830 9.3005
R11658 gnd.n6603 gnd.n829 9.3005
R11659 gnd.n6604 gnd.n828 9.3005
R11660 gnd.n6605 gnd.n827 9.3005
R11661 gnd.n826 gnd.n822 9.3005
R11662 gnd.n6611 gnd.n821 9.3005
R11663 gnd.n6612 gnd.n820 9.3005
R11664 gnd.n6613 gnd.n819 9.3005
R11665 gnd.n818 gnd.n814 9.3005
R11666 gnd.n6619 gnd.n813 9.3005
R11667 gnd.n6620 gnd.n812 9.3005
R11668 gnd.n6621 gnd.n811 9.3005
R11669 gnd.n810 gnd.n806 9.3005
R11670 gnd.n6627 gnd.n805 9.3005
R11671 gnd.n6628 gnd.n804 9.3005
R11672 gnd.n6629 gnd.n803 9.3005
R11673 gnd.n2788 gnd.n2787 9.3005
R11674 gnd.n3930 gnd.n3929 9.3005
R11675 gnd.n3148 gnd.n2329 9.3005
R11676 gnd.n3151 gnd.n3150 9.3005
R11677 gnd.n3149 gnd.n2330 9.3005
R11678 gnd.n2306 gnd.n2305 9.3005
R11679 gnd.n3177 gnd.n3176 9.3005
R11680 gnd.n3178 gnd.n2303 9.3005
R11681 gnd.n3181 gnd.n3180 9.3005
R11682 gnd.n3179 gnd.n2304 9.3005
R11683 gnd.n2282 gnd.n2281 9.3005
R11684 gnd.n3207 gnd.n3206 9.3005
R11685 gnd.n3208 gnd.n2279 9.3005
R11686 gnd.n3211 gnd.n3210 9.3005
R11687 gnd.n3209 gnd.n2280 9.3005
R11688 gnd.n2257 gnd.n2256 9.3005
R11689 gnd.n3247 gnd.n3246 9.3005
R11690 gnd.n3248 gnd.n2254 9.3005
R11691 gnd.n3254 gnd.n3253 9.3005
R11692 gnd.n3252 gnd.n2255 9.3005
R11693 gnd.n3251 gnd.n3250 9.3005
R11694 gnd.n2173 gnd.n2172 9.3005
R11695 gnd.n3303 gnd.n3302 9.3005
R11696 gnd.n3304 gnd.n2170 9.3005
R11697 gnd.n3326 gnd.n3325 9.3005
R11698 gnd.n3324 gnd.n2171 9.3005
R11699 gnd.n3323 gnd.n3322 9.3005
R11700 gnd.n3321 gnd.n3305 9.3005
R11701 gnd.n3320 gnd.n3319 9.3005
R11702 gnd.n3318 gnd.n3312 9.3005
R11703 gnd.n3317 gnd.n3316 9.3005
R11704 gnd.n3315 gnd.n3314 9.3005
R11705 gnd.n3313 gnd.n2123 9.3005
R11706 gnd.n2121 gnd.n2120 9.3005
R11707 gnd.n3405 gnd.n3404 9.3005
R11708 gnd.n3406 gnd.n2119 9.3005
R11709 gnd.n3408 gnd.n3407 9.3005
R11710 gnd.n2096 gnd.n2094 9.3005
R11711 gnd.n3456 gnd.n3455 9.3005
R11712 gnd.n3454 gnd.n2095 9.3005
R11713 gnd.n3453 gnd.n3452 9.3005
R11714 gnd.n2073 gnd.n2071 9.3005
R11715 gnd.n3514 gnd.n3513 9.3005
R11716 gnd.n3512 gnd.n2072 9.3005
R11717 gnd.n3511 gnd.n3510 9.3005
R11718 gnd.n3509 gnd.n2074 9.3005
R11719 gnd.n3508 gnd.n3507 9.3005
R11720 gnd.n3506 gnd.n3495 9.3005
R11721 gnd.n3505 gnd.n3504 9.3005
R11722 gnd.n3503 gnd.n3496 9.3005
R11723 gnd.n3502 gnd.n3501 9.3005
R11724 gnd.n2013 gnd.n2012 9.3005
R11725 gnd.n3623 gnd.n3622 9.3005
R11726 gnd.n3624 gnd.n2010 9.3005
R11727 gnd.n3627 gnd.n3626 9.3005
R11728 gnd.n3625 gnd.n2011 9.3005
R11729 gnd.n1984 gnd.n1983 9.3005
R11730 gnd.n3662 gnd.n3661 9.3005
R11731 gnd.n3663 gnd.n1981 9.3005
R11732 gnd.n3672 gnd.n3671 9.3005
R11733 gnd.n3670 gnd.n1982 9.3005
R11734 gnd.n3669 gnd.n3668 9.3005
R11735 gnd.n3667 gnd.n3664 9.3005
R11736 gnd.n1949 gnd.n1948 9.3005
R11737 gnd.n3719 gnd.n3718 9.3005
R11738 gnd.n3720 gnd.n1947 9.3005
R11739 gnd.n3722 gnd.n3721 9.3005
R11740 gnd.n3725 gnd.n1946 9.3005
R11741 gnd.n3727 gnd.n3726 9.3005
R11742 gnd.n3728 gnd.n1945 9.3005
R11743 gnd.n3730 gnd.n3729 9.3005
R11744 gnd.n3733 gnd.n1944 9.3005
R11745 gnd.n3735 gnd.n3734 9.3005
R11746 gnd.n3736 gnd.n1943 9.3005
R11747 gnd.n3738 gnd.n3737 9.3005
R11748 gnd.n3741 gnd.n1942 9.3005
R11749 gnd.n3743 gnd.n3742 9.3005
R11750 gnd.n3744 gnd.n1941 9.3005
R11751 gnd.n3746 gnd.n3745 9.3005
R11752 gnd.n3749 gnd.n1940 9.3005
R11753 gnd.n3751 gnd.n3750 9.3005
R11754 gnd.n3752 gnd.n1938 9.3005
R11755 gnd.n3933 gnd.n3932 9.3005
R11756 gnd.n3931 gnd.n1939 9.3005
R11757 gnd.n3147 gnd.n3146 9.3005
R11758 gnd.n3073 gnd.n2331 9.3005
R11759 gnd.n2894 gnd.n2616 9.3005
R11760 gnd.n2896 gnd.n2895 9.3005
R11761 gnd.n2602 gnd.n2600 9.3005
R11762 gnd.n2937 gnd.n2936 9.3005
R11763 gnd.n2935 gnd.n2601 9.3005
R11764 gnd.n2934 gnd.n2933 9.3005
R11765 gnd.n2932 gnd.n2603 9.3005
R11766 gnd.n2931 gnd.n2930 9.3005
R11767 gnd.n2929 gnd.n2606 9.3005
R11768 gnd.n2928 gnd.n2927 9.3005
R11769 gnd.n2584 gnd.n2583 9.3005
R11770 gnd.n2982 gnd.n2981 9.3005
R11771 gnd.n2983 gnd.n2582 9.3005
R11772 gnd.n2985 gnd.n2984 9.3005
R11773 gnd.n2579 gnd.n2578 9.3005
R11774 gnd.n2997 gnd.n2996 9.3005
R11775 gnd.n2998 gnd.n2577 9.3005
R11776 gnd.n3000 gnd.n2999 9.3005
R11777 gnd.n2570 gnd.n2568 9.3005
R11778 gnd.n3034 gnd.n3033 9.3005
R11779 gnd.n3032 gnd.n2569 9.3005
R11780 gnd.n3031 gnd.n3030 9.3005
R11781 gnd.n3029 gnd.n2571 9.3005
R11782 gnd.n3028 gnd.n3027 9.3005
R11783 gnd.n3026 gnd.n2574 9.3005
R11784 gnd.n3025 gnd.n3024 9.3005
R11785 gnd.n3023 gnd.n2575 9.3005
R11786 gnd.n3122 gnd.n3121 9.3005
R11787 gnd.n3120 gnd.n3119 9.3005
R11788 gnd.n2470 gnd.n2469 9.3005
R11789 gnd.n3114 gnd.n3113 9.3005
R11790 gnd.n3112 gnd.n3111 9.3005
R11791 gnd.n2480 gnd.n2479 9.3005
R11792 gnd.n3106 gnd.n3105 9.3005
R11793 gnd.n3104 gnd.n3103 9.3005
R11794 gnd.n2491 gnd.n2490 9.3005
R11795 gnd.n3098 gnd.n3097 9.3005
R11796 gnd.n3096 gnd.n3095 9.3005
R11797 gnd.n2501 gnd.n2500 9.3005
R11798 gnd.n3090 gnd.n3089 9.3005
R11799 gnd.n3088 gnd.n3087 9.3005
R11800 gnd.n2512 gnd.n2511 9.3005
R11801 gnd.n3082 gnd.n3081 9.3005
R11802 gnd.n3080 gnd.n2524 9.3005
R11803 gnd.n3079 gnd.n3076 9.3005
R11804 gnd.n2465 gnd.n2460 9.3005
R11805 gnd.n3075 gnd.n3074 9.3005
R11806 gnd.n2528 gnd.n2526 9.3005
R11807 gnd.n2549 gnd.n2518 9.3005
R11808 gnd.n3084 gnd.n3083 9.3005
R11809 gnd.n3086 gnd.n3085 9.3005
R11810 gnd.n2505 gnd.n2504 9.3005
R11811 gnd.n3092 gnd.n3091 9.3005
R11812 gnd.n3094 gnd.n3093 9.3005
R11813 gnd.n2495 gnd.n2494 9.3005
R11814 gnd.n3100 gnd.n3099 9.3005
R11815 gnd.n3102 gnd.n3101 9.3005
R11816 gnd.n2484 gnd.n2483 9.3005
R11817 gnd.n3108 gnd.n3107 9.3005
R11818 gnd.n3110 gnd.n3109 9.3005
R11819 gnd.n2474 gnd.n2473 9.3005
R11820 gnd.n3116 gnd.n3115 9.3005
R11821 gnd.n3118 gnd.n3117 9.3005
R11822 gnd.n2464 gnd.n2463 9.3005
R11823 gnd.n3124 gnd.n3123 9.3005
R11824 gnd.n3126 gnd.n3125 9.3005
R11825 gnd.n3127 gnd.n2346 9.3005
R11826 gnd.n3130 gnd.n3129 9.3005
R11827 gnd.n3131 gnd.n2342 9.3005
R11828 gnd.n3133 gnd.n3132 9.3005
R11829 gnd.n3134 gnd.n2341 9.3005
R11830 gnd.n3136 gnd.n3135 9.3005
R11831 gnd.n3137 gnd.n2338 9.3005
R11832 gnd.n3139 gnd.n3138 9.3005
R11833 gnd.n3140 gnd.n2337 9.3005
R11834 gnd.n2316 gnd.n2315 9.3005
R11835 gnd.n3168 gnd.n3167 9.3005
R11836 gnd.n3169 gnd.n2313 9.3005
R11837 gnd.n3172 gnd.n3171 9.3005
R11838 gnd.n3170 gnd.n2314 9.3005
R11839 gnd.n2291 gnd.n2290 9.3005
R11840 gnd.n3198 gnd.n3197 9.3005
R11841 gnd.n3199 gnd.n2288 9.3005
R11842 gnd.n3202 gnd.n3201 9.3005
R11843 gnd.n3200 gnd.n2289 9.3005
R11844 gnd.n2266 gnd.n2265 9.3005
R11845 gnd.n3238 gnd.n3237 9.3005
R11846 gnd.n3239 gnd.n2263 9.3005
R11847 gnd.n3242 gnd.n3241 9.3005
R11848 gnd.n3240 gnd.n2264 9.3005
R11849 gnd.n1498 gnd.n1496 9.3005
R11850 gnd.n4660 gnd.n4659 9.3005
R11851 gnd.n4658 gnd.n1497 9.3005
R11852 gnd.n4657 gnd.n4656 9.3005
R11853 gnd.n4655 gnd.n1499 9.3005
R11854 gnd.n4654 gnd.n4653 9.3005
R11855 gnd.n4652 gnd.n1503 9.3005
R11856 gnd.n4651 gnd.n4650 9.3005
R11857 gnd.n4649 gnd.n1504 9.3005
R11858 gnd.n4648 gnd.n4647 9.3005
R11859 gnd.n4646 gnd.n1508 9.3005
R11860 gnd.n4645 gnd.n4644 9.3005
R11861 gnd.n4643 gnd.n1509 9.3005
R11862 gnd.n4642 gnd.n4641 9.3005
R11863 gnd.n4640 gnd.n1513 9.3005
R11864 gnd.n4639 gnd.n4638 9.3005
R11865 gnd.n4637 gnd.n1514 9.3005
R11866 gnd.n4636 gnd.n4635 9.3005
R11867 gnd.n4634 gnd.n1518 9.3005
R11868 gnd.n4633 gnd.n4632 9.3005
R11869 gnd.n4631 gnd.n1519 9.3005
R11870 gnd.n4630 gnd.n4629 9.3005
R11871 gnd.n4628 gnd.n1523 9.3005
R11872 gnd.n4627 gnd.n4626 9.3005
R11873 gnd.n4625 gnd.n1524 9.3005
R11874 gnd.n4624 gnd.n4623 9.3005
R11875 gnd.n4622 gnd.n1528 9.3005
R11876 gnd.n4621 gnd.n4620 9.3005
R11877 gnd.n4619 gnd.n1529 9.3005
R11878 gnd.n4618 gnd.n4617 9.3005
R11879 gnd.n4616 gnd.n1533 9.3005
R11880 gnd.n4615 gnd.n4614 9.3005
R11881 gnd.n4613 gnd.n1534 9.3005
R11882 gnd.n4612 gnd.n4611 9.3005
R11883 gnd.n4610 gnd.n1538 9.3005
R11884 gnd.n4609 gnd.n4608 9.3005
R11885 gnd.n4607 gnd.n1539 9.3005
R11886 gnd.n4606 gnd.n4605 9.3005
R11887 gnd.n4604 gnd.n1543 9.3005
R11888 gnd.n4603 gnd.n4602 9.3005
R11889 gnd.n4601 gnd.n1544 9.3005
R11890 gnd.n4600 gnd.n4599 9.3005
R11891 gnd.n4598 gnd.n1548 9.3005
R11892 gnd.n4597 gnd.n4596 9.3005
R11893 gnd.n4595 gnd.n1549 9.3005
R11894 gnd.n4594 gnd.n4593 9.3005
R11895 gnd.n4592 gnd.n1553 9.3005
R11896 gnd.n4591 gnd.n4590 9.3005
R11897 gnd.n4589 gnd.n1554 9.3005
R11898 gnd.n4588 gnd.n4587 9.3005
R11899 gnd.n4586 gnd.n1558 9.3005
R11900 gnd.n4585 gnd.n4584 9.3005
R11901 gnd.n4583 gnd.n1559 9.3005
R11902 gnd.n4582 gnd.n4581 9.3005
R11903 gnd.n4580 gnd.n1563 9.3005
R11904 gnd.n4579 gnd.n4578 9.3005
R11905 gnd.n4577 gnd.n1564 9.3005
R11906 gnd.n4576 gnd.n4575 9.3005
R11907 gnd.n4574 gnd.n1568 9.3005
R11908 gnd.n4573 gnd.n4572 9.3005
R11909 gnd.n4571 gnd.n1569 9.3005
R11910 gnd.n4570 gnd.n4569 9.3005
R11911 gnd.n4568 gnd.n1573 9.3005
R11912 gnd.n4567 gnd.n4566 9.3005
R11913 gnd.n4565 gnd.n1574 9.3005
R11914 gnd.n4564 gnd.n1577 9.3005
R11915 gnd.n3142 gnd.n3141 9.3005
R11916 gnd.n3819 gnd.n3818 9.3005
R11917 gnd.n3814 gnd.n3813 9.3005
R11918 gnd.n3826 gnd.n3825 9.3005
R11919 gnd.n3827 gnd.n3812 9.3005
R11920 gnd.n3830 gnd.n3829 9.3005
R11921 gnd.n3828 gnd.n3810 9.3005
R11922 gnd.n3817 gnd.n3816 9.3005
R11923 gnd.n3918 gnd.n3766 9.3005
R11924 gnd.n3779 gnd.n3775 9.3005
R11925 gnd.n3912 gnd.n3911 9.3005
R11926 gnd.n3900 gnd.n3777 9.3005
R11927 gnd.n3899 gnd.n3898 9.3005
R11928 gnd.n3788 gnd.n3784 9.3005
R11929 gnd.n3892 gnd.n3891 9.3005
R11930 gnd.n3881 gnd.n3786 9.3005
R11931 gnd.n3880 gnd.n3879 9.3005
R11932 gnd.n3797 gnd.n3793 9.3005
R11933 gnd.n3873 gnd.n3872 9.3005
R11934 gnd.n3862 gnd.n3795 9.3005
R11935 gnd.n3861 gnd.n3860 9.3005
R11936 gnd.n3806 gnd.n3802 9.3005
R11937 gnd.n3854 gnd.n3853 9.3005
R11938 gnd.n3843 gnd.n3804 9.3005
R11939 gnd.n3842 gnd.n3841 9.3005
R11940 gnd.n3920 gnd.n3919 9.3005
R11941 gnd.n3770 gnd.n3769 9.3005
R11942 gnd.n3837 gnd.n3836 9.3005
R11943 gnd.n3838 gnd.n3809 9.3005
R11944 gnd.n3845 gnd.n3844 9.3005
R11945 gnd.n3807 gnd.n3805 9.3005
R11946 gnd.n3852 gnd.n3851 9.3005
R11947 gnd.n3801 gnd.n3800 9.3005
R11948 gnd.n3864 gnd.n3863 9.3005
R11949 gnd.n3798 gnd.n3796 9.3005
R11950 gnd.n3871 gnd.n3870 9.3005
R11951 gnd.n3792 gnd.n3791 9.3005
R11952 gnd.n3883 gnd.n3882 9.3005
R11953 gnd.n3789 gnd.n3787 9.3005
R11954 gnd.n3890 gnd.n3889 9.3005
R11955 gnd.n3783 gnd.n3782 9.3005
R11956 gnd.n3902 gnd.n3901 9.3005
R11957 gnd.n3780 gnd.n3778 9.3005
R11958 gnd.n3910 gnd.n3909 9.3005
R11959 gnd.n3908 gnd.n3907 9.3005
R11960 gnd.n3922 gnd.n3921 9.3005
R11961 gnd.n3767 gnd.n3761 9.3005
R11962 gnd.n3768 gnd.n3760 9.3005
R11963 gnd.n3756 gnd.n3753 9.3005
R11964 gnd.n1805 gnd.n1804 9.3005
R11965 gnd.n4336 gnd.n4335 9.3005
R11966 gnd.n4337 gnd.n1803 9.3005
R11967 gnd.n4339 gnd.n4338 9.3005
R11968 gnd.n1768 gnd.n1767 9.3005
R11969 gnd.n4350 gnd.n4349 9.3005
R11970 gnd.n4351 gnd.n1766 9.3005
R11971 gnd.n4353 gnd.n4352 9.3005
R11972 gnd.n1758 gnd.n1756 9.3005
R11973 gnd.n4389 gnd.n4388 9.3005
R11974 gnd.n4387 gnd.n1757 9.3005
R11975 gnd.n4386 gnd.n4385 9.3005
R11976 gnd.n4384 gnd.n1759 9.3005
R11977 gnd.n4383 gnd.n4382 9.3005
R11978 gnd.n4381 gnd.n1762 9.3005
R11979 gnd.n4380 gnd.n4379 9.3005
R11980 gnd.n4378 gnd.n1763 9.3005
R11981 gnd.n4377 gnd.n4376 9.3005
R11982 gnd.n1741 gnd.n1740 9.3005
R11983 gnd.n4448 gnd.n4447 9.3005
R11984 gnd.n4449 gnd.n1738 9.3005
R11985 gnd.n4454 gnd.n4453 9.3005
R11986 gnd.n4452 gnd.n1739 9.3005
R11987 gnd.n4451 gnd.n4450 9.3005
R11988 gnd.n81 gnd.n79 9.3005
R11989 gnd.n3758 gnd.n3757 9.3005
R11990 gnd.t345 gnd.n5182 9.24152
R11991 gnd.n6435 gnd.t81 9.24152
R11992 gnd.t179 gnd.n1019 9.24152
R11993 gnd.n1152 gnd.t93 9.24152
R11994 gnd.n3037 gnd.t2 9.24152
R11995 gnd.n4733 gnd.n1464 9.24152
R11996 gnd.n4145 gnd.n1846 9.24152
R11997 gnd.n1800 gnd.t16 9.24152
R11998 gnd.n7563 gnd.t103 9.24152
R11999 gnd.t276 gnd.t345 8.92286
R12000 gnd.n3391 gnd.n2130 8.92286
R12001 gnd.n3437 gnd.n2100 8.92286
R12002 gnd.n3562 gnd.n2034 8.92286
R12003 gnd.n3632 gnd.n3631 8.92286
R12004 gnd.n3988 gnd.n1889 8.92286
R12005 gnd.n3985 gnd.t148 8.92286
R12006 gnd.n6289 gnd.n6264 8.92171
R12007 gnd.n6257 gnd.n6232 8.92171
R12008 gnd.n6225 gnd.n6200 8.92171
R12009 gnd.n6194 gnd.n6169 8.92171
R12010 gnd.n6162 gnd.n6137 8.92171
R12011 gnd.n6130 gnd.n6105 8.92171
R12012 gnd.n6098 gnd.n6073 8.92171
R12013 gnd.n6067 gnd.n6042 8.92171
R12014 gnd.n4010 gnd.n3992 8.72777
R12015 gnd.t321 gnd.n5293 8.60421
R12016 gnd.n5245 gnd.n5229 8.43656
R12017 gnd.n46 gnd.n30 8.43656
R12018 gnd.n3367 gnd.n2145 8.28555
R12019 gnd.n3458 gnd.n2083 8.28555
R12020 gnd.n3541 gnd.n2048 8.28555
R12021 gnd.n3597 gnd.n2001 8.28555
R12022 gnd.n6290 gnd.n6262 8.14595
R12023 gnd.n6258 gnd.n6230 8.14595
R12024 gnd.n6226 gnd.n6198 8.14595
R12025 gnd.n6195 gnd.n6167 8.14595
R12026 gnd.n6163 gnd.n6135 8.14595
R12027 gnd.n6131 gnd.n6103 8.14595
R12028 gnd.n6099 gnd.n6071 8.14595
R12029 gnd.n6068 gnd.n6040 8.14595
R12030 gnd.n2893 gnd.n0 8.10675
R12031 gnd.n7637 gnd.n7636 8.10675
R12032 gnd.n6295 gnd.n6294 7.97301
R12033 gnd.n5786 gnd.t319 7.9669
R12034 gnd.n7637 gnd.n78 7.86902
R12035 gnd.n3919 gnd.n3770 7.75808
R12036 gnd.n3080 gnd.n3079 7.75808
R12037 gnd.n7413 gnd.n349 7.75808
R12038 gnd.n2741 gnd.n2740 7.75808
R12039 gnd.n3274 gnd.n3273 7.64824
R12040 gnd.n3367 gnd.n2144 7.64824
R12041 gnd.t288 gnd.n3411 7.64824
R12042 gnd.n3459 gnd.t243 7.64824
R12043 gnd.n3469 gnd.n2083 7.64824
R12044 gnd.n3541 gnd.n2047 7.64824
R12045 gnd.t37 gnd.n2042 7.64824
R12046 gnd.n3561 gnd.t272 7.64824
R12047 gnd.n3597 gnd.n1992 7.64824
R12048 gnd.n3706 gnd.n1955 7.64824
R12049 gnd.n5278 gnd.n5277 7.53171
R12050 gnd.t305 gnd.n5379 7.32958
R12051 gnd.n1486 gnd.n1485 7.30353
R12052 gnd.n4009 gnd.n4008 7.30353
R12053 gnd.n5688 gnd.n5687 7.01093
R12054 gnd.n5698 gnd.n5408 7.01093
R12055 gnd.n5697 gnd.n5411 7.01093
R12056 gnd.n5706 gnd.n5402 7.01093
R12057 gnd.n5710 gnd.n5709 7.01093
R12058 gnd.n5728 gnd.n5387 7.01093
R12059 gnd.n5727 gnd.n5390 7.01093
R12060 gnd.n5738 gnd.n5379 7.01093
R12061 gnd.n5380 gnd.n5368 7.01093
R12062 gnd.n5751 gnd.n5369 7.01093
R12063 gnd.n5762 gnd.n5361 7.01093
R12064 gnd.n5761 gnd.n5352 7.01093
R12065 gnd.n5354 gnd.n5336 7.01093
R12066 gnd.n5798 gnd.n5337 7.01093
R12067 gnd.n5787 gnd.n5786 7.01093
R12068 gnd.n5823 gnd.n5328 7.01093
R12069 gnd.n5834 gnd.n5833 7.01093
R12070 gnd.n5321 gnd.n5313 7.01093
R12071 gnd.n5863 gnd.n5301 7.01093
R12072 gnd.n5862 gnd.n5304 7.01093
R12073 gnd.n5873 gnd.n5293 7.01093
R12074 gnd.n5294 gnd.n5282 7.01093
R12075 gnd.n5884 gnd.n5283 7.01093
R12076 gnd.n5908 gnd.n5210 7.01093
R12077 gnd.n5907 gnd.n5201 7.01093
R12078 gnd.n5203 gnd.n5194 7.01093
R12079 gnd.n5930 gnd.n5929 7.01093
R12080 gnd.n5947 gnd.n5182 7.01093
R12081 gnd.n5946 gnd.n5185 7.01093
R12082 gnd.n5960 gnd.n5174 7.01093
R12083 gnd.n5175 gnd.n5164 7.01093
R12084 gnd.n5970 gnd.n5166 7.01093
R12085 gnd.n6003 gnd.n6002 7.01093
R12086 gnd.n6019 gnd.n6018 7.01093
R12087 gnd.n5145 gnd.n968 7.01093
R12088 gnd.n6462 gnd.n970 7.01093
R12089 gnd.n5983 gnd.n979 7.01093
R12090 gnd.n6456 gnd.n6455 7.01093
R12091 gnd.n6449 gnd.n990 7.01093
R12092 gnd.n6448 gnd.n993 7.01093
R12093 gnd.n6327 gnd.n1002 7.01093
R12094 gnd.n6442 gnd.n6441 7.01093
R12095 gnd.n6308 gnd.n1005 7.01093
R12096 gnd.n6435 gnd.n1016 7.01093
R12097 gnd.n6434 gnd.n1019 7.01093
R12098 gnd.n6338 gnd.n1027 7.01093
R12099 gnd.n6428 gnd.n6427 7.01093
R12100 gnd.n4662 gnd.n1493 7.01093
R12101 gnd.n3391 gnd.n3390 7.01093
R12102 gnd.n3412 gnd.t288 7.01093
R12103 gnd.n3411 gnd.n2100 7.01093
R12104 gnd.n3562 gnd.n3561 7.01093
R12105 gnd.t272 gnd.n3559 7.01093
R12106 gnd.n3632 gnd.n2005 7.01093
R12107 gnd.n3988 gnd.n3987 7.01093
R12108 gnd.t148 gnd.n1883 7.01093
R12109 gnd.n5369 gnd.t324 6.69227
R12110 gnd.n5929 gnd.t276 6.69227
R12111 gnd.t322 gnd.n6319 6.69227
R12112 gnd.n4898 gnd.t18 6.69227
R12113 gnd.n3002 gnd.t61 6.69227
R12114 gnd.n1957 gnd.t285 6.69227
R12115 gnd.n4355 gnd.t44 6.69227
R12116 gnd.n7392 gnd.t38 6.69227
R12117 gnd.n4139 gnd.n4138 6.5566
R12118 gnd.n2194 gnd.n2193 6.5566
R12119 gnd.n4674 gnd.n4670 6.5566
R12120 gnd.n4017 gnd.n4016 6.5566
R12121 gnd.n6463 gnd.n6462 6.37362
R12122 gnd.n3227 gnd.t121 6.37362
R12123 gnd.n3280 gnd.n2168 6.37362
R12124 gnd.n3335 gnd.n2159 6.37362
R12125 gnd.n3419 gnd.t36 6.37362
R12126 gnd.n3477 gnd.n2077 6.37362
R12127 gnd.n3489 gnd.n2064 6.37362
R12128 gnd.n3610 gnd.t34 6.37362
R12129 gnd.n3658 gnd.n1988 6.37362
R12130 gnd.n3581 gnd.n1975 6.37362
R12131 gnd.t100 gnd.n1962 6.37362
R12132 gnd.n2549 gnd.n2517 6.20656
R12133 gnd.n3922 gnd.n3765 6.20656
R12134 gnd.n5822 gnd.t351 6.05496
R12135 gnd.n5821 gnd.t325 6.05496
R12136 gnd.t235 gnd.n5294 6.05496
R12137 gnd.t328 gnd.n5158 6.05496
R12138 gnd.n2925 gnd.t48 6.05496
R12139 gnd.t210 gnd.t128 6.05496
R12140 gnd.t287 gnd.t268 6.05496
R12141 gnd.t223 gnd.t300 6.05496
R12142 gnd.n4374 gnd.t20 6.05496
R12143 gnd.n6292 gnd.n6262 5.81868
R12144 gnd.n6260 gnd.n6230 5.81868
R12145 gnd.n6228 gnd.n6198 5.81868
R12146 gnd.n6197 gnd.n6167 5.81868
R12147 gnd.n6165 gnd.n6135 5.81868
R12148 gnd.n6133 gnd.n6103 5.81868
R12149 gnd.n6101 gnd.n6071 5.81868
R12150 gnd.n6070 gnd.n6040 5.81868
R12151 gnd.n2125 gnd.n2113 5.73631
R12152 gnd.n3402 gnd.n2106 5.73631
R12153 gnd.t243 gnd.n3458 5.73631
R12154 gnd.n2048 gnd.t37 5.73631
R12155 gnd.n3499 gnd.n3498 5.73631
R12156 gnd.n3569 gnd.n2023 5.73631
R12157 gnd.n4148 gnd.n1842 5.62001
R12158 gnd.n4736 gnd.n1429 5.62001
R12159 gnd.n4736 gnd.n1430 5.62001
R12160 gnd.n4148 gnd.n1843 5.62001
R12161 gnd.n5506 gnd.n5505 5.4308
R12162 gnd.n5125 gnd.n5123 5.4308
R12163 gnd.n5283 gnd.t318 5.41765
R12164 gnd.t306 gnd.n5918 5.41765
R12165 gnd.n6004 gnd.t358 5.41765
R12166 gnd.n2898 gnd.t24 5.41765
R12167 gnd.t40 gnd.n3350 5.41765
R12168 gnd.n3589 gnd.t348 5.41765
R12169 gnd.n4471 gnd.t8 5.41765
R12170 gnd.n2766 gnd.n1194 5.09899
R12171 gnd.n4892 gnd.n1197 5.09899
R12172 gnd.n2772 gnd.n1204 5.09899
R12173 gnd.n4886 gnd.n1207 5.09899
R12174 gnd.n2819 gnd.n2818 5.09899
R12175 gnd.n4880 gnd.n1217 5.09899
R12176 gnd.n2825 gnd.n1224 5.09899
R12177 gnd.n4874 gnd.n1227 5.09899
R12178 gnd.n2834 gnd.n1235 5.09899
R12179 gnd.n4868 gnd.n1238 5.09899
R12180 gnd.n2841 gnd.n1245 5.09899
R12181 gnd.n4862 gnd.n1248 5.09899
R12182 gnd.n2861 gnd.n2640 5.09899
R12183 gnd.n2860 gnd.n2643 5.09899
R12184 gnd.n2852 gnd.n2625 5.09899
R12185 gnd.n2884 gnd.n2627 5.09899
R12186 gnd.n2889 gnd.n2621 5.09899
R12187 gnd.n2878 gnd.n2877 5.09899
R12188 gnd.n2898 gnd.n2611 5.09899
R12189 gnd.n2903 gnd.n2597 5.09899
R12190 gnd.n2940 gnd.n2939 5.09899
R12191 gnd.n4854 gnd.n1265 5.09899
R12192 gnd.n2910 gnd.n1274 5.09899
R12193 gnd.n2916 gnd.n1283 5.09899
R12194 gnd.n4842 gnd.n1286 5.09899
R12195 gnd.n2925 gnd.n1293 5.09899
R12196 gnd.n4836 gnd.n1296 5.09899
R12197 gnd.n2979 gnd.n2978 5.09899
R12198 gnd.n4830 gnd.n1306 5.09899
R12199 gnd.n2987 gnd.n1313 5.09899
R12200 gnd.n2994 gnd.n1323 5.09899
R12201 gnd.n4818 gnd.n1326 5.09899
R12202 gnd.n3002 gnd.n1333 5.09899
R12203 gnd.n4812 gnd.n1336 5.09899
R12204 gnd.n3037 gnd.n3036 5.09899
R12205 gnd.n4806 gnd.n1346 5.09899
R12206 gnd.n3009 gnd.n1353 5.09899
R12207 gnd.n4800 gnd.n1356 5.09899
R12208 gnd.n3014 gnd.n1364 5.09899
R12209 gnd.n4794 gnd.n1367 5.09899
R12210 gnd.n3021 gnd.n1373 5.09899
R12211 gnd.n4788 gnd.n1376 5.09899
R12212 gnd.n3257 gnd.t121 5.09899
R12213 gnd.t158 gnd.n2163 5.09899
R12214 gnd.n3343 gnd.n2163 5.09899
R12215 gnd.n3517 gnd.n2068 5.09899
R12216 gnd.n3525 gnd.n2061 5.09899
R12217 gnd.n3684 gnd.n1972 5.09899
R12218 gnd.n4547 gnd.n4546 5.09899
R12219 gnd.n3754 gnd.n1602 5.09899
R12220 gnd.n4540 gnd.n1611 5.09899
R12221 gnd.n4333 gnd.n1614 5.09899
R12222 gnd.n4534 gnd.n1623 5.09899
R12223 gnd.n4341 gnd.n1626 5.09899
R12224 gnd.n4528 gnd.n1634 5.09899
R12225 gnd.n4347 gnd.n1800 5.09899
R12226 gnd.n4522 gnd.n1643 5.09899
R12227 gnd.n4355 gnd.n1646 5.09899
R12228 gnd.n4516 gnd.n1654 5.09899
R12229 gnd.n4391 gnd.n1657 5.09899
R12230 gnd.n4362 gnd.n1666 5.09899
R12231 gnd.n4504 gnd.n1674 5.09899
R12232 gnd.n4367 gnd.n4366 5.09899
R12233 gnd.n4498 gnd.n1683 5.09899
R12234 gnd.n4374 gnd.n1686 5.09899
R12235 gnd.n4492 gnd.n1694 5.09899
R12236 gnd.n4415 gnd.n1697 5.09899
R12237 gnd.n4445 gnd.n1706 5.09899
R12238 gnd.n4480 gnd.n1712 5.09899
R12239 gnd.n4457 gnd.n4456 5.09899
R12240 gnd.n4474 gnd.n1721 5.09899
R12241 gnd.n4471 gnd.n1724 5.09899
R12242 gnd.n4470 gnd.n1732 5.09899
R12243 gnd.n4435 gnd.n4423 5.09899
R12244 gnd.n7631 gnd.n85 5.09899
R12245 gnd.n381 gnd.n87 5.09899
R12246 gnd.n7328 gnd.n7323 5.09899
R12247 gnd.n7623 gnd.n102 5.09899
R12248 gnd.n7334 gnd.n105 5.09899
R12249 gnd.n7617 gnd.n114 5.09899
R12250 gnd.n7342 gnd.n374 5.09899
R12251 gnd.n7611 gnd.n123 5.09899
R12252 gnd.n7348 gnd.n371 5.09899
R12253 gnd.n7605 gnd.n132 5.09899
R12254 gnd.n7356 gnd.n135 5.09899
R12255 gnd.n7599 gnd.n143 5.09899
R12256 gnd.n7362 gnd.n146 5.09899
R12257 gnd.n7593 gnd.n153 5.09899
R12258 gnd.n7371 gnd.n362 5.09899
R12259 gnd.n7587 gnd.n163 5.09899
R12260 gnd.n6290 gnd.n6289 5.04292
R12261 gnd.n6258 gnd.n6257 5.04292
R12262 gnd.n6226 gnd.n6225 5.04292
R12263 gnd.n6195 gnd.n6194 5.04292
R12264 gnd.n6163 gnd.n6162 5.04292
R12265 gnd.n6131 gnd.n6130 5.04292
R12266 gnd.n6099 gnd.n6098 5.04292
R12267 gnd.n6068 gnd.n6067 5.04292
R12268 gnd.t326 gnd.n5844 4.78034
R12269 gnd.n5960 gnd.t293 4.78034
R12270 gnd.n2841 gnd.t4 4.78034
R12271 gnd.n4848 gnd.t12 4.78034
R12272 gnd.n3184 gnd.t262 4.78034
R12273 gnd.n3954 gnd.t50 4.78034
R12274 gnd.n4486 gnd.t42 4.78034
R12275 gnd.n7617 gnd.t46 4.78034
R12276 gnd.n5818 gnd.n5817 4.74817
R12277 gnd.n5813 gnd.n5812 4.74817
R12278 gnd.n5809 gnd.n5808 4.74817
R12279 gnd.n5805 gnd.n5280 4.74817
R12280 gnd.n5817 gnd.n5816 4.74817
R12281 gnd.n5815 gnd.n5813 4.74817
R12282 gnd.n5811 gnd.n5809 4.74817
R12283 gnd.n5807 gnd.n5805 4.74817
R12284 gnd.n4482 gnd.n98 4.74817
R12285 gnd.n1726 gnd.n96 4.74817
R12286 gnd.n7629 gnd.n91 4.74817
R12287 gnd.n7627 gnd.n92 4.74817
R12288 gnd.n1710 gnd.n98 4.74817
R12289 gnd.n1728 gnd.n96 4.74817
R12290 gnd.n1725 gnd.n91 4.74817
R12291 gnd.n7628 gnd.n7627 4.74817
R12292 gnd.n2864 gnd.n2863 4.74817
R12293 gnd.n2869 gnd.n2636 4.74817
R12294 gnd.n2875 gnd.n2871 4.74817
R12295 gnd.n2873 gnd.n2872 4.74817
R12296 gnd.n2595 gnd.n2593 4.74817
R12297 gnd.n4409 gnd.n1735 4.74817
R12298 gnd.n4462 gnd.n4461 4.74817
R12299 gnd.n4467 gnd.n4466 4.74817
R12300 gnd.n4463 gnd.n384 4.74817
R12301 gnd.n7320 gnd.n7319 4.74817
R12302 gnd.n4410 gnd.n4409 4.74817
R12303 gnd.n4461 gnd.n4460 4.74817
R12304 gnd.n4468 gnd.n4467 4.74817
R12305 gnd.n4465 gnd.n4463 4.74817
R12306 gnd.n7321 gnd.n7320 4.74817
R12307 gnd.n4859 gnd.n4858 4.74817
R12308 gnd.n2887 gnd.n1257 4.74817
R12309 gnd.n2900 gnd.n1256 4.74817
R12310 gnd.n1259 gnd.n1255 4.74817
R12311 gnd.n4858 gnd.n1252 4.74817
R12312 gnd.n2624 gnd.n1257 4.74817
R12313 gnd.n2886 gnd.n1256 4.74817
R12314 gnd.n2901 gnd.n1255 4.74817
R12315 gnd.n2865 gnd.n2864 4.74817
R12316 gnd.n2866 gnd.n2636 4.74817
R12317 gnd.n2871 gnd.n2870 4.74817
R12318 gnd.n2874 gnd.n2873 4.74817
R12319 gnd.n2596 gnd.n2595 4.74817
R12320 gnd.n5277 gnd.n5276 4.74296
R12321 gnd.n78 gnd.n77 4.74296
R12322 gnd.n5245 gnd.n5244 4.7074
R12323 gnd.n5261 gnd.n5260 4.7074
R12324 gnd.n46 gnd.n45 4.7074
R12325 gnd.n62 gnd.n61 4.7074
R12326 gnd.n5277 gnd.n5261 4.65959
R12327 gnd.n78 gnd.n62 4.65959
R12328 gnd.n4239 gnd.n4149 4.6132
R12329 gnd.n4737 gnd.n1428 4.6132
R12330 gnd.n3257 gnd.n3256 4.46168
R12331 gnd.t78 gnd.n1493 4.46168
R12332 gnd.n3263 gnd.t78 4.46168
R12333 gnd.n3388 gnd.t266 4.46168
R12334 gnd.n3399 gnd.n3397 4.46168
R12335 gnd.n3428 gnd.n2108 4.46168
R12336 gnd.n3576 gnd.n2028 4.46168
R12337 gnd.n3620 gnd.n2015 4.46168
R12338 gnd.t314 gnd.n3618 4.46168
R12339 gnd.n4078 gnd.n1883 4.46168
R12340 gnd.n4005 gnd.n3992 4.46111
R12341 gnd.n6275 gnd.n6271 4.38594
R12342 gnd.n6243 gnd.n6239 4.38594
R12343 gnd.n6211 gnd.n6207 4.38594
R12344 gnd.n6180 gnd.n6176 4.38594
R12345 gnd.n6148 gnd.n6144 4.38594
R12346 gnd.n6116 gnd.n6112 4.38594
R12347 gnd.n6084 gnd.n6080 4.38594
R12348 gnd.n6053 gnd.n6049 4.38594
R12349 gnd.n6286 gnd.n6264 4.26717
R12350 gnd.n6254 gnd.n6232 4.26717
R12351 gnd.n6222 gnd.n6200 4.26717
R12352 gnd.n6191 gnd.n6169 4.26717
R12353 gnd.n6159 gnd.n6137 4.26717
R12354 gnd.n6127 gnd.n6105 4.26717
R12355 gnd.n6095 gnd.n6073 4.26717
R12356 gnd.n6064 gnd.n6042 4.26717
R12357 gnd.t344 gnd.n5775 4.14303
R12358 gnd.t295 gnd.n970 4.14303
R12359 gnd.n2772 gnd.t200 4.14303
R12360 gnd.n4824 gnd.t69 4.14303
R12361 gnd.t111 gnd.n1367 4.14303
R12362 gnd.t89 gnd.n1611 4.14303
R12363 gnd.n4510 gnd.t14 4.14303
R12364 gnd.n7593 gnd.t241 4.14303
R12365 gnd.n6294 gnd.n6293 4.08274
R12366 gnd.n4138 gnd.n4137 4.05904
R12367 gnd.n2195 gnd.n2194 4.05904
R12368 gnd.n4677 gnd.n4670 4.05904
R12369 gnd.n4018 gnd.n4017 4.05904
R12370 gnd.n15 gnd.n7 3.99943
R12371 gnd.n4733 gnd.t10 3.82437
R12372 gnd.n3299 gnd.n2176 3.82437
R12373 gnd.n3341 gnd.t33 3.82437
R12374 gnd.n3360 gnd.n3359 3.82437
R12375 gnd.n3448 gnd.n2097 3.82437
R12376 gnd.n3450 gnd.t287 3.82437
R12377 gnd.n3491 gnd.t223 3.82437
R12378 gnd.n3534 gnd.n3533 3.82437
R12379 gnd.n3649 gnd.n1986 3.82437
R12380 gnd.n3675 gnd.t65 3.82437
R12381 gnd.n3699 gnd.n3698 3.82437
R12382 gnd.n4145 gnd.t356 3.82437
R12383 gnd.n5279 gnd.n5278 3.81325
R12384 gnd.n5261 gnd.n5245 3.72967
R12385 gnd.n62 gnd.n46 3.72967
R12386 gnd.n6294 gnd.n6166 3.70378
R12387 gnd.n15 gnd.n14 3.60163
R12388 gnd.n6285 gnd.n6266 3.49141
R12389 gnd.n6253 gnd.n6234 3.49141
R12390 gnd.n6221 gnd.n6202 3.49141
R12391 gnd.n6190 gnd.n6171 3.49141
R12392 gnd.n6158 gnd.n6139 3.49141
R12393 gnd.n6126 gnd.n6107 3.49141
R12394 gnd.n6094 gnd.n6075 3.49141
R12395 gnd.n6063 gnd.n6044 3.49141
R12396 gnd.n4220 gnd.n4219 3.29747
R12397 gnd.n4219 gnd.n4157 3.29747
R12398 gnd.n7522 gnd.n7519 3.29747
R12399 gnd.n7523 gnd.n7522 3.29747
R12400 gnd.n5011 gnd.n5010 3.29747
R12401 gnd.n5010 gnd.n5009 3.29747
R12402 gnd.n4753 gnd.n4752 3.29747
R12403 gnd.n4752 gnd.n4751 3.29747
R12404 gnd.n3264 gnd.n2183 3.18706
R12405 gnd.n3377 gnd.n3376 3.18706
R12406 gnd.n3439 gnd.n3438 3.18706
R12407 gnd.n3549 gnd.n3548 3.18706
R12408 gnd.n3630 gnd.n3629 3.18706
R12409 gnd.n3581 gnd.t100 3.18706
R12410 gnd.n3716 gnd.n3714 3.18706
R12411 gnd.n5776 gnd.t344 2.8684
R12412 gnd.n2260 gnd.t10 2.8684
R12413 gnd.n5262 gnd.t76 2.82907
R12414 gnd.n5262 gnd.t267 2.82907
R12415 gnd.n5264 gnd.t55 2.82907
R12416 gnd.n5264 gnd.t218 2.82907
R12417 gnd.n5266 gnd.t291 2.82907
R12418 gnd.n5266 gnd.t13 2.82907
R12419 gnd.n5268 gnd.t313 2.82907
R12420 gnd.n5268 gnd.t292 2.82907
R12421 gnd.n5270 gnd.t5 2.82907
R12422 gnd.n5270 gnd.t323 2.82907
R12423 gnd.n5272 gnd.t57 2.82907
R12424 gnd.n5272 gnd.t7 2.82907
R12425 gnd.n5274 gnd.t198 2.82907
R12426 gnd.n5274 gnd.t201 2.82907
R12427 gnd.n5215 gnd.t250 2.82907
R12428 gnd.n5215 gnd.t308 2.82907
R12429 gnd.n5217 gnd.t339 2.82907
R12430 gnd.n5217 gnd.t247 2.82907
R12431 gnd.n5219 gnd.t333 2.82907
R12432 gnd.n5219 gnd.t237 2.82907
R12433 gnd.n5221 gnd.t275 2.82907
R12434 gnd.n5221 gnd.t73 2.82907
R12435 gnd.n5223 gnd.t311 2.82907
R12436 gnd.n5223 gnd.t342 2.82907
R12437 gnd.n5225 gnd.t203 2.82907
R12438 gnd.n5225 gnd.t317 2.82907
R12439 gnd.n5227 gnd.t68 2.82907
R12440 gnd.n5227 gnd.t331 2.82907
R12441 gnd.n5230 gnd.t70 2.82907
R12442 gnd.n5230 gnd.t62 2.82907
R12443 gnd.n5232 gnd.t49 2.82907
R12444 gnd.n5232 gnd.t207 2.82907
R12445 gnd.n5234 gnd.t278 2.82907
R12446 gnd.n5234 gnd.t199 2.82907
R12447 gnd.n5236 gnd.t240 2.82907
R12448 gnd.n5236 gnd.t25 2.82907
R12449 gnd.n5238 gnd.t279 2.82907
R12450 gnd.n5238 gnd.t283 2.82907
R12451 gnd.n5240 gnd.t216 2.82907
R12452 gnd.n5240 gnd.t284 2.82907
R12453 gnd.n5242 gnd.t251 2.82907
R12454 gnd.n5242 gnd.t289 2.82907
R12455 gnd.n5246 gnd.t310 2.82907
R12456 gnd.n5246 gnd.t227 2.82907
R12457 gnd.n5248 gnd.t281 2.82907
R12458 gnd.n5248 gnd.t217 2.82907
R12459 gnd.n5250 gnd.t64 2.82907
R12460 gnd.n5250 gnd.t212 2.82907
R12461 gnd.n5252 gnd.t234 2.82907
R12462 gnd.n5252 gnd.t52 2.82907
R12463 gnd.n5254 gnd.t27 2.82907
R12464 gnd.n5254 gnd.t249 2.82907
R12465 gnd.n5256 gnd.t226 2.82907
R12466 gnd.n5256 gnd.t327 2.82907
R12467 gnd.n5258 gnd.t19 2.82907
R12468 gnd.n5258 gnd.t246 2.82907
R12469 gnd.n75 gnd.t336 2.82907
R12470 gnd.n75 gnd.t225 2.82907
R12471 gnd.n73 gnd.t260 2.82907
R12472 gnd.n73 gnd.t329 2.82907
R12473 gnd.n71 gnd.t238 2.82907
R12474 gnd.n71 gnd.t60 2.82907
R12475 gnd.n69 gnd.t28 2.82907
R12476 gnd.n69 gnd.t290 2.82907
R12477 gnd.n67 gnd.t67 2.82907
R12478 gnd.n67 gnd.t1 2.82907
R12479 gnd.n65 gnd.t280 2.82907
R12480 gnd.n65 gnd.t350 2.82907
R12481 gnd.n63 gnd.t45 2.82907
R12482 gnd.n63 gnd.t219 2.82907
R12483 gnd.n28 gnd.t304 2.82907
R12484 gnd.n28 gnd.t39 2.82907
R12485 gnd.n26 gnd.t299 2.82907
R12486 gnd.n26 gnd.t59 2.82907
R12487 gnd.n24 gnd.t30 2.82907
R12488 gnd.n24 gnd.t47 2.82907
R12489 gnd.n22 gnd.t75 2.82907
R12490 gnd.n22 gnd.t23 2.82907
R12491 gnd.n20 gnd.t43 2.82907
R12492 gnd.n20 gnd.t346 2.82907
R12493 gnd.n18 gnd.t245 2.82907
R12494 gnd.n18 gnd.t337 2.82907
R12495 gnd.n16 gnd.t202 2.82907
R12496 gnd.n16 gnd.t15 2.82907
R12497 gnd.n43 gnd.t343 2.82907
R12498 gnd.n43 gnd.t230 2.82907
R12499 gnd.n41 gnd.t274 2.82907
R12500 gnd.n41 gnd.t334 2.82907
R12501 gnd.n39 gnd.t338 2.82907
R12502 gnd.n39 gnd.t335 2.82907
R12503 gnd.n37 gnd.t332 2.82907
R12504 gnd.n37 gnd.t239 2.82907
R12505 gnd.n35 gnd.t347 2.82907
R12506 gnd.n35 gnd.t204 2.82907
R12507 gnd.n33 gnd.t72 2.82907
R12508 gnd.n33 gnd.t74 2.82907
R12509 gnd.n31 gnd.t330 2.82907
R12510 gnd.n31 gnd.t244 2.82907
R12511 gnd.n59 gnd.t242 2.82907
R12512 gnd.n59 gnd.t320 2.82907
R12513 gnd.n57 gnd.t273 2.82907
R12514 gnd.n57 gnd.t228 2.82907
R12515 gnd.n55 gnd.t254 2.82907
R12516 gnd.n55 gnd.t312 2.82907
R12517 gnd.n53 gnd.t9 2.82907
R12518 gnd.n53 gnd.t341 2.82907
R12519 gnd.n51 gnd.t353 2.82907
R12520 gnd.n51 gnd.t340 2.82907
R12521 gnd.n49 gnd.t197 2.82907
R12522 gnd.n49 gnd.t21 2.82907
R12523 gnd.n47 gnd.t282 2.82907
R12524 gnd.n47 gnd.t296 2.82907
R12525 gnd.n6282 gnd.n6281 2.71565
R12526 gnd.n6250 gnd.n6249 2.71565
R12527 gnd.n6218 gnd.n6217 2.71565
R12528 gnd.n6187 gnd.n6186 2.71565
R12529 gnd.n6155 gnd.n6154 2.71565
R12530 gnd.n6123 gnd.n6122 2.71565
R12531 gnd.n6091 gnd.n6090 2.71565
R12532 gnd.n6060 gnd.n6059 2.71565
R12533 gnd.n3289 gnd.n3288 2.54975
R12534 gnd.n3378 gnd.n2139 2.54975
R12535 gnd.n3378 gnd.t315 2.54975
R12536 gnd.n3459 gnd.n2090 2.54975
R12537 gnd.n3550 gnd.n2042 2.54975
R12538 gnd.n3639 gnd.t35 2.54975
R12539 gnd.n3639 gnd.n3638 2.54975
R12540 gnd.n1958 gnd.n1951 2.54975
R12541 gnd.n5817 gnd.n5279 2.27742
R12542 gnd.n5813 gnd.n5279 2.27742
R12543 gnd.n5809 gnd.n5279 2.27742
R12544 gnd.n5805 gnd.n5279 2.27742
R12545 gnd.n7626 gnd.n98 2.27742
R12546 gnd.n7626 gnd.n96 2.27742
R12547 gnd.n7626 gnd.n91 2.27742
R12548 gnd.n7627 gnd.n7626 2.27742
R12549 gnd.n4409 gnd.n95 2.27742
R12550 gnd.n4461 gnd.n95 2.27742
R12551 gnd.n4467 gnd.n95 2.27742
R12552 gnd.n4463 gnd.n95 2.27742
R12553 gnd.n7320 gnd.n95 2.27742
R12554 gnd.n4858 gnd.n4857 2.27742
R12555 gnd.n4857 gnd.n1257 2.27742
R12556 gnd.n4857 gnd.n1256 2.27742
R12557 gnd.n4857 gnd.n1255 2.27742
R12558 gnd.n2864 gnd.n1254 2.27742
R12559 gnd.n2636 gnd.n1254 2.27742
R12560 gnd.n2871 gnd.n1254 2.27742
R12561 gnd.n2873 gnd.n1254 2.27742
R12562 gnd.n2595 gnd.n1254 2.27742
R12563 gnd.t151 gnd.n5697 2.23109
R12564 gnd.n5845 gnd.t326 2.23109
R12565 gnd.t208 gnd.n2108 2.23109
R12566 gnd.t268 gnd.n3448 2.23109
R12567 gnd.n3534 gnd.t300 2.23109
R12568 gnd.t231 gnd.n2028 2.23109
R12569 gnd.n6278 gnd.n6268 1.93989
R12570 gnd.n6246 gnd.n6236 1.93989
R12571 gnd.n6214 gnd.n6204 1.93989
R12572 gnd.n6183 gnd.n6173 1.93989
R12573 gnd.n6151 gnd.n6141 1.93989
R12574 gnd.n6119 gnd.n6109 1.93989
R12575 gnd.n6087 gnd.n6077 1.93989
R12576 gnd.n6056 gnd.n6046 1.93989
R12577 gnd.n3300 gnd.n2175 1.91244
R12578 gnd.t195 gnd.n2176 1.91244
R12579 gnd.n3309 gnd.n3307 1.91244
R12580 gnd.n3468 gnd.n2085 1.91244
R12581 gnd.n2055 gnd.n2054 1.91244
R12582 gnd.n3652 gnd.n3651 1.91244
R12583 gnd.n1965 gnd.n1964 1.91244
R12584 gnd.n3979 gnd.t186 1.91244
R12585 gnd.n5710 gnd.t252 1.59378
R12586 gnd.n5919 gnd.t306 1.59378
R12587 gnd.n5993 gnd.t358 1.59378
R12588 gnd.t354 gnd.n2130 1.59378
R12589 gnd.n3631 gnd.t264 1.59378
R12590 gnd.n4663 gnd.n1490 1.27512
R12591 gnd.n3274 gnd.t107 1.27512
R12592 gnd.n3351 gnd.t33 1.27512
R12593 gnd.n3389 gnd.n3388 1.27512
R12594 gnd.n3412 gnd.n2117 1.27512
R12595 gnd.n3559 gnd.n3558 1.27512
R12596 gnd.n3618 gnd.n2016 1.27512
R12597 gnd.n3588 gnd.t65 1.27512
R12598 gnd.t97 gnd.n1955 1.27512
R12599 gnd.n3706 gnd.t131 1.27512
R12600 gnd.n3986 gnd.n3985 1.27512
R12601 gnd.n5507 gnd.n5506 1.16414
R12602 gnd.n6353 gnd.n5123 1.16414
R12603 gnd.n6277 gnd.n6270 1.16414
R12604 gnd.n6245 gnd.n6238 1.16414
R12605 gnd.n6213 gnd.n6206 1.16414
R12606 gnd.n6182 gnd.n6175 1.16414
R12607 gnd.n6150 gnd.n6143 1.16414
R12608 gnd.n6118 gnd.n6111 1.16414
R12609 gnd.n6086 gnd.n6079 1.16414
R12610 gnd.n6055 gnd.n6048 1.16414
R12611 gnd.n4149 gnd.n1841 0.970197
R12612 gnd.n4737 gnd.n1425 0.970197
R12613 gnd.n6261 gnd.n6229 0.962709
R12614 gnd.n6293 gnd.n6261 0.962709
R12615 gnd.n6134 gnd.n6102 0.962709
R12616 gnd.n6166 gnd.n6134 0.962709
R12617 gnd.t351 gnd.n5821 0.956468
R12618 gnd.n5165 gnd.t328 0.956468
R12619 gnd.t6 gnd.n1227 0.956468
R12620 gnd.n2580 gnd.t69 0.956468
R12621 gnd.t255 gnd.n2277 0.956468
R12622 gnd.t186 gnd.t356 0.956468
R12623 gnd.n3967 gnd.t31 0.956468
R12624 gnd.n4392 gnd.t14 0.956468
R12625 gnd.n371 gnd.t259 0.956468
R12626 gnd.n2 gnd.n1 0.672012
R12627 gnd.n3 gnd.n2 0.672012
R12628 gnd.n4 gnd.n3 0.672012
R12629 gnd.n5 gnd.n4 0.672012
R12630 gnd.n6 gnd.n5 0.672012
R12631 gnd.n7 gnd.n6 0.672012
R12632 gnd.n9 gnd.n8 0.672012
R12633 gnd.n10 gnd.n9 0.672012
R12634 gnd.n11 gnd.n10 0.672012
R12635 gnd.n12 gnd.n11 0.672012
R12636 gnd.n13 gnd.n12 0.672012
R12637 gnd.n14 gnd.n13 0.672012
R12638 gnd.t128 gnd.n2185 0.637812
R12639 gnd.n3330 gnd.n3329 0.637812
R12640 gnd.n3350 gnd.n3349 0.637812
R12641 gnd.n3359 gnd.t316 0.637812
R12642 gnd.n3479 gnd.n3478 0.637812
R12643 gnd.n3524 gnd.n3523 0.637812
R12644 gnd.t66 gnd.n3649 0.637812
R12645 gnd.n3590 gnd.n3589 0.637812
R12646 gnd.n3683 gnd.n3681 0.637812
R12647 gnd.n3714 gnd.t170 0.637812
R12648 gnd gnd.n0 0.59317
R12649 gnd.n5276 gnd.n5275 0.573776
R12650 gnd.n5275 gnd.n5273 0.573776
R12651 gnd.n5273 gnd.n5271 0.573776
R12652 gnd.n5271 gnd.n5269 0.573776
R12653 gnd.n5269 gnd.n5267 0.573776
R12654 gnd.n5267 gnd.n5265 0.573776
R12655 gnd.n5265 gnd.n5263 0.573776
R12656 gnd.n5229 gnd.n5228 0.573776
R12657 gnd.n5228 gnd.n5226 0.573776
R12658 gnd.n5226 gnd.n5224 0.573776
R12659 gnd.n5224 gnd.n5222 0.573776
R12660 gnd.n5222 gnd.n5220 0.573776
R12661 gnd.n5220 gnd.n5218 0.573776
R12662 gnd.n5218 gnd.n5216 0.573776
R12663 gnd.n5244 gnd.n5243 0.573776
R12664 gnd.n5243 gnd.n5241 0.573776
R12665 gnd.n5241 gnd.n5239 0.573776
R12666 gnd.n5239 gnd.n5237 0.573776
R12667 gnd.n5237 gnd.n5235 0.573776
R12668 gnd.n5235 gnd.n5233 0.573776
R12669 gnd.n5233 gnd.n5231 0.573776
R12670 gnd.n5260 gnd.n5259 0.573776
R12671 gnd.n5259 gnd.n5257 0.573776
R12672 gnd.n5257 gnd.n5255 0.573776
R12673 gnd.n5255 gnd.n5253 0.573776
R12674 gnd.n5253 gnd.n5251 0.573776
R12675 gnd.n5251 gnd.n5249 0.573776
R12676 gnd.n5249 gnd.n5247 0.573776
R12677 gnd.n66 gnd.n64 0.573776
R12678 gnd.n68 gnd.n66 0.573776
R12679 gnd.n70 gnd.n68 0.573776
R12680 gnd.n72 gnd.n70 0.573776
R12681 gnd.n74 gnd.n72 0.573776
R12682 gnd.n76 gnd.n74 0.573776
R12683 gnd.n77 gnd.n76 0.573776
R12684 gnd.n19 gnd.n17 0.573776
R12685 gnd.n21 gnd.n19 0.573776
R12686 gnd.n23 gnd.n21 0.573776
R12687 gnd.n25 gnd.n23 0.573776
R12688 gnd.n27 gnd.n25 0.573776
R12689 gnd.n29 gnd.n27 0.573776
R12690 gnd.n30 gnd.n29 0.573776
R12691 gnd.n34 gnd.n32 0.573776
R12692 gnd.n36 gnd.n34 0.573776
R12693 gnd.n38 gnd.n36 0.573776
R12694 gnd.n40 gnd.n38 0.573776
R12695 gnd.n42 gnd.n40 0.573776
R12696 gnd.n44 gnd.n42 0.573776
R12697 gnd.n45 gnd.n44 0.573776
R12698 gnd.n50 gnd.n48 0.573776
R12699 gnd.n52 gnd.n50 0.573776
R12700 gnd.n54 gnd.n52 0.573776
R12701 gnd.n56 gnd.n54 0.573776
R12702 gnd.n58 gnd.n56 0.573776
R12703 gnd.n60 gnd.n58 0.573776
R12704 gnd.n61 gnd.n60 0.573776
R12705 gnd.n7638 gnd.n7637 0.553533
R12706 gnd.n7411 gnd.n7410 0.505073
R12707 gnd.n2745 gnd.n2742 0.505073
R12708 gnd.n3931 gnd.n3930 0.489829
R12709 gnd.n3147 gnd.n2331 0.489829
R12710 gnd.n3141 gnd.n3139 0.489829
R12711 gnd.n3817 gnd.n1577 0.489829
R12712 gnd.n6343 gnd.n6342 0.486781
R12713 gnd.n5559 gnd.n5455 0.48678
R12714 gnd.n6424 gnd.n6423 0.480683
R12715 gnd.n5627 gnd.n5405 0.480683
R12716 gnd.n7554 gnd.n7553 0.470012
R12717 gnd.n4175 gnd.n1606 0.470012
R12718 gnd.n4785 gnd.n4784 0.470012
R12719 gnd.n1146 gnd.n1072 0.470012
R12720 gnd.n803 gnd.n798 0.425805
R12721 gnd.n7087 gnd.n7086 0.425805
R12722 gnd.n7300 gnd.n7299 0.425805
R12723 gnd.n2789 gnd.n2788 0.425805
R12724 gnd.n7626 gnd.n95 0.4255
R12725 gnd.n4857 gnd.n1254 0.4255
R12726 gnd.n3084 gnd.n2517 0.388379
R12727 gnd.n6274 gnd.n6273 0.388379
R12728 gnd.n6242 gnd.n6241 0.388379
R12729 gnd.n6210 gnd.n6209 0.388379
R12730 gnd.n6179 gnd.n6178 0.388379
R12731 gnd.n6147 gnd.n6146 0.388379
R12732 gnd.n6115 gnd.n6114 0.388379
R12733 gnd.n6083 gnd.n6082 0.388379
R12734 gnd.n6052 gnd.n6051 0.388379
R12735 gnd.n3908 gnd.n3765 0.388379
R12736 gnd.n7638 gnd.n15 0.374463
R12737 gnd.n6320 gnd.t322 0.319156
R12738 gnd.n2627 gnd.t233 0.319156
R12739 gnd.n2915 gnd.t12 0.319156
R12740 gnd.n3154 gnd.t141 0.319156
R12741 gnd.t107 gnd.t210 0.319156
R12742 gnd.t285 gnd.t131 0.319156
R12743 gnd.t124 gnd.n3941 0.319156
R12744 gnd.n4414 gnd.t42 0.319156
R12745 gnd.t22 gnd.n85 0.319156
R12746 gnd.n5553 gnd.n5552 0.311721
R12747 gnd gnd.n7638 0.295112
R12748 gnd.n7444 gnd.n7443 0.293183
R12749 gnd.n4927 gnd.n1136 0.293183
R12750 gnd.n2575 gnd.n2527 0.27489
R12751 gnd.n3759 gnd.n3758 0.27489
R12752 gnd.n6393 gnd.n6392 0.268793
R12753 gnd.n7445 gnd.n7444 0.258122
R12754 gnd.n4325 gnd.n4324 0.258122
R12755 gnd.n2459 gnd.n2458 0.258122
R12756 gnd.n4928 gnd.n4927 0.258122
R12757 gnd.n6392 gnd.n6391 0.241354
R12758 gnd.n4240 gnd.n4239 0.229039
R12759 gnd.n4239 gnd.n1840 0.229039
R12760 gnd.n1428 gnd.n1424 0.229039
R12761 gnd.n2379 gnd.n1428 0.229039
R12762 gnd.n5682 gnd.n5423 0.206293
R12763 gnd.n5278 gnd.n0 0.169152
R12764 gnd.n6291 gnd.n6263 0.155672
R12765 gnd.n6284 gnd.n6263 0.155672
R12766 gnd.n6284 gnd.n6283 0.155672
R12767 gnd.n6283 gnd.n6267 0.155672
R12768 gnd.n6276 gnd.n6267 0.155672
R12769 gnd.n6276 gnd.n6275 0.155672
R12770 gnd.n6259 gnd.n6231 0.155672
R12771 gnd.n6252 gnd.n6231 0.155672
R12772 gnd.n6252 gnd.n6251 0.155672
R12773 gnd.n6251 gnd.n6235 0.155672
R12774 gnd.n6244 gnd.n6235 0.155672
R12775 gnd.n6244 gnd.n6243 0.155672
R12776 gnd.n6227 gnd.n6199 0.155672
R12777 gnd.n6220 gnd.n6199 0.155672
R12778 gnd.n6220 gnd.n6219 0.155672
R12779 gnd.n6219 gnd.n6203 0.155672
R12780 gnd.n6212 gnd.n6203 0.155672
R12781 gnd.n6212 gnd.n6211 0.155672
R12782 gnd.n6196 gnd.n6168 0.155672
R12783 gnd.n6189 gnd.n6168 0.155672
R12784 gnd.n6189 gnd.n6188 0.155672
R12785 gnd.n6188 gnd.n6172 0.155672
R12786 gnd.n6181 gnd.n6172 0.155672
R12787 gnd.n6181 gnd.n6180 0.155672
R12788 gnd.n6164 gnd.n6136 0.155672
R12789 gnd.n6157 gnd.n6136 0.155672
R12790 gnd.n6157 gnd.n6156 0.155672
R12791 gnd.n6156 gnd.n6140 0.155672
R12792 gnd.n6149 gnd.n6140 0.155672
R12793 gnd.n6149 gnd.n6148 0.155672
R12794 gnd.n6132 gnd.n6104 0.155672
R12795 gnd.n6125 gnd.n6104 0.155672
R12796 gnd.n6125 gnd.n6124 0.155672
R12797 gnd.n6124 gnd.n6108 0.155672
R12798 gnd.n6117 gnd.n6108 0.155672
R12799 gnd.n6117 gnd.n6116 0.155672
R12800 gnd.n6100 gnd.n6072 0.155672
R12801 gnd.n6093 gnd.n6072 0.155672
R12802 gnd.n6093 gnd.n6092 0.155672
R12803 gnd.n6092 gnd.n6076 0.155672
R12804 gnd.n6085 gnd.n6076 0.155672
R12805 gnd.n6085 gnd.n6084 0.155672
R12806 gnd.n6069 gnd.n6041 0.155672
R12807 gnd.n6062 gnd.n6041 0.155672
R12808 gnd.n6062 gnd.n6061 0.155672
R12809 gnd.n6061 gnd.n6045 0.155672
R12810 gnd.n6054 gnd.n6045 0.155672
R12811 gnd.n6054 gnd.n6053 0.155672
R12812 gnd.n6423 gnd.n5053 0.152939
R12813 gnd.n5055 gnd.n5053 0.152939
R12814 gnd.n5059 gnd.n5055 0.152939
R12815 gnd.n5060 gnd.n5059 0.152939
R12816 gnd.n5061 gnd.n5060 0.152939
R12817 gnd.n5062 gnd.n5061 0.152939
R12818 gnd.n5066 gnd.n5062 0.152939
R12819 gnd.n5067 gnd.n5066 0.152939
R12820 gnd.n5068 gnd.n5067 0.152939
R12821 gnd.n5069 gnd.n5068 0.152939
R12822 gnd.n5073 gnd.n5069 0.152939
R12823 gnd.n5074 gnd.n5073 0.152939
R12824 gnd.n5075 gnd.n5074 0.152939
R12825 gnd.n5076 gnd.n5075 0.152939
R12826 gnd.n5081 gnd.n5076 0.152939
R12827 gnd.n6393 gnd.n5081 0.152939
R12828 gnd.n5701 gnd.n5405 0.152939
R12829 gnd.n5702 gnd.n5701 0.152939
R12830 gnd.n5703 gnd.n5702 0.152939
R12831 gnd.n5703 gnd.n5384 0.152939
R12832 gnd.n5731 gnd.n5384 0.152939
R12833 gnd.n5732 gnd.n5731 0.152939
R12834 gnd.n5733 gnd.n5732 0.152939
R12835 gnd.n5734 gnd.n5733 0.152939
R12836 gnd.n5734 gnd.n5358 0.152939
R12837 gnd.n5765 gnd.n5358 0.152939
R12838 gnd.n5766 gnd.n5765 0.152939
R12839 gnd.n5767 gnd.n5766 0.152939
R12840 gnd.n5768 gnd.n5767 0.152939
R12841 gnd.n5769 gnd.n5768 0.152939
R12842 gnd.n5769 gnd.n5325 0.152939
R12843 gnd.n5826 gnd.n5325 0.152939
R12844 gnd.n5827 gnd.n5826 0.152939
R12845 gnd.n5828 gnd.n5827 0.152939
R12846 gnd.n5829 gnd.n5828 0.152939
R12847 gnd.n5829 gnd.n5298 0.152939
R12848 gnd.n5866 gnd.n5298 0.152939
R12849 gnd.n5867 gnd.n5866 0.152939
R12850 gnd.n5868 gnd.n5867 0.152939
R12851 gnd.n5869 gnd.n5868 0.152939
R12852 gnd.n5869 gnd.n5207 0.152939
R12853 gnd.n5911 gnd.n5207 0.152939
R12854 gnd.n5912 gnd.n5911 0.152939
R12855 gnd.n5913 gnd.n5912 0.152939
R12856 gnd.n5914 gnd.n5913 0.152939
R12857 gnd.n5914 gnd.n5179 0.152939
R12858 gnd.n5950 gnd.n5179 0.152939
R12859 gnd.n5951 gnd.n5950 0.152939
R12860 gnd.n5952 gnd.n5951 0.152939
R12861 gnd.n5953 gnd.n5952 0.152939
R12862 gnd.n5954 gnd.n5953 0.152939
R12863 gnd.n5954 gnd.n5149 0.152939
R12864 gnd.n6007 gnd.n5149 0.152939
R12865 gnd.n6008 gnd.n6007 0.152939
R12866 gnd.n6009 gnd.n6008 0.152939
R12867 gnd.n6010 gnd.n6009 0.152939
R12868 gnd.n6012 gnd.n6010 0.152939
R12869 gnd.n6012 gnd.n6011 0.152939
R12870 gnd.n6011 gnd.n985 0.152939
R12871 gnd.n986 gnd.n985 0.152939
R12872 gnd.n987 gnd.n986 0.152939
R12873 gnd.n1009 gnd.n987 0.152939
R12874 gnd.n1010 gnd.n1009 0.152939
R12875 gnd.n1011 gnd.n1010 0.152939
R12876 gnd.n1012 gnd.n1011 0.152939
R12877 gnd.n1013 gnd.n1012 0.152939
R12878 gnd.n5051 gnd.n1013 0.152939
R12879 gnd.n5052 gnd.n5051 0.152939
R12880 gnd.n6424 gnd.n5052 0.152939
R12881 gnd.n5628 gnd.n5627 0.152939
R12882 gnd.n5629 gnd.n5628 0.152939
R12883 gnd.n5630 gnd.n5629 0.152939
R12884 gnd.n5631 gnd.n5630 0.152939
R12885 gnd.n5632 gnd.n5631 0.152939
R12886 gnd.n5633 gnd.n5632 0.152939
R12887 gnd.n5634 gnd.n5633 0.152939
R12888 gnd.n5635 gnd.n5634 0.152939
R12889 gnd.n5636 gnd.n5635 0.152939
R12890 gnd.n5637 gnd.n5636 0.152939
R12891 gnd.n5638 gnd.n5637 0.152939
R12892 gnd.n5639 gnd.n5638 0.152939
R12893 gnd.n5640 gnd.n5639 0.152939
R12894 gnd.n5641 gnd.n5640 0.152939
R12895 gnd.n5645 gnd.n5641 0.152939
R12896 gnd.n5645 gnd.n5423 0.152939
R12897 gnd.n6391 gnd.n5083 0.152939
R12898 gnd.n5085 gnd.n5083 0.152939
R12899 gnd.n5089 gnd.n5085 0.152939
R12900 gnd.n5090 gnd.n5089 0.152939
R12901 gnd.n5091 gnd.n5090 0.152939
R12902 gnd.n5092 gnd.n5091 0.152939
R12903 gnd.n5096 gnd.n5092 0.152939
R12904 gnd.n5097 gnd.n5096 0.152939
R12905 gnd.n5098 gnd.n5097 0.152939
R12906 gnd.n5099 gnd.n5098 0.152939
R12907 gnd.n5103 gnd.n5099 0.152939
R12908 gnd.n5104 gnd.n5103 0.152939
R12909 gnd.n5105 gnd.n5104 0.152939
R12910 gnd.n5106 gnd.n5105 0.152939
R12911 gnd.n5110 gnd.n5106 0.152939
R12912 gnd.n5111 gnd.n5110 0.152939
R12913 gnd.n5112 gnd.n5111 0.152939
R12914 gnd.n5113 gnd.n5112 0.152939
R12915 gnd.n5117 gnd.n5113 0.152939
R12916 gnd.n5118 gnd.n5117 0.152939
R12917 gnd.n5119 gnd.n5118 0.152939
R12918 gnd.n5120 gnd.n5119 0.152939
R12919 gnd.n5127 gnd.n5120 0.152939
R12920 gnd.n5128 gnd.n5127 0.152939
R12921 gnd.n5129 gnd.n5128 0.152939
R12922 gnd.n6343 gnd.n5129 0.152939
R12923 gnd.n5888 gnd.n5887 0.152939
R12924 gnd.n5889 gnd.n5888 0.152939
R12925 gnd.n5890 gnd.n5889 0.152939
R12926 gnd.n5891 gnd.n5890 0.152939
R12927 gnd.n5892 gnd.n5891 0.152939
R12928 gnd.n5893 gnd.n5892 0.152939
R12929 gnd.n5894 gnd.n5893 0.152939
R12930 gnd.n5895 gnd.n5894 0.152939
R12931 gnd.n5895 gnd.n5161 0.152939
R12932 gnd.n5973 gnd.n5161 0.152939
R12933 gnd.n5974 gnd.n5973 0.152939
R12934 gnd.n5975 gnd.n5974 0.152939
R12935 gnd.n5976 gnd.n5975 0.152939
R12936 gnd.n5977 gnd.n5976 0.152939
R12937 gnd.n5978 gnd.n5977 0.152939
R12938 gnd.n5979 gnd.n5978 0.152939
R12939 gnd.n5980 gnd.n5979 0.152939
R12940 gnd.n5981 gnd.n5980 0.152939
R12941 gnd.n5981 gnd.n5134 0.152939
R12942 gnd.n6324 gnd.n5134 0.152939
R12943 gnd.n6325 gnd.n6324 0.152939
R12944 gnd.n6326 gnd.n6325 0.152939
R12945 gnd.n6326 gnd.n5132 0.152939
R12946 gnd.n6334 gnd.n5132 0.152939
R12947 gnd.n6335 gnd.n6334 0.152939
R12948 gnd.n6336 gnd.n6335 0.152939
R12949 gnd.n6336 gnd.n5130 0.152939
R12950 gnd.n6342 gnd.n5130 0.152939
R12951 gnd.n5560 gnd.n5559 0.152939
R12952 gnd.n5561 gnd.n5560 0.152939
R12953 gnd.n5561 gnd.n5443 0.152939
R12954 gnd.n5575 gnd.n5443 0.152939
R12955 gnd.n5576 gnd.n5575 0.152939
R12956 gnd.n5577 gnd.n5576 0.152939
R12957 gnd.n5577 gnd.n5430 0.152939
R12958 gnd.n5591 gnd.n5430 0.152939
R12959 gnd.n5592 gnd.n5591 0.152939
R12960 gnd.n5593 gnd.n5592 0.152939
R12961 gnd.n5594 gnd.n5593 0.152939
R12962 gnd.n5595 gnd.n5594 0.152939
R12963 gnd.n5596 gnd.n5595 0.152939
R12964 gnd.n5597 gnd.n5596 0.152939
R12965 gnd.n5598 gnd.n5597 0.152939
R12966 gnd.n5599 gnd.n5598 0.152939
R12967 gnd.n5600 gnd.n5599 0.152939
R12968 gnd.n5601 gnd.n5600 0.152939
R12969 gnd.n5602 gnd.n5601 0.152939
R12970 gnd.n5602 gnd.n5365 0.152939
R12971 gnd.n5754 gnd.n5365 0.152939
R12972 gnd.n5755 gnd.n5754 0.152939
R12973 gnd.n5756 gnd.n5755 0.152939
R12974 gnd.n5757 gnd.n5756 0.152939
R12975 gnd.n5757 gnd.n5332 0.152939
R12976 gnd.n5801 gnd.n5332 0.152939
R12977 gnd.n5802 gnd.n5801 0.152939
R12978 gnd.n5803 gnd.n5802 0.152939
R12979 gnd.n5552 gnd.n5459 0.152939
R12980 gnd.n5462 gnd.n5459 0.152939
R12981 gnd.n5463 gnd.n5462 0.152939
R12982 gnd.n5464 gnd.n5463 0.152939
R12983 gnd.n5467 gnd.n5464 0.152939
R12984 gnd.n5468 gnd.n5467 0.152939
R12985 gnd.n5469 gnd.n5468 0.152939
R12986 gnd.n5470 gnd.n5469 0.152939
R12987 gnd.n5473 gnd.n5470 0.152939
R12988 gnd.n5474 gnd.n5473 0.152939
R12989 gnd.n5475 gnd.n5474 0.152939
R12990 gnd.n5476 gnd.n5475 0.152939
R12991 gnd.n5479 gnd.n5476 0.152939
R12992 gnd.n5480 gnd.n5479 0.152939
R12993 gnd.n5481 gnd.n5480 0.152939
R12994 gnd.n5482 gnd.n5481 0.152939
R12995 gnd.n5485 gnd.n5482 0.152939
R12996 gnd.n5486 gnd.n5485 0.152939
R12997 gnd.n5487 gnd.n5486 0.152939
R12998 gnd.n5488 gnd.n5487 0.152939
R12999 gnd.n5491 gnd.n5488 0.152939
R13000 gnd.n5492 gnd.n5491 0.152939
R13001 gnd.n5495 gnd.n5492 0.152939
R13002 gnd.n5496 gnd.n5495 0.152939
R13003 gnd.n5498 gnd.n5496 0.152939
R13004 gnd.n5498 gnd.n5455 0.152939
R13005 gnd.n6636 gnd.n798 0.152939
R13006 gnd.n6637 gnd.n6636 0.152939
R13007 gnd.n6638 gnd.n6637 0.152939
R13008 gnd.n6638 gnd.n792 0.152939
R13009 gnd.n6646 gnd.n792 0.152939
R13010 gnd.n6647 gnd.n6646 0.152939
R13011 gnd.n6648 gnd.n6647 0.152939
R13012 gnd.n6648 gnd.n786 0.152939
R13013 gnd.n6656 gnd.n786 0.152939
R13014 gnd.n6657 gnd.n6656 0.152939
R13015 gnd.n6658 gnd.n6657 0.152939
R13016 gnd.n6658 gnd.n780 0.152939
R13017 gnd.n6666 gnd.n780 0.152939
R13018 gnd.n6667 gnd.n6666 0.152939
R13019 gnd.n6668 gnd.n6667 0.152939
R13020 gnd.n6668 gnd.n774 0.152939
R13021 gnd.n6676 gnd.n774 0.152939
R13022 gnd.n6677 gnd.n6676 0.152939
R13023 gnd.n6678 gnd.n6677 0.152939
R13024 gnd.n6678 gnd.n768 0.152939
R13025 gnd.n6686 gnd.n768 0.152939
R13026 gnd.n6687 gnd.n6686 0.152939
R13027 gnd.n6688 gnd.n6687 0.152939
R13028 gnd.n6688 gnd.n762 0.152939
R13029 gnd.n6696 gnd.n762 0.152939
R13030 gnd.n6697 gnd.n6696 0.152939
R13031 gnd.n6698 gnd.n6697 0.152939
R13032 gnd.n6698 gnd.n756 0.152939
R13033 gnd.n6706 gnd.n756 0.152939
R13034 gnd.n6707 gnd.n6706 0.152939
R13035 gnd.n6708 gnd.n6707 0.152939
R13036 gnd.n6708 gnd.n750 0.152939
R13037 gnd.n6716 gnd.n750 0.152939
R13038 gnd.n6717 gnd.n6716 0.152939
R13039 gnd.n6718 gnd.n6717 0.152939
R13040 gnd.n6718 gnd.n744 0.152939
R13041 gnd.n6726 gnd.n744 0.152939
R13042 gnd.n6727 gnd.n6726 0.152939
R13043 gnd.n6728 gnd.n6727 0.152939
R13044 gnd.n6728 gnd.n738 0.152939
R13045 gnd.n6736 gnd.n738 0.152939
R13046 gnd.n6737 gnd.n6736 0.152939
R13047 gnd.n6738 gnd.n6737 0.152939
R13048 gnd.n6738 gnd.n732 0.152939
R13049 gnd.n6746 gnd.n732 0.152939
R13050 gnd.n6747 gnd.n6746 0.152939
R13051 gnd.n6748 gnd.n6747 0.152939
R13052 gnd.n6748 gnd.n726 0.152939
R13053 gnd.n6756 gnd.n726 0.152939
R13054 gnd.n6757 gnd.n6756 0.152939
R13055 gnd.n6758 gnd.n6757 0.152939
R13056 gnd.n6758 gnd.n720 0.152939
R13057 gnd.n6766 gnd.n720 0.152939
R13058 gnd.n6767 gnd.n6766 0.152939
R13059 gnd.n6768 gnd.n6767 0.152939
R13060 gnd.n6768 gnd.n714 0.152939
R13061 gnd.n6776 gnd.n714 0.152939
R13062 gnd.n6777 gnd.n6776 0.152939
R13063 gnd.n6778 gnd.n6777 0.152939
R13064 gnd.n6778 gnd.n708 0.152939
R13065 gnd.n6786 gnd.n708 0.152939
R13066 gnd.n6787 gnd.n6786 0.152939
R13067 gnd.n6788 gnd.n6787 0.152939
R13068 gnd.n6788 gnd.n702 0.152939
R13069 gnd.n6796 gnd.n702 0.152939
R13070 gnd.n6797 gnd.n6796 0.152939
R13071 gnd.n6798 gnd.n6797 0.152939
R13072 gnd.n6798 gnd.n696 0.152939
R13073 gnd.n6806 gnd.n696 0.152939
R13074 gnd.n6807 gnd.n6806 0.152939
R13075 gnd.n6808 gnd.n6807 0.152939
R13076 gnd.n6808 gnd.n690 0.152939
R13077 gnd.n6816 gnd.n690 0.152939
R13078 gnd.n6817 gnd.n6816 0.152939
R13079 gnd.n6818 gnd.n6817 0.152939
R13080 gnd.n6818 gnd.n684 0.152939
R13081 gnd.n6826 gnd.n684 0.152939
R13082 gnd.n6827 gnd.n6826 0.152939
R13083 gnd.n6828 gnd.n6827 0.152939
R13084 gnd.n6828 gnd.n678 0.152939
R13085 gnd.n6836 gnd.n678 0.152939
R13086 gnd.n6837 gnd.n6836 0.152939
R13087 gnd.n6838 gnd.n6837 0.152939
R13088 gnd.n6838 gnd.n672 0.152939
R13089 gnd.n6846 gnd.n672 0.152939
R13090 gnd.n6847 gnd.n6846 0.152939
R13091 gnd.n6848 gnd.n6847 0.152939
R13092 gnd.n6848 gnd.n666 0.152939
R13093 gnd.n6856 gnd.n666 0.152939
R13094 gnd.n6857 gnd.n6856 0.152939
R13095 gnd.n6858 gnd.n6857 0.152939
R13096 gnd.n6858 gnd.n660 0.152939
R13097 gnd.n6866 gnd.n660 0.152939
R13098 gnd.n6867 gnd.n6866 0.152939
R13099 gnd.n6868 gnd.n6867 0.152939
R13100 gnd.n6868 gnd.n654 0.152939
R13101 gnd.n6876 gnd.n654 0.152939
R13102 gnd.n6877 gnd.n6876 0.152939
R13103 gnd.n6878 gnd.n6877 0.152939
R13104 gnd.n6878 gnd.n648 0.152939
R13105 gnd.n6886 gnd.n648 0.152939
R13106 gnd.n6887 gnd.n6886 0.152939
R13107 gnd.n6888 gnd.n6887 0.152939
R13108 gnd.n6888 gnd.n642 0.152939
R13109 gnd.n6896 gnd.n642 0.152939
R13110 gnd.n6897 gnd.n6896 0.152939
R13111 gnd.n6898 gnd.n6897 0.152939
R13112 gnd.n6898 gnd.n636 0.152939
R13113 gnd.n6906 gnd.n636 0.152939
R13114 gnd.n6907 gnd.n6906 0.152939
R13115 gnd.n6908 gnd.n6907 0.152939
R13116 gnd.n6908 gnd.n630 0.152939
R13117 gnd.n6916 gnd.n630 0.152939
R13118 gnd.n6917 gnd.n6916 0.152939
R13119 gnd.n6918 gnd.n6917 0.152939
R13120 gnd.n6918 gnd.n624 0.152939
R13121 gnd.n6926 gnd.n624 0.152939
R13122 gnd.n6927 gnd.n6926 0.152939
R13123 gnd.n6928 gnd.n6927 0.152939
R13124 gnd.n6928 gnd.n618 0.152939
R13125 gnd.n6936 gnd.n618 0.152939
R13126 gnd.n6937 gnd.n6936 0.152939
R13127 gnd.n6938 gnd.n6937 0.152939
R13128 gnd.n6938 gnd.n612 0.152939
R13129 gnd.n6946 gnd.n612 0.152939
R13130 gnd.n6947 gnd.n6946 0.152939
R13131 gnd.n6948 gnd.n6947 0.152939
R13132 gnd.n6948 gnd.n606 0.152939
R13133 gnd.n6956 gnd.n606 0.152939
R13134 gnd.n6957 gnd.n6956 0.152939
R13135 gnd.n6958 gnd.n6957 0.152939
R13136 gnd.n6958 gnd.n600 0.152939
R13137 gnd.n6966 gnd.n600 0.152939
R13138 gnd.n6967 gnd.n6966 0.152939
R13139 gnd.n6968 gnd.n6967 0.152939
R13140 gnd.n6968 gnd.n594 0.152939
R13141 gnd.n6976 gnd.n594 0.152939
R13142 gnd.n6977 gnd.n6976 0.152939
R13143 gnd.n6978 gnd.n6977 0.152939
R13144 gnd.n6978 gnd.n588 0.152939
R13145 gnd.n6986 gnd.n588 0.152939
R13146 gnd.n6987 gnd.n6986 0.152939
R13147 gnd.n6988 gnd.n6987 0.152939
R13148 gnd.n6988 gnd.n582 0.152939
R13149 gnd.n6996 gnd.n582 0.152939
R13150 gnd.n6997 gnd.n6996 0.152939
R13151 gnd.n6998 gnd.n6997 0.152939
R13152 gnd.n6998 gnd.n576 0.152939
R13153 gnd.n7006 gnd.n576 0.152939
R13154 gnd.n7007 gnd.n7006 0.152939
R13155 gnd.n7008 gnd.n7007 0.152939
R13156 gnd.n7008 gnd.n570 0.152939
R13157 gnd.n7016 gnd.n570 0.152939
R13158 gnd.n7017 gnd.n7016 0.152939
R13159 gnd.n7018 gnd.n7017 0.152939
R13160 gnd.n7018 gnd.n564 0.152939
R13161 gnd.n7026 gnd.n564 0.152939
R13162 gnd.n7027 gnd.n7026 0.152939
R13163 gnd.n7028 gnd.n7027 0.152939
R13164 gnd.n7028 gnd.n558 0.152939
R13165 gnd.n7036 gnd.n558 0.152939
R13166 gnd.n7037 gnd.n7036 0.152939
R13167 gnd.n7038 gnd.n7037 0.152939
R13168 gnd.n7038 gnd.n552 0.152939
R13169 gnd.n7046 gnd.n552 0.152939
R13170 gnd.n7047 gnd.n7046 0.152939
R13171 gnd.n7048 gnd.n7047 0.152939
R13172 gnd.n7048 gnd.n546 0.152939
R13173 gnd.n7056 gnd.n546 0.152939
R13174 gnd.n7057 gnd.n7056 0.152939
R13175 gnd.n7058 gnd.n7057 0.152939
R13176 gnd.n7058 gnd.n540 0.152939
R13177 gnd.n7066 gnd.n540 0.152939
R13178 gnd.n7067 gnd.n7066 0.152939
R13179 gnd.n7068 gnd.n7067 0.152939
R13180 gnd.n7068 gnd.n534 0.152939
R13181 gnd.n7076 gnd.n534 0.152939
R13182 gnd.n7077 gnd.n7076 0.152939
R13183 gnd.n7078 gnd.n7077 0.152939
R13184 gnd.n7078 gnd.n528 0.152939
R13185 gnd.n7086 gnd.n528 0.152939
R13186 gnd.n7088 gnd.n7087 0.152939
R13187 gnd.n7088 gnd.n522 0.152939
R13188 gnd.n7096 gnd.n522 0.152939
R13189 gnd.n7097 gnd.n7096 0.152939
R13190 gnd.n7098 gnd.n7097 0.152939
R13191 gnd.n7098 gnd.n516 0.152939
R13192 gnd.n7106 gnd.n516 0.152939
R13193 gnd.n7107 gnd.n7106 0.152939
R13194 gnd.n7108 gnd.n7107 0.152939
R13195 gnd.n7108 gnd.n510 0.152939
R13196 gnd.n7116 gnd.n510 0.152939
R13197 gnd.n7117 gnd.n7116 0.152939
R13198 gnd.n7118 gnd.n7117 0.152939
R13199 gnd.n7118 gnd.n504 0.152939
R13200 gnd.n7126 gnd.n504 0.152939
R13201 gnd.n7127 gnd.n7126 0.152939
R13202 gnd.n7128 gnd.n7127 0.152939
R13203 gnd.n7128 gnd.n498 0.152939
R13204 gnd.n7136 gnd.n498 0.152939
R13205 gnd.n7137 gnd.n7136 0.152939
R13206 gnd.n7138 gnd.n7137 0.152939
R13207 gnd.n7138 gnd.n492 0.152939
R13208 gnd.n7146 gnd.n492 0.152939
R13209 gnd.n7147 gnd.n7146 0.152939
R13210 gnd.n7148 gnd.n7147 0.152939
R13211 gnd.n7148 gnd.n486 0.152939
R13212 gnd.n7156 gnd.n486 0.152939
R13213 gnd.n7157 gnd.n7156 0.152939
R13214 gnd.n7158 gnd.n7157 0.152939
R13215 gnd.n7158 gnd.n480 0.152939
R13216 gnd.n7166 gnd.n480 0.152939
R13217 gnd.n7167 gnd.n7166 0.152939
R13218 gnd.n7168 gnd.n7167 0.152939
R13219 gnd.n7168 gnd.n474 0.152939
R13220 gnd.n7176 gnd.n474 0.152939
R13221 gnd.n7177 gnd.n7176 0.152939
R13222 gnd.n7178 gnd.n7177 0.152939
R13223 gnd.n7178 gnd.n468 0.152939
R13224 gnd.n7186 gnd.n468 0.152939
R13225 gnd.n7187 gnd.n7186 0.152939
R13226 gnd.n7188 gnd.n7187 0.152939
R13227 gnd.n7188 gnd.n462 0.152939
R13228 gnd.n7196 gnd.n462 0.152939
R13229 gnd.n7197 gnd.n7196 0.152939
R13230 gnd.n7198 gnd.n7197 0.152939
R13231 gnd.n7198 gnd.n456 0.152939
R13232 gnd.n7206 gnd.n456 0.152939
R13233 gnd.n7207 gnd.n7206 0.152939
R13234 gnd.n7208 gnd.n7207 0.152939
R13235 gnd.n7208 gnd.n450 0.152939
R13236 gnd.n7216 gnd.n450 0.152939
R13237 gnd.n7217 gnd.n7216 0.152939
R13238 gnd.n7218 gnd.n7217 0.152939
R13239 gnd.n7218 gnd.n444 0.152939
R13240 gnd.n7226 gnd.n444 0.152939
R13241 gnd.n7227 gnd.n7226 0.152939
R13242 gnd.n7228 gnd.n7227 0.152939
R13243 gnd.n7228 gnd.n438 0.152939
R13244 gnd.n7236 gnd.n438 0.152939
R13245 gnd.n7237 gnd.n7236 0.152939
R13246 gnd.n7238 gnd.n7237 0.152939
R13247 gnd.n7238 gnd.n432 0.152939
R13248 gnd.n7246 gnd.n432 0.152939
R13249 gnd.n7247 gnd.n7246 0.152939
R13250 gnd.n7248 gnd.n7247 0.152939
R13251 gnd.n7248 gnd.n426 0.152939
R13252 gnd.n7256 gnd.n426 0.152939
R13253 gnd.n7257 gnd.n7256 0.152939
R13254 gnd.n7258 gnd.n7257 0.152939
R13255 gnd.n7258 gnd.n420 0.152939
R13256 gnd.n7266 gnd.n420 0.152939
R13257 gnd.n7267 gnd.n7266 0.152939
R13258 gnd.n7268 gnd.n7267 0.152939
R13259 gnd.n7268 gnd.n414 0.152939
R13260 gnd.n7276 gnd.n414 0.152939
R13261 gnd.n7277 gnd.n7276 0.152939
R13262 gnd.n7278 gnd.n7277 0.152939
R13263 gnd.n7278 gnd.n408 0.152939
R13264 gnd.n7286 gnd.n408 0.152939
R13265 gnd.n7287 gnd.n7286 0.152939
R13266 gnd.n7288 gnd.n7287 0.152939
R13267 gnd.n7289 gnd.n7288 0.152939
R13268 gnd.n7289 gnd.n402 0.152939
R13269 gnd.n7299 gnd.n402 0.152939
R13270 gnd.n388 gnd.n385 0.152939
R13271 gnd.n389 gnd.n388 0.152939
R13272 gnd.n390 gnd.n389 0.152939
R13273 gnd.n391 gnd.n390 0.152939
R13274 gnd.n394 gnd.n391 0.152939
R13275 gnd.n395 gnd.n394 0.152939
R13276 gnd.n396 gnd.n395 0.152939
R13277 gnd.n397 gnd.n396 0.152939
R13278 gnd.n400 gnd.n397 0.152939
R13279 gnd.n401 gnd.n400 0.152939
R13280 gnd.n7300 gnd.n401 0.152939
R13281 gnd.n118 gnd.n93 0.152939
R13282 gnd.n119 gnd.n118 0.152939
R13283 gnd.n120 gnd.n119 0.152939
R13284 gnd.n137 gnd.n120 0.152939
R13285 gnd.n138 gnd.n137 0.152939
R13286 gnd.n139 gnd.n138 0.152939
R13287 gnd.n140 gnd.n139 0.152939
R13288 gnd.n157 gnd.n140 0.152939
R13289 gnd.n158 gnd.n157 0.152939
R13290 gnd.n159 gnd.n158 0.152939
R13291 gnd.n160 gnd.n159 0.152939
R13292 gnd.n177 gnd.n160 0.152939
R13293 gnd.n178 gnd.n177 0.152939
R13294 gnd.n179 gnd.n178 0.152939
R13295 gnd.n180 gnd.n179 0.152939
R13296 gnd.n196 gnd.n180 0.152939
R13297 gnd.n197 gnd.n196 0.152939
R13298 gnd.n198 gnd.n197 0.152939
R13299 gnd.n199 gnd.n198 0.152939
R13300 gnd.n214 gnd.n199 0.152939
R13301 gnd.n7554 gnd.n214 0.152939
R13302 gnd.n7635 gnd.n80 0.152939
R13303 gnd.n7324 gnd.n80 0.152939
R13304 gnd.n7325 gnd.n7324 0.152939
R13305 gnd.n7325 gnd.n376 0.152939
R13306 gnd.n7337 gnd.n376 0.152939
R13307 gnd.n7338 gnd.n7337 0.152939
R13308 gnd.n7339 gnd.n7338 0.152939
R13309 gnd.n7339 gnd.n369 0.152939
R13310 gnd.n7351 gnd.n369 0.152939
R13311 gnd.n7352 gnd.n7351 0.152939
R13312 gnd.n7353 gnd.n7352 0.152939
R13313 gnd.n7353 gnd.n364 0.152939
R13314 gnd.n7365 gnd.n364 0.152939
R13315 gnd.n7366 gnd.n7365 0.152939
R13316 gnd.n7368 gnd.n7366 0.152939
R13317 gnd.n7368 gnd.n7367 0.152939
R13318 gnd.n7367 gnd.n358 0.152939
R13319 gnd.n7396 gnd.n358 0.152939
R13320 gnd.n7397 gnd.n7396 0.152939
R13321 gnd.n7398 gnd.n7397 0.152939
R13322 gnd.n7398 gnd.n355 0.152939
R13323 gnd.n7403 gnd.n355 0.152939
R13324 gnd.n7404 gnd.n7403 0.152939
R13325 gnd.n7405 gnd.n7404 0.152939
R13326 gnd.n7405 gnd.n352 0.152939
R13327 gnd.n7410 gnd.n352 0.152939
R13328 gnd.n7443 gnd.n318 0.152939
R13329 gnd.n320 gnd.n318 0.152939
R13330 gnd.n324 gnd.n320 0.152939
R13331 gnd.n325 gnd.n324 0.152939
R13332 gnd.n326 gnd.n325 0.152939
R13333 gnd.n327 gnd.n326 0.152939
R13334 gnd.n331 gnd.n327 0.152939
R13335 gnd.n332 gnd.n331 0.152939
R13336 gnd.n333 gnd.n332 0.152939
R13337 gnd.n334 gnd.n333 0.152939
R13338 gnd.n338 gnd.n334 0.152939
R13339 gnd.n339 gnd.n338 0.152939
R13340 gnd.n340 gnd.n339 0.152939
R13341 gnd.n341 gnd.n340 0.152939
R13342 gnd.n345 gnd.n341 0.152939
R13343 gnd.n346 gnd.n345 0.152939
R13344 gnd.n7412 gnd.n346 0.152939
R13345 gnd.n7412 gnd.n7411 0.152939
R13346 gnd.n7553 gnd.n215 0.152939
R13347 gnd.n217 gnd.n215 0.152939
R13348 gnd.n221 gnd.n217 0.152939
R13349 gnd.n222 gnd.n221 0.152939
R13350 gnd.n223 gnd.n222 0.152939
R13351 gnd.n224 gnd.n223 0.152939
R13352 gnd.n228 gnd.n224 0.152939
R13353 gnd.n229 gnd.n228 0.152939
R13354 gnd.n230 gnd.n229 0.152939
R13355 gnd.n231 gnd.n230 0.152939
R13356 gnd.n235 gnd.n231 0.152939
R13357 gnd.n236 gnd.n235 0.152939
R13358 gnd.n237 gnd.n236 0.152939
R13359 gnd.n238 gnd.n237 0.152939
R13360 gnd.n242 gnd.n238 0.152939
R13361 gnd.n243 gnd.n242 0.152939
R13362 gnd.n244 gnd.n243 0.152939
R13363 gnd.n245 gnd.n244 0.152939
R13364 gnd.n249 gnd.n245 0.152939
R13365 gnd.n250 gnd.n249 0.152939
R13366 gnd.n251 gnd.n250 0.152939
R13367 gnd.n252 gnd.n251 0.152939
R13368 gnd.n256 gnd.n252 0.152939
R13369 gnd.n257 gnd.n256 0.152939
R13370 gnd.n258 gnd.n257 0.152939
R13371 gnd.n259 gnd.n258 0.152939
R13372 gnd.n263 gnd.n259 0.152939
R13373 gnd.n264 gnd.n263 0.152939
R13374 gnd.n265 gnd.n264 0.152939
R13375 gnd.n266 gnd.n265 0.152939
R13376 gnd.n270 gnd.n266 0.152939
R13377 gnd.n271 gnd.n270 0.152939
R13378 gnd.n272 gnd.n271 0.152939
R13379 gnd.n273 gnd.n272 0.152939
R13380 gnd.n277 gnd.n273 0.152939
R13381 gnd.n278 gnd.n277 0.152939
R13382 gnd.n7484 gnd.n278 0.152939
R13383 gnd.n7484 gnd.n7483 0.152939
R13384 gnd.n7483 gnd.n7482 0.152939
R13385 gnd.n7482 gnd.n282 0.152939
R13386 gnd.n288 gnd.n282 0.152939
R13387 gnd.n289 gnd.n288 0.152939
R13388 gnd.n290 gnd.n289 0.152939
R13389 gnd.n291 gnd.n290 0.152939
R13390 gnd.n295 gnd.n291 0.152939
R13391 gnd.n296 gnd.n295 0.152939
R13392 gnd.n297 gnd.n296 0.152939
R13393 gnd.n298 gnd.n297 0.152939
R13394 gnd.n302 gnd.n298 0.152939
R13395 gnd.n303 gnd.n302 0.152939
R13396 gnd.n304 gnd.n303 0.152939
R13397 gnd.n305 gnd.n304 0.152939
R13398 gnd.n309 gnd.n305 0.152939
R13399 gnd.n310 gnd.n309 0.152939
R13400 gnd.n311 gnd.n310 0.152939
R13401 gnd.n312 gnd.n311 0.152939
R13402 gnd.n317 gnd.n312 0.152939
R13403 gnd.n7445 gnd.n317 0.152939
R13404 gnd.n4176 gnd.n4175 0.152939
R13405 gnd.n4176 gnd.n4172 0.152939
R13406 gnd.n4184 gnd.n4172 0.152939
R13407 gnd.n4185 gnd.n4184 0.152939
R13408 gnd.n4186 gnd.n4185 0.152939
R13409 gnd.n4186 gnd.n4168 0.152939
R13410 gnd.n4194 gnd.n4168 0.152939
R13411 gnd.n4195 gnd.n4194 0.152939
R13412 gnd.n4196 gnd.n4195 0.152939
R13413 gnd.n4196 gnd.n4164 0.152939
R13414 gnd.n4204 gnd.n4164 0.152939
R13415 gnd.n4205 gnd.n4204 0.152939
R13416 gnd.n4206 gnd.n4205 0.152939
R13417 gnd.n4206 gnd.n4160 0.152939
R13418 gnd.n4214 gnd.n4160 0.152939
R13419 gnd.n4215 gnd.n4214 0.152939
R13420 gnd.n4216 gnd.n4215 0.152939
R13421 gnd.n4216 gnd.n4156 0.152939
R13422 gnd.n4227 gnd.n4156 0.152939
R13423 gnd.n4228 gnd.n4227 0.152939
R13424 gnd.n4229 gnd.n4228 0.152939
R13425 gnd.n4229 gnd.n4152 0.152939
R13426 gnd.n4237 gnd.n4152 0.152939
R13427 gnd.n4238 gnd.n4237 0.152939
R13428 gnd.n4240 gnd.n4238 0.152939
R13429 gnd.n4250 gnd.n1840 0.152939
R13430 gnd.n4251 gnd.n4250 0.152939
R13431 gnd.n4252 gnd.n4251 0.152939
R13432 gnd.n4252 gnd.n1836 0.152939
R13433 gnd.n4260 gnd.n1836 0.152939
R13434 gnd.n4261 gnd.n4260 0.152939
R13435 gnd.n4262 gnd.n4261 0.152939
R13436 gnd.n4262 gnd.n1832 0.152939
R13437 gnd.n4272 gnd.n1832 0.152939
R13438 gnd.n4273 gnd.n4272 0.152939
R13439 gnd.n4274 gnd.n4273 0.152939
R13440 gnd.n4274 gnd.n1828 0.152939
R13441 gnd.n4282 gnd.n1828 0.152939
R13442 gnd.n4283 gnd.n4282 0.152939
R13443 gnd.n4284 gnd.n4283 0.152939
R13444 gnd.n4284 gnd.n1824 0.152939
R13445 gnd.n4292 gnd.n1824 0.152939
R13446 gnd.n4293 gnd.n4292 0.152939
R13447 gnd.n4294 gnd.n4293 0.152939
R13448 gnd.n4294 gnd.n1820 0.152939
R13449 gnd.n4302 gnd.n1820 0.152939
R13450 gnd.n4303 gnd.n4302 0.152939
R13451 gnd.n4304 gnd.n4303 0.152939
R13452 gnd.n4304 gnd.n1816 0.152939
R13453 gnd.n4312 gnd.n1816 0.152939
R13454 gnd.n4313 gnd.n4312 0.152939
R13455 gnd.n4315 gnd.n4313 0.152939
R13456 gnd.n4315 gnd.n4314 0.152939
R13457 gnd.n4314 gnd.n1809 0.152939
R13458 gnd.n4324 gnd.n1809 0.152939
R13459 gnd.n1607 gnd.n1606 0.152939
R13460 gnd.n1608 gnd.n1607 0.152939
R13461 gnd.n1628 gnd.n1608 0.152939
R13462 gnd.n1629 gnd.n1628 0.152939
R13463 gnd.n1630 gnd.n1629 0.152939
R13464 gnd.n1631 gnd.n1630 0.152939
R13465 gnd.n1648 gnd.n1631 0.152939
R13466 gnd.n1649 gnd.n1648 0.152939
R13467 gnd.n1650 gnd.n1649 0.152939
R13468 gnd.n1651 gnd.n1650 0.152939
R13469 gnd.n1668 gnd.n1651 0.152939
R13470 gnd.n1669 gnd.n1668 0.152939
R13471 gnd.n1670 gnd.n1669 0.152939
R13472 gnd.n1671 gnd.n1670 0.152939
R13473 gnd.n1688 gnd.n1671 0.152939
R13474 gnd.n1689 gnd.n1688 0.152939
R13475 gnd.n1690 gnd.n1689 0.152939
R13476 gnd.n1691 gnd.n1690 0.152939
R13477 gnd.n1708 gnd.n1691 0.152939
R13478 gnd.n1709 gnd.n1708 0.152939
R13479 gnd.n1709 gnd.n94 0.152939
R13480 gnd.n2946 gnd.n2945 0.152939
R13481 gnd.n2947 gnd.n2946 0.152939
R13482 gnd.n2947 gnd.n2589 0.152939
R13483 gnd.n2953 gnd.n2589 0.152939
R13484 gnd.n2954 gnd.n2953 0.152939
R13485 gnd.n2955 gnd.n2954 0.152939
R13486 gnd.n2956 gnd.n2955 0.152939
R13487 gnd.n2957 gnd.n2956 0.152939
R13488 gnd.n2960 gnd.n2957 0.152939
R13489 gnd.n2961 gnd.n2960 0.152939
R13490 gnd.n2962 gnd.n2961 0.152939
R13491 gnd.n2963 gnd.n2962 0.152939
R13492 gnd.n2965 gnd.n2963 0.152939
R13493 gnd.n2965 gnd.n2964 0.152939
R13494 gnd.n2964 gnd.n2563 0.152939
R13495 gnd.n3042 gnd.n2563 0.152939
R13496 gnd.n3043 gnd.n3042 0.152939
R13497 gnd.n3044 gnd.n3043 0.152939
R13498 gnd.n3044 gnd.n2559 0.152939
R13499 gnd.n3050 gnd.n2559 0.152939
R13500 gnd.n3051 gnd.n3050 0.152939
R13501 gnd.n3052 gnd.n3051 0.152939
R13502 gnd.n3052 gnd.n2555 0.152939
R13503 gnd.n3061 gnd.n2555 0.152939
R13504 gnd.n3062 gnd.n3061 0.152939
R13505 gnd.n3063 gnd.n3062 0.152939
R13506 gnd.n3064 gnd.n3063 0.152939
R13507 gnd.n3064 gnd.n2324 0.152939
R13508 gnd.n3157 gnd.n2324 0.152939
R13509 gnd.n3158 gnd.n3157 0.152939
R13510 gnd.n3159 gnd.n3158 0.152939
R13511 gnd.n3160 gnd.n3159 0.152939
R13512 gnd.n3160 gnd.n2299 0.152939
R13513 gnd.n3187 gnd.n2299 0.152939
R13514 gnd.n3188 gnd.n3187 0.152939
R13515 gnd.n3189 gnd.n3188 0.152939
R13516 gnd.n3190 gnd.n3189 0.152939
R13517 gnd.n3190 gnd.n2274 0.152939
R13518 gnd.n3217 gnd.n2274 0.152939
R13519 gnd.n3218 gnd.n3217 0.152939
R13520 gnd.n3219 gnd.n3218 0.152939
R13521 gnd.n3220 gnd.n3219 0.152939
R13522 gnd.n3221 gnd.n3220 0.152939
R13523 gnd.n3223 gnd.n3221 0.152939
R13524 gnd.n3224 gnd.n3223 0.152939
R13525 gnd.n3224 gnd.n2180 0.152939
R13526 gnd.n3292 gnd.n2180 0.152939
R13527 gnd.n3293 gnd.n3292 0.152939
R13528 gnd.n3294 gnd.n3293 0.152939
R13529 gnd.n3295 gnd.n3294 0.152939
R13530 gnd.n3295 gnd.n2154 0.152939
R13531 gnd.n3354 gnd.n2154 0.152939
R13532 gnd.n3355 gnd.n3354 0.152939
R13533 gnd.n3356 gnd.n3355 0.152939
R13534 gnd.n3356 gnd.n2136 0.152939
R13535 gnd.n3381 gnd.n2136 0.152939
R13536 gnd.n3382 gnd.n3381 0.152939
R13537 gnd.n3383 gnd.n3382 0.152939
R13538 gnd.n3384 gnd.n3383 0.152939
R13539 gnd.n3384 gnd.n2103 0.152939
R13540 gnd.n3432 gnd.n2103 0.152939
R13541 gnd.n3433 gnd.n3432 0.152939
R13542 gnd.n3434 gnd.n3433 0.152939
R13543 gnd.n3434 gnd.n2080 0.152939
R13544 gnd.n3472 gnd.n2080 0.152939
R13545 gnd.n3473 gnd.n3472 0.152939
R13546 gnd.n3474 gnd.n3473 0.152939
R13547 gnd.n3474 gnd.n2058 0.152939
R13548 gnd.n3528 gnd.n2058 0.152939
R13549 gnd.n3529 gnd.n3528 0.152939
R13550 gnd.n3530 gnd.n3529 0.152939
R13551 gnd.n3530 gnd.n2039 0.152939
R13552 gnd.n3553 gnd.n2039 0.152939
R13553 gnd.n3554 gnd.n3553 0.152939
R13554 gnd.n3555 gnd.n3554 0.152939
R13555 gnd.n3555 gnd.n2019 0.152939
R13556 gnd.n3613 gnd.n2019 0.152939
R13557 gnd.n3614 gnd.n3613 0.152939
R13558 gnd.n3615 gnd.n3614 0.152939
R13559 gnd.n3615 gnd.n1997 0.152939
R13560 gnd.n3642 gnd.n1997 0.152939
R13561 gnd.n3643 gnd.n3642 0.152939
R13562 gnd.n3644 gnd.n3643 0.152939
R13563 gnd.n3645 gnd.n3644 0.152939
R13564 gnd.n3645 gnd.n1969 0.152939
R13565 gnd.n3687 gnd.n1969 0.152939
R13566 gnd.n3688 gnd.n3687 0.152939
R13567 gnd.n3689 gnd.n3688 0.152939
R13568 gnd.n3690 gnd.n3689 0.152939
R13569 gnd.n3692 gnd.n3690 0.152939
R13570 gnd.n3692 gnd.n3691 0.152939
R13571 gnd.n3691 gnd.n1895 0.152939
R13572 gnd.n1896 gnd.n1895 0.152939
R13573 gnd.n1897 gnd.n1896 0.152939
R13574 gnd.n1904 gnd.n1897 0.152939
R13575 gnd.n1905 gnd.n1904 0.152939
R13576 gnd.n1906 gnd.n1905 0.152939
R13577 gnd.n1907 gnd.n1906 0.152939
R13578 gnd.n1916 gnd.n1907 0.152939
R13579 gnd.n1917 gnd.n1916 0.152939
R13580 gnd.n1918 gnd.n1917 0.152939
R13581 gnd.n1919 gnd.n1918 0.152939
R13582 gnd.n1928 gnd.n1919 0.152939
R13583 gnd.n1929 gnd.n1928 0.152939
R13584 gnd.n1930 gnd.n1929 0.152939
R13585 gnd.n1931 gnd.n1930 0.152939
R13586 gnd.n3936 gnd.n1931 0.152939
R13587 gnd.n3938 gnd.n3936 0.152939
R13588 gnd.n3938 gnd.n3937 0.152939
R13589 gnd.n3937 gnd.n1585 0.152939
R13590 gnd.n1586 gnd.n1585 0.152939
R13591 gnd.n1587 gnd.n1586 0.152939
R13592 gnd.n1593 gnd.n1587 0.152939
R13593 gnd.n1594 gnd.n1593 0.152939
R13594 gnd.n1595 gnd.n1594 0.152939
R13595 gnd.n1596 gnd.n1595 0.152939
R13596 gnd.n1776 gnd.n1596 0.152939
R13597 gnd.n1777 gnd.n1776 0.152939
R13598 gnd.n1778 gnd.n1777 0.152939
R13599 gnd.n1778 gnd.n1772 0.152939
R13600 gnd.n1784 gnd.n1772 0.152939
R13601 gnd.n1785 gnd.n1784 0.152939
R13602 gnd.n1786 gnd.n1785 0.152939
R13603 gnd.n1787 gnd.n1786 0.152939
R13604 gnd.n1788 gnd.n1787 0.152939
R13605 gnd.n1789 gnd.n1788 0.152939
R13606 gnd.n1791 gnd.n1789 0.152939
R13607 gnd.n1791 gnd.n1790 0.152939
R13608 gnd.n1790 gnd.n1751 0.152939
R13609 gnd.n4397 gnd.n1751 0.152939
R13610 gnd.n4398 gnd.n4397 0.152939
R13611 gnd.n4399 gnd.n4398 0.152939
R13612 gnd.n4399 gnd.n1747 0.152939
R13613 gnd.n4405 gnd.n1747 0.152939
R13614 gnd.n4406 gnd.n4405 0.152939
R13615 gnd.n4407 gnd.n4406 0.152939
R13616 gnd.n4408 gnd.n4407 0.152939
R13617 gnd.n2746 gnd.n2745 0.152939
R13618 gnd.n2747 gnd.n2746 0.152939
R13619 gnd.n2747 gnd.n2683 0.152939
R13620 gnd.n2753 gnd.n2683 0.152939
R13621 gnd.n2754 gnd.n2753 0.152939
R13622 gnd.n2755 gnd.n2754 0.152939
R13623 gnd.n2755 gnd.n2681 0.152939
R13624 gnd.n2761 gnd.n2681 0.152939
R13625 gnd.n2762 gnd.n2761 0.152939
R13626 gnd.n2763 gnd.n2762 0.152939
R13627 gnd.n2763 gnd.n2664 0.152939
R13628 gnd.n2775 gnd.n2664 0.152939
R13629 gnd.n2776 gnd.n2775 0.152939
R13630 gnd.n2777 gnd.n2776 0.152939
R13631 gnd.n2777 gnd.n2659 0.152939
R13632 gnd.n2828 gnd.n2659 0.152939
R13633 gnd.n2829 gnd.n2828 0.152939
R13634 gnd.n2831 gnd.n2829 0.152939
R13635 gnd.n2831 gnd.n2830 0.152939
R13636 gnd.n2830 gnd.n2655 0.152939
R13637 gnd.n2655 gnd.n2653 0.152939
R13638 gnd.n2847 gnd.n2653 0.152939
R13639 gnd.n2848 gnd.n2847 0.152939
R13640 gnd.n2849 gnd.n2848 0.152939
R13641 gnd.n2849 gnd.n2617 0.152939
R13642 gnd.n2892 gnd.n2617 0.152939
R13643 gnd.n2698 gnd.n1136 0.152939
R13644 gnd.n2706 gnd.n2698 0.152939
R13645 gnd.n2707 gnd.n2706 0.152939
R13646 gnd.n2708 gnd.n2707 0.152939
R13647 gnd.n2708 gnd.n2696 0.152939
R13648 gnd.n2716 gnd.n2696 0.152939
R13649 gnd.n2717 gnd.n2716 0.152939
R13650 gnd.n2718 gnd.n2717 0.152939
R13651 gnd.n2718 gnd.n2694 0.152939
R13652 gnd.n2726 gnd.n2694 0.152939
R13653 gnd.n2727 gnd.n2726 0.152939
R13654 gnd.n2728 gnd.n2727 0.152939
R13655 gnd.n2728 gnd.n2692 0.152939
R13656 gnd.n2736 gnd.n2692 0.152939
R13657 gnd.n2737 gnd.n2736 0.152939
R13658 gnd.n2738 gnd.n2737 0.152939
R13659 gnd.n2738 gnd.n2685 0.152939
R13660 gnd.n2742 gnd.n2685 0.152939
R13661 gnd.n1278 gnd.n1253 0.152939
R13662 gnd.n1279 gnd.n1278 0.152939
R13663 gnd.n1280 gnd.n1279 0.152939
R13664 gnd.n1298 gnd.n1280 0.152939
R13665 gnd.n1299 gnd.n1298 0.152939
R13666 gnd.n1300 gnd.n1299 0.152939
R13667 gnd.n1301 gnd.n1300 0.152939
R13668 gnd.n1317 gnd.n1301 0.152939
R13669 gnd.n1318 gnd.n1317 0.152939
R13670 gnd.n1319 gnd.n1318 0.152939
R13671 gnd.n1320 gnd.n1319 0.152939
R13672 gnd.n1338 gnd.n1320 0.152939
R13673 gnd.n1339 gnd.n1338 0.152939
R13674 gnd.n1340 gnd.n1339 0.152939
R13675 gnd.n1341 gnd.n1340 0.152939
R13676 gnd.n1358 gnd.n1341 0.152939
R13677 gnd.n1359 gnd.n1358 0.152939
R13678 gnd.n1360 gnd.n1359 0.152939
R13679 gnd.n1361 gnd.n1360 0.152939
R13680 gnd.n1378 gnd.n1361 0.152939
R13681 gnd.n4785 gnd.n1378 0.152939
R13682 gnd.n4784 gnd.n1379 0.152939
R13683 gnd.n1384 gnd.n1379 0.152939
R13684 gnd.n1385 gnd.n1384 0.152939
R13685 gnd.n1386 gnd.n1385 0.152939
R13686 gnd.n1387 gnd.n1386 0.152939
R13687 gnd.n1388 gnd.n1387 0.152939
R13688 gnd.n1392 gnd.n1388 0.152939
R13689 gnd.n1393 gnd.n1392 0.152939
R13690 gnd.n1394 gnd.n1393 0.152939
R13691 gnd.n1395 gnd.n1394 0.152939
R13692 gnd.n1399 gnd.n1395 0.152939
R13693 gnd.n1400 gnd.n1399 0.152939
R13694 gnd.n1401 gnd.n1400 0.152939
R13695 gnd.n1402 gnd.n1401 0.152939
R13696 gnd.n1406 gnd.n1402 0.152939
R13697 gnd.n1407 gnd.n1406 0.152939
R13698 gnd.n1408 gnd.n1407 0.152939
R13699 gnd.n1411 gnd.n1408 0.152939
R13700 gnd.n1415 gnd.n1411 0.152939
R13701 gnd.n1416 gnd.n1415 0.152939
R13702 gnd.n1417 gnd.n1416 0.152939
R13703 gnd.n1418 gnd.n1417 0.152939
R13704 gnd.n1422 gnd.n1418 0.152939
R13705 gnd.n1423 gnd.n1422 0.152939
R13706 gnd.n1424 gnd.n1423 0.152939
R13707 gnd.n2380 gnd.n2379 0.152939
R13708 gnd.n2389 gnd.n2380 0.152939
R13709 gnd.n2390 gnd.n2389 0.152939
R13710 gnd.n2391 gnd.n2390 0.152939
R13711 gnd.n2391 gnd.n2375 0.152939
R13712 gnd.n2399 gnd.n2375 0.152939
R13713 gnd.n2400 gnd.n2399 0.152939
R13714 gnd.n2401 gnd.n2400 0.152939
R13715 gnd.n2401 gnd.n2369 0.152939
R13716 gnd.n2409 gnd.n2369 0.152939
R13717 gnd.n2410 gnd.n2409 0.152939
R13718 gnd.n2411 gnd.n2410 0.152939
R13719 gnd.n2411 gnd.n2365 0.152939
R13720 gnd.n2419 gnd.n2365 0.152939
R13721 gnd.n2420 gnd.n2419 0.152939
R13722 gnd.n2421 gnd.n2420 0.152939
R13723 gnd.n2421 gnd.n2361 0.152939
R13724 gnd.n2429 gnd.n2361 0.152939
R13725 gnd.n2430 gnd.n2429 0.152939
R13726 gnd.n2431 gnd.n2430 0.152939
R13727 gnd.n2431 gnd.n2357 0.152939
R13728 gnd.n2439 gnd.n2357 0.152939
R13729 gnd.n2440 gnd.n2439 0.152939
R13730 gnd.n2441 gnd.n2440 0.152939
R13731 gnd.n2441 gnd.n2353 0.152939
R13732 gnd.n2449 gnd.n2353 0.152939
R13733 gnd.n2450 gnd.n2449 0.152939
R13734 gnd.n2451 gnd.n2450 0.152939
R13735 gnd.n2451 gnd.n2347 0.152939
R13736 gnd.n2458 gnd.n2347 0.152939
R13737 gnd.n1073 gnd.n1072 0.152939
R13738 gnd.n1074 gnd.n1073 0.152939
R13739 gnd.n1075 gnd.n1074 0.152939
R13740 gnd.n1076 gnd.n1075 0.152939
R13741 gnd.n1077 gnd.n1076 0.152939
R13742 gnd.n1078 gnd.n1077 0.152939
R13743 gnd.n1079 gnd.n1078 0.152939
R13744 gnd.n1080 gnd.n1079 0.152939
R13745 gnd.n1081 gnd.n1080 0.152939
R13746 gnd.n1082 gnd.n1081 0.152939
R13747 gnd.n1083 gnd.n1082 0.152939
R13748 gnd.n1084 gnd.n1083 0.152939
R13749 gnd.n1085 gnd.n1084 0.152939
R13750 gnd.n1086 gnd.n1085 0.152939
R13751 gnd.n1087 gnd.n1086 0.152939
R13752 gnd.n1088 gnd.n1087 0.152939
R13753 gnd.n1089 gnd.n1088 0.152939
R13754 gnd.n1092 gnd.n1089 0.152939
R13755 gnd.n1093 gnd.n1092 0.152939
R13756 gnd.n1094 gnd.n1093 0.152939
R13757 gnd.n1095 gnd.n1094 0.152939
R13758 gnd.n1096 gnd.n1095 0.152939
R13759 gnd.n1097 gnd.n1096 0.152939
R13760 gnd.n1098 gnd.n1097 0.152939
R13761 gnd.n1099 gnd.n1098 0.152939
R13762 gnd.n1100 gnd.n1099 0.152939
R13763 gnd.n1101 gnd.n1100 0.152939
R13764 gnd.n1102 gnd.n1101 0.152939
R13765 gnd.n1103 gnd.n1102 0.152939
R13766 gnd.n1104 gnd.n1103 0.152939
R13767 gnd.n1105 gnd.n1104 0.152939
R13768 gnd.n1106 gnd.n1105 0.152939
R13769 gnd.n1107 gnd.n1106 0.152939
R13770 gnd.n1108 gnd.n1107 0.152939
R13771 gnd.n1109 gnd.n1108 0.152939
R13772 gnd.n1110 gnd.n1109 0.152939
R13773 gnd.n1111 gnd.n1110 0.152939
R13774 gnd.n1114 gnd.n1111 0.152939
R13775 gnd.n1115 gnd.n1114 0.152939
R13776 gnd.n1116 gnd.n1115 0.152939
R13777 gnd.n1117 gnd.n1116 0.152939
R13778 gnd.n1118 gnd.n1117 0.152939
R13779 gnd.n1119 gnd.n1118 0.152939
R13780 gnd.n1120 gnd.n1119 0.152939
R13781 gnd.n1121 gnd.n1120 0.152939
R13782 gnd.n1122 gnd.n1121 0.152939
R13783 gnd.n1123 gnd.n1122 0.152939
R13784 gnd.n1124 gnd.n1123 0.152939
R13785 gnd.n1125 gnd.n1124 0.152939
R13786 gnd.n1126 gnd.n1125 0.152939
R13787 gnd.n1127 gnd.n1126 0.152939
R13788 gnd.n1128 gnd.n1127 0.152939
R13789 gnd.n1129 gnd.n1128 0.152939
R13790 gnd.n1130 gnd.n1129 0.152939
R13791 gnd.n1131 gnd.n1130 0.152939
R13792 gnd.n1132 gnd.n1131 0.152939
R13793 gnd.n4929 gnd.n1132 0.152939
R13794 gnd.n4929 gnd.n4928 0.152939
R13795 gnd.n1147 gnd.n1146 0.152939
R13796 gnd.n1148 gnd.n1147 0.152939
R13797 gnd.n1149 gnd.n1148 0.152939
R13798 gnd.n1169 gnd.n1149 0.152939
R13799 gnd.n1170 gnd.n1169 0.152939
R13800 gnd.n1171 gnd.n1170 0.152939
R13801 gnd.n1172 gnd.n1171 0.152939
R13802 gnd.n1188 gnd.n1172 0.152939
R13803 gnd.n1189 gnd.n1188 0.152939
R13804 gnd.n1190 gnd.n1189 0.152939
R13805 gnd.n1191 gnd.n1190 0.152939
R13806 gnd.n1209 gnd.n1191 0.152939
R13807 gnd.n1210 gnd.n1209 0.152939
R13808 gnd.n1211 gnd.n1210 0.152939
R13809 gnd.n1212 gnd.n1211 0.152939
R13810 gnd.n1229 gnd.n1212 0.152939
R13811 gnd.n1230 gnd.n1229 0.152939
R13812 gnd.n1231 gnd.n1230 0.152939
R13813 gnd.n1232 gnd.n1231 0.152939
R13814 gnd.n1250 gnd.n1232 0.152939
R13815 gnd.n1251 gnd.n1250 0.152939
R13816 gnd.n2789 gnd.n2783 0.152939
R13817 gnd.n2795 gnd.n2783 0.152939
R13818 gnd.n2796 gnd.n2795 0.152939
R13819 gnd.n2797 gnd.n2796 0.152939
R13820 gnd.n2798 gnd.n2797 0.152939
R13821 gnd.n2799 gnd.n2798 0.152939
R13822 gnd.n2802 gnd.n2799 0.152939
R13823 gnd.n2803 gnd.n2802 0.152939
R13824 gnd.n2804 gnd.n2803 0.152939
R13825 gnd.n2806 gnd.n2804 0.152939
R13826 gnd.n2806 gnd.n2805 0.152939
R13827 gnd.n804 gnd.n803 0.152939
R13828 gnd.n805 gnd.n804 0.152939
R13829 gnd.n810 gnd.n805 0.152939
R13830 gnd.n811 gnd.n810 0.152939
R13831 gnd.n812 gnd.n811 0.152939
R13832 gnd.n813 gnd.n812 0.152939
R13833 gnd.n818 gnd.n813 0.152939
R13834 gnd.n819 gnd.n818 0.152939
R13835 gnd.n820 gnd.n819 0.152939
R13836 gnd.n821 gnd.n820 0.152939
R13837 gnd.n826 gnd.n821 0.152939
R13838 gnd.n827 gnd.n826 0.152939
R13839 gnd.n828 gnd.n827 0.152939
R13840 gnd.n829 gnd.n828 0.152939
R13841 gnd.n834 gnd.n829 0.152939
R13842 gnd.n835 gnd.n834 0.152939
R13843 gnd.n836 gnd.n835 0.152939
R13844 gnd.n837 gnd.n836 0.152939
R13845 gnd.n842 gnd.n837 0.152939
R13846 gnd.n843 gnd.n842 0.152939
R13847 gnd.n844 gnd.n843 0.152939
R13848 gnd.n845 gnd.n844 0.152939
R13849 gnd.n850 gnd.n845 0.152939
R13850 gnd.n851 gnd.n850 0.152939
R13851 gnd.n852 gnd.n851 0.152939
R13852 gnd.n853 gnd.n852 0.152939
R13853 gnd.n858 gnd.n853 0.152939
R13854 gnd.n859 gnd.n858 0.152939
R13855 gnd.n860 gnd.n859 0.152939
R13856 gnd.n861 gnd.n860 0.152939
R13857 gnd.n866 gnd.n861 0.152939
R13858 gnd.n867 gnd.n866 0.152939
R13859 gnd.n868 gnd.n867 0.152939
R13860 gnd.n869 gnd.n868 0.152939
R13861 gnd.n874 gnd.n869 0.152939
R13862 gnd.n875 gnd.n874 0.152939
R13863 gnd.n876 gnd.n875 0.152939
R13864 gnd.n877 gnd.n876 0.152939
R13865 gnd.n882 gnd.n877 0.152939
R13866 gnd.n883 gnd.n882 0.152939
R13867 gnd.n884 gnd.n883 0.152939
R13868 gnd.n885 gnd.n884 0.152939
R13869 gnd.n890 gnd.n885 0.152939
R13870 gnd.n891 gnd.n890 0.152939
R13871 gnd.n892 gnd.n891 0.152939
R13872 gnd.n893 gnd.n892 0.152939
R13873 gnd.n898 gnd.n893 0.152939
R13874 gnd.n899 gnd.n898 0.152939
R13875 gnd.n900 gnd.n899 0.152939
R13876 gnd.n901 gnd.n900 0.152939
R13877 gnd.n906 gnd.n901 0.152939
R13878 gnd.n907 gnd.n906 0.152939
R13879 gnd.n908 gnd.n907 0.152939
R13880 gnd.n909 gnd.n908 0.152939
R13881 gnd.n914 gnd.n909 0.152939
R13882 gnd.n915 gnd.n914 0.152939
R13883 gnd.n916 gnd.n915 0.152939
R13884 gnd.n917 gnd.n916 0.152939
R13885 gnd.n922 gnd.n917 0.152939
R13886 gnd.n923 gnd.n922 0.152939
R13887 gnd.n924 gnd.n923 0.152939
R13888 gnd.n925 gnd.n924 0.152939
R13889 gnd.n930 gnd.n925 0.152939
R13890 gnd.n931 gnd.n930 0.152939
R13891 gnd.n932 gnd.n931 0.152939
R13892 gnd.n933 gnd.n932 0.152939
R13893 gnd.n938 gnd.n933 0.152939
R13894 gnd.n939 gnd.n938 0.152939
R13895 gnd.n940 gnd.n939 0.152939
R13896 gnd.n941 gnd.n940 0.152939
R13897 gnd.n946 gnd.n941 0.152939
R13898 gnd.n947 gnd.n946 0.152939
R13899 gnd.n948 gnd.n947 0.152939
R13900 gnd.n949 gnd.n948 0.152939
R13901 gnd.n954 gnd.n949 0.152939
R13902 gnd.n955 gnd.n954 0.152939
R13903 gnd.n956 gnd.n955 0.152939
R13904 gnd.n957 gnd.n956 0.152939
R13905 gnd.n962 gnd.n957 0.152939
R13906 gnd.n963 gnd.n962 0.152939
R13907 gnd.n964 gnd.n963 0.152939
R13908 gnd.n965 gnd.n964 0.152939
R13909 gnd.n2786 gnd.n965 0.152939
R13910 gnd.n2788 gnd.n2786 0.152939
R13911 gnd.n3148 gnd.n3147 0.152939
R13912 gnd.n3150 gnd.n3148 0.152939
R13913 gnd.n3150 gnd.n3149 0.152939
R13914 gnd.n3149 gnd.n2305 0.152939
R13915 gnd.n3177 gnd.n2305 0.152939
R13916 gnd.n3178 gnd.n3177 0.152939
R13917 gnd.n3180 gnd.n3178 0.152939
R13918 gnd.n3180 gnd.n3179 0.152939
R13919 gnd.n3179 gnd.n2281 0.152939
R13920 gnd.n3207 gnd.n2281 0.152939
R13921 gnd.n3208 gnd.n3207 0.152939
R13922 gnd.n3210 gnd.n3208 0.152939
R13923 gnd.n3210 gnd.n3209 0.152939
R13924 gnd.n3209 gnd.n2256 0.152939
R13925 gnd.n3247 gnd.n2256 0.152939
R13926 gnd.n3248 gnd.n3247 0.152939
R13927 gnd.n3253 gnd.n3248 0.152939
R13928 gnd.n3253 gnd.n3252 0.152939
R13929 gnd.n3252 gnd.n3251 0.152939
R13930 gnd.n3251 gnd.n2172 0.152939
R13931 gnd.n3303 gnd.n2172 0.152939
R13932 gnd.n3304 gnd.n3303 0.152939
R13933 gnd.n3325 gnd.n3304 0.152939
R13934 gnd.n3325 gnd.n3324 0.152939
R13935 gnd.n3324 gnd.n3323 0.152939
R13936 gnd.n3323 gnd.n3305 0.152939
R13937 gnd.n3319 gnd.n3305 0.152939
R13938 gnd.n3319 gnd.n3318 0.152939
R13939 gnd.n3318 gnd.n3317 0.152939
R13940 gnd.n3317 gnd.n3314 0.152939
R13941 gnd.n3314 gnd.n3313 0.152939
R13942 gnd.n3313 gnd.n2120 0.152939
R13943 gnd.n3405 gnd.n2120 0.152939
R13944 gnd.n3406 gnd.n3405 0.152939
R13945 gnd.n3407 gnd.n3406 0.152939
R13946 gnd.n3407 gnd.n2096 0.152939
R13947 gnd.n3455 gnd.n2096 0.152939
R13948 gnd.n3455 gnd.n3454 0.152939
R13949 gnd.n3454 gnd.n3453 0.152939
R13950 gnd.n3453 gnd.n2073 0.152939
R13951 gnd.n3513 gnd.n2073 0.152939
R13952 gnd.n3513 gnd.n3512 0.152939
R13953 gnd.n3512 gnd.n3511 0.152939
R13954 gnd.n3511 gnd.n2074 0.152939
R13955 gnd.n3507 gnd.n2074 0.152939
R13956 gnd.n3507 gnd.n3506 0.152939
R13957 gnd.n3506 gnd.n3505 0.152939
R13958 gnd.n3505 gnd.n3496 0.152939
R13959 gnd.n3501 gnd.n3496 0.152939
R13960 gnd.n3501 gnd.n2012 0.152939
R13961 gnd.n3623 gnd.n2012 0.152939
R13962 gnd.n3624 gnd.n3623 0.152939
R13963 gnd.n3626 gnd.n3624 0.152939
R13964 gnd.n3626 gnd.n3625 0.152939
R13965 gnd.n3625 gnd.n1983 0.152939
R13966 gnd.n3662 gnd.n1983 0.152939
R13967 gnd.n3663 gnd.n3662 0.152939
R13968 gnd.n3671 gnd.n3663 0.152939
R13969 gnd.n3671 gnd.n3670 0.152939
R13970 gnd.n3670 gnd.n3669 0.152939
R13971 gnd.n3669 gnd.n3664 0.152939
R13972 gnd.n3664 gnd.n1948 0.152939
R13973 gnd.n3719 gnd.n1948 0.152939
R13974 gnd.n3720 gnd.n3719 0.152939
R13975 gnd.n3721 gnd.n3720 0.152939
R13976 gnd.n3721 gnd.n1946 0.152939
R13977 gnd.n3727 gnd.n1946 0.152939
R13978 gnd.n3728 gnd.n3727 0.152939
R13979 gnd.n3729 gnd.n3728 0.152939
R13980 gnd.n3729 gnd.n1944 0.152939
R13981 gnd.n3735 gnd.n1944 0.152939
R13982 gnd.n3736 gnd.n3735 0.152939
R13983 gnd.n3737 gnd.n3736 0.152939
R13984 gnd.n3737 gnd.n1942 0.152939
R13985 gnd.n3743 gnd.n1942 0.152939
R13986 gnd.n3744 gnd.n3743 0.152939
R13987 gnd.n3745 gnd.n3744 0.152939
R13988 gnd.n3745 gnd.n1940 0.152939
R13989 gnd.n3751 gnd.n1940 0.152939
R13990 gnd.n3752 gnd.n3751 0.152939
R13991 gnd.n3932 gnd.n3752 0.152939
R13992 gnd.n3932 gnd.n3931 0.152939
R13993 gnd.n2895 gnd.n2894 0.152939
R13994 gnd.n2895 gnd.n2602 0.152939
R13995 gnd.n2936 gnd.n2602 0.152939
R13996 gnd.n2936 gnd.n2935 0.152939
R13997 gnd.n2935 gnd.n2934 0.152939
R13998 gnd.n2934 gnd.n2603 0.152939
R13999 gnd.n2930 gnd.n2603 0.152939
R14000 gnd.n2930 gnd.n2929 0.152939
R14001 gnd.n2929 gnd.n2928 0.152939
R14002 gnd.n2928 gnd.n2583 0.152939
R14003 gnd.n2982 gnd.n2583 0.152939
R14004 gnd.n2983 gnd.n2982 0.152939
R14005 gnd.n2984 gnd.n2983 0.152939
R14006 gnd.n2984 gnd.n2578 0.152939
R14007 gnd.n2997 gnd.n2578 0.152939
R14008 gnd.n2998 gnd.n2997 0.152939
R14009 gnd.n2999 gnd.n2998 0.152939
R14010 gnd.n2999 gnd.n2570 0.152939
R14011 gnd.n3033 gnd.n2570 0.152939
R14012 gnd.n3033 gnd.n3032 0.152939
R14013 gnd.n3032 gnd.n3031 0.152939
R14014 gnd.n3031 gnd.n2571 0.152939
R14015 gnd.n3027 gnd.n2571 0.152939
R14016 gnd.n3027 gnd.n3026 0.152939
R14017 gnd.n3026 gnd.n3025 0.152939
R14018 gnd.n3025 gnd.n2575 0.152939
R14019 gnd.n3139 gnd.n2338 0.152939
R14020 gnd.n3135 gnd.n2338 0.152939
R14021 gnd.n3135 gnd.n3134 0.152939
R14022 gnd.n3134 gnd.n3133 0.152939
R14023 gnd.n3133 gnd.n2342 0.152939
R14024 gnd.n3129 gnd.n2342 0.152939
R14025 gnd.n3141 gnd.n3140 0.152939
R14026 gnd.n3140 gnd.n2315 0.152939
R14027 gnd.n3168 gnd.n2315 0.152939
R14028 gnd.n3169 gnd.n3168 0.152939
R14029 gnd.n3171 gnd.n3169 0.152939
R14030 gnd.n3171 gnd.n3170 0.152939
R14031 gnd.n3170 gnd.n2290 0.152939
R14032 gnd.n3198 gnd.n2290 0.152939
R14033 gnd.n3199 gnd.n3198 0.152939
R14034 gnd.n3201 gnd.n3199 0.152939
R14035 gnd.n3201 gnd.n3200 0.152939
R14036 gnd.n3200 gnd.n2265 0.152939
R14037 gnd.n3238 gnd.n2265 0.152939
R14038 gnd.n3239 gnd.n3238 0.152939
R14039 gnd.n3241 gnd.n3239 0.152939
R14040 gnd.n3241 gnd.n3240 0.152939
R14041 gnd.n3240 gnd.n1498 0.152939
R14042 gnd.n4659 gnd.n1498 0.152939
R14043 gnd.n4659 gnd.n4658 0.152939
R14044 gnd.n4658 gnd.n4657 0.152939
R14045 gnd.n4657 gnd.n1499 0.152939
R14046 gnd.n4653 gnd.n1499 0.152939
R14047 gnd.n4653 gnd.n4652 0.152939
R14048 gnd.n4652 gnd.n4651 0.152939
R14049 gnd.n4651 gnd.n1504 0.152939
R14050 gnd.n4647 gnd.n1504 0.152939
R14051 gnd.n4647 gnd.n4646 0.152939
R14052 gnd.n4646 gnd.n4645 0.152939
R14053 gnd.n4645 gnd.n1509 0.152939
R14054 gnd.n4641 gnd.n1509 0.152939
R14055 gnd.n4641 gnd.n4640 0.152939
R14056 gnd.n4640 gnd.n4639 0.152939
R14057 gnd.n4639 gnd.n1514 0.152939
R14058 gnd.n4635 gnd.n1514 0.152939
R14059 gnd.n4635 gnd.n4634 0.152939
R14060 gnd.n4634 gnd.n4633 0.152939
R14061 gnd.n4633 gnd.n1519 0.152939
R14062 gnd.n4629 gnd.n1519 0.152939
R14063 gnd.n4629 gnd.n4628 0.152939
R14064 gnd.n4628 gnd.n4627 0.152939
R14065 gnd.n4627 gnd.n1524 0.152939
R14066 gnd.n4623 gnd.n1524 0.152939
R14067 gnd.n4623 gnd.n4622 0.152939
R14068 gnd.n4622 gnd.n4621 0.152939
R14069 gnd.n4621 gnd.n1529 0.152939
R14070 gnd.n4617 gnd.n1529 0.152939
R14071 gnd.n4617 gnd.n4616 0.152939
R14072 gnd.n4616 gnd.n4615 0.152939
R14073 gnd.n4615 gnd.n1534 0.152939
R14074 gnd.n4611 gnd.n1534 0.152939
R14075 gnd.n4611 gnd.n4610 0.152939
R14076 gnd.n4610 gnd.n4609 0.152939
R14077 gnd.n4609 gnd.n1539 0.152939
R14078 gnd.n4605 gnd.n1539 0.152939
R14079 gnd.n4605 gnd.n4604 0.152939
R14080 gnd.n4604 gnd.n4603 0.152939
R14081 gnd.n4603 gnd.n1544 0.152939
R14082 gnd.n4599 gnd.n1544 0.152939
R14083 gnd.n4599 gnd.n4598 0.152939
R14084 gnd.n4598 gnd.n4597 0.152939
R14085 gnd.n4597 gnd.n1549 0.152939
R14086 gnd.n4593 gnd.n1549 0.152939
R14087 gnd.n4593 gnd.n4592 0.152939
R14088 gnd.n4592 gnd.n4591 0.152939
R14089 gnd.n4591 gnd.n1554 0.152939
R14090 gnd.n4587 gnd.n1554 0.152939
R14091 gnd.n4587 gnd.n4586 0.152939
R14092 gnd.n4586 gnd.n4585 0.152939
R14093 gnd.n4585 gnd.n1559 0.152939
R14094 gnd.n4581 gnd.n1559 0.152939
R14095 gnd.n4581 gnd.n4580 0.152939
R14096 gnd.n4580 gnd.n4579 0.152939
R14097 gnd.n4579 gnd.n1564 0.152939
R14098 gnd.n4575 gnd.n1564 0.152939
R14099 gnd.n4575 gnd.n4574 0.152939
R14100 gnd.n4574 gnd.n4573 0.152939
R14101 gnd.n4573 gnd.n1569 0.152939
R14102 gnd.n4569 gnd.n1569 0.152939
R14103 gnd.n4569 gnd.n4568 0.152939
R14104 gnd.n4568 gnd.n4567 0.152939
R14105 gnd.n4567 gnd.n1574 0.152939
R14106 gnd.n1577 gnd.n1574 0.152939
R14107 gnd.n3818 gnd.n3817 0.152939
R14108 gnd.n3818 gnd.n3813 0.152939
R14109 gnd.n3826 gnd.n3813 0.152939
R14110 gnd.n3827 gnd.n3826 0.152939
R14111 gnd.n3829 gnd.n3827 0.152939
R14112 gnd.n3829 gnd.n3828 0.152939
R14113 gnd.n3758 gnd.n3753 0.152939
R14114 gnd.n3753 gnd.n1804 0.152939
R14115 gnd.n4336 gnd.n1804 0.152939
R14116 gnd.n4337 gnd.n4336 0.152939
R14117 gnd.n4338 gnd.n4337 0.152939
R14118 gnd.n4338 gnd.n1767 0.152939
R14119 gnd.n4350 gnd.n1767 0.152939
R14120 gnd.n4351 gnd.n4350 0.152939
R14121 gnd.n4352 gnd.n4351 0.152939
R14122 gnd.n4352 gnd.n1758 0.152939
R14123 gnd.n4388 gnd.n1758 0.152939
R14124 gnd.n4388 gnd.n4387 0.152939
R14125 gnd.n4387 gnd.n4386 0.152939
R14126 gnd.n4386 gnd.n1759 0.152939
R14127 gnd.n4382 gnd.n1759 0.152939
R14128 gnd.n4382 gnd.n4381 0.152939
R14129 gnd.n4381 gnd.n4380 0.152939
R14130 gnd.n4380 gnd.n1763 0.152939
R14131 gnd.n4376 gnd.n1763 0.152939
R14132 gnd.n4376 gnd.n1740 0.152939
R14133 gnd.n4448 gnd.n1740 0.152939
R14134 gnd.n4449 gnd.n4448 0.152939
R14135 gnd.n4453 gnd.n4449 0.152939
R14136 gnd.n4453 gnd.n4452 0.152939
R14137 gnd.n4452 gnd.n4451 0.152939
R14138 gnd.n4451 gnd.n79 0.152939
R14139 gnd.n3129 gnd.n3128 0.128549
R14140 gnd.n3828 gnd.n1808 0.128549
R14141 gnd.n2945 gnd.n1254 0.10111
R14142 gnd.n4408 gnd.n95 0.10111
R14143 gnd.n5887 gnd.n5279 0.0767195
R14144 gnd.n5803 gnd.n5279 0.0767195
R14145 gnd.n7626 gnd.n93 0.0767195
R14146 gnd.n7626 gnd.n94 0.0767195
R14147 gnd.n4857 gnd.n1253 0.0767195
R14148 gnd.n4857 gnd.n1251 0.0767195
R14149 gnd.n7636 gnd.n7635 0.0695946
R14150 gnd.n2893 gnd.n2892 0.0695946
R14151 gnd.n2894 gnd.n2893 0.0695946
R14152 gnd.n7636 gnd.n79 0.0695946
R14153 gnd.n3128 gnd.n2459 0.063
R14154 gnd.n4325 gnd.n1808 0.063
R14155 gnd.n385 gnd.n95 0.0523293
R14156 gnd.n2805 gnd.n1254 0.0523293
R14157 gnd.n6392 gnd.n5082 0.0477147
R14158 gnd.n4327 gnd.n4325 0.0477147
R14159 gnd.n7444 gnd.n207 0.0477147
R14160 gnd.n4927 gnd.n4926 0.0477147
R14161 gnd.n2459 gnd.n1371 0.0477147
R14162 gnd.n5553 gnd.n5449 0.0442063
R14163 gnd.n5567 gnd.n5449 0.0442063
R14164 gnd.n5568 gnd.n5567 0.0442063
R14165 gnd.n5569 gnd.n5568 0.0442063
R14166 gnd.n5569 gnd.n5437 0.0442063
R14167 gnd.n5583 gnd.n5437 0.0442063
R14168 gnd.n5584 gnd.n5583 0.0442063
R14169 gnd.n5585 gnd.n5584 0.0442063
R14170 gnd.n5585 gnd.n5424 0.0442063
R14171 gnd.n5681 gnd.n5424 0.0442063
R14172 gnd.n5684 gnd.n5683 0.0344674
R14173 gnd.n4328 gnd.n4327 0.0344674
R14174 gnd.n4328 gnd.n1618 0.0344674
R14175 gnd.n1619 gnd.n1618 0.0344674
R14176 gnd.n1620 gnd.n1619 0.0344674
R14177 gnd.n1802 gnd.n1620 0.0344674
R14178 gnd.n1802 gnd.n1638 0.0344674
R14179 gnd.n1639 gnd.n1638 0.0344674
R14180 gnd.n1640 gnd.n1639 0.0344674
R14181 gnd.n1765 gnd.n1640 0.0344674
R14182 gnd.n1765 gnd.n1659 0.0344674
R14183 gnd.n1660 gnd.n1659 0.0344674
R14184 gnd.n1661 gnd.n1660 0.0344674
R14185 gnd.n4361 gnd.n1661 0.0344674
R14186 gnd.n4361 gnd.n1678 0.0344674
R14187 gnd.n1679 gnd.n1678 0.0344674
R14188 gnd.n1680 gnd.n1679 0.0344674
R14189 gnd.n4371 gnd.n1680 0.0344674
R14190 gnd.n4371 gnd.n1699 0.0344674
R14191 gnd.n1700 gnd.n1699 0.0344674
R14192 gnd.n1701 gnd.n1700 0.0344674
R14193 gnd.n4419 gnd.n1701 0.0344674
R14194 gnd.n4419 gnd.n1716 0.0344674
R14195 gnd.n1717 gnd.n1716 0.0344674
R14196 gnd.n1718 gnd.n1717 0.0344674
R14197 gnd.n4420 gnd.n1718 0.0344674
R14198 gnd.n4421 gnd.n4420 0.0344674
R14199 gnd.n4426 gnd.n4421 0.0344674
R14200 gnd.n4428 gnd.n4426 0.0344674
R14201 gnd.n4429 gnd.n4428 0.0344674
R14202 gnd.n4429 gnd.n379 0.0344674
R14203 gnd.n379 gnd.n109 0.0344674
R14204 gnd.n110 gnd.n109 0.0344674
R14205 gnd.n111 gnd.n110 0.0344674
R14206 gnd.n373 gnd.n111 0.0344674
R14207 gnd.n373 gnd.n127 0.0344674
R14208 gnd.n128 gnd.n127 0.0344674
R14209 gnd.n129 gnd.n128 0.0344674
R14210 gnd.n367 gnd.n129 0.0344674
R14211 gnd.n367 gnd.n148 0.0344674
R14212 gnd.n149 gnd.n148 0.0344674
R14213 gnd.n150 gnd.n149 0.0344674
R14214 gnd.n361 gnd.n150 0.0344674
R14215 gnd.n361 gnd.n167 0.0344674
R14216 gnd.n168 gnd.n167 0.0344674
R14217 gnd.n169 gnd.n168 0.0344674
R14218 gnd.n7375 gnd.n169 0.0344674
R14219 gnd.n7375 gnd.n187 0.0344674
R14220 gnd.n188 gnd.n187 0.0344674
R14221 gnd.n189 gnd.n188 0.0344674
R14222 gnd.n7376 gnd.n189 0.0344674
R14223 gnd.n7376 gnd.n205 0.0344674
R14224 gnd.n206 gnd.n205 0.0344674
R14225 gnd.n207 gnd.n206 0.0344674
R14226 gnd.n4926 gnd.n1138 0.0344674
R14227 gnd.n2666 gnd.n1138 0.0344674
R14228 gnd.n2666 gnd.n1160 0.0344674
R14229 gnd.n1161 gnd.n1160 0.0344674
R14230 gnd.n1162 gnd.n1161 0.0344674
R14231 gnd.n2672 gnd.n1162 0.0344674
R14232 gnd.n2672 gnd.n1179 0.0344674
R14233 gnd.n1180 gnd.n1179 0.0344674
R14234 gnd.n1181 gnd.n1180 0.0344674
R14235 gnd.n2679 gnd.n1181 0.0344674
R14236 gnd.n2679 gnd.n1199 0.0344674
R14237 gnd.n1200 gnd.n1199 0.0344674
R14238 gnd.n1201 gnd.n1200 0.0344674
R14239 gnd.n2662 gnd.n1201 0.0344674
R14240 gnd.n2662 gnd.n1219 0.0344674
R14241 gnd.n1220 gnd.n1219 0.0344674
R14242 gnd.n1221 gnd.n1220 0.0344674
R14243 gnd.n2657 gnd.n1221 0.0344674
R14244 gnd.n2657 gnd.n1240 0.0344674
R14245 gnd.n1241 gnd.n1240 0.0344674
R14246 gnd.n1242 gnd.n1241 0.0344674
R14247 gnd.n2644 gnd.n1242 0.0344674
R14248 gnd.n2856 gnd.n2644 0.0344674
R14249 gnd.n2856 gnd.n2645 0.0344674
R14250 gnd.n2645 gnd.n2630 0.0344674
R14251 gnd.n2631 gnd.n2630 0.0344674
R14252 gnd.n2632 gnd.n2631 0.0344674
R14253 gnd.n2632 gnd.n2608 0.0344674
R14254 gnd.n2906 gnd.n2608 0.0344674
R14255 gnd.n2907 gnd.n2906 0.0344674
R14256 gnd.n2907 gnd.n1269 0.0344674
R14257 gnd.n1270 gnd.n1269 0.0344674
R14258 gnd.n1271 gnd.n1270 0.0344674
R14259 gnd.n2914 gnd.n1271 0.0344674
R14260 gnd.n2914 gnd.n1288 0.0344674
R14261 gnd.n1289 gnd.n1288 0.0344674
R14262 gnd.n1290 gnd.n1289 0.0344674
R14263 gnd.n2920 gnd.n1290 0.0344674
R14264 gnd.n2920 gnd.n1308 0.0344674
R14265 gnd.n1309 gnd.n1308 0.0344674
R14266 gnd.n1310 gnd.n1309 0.0344674
R14267 gnd.n2991 gnd.n1310 0.0344674
R14268 gnd.n2991 gnd.n1328 0.0344674
R14269 gnd.n1329 gnd.n1328 0.0344674
R14270 gnd.n1330 gnd.n1329 0.0344674
R14271 gnd.n3006 gnd.n1330 0.0344674
R14272 gnd.n3006 gnd.n1348 0.0344674
R14273 gnd.n1349 gnd.n1348 0.0344674
R14274 gnd.n1350 gnd.n1349 0.0344674
R14275 gnd.n3013 gnd.n1350 0.0344674
R14276 gnd.n3013 gnd.n1369 0.0344674
R14277 gnd.n1370 gnd.n1369 0.0344674
R14278 gnd.n1371 gnd.n1370 0.0344674
R14279 gnd.n3127 gnd.n3126 0.0344674
R14280 gnd.n3838 gnd.n3837 0.0344674
R14281 gnd.n3075 gnd.n2527 0.029712
R14282 gnd.n3768 gnd.n3759 0.029712
R14283 gnd.n5417 gnd.n5416 0.0269946
R14284 gnd.n5694 gnd.n5414 0.0269946
R14285 gnd.n5693 gnd.n5415 0.0269946
R14286 gnd.n5713 gnd.n5396 0.0269946
R14287 gnd.n5715 gnd.n5714 0.0269946
R14288 gnd.n5716 gnd.n5394 0.0269946
R14289 gnd.n5723 gnd.n5719 0.0269946
R14290 gnd.n5722 gnd.n5721 0.0269946
R14291 gnd.n5720 gnd.n5373 0.0269946
R14292 gnd.n5747 gnd.n5374 0.0269946
R14293 gnd.n5746 gnd.n5375 0.0269946
R14294 gnd.n5779 gnd.n5349 0.0269946
R14295 gnd.n5781 gnd.n5780 0.0269946
R14296 gnd.n5782 gnd.n5341 0.0269946
R14297 gnd.n5345 gnd.n5342 0.0269946
R14298 gnd.n5792 gnd.n5343 0.0269946
R14299 gnd.n5791 gnd.n5344 0.0269946
R14300 gnd.n5837 gnd.n5317 0.0269946
R14301 gnd.n5839 gnd.n5838 0.0269946
R14302 gnd.n5848 gnd.n5310 0.0269946
R14303 gnd.n5850 gnd.n5849 0.0269946
R14304 gnd.n5851 gnd.n5308 0.0269946
R14305 gnd.n5858 gnd.n5854 0.0269946
R14306 gnd.n5857 gnd.n5856 0.0269946
R14307 gnd.n5855 gnd.n5287 0.0269946
R14308 gnd.n5880 gnd.n5288 0.0269946
R14309 gnd.n5879 gnd.n5289 0.0269946
R14310 gnd.n5922 gnd.n5198 0.0269946
R14311 gnd.n5924 gnd.n5923 0.0269946
R14312 gnd.n5933 gnd.n5191 0.0269946
R14313 gnd.n5935 gnd.n5934 0.0269946
R14314 gnd.n5936 gnd.n5189 0.0269946
R14315 gnd.n5942 gnd.n5939 0.0269946
R14316 gnd.n5941 gnd.n5940 0.0269946
R14317 gnd.n5967 gnd.n5169 0.0269946
R14318 gnd.n5966 gnd.n5170 0.0269946
R14319 gnd.n5996 gnd.n5155 0.0269946
R14320 gnd.n5998 gnd.n5997 0.0269946
R14321 gnd.n6022 gnd.n5141 0.0269946
R14322 gnd.n6024 gnd.n6023 0.0269946
R14323 gnd.n6025 gnd.n974 0.0269946
R14324 gnd.n5136 gnd.n975 0.0269946
R14325 gnd.n5138 gnd.n976 0.0269946
R14326 gnd.n6033 gnd.n6032 0.0269946
R14327 gnd.n6035 gnd.n6034 0.0269946
R14328 gnd.n6036 gnd.n997 0.0269946
R14329 gnd.n6037 gnd.n998 0.0269946
R14330 gnd.n6038 gnd.n999 0.0269946
R14331 gnd.n6298 gnd.n6297 0.0269946
R14332 gnd.n6299 gnd.n1023 0.0269946
R14333 gnd.n6300 gnd.n1024 0.0269946
R14334 gnd.n6301 gnd.n1025 0.0269946
R14335 gnd.n3123 gnd.n2460 0.0225788
R14336 gnd.n3122 gnd.n2464 0.0225788
R14337 gnd.n3119 gnd.n3118 0.0225788
R14338 gnd.n3115 gnd.n2470 0.0225788
R14339 gnd.n3114 gnd.n2474 0.0225788
R14340 gnd.n3111 gnd.n3110 0.0225788
R14341 gnd.n3107 gnd.n2480 0.0225788
R14342 gnd.n3106 gnd.n2484 0.0225788
R14343 gnd.n3103 gnd.n3102 0.0225788
R14344 gnd.n3099 gnd.n2491 0.0225788
R14345 gnd.n3098 gnd.n2495 0.0225788
R14346 gnd.n3095 gnd.n3094 0.0225788
R14347 gnd.n3091 gnd.n2501 0.0225788
R14348 gnd.n3090 gnd.n2505 0.0225788
R14349 gnd.n3087 gnd.n3086 0.0225788
R14350 gnd.n3083 gnd.n2512 0.0225788
R14351 gnd.n3082 gnd.n2518 0.0225788
R14352 gnd.n2526 gnd.n2524 0.0225788
R14353 gnd.n3076 gnd.n3075 0.0225788
R14354 gnd.n3844 gnd.n3842 0.0225788
R14355 gnd.n3843 gnd.n3805 0.0225788
R14356 gnd.n3853 gnd.n3852 0.0225788
R14357 gnd.n3806 gnd.n3801 0.0225788
R14358 gnd.n3863 gnd.n3861 0.0225788
R14359 gnd.n3862 gnd.n3796 0.0225788
R14360 gnd.n3872 gnd.n3871 0.0225788
R14361 gnd.n3797 gnd.n3792 0.0225788
R14362 gnd.n3882 gnd.n3880 0.0225788
R14363 gnd.n3881 gnd.n3787 0.0225788
R14364 gnd.n3891 gnd.n3890 0.0225788
R14365 gnd.n3788 gnd.n3783 0.0225788
R14366 gnd.n3901 gnd.n3899 0.0225788
R14367 gnd.n3900 gnd.n3778 0.0225788
R14368 gnd.n3911 gnd.n3910 0.0225788
R14369 gnd.n3907 gnd.n3779 0.0225788
R14370 gnd.n3921 gnd.n3766 0.0225788
R14371 gnd.n3920 gnd.n3767 0.0225788
R14372 gnd.n3769 gnd.n3768 0.0225788
R14373 gnd.n3930 gnd.n3759 0.0218415
R14374 gnd.n2527 gnd.n2331 0.0218415
R14375 gnd.n5683 gnd.n5682 0.0202011
R14376 gnd.n5682 gnd.n5681 0.0148637
R14377 gnd.n6295 gnd.n6039 0.0144266
R14378 gnd.n6296 gnd.n6295 0.0130679
R14379 gnd.n3126 gnd.n2460 0.0123886
R14380 gnd.n3123 gnd.n3122 0.0123886
R14381 gnd.n3119 gnd.n2464 0.0123886
R14382 gnd.n3118 gnd.n2470 0.0123886
R14383 gnd.n3115 gnd.n3114 0.0123886
R14384 gnd.n3111 gnd.n2474 0.0123886
R14385 gnd.n3110 gnd.n2480 0.0123886
R14386 gnd.n3107 gnd.n3106 0.0123886
R14387 gnd.n3103 gnd.n2484 0.0123886
R14388 gnd.n3102 gnd.n2491 0.0123886
R14389 gnd.n3099 gnd.n3098 0.0123886
R14390 gnd.n3095 gnd.n2495 0.0123886
R14391 gnd.n3094 gnd.n2501 0.0123886
R14392 gnd.n3091 gnd.n3090 0.0123886
R14393 gnd.n3087 gnd.n2505 0.0123886
R14394 gnd.n3086 gnd.n2512 0.0123886
R14395 gnd.n3083 gnd.n3082 0.0123886
R14396 gnd.n2524 gnd.n2518 0.0123886
R14397 gnd.n3076 gnd.n2526 0.0123886
R14398 gnd.n3842 gnd.n3838 0.0123886
R14399 gnd.n3844 gnd.n3843 0.0123886
R14400 gnd.n3853 gnd.n3805 0.0123886
R14401 gnd.n3852 gnd.n3806 0.0123886
R14402 gnd.n3861 gnd.n3801 0.0123886
R14403 gnd.n3863 gnd.n3862 0.0123886
R14404 gnd.n3872 gnd.n3796 0.0123886
R14405 gnd.n3871 gnd.n3797 0.0123886
R14406 gnd.n3880 gnd.n3792 0.0123886
R14407 gnd.n3882 gnd.n3881 0.0123886
R14408 gnd.n3891 gnd.n3787 0.0123886
R14409 gnd.n3890 gnd.n3788 0.0123886
R14410 gnd.n3899 gnd.n3783 0.0123886
R14411 gnd.n3901 gnd.n3900 0.0123886
R14412 gnd.n3911 gnd.n3778 0.0123886
R14413 gnd.n3910 gnd.n3779 0.0123886
R14414 gnd.n3907 gnd.n3766 0.0123886
R14415 gnd.n3921 gnd.n3920 0.0123886
R14416 gnd.n3769 gnd.n3767 0.0123886
R14417 gnd.n5684 gnd.n5417 0.00797283
R14418 gnd.n5416 gnd.n5414 0.00797283
R14419 gnd.n5694 gnd.n5693 0.00797283
R14420 gnd.n5415 gnd.n5396 0.00797283
R14421 gnd.n5714 gnd.n5713 0.00797283
R14422 gnd.n5716 gnd.n5715 0.00797283
R14423 gnd.n5719 gnd.n5394 0.00797283
R14424 gnd.n5723 gnd.n5722 0.00797283
R14425 gnd.n5721 gnd.n5720 0.00797283
R14426 gnd.n5374 gnd.n5373 0.00797283
R14427 gnd.n5747 gnd.n5746 0.00797283
R14428 gnd.n5375 gnd.n5349 0.00797283
R14429 gnd.n5780 gnd.n5779 0.00797283
R14430 gnd.n5782 gnd.n5781 0.00797283
R14431 gnd.n5345 gnd.n5341 0.00797283
R14432 gnd.n5343 gnd.n5342 0.00797283
R14433 gnd.n5792 gnd.n5791 0.00797283
R14434 gnd.n5344 gnd.n5317 0.00797283
R14435 gnd.n5839 gnd.n5837 0.00797283
R14436 gnd.n5838 gnd.n5310 0.00797283
R14437 gnd.n5849 gnd.n5848 0.00797283
R14438 gnd.n5851 gnd.n5850 0.00797283
R14439 gnd.n5854 gnd.n5308 0.00797283
R14440 gnd.n5858 gnd.n5857 0.00797283
R14441 gnd.n5856 gnd.n5855 0.00797283
R14442 gnd.n5288 gnd.n5287 0.00797283
R14443 gnd.n5880 gnd.n5879 0.00797283
R14444 gnd.n5289 gnd.n5198 0.00797283
R14445 gnd.n5924 gnd.n5922 0.00797283
R14446 gnd.n5923 gnd.n5191 0.00797283
R14447 gnd.n5934 gnd.n5933 0.00797283
R14448 gnd.n5936 gnd.n5935 0.00797283
R14449 gnd.n5939 gnd.n5189 0.00797283
R14450 gnd.n5942 gnd.n5941 0.00797283
R14451 gnd.n5940 gnd.n5169 0.00797283
R14452 gnd.n5967 gnd.n5966 0.00797283
R14453 gnd.n5170 gnd.n5155 0.00797283
R14454 gnd.n5998 gnd.n5996 0.00797283
R14455 gnd.n5997 gnd.n5141 0.00797283
R14456 gnd.n6023 gnd.n6022 0.00797283
R14457 gnd.n6025 gnd.n6024 0.00797283
R14458 gnd.n5136 gnd.n974 0.00797283
R14459 gnd.n5138 gnd.n975 0.00797283
R14460 gnd.n6032 gnd.n976 0.00797283
R14461 gnd.n6034 gnd.n6033 0.00797283
R14462 gnd.n6036 gnd.n6035 0.00797283
R14463 gnd.n6037 gnd.n997 0.00797283
R14464 gnd.n6038 gnd.n998 0.00797283
R14465 gnd.n6039 gnd.n999 0.00797283
R14466 gnd.n6297 gnd.n6296 0.00797283
R14467 gnd.n6299 gnd.n6298 0.00797283
R14468 gnd.n6300 gnd.n1023 0.00797283
R14469 gnd.n6301 gnd.n1024 0.00797283
R14470 gnd.n5082 gnd.n1025 0.00797283
R14471 gnd.n3128 gnd.n3127 0.00593478
R14472 gnd.n3837 gnd.n1808 0.00593478
R14473 commonsourceibias.n35 commonsourceibias.t0 223.028
R14474 commonsourceibias.n128 commonsourceibias.t129 223.028
R14475 commonsourceibias.n307 commonsourceibias.t140 223.028
R14476 commonsourceibias.n217 commonsourceibias.t112 223.028
R14477 commonsourceibias.n454 commonsourceibias.t22 223.028
R14478 commonsourceibias.n395 commonsourceibias.t108 223.028
R14479 commonsourceibias.n679 commonsourceibias.t74 223.028
R14480 commonsourceibias.n589 commonsourceibias.t97 223.028
R14481 commonsourceibias.n99 commonsourceibias.t12 207.983
R14482 commonsourceibias.n192 commonsourceibias.t120 207.983
R14483 commonsourceibias.n371 commonsourceibias.t147 207.983
R14484 commonsourceibias.n281 commonsourceibias.t71 207.983
R14485 commonsourceibias.n520 commonsourceibias.t34 207.983
R14486 commonsourceibias.n566 commonsourceibias.t91 207.983
R14487 commonsourceibias.n745 commonsourceibias.t82 207.983
R14488 commonsourceibias.n655 commonsourceibias.t151 207.983
R14489 commonsourceibias.n97 commonsourceibias.t48 168.701
R14490 commonsourceibias.n91 commonsourceibias.t4 168.701
R14491 commonsourceibias.n17 commonsourceibias.t10 168.701
R14492 commonsourceibias.n83 commonsourceibias.t58 168.701
R14493 commonsourceibias.n77 commonsourceibias.t16 168.701
R14494 commonsourceibias.n22 commonsourceibias.t28 168.701
R14495 commonsourceibias.n69 commonsourceibias.t6 168.701
R14496 commonsourceibias.n63 commonsourceibias.t14 168.701
R14497 commonsourceibias.n25 commonsourceibias.t44 168.701
R14498 commonsourceibias.n27 commonsourceibias.t24 168.701
R14499 commonsourceibias.n29 commonsourceibias.t30 168.701
R14500 commonsourceibias.n46 commonsourceibias.t54 168.701
R14501 commonsourceibias.n40 commonsourceibias.t18 168.701
R14502 commonsourceibias.n34 commonsourceibias.t50 168.701
R14503 commonsourceibias.n190 commonsourceibias.t67 168.701
R14504 commonsourceibias.n184 commonsourceibias.t126 168.701
R14505 commonsourceibias.n5 commonsourceibias.t121 168.701
R14506 commonsourceibias.n176 commonsourceibias.t136 168.701
R14507 commonsourceibias.n170 commonsourceibias.t117 168.701
R14508 commonsourceibias.n10 commonsourceibias.t102 168.701
R14509 commonsourceibias.n162 commonsourceibias.t125 168.701
R14510 commonsourceibias.n156 commonsourceibias.t118 168.701
R14511 commonsourceibias.n118 commonsourceibias.t76 168.701
R14512 commonsourceibias.n120 commonsourceibias.t106 168.701
R14513 commonsourceibias.n122 commonsourceibias.t96 168.701
R14514 commonsourceibias.n139 commonsourceibias.t141 168.701
R14515 commonsourceibias.n133 commonsourceibias.t116 168.701
R14516 commonsourceibias.n127 commonsourceibias.t152 168.701
R14517 commonsourceibias.n306 commonsourceibias.t130 168.701
R14518 commonsourceibias.n312 commonsourceibias.t79 168.701
R14519 commonsourceibias.n318 commonsourceibias.t149 168.701
R14520 commonsourceibias.n301 commonsourceibias.t133 168.701
R14521 commonsourceibias.n299 commonsourceibias.t137 168.701
R14522 commonsourceibias.n297 commonsourceibias.t64 168.701
R14523 commonsourceibias.n335 commonsourceibias.t138 168.701
R14524 commonsourceibias.n341 commonsourceibias.t146 168.701
R14525 commonsourceibias.n294 commonsourceibias.t119 168.701
R14526 commonsourceibias.n349 commonsourceibias.t90 168.701
R14527 commonsourceibias.n355 commonsourceibias.t155 168.701
R14528 commonsourceibias.n289 commonsourceibias.t124 168.701
R14529 commonsourceibias.n363 commonsourceibias.t128 168.701
R14530 commonsourceibias.n369 commonsourceibias.t75 168.701
R14531 commonsourceibias.n279 commonsourceibias.t159 168.701
R14532 commonsourceibias.n273 commonsourceibias.t148 168.701
R14533 commonsourceibias.n199 commonsourceibias.t78 168.701
R14534 commonsourceibias.n265 commonsourceibias.t157 168.701
R14535 commonsourceibias.n259 commonsourceibias.t85 168.701
R14536 commonsourceibias.n204 commonsourceibias.t77 168.701
R14537 commonsourceibias.n251 commonsourceibias.t158 168.701
R14538 commonsourceibias.n245 commonsourceibias.t94 168.701
R14539 commonsourceibias.n207 commonsourceibias.t113 168.701
R14540 commonsourceibias.n209 commonsourceibias.t156 168.701
R14541 commonsourceibias.n211 commonsourceibias.t92 168.701
R14542 commonsourceibias.n228 commonsourceibias.t111 168.701
R14543 commonsourceibias.n222 commonsourceibias.t105 168.701
R14544 commonsourceibias.n216 commonsourceibias.t93 168.701
R14545 commonsourceibias.n453 commonsourceibias.t62 168.701
R14546 commonsourceibias.n459 commonsourceibias.t40 168.701
R14547 commonsourceibias.n465 commonsourceibias.t2 168.701
R14548 commonsourceibias.n448 commonsourceibias.t52 168.701
R14549 commonsourceibias.n446 commonsourceibias.t42 168.701
R14550 commonsourceibias.n444 commonsourceibias.t56 168.701
R14551 commonsourceibias.n482 commonsourceibias.t36 168.701
R14552 commonsourceibias.n488 commonsourceibias.t26 168.701
R14553 commonsourceibias.n490 commonsourceibias.t46 168.701
R14554 commonsourceibias.n497 commonsourceibias.t38 168.701
R14555 commonsourceibias.n503 commonsourceibias.t8 168.701
R14556 commonsourceibias.n505 commonsourceibias.t32 168.701
R14557 commonsourceibias.n512 commonsourceibias.t20 168.701
R14558 commonsourceibias.n518 commonsourceibias.t60 168.701
R14559 commonsourceibias.n564 commonsourceibias.t134 168.701
R14560 commonsourceibias.n558 commonsourceibias.t114 168.701
R14561 commonsourceibias.n551 commonsourceibias.t95 168.701
R14562 commonsourceibias.n549 commonsourceibias.t123 168.701
R14563 commonsourceibias.n543 commonsourceibias.t88 168.701
R14564 commonsourceibias.n536 commonsourceibias.t73 168.701
R14565 commonsourceibias.n534 commonsourceibias.t104 168.701
R14566 commonsourceibias.n394 commonsourceibias.t131 168.701
R14567 commonsourceibias.n400 commonsourceibias.t84 168.701
R14568 commonsourceibias.n406 commonsourceibias.t127 168.701
R14569 commonsourceibias.n389 commonsourceibias.t150 168.701
R14570 commonsourceibias.n387 commonsourceibias.t83 168.701
R14571 commonsourceibias.n385 commonsourceibias.t139 168.701
R14572 commonsourceibias.n423 commonsourceibias.t89 168.701
R14573 commonsourceibias.n678 commonsourceibias.t145 168.701
R14574 commonsourceibias.n684 commonsourceibias.t109 168.701
R14575 commonsourceibias.n690 commonsourceibias.t87 168.701
R14576 commonsourceibias.n673 commonsourceibias.t153 168.701
R14577 commonsourceibias.n671 commonsourceibias.t132 168.701
R14578 commonsourceibias.n669 commonsourceibias.t103 168.701
R14579 commonsourceibias.n707 commonsourceibias.t70 168.701
R14580 commonsourceibias.n713 commonsourceibias.t81 168.701
R14581 commonsourceibias.n715 commonsourceibias.t110 168.701
R14582 commonsourceibias.n722 commonsourceibias.t115 168.701
R14583 commonsourceibias.n728 commonsourceibias.t101 168.701
R14584 commonsourceibias.n730 commonsourceibias.t135 168.701
R14585 commonsourceibias.n737 commonsourceibias.t122 168.701
R14586 commonsourceibias.n743 commonsourceibias.t107 168.701
R14587 commonsourceibias.n588 commonsourceibias.t68 168.701
R14588 commonsourceibias.n594 commonsourceibias.t86 168.701
R14589 commonsourceibias.n600 commonsourceibias.t98 168.701
R14590 commonsourceibias.n583 commonsourceibias.t69 168.701
R14591 commonsourceibias.n581 commonsourceibias.t80 168.701
R14592 commonsourceibias.n579 commonsourceibias.t99 168.701
R14593 commonsourceibias.n617 commonsourceibias.t72 168.701
R14594 commonsourceibias.n623 commonsourceibias.t142 168.701
R14595 commonsourceibias.n625 commonsourceibias.t100 168.701
R14596 commonsourceibias.n632 commonsourceibias.t65 168.701
R14597 commonsourceibias.n638 commonsourceibias.t143 168.701
R14598 commonsourceibias.n640 commonsourceibias.t154 168.701
R14599 commonsourceibias.n647 commonsourceibias.t66 168.701
R14600 commonsourceibias.n653 commonsourceibias.t144 168.701
R14601 commonsourceibias.n36 commonsourceibias.n33 161.3
R14602 commonsourceibias.n38 commonsourceibias.n37 161.3
R14603 commonsourceibias.n39 commonsourceibias.n32 161.3
R14604 commonsourceibias.n42 commonsourceibias.n41 161.3
R14605 commonsourceibias.n43 commonsourceibias.n31 161.3
R14606 commonsourceibias.n45 commonsourceibias.n44 161.3
R14607 commonsourceibias.n47 commonsourceibias.n30 161.3
R14608 commonsourceibias.n49 commonsourceibias.n48 161.3
R14609 commonsourceibias.n51 commonsourceibias.n50 161.3
R14610 commonsourceibias.n52 commonsourceibias.n28 161.3
R14611 commonsourceibias.n54 commonsourceibias.n53 161.3
R14612 commonsourceibias.n56 commonsourceibias.n55 161.3
R14613 commonsourceibias.n57 commonsourceibias.n26 161.3
R14614 commonsourceibias.n59 commonsourceibias.n58 161.3
R14615 commonsourceibias.n61 commonsourceibias.n60 161.3
R14616 commonsourceibias.n62 commonsourceibias.n24 161.3
R14617 commonsourceibias.n65 commonsourceibias.n64 161.3
R14618 commonsourceibias.n66 commonsourceibias.n23 161.3
R14619 commonsourceibias.n68 commonsourceibias.n67 161.3
R14620 commonsourceibias.n70 commonsourceibias.n21 161.3
R14621 commonsourceibias.n72 commonsourceibias.n71 161.3
R14622 commonsourceibias.n73 commonsourceibias.n20 161.3
R14623 commonsourceibias.n75 commonsourceibias.n74 161.3
R14624 commonsourceibias.n76 commonsourceibias.n19 161.3
R14625 commonsourceibias.n79 commonsourceibias.n78 161.3
R14626 commonsourceibias.n80 commonsourceibias.n18 161.3
R14627 commonsourceibias.n82 commonsourceibias.n81 161.3
R14628 commonsourceibias.n84 commonsourceibias.n16 161.3
R14629 commonsourceibias.n86 commonsourceibias.n85 161.3
R14630 commonsourceibias.n87 commonsourceibias.n15 161.3
R14631 commonsourceibias.n89 commonsourceibias.n88 161.3
R14632 commonsourceibias.n90 commonsourceibias.n14 161.3
R14633 commonsourceibias.n93 commonsourceibias.n92 161.3
R14634 commonsourceibias.n94 commonsourceibias.n13 161.3
R14635 commonsourceibias.n96 commonsourceibias.n95 161.3
R14636 commonsourceibias.n98 commonsourceibias.n12 161.3
R14637 commonsourceibias.n129 commonsourceibias.n126 161.3
R14638 commonsourceibias.n131 commonsourceibias.n130 161.3
R14639 commonsourceibias.n132 commonsourceibias.n125 161.3
R14640 commonsourceibias.n135 commonsourceibias.n134 161.3
R14641 commonsourceibias.n136 commonsourceibias.n124 161.3
R14642 commonsourceibias.n138 commonsourceibias.n137 161.3
R14643 commonsourceibias.n140 commonsourceibias.n123 161.3
R14644 commonsourceibias.n142 commonsourceibias.n141 161.3
R14645 commonsourceibias.n144 commonsourceibias.n143 161.3
R14646 commonsourceibias.n145 commonsourceibias.n121 161.3
R14647 commonsourceibias.n147 commonsourceibias.n146 161.3
R14648 commonsourceibias.n149 commonsourceibias.n148 161.3
R14649 commonsourceibias.n150 commonsourceibias.n119 161.3
R14650 commonsourceibias.n152 commonsourceibias.n151 161.3
R14651 commonsourceibias.n154 commonsourceibias.n153 161.3
R14652 commonsourceibias.n155 commonsourceibias.n117 161.3
R14653 commonsourceibias.n158 commonsourceibias.n157 161.3
R14654 commonsourceibias.n159 commonsourceibias.n11 161.3
R14655 commonsourceibias.n161 commonsourceibias.n160 161.3
R14656 commonsourceibias.n163 commonsourceibias.n9 161.3
R14657 commonsourceibias.n165 commonsourceibias.n164 161.3
R14658 commonsourceibias.n166 commonsourceibias.n8 161.3
R14659 commonsourceibias.n168 commonsourceibias.n167 161.3
R14660 commonsourceibias.n169 commonsourceibias.n7 161.3
R14661 commonsourceibias.n172 commonsourceibias.n171 161.3
R14662 commonsourceibias.n173 commonsourceibias.n6 161.3
R14663 commonsourceibias.n175 commonsourceibias.n174 161.3
R14664 commonsourceibias.n177 commonsourceibias.n4 161.3
R14665 commonsourceibias.n179 commonsourceibias.n178 161.3
R14666 commonsourceibias.n180 commonsourceibias.n3 161.3
R14667 commonsourceibias.n182 commonsourceibias.n181 161.3
R14668 commonsourceibias.n183 commonsourceibias.n2 161.3
R14669 commonsourceibias.n186 commonsourceibias.n185 161.3
R14670 commonsourceibias.n187 commonsourceibias.n1 161.3
R14671 commonsourceibias.n189 commonsourceibias.n188 161.3
R14672 commonsourceibias.n191 commonsourceibias.n0 161.3
R14673 commonsourceibias.n370 commonsourceibias.n284 161.3
R14674 commonsourceibias.n368 commonsourceibias.n367 161.3
R14675 commonsourceibias.n366 commonsourceibias.n285 161.3
R14676 commonsourceibias.n365 commonsourceibias.n364 161.3
R14677 commonsourceibias.n362 commonsourceibias.n286 161.3
R14678 commonsourceibias.n361 commonsourceibias.n360 161.3
R14679 commonsourceibias.n359 commonsourceibias.n287 161.3
R14680 commonsourceibias.n358 commonsourceibias.n357 161.3
R14681 commonsourceibias.n356 commonsourceibias.n288 161.3
R14682 commonsourceibias.n354 commonsourceibias.n353 161.3
R14683 commonsourceibias.n352 commonsourceibias.n290 161.3
R14684 commonsourceibias.n351 commonsourceibias.n350 161.3
R14685 commonsourceibias.n348 commonsourceibias.n291 161.3
R14686 commonsourceibias.n347 commonsourceibias.n346 161.3
R14687 commonsourceibias.n345 commonsourceibias.n292 161.3
R14688 commonsourceibias.n344 commonsourceibias.n343 161.3
R14689 commonsourceibias.n342 commonsourceibias.n293 161.3
R14690 commonsourceibias.n340 commonsourceibias.n339 161.3
R14691 commonsourceibias.n338 commonsourceibias.n295 161.3
R14692 commonsourceibias.n337 commonsourceibias.n336 161.3
R14693 commonsourceibias.n334 commonsourceibias.n296 161.3
R14694 commonsourceibias.n333 commonsourceibias.n332 161.3
R14695 commonsourceibias.n331 commonsourceibias.n330 161.3
R14696 commonsourceibias.n329 commonsourceibias.n298 161.3
R14697 commonsourceibias.n328 commonsourceibias.n327 161.3
R14698 commonsourceibias.n326 commonsourceibias.n325 161.3
R14699 commonsourceibias.n324 commonsourceibias.n300 161.3
R14700 commonsourceibias.n323 commonsourceibias.n322 161.3
R14701 commonsourceibias.n321 commonsourceibias.n320 161.3
R14702 commonsourceibias.n319 commonsourceibias.n302 161.3
R14703 commonsourceibias.n317 commonsourceibias.n316 161.3
R14704 commonsourceibias.n315 commonsourceibias.n303 161.3
R14705 commonsourceibias.n314 commonsourceibias.n313 161.3
R14706 commonsourceibias.n311 commonsourceibias.n304 161.3
R14707 commonsourceibias.n310 commonsourceibias.n309 161.3
R14708 commonsourceibias.n308 commonsourceibias.n305 161.3
R14709 commonsourceibias.n218 commonsourceibias.n215 161.3
R14710 commonsourceibias.n220 commonsourceibias.n219 161.3
R14711 commonsourceibias.n221 commonsourceibias.n214 161.3
R14712 commonsourceibias.n224 commonsourceibias.n223 161.3
R14713 commonsourceibias.n225 commonsourceibias.n213 161.3
R14714 commonsourceibias.n227 commonsourceibias.n226 161.3
R14715 commonsourceibias.n229 commonsourceibias.n212 161.3
R14716 commonsourceibias.n231 commonsourceibias.n230 161.3
R14717 commonsourceibias.n233 commonsourceibias.n232 161.3
R14718 commonsourceibias.n234 commonsourceibias.n210 161.3
R14719 commonsourceibias.n236 commonsourceibias.n235 161.3
R14720 commonsourceibias.n238 commonsourceibias.n237 161.3
R14721 commonsourceibias.n239 commonsourceibias.n208 161.3
R14722 commonsourceibias.n241 commonsourceibias.n240 161.3
R14723 commonsourceibias.n243 commonsourceibias.n242 161.3
R14724 commonsourceibias.n244 commonsourceibias.n206 161.3
R14725 commonsourceibias.n247 commonsourceibias.n246 161.3
R14726 commonsourceibias.n248 commonsourceibias.n205 161.3
R14727 commonsourceibias.n250 commonsourceibias.n249 161.3
R14728 commonsourceibias.n252 commonsourceibias.n203 161.3
R14729 commonsourceibias.n254 commonsourceibias.n253 161.3
R14730 commonsourceibias.n255 commonsourceibias.n202 161.3
R14731 commonsourceibias.n257 commonsourceibias.n256 161.3
R14732 commonsourceibias.n258 commonsourceibias.n201 161.3
R14733 commonsourceibias.n261 commonsourceibias.n260 161.3
R14734 commonsourceibias.n262 commonsourceibias.n200 161.3
R14735 commonsourceibias.n264 commonsourceibias.n263 161.3
R14736 commonsourceibias.n266 commonsourceibias.n198 161.3
R14737 commonsourceibias.n268 commonsourceibias.n267 161.3
R14738 commonsourceibias.n269 commonsourceibias.n197 161.3
R14739 commonsourceibias.n271 commonsourceibias.n270 161.3
R14740 commonsourceibias.n272 commonsourceibias.n196 161.3
R14741 commonsourceibias.n275 commonsourceibias.n274 161.3
R14742 commonsourceibias.n276 commonsourceibias.n195 161.3
R14743 commonsourceibias.n278 commonsourceibias.n277 161.3
R14744 commonsourceibias.n280 commonsourceibias.n194 161.3
R14745 commonsourceibias.n519 commonsourceibias.n433 161.3
R14746 commonsourceibias.n517 commonsourceibias.n516 161.3
R14747 commonsourceibias.n515 commonsourceibias.n434 161.3
R14748 commonsourceibias.n514 commonsourceibias.n513 161.3
R14749 commonsourceibias.n511 commonsourceibias.n435 161.3
R14750 commonsourceibias.n510 commonsourceibias.n509 161.3
R14751 commonsourceibias.n508 commonsourceibias.n436 161.3
R14752 commonsourceibias.n507 commonsourceibias.n506 161.3
R14753 commonsourceibias.n504 commonsourceibias.n437 161.3
R14754 commonsourceibias.n502 commonsourceibias.n501 161.3
R14755 commonsourceibias.n500 commonsourceibias.n438 161.3
R14756 commonsourceibias.n499 commonsourceibias.n498 161.3
R14757 commonsourceibias.n496 commonsourceibias.n439 161.3
R14758 commonsourceibias.n495 commonsourceibias.n494 161.3
R14759 commonsourceibias.n493 commonsourceibias.n440 161.3
R14760 commonsourceibias.n492 commonsourceibias.n491 161.3
R14761 commonsourceibias.n489 commonsourceibias.n441 161.3
R14762 commonsourceibias.n487 commonsourceibias.n486 161.3
R14763 commonsourceibias.n485 commonsourceibias.n442 161.3
R14764 commonsourceibias.n484 commonsourceibias.n483 161.3
R14765 commonsourceibias.n481 commonsourceibias.n443 161.3
R14766 commonsourceibias.n480 commonsourceibias.n479 161.3
R14767 commonsourceibias.n478 commonsourceibias.n477 161.3
R14768 commonsourceibias.n476 commonsourceibias.n445 161.3
R14769 commonsourceibias.n475 commonsourceibias.n474 161.3
R14770 commonsourceibias.n473 commonsourceibias.n472 161.3
R14771 commonsourceibias.n471 commonsourceibias.n447 161.3
R14772 commonsourceibias.n470 commonsourceibias.n469 161.3
R14773 commonsourceibias.n468 commonsourceibias.n467 161.3
R14774 commonsourceibias.n466 commonsourceibias.n449 161.3
R14775 commonsourceibias.n464 commonsourceibias.n463 161.3
R14776 commonsourceibias.n462 commonsourceibias.n450 161.3
R14777 commonsourceibias.n461 commonsourceibias.n460 161.3
R14778 commonsourceibias.n458 commonsourceibias.n451 161.3
R14779 commonsourceibias.n457 commonsourceibias.n456 161.3
R14780 commonsourceibias.n455 commonsourceibias.n452 161.3
R14781 commonsourceibias.n425 commonsourceibias.n424 161.3
R14782 commonsourceibias.n422 commonsourceibias.n384 161.3
R14783 commonsourceibias.n421 commonsourceibias.n420 161.3
R14784 commonsourceibias.n419 commonsourceibias.n418 161.3
R14785 commonsourceibias.n417 commonsourceibias.n386 161.3
R14786 commonsourceibias.n416 commonsourceibias.n415 161.3
R14787 commonsourceibias.n414 commonsourceibias.n413 161.3
R14788 commonsourceibias.n412 commonsourceibias.n388 161.3
R14789 commonsourceibias.n411 commonsourceibias.n410 161.3
R14790 commonsourceibias.n409 commonsourceibias.n408 161.3
R14791 commonsourceibias.n407 commonsourceibias.n390 161.3
R14792 commonsourceibias.n405 commonsourceibias.n404 161.3
R14793 commonsourceibias.n403 commonsourceibias.n391 161.3
R14794 commonsourceibias.n402 commonsourceibias.n401 161.3
R14795 commonsourceibias.n399 commonsourceibias.n392 161.3
R14796 commonsourceibias.n398 commonsourceibias.n397 161.3
R14797 commonsourceibias.n396 commonsourceibias.n393 161.3
R14798 commonsourceibias.n531 commonsourceibias.n383 161.3
R14799 commonsourceibias.n565 commonsourceibias.n374 161.3
R14800 commonsourceibias.n563 commonsourceibias.n562 161.3
R14801 commonsourceibias.n561 commonsourceibias.n375 161.3
R14802 commonsourceibias.n560 commonsourceibias.n559 161.3
R14803 commonsourceibias.n557 commonsourceibias.n376 161.3
R14804 commonsourceibias.n556 commonsourceibias.n555 161.3
R14805 commonsourceibias.n554 commonsourceibias.n377 161.3
R14806 commonsourceibias.n553 commonsourceibias.n552 161.3
R14807 commonsourceibias.n550 commonsourceibias.n378 161.3
R14808 commonsourceibias.n548 commonsourceibias.n547 161.3
R14809 commonsourceibias.n546 commonsourceibias.n379 161.3
R14810 commonsourceibias.n545 commonsourceibias.n544 161.3
R14811 commonsourceibias.n542 commonsourceibias.n380 161.3
R14812 commonsourceibias.n541 commonsourceibias.n540 161.3
R14813 commonsourceibias.n539 commonsourceibias.n381 161.3
R14814 commonsourceibias.n538 commonsourceibias.n537 161.3
R14815 commonsourceibias.n535 commonsourceibias.n382 161.3
R14816 commonsourceibias.n533 commonsourceibias.n532 161.3
R14817 commonsourceibias.n744 commonsourceibias.n658 161.3
R14818 commonsourceibias.n742 commonsourceibias.n741 161.3
R14819 commonsourceibias.n740 commonsourceibias.n659 161.3
R14820 commonsourceibias.n739 commonsourceibias.n738 161.3
R14821 commonsourceibias.n736 commonsourceibias.n660 161.3
R14822 commonsourceibias.n735 commonsourceibias.n734 161.3
R14823 commonsourceibias.n733 commonsourceibias.n661 161.3
R14824 commonsourceibias.n732 commonsourceibias.n731 161.3
R14825 commonsourceibias.n729 commonsourceibias.n662 161.3
R14826 commonsourceibias.n727 commonsourceibias.n726 161.3
R14827 commonsourceibias.n725 commonsourceibias.n663 161.3
R14828 commonsourceibias.n724 commonsourceibias.n723 161.3
R14829 commonsourceibias.n721 commonsourceibias.n664 161.3
R14830 commonsourceibias.n720 commonsourceibias.n719 161.3
R14831 commonsourceibias.n718 commonsourceibias.n665 161.3
R14832 commonsourceibias.n717 commonsourceibias.n716 161.3
R14833 commonsourceibias.n714 commonsourceibias.n666 161.3
R14834 commonsourceibias.n712 commonsourceibias.n711 161.3
R14835 commonsourceibias.n710 commonsourceibias.n667 161.3
R14836 commonsourceibias.n709 commonsourceibias.n708 161.3
R14837 commonsourceibias.n706 commonsourceibias.n668 161.3
R14838 commonsourceibias.n705 commonsourceibias.n704 161.3
R14839 commonsourceibias.n703 commonsourceibias.n702 161.3
R14840 commonsourceibias.n701 commonsourceibias.n670 161.3
R14841 commonsourceibias.n700 commonsourceibias.n699 161.3
R14842 commonsourceibias.n698 commonsourceibias.n697 161.3
R14843 commonsourceibias.n696 commonsourceibias.n672 161.3
R14844 commonsourceibias.n695 commonsourceibias.n694 161.3
R14845 commonsourceibias.n693 commonsourceibias.n692 161.3
R14846 commonsourceibias.n691 commonsourceibias.n674 161.3
R14847 commonsourceibias.n689 commonsourceibias.n688 161.3
R14848 commonsourceibias.n687 commonsourceibias.n675 161.3
R14849 commonsourceibias.n686 commonsourceibias.n685 161.3
R14850 commonsourceibias.n683 commonsourceibias.n676 161.3
R14851 commonsourceibias.n682 commonsourceibias.n681 161.3
R14852 commonsourceibias.n680 commonsourceibias.n677 161.3
R14853 commonsourceibias.n654 commonsourceibias.n568 161.3
R14854 commonsourceibias.n652 commonsourceibias.n651 161.3
R14855 commonsourceibias.n650 commonsourceibias.n569 161.3
R14856 commonsourceibias.n649 commonsourceibias.n648 161.3
R14857 commonsourceibias.n646 commonsourceibias.n570 161.3
R14858 commonsourceibias.n645 commonsourceibias.n644 161.3
R14859 commonsourceibias.n643 commonsourceibias.n571 161.3
R14860 commonsourceibias.n642 commonsourceibias.n641 161.3
R14861 commonsourceibias.n639 commonsourceibias.n572 161.3
R14862 commonsourceibias.n637 commonsourceibias.n636 161.3
R14863 commonsourceibias.n635 commonsourceibias.n573 161.3
R14864 commonsourceibias.n634 commonsourceibias.n633 161.3
R14865 commonsourceibias.n631 commonsourceibias.n574 161.3
R14866 commonsourceibias.n630 commonsourceibias.n629 161.3
R14867 commonsourceibias.n628 commonsourceibias.n575 161.3
R14868 commonsourceibias.n627 commonsourceibias.n626 161.3
R14869 commonsourceibias.n624 commonsourceibias.n576 161.3
R14870 commonsourceibias.n622 commonsourceibias.n621 161.3
R14871 commonsourceibias.n620 commonsourceibias.n577 161.3
R14872 commonsourceibias.n619 commonsourceibias.n618 161.3
R14873 commonsourceibias.n616 commonsourceibias.n578 161.3
R14874 commonsourceibias.n615 commonsourceibias.n614 161.3
R14875 commonsourceibias.n613 commonsourceibias.n612 161.3
R14876 commonsourceibias.n611 commonsourceibias.n580 161.3
R14877 commonsourceibias.n610 commonsourceibias.n609 161.3
R14878 commonsourceibias.n608 commonsourceibias.n607 161.3
R14879 commonsourceibias.n606 commonsourceibias.n582 161.3
R14880 commonsourceibias.n605 commonsourceibias.n604 161.3
R14881 commonsourceibias.n603 commonsourceibias.n602 161.3
R14882 commonsourceibias.n601 commonsourceibias.n584 161.3
R14883 commonsourceibias.n599 commonsourceibias.n598 161.3
R14884 commonsourceibias.n597 commonsourceibias.n585 161.3
R14885 commonsourceibias.n596 commonsourceibias.n595 161.3
R14886 commonsourceibias.n593 commonsourceibias.n586 161.3
R14887 commonsourceibias.n592 commonsourceibias.n591 161.3
R14888 commonsourceibias.n590 commonsourceibias.n587 161.3
R14889 commonsourceibias.n111 commonsourceibias.n109 81.5057
R14890 commonsourceibias.n428 commonsourceibias.n426 81.5057
R14891 commonsourceibias.n111 commonsourceibias.n110 80.9324
R14892 commonsourceibias.n113 commonsourceibias.n112 80.9324
R14893 commonsourceibias.n115 commonsourceibias.n114 80.9324
R14894 commonsourceibias.n108 commonsourceibias.n107 80.9324
R14895 commonsourceibias.n106 commonsourceibias.n105 80.9324
R14896 commonsourceibias.n104 commonsourceibias.n103 80.9324
R14897 commonsourceibias.n102 commonsourceibias.n101 80.9324
R14898 commonsourceibias.n523 commonsourceibias.n522 80.9324
R14899 commonsourceibias.n525 commonsourceibias.n524 80.9324
R14900 commonsourceibias.n527 commonsourceibias.n526 80.9324
R14901 commonsourceibias.n529 commonsourceibias.n528 80.9324
R14902 commonsourceibias.n432 commonsourceibias.n431 80.9324
R14903 commonsourceibias.n430 commonsourceibias.n429 80.9324
R14904 commonsourceibias.n428 commonsourceibias.n427 80.9324
R14905 commonsourceibias.n100 commonsourceibias.n99 80.6037
R14906 commonsourceibias.n193 commonsourceibias.n192 80.6037
R14907 commonsourceibias.n372 commonsourceibias.n371 80.6037
R14908 commonsourceibias.n282 commonsourceibias.n281 80.6037
R14909 commonsourceibias.n521 commonsourceibias.n520 80.6037
R14910 commonsourceibias.n567 commonsourceibias.n566 80.6037
R14911 commonsourceibias.n746 commonsourceibias.n745 80.6037
R14912 commonsourceibias.n656 commonsourceibias.n655 80.6037
R14913 commonsourceibias.n85 commonsourceibias.n84 56.5617
R14914 commonsourceibias.n71 commonsourceibias.n70 56.5617
R14915 commonsourceibias.n62 commonsourceibias.n61 56.5617
R14916 commonsourceibias.n48 commonsourceibias.n47 56.5617
R14917 commonsourceibias.n178 commonsourceibias.n177 56.5617
R14918 commonsourceibias.n164 commonsourceibias.n163 56.5617
R14919 commonsourceibias.n155 commonsourceibias.n154 56.5617
R14920 commonsourceibias.n141 commonsourceibias.n140 56.5617
R14921 commonsourceibias.n320 commonsourceibias.n319 56.5617
R14922 commonsourceibias.n334 commonsourceibias.n333 56.5617
R14923 commonsourceibias.n343 commonsourceibias.n342 56.5617
R14924 commonsourceibias.n357 commonsourceibias.n356 56.5617
R14925 commonsourceibias.n267 commonsourceibias.n266 56.5617
R14926 commonsourceibias.n253 commonsourceibias.n252 56.5617
R14927 commonsourceibias.n244 commonsourceibias.n243 56.5617
R14928 commonsourceibias.n230 commonsourceibias.n229 56.5617
R14929 commonsourceibias.n467 commonsourceibias.n466 56.5617
R14930 commonsourceibias.n481 commonsourceibias.n480 56.5617
R14931 commonsourceibias.n491 commonsourceibias.n489 56.5617
R14932 commonsourceibias.n506 commonsourceibias.n504 56.5617
R14933 commonsourceibias.n552 commonsourceibias.n550 56.5617
R14934 commonsourceibias.n537 commonsourceibias.n535 56.5617
R14935 commonsourceibias.n408 commonsourceibias.n407 56.5617
R14936 commonsourceibias.n422 commonsourceibias.n421 56.5617
R14937 commonsourceibias.n692 commonsourceibias.n691 56.5617
R14938 commonsourceibias.n706 commonsourceibias.n705 56.5617
R14939 commonsourceibias.n716 commonsourceibias.n714 56.5617
R14940 commonsourceibias.n731 commonsourceibias.n729 56.5617
R14941 commonsourceibias.n602 commonsourceibias.n601 56.5617
R14942 commonsourceibias.n616 commonsourceibias.n615 56.5617
R14943 commonsourceibias.n626 commonsourceibias.n624 56.5617
R14944 commonsourceibias.n641 commonsourceibias.n639 56.5617
R14945 commonsourceibias.n76 commonsourceibias.n75 56.0773
R14946 commonsourceibias.n57 commonsourceibias.n56 56.0773
R14947 commonsourceibias.n169 commonsourceibias.n168 56.0773
R14948 commonsourceibias.n150 commonsourceibias.n149 56.0773
R14949 commonsourceibias.n329 commonsourceibias.n328 56.0773
R14950 commonsourceibias.n348 commonsourceibias.n347 56.0773
R14951 commonsourceibias.n258 commonsourceibias.n257 56.0773
R14952 commonsourceibias.n239 commonsourceibias.n238 56.0773
R14953 commonsourceibias.n476 commonsourceibias.n475 56.0773
R14954 commonsourceibias.n496 commonsourceibias.n495 56.0773
R14955 commonsourceibias.n542 commonsourceibias.n541 56.0773
R14956 commonsourceibias.n417 commonsourceibias.n416 56.0773
R14957 commonsourceibias.n701 commonsourceibias.n700 56.0773
R14958 commonsourceibias.n721 commonsourceibias.n720 56.0773
R14959 commonsourceibias.n611 commonsourceibias.n610 56.0773
R14960 commonsourceibias.n631 commonsourceibias.n630 56.0773
R14961 commonsourceibias.n99 commonsourceibias.n98 55.3321
R14962 commonsourceibias.n192 commonsourceibias.n191 55.3321
R14963 commonsourceibias.n371 commonsourceibias.n370 55.3321
R14964 commonsourceibias.n281 commonsourceibias.n280 55.3321
R14965 commonsourceibias.n520 commonsourceibias.n519 55.3321
R14966 commonsourceibias.n566 commonsourceibias.n565 55.3321
R14967 commonsourceibias.n745 commonsourceibias.n744 55.3321
R14968 commonsourceibias.n655 commonsourceibias.n654 55.3321
R14969 commonsourceibias.n90 commonsourceibias.n89 55.1086
R14970 commonsourceibias.n41 commonsourceibias.n31 55.1086
R14971 commonsourceibias.n183 commonsourceibias.n182 55.1086
R14972 commonsourceibias.n134 commonsourceibias.n124 55.1086
R14973 commonsourceibias.n313 commonsourceibias.n303 55.1086
R14974 commonsourceibias.n362 commonsourceibias.n361 55.1086
R14975 commonsourceibias.n272 commonsourceibias.n271 55.1086
R14976 commonsourceibias.n223 commonsourceibias.n213 55.1086
R14977 commonsourceibias.n460 commonsourceibias.n450 55.1086
R14978 commonsourceibias.n511 commonsourceibias.n510 55.1086
R14979 commonsourceibias.n557 commonsourceibias.n556 55.1086
R14980 commonsourceibias.n401 commonsourceibias.n391 55.1086
R14981 commonsourceibias.n685 commonsourceibias.n675 55.1086
R14982 commonsourceibias.n736 commonsourceibias.n735 55.1086
R14983 commonsourceibias.n595 commonsourceibias.n585 55.1086
R14984 commonsourceibias.n646 commonsourceibias.n645 55.1086
R14985 commonsourceibias.n35 commonsourceibias.n34 47.4592
R14986 commonsourceibias.n128 commonsourceibias.n127 47.4592
R14987 commonsourceibias.n307 commonsourceibias.n306 47.4592
R14988 commonsourceibias.n217 commonsourceibias.n216 47.4592
R14989 commonsourceibias.n454 commonsourceibias.n453 47.4592
R14990 commonsourceibias.n395 commonsourceibias.n394 47.4592
R14991 commonsourceibias.n679 commonsourceibias.n678 47.4592
R14992 commonsourceibias.n589 commonsourceibias.n588 47.4592
R14993 commonsourceibias.n308 commonsourceibias.n307 44.0436
R14994 commonsourceibias.n455 commonsourceibias.n454 44.0436
R14995 commonsourceibias.n396 commonsourceibias.n395 44.0436
R14996 commonsourceibias.n680 commonsourceibias.n679 44.0436
R14997 commonsourceibias.n590 commonsourceibias.n589 44.0436
R14998 commonsourceibias.n36 commonsourceibias.n35 44.0436
R14999 commonsourceibias.n129 commonsourceibias.n128 44.0436
R15000 commonsourceibias.n218 commonsourceibias.n217 44.0436
R15001 commonsourceibias.n92 commonsourceibias.n13 42.5146
R15002 commonsourceibias.n39 commonsourceibias.n38 42.5146
R15003 commonsourceibias.n185 commonsourceibias.n1 42.5146
R15004 commonsourceibias.n132 commonsourceibias.n131 42.5146
R15005 commonsourceibias.n311 commonsourceibias.n310 42.5146
R15006 commonsourceibias.n364 commonsourceibias.n285 42.5146
R15007 commonsourceibias.n274 commonsourceibias.n195 42.5146
R15008 commonsourceibias.n221 commonsourceibias.n220 42.5146
R15009 commonsourceibias.n458 commonsourceibias.n457 42.5146
R15010 commonsourceibias.n513 commonsourceibias.n434 42.5146
R15011 commonsourceibias.n559 commonsourceibias.n375 42.5146
R15012 commonsourceibias.n399 commonsourceibias.n398 42.5146
R15013 commonsourceibias.n683 commonsourceibias.n682 42.5146
R15014 commonsourceibias.n738 commonsourceibias.n659 42.5146
R15015 commonsourceibias.n593 commonsourceibias.n592 42.5146
R15016 commonsourceibias.n648 commonsourceibias.n569 42.5146
R15017 commonsourceibias.n78 commonsourceibias.n18 41.5458
R15018 commonsourceibias.n53 commonsourceibias.n52 41.5458
R15019 commonsourceibias.n171 commonsourceibias.n6 41.5458
R15020 commonsourceibias.n146 commonsourceibias.n145 41.5458
R15021 commonsourceibias.n325 commonsourceibias.n324 41.5458
R15022 commonsourceibias.n350 commonsourceibias.n290 41.5458
R15023 commonsourceibias.n260 commonsourceibias.n200 41.5458
R15024 commonsourceibias.n235 commonsourceibias.n234 41.5458
R15025 commonsourceibias.n472 commonsourceibias.n471 41.5458
R15026 commonsourceibias.n498 commonsourceibias.n438 41.5458
R15027 commonsourceibias.n544 commonsourceibias.n379 41.5458
R15028 commonsourceibias.n413 commonsourceibias.n412 41.5458
R15029 commonsourceibias.n697 commonsourceibias.n696 41.5458
R15030 commonsourceibias.n723 commonsourceibias.n663 41.5458
R15031 commonsourceibias.n607 commonsourceibias.n606 41.5458
R15032 commonsourceibias.n633 commonsourceibias.n573 41.5458
R15033 commonsourceibias.n68 commonsourceibias.n23 40.577
R15034 commonsourceibias.n64 commonsourceibias.n23 40.577
R15035 commonsourceibias.n161 commonsourceibias.n11 40.577
R15036 commonsourceibias.n157 commonsourceibias.n11 40.577
R15037 commonsourceibias.n336 commonsourceibias.n295 40.577
R15038 commonsourceibias.n340 commonsourceibias.n295 40.577
R15039 commonsourceibias.n250 commonsourceibias.n205 40.577
R15040 commonsourceibias.n246 commonsourceibias.n205 40.577
R15041 commonsourceibias.n483 commonsourceibias.n442 40.577
R15042 commonsourceibias.n487 commonsourceibias.n442 40.577
R15043 commonsourceibias.n533 commonsourceibias.n383 40.577
R15044 commonsourceibias.n424 commonsourceibias.n383 40.577
R15045 commonsourceibias.n708 commonsourceibias.n667 40.577
R15046 commonsourceibias.n712 commonsourceibias.n667 40.577
R15047 commonsourceibias.n618 commonsourceibias.n577 40.577
R15048 commonsourceibias.n622 commonsourceibias.n577 40.577
R15049 commonsourceibias.n82 commonsourceibias.n18 39.6083
R15050 commonsourceibias.n52 commonsourceibias.n51 39.6083
R15051 commonsourceibias.n175 commonsourceibias.n6 39.6083
R15052 commonsourceibias.n145 commonsourceibias.n144 39.6083
R15053 commonsourceibias.n324 commonsourceibias.n323 39.6083
R15054 commonsourceibias.n354 commonsourceibias.n290 39.6083
R15055 commonsourceibias.n264 commonsourceibias.n200 39.6083
R15056 commonsourceibias.n234 commonsourceibias.n233 39.6083
R15057 commonsourceibias.n471 commonsourceibias.n470 39.6083
R15058 commonsourceibias.n502 commonsourceibias.n438 39.6083
R15059 commonsourceibias.n548 commonsourceibias.n379 39.6083
R15060 commonsourceibias.n412 commonsourceibias.n411 39.6083
R15061 commonsourceibias.n696 commonsourceibias.n695 39.6083
R15062 commonsourceibias.n727 commonsourceibias.n663 39.6083
R15063 commonsourceibias.n606 commonsourceibias.n605 39.6083
R15064 commonsourceibias.n637 commonsourceibias.n573 39.6083
R15065 commonsourceibias.n96 commonsourceibias.n13 38.6395
R15066 commonsourceibias.n38 commonsourceibias.n33 38.6395
R15067 commonsourceibias.n189 commonsourceibias.n1 38.6395
R15068 commonsourceibias.n131 commonsourceibias.n126 38.6395
R15069 commonsourceibias.n310 commonsourceibias.n305 38.6395
R15070 commonsourceibias.n368 commonsourceibias.n285 38.6395
R15071 commonsourceibias.n278 commonsourceibias.n195 38.6395
R15072 commonsourceibias.n220 commonsourceibias.n215 38.6395
R15073 commonsourceibias.n457 commonsourceibias.n452 38.6395
R15074 commonsourceibias.n517 commonsourceibias.n434 38.6395
R15075 commonsourceibias.n563 commonsourceibias.n375 38.6395
R15076 commonsourceibias.n398 commonsourceibias.n393 38.6395
R15077 commonsourceibias.n682 commonsourceibias.n677 38.6395
R15078 commonsourceibias.n742 commonsourceibias.n659 38.6395
R15079 commonsourceibias.n592 commonsourceibias.n587 38.6395
R15080 commonsourceibias.n652 commonsourceibias.n569 38.6395
R15081 commonsourceibias.n89 commonsourceibias.n15 26.0455
R15082 commonsourceibias.n45 commonsourceibias.n31 26.0455
R15083 commonsourceibias.n182 commonsourceibias.n3 26.0455
R15084 commonsourceibias.n138 commonsourceibias.n124 26.0455
R15085 commonsourceibias.n317 commonsourceibias.n303 26.0455
R15086 commonsourceibias.n361 commonsourceibias.n287 26.0455
R15087 commonsourceibias.n271 commonsourceibias.n197 26.0455
R15088 commonsourceibias.n227 commonsourceibias.n213 26.0455
R15089 commonsourceibias.n464 commonsourceibias.n450 26.0455
R15090 commonsourceibias.n510 commonsourceibias.n436 26.0455
R15091 commonsourceibias.n556 commonsourceibias.n377 26.0455
R15092 commonsourceibias.n405 commonsourceibias.n391 26.0455
R15093 commonsourceibias.n689 commonsourceibias.n675 26.0455
R15094 commonsourceibias.n735 commonsourceibias.n661 26.0455
R15095 commonsourceibias.n599 commonsourceibias.n585 26.0455
R15096 commonsourceibias.n645 commonsourceibias.n571 26.0455
R15097 commonsourceibias.n75 commonsourceibias.n20 25.0767
R15098 commonsourceibias.n58 commonsourceibias.n57 25.0767
R15099 commonsourceibias.n168 commonsourceibias.n8 25.0767
R15100 commonsourceibias.n151 commonsourceibias.n150 25.0767
R15101 commonsourceibias.n330 commonsourceibias.n329 25.0767
R15102 commonsourceibias.n347 commonsourceibias.n292 25.0767
R15103 commonsourceibias.n257 commonsourceibias.n202 25.0767
R15104 commonsourceibias.n240 commonsourceibias.n239 25.0767
R15105 commonsourceibias.n477 commonsourceibias.n476 25.0767
R15106 commonsourceibias.n495 commonsourceibias.n440 25.0767
R15107 commonsourceibias.n541 commonsourceibias.n381 25.0767
R15108 commonsourceibias.n418 commonsourceibias.n417 25.0767
R15109 commonsourceibias.n702 commonsourceibias.n701 25.0767
R15110 commonsourceibias.n720 commonsourceibias.n665 25.0767
R15111 commonsourceibias.n612 commonsourceibias.n611 25.0767
R15112 commonsourceibias.n630 commonsourceibias.n575 25.0767
R15113 commonsourceibias.n71 commonsourceibias.n22 24.3464
R15114 commonsourceibias.n61 commonsourceibias.n25 24.3464
R15115 commonsourceibias.n164 commonsourceibias.n10 24.3464
R15116 commonsourceibias.n154 commonsourceibias.n118 24.3464
R15117 commonsourceibias.n333 commonsourceibias.n297 24.3464
R15118 commonsourceibias.n343 commonsourceibias.n294 24.3464
R15119 commonsourceibias.n253 commonsourceibias.n204 24.3464
R15120 commonsourceibias.n243 commonsourceibias.n207 24.3464
R15121 commonsourceibias.n480 commonsourceibias.n444 24.3464
R15122 commonsourceibias.n491 commonsourceibias.n490 24.3464
R15123 commonsourceibias.n537 commonsourceibias.n536 24.3464
R15124 commonsourceibias.n421 commonsourceibias.n385 24.3464
R15125 commonsourceibias.n705 commonsourceibias.n669 24.3464
R15126 commonsourceibias.n716 commonsourceibias.n715 24.3464
R15127 commonsourceibias.n615 commonsourceibias.n579 24.3464
R15128 commonsourceibias.n626 commonsourceibias.n625 24.3464
R15129 commonsourceibias.n85 commonsourceibias.n17 23.8546
R15130 commonsourceibias.n47 commonsourceibias.n46 23.8546
R15131 commonsourceibias.n178 commonsourceibias.n5 23.8546
R15132 commonsourceibias.n140 commonsourceibias.n139 23.8546
R15133 commonsourceibias.n319 commonsourceibias.n318 23.8546
R15134 commonsourceibias.n357 commonsourceibias.n289 23.8546
R15135 commonsourceibias.n267 commonsourceibias.n199 23.8546
R15136 commonsourceibias.n229 commonsourceibias.n228 23.8546
R15137 commonsourceibias.n466 commonsourceibias.n465 23.8546
R15138 commonsourceibias.n506 commonsourceibias.n505 23.8546
R15139 commonsourceibias.n552 commonsourceibias.n551 23.8546
R15140 commonsourceibias.n407 commonsourceibias.n406 23.8546
R15141 commonsourceibias.n691 commonsourceibias.n690 23.8546
R15142 commonsourceibias.n731 commonsourceibias.n730 23.8546
R15143 commonsourceibias.n601 commonsourceibias.n600 23.8546
R15144 commonsourceibias.n641 commonsourceibias.n640 23.8546
R15145 commonsourceibias.n98 commonsourceibias.n97 17.4607
R15146 commonsourceibias.n191 commonsourceibias.n190 17.4607
R15147 commonsourceibias.n370 commonsourceibias.n369 17.4607
R15148 commonsourceibias.n280 commonsourceibias.n279 17.4607
R15149 commonsourceibias.n519 commonsourceibias.n518 17.4607
R15150 commonsourceibias.n565 commonsourceibias.n564 17.4607
R15151 commonsourceibias.n744 commonsourceibias.n743 17.4607
R15152 commonsourceibias.n654 commonsourceibias.n653 17.4607
R15153 commonsourceibias.n84 commonsourceibias.n83 16.9689
R15154 commonsourceibias.n48 commonsourceibias.n29 16.9689
R15155 commonsourceibias.n177 commonsourceibias.n176 16.9689
R15156 commonsourceibias.n141 commonsourceibias.n122 16.9689
R15157 commonsourceibias.n320 commonsourceibias.n301 16.9689
R15158 commonsourceibias.n356 commonsourceibias.n355 16.9689
R15159 commonsourceibias.n266 commonsourceibias.n265 16.9689
R15160 commonsourceibias.n230 commonsourceibias.n211 16.9689
R15161 commonsourceibias.n467 commonsourceibias.n448 16.9689
R15162 commonsourceibias.n504 commonsourceibias.n503 16.9689
R15163 commonsourceibias.n550 commonsourceibias.n549 16.9689
R15164 commonsourceibias.n408 commonsourceibias.n389 16.9689
R15165 commonsourceibias.n692 commonsourceibias.n673 16.9689
R15166 commonsourceibias.n729 commonsourceibias.n728 16.9689
R15167 commonsourceibias.n602 commonsourceibias.n583 16.9689
R15168 commonsourceibias.n639 commonsourceibias.n638 16.9689
R15169 commonsourceibias.n70 commonsourceibias.n69 16.477
R15170 commonsourceibias.n63 commonsourceibias.n62 16.477
R15171 commonsourceibias.n163 commonsourceibias.n162 16.477
R15172 commonsourceibias.n156 commonsourceibias.n155 16.477
R15173 commonsourceibias.n335 commonsourceibias.n334 16.477
R15174 commonsourceibias.n342 commonsourceibias.n341 16.477
R15175 commonsourceibias.n252 commonsourceibias.n251 16.477
R15176 commonsourceibias.n245 commonsourceibias.n244 16.477
R15177 commonsourceibias.n482 commonsourceibias.n481 16.477
R15178 commonsourceibias.n489 commonsourceibias.n488 16.477
R15179 commonsourceibias.n535 commonsourceibias.n534 16.477
R15180 commonsourceibias.n423 commonsourceibias.n422 16.477
R15181 commonsourceibias.n707 commonsourceibias.n706 16.477
R15182 commonsourceibias.n714 commonsourceibias.n713 16.477
R15183 commonsourceibias.n617 commonsourceibias.n616 16.477
R15184 commonsourceibias.n624 commonsourceibias.n623 16.477
R15185 commonsourceibias.n77 commonsourceibias.n76 15.9852
R15186 commonsourceibias.n56 commonsourceibias.n27 15.9852
R15187 commonsourceibias.n170 commonsourceibias.n169 15.9852
R15188 commonsourceibias.n149 commonsourceibias.n120 15.9852
R15189 commonsourceibias.n328 commonsourceibias.n299 15.9852
R15190 commonsourceibias.n349 commonsourceibias.n348 15.9852
R15191 commonsourceibias.n259 commonsourceibias.n258 15.9852
R15192 commonsourceibias.n238 commonsourceibias.n209 15.9852
R15193 commonsourceibias.n475 commonsourceibias.n446 15.9852
R15194 commonsourceibias.n497 commonsourceibias.n496 15.9852
R15195 commonsourceibias.n543 commonsourceibias.n542 15.9852
R15196 commonsourceibias.n416 commonsourceibias.n387 15.9852
R15197 commonsourceibias.n700 commonsourceibias.n671 15.9852
R15198 commonsourceibias.n722 commonsourceibias.n721 15.9852
R15199 commonsourceibias.n610 commonsourceibias.n581 15.9852
R15200 commonsourceibias.n632 commonsourceibias.n631 15.9852
R15201 commonsourceibias.n91 commonsourceibias.n90 15.4934
R15202 commonsourceibias.n41 commonsourceibias.n40 15.4934
R15203 commonsourceibias.n184 commonsourceibias.n183 15.4934
R15204 commonsourceibias.n134 commonsourceibias.n133 15.4934
R15205 commonsourceibias.n313 commonsourceibias.n312 15.4934
R15206 commonsourceibias.n363 commonsourceibias.n362 15.4934
R15207 commonsourceibias.n273 commonsourceibias.n272 15.4934
R15208 commonsourceibias.n223 commonsourceibias.n222 15.4934
R15209 commonsourceibias.n460 commonsourceibias.n459 15.4934
R15210 commonsourceibias.n512 commonsourceibias.n511 15.4934
R15211 commonsourceibias.n558 commonsourceibias.n557 15.4934
R15212 commonsourceibias.n401 commonsourceibias.n400 15.4934
R15213 commonsourceibias.n685 commonsourceibias.n684 15.4934
R15214 commonsourceibias.n737 commonsourceibias.n736 15.4934
R15215 commonsourceibias.n595 commonsourceibias.n594 15.4934
R15216 commonsourceibias.n647 commonsourceibias.n646 15.4934
R15217 commonsourceibias.n102 commonsourceibias.n100 13.2663
R15218 commonsourceibias.n523 commonsourceibias.n521 13.2663
R15219 commonsourceibias.n748 commonsourceibias.n373 10.122
R15220 commonsourceibias.n159 commonsourceibias.n116 9.50363
R15221 commonsourceibias.n531 commonsourceibias.n530 9.50363
R15222 commonsourceibias.n92 commonsourceibias.n91 9.09948
R15223 commonsourceibias.n40 commonsourceibias.n39 9.09948
R15224 commonsourceibias.n185 commonsourceibias.n184 9.09948
R15225 commonsourceibias.n133 commonsourceibias.n132 9.09948
R15226 commonsourceibias.n312 commonsourceibias.n311 9.09948
R15227 commonsourceibias.n364 commonsourceibias.n363 9.09948
R15228 commonsourceibias.n274 commonsourceibias.n273 9.09948
R15229 commonsourceibias.n222 commonsourceibias.n221 9.09948
R15230 commonsourceibias.n459 commonsourceibias.n458 9.09948
R15231 commonsourceibias.n513 commonsourceibias.n512 9.09948
R15232 commonsourceibias.n559 commonsourceibias.n558 9.09948
R15233 commonsourceibias.n400 commonsourceibias.n399 9.09948
R15234 commonsourceibias.n684 commonsourceibias.n683 9.09948
R15235 commonsourceibias.n738 commonsourceibias.n737 9.09948
R15236 commonsourceibias.n594 commonsourceibias.n593 9.09948
R15237 commonsourceibias.n648 commonsourceibias.n647 9.09948
R15238 commonsourceibias.n283 commonsourceibias.n193 8.79451
R15239 commonsourceibias.n657 commonsourceibias.n567 8.79451
R15240 commonsourceibias.n78 commonsourceibias.n77 8.60764
R15241 commonsourceibias.n53 commonsourceibias.n27 8.60764
R15242 commonsourceibias.n171 commonsourceibias.n170 8.60764
R15243 commonsourceibias.n146 commonsourceibias.n120 8.60764
R15244 commonsourceibias.n325 commonsourceibias.n299 8.60764
R15245 commonsourceibias.n350 commonsourceibias.n349 8.60764
R15246 commonsourceibias.n260 commonsourceibias.n259 8.60764
R15247 commonsourceibias.n235 commonsourceibias.n209 8.60764
R15248 commonsourceibias.n472 commonsourceibias.n446 8.60764
R15249 commonsourceibias.n498 commonsourceibias.n497 8.60764
R15250 commonsourceibias.n544 commonsourceibias.n543 8.60764
R15251 commonsourceibias.n413 commonsourceibias.n387 8.60764
R15252 commonsourceibias.n697 commonsourceibias.n671 8.60764
R15253 commonsourceibias.n723 commonsourceibias.n722 8.60764
R15254 commonsourceibias.n607 commonsourceibias.n581 8.60764
R15255 commonsourceibias.n633 commonsourceibias.n632 8.60764
R15256 commonsourceibias.n748 commonsourceibias.n747 8.46921
R15257 commonsourceibias.n69 commonsourceibias.n68 8.11581
R15258 commonsourceibias.n64 commonsourceibias.n63 8.11581
R15259 commonsourceibias.n162 commonsourceibias.n161 8.11581
R15260 commonsourceibias.n157 commonsourceibias.n156 8.11581
R15261 commonsourceibias.n336 commonsourceibias.n335 8.11581
R15262 commonsourceibias.n341 commonsourceibias.n340 8.11581
R15263 commonsourceibias.n251 commonsourceibias.n250 8.11581
R15264 commonsourceibias.n246 commonsourceibias.n245 8.11581
R15265 commonsourceibias.n483 commonsourceibias.n482 8.11581
R15266 commonsourceibias.n488 commonsourceibias.n487 8.11581
R15267 commonsourceibias.n534 commonsourceibias.n533 8.11581
R15268 commonsourceibias.n424 commonsourceibias.n423 8.11581
R15269 commonsourceibias.n708 commonsourceibias.n707 8.11581
R15270 commonsourceibias.n713 commonsourceibias.n712 8.11581
R15271 commonsourceibias.n618 commonsourceibias.n617 8.11581
R15272 commonsourceibias.n623 commonsourceibias.n622 8.11581
R15273 commonsourceibias.n83 commonsourceibias.n82 7.62397
R15274 commonsourceibias.n51 commonsourceibias.n29 7.62397
R15275 commonsourceibias.n176 commonsourceibias.n175 7.62397
R15276 commonsourceibias.n144 commonsourceibias.n122 7.62397
R15277 commonsourceibias.n323 commonsourceibias.n301 7.62397
R15278 commonsourceibias.n355 commonsourceibias.n354 7.62397
R15279 commonsourceibias.n265 commonsourceibias.n264 7.62397
R15280 commonsourceibias.n233 commonsourceibias.n211 7.62397
R15281 commonsourceibias.n470 commonsourceibias.n448 7.62397
R15282 commonsourceibias.n503 commonsourceibias.n502 7.62397
R15283 commonsourceibias.n549 commonsourceibias.n548 7.62397
R15284 commonsourceibias.n411 commonsourceibias.n389 7.62397
R15285 commonsourceibias.n695 commonsourceibias.n673 7.62397
R15286 commonsourceibias.n728 commonsourceibias.n727 7.62397
R15287 commonsourceibias.n605 commonsourceibias.n583 7.62397
R15288 commonsourceibias.n638 commonsourceibias.n637 7.62397
R15289 commonsourceibias.n97 commonsourceibias.n96 7.13213
R15290 commonsourceibias.n34 commonsourceibias.n33 7.13213
R15291 commonsourceibias.n190 commonsourceibias.n189 7.13213
R15292 commonsourceibias.n127 commonsourceibias.n126 7.13213
R15293 commonsourceibias.n306 commonsourceibias.n305 7.13213
R15294 commonsourceibias.n369 commonsourceibias.n368 7.13213
R15295 commonsourceibias.n279 commonsourceibias.n278 7.13213
R15296 commonsourceibias.n216 commonsourceibias.n215 7.13213
R15297 commonsourceibias.n453 commonsourceibias.n452 7.13213
R15298 commonsourceibias.n518 commonsourceibias.n517 7.13213
R15299 commonsourceibias.n564 commonsourceibias.n563 7.13213
R15300 commonsourceibias.n394 commonsourceibias.n393 7.13213
R15301 commonsourceibias.n678 commonsourceibias.n677 7.13213
R15302 commonsourceibias.n743 commonsourceibias.n742 7.13213
R15303 commonsourceibias.n588 commonsourceibias.n587 7.13213
R15304 commonsourceibias.n653 commonsourceibias.n652 7.13213
R15305 commonsourceibias.n373 commonsourceibias.n372 5.06534
R15306 commonsourceibias.n283 commonsourceibias.n282 5.06534
R15307 commonsourceibias.n747 commonsourceibias.n746 5.06534
R15308 commonsourceibias.n657 commonsourceibias.n656 5.06534
R15309 commonsourceibias commonsourceibias.n748 4.04308
R15310 commonsourceibias.n373 commonsourceibias.n283 3.72967
R15311 commonsourceibias.n747 commonsourceibias.n657 3.72967
R15312 commonsourceibias.n109 commonsourceibias.t51 2.82907
R15313 commonsourceibias.n109 commonsourceibias.t1 2.82907
R15314 commonsourceibias.n110 commonsourceibias.t55 2.82907
R15315 commonsourceibias.n110 commonsourceibias.t19 2.82907
R15316 commonsourceibias.n112 commonsourceibias.t25 2.82907
R15317 commonsourceibias.n112 commonsourceibias.t31 2.82907
R15318 commonsourceibias.n114 commonsourceibias.t15 2.82907
R15319 commonsourceibias.n114 commonsourceibias.t45 2.82907
R15320 commonsourceibias.n107 commonsourceibias.t29 2.82907
R15321 commonsourceibias.n107 commonsourceibias.t7 2.82907
R15322 commonsourceibias.n105 commonsourceibias.t59 2.82907
R15323 commonsourceibias.n105 commonsourceibias.t17 2.82907
R15324 commonsourceibias.n103 commonsourceibias.t5 2.82907
R15325 commonsourceibias.n103 commonsourceibias.t11 2.82907
R15326 commonsourceibias.n101 commonsourceibias.t13 2.82907
R15327 commonsourceibias.n101 commonsourceibias.t49 2.82907
R15328 commonsourceibias.n522 commonsourceibias.t61 2.82907
R15329 commonsourceibias.n522 commonsourceibias.t35 2.82907
R15330 commonsourceibias.n524 commonsourceibias.t33 2.82907
R15331 commonsourceibias.n524 commonsourceibias.t21 2.82907
R15332 commonsourceibias.n526 commonsourceibias.t39 2.82907
R15333 commonsourceibias.n526 commonsourceibias.t9 2.82907
R15334 commonsourceibias.n528 commonsourceibias.t27 2.82907
R15335 commonsourceibias.n528 commonsourceibias.t47 2.82907
R15336 commonsourceibias.n431 commonsourceibias.t57 2.82907
R15337 commonsourceibias.n431 commonsourceibias.t37 2.82907
R15338 commonsourceibias.n429 commonsourceibias.t53 2.82907
R15339 commonsourceibias.n429 commonsourceibias.t43 2.82907
R15340 commonsourceibias.n427 commonsourceibias.t41 2.82907
R15341 commonsourceibias.n427 commonsourceibias.t3 2.82907
R15342 commonsourceibias.n426 commonsourceibias.t23 2.82907
R15343 commonsourceibias.n426 commonsourceibias.t63 2.82907
R15344 commonsourceibias.n17 commonsourceibias.n15 0.738255
R15345 commonsourceibias.n46 commonsourceibias.n45 0.738255
R15346 commonsourceibias.n5 commonsourceibias.n3 0.738255
R15347 commonsourceibias.n139 commonsourceibias.n138 0.738255
R15348 commonsourceibias.n318 commonsourceibias.n317 0.738255
R15349 commonsourceibias.n289 commonsourceibias.n287 0.738255
R15350 commonsourceibias.n199 commonsourceibias.n197 0.738255
R15351 commonsourceibias.n228 commonsourceibias.n227 0.738255
R15352 commonsourceibias.n465 commonsourceibias.n464 0.738255
R15353 commonsourceibias.n505 commonsourceibias.n436 0.738255
R15354 commonsourceibias.n551 commonsourceibias.n377 0.738255
R15355 commonsourceibias.n406 commonsourceibias.n405 0.738255
R15356 commonsourceibias.n690 commonsourceibias.n689 0.738255
R15357 commonsourceibias.n730 commonsourceibias.n661 0.738255
R15358 commonsourceibias.n600 commonsourceibias.n599 0.738255
R15359 commonsourceibias.n640 commonsourceibias.n571 0.738255
R15360 commonsourceibias.n104 commonsourceibias.n102 0.573776
R15361 commonsourceibias.n106 commonsourceibias.n104 0.573776
R15362 commonsourceibias.n108 commonsourceibias.n106 0.573776
R15363 commonsourceibias.n115 commonsourceibias.n113 0.573776
R15364 commonsourceibias.n113 commonsourceibias.n111 0.573776
R15365 commonsourceibias.n430 commonsourceibias.n428 0.573776
R15366 commonsourceibias.n432 commonsourceibias.n430 0.573776
R15367 commonsourceibias.n529 commonsourceibias.n527 0.573776
R15368 commonsourceibias.n527 commonsourceibias.n525 0.573776
R15369 commonsourceibias.n525 commonsourceibias.n523 0.573776
R15370 commonsourceibias.n116 commonsourceibias.n108 0.287138
R15371 commonsourceibias.n116 commonsourceibias.n115 0.287138
R15372 commonsourceibias.n530 commonsourceibias.n432 0.287138
R15373 commonsourceibias.n530 commonsourceibias.n529 0.287138
R15374 commonsourceibias.n100 commonsourceibias.n12 0.285035
R15375 commonsourceibias.n193 commonsourceibias.n0 0.285035
R15376 commonsourceibias.n372 commonsourceibias.n284 0.285035
R15377 commonsourceibias.n282 commonsourceibias.n194 0.285035
R15378 commonsourceibias.n521 commonsourceibias.n433 0.285035
R15379 commonsourceibias.n567 commonsourceibias.n374 0.285035
R15380 commonsourceibias.n746 commonsourceibias.n658 0.285035
R15381 commonsourceibias.n656 commonsourceibias.n568 0.285035
R15382 commonsourceibias.n22 commonsourceibias.n20 0.246418
R15383 commonsourceibias.n58 commonsourceibias.n25 0.246418
R15384 commonsourceibias.n10 commonsourceibias.n8 0.246418
R15385 commonsourceibias.n151 commonsourceibias.n118 0.246418
R15386 commonsourceibias.n330 commonsourceibias.n297 0.246418
R15387 commonsourceibias.n294 commonsourceibias.n292 0.246418
R15388 commonsourceibias.n204 commonsourceibias.n202 0.246418
R15389 commonsourceibias.n240 commonsourceibias.n207 0.246418
R15390 commonsourceibias.n477 commonsourceibias.n444 0.246418
R15391 commonsourceibias.n490 commonsourceibias.n440 0.246418
R15392 commonsourceibias.n536 commonsourceibias.n381 0.246418
R15393 commonsourceibias.n418 commonsourceibias.n385 0.246418
R15394 commonsourceibias.n702 commonsourceibias.n669 0.246418
R15395 commonsourceibias.n715 commonsourceibias.n665 0.246418
R15396 commonsourceibias.n612 commonsourceibias.n579 0.246418
R15397 commonsourceibias.n625 commonsourceibias.n575 0.246418
R15398 commonsourceibias.n95 commonsourceibias.n12 0.189894
R15399 commonsourceibias.n95 commonsourceibias.n94 0.189894
R15400 commonsourceibias.n94 commonsourceibias.n93 0.189894
R15401 commonsourceibias.n93 commonsourceibias.n14 0.189894
R15402 commonsourceibias.n88 commonsourceibias.n14 0.189894
R15403 commonsourceibias.n88 commonsourceibias.n87 0.189894
R15404 commonsourceibias.n87 commonsourceibias.n86 0.189894
R15405 commonsourceibias.n86 commonsourceibias.n16 0.189894
R15406 commonsourceibias.n81 commonsourceibias.n16 0.189894
R15407 commonsourceibias.n81 commonsourceibias.n80 0.189894
R15408 commonsourceibias.n80 commonsourceibias.n79 0.189894
R15409 commonsourceibias.n79 commonsourceibias.n19 0.189894
R15410 commonsourceibias.n74 commonsourceibias.n19 0.189894
R15411 commonsourceibias.n74 commonsourceibias.n73 0.189894
R15412 commonsourceibias.n73 commonsourceibias.n72 0.189894
R15413 commonsourceibias.n72 commonsourceibias.n21 0.189894
R15414 commonsourceibias.n67 commonsourceibias.n21 0.189894
R15415 commonsourceibias.n67 commonsourceibias.n66 0.189894
R15416 commonsourceibias.n66 commonsourceibias.n65 0.189894
R15417 commonsourceibias.n65 commonsourceibias.n24 0.189894
R15418 commonsourceibias.n60 commonsourceibias.n24 0.189894
R15419 commonsourceibias.n60 commonsourceibias.n59 0.189894
R15420 commonsourceibias.n59 commonsourceibias.n26 0.189894
R15421 commonsourceibias.n55 commonsourceibias.n26 0.189894
R15422 commonsourceibias.n55 commonsourceibias.n54 0.189894
R15423 commonsourceibias.n54 commonsourceibias.n28 0.189894
R15424 commonsourceibias.n50 commonsourceibias.n28 0.189894
R15425 commonsourceibias.n50 commonsourceibias.n49 0.189894
R15426 commonsourceibias.n49 commonsourceibias.n30 0.189894
R15427 commonsourceibias.n44 commonsourceibias.n30 0.189894
R15428 commonsourceibias.n44 commonsourceibias.n43 0.189894
R15429 commonsourceibias.n43 commonsourceibias.n42 0.189894
R15430 commonsourceibias.n42 commonsourceibias.n32 0.189894
R15431 commonsourceibias.n37 commonsourceibias.n32 0.189894
R15432 commonsourceibias.n37 commonsourceibias.n36 0.189894
R15433 commonsourceibias.n158 commonsourceibias.n117 0.189894
R15434 commonsourceibias.n153 commonsourceibias.n117 0.189894
R15435 commonsourceibias.n153 commonsourceibias.n152 0.189894
R15436 commonsourceibias.n152 commonsourceibias.n119 0.189894
R15437 commonsourceibias.n148 commonsourceibias.n119 0.189894
R15438 commonsourceibias.n148 commonsourceibias.n147 0.189894
R15439 commonsourceibias.n147 commonsourceibias.n121 0.189894
R15440 commonsourceibias.n143 commonsourceibias.n121 0.189894
R15441 commonsourceibias.n143 commonsourceibias.n142 0.189894
R15442 commonsourceibias.n142 commonsourceibias.n123 0.189894
R15443 commonsourceibias.n137 commonsourceibias.n123 0.189894
R15444 commonsourceibias.n137 commonsourceibias.n136 0.189894
R15445 commonsourceibias.n136 commonsourceibias.n135 0.189894
R15446 commonsourceibias.n135 commonsourceibias.n125 0.189894
R15447 commonsourceibias.n130 commonsourceibias.n125 0.189894
R15448 commonsourceibias.n130 commonsourceibias.n129 0.189894
R15449 commonsourceibias.n188 commonsourceibias.n0 0.189894
R15450 commonsourceibias.n188 commonsourceibias.n187 0.189894
R15451 commonsourceibias.n187 commonsourceibias.n186 0.189894
R15452 commonsourceibias.n186 commonsourceibias.n2 0.189894
R15453 commonsourceibias.n181 commonsourceibias.n2 0.189894
R15454 commonsourceibias.n181 commonsourceibias.n180 0.189894
R15455 commonsourceibias.n180 commonsourceibias.n179 0.189894
R15456 commonsourceibias.n179 commonsourceibias.n4 0.189894
R15457 commonsourceibias.n174 commonsourceibias.n4 0.189894
R15458 commonsourceibias.n174 commonsourceibias.n173 0.189894
R15459 commonsourceibias.n173 commonsourceibias.n172 0.189894
R15460 commonsourceibias.n172 commonsourceibias.n7 0.189894
R15461 commonsourceibias.n167 commonsourceibias.n7 0.189894
R15462 commonsourceibias.n167 commonsourceibias.n166 0.189894
R15463 commonsourceibias.n166 commonsourceibias.n165 0.189894
R15464 commonsourceibias.n165 commonsourceibias.n9 0.189894
R15465 commonsourceibias.n160 commonsourceibias.n9 0.189894
R15466 commonsourceibias.n367 commonsourceibias.n284 0.189894
R15467 commonsourceibias.n367 commonsourceibias.n366 0.189894
R15468 commonsourceibias.n366 commonsourceibias.n365 0.189894
R15469 commonsourceibias.n365 commonsourceibias.n286 0.189894
R15470 commonsourceibias.n360 commonsourceibias.n286 0.189894
R15471 commonsourceibias.n360 commonsourceibias.n359 0.189894
R15472 commonsourceibias.n359 commonsourceibias.n358 0.189894
R15473 commonsourceibias.n358 commonsourceibias.n288 0.189894
R15474 commonsourceibias.n353 commonsourceibias.n288 0.189894
R15475 commonsourceibias.n353 commonsourceibias.n352 0.189894
R15476 commonsourceibias.n352 commonsourceibias.n351 0.189894
R15477 commonsourceibias.n351 commonsourceibias.n291 0.189894
R15478 commonsourceibias.n346 commonsourceibias.n291 0.189894
R15479 commonsourceibias.n346 commonsourceibias.n345 0.189894
R15480 commonsourceibias.n345 commonsourceibias.n344 0.189894
R15481 commonsourceibias.n344 commonsourceibias.n293 0.189894
R15482 commonsourceibias.n339 commonsourceibias.n293 0.189894
R15483 commonsourceibias.n339 commonsourceibias.n338 0.189894
R15484 commonsourceibias.n338 commonsourceibias.n337 0.189894
R15485 commonsourceibias.n337 commonsourceibias.n296 0.189894
R15486 commonsourceibias.n332 commonsourceibias.n296 0.189894
R15487 commonsourceibias.n332 commonsourceibias.n331 0.189894
R15488 commonsourceibias.n331 commonsourceibias.n298 0.189894
R15489 commonsourceibias.n327 commonsourceibias.n298 0.189894
R15490 commonsourceibias.n327 commonsourceibias.n326 0.189894
R15491 commonsourceibias.n326 commonsourceibias.n300 0.189894
R15492 commonsourceibias.n322 commonsourceibias.n300 0.189894
R15493 commonsourceibias.n322 commonsourceibias.n321 0.189894
R15494 commonsourceibias.n321 commonsourceibias.n302 0.189894
R15495 commonsourceibias.n316 commonsourceibias.n302 0.189894
R15496 commonsourceibias.n316 commonsourceibias.n315 0.189894
R15497 commonsourceibias.n315 commonsourceibias.n314 0.189894
R15498 commonsourceibias.n314 commonsourceibias.n304 0.189894
R15499 commonsourceibias.n309 commonsourceibias.n304 0.189894
R15500 commonsourceibias.n309 commonsourceibias.n308 0.189894
R15501 commonsourceibias.n277 commonsourceibias.n194 0.189894
R15502 commonsourceibias.n277 commonsourceibias.n276 0.189894
R15503 commonsourceibias.n276 commonsourceibias.n275 0.189894
R15504 commonsourceibias.n275 commonsourceibias.n196 0.189894
R15505 commonsourceibias.n270 commonsourceibias.n196 0.189894
R15506 commonsourceibias.n270 commonsourceibias.n269 0.189894
R15507 commonsourceibias.n269 commonsourceibias.n268 0.189894
R15508 commonsourceibias.n268 commonsourceibias.n198 0.189894
R15509 commonsourceibias.n263 commonsourceibias.n198 0.189894
R15510 commonsourceibias.n263 commonsourceibias.n262 0.189894
R15511 commonsourceibias.n262 commonsourceibias.n261 0.189894
R15512 commonsourceibias.n261 commonsourceibias.n201 0.189894
R15513 commonsourceibias.n256 commonsourceibias.n201 0.189894
R15514 commonsourceibias.n256 commonsourceibias.n255 0.189894
R15515 commonsourceibias.n255 commonsourceibias.n254 0.189894
R15516 commonsourceibias.n254 commonsourceibias.n203 0.189894
R15517 commonsourceibias.n249 commonsourceibias.n203 0.189894
R15518 commonsourceibias.n249 commonsourceibias.n248 0.189894
R15519 commonsourceibias.n248 commonsourceibias.n247 0.189894
R15520 commonsourceibias.n247 commonsourceibias.n206 0.189894
R15521 commonsourceibias.n242 commonsourceibias.n206 0.189894
R15522 commonsourceibias.n242 commonsourceibias.n241 0.189894
R15523 commonsourceibias.n241 commonsourceibias.n208 0.189894
R15524 commonsourceibias.n237 commonsourceibias.n208 0.189894
R15525 commonsourceibias.n237 commonsourceibias.n236 0.189894
R15526 commonsourceibias.n236 commonsourceibias.n210 0.189894
R15527 commonsourceibias.n232 commonsourceibias.n210 0.189894
R15528 commonsourceibias.n232 commonsourceibias.n231 0.189894
R15529 commonsourceibias.n231 commonsourceibias.n212 0.189894
R15530 commonsourceibias.n226 commonsourceibias.n212 0.189894
R15531 commonsourceibias.n226 commonsourceibias.n225 0.189894
R15532 commonsourceibias.n225 commonsourceibias.n224 0.189894
R15533 commonsourceibias.n224 commonsourceibias.n214 0.189894
R15534 commonsourceibias.n219 commonsourceibias.n214 0.189894
R15535 commonsourceibias.n219 commonsourceibias.n218 0.189894
R15536 commonsourceibias.n456 commonsourceibias.n455 0.189894
R15537 commonsourceibias.n456 commonsourceibias.n451 0.189894
R15538 commonsourceibias.n461 commonsourceibias.n451 0.189894
R15539 commonsourceibias.n462 commonsourceibias.n461 0.189894
R15540 commonsourceibias.n463 commonsourceibias.n462 0.189894
R15541 commonsourceibias.n463 commonsourceibias.n449 0.189894
R15542 commonsourceibias.n468 commonsourceibias.n449 0.189894
R15543 commonsourceibias.n469 commonsourceibias.n468 0.189894
R15544 commonsourceibias.n469 commonsourceibias.n447 0.189894
R15545 commonsourceibias.n473 commonsourceibias.n447 0.189894
R15546 commonsourceibias.n474 commonsourceibias.n473 0.189894
R15547 commonsourceibias.n474 commonsourceibias.n445 0.189894
R15548 commonsourceibias.n478 commonsourceibias.n445 0.189894
R15549 commonsourceibias.n479 commonsourceibias.n478 0.189894
R15550 commonsourceibias.n479 commonsourceibias.n443 0.189894
R15551 commonsourceibias.n484 commonsourceibias.n443 0.189894
R15552 commonsourceibias.n485 commonsourceibias.n484 0.189894
R15553 commonsourceibias.n486 commonsourceibias.n485 0.189894
R15554 commonsourceibias.n486 commonsourceibias.n441 0.189894
R15555 commonsourceibias.n492 commonsourceibias.n441 0.189894
R15556 commonsourceibias.n493 commonsourceibias.n492 0.189894
R15557 commonsourceibias.n494 commonsourceibias.n493 0.189894
R15558 commonsourceibias.n494 commonsourceibias.n439 0.189894
R15559 commonsourceibias.n499 commonsourceibias.n439 0.189894
R15560 commonsourceibias.n500 commonsourceibias.n499 0.189894
R15561 commonsourceibias.n501 commonsourceibias.n500 0.189894
R15562 commonsourceibias.n501 commonsourceibias.n437 0.189894
R15563 commonsourceibias.n507 commonsourceibias.n437 0.189894
R15564 commonsourceibias.n508 commonsourceibias.n507 0.189894
R15565 commonsourceibias.n509 commonsourceibias.n508 0.189894
R15566 commonsourceibias.n509 commonsourceibias.n435 0.189894
R15567 commonsourceibias.n514 commonsourceibias.n435 0.189894
R15568 commonsourceibias.n515 commonsourceibias.n514 0.189894
R15569 commonsourceibias.n516 commonsourceibias.n515 0.189894
R15570 commonsourceibias.n516 commonsourceibias.n433 0.189894
R15571 commonsourceibias.n397 commonsourceibias.n396 0.189894
R15572 commonsourceibias.n397 commonsourceibias.n392 0.189894
R15573 commonsourceibias.n402 commonsourceibias.n392 0.189894
R15574 commonsourceibias.n403 commonsourceibias.n402 0.189894
R15575 commonsourceibias.n404 commonsourceibias.n403 0.189894
R15576 commonsourceibias.n404 commonsourceibias.n390 0.189894
R15577 commonsourceibias.n409 commonsourceibias.n390 0.189894
R15578 commonsourceibias.n410 commonsourceibias.n409 0.189894
R15579 commonsourceibias.n410 commonsourceibias.n388 0.189894
R15580 commonsourceibias.n414 commonsourceibias.n388 0.189894
R15581 commonsourceibias.n415 commonsourceibias.n414 0.189894
R15582 commonsourceibias.n415 commonsourceibias.n386 0.189894
R15583 commonsourceibias.n419 commonsourceibias.n386 0.189894
R15584 commonsourceibias.n420 commonsourceibias.n419 0.189894
R15585 commonsourceibias.n420 commonsourceibias.n384 0.189894
R15586 commonsourceibias.n425 commonsourceibias.n384 0.189894
R15587 commonsourceibias.n532 commonsourceibias.n382 0.189894
R15588 commonsourceibias.n538 commonsourceibias.n382 0.189894
R15589 commonsourceibias.n539 commonsourceibias.n538 0.189894
R15590 commonsourceibias.n540 commonsourceibias.n539 0.189894
R15591 commonsourceibias.n540 commonsourceibias.n380 0.189894
R15592 commonsourceibias.n545 commonsourceibias.n380 0.189894
R15593 commonsourceibias.n546 commonsourceibias.n545 0.189894
R15594 commonsourceibias.n547 commonsourceibias.n546 0.189894
R15595 commonsourceibias.n547 commonsourceibias.n378 0.189894
R15596 commonsourceibias.n553 commonsourceibias.n378 0.189894
R15597 commonsourceibias.n554 commonsourceibias.n553 0.189894
R15598 commonsourceibias.n555 commonsourceibias.n554 0.189894
R15599 commonsourceibias.n555 commonsourceibias.n376 0.189894
R15600 commonsourceibias.n560 commonsourceibias.n376 0.189894
R15601 commonsourceibias.n561 commonsourceibias.n560 0.189894
R15602 commonsourceibias.n562 commonsourceibias.n561 0.189894
R15603 commonsourceibias.n562 commonsourceibias.n374 0.189894
R15604 commonsourceibias.n681 commonsourceibias.n680 0.189894
R15605 commonsourceibias.n681 commonsourceibias.n676 0.189894
R15606 commonsourceibias.n686 commonsourceibias.n676 0.189894
R15607 commonsourceibias.n687 commonsourceibias.n686 0.189894
R15608 commonsourceibias.n688 commonsourceibias.n687 0.189894
R15609 commonsourceibias.n688 commonsourceibias.n674 0.189894
R15610 commonsourceibias.n693 commonsourceibias.n674 0.189894
R15611 commonsourceibias.n694 commonsourceibias.n693 0.189894
R15612 commonsourceibias.n694 commonsourceibias.n672 0.189894
R15613 commonsourceibias.n698 commonsourceibias.n672 0.189894
R15614 commonsourceibias.n699 commonsourceibias.n698 0.189894
R15615 commonsourceibias.n699 commonsourceibias.n670 0.189894
R15616 commonsourceibias.n703 commonsourceibias.n670 0.189894
R15617 commonsourceibias.n704 commonsourceibias.n703 0.189894
R15618 commonsourceibias.n704 commonsourceibias.n668 0.189894
R15619 commonsourceibias.n709 commonsourceibias.n668 0.189894
R15620 commonsourceibias.n710 commonsourceibias.n709 0.189894
R15621 commonsourceibias.n711 commonsourceibias.n710 0.189894
R15622 commonsourceibias.n711 commonsourceibias.n666 0.189894
R15623 commonsourceibias.n717 commonsourceibias.n666 0.189894
R15624 commonsourceibias.n718 commonsourceibias.n717 0.189894
R15625 commonsourceibias.n719 commonsourceibias.n718 0.189894
R15626 commonsourceibias.n719 commonsourceibias.n664 0.189894
R15627 commonsourceibias.n724 commonsourceibias.n664 0.189894
R15628 commonsourceibias.n725 commonsourceibias.n724 0.189894
R15629 commonsourceibias.n726 commonsourceibias.n725 0.189894
R15630 commonsourceibias.n726 commonsourceibias.n662 0.189894
R15631 commonsourceibias.n732 commonsourceibias.n662 0.189894
R15632 commonsourceibias.n733 commonsourceibias.n732 0.189894
R15633 commonsourceibias.n734 commonsourceibias.n733 0.189894
R15634 commonsourceibias.n734 commonsourceibias.n660 0.189894
R15635 commonsourceibias.n739 commonsourceibias.n660 0.189894
R15636 commonsourceibias.n740 commonsourceibias.n739 0.189894
R15637 commonsourceibias.n741 commonsourceibias.n740 0.189894
R15638 commonsourceibias.n741 commonsourceibias.n658 0.189894
R15639 commonsourceibias.n591 commonsourceibias.n590 0.189894
R15640 commonsourceibias.n591 commonsourceibias.n586 0.189894
R15641 commonsourceibias.n596 commonsourceibias.n586 0.189894
R15642 commonsourceibias.n597 commonsourceibias.n596 0.189894
R15643 commonsourceibias.n598 commonsourceibias.n597 0.189894
R15644 commonsourceibias.n598 commonsourceibias.n584 0.189894
R15645 commonsourceibias.n603 commonsourceibias.n584 0.189894
R15646 commonsourceibias.n604 commonsourceibias.n603 0.189894
R15647 commonsourceibias.n604 commonsourceibias.n582 0.189894
R15648 commonsourceibias.n608 commonsourceibias.n582 0.189894
R15649 commonsourceibias.n609 commonsourceibias.n608 0.189894
R15650 commonsourceibias.n609 commonsourceibias.n580 0.189894
R15651 commonsourceibias.n613 commonsourceibias.n580 0.189894
R15652 commonsourceibias.n614 commonsourceibias.n613 0.189894
R15653 commonsourceibias.n614 commonsourceibias.n578 0.189894
R15654 commonsourceibias.n619 commonsourceibias.n578 0.189894
R15655 commonsourceibias.n620 commonsourceibias.n619 0.189894
R15656 commonsourceibias.n621 commonsourceibias.n620 0.189894
R15657 commonsourceibias.n621 commonsourceibias.n576 0.189894
R15658 commonsourceibias.n627 commonsourceibias.n576 0.189894
R15659 commonsourceibias.n628 commonsourceibias.n627 0.189894
R15660 commonsourceibias.n629 commonsourceibias.n628 0.189894
R15661 commonsourceibias.n629 commonsourceibias.n574 0.189894
R15662 commonsourceibias.n634 commonsourceibias.n574 0.189894
R15663 commonsourceibias.n635 commonsourceibias.n634 0.189894
R15664 commonsourceibias.n636 commonsourceibias.n635 0.189894
R15665 commonsourceibias.n636 commonsourceibias.n572 0.189894
R15666 commonsourceibias.n642 commonsourceibias.n572 0.189894
R15667 commonsourceibias.n643 commonsourceibias.n642 0.189894
R15668 commonsourceibias.n644 commonsourceibias.n643 0.189894
R15669 commonsourceibias.n644 commonsourceibias.n570 0.189894
R15670 commonsourceibias.n649 commonsourceibias.n570 0.189894
R15671 commonsourceibias.n650 commonsourceibias.n649 0.189894
R15672 commonsourceibias.n651 commonsourceibias.n650 0.189894
R15673 commonsourceibias.n651 commonsourceibias.n568 0.189894
R15674 commonsourceibias.n159 commonsourceibias.n158 0.170955
R15675 commonsourceibias.n160 commonsourceibias.n159 0.170955
R15676 commonsourceibias.n531 commonsourceibias.n425 0.170955
R15677 commonsourceibias.n532 commonsourceibias.n531 0.170955
R15678 CSoutput.n19 CSoutput.t185 184.661
R15679 CSoutput.n78 CSoutput.n77 165.8
R15680 CSoutput.n76 CSoutput.n0 165.8
R15681 CSoutput.n75 CSoutput.n74 165.8
R15682 CSoutput.n73 CSoutput.n72 165.8
R15683 CSoutput.n71 CSoutput.n2 165.8
R15684 CSoutput.n69 CSoutput.n68 165.8
R15685 CSoutput.n67 CSoutput.n3 165.8
R15686 CSoutput.n66 CSoutput.n65 165.8
R15687 CSoutput.n63 CSoutput.n4 165.8
R15688 CSoutput.n61 CSoutput.n60 165.8
R15689 CSoutput.n59 CSoutput.n5 165.8
R15690 CSoutput.n58 CSoutput.n57 165.8
R15691 CSoutput.n55 CSoutput.n6 165.8
R15692 CSoutput.n54 CSoutput.n53 165.8
R15693 CSoutput.n52 CSoutput.n51 165.8
R15694 CSoutput.n50 CSoutput.n8 165.8
R15695 CSoutput.n48 CSoutput.n47 165.8
R15696 CSoutput.n46 CSoutput.n9 165.8
R15697 CSoutput.n45 CSoutput.n44 165.8
R15698 CSoutput.n42 CSoutput.n10 165.8
R15699 CSoutput.n41 CSoutput.n40 165.8
R15700 CSoutput.n39 CSoutput.n38 165.8
R15701 CSoutput.n37 CSoutput.n12 165.8
R15702 CSoutput.n35 CSoutput.n34 165.8
R15703 CSoutput.n33 CSoutput.n13 165.8
R15704 CSoutput.n32 CSoutput.n31 165.8
R15705 CSoutput.n29 CSoutput.n14 165.8
R15706 CSoutput.n28 CSoutput.n27 165.8
R15707 CSoutput.n26 CSoutput.n25 165.8
R15708 CSoutput.n24 CSoutput.n16 165.8
R15709 CSoutput.n22 CSoutput.n21 165.8
R15710 CSoutput.n20 CSoutput.n17 165.8
R15711 CSoutput.n77 CSoutput.t187 162.194
R15712 CSoutput.n18 CSoutput.t182 120.501
R15713 CSoutput.n23 CSoutput.t176 120.501
R15714 CSoutput.n15 CSoutput.t171 120.501
R15715 CSoutput.n30 CSoutput.t183 120.501
R15716 CSoutput.n36 CSoutput.t184 120.501
R15717 CSoutput.n11 CSoutput.t173 120.501
R15718 CSoutput.n43 CSoutput.t169 120.501
R15719 CSoutput.n49 CSoutput.t186 120.501
R15720 CSoutput.n7 CSoutput.t177 120.501
R15721 CSoutput.n56 CSoutput.t179 120.501
R15722 CSoutput.n62 CSoutput.t188 120.501
R15723 CSoutput.n64 CSoutput.t180 120.501
R15724 CSoutput.n70 CSoutput.t181 120.501
R15725 CSoutput.n1 CSoutput.t174 120.501
R15726 CSoutput.n290 CSoutput.n288 103.469
R15727 CSoutput.n278 CSoutput.n276 103.469
R15728 CSoutput.n267 CSoutput.n265 103.469
R15729 CSoutput.n104 CSoutput.n102 103.469
R15730 CSoutput.n92 CSoutput.n90 103.469
R15731 CSoutput.n81 CSoutput.n79 103.469
R15732 CSoutput.n296 CSoutput.n295 103.111
R15733 CSoutput.n294 CSoutput.n293 103.111
R15734 CSoutput.n292 CSoutput.n291 103.111
R15735 CSoutput.n290 CSoutput.n289 103.111
R15736 CSoutput.n286 CSoutput.n285 103.111
R15737 CSoutput.n284 CSoutput.n283 103.111
R15738 CSoutput.n282 CSoutput.n281 103.111
R15739 CSoutput.n280 CSoutput.n279 103.111
R15740 CSoutput.n278 CSoutput.n277 103.111
R15741 CSoutput.n275 CSoutput.n274 103.111
R15742 CSoutput.n273 CSoutput.n272 103.111
R15743 CSoutput.n271 CSoutput.n270 103.111
R15744 CSoutput.n269 CSoutput.n268 103.111
R15745 CSoutput.n267 CSoutput.n266 103.111
R15746 CSoutput.n104 CSoutput.n103 103.111
R15747 CSoutput.n106 CSoutput.n105 103.111
R15748 CSoutput.n108 CSoutput.n107 103.111
R15749 CSoutput.n110 CSoutput.n109 103.111
R15750 CSoutput.n112 CSoutput.n111 103.111
R15751 CSoutput.n92 CSoutput.n91 103.111
R15752 CSoutput.n94 CSoutput.n93 103.111
R15753 CSoutput.n96 CSoutput.n95 103.111
R15754 CSoutput.n98 CSoutput.n97 103.111
R15755 CSoutput.n100 CSoutput.n99 103.111
R15756 CSoutput.n81 CSoutput.n80 103.111
R15757 CSoutput.n83 CSoutput.n82 103.111
R15758 CSoutput.n85 CSoutput.n84 103.111
R15759 CSoutput.n87 CSoutput.n86 103.111
R15760 CSoutput.n89 CSoutput.n88 103.111
R15761 CSoutput.n298 CSoutput.n297 103.111
R15762 CSoutput.n334 CSoutput.n332 81.5057
R15763 CSoutput.n318 CSoutput.n316 81.5057
R15764 CSoutput.n303 CSoutput.n301 81.5057
R15765 CSoutput.n382 CSoutput.n380 81.5057
R15766 CSoutput.n366 CSoutput.n364 81.5057
R15767 CSoutput.n351 CSoutput.n349 81.5057
R15768 CSoutput.n346 CSoutput.n345 80.9324
R15769 CSoutput.n344 CSoutput.n343 80.9324
R15770 CSoutput.n342 CSoutput.n341 80.9324
R15771 CSoutput.n340 CSoutput.n339 80.9324
R15772 CSoutput.n338 CSoutput.n337 80.9324
R15773 CSoutput.n336 CSoutput.n335 80.9324
R15774 CSoutput.n334 CSoutput.n333 80.9324
R15775 CSoutput.n330 CSoutput.n329 80.9324
R15776 CSoutput.n328 CSoutput.n327 80.9324
R15777 CSoutput.n326 CSoutput.n325 80.9324
R15778 CSoutput.n324 CSoutput.n323 80.9324
R15779 CSoutput.n322 CSoutput.n321 80.9324
R15780 CSoutput.n320 CSoutput.n319 80.9324
R15781 CSoutput.n318 CSoutput.n317 80.9324
R15782 CSoutput.n315 CSoutput.n314 80.9324
R15783 CSoutput.n313 CSoutput.n312 80.9324
R15784 CSoutput.n311 CSoutput.n310 80.9324
R15785 CSoutput.n309 CSoutput.n308 80.9324
R15786 CSoutput.n307 CSoutput.n306 80.9324
R15787 CSoutput.n305 CSoutput.n304 80.9324
R15788 CSoutput.n303 CSoutput.n302 80.9324
R15789 CSoutput.n382 CSoutput.n381 80.9324
R15790 CSoutput.n384 CSoutput.n383 80.9324
R15791 CSoutput.n386 CSoutput.n385 80.9324
R15792 CSoutput.n388 CSoutput.n387 80.9324
R15793 CSoutput.n390 CSoutput.n389 80.9324
R15794 CSoutput.n392 CSoutput.n391 80.9324
R15795 CSoutput.n394 CSoutput.n393 80.9324
R15796 CSoutput.n366 CSoutput.n365 80.9324
R15797 CSoutput.n368 CSoutput.n367 80.9324
R15798 CSoutput.n370 CSoutput.n369 80.9324
R15799 CSoutput.n372 CSoutput.n371 80.9324
R15800 CSoutput.n374 CSoutput.n373 80.9324
R15801 CSoutput.n376 CSoutput.n375 80.9324
R15802 CSoutput.n378 CSoutput.n377 80.9324
R15803 CSoutput.n351 CSoutput.n350 80.9324
R15804 CSoutput.n353 CSoutput.n352 80.9324
R15805 CSoutput.n355 CSoutput.n354 80.9324
R15806 CSoutput.n357 CSoutput.n356 80.9324
R15807 CSoutput.n359 CSoutput.n358 80.9324
R15808 CSoutput.n361 CSoutput.n360 80.9324
R15809 CSoutput.n363 CSoutput.n362 80.9324
R15810 CSoutput.n25 CSoutput.n24 48.1486
R15811 CSoutput.n69 CSoutput.n3 48.1486
R15812 CSoutput.n38 CSoutput.n37 48.1486
R15813 CSoutput.n42 CSoutput.n41 48.1486
R15814 CSoutput.n51 CSoutput.n50 48.1486
R15815 CSoutput.n55 CSoutput.n54 48.1486
R15816 CSoutput.n22 CSoutput.n17 46.462
R15817 CSoutput.n72 CSoutput.n71 46.462
R15818 CSoutput.n20 CSoutput.n19 44.9055
R15819 CSoutput.n29 CSoutput.n28 43.7635
R15820 CSoutput.n65 CSoutput.n63 43.7635
R15821 CSoutput.n35 CSoutput.n13 41.7396
R15822 CSoutput.n57 CSoutput.n5 41.7396
R15823 CSoutput.n44 CSoutput.n9 37.0171
R15824 CSoutput.n48 CSoutput.n9 37.0171
R15825 CSoutput.n76 CSoutput.n75 34.9932
R15826 CSoutput.n31 CSoutput.n13 32.2947
R15827 CSoutput.n61 CSoutput.n5 32.2947
R15828 CSoutput.n30 CSoutput.n29 29.6014
R15829 CSoutput.n63 CSoutput.n62 29.6014
R15830 CSoutput.n19 CSoutput.n18 28.4085
R15831 CSoutput.n18 CSoutput.n17 25.1176
R15832 CSoutput.n72 CSoutput.n1 25.1176
R15833 CSoutput.n43 CSoutput.n42 22.0922
R15834 CSoutput.n50 CSoutput.n49 22.0922
R15835 CSoutput.n77 CSoutput.n76 21.8586
R15836 CSoutput.n37 CSoutput.n36 18.9681
R15837 CSoutput.n56 CSoutput.n55 18.9681
R15838 CSoutput.n25 CSoutput.n15 17.6292
R15839 CSoutput.n64 CSoutput.n3 17.6292
R15840 CSoutput.n24 CSoutput.n23 15.844
R15841 CSoutput.n70 CSoutput.n69 15.844
R15842 CSoutput.n38 CSoutput.n11 14.5051
R15843 CSoutput.n54 CSoutput.n7 14.5051
R15844 CSoutput.n397 CSoutput.n78 11.4982
R15845 CSoutput.n41 CSoutput.n11 11.3811
R15846 CSoutput.n51 CSoutput.n7 11.3811
R15847 CSoutput.n23 CSoutput.n22 10.0422
R15848 CSoutput.n71 CSoutput.n70 10.0422
R15849 CSoutput.n287 CSoutput.n275 9.25285
R15850 CSoutput.n101 CSoutput.n89 9.25285
R15851 CSoutput.n331 CSoutput.n315 8.98182
R15852 CSoutput.n379 CSoutput.n363 8.98182
R15853 CSoutput.n348 CSoutput.n300 8.67888
R15854 CSoutput.n28 CSoutput.n15 8.25698
R15855 CSoutput.n65 CSoutput.n64 8.25698
R15856 CSoutput.n300 CSoutput.n299 7.12641
R15857 CSoutput.n114 CSoutput.n113 7.12641
R15858 CSoutput.n36 CSoutput.n35 6.91809
R15859 CSoutput.n57 CSoutput.n56 6.91809
R15860 CSoutput.n348 CSoutput.n347 6.02792
R15861 CSoutput.n396 CSoutput.n395 6.02792
R15862 CSoutput.n347 CSoutput.n346 5.25266
R15863 CSoutput.n331 CSoutput.n330 5.25266
R15864 CSoutput.n395 CSoutput.n394 5.25266
R15865 CSoutput.n379 CSoutput.n378 5.25266
R15866 CSoutput.n299 CSoutput.n298 5.1449
R15867 CSoutput.n287 CSoutput.n286 5.1449
R15868 CSoutput.n113 CSoutput.n112 5.1449
R15869 CSoutput.n101 CSoutput.n100 5.1449
R15870 CSoutput.n397 CSoutput.n114 5.08644
R15871 CSoutput.n205 CSoutput.n158 4.5005
R15872 CSoutput.n174 CSoutput.n158 4.5005
R15873 CSoutput.n169 CSoutput.n153 4.5005
R15874 CSoutput.n169 CSoutput.n155 4.5005
R15875 CSoutput.n169 CSoutput.n152 4.5005
R15876 CSoutput.n169 CSoutput.n156 4.5005
R15877 CSoutput.n169 CSoutput.n151 4.5005
R15878 CSoutput.n169 CSoutput.t189 4.5005
R15879 CSoutput.n169 CSoutput.n150 4.5005
R15880 CSoutput.n169 CSoutput.n157 4.5005
R15881 CSoutput.n169 CSoutput.n158 4.5005
R15882 CSoutput.n167 CSoutput.n153 4.5005
R15883 CSoutput.n167 CSoutput.n155 4.5005
R15884 CSoutput.n167 CSoutput.n152 4.5005
R15885 CSoutput.n167 CSoutput.n156 4.5005
R15886 CSoutput.n167 CSoutput.n151 4.5005
R15887 CSoutput.n167 CSoutput.t189 4.5005
R15888 CSoutput.n167 CSoutput.n150 4.5005
R15889 CSoutput.n167 CSoutput.n157 4.5005
R15890 CSoutput.n167 CSoutput.n158 4.5005
R15891 CSoutput.n166 CSoutput.n153 4.5005
R15892 CSoutput.n166 CSoutput.n155 4.5005
R15893 CSoutput.n166 CSoutput.n152 4.5005
R15894 CSoutput.n166 CSoutput.n156 4.5005
R15895 CSoutput.n166 CSoutput.n151 4.5005
R15896 CSoutput.n166 CSoutput.t189 4.5005
R15897 CSoutput.n166 CSoutput.n150 4.5005
R15898 CSoutput.n166 CSoutput.n157 4.5005
R15899 CSoutput.n166 CSoutput.n158 4.5005
R15900 CSoutput.n251 CSoutput.n153 4.5005
R15901 CSoutput.n251 CSoutput.n155 4.5005
R15902 CSoutput.n251 CSoutput.n152 4.5005
R15903 CSoutput.n251 CSoutput.n156 4.5005
R15904 CSoutput.n251 CSoutput.n151 4.5005
R15905 CSoutput.n251 CSoutput.t189 4.5005
R15906 CSoutput.n251 CSoutput.n150 4.5005
R15907 CSoutput.n251 CSoutput.n157 4.5005
R15908 CSoutput.n251 CSoutput.n158 4.5005
R15909 CSoutput.n249 CSoutput.n153 4.5005
R15910 CSoutput.n249 CSoutput.n155 4.5005
R15911 CSoutput.n249 CSoutput.n152 4.5005
R15912 CSoutput.n249 CSoutput.n156 4.5005
R15913 CSoutput.n249 CSoutput.n151 4.5005
R15914 CSoutput.n249 CSoutput.t189 4.5005
R15915 CSoutput.n249 CSoutput.n150 4.5005
R15916 CSoutput.n249 CSoutput.n157 4.5005
R15917 CSoutput.n247 CSoutput.n153 4.5005
R15918 CSoutput.n247 CSoutput.n155 4.5005
R15919 CSoutput.n247 CSoutput.n152 4.5005
R15920 CSoutput.n247 CSoutput.n156 4.5005
R15921 CSoutput.n247 CSoutput.n151 4.5005
R15922 CSoutput.n247 CSoutput.t189 4.5005
R15923 CSoutput.n247 CSoutput.n150 4.5005
R15924 CSoutput.n247 CSoutput.n157 4.5005
R15925 CSoutput.n177 CSoutput.n153 4.5005
R15926 CSoutput.n177 CSoutput.n155 4.5005
R15927 CSoutput.n177 CSoutput.n152 4.5005
R15928 CSoutput.n177 CSoutput.n156 4.5005
R15929 CSoutput.n177 CSoutput.n151 4.5005
R15930 CSoutput.n177 CSoutput.t189 4.5005
R15931 CSoutput.n177 CSoutput.n150 4.5005
R15932 CSoutput.n177 CSoutput.n157 4.5005
R15933 CSoutput.n177 CSoutput.n158 4.5005
R15934 CSoutput.n176 CSoutput.n153 4.5005
R15935 CSoutput.n176 CSoutput.n155 4.5005
R15936 CSoutput.n176 CSoutput.n152 4.5005
R15937 CSoutput.n176 CSoutput.n156 4.5005
R15938 CSoutput.n176 CSoutput.n151 4.5005
R15939 CSoutput.n176 CSoutput.t189 4.5005
R15940 CSoutput.n176 CSoutput.n150 4.5005
R15941 CSoutput.n176 CSoutput.n157 4.5005
R15942 CSoutput.n176 CSoutput.n158 4.5005
R15943 CSoutput.n180 CSoutput.n153 4.5005
R15944 CSoutput.n180 CSoutput.n155 4.5005
R15945 CSoutput.n180 CSoutput.n152 4.5005
R15946 CSoutput.n180 CSoutput.n156 4.5005
R15947 CSoutput.n180 CSoutput.n151 4.5005
R15948 CSoutput.n180 CSoutput.t189 4.5005
R15949 CSoutput.n180 CSoutput.n150 4.5005
R15950 CSoutput.n180 CSoutput.n157 4.5005
R15951 CSoutput.n180 CSoutput.n158 4.5005
R15952 CSoutput.n179 CSoutput.n153 4.5005
R15953 CSoutput.n179 CSoutput.n155 4.5005
R15954 CSoutput.n179 CSoutput.n152 4.5005
R15955 CSoutput.n179 CSoutput.n156 4.5005
R15956 CSoutput.n179 CSoutput.n151 4.5005
R15957 CSoutput.n179 CSoutput.t189 4.5005
R15958 CSoutput.n179 CSoutput.n150 4.5005
R15959 CSoutput.n179 CSoutput.n157 4.5005
R15960 CSoutput.n179 CSoutput.n158 4.5005
R15961 CSoutput.n162 CSoutput.n153 4.5005
R15962 CSoutput.n162 CSoutput.n155 4.5005
R15963 CSoutput.n162 CSoutput.n152 4.5005
R15964 CSoutput.n162 CSoutput.n156 4.5005
R15965 CSoutput.n162 CSoutput.n151 4.5005
R15966 CSoutput.n162 CSoutput.t189 4.5005
R15967 CSoutput.n162 CSoutput.n150 4.5005
R15968 CSoutput.n162 CSoutput.n157 4.5005
R15969 CSoutput.n162 CSoutput.n158 4.5005
R15970 CSoutput.n254 CSoutput.n153 4.5005
R15971 CSoutput.n254 CSoutput.n155 4.5005
R15972 CSoutput.n254 CSoutput.n152 4.5005
R15973 CSoutput.n254 CSoutput.n156 4.5005
R15974 CSoutput.n254 CSoutput.n151 4.5005
R15975 CSoutput.n254 CSoutput.t189 4.5005
R15976 CSoutput.n254 CSoutput.n150 4.5005
R15977 CSoutput.n254 CSoutput.n157 4.5005
R15978 CSoutput.n254 CSoutput.n158 4.5005
R15979 CSoutput.n241 CSoutput.n212 4.5005
R15980 CSoutput.n241 CSoutput.n218 4.5005
R15981 CSoutput.n199 CSoutput.n188 4.5005
R15982 CSoutput.n199 CSoutput.n190 4.5005
R15983 CSoutput.n199 CSoutput.n187 4.5005
R15984 CSoutput.n199 CSoutput.n191 4.5005
R15985 CSoutput.n199 CSoutput.n186 4.5005
R15986 CSoutput.n199 CSoutput.t168 4.5005
R15987 CSoutput.n199 CSoutput.n185 4.5005
R15988 CSoutput.n199 CSoutput.n192 4.5005
R15989 CSoutput.n241 CSoutput.n199 4.5005
R15990 CSoutput.n220 CSoutput.n188 4.5005
R15991 CSoutput.n220 CSoutput.n190 4.5005
R15992 CSoutput.n220 CSoutput.n187 4.5005
R15993 CSoutput.n220 CSoutput.n191 4.5005
R15994 CSoutput.n220 CSoutput.n186 4.5005
R15995 CSoutput.n220 CSoutput.t168 4.5005
R15996 CSoutput.n220 CSoutput.n185 4.5005
R15997 CSoutput.n220 CSoutput.n192 4.5005
R15998 CSoutput.n241 CSoutput.n220 4.5005
R15999 CSoutput.n198 CSoutput.n188 4.5005
R16000 CSoutput.n198 CSoutput.n190 4.5005
R16001 CSoutput.n198 CSoutput.n187 4.5005
R16002 CSoutput.n198 CSoutput.n191 4.5005
R16003 CSoutput.n198 CSoutput.n186 4.5005
R16004 CSoutput.n198 CSoutput.t168 4.5005
R16005 CSoutput.n198 CSoutput.n185 4.5005
R16006 CSoutput.n198 CSoutput.n192 4.5005
R16007 CSoutput.n241 CSoutput.n198 4.5005
R16008 CSoutput.n222 CSoutput.n188 4.5005
R16009 CSoutput.n222 CSoutput.n190 4.5005
R16010 CSoutput.n222 CSoutput.n187 4.5005
R16011 CSoutput.n222 CSoutput.n191 4.5005
R16012 CSoutput.n222 CSoutput.n186 4.5005
R16013 CSoutput.n222 CSoutput.t168 4.5005
R16014 CSoutput.n222 CSoutput.n185 4.5005
R16015 CSoutput.n222 CSoutput.n192 4.5005
R16016 CSoutput.n241 CSoutput.n222 4.5005
R16017 CSoutput.n188 CSoutput.n183 4.5005
R16018 CSoutput.n190 CSoutput.n183 4.5005
R16019 CSoutput.n187 CSoutput.n183 4.5005
R16020 CSoutput.n191 CSoutput.n183 4.5005
R16021 CSoutput.n186 CSoutput.n183 4.5005
R16022 CSoutput.t168 CSoutput.n183 4.5005
R16023 CSoutput.n185 CSoutput.n183 4.5005
R16024 CSoutput.n192 CSoutput.n183 4.5005
R16025 CSoutput.n244 CSoutput.n188 4.5005
R16026 CSoutput.n244 CSoutput.n190 4.5005
R16027 CSoutput.n244 CSoutput.n187 4.5005
R16028 CSoutput.n244 CSoutput.n191 4.5005
R16029 CSoutput.n244 CSoutput.n186 4.5005
R16030 CSoutput.n244 CSoutput.t168 4.5005
R16031 CSoutput.n244 CSoutput.n185 4.5005
R16032 CSoutput.n244 CSoutput.n192 4.5005
R16033 CSoutput.n242 CSoutput.n188 4.5005
R16034 CSoutput.n242 CSoutput.n190 4.5005
R16035 CSoutput.n242 CSoutput.n187 4.5005
R16036 CSoutput.n242 CSoutput.n191 4.5005
R16037 CSoutput.n242 CSoutput.n186 4.5005
R16038 CSoutput.n242 CSoutput.t168 4.5005
R16039 CSoutput.n242 CSoutput.n185 4.5005
R16040 CSoutput.n242 CSoutput.n192 4.5005
R16041 CSoutput.n242 CSoutput.n241 4.5005
R16042 CSoutput.n224 CSoutput.n188 4.5005
R16043 CSoutput.n224 CSoutput.n190 4.5005
R16044 CSoutput.n224 CSoutput.n187 4.5005
R16045 CSoutput.n224 CSoutput.n191 4.5005
R16046 CSoutput.n224 CSoutput.n186 4.5005
R16047 CSoutput.n224 CSoutput.t168 4.5005
R16048 CSoutput.n224 CSoutput.n185 4.5005
R16049 CSoutput.n224 CSoutput.n192 4.5005
R16050 CSoutput.n241 CSoutput.n224 4.5005
R16051 CSoutput.n196 CSoutput.n188 4.5005
R16052 CSoutput.n196 CSoutput.n190 4.5005
R16053 CSoutput.n196 CSoutput.n187 4.5005
R16054 CSoutput.n196 CSoutput.n191 4.5005
R16055 CSoutput.n196 CSoutput.n186 4.5005
R16056 CSoutput.n196 CSoutput.t168 4.5005
R16057 CSoutput.n196 CSoutput.n185 4.5005
R16058 CSoutput.n196 CSoutput.n192 4.5005
R16059 CSoutput.n241 CSoutput.n196 4.5005
R16060 CSoutput.n226 CSoutput.n188 4.5005
R16061 CSoutput.n226 CSoutput.n190 4.5005
R16062 CSoutput.n226 CSoutput.n187 4.5005
R16063 CSoutput.n226 CSoutput.n191 4.5005
R16064 CSoutput.n226 CSoutput.n186 4.5005
R16065 CSoutput.n226 CSoutput.t168 4.5005
R16066 CSoutput.n226 CSoutput.n185 4.5005
R16067 CSoutput.n226 CSoutput.n192 4.5005
R16068 CSoutput.n241 CSoutput.n226 4.5005
R16069 CSoutput.n195 CSoutput.n188 4.5005
R16070 CSoutput.n195 CSoutput.n190 4.5005
R16071 CSoutput.n195 CSoutput.n187 4.5005
R16072 CSoutput.n195 CSoutput.n191 4.5005
R16073 CSoutput.n195 CSoutput.n186 4.5005
R16074 CSoutput.n195 CSoutput.t168 4.5005
R16075 CSoutput.n195 CSoutput.n185 4.5005
R16076 CSoutput.n195 CSoutput.n192 4.5005
R16077 CSoutput.n241 CSoutput.n195 4.5005
R16078 CSoutput.n240 CSoutput.n188 4.5005
R16079 CSoutput.n240 CSoutput.n190 4.5005
R16080 CSoutput.n240 CSoutput.n187 4.5005
R16081 CSoutput.n240 CSoutput.n191 4.5005
R16082 CSoutput.n240 CSoutput.n186 4.5005
R16083 CSoutput.n240 CSoutput.t168 4.5005
R16084 CSoutput.n240 CSoutput.n185 4.5005
R16085 CSoutput.n240 CSoutput.n192 4.5005
R16086 CSoutput.n241 CSoutput.n240 4.5005
R16087 CSoutput.n239 CSoutput.n124 4.5005
R16088 CSoutput.n140 CSoutput.n124 4.5005
R16089 CSoutput.n135 CSoutput.n119 4.5005
R16090 CSoutput.n135 CSoutput.n121 4.5005
R16091 CSoutput.n135 CSoutput.n118 4.5005
R16092 CSoutput.n135 CSoutput.n122 4.5005
R16093 CSoutput.n135 CSoutput.n117 4.5005
R16094 CSoutput.n135 CSoutput.t175 4.5005
R16095 CSoutput.n135 CSoutput.n116 4.5005
R16096 CSoutput.n135 CSoutput.n123 4.5005
R16097 CSoutput.n135 CSoutput.n124 4.5005
R16098 CSoutput.n133 CSoutput.n119 4.5005
R16099 CSoutput.n133 CSoutput.n121 4.5005
R16100 CSoutput.n133 CSoutput.n118 4.5005
R16101 CSoutput.n133 CSoutput.n122 4.5005
R16102 CSoutput.n133 CSoutput.n117 4.5005
R16103 CSoutput.n133 CSoutput.t175 4.5005
R16104 CSoutput.n133 CSoutput.n116 4.5005
R16105 CSoutput.n133 CSoutput.n123 4.5005
R16106 CSoutput.n133 CSoutput.n124 4.5005
R16107 CSoutput.n132 CSoutput.n119 4.5005
R16108 CSoutput.n132 CSoutput.n121 4.5005
R16109 CSoutput.n132 CSoutput.n118 4.5005
R16110 CSoutput.n132 CSoutput.n122 4.5005
R16111 CSoutput.n132 CSoutput.n117 4.5005
R16112 CSoutput.n132 CSoutput.t175 4.5005
R16113 CSoutput.n132 CSoutput.n116 4.5005
R16114 CSoutput.n132 CSoutput.n123 4.5005
R16115 CSoutput.n132 CSoutput.n124 4.5005
R16116 CSoutput.n261 CSoutput.n119 4.5005
R16117 CSoutput.n261 CSoutput.n121 4.5005
R16118 CSoutput.n261 CSoutput.n118 4.5005
R16119 CSoutput.n261 CSoutput.n122 4.5005
R16120 CSoutput.n261 CSoutput.n117 4.5005
R16121 CSoutput.n261 CSoutput.t175 4.5005
R16122 CSoutput.n261 CSoutput.n116 4.5005
R16123 CSoutput.n261 CSoutput.n123 4.5005
R16124 CSoutput.n261 CSoutput.n124 4.5005
R16125 CSoutput.n259 CSoutput.n119 4.5005
R16126 CSoutput.n259 CSoutput.n121 4.5005
R16127 CSoutput.n259 CSoutput.n118 4.5005
R16128 CSoutput.n259 CSoutput.n122 4.5005
R16129 CSoutput.n259 CSoutput.n117 4.5005
R16130 CSoutput.n259 CSoutput.t175 4.5005
R16131 CSoutput.n259 CSoutput.n116 4.5005
R16132 CSoutput.n259 CSoutput.n123 4.5005
R16133 CSoutput.n257 CSoutput.n119 4.5005
R16134 CSoutput.n257 CSoutput.n121 4.5005
R16135 CSoutput.n257 CSoutput.n118 4.5005
R16136 CSoutput.n257 CSoutput.n122 4.5005
R16137 CSoutput.n257 CSoutput.n117 4.5005
R16138 CSoutput.n257 CSoutput.t175 4.5005
R16139 CSoutput.n257 CSoutput.n116 4.5005
R16140 CSoutput.n257 CSoutput.n123 4.5005
R16141 CSoutput.n143 CSoutput.n119 4.5005
R16142 CSoutput.n143 CSoutput.n121 4.5005
R16143 CSoutput.n143 CSoutput.n118 4.5005
R16144 CSoutput.n143 CSoutput.n122 4.5005
R16145 CSoutput.n143 CSoutput.n117 4.5005
R16146 CSoutput.n143 CSoutput.t175 4.5005
R16147 CSoutput.n143 CSoutput.n116 4.5005
R16148 CSoutput.n143 CSoutput.n123 4.5005
R16149 CSoutput.n143 CSoutput.n124 4.5005
R16150 CSoutput.n142 CSoutput.n119 4.5005
R16151 CSoutput.n142 CSoutput.n121 4.5005
R16152 CSoutput.n142 CSoutput.n118 4.5005
R16153 CSoutput.n142 CSoutput.n122 4.5005
R16154 CSoutput.n142 CSoutput.n117 4.5005
R16155 CSoutput.n142 CSoutput.t175 4.5005
R16156 CSoutput.n142 CSoutput.n116 4.5005
R16157 CSoutput.n142 CSoutput.n123 4.5005
R16158 CSoutput.n142 CSoutput.n124 4.5005
R16159 CSoutput.n146 CSoutput.n119 4.5005
R16160 CSoutput.n146 CSoutput.n121 4.5005
R16161 CSoutput.n146 CSoutput.n118 4.5005
R16162 CSoutput.n146 CSoutput.n122 4.5005
R16163 CSoutput.n146 CSoutput.n117 4.5005
R16164 CSoutput.n146 CSoutput.t175 4.5005
R16165 CSoutput.n146 CSoutput.n116 4.5005
R16166 CSoutput.n146 CSoutput.n123 4.5005
R16167 CSoutput.n146 CSoutput.n124 4.5005
R16168 CSoutput.n145 CSoutput.n119 4.5005
R16169 CSoutput.n145 CSoutput.n121 4.5005
R16170 CSoutput.n145 CSoutput.n118 4.5005
R16171 CSoutput.n145 CSoutput.n122 4.5005
R16172 CSoutput.n145 CSoutput.n117 4.5005
R16173 CSoutput.n145 CSoutput.t175 4.5005
R16174 CSoutput.n145 CSoutput.n116 4.5005
R16175 CSoutput.n145 CSoutput.n123 4.5005
R16176 CSoutput.n145 CSoutput.n124 4.5005
R16177 CSoutput.n128 CSoutput.n119 4.5005
R16178 CSoutput.n128 CSoutput.n121 4.5005
R16179 CSoutput.n128 CSoutput.n118 4.5005
R16180 CSoutput.n128 CSoutput.n122 4.5005
R16181 CSoutput.n128 CSoutput.n117 4.5005
R16182 CSoutput.n128 CSoutput.t175 4.5005
R16183 CSoutput.n128 CSoutput.n116 4.5005
R16184 CSoutput.n128 CSoutput.n123 4.5005
R16185 CSoutput.n128 CSoutput.n124 4.5005
R16186 CSoutput.n264 CSoutput.n119 4.5005
R16187 CSoutput.n264 CSoutput.n121 4.5005
R16188 CSoutput.n264 CSoutput.n118 4.5005
R16189 CSoutput.n264 CSoutput.n122 4.5005
R16190 CSoutput.n264 CSoutput.n117 4.5005
R16191 CSoutput.n264 CSoutput.t175 4.5005
R16192 CSoutput.n264 CSoutput.n116 4.5005
R16193 CSoutput.n264 CSoutput.n123 4.5005
R16194 CSoutput.n264 CSoutput.n124 4.5005
R16195 CSoutput.n299 CSoutput.n287 4.10845
R16196 CSoutput.n113 CSoutput.n101 4.10845
R16197 CSoutput.n297 CSoutput.t146 4.06363
R16198 CSoutput.n297 CSoutput.t140 4.06363
R16199 CSoutput.n295 CSoutput.t130 4.06363
R16200 CSoutput.n295 CSoutput.t165 4.06363
R16201 CSoutput.n293 CSoutput.t123 4.06363
R16202 CSoutput.n293 CSoutput.t148 4.06363
R16203 CSoutput.n291 CSoutput.t122 4.06363
R16204 CSoutput.n291 CSoutput.t102 4.06363
R16205 CSoutput.n289 CSoutput.t150 4.06363
R16206 CSoutput.n289 CSoutput.t96 4.06363
R16207 CSoutput.n288 CSoutput.t161 4.06363
R16208 CSoutput.n288 CSoutput.t162 4.06363
R16209 CSoutput.n285 CSoutput.t113 4.06363
R16210 CSoutput.n285 CSoutput.t133 4.06363
R16211 CSoutput.n283 CSoutput.t160 4.06363
R16212 CSoutput.n283 CSoutput.t99 4.06363
R16213 CSoutput.n281 CSoutput.t137 4.06363
R16214 CSoutput.n281 CSoutput.t114 4.06363
R16215 CSoutput.n279 CSoutput.t97 4.06363
R16216 CSoutput.n279 CSoutput.t139 4.06363
R16217 CSoutput.n277 CSoutput.t116 4.06363
R16218 CSoutput.n277 CSoutput.t109 4.06363
R16219 CSoutput.n276 CSoutput.t144 4.06363
R16220 CSoutput.n276 CSoutput.t145 4.06363
R16221 CSoutput.n274 CSoutput.t115 4.06363
R16222 CSoutput.n274 CSoutput.t153 4.06363
R16223 CSoutput.n272 CSoutput.t120 4.06363
R16224 CSoutput.n272 CSoutput.t107 4.06363
R16225 CSoutput.n270 CSoutput.t147 4.06363
R16226 CSoutput.n270 CSoutput.t126 4.06363
R16227 CSoutput.n268 CSoutput.t136 4.06363
R16228 CSoutput.n268 CSoutput.t101 4.06363
R16229 CSoutput.n266 CSoutput.t98 4.06363
R16230 CSoutput.n266 CSoutput.t111 4.06363
R16231 CSoutput.n265 CSoutput.t138 4.06363
R16232 CSoutput.n265 CSoutput.t103 4.06363
R16233 CSoutput.n102 CSoutput.t125 4.06363
R16234 CSoutput.n102 CSoutput.t142 4.06363
R16235 CSoutput.n103 CSoutput.t157 4.06363
R16236 CSoutput.n103 CSoutput.t135 4.06363
R16237 CSoutput.n105 CSoutput.t124 4.06363
R16238 CSoutput.n105 CSoutput.t100 4.06363
R16239 CSoutput.n107 CSoutput.t156 4.06363
R16240 CSoutput.n107 CSoutput.t155 4.06363
R16241 CSoutput.n109 CSoutput.t110 4.06363
R16242 CSoutput.n109 CSoutput.t166 4.06363
R16243 CSoutput.n111 CSoutput.t128 4.06363
R16244 CSoutput.n111 CSoutput.t117 4.06363
R16245 CSoutput.n90 CSoutput.t119 4.06363
R16246 CSoutput.n90 CSoutput.t149 4.06363
R16247 CSoutput.n91 CSoutput.t132 4.06363
R16248 CSoutput.n91 CSoutput.t163 4.06363
R16249 CSoutput.n93 CSoutput.t106 4.06363
R16250 CSoutput.n93 CSoutput.t151 4.06363
R16251 CSoutput.n95 CSoutput.t131 4.06363
R16252 CSoutput.n95 CSoutput.t129 4.06363
R16253 CSoutput.n97 CSoutput.t159 4.06363
R16254 CSoutput.n97 CSoutput.t141 4.06363
R16255 CSoutput.n99 CSoutput.t154 4.06363
R16256 CSoutput.n99 CSoutput.t167 4.06363
R16257 CSoutput.n79 CSoutput.t134 4.06363
R16258 CSoutput.n79 CSoutput.t105 4.06363
R16259 CSoutput.n80 CSoutput.t112 4.06363
R16260 CSoutput.n80 CSoutput.t143 4.06363
R16261 CSoutput.n82 CSoutput.t152 4.06363
R16262 CSoutput.n82 CSoutput.t158 4.06363
R16263 CSoutput.n84 CSoutput.t127 4.06363
R16264 CSoutput.n84 CSoutput.t164 4.06363
R16265 CSoutput.n86 CSoutput.t118 4.06363
R16266 CSoutput.n86 CSoutput.t121 4.06363
R16267 CSoutput.n88 CSoutput.t104 4.06363
R16268 CSoutput.n88 CSoutput.t108 4.06363
R16269 CSoutput.n44 CSoutput.n43 3.79402
R16270 CSoutput.n49 CSoutput.n48 3.79402
R16271 CSoutput.n347 CSoutput.n331 3.72967
R16272 CSoutput.n395 CSoutput.n379 3.72967
R16273 CSoutput.n397 CSoutput.n396 3.57343
R16274 CSoutput.n396 CSoutput.n348 3.08965
R16275 CSoutput.n345 CSoutput.t29 2.82907
R16276 CSoutput.n345 CSoutput.t19 2.82907
R16277 CSoutput.n343 CSoutput.t10 2.82907
R16278 CSoutput.n343 CSoutput.t80 2.82907
R16279 CSoutput.n341 CSoutput.t22 2.82907
R16280 CSoutput.n341 CSoutput.t26 2.82907
R16281 CSoutput.n339 CSoutput.t21 2.82907
R16282 CSoutput.n339 CSoutput.t95 2.82907
R16283 CSoutput.n337 CSoutput.t40 2.82907
R16284 CSoutput.n337 CSoutput.t13 2.82907
R16285 CSoutput.n335 CSoutput.t4 2.82907
R16286 CSoutput.n335 CSoutput.t69 2.82907
R16287 CSoutput.n333 CSoutput.t31 2.82907
R16288 CSoutput.n333 CSoutput.t35 2.82907
R16289 CSoutput.n332 CSoutput.t12 2.82907
R16290 CSoutput.n332 CSoutput.t84 2.82907
R16291 CSoutput.n329 CSoutput.t66 2.82907
R16292 CSoutput.n329 CSoutput.t47 2.82907
R16293 CSoutput.n327 CSoutput.t48 2.82907
R16294 CSoutput.n327 CSoutput.t54 2.82907
R16295 CSoutput.n325 CSoutput.t3 2.82907
R16296 CSoutput.n325 CSoutput.t67 2.82907
R16297 CSoutput.n323 CSoutput.t65 2.82907
R16298 CSoutput.n323 CSoutput.t46 2.82907
R16299 CSoutput.n321 CSoutput.t82 2.82907
R16300 CSoutput.n321 CSoutput.t1 2.82907
R16301 CSoutput.n319 CSoutput.t2 2.82907
R16302 CSoutput.n319 CSoutput.t74 2.82907
R16303 CSoutput.n317 CSoutput.t11 2.82907
R16304 CSoutput.n317 CSoutput.t81 2.82907
R16305 CSoutput.n316 CSoutput.t88 2.82907
R16306 CSoutput.n316 CSoutput.t0 2.82907
R16307 CSoutput.n314 CSoutput.t7 2.82907
R16308 CSoutput.n314 CSoutput.t30 2.82907
R16309 CSoutput.n312 CSoutput.t18 2.82907
R16310 CSoutput.n312 CSoutput.t43 2.82907
R16311 CSoutput.n310 CSoutput.t53 2.82907
R16312 CSoutput.n310 CSoutput.t63 2.82907
R16313 CSoutput.n308 CSoutput.t41 2.82907
R16314 CSoutput.n308 CSoutput.t83 2.82907
R16315 CSoutput.n306 CSoutput.t57 2.82907
R16316 CSoutput.n306 CSoutput.t34 2.82907
R16317 CSoutput.n304 CSoutput.t23 2.82907
R16318 CSoutput.n304 CSoutput.t42 2.82907
R16319 CSoutput.n302 CSoutput.t33 2.82907
R16320 CSoutput.n302 CSoutput.t38 2.82907
R16321 CSoutput.n301 CSoutput.t39 2.82907
R16322 CSoutput.n301 CSoutput.t92 2.82907
R16323 CSoutput.n380 CSoutput.t52 2.82907
R16324 CSoutput.n380 CSoutput.t77 2.82907
R16325 CSoutput.n381 CSoutput.t24 2.82907
R16326 CSoutput.n381 CSoutput.t37 2.82907
R16327 CSoutput.n383 CSoutput.t44 2.82907
R16328 CSoutput.n383 CSoutput.t58 2.82907
R16329 CSoutput.n385 CSoutput.t78 2.82907
R16330 CSoutput.n385 CSoutput.t49 2.82907
R16331 CSoutput.n387 CSoutput.t56 2.82907
R16332 CSoutput.n387 CSoutput.t89 2.82907
R16333 CSoutput.n389 CSoutput.t6 2.82907
R16334 CSoutput.n389 CSoutput.t27 2.82907
R16335 CSoutput.n391 CSoutput.t50 2.82907
R16336 CSoutput.n391 CSoutput.t72 2.82907
R16337 CSoutput.n393 CSoutput.t85 2.82907
R16338 CSoutput.n393 CSoutput.t14 2.82907
R16339 CSoutput.n364 CSoutput.t15 2.82907
R16340 CSoutput.n364 CSoutput.t8 2.82907
R16341 CSoutput.n365 CSoutput.t5 2.82907
R16342 CSoutput.n365 CSoutput.t93 2.82907
R16343 CSoutput.n367 CSoutput.t94 2.82907
R16344 CSoutput.n367 CSoutput.t16 2.82907
R16345 CSoutput.n369 CSoutput.t17 2.82907
R16346 CSoutput.n369 CSoutput.t59 2.82907
R16347 CSoutput.n371 CSoutput.t60 2.82907
R16348 CSoutput.n371 CSoutput.t87 2.82907
R16349 CSoutput.n373 CSoutput.t90 2.82907
R16350 CSoutput.n373 CSoutput.t79 2.82907
R16351 CSoutput.n375 CSoutput.t73 2.82907
R16352 CSoutput.n375 CSoutput.t61 2.82907
R16353 CSoutput.n377 CSoutput.t62 2.82907
R16354 CSoutput.n377 CSoutput.t91 2.82907
R16355 CSoutput.n349 CSoutput.t25 2.82907
R16356 CSoutput.n349 CSoutput.t68 2.82907
R16357 CSoutput.n350 CSoutput.t64 2.82907
R16358 CSoutput.n350 CSoutput.t45 2.82907
R16359 CSoutput.n352 CSoutput.t71 2.82907
R16360 CSoutput.n352 CSoutput.t36 2.82907
R16361 CSoutput.n354 CSoutput.t55 2.82907
R16362 CSoutput.n354 CSoutput.t86 2.82907
R16363 CSoutput.n356 CSoutput.t20 2.82907
R16364 CSoutput.n356 CSoutput.t70 2.82907
R16365 CSoutput.n358 CSoutput.t9 2.82907
R16366 CSoutput.n358 CSoutput.t76 2.82907
R16367 CSoutput.n360 CSoutput.t75 2.82907
R16368 CSoutput.n360 CSoutput.t32 2.82907
R16369 CSoutput.n362 CSoutput.t51 2.82907
R16370 CSoutput.n362 CSoutput.t28 2.82907
R16371 CSoutput.n300 CSoutput.n114 2.78353
R16372 CSoutput.n75 CSoutput.n1 2.45513
R16373 CSoutput.n205 CSoutput.n203 2.251
R16374 CSoutput.n205 CSoutput.n202 2.251
R16375 CSoutput.n205 CSoutput.n201 2.251
R16376 CSoutput.n205 CSoutput.n200 2.251
R16377 CSoutput.n174 CSoutput.n173 2.251
R16378 CSoutput.n174 CSoutput.n172 2.251
R16379 CSoutput.n174 CSoutput.n171 2.251
R16380 CSoutput.n174 CSoutput.n170 2.251
R16381 CSoutput.n247 CSoutput.n246 2.251
R16382 CSoutput.n212 CSoutput.n210 2.251
R16383 CSoutput.n212 CSoutput.n209 2.251
R16384 CSoutput.n212 CSoutput.n208 2.251
R16385 CSoutput.n230 CSoutput.n212 2.251
R16386 CSoutput.n218 CSoutput.n217 2.251
R16387 CSoutput.n218 CSoutput.n216 2.251
R16388 CSoutput.n218 CSoutput.n215 2.251
R16389 CSoutput.n218 CSoutput.n214 2.251
R16390 CSoutput.n244 CSoutput.n184 2.251
R16391 CSoutput.n239 CSoutput.n237 2.251
R16392 CSoutput.n239 CSoutput.n236 2.251
R16393 CSoutput.n239 CSoutput.n235 2.251
R16394 CSoutput.n239 CSoutput.n234 2.251
R16395 CSoutput.n140 CSoutput.n139 2.251
R16396 CSoutput.n140 CSoutput.n138 2.251
R16397 CSoutput.n140 CSoutput.n137 2.251
R16398 CSoutput.n140 CSoutput.n136 2.251
R16399 CSoutput.n257 CSoutput.n256 2.251
R16400 CSoutput.n174 CSoutput.n154 2.2505
R16401 CSoutput.n169 CSoutput.n154 2.2505
R16402 CSoutput.n167 CSoutput.n154 2.2505
R16403 CSoutput.n166 CSoutput.n154 2.2505
R16404 CSoutput.n251 CSoutput.n154 2.2505
R16405 CSoutput.n249 CSoutput.n154 2.2505
R16406 CSoutput.n247 CSoutput.n154 2.2505
R16407 CSoutput.n177 CSoutput.n154 2.2505
R16408 CSoutput.n176 CSoutput.n154 2.2505
R16409 CSoutput.n180 CSoutput.n154 2.2505
R16410 CSoutput.n179 CSoutput.n154 2.2505
R16411 CSoutput.n162 CSoutput.n154 2.2505
R16412 CSoutput.n254 CSoutput.n154 2.2505
R16413 CSoutput.n254 CSoutput.n253 2.2505
R16414 CSoutput.n218 CSoutput.n189 2.2505
R16415 CSoutput.n199 CSoutput.n189 2.2505
R16416 CSoutput.n220 CSoutput.n189 2.2505
R16417 CSoutput.n198 CSoutput.n189 2.2505
R16418 CSoutput.n222 CSoutput.n189 2.2505
R16419 CSoutput.n189 CSoutput.n183 2.2505
R16420 CSoutput.n244 CSoutput.n189 2.2505
R16421 CSoutput.n242 CSoutput.n189 2.2505
R16422 CSoutput.n224 CSoutput.n189 2.2505
R16423 CSoutput.n196 CSoutput.n189 2.2505
R16424 CSoutput.n226 CSoutput.n189 2.2505
R16425 CSoutput.n195 CSoutput.n189 2.2505
R16426 CSoutput.n240 CSoutput.n189 2.2505
R16427 CSoutput.n240 CSoutput.n193 2.2505
R16428 CSoutput.n140 CSoutput.n120 2.2505
R16429 CSoutput.n135 CSoutput.n120 2.2505
R16430 CSoutput.n133 CSoutput.n120 2.2505
R16431 CSoutput.n132 CSoutput.n120 2.2505
R16432 CSoutput.n261 CSoutput.n120 2.2505
R16433 CSoutput.n259 CSoutput.n120 2.2505
R16434 CSoutput.n257 CSoutput.n120 2.2505
R16435 CSoutput.n143 CSoutput.n120 2.2505
R16436 CSoutput.n142 CSoutput.n120 2.2505
R16437 CSoutput.n146 CSoutput.n120 2.2505
R16438 CSoutput.n145 CSoutput.n120 2.2505
R16439 CSoutput.n128 CSoutput.n120 2.2505
R16440 CSoutput.n264 CSoutput.n120 2.2505
R16441 CSoutput.n264 CSoutput.n263 2.2505
R16442 CSoutput.n182 CSoutput.n175 2.25024
R16443 CSoutput.n182 CSoutput.n168 2.25024
R16444 CSoutput.n250 CSoutput.n182 2.25024
R16445 CSoutput.n182 CSoutput.n178 2.25024
R16446 CSoutput.n182 CSoutput.n181 2.25024
R16447 CSoutput.n182 CSoutput.n149 2.25024
R16448 CSoutput.n232 CSoutput.n229 2.25024
R16449 CSoutput.n232 CSoutput.n228 2.25024
R16450 CSoutput.n232 CSoutput.n227 2.25024
R16451 CSoutput.n232 CSoutput.n194 2.25024
R16452 CSoutput.n232 CSoutput.n231 2.25024
R16453 CSoutput.n233 CSoutput.n232 2.25024
R16454 CSoutput.n148 CSoutput.n141 2.25024
R16455 CSoutput.n148 CSoutput.n134 2.25024
R16456 CSoutput.n260 CSoutput.n148 2.25024
R16457 CSoutput.n148 CSoutput.n144 2.25024
R16458 CSoutput.n148 CSoutput.n147 2.25024
R16459 CSoutput.n148 CSoutput.n115 2.25024
R16460 CSoutput.n249 CSoutput.n159 1.50111
R16461 CSoutput.n197 CSoutput.n183 1.50111
R16462 CSoutput.n259 CSoutput.n125 1.50111
R16463 CSoutput.n205 CSoutput.n204 1.501
R16464 CSoutput.n212 CSoutput.n211 1.501
R16465 CSoutput.n239 CSoutput.n238 1.501
R16466 CSoutput.n253 CSoutput.n164 1.12536
R16467 CSoutput.n253 CSoutput.n165 1.12536
R16468 CSoutput.n253 CSoutput.n252 1.12536
R16469 CSoutput.n213 CSoutput.n193 1.12536
R16470 CSoutput.n219 CSoutput.n193 1.12536
R16471 CSoutput.n221 CSoutput.n193 1.12536
R16472 CSoutput.n263 CSoutput.n130 1.12536
R16473 CSoutput.n263 CSoutput.n131 1.12536
R16474 CSoutput.n263 CSoutput.n262 1.12536
R16475 CSoutput.n253 CSoutput.n160 1.12536
R16476 CSoutput.n253 CSoutput.n161 1.12536
R16477 CSoutput.n253 CSoutput.n163 1.12536
R16478 CSoutput.n243 CSoutput.n193 1.12536
R16479 CSoutput.n223 CSoutput.n193 1.12536
R16480 CSoutput.n225 CSoutput.n193 1.12536
R16481 CSoutput.n263 CSoutput.n126 1.12536
R16482 CSoutput.n263 CSoutput.n127 1.12536
R16483 CSoutput.n263 CSoutput.n129 1.12536
R16484 CSoutput.n31 CSoutput.n30 0.669944
R16485 CSoutput.n62 CSoutput.n61 0.669944
R16486 CSoutput.n336 CSoutput.n334 0.573776
R16487 CSoutput.n338 CSoutput.n336 0.573776
R16488 CSoutput.n340 CSoutput.n338 0.573776
R16489 CSoutput.n342 CSoutput.n340 0.573776
R16490 CSoutput.n344 CSoutput.n342 0.573776
R16491 CSoutput.n346 CSoutput.n344 0.573776
R16492 CSoutput.n320 CSoutput.n318 0.573776
R16493 CSoutput.n322 CSoutput.n320 0.573776
R16494 CSoutput.n324 CSoutput.n322 0.573776
R16495 CSoutput.n326 CSoutput.n324 0.573776
R16496 CSoutput.n328 CSoutput.n326 0.573776
R16497 CSoutput.n330 CSoutput.n328 0.573776
R16498 CSoutput.n305 CSoutput.n303 0.573776
R16499 CSoutput.n307 CSoutput.n305 0.573776
R16500 CSoutput.n309 CSoutput.n307 0.573776
R16501 CSoutput.n311 CSoutput.n309 0.573776
R16502 CSoutput.n313 CSoutput.n311 0.573776
R16503 CSoutput.n315 CSoutput.n313 0.573776
R16504 CSoutput.n394 CSoutput.n392 0.573776
R16505 CSoutput.n392 CSoutput.n390 0.573776
R16506 CSoutput.n390 CSoutput.n388 0.573776
R16507 CSoutput.n388 CSoutput.n386 0.573776
R16508 CSoutput.n386 CSoutput.n384 0.573776
R16509 CSoutput.n384 CSoutput.n382 0.573776
R16510 CSoutput.n378 CSoutput.n376 0.573776
R16511 CSoutput.n376 CSoutput.n374 0.573776
R16512 CSoutput.n374 CSoutput.n372 0.573776
R16513 CSoutput.n372 CSoutput.n370 0.573776
R16514 CSoutput.n370 CSoutput.n368 0.573776
R16515 CSoutput.n368 CSoutput.n366 0.573776
R16516 CSoutput.n363 CSoutput.n361 0.573776
R16517 CSoutput.n361 CSoutput.n359 0.573776
R16518 CSoutput.n359 CSoutput.n357 0.573776
R16519 CSoutput.n357 CSoutput.n355 0.573776
R16520 CSoutput.n355 CSoutput.n353 0.573776
R16521 CSoutput.n353 CSoutput.n351 0.573776
R16522 CSoutput.n397 CSoutput.n264 0.53442
R16523 CSoutput.n292 CSoutput.n290 0.358259
R16524 CSoutput.n294 CSoutput.n292 0.358259
R16525 CSoutput.n296 CSoutput.n294 0.358259
R16526 CSoutput.n298 CSoutput.n296 0.358259
R16527 CSoutput.n280 CSoutput.n278 0.358259
R16528 CSoutput.n282 CSoutput.n280 0.358259
R16529 CSoutput.n284 CSoutput.n282 0.358259
R16530 CSoutput.n286 CSoutput.n284 0.358259
R16531 CSoutput.n269 CSoutput.n267 0.358259
R16532 CSoutput.n271 CSoutput.n269 0.358259
R16533 CSoutput.n273 CSoutput.n271 0.358259
R16534 CSoutput.n275 CSoutput.n273 0.358259
R16535 CSoutput.n112 CSoutput.n110 0.358259
R16536 CSoutput.n110 CSoutput.n108 0.358259
R16537 CSoutput.n108 CSoutput.n106 0.358259
R16538 CSoutput.n106 CSoutput.n104 0.358259
R16539 CSoutput.n100 CSoutput.n98 0.358259
R16540 CSoutput.n98 CSoutput.n96 0.358259
R16541 CSoutput.n96 CSoutput.n94 0.358259
R16542 CSoutput.n94 CSoutput.n92 0.358259
R16543 CSoutput.n89 CSoutput.n87 0.358259
R16544 CSoutput.n87 CSoutput.n85 0.358259
R16545 CSoutput.n85 CSoutput.n83 0.358259
R16546 CSoutput.n83 CSoutput.n81 0.358259
R16547 CSoutput.n21 CSoutput.n20 0.169105
R16548 CSoutput.n21 CSoutput.n16 0.169105
R16549 CSoutput.n26 CSoutput.n16 0.169105
R16550 CSoutput.n27 CSoutput.n26 0.169105
R16551 CSoutput.n27 CSoutput.n14 0.169105
R16552 CSoutput.n32 CSoutput.n14 0.169105
R16553 CSoutput.n33 CSoutput.n32 0.169105
R16554 CSoutput.n34 CSoutput.n33 0.169105
R16555 CSoutput.n34 CSoutput.n12 0.169105
R16556 CSoutput.n39 CSoutput.n12 0.169105
R16557 CSoutput.n40 CSoutput.n39 0.169105
R16558 CSoutput.n40 CSoutput.n10 0.169105
R16559 CSoutput.n45 CSoutput.n10 0.169105
R16560 CSoutput.n46 CSoutput.n45 0.169105
R16561 CSoutput.n47 CSoutput.n46 0.169105
R16562 CSoutput.n47 CSoutput.n8 0.169105
R16563 CSoutput.n52 CSoutput.n8 0.169105
R16564 CSoutput.n53 CSoutput.n52 0.169105
R16565 CSoutput.n53 CSoutput.n6 0.169105
R16566 CSoutput.n58 CSoutput.n6 0.169105
R16567 CSoutput.n59 CSoutput.n58 0.169105
R16568 CSoutput.n60 CSoutput.n59 0.169105
R16569 CSoutput.n60 CSoutput.n4 0.169105
R16570 CSoutput.n66 CSoutput.n4 0.169105
R16571 CSoutput.n67 CSoutput.n66 0.169105
R16572 CSoutput.n68 CSoutput.n67 0.169105
R16573 CSoutput.n68 CSoutput.n2 0.169105
R16574 CSoutput.n73 CSoutput.n2 0.169105
R16575 CSoutput.n74 CSoutput.n73 0.169105
R16576 CSoutput.n74 CSoutput.n0 0.169105
R16577 CSoutput.n78 CSoutput.n0 0.169105
R16578 CSoutput.n207 CSoutput.n206 0.0910737
R16579 CSoutput.n258 CSoutput.n255 0.0723685
R16580 CSoutput.n212 CSoutput.n207 0.0522944
R16581 CSoutput.n255 CSoutput.n254 0.0499135
R16582 CSoutput.n206 CSoutput.n205 0.0499135
R16583 CSoutput.n240 CSoutput.n239 0.0464294
R16584 CSoutput.n248 CSoutput.n245 0.0391444
R16585 CSoutput.n207 CSoutput.t178 0.023435
R16586 CSoutput.n255 CSoutput.t170 0.02262
R16587 CSoutput.n206 CSoutput.t172 0.02262
R16588 CSoutput CSoutput.n397 0.0052
R16589 CSoutput.n177 CSoutput.n160 0.00365111
R16590 CSoutput.n180 CSoutput.n161 0.00365111
R16591 CSoutput.n163 CSoutput.n162 0.00365111
R16592 CSoutput.n205 CSoutput.n164 0.00365111
R16593 CSoutput.n169 CSoutput.n165 0.00365111
R16594 CSoutput.n252 CSoutput.n166 0.00365111
R16595 CSoutput.n243 CSoutput.n242 0.00365111
R16596 CSoutput.n223 CSoutput.n196 0.00365111
R16597 CSoutput.n225 CSoutput.n195 0.00365111
R16598 CSoutput.n213 CSoutput.n212 0.00365111
R16599 CSoutput.n219 CSoutput.n199 0.00365111
R16600 CSoutput.n221 CSoutput.n198 0.00365111
R16601 CSoutput.n143 CSoutput.n126 0.00365111
R16602 CSoutput.n146 CSoutput.n127 0.00365111
R16603 CSoutput.n129 CSoutput.n128 0.00365111
R16604 CSoutput.n239 CSoutput.n130 0.00365111
R16605 CSoutput.n135 CSoutput.n131 0.00365111
R16606 CSoutput.n262 CSoutput.n132 0.00365111
R16607 CSoutput.n174 CSoutput.n164 0.00340054
R16608 CSoutput.n167 CSoutput.n165 0.00340054
R16609 CSoutput.n252 CSoutput.n251 0.00340054
R16610 CSoutput.n247 CSoutput.n160 0.00340054
R16611 CSoutput.n176 CSoutput.n161 0.00340054
R16612 CSoutput.n179 CSoutput.n163 0.00340054
R16613 CSoutput.n218 CSoutput.n213 0.00340054
R16614 CSoutput.n220 CSoutput.n219 0.00340054
R16615 CSoutput.n222 CSoutput.n221 0.00340054
R16616 CSoutput.n244 CSoutput.n243 0.00340054
R16617 CSoutput.n224 CSoutput.n223 0.00340054
R16618 CSoutput.n226 CSoutput.n225 0.00340054
R16619 CSoutput.n140 CSoutput.n130 0.00340054
R16620 CSoutput.n133 CSoutput.n131 0.00340054
R16621 CSoutput.n262 CSoutput.n261 0.00340054
R16622 CSoutput.n257 CSoutput.n126 0.00340054
R16623 CSoutput.n142 CSoutput.n127 0.00340054
R16624 CSoutput.n145 CSoutput.n129 0.00340054
R16625 CSoutput.n175 CSoutput.n169 0.00252698
R16626 CSoutput.n168 CSoutput.n166 0.00252698
R16627 CSoutput.n250 CSoutput.n249 0.00252698
R16628 CSoutput.n178 CSoutput.n176 0.00252698
R16629 CSoutput.n181 CSoutput.n179 0.00252698
R16630 CSoutput.n254 CSoutput.n149 0.00252698
R16631 CSoutput.n175 CSoutput.n174 0.00252698
R16632 CSoutput.n168 CSoutput.n167 0.00252698
R16633 CSoutput.n251 CSoutput.n250 0.00252698
R16634 CSoutput.n178 CSoutput.n177 0.00252698
R16635 CSoutput.n181 CSoutput.n180 0.00252698
R16636 CSoutput.n162 CSoutput.n149 0.00252698
R16637 CSoutput.n229 CSoutput.n199 0.00252698
R16638 CSoutput.n228 CSoutput.n198 0.00252698
R16639 CSoutput.n227 CSoutput.n183 0.00252698
R16640 CSoutput.n224 CSoutput.n194 0.00252698
R16641 CSoutput.n231 CSoutput.n226 0.00252698
R16642 CSoutput.n240 CSoutput.n233 0.00252698
R16643 CSoutput.n229 CSoutput.n218 0.00252698
R16644 CSoutput.n228 CSoutput.n220 0.00252698
R16645 CSoutput.n227 CSoutput.n222 0.00252698
R16646 CSoutput.n242 CSoutput.n194 0.00252698
R16647 CSoutput.n231 CSoutput.n196 0.00252698
R16648 CSoutput.n233 CSoutput.n195 0.00252698
R16649 CSoutput.n141 CSoutput.n135 0.00252698
R16650 CSoutput.n134 CSoutput.n132 0.00252698
R16651 CSoutput.n260 CSoutput.n259 0.00252698
R16652 CSoutput.n144 CSoutput.n142 0.00252698
R16653 CSoutput.n147 CSoutput.n145 0.00252698
R16654 CSoutput.n264 CSoutput.n115 0.00252698
R16655 CSoutput.n141 CSoutput.n140 0.00252698
R16656 CSoutput.n134 CSoutput.n133 0.00252698
R16657 CSoutput.n261 CSoutput.n260 0.00252698
R16658 CSoutput.n144 CSoutput.n143 0.00252698
R16659 CSoutput.n147 CSoutput.n146 0.00252698
R16660 CSoutput.n128 CSoutput.n115 0.00252698
R16661 CSoutput.n249 CSoutput.n248 0.0020275
R16662 CSoutput.n248 CSoutput.n247 0.0020275
R16663 CSoutput.n245 CSoutput.n183 0.0020275
R16664 CSoutput.n245 CSoutput.n244 0.0020275
R16665 CSoutput.n259 CSoutput.n258 0.0020275
R16666 CSoutput.n258 CSoutput.n257 0.0020275
R16667 CSoutput.n159 CSoutput.n158 0.00166668
R16668 CSoutput.n241 CSoutput.n197 0.00166668
R16669 CSoutput.n125 CSoutput.n124 0.00166668
R16670 CSoutput.n263 CSoutput.n125 0.00133328
R16671 CSoutput.n197 CSoutput.n193 0.00133328
R16672 CSoutput.n253 CSoutput.n159 0.00133328
R16673 CSoutput.n256 CSoutput.n148 0.001
R16674 CSoutput.n234 CSoutput.n148 0.001
R16675 CSoutput.n136 CSoutput.n116 0.001
R16676 CSoutput.n235 CSoutput.n116 0.001
R16677 CSoutput.n137 CSoutput.n117 0.001
R16678 CSoutput.n236 CSoutput.n117 0.001
R16679 CSoutput.n138 CSoutput.n118 0.001
R16680 CSoutput.n237 CSoutput.n118 0.001
R16681 CSoutput.n139 CSoutput.n119 0.001
R16682 CSoutput.n238 CSoutput.n119 0.001
R16683 CSoutput.n232 CSoutput.n184 0.001
R16684 CSoutput.n232 CSoutput.n230 0.001
R16685 CSoutput.n214 CSoutput.n185 0.001
R16686 CSoutput.n208 CSoutput.n185 0.001
R16687 CSoutput.n215 CSoutput.n186 0.001
R16688 CSoutput.n209 CSoutput.n186 0.001
R16689 CSoutput.n216 CSoutput.n187 0.001
R16690 CSoutput.n210 CSoutput.n187 0.001
R16691 CSoutput.n217 CSoutput.n188 0.001
R16692 CSoutput.n211 CSoutput.n188 0.001
R16693 CSoutput.n246 CSoutput.n182 0.001
R16694 CSoutput.n200 CSoutput.n182 0.001
R16695 CSoutput.n170 CSoutput.n150 0.001
R16696 CSoutput.n201 CSoutput.n150 0.001
R16697 CSoutput.n171 CSoutput.n151 0.001
R16698 CSoutput.n202 CSoutput.n151 0.001
R16699 CSoutput.n172 CSoutput.n152 0.001
R16700 CSoutput.n203 CSoutput.n152 0.001
R16701 CSoutput.n173 CSoutput.n153 0.001
R16702 CSoutput.n204 CSoutput.n153 0.001
R16703 CSoutput.n204 CSoutput.n154 0.001
R16704 CSoutput.n203 CSoutput.n155 0.001
R16705 CSoutput.n202 CSoutput.n156 0.001
R16706 CSoutput.n201 CSoutput.t189 0.001
R16707 CSoutput.n200 CSoutput.n157 0.001
R16708 CSoutput.n173 CSoutput.n155 0.001
R16709 CSoutput.n172 CSoutput.n156 0.001
R16710 CSoutput.n171 CSoutput.t189 0.001
R16711 CSoutput.n170 CSoutput.n157 0.001
R16712 CSoutput.n246 CSoutput.n158 0.001
R16713 CSoutput.n211 CSoutput.n189 0.001
R16714 CSoutput.n210 CSoutput.n190 0.001
R16715 CSoutput.n209 CSoutput.n191 0.001
R16716 CSoutput.n208 CSoutput.t168 0.001
R16717 CSoutput.n230 CSoutput.n192 0.001
R16718 CSoutput.n217 CSoutput.n190 0.001
R16719 CSoutput.n216 CSoutput.n191 0.001
R16720 CSoutput.n215 CSoutput.t168 0.001
R16721 CSoutput.n214 CSoutput.n192 0.001
R16722 CSoutput.n241 CSoutput.n184 0.001
R16723 CSoutput.n238 CSoutput.n120 0.001
R16724 CSoutput.n237 CSoutput.n121 0.001
R16725 CSoutput.n236 CSoutput.n122 0.001
R16726 CSoutput.n235 CSoutput.t175 0.001
R16727 CSoutput.n234 CSoutput.n123 0.001
R16728 CSoutput.n139 CSoutput.n121 0.001
R16729 CSoutput.n138 CSoutput.n122 0.001
R16730 CSoutput.n137 CSoutput.t175 0.001
R16731 CSoutput.n136 CSoutput.n123 0.001
R16732 CSoutput.n256 CSoutput.n124 0.001
R16733 a_n2982_13878.n8 a_n2982_13878.t102 538.698
R16734 a_n2982_13878.n104 a_n2982_13878.t79 512.366
R16735 a_n2982_13878.n103 a_n2982_13878.t84 512.366
R16736 a_n2982_13878.n95 a_n2982_13878.t72 512.366
R16737 a_n2982_13878.n102 a_n2982_13878.t89 512.366
R16738 a_n2982_13878.n101 a_n2982_13878.t98 512.366
R16739 a_n2982_13878.n96 a_n2982_13878.t99 512.366
R16740 a_n2982_13878.n100 a_n2982_13878.t66 512.366
R16741 a_n2982_13878.n99 a_n2982_13878.t81 512.366
R16742 a_n2982_13878.n97 a_n2982_13878.t69 512.366
R16743 a_n2982_13878.n98 a_n2982_13878.t76 512.366
R16744 a_n2982_13878.n66 a_n2982_13878.t49 532.5
R16745 a_n2982_13878.n119 a_n2982_13878.t15 512.366
R16746 a_n2982_13878.n118 a_n2982_13878.t33 512.366
R16747 a_n2982_13878.n92 a_n2982_13878.t45 512.366
R16748 a_n2982_13878.n117 a_n2982_13878.t37 512.366
R16749 a_n2982_13878.n116 a_n2982_13878.t51 512.366
R16750 a_n2982_13878.n93 a_n2982_13878.t29 512.366
R16751 a_n2982_13878.n115 a_n2982_13878.t23 512.366
R16752 a_n2982_13878.n114 a_n2982_13878.t53 512.366
R16753 a_n2982_13878.n94 a_n2982_13878.t25 512.366
R16754 a_n2982_13878.n113 a_n2982_13878.t35 512.366
R16755 a_n2982_13878.n26 a_n2982_13878.t39 538.698
R16756 a_n2982_13878.n145 a_n2982_13878.t55 512.366
R16757 a_n2982_13878.n87 a_n2982_13878.t47 512.366
R16758 a_n2982_13878.n146 a_n2982_13878.t43 512.366
R16759 a_n2982_13878.n86 a_n2982_13878.t13 512.366
R16760 a_n2982_13878.n147 a_n2982_13878.t59 512.366
R16761 a_n2982_13878.n148 a_n2982_13878.t27 512.366
R16762 a_n2982_13878.n85 a_n2982_13878.t19 512.366
R16763 a_n2982_13878.n149 a_n2982_13878.t41 512.366
R16764 a_n2982_13878.n84 a_n2982_13878.t57 512.366
R16765 a_n2982_13878.n150 a_n2982_13878.t17 512.366
R16766 a_n2982_13878.n32 a_n2982_13878.t101 538.698
R16767 a_n2982_13878.n139 a_n2982_13878.t70 512.366
R16768 a_n2982_13878.n91 a_n2982_13878.t71 512.366
R16769 a_n2982_13878.n140 a_n2982_13878.t96 512.366
R16770 a_n2982_13878.n90 a_n2982_13878.t97 512.366
R16771 a_n2982_13878.n141 a_n2982_13878.t68 512.366
R16772 a_n2982_13878.n142 a_n2982_13878.t92 512.366
R16773 a_n2982_13878.n89 a_n2982_13878.t93 512.366
R16774 a_n2982_13878.n143 a_n2982_13878.t65 512.366
R16775 a_n2982_13878.n88 a_n2982_13878.t78 512.366
R16776 a_n2982_13878.n144 a_n2982_13878.t88 512.366
R16777 a_n2982_13878.n131 a_n2982_13878.t86 512.366
R16778 a_n2982_13878.n130 a_n2982_13878.t75 512.366
R16779 a_n2982_13878.n129 a_n2982_13878.t64 512.366
R16780 a_n2982_13878.n133 a_n2982_13878.t94 512.366
R16781 a_n2982_13878.n132 a_n2982_13878.t83 512.366
R16782 a_n2982_13878.n128 a_n2982_13878.t82 512.366
R16783 a_n2982_13878.n135 a_n2982_13878.t90 512.366
R16784 a_n2982_13878.n134 a_n2982_13878.t73 512.366
R16785 a_n2982_13878.n127 a_n2982_13878.t74 512.366
R16786 a_n2982_13878.n137 a_n2982_13878.t77 512.366
R16787 a_n2982_13878.n136 a_n2982_13878.t87 512.366
R16788 a_n2982_13878.n126 a_n2982_13878.t103 512.366
R16789 a_n2982_13878.n82 a_n2982_13878.n3 70.5844
R16790 a_n2982_13878.n34 a_n2982_13878.n33 44.7878
R16791 a_n2982_13878.n22 a_n2982_13878.n56 70.5844
R16792 a_n2982_13878.n28 a_n2982_13878.n48 70.5844
R16793 a_n2982_13878.n47 a_n2982_13878.n28 70.1674
R16794 a_n2982_13878.n47 a_n2982_13878.n88 20.9683
R16795 a_n2982_13878.n27 a_n2982_13878.n46 74.73
R16796 a_n2982_13878.n143 a_n2982_13878.n46 11.843
R16797 a_n2982_13878.n45 a_n2982_13878.n27 80.4688
R16798 a_n2982_13878.n45 a_n2982_13878.n89 0.365327
R16799 a_n2982_13878.n29 a_n2982_13878.n44 75.0448
R16800 a_n2982_13878.n43 a_n2982_13878.n29 70.1674
R16801 a_n2982_13878.n43 a_n2982_13878.n90 20.9683
R16802 a_n2982_13878.n30 a_n2982_13878.n42 70.3058
R16803 a_n2982_13878.n140 a_n2982_13878.n42 20.6913
R16804 a_n2982_13878.n41 a_n2982_13878.n30 75.3623
R16805 a_n2982_13878.n41 a_n2982_13878.n91 10.5784
R16806 a_n2982_13878.n32 a_n2982_13878.n31 44.7878
R16807 a_n2982_13878.n55 a_n2982_13878.n22 70.1674
R16808 a_n2982_13878.n55 a_n2982_13878.n84 20.9683
R16809 a_n2982_13878.n21 a_n2982_13878.n54 74.73
R16810 a_n2982_13878.n149 a_n2982_13878.n54 11.843
R16811 a_n2982_13878.n53 a_n2982_13878.n21 80.4688
R16812 a_n2982_13878.n53 a_n2982_13878.n85 0.365327
R16813 a_n2982_13878.n23 a_n2982_13878.n52 75.0448
R16814 a_n2982_13878.n51 a_n2982_13878.n23 70.1674
R16815 a_n2982_13878.n51 a_n2982_13878.n86 20.9683
R16816 a_n2982_13878.n24 a_n2982_13878.n50 70.3058
R16817 a_n2982_13878.n146 a_n2982_13878.n50 20.6913
R16818 a_n2982_13878.n49 a_n2982_13878.n24 75.3623
R16819 a_n2982_13878.n49 a_n2982_13878.n87 10.5784
R16820 a_n2982_13878.n26 a_n2982_13878.n25 44.7878
R16821 a_n2982_13878.n13 a_n2982_13878.n65 70.1674
R16822 a_n2982_13878.n15 a_n2982_13878.n62 70.1674
R16823 a_n2982_13878.n17 a_n2982_13878.n60 70.1674
R16824 a_n2982_13878.n19 a_n2982_13878.n58 70.1674
R16825 a_n2982_13878.n58 a_n2982_13878.n126 20.9683
R16826 a_n2982_13878.n57 a_n2982_13878.n20 75.0448
R16827 a_n2982_13878.n136 a_n2982_13878.n57 11.2134
R16828 a_n2982_13878.n20 a_n2982_13878.n137 161.3
R16829 a_n2982_13878.n60 a_n2982_13878.n127 20.9683
R16830 a_n2982_13878.n59 a_n2982_13878.n18 75.0448
R16831 a_n2982_13878.n134 a_n2982_13878.n59 11.2134
R16832 a_n2982_13878.n18 a_n2982_13878.n135 161.3
R16833 a_n2982_13878.n62 a_n2982_13878.n128 20.9683
R16834 a_n2982_13878.n61 a_n2982_13878.n16 75.0448
R16835 a_n2982_13878.n132 a_n2982_13878.n61 11.2134
R16836 a_n2982_13878.n16 a_n2982_13878.n133 161.3
R16837 a_n2982_13878.n65 a_n2982_13878.n129 20.9683
R16838 a_n2982_13878.n63 a_n2982_13878.n14 75.0448
R16839 a_n2982_13878.n130 a_n2982_13878.n63 11.2134
R16840 a_n2982_13878.n14 a_n2982_13878.n131 161.3
R16841 a_n2982_13878.n34 a_n2982_13878.n113 14.1668
R16842 a_n2982_13878.n74 a_n2982_13878.n73 75.3623
R16843 a_n2982_13878.n72 a_n2982_13878.n9 70.3058
R16844 a_n2982_13878.n9 a_n2982_13878.n71 70.1674
R16845 a_n2982_13878.n71 a_n2982_13878.n93 20.9683
R16846 a_n2982_13878.n70 a_n2982_13878.n10 75.0448
R16847 a_n2982_13878.n116 a_n2982_13878.n70 11.2134
R16848 a_n2982_13878.n69 a_n2982_13878.n10 80.4688
R16849 a_n2982_13878.n12 a_n2982_13878.n68 74.73
R16850 a_n2982_13878.n67 a_n2982_13878.n12 70.1674
R16851 a_n2982_13878.n119 a_n2982_13878.n67 20.9683
R16852 a_n2982_13878.n11 a_n2982_13878.n66 70.5844
R16853 a_n2982_13878.n3 a_n2982_13878.n81 70.1674
R16854 a_n2982_13878.n81 a_n2982_13878.n97 20.9683
R16855 a_n2982_13878.n80 a_n2982_13878.n4 74.73
R16856 a_n2982_13878.n99 a_n2982_13878.n80 11.843
R16857 a_n2982_13878.n79 a_n2982_13878.n4 80.4688
R16858 a_n2982_13878.n79 a_n2982_13878.n100 0.365327
R16859 a_n2982_13878.n5 a_n2982_13878.n78 75.0448
R16860 a_n2982_13878.n77 a_n2982_13878.n5 70.1674
R16861 a_n2982_13878.n102 a_n2982_13878.n77 20.9683
R16862 a_n2982_13878.n7 a_n2982_13878.n76 70.3058
R16863 a_n2982_13878.n76 a_n2982_13878.n95 20.6913
R16864 a_n2982_13878.n75 a_n2982_13878.n7 75.3623
R16865 a_n2982_13878.n103 a_n2982_13878.n75 10.5784
R16866 a_n2982_13878.n6 a_n2982_13878.n8 44.7878
R16867 a_n2982_13878.n1 a_n2982_13878.n111 81.3764
R16868 a_n2982_13878.n2 a_n2982_13878.n107 81.3764
R16869 a_n2982_13878.n2 a_n2982_13878.n105 81.3764
R16870 a_n2982_13878.n1 a_n2982_13878.n112 80.9324
R16871 a_n2982_13878.n1 a_n2982_13878.n110 80.9324
R16872 a_n2982_13878.n0 a_n2982_13878.n109 80.9324
R16873 a_n2982_13878.n2 a_n2982_13878.n108 80.9324
R16874 a_n2982_13878.n2 a_n2982_13878.n106 80.9324
R16875 a_n2982_13878.n39 a_n2982_13878.t40 74.6477
R16876 a_n2982_13878.n37 a_n2982_13878.t22 74.6477
R16877 a_n2982_13878.n36 a_n2982_13878.t50 74.2899
R16878 a_n2982_13878.n40 a_n2982_13878.t32 74.2897
R16879 a_n2982_13878.n40 a_n2982_13878.n152 70.6783
R16880 a_n2982_13878.n38 a_n2982_13878.n153 70.6783
R16881 a_n2982_13878.n38 a_n2982_13878.n154 70.6783
R16882 a_n2982_13878.n39 a_n2982_13878.n83 70.6783
R16883 a_n2982_13878.n37 a_n2982_13878.n120 70.6783
R16884 a_n2982_13878.n37 a_n2982_13878.n121 70.6783
R16885 a_n2982_13878.n35 a_n2982_13878.n122 70.6783
R16886 a_n2982_13878.n35 a_n2982_13878.n123 70.6783
R16887 a_n2982_13878.n36 a_n2982_13878.n124 70.6783
R16888 a_n2982_13878.n155 a_n2982_13878.n39 70.6782
R16889 a_n2982_13878.n104 a_n2982_13878.n103 48.2005
R16890 a_n2982_13878.n77 a_n2982_13878.n101 20.9683
R16891 a_n2982_13878.n100 a_n2982_13878.n96 48.2005
R16892 a_n2982_13878.n98 a_n2982_13878.n81 20.9683
R16893 a_n2982_13878.n67 a_n2982_13878.n118 20.9683
R16894 a_n2982_13878.n117 a_n2982_13878.n116 48.2005
R16895 a_n2982_13878.n115 a_n2982_13878.n71 20.9683
R16896 a_n2982_13878.n113 a_n2982_13878.n94 48.2005
R16897 a_n2982_13878.n145 a_n2982_13878.n87 48.2005
R16898 a_n2982_13878.n147 a_n2982_13878.n51 20.9683
R16899 a_n2982_13878.n148 a_n2982_13878.n85 48.2005
R16900 a_n2982_13878.n150 a_n2982_13878.n55 20.9683
R16901 a_n2982_13878.n139 a_n2982_13878.n91 48.2005
R16902 a_n2982_13878.n141 a_n2982_13878.n43 20.9683
R16903 a_n2982_13878.n142 a_n2982_13878.n89 48.2005
R16904 a_n2982_13878.n144 a_n2982_13878.n47 20.9683
R16905 a_n2982_13878.n131 a_n2982_13878.n130 48.2005
R16906 a_n2982_13878.t91 a_n2982_13878.n65 533.335
R16907 a_n2982_13878.n133 a_n2982_13878.n132 48.2005
R16908 a_n2982_13878.t100 a_n2982_13878.n62 533.335
R16909 a_n2982_13878.n135 a_n2982_13878.n134 48.2005
R16910 a_n2982_13878.t85 a_n2982_13878.n60 533.335
R16911 a_n2982_13878.n137 a_n2982_13878.n136 48.2005
R16912 a_n2982_13878.t80 a_n2982_13878.n58 533.335
R16913 a_n2982_13878.n102 a_n2982_13878.n76 21.4216
R16914 a_n2982_13878.n69 a_n2982_13878.n92 47.835
R16915 a_n2982_13878.n72 a_n2982_13878.n114 20.6913
R16916 a_n2982_13878.n86 a_n2982_13878.n50 21.4216
R16917 a_n2982_13878.n90 a_n2982_13878.n42 21.4216
R16918 a_n2982_13878.n82 a_n2982_13878.t95 532.5
R16919 a_n2982_13878.t31 a_n2982_13878.n56 532.5
R16920 a_n2982_13878.t67 a_n2982_13878.n48 532.5
R16921 a_n2982_13878.n80 a_n2982_13878.n97 34.4824
R16922 a_n2982_13878.n68 a_n2982_13878.n92 11.843
R16923 a_n2982_13878.n114 a_n2982_13878.n73 36.139
R16924 a_n2982_13878.n84 a_n2982_13878.n54 34.4824
R16925 a_n2982_13878.n88 a_n2982_13878.n46 34.4824
R16926 a_n2982_13878.n101 a_n2982_13878.n78 35.3134
R16927 a_n2982_13878.n78 a_n2982_13878.n96 11.2134
R16928 a_n2982_13878.n70 a_n2982_13878.n93 35.3134
R16929 a_n2982_13878.n52 a_n2982_13878.n147 35.3134
R16930 a_n2982_13878.n148 a_n2982_13878.n52 11.2134
R16931 a_n2982_13878.n44 a_n2982_13878.n141 35.3134
R16932 a_n2982_13878.n142 a_n2982_13878.n44 11.2134
R16933 a_n2982_13878.n63 a_n2982_13878.n129 35.3134
R16934 a_n2982_13878.n61 a_n2982_13878.n128 35.3134
R16935 a_n2982_13878.n59 a_n2982_13878.n127 35.3134
R16936 a_n2982_13878.n57 a_n2982_13878.n126 35.3134
R16937 a_n2982_13878.n33 a_n2982_13878.n1 23.891
R16938 a_n2982_13878.n75 a_n2982_13878.n95 36.139
R16939 a_n2982_13878.n118 a_n2982_13878.n68 34.4824
R16940 a_n2982_13878.n73 a_n2982_13878.n94 10.5784
R16941 a_n2982_13878.n146 a_n2982_13878.n49 36.139
R16942 a_n2982_13878.n140 a_n2982_13878.n41 36.139
R16943 a_n2982_13878.n31 a_n2982_13878.n138 13.9285
R16944 a_n2982_13878.n3 a_n2982_13878.n64 13.724
R16945 a_n2982_13878.n125 a_n2982_13878.n11 12.4191
R16946 a_n2982_13878.n13 a_n2982_13878.n64 11.2486
R16947 a_n2982_13878.n138 a_n2982_13878.n20 11.2486
R16948 a_n2982_13878.n40 a_n2982_13878.n151 10.5745
R16949 a_n2982_13878.n151 a_n2982_13878.n22 8.58383
R16950 a_n2982_13878.n125 a_n2982_13878.n36 6.7311
R16951 a_n2982_13878.n151 a_n2982_13878.n64 5.3452
R16952 a_n2982_13878.n25 a_n2982_13878.n28 3.94368
R16953 a_n2982_13878.n33 a_n2982_13878.n6 3.7202
R16954 a_n2982_13878.n152 a_n2982_13878.t58 3.61217
R16955 a_n2982_13878.n152 a_n2982_13878.t18 3.61217
R16956 a_n2982_13878.n153 a_n2982_13878.t20 3.61217
R16957 a_n2982_13878.n153 a_n2982_13878.t42 3.61217
R16958 a_n2982_13878.n154 a_n2982_13878.t60 3.61217
R16959 a_n2982_13878.n154 a_n2982_13878.t28 3.61217
R16960 a_n2982_13878.n83 a_n2982_13878.t56 3.61217
R16961 a_n2982_13878.n83 a_n2982_13878.t48 3.61217
R16962 a_n2982_13878.n120 a_n2982_13878.t26 3.61217
R16963 a_n2982_13878.n120 a_n2982_13878.t36 3.61217
R16964 a_n2982_13878.n121 a_n2982_13878.t24 3.61217
R16965 a_n2982_13878.n121 a_n2982_13878.t54 3.61217
R16966 a_n2982_13878.n122 a_n2982_13878.t52 3.61217
R16967 a_n2982_13878.n122 a_n2982_13878.t30 3.61217
R16968 a_n2982_13878.n123 a_n2982_13878.t46 3.61217
R16969 a_n2982_13878.n123 a_n2982_13878.t38 3.61217
R16970 a_n2982_13878.n124 a_n2982_13878.t16 3.61217
R16971 a_n2982_13878.n124 a_n2982_13878.t34 3.61217
R16972 a_n2982_13878.n155 a_n2982_13878.t44 3.61217
R16973 a_n2982_13878.t14 a_n2982_13878.n155 3.61217
R16974 a_n2982_13878.n111 a_n2982_13878.t8 2.82907
R16975 a_n2982_13878.n111 a_n2982_13878.t11 2.82907
R16976 a_n2982_13878.n112 a_n2982_13878.t3 2.82907
R16977 a_n2982_13878.n112 a_n2982_13878.t12 2.82907
R16978 a_n2982_13878.n110 a_n2982_13878.t63 2.82907
R16979 a_n2982_13878.n110 a_n2982_13878.t9 2.82907
R16980 a_n2982_13878.n109 a_n2982_13878.t0 2.82907
R16981 a_n2982_13878.n109 a_n2982_13878.t62 2.82907
R16982 a_n2982_13878.n107 a_n2982_13878.t6 2.82907
R16983 a_n2982_13878.n107 a_n2982_13878.t5 2.82907
R16984 a_n2982_13878.n108 a_n2982_13878.t61 2.82907
R16985 a_n2982_13878.n108 a_n2982_13878.t2 2.82907
R16986 a_n2982_13878.n106 a_n2982_13878.t10 2.82907
R16987 a_n2982_13878.n106 a_n2982_13878.t1 2.82907
R16988 a_n2982_13878.n105 a_n2982_13878.t7 2.82907
R16989 a_n2982_13878.n105 a_n2982_13878.t4 2.82907
R16990 a_n2982_13878.n8 a_n2982_13878.n104 14.1668
R16991 a_n2982_13878.n98 a_n2982_13878.n82 22.3251
R16992 a_n2982_13878.n66 a_n2982_13878.n119 22.3251
R16993 a_n2982_13878.n34 a_n2982_13878.t21 538.698
R16994 a_n2982_13878.n145 a_n2982_13878.n26 14.1668
R16995 a_n2982_13878.n56 a_n2982_13878.n150 22.3251
R16996 a_n2982_13878.n139 a_n2982_13878.n32 14.1668
R16997 a_n2982_13878.n48 a_n2982_13878.n144 22.3251
R16998 a_n2982_13878.n138 a_n2982_13878.n125 1.30542
R16999 a_n2982_13878.n17 a_n2982_13878.n16 1.04595
R17000 a_n2982_13878.n79 a_n2982_13878.n99 47.835
R17001 a_n2982_13878.n69 a_n2982_13878.n117 0.365327
R17002 a_n2982_13878.n115 a_n2982_13878.n72 21.4216
R17003 a_n2982_13878.n149 a_n2982_13878.n53 47.835
R17004 a_n2982_13878.n143 a_n2982_13878.n45 47.835
R17005 a_n2982_13878.n0 a_n2982_13878.n2 31.7919
R17006 a_n2982_13878.n28 a_n2982_13878.n27 1.13686
R17007 a_n2982_13878.n22 a_n2982_13878.n21 1.13686
R17008 a_n2982_13878.n4 a_n2982_13878.n3 1.13686
R17009 a_n2982_13878.n39 a_n2982_13878.n38 1.07378
R17010 a_n2982_13878.n36 a_n2982_13878.n35 1.07378
R17011 a_n2982_13878.n1 a_n2982_13878.n0 0.888431
R17012 a_n2982_13878.n30 a_n2982_13878.n31 0.758076
R17013 a_n2982_13878.n29 a_n2982_13878.n30 0.758076
R17014 a_n2982_13878.n27 a_n2982_13878.n29 0.758076
R17015 a_n2982_13878.n24 a_n2982_13878.n25 0.758076
R17016 a_n2982_13878.n23 a_n2982_13878.n24 0.758076
R17017 a_n2982_13878.n21 a_n2982_13878.n23 0.758076
R17018 a_n2982_13878.n20 a_n2982_13878.n19 0.758076
R17019 a_n2982_13878.n18 a_n2982_13878.n17 0.758076
R17020 a_n2982_13878.n16 a_n2982_13878.n15 0.758076
R17021 a_n2982_13878.n14 a_n2982_13878.n13 0.758076
R17022 a_n2982_13878.n12 a_n2982_13878.n10 0.758076
R17023 a_n2982_13878.n10 a_n2982_13878.n9 0.758076
R17024 a_n2982_13878.n74 a_n2982_13878.n9 0.758076
R17025 a_n2982_13878.n7 a_n2982_13878.n6 0.758076
R17026 a_n2982_13878.n7 a_n2982_13878.n5 0.758076
R17027 a_n2982_13878.n5 a_n2982_13878.n4 0.758076
R17028 a_n2982_13878.n74 a_n2982_13878.n33 0.754288
R17029 a_n2982_13878.n38 a_n2982_13878.n40 0.716017
R17030 a_n2982_13878.n35 a_n2982_13878.n37 0.716017
R17031 a_n2982_13878.n19 a_n2982_13878.n18 0.67853
R17032 a_n2982_13878.n15 a_n2982_13878.n14 0.67853
R17033 a_n2982_13878.n12 a_n2982_13878.n11 0.568682
R17034 vdd.n303 vdd.n267 756.745
R17035 vdd.n252 vdd.n216 756.745
R17036 vdd.n209 vdd.n173 756.745
R17037 vdd.n158 vdd.n122 756.745
R17038 vdd.n116 vdd.n80 756.745
R17039 vdd.n65 vdd.n29 756.745
R17040 vdd.n1953 vdd.n1917 756.745
R17041 vdd.n2004 vdd.n1968 756.745
R17042 vdd.n1859 vdd.n1823 756.745
R17043 vdd.n1910 vdd.n1874 756.745
R17044 vdd.n1766 vdd.n1730 756.745
R17045 vdd.n1817 vdd.n1781 756.745
R17046 vdd.n1143 vdd.t4 640.208
R17047 vdd.n838 vdd.t49 640.208
R17048 vdd.n1147 vdd.t46 640.208
R17049 vdd.n829 vdd.t73 640.208
R17050 vdd.n724 vdd.t26 640.208
R17051 vdd.n2535 vdd.t67 640.208
R17052 vdd.n661 vdd.t15 640.208
R17053 vdd.n2532 vdd.t56 640.208
R17054 vdd.n625 vdd.t0 640.208
R17055 vdd.n899 vdd.t63 640.208
R17056 vdd.n1565 vdd.t36 592.009
R17057 vdd.n1602 vdd.t60 592.009
R17058 vdd.n1476 vdd.t70 592.009
R17059 vdd.n2074 vdd.t30 592.009
R17060 vdd.n1076 vdd.t8 592.009
R17061 vdd.n1036 vdd.t12 592.009
R17062 vdd.n3293 vdd.t33 592.009
R17063 vdd.n427 vdd.t22 592.009
R17064 vdd.n387 vdd.t40 592.009
R17065 vdd.n580 vdd.t43 592.009
R17066 vdd.n543 vdd.t53 592.009
R17067 vdd.n3080 vdd.t18 592.009
R17068 vdd.n304 vdd.n303 585
R17069 vdd.n302 vdd.n269 585
R17070 vdd.n301 vdd.n300 585
R17071 vdd.n272 vdd.n270 585
R17072 vdd.n295 vdd.n294 585
R17073 vdd.n293 vdd.n292 585
R17074 vdd.n276 vdd.n275 585
R17075 vdd.n287 vdd.n286 585
R17076 vdd.n285 vdd.n284 585
R17077 vdd.n280 vdd.n279 585
R17078 vdd.n253 vdd.n252 585
R17079 vdd.n251 vdd.n218 585
R17080 vdd.n250 vdd.n249 585
R17081 vdd.n221 vdd.n219 585
R17082 vdd.n244 vdd.n243 585
R17083 vdd.n242 vdd.n241 585
R17084 vdd.n225 vdd.n224 585
R17085 vdd.n236 vdd.n235 585
R17086 vdd.n234 vdd.n233 585
R17087 vdd.n229 vdd.n228 585
R17088 vdd.n210 vdd.n209 585
R17089 vdd.n208 vdd.n175 585
R17090 vdd.n207 vdd.n206 585
R17091 vdd.n178 vdd.n176 585
R17092 vdd.n201 vdd.n200 585
R17093 vdd.n199 vdd.n198 585
R17094 vdd.n182 vdd.n181 585
R17095 vdd.n193 vdd.n192 585
R17096 vdd.n191 vdd.n190 585
R17097 vdd.n186 vdd.n185 585
R17098 vdd.n159 vdd.n158 585
R17099 vdd.n157 vdd.n124 585
R17100 vdd.n156 vdd.n155 585
R17101 vdd.n127 vdd.n125 585
R17102 vdd.n150 vdd.n149 585
R17103 vdd.n148 vdd.n147 585
R17104 vdd.n131 vdd.n130 585
R17105 vdd.n142 vdd.n141 585
R17106 vdd.n140 vdd.n139 585
R17107 vdd.n135 vdd.n134 585
R17108 vdd.n117 vdd.n116 585
R17109 vdd.n115 vdd.n82 585
R17110 vdd.n114 vdd.n113 585
R17111 vdd.n85 vdd.n83 585
R17112 vdd.n108 vdd.n107 585
R17113 vdd.n106 vdd.n105 585
R17114 vdd.n89 vdd.n88 585
R17115 vdd.n100 vdd.n99 585
R17116 vdd.n98 vdd.n97 585
R17117 vdd.n93 vdd.n92 585
R17118 vdd.n66 vdd.n65 585
R17119 vdd.n64 vdd.n31 585
R17120 vdd.n63 vdd.n62 585
R17121 vdd.n34 vdd.n32 585
R17122 vdd.n57 vdd.n56 585
R17123 vdd.n55 vdd.n54 585
R17124 vdd.n38 vdd.n37 585
R17125 vdd.n49 vdd.n48 585
R17126 vdd.n47 vdd.n46 585
R17127 vdd.n42 vdd.n41 585
R17128 vdd.n1954 vdd.n1953 585
R17129 vdd.n1952 vdd.n1919 585
R17130 vdd.n1951 vdd.n1950 585
R17131 vdd.n1922 vdd.n1920 585
R17132 vdd.n1945 vdd.n1944 585
R17133 vdd.n1943 vdd.n1942 585
R17134 vdd.n1926 vdd.n1925 585
R17135 vdd.n1937 vdd.n1936 585
R17136 vdd.n1935 vdd.n1934 585
R17137 vdd.n1930 vdd.n1929 585
R17138 vdd.n2005 vdd.n2004 585
R17139 vdd.n2003 vdd.n1970 585
R17140 vdd.n2002 vdd.n2001 585
R17141 vdd.n1973 vdd.n1971 585
R17142 vdd.n1996 vdd.n1995 585
R17143 vdd.n1994 vdd.n1993 585
R17144 vdd.n1977 vdd.n1976 585
R17145 vdd.n1988 vdd.n1987 585
R17146 vdd.n1986 vdd.n1985 585
R17147 vdd.n1981 vdd.n1980 585
R17148 vdd.n1860 vdd.n1859 585
R17149 vdd.n1858 vdd.n1825 585
R17150 vdd.n1857 vdd.n1856 585
R17151 vdd.n1828 vdd.n1826 585
R17152 vdd.n1851 vdd.n1850 585
R17153 vdd.n1849 vdd.n1848 585
R17154 vdd.n1832 vdd.n1831 585
R17155 vdd.n1843 vdd.n1842 585
R17156 vdd.n1841 vdd.n1840 585
R17157 vdd.n1836 vdd.n1835 585
R17158 vdd.n1911 vdd.n1910 585
R17159 vdd.n1909 vdd.n1876 585
R17160 vdd.n1908 vdd.n1907 585
R17161 vdd.n1879 vdd.n1877 585
R17162 vdd.n1902 vdd.n1901 585
R17163 vdd.n1900 vdd.n1899 585
R17164 vdd.n1883 vdd.n1882 585
R17165 vdd.n1894 vdd.n1893 585
R17166 vdd.n1892 vdd.n1891 585
R17167 vdd.n1887 vdd.n1886 585
R17168 vdd.n1767 vdd.n1766 585
R17169 vdd.n1765 vdd.n1732 585
R17170 vdd.n1764 vdd.n1763 585
R17171 vdd.n1735 vdd.n1733 585
R17172 vdd.n1758 vdd.n1757 585
R17173 vdd.n1756 vdd.n1755 585
R17174 vdd.n1739 vdd.n1738 585
R17175 vdd.n1750 vdd.n1749 585
R17176 vdd.n1748 vdd.n1747 585
R17177 vdd.n1743 vdd.n1742 585
R17178 vdd.n1818 vdd.n1817 585
R17179 vdd.n1816 vdd.n1783 585
R17180 vdd.n1815 vdd.n1814 585
R17181 vdd.n1786 vdd.n1784 585
R17182 vdd.n1809 vdd.n1808 585
R17183 vdd.n1807 vdd.n1806 585
R17184 vdd.n1790 vdd.n1789 585
R17185 vdd.n1801 vdd.n1800 585
R17186 vdd.n1799 vdd.n1798 585
R17187 vdd.n1794 vdd.n1793 585
R17188 vdd.n3409 vdd.n352 488.781
R17189 vdd.n3291 vdd.n350 488.781
R17190 vdd.n3213 vdd.n515 488.781
R17191 vdd.n3211 vdd.n517 488.781
R17192 vdd.n2069 vdd.n1358 488.781
R17193 vdd.n2072 vdd.n2071 488.781
R17194 vdd.n1671 vdd.n1436 488.781
R17195 vdd.n1669 vdd.n1439 488.781
R17196 vdd.n281 vdd.t161 329.043
R17197 vdd.n230 vdd.t240 329.043
R17198 vdd.n187 vdd.t242 329.043
R17199 vdd.n136 vdd.t234 329.043
R17200 vdd.n94 vdd.t184 329.043
R17201 vdd.n43 vdd.t201 329.043
R17202 vdd.n1931 vdd.t191 329.043
R17203 vdd.n1982 vdd.t195 329.043
R17204 vdd.n1837 vdd.t178 329.043
R17205 vdd.n1888 vdd.t185 329.043
R17206 vdd.n1744 vdd.t202 329.043
R17207 vdd.n1795 vdd.t183 329.043
R17208 vdd.n1565 vdd.t39 319.788
R17209 vdd.n1602 vdd.t62 319.788
R17210 vdd.n1476 vdd.t72 319.788
R17211 vdd.n2074 vdd.t31 319.788
R17212 vdd.n1076 vdd.t10 319.788
R17213 vdd.n1036 vdd.t13 319.788
R17214 vdd.n3293 vdd.t34 319.788
R17215 vdd.n427 vdd.t24 319.788
R17216 vdd.n387 vdd.t41 319.788
R17217 vdd.n580 vdd.t45 319.788
R17218 vdd.n543 vdd.t55 319.788
R17219 vdd.n3080 vdd.t21 319.788
R17220 vdd.n1566 vdd.t38 303.69
R17221 vdd.n1603 vdd.t61 303.69
R17222 vdd.n1477 vdd.t71 303.69
R17223 vdd.n2075 vdd.t32 303.69
R17224 vdd.n1077 vdd.t11 303.69
R17225 vdd.n1037 vdd.t14 303.69
R17226 vdd.n3294 vdd.t35 303.69
R17227 vdd.n428 vdd.t25 303.69
R17228 vdd.n388 vdd.t42 303.69
R17229 vdd.n581 vdd.t44 303.69
R17230 vdd.n544 vdd.t54 303.69
R17231 vdd.n3081 vdd.t20 303.69
R17232 vdd.n2802 vdd.n788 279.512
R17233 vdd.n3042 vdd.n635 279.512
R17234 vdd.n2979 vdd.n632 279.512
R17235 vdd.n2734 vdd.n2733 279.512
R17236 vdd.n2495 vdd.n826 279.512
R17237 vdd.n2426 vdd.n2425 279.512
R17238 vdd.n1183 vdd.n1182 279.512
R17239 vdd.n2220 vdd.n966 279.512
R17240 vdd.n2958 vdd.n633 279.512
R17241 vdd.n3045 vdd.n3044 279.512
R17242 vdd.n2607 vdd.n2530 279.512
R17243 vdd.n2538 vdd.n784 279.512
R17244 vdd.n2423 vdd.n836 279.512
R17245 vdd.n834 vdd.n808 279.512
R17246 vdd.n1308 vdd.n1003 279.512
R17247 vdd.n1108 vdd.n961 279.512
R17248 vdd.n2218 vdd.n969 254.619
R17249 vdd.n613 vdd.n516 254.619
R17250 vdd.n2960 vdd.n633 185
R17251 vdd.n3043 vdd.n633 185
R17252 vdd.n2962 vdd.n2961 185
R17253 vdd.n2961 vdd.n631 185
R17254 vdd.n2963 vdd.n667 185
R17255 vdd.n2973 vdd.n667 185
R17256 vdd.n2964 vdd.n676 185
R17257 vdd.n676 vdd.n674 185
R17258 vdd.n2966 vdd.n2965 185
R17259 vdd.n2967 vdd.n2966 185
R17260 vdd.n2919 vdd.n675 185
R17261 vdd.n675 vdd.n671 185
R17262 vdd.n2918 vdd.n2917 185
R17263 vdd.n2917 vdd.n2916 185
R17264 vdd.n678 vdd.n677 185
R17265 vdd.n679 vdd.n678 185
R17266 vdd.n2909 vdd.n2908 185
R17267 vdd.n2910 vdd.n2909 185
R17268 vdd.n2907 vdd.n687 185
R17269 vdd.n692 vdd.n687 185
R17270 vdd.n2906 vdd.n2905 185
R17271 vdd.n2905 vdd.n2904 185
R17272 vdd.n689 vdd.n688 185
R17273 vdd.n698 vdd.n689 185
R17274 vdd.n2897 vdd.n2896 185
R17275 vdd.n2898 vdd.n2897 185
R17276 vdd.n2895 vdd.n699 185
R17277 vdd.n705 vdd.n699 185
R17278 vdd.n2894 vdd.n2893 185
R17279 vdd.n2893 vdd.n2892 185
R17280 vdd.n701 vdd.n700 185
R17281 vdd.n702 vdd.n701 185
R17282 vdd.n2885 vdd.n2884 185
R17283 vdd.n2886 vdd.n2885 185
R17284 vdd.n2883 vdd.n712 185
R17285 vdd.n712 vdd.n709 185
R17286 vdd.n2882 vdd.n2881 185
R17287 vdd.n2881 vdd.n2880 185
R17288 vdd.n714 vdd.n713 185
R17289 vdd.n715 vdd.n714 185
R17290 vdd.n2873 vdd.n2872 185
R17291 vdd.n2874 vdd.n2873 185
R17292 vdd.n2871 vdd.n723 185
R17293 vdd.n729 vdd.n723 185
R17294 vdd.n2870 vdd.n2869 185
R17295 vdd.n2869 vdd.n2868 185
R17296 vdd.n2859 vdd.n726 185
R17297 vdd.n736 vdd.n726 185
R17298 vdd.n2861 vdd.n2860 185
R17299 vdd.n2862 vdd.n2861 185
R17300 vdd.n2858 vdd.n737 185
R17301 vdd.n737 vdd.n733 185
R17302 vdd.n2857 vdd.n2856 185
R17303 vdd.n2856 vdd.n2855 185
R17304 vdd.n739 vdd.n738 185
R17305 vdd.n740 vdd.n739 185
R17306 vdd.n2848 vdd.n2847 185
R17307 vdd.n2849 vdd.n2848 185
R17308 vdd.n2846 vdd.n748 185
R17309 vdd.n753 vdd.n748 185
R17310 vdd.n2845 vdd.n2844 185
R17311 vdd.n2844 vdd.n2843 185
R17312 vdd.n750 vdd.n749 185
R17313 vdd.n759 vdd.n750 185
R17314 vdd.n2836 vdd.n2835 185
R17315 vdd.n2837 vdd.n2836 185
R17316 vdd.n2834 vdd.n760 185
R17317 vdd.n2710 vdd.n760 185
R17318 vdd.n2833 vdd.n2832 185
R17319 vdd.n2832 vdd.n2831 185
R17320 vdd.n762 vdd.n761 185
R17321 vdd.n2716 vdd.n762 185
R17322 vdd.n2824 vdd.n2823 185
R17323 vdd.n2825 vdd.n2824 185
R17324 vdd.n2822 vdd.n771 185
R17325 vdd.n771 vdd.n768 185
R17326 vdd.n2821 vdd.n2820 185
R17327 vdd.n2820 vdd.n2819 185
R17328 vdd.n773 vdd.n772 185
R17329 vdd.n774 vdd.n773 185
R17330 vdd.n2812 vdd.n2811 185
R17331 vdd.n2813 vdd.n2812 185
R17332 vdd.n2810 vdd.n782 185
R17333 vdd.n2728 vdd.n782 185
R17334 vdd.n2809 vdd.n2808 185
R17335 vdd.n2808 vdd.n2807 185
R17336 vdd.n784 vdd.n783 185
R17337 vdd.n785 vdd.n784 185
R17338 vdd.n2539 vdd.n2538 185
R17339 vdd.n2541 vdd.n2540 185
R17340 vdd.n2543 vdd.n2542 185
R17341 vdd.n2545 vdd.n2544 185
R17342 vdd.n2547 vdd.n2546 185
R17343 vdd.n2549 vdd.n2548 185
R17344 vdd.n2551 vdd.n2550 185
R17345 vdd.n2553 vdd.n2552 185
R17346 vdd.n2555 vdd.n2554 185
R17347 vdd.n2557 vdd.n2556 185
R17348 vdd.n2559 vdd.n2558 185
R17349 vdd.n2561 vdd.n2560 185
R17350 vdd.n2563 vdd.n2562 185
R17351 vdd.n2565 vdd.n2564 185
R17352 vdd.n2567 vdd.n2566 185
R17353 vdd.n2569 vdd.n2568 185
R17354 vdd.n2571 vdd.n2570 185
R17355 vdd.n2573 vdd.n2572 185
R17356 vdd.n2575 vdd.n2574 185
R17357 vdd.n2577 vdd.n2576 185
R17358 vdd.n2579 vdd.n2578 185
R17359 vdd.n2581 vdd.n2580 185
R17360 vdd.n2583 vdd.n2582 185
R17361 vdd.n2585 vdd.n2584 185
R17362 vdd.n2587 vdd.n2586 185
R17363 vdd.n2589 vdd.n2588 185
R17364 vdd.n2591 vdd.n2590 185
R17365 vdd.n2593 vdd.n2592 185
R17366 vdd.n2595 vdd.n2594 185
R17367 vdd.n2597 vdd.n2596 185
R17368 vdd.n2599 vdd.n2598 185
R17369 vdd.n2601 vdd.n2600 185
R17370 vdd.n2603 vdd.n2602 185
R17371 vdd.n2605 vdd.n2604 185
R17372 vdd.n2606 vdd.n2530 185
R17373 vdd.n2800 vdd.n2530 185
R17374 vdd.n3046 vdd.n3045 185
R17375 vdd.n3047 vdd.n624 185
R17376 vdd.n3049 vdd.n3048 185
R17377 vdd.n3051 vdd.n622 185
R17378 vdd.n3053 vdd.n3052 185
R17379 vdd.n3054 vdd.n621 185
R17380 vdd.n3056 vdd.n3055 185
R17381 vdd.n3058 vdd.n619 185
R17382 vdd.n3060 vdd.n3059 185
R17383 vdd.n3061 vdd.n618 185
R17384 vdd.n3063 vdd.n3062 185
R17385 vdd.n3065 vdd.n616 185
R17386 vdd.n3067 vdd.n3066 185
R17387 vdd.n3068 vdd.n615 185
R17388 vdd.n3070 vdd.n3069 185
R17389 vdd.n3072 vdd.n614 185
R17390 vdd.n3073 vdd.n611 185
R17391 vdd.n3076 vdd.n3075 185
R17392 vdd.n612 vdd.n610 185
R17393 vdd.n2932 vdd.n2931 185
R17394 vdd.n2934 vdd.n2933 185
R17395 vdd.n2936 vdd.n2928 185
R17396 vdd.n2938 vdd.n2937 185
R17397 vdd.n2939 vdd.n2927 185
R17398 vdd.n2941 vdd.n2940 185
R17399 vdd.n2943 vdd.n2925 185
R17400 vdd.n2945 vdd.n2944 185
R17401 vdd.n2946 vdd.n2924 185
R17402 vdd.n2948 vdd.n2947 185
R17403 vdd.n2950 vdd.n2922 185
R17404 vdd.n2952 vdd.n2951 185
R17405 vdd.n2953 vdd.n2921 185
R17406 vdd.n2955 vdd.n2954 185
R17407 vdd.n2957 vdd.n2920 185
R17408 vdd.n2959 vdd.n2958 185
R17409 vdd.n2958 vdd.n613 185
R17410 vdd.n3044 vdd.n628 185
R17411 vdd.n3044 vdd.n3043 185
R17412 vdd.n2661 vdd.n630 185
R17413 vdd.n631 vdd.n630 185
R17414 vdd.n2662 vdd.n666 185
R17415 vdd.n2973 vdd.n666 185
R17416 vdd.n2664 vdd.n2663 185
R17417 vdd.n2663 vdd.n674 185
R17418 vdd.n2665 vdd.n673 185
R17419 vdd.n2967 vdd.n673 185
R17420 vdd.n2667 vdd.n2666 185
R17421 vdd.n2666 vdd.n671 185
R17422 vdd.n2668 vdd.n681 185
R17423 vdd.n2916 vdd.n681 185
R17424 vdd.n2670 vdd.n2669 185
R17425 vdd.n2669 vdd.n679 185
R17426 vdd.n2671 vdd.n686 185
R17427 vdd.n2910 vdd.n686 185
R17428 vdd.n2673 vdd.n2672 185
R17429 vdd.n2672 vdd.n692 185
R17430 vdd.n2674 vdd.n691 185
R17431 vdd.n2904 vdd.n691 185
R17432 vdd.n2676 vdd.n2675 185
R17433 vdd.n2675 vdd.n698 185
R17434 vdd.n2677 vdd.n697 185
R17435 vdd.n2898 vdd.n697 185
R17436 vdd.n2679 vdd.n2678 185
R17437 vdd.n2678 vdd.n705 185
R17438 vdd.n2680 vdd.n704 185
R17439 vdd.n2892 vdd.n704 185
R17440 vdd.n2682 vdd.n2681 185
R17441 vdd.n2681 vdd.n702 185
R17442 vdd.n2683 vdd.n711 185
R17443 vdd.n2886 vdd.n711 185
R17444 vdd.n2685 vdd.n2684 185
R17445 vdd.n2684 vdd.n709 185
R17446 vdd.n2686 vdd.n717 185
R17447 vdd.n2880 vdd.n717 185
R17448 vdd.n2688 vdd.n2687 185
R17449 vdd.n2687 vdd.n715 185
R17450 vdd.n2689 vdd.n722 185
R17451 vdd.n2874 vdd.n722 185
R17452 vdd.n2691 vdd.n2690 185
R17453 vdd.n2690 vdd.n729 185
R17454 vdd.n2692 vdd.n728 185
R17455 vdd.n2868 vdd.n728 185
R17456 vdd.n2694 vdd.n2693 185
R17457 vdd.n2693 vdd.n736 185
R17458 vdd.n2695 vdd.n735 185
R17459 vdd.n2862 vdd.n735 185
R17460 vdd.n2697 vdd.n2696 185
R17461 vdd.n2696 vdd.n733 185
R17462 vdd.n2698 vdd.n742 185
R17463 vdd.n2855 vdd.n742 185
R17464 vdd.n2700 vdd.n2699 185
R17465 vdd.n2699 vdd.n740 185
R17466 vdd.n2701 vdd.n747 185
R17467 vdd.n2849 vdd.n747 185
R17468 vdd.n2703 vdd.n2702 185
R17469 vdd.n2702 vdd.n753 185
R17470 vdd.n2704 vdd.n752 185
R17471 vdd.n2843 vdd.n752 185
R17472 vdd.n2706 vdd.n2705 185
R17473 vdd.n2705 vdd.n759 185
R17474 vdd.n2707 vdd.n758 185
R17475 vdd.n2837 vdd.n758 185
R17476 vdd.n2709 vdd.n2708 185
R17477 vdd.n2710 vdd.n2709 185
R17478 vdd.n2610 vdd.n764 185
R17479 vdd.n2831 vdd.n764 185
R17480 vdd.n2718 vdd.n2717 185
R17481 vdd.n2717 vdd.n2716 185
R17482 vdd.n2719 vdd.n770 185
R17483 vdd.n2825 vdd.n770 185
R17484 vdd.n2721 vdd.n2720 185
R17485 vdd.n2720 vdd.n768 185
R17486 vdd.n2722 vdd.n776 185
R17487 vdd.n2819 vdd.n776 185
R17488 vdd.n2724 vdd.n2723 185
R17489 vdd.n2723 vdd.n774 185
R17490 vdd.n2725 vdd.n781 185
R17491 vdd.n2813 vdd.n781 185
R17492 vdd.n2727 vdd.n2726 185
R17493 vdd.n2728 vdd.n2727 185
R17494 vdd.n2609 vdd.n787 185
R17495 vdd.n2807 vdd.n787 185
R17496 vdd.n2608 vdd.n2607 185
R17497 vdd.n2607 vdd.n785 185
R17498 vdd.n2069 vdd.n2068 185
R17499 vdd.n2070 vdd.n2069 185
R17500 vdd.n1359 vdd.n1357 185
R17501 vdd.n2061 vdd.n1357 185
R17502 vdd.n2064 vdd.n2063 185
R17503 vdd.n2063 vdd.n2062 185
R17504 vdd.n1362 vdd.n1361 185
R17505 vdd.n1363 vdd.n1362 185
R17506 vdd.n2050 vdd.n2049 185
R17507 vdd.n2051 vdd.n2050 185
R17508 vdd.n1371 vdd.n1370 185
R17509 vdd.n2042 vdd.n1370 185
R17510 vdd.n2045 vdd.n2044 185
R17511 vdd.n2044 vdd.n2043 185
R17512 vdd.n1374 vdd.n1373 185
R17513 vdd.n1380 vdd.n1374 185
R17514 vdd.n2033 vdd.n2032 185
R17515 vdd.n2034 vdd.n2033 185
R17516 vdd.n1382 vdd.n1381 185
R17517 vdd.n2025 vdd.n1381 185
R17518 vdd.n2028 vdd.n2027 185
R17519 vdd.n2027 vdd.n2026 185
R17520 vdd.n1385 vdd.n1384 185
R17521 vdd.n1386 vdd.n1385 185
R17522 vdd.n2016 vdd.n2015 185
R17523 vdd.n2017 vdd.n2016 185
R17524 vdd.n1394 vdd.n1393 185
R17525 vdd.n1393 vdd.n1392 185
R17526 vdd.n1729 vdd.n1728 185
R17527 vdd.n1728 vdd.n1727 185
R17528 vdd.n1397 vdd.n1396 185
R17529 vdd.n1403 vdd.n1397 185
R17530 vdd.n1718 vdd.n1717 185
R17531 vdd.n1719 vdd.n1718 185
R17532 vdd.n1405 vdd.n1404 185
R17533 vdd.n1710 vdd.n1404 185
R17534 vdd.n1713 vdd.n1712 185
R17535 vdd.n1712 vdd.n1711 185
R17536 vdd.n1408 vdd.n1407 185
R17537 vdd.n1415 vdd.n1408 185
R17538 vdd.n1701 vdd.n1700 185
R17539 vdd.n1702 vdd.n1701 185
R17540 vdd.n1417 vdd.n1416 185
R17541 vdd.n1416 vdd.n1414 185
R17542 vdd.n1696 vdd.n1695 185
R17543 vdd.n1695 vdd.n1694 185
R17544 vdd.n1420 vdd.n1419 185
R17545 vdd.n1421 vdd.n1420 185
R17546 vdd.n1685 vdd.n1684 185
R17547 vdd.n1686 vdd.n1685 185
R17548 vdd.n1429 vdd.n1428 185
R17549 vdd.n1428 vdd.n1427 185
R17550 vdd.n1680 vdd.n1679 185
R17551 vdd.n1679 vdd.n1678 185
R17552 vdd.n1432 vdd.n1431 185
R17553 vdd.n1438 vdd.n1432 185
R17554 vdd.n1669 vdd.n1668 185
R17555 vdd.n1670 vdd.n1669 185
R17556 vdd.n1665 vdd.n1439 185
R17557 vdd.n1664 vdd.n1442 185
R17558 vdd.n1663 vdd.n1443 185
R17559 vdd.n1443 vdd.n1437 185
R17560 vdd.n1446 vdd.n1444 185
R17561 vdd.n1659 vdd.n1448 185
R17562 vdd.n1658 vdd.n1449 185
R17563 vdd.n1657 vdd.n1451 185
R17564 vdd.n1454 vdd.n1452 185
R17565 vdd.n1653 vdd.n1456 185
R17566 vdd.n1652 vdd.n1457 185
R17567 vdd.n1651 vdd.n1459 185
R17568 vdd.n1462 vdd.n1460 185
R17569 vdd.n1647 vdd.n1464 185
R17570 vdd.n1646 vdd.n1465 185
R17571 vdd.n1645 vdd.n1467 185
R17572 vdd.n1470 vdd.n1468 185
R17573 vdd.n1641 vdd.n1472 185
R17574 vdd.n1640 vdd.n1473 185
R17575 vdd.n1639 vdd.n1475 185
R17576 vdd.n1480 vdd.n1478 185
R17577 vdd.n1635 vdd.n1482 185
R17578 vdd.n1634 vdd.n1483 185
R17579 vdd.n1633 vdd.n1485 185
R17580 vdd.n1488 vdd.n1486 185
R17581 vdd.n1629 vdd.n1490 185
R17582 vdd.n1628 vdd.n1491 185
R17583 vdd.n1627 vdd.n1493 185
R17584 vdd.n1496 vdd.n1494 185
R17585 vdd.n1623 vdd.n1498 185
R17586 vdd.n1622 vdd.n1499 185
R17587 vdd.n1621 vdd.n1501 185
R17588 vdd.n1504 vdd.n1502 185
R17589 vdd.n1617 vdd.n1506 185
R17590 vdd.n1616 vdd.n1507 185
R17591 vdd.n1615 vdd.n1509 185
R17592 vdd.n1512 vdd.n1510 185
R17593 vdd.n1611 vdd.n1514 185
R17594 vdd.n1610 vdd.n1515 185
R17595 vdd.n1609 vdd.n1517 185
R17596 vdd.n1520 vdd.n1518 185
R17597 vdd.n1605 vdd.n1522 185
R17598 vdd.n1604 vdd.n1601 185
R17599 vdd.n1599 vdd.n1523 185
R17600 vdd.n1598 vdd.n1597 185
R17601 vdd.n1528 vdd.n1525 185
R17602 vdd.n1593 vdd.n1529 185
R17603 vdd.n1592 vdd.n1531 185
R17604 vdd.n1591 vdd.n1532 185
R17605 vdd.n1536 vdd.n1533 185
R17606 vdd.n1587 vdd.n1537 185
R17607 vdd.n1586 vdd.n1539 185
R17608 vdd.n1585 vdd.n1540 185
R17609 vdd.n1544 vdd.n1541 185
R17610 vdd.n1581 vdd.n1545 185
R17611 vdd.n1580 vdd.n1547 185
R17612 vdd.n1579 vdd.n1548 185
R17613 vdd.n1552 vdd.n1549 185
R17614 vdd.n1575 vdd.n1553 185
R17615 vdd.n1574 vdd.n1555 185
R17616 vdd.n1573 vdd.n1556 185
R17617 vdd.n1560 vdd.n1557 185
R17618 vdd.n1569 vdd.n1561 185
R17619 vdd.n1568 vdd.n1563 185
R17620 vdd.n1564 vdd.n1436 185
R17621 vdd.n1437 vdd.n1436 185
R17622 vdd.n2073 vdd.n2072 185
R17623 vdd.n2077 vdd.n1353 185
R17624 vdd.n1352 vdd.n1346 185
R17625 vdd.n1350 vdd.n1349 185
R17626 vdd.n1348 vdd.n1107 185
R17627 vdd.n2081 vdd.n1104 185
R17628 vdd.n2083 vdd.n2082 185
R17629 vdd.n2085 vdd.n1102 185
R17630 vdd.n2087 vdd.n2086 185
R17631 vdd.n2088 vdd.n1097 185
R17632 vdd.n2090 vdd.n2089 185
R17633 vdd.n2092 vdd.n1095 185
R17634 vdd.n2094 vdd.n2093 185
R17635 vdd.n2095 vdd.n1090 185
R17636 vdd.n2097 vdd.n2096 185
R17637 vdd.n2099 vdd.n1088 185
R17638 vdd.n2101 vdd.n2100 185
R17639 vdd.n2102 vdd.n1084 185
R17640 vdd.n2104 vdd.n2103 185
R17641 vdd.n2106 vdd.n1081 185
R17642 vdd.n2108 vdd.n2107 185
R17643 vdd.n1082 vdd.n1075 185
R17644 vdd.n2112 vdd.n1079 185
R17645 vdd.n2113 vdd.n1071 185
R17646 vdd.n2115 vdd.n2114 185
R17647 vdd.n2117 vdd.n1069 185
R17648 vdd.n2119 vdd.n2118 185
R17649 vdd.n2120 vdd.n1064 185
R17650 vdd.n2122 vdd.n2121 185
R17651 vdd.n2124 vdd.n1062 185
R17652 vdd.n2126 vdd.n2125 185
R17653 vdd.n2127 vdd.n1057 185
R17654 vdd.n2129 vdd.n2128 185
R17655 vdd.n2131 vdd.n1055 185
R17656 vdd.n2133 vdd.n2132 185
R17657 vdd.n2134 vdd.n1050 185
R17658 vdd.n2136 vdd.n2135 185
R17659 vdd.n2138 vdd.n1048 185
R17660 vdd.n2140 vdd.n2139 185
R17661 vdd.n2141 vdd.n1044 185
R17662 vdd.n2143 vdd.n2142 185
R17663 vdd.n2145 vdd.n1041 185
R17664 vdd.n2147 vdd.n2146 185
R17665 vdd.n1042 vdd.n1035 185
R17666 vdd.n2151 vdd.n1039 185
R17667 vdd.n2152 vdd.n1031 185
R17668 vdd.n2154 vdd.n2153 185
R17669 vdd.n2156 vdd.n1029 185
R17670 vdd.n2158 vdd.n2157 185
R17671 vdd.n2159 vdd.n1024 185
R17672 vdd.n2161 vdd.n2160 185
R17673 vdd.n2163 vdd.n1022 185
R17674 vdd.n2165 vdd.n2164 185
R17675 vdd.n2166 vdd.n1017 185
R17676 vdd.n2168 vdd.n2167 185
R17677 vdd.n2170 vdd.n1015 185
R17678 vdd.n2172 vdd.n2171 185
R17679 vdd.n2173 vdd.n1013 185
R17680 vdd.n2175 vdd.n2174 185
R17681 vdd.n2178 vdd.n2177 185
R17682 vdd.n2180 vdd.n2179 185
R17683 vdd.n2182 vdd.n1011 185
R17684 vdd.n2184 vdd.n2183 185
R17685 vdd.n1358 vdd.n1010 185
R17686 vdd.n2071 vdd.n1356 185
R17687 vdd.n2071 vdd.n2070 185
R17688 vdd.n1366 vdd.n1355 185
R17689 vdd.n2061 vdd.n1355 185
R17690 vdd.n2060 vdd.n2059 185
R17691 vdd.n2062 vdd.n2060 185
R17692 vdd.n1365 vdd.n1364 185
R17693 vdd.n1364 vdd.n1363 185
R17694 vdd.n2053 vdd.n2052 185
R17695 vdd.n2052 vdd.n2051 185
R17696 vdd.n1369 vdd.n1368 185
R17697 vdd.n2042 vdd.n1369 185
R17698 vdd.n2041 vdd.n2040 185
R17699 vdd.n2043 vdd.n2041 185
R17700 vdd.n1376 vdd.n1375 185
R17701 vdd.n1380 vdd.n1375 185
R17702 vdd.n2036 vdd.n2035 185
R17703 vdd.n2035 vdd.n2034 185
R17704 vdd.n1379 vdd.n1378 185
R17705 vdd.n2025 vdd.n1379 185
R17706 vdd.n2024 vdd.n2023 185
R17707 vdd.n2026 vdd.n2024 185
R17708 vdd.n1388 vdd.n1387 185
R17709 vdd.n1387 vdd.n1386 185
R17710 vdd.n2019 vdd.n2018 185
R17711 vdd.n2018 vdd.n2017 185
R17712 vdd.n1391 vdd.n1390 185
R17713 vdd.n1392 vdd.n1391 185
R17714 vdd.n1726 vdd.n1725 185
R17715 vdd.n1727 vdd.n1726 185
R17716 vdd.n1399 vdd.n1398 185
R17717 vdd.n1403 vdd.n1398 185
R17718 vdd.n1721 vdd.n1720 185
R17719 vdd.n1720 vdd.n1719 185
R17720 vdd.n1402 vdd.n1401 185
R17721 vdd.n1710 vdd.n1402 185
R17722 vdd.n1709 vdd.n1708 185
R17723 vdd.n1711 vdd.n1709 185
R17724 vdd.n1410 vdd.n1409 185
R17725 vdd.n1415 vdd.n1409 185
R17726 vdd.n1704 vdd.n1703 185
R17727 vdd.n1703 vdd.n1702 185
R17728 vdd.n1413 vdd.n1412 185
R17729 vdd.n1414 vdd.n1413 185
R17730 vdd.n1693 vdd.n1692 185
R17731 vdd.n1694 vdd.n1693 185
R17732 vdd.n1423 vdd.n1422 185
R17733 vdd.n1422 vdd.n1421 185
R17734 vdd.n1688 vdd.n1687 185
R17735 vdd.n1687 vdd.n1686 185
R17736 vdd.n1426 vdd.n1425 185
R17737 vdd.n1427 vdd.n1426 185
R17738 vdd.n1677 vdd.n1676 185
R17739 vdd.n1678 vdd.n1677 185
R17740 vdd.n1434 vdd.n1433 185
R17741 vdd.n1438 vdd.n1433 185
R17742 vdd.n1672 vdd.n1671 185
R17743 vdd.n1671 vdd.n1670 185
R17744 vdd.n828 vdd.n826 185
R17745 vdd.n2424 vdd.n826 185
R17746 vdd.n2346 vdd.n846 185
R17747 vdd.n846 vdd.n833 185
R17748 vdd.n2348 vdd.n2347 185
R17749 vdd.n2349 vdd.n2348 185
R17750 vdd.n2345 vdd.n845 185
R17751 vdd.n1227 vdd.n845 185
R17752 vdd.n2344 vdd.n2343 185
R17753 vdd.n2343 vdd.n2342 185
R17754 vdd.n848 vdd.n847 185
R17755 vdd.n849 vdd.n848 185
R17756 vdd.n2333 vdd.n2332 185
R17757 vdd.n2334 vdd.n2333 185
R17758 vdd.n2331 vdd.n859 185
R17759 vdd.n859 vdd.n856 185
R17760 vdd.n2330 vdd.n2329 185
R17761 vdd.n2329 vdd.n2328 185
R17762 vdd.n861 vdd.n860 185
R17763 vdd.n1253 vdd.n861 185
R17764 vdd.n2321 vdd.n2320 185
R17765 vdd.n2322 vdd.n2321 185
R17766 vdd.n2319 vdd.n869 185
R17767 vdd.n874 vdd.n869 185
R17768 vdd.n2318 vdd.n2317 185
R17769 vdd.n2317 vdd.n2316 185
R17770 vdd.n871 vdd.n870 185
R17771 vdd.n880 vdd.n871 185
R17772 vdd.n2309 vdd.n2308 185
R17773 vdd.n2310 vdd.n2309 185
R17774 vdd.n2307 vdd.n881 185
R17775 vdd.n1265 vdd.n881 185
R17776 vdd.n2306 vdd.n2305 185
R17777 vdd.n2305 vdd.n2304 185
R17778 vdd.n883 vdd.n882 185
R17779 vdd.n884 vdd.n883 185
R17780 vdd.n2297 vdd.n2296 185
R17781 vdd.n2298 vdd.n2297 185
R17782 vdd.n2295 vdd.n893 185
R17783 vdd.n893 vdd.n890 185
R17784 vdd.n2294 vdd.n2293 185
R17785 vdd.n2293 vdd.n2292 185
R17786 vdd.n895 vdd.n894 185
R17787 vdd.n904 vdd.n895 185
R17788 vdd.n2284 vdd.n2283 185
R17789 vdd.n2285 vdd.n2284 185
R17790 vdd.n2282 vdd.n905 185
R17791 vdd.n911 vdd.n905 185
R17792 vdd.n2281 vdd.n2280 185
R17793 vdd.n2280 vdd.n2279 185
R17794 vdd.n907 vdd.n906 185
R17795 vdd.n908 vdd.n907 185
R17796 vdd.n2272 vdd.n2271 185
R17797 vdd.n2273 vdd.n2272 185
R17798 vdd.n2270 vdd.n918 185
R17799 vdd.n918 vdd.n915 185
R17800 vdd.n2269 vdd.n2268 185
R17801 vdd.n2268 vdd.n2267 185
R17802 vdd.n920 vdd.n919 185
R17803 vdd.n921 vdd.n920 185
R17804 vdd.n2260 vdd.n2259 185
R17805 vdd.n2261 vdd.n2260 185
R17806 vdd.n2258 vdd.n929 185
R17807 vdd.n934 vdd.n929 185
R17808 vdd.n2257 vdd.n2256 185
R17809 vdd.n2256 vdd.n2255 185
R17810 vdd.n931 vdd.n930 185
R17811 vdd.n940 vdd.n931 185
R17812 vdd.n2248 vdd.n2247 185
R17813 vdd.n2249 vdd.n2248 185
R17814 vdd.n2246 vdd.n941 185
R17815 vdd.n947 vdd.n941 185
R17816 vdd.n2245 vdd.n2244 185
R17817 vdd.n2244 vdd.n2243 185
R17818 vdd.n943 vdd.n942 185
R17819 vdd.n944 vdd.n943 185
R17820 vdd.n2236 vdd.n2235 185
R17821 vdd.n2237 vdd.n2236 185
R17822 vdd.n2234 vdd.n954 185
R17823 vdd.n954 vdd.n951 185
R17824 vdd.n2233 vdd.n2232 185
R17825 vdd.n2232 vdd.n2231 185
R17826 vdd.n956 vdd.n955 185
R17827 vdd.n965 vdd.n956 185
R17828 vdd.n2224 vdd.n2223 185
R17829 vdd.n2225 vdd.n2224 185
R17830 vdd.n2222 vdd.n966 185
R17831 vdd.n966 vdd.n962 185
R17832 vdd.n2221 vdd.n2220 185
R17833 vdd.n968 vdd.n967 185
R17834 vdd.n2217 vdd.n2216 185
R17835 vdd.n2218 vdd.n2217 185
R17836 vdd.n2215 vdd.n1004 185
R17837 vdd.n2214 vdd.n2213 185
R17838 vdd.n2212 vdd.n2211 185
R17839 vdd.n2210 vdd.n2209 185
R17840 vdd.n2208 vdd.n2207 185
R17841 vdd.n2206 vdd.n2205 185
R17842 vdd.n2204 vdd.n2203 185
R17843 vdd.n2202 vdd.n2201 185
R17844 vdd.n2200 vdd.n2199 185
R17845 vdd.n2198 vdd.n2197 185
R17846 vdd.n2196 vdd.n2195 185
R17847 vdd.n2194 vdd.n2193 185
R17848 vdd.n2192 vdd.n2191 185
R17849 vdd.n2190 vdd.n2189 185
R17850 vdd.n2188 vdd.n2187 185
R17851 vdd.n1149 vdd.n1005 185
R17852 vdd.n1151 vdd.n1150 185
R17853 vdd.n1153 vdd.n1152 185
R17854 vdd.n1155 vdd.n1154 185
R17855 vdd.n1157 vdd.n1156 185
R17856 vdd.n1159 vdd.n1158 185
R17857 vdd.n1161 vdd.n1160 185
R17858 vdd.n1163 vdd.n1162 185
R17859 vdd.n1165 vdd.n1164 185
R17860 vdd.n1167 vdd.n1166 185
R17861 vdd.n1169 vdd.n1168 185
R17862 vdd.n1171 vdd.n1170 185
R17863 vdd.n1173 vdd.n1172 185
R17864 vdd.n1175 vdd.n1174 185
R17865 vdd.n1178 vdd.n1177 185
R17866 vdd.n1180 vdd.n1179 185
R17867 vdd.n1182 vdd.n1181 185
R17868 vdd.n2427 vdd.n2426 185
R17869 vdd.n2429 vdd.n2428 185
R17870 vdd.n2431 vdd.n2430 185
R17871 vdd.n2434 vdd.n2433 185
R17872 vdd.n2436 vdd.n2435 185
R17873 vdd.n2438 vdd.n2437 185
R17874 vdd.n2440 vdd.n2439 185
R17875 vdd.n2442 vdd.n2441 185
R17876 vdd.n2444 vdd.n2443 185
R17877 vdd.n2446 vdd.n2445 185
R17878 vdd.n2448 vdd.n2447 185
R17879 vdd.n2450 vdd.n2449 185
R17880 vdd.n2452 vdd.n2451 185
R17881 vdd.n2454 vdd.n2453 185
R17882 vdd.n2456 vdd.n2455 185
R17883 vdd.n2458 vdd.n2457 185
R17884 vdd.n2460 vdd.n2459 185
R17885 vdd.n2462 vdd.n2461 185
R17886 vdd.n2464 vdd.n2463 185
R17887 vdd.n2466 vdd.n2465 185
R17888 vdd.n2468 vdd.n2467 185
R17889 vdd.n2470 vdd.n2469 185
R17890 vdd.n2472 vdd.n2471 185
R17891 vdd.n2474 vdd.n2473 185
R17892 vdd.n2476 vdd.n2475 185
R17893 vdd.n2478 vdd.n2477 185
R17894 vdd.n2480 vdd.n2479 185
R17895 vdd.n2482 vdd.n2481 185
R17896 vdd.n2484 vdd.n2483 185
R17897 vdd.n2486 vdd.n2485 185
R17898 vdd.n2488 vdd.n2487 185
R17899 vdd.n2490 vdd.n2489 185
R17900 vdd.n2492 vdd.n2491 185
R17901 vdd.n2493 vdd.n827 185
R17902 vdd.n2495 vdd.n2494 185
R17903 vdd.n2496 vdd.n2495 185
R17904 vdd.n2425 vdd.n831 185
R17905 vdd.n2425 vdd.n2424 185
R17906 vdd.n1225 vdd.n832 185
R17907 vdd.n833 vdd.n832 185
R17908 vdd.n1226 vdd.n843 185
R17909 vdd.n2349 vdd.n843 185
R17910 vdd.n1229 vdd.n1228 185
R17911 vdd.n1228 vdd.n1227 185
R17912 vdd.n1230 vdd.n850 185
R17913 vdd.n2342 vdd.n850 185
R17914 vdd.n1232 vdd.n1231 185
R17915 vdd.n1231 vdd.n849 185
R17916 vdd.n1233 vdd.n857 185
R17917 vdd.n2334 vdd.n857 185
R17918 vdd.n1235 vdd.n1234 185
R17919 vdd.n1234 vdd.n856 185
R17920 vdd.n1236 vdd.n862 185
R17921 vdd.n2328 vdd.n862 185
R17922 vdd.n1255 vdd.n1254 185
R17923 vdd.n1254 vdd.n1253 185
R17924 vdd.n1256 vdd.n867 185
R17925 vdd.n2322 vdd.n867 185
R17926 vdd.n1258 vdd.n1257 185
R17927 vdd.n1257 vdd.n874 185
R17928 vdd.n1259 vdd.n872 185
R17929 vdd.n2316 vdd.n872 185
R17930 vdd.n1261 vdd.n1260 185
R17931 vdd.n1260 vdd.n880 185
R17932 vdd.n1262 vdd.n878 185
R17933 vdd.n2310 vdd.n878 185
R17934 vdd.n1264 vdd.n1263 185
R17935 vdd.n1265 vdd.n1264 185
R17936 vdd.n1224 vdd.n885 185
R17937 vdd.n2304 vdd.n885 185
R17938 vdd.n1223 vdd.n1222 185
R17939 vdd.n1222 vdd.n884 185
R17940 vdd.n1221 vdd.n891 185
R17941 vdd.n2298 vdd.n891 185
R17942 vdd.n1220 vdd.n1219 185
R17943 vdd.n1219 vdd.n890 185
R17944 vdd.n1218 vdd.n896 185
R17945 vdd.n2292 vdd.n896 185
R17946 vdd.n1217 vdd.n1216 185
R17947 vdd.n1216 vdd.n904 185
R17948 vdd.n1215 vdd.n902 185
R17949 vdd.n2285 vdd.n902 185
R17950 vdd.n1214 vdd.n1213 185
R17951 vdd.n1213 vdd.n911 185
R17952 vdd.n1212 vdd.n909 185
R17953 vdd.n2279 vdd.n909 185
R17954 vdd.n1211 vdd.n1210 185
R17955 vdd.n1210 vdd.n908 185
R17956 vdd.n1209 vdd.n916 185
R17957 vdd.n2273 vdd.n916 185
R17958 vdd.n1208 vdd.n1207 185
R17959 vdd.n1207 vdd.n915 185
R17960 vdd.n1206 vdd.n922 185
R17961 vdd.n2267 vdd.n922 185
R17962 vdd.n1205 vdd.n1204 185
R17963 vdd.n1204 vdd.n921 185
R17964 vdd.n1203 vdd.n927 185
R17965 vdd.n2261 vdd.n927 185
R17966 vdd.n1202 vdd.n1201 185
R17967 vdd.n1201 vdd.n934 185
R17968 vdd.n1200 vdd.n932 185
R17969 vdd.n2255 vdd.n932 185
R17970 vdd.n1199 vdd.n1198 185
R17971 vdd.n1198 vdd.n940 185
R17972 vdd.n1197 vdd.n938 185
R17973 vdd.n2249 vdd.n938 185
R17974 vdd.n1196 vdd.n1195 185
R17975 vdd.n1195 vdd.n947 185
R17976 vdd.n1194 vdd.n945 185
R17977 vdd.n2243 vdd.n945 185
R17978 vdd.n1193 vdd.n1192 185
R17979 vdd.n1192 vdd.n944 185
R17980 vdd.n1191 vdd.n952 185
R17981 vdd.n2237 vdd.n952 185
R17982 vdd.n1190 vdd.n1189 185
R17983 vdd.n1189 vdd.n951 185
R17984 vdd.n1188 vdd.n957 185
R17985 vdd.n2231 vdd.n957 185
R17986 vdd.n1187 vdd.n1186 185
R17987 vdd.n1186 vdd.n965 185
R17988 vdd.n1185 vdd.n963 185
R17989 vdd.n2225 vdd.n963 185
R17990 vdd.n1184 vdd.n1183 185
R17991 vdd.n1183 vdd.n962 185
R17992 vdd.n3409 vdd.n3408 185
R17993 vdd.n3410 vdd.n3409 185
R17994 vdd.n347 vdd.n346 185
R17995 vdd.n3411 vdd.n347 185
R17996 vdd.n3414 vdd.n3413 185
R17997 vdd.n3413 vdd.n3412 185
R17998 vdd.n3415 vdd.n341 185
R17999 vdd.n341 vdd.n340 185
R18000 vdd.n3417 vdd.n3416 185
R18001 vdd.n3418 vdd.n3417 185
R18002 vdd.n336 vdd.n335 185
R18003 vdd.n3419 vdd.n336 185
R18004 vdd.n3422 vdd.n3421 185
R18005 vdd.n3421 vdd.n3420 185
R18006 vdd.n3423 vdd.n330 185
R18007 vdd.n330 vdd.n329 185
R18008 vdd.n3425 vdd.n3424 185
R18009 vdd.n3426 vdd.n3425 185
R18010 vdd.n324 vdd.n323 185
R18011 vdd.n3427 vdd.n324 185
R18012 vdd.n3430 vdd.n3429 185
R18013 vdd.n3429 vdd.n3428 185
R18014 vdd.n3431 vdd.n319 185
R18015 vdd.n325 vdd.n319 185
R18016 vdd.n3433 vdd.n3432 185
R18017 vdd.n3434 vdd.n3433 185
R18018 vdd.n315 vdd.n313 185
R18019 vdd.n3435 vdd.n315 185
R18020 vdd.n3438 vdd.n3437 185
R18021 vdd.n3437 vdd.n3436 185
R18022 vdd.n314 vdd.n312 185
R18023 vdd.n481 vdd.n314 185
R18024 vdd.n3260 vdd.n3259 185
R18025 vdd.n3261 vdd.n3260 185
R18026 vdd.n483 vdd.n482 185
R18027 vdd.n3252 vdd.n482 185
R18028 vdd.n3255 vdd.n3254 185
R18029 vdd.n3254 vdd.n3253 185
R18030 vdd.n486 vdd.n485 185
R18031 vdd.n493 vdd.n486 185
R18032 vdd.n3243 vdd.n3242 185
R18033 vdd.n3244 vdd.n3243 185
R18034 vdd.n495 vdd.n494 185
R18035 vdd.n494 vdd.n492 185
R18036 vdd.n3238 vdd.n3237 185
R18037 vdd.n3237 vdd.n3236 185
R18038 vdd.n498 vdd.n497 185
R18039 vdd.n499 vdd.n498 185
R18040 vdd.n3227 vdd.n3226 185
R18041 vdd.n3228 vdd.n3227 185
R18042 vdd.n507 vdd.n506 185
R18043 vdd.n506 vdd.n505 185
R18044 vdd.n3222 vdd.n3221 185
R18045 vdd.n3221 vdd.n3220 185
R18046 vdd.n510 vdd.n509 185
R18047 vdd.n511 vdd.n510 185
R18048 vdd.n3211 vdd.n3210 185
R18049 vdd.n3212 vdd.n3211 185
R18050 vdd.n3207 vdd.n517 185
R18051 vdd.n3206 vdd.n3205 185
R18052 vdd.n3203 vdd.n519 185
R18053 vdd.n3203 vdd.n516 185
R18054 vdd.n3202 vdd.n3201 185
R18055 vdd.n3200 vdd.n3199 185
R18056 vdd.n3198 vdd.n3197 185
R18057 vdd.n3196 vdd.n3195 185
R18058 vdd.n3194 vdd.n525 185
R18059 vdd.n3192 vdd.n3191 185
R18060 vdd.n3190 vdd.n526 185
R18061 vdd.n3189 vdd.n3188 185
R18062 vdd.n3186 vdd.n531 185
R18063 vdd.n3184 vdd.n3183 185
R18064 vdd.n3182 vdd.n532 185
R18065 vdd.n3181 vdd.n3180 185
R18066 vdd.n3178 vdd.n537 185
R18067 vdd.n3176 vdd.n3175 185
R18068 vdd.n3174 vdd.n538 185
R18069 vdd.n3173 vdd.n3172 185
R18070 vdd.n3170 vdd.n545 185
R18071 vdd.n3168 vdd.n3167 185
R18072 vdd.n3166 vdd.n546 185
R18073 vdd.n3165 vdd.n3164 185
R18074 vdd.n3162 vdd.n551 185
R18075 vdd.n3160 vdd.n3159 185
R18076 vdd.n3158 vdd.n552 185
R18077 vdd.n3157 vdd.n3156 185
R18078 vdd.n3154 vdd.n557 185
R18079 vdd.n3152 vdd.n3151 185
R18080 vdd.n3150 vdd.n558 185
R18081 vdd.n3149 vdd.n3148 185
R18082 vdd.n3146 vdd.n563 185
R18083 vdd.n3144 vdd.n3143 185
R18084 vdd.n3142 vdd.n564 185
R18085 vdd.n3141 vdd.n3140 185
R18086 vdd.n3138 vdd.n569 185
R18087 vdd.n3136 vdd.n3135 185
R18088 vdd.n3134 vdd.n570 185
R18089 vdd.n3133 vdd.n3132 185
R18090 vdd.n3130 vdd.n575 185
R18091 vdd.n3128 vdd.n3127 185
R18092 vdd.n3126 vdd.n576 185
R18093 vdd.n585 vdd.n579 185
R18094 vdd.n3122 vdd.n3121 185
R18095 vdd.n3119 vdd.n583 185
R18096 vdd.n3118 vdd.n3117 185
R18097 vdd.n3116 vdd.n3115 185
R18098 vdd.n3114 vdd.n589 185
R18099 vdd.n3112 vdd.n3111 185
R18100 vdd.n3110 vdd.n590 185
R18101 vdd.n3109 vdd.n3108 185
R18102 vdd.n3106 vdd.n595 185
R18103 vdd.n3104 vdd.n3103 185
R18104 vdd.n3102 vdd.n596 185
R18105 vdd.n3101 vdd.n3100 185
R18106 vdd.n3098 vdd.n601 185
R18107 vdd.n3096 vdd.n3095 185
R18108 vdd.n3094 vdd.n602 185
R18109 vdd.n3093 vdd.n3092 185
R18110 vdd.n3090 vdd.n3089 185
R18111 vdd.n3088 vdd.n3087 185
R18112 vdd.n3086 vdd.n3085 185
R18113 vdd.n3084 vdd.n3083 185
R18114 vdd.n3079 vdd.n515 185
R18115 vdd.n516 vdd.n515 185
R18116 vdd.n3292 vdd.n3291 185
R18117 vdd.n3296 vdd.n462 185
R18118 vdd.n3298 vdd.n3297 185
R18119 vdd.n3300 vdd.n460 185
R18120 vdd.n3302 vdd.n3301 185
R18121 vdd.n3303 vdd.n455 185
R18122 vdd.n3305 vdd.n3304 185
R18123 vdd.n3307 vdd.n453 185
R18124 vdd.n3309 vdd.n3308 185
R18125 vdd.n3310 vdd.n448 185
R18126 vdd.n3312 vdd.n3311 185
R18127 vdd.n3314 vdd.n446 185
R18128 vdd.n3316 vdd.n3315 185
R18129 vdd.n3317 vdd.n441 185
R18130 vdd.n3319 vdd.n3318 185
R18131 vdd.n3321 vdd.n439 185
R18132 vdd.n3323 vdd.n3322 185
R18133 vdd.n3324 vdd.n435 185
R18134 vdd.n3326 vdd.n3325 185
R18135 vdd.n3328 vdd.n432 185
R18136 vdd.n3330 vdd.n3329 185
R18137 vdd.n433 vdd.n426 185
R18138 vdd.n3334 vdd.n430 185
R18139 vdd.n3335 vdd.n422 185
R18140 vdd.n3337 vdd.n3336 185
R18141 vdd.n3339 vdd.n420 185
R18142 vdd.n3341 vdd.n3340 185
R18143 vdd.n3342 vdd.n415 185
R18144 vdd.n3344 vdd.n3343 185
R18145 vdd.n3346 vdd.n413 185
R18146 vdd.n3348 vdd.n3347 185
R18147 vdd.n3349 vdd.n408 185
R18148 vdd.n3351 vdd.n3350 185
R18149 vdd.n3353 vdd.n406 185
R18150 vdd.n3355 vdd.n3354 185
R18151 vdd.n3356 vdd.n401 185
R18152 vdd.n3358 vdd.n3357 185
R18153 vdd.n3360 vdd.n399 185
R18154 vdd.n3362 vdd.n3361 185
R18155 vdd.n3363 vdd.n395 185
R18156 vdd.n3365 vdd.n3364 185
R18157 vdd.n3367 vdd.n392 185
R18158 vdd.n3369 vdd.n3368 185
R18159 vdd.n393 vdd.n386 185
R18160 vdd.n3373 vdd.n390 185
R18161 vdd.n3374 vdd.n382 185
R18162 vdd.n3376 vdd.n3375 185
R18163 vdd.n3378 vdd.n380 185
R18164 vdd.n3380 vdd.n3379 185
R18165 vdd.n3381 vdd.n375 185
R18166 vdd.n3383 vdd.n3382 185
R18167 vdd.n3385 vdd.n373 185
R18168 vdd.n3387 vdd.n3386 185
R18169 vdd.n3388 vdd.n368 185
R18170 vdd.n3390 vdd.n3389 185
R18171 vdd.n3392 vdd.n366 185
R18172 vdd.n3394 vdd.n3393 185
R18173 vdd.n3395 vdd.n360 185
R18174 vdd.n3397 vdd.n3396 185
R18175 vdd.n3399 vdd.n359 185
R18176 vdd.n3400 vdd.n358 185
R18177 vdd.n3403 vdd.n3402 185
R18178 vdd.n3404 vdd.n356 185
R18179 vdd.n3405 vdd.n352 185
R18180 vdd.n3287 vdd.n350 185
R18181 vdd.n3410 vdd.n350 185
R18182 vdd.n3286 vdd.n349 185
R18183 vdd.n3411 vdd.n349 185
R18184 vdd.n3285 vdd.n348 185
R18185 vdd.n3412 vdd.n348 185
R18186 vdd.n468 vdd.n467 185
R18187 vdd.n467 vdd.n340 185
R18188 vdd.n3281 vdd.n339 185
R18189 vdd.n3418 vdd.n339 185
R18190 vdd.n3280 vdd.n338 185
R18191 vdd.n3419 vdd.n338 185
R18192 vdd.n3279 vdd.n337 185
R18193 vdd.n3420 vdd.n337 185
R18194 vdd.n471 vdd.n470 185
R18195 vdd.n470 vdd.n329 185
R18196 vdd.n3275 vdd.n328 185
R18197 vdd.n3426 vdd.n328 185
R18198 vdd.n3274 vdd.n327 185
R18199 vdd.n3427 vdd.n327 185
R18200 vdd.n3273 vdd.n326 185
R18201 vdd.n3428 vdd.n326 185
R18202 vdd.n474 vdd.n473 185
R18203 vdd.n473 vdd.n325 185
R18204 vdd.n3269 vdd.n318 185
R18205 vdd.n3434 vdd.n318 185
R18206 vdd.n3268 vdd.n317 185
R18207 vdd.n3435 vdd.n317 185
R18208 vdd.n3267 vdd.n316 185
R18209 vdd.n3436 vdd.n316 185
R18210 vdd.n480 vdd.n476 185
R18211 vdd.n481 vdd.n480 185
R18212 vdd.n3263 vdd.n3262 185
R18213 vdd.n3262 vdd.n3261 185
R18214 vdd.n479 vdd.n478 185
R18215 vdd.n3252 vdd.n479 185
R18216 vdd.n3251 vdd.n3250 185
R18217 vdd.n3253 vdd.n3251 185
R18218 vdd.n488 vdd.n487 185
R18219 vdd.n493 vdd.n487 185
R18220 vdd.n3246 vdd.n3245 185
R18221 vdd.n3245 vdd.n3244 185
R18222 vdd.n491 vdd.n490 185
R18223 vdd.n492 vdd.n491 185
R18224 vdd.n3235 vdd.n3234 185
R18225 vdd.n3236 vdd.n3235 185
R18226 vdd.n501 vdd.n500 185
R18227 vdd.n500 vdd.n499 185
R18228 vdd.n3230 vdd.n3229 185
R18229 vdd.n3229 vdd.n3228 185
R18230 vdd.n504 vdd.n503 185
R18231 vdd.n505 vdd.n504 185
R18232 vdd.n3219 vdd.n3218 185
R18233 vdd.n3220 vdd.n3219 185
R18234 vdd.n513 vdd.n512 185
R18235 vdd.n512 vdd.n511 185
R18236 vdd.n3214 vdd.n3213 185
R18237 vdd.n3213 vdd.n3212 185
R18238 vdd.n2803 vdd.n2802 185
R18239 vdd.n790 vdd.n789 185
R18240 vdd.n2799 vdd.n2798 185
R18241 vdd.n2800 vdd.n2799 185
R18242 vdd.n2797 vdd.n2531 185
R18243 vdd.n2796 vdd.n2795 185
R18244 vdd.n2794 vdd.n2793 185
R18245 vdd.n2792 vdd.n2791 185
R18246 vdd.n2790 vdd.n2789 185
R18247 vdd.n2788 vdd.n2787 185
R18248 vdd.n2786 vdd.n2785 185
R18249 vdd.n2784 vdd.n2783 185
R18250 vdd.n2782 vdd.n2781 185
R18251 vdd.n2780 vdd.n2779 185
R18252 vdd.n2778 vdd.n2777 185
R18253 vdd.n2776 vdd.n2775 185
R18254 vdd.n2774 vdd.n2773 185
R18255 vdd.n2772 vdd.n2771 185
R18256 vdd.n2770 vdd.n2769 185
R18257 vdd.n2768 vdd.n2767 185
R18258 vdd.n2766 vdd.n2765 185
R18259 vdd.n2764 vdd.n2763 185
R18260 vdd.n2762 vdd.n2761 185
R18261 vdd.n2760 vdd.n2759 185
R18262 vdd.n2758 vdd.n2757 185
R18263 vdd.n2756 vdd.n2755 185
R18264 vdd.n2754 vdd.n2753 185
R18265 vdd.n2752 vdd.n2751 185
R18266 vdd.n2750 vdd.n2749 185
R18267 vdd.n2748 vdd.n2747 185
R18268 vdd.n2746 vdd.n2745 185
R18269 vdd.n2744 vdd.n2743 185
R18270 vdd.n2742 vdd.n2741 185
R18271 vdd.n2739 vdd.n2738 185
R18272 vdd.n2737 vdd.n2736 185
R18273 vdd.n2735 vdd.n2734 185
R18274 vdd.n2980 vdd.n2979 185
R18275 vdd.n2981 vdd.n660 185
R18276 vdd.n2983 vdd.n2982 185
R18277 vdd.n2985 vdd.n658 185
R18278 vdd.n2987 vdd.n2986 185
R18279 vdd.n2988 vdd.n657 185
R18280 vdd.n2990 vdd.n2989 185
R18281 vdd.n2992 vdd.n655 185
R18282 vdd.n2994 vdd.n2993 185
R18283 vdd.n2995 vdd.n654 185
R18284 vdd.n2997 vdd.n2996 185
R18285 vdd.n2999 vdd.n652 185
R18286 vdd.n3001 vdd.n3000 185
R18287 vdd.n3002 vdd.n651 185
R18288 vdd.n3004 vdd.n3003 185
R18289 vdd.n3006 vdd.n649 185
R18290 vdd.n3008 vdd.n3007 185
R18291 vdd.n3010 vdd.n648 185
R18292 vdd.n3012 vdd.n3011 185
R18293 vdd.n3014 vdd.n646 185
R18294 vdd.n3016 vdd.n3015 185
R18295 vdd.n3017 vdd.n645 185
R18296 vdd.n3019 vdd.n3018 185
R18297 vdd.n3021 vdd.n643 185
R18298 vdd.n3023 vdd.n3022 185
R18299 vdd.n3024 vdd.n642 185
R18300 vdd.n3026 vdd.n3025 185
R18301 vdd.n3028 vdd.n640 185
R18302 vdd.n3030 vdd.n3029 185
R18303 vdd.n3031 vdd.n639 185
R18304 vdd.n3033 vdd.n3032 185
R18305 vdd.n3035 vdd.n638 185
R18306 vdd.n3036 vdd.n637 185
R18307 vdd.n3039 vdd.n3038 185
R18308 vdd.n3040 vdd.n635 185
R18309 vdd.n635 vdd.n613 185
R18310 vdd.n2977 vdd.n632 185
R18311 vdd.n3043 vdd.n632 185
R18312 vdd.n2976 vdd.n2975 185
R18313 vdd.n2975 vdd.n631 185
R18314 vdd.n2974 vdd.n664 185
R18315 vdd.n2974 vdd.n2973 185
R18316 vdd.n2617 vdd.n665 185
R18317 vdd.n674 vdd.n665 185
R18318 vdd.n2618 vdd.n672 185
R18319 vdd.n2967 vdd.n672 185
R18320 vdd.n2620 vdd.n2619 185
R18321 vdd.n2619 vdd.n671 185
R18322 vdd.n2621 vdd.n680 185
R18323 vdd.n2916 vdd.n680 185
R18324 vdd.n2623 vdd.n2622 185
R18325 vdd.n2622 vdd.n679 185
R18326 vdd.n2624 vdd.n685 185
R18327 vdd.n2910 vdd.n685 185
R18328 vdd.n2626 vdd.n2625 185
R18329 vdd.n2625 vdd.n692 185
R18330 vdd.n2627 vdd.n690 185
R18331 vdd.n2904 vdd.n690 185
R18332 vdd.n2629 vdd.n2628 185
R18333 vdd.n2628 vdd.n698 185
R18334 vdd.n2630 vdd.n696 185
R18335 vdd.n2898 vdd.n696 185
R18336 vdd.n2632 vdd.n2631 185
R18337 vdd.n2631 vdd.n705 185
R18338 vdd.n2633 vdd.n703 185
R18339 vdd.n2892 vdd.n703 185
R18340 vdd.n2635 vdd.n2634 185
R18341 vdd.n2634 vdd.n702 185
R18342 vdd.n2636 vdd.n710 185
R18343 vdd.n2886 vdd.n710 185
R18344 vdd.n2638 vdd.n2637 185
R18345 vdd.n2637 vdd.n709 185
R18346 vdd.n2639 vdd.n716 185
R18347 vdd.n2880 vdd.n716 185
R18348 vdd.n2641 vdd.n2640 185
R18349 vdd.n2640 vdd.n715 185
R18350 vdd.n2642 vdd.n721 185
R18351 vdd.n2874 vdd.n721 185
R18352 vdd.n2644 vdd.n2643 185
R18353 vdd.n2643 vdd.n729 185
R18354 vdd.n2645 vdd.n727 185
R18355 vdd.n2868 vdd.n727 185
R18356 vdd.n2647 vdd.n2646 185
R18357 vdd.n2646 vdd.n736 185
R18358 vdd.n2648 vdd.n734 185
R18359 vdd.n2862 vdd.n734 185
R18360 vdd.n2650 vdd.n2649 185
R18361 vdd.n2649 vdd.n733 185
R18362 vdd.n2651 vdd.n741 185
R18363 vdd.n2855 vdd.n741 185
R18364 vdd.n2653 vdd.n2652 185
R18365 vdd.n2652 vdd.n740 185
R18366 vdd.n2654 vdd.n746 185
R18367 vdd.n2849 vdd.n746 185
R18368 vdd.n2656 vdd.n2655 185
R18369 vdd.n2655 vdd.n753 185
R18370 vdd.n2657 vdd.n751 185
R18371 vdd.n2843 vdd.n751 185
R18372 vdd.n2659 vdd.n2658 185
R18373 vdd.n2658 vdd.n759 185
R18374 vdd.n2660 vdd.n757 185
R18375 vdd.n2837 vdd.n757 185
R18376 vdd.n2712 vdd.n2711 185
R18377 vdd.n2711 vdd.n2710 185
R18378 vdd.n2713 vdd.n763 185
R18379 vdd.n2831 vdd.n763 185
R18380 vdd.n2715 vdd.n2714 185
R18381 vdd.n2716 vdd.n2715 185
R18382 vdd.n2616 vdd.n769 185
R18383 vdd.n2825 vdd.n769 185
R18384 vdd.n2615 vdd.n2614 185
R18385 vdd.n2614 vdd.n768 185
R18386 vdd.n2613 vdd.n775 185
R18387 vdd.n2819 vdd.n775 185
R18388 vdd.n2612 vdd.n2611 185
R18389 vdd.n2611 vdd.n774 185
R18390 vdd.n2534 vdd.n780 185
R18391 vdd.n2813 vdd.n780 185
R18392 vdd.n2730 vdd.n2729 185
R18393 vdd.n2729 vdd.n2728 185
R18394 vdd.n2731 vdd.n786 185
R18395 vdd.n2807 vdd.n786 185
R18396 vdd.n2733 vdd.n2732 185
R18397 vdd.n2733 vdd.n785 185
R18398 vdd.n2804 vdd.n788 185
R18399 vdd.n788 vdd.n785 185
R18400 vdd.n2806 vdd.n2805 185
R18401 vdd.n2807 vdd.n2806 185
R18402 vdd.n779 vdd.n778 185
R18403 vdd.n2728 vdd.n779 185
R18404 vdd.n2815 vdd.n2814 185
R18405 vdd.n2814 vdd.n2813 185
R18406 vdd.n2816 vdd.n777 185
R18407 vdd.n777 vdd.n774 185
R18408 vdd.n2818 vdd.n2817 185
R18409 vdd.n2819 vdd.n2818 185
R18410 vdd.n767 vdd.n766 185
R18411 vdd.n768 vdd.n767 185
R18412 vdd.n2827 vdd.n2826 185
R18413 vdd.n2826 vdd.n2825 185
R18414 vdd.n2828 vdd.n765 185
R18415 vdd.n2716 vdd.n765 185
R18416 vdd.n2830 vdd.n2829 185
R18417 vdd.n2831 vdd.n2830 185
R18418 vdd.n756 vdd.n755 185
R18419 vdd.n2710 vdd.n756 185
R18420 vdd.n2839 vdd.n2838 185
R18421 vdd.n2838 vdd.n2837 185
R18422 vdd.n2840 vdd.n754 185
R18423 vdd.n759 vdd.n754 185
R18424 vdd.n2842 vdd.n2841 185
R18425 vdd.n2843 vdd.n2842 185
R18426 vdd.n745 vdd.n744 185
R18427 vdd.n753 vdd.n745 185
R18428 vdd.n2851 vdd.n2850 185
R18429 vdd.n2850 vdd.n2849 185
R18430 vdd.n2852 vdd.n743 185
R18431 vdd.n743 vdd.n740 185
R18432 vdd.n2854 vdd.n2853 185
R18433 vdd.n2855 vdd.n2854 185
R18434 vdd.n732 vdd.n731 185
R18435 vdd.n733 vdd.n732 185
R18436 vdd.n2864 vdd.n2863 185
R18437 vdd.n2863 vdd.n2862 185
R18438 vdd.n2865 vdd.n730 185
R18439 vdd.n736 vdd.n730 185
R18440 vdd.n2867 vdd.n2866 185
R18441 vdd.n2868 vdd.n2867 185
R18442 vdd.n720 vdd.n719 185
R18443 vdd.n729 vdd.n720 185
R18444 vdd.n2876 vdd.n2875 185
R18445 vdd.n2875 vdd.n2874 185
R18446 vdd.n2877 vdd.n718 185
R18447 vdd.n718 vdd.n715 185
R18448 vdd.n2879 vdd.n2878 185
R18449 vdd.n2880 vdd.n2879 185
R18450 vdd.n708 vdd.n707 185
R18451 vdd.n709 vdd.n708 185
R18452 vdd.n2888 vdd.n2887 185
R18453 vdd.n2887 vdd.n2886 185
R18454 vdd.n2889 vdd.n706 185
R18455 vdd.n706 vdd.n702 185
R18456 vdd.n2891 vdd.n2890 185
R18457 vdd.n2892 vdd.n2891 185
R18458 vdd.n695 vdd.n694 185
R18459 vdd.n705 vdd.n695 185
R18460 vdd.n2900 vdd.n2899 185
R18461 vdd.n2899 vdd.n2898 185
R18462 vdd.n2901 vdd.n693 185
R18463 vdd.n698 vdd.n693 185
R18464 vdd.n2903 vdd.n2902 185
R18465 vdd.n2904 vdd.n2903 185
R18466 vdd.n684 vdd.n683 185
R18467 vdd.n692 vdd.n684 185
R18468 vdd.n2912 vdd.n2911 185
R18469 vdd.n2911 vdd.n2910 185
R18470 vdd.n2913 vdd.n682 185
R18471 vdd.n682 vdd.n679 185
R18472 vdd.n2915 vdd.n2914 185
R18473 vdd.n2916 vdd.n2915 185
R18474 vdd.n670 vdd.n669 185
R18475 vdd.n671 vdd.n670 185
R18476 vdd.n2969 vdd.n2968 185
R18477 vdd.n2968 vdd.n2967 185
R18478 vdd.n2970 vdd.n668 185
R18479 vdd.n674 vdd.n668 185
R18480 vdd.n2972 vdd.n2971 185
R18481 vdd.n2973 vdd.n2972 185
R18482 vdd.n636 vdd.n634 185
R18483 vdd.n634 vdd.n631 185
R18484 vdd.n3042 vdd.n3041 185
R18485 vdd.n3043 vdd.n3042 185
R18486 vdd.n2423 vdd.n2422 185
R18487 vdd.n2424 vdd.n2423 185
R18488 vdd.n837 vdd.n835 185
R18489 vdd.n835 vdd.n833 185
R18490 vdd.n2338 vdd.n844 185
R18491 vdd.n2349 vdd.n844 185
R18492 vdd.n2339 vdd.n853 185
R18493 vdd.n1227 vdd.n853 185
R18494 vdd.n2341 vdd.n2340 185
R18495 vdd.n2342 vdd.n2341 185
R18496 vdd.n2337 vdd.n852 185
R18497 vdd.n852 vdd.n849 185
R18498 vdd.n2336 vdd.n2335 185
R18499 vdd.n2335 vdd.n2334 185
R18500 vdd.n855 vdd.n854 185
R18501 vdd.n856 vdd.n855 185
R18502 vdd.n2327 vdd.n2326 185
R18503 vdd.n2328 vdd.n2327 185
R18504 vdd.n2325 vdd.n864 185
R18505 vdd.n1253 vdd.n864 185
R18506 vdd.n2324 vdd.n2323 185
R18507 vdd.n2323 vdd.n2322 185
R18508 vdd.n866 vdd.n865 185
R18509 vdd.n874 vdd.n866 185
R18510 vdd.n2315 vdd.n2314 185
R18511 vdd.n2316 vdd.n2315 185
R18512 vdd.n2313 vdd.n875 185
R18513 vdd.n880 vdd.n875 185
R18514 vdd.n2312 vdd.n2311 185
R18515 vdd.n2311 vdd.n2310 185
R18516 vdd.n877 vdd.n876 185
R18517 vdd.n1265 vdd.n877 185
R18518 vdd.n2303 vdd.n2302 185
R18519 vdd.n2304 vdd.n2303 185
R18520 vdd.n2301 vdd.n887 185
R18521 vdd.n887 vdd.n884 185
R18522 vdd.n2300 vdd.n2299 185
R18523 vdd.n2299 vdd.n2298 185
R18524 vdd.n889 vdd.n888 185
R18525 vdd.n890 vdd.n889 185
R18526 vdd.n2291 vdd.n2290 185
R18527 vdd.n2292 vdd.n2291 185
R18528 vdd.n2288 vdd.n898 185
R18529 vdd.n904 vdd.n898 185
R18530 vdd.n2287 vdd.n2286 185
R18531 vdd.n2286 vdd.n2285 185
R18532 vdd.n901 vdd.n900 185
R18533 vdd.n911 vdd.n901 185
R18534 vdd.n2278 vdd.n2277 185
R18535 vdd.n2279 vdd.n2278 185
R18536 vdd.n2276 vdd.n912 185
R18537 vdd.n912 vdd.n908 185
R18538 vdd.n2275 vdd.n2274 185
R18539 vdd.n2274 vdd.n2273 185
R18540 vdd.n914 vdd.n913 185
R18541 vdd.n915 vdd.n914 185
R18542 vdd.n2266 vdd.n2265 185
R18543 vdd.n2267 vdd.n2266 185
R18544 vdd.n2264 vdd.n924 185
R18545 vdd.n924 vdd.n921 185
R18546 vdd.n2263 vdd.n2262 185
R18547 vdd.n2262 vdd.n2261 185
R18548 vdd.n926 vdd.n925 185
R18549 vdd.n934 vdd.n926 185
R18550 vdd.n2254 vdd.n2253 185
R18551 vdd.n2255 vdd.n2254 185
R18552 vdd.n2252 vdd.n935 185
R18553 vdd.n940 vdd.n935 185
R18554 vdd.n2251 vdd.n2250 185
R18555 vdd.n2250 vdd.n2249 185
R18556 vdd.n937 vdd.n936 185
R18557 vdd.n947 vdd.n937 185
R18558 vdd.n2242 vdd.n2241 185
R18559 vdd.n2243 vdd.n2242 185
R18560 vdd.n2240 vdd.n948 185
R18561 vdd.n948 vdd.n944 185
R18562 vdd.n2239 vdd.n2238 185
R18563 vdd.n2238 vdd.n2237 185
R18564 vdd.n950 vdd.n949 185
R18565 vdd.n951 vdd.n950 185
R18566 vdd.n2230 vdd.n2229 185
R18567 vdd.n2231 vdd.n2230 185
R18568 vdd.n2228 vdd.n959 185
R18569 vdd.n965 vdd.n959 185
R18570 vdd.n2227 vdd.n2226 185
R18571 vdd.n2226 vdd.n2225 185
R18572 vdd.n961 vdd.n960 185
R18573 vdd.n962 vdd.n961 185
R18574 vdd.n2354 vdd.n808 185
R18575 vdd.n2496 vdd.n808 185
R18576 vdd.n2356 vdd.n2355 185
R18577 vdd.n2358 vdd.n2357 185
R18578 vdd.n2360 vdd.n2359 185
R18579 vdd.n2362 vdd.n2361 185
R18580 vdd.n2364 vdd.n2363 185
R18581 vdd.n2366 vdd.n2365 185
R18582 vdd.n2368 vdd.n2367 185
R18583 vdd.n2370 vdd.n2369 185
R18584 vdd.n2372 vdd.n2371 185
R18585 vdd.n2374 vdd.n2373 185
R18586 vdd.n2376 vdd.n2375 185
R18587 vdd.n2378 vdd.n2377 185
R18588 vdd.n2380 vdd.n2379 185
R18589 vdd.n2382 vdd.n2381 185
R18590 vdd.n2384 vdd.n2383 185
R18591 vdd.n2386 vdd.n2385 185
R18592 vdd.n2388 vdd.n2387 185
R18593 vdd.n2390 vdd.n2389 185
R18594 vdd.n2392 vdd.n2391 185
R18595 vdd.n2394 vdd.n2393 185
R18596 vdd.n2396 vdd.n2395 185
R18597 vdd.n2398 vdd.n2397 185
R18598 vdd.n2400 vdd.n2399 185
R18599 vdd.n2402 vdd.n2401 185
R18600 vdd.n2404 vdd.n2403 185
R18601 vdd.n2406 vdd.n2405 185
R18602 vdd.n2408 vdd.n2407 185
R18603 vdd.n2410 vdd.n2409 185
R18604 vdd.n2412 vdd.n2411 185
R18605 vdd.n2414 vdd.n2413 185
R18606 vdd.n2416 vdd.n2415 185
R18607 vdd.n2418 vdd.n2417 185
R18608 vdd.n2420 vdd.n2419 185
R18609 vdd.n2421 vdd.n836 185
R18610 vdd.n2353 vdd.n834 185
R18611 vdd.n2424 vdd.n834 185
R18612 vdd.n2352 vdd.n2351 185
R18613 vdd.n2351 vdd.n833 185
R18614 vdd.n2350 vdd.n841 185
R18615 vdd.n2350 vdd.n2349 185
R18616 vdd.n1243 vdd.n842 185
R18617 vdd.n1227 vdd.n842 185
R18618 vdd.n1244 vdd.n851 185
R18619 vdd.n2342 vdd.n851 185
R18620 vdd.n1246 vdd.n1245 185
R18621 vdd.n1245 vdd.n849 185
R18622 vdd.n1247 vdd.n858 185
R18623 vdd.n2334 vdd.n858 185
R18624 vdd.n1249 vdd.n1248 185
R18625 vdd.n1248 vdd.n856 185
R18626 vdd.n1250 vdd.n863 185
R18627 vdd.n2328 vdd.n863 185
R18628 vdd.n1252 vdd.n1251 185
R18629 vdd.n1253 vdd.n1252 185
R18630 vdd.n1242 vdd.n868 185
R18631 vdd.n2322 vdd.n868 185
R18632 vdd.n1241 vdd.n1240 185
R18633 vdd.n1240 vdd.n874 185
R18634 vdd.n1239 vdd.n873 185
R18635 vdd.n2316 vdd.n873 185
R18636 vdd.n1238 vdd.n1237 185
R18637 vdd.n1237 vdd.n880 185
R18638 vdd.n1146 vdd.n879 185
R18639 vdd.n2310 vdd.n879 185
R18640 vdd.n1267 vdd.n1266 185
R18641 vdd.n1266 vdd.n1265 185
R18642 vdd.n1268 vdd.n886 185
R18643 vdd.n2304 vdd.n886 185
R18644 vdd.n1270 vdd.n1269 185
R18645 vdd.n1269 vdd.n884 185
R18646 vdd.n1271 vdd.n892 185
R18647 vdd.n2298 vdd.n892 185
R18648 vdd.n1273 vdd.n1272 185
R18649 vdd.n1272 vdd.n890 185
R18650 vdd.n1274 vdd.n897 185
R18651 vdd.n2292 vdd.n897 185
R18652 vdd.n1276 vdd.n1275 185
R18653 vdd.n1275 vdd.n904 185
R18654 vdd.n1277 vdd.n903 185
R18655 vdd.n2285 vdd.n903 185
R18656 vdd.n1279 vdd.n1278 185
R18657 vdd.n1278 vdd.n911 185
R18658 vdd.n1280 vdd.n910 185
R18659 vdd.n2279 vdd.n910 185
R18660 vdd.n1282 vdd.n1281 185
R18661 vdd.n1281 vdd.n908 185
R18662 vdd.n1283 vdd.n917 185
R18663 vdd.n2273 vdd.n917 185
R18664 vdd.n1285 vdd.n1284 185
R18665 vdd.n1284 vdd.n915 185
R18666 vdd.n1286 vdd.n923 185
R18667 vdd.n2267 vdd.n923 185
R18668 vdd.n1288 vdd.n1287 185
R18669 vdd.n1287 vdd.n921 185
R18670 vdd.n1289 vdd.n928 185
R18671 vdd.n2261 vdd.n928 185
R18672 vdd.n1291 vdd.n1290 185
R18673 vdd.n1290 vdd.n934 185
R18674 vdd.n1292 vdd.n933 185
R18675 vdd.n2255 vdd.n933 185
R18676 vdd.n1294 vdd.n1293 185
R18677 vdd.n1293 vdd.n940 185
R18678 vdd.n1295 vdd.n939 185
R18679 vdd.n2249 vdd.n939 185
R18680 vdd.n1297 vdd.n1296 185
R18681 vdd.n1296 vdd.n947 185
R18682 vdd.n1298 vdd.n946 185
R18683 vdd.n2243 vdd.n946 185
R18684 vdd.n1300 vdd.n1299 185
R18685 vdd.n1299 vdd.n944 185
R18686 vdd.n1301 vdd.n953 185
R18687 vdd.n2237 vdd.n953 185
R18688 vdd.n1303 vdd.n1302 185
R18689 vdd.n1302 vdd.n951 185
R18690 vdd.n1304 vdd.n958 185
R18691 vdd.n2231 vdd.n958 185
R18692 vdd.n1306 vdd.n1305 185
R18693 vdd.n1305 vdd.n965 185
R18694 vdd.n1307 vdd.n964 185
R18695 vdd.n2225 vdd.n964 185
R18696 vdd.n1309 vdd.n1308 185
R18697 vdd.n1308 vdd.n962 185
R18698 vdd.n1109 vdd.n1108 185
R18699 vdd.n1111 vdd.n1110 185
R18700 vdd.n1113 vdd.n1112 185
R18701 vdd.n1115 vdd.n1114 185
R18702 vdd.n1117 vdd.n1116 185
R18703 vdd.n1119 vdd.n1118 185
R18704 vdd.n1121 vdd.n1120 185
R18705 vdd.n1123 vdd.n1122 185
R18706 vdd.n1125 vdd.n1124 185
R18707 vdd.n1127 vdd.n1126 185
R18708 vdd.n1129 vdd.n1128 185
R18709 vdd.n1131 vdd.n1130 185
R18710 vdd.n1133 vdd.n1132 185
R18711 vdd.n1135 vdd.n1134 185
R18712 vdd.n1137 vdd.n1136 185
R18713 vdd.n1139 vdd.n1138 185
R18714 vdd.n1141 vdd.n1140 185
R18715 vdd.n1343 vdd.n1142 185
R18716 vdd.n1342 vdd.n1341 185
R18717 vdd.n1340 vdd.n1339 185
R18718 vdd.n1338 vdd.n1337 185
R18719 vdd.n1336 vdd.n1335 185
R18720 vdd.n1334 vdd.n1333 185
R18721 vdd.n1332 vdd.n1331 185
R18722 vdd.n1330 vdd.n1329 185
R18723 vdd.n1328 vdd.n1327 185
R18724 vdd.n1326 vdd.n1325 185
R18725 vdd.n1324 vdd.n1323 185
R18726 vdd.n1322 vdd.n1321 185
R18727 vdd.n1320 vdd.n1319 185
R18728 vdd.n1318 vdd.n1317 185
R18729 vdd.n1316 vdd.n1315 185
R18730 vdd.n1314 vdd.n1313 185
R18731 vdd.n1312 vdd.n1311 185
R18732 vdd.n1310 vdd.n1003 185
R18733 vdd.n2218 vdd.n1003 185
R18734 vdd.n303 vdd.n302 171.744
R18735 vdd.n302 vdd.n301 171.744
R18736 vdd.n301 vdd.n270 171.744
R18737 vdd.n294 vdd.n270 171.744
R18738 vdd.n294 vdd.n293 171.744
R18739 vdd.n293 vdd.n275 171.744
R18740 vdd.n286 vdd.n275 171.744
R18741 vdd.n286 vdd.n285 171.744
R18742 vdd.n285 vdd.n279 171.744
R18743 vdd.n252 vdd.n251 171.744
R18744 vdd.n251 vdd.n250 171.744
R18745 vdd.n250 vdd.n219 171.744
R18746 vdd.n243 vdd.n219 171.744
R18747 vdd.n243 vdd.n242 171.744
R18748 vdd.n242 vdd.n224 171.744
R18749 vdd.n235 vdd.n224 171.744
R18750 vdd.n235 vdd.n234 171.744
R18751 vdd.n234 vdd.n228 171.744
R18752 vdd.n209 vdd.n208 171.744
R18753 vdd.n208 vdd.n207 171.744
R18754 vdd.n207 vdd.n176 171.744
R18755 vdd.n200 vdd.n176 171.744
R18756 vdd.n200 vdd.n199 171.744
R18757 vdd.n199 vdd.n181 171.744
R18758 vdd.n192 vdd.n181 171.744
R18759 vdd.n192 vdd.n191 171.744
R18760 vdd.n191 vdd.n185 171.744
R18761 vdd.n158 vdd.n157 171.744
R18762 vdd.n157 vdd.n156 171.744
R18763 vdd.n156 vdd.n125 171.744
R18764 vdd.n149 vdd.n125 171.744
R18765 vdd.n149 vdd.n148 171.744
R18766 vdd.n148 vdd.n130 171.744
R18767 vdd.n141 vdd.n130 171.744
R18768 vdd.n141 vdd.n140 171.744
R18769 vdd.n140 vdd.n134 171.744
R18770 vdd.n116 vdd.n115 171.744
R18771 vdd.n115 vdd.n114 171.744
R18772 vdd.n114 vdd.n83 171.744
R18773 vdd.n107 vdd.n83 171.744
R18774 vdd.n107 vdd.n106 171.744
R18775 vdd.n106 vdd.n88 171.744
R18776 vdd.n99 vdd.n88 171.744
R18777 vdd.n99 vdd.n98 171.744
R18778 vdd.n98 vdd.n92 171.744
R18779 vdd.n65 vdd.n64 171.744
R18780 vdd.n64 vdd.n63 171.744
R18781 vdd.n63 vdd.n32 171.744
R18782 vdd.n56 vdd.n32 171.744
R18783 vdd.n56 vdd.n55 171.744
R18784 vdd.n55 vdd.n37 171.744
R18785 vdd.n48 vdd.n37 171.744
R18786 vdd.n48 vdd.n47 171.744
R18787 vdd.n47 vdd.n41 171.744
R18788 vdd.n1953 vdd.n1952 171.744
R18789 vdd.n1952 vdd.n1951 171.744
R18790 vdd.n1951 vdd.n1920 171.744
R18791 vdd.n1944 vdd.n1920 171.744
R18792 vdd.n1944 vdd.n1943 171.744
R18793 vdd.n1943 vdd.n1925 171.744
R18794 vdd.n1936 vdd.n1925 171.744
R18795 vdd.n1936 vdd.n1935 171.744
R18796 vdd.n1935 vdd.n1929 171.744
R18797 vdd.n2004 vdd.n2003 171.744
R18798 vdd.n2003 vdd.n2002 171.744
R18799 vdd.n2002 vdd.n1971 171.744
R18800 vdd.n1995 vdd.n1971 171.744
R18801 vdd.n1995 vdd.n1994 171.744
R18802 vdd.n1994 vdd.n1976 171.744
R18803 vdd.n1987 vdd.n1976 171.744
R18804 vdd.n1987 vdd.n1986 171.744
R18805 vdd.n1986 vdd.n1980 171.744
R18806 vdd.n1859 vdd.n1858 171.744
R18807 vdd.n1858 vdd.n1857 171.744
R18808 vdd.n1857 vdd.n1826 171.744
R18809 vdd.n1850 vdd.n1826 171.744
R18810 vdd.n1850 vdd.n1849 171.744
R18811 vdd.n1849 vdd.n1831 171.744
R18812 vdd.n1842 vdd.n1831 171.744
R18813 vdd.n1842 vdd.n1841 171.744
R18814 vdd.n1841 vdd.n1835 171.744
R18815 vdd.n1910 vdd.n1909 171.744
R18816 vdd.n1909 vdd.n1908 171.744
R18817 vdd.n1908 vdd.n1877 171.744
R18818 vdd.n1901 vdd.n1877 171.744
R18819 vdd.n1901 vdd.n1900 171.744
R18820 vdd.n1900 vdd.n1882 171.744
R18821 vdd.n1893 vdd.n1882 171.744
R18822 vdd.n1893 vdd.n1892 171.744
R18823 vdd.n1892 vdd.n1886 171.744
R18824 vdd.n1766 vdd.n1765 171.744
R18825 vdd.n1765 vdd.n1764 171.744
R18826 vdd.n1764 vdd.n1733 171.744
R18827 vdd.n1757 vdd.n1733 171.744
R18828 vdd.n1757 vdd.n1756 171.744
R18829 vdd.n1756 vdd.n1738 171.744
R18830 vdd.n1749 vdd.n1738 171.744
R18831 vdd.n1749 vdd.n1748 171.744
R18832 vdd.n1748 vdd.n1742 171.744
R18833 vdd.n1817 vdd.n1816 171.744
R18834 vdd.n1816 vdd.n1815 171.744
R18835 vdd.n1815 vdd.n1784 171.744
R18836 vdd.n1808 vdd.n1784 171.744
R18837 vdd.n1808 vdd.n1807 171.744
R18838 vdd.n1807 vdd.n1789 171.744
R18839 vdd.n1800 vdd.n1789 171.744
R18840 vdd.n1800 vdd.n1799 171.744
R18841 vdd.n1799 vdd.n1793 171.744
R18842 vdd.n3402 vdd.n356 146.341
R18843 vdd.n3400 vdd.n3399 146.341
R18844 vdd.n3397 vdd.n360 146.341
R18845 vdd.n3393 vdd.n3392 146.341
R18846 vdd.n3390 vdd.n368 146.341
R18847 vdd.n3386 vdd.n3385 146.341
R18848 vdd.n3383 vdd.n375 146.341
R18849 vdd.n3379 vdd.n3378 146.341
R18850 vdd.n3376 vdd.n382 146.341
R18851 vdd.n393 vdd.n390 146.341
R18852 vdd.n3368 vdd.n3367 146.341
R18853 vdd.n3365 vdd.n395 146.341
R18854 vdd.n3361 vdd.n3360 146.341
R18855 vdd.n3358 vdd.n401 146.341
R18856 vdd.n3354 vdd.n3353 146.341
R18857 vdd.n3351 vdd.n408 146.341
R18858 vdd.n3347 vdd.n3346 146.341
R18859 vdd.n3344 vdd.n415 146.341
R18860 vdd.n3340 vdd.n3339 146.341
R18861 vdd.n3337 vdd.n422 146.341
R18862 vdd.n433 vdd.n430 146.341
R18863 vdd.n3329 vdd.n3328 146.341
R18864 vdd.n3326 vdd.n435 146.341
R18865 vdd.n3322 vdd.n3321 146.341
R18866 vdd.n3319 vdd.n441 146.341
R18867 vdd.n3315 vdd.n3314 146.341
R18868 vdd.n3312 vdd.n448 146.341
R18869 vdd.n3308 vdd.n3307 146.341
R18870 vdd.n3305 vdd.n455 146.341
R18871 vdd.n3301 vdd.n3300 146.341
R18872 vdd.n3298 vdd.n462 146.341
R18873 vdd.n3213 vdd.n512 146.341
R18874 vdd.n3219 vdd.n512 146.341
R18875 vdd.n3219 vdd.n504 146.341
R18876 vdd.n3229 vdd.n504 146.341
R18877 vdd.n3229 vdd.n500 146.341
R18878 vdd.n3235 vdd.n500 146.341
R18879 vdd.n3235 vdd.n491 146.341
R18880 vdd.n3245 vdd.n491 146.341
R18881 vdd.n3245 vdd.n487 146.341
R18882 vdd.n3251 vdd.n487 146.341
R18883 vdd.n3251 vdd.n479 146.341
R18884 vdd.n3262 vdd.n479 146.341
R18885 vdd.n3262 vdd.n480 146.341
R18886 vdd.n480 vdd.n316 146.341
R18887 vdd.n317 vdd.n316 146.341
R18888 vdd.n318 vdd.n317 146.341
R18889 vdd.n473 vdd.n318 146.341
R18890 vdd.n473 vdd.n326 146.341
R18891 vdd.n327 vdd.n326 146.341
R18892 vdd.n328 vdd.n327 146.341
R18893 vdd.n470 vdd.n328 146.341
R18894 vdd.n470 vdd.n337 146.341
R18895 vdd.n338 vdd.n337 146.341
R18896 vdd.n339 vdd.n338 146.341
R18897 vdd.n467 vdd.n339 146.341
R18898 vdd.n467 vdd.n348 146.341
R18899 vdd.n349 vdd.n348 146.341
R18900 vdd.n350 vdd.n349 146.341
R18901 vdd.n3205 vdd.n3203 146.341
R18902 vdd.n3203 vdd.n3202 146.341
R18903 vdd.n3199 vdd.n3198 146.341
R18904 vdd.n3195 vdd.n3194 146.341
R18905 vdd.n3192 vdd.n526 146.341
R18906 vdd.n3188 vdd.n3186 146.341
R18907 vdd.n3184 vdd.n532 146.341
R18908 vdd.n3180 vdd.n3178 146.341
R18909 vdd.n3176 vdd.n538 146.341
R18910 vdd.n3172 vdd.n3170 146.341
R18911 vdd.n3168 vdd.n546 146.341
R18912 vdd.n3164 vdd.n3162 146.341
R18913 vdd.n3160 vdd.n552 146.341
R18914 vdd.n3156 vdd.n3154 146.341
R18915 vdd.n3152 vdd.n558 146.341
R18916 vdd.n3148 vdd.n3146 146.341
R18917 vdd.n3144 vdd.n564 146.341
R18918 vdd.n3140 vdd.n3138 146.341
R18919 vdd.n3136 vdd.n570 146.341
R18920 vdd.n3132 vdd.n3130 146.341
R18921 vdd.n3128 vdd.n576 146.341
R18922 vdd.n3121 vdd.n585 146.341
R18923 vdd.n3119 vdd.n3118 146.341
R18924 vdd.n3115 vdd.n3114 146.341
R18925 vdd.n3112 vdd.n590 146.341
R18926 vdd.n3108 vdd.n3106 146.341
R18927 vdd.n3104 vdd.n596 146.341
R18928 vdd.n3100 vdd.n3098 146.341
R18929 vdd.n3096 vdd.n602 146.341
R18930 vdd.n3092 vdd.n3090 146.341
R18931 vdd.n3087 vdd.n3086 146.341
R18932 vdd.n3083 vdd.n515 146.341
R18933 vdd.n3211 vdd.n510 146.341
R18934 vdd.n3221 vdd.n510 146.341
R18935 vdd.n3221 vdd.n506 146.341
R18936 vdd.n3227 vdd.n506 146.341
R18937 vdd.n3227 vdd.n498 146.341
R18938 vdd.n3237 vdd.n498 146.341
R18939 vdd.n3237 vdd.n494 146.341
R18940 vdd.n3243 vdd.n494 146.341
R18941 vdd.n3243 vdd.n486 146.341
R18942 vdd.n3254 vdd.n486 146.341
R18943 vdd.n3254 vdd.n482 146.341
R18944 vdd.n3260 vdd.n482 146.341
R18945 vdd.n3260 vdd.n314 146.341
R18946 vdd.n3437 vdd.n314 146.341
R18947 vdd.n3437 vdd.n315 146.341
R18948 vdd.n3433 vdd.n315 146.341
R18949 vdd.n3433 vdd.n319 146.341
R18950 vdd.n3429 vdd.n319 146.341
R18951 vdd.n3429 vdd.n324 146.341
R18952 vdd.n3425 vdd.n324 146.341
R18953 vdd.n3425 vdd.n330 146.341
R18954 vdd.n3421 vdd.n330 146.341
R18955 vdd.n3421 vdd.n336 146.341
R18956 vdd.n3417 vdd.n336 146.341
R18957 vdd.n3417 vdd.n341 146.341
R18958 vdd.n3413 vdd.n341 146.341
R18959 vdd.n3413 vdd.n347 146.341
R18960 vdd.n3409 vdd.n347 146.341
R18961 vdd.n2183 vdd.n2182 146.341
R18962 vdd.n2180 vdd.n2177 146.341
R18963 vdd.n2175 vdd.n1013 146.341
R18964 vdd.n2171 vdd.n2170 146.341
R18965 vdd.n2168 vdd.n1017 146.341
R18966 vdd.n2164 vdd.n2163 146.341
R18967 vdd.n2161 vdd.n1024 146.341
R18968 vdd.n2157 vdd.n2156 146.341
R18969 vdd.n2154 vdd.n1031 146.341
R18970 vdd.n1042 vdd.n1039 146.341
R18971 vdd.n2146 vdd.n2145 146.341
R18972 vdd.n2143 vdd.n1044 146.341
R18973 vdd.n2139 vdd.n2138 146.341
R18974 vdd.n2136 vdd.n1050 146.341
R18975 vdd.n2132 vdd.n2131 146.341
R18976 vdd.n2129 vdd.n1057 146.341
R18977 vdd.n2125 vdd.n2124 146.341
R18978 vdd.n2122 vdd.n1064 146.341
R18979 vdd.n2118 vdd.n2117 146.341
R18980 vdd.n2115 vdd.n1071 146.341
R18981 vdd.n1082 vdd.n1079 146.341
R18982 vdd.n2107 vdd.n2106 146.341
R18983 vdd.n2104 vdd.n1084 146.341
R18984 vdd.n2100 vdd.n2099 146.341
R18985 vdd.n2097 vdd.n1090 146.341
R18986 vdd.n2093 vdd.n2092 146.341
R18987 vdd.n2090 vdd.n1097 146.341
R18988 vdd.n2086 vdd.n2085 146.341
R18989 vdd.n2083 vdd.n1104 146.341
R18990 vdd.n1350 vdd.n1348 146.341
R18991 vdd.n1353 vdd.n1352 146.341
R18992 vdd.n1671 vdd.n1433 146.341
R18993 vdd.n1677 vdd.n1433 146.341
R18994 vdd.n1677 vdd.n1426 146.341
R18995 vdd.n1687 vdd.n1426 146.341
R18996 vdd.n1687 vdd.n1422 146.341
R18997 vdd.n1693 vdd.n1422 146.341
R18998 vdd.n1693 vdd.n1413 146.341
R18999 vdd.n1703 vdd.n1413 146.341
R19000 vdd.n1703 vdd.n1409 146.341
R19001 vdd.n1709 vdd.n1409 146.341
R19002 vdd.n1709 vdd.n1402 146.341
R19003 vdd.n1720 vdd.n1402 146.341
R19004 vdd.n1720 vdd.n1398 146.341
R19005 vdd.n1726 vdd.n1398 146.341
R19006 vdd.n1726 vdd.n1391 146.341
R19007 vdd.n2018 vdd.n1391 146.341
R19008 vdd.n2018 vdd.n1387 146.341
R19009 vdd.n2024 vdd.n1387 146.341
R19010 vdd.n2024 vdd.n1379 146.341
R19011 vdd.n2035 vdd.n1379 146.341
R19012 vdd.n2035 vdd.n1375 146.341
R19013 vdd.n2041 vdd.n1375 146.341
R19014 vdd.n2041 vdd.n1369 146.341
R19015 vdd.n2052 vdd.n1369 146.341
R19016 vdd.n2052 vdd.n1364 146.341
R19017 vdd.n2060 vdd.n1364 146.341
R19018 vdd.n2060 vdd.n1355 146.341
R19019 vdd.n2071 vdd.n1355 146.341
R19020 vdd.n1443 vdd.n1442 146.341
R19021 vdd.n1446 vdd.n1443 146.341
R19022 vdd.n1449 vdd.n1448 146.341
R19023 vdd.n1454 vdd.n1451 146.341
R19024 vdd.n1457 vdd.n1456 146.341
R19025 vdd.n1462 vdd.n1459 146.341
R19026 vdd.n1465 vdd.n1464 146.341
R19027 vdd.n1470 vdd.n1467 146.341
R19028 vdd.n1473 vdd.n1472 146.341
R19029 vdd.n1480 vdd.n1475 146.341
R19030 vdd.n1483 vdd.n1482 146.341
R19031 vdd.n1488 vdd.n1485 146.341
R19032 vdd.n1491 vdd.n1490 146.341
R19033 vdd.n1496 vdd.n1493 146.341
R19034 vdd.n1499 vdd.n1498 146.341
R19035 vdd.n1504 vdd.n1501 146.341
R19036 vdd.n1507 vdd.n1506 146.341
R19037 vdd.n1512 vdd.n1509 146.341
R19038 vdd.n1515 vdd.n1514 146.341
R19039 vdd.n1520 vdd.n1517 146.341
R19040 vdd.n1601 vdd.n1522 146.341
R19041 vdd.n1599 vdd.n1598 146.341
R19042 vdd.n1529 vdd.n1528 146.341
R19043 vdd.n1532 vdd.n1531 146.341
R19044 vdd.n1537 vdd.n1536 146.341
R19045 vdd.n1540 vdd.n1539 146.341
R19046 vdd.n1545 vdd.n1544 146.341
R19047 vdd.n1548 vdd.n1547 146.341
R19048 vdd.n1553 vdd.n1552 146.341
R19049 vdd.n1556 vdd.n1555 146.341
R19050 vdd.n1561 vdd.n1560 146.341
R19051 vdd.n1563 vdd.n1436 146.341
R19052 vdd.n1669 vdd.n1432 146.341
R19053 vdd.n1679 vdd.n1432 146.341
R19054 vdd.n1679 vdd.n1428 146.341
R19055 vdd.n1685 vdd.n1428 146.341
R19056 vdd.n1685 vdd.n1420 146.341
R19057 vdd.n1695 vdd.n1420 146.341
R19058 vdd.n1695 vdd.n1416 146.341
R19059 vdd.n1701 vdd.n1416 146.341
R19060 vdd.n1701 vdd.n1408 146.341
R19061 vdd.n1712 vdd.n1408 146.341
R19062 vdd.n1712 vdd.n1404 146.341
R19063 vdd.n1718 vdd.n1404 146.341
R19064 vdd.n1718 vdd.n1397 146.341
R19065 vdd.n1728 vdd.n1397 146.341
R19066 vdd.n1728 vdd.n1393 146.341
R19067 vdd.n2016 vdd.n1393 146.341
R19068 vdd.n2016 vdd.n1385 146.341
R19069 vdd.n2027 vdd.n1385 146.341
R19070 vdd.n2027 vdd.n1381 146.341
R19071 vdd.n2033 vdd.n1381 146.341
R19072 vdd.n2033 vdd.n1374 146.341
R19073 vdd.n2044 vdd.n1374 146.341
R19074 vdd.n2044 vdd.n1370 146.341
R19075 vdd.n2050 vdd.n1370 146.341
R19076 vdd.n2050 vdd.n1362 146.341
R19077 vdd.n2063 vdd.n1362 146.341
R19078 vdd.n2063 vdd.n1357 146.341
R19079 vdd.n2069 vdd.n1357 146.341
R19080 vdd.n1143 vdd.t7 127.284
R19081 vdd.n838 vdd.t51 127.284
R19082 vdd.n1147 vdd.t48 127.284
R19083 vdd.n829 vdd.t74 127.284
R19084 vdd.n724 vdd.t28 127.284
R19085 vdd.n724 vdd.t29 127.284
R19086 vdd.n2535 vdd.t69 127.284
R19087 vdd.n661 vdd.t16 127.284
R19088 vdd.n2532 vdd.t59 127.284
R19089 vdd.n625 vdd.t2 127.284
R19090 vdd.n899 vdd.t65 127.284
R19091 vdd.n899 vdd.t66 127.284
R19092 vdd.n22 vdd.n20 117.314
R19093 vdd.n17 vdd.n15 117.314
R19094 vdd.n27 vdd.n26 116.927
R19095 vdd.n24 vdd.n23 116.927
R19096 vdd.n22 vdd.n21 116.927
R19097 vdd.n17 vdd.n16 116.927
R19098 vdd.n19 vdd.n18 116.927
R19099 vdd.n27 vdd.n25 116.927
R19100 vdd.n1144 vdd.t6 111.188
R19101 vdd.n839 vdd.t52 111.188
R19102 vdd.n1148 vdd.t47 111.188
R19103 vdd.n830 vdd.t75 111.188
R19104 vdd.n2536 vdd.t68 111.188
R19105 vdd.n662 vdd.t17 111.188
R19106 vdd.n2533 vdd.t58 111.188
R19107 vdd.n626 vdd.t3 111.188
R19108 vdd.n2806 vdd.n788 99.5127
R19109 vdd.n2806 vdd.n779 99.5127
R19110 vdd.n2814 vdd.n779 99.5127
R19111 vdd.n2814 vdd.n777 99.5127
R19112 vdd.n2818 vdd.n777 99.5127
R19113 vdd.n2818 vdd.n767 99.5127
R19114 vdd.n2826 vdd.n767 99.5127
R19115 vdd.n2826 vdd.n765 99.5127
R19116 vdd.n2830 vdd.n765 99.5127
R19117 vdd.n2830 vdd.n756 99.5127
R19118 vdd.n2838 vdd.n756 99.5127
R19119 vdd.n2838 vdd.n754 99.5127
R19120 vdd.n2842 vdd.n754 99.5127
R19121 vdd.n2842 vdd.n745 99.5127
R19122 vdd.n2850 vdd.n745 99.5127
R19123 vdd.n2850 vdd.n743 99.5127
R19124 vdd.n2854 vdd.n743 99.5127
R19125 vdd.n2854 vdd.n732 99.5127
R19126 vdd.n2863 vdd.n732 99.5127
R19127 vdd.n2863 vdd.n730 99.5127
R19128 vdd.n2867 vdd.n730 99.5127
R19129 vdd.n2867 vdd.n720 99.5127
R19130 vdd.n2875 vdd.n720 99.5127
R19131 vdd.n2875 vdd.n718 99.5127
R19132 vdd.n2879 vdd.n718 99.5127
R19133 vdd.n2879 vdd.n708 99.5127
R19134 vdd.n2887 vdd.n708 99.5127
R19135 vdd.n2887 vdd.n706 99.5127
R19136 vdd.n2891 vdd.n706 99.5127
R19137 vdd.n2891 vdd.n695 99.5127
R19138 vdd.n2899 vdd.n695 99.5127
R19139 vdd.n2899 vdd.n693 99.5127
R19140 vdd.n2903 vdd.n693 99.5127
R19141 vdd.n2903 vdd.n684 99.5127
R19142 vdd.n2911 vdd.n684 99.5127
R19143 vdd.n2911 vdd.n682 99.5127
R19144 vdd.n2915 vdd.n682 99.5127
R19145 vdd.n2915 vdd.n670 99.5127
R19146 vdd.n2968 vdd.n670 99.5127
R19147 vdd.n2968 vdd.n668 99.5127
R19148 vdd.n2972 vdd.n668 99.5127
R19149 vdd.n2972 vdd.n634 99.5127
R19150 vdd.n3042 vdd.n634 99.5127
R19151 vdd.n3038 vdd.n635 99.5127
R19152 vdd.n3036 vdd.n3035 99.5127
R19153 vdd.n3033 vdd.n639 99.5127
R19154 vdd.n3029 vdd.n3028 99.5127
R19155 vdd.n3026 vdd.n642 99.5127
R19156 vdd.n3022 vdd.n3021 99.5127
R19157 vdd.n3019 vdd.n645 99.5127
R19158 vdd.n3015 vdd.n3014 99.5127
R19159 vdd.n3012 vdd.n648 99.5127
R19160 vdd.n3007 vdd.n3006 99.5127
R19161 vdd.n3004 vdd.n651 99.5127
R19162 vdd.n3000 vdd.n2999 99.5127
R19163 vdd.n2997 vdd.n654 99.5127
R19164 vdd.n2993 vdd.n2992 99.5127
R19165 vdd.n2990 vdd.n657 99.5127
R19166 vdd.n2986 vdd.n2985 99.5127
R19167 vdd.n2983 vdd.n660 99.5127
R19168 vdd.n2733 vdd.n786 99.5127
R19169 vdd.n2729 vdd.n786 99.5127
R19170 vdd.n2729 vdd.n780 99.5127
R19171 vdd.n2611 vdd.n780 99.5127
R19172 vdd.n2611 vdd.n775 99.5127
R19173 vdd.n2614 vdd.n775 99.5127
R19174 vdd.n2614 vdd.n769 99.5127
R19175 vdd.n2715 vdd.n769 99.5127
R19176 vdd.n2715 vdd.n763 99.5127
R19177 vdd.n2711 vdd.n763 99.5127
R19178 vdd.n2711 vdd.n757 99.5127
R19179 vdd.n2658 vdd.n757 99.5127
R19180 vdd.n2658 vdd.n751 99.5127
R19181 vdd.n2655 vdd.n751 99.5127
R19182 vdd.n2655 vdd.n746 99.5127
R19183 vdd.n2652 vdd.n746 99.5127
R19184 vdd.n2652 vdd.n741 99.5127
R19185 vdd.n2649 vdd.n741 99.5127
R19186 vdd.n2649 vdd.n734 99.5127
R19187 vdd.n2646 vdd.n734 99.5127
R19188 vdd.n2646 vdd.n727 99.5127
R19189 vdd.n2643 vdd.n727 99.5127
R19190 vdd.n2643 vdd.n721 99.5127
R19191 vdd.n2640 vdd.n721 99.5127
R19192 vdd.n2640 vdd.n716 99.5127
R19193 vdd.n2637 vdd.n716 99.5127
R19194 vdd.n2637 vdd.n710 99.5127
R19195 vdd.n2634 vdd.n710 99.5127
R19196 vdd.n2634 vdd.n703 99.5127
R19197 vdd.n2631 vdd.n703 99.5127
R19198 vdd.n2631 vdd.n696 99.5127
R19199 vdd.n2628 vdd.n696 99.5127
R19200 vdd.n2628 vdd.n690 99.5127
R19201 vdd.n2625 vdd.n690 99.5127
R19202 vdd.n2625 vdd.n685 99.5127
R19203 vdd.n2622 vdd.n685 99.5127
R19204 vdd.n2622 vdd.n680 99.5127
R19205 vdd.n2619 vdd.n680 99.5127
R19206 vdd.n2619 vdd.n672 99.5127
R19207 vdd.n672 vdd.n665 99.5127
R19208 vdd.n2974 vdd.n665 99.5127
R19209 vdd.n2975 vdd.n2974 99.5127
R19210 vdd.n2975 vdd.n632 99.5127
R19211 vdd.n2799 vdd.n790 99.5127
R19212 vdd.n2799 vdd.n2531 99.5127
R19213 vdd.n2795 vdd.n2794 99.5127
R19214 vdd.n2791 vdd.n2790 99.5127
R19215 vdd.n2787 vdd.n2786 99.5127
R19216 vdd.n2783 vdd.n2782 99.5127
R19217 vdd.n2779 vdd.n2778 99.5127
R19218 vdd.n2775 vdd.n2774 99.5127
R19219 vdd.n2771 vdd.n2770 99.5127
R19220 vdd.n2767 vdd.n2766 99.5127
R19221 vdd.n2763 vdd.n2762 99.5127
R19222 vdd.n2759 vdd.n2758 99.5127
R19223 vdd.n2755 vdd.n2754 99.5127
R19224 vdd.n2751 vdd.n2750 99.5127
R19225 vdd.n2747 vdd.n2746 99.5127
R19226 vdd.n2743 vdd.n2742 99.5127
R19227 vdd.n2738 vdd.n2737 99.5127
R19228 vdd.n2495 vdd.n827 99.5127
R19229 vdd.n2491 vdd.n2490 99.5127
R19230 vdd.n2487 vdd.n2486 99.5127
R19231 vdd.n2483 vdd.n2482 99.5127
R19232 vdd.n2479 vdd.n2478 99.5127
R19233 vdd.n2475 vdd.n2474 99.5127
R19234 vdd.n2471 vdd.n2470 99.5127
R19235 vdd.n2467 vdd.n2466 99.5127
R19236 vdd.n2463 vdd.n2462 99.5127
R19237 vdd.n2459 vdd.n2458 99.5127
R19238 vdd.n2455 vdd.n2454 99.5127
R19239 vdd.n2451 vdd.n2450 99.5127
R19240 vdd.n2447 vdd.n2446 99.5127
R19241 vdd.n2443 vdd.n2442 99.5127
R19242 vdd.n2439 vdd.n2438 99.5127
R19243 vdd.n2435 vdd.n2434 99.5127
R19244 vdd.n2430 vdd.n2429 99.5127
R19245 vdd.n1183 vdd.n963 99.5127
R19246 vdd.n1186 vdd.n963 99.5127
R19247 vdd.n1186 vdd.n957 99.5127
R19248 vdd.n1189 vdd.n957 99.5127
R19249 vdd.n1189 vdd.n952 99.5127
R19250 vdd.n1192 vdd.n952 99.5127
R19251 vdd.n1192 vdd.n945 99.5127
R19252 vdd.n1195 vdd.n945 99.5127
R19253 vdd.n1195 vdd.n938 99.5127
R19254 vdd.n1198 vdd.n938 99.5127
R19255 vdd.n1198 vdd.n932 99.5127
R19256 vdd.n1201 vdd.n932 99.5127
R19257 vdd.n1201 vdd.n927 99.5127
R19258 vdd.n1204 vdd.n927 99.5127
R19259 vdd.n1204 vdd.n922 99.5127
R19260 vdd.n1207 vdd.n922 99.5127
R19261 vdd.n1207 vdd.n916 99.5127
R19262 vdd.n1210 vdd.n916 99.5127
R19263 vdd.n1210 vdd.n909 99.5127
R19264 vdd.n1213 vdd.n909 99.5127
R19265 vdd.n1213 vdd.n902 99.5127
R19266 vdd.n1216 vdd.n902 99.5127
R19267 vdd.n1216 vdd.n896 99.5127
R19268 vdd.n1219 vdd.n896 99.5127
R19269 vdd.n1219 vdd.n891 99.5127
R19270 vdd.n1222 vdd.n891 99.5127
R19271 vdd.n1222 vdd.n885 99.5127
R19272 vdd.n1264 vdd.n885 99.5127
R19273 vdd.n1264 vdd.n878 99.5127
R19274 vdd.n1260 vdd.n878 99.5127
R19275 vdd.n1260 vdd.n872 99.5127
R19276 vdd.n1257 vdd.n872 99.5127
R19277 vdd.n1257 vdd.n867 99.5127
R19278 vdd.n1254 vdd.n867 99.5127
R19279 vdd.n1254 vdd.n862 99.5127
R19280 vdd.n1234 vdd.n862 99.5127
R19281 vdd.n1234 vdd.n857 99.5127
R19282 vdd.n1231 vdd.n857 99.5127
R19283 vdd.n1231 vdd.n850 99.5127
R19284 vdd.n1228 vdd.n850 99.5127
R19285 vdd.n1228 vdd.n843 99.5127
R19286 vdd.n843 vdd.n832 99.5127
R19287 vdd.n2425 vdd.n832 99.5127
R19288 vdd.n2217 vdd.n968 99.5127
R19289 vdd.n2217 vdd.n1004 99.5127
R19290 vdd.n2213 vdd.n2212 99.5127
R19291 vdd.n2209 vdd.n2208 99.5127
R19292 vdd.n2205 vdd.n2204 99.5127
R19293 vdd.n2201 vdd.n2200 99.5127
R19294 vdd.n2197 vdd.n2196 99.5127
R19295 vdd.n2193 vdd.n2192 99.5127
R19296 vdd.n2189 vdd.n2188 99.5127
R19297 vdd.n1150 vdd.n1149 99.5127
R19298 vdd.n1154 vdd.n1153 99.5127
R19299 vdd.n1158 vdd.n1157 99.5127
R19300 vdd.n1162 vdd.n1161 99.5127
R19301 vdd.n1166 vdd.n1165 99.5127
R19302 vdd.n1170 vdd.n1169 99.5127
R19303 vdd.n1174 vdd.n1173 99.5127
R19304 vdd.n1179 vdd.n1178 99.5127
R19305 vdd.n2224 vdd.n966 99.5127
R19306 vdd.n2224 vdd.n956 99.5127
R19307 vdd.n2232 vdd.n956 99.5127
R19308 vdd.n2232 vdd.n954 99.5127
R19309 vdd.n2236 vdd.n954 99.5127
R19310 vdd.n2236 vdd.n943 99.5127
R19311 vdd.n2244 vdd.n943 99.5127
R19312 vdd.n2244 vdd.n941 99.5127
R19313 vdd.n2248 vdd.n941 99.5127
R19314 vdd.n2248 vdd.n931 99.5127
R19315 vdd.n2256 vdd.n931 99.5127
R19316 vdd.n2256 vdd.n929 99.5127
R19317 vdd.n2260 vdd.n929 99.5127
R19318 vdd.n2260 vdd.n920 99.5127
R19319 vdd.n2268 vdd.n920 99.5127
R19320 vdd.n2268 vdd.n918 99.5127
R19321 vdd.n2272 vdd.n918 99.5127
R19322 vdd.n2272 vdd.n907 99.5127
R19323 vdd.n2280 vdd.n907 99.5127
R19324 vdd.n2280 vdd.n905 99.5127
R19325 vdd.n2284 vdd.n905 99.5127
R19326 vdd.n2284 vdd.n895 99.5127
R19327 vdd.n2293 vdd.n895 99.5127
R19328 vdd.n2293 vdd.n893 99.5127
R19329 vdd.n2297 vdd.n893 99.5127
R19330 vdd.n2297 vdd.n883 99.5127
R19331 vdd.n2305 vdd.n883 99.5127
R19332 vdd.n2305 vdd.n881 99.5127
R19333 vdd.n2309 vdd.n881 99.5127
R19334 vdd.n2309 vdd.n871 99.5127
R19335 vdd.n2317 vdd.n871 99.5127
R19336 vdd.n2317 vdd.n869 99.5127
R19337 vdd.n2321 vdd.n869 99.5127
R19338 vdd.n2321 vdd.n861 99.5127
R19339 vdd.n2329 vdd.n861 99.5127
R19340 vdd.n2329 vdd.n859 99.5127
R19341 vdd.n2333 vdd.n859 99.5127
R19342 vdd.n2333 vdd.n848 99.5127
R19343 vdd.n2343 vdd.n848 99.5127
R19344 vdd.n2343 vdd.n845 99.5127
R19345 vdd.n2348 vdd.n845 99.5127
R19346 vdd.n2348 vdd.n846 99.5127
R19347 vdd.n846 vdd.n826 99.5127
R19348 vdd.n2958 vdd.n2957 99.5127
R19349 vdd.n2955 vdd.n2921 99.5127
R19350 vdd.n2951 vdd.n2950 99.5127
R19351 vdd.n2948 vdd.n2924 99.5127
R19352 vdd.n2944 vdd.n2943 99.5127
R19353 vdd.n2941 vdd.n2927 99.5127
R19354 vdd.n2937 vdd.n2936 99.5127
R19355 vdd.n2934 vdd.n2931 99.5127
R19356 vdd.n3075 vdd.n612 99.5127
R19357 vdd.n3073 vdd.n3072 99.5127
R19358 vdd.n3070 vdd.n615 99.5127
R19359 vdd.n3066 vdd.n3065 99.5127
R19360 vdd.n3063 vdd.n618 99.5127
R19361 vdd.n3059 vdd.n3058 99.5127
R19362 vdd.n3056 vdd.n621 99.5127
R19363 vdd.n3052 vdd.n3051 99.5127
R19364 vdd.n3049 vdd.n624 99.5127
R19365 vdd.n2607 vdd.n787 99.5127
R19366 vdd.n2727 vdd.n787 99.5127
R19367 vdd.n2727 vdd.n781 99.5127
R19368 vdd.n2723 vdd.n781 99.5127
R19369 vdd.n2723 vdd.n776 99.5127
R19370 vdd.n2720 vdd.n776 99.5127
R19371 vdd.n2720 vdd.n770 99.5127
R19372 vdd.n2717 vdd.n770 99.5127
R19373 vdd.n2717 vdd.n764 99.5127
R19374 vdd.n2709 vdd.n764 99.5127
R19375 vdd.n2709 vdd.n758 99.5127
R19376 vdd.n2705 vdd.n758 99.5127
R19377 vdd.n2705 vdd.n752 99.5127
R19378 vdd.n2702 vdd.n752 99.5127
R19379 vdd.n2702 vdd.n747 99.5127
R19380 vdd.n2699 vdd.n747 99.5127
R19381 vdd.n2699 vdd.n742 99.5127
R19382 vdd.n2696 vdd.n742 99.5127
R19383 vdd.n2696 vdd.n735 99.5127
R19384 vdd.n2693 vdd.n735 99.5127
R19385 vdd.n2693 vdd.n728 99.5127
R19386 vdd.n2690 vdd.n728 99.5127
R19387 vdd.n2690 vdd.n722 99.5127
R19388 vdd.n2687 vdd.n722 99.5127
R19389 vdd.n2687 vdd.n717 99.5127
R19390 vdd.n2684 vdd.n717 99.5127
R19391 vdd.n2684 vdd.n711 99.5127
R19392 vdd.n2681 vdd.n711 99.5127
R19393 vdd.n2681 vdd.n704 99.5127
R19394 vdd.n2678 vdd.n704 99.5127
R19395 vdd.n2678 vdd.n697 99.5127
R19396 vdd.n2675 vdd.n697 99.5127
R19397 vdd.n2675 vdd.n691 99.5127
R19398 vdd.n2672 vdd.n691 99.5127
R19399 vdd.n2672 vdd.n686 99.5127
R19400 vdd.n2669 vdd.n686 99.5127
R19401 vdd.n2669 vdd.n681 99.5127
R19402 vdd.n2666 vdd.n681 99.5127
R19403 vdd.n2666 vdd.n673 99.5127
R19404 vdd.n2663 vdd.n673 99.5127
R19405 vdd.n2663 vdd.n666 99.5127
R19406 vdd.n666 vdd.n630 99.5127
R19407 vdd.n3044 vdd.n630 99.5127
R19408 vdd.n2542 vdd.n2541 99.5127
R19409 vdd.n2546 vdd.n2545 99.5127
R19410 vdd.n2550 vdd.n2549 99.5127
R19411 vdd.n2554 vdd.n2553 99.5127
R19412 vdd.n2558 vdd.n2557 99.5127
R19413 vdd.n2562 vdd.n2561 99.5127
R19414 vdd.n2566 vdd.n2565 99.5127
R19415 vdd.n2570 vdd.n2569 99.5127
R19416 vdd.n2574 vdd.n2573 99.5127
R19417 vdd.n2578 vdd.n2577 99.5127
R19418 vdd.n2582 vdd.n2581 99.5127
R19419 vdd.n2586 vdd.n2585 99.5127
R19420 vdd.n2590 vdd.n2589 99.5127
R19421 vdd.n2594 vdd.n2593 99.5127
R19422 vdd.n2598 vdd.n2597 99.5127
R19423 vdd.n2602 vdd.n2601 99.5127
R19424 vdd.n2604 vdd.n2530 99.5127
R19425 vdd.n2808 vdd.n784 99.5127
R19426 vdd.n2808 vdd.n782 99.5127
R19427 vdd.n2812 vdd.n782 99.5127
R19428 vdd.n2812 vdd.n773 99.5127
R19429 vdd.n2820 vdd.n773 99.5127
R19430 vdd.n2820 vdd.n771 99.5127
R19431 vdd.n2824 vdd.n771 99.5127
R19432 vdd.n2824 vdd.n762 99.5127
R19433 vdd.n2832 vdd.n762 99.5127
R19434 vdd.n2832 vdd.n760 99.5127
R19435 vdd.n2836 vdd.n760 99.5127
R19436 vdd.n2836 vdd.n750 99.5127
R19437 vdd.n2844 vdd.n750 99.5127
R19438 vdd.n2844 vdd.n748 99.5127
R19439 vdd.n2848 vdd.n748 99.5127
R19440 vdd.n2848 vdd.n739 99.5127
R19441 vdd.n2856 vdd.n739 99.5127
R19442 vdd.n2856 vdd.n737 99.5127
R19443 vdd.n2861 vdd.n737 99.5127
R19444 vdd.n2861 vdd.n726 99.5127
R19445 vdd.n2869 vdd.n726 99.5127
R19446 vdd.n2869 vdd.n723 99.5127
R19447 vdd.n2873 vdd.n723 99.5127
R19448 vdd.n2873 vdd.n714 99.5127
R19449 vdd.n2881 vdd.n714 99.5127
R19450 vdd.n2881 vdd.n712 99.5127
R19451 vdd.n2885 vdd.n712 99.5127
R19452 vdd.n2885 vdd.n701 99.5127
R19453 vdd.n2893 vdd.n701 99.5127
R19454 vdd.n2893 vdd.n699 99.5127
R19455 vdd.n2897 vdd.n699 99.5127
R19456 vdd.n2897 vdd.n689 99.5127
R19457 vdd.n2905 vdd.n689 99.5127
R19458 vdd.n2905 vdd.n687 99.5127
R19459 vdd.n2909 vdd.n687 99.5127
R19460 vdd.n2909 vdd.n678 99.5127
R19461 vdd.n2917 vdd.n678 99.5127
R19462 vdd.n2917 vdd.n675 99.5127
R19463 vdd.n2966 vdd.n675 99.5127
R19464 vdd.n2966 vdd.n676 99.5127
R19465 vdd.n676 vdd.n667 99.5127
R19466 vdd.n2961 vdd.n667 99.5127
R19467 vdd.n2961 vdd.n633 99.5127
R19468 vdd.n2419 vdd.n2418 99.5127
R19469 vdd.n2415 vdd.n2414 99.5127
R19470 vdd.n2411 vdd.n2410 99.5127
R19471 vdd.n2407 vdd.n2406 99.5127
R19472 vdd.n2403 vdd.n2402 99.5127
R19473 vdd.n2399 vdd.n2398 99.5127
R19474 vdd.n2395 vdd.n2394 99.5127
R19475 vdd.n2391 vdd.n2390 99.5127
R19476 vdd.n2387 vdd.n2386 99.5127
R19477 vdd.n2383 vdd.n2382 99.5127
R19478 vdd.n2379 vdd.n2378 99.5127
R19479 vdd.n2375 vdd.n2374 99.5127
R19480 vdd.n2371 vdd.n2370 99.5127
R19481 vdd.n2367 vdd.n2366 99.5127
R19482 vdd.n2363 vdd.n2362 99.5127
R19483 vdd.n2359 vdd.n2358 99.5127
R19484 vdd.n2355 vdd.n808 99.5127
R19485 vdd.n1308 vdd.n964 99.5127
R19486 vdd.n1305 vdd.n964 99.5127
R19487 vdd.n1305 vdd.n958 99.5127
R19488 vdd.n1302 vdd.n958 99.5127
R19489 vdd.n1302 vdd.n953 99.5127
R19490 vdd.n1299 vdd.n953 99.5127
R19491 vdd.n1299 vdd.n946 99.5127
R19492 vdd.n1296 vdd.n946 99.5127
R19493 vdd.n1296 vdd.n939 99.5127
R19494 vdd.n1293 vdd.n939 99.5127
R19495 vdd.n1293 vdd.n933 99.5127
R19496 vdd.n1290 vdd.n933 99.5127
R19497 vdd.n1290 vdd.n928 99.5127
R19498 vdd.n1287 vdd.n928 99.5127
R19499 vdd.n1287 vdd.n923 99.5127
R19500 vdd.n1284 vdd.n923 99.5127
R19501 vdd.n1284 vdd.n917 99.5127
R19502 vdd.n1281 vdd.n917 99.5127
R19503 vdd.n1281 vdd.n910 99.5127
R19504 vdd.n1278 vdd.n910 99.5127
R19505 vdd.n1278 vdd.n903 99.5127
R19506 vdd.n1275 vdd.n903 99.5127
R19507 vdd.n1275 vdd.n897 99.5127
R19508 vdd.n1272 vdd.n897 99.5127
R19509 vdd.n1272 vdd.n892 99.5127
R19510 vdd.n1269 vdd.n892 99.5127
R19511 vdd.n1269 vdd.n886 99.5127
R19512 vdd.n1266 vdd.n886 99.5127
R19513 vdd.n1266 vdd.n879 99.5127
R19514 vdd.n1237 vdd.n879 99.5127
R19515 vdd.n1237 vdd.n873 99.5127
R19516 vdd.n1240 vdd.n873 99.5127
R19517 vdd.n1240 vdd.n868 99.5127
R19518 vdd.n1252 vdd.n868 99.5127
R19519 vdd.n1252 vdd.n863 99.5127
R19520 vdd.n1248 vdd.n863 99.5127
R19521 vdd.n1248 vdd.n858 99.5127
R19522 vdd.n1245 vdd.n858 99.5127
R19523 vdd.n1245 vdd.n851 99.5127
R19524 vdd.n851 vdd.n842 99.5127
R19525 vdd.n2350 vdd.n842 99.5127
R19526 vdd.n2351 vdd.n2350 99.5127
R19527 vdd.n2351 vdd.n834 99.5127
R19528 vdd.n1112 vdd.n1111 99.5127
R19529 vdd.n1116 vdd.n1115 99.5127
R19530 vdd.n1120 vdd.n1119 99.5127
R19531 vdd.n1124 vdd.n1123 99.5127
R19532 vdd.n1128 vdd.n1127 99.5127
R19533 vdd.n1132 vdd.n1131 99.5127
R19534 vdd.n1136 vdd.n1135 99.5127
R19535 vdd.n1140 vdd.n1139 99.5127
R19536 vdd.n1341 vdd.n1142 99.5127
R19537 vdd.n1339 vdd.n1338 99.5127
R19538 vdd.n1335 vdd.n1334 99.5127
R19539 vdd.n1331 vdd.n1330 99.5127
R19540 vdd.n1327 vdd.n1326 99.5127
R19541 vdd.n1323 vdd.n1322 99.5127
R19542 vdd.n1319 vdd.n1318 99.5127
R19543 vdd.n1315 vdd.n1314 99.5127
R19544 vdd.n1311 vdd.n1003 99.5127
R19545 vdd.n2226 vdd.n961 99.5127
R19546 vdd.n2226 vdd.n959 99.5127
R19547 vdd.n2230 vdd.n959 99.5127
R19548 vdd.n2230 vdd.n950 99.5127
R19549 vdd.n2238 vdd.n950 99.5127
R19550 vdd.n2238 vdd.n948 99.5127
R19551 vdd.n2242 vdd.n948 99.5127
R19552 vdd.n2242 vdd.n937 99.5127
R19553 vdd.n2250 vdd.n937 99.5127
R19554 vdd.n2250 vdd.n935 99.5127
R19555 vdd.n2254 vdd.n935 99.5127
R19556 vdd.n2254 vdd.n926 99.5127
R19557 vdd.n2262 vdd.n926 99.5127
R19558 vdd.n2262 vdd.n924 99.5127
R19559 vdd.n2266 vdd.n924 99.5127
R19560 vdd.n2266 vdd.n914 99.5127
R19561 vdd.n2274 vdd.n914 99.5127
R19562 vdd.n2274 vdd.n912 99.5127
R19563 vdd.n2278 vdd.n912 99.5127
R19564 vdd.n2278 vdd.n901 99.5127
R19565 vdd.n2286 vdd.n901 99.5127
R19566 vdd.n2286 vdd.n898 99.5127
R19567 vdd.n2291 vdd.n898 99.5127
R19568 vdd.n2291 vdd.n889 99.5127
R19569 vdd.n2299 vdd.n889 99.5127
R19570 vdd.n2299 vdd.n887 99.5127
R19571 vdd.n2303 vdd.n887 99.5127
R19572 vdd.n2303 vdd.n877 99.5127
R19573 vdd.n2311 vdd.n877 99.5127
R19574 vdd.n2311 vdd.n875 99.5127
R19575 vdd.n2315 vdd.n875 99.5127
R19576 vdd.n2315 vdd.n866 99.5127
R19577 vdd.n2323 vdd.n866 99.5127
R19578 vdd.n2323 vdd.n864 99.5127
R19579 vdd.n2327 vdd.n864 99.5127
R19580 vdd.n2327 vdd.n855 99.5127
R19581 vdd.n2335 vdd.n855 99.5127
R19582 vdd.n2335 vdd.n852 99.5127
R19583 vdd.n2341 vdd.n852 99.5127
R19584 vdd.n2341 vdd.n853 99.5127
R19585 vdd.n853 vdd.n844 99.5127
R19586 vdd.n844 vdd.n835 99.5127
R19587 vdd.n2423 vdd.n835 99.5127
R19588 vdd.n9 vdd.n7 98.9633
R19589 vdd.n2 vdd.n0 98.9633
R19590 vdd.n9 vdd.n8 98.6055
R19591 vdd.n11 vdd.n10 98.6055
R19592 vdd.n13 vdd.n12 98.6055
R19593 vdd.n6 vdd.n5 98.6055
R19594 vdd.n4 vdd.n3 98.6055
R19595 vdd.n2 vdd.n1 98.6055
R19596 vdd.t161 vdd.n279 85.8723
R19597 vdd.t240 vdd.n228 85.8723
R19598 vdd.t242 vdd.n185 85.8723
R19599 vdd.t234 vdd.n134 85.8723
R19600 vdd.t184 vdd.n92 85.8723
R19601 vdd.t201 vdd.n41 85.8723
R19602 vdd.t191 vdd.n1929 85.8723
R19603 vdd.t195 vdd.n1980 85.8723
R19604 vdd.t178 vdd.n1835 85.8723
R19605 vdd.t185 vdd.n1886 85.8723
R19606 vdd.t202 vdd.n1742 85.8723
R19607 vdd.t183 vdd.n1793 85.8723
R19608 vdd.n725 vdd.n724 78.546
R19609 vdd.n2289 vdd.n899 78.546
R19610 vdd.n266 vdd.n265 75.1835
R19611 vdd.n264 vdd.n263 75.1835
R19612 vdd.n262 vdd.n261 75.1835
R19613 vdd.n260 vdd.n259 75.1835
R19614 vdd.n258 vdd.n257 75.1835
R19615 vdd.n172 vdd.n171 75.1835
R19616 vdd.n170 vdd.n169 75.1835
R19617 vdd.n168 vdd.n167 75.1835
R19618 vdd.n166 vdd.n165 75.1835
R19619 vdd.n164 vdd.n163 75.1835
R19620 vdd.n79 vdd.n78 75.1835
R19621 vdd.n77 vdd.n76 75.1835
R19622 vdd.n75 vdd.n74 75.1835
R19623 vdd.n73 vdd.n72 75.1835
R19624 vdd.n71 vdd.n70 75.1835
R19625 vdd.n1959 vdd.n1958 75.1835
R19626 vdd.n1961 vdd.n1960 75.1835
R19627 vdd.n1963 vdd.n1962 75.1835
R19628 vdd.n1965 vdd.n1964 75.1835
R19629 vdd.n1967 vdd.n1966 75.1835
R19630 vdd.n1865 vdd.n1864 75.1835
R19631 vdd.n1867 vdd.n1866 75.1835
R19632 vdd.n1869 vdd.n1868 75.1835
R19633 vdd.n1871 vdd.n1870 75.1835
R19634 vdd.n1873 vdd.n1872 75.1835
R19635 vdd.n1772 vdd.n1771 75.1835
R19636 vdd.n1774 vdd.n1773 75.1835
R19637 vdd.n1776 vdd.n1775 75.1835
R19638 vdd.n1778 vdd.n1777 75.1835
R19639 vdd.n1780 vdd.n1779 75.1835
R19640 vdd.n2800 vdd.n2513 72.8958
R19641 vdd.n2800 vdd.n2514 72.8958
R19642 vdd.n2800 vdd.n2515 72.8958
R19643 vdd.n2800 vdd.n2516 72.8958
R19644 vdd.n2800 vdd.n2517 72.8958
R19645 vdd.n2800 vdd.n2518 72.8958
R19646 vdd.n2800 vdd.n2519 72.8958
R19647 vdd.n2800 vdd.n2520 72.8958
R19648 vdd.n2800 vdd.n2521 72.8958
R19649 vdd.n2800 vdd.n2522 72.8958
R19650 vdd.n2800 vdd.n2523 72.8958
R19651 vdd.n2800 vdd.n2524 72.8958
R19652 vdd.n2800 vdd.n2525 72.8958
R19653 vdd.n2800 vdd.n2526 72.8958
R19654 vdd.n2800 vdd.n2527 72.8958
R19655 vdd.n2800 vdd.n2528 72.8958
R19656 vdd.n2800 vdd.n2529 72.8958
R19657 vdd.n629 vdd.n613 72.8958
R19658 vdd.n3050 vdd.n613 72.8958
R19659 vdd.n623 vdd.n613 72.8958
R19660 vdd.n3057 vdd.n613 72.8958
R19661 vdd.n620 vdd.n613 72.8958
R19662 vdd.n3064 vdd.n613 72.8958
R19663 vdd.n617 vdd.n613 72.8958
R19664 vdd.n3071 vdd.n613 72.8958
R19665 vdd.n3074 vdd.n613 72.8958
R19666 vdd.n2930 vdd.n613 72.8958
R19667 vdd.n2935 vdd.n613 72.8958
R19668 vdd.n2929 vdd.n613 72.8958
R19669 vdd.n2942 vdd.n613 72.8958
R19670 vdd.n2926 vdd.n613 72.8958
R19671 vdd.n2949 vdd.n613 72.8958
R19672 vdd.n2923 vdd.n613 72.8958
R19673 vdd.n2956 vdd.n613 72.8958
R19674 vdd.n2219 vdd.n2218 72.8958
R19675 vdd.n2218 vdd.n970 72.8958
R19676 vdd.n2218 vdd.n971 72.8958
R19677 vdd.n2218 vdd.n972 72.8958
R19678 vdd.n2218 vdd.n973 72.8958
R19679 vdd.n2218 vdd.n974 72.8958
R19680 vdd.n2218 vdd.n975 72.8958
R19681 vdd.n2218 vdd.n976 72.8958
R19682 vdd.n2218 vdd.n977 72.8958
R19683 vdd.n2218 vdd.n978 72.8958
R19684 vdd.n2218 vdd.n979 72.8958
R19685 vdd.n2218 vdd.n980 72.8958
R19686 vdd.n2218 vdd.n981 72.8958
R19687 vdd.n2218 vdd.n982 72.8958
R19688 vdd.n2218 vdd.n983 72.8958
R19689 vdd.n2218 vdd.n984 72.8958
R19690 vdd.n2218 vdd.n985 72.8958
R19691 vdd.n2496 vdd.n809 72.8958
R19692 vdd.n2496 vdd.n810 72.8958
R19693 vdd.n2496 vdd.n811 72.8958
R19694 vdd.n2496 vdd.n812 72.8958
R19695 vdd.n2496 vdd.n813 72.8958
R19696 vdd.n2496 vdd.n814 72.8958
R19697 vdd.n2496 vdd.n815 72.8958
R19698 vdd.n2496 vdd.n816 72.8958
R19699 vdd.n2496 vdd.n817 72.8958
R19700 vdd.n2496 vdd.n818 72.8958
R19701 vdd.n2496 vdd.n819 72.8958
R19702 vdd.n2496 vdd.n820 72.8958
R19703 vdd.n2496 vdd.n821 72.8958
R19704 vdd.n2496 vdd.n822 72.8958
R19705 vdd.n2496 vdd.n823 72.8958
R19706 vdd.n2496 vdd.n824 72.8958
R19707 vdd.n2496 vdd.n825 72.8958
R19708 vdd.n2801 vdd.n2800 72.8958
R19709 vdd.n2800 vdd.n2497 72.8958
R19710 vdd.n2800 vdd.n2498 72.8958
R19711 vdd.n2800 vdd.n2499 72.8958
R19712 vdd.n2800 vdd.n2500 72.8958
R19713 vdd.n2800 vdd.n2501 72.8958
R19714 vdd.n2800 vdd.n2502 72.8958
R19715 vdd.n2800 vdd.n2503 72.8958
R19716 vdd.n2800 vdd.n2504 72.8958
R19717 vdd.n2800 vdd.n2505 72.8958
R19718 vdd.n2800 vdd.n2506 72.8958
R19719 vdd.n2800 vdd.n2507 72.8958
R19720 vdd.n2800 vdd.n2508 72.8958
R19721 vdd.n2800 vdd.n2509 72.8958
R19722 vdd.n2800 vdd.n2510 72.8958
R19723 vdd.n2800 vdd.n2511 72.8958
R19724 vdd.n2800 vdd.n2512 72.8958
R19725 vdd.n2978 vdd.n613 72.8958
R19726 vdd.n2984 vdd.n613 72.8958
R19727 vdd.n659 vdd.n613 72.8958
R19728 vdd.n2991 vdd.n613 72.8958
R19729 vdd.n656 vdd.n613 72.8958
R19730 vdd.n2998 vdd.n613 72.8958
R19731 vdd.n653 vdd.n613 72.8958
R19732 vdd.n3005 vdd.n613 72.8958
R19733 vdd.n650 vdd.n613 72.8958
R19734 vdd.n3013 vdd.n613 72.8958
R19735 vdd.n647 vdd.n613 72.8958
R19736 vdd.n3020 vdd.n613 72.8958
R19737 vdd.n644 vdd.n613 72.8958
R19738 vdd.n3027 vdd.n613 72.8958
R19739 vdd.n641 vdd.n613 72.8958
R19740 vdd.n3034 vdd.n613 72.8958
R19741 vdd.n3037 vdd.n613 72.8958
R19742 vdd.n2496 vdd.n807 72.8958
R19743 vdd.n2496 vdd.n806 72.8958
R19744 vdd.n2496 vdd.n805 72.8958
R19745 vdd.n2496 vdd.n804 72.8958
R19746 vdd.n2496 vdd.n803 72.8958
R19747 vdd.n2496 vdd.n802 72.8958
R19748 vdd.n2496 vdd.n801 72.8958
R19749 vdd.n2496 vdd.n800 72.8958
R19750 vdd.n2496 vdd.n799 72.8958
R19751 vdd.n2496 vdd.n798 72.8958
R19752 vdd.n2496 vdd.n797 72.8958
R19753 vdd.n2496 vdd.n796 72.8958
R19754 vdd.n2496 vdd.n795 72.8958
R19755 vdd.n2496 vdd.n794 72.8958
R19756 vdd.n2496 vdd.n793 72.8958
R19757 vdd.n2496 vdd.n792 72.8958
R19758 vdd.n2496 vdd.n791 72.8958
R19759 vdd.n2218 vdd.n986 72.8958
R19760 vdd.n2218 vdd.n987 72.8958
R19761 vdd.n2218 vdd.n988 72.8958
R19762 vdd.n2218 vdd.n989 72.8958
R19763 vdd.n2218 vdd.n990 72.8958
R19764 vdd.n2218 vdd.n991 72.8958
R19765 vdd.n2218 vdd.n992 72.8958
R19766 vdd.n2218 vdd.n993 72.8958
R19767 vdd.n2218 vdd.n994 72.8958
R19768 vdd.n2218 vdd.n995 72.8958
R19769 vdd.n2218 vdd.n996 72.8958
R19770 vdd.n2218 vdd.n997 72.8958
R19771 vdd.n2218 vdd.n998 72.8958
R19772 vdd.n2218 vdd.n999 72.8958
R19773 vdd.n2218 vdd.n1000 72.8958
R19774 vdd.n2218 vdd.n1001 72.8958
R19775 vdd.n2218 vdd.n1002 72.8958
R19776 vdd.n1441 vdd.n1437 66.2847
R19777 vdd.n1447 vdd.n1437 66.2847
R19778 vdd.n1450 vdd.n1437 66.2847
R19779 vdd.n1455 vdd.n1437 66.2847
R19780 vdd.n1458 vdd.n1437 66.2847
R19781 vdd.n1463 vdd.n1437 66.2847
R19782 vdd.n1466 vdd.n1437 66.2847
R19783 vdd.n1471 vdd.n1437 66.2847
R19784 vdd.n1474 vdd.n1437 66.2847
R19785 vdd.n1481 vdd.n1437 66.2847
R19786 vdd.n1484 vdd.n1437 66.2847
R19787 vdd.n1489 vdd.n1437 66.2847
R19788 vdd.n1492 vdd.n1437 66.2847
R19789 vdd.n1497 vdd.n1437 66.2847
R19790 vdd.n1500 vdd.n1437 66.2847
R19791 vdd.n1505 vdd.n1437 66.2847
R19792 vdd.n1508 vdd.n1437 66.2847
R19793 vdd.n1513 vdd.n1437 66.2847
R19794 vdd.n1516 vdd.n1437 66.2847
R19795 vdd.n1521 vdd.n1437 66.2847
R19796 vdd.n1600 vdd.n1437 66.2847
R19797 vdd.n1524 vdd.n1437 66.2847
R19798 vdd.n1530 vdd.n1437 66.2847
R19799 vdd.n1535 vdd.n1437 66.2847
R19800 vdd.n1538 vdd.n1437 66.2847
R19801 vdd.n1543 vdd.n1437 66.2847
R19802 vdd.n1546 vdd.n1437 66.2847
R19803 vdd.n1551 vdd.n1437 66.2847
R19804 vdd.n1554 vdd.n1437 66.2847
R19805 vdd.n1559 vdd.n1437 66.2847
R19806 vdd.n1562 vdd.n1437 66.2847
R19807 vdd.n1354 vdd.n969 66.2847
R19808 vdd.n1351 vdd.n969 66.2847
R19809 vdd.n1347 vdd.n969 66.2847
R19810 vdd.n2084 vdd.n969 66.2847
R19811 vdd.n1103 vdd.n969 66.2847
R19812 vdd.n2091 vdd.n969 66.2847
R19813 vdd.n1096 vdd.n969 66.2847
R19814 vdd.n2098 vdd.n969 66.2847
R19815 vdd.n1089 vdd.n969 66.2847
R19816 vdd.n2105 vdd.n969 66.2847
R19817 vdd.n1083 vdd.n969 66.2847
R19818 vdd.n1078 vdd.n969 66.2847
R19819 vdd.n2116 vdd.n969 66.2847
R19820 vdd.n1070 vdd.n969 66.2847
R19821 vdd.n2123 vdd.n969 66.2847
R19822 vdd.n1063 vdd.n969 66.2847
R19823 vdd.n2130 vdd.n969 66.2847
R19824 vdd.n1056 vdd.n969 66.2847
R19825 vdd.n2137 vdd.n969 66.2847
R19826 vdd.n1049 vdd.n969 66.2847
R19827 vdd.n2144 vdd.n969 66.2847
R19828 vdd.n1043 vdd.n969 66.2847
R19829 vdd.n1038 vdd.n969 66.2847
R19830 vdd.n2155 vdd.n969 66.2847
R19831 vdd.n1030 vdd.n969 66.2847
R19832 vdd.n2162 vdd.n969 66.2847
R19833 vdd.n1023 vdd.n969 66.2847
R19834 vdd.n2169 vdd.n969 66.2847
R19835 vdd.n1016 vdd.n969 66.2847
R19836 vdd.n2176 vdd.n969 66.2847
R19837 vdd.n2181 vdd.n969 66.2847
R19838 vdd.n1012 vdd.n969 66.2847
R19839 vdd.n3204 vdd.n516 66.2847
R19840 vdd.n520 vdd.n516 66.2847
R19841 vdd.n523 vdd.n516 66.2847
R19842 vdd.n3193 vdd.n516 66.2847
R19843 vdd.n3187 vdd.n516 66.2847
R19844 vdd.n3185 vdd.n516 66.2847
R19845 vdd.n3179 vdd.n516 66.2847
R19846 vdd.n3177 vdd.n516 66.2847
R19847 vdd.n3171 vdd.n516 66.2847
R19848 vdd.n3169 vdd.n516 66.2847
R19849 vdd.n3163 vdd.n516 66.2847
R19850 vdd.n3161 vdd.n516 66.2847
R19851 vdd.n3155 vdd.n516 66.2847
R19852 vdd.n3153 vdd.n516 66.2847
R19853 vdd.n3147 vdd.n516 66.2847
R19854 vdd.n3145 vdd.n516 66.2847
R19855 vdd.n3139 vdd.n516 66.2847
R19856 vdd.n3137 vdd.n516 66.2847
R19857 vdd.n3131 vdd.n516 66.2847
R19858 vdd.n3129 vdd.n516 66.2847
R19859 vdd.n584 vdd.n516 66.2847
R19860 vdd.n3120 vdd.n516 66.2847
R19861 vdd.n586 vdd.n516 66.2847
R19862 vdd.n3113 vdd.n516 66.2847
R19863 vdd.n3107 vdd.n516 66.2847
R19864 vdd.n3105 vdd.n516 66.2847
R19865 vdd.n3099 vdd.n516 66.2847
R19866 vdd.n3097 vdd.n516 66.2847
R19867 vdd.n3091 vdd.n516 66.2847
R19868 vdd.n607 vdd.n516 66.2847
R19869 vdd.n609 vdd.n516 66.2847
R19870 vdd.n3290 vdd.n351 66.2847
R19871 vdd.n3299 vdd.n351 66.2847
R19872 vdd.n461 vdd.n351 66.2847
R19873 vdd.n3306 vdd.n351 66.2847
R19874 vdd.n454 vdd.n351 66.2847
R19875 vdd.n3313 vdd.n351 66.2847
R19876 vdd.n447 vdd.n351 66.2847
R19877 vdd.n3320 vdd.n351 66.2847
R19878 vdd.n440 vdd.n351 66.2847
R19879 vdd.n3327 vdd.n351 66.2847
R19880 vdd.n434 vdd.n351 66.2847
R19881 vdd.n429 vdd.n351 66.2847
R19882 vdd.n3338 vdd.n351 66.2847
R19883 vdd.n421 vdd.n351 66.2847
R19884 vdd.n3345 vdd.n351 66.2847
R19885 vdd.n414 vdd.n351 66.2847
R19886 vdd.n3352 vdd.n351 66.2847
R19887 vdd.n407 vdd.n351 66.2847
R19888 vdd.n3359 vdd.n351 66.2847
R19889 vdd.n400 vdd.n351 66.2847
R19890 vdd.n3366 vdd.n351 66.2847
R19891 vdd.n394 vdd.n351 66.2847
R19892 vdd.n389 vdd.n351 66.2847
R19893 vdd.n3377 vdd.n351 66.2847
R19894 vdd.n381 vdd.n351 66.2847
R19895 vdd.n3384 vdd.n351 66.2847
R19896 vdd.n374 vdd.n351 66.2847
R19897 vdd.n3391 vdd.n351 66.2847
R19898 vdd.n367 vdd.n351 66.2847
R19899 vdd.n3398 vdd.n351 66.2847
R19900 vdd.n3401 vdd.n351 66.2847
R19901 vdd.n355 vdd.n351 66.2847
R19902 vdd.n356 vdd.n355 52.4337
R19903 vdd.n3401 vdd.n3400 52.4337
R19904 vdd.n3398 vdd.n3397 52.4337
R19905 vdd.n3393 vdd.n367 52.4337
R19906 vdd.n3391 vdd.n3390 52.4337
R19907 vdd.n3386 vdd.n374 52.4337
R19908 vdd.n3384 vdd.n3383 52.4337
R19909 vdd.n3379 vdd.n381 52.4337
R19910 vdd.n3377 vdd.n3376 52.4337
R19911 vdd.n390 vdd.n389 52.4337
R19912 vdd.n3368 vdd.n394 52.4337
R19913 vdd.n3366 vdd.n3365 52.4337
R19914 vdd.n3361 vdd.n400 52.4337
R19915 vdd.n3359 vdd.n3358 52.4337
R19916 vdd.n3354 vdd.n407 52.4337
R19917 vdd.n3352 vdd.n3351 52.4337
R19918 vdd.n3347 vdd.n414 52.4337
R19919 vdd.n3345 vdd.n3344 52.4337
R19920 vdd.n3340 vdd.n421 52.4337
R19921 vdd.n3338 vdd.n3337 52.4337
R19922 vdd.n430 vdd.n429 52.4337
R19923 vdd.n3329 vdd.n434 52.4337
R19924 vdd.n3327 vdd.n3326 52.4337
R19925 vdd.n3322 vdd.n440 52.4337
R19926 vdd.n3320 vdd.n3319 52.4337
R19927 vdd.n3315 vdd.n447 52.4337
R19928 vdd.n3313 vdd.n3312 52.4337
R19929 vdd.n3308 vdd.n454 52.4337
R19930 vdd.n3306 vdd.n3305 52.4337
R19931 vdd.n3301 vdd.n461 52.4337
R19932 vdd.n3299 vdd.n3298 52.4337
R19933 vdd.n3291 vdd.n3290 52.4337
R19934 vdd.n3204 vdd.n517 52.4337
R19935 vdd.n3202 vdd.n520 52.4337
R19936 vdd.n3198 vdd.n523 52.4337
R19937 vdd.n3194 vdd.n3193 52.4337
R19938 vdd.n3187 vdd.n526 52.4337
R19939 vdd.n3186 vdd.n3185 52.4337
R19940 vdd.n3179 vdd.n532 52.4337
R19941 vdd.n3178 vdd.n3177 52.4337
R19942 vdd.n3171 vdd.n538 52.4337
R19943 vdd.n3170 vdd.n3169 52.4337
R19944 vdd.n3163 vdd.n546 52.4337
R19945 vdd.n3162 vdd.n3161 52.4337
R19946 vdd.n3155 vdd.n552 52.4337
R19947 vdd.n3154 vdd.n3153 52.4337
R19948 vdd.n3147 vdd.n558 52.4337
R19949 vdd.n3146 vdd.n3145 52.4337
R19950 vdd.n3139 vdd.n564 52.4337
R19951 vdd.n3138 vdd.n3137 52.4337
R19952 vdd.n3131 vdd.n570 52.4337
R19953 vdd.n3130 vdd.n3129 52.4337
R19954 vdd.n584 vdd.n576 52.4337
R19955 vdd.n3121 vdd.n3120 52.4337
R19956 vdd.n3118 vdd.n586 52.4337
R19957 vdd.n3114 vdd.n3113 52.4337
R19958 vdd.n3107 vdd.n590 52.4337
R19959 vdd.n3106 vdd.n3105 52.4337
R19960 vdd.n3099 vdd.n596 52.4337
R19961 vdd.n3098 vdd.n3097 52.4337
R19962 vdd.n3091 vdd.n602 52.4337
R19963 vdd.n3090 vdd.n607 52.4337
R19964 vdd.n3086 vdd.n609 52.4337
R19965 vdd.n2183 vdd.n1012 52.4337
R19966 vdd.n2181 vdd.n2180 52.4337
R19967 vdd.n2176 vdd.n2175 52.4337
R19968 vdd.n2171 vdd.n1016 52.4337
R19969 vdd.n2169 vdd.n2168 52.4337
R19970 vdd.n2164 vdd.n1023 52.4337
R19971 vdd.n2162 vdd.n2161 52.4337
R19972 vdd.n2157 vdd.n1030 52.4337
R19973 vdd.n2155 vdd.n2154 52.4337
R19974 vdd.n1039 vdd.n1038 52.4337
R19975 vdd.n2146 vdd.n1043 52.4337
R19976 vdd.n2144 vdd.n2143 52.4337
R19977 vdd.n2139 vdd.n1049 52.4337
R19978 vdd.n2137 vdd.n2136 52.4337
R19979 vdd.n2132 vdd.n1056 52.4337
R19980 vdd.n2130 vdd.n2129 52.4337
R19981 vdd.n2125 vdd.n1063 52.4337
R19982 vdd.n2123 vdd.n2122 52.4337
R19983 vdd.n2118 vdd.n1070 52.4337
R19984 vdd.n2116 vdd.n2115 52.4337
R19985 vdd.n1079 vdd.n1078 52.4337
R19986 vdd.n2107 vdd.n1083 52.4337
R19987 vdd.n2105 vdd.n2104 52.4337
R19988 vdd.n2100 vdd.n1089 52.4337
R19989 vdd.n2098 vdd.n2097 52.4337
R19990 vdd.n2093 vdd.n1096 52.4337
R19991 vdd.n2091 vdd.n2090 52.4337
R19992 vdd.n2086 vdd.n1103 52.4337
R19993 vdd.n2084 vdd.n2083 52.4337
R19994 vdd.n1348 vdd.n1347 52.4337
R19995 vdd.n1352 vdd.n1351 52.4337
R19996 vdd.n2072 vdd.n1354 52.4337
R19997 vdd.n1441 vdd.n1439 52.4337
R19998 vdd.n1447 vdd.n1446 52.4337
R19999 vdd.n1450 vdd.n1449 52.4337
R20000 vdd.n1455 vdd.n1454 52.4337
R20001 vdd.n1458 vdd.n1457 52.4337
R20002 vdd.n1463 vdd.n1462 52.4337
R20003 vdd.n1466 vdd.n1465 52.4337
R20004 vdd.n1471 vdd.n1470 52.4337
R20005 vdd.n1474 vdd.n1473 52.4337
R20006 vdd.n1481 vdd.n1480 52.4337
R20007 vdd.n1484 vdd.n1483 52.4337
R20008 vdd.n1489 vdd.n1488 52.4337
R20009 vdd.n1492 vdd.n1491 52.4337
R20010 vdd.n1497 vdd.n1496 52.4337
R20011 vdd.n1500 vdd.n1499 52.4337
R20012 vdd.n1505 vdd.n1504 52.4337
R20013 vdd.n1508 vdd.n1507 52.4337
R20014 vdd.n1513 vdd.n1512 52.4337
R20015 vdd.n1516 vdd.n1515 52.4337
R20016 vdd.n1521 vdd.n1520 52.4337
R20017 vdd.n1601 vdd.n1600 52.4337
R20018 vdd.n1598 vdd.n1524 52.4337
R20019 vdd.n1530 vdd.n1529 52.4337
R20020 vdd.n1535 vdd.n1532 52.4337
R20021 vdd.n1538 vdd.n1537 52.4337
R20022 vdd.n1543 vdd.n1540 52.4337
R20023 vdd.n1546 vdd.n1545 52.4337
R20024 vdd.n1551 vdd.n1548 52.4337
R20025 vdd.n1554 vdd.n1553 52.4337
R20026 vdd.n1559 vdd.n1556 52.4337
R20027 vdd.n1562 vdd.n1561 52.4337
R20028 vdd.n1442 vdd.n1441 52.4337
R20029 vdd.n1448 vdd.n1447 52.4337
R20030 vdd.n1451 vdd.n1450 52.4337
R20031 vdd.n1456 vdd.n1455 52.4337
R20032 vdd.n1459 vdd.n1458 52.4337
R20033 vdd.n1464 vdd.n1463 52.4337
R20034 vdd.n1467 vdd.n1466 52.4337
R20035 vdd.n1472 vdd.n1471 52.4337
R20036 vdd.n1475 vdd.n1474 52.4337
R20037 vdd.n1482 vdd.n1481 52.4337
R20038 vdd.n1485 vdd.n1484 52.4337
R20039 vdd.n1490 vdd.n1489 52.4337
R20040 vdd.n1493 vdd.n1492 52.4337
R20041 vdd.n1498 vdd.n1497 52.4337
R20042 vdd.n1501 vdd.n1500 52.4337
R20043 vdd.n1506 vdd.n1505 52.4337
R20044 vdd.n1509 vdd.n1508 52.4337
R20045 vdd.n1514 vdd.n1513 52.4337
R20046 vdd.n1517 vdd.n1516 52.4337
R20047 vdd.n1522 vdd.n1521 52.4337
R20048 vdd.n1600 vdd.n1599 52.4337
R20049 vdd.n1528 vdd.n1524 52.4337
R20050 vdd.n1531 vdd.n1530 52.4337
R20051 vdd.n1536 vdd.n1535 52.4337
R20052 vdd.n1539 vdd.n1538 52.4337
R20053 vdd.n1544 vdd.n1543 52.4337
R20054 vdd.n1547 vdd.n1546 52.4337
R20055 vdd.n1552 vdd.n1551 52.4337
R20056 vdd.n1555 vdd.n1554 52.4337
R20057 vdd.n1560 vdd.n1559 52.4337
R20058 vdd.n1563 vdd.n1562 52.4337
R20059 vdd.n1354 vdd.n1353 52.4337
R20060 vdd.n1351 vdd.n1350 52.4337
R20061 vdd.n1347 vdd.n1104 52.4337
R20062 vdd.n2085 vdd.n2084 52.4337
R20063 vdd.n1103 vdd.n1097 52.4337
R20064 vdd.n2092 vdd.n2091 52.4337
R20065 vdd.n1096 vdd.n1090 52.4337
R20066 vdd.n2099 vdd.n2098 52.4337
R20067 vdd.n1089 vdd.n1084 52.4337
R20068 vdd.n2106 vdd.n2105 52.4337
R20069 vdd.n1083 vdd.n1082 52.4337
R20070 vdd.n1078 vdd.n1071 52.4337
R20071 vdd.n2117 vdd.n2116 52.4337
R20072 vdd.n1070 vdd.n1064 52.4337
R20073 vdd.n2124 vdd.n2123 52.4337
R20074 vdd.n1063 vdd.n1057 52.4337
R20075 vdd.n2131 vdd.n2130 52.4337
R20076 vdd.n1056 vdd.n1050 52.4337
R20077 vdd.n2138 vdd.n2137 52.4337
R20078 vdd.n1049 vdd.n1044 52.4337
R20079 vdd.n2145 vdd.n2144 52.4337
R20080 vdd.n1043 vdd.n1042 52.4337
R20081 vdd.n1038 vdd.n1031 52.4337
R20082 vdd.n2156 vdd.n2155 52.4337
R20083 vdd.n1030 vdd.n1024 52.4337
R20084 vdd.n2163 vdd.n2162 52.4337
R20085 vdd.n1023 vdd.n1017 52.4337
R20086 vdd.n2170 vdd.n2169 52.4337
R20087 vdd.n1016 vdd.n1013 52.4337
R20088 vdd.n2177 vdd.n2176 52.4337
R20089 vdd.n2182 vdd.n2181 52.4337
R20090 vdd.n1358 vdd.n1012 52.4337
R20091 vdd.n3205 vdd.n3204 52.4337
R20092 vdd.n3199 vdd.n520 52.4337
R20093 vdd.n3195 vdd.n523 52.4337
R20094 vdd.n3193 vdd.n3192 52.4337
R20095 vdd.n3188 vdd.n3187 52.4337
R20096 vdd.n3185 vdd.n3184 52.4337
R20097 vdd.n3180 vdd.n3179 52.4337
R20098 vdd.n3177 vdd.n3176 52.4337
R20099 vdd.n3172 vdd.n3171 52.4337
R20100 vdd.n3169 vdd.n3168 52.4337
R20101 vdd.n3164 vdd.n3163 52.4337
R20102 vdd.n3161 vdd.n3160 52.4337
R20103 vdd.n3156 vdd.n3155 52.4337
R20104 vdd.n3153 vdd.n3152 52.4337
R20105 vdd.n3148 vdd.n3147 52.4337
R20106 vdd.n3145 vdd.n3144 52.4337
R20107 vdd.n3140 vdd.n3139 52.4337
R20108 vdd.n3137 vdd.n3136 52.4337
R20109 vdd.n3132 vdd.n3131 52.4337
R20110 vdd.n3129 vdd.n3128 52.4337
R20111 vdd.n585 vdd.n584 52.4337
R20112 vdd.n3120 vdd.n3119 52.4337
R20113 vdd.n3115 vdd.n586 52.4337
R20114 vdd.n3113 vdd.n3112 52.4337
R20115 vdd.n3108 vdd.n3107 52.4337
R20116 vdd.n3105 vdd.n3104 52.4337
R20117 vdd.n3100 vdd.n3099 52.4337
R20118 vdd.n3097 vdd.n3096 52.4337
R20119 vdd.n3092 vdd.n3091 52.4337
R20120 vdd.n3087 vdd.n607 52.4337
R20121 vdd.n3083 vdd.n609 52.4337
R20122 vdd.n3290 vdd.n462 52.4337
R20123 vdd.n3300 vdd.n3299 52.4337
R20124 vdd.n461 vdd.n455 52.4337
R20125 vdd.n3307 vdd.n3306 52.4337
R20126 vdd.n454 vdd.n448 52.4337
R20127 vdd.n3314 vdd.n3313 52.4337
R20128 vdd.n447 vdd.n441 52.4337
R20129 vdd.n3321 vdd.n3320 52.4337
R20130 vdd.n440 vdd.n435 52.4337
R20131 vdd.n3328 vdd.n3327 52.4337
R20132 vdd.n434 vdd.n433 52.4337
R20133 vdd.n429 vdd.n422 52.4337
R20134 vdd.n3339 vdd.n3338 52.4337
R20135 vdd.n421 vdd.n415 52.4337
R20136 vdd.n3346 vdd.n3345 52.4337
R20137 vdd.n414 vdd.n408 52.4337
R20138 vdd.n3353 vdd.n3352 52.4337
R20139 vdd.n407 vdd.n401 52.4337
R20140 vdd.n3360 vdd.n3359 52.4337
R20141 vdd.n400 vdd.n395 52.4337
R20142 vdd.n3367 vdd.n3366 52.4337
R20143 vdd.n394 vdd.n393 52.4337
R20144 vdd.n389 vdd.n382 52.4337
R20145 vdd.n3378 vdd.n3377 52.4337
R20146 vdd.n381 vdd.n375 52.4337
R20147 vdd.n3385 vdd.n3384 52.4337
R20148 vdd.n374 vdd.n368 52.4337
R20149 vdd.n3392 vdd.n3391 52.4337
R20150 vdd.n367 vdd.n360 52.4337
R20151 vdd.n3399 vdd.n3398 52.4337
R20152 vdd.n3402 vdd.n3401 52.4337
R20153 vdd.n355 vdd.n352 52.4337
R20154 vdd.t91 vdd.t104 51.4683
R20155 vdd.n258 vdd.n256 42.0461
R20156 vdd.n164 vdd.n162 42.0461
R20157 vdd.n71 vdd.n69 42.0461
R20158 vdd.n1959 vdd.n1957 42.0461
R20159 vdd.n1865 vdd.n1863 42.0461
R20160 vdd.n1772 vdd.n1770 42.0461
R20161 vdd.n308 vdd.n307 41.6884
R20162 vdd.n214 vdd.n213 41.6884
R20163 vdd.n121 vdd.n120 41.6884
R20164 vdd.n2009 vdd.n2008 41.6884
R20165 vdd.n1915 vdd.n1914 41.6884
R20166 vdd.n1822 vdd.n1821 41.6884
R20167 vdd.n1567 vdd.n1566 41.1157
R20168 vdd.n1604 vdd.n1603 41.1157
R20169 vdd.n1478 vdd.n1477 41.1157
R20170 vdd.n3295 vdd.n3294 41.1157
R20171 vdd.n3334 vdd.n428 41.1157
R20172 vdd.n3373 vdd.n388 41.1157
R20173 vdd.n3037 vdd.n3036 39.2114
R20174 vdd.n3034 vdd.n3033 39.2114
R20175 vdd.n3029 vdd.n641 39.2114
R20176 vdd.n3027 vdd.n3026 39.2114
R20177 vdd.n3022 vdd.n644 39.2114
R20178 vdd.n3020 vdd.n3019 39.2114
R20179 vdd.n3015 vdd.n647 39.2114
R20180 vdd.n3013 vdd.n3012 39.2114
R20181 vdd.n3007 vdd.n650 39.2114
R20182 vdd.n3005 vdd.n3004 39.2114
R20183 vdd.n3000 vdd.n653 39.2114
R20184 vdd.n2998 vdd.n2997 39.2114
R20185 vdd.n2993 vdd.n656 39.2114
R20186 vdd.n2991 vdd.n2990 39.2114
R20187 vdd.n2986 vdd.n659 39.2114
R20188 vdd.n2984 vdd.n2983 39.2114
R20189 vdd.n2979 vdd.n2978 39.2114
R20190 vdd.n2802 vdd.n2801 39.2114
R20191 vdd.n2531 vdd.n2497 39.2114
R20192 vdd.n2794 vdd.n2498 39.2114
R20193 vdd.n2790 vdd.n2499 39.2114
R20194 vdd.n2786 vdd.n2500 39.2114
R20195 vdd.n2782 vdd.n2501 39.2114
R20196 vdd.n2778 vdd.n2502 39.2114
R20197 vdd.n2774 vdd.n2503 39.2114
R20198 vdd.n2770 vdd.n2504 39.2114
R20199 vdd.n2766 vdd.n2505 39.2114
R20200 vdd.n2762 vdd.n2506 39.2114
R20201 vdd.n2758 vdd.n2507 39.2114
R20202 vdd.n2754 vdd.n2508 39.2114
R20203 vdd.n2750 vdd.n2509 39.2114
R20204 vdd.n2746 vdd.n2510 39.2114
R20205 vdd.n2742 vdd.n2511 39.2114
R20206 vdd.n2737 vdd.n2512 39.2114
R20207 vdd.n2491 vdd.n825 39.2114
R20208 vdd.n2487 vdd.n824 39.2114
R20209 vdd.n2483 vdd.n823 39.2114
R20210 vdd.n2479 vdd.n822 39.2114
R20211 vdd.n2475 vdd.n821 39.2114
R20212 vdd.n2471 vdd.n820 39.2114
R20213 vdd.n2467 vdd.n819 39.2114
R20214 vdd.n2463 vdd.n818 39.2114
R20215 vdd.n2459 vdd.n817 39.2114
R20216 vdd.n2455 vdd.n816 39.2114
R20217 vdd.n2451 vdd.n815 39.2114
R20218 vdd.n2447 vdd.n814 39.2114
R20219 vdd.n2443 vdd.n813 39.2114
R20220 vdd.n2439 vdd.n812 39.2114
R20221 vdd.n2435 vdd.n811 39.2114
R20222 vdd.n2430 vdd.n810 39.2114
R20223 vdd.n2426 vdd.n809 39.2114
R20224 vdd.n2220 vdd.n2219 39.2114
R20225 vdd.n1004 vdd.n970 39.2114
R20226 vdd.n2212 vdd.n971 39.2114
R20227 vdd.n2208 vdd.n972 39.2114
R20228 vdd.n2204 vdd.n973 39.2114
R20229 vdd.n2200 vdd.n974 39.2114
R20230 vdd.n2196 vdd.n975 39.2114
R20231 vdd.n2192 vdd.n976 39.2114
R20232 vdd.n2188 vdd.n977 39.2114
R20233 vdd.n1150 vdd.n978 39.2114
R20234 vdd.n1154 vdd.n979 39.2114
R20235 vdd.n1158 vdd.n980 39.2114
R20236 vdd.n1162 vdd.n981 39.2114
R20237 vdd.n1166 vdd.n982 39.2114
R20238 vdd.n1170 vdd.n983 39.2114
R20239 vdd.n1174 vdd.n984 39.2114
R20240 vdd.n1179 vdd.n985 39.2114
R20241 vdd.n2956 vdd.n2955 39.2114
R20242 vdd.n2951 vdd.n2923 39.2114
R20243 vdd.n2949 vdd.n2948 39.2114
R20244 vdd.n2944 vdd.n2926 39.2114
R20245 vdd.n2942 vdd.n2941 39.2114
R20246 vdd.n2937 vdd.n2929 39.2114
R20247 vdd.n2935 vdd.n2934 39.2114
R20248 vdd.n2930 vdd.n612 39.2114
R20249 vdd.n3074 vdd.n3073 39.2114
R20250 vdd.n3071 vdd.n3070 39.2114
R20251 vdd.n3066 vdd.n617 39.2114
R20252 vdd.n3064 vdd.n3063 39.2114
R20253 vdd.n3059 vdd.n620 39.2114
R20254 vdd.n3057 vdd.n3056 39.2114
R20255 vdd.n3052 vdd.n623 39.2114
R20256 vdd.n3050 vdd.n3049 39.2114
R20257 vdd.n3045 vdd.n629 39.2114
R20258 vdd.n2538 vdd.n2513 39.2114
R20259 vdd.n2542 vdd.n2514 39.2114
R20260 vdd.n2546 vdd.n2515 39.2114
R20261 vdd.n2550 vdd.n2516 39.2114
R20262 vdd.n2554 vdd.n2517 39.2114
R20263 vdd.n2558 vdd.n2518 39.2114
R20264 vdd.n2562 vdd.n2519 39.2114
R20265 vdd.n2566 vdd.n2520 39.2114
R20266 vdd.n2570 vdd.n2521 39.2114
R20267 vdd.n2574 vdd.n2522 39.2114
R20268 vdd.n2578 vdd.n2523 39.2114
R20269 vdd.n2582 vdd.n2524 39.2114
R20270 vdd.n2586 vdd.n2525 39.2114
R20271 vdd.n2590 vdd.n2526 39.2114
R20272 vdd.n2594 vdd.n2527 39.2114
R20273 vdd.n2598 vdd.n2528 39.2114
R20274 vdd.n2602 vdd.n2529 39.2114
R20275 vdd.n2541 vdd.n2513 39.2114
R20276 vdd.n2545 vdd.n2514 39.2114
R20277 vdd.n2549 vdd.n2515 39.2114
R20278 vdd.n2553 vdd.n2516 39.2114
R20279 vdd.n2557 vdd.n2517 39.2114
R20280 vdd.n2561 vdd.n2518 39.2114
R20281 vdd.n2565 vdd.n2519 39.2114
R20282 vdd.n2569 vdd.n2520 39.2114
R20283 vdd.n2573 vdd.n2521 39.2114
R20284 vdd.n2577 vdd.n2522 39.2114
R20285 vdd.n2581 vdd.n2523 39.2114
R20286 vdd.n2585 vdd.n2524 39.2114
R20287 vdd.n2589 vdd.n2525 39.2114
R20288 vdd.n2593 vdd.n2526 39.2114
R20289 vdd.n2597 vdd.n2527 39.2114
R20290 vdd.n2601 vdd.n2528 39.2114
R20291 vdd.n2604 vdd.n2529 39.2114
R20292 vdd.n629 vdd.n624 39.2114
R20293 vdd.n3051 vdd.n3050 39.2114
R20294 vdd.n623 vdd.n621 39.2114
R20295 vdd.n3058 vdd.n3057 39.2114
R20296 vdd.n620 vdd.n618 39.2114
R20297 vdd.n3065 vdd.n3064 39.2114
R20298 vdd.n617 vdd.n615 39.2114
R20299 vdd.n3072 vdd.n3071 39.2114
R20300 vdd.n3075 vdd.n3074 39.2114
R20301 vdd.n2931 vdd.n2930 39.2114
R20302 vdd.n2936 vdd.n2935 39.2114
R20303 vdd.n2929 vdd.n2927 39.2114
R20304 vdd.n2943 vdd.n2942 39.2114
R20305 vdd.n2926 vdd.n2924 39.2114
R20306 vdd.n2950 vdd.n2949 39.2114
R20307 vdd.n2923 vdd.n2921 39.2114
R20308 vdd.n2957 vdd.n2956 39.2114
R20309 vdd.n2219 vdd.n968 39.2114
R20310 vdd.n2213 vdd.n970 39.2114
R20311 vdd.n2209 vdd.n971 39.2114
R20312 vdd.n2205 vdd.n972 39.2114
R20313 vdd.n2201 vdd.n973 39.2114
R20314 vdd.n2197 vdd.n974 39.2114
R20315 vdd.n2193 vdd.n975 39.2114
R20316 vdd.n2189 vdd.n976 39.2114
R20317 vdd.n1149 vdd.n977 39.2114
R20318 vdd.n1153 vdd.n978 39.2114
R20319 vdd.n1157 vdd.n979 39.2114
R20320 vdd.n1161 vdd.n980 39.2114
R20321 vdd.n1165 vdd.n981 39.2114
R20322 vdd.n1169 vdd.n982 39.2114
R20323 vdd.n1173 vdd.n983 39.2114
R20324 vdd.n1178 vdd.n984 39.2114
R20325 vdd.n1182 vdd.n985 39.2114
R20326 vdd.n2429 vdd.n809 39.2114
R20327 vdd.n2434 vdd.n810 39.2114
R20328 vdd.n2438 vdd.n811 39.2114
R20329 vdd.n2442 vdd.n812 39.2114
R20330 vdd.n2446 vdd.n813 39.2114
R20331 vdd.n2450 vdd.n814 39.2114
R20332 vdd.n2454 vdd.n815 39.2114
R20333 vdd.n2458 vdd.n816 39.2114
R20334 vdd.n2462 vdd.n817 39.2114
R20335 vdd.n2466 vdd.n818 39.2114
R20336 vdd.n2470 vdd.n819 39.2114
R20337 vdd.n2474 vdd.n820 39.2114
R20338 vdd.n2478 vdd.n821 39.2114
R20339 vdd.n2482 vdd.n822 39.2114
R20340 vdd.n2486 vdd.n823 39.2114
R20341 vdd.n2490 vdd.n824 39.2114
R20342 vdd.n827 vdd.n825 39.2114
R20343 vdd.n2801 vdd.n790 39.2114
R20344 vdd.n2795 vdd.n2497 39.2114
R20345 vdd.n2791 vdd.n2498 39.2114
R20346 vdd.n2787 vdd.n2499 39.2114
R20347 vdd.n2783 vdd.n2500 39.2114
R20348 vdd.n2779 vdd.n2501 39.2114
R20349 vdd.n2775 vdd.n2502 39.2114
R20350 vdd.n2771 vdd.n2503 39.2114
R20351 vdd.n2767 vdd.n2504 39.2114
R20352 vdd.n2763 vdd.n2505 39.2114
R20353 vdd.n2759 vdd.n2506 39.2114
R20354 vdd.n2755 vdd.n2507 39.2114
R20355 vdd.n2751 vdd.n2508 39.2114
R20356 vdd.n2747 vdd.n2509 39.2114
R20357 vdd.n2743 vdd.n2510 39.2114
R20358 vdd.n2738 vdd.n2511 39.2114
R20359 vdd.n2734 vdd.n2512 39.2114
R20360 vdd.n2978 vdd.n660 39.2114
R20361 vdd.n2985 vdd.n2984 39.2114
R20362 vdd.n659 vdd.n657 39.2114
R20363 vdd.n2992 vdd.n2991 39.2114
R20364 vdd.n656 vdd.n654 39.2114
R20365 vdd.n2999 vdd.n2998 39.2114
R20366 vdd.n653 vdd.n651 39.2114
R20367 vdd.n3006 vdd.n3005 39.2114
R20368 vdd.n650 vdd.n648 39.2114
R20369 vdd.n3014 vdd.n3013 39.2114
R20370 vdd.n647 vdd.n645 39.2114
R20371 vdd.n3021 vdd.n3020 39.2114
R20372 vdd.n644 vdd.n642 39.2114
R20373 vdd.n3028 vdd.n3027 39.2114
R20374 vdd.n641 vdd.n639 39.2114
R20375 vdd.n3035 vdd.n3034 39.2114
R20376 vdd.n3038 vdd.n3037 39.2114
R20377 vdd.n836 vdd.n791 39.2114
R20378 vdd.n2418 vdd.n792 39.2114
R20379 vdd.n2414 vdd.n793 39.2114
R20380 vdd.n2410 vdd.n794 39.2114
R20381 vdd.n2406 vdd.n795 39.2114
R20382 vdd.n2402 vdd.n796 39.2114
R20383 vdd.n2398 vdd.n797 39.2114
R20384 vdd.n2394 vdd.n798 39.2114
R20385 vdd.n2390 vdd.n799 39.2114
R20386 vdd.n2386 vdd.n800 39.2114
R20387 vdd.n2382 vdd.n801 39.2114
R20388 vdd.n2378 vdd.n802 39.2114
R20389 vdd.n2374 vdd.n803 39.2114
R20390 vdd.n2370 vdd.n804 39.2114
R20391 vdd.n2366 vdd.n805 39.2114
R20392 vdd.n2362 vdd.n806 39.2114
R20393 vdd.n2358 vdd.n807 39.2114
R20394 vdd.n1108 vdd.n986 39.2114
R20395 vdd.n1112 vdd.n987 39.2114
R20396 vdd.n1116 vdd.n988 39.2114
R20397 vdd.n1120 vdd.n989 39.2114
R20398 vdd.n1124 vdd.n990 39.2114
R20399 vdd.n1128 vdd.n991 39.2114
R20400 vdd.n1132 vdd.n992 39.2114
R20401 vdd.n1136 vdd.n993 39.2114
R20402 vdd.n1140 vdd.n994 39.2114
R20403 vdd.n1341 vdd.n995 39.2114
R20404 vdd.n1338 vdd.n996 39.2114
R20405 vdd.n1334 vdd.n997 39.2114
R20406 vdd.n1330 vdd.n998 39.2114
R20407 vdd.n1326 vdd.n999 39.2114
R20408 vdd.n1322 vdd.n1000 39.2114
R20409 vdd.n1318 vdd.n1001 39.2114
R20410 vdd.n1314 vdd.n1002 39.2114
R20411 vdd.n2355 vdd.n807 39.2114
R20412 vdd.n2359 vdd.n806 39.2114
R20413 vdd.n2363 vdd.n805 39.2114
R20414 vdd.n2367 vdd.n804 39.2114
R20415 vdd.n2371 vdd.n803 39.2114
R20416 vdd.n2375 vdd.n802 39.2114
R20417 vdd.n2379 vdd.n801 39.2114
R20418 vdd.n2383 vdd.n800 39.2114
R20419 vdd.n2387 vdd.n799 39.2114
R20420 vdd.n2391 vdd.n798 39.2114
R20421 vdd.n2395 vdd.n797 39.2114
R20422 vdd.n2399 vdd.n796 39.2114
R20423 vdd.n2403 vdd.n795 39.2114
R20424 vdd.n2407 vdd.n794 39.2114
R20425 vdd.n2411 vdd.n793 39.2114
R20426 vdd.n2415 vdd.n792 39.2114
R20427 vdd.n2419 vdd.n791 39.2114
R20428 vdd.n1111 vdd.n986 39.2114
R20429 vdd.n1115 vdd.n987 39.2114
R20430 vdd.n1119 vdd.n988 39.2114
R20431 vdd.n1123 vdd.n989 39.2114
R20432 vdd.n1127 vdd.n990 39.2114
R20433 vdd.n1131 vdd.n991 39.2114
R20434 vdd.n1135 vdd.n992 39.2114
R20435 vdd.n1139 vdd.n993 39.2114
R20436 vdd.n1142 vdd.n994 39.2114
R20437 vdd.n1339 vdd.n995 39.2114
R20438 vdd.n1335 vdd.n996 39.2114
R20439 vdd.n1331 vdd.n997 39.2114
R20440 vdd.n1327 vdd.n998 39.2114
R20441 vdd.n1323 vdd.n999 39.2114
R20442 vdd.n1319 vdd.n1000 39.2114
R20443 vdd.n1315 vdd.n1001 39.2114
R20444 vdd.n1311 vdd.n1002 39.2114
R20445 vdd.n2076 vdd.n2075 37.2369
R20446 vdd.n2112 vdd.n1077 37.2369
R20447 vdd.n2151 vdd.n1037 37.2369
R20448 vdd.n3126 vdd.n581 37.2369
R20449 vdd.n545 vdd.n544 37.2369
R20450 vdd.n3082 vdd.n3081 37.2369
R20451 vdd.n1145 vdd.n1144 30.449
R20452 vdd.n840 vdd.n839 30.449
R20453 vdd.n1176 vdd.n1148 30.449
R20454 vdd.n2432 vdd.n830 30.449
R20455 vdd.n2537 vdd.n2536 30.449
R20456 vdd.n663 vdd.n662 30.449
R20457 vdd.n2740 vdd.n2533 30.449
R20458 vdd.n627 vdd.n626 30.449
R20459 vdd.n2222 vdd.n2221 29.8151
R20460 vdd.n2494 vdd.n828 29.8151
R20461 vdd.n2427 vdd.n831 29.8151
R20462 vdd.n1184 vdd.n1181 29.8151
R20463 vdd.n2735 vdd.n2732 29.8151
R20464 vdd.n2980 vdd.n2977 29.8151
R20465 vdd.n2804 vdd.n2803 29.8151
R20466 vdd.n3041 vdd.n3040 29.8151
R20467 vdd.n2960 vdd.n2959 29.8151
R20468 vdd.n3046 vdd.n628 29.8151
R20469 vdd.n2608 vdd.n2606 29.8151
R20470 vdd.n2539 vdd.n783 29.8151
R20471 vdd.n1109 vdd.n960 29.8151
R20472 vdd.n2422 vdd.n2421 29.8151
R20473 vdd.n2354 vdd.n2353 29.8151
R20474 vdd.n1310 vdd.n1309 29.8151
R20475 vdd.n1670 vdd.n1437 20.633
R20476 vdd.n2070 vdd.n969 20.633
R20477 vdd.n3212 vdd.n516 20.633
R20478 vdd.n3410 vdd.n351 20.633
R20479 vdd.n1672 vdd.n1434 19.3944
R20480 vdd.n1676 vdd.n1434 19.3944
R20481 vdd.n1676 vdd.n1425 19.3944
R20482 vdd.n1688 vdd.n1425 19.3944
R20483 vdd.n1688 vdd.n1423 19.3944
R20484 vdd.n1692 vdd.n1423 19.3944
R20485 vdd.n1692 vdd.n1412 19.3944
R20486 vdd.n1704 vdd.n1412 19.3944
R20487 vdd.n1704 vdd.n1410 19.3944
R20488 vdd.n1708 vdd.n1410 19.3944
R20489 vdd.n1708 vdd.n1401 19.3944
R20490 vdd.n1721 vdd.n1401 19.3944
R20491 vdd.n1721 vdd.n1399 19.3944
R20492 vdd.n1725 vdd.n1399 19.3944
R20493 vdd.n1725 vdd.n1390 19.3944
R20494 vdd.n2019 vdd.n1390 19.3944
R20495 vdd.n2019 vdd.n1388 19.3944
R20496 vdd.n2023 vdd.n1388 19.3944
R20497 vdd.n2023 vdd.n1378 19.3944
R20498 vdd.n2036 vdd.n1378 19.3944
R20499 vdd.n2036 vdd.n1376 19.3944
R20500 vdd.n2040 vdd.n1376 19.3944
R20501 vdd.n2040 vdd.n1368 19.3944
R20502 vdd.n2053 vdd.n1368 19.3944
R20503 vdd.n2053 vdd.n1365 19.3944
R20504 vdd.n2059 vdd.n1365 19.3944
R20505 vdd.n2059 vdd.n1366 19.3944
R20506 vdd.n1366 vdd.n1356 19.3944
R20507 vdd.n1597 vdd.n1523 19.3944
R20508 vdd.n1597 vdd.n1525 19.3944
R20509 vdd.n1593 vdd.n1525 19.3944
R20510 vdd.n1593 vdd.n1592 19.3944
R20511 vdd.n1592 vdd.n1591 19.3944
R20512 vdd.n1591 vdd.n1533 19.3944
R20513 vdd.n1587 vdd.n1533 19.3944
R20514 vdd.n1587 vdd.n1586 19.3944
R20515 vdd.n1586 vdd.n1585 19.3944
R20516 vdd.n1585 vdd.n1541 19.3944
R20517 vdd.n1581 vdd.n1541 19.3944
R20518 vdd.n1581 vdd.n1580 19.3944
R20519 vdd.n1580 vdd.n1579 19.3944
R20520 vdd.n1579 vdd.n1549 19.3944
R20521 vdd.n1575 vdd.n1549 19.3944
R20522 vdd.n1575 vdd.n1574 19.3944
R20523 vdd.n1574 vdd.n1573 19.3944
R20524 vdd.n1573 vdd.n1557 19.3944
R20525 vdd.n1569 vdd.n1557 19.3944
R20526 vdd.n1569 vdd.n1568 19.3944
R20527 vdd.n1635 vdd.n1634 19.3944
R20528 vdd.n1634 vdd.n1633 19.3944
R20529 vdd.n1633 vdd.n1486 19.3944
R20530 vdd.n1629 vdd.n1486 19.3944
R20531 vdd.n1629 vdd.n1628 19.3944
R20532 vdd.n1628 vdd.n1627 19.3944
R20533 vdd.n1627 vdd.n1494 19.3944
R20534 vdd.n1623 vdd.n1494 19.3944
R20535 vdd.n1623 vdd.n1622 19.3944
R20536 vdd.n1622 vdd.n1621 19.3944
R20537 vdd.n1621 vdd.n1502 19.3944
R20538 vdd.n1617 vdd.n1502 19.3944
R20539 vdd.n1617 vdd.n1616 19.3944
R20540 vdd.n1616 vdd.n1615 19.3944
R20541 vdd.n1615 vdd.n1510 19.3944
R20542 vdd.n1611 vdd.n1510 19.3944
R20543 vdd.n1611 vdd.n1610 19.3944
R20544 vdd.n1610 vdd.n1609 19.3944
R20545 vdd.n1609 vdd.n1518 19.3944
R20546 vdd.n1605 vdd.n1518 19.3944
R20547 vdd.n1665 vdd.n1664 19.3944
R20548 vdd.n1664 vdd.n1663 19.3944
R20549 vdd.n1663 vdd.n1444 19.3944
R20550 vdd.n1659 vdd.n1444 19.3944
R20551 vdd.n1659 vdd.n1658 19.3944
R20552 vdd.n1658 vdd.n1657 19.3944
R20553 vdd.n1657 vdd.n1452 19.3944
R20554 vdd.n1653 vdd.n1452 19.3944
R20555 vdd.n1653 vdd.n1652 19.3944
R20556 vdd.n1652 vdd.n1651 19.3944
R20557 vdd.n1651 vdd.n1460 19.3944
R20558 vdd.n1647 vdd.n1460 19.3944
R20559 vdd.n1647 vdd.n1646 19.3944
R20560 vdd.n1646 vdd.n1645 19.3944
R20561 vdd.n1645 vdd.n1468 19.3944
R20562 vdd.n1641 vdd.n1468 19.3944
R20563 vdd.n1641 vdd.n1640 19.3944
R20564 vdd.n1640 vdd.n1639 19.3944
R20565 vdd.n2108 vdd.n1075 19.3944
R20566 vdd.n2108 vdd.n1081 19.3944
R20567 vdd.n2103 vdd.n1081 19.3944
R20568 vdd.n2103 vdd.n2102 19.3944
R20569 vdd.n2102 vdd.n2101 19.3944
R20570 vdd.n2101 vdd.n1088 19.3944
R20571 vdd.n2096 vdd.n1088 19.3944
R20572 vdd.n2096 vdd.n2095 19.3944
R20573 vdd.n2095 vdd.n2094 19.3944
R20574 vdd.n2094 vdd.n1095 19.3944
R20575 vdd.n2089 vdd.n1095 19.3944
R20576 vdd.n2089 vdd.n2088 19.3944
R20577 vdd.n2088 vdd.n2087 19.3944
R20578 vdd.n2087 vdd.n1102 19.3944
R20579 vdd.n2082 vdd.n1102 19.3944
R20580 vdd.n2082 vdd.n2081 19.3944
R20581 vdd.n1349 vdd.n1107 19.3944
R20582 vdd.n2077 vdd.n1346 19.3944
R20583 vdd.n2147 vdd.n1035 19.3944
R20584 vdd.n2147 vdd.n1041 19.3944
R20585 vdd.n2142 vdd.n1041 19.3944
R20586 vdd.n2142 vdd.n2141 19.3944
R20587 vdd.n2141 vdd.n2140 19.3944
R20588 vdd.n2140 vdd.n1048 19.3944
R20589 vdd.n2135 vdd.n1048 19.3944
R20590 vdd.n2135 vdd.n2134 19.3944
R20591 vdd.n2134 vdd.n2133 19.3944
R20592 vdd.n2133 vdd.n1055 19.3944
R20593 vdd.n2128 vdd.n1055 19.3944
R20594 vdd.n2128 vdd.n2127 19.3944
R20595 vdd.n2127 vdd.n2126 19.3944
R20596 vdd.n2126 vdd.n1062 19.3944
R20597 vdd.n2121 vdd.n1062 19.3944
R20598 vdd.n2121 vdd.n2120 19.3944
R20599 vdd.n2120 vdd.n2119 19.3944
R20600 vdd.n2119 vdd.n1069 19.3944
R20601 vdd.n2114 vdd.n1069 19.3944
R20602 vdd.n2114 vdd.n2113 19.3944
R20603 vdd.n2184 vdd.n1010 19.3944
R20604 vdd.n2184 vdd.n1011 19.3944
R20605 vdd.n2179 vdd.n2178 19.3944
R20606 vdd.n2174 vdd.n2173 19.3944
R20607 vdd.n2173 vdd.n2172 19.3944
R20608 vdd.n2172 vdd.n1015 19.3944
R20609 vdd.n2167 vdd.n1015 19.3944
R20610 vdd.n2167 vdd.n2166 19.3944
R20611 vdd.n2166 vdd.n2165 19.3944
R20612 vdd.n2165 vdd.n1022 19.3944
R20613 vdd.n2160 vdd.n1022 19.3944
R20614 vdd.n2160 vdd.n2159 19.3944
R20615 vdd.n2159 vdd.n2158 19.3944
R20616 vdd.n2158 vdd.n1029 19.3944
R20617 vdd.n2153 vdd.n1029 19.3944
R20618 vdd.n2153 vdd.n2152 19.3944
R20619 vdd.n1668 vdd.n1431 19.3944
R20620 vdd.n1680 vdd.n1431 19.3944
R20621 vdd.n1680 vdd.n1429 19.3944
R20622 vdd.n1684 vdd.n1429 19.3944
R20623 vdd.n1684 vdd.n1419 19.3944
R20624 vdd.n1696 vdd.n1419 19.3944
R20625 vdd.n1696 vdd.n1417 19.3944
R20626 vdd.n1700 vdd.n1417 19.3944
R20627 vdd.n1700 vdd.n1407 19.3944
R20628 vdd.n1713 vdd.n1407 19.3944
R20629 vdd.n1713 vdd.n1405 19.3944
R20630 vdd.n1717 vdd.n1405 19.3944
R20631 vdd.n1717 vdd.n1396 19.3944
R20632 vdd.n1729 vdd.n1396 19.3944
R20633 vdd.n1729 vdd.n1394 19.3944
R20634 vdd.n2015 vdd.n1394 19.3944
R20635 vdd.n2015 vdd.n1384 19.3944
R20636 vdd.n2028 vdd.n1384 19.3944
R20637 vdd.n2028 vdd.n1382 19.3944
R20638 vdd.n2032 vdd.n1382 19.3944
R20639 vdd.n2032 vdd.n1373 19.3944
R20640 vdd.n2045 vdd.n1373 19.3944
R20641 vdd.n2045 vdd.n1371 19.3944
R20642 vdd.n2049 vdd.n1371 19.3944
R20643 vdd.n2049 vdd.n1361 19.3944
R20644 vdd.n2064 vdd.n1361 19.3944
R20645 vdd.n2064 vdd.n1359 19.3944
R20646 vdd.n2068 vdd.n1359 19.3944
R20647 vdd.n3214 vdd.n513 19.3944
R20648 vdd.n3218 vdd.n513 19.3944
R20649 vdd.n3218 vdd.n503 19.3944
R20650 vdd.n3230 vdd.n503 19.3944
R20651 vdd.n3230 vdd.n501 19.3944
R20652 vdd.n3234 vdd.n501 19.3944
R20653 vdd.n3234 vdd.n490 19.3944
R20654 vdd.n3246 vdd.n490 19.3944
R20655 vdd.n3246 vdd.n488 19.3944
R20656 vdd.n3250 vdd.n488 19.3944
R20657 vdd.n3250 vdd.n478 19.3944
R20658 vdd.n3263 vdd.n478 19.3944
R20659 vdd.n3263 vdd.n476 19.3944
R20660 vdd.n3267 vdd.n476 19.3944
R20661 vdd.n3268 vdd.n3267 19.3944
R20662 vdd.n3269 vdd.n3268 19.3944
R20663 vdd.n3269 vdd.n474 19.3944
R20664 vdd.n3273 vdd.n474 19.3944
R20665 vdd.n3274 vdd.n3273 19.3944
R20666 vdd.n3275 vdd.n3274 19.3944
R20667 vdd.n3275 vdd.n471 19.3944
R20668 vdd.n3279 vdd.n471 19.3944
R20669 vdd.n3280 vdd.n3279 19.3944
R20670 vdd.n3281 vdd.n3280 19.3944
R20671 vdd.n3281 vdd.n468 19.3944
R20672 vdd.n3285 vdd.n468 19.3944
R20673 vdd.n3286 vdd.n3285 19.3944
R20674 vdd.n3287 vdd.n3286 19.3944
R20675 vdd.n3330 vdd.n426 19.3944
R20676 vdd.n3330 vdd.n432 19.3944
R20677 vdd.n3325 vdd.n432 19.3944
R20678 vdd.n3325 vdd.n3324 19.3944
R20679 vdd.n3324 vdd.n3323 19.3944
R20680 vdd.n3323 vdd.n439 19.3944
R20681 vdd.n3318 vdd.n439 19.3944
R20682 vdd.n3318 vdd.n3317 19.3944
R20683 vdd.n3317 vdd.n3316 19.3944
R20684 vdd.n3316 vdd.n446 19.3944
R20685 vdd.n3311 vdd.n446 19.3944
R20686 vdd.n3311 vdd.n3310 19.3944
R20687 vdd.n3310 vdd.n3309 19.3944
R20688 vdd.n3309 vdd.n453 19.3944
R20689 vdd.n3304 vdd.n453 19.3944
R20690 vdd.n3304 vdd.n3303 19.3944
R20691 vdd.n3303 vdd.n3302 19.3944
R20692 vdd.n3302 vdd.n460 19.3944
R20693 vdd.n3297 vdd.n460 19.3944
R20694 vdd.n3297 vdd.n3296 19.3944
R20695 vdd.n3369 vdd.n386 19.3944
R20696 vdd.n3369 vdd.n392 19.3944
R20697 vdd.n3364 vdd.n392 19.3944
R20698 vdd.n3364 vdd.n3363 19.3944
R20699 vdd.n3363 vdd.n3362 19.3944
R20700 vdd.n3362 vdd.n399 19.3944
R20701 vdd.n3357 vdd.n399 19.3944
R20702 vdd.n3357 vdd.n3356 19.3944
R20703 vdd.n3356 vdd.n3355 19.3944
R20704 vdd.n3355 vdd.n406 19.3944
R20705 vdd.n3350 vdd.n406 19.3944
R20706 vdd.n3350 vdd.n3349 19.3944
R20707 vdd.n3349 vdd.n3348 19.3944
R20708 vdd.n3348 vdd.n413 19.3944
R20709 vdd.n3343 vdd.n413 19.3944
R20710 vdd.n3343 vdd.n3342 19.3944
R20711 vdd.n3342 vdd.n3341 19.3944
R20712 vdd.n3341 vdd.n420 19.3944
R20713 vdd.n3336 vdd.n420 19.3944
R20714 vdd.n3336 vdd.n3335 19.3944
R20715 vdd.n3405 vdd.n3404 19.3944
R20716 vdd.n3404 vdd.n3403 19.3944
R20717 vdd.n3403 vdd.n358 19.3944
R20718 vdd.n359 vdd.n358 19.3944
R20719 vdd.n3396 vdd.n359 19.3944
R20720 vdd.n3396 vdd.n3395 19.3944
R20721 vdd.n3395 vdd.n3394 19.3944
R20722 vdd.n3394 vdd.n366 19.3944
R20723 vdd.n3389 vdd.n366 19.3944
R20724 vdd.n3389 vdd.n3388 19.3944
R20725 vdd.n3388 vdd.n3387 19.3944
R20726 vdd.n3387 vdd.n373 19.3944
R20727 vdd.n3382 vdd.n373 19.3944
R20728 vdd.n3382 vdd.n3381 19.3944
R20729 vdd.n3381 vdd.n3380 19.3944
R20730 vdd.n3380 vdd.n380 19.3944
R20731 vdd.n3375 vdd.n380 19.3944
R20732 vdd.n3375 vdd.n3374 19.3944
R20733 vdd.n3210 vdd.n509 19.3944
R20734 vdd.n3222 vdd.n509 19.3944
R20735 vdd.n3222 vdd.n507 19.3944
R20736 vdd.n3226 vdd.n507 19.3944
R20737 vdd.n3226 vdd.n497 19.3944
R20738 vdd.n3238 vdd.n497 19.3944
R20739 vdd.n3238 vdd.n495 19.3944
R20740 vdd.n3242 vdd.n495 19.3944
R20741 vdd.n3242 vdd.n485 19.3944
R20742 vdd.n3255 vdd.n485 19.3944
R20743 vdd.n3255 vdd.n483 19.3944
R20744 vdd.n3259 vdd.n483 19.3944
R20745 vdd.n3259 vdd.n312 19.3944
R20746 vdd.n3438 vdd.n312 19.3944
R20747 vdd.n3438 vdd.n313 19.3944
R20748 vdd.n3432 vdd.n313 19.3944
R20749 vdd.n3432 vdd.n3431 19.3944
R20750 vdd.n3431 vdd.n3430 19.3944
R20751 vdd.n3430 vdd.n323 19.3944
R20752 vdd.n3424 vdd.n323 19.3944
R20753 vdd.n3424 vdd.n3423 19.3944
R20754 vdd.n3423 vdd.n3422 19.3944
R20755 vdd.n3422 vdd.n335 19.3944
R20756 vdd.n3416 vdd.n335 19.3944
R20757 vdd.n3416 vdd.n3415 19.3944
R20758 vdd.n3415 vdd.n3414 19.3944
R20759 vdd.n3414 vdd.n346 19.3944
R20760 vdd.n3408 vdd.n346 19.3944
R20761 vdd.n3167 vdd.n3166 19.3944
R20762 vdd.n3166 vdd.n3165 19.3944
R20763 vdd.n3165 vdd.n551 19.3944
R20764 vdd.n3159 vdd.n551 19.3944
R20765 vdd.n3159 vdd.n3158 19.3944
R20766 vdd.n3158 vdd.n3157 19.3944
R20767 vdd.n3157 vdd.n557 19.3944
R20768 vdd.n3151 vdd.n557 19.3944
R20769 vdd.n3151 vdd.n3150 19.3944
R20770 vdd.n3150 vdd.n3149 19.3944
R20771 vdd.n3149 vdd.n563 19.3944
R20772 vdd.n3143 vdd.n563 19.3944
R20773 vdd.n3143 vdd.n3142 19.3944
R20774 vdd.n3142 vdd.n3141 19.3944
R20775 vdd.n3141 vdd.n569 19.3944
R20776 vdd.n3135 vdd.n569 19.3944
R20777 vdd.n3135 vdd.n3134 19.3944
R20778 vdd.n3134 vdd.n3133 19.3944
R20779 vdd.n3133 vdd.n575 19.3944
R20780 vdd.n3127 vdd.n575 19.3944
R20781 vdd.n3207 vdd.n3206 19.3944
R20782 vdd.n3206 vdd.n519 19.3944
R20783 vdd.n3201 vdd.n3200 19.3944
R20784 vdd.n3197 vdd.n3196 19.3944
R20785 vdd.n3196 vdd.n525 19.3944
R20786 vdd.n3191 vdd.n525 19.3944
R20787 vdd.n3191 vdd.n3190 19.3944
R20788 vdd.n3190 vdd.n3189 19.3944
R20789 vdd.n3189 vdd.n531 19.3944
R20790 vdd.n3183 vdd.n531 19.3944
R20791 vdd.n3183 vdd.n3182 19.3944
R20792 vdd.n3182 vdd.n3181 19.3944
R20793 vdd.n3181 vdd.n537 19.3944
R20794 vdd.n3175 vdd.n537 19.3944
R20795 vdd.n3175 vdd.n3174 19.3944
R20796 vdd.n3174 vdd.n3173 19.3944
R20797 vdd.n3122 vdd.n579 19.3944
R20798 vdd.n3122 vdd.n583 19.3944
R20799 vdd.n3117 vdd.n583 19.3944
R20800 vdd.n3117 vdd.n3116 19.3944
R20801 vdd.n3116 vdd.n589 19.3944
R20802 vdd.n3111 vdd.n589 19.3944
R20803 vdd.n3111 vdd.n3110 19.3944
R20804 vdd.n3110 vdd.n3109 19.3944
R20805 vdd.n3109 vdd.n595 19.3944
R20806 vdd.n3103 vdd.n595 19.3944
R20807 vdd.n3103 vdd.n3102 19.3944
R20808 vdd.n3102 vdd.n3101 19.3944
R20809 vdd.n3101 vdd.n601 19.3944
R20810 vdd.n3095 vdd.n601 19.3944
R20811 vdd.n3095 vdd.n3094 19.3944
R20812 vdd.n3094 vdd.n3093 19.3944
R20813 vdd.n3089 vdd.n3088 19.3944
R20814 vdd.n3085 vdd.n3084 19.3944
R20815 vdd.n1604 vdd.n1523 19.0066
R20816 vdd.n2112 vdd.n1075 19.0066
R20817 vdd.n3334 vdd.n426 19.0066
R20818 vdd.n3126 vdd.n579 19.0066
R20819 vdd.n1144 vdd.n1143 16.0975
R20820 vdd.n839 vdd.n838 16.0975
R20821 vdd.n1566 vdd.n1565 16.0975
R20822 vdd.n1603 vdd.n1602 16.0975
R20823 vdd.n1477 vdd.n1476 16.0975
R20824 vdd.n2075 vdd.n2074 16.0975
R20825 vdd.n1077 vdd.n1076 16.0975
R20826 vdd.n1037 vdd.n1036 16.0975
R20827 vdd.n1148 vdd.n1147 16.0975
R20828 vdd.n830 vdd.n829 16.0975
R20829 vdd.n2536 vdd.n2535 16.0975
R20830 vdd.n3294 vdd.n3293 16.0975
R20831 vdd.n428 vdd.n427 16.0975
R20832 vdd.n388 vdd.n387 16.0975
R20833 vdd.n581 vdd.n580 16.0975
R20834 vdd.n544 vdd.n543 16.0975
R20835 vdd.n662 vdd.n661 16.0975
R20836 vdd.n2533 vdd.n2532 16.0975
R20837 vdd.n3081 vdd.n3080 16.0975
R20838 vdd.n626 vdd.n625 16.0975
R20839 vdd.t104 vdd.n2496 15.4182
R20840 vdd.n2800 vdd.t91 15.4182
R20841 vdd.n28 vdd.n27 14.5674
R20842 vdd.n304 vdd.n269 13.1884
R20843 vdd.n253 vdd.n218 13.1884
R20844 vdd.n210 vdd.n175 13.1884
R20845 vdd.n159 vdd.n124 13.1884
R20846 vdd.n117 vdd.n82 13.1884
R20847 vdd.n66 vdd.n31 13.1884
R20848 vdd.n1954 vdd.n1919 13.1884
R20849 vdd.n2005 vdd.n1970 13.1884
R20850 vdd.n1860 vdd.n1825 13.1884
R20851 vdd.n1911 vdd.n1876 13.1884
R20852 vdd.n1767 vdd.n1732 13.1884
R20853 vdd.n1818 vdd.n1783 13.1884
R20854 vdd.n2218 vdd.n962 13.1509
R20855 vdd.n3043 vdd.n613 13.1509
R20856 vdd.n1635 vdd.n1478 12.9944
R20857 vdd.n1639 vdd.n1478 12.9944
R20858 vdd.n2151 vdd.n1035 12.9944
R20859 vdd.n2152 vdd.n2151 12.9944
R20860 vdd.n3373 vdd.n386 12.9944
R20861 vdd.n3374 vdd.n3373 12.9944
R20862 vdd.n3167 vdd.n545 12.9944
R20863 vdd.n3173 vdd.n545 12.9944
R20864 vdd.n305 vdd.n267 12.8005
R20865 vdd.n300 vdd.n271 12.8005
R20866 vdd.n254 vdd.n216 12.8005
R20867 vdd.n249 vdd.n220 12.8005
R20868 vdd.n211 vdd.n173 12.8005
R20869 vdd.n206 vdd.n177 12.8005
R20870 vdd.n160 vdd.n122 12.8005
R20871 vdd.n155 vdd.n126 12.8005
R20872 vdd.n118 vdd.n80 12.8005
R20873 vdd.n113 vdd.n84 12.8005
R20874 vdd.n67 vdd.n29 12.8005
R20875 vdd.n62 vdd.n33 12.8005
R20876 vdd.n1955 vdd.n1917 12.8005
R20877 vdd.n1950 vdd.n1921 12.8005
R20878 vdd.n2006 vdd.n1968 12.8005
R20879 vdd.n2001 vdd.n1972 12.8005
R20880 vdd.n1861 vdd.n1823 12.8005
R20881 vdd.n1856 vdd.n1827 12.8005
R20882 vdd.n1912 vdd.n1874 12.8005
R20883 vdd.n1907 vdd.n1878 12.8005
R20884 vdd.n1768 vdd.n1730 12.8005
R20885 vdd.n1763 vdd.n1734 12.8005
R20886 vdd.n1819 vdd.n1781 12.8005
R20887 vdd.n1814 vdd.n1785 12.8005
R20888 vdd.n299 vdd.n272 12.0247
R20889 vdd.n248 vdd.n221 12.0247
R20890 vdd.n205 vdd.n178 12.0247
R20891 vdd.n154 vdd.n127 12.0247
R20892 vdd.n112 vdd.n85 12.0247
R20893 vdd.n61 vdd.n34 12.0247
R20894 vdd.n1949 vdd.n1922 12.0247
R20895 vdd.n2000 vdd.n1973 12.0247
R20896 vdd.n1855 vdd.n1828 12.0247
R20897 vdd.n1906 vdd.n1879 12.0247
R20898 vdd.n1762 vdd.n1735 12.0247
R20899 vdd.n1813 vdd.n1786 12.0247
R20900 vdd.n1670 vdd.n1438 11.337
R20901 vdd.n1678 vdd.n1427 11.337
R20902 vdd.n1686 vdd.n1427 11.337
R20903 vdd.n1694 vdd.n1421 11.337
R20904 vdd.n1702 vdd.n1414 11.337
R20905 vdd.n1711 vdd.n1710 11.337
R20906 vdd.n1719 vdd.n1403 11.337
R20907 vdd.n2017 vdd.n1392 11.337
R20908 vdd.n2026 vdd.n1386 11.337
R20909 vdd.n2034 vdd.n1380 11.337
R20910 vdd.n2043 vdd.n2042 11.337
R20911 vdd.n2051 vdd.n1363 11.337
R20912 vdd.n2062 vdd.n1363 11.337
R20913 vdd.n2062 vdd.n2061 11.337
R20914 vdd.n3220 vdd.n511 11.337
R20915 vdd.n3220 vdd.n505 11.337
R20916 vdd.n3228 vdd.n505 11.337
R20917 vdd.n3236 vdd.n499 11.337
R20918 vdd.n3244 vdd.n492 11.337
R20919 vdd.n3253 vdd.n3252 11.337
R20920 vdd.n3261 vdd.n481 11.337
R20921 vdd.n3435 vdd.n3434 11.337
R20922 vdd.n3428 vdd.n325 11.337
R20923 vdd.n3426 vdd.n329 11.337
R20924 vdd.n3420 vdd.n3419 11.337
R20925 vdd.n3418 vdd.n340 11.337
R20926 vdd.n3412 vdd.n340 11.337
R20927 vdd.n3411 vdd.n3410 11.337
R20928 vdd.n296 vdd.n295 11.249
R20929 vdd.n245 vdd.n244 11.249
R20930 vdd.n202 vdd.n201 11.249
R20931 vdd.n151 vdd.n150 11.249
R20932 vdd.n109 vdd.n108 11.249
R20933 vdd.n58 vdd.n57 11.249
R20934 vdd.n1946 vdd.n1945 11.249
R20935 vdd.n1997 vdd.n1996 11.249
R20936 vdd.n1852 vdd.n1851 11.249
R20937 vdd.n1903 vdd.n1902 11.249
R20938 vdd.n1759 vdd.n1758 11.249
R20939 vdd.n1810 vdd.n1809 11.249
R20940 vdd.n1686 vdd.t182 10.9969
R20941 vdd.t160 vdd.n3418 10.9969
R20942 vdd.n1415 vdd.t189 10.7702
R20943 vdd.t152 vdd.n3427 10.7702
R20944 vdd.n281 vdd.n280 10.7238
R20945 vdd.n230 vdd.n229 10.7238
R20946 vdd.n187 vdd.n186 10.7238
R20947 vdd.n136 vdd.n135 10.7238
R20948 vdd.n94 vdd.n93 10.7238
R20949 vdd.n43 vdd.n42 10.7238
R20950 vdd.n1931 vdd.n1930 10.7238
R20951 vdd.n1982 vdd.n1981 10.7238
R20952 vdd.n1837 vdd.n1836 10.7238
R20953 vdd.n1888 vdd.n1887 10.7238
R20954 vdd.n1744 vdd.n1743 10.7238
R20955 vdd.n1795 vdd.n1794 10.7238
R20956 vdd.n2223 vdd.n2222 10.6151
R20957 vdd.n2223 vdd.n955 10.6151
R20958 vdd.n2233 vdd.n955 10.6151
R20959 vdd.n2234 vdd.n2233 10.6151
R20960 vdd.n2235 vdd.n2234 10.6151
R20961 vdd.n2235 vdd.n942 10.6151
R20962 vdd.n2245 vdd.n942 10.6151
R20963 vdd.n2246 vdd.n2245 10.6151
R20964 vdd.n2247 vdd.n2246 10.6151
R20965 vdd.n2247 vdd.n930 10.6151
R20966 vdd.n2257 vdd.n930 10.6151
R20967 vdd.n2258 vdd.n2257 10.6151
R20968 vdd.n2259 vdd.n2258 10.6151
R20969 vdd.n2259 vdd.n919 10.6151
R20970 vdd.n2269 vdd.n919 10.6151
R20971 vdd.n2270 vdd.n2269 10.6151
R20972 vdd.n2271 vdd.n2270 10.6151
R20973 vdd.n2271 vdd.n906 10.6151
R20974 vdd.n2281 vdd.n906 10.6151
R20975 vdd.n2282 vdd.n2281 10.6151
R20976 vdd.n2283 vdd.n2282 10.6151
R20977 vdd.n2283 vdd.n894 10.6151
R20978 vdd.n2294 vdd.n894 10.6151
R20979 vdd.n2295 vdd.n2294 10.6151
R20980 vdd.n2296 vdd.n2295 10.6151
R20981 vdd.n2296 vdd.n882 10.6151
R20982 vdd.n2306 vdd.n882 10.6151
R20983 vdd.n2307 vdd.n2306 10.6151
R20984 vdd.n2308 vdd.n2307 10.6151
R20985 vdd.n2308 vdd.n870 10.6151
R20986 vdd.n2318 vdd.n870 10.6151
R20987 vdd.n2319 vdd.n2318 10.6151
R20988 vdd.n2320 vdd.n2319 10.6151
R20989 vdd.n2320 vdd.n860 10.6151
R20990 vdd.n2330 vdd.n860 10.6151
R20991 vdd.n2331 vdd.n2330 10.6151
R20992 vdd.n2332 vdd.n2331 10.6151
R20993 vdd.n2332 vdd.n847 10.6151
R20994 vdd.n2344 vdd.n847 10.6151
R20995 vdd.n2345 vdd.n2344 10.6151
R20996 vdd.n2347 vdd.n2345 10.6151
R20997 vdd.n2347 vdd.n2346 10.6151
R20998 vdd.n2346 vdd.n828 10.6151
R20999 vdd.n2494 vdd.n2493 10.6151
R21000 vdd.n2493 vdd.n2492 10.6151
R21001 vdd.n2492 vdd.n2489 10.6151
R21002 vdd.n2489 vdd.n2488 10.6151
R21003 vdd.n2488 vdd.n2485 10.6151
R21004 vdd.n2485 vdd.n2484 10.6151
R21005 vdd.n2484 vdd.n2481 10.6151
R21006 vdd.n2481 vdd.n2480 10.6151
R21007 vdd.n2480 vdd.n2477 10.6151
R21008 vdd.n2477 vdd.n2476 10.6151
R21009 vdd.n2476 vdd.n2473 10.6151
R21010 vdd.n2473 vdd.n2472 10.6151
R21011 vdd.n2472 vdd.n2469 10.6151
R21012 vdd.n2469 vdd.n2468 10.6151
R21013 vdd.n2468 vdd.n2465 10.6151
R21014 vdd.n2465 vdd.n2464 10.6151
R21015 vdd.n2464 vdd.n2461 10.6151
R21016 vdd.n2461 vdd.n2460 10.6151
R21017 vdd.n2460 vdd.n2457 10.6151
R21018 vdd.n2457 vdd.n2456 10.6151
R21019 vdd.n2456 vdd.n2453 10.6151
R21020 vdd.n2453 vdd.n2452 10.6151
R21021 vdd.n2452 vdd.n2449 10.6151
R21022 vdd.n2449 vdd.n2448 10.6151
R21023 vdd.n2448 vdd.n2445 10.6151
R21024 vdd.n2445 vdd.n2444 10.6151
R21025 vdd.n2444 vdd.n2441 10.6151
R21026 vdd.n2441 vdd.n2440 10.6151
R21027 vdd.n2440 vdd.n2437 10.6151
R21028 vdd.n2437 vdd.n2436 10.6151
R21029 vdd.n2436 vdd.n2433 10.6151
R21030 vdd.n2431 vdd.n2428 10.6151
R21031 vdd.n2428 vdd.n2427 10.6151
R21032 vdd.n1185 vdd.n1184 10.6151
R21033 vdd.n1187 vdd.n1185 10.6151
R21034 vdd.n1188 vdd.n1187 10.6151
R21035 vdd.n1190 vdd.n1188 10.6151
R21036 vdd.n1191 vdd.n1190 10.6151
R21037 vdd.n1193 vdd.n1191 10.6151
R21038 vdd.n1194 vdd.n1193 10.6151
R21039 vdd.n1196 vdd.n1194 10.6151
R21040 vdd.n1197 vdd.n1196 10.6151
R21041 vdd.n1199 vdd.n1197 10.6151
R21042 vdd.n1200 vdd.n1199 10.6151
R21043 vdd.n1202 vdd.n1200 10.6151
R21044 vdd.n1203 vdd.n1202 10.6151
R21045 vdd.n1205 vdd.n1203 10.6151
R21046 vdd.n1206 vdd.n1205 10.6151
R21047 vdd.n1208 vdd.n1206 10.6151
R21048 vdd.n1209 vdd.n1208 10.6151
R21049 vdd.n1211 vdd.n1209 10.6151
R21050 vdd.n1212 vdd.n1211 10.6151
R21051 vdd.n1214 vdd.n1212 10.6151
R21052 vdd.n1215 vdd.n1214 10.6151
R21053 vdd.n1217 vdd.n1215 10.6151
R21054 vdd.n1218 vdd.n1217 10.6151
R21055 vdd.n1220 vdd.n1218 10.6151
R21056 vdd.n1221 vdd.n1220 10.6151
R21057 vdd.n1223 vdd.n1221 10.6151
R21058 vdd.n1224 vdd.n1223 10.6151
R21059 vdd.n1263 vdd.n1224 10.6151
R21060 vdd.n1263 vdd.n1262 10.6151
R21061 vdd.n1262 vdd.n1261 10.6151
R21062 vdd.n1261 vdd.n1259 10.6151
R21063 vdd.n1259 vdd.n1258 10.6151
R21064 vdd.n1258 vdd.n1256 10.6151
R21065 vdd.n1256 vdd.n1255 10.6151
R21066 vdd.n1255 vdd.n1236 10.6151
R21067 vdd.n1236 vdd.n1235 10.6151
R21068 vdd.n1235 vdd.n1233 10.6151
R21069 vdd.n1233 vdd.n1232 10.6151
R21070 vdd.n1232 vdd.n1230 10.6151
R21071 vdd.n1230 vdd.n1229 10.6151
R21072 vdd.n1229 vdd.n1226 10.6151
R21073 vdd.n1226 vdd.n1225 10.6151
R21074 vdd.n1225 vdd.n831 10.6151
R21075 vdd.n2221 vdd.n967 10.6151
R21076 vdd.n2216 vdd.n967 10.6151
R21077 vdd.n2216 vdd.n2215 10.6151
R21078 vdd.n2215 vdd.n2214 10.6151
R21079 vdd.n2214 vdd.n2211 10.6151
R21080 vdd.n2211 vdd.n2210 10.6151
R21081 vdd.n2210 vdd.n2207 10.6151
R21082 vdd.n2207 vdd.n2206 10.6151
R21083 vdd.n2206 vdd.n2203 10.6151
R21084 vdd.n2203 vdd.n2202 10.6151
R21085 vdd.n2202 vdd.n2199 10.6151
R21086 vdd.n2199 vdd.n2198 10.6151
R21087 vdd.n2198 vdd.n2195 10.6151
R21088 vdd.n2195 vdd.n2194 10.6151
R21089 vdd.n2194 vdd.n2191 10.6151
R21090 vdd.n2191 vdd.n2190 10.6151
R21091 vdd.n2190 vdd.n2187 10.6151
R21092 vdd.n2187 vdd.n1005 10.6151
R21093 vdd.n1151 vdd.n1005 10.6151
R21094 vdd.n1152 vdd.n1151 10.6151
R21095 vdd.n1155 vdd.n1152 10.6151
R21096 vdd.n1156 vdd.n1155 10.6151
R21097 vdd.n1159 vdd.n1156 10.6151
R21098 vdd.n1160 vdd.n1159 10.6151
R21099 vdd.n1163 vdd.n1160 10.6151
R21100 vdd.n1164 vdd.n1163 10.6151
R21101 vdd.n1167 vdd.n1164 10.6151
R21102 vdd.n1168 vdd.n1167 10.6151
R21103 vdd.n1171 vdd.n1168 10.6151
R21104 vdd.n1172 vdd.n1171 10.6151
R21105 vdd.n1175 vdd.n1172 10.6151
R21106 vdd.n1180 vdd.n1177 10.6151
R21107 vdd.n1181 vdd.n1180 10.6151
R21108 vdd.n2732 vdd.n2731 10.6151
R21109 vdd.n2731 vdd.n2730 10.6151
R21110 vdd.n2730 vdd.n2534 10.6151
R21111 vdd.n2612 vdd.n2534 10.6151
R21112 vdd.n2613 vdd.n2612 10.6151
R21113 vdd.n2615 vdd.n2613 10.6151
R21114 vdd.n2616 vdd.n2615 10.6151
R21115 vdd.n2714 vdd.n2616 10.6151
R21116 vdd.n2714 vdd.n2713 10.6151
R21117 vdd.n2713 vdd.n2712 10.6151
R21118 vdd.n2712 vdd.n2660 10.6151
R21119 vdd.n2660 vdd.n2659 10.6151
R21120 vdd.n2659 vdd.n2657 10.6151
R21121 vdd.n2657 vdd.n2656 10.6151
R21122 vdd.n2656 vdd.n2654 10.6151
R21123 vdd.n2654 vdd.n2653 10.6151
R21124 vdd.n2653 vdd.n2651 10.6151
R21125 vdd.n2651 vdd.n2650 10.6151
R21126 vdd.n2650 vdd.n2648 10.6151
R21127 vdd.n2648 vdd.n2647 10.6151
R21128 vdd.n2647 vdd.n2645 10.6151
R21129 vdd.n2645 vdd.n2644 10.6151
R21130 vdd.n2644 vdd.n2642 10.6151
R21131 vdd.n2642 vdd.n2641 10.6151
R21132 vdd.n2641 vdd.n2639 10.6151
R21133 vdd.n2639 vdd.n2638 10.6151
R21134 vdd.n2638 vdd.n2636 10.6151
R21135 vdd.n2636 vdd.n2635 10.6151
R21136 vdd.n2635 vdd.n2633 10.6151
R21137 vdd.n2633 vdd.n2632 10.6151
R21138 vdd.n2632 vdd.n2630 10.6151
R21139 vdd.n2630 vdd.n2629 10.6151
R21140 vdd.n2629 vdd.n2627 10.6151
R21141 vdd.n2627 vdd.n2626 10.6151
R21142 vdd.n2626 vdd.n2624 10.6151
R21143 vdd.n2624 vdd.n2623 10.6151
R21144 vdd.n2623 vdd.n2621 10.6151
R21145 vdd.n2621 vdd.n2620 10.6151
R21146 vdd.n2620 vdd.n2618 10.6151
R21147 vdd.n2618 vdd.n2617 10.6151
R21148 vdd.n2617 vdd.n664 10.6151
R21149 vdd.n2976 vdd.n664 10.6151
R21150 vdd.n2977 vdd.n2976 10.6151
R21151 vdd.n2803 vdd.n789 10.6151
R21152 vdd.n2798 vdd.n789 10.6151
R21153 vdd.n2798 vdd.n2797 10.6151
R21154 vdd.n2797 vdd.n2796 10.6151
R21155 vdd.n2796 vdd.n2793 10.6151
R21156 vdd.n2793 vdd.n2792 10.6151
R21157 vdd.n2792 vdd.n2789 10.6151
R21158 vdd.n2789 vdd.n2788 10.6151
R21159 vdd.n2788 vdd.n2785 10.6151
R21160 vdd.n2785 vdd.n2784 10.6151
R21161 vdd.n2784 vdd.n2781 10.6151
R21162 vdd.n2781 vdd.n2780 10.6151
R21163 vdd.n2780 vdd.n2777 10.6151
R21164 vdd.n2777 vdd.n2776 10.6151
R21165 vdd.n2776 vdd.n2773 10.6151
R21166 vdd.n2773 vdd.n2772 10.6151
R21167 vdd.n2772 vdd.n2769 10.6151
R21168 vdd.n2769 vdd.n2768 10.6151
R21169 vdd.n2768 vdd.n2765 10.6151
R21170 vdd.n2765 vdd.n2764 10.6151
R21171 vdd.n2764 vdd.n2761 10.6151
R21172 vdd.n2761 vdd.n2760 10.6151
R21173 vdd.n2760 vdd.n2757 10.6151
R21174 vdd.n2757 vdd.n2756 10.6151
R21175 vdd.n2756 vdd.n2753 10.6151
R21176 vdd.n2753 vdd.n2752 10.6151
R21177 vdd.n2752 vdd.n2749 10.6151
R21178 vdd.n2749 vdd.n2748 10.6151
R21179 vdd.n2748 vdd.n2745 10.6151
R21180 vdd.n2745 vdd.n2744 10.6151
R21181 vdd.n2744 vdd.n2741 10.6151
R21182 vdd.n2739 vdd.n2736 10.6151
R21183 vdd.n2736 vdd.n2735 10.6151
R21184 vdd.n2805 vdd.n2804 10.6151
R21185 vdd.n2805 vdd.n778 10.6151
R21186 vdd.n2815 vdd.n778 10.6151
R21187 vdd.n2816 vdd.n2815 10.6151
R21188 vdd.n2817 vdd.n2816 10.6151
R21189 vdd.n2817 vdd.n766 10.6151
R21190 vdd.n2827 vdd.n766 10.6151
R21191 vdd.n2828 vdd.n2827 10.6151
R21192 vdd.n2829 vdd.n2828 10.6151
R21193 vdd.n2829 vdd.n755 10.6151
R21194 vdd.n2839 vdd.n755 10.6151
R21195 vdd.n2840 vdd.n2839 10.6151
R21196 vdd.n2841 vdd.n2840 10.6151
R21197 vdd.n2841 vdd.n744 10.6151
R21198 vdd.n2851 vdd.n744 10.6151
R21199 vdd.n2852 vdd.n2851 10.6151
R21200 vdd.n2853 vdd.n2852 10.6151
R21201 vdd.n2853 vdd.n731 10.6151
R21202 vdd.n2864 vdd.n731 10.6151
R21203 vdd.n2865 vdd.n2864 10.6151
R21204 vdd.n2866 vdd.n2865 10.6151
R21205 vdd.n2866 vdd.n719 10.6151
R21206 vdd.n2876 vdd.n719 10.6151
R21207 vdd.n2877 vdd.n2876 10.6151
R21208 vdd.n2878 vdd.n2877 10.6151
R21209 vdd.n2878 vdd.n707 10.6151
R21210 vdd.n2888 vdd.n707 10.6151
R21211 vdd.n2889 vdd.n2888 10.6151
R21212 vdd.n2890 vdd.n2889 10.6151
R21213 vdd.n2890 vdd.n694 10.6151
R21214 vdd.n2900 vdd.n694 10.6151
R21215 vdd.n2901 vdd.n2900 10.6151
R21216 vdd.n2902 vdd.n2901 10.6151
R21217 vdd.n2902 vdd.n683 10.6151
R21218 vdd.n2912 vdd.n683 10.6151
R21219 vdd.n2913 vdd.n2912 10.6151
R21220 vdd.n2914 vdd.n2913 10.6151
R21221 vdd.n2914 vdd.n669 10.6151
R21222 vdd.n2969 vdd.n669 10.6151
R21223 vdd.n2970 vdd.n2969 10.6151
R21224 vdd.n2971 vdd.n2970 10.6151
R21225 vdd.n2971 vdd.n636 10.6151
R21226 vdd.n3041 vdd.n636 10.6151
R21227 vdd.n3040 vdd.n3039 10.6151
R21228 vdd.n3039 vdd.n637 10.6151
R21229 vdd.n638 vdd.n637 10.6151
R21230 vdd.n3032 vdd.n638 10.6151
R21231 vdd.n3032 vdd.n3031 10.6151
R21232 vdd.n3031 vdd.n3030 10.6151
R21233 vdd.n3030 vdd.n640 10.6151
R21234 vdd.n3025 vdd.n640 10.6151
R21235 vdd.n3025 vdd.n3024 10.6151
R21236 vdd.n3024 vdd.n3023 10.6151
R21237 vdd.n3023 vdd.n643 10.6151
R21238 vdd.n3018 vdd.n643 10.6151
R21239 vdd.n3018 vdd.n3017 10.6151
R21240 vdd.n3017 vdd.n3016 10.6151
R21241 vdd.n3016 vdd.n646 10.6151
R21242 vdd.n3011 vdd.n646 10.6151
R21243 vdd.n3011 vdd.n3010 10.6151
R21244 vdd.n3010 vdd.n3008 10.6151
R21245 vdd.n3008 vdd.n649 10.6151
R21246 vdd.n3003 vdd.n649 10.6151
R21247 vdd.n3003 vdd.n3002 10.6151
R21248 vdd.n3002 vdd.n3001 10.6151
R21249 vdd.n3001 vdd.n652 10.6151
R21250 vdd.n2996 vdd.n652 10.6151
R21251 vdd.n2996 vdd.n2995 10.6151
R21252 vdd.n2995 vdd.n2994 10.6151
R21253 vdd.n2994 vdd.n655 10.6151
R21254 vdd.n2989 vdd.n655 10.6151
R21255 vdd.n2989 vdd.n2988 10.6151
R21256 vdd.n2988 vdd.n2987 10.6151
R21257 vdd.n2987 vdd.n658 10.6151
R21258 vdd.n2982 vdd.n2981 10.6151
R21259 vdd.n2981 vdd.n2980 10.6151
R21260 vdd.n2959 vdd.n2920 10.6151
R21261 vdd.n2954 vdd.n2920 10.6151
R21262 vdd.n2954 vdd.n2953 10.6151
R21263 vdd.n2953 vdd.n2952 10.6151
R21264 vdd.n2952 vdd.n2922 10.6151
R21265 vdd.n2947 vdd.n2922 10.6151
R21266 vdd.n2947 vdd.n2946 10.6151
R21267 vdd.n2946 vdd.n2945 10.6151
R21268 vdd.n2945 vdd.n2925 10.6151
R21269 vdd.n2940 vdd.n2925 10.6151
R21270 vdd.n2940 vdd.n2939 10.6151
R21271 vdd.n2939 vdd.n2938 10.6151
R21272 vdd.n2938 vdd.n2928 10.6151
R21273 vdd.n2933 vdd.n2928 10.6151
R21274 vdd.n2933 vdd.n2932 10.6151
R21275 vdd.n2932 vdd.n610 10.6151
R21276 vdd.n3076 vdd.n610 10.6151
R21277 vdd.n3076 vdd.n611 10.6151
R21278 vdd.n614 vdd.n611 10.6151
R21279 vdd.n3069 vdd.n614 10.6151
R21280 vdd.n3069 vdd.n3068 10.6151
R21281 vdd.n3068 vdd.n3067 10.6151
R21282 vdd.n3067 vdd.n616 10.6151
R21283 vdd.n3062 vdd.n616 10.6151
R21284 vdd.n3062 vdd.n3061 10.6151
R21285 vdd.n3061 vdd.n3060 10.6151
R21286 vdd.n3060 vdd.n619 10.6151
R21287 vdd.n3055 vdd.n619 10.6151
R21288 vdd.n3055 vdd.n3054 10.6151
R21289 vdd.n3054 vdd.n3053 10.6151
R21290 vdd.n3053 vdd.n622 10.6151
R21291 vdd.n3048 vdd.n3047 10.6151
R21292 vdd.n3047 vdd.n3046 10.6151
R21293 vdd.n2609 vdd.n2608 10.6151
R21294 vdd.n2726 vdd.n2609 10.6151
R21295 vdd.n2726 vdd.n2725 10.6151
R21296 vdd.n2725 vdd.n2724 10.6151
R21297 vdd.n2724 vdd.n2722 10.6151
R21298 vdd.n2722 vdd.n2721 10.6151
R21299 vdd.n2721 vdd.n2719 10.6151
R21300 vdd.n2719 vdd.n2718 10.6151
R21301 vdd.n2718 vdd.n2610 10.6151
R21302 vdd.n2708 vdd.n2610 10.6151
R21303 vdd.n2708 vdd.n2707 10.6151
R21304 vdd.n2707 vdd.n2706 10.6151
R21305 vdd.n2706 vdd.n2704 10.6151
R21306 vdd.n2704 vdd.n2703 10.6151
R21307 vdd.n2703 vdd.n2701 10.6151
R21308 vdd.n2701 vdd.n2700 10.6151
R21309 vdd.n2700 vdd.n2698 10.6151
R21310 vdd.n2698 vdd.n2697 10.6151
R21311 vdd.n2697 vdd.n2695 10.6151
R21312 vdd.n2695 vdd.n2694 10.6151
R21313 vdd.n2694 vdd.n2692 10.6151
R21314 vdd.n2692 vdd.n2691 10.6151
R21315 vdd.n2691 vdd.n2689 10.6151
R21316 vdd.n2689 vdd.n2688 10.6151
R21317 vdd.n2688 vdd.n2686 10.6151
R21318 vdd.n2686 vdd.n2685 10.6151
R21319 vdd.n2685 vdd.n2683 10.6151
R21320 vdd.n2683 vdd.n2682 10.6151
R21321 vdd.n2682 vdd.n2680 10.6151
R21322 vdd.n2680 vdd.n2679 10.6151
R21323 vdd.n2679 vdd.n2677 10.6151
R21324 vdd.n2677 vdd.n2676 10.6151
R21325 vdd.n2676 vdd.n2674 10.6151
R21326 vdd.n2674 vdd.n2673 10.6151
R21327 vdd.n2673 vdd.n2671 10.6151
R21328 vdd.n2671 vdd.n2670 10.6151
R21329 vdd.n2670 vdd.n2668 10.6151
R21330 vdd.n2668 vdd.n2667 10.6151
R21331 vdd.n2667 vdd.n2665 10.6151
R21332 vdd.n2665 vdd.n2664 10.6151
R21333 vdd.n2664 vdd.n2662 10.6151
R21334 vdd.n2662 vdd.n2661 10.6151
R21335 vdd.n2661 vdd.n628 10.6151
R21336 vdd.n2540 vdd.n2539 10.6151
R21337 vdd.n2543 vdd.n2540 10.6151
R21338 vdd.n2544 vdd.n2543 10.6151
R21339 vdd.n2547 vdd.n2544 10.6151
R21340 vdd.n2548 vdd.n2547 10.6151
R21341 vdd.n2551 vdd.n2548 10.6151
R21342 vdd.n2552 vdd.n2551 10.6151
R21343 vdd.n2555 vdd.n2552 10.6151
R21344 vdd.n2556 vdd.n2555 10.6151
R21345 vdd.n2559 vdd.n2556 10.6151
R21346 vdd.n2560 vdd.n2559 10.6151
R21347 vdd.n2563 vdd.n2560 10.6151
R21348 vdd.n2564 vdd.n2563 10.6151
R21349 vdd.n2567 vdd.n2564 10.6151
R21350 vdd.n2568 vdd.n2567 10.6151
R21351 vdd.n2571 vdd.n2568 10.6151
R21352 vdd.n2572 vdd.n2571 10.6151
R21353 vdd.n2575 vdd.n2572 10.6151
R21354 vdd.n2576 vdd.n2575 10.6151
R21355 vdd.n2579 vdd.n2576 10.6151
R21356 vdd.n2580 vdd.n2579 10.6151
R21357 vdd.n2583 vdd.n2580 10.6151
R21358 vdd.n2584 vdd.n2583 10.6151
R21359 vdd.n2587 vdd.n2584 10.6151
R21360 vdd.n2588 vdd.n2587 10.6151
R21361 vdd.n2591 vdd.n2588 10.6151
R21362 vdd.n2592 vdd.n2591 10.6151
R21363 vdd.n2595 vdd.n2592 10.6151
R21364 vdd.n2596 vdd.n2595 10.6151
R21365 vdd.n2599 vdd.n2596 10.6151
R21366 vdd.n2600 vdd.n2599 10.6151
R21367 vdd.n2605 vdd.n2603 10.6151
R21368 vdd.n2606 vdd.n2605 10.6151
R21369 vdd.n2809 vdd.n783 10.6151
R21370 vdd.n2810 vdd.n2809 10.6151
R21371 vdd.n2811 vdd.n2810 10.6151
R21372 vdd.n2811 vdd.n772 10.6151
R21373 vdd.n2821 vdd.n772 10.6151
R21374 vdd.n2822 vdd.n2821 10.6151
R21375 vdd.n2823 vdd.n2822 10.6151
R21376 vdd.n2823 vdd.n761 10.6151
R21377 vdd.n2833 vdd.n761 10.6151
R21378 vdd.n2834 vdd.n2833 10.6151
R21379 vdd.n2835 vdd.n2834 10.6151
R21380 vdd.n2835 vdd.n749 10.6151
R21381 vdd.n2845 vdd.n749 10.6151
R21382 vdd.n2846 vdd.n2845 10.6151
R21383 vdd.n2847 vdd.n2846 10.6151
R21384 vdd.n2847 vdd.n738 10.6151
R21385 vdd.n2857 vdd.n738 10.6151
R21386 vdd.n2858 vdd.n2857 10.6151
R21387 vdd.n2860 vdd.n2858 10.6151
R21388 vdd.n2860 vdd.n2859 10.6151
R21389 vdd.n2871 vdd.n2870 10.6151
R21390 vdd.n2872 vdd.n2871 10.6151
R21391 vdd.n2872 vdd.n713 10.6151
R21392 vdd.n2882 vdd.n713 10.6151
R21393 vdd.n2883 vdd.n2882 10.6151
R21394 vdd.n2884 vdd.n2883 10.6151
R21395 vdd.n2884 vdd.n700 10.6151
R21396 vdd.n2894 vdd.n700 10.6151
R21397 vdd.n2895 vdd.n2894 10.6151
R21398 vdd.n2896 vdd.n2895 10.6151
R21399 vdd.n2896 vdd.n688 10.6151
R21400 vdd.n2906 vdd.n688 10.6151
R21401 vdd.n2907 vdd.n2906 10.6151
R21402 vdd.n2908 vdd.n2907 10.6151
R21403 vdd.n2908 vdd.n677 10.6151
R21404 vdd.n2918 vdd.n677 10.6151
R21405 vdd.n2919 vdd.n2918 10.6151
R21406 vdd.n2965 vdd.n2919 10.6151
R21407 vdd.n2965 vdd.n2964 10.6151
R21408 vdd.n2964 vdd.n2963 10.6151
R21409 vdd.n2963 vdd.n2962 10.6151
R21410 vdd.n2962 vdd.n2960 10.6151
R21411 vdd.n2227 vdd.n960 10.6151
R21412 vdd.n2228 vdd.n2227 10.6151
R21413 vdd.n2229 vdd.n2228 10.6151
R21414 vdd.n2229 vdd.n949 10.6151
R21415 vdd.n2239 vdd.n949 10.6151
R21416 vdd.n2240 vdd.n2239 10.6151
R21417 vdd.n2241 vdd.n2240 10.6151
R21418 vdd.n2241 vdd.n936 10.6151
R21419 vdd.n2251 vdd.n936 10.6151
R21420 vdd.n2252 vdd.n2251 10.6151
R21421 vdd.n2253 vdd.n2252 10.6151
R21422 vdd.n2253 vdd.n925 10.6151
R21423 vdd.n2263 vdd.n925 10.6151
R21424 vdd.n2264 vdd.n2263 10.6151
R21425 vdd.n2265 vdd.n2264 10.6151
R21426 vdd.n2265 vdd.n913 10.6151
R21427 vdd.n2275 vdd.n913 10.6151
R21428 vdd.n2276 vdd.n2275 10.6151
R21429 vdd.n2277 vdd.n2276 10.6151
R21430 vdd.n2277 vdd.n900 10.6151
R21431 vdd.n2287 vdd.n900 10.6151
R21432 vdd.n2288 vdd.n2287 10.6151
R21433 vdd.n2290 vdd.n888 10.6151
R21434 vdd.n2300 vdd.n888 10.6151
R21435 vdd.n2301 vdd.n2300 10.6151
R21436 vdd.n2302 vdd.n2301 10.6151
R21437 vdd.n2302 vdd.n876 10.6151
R21438 vdd.n2312 vdd.n876 10.6151
R21439 vdd.n2313 vdd.n2312 10.6151
R21440 vdd.n2314 vdd.n2313 10.6151
R21441 vdd.n2314 vdd.n865 10.6151
R21442 vdd.n2324 vdd.n865 10.6151
R21443 vdd.n2325 vdd.n2324 10.6151
R21444 vdd.n2326 vdd.n2325 10.6151
R21445 vdd.n2326 vdd.n854 10.6151
R21446 vdd.n2336 vdd.n854 10.6151
R21447 vdd.n2337 vdd.n2336 10.6151
R21448 vdd.n2340 vdd.n2337 10.6151
R21449 vdd.n2340 vdd.n2339 10.6151
R21450 vdd.n2339 vdd.n2338 10.6151
R21451 vdd.n2338 vdd.n837 10.6151
R21452 vdd.n2422 vdd.n837 10.6151
R21453 vdd.n2421 vdd.n2420 10.6151
R21454 vdd.n2420 vdd.n2417 10.6151
R21455 vdd.n2417 vdd.n2416 10.6151
R21456 vdd.n2416 vdd.n2413 10.6151
R21457 vdd.n2413 vdd.n2412 10.6151
R21458 vdd.n2412 vdd.n2409 10.6151
R21459 vdd.n2409 vdd.n2408 10.6151
R21460 vdd.n2408 vdd.n2405 10.6151
R21461 vdd.n2405 vdd.n2404 10.6151
R21462 vdd.n2404 vdd.n2401 10.6151
R21463 vdd.n2401 vdd.n2400 10.6151
R21464 vdd.n2400 vdd.n2397 10.6151
R21465 vdd.n2397 vdd.n2396 10.6151
R21466 vdd.n2396 vdd.n2393 10.6151
R21467 vdd.n2393 vdd.n2392 10.6151
R21468 vdd.n2392 vdd.n2389 10.6151
R21469 vdd.n2389 vdd.n2388 10.6151
R21470 vdd.n2388 vdd.n2385 10.6151
R21471 vdd.n2385 vdd.n2384 10.6151
R21472 vdd.n2384 vdd.n2381 10.6151
R21473 vdd.n2381 vdd.n2380 10.6151
R21474 vdd.n2380 vdd.n2377 10.6151
R21475 vdd.n2377 vdd.n2376 10.6151
R21476 vdd.n2376 vdd.n2373 10.6151
R21477 vdd.n2373 vdd.n2372 10.6151
R21478 vdd.n2372 vdd.n2369 10.6151
R21479 vdd.n2369 vdd.n2368 10.6151
R21480 vdd.n2368 vdd.n2365 10.6151
R21481 vdd.n2365 vdd.n2364 10.6151
R21482 vdd.n2364 vdd.n2361 10.6151
R21483 vdd.n2361 vdd.n2360 10.6151
R21484 vdd.n2357 vdd.n2356 10.6151
R21485 vdd.n2356 vdd.n2354 10.6151
R21486 vdd.n1309 vdd.n1307 10.6151
R21487 vdd.n1307 vdd.n1306 10.6151
R21488 vdd.n1306 vdd.n1304 10.6151
R21489 vdd.n1304 vdd.n1303 10.6151
R21490 vdd.n1303 vdd.n1301 10.6151
R21491 vdd.n1301 vdd.n1300 10.6151
R21492 vdd.n1300 vdd.n1298 10.6151
R21493 vdd.n1298 vdd.n1297 10.6151
R21494 vdd.n1297 vdd.n1295 10.6151
R21495 vdd.n1295 vdd.n1294 10.6151
R21496 vdd.n1294 vdd.n1292 10.6151
R21497 vdd.n1292 vdd.n1291 10.6151
R21498 vdd.n1291 vdd.n1289 10.6151
R21499 vdd.n1289 vdd.n1288 10.6151
R21500 vdd.n1288 vdd.n1286 10.6151
R21501 vdd.n1286 vdd.n1285 10.6151
R21502 vdd.n1285 vdd.n1283 10.6151
R21503 vdd.n1283 vdd.n1282 10.6151
R21504 vdd.n1282 vdd.n1280 10.6151
R21505 vdd.n1280 vdd.n1279 10.6151
R21506 vdd.n1279 vdd.n1277 10.6151
R21507 vdd.n1277 vdd.n1276 10.6151
R21508 vdd.n1276 vdd.n1274 10.6151
R21509 vdd.n1274 vdd.n1273 10.6151
R21510 vdd.n1273 vdd.n1271 10.6151
R21511 vdd.n1271 vdd.n1270 10.6151
R21512 vdd.n1270 vdd.n1268 10.6151
R21513 vdd.n1268 vdd.n1267 10.6151
R21514 vdd.n1267 vdd.n1146 10.6151
R21515 vdd.n1238 vdd.n1146 10.6151
R21516 vdd.n1239 vdd.n1238 10.6151
R21517 vdd.n1241 vdd.n1239 10.6151
R21518 vdd.n1242 vdd.n1241 10.6151
R21519 vdd.n1251 vdd.n1242 10.6151
R21520 vdd.n1251 vdd.n1250 10.6151
R21521 vdd.n1250 vdd.n1249 10.6151
R21522 vdd.n1249 vdd.n1247 10.6151
R21523 vdd.n1247 vdd.n1246 10.6151
R21524 vdd.n1246 vdd.n1244 10.6151
R21525 vdd.n1244 vdd.n1243 10.6151
R21526 vdd.n1243 vdd.n841 10.6151
R21527 vdd.n2352 vdd.n841 10.6151
R21528 vdd.n2353 vdd.n2352 10.6151
R21529 vdd.n1110 vdd.n1109 10.6151
R21530 vdd.n1113 vdd.n1110 10.6151
R21531 vdd.n1114 vdd.n1113 10.6151
R21532 vdd.n1117 vdd.n1114 10.6151
R21533 vdd.n1118 vdd.n1117 10.6151
R21534 vdd.n1121 vdd.n1118 10.6151
R21535 vdd.n1122 vdd.n1121 10.6151
R21536 vdd.n1125 vdd.n1122 10.6151
R21537 vdd.n1126 vdd.n1125 10.6151
R21538 vdd.n1129 vdd.n1126 10.6151
R21539 vdd.n1130 vdd.n1129 10.6151
R21540 vdd.n1133 vdd.n1130 10.6151
R21541 vdd.n1134 vdd.n1133 10.6151
R21542 vdd.n1137 vdd.n1134 10.6151
R21543 vdd.n1138 vdd.n1137 10.6151
R21544 vdd.n1141 vdd.n1138 10.6151
R21545 vdd.n1343 vdd.n1141 10.6151
R21546 vdd.n1343 vdd.n1342 10.6151
R21547 vdd.n1342 vdd.n1340 10.6151
R21548 vdd.n1340 vdd.n1337 10.6151
R21549 vdd.n1337 vdd.n1336 10.6151
R21550 vdd.n1336 vdd.n1333 10.6151
R21551 vdd.n1333 vdd.n1332 10.6151
R21552 vdd.n1332 vdd.n1329 10.6151
R21553 vdd.n1329 vdd.n1328 10.6151
R21554 vdd.n1328 vdd.n1325 10.6151
R21555 vdd.n1325 vdd.n1324 10.6151
R21556 vdd.n1324 vdd.n1321 10.6151
R21557 vdd.n1321 vdd.n1320 10.6151
R21558 vdd.n1320 vdd.n1317 10.6151
R21559 vdd.n1317 vdd.n1316 10.6151
R21560 vdd.n1313 vdd.n1312 10.6151
R21561 vdd.n1312 vdd.n1310 10.6151
R21562 vdd.n1727 vdd.t175 10.5435
R21563 vdd.n2070 vdd.t9 10.5435
R21564 vdd.n3212 vdd.t19 10.5435
R21565 vdd.n3436 vdd.t158 10.5435
R21566 vdd.n292 vdd.n274 10.4732
R21567 vdd.n241 vdd.n223 10.4732
R21568 vdd.n198 vdd.n180 10.4732
R21569 vdd.n147 vdd.n129 10.4732
R21570 vdd.n105 vdd.n87 10.4732
R21571 vdd.n54 vdd.n36 10.4732
R21572 vdd.n1942 vdd.n1924 10.4732
R21573 vdd.n1993 vdd.n1975 10.4732
R21574 vdd.n1848 vdd.n1830 10.4732
R21575 vdd.n1899 vdd.n1881 10.4732
R21576 vdd.n1755 vdd.n1737 10.4732
R21577 vdd.n1806 vdd.n1788 10.4732
R21578 vdd.n2025 vdd.t209 10.3167
R21579 vdd.t162 vdd.n493 10.3167
R21580 vdd.n2187 vdd.n2186 9.98956
R21581 vdd.n3010 vdd.n3009 9.98956
R21582 vdd.n3077 vdd.n3076 9.98956
R21583 vdd.n2079 vdd.n1343 9.98956
R21584 vdd.n1678 vdd.t37 9.86327
R21585 vdd.n3412 vdd.t23 9.86327
R21586 vdd.n2424 vdd.t124 9.7499
R21587 vdd.t109 vdd.n785 9.7499
R21588 vdd.n291 vdd.n276 9.69747
R21589 vdd.n240 vdd.n225 9.69747
R21590 vdd.n197 vdd.n182 9.69747
R21591 vdd.n146 vdd.n131 9.69747
R21592 vdd.n104 vdd.n89 9.69747
R21593 vdd.n53 vdd.n38 9.69747
R21594 vdd.n1941 vdd.n1926 9.69747
R21595 vdd.n1992 vdd.n1977 9.69747
R21596 vdd.n1847 vdd.n1832 9.69747
R21597 vdd.n1898 vdd.n1883 9.69747
R21598 vdd.n1754 vdd.n1739 9.69747
R21599 vdd.n1805 vdd.n1790 9.69747
R21600 vdd.n307 vdd.n306 9.45567
R21601 vdd.n256 vdd.n255 9.45567
R21602 vdd.n213 vdd.n212 9.45567
R21603 vdd.n162 vdd.n161 9.45567
R21604 vdd.n120 vdd.n119 9.45567
R21605 vdd.n69 vdd.n68 9.45567
R21606 vdd.n1957 vdd.n1956 9.45567
R21607 vdd.n2008 vdd.n2007 9.45567
R21608 vdd.n1863 vdd.n1862 9.45567
R21609 vdd.n1914 vdd.n1913 9.45567
R21610 vdd.n1770 vdd.n1769 9.45567
R21611 vdd.n1821 vdd.n1820 9.45567
R21612 vdd.n2149 vdd.n1035 9.3005
R21613 vdd.n2148 vdd.n2147 9.3005
R21614 vdd.n1041 vdd.n1040 9.3005
R21615 vdd.n2142 vdd.n1045 9.3005
R21616 vdd.n2141 vdd.n1046 9.3005
R21617 vdd.n2140 vdd.n1047 9.3005
R21618 vdd.n1051 vdd.n1048 9.3005
R21619 vdd.n2135 vdd.n1052 9.3005
R21620 vdd.n2134 vdd.n1053 9.3005
R21621 vdd.n2133 vdd.n1054 9.3005
R21622 vdd.n1058 vdd.n1055 9.3005
R21623 vdd.n2128 vdd.n1059 9.3005
R21624 vdd.n2127 vdd.n1060 9.3005
R21625 vdd.n2126 vdd.n1061 9.3005
R21626 vdd.n1065 vdd.n1062 9.3005
R21627 vdd.n2121 vdd.n1066 9.3005
R21628 vdd.n2120 vdd.n1067 9.3005
R21629 vdd.n2119 vdd.n1068 9.3005
R21630 vdd.n1072 vdd.n1069 9.3005
R21631 vdd.n2114 vdd.n1073 9.3005
R21632 vdd.n2113 vdd.n1074 9.3005
R21633 vdd.n2112 vdd.n2111 9.3005
R21634 vdd.n2110 vdd.n1075 9.3005
R21635 vdd.n2109 vdd.n2108 9.3005
R21636 vdd.n1081 vdd.n1080 9.3005
R21637 vdd.n2103 vdd.n1085 9.3005
R21638 vdd.n2102 vdd.n1086 9.3005
R21639 vdd.n2101 vdd.n1087 9.3005
R21640 vdd.n1091 vdd.n1088 9.3005
R21641 vdd.n2096 vdd.n1092 9.3005
R21642 vdd.n2095 vdd.n1093 9.3005
R21643 vdd.n2094 vdd.n1094 9.3005
R21644 vdd.n1098 vdd.n1095 9.3005
R21645 vdd.n2089 vdd.n1099 9.3005
R21646 vdd.n2088 vdd.n1100 9.3005
R21647 vdd.n2087 vdd.n1101 9.3005
R21648 vdd.n1105 vdd.n1102 9.3005
R21649 vdd.n2082 vdd.n1106 9.3005
R21650 vdd.n2151 vdd.n2150 9.3005
R21651 vdd.n2173 vdd.n1006 9.3005
R21652 vdd.n2172 vdd.n1014 9.3005
R21653 vdd.n1018 vdd.n1015 9.3005
R21654 vdd.n2167 vdd.n1019 9.3005
R21655 vdd.n2166 vdd.n1020 9.3005
R21656 vdd.n2165 vdd.n1021 9.3005
R21657 vdd.n1025 vdd.n1022 9.3005
R21658 vdd.n2160 vdd.n1026 9.3005
R21659 vdd.n2159 vdd.n1027 9.3005
R21660 vdd.n2158 vdd.n1028 9.3005
R21661 vdd.n1032 vdd.n1029 9.3005
R21662 vdd.n2153 vdd.n1033 9.3005
R21663 vdd.n2152 vdd.n1034 9.3005
R21664 vdd.n2185 vdd.n2184 9.3005
R21665 vdd.n1010 vdd.n1009 9.3005
R21666 vdd.n2013 vdd.n1394 9.3005
R21667 vdd.n2015 vdd.n2014 9.3005
R21668 vdd.n1384 vdd.n1383 9.3005
R21669 vdd.n2029 vdd.n2028 9.3005
R21670 vdd.n2030 vdd.n1382 9.3005
R21671 vdd.n2032 vdd.n2031 9.3005
R21672 vdd.n1373 vdd.n1372 9.3005
R21673 vdd.n2046 vdd.n2045 9.3005
R21674 vdd.n2047 vdd.n1371 9.3005
R21675 vdd.n2049 vdd.n2048 9.3005
R21676 vdd.n1361 vdd.n1360 9.3005
R21677 vdd.n2065 vdd.n2064 9.3005
R21678 vdd.n2066 vdd.n1359 9.3005
R21679 vdd.n2068 vdd.n2067 9.3005
R21680 vdd.n283 vdd.n282 9.3005
R21681 vdd.n278 vdd.n277 9.3005
R21682 vdd.n289 vdd.n288 9.3005
R21683 vdd.n291 vdd.n290 9.3005
R21684 vdd.n274 vdd.n273 9.3005
R21685 vdd.n297 vdd.n296 9.3005
R21686 vdd.n299 vdd.n298 9.3005
R21687 vdd.n271 vdd.n268 9.3005
R21688 vdd.n306 vdd.n305 9.3005
R21689 vdd.n232 vdd.n231 9.3005
R21690 vdd.n227 vdd.n226 9.3005
R21691 vdd.n238 vdd.n237 9.3005
R21692 vdd.n240 vdd.n239 9.3005
R21693 vdd.n223 vdd.n222 9.3005
R21694 vdd.n246 vdd.n245 9.3005
R21695 vdd.n248 vdd.n247 9.3005
R21696 vdd.n220 vdd.n217 9.3005
R21697 vdd.n255 vdd.n254 9.3005
R21698 vdd.n189 vdd.n188 9.3005
R21699 vdd.n184 vdd.n183 9.3005
R21700 vdd.n195 vdd.n194 9.3005
R21701 vdd.n197 vdd.n196 9.3005
R21702 vdd.n180 vdd.n179 9.3005
R21703 vdd.n203 vdd.n202 9.3005
R21704 vdd.n205 vdd.n204 9.3005
R21705 vdd.n177 vdd.n174 9.3005
R21706 vdd.n212 vdd.n211 9.3005
R21707 vdd.n138 vdd.n137 9.3005
R21708 vdd.n133 vdd.n132 9.3005
R21709 vdd.n144 vdd.n143 9.3005
R21710 vdd.n146 vdd.n145 9.3005
R21711 vdd.n129 vdd.n128 9.3005
R21712 vdd.n152 vdd.n151 9.3005
R21713 vdd.n154 vdd.n153 9.3005
R21714 vdd.n126 vdd.n123 9.3005
R21715 vdd.n161 vdd.n160 9.3005
R21716 vdd.n96 vdd.n95 9.3005
R21717 vdd.n91 vdd.n90 9.3005
R21718 vdd.n102 vdd.n101 9.3005
R21719 vdd.n104 vdd.n103 9.3005
R21720 vdd.n87 vdd.n86 9.3005
R21721 vdd.n110 vdd.n109 9.3005
R21722 vdd.n112 vdd.n111 9.3005
R21723 vdd.n84 vdd.n81 9.3005
R21724 vdd.n119 vdd.n118 9.3005
R21725 vdd.n45 vdd.n44 9.3005
R21726 vdd.n40 vdd.n39 9.3005
R21727 vdd.n51 vdd.n50 9.3005
R21728 vdd.n53 vdd.n52 9.3005
R21729 vdd.n36 vdd.n35 9.3005
R21730 vdd.n59 vdd.n58 9.3005
R21731 vdd.n61 vdd.n60 9.3005
R21732 vdd.n33 vdd.n30 9.3005
R21733 vdd.n68 vdd.n67 9.3005
R21734 vdd.n3126 vdd.n3125 9.3005
R21735 vdd.n3127 vdd.n578 9.3005
R21736 vdd.n577 vdd.n575 9.3005
R21737 vdd.n3133 vdd.n574 9.3005
R21738 vdd.n3134 vdd.n573 9.3005
R21739 vdd.n3135 vdd.n572 9.3005
R21740 vdd.n571 vdd.n569 9.3005
R21741 vdd.n3141 vdd.n568 9.3005
R21742 vdd.n3142 vdd.n567 9.3005
R21743 vdd.n3143 vdd.n566 9.3005
R21744 vdd.n565 vdd.n563 9.3005
R21745 vdd.n3149 vdd.n562 9.3005
R21746 vdd.n3150 vdd.n561 9.3005
R21747 vdd.n3151 vdd.n560 9.3005
R21748 vdd.n559 vdd.n557 9.3005
R21749 vdd.n3157 vdd.n556 9.3005
R21750 vdd.n3158 vdd.n555 9.3005
R21751 vdd.n3159 vdd.n554 9.3005
R21752 vdd.n553 vdd.n551 9.3005
R21753 vdd.n3165 vdd.n550 9.3005
R21754 vdd.n3166 vdd.n549 9.3005
R21755 vdd.n3167 vdd.n548 9.3005
R21756 vdd.n547 vdd.n545 9.3005
R21757 vdd.n3173 vdd.n542 9.3005
R21758 vdd.n3174 vdd.n541 9.3005
R21759 vdd.n3175 vdd.n540 9.3005
R21760 vdd.n539 vdd.n537 9.3005
R21761 vdd.n3181 vdd.n536 9.3005
R21762 vdd.n3182 vdd.n535 9.3005
R21763 vdd.n3183 vdd.n534 9.3005
R21764 vdd.n533 vdd.n531 9.3005
R21765 vdd.n3189 vdd.n530 9.3005
R21766 vdd.n3190 vdd.n529 9.3005
R21767 vdd.n3191 vdd.n528 9.3005
R21768 vdd.n527 vdd.n525 9.3005
R21769 vdd.n3196 vdd.n524 9.3005
R21770 vdd.n3206 vdd.n518 9.3005
R21771 vdd.n3208 vdd.n3207 9.3005
R21772 vdd.n509 vdd.n508 9.3005
R21773 vdd.n3223 vdd.n3222 9.3005
R21774 vdd.n3224 vdd.n507 9.3005
R21775 vdd.n3226 vdd.n3225 9.3005
R21776 vdd.n497 vdd.n496 9.3005
R21777 vdd.n3239 vdd.n3238 9.3005
R21778 vdd.n3240 vdd.n495 9.3005
R21779 vdd.n3242 vdd.n3241 9.3005
R21780 vdd.n485 vdd.n484 9.3005
R21781 vdd.n3256 vdd.n3255 9.3005
R21782 vdd.n3257 vdd.n483 9.3005
R21783 vdd.n3259 vdd.n3258 9.3005
R21784 vdd.n312 vdd.n310 9.3005
R21785 vdd.n3210 vdd.n3209 9.3005
R21786 vdd.n3439 vdd.n3438 9.3005
R21787 vdd.n313 vdd.n311 9.3005
R21788 vdd.n3432 vdd.n320 9.3005
R21789 vdd.n3431 vdd.n321 9.3005
R21790 vdd.n3430 vdd.n322 9.3005
R21791 vdd.n331 vdd.n323 9.3005
R21792 vdd.n3424 vdd.n332 9.3005
R21793 vdd.n3423 vdd.n333 9.3005
R21794 vdd.n3422 vdd.n334 9.3005
R21795 vdd.n342 vdd.n335 9.3005
R21796 vdd.n3416 vdd.n343 9.3005
R21797 vdd.n3415 vdd.n344 9.3005
R21798 vdd.n3414 vdd.n345 9.3005
R21799 vdd.n353 vdd.n346 9.3005
R21800 vdd.n3408 vdd.n3407 9.3005
R21801 vdd.n3404 vdd.n354 9.3005
R21802 vdd.n3403 vdd.n357 9.3005
R21803 vdd.n361 vdd.n358 9.3005
R21804 vdd.n362 vdd.n359 9.3005
R21805 vdd.n3396 vdd.n363 9.3005
R21806 vdd.n3395 vdd.n364 9.3005
R21807 vdd.n3394 vdd.n365 9.3005
R21808 vdd.n369 vdd.n366 9.3005
R21809 vdd.n3389 vdd.n370 9.3005
R21810 vdd.n3388 vdd.n371 9.3005
R21811 vdd.n3387 vdd.n372 9.3005
R21812 vdd.n376 vdd.n373 9.3005
R21813 vdd.n3382 vdd.n377 9.3005
R21814 vdd.n3381 vdd.n378 9.3005
R21815 vdd.n3380 vdd.n379 9.3005
R21816 vdd.n383 vdd.n380 9.3005
R21817 vdd.n3375 vdd.n384 9.3005
R21818 vdd.n3374 vdd.n385 9.3005
R21819 vdd.n3373 vdd.n3372 9.3005
R21820 vdd.n3371 vdd.n386 9.3005
R21821 vdd.n3370 vdd.n3369 9.3005
R21822 vdd.n392 vdd.n391 9.3005
R21823 vdd.n3364 vdd.n396 9.3005
R21824 vdd.n3363 vdd.n397 9.3005
R21825 vdd.n3362 vdd.n398 9.3005
R21826 vdd.n402 vdd.n399 9.3005
R21827 vdd.n3357 vdd.n403 9.3005
R21828 vdd.n3356 vdd.n404 9.3005
R21829 vdd.n3355 vdd.n405 9.3005
R21830 vdd.n409 vdd.n406 9.3005
R21831 vdd.n3350 vdd.n410 9.3005
R21832 vdd.n3349 vdd.n411 9.3005
R21833 vdd.n3348 vdd.n412 9.3005
R21834 vdd.n416 vdd.n413 9.3005
R21835 vdd.n3343 vdd.n417 9.3005
R21836 vdd.n3342 vdd.n418 9.3005
R21837 vdd.n3341 vdd.n419 9.3005
R21838 vdd.n423 vdd.n420 9.3005
R21839 vdd.n3336 vdd.n424 9.3005
R21840 vdd.n3335 vdd.n425 9.3005
R21841 vdd.n3334 vdd.n3333 9.3005
R21842 vdd.n3332 vdd.n426 9.3005
R21843 vdd.n3331 vdd.n3330 9.3005
R21844 vdd.n432 vdd.n431 9.3005
R21845 vdd.n3325 vdd.n436 9.3005
R21846 vdd.n3324 vdd.n437 9.3005
R21847 vdd.n3323 vdd.n438 9.3005
R21848 vdd.n442 vdd.n439 9.3005
R21849 vdd.n3318 vdd.n443 9.3005
R21850 vdd.n3317 vdd.n444 9.3005
R21851 vdd.n3316 vdd.n445 9.3005
R21852 vdd.n449 vdd.n446 9.3005
R21853 vdd.n3311 vdd.n450 9.3005
R21854 vdd.n3310 vdd.n451 9.3005
R21855 vdd.n3309 vdd.n452 9.3005
R21856 vdd.n456 vdd.n453 9.3005
R21857 vdd.n3304 vdd.n457 9.3005
R21858 vdd.n3303 vdd.n458 9.3005
R21859 vdd.n3302 vdd.n459 9.3005
R21860 vdd.n463 vdd.n460 9.3005
R21861 vdd.n3297 vdd.n464 9.3005
R21862 vdd.n3296 vdd.n465 9.3005
R21863 vdd.n3292 vdd.n3289 9.3005
R21864 vdd.n3406 vdd.n3405 9.3005
R21865 vdd.n3216 vdd.n513 9.3005
R21866 vdd.n3218 vdd.n3217 9.3005
R21867 vdd.n503 vdd.n502 9.3005
R21868 vdd.n3231 vdd.n3230 9.3005
R21869 vdd.n3232 vdd.n501 9.3005
R21870 vdd.n3234 vdd.n3233 9.3005
R21871 vdd.n490 vdd.n489 9.3005
R21872 vdd.n3247 vdd.n3246 9.3005
R21873 vdd.n3248 vdd.n488 9.3005
R21874 vdd.n3250 vdd.n3249 9.3005
R21875 vdd.n478 vdd.n477 9.3005
R21876 vdd.n3264 vdd.n3263 9.3005
R21877 vdd.n3265 vdd.n476 9.3005
R21878 vdd.n3267 vdd.n3266 9.3005
R21879 vdd.n3268 vdd.n475 9.3005
R21880 vdd.n3270 vdd.n3269 9.3005
R21881 vdd.n3271 vdd.n474 9.3005
R21882 vdd.n3273 vdd.n3272 9.3005
R21883 vdd.n3274 vdd.n472 9.3005
R21884 vdd.n3276 vdd.n3275 9.3005
R21885 vdd.n3277 vdd.n471 9.3005
R21886 vdd.n3279 vdd.n3278 9.3005
R21887 vdd.n3280 vdd.n469 9.3005
R21888 vdd.n3282 vdd.n3281 9.3005
R21889 vdd.n3283 vdd.n468 9.3005
R21890 vdd.n3285 vdd.n3284 9.3005
R21891 vdd.n3286 vdd.n466 9.3005
R21892 vdd.n3288 vdd.n3287 9.3005
R21893 vdd.n3215 vdd.n3214 9.3005
R21894 vdd.n3079 vdd.n514 9.3005
R21895 vdd.n3084 vdd.n3078 9.3005
R21896 vdd.n3094 vdd.n605 9.3005
R21897 vdd.n3095 vdd.n604 9.3005
R21898 vdd.n603 vdd.n601 9.3005
R21899 vdd.n3101 vdd.n600 9.3005
R21900 vdd.n3102 vdd.n599 9.3005
R21901 vdd.n3103 vdd.n598 9.3005
R21902 vdd.n597 vdd.n595 9.3005
R21903 vdd.n3109 vdd.n594 9.3005
R21904 vdd.n3110 vdd.n593 9.3005
R21905 vdd.n3111 vdd.n592 9.3005
R21906 vdd.n591 vdd.n589 9.3005
R21907 vdd.n3116 vdd.n588 9.3005
R21908 vdd.n3117 vdd.n587 9.3005
R21909 vdd.n583 vdd.n582 9.3005
R21910 vdd.n3123 vdd.n3122 9.3005
R21911 vdd.n3124 vdd.n579 9.3005
R21912 vdd.n2078 vdd.n2077 9.3005
R21913 vdd.n2073 vdd.n1345 9.3005
R21914 vdd.n1674 vdd.n1434 9.3005
R21915 vdd.n1676 vdd.n1675 9.3005
R21916 vdd.n1425 vdd.n1424 9.3005
R21917 vdd.n1689 vdd.n1688 9.3005
R21918 vdd.n1690 vdd.n1423 9.3005
R21919 vdd.n1692 vdd.n1691 9.3005
R21920 vdd.n1412 vdd.n1411 9.3005
R21921 vdd.n1705 vdd.n1704 9.3005
R21922 vdd.n1706 vdd.n1410 9.3005
R21923 vdd.n1708 vdd.n1707 9.3005
R21924 vdd.n1401 vdd.n1400 9.3005
R21925 vdd.n1722 vdd.n1721 9.3005
R21926 vdd.n1723 vdd.n1399 9.3005
R21927 vdd.n1725 vdd.n1724 9.3005
R21928 vdd.n1390 vdd.n1389 9.3005
R21929 vdd.n2020 vdd.n2019 9.3005
R21930 vdd.n2021 vdd.n1388 9.3005
R21931 vdd.n2023 vdd.n2022 9.3005
R21932 vdd.n1378 vdd.n1377 9.3005
R21933 vdd.n2037 vdd.n2036 9.3005
R21934 vdd.n2038 vdd.n1376 9.3005
R21935 vdd.n2040 vdd.n2039 9.3005
R21936 vdd.n1368 vdd.n1367 9.3005
R21937 vdd.n2054 vdd.n2053 9.3005
R21938 vdd.n2055 vdd.n1365 9.3005
R21939 vdd.n2059 vdd.n2058 9.3005
R21940 vdd.n2057 vdd.n1366 9.3005
R21941 vdd.n2056 vdd.n1356 9.3005
R21942 vdd.n1673 vdd.n1672 9.3005
R21943 vdd.n1568 vdd.n1558 9.3005
R21944 vdd.n1570 vdd.n1569 9.3005
R21945 vdd.n1571 vdd.n1557 9.3005
R21946 vdd.n1573 vdd.n1572 9.3005
R21947 vdd.n1574 vdd.n1550 9.3005
R21948 vdd.n1576 vdd.n1575 9.3005
R21949 vdd.n1577 vdd.n1549 9.3005
R21950 vdd.n1579 vdd.n1578 9.3005
R21951 vdd.n1580 vdd.n1542 9.3005
R21952 vdd.n1582 vdd.n1581 9.3005
R21953 vdd.n1583 vdd.n1541 9.3005
R21954 vdd.n1585 vdd.n1584 9.3005
R21955 vdd.n1586 vdd.n1534 9.3005
R21956 vdd.n1588 vdd.n1587 9.3005
R21957 vdd.n1589 vdd.n1533 9.3005
R21958 vdd.n1591 vdd.n1590 9.3005
R21959 vdd.n1592 vdd.n1527 9.3005
R21960 vdd.n1594 vdd.n1593 9.3005
R21961 vdd.n1595 vdd.n1525 9.3005
R21962 vdd.n1597 vdd.n1596 9.3005
R21963 vdd.n1526 vdd.n1523 9.3005
R21964 vdd.n1604 vdd.n1519 9.3005
R21965 vdd.n1606 vdd.n1605 9.3005
R21966 vdd.n1607 vdd.n1518 9.3005
R21967 vdd.n1609 vdd.n1608 9.3005
R21968 vdd.n1610 vdd.n1511 9.3005
R21969 vdd.n1612 vdd.n1611 9.3005
R21970 vdd.n1613 vdd.n1510 9.3005
R21971 vdd.n1615 vdd.n1614 9.3005
R21972 vdd.n1616 vdd.n1503 9.3005
R21973 vdd.n1618 vdd.n1617 9.3005
R21974 vdd.n1619 vdd.n1502 9.3005
R21975 vdd.n1621 vdd.n1620 9.3005
R21976 vdd.n1622 vdd.n1495 9.3005
R21977 vdd.n1624 vdd.n1623 9.3005
R21978 vdd.n1625 vdd.n1494 9.3005
R21979 vdd.n1627 vdd.n1626 9.3005
R21980 vdd.n1628 vdd.n1487 9.3005
R21981 vdd.n1630 vdd.n1629 9.3005
R21982 vdd.n1631 vdd.n1486 9.3005
R21983 vdd.n1633 vdd.n1632 9.3005
R21984 vdd.n1634 vdd.n1479 9.3005
R21985 vdd.n1636 vdd.n1635 9.3005
R21986 vdd.n1637 vdd.n1478 9.3005
R21987 vdd.n1639 vdd.n1638 9.3005
R21988 vdd.n1640 vdd.n1469 9.3005
R21989 vdd.n1642 vdd.n1641 9.3005
R21990 vdd.n1643 vdd.n1468 9.3005
R21991 vdd.n1645 vdd.n1644 9.3005
R21992 vdd.n1646 vdd.n1461 9.3005
R21993 vdd.n1648 vdd.n1647 9.3005
R21994 vdd.n1649 vdd.n1460 9.3005
R21995 vdd.n1651 vdd.n1650 9.3005
R21996 vdd.n1652 vdd.n1453 9.3005
R21997 vdd.n1654 vdd.n1653 9.3005
R21998 vdd.n1655 vdd.n1452 9.3005
R21999 vdd.n1657 vdd.n1656 9.3005
R22000 vdd.n1658 vdd.n1445 9.3005
R22001 vdd.n1660 vdd.n1659 9.3005
R22002 vdd.n1661 vdd.n1444 9.3005
R22003 vdd.n1663 vdd.n1662 9.3005
R22004 vdd.n1664 vdd.n1440 9.3005
R22005 vdd.n1666 vdd.n1665 9.3005
R22006 vdd.n1564 vdd.n1435 9.3005
R22007 vdd.n1431 vdd.n1430 9.3005
R22008 vdd.n1681 vdd.n1680 9.3005
R22009 vdd.n1682 vdd.n1429 9.3005
R22010 vdd.n1684 vdd.n1683 9.3005
R22011 vdd.n1419 vdd.n1418 9.3005
R22012 vdd.n1697 vdd.n1696 9.3005
R22013 vdd.n1698 vdd.n1417 9.3005
R22014 vdd.n1700 vdd.n1699 9.3005
R22015 vdd.n1407 vdd.n1406 9.3005
R22016 vdd.n1714 vdd.n1713 9.3005
R22017 vdd.n1715 vdd.n1405 9.3005
R22018 vdd.n1717 vdd.n1716 9.3005
R22019 vdd.n1396 vdd.n1395 9.3005
R22020 vdd.n1668 vdd.n1667 9.3005
R22021 vdd.n2012 vdd.n1729 9.3005
R22022 vdd.n1933 vdd.n1932 9.3005
R22023 vdd.n1928 vdd.n1927 9.3005
R22024 vdd.n1939 vdd.n1938 9.3005
R22025 vdd.n1941 vdd.n1940 9.3005
R22026 vdd.n1924 vdd.n1923 9.3005
R22027 vdd.n1947 vdd.n1946 9.3005
R22028 vdd.n1949 vdd.n1948 9.3005
R22029 vdd.n1921 vdd.n1918 9.3005
R22030 vdd.n1956 vdd.n1955 9.3005
R22031 vdd.n1984 vdd.n1983 9.3005
R22032 vdd.n1979 vdd.n1978 9.3005
R22033 vdd.n1990 vdd.n1989 9.3005
R22034 vdd.n1992 vdd.n1991 9.3005
R22035 vdd.n1975 vdd.n1974 9.3005
R22036 vdd.n1998 vdd.n1997 9.3005
R22037 vdd.n2000 vdd.n1999 9.3005
R22038 vdd.n1972 vdd.n1969 9.3005
R22039 vdd.n2007 vdd.n2006 9.3005
R22040 vdd.n1839 vdd.n1838 9.3005
R22041 vdd.n1834 vdd.n1833 9.3005
R22042 vdd.n1845 vdd.n1844 9.3005
R22043 vdd.n1847 vdd.n1846 9.3005
R22044 vdd.n1830 vdd.n1829 9.3005
R22045 vdd.n1853 vdd.n1852 9.3005
R22046 vdd.n1855 vdd.n1854 9.3005
R22047 vdd.n1827 vdd.n1824 9.3005
R22048 vdd.n1862 vdd.n1861 9.3005
R22049 vdd.n1890 vdd.n1889 9.3005
R22050 vdd.n1885 vdd.n1884 9.3005
R22051 vdd.n1896 vdd.n1895 9.3005
R22052 vdd.n1898 vdd.n1897 9.3005
R22053 vdd.n1881 vdd.n1880 9.3005
R22054 vdd.n1904 vdd.n1903 9.3005
R22055 vdd.n1906 vdd.n1905 9.3005
R22056 vdd.n1878 vdd.n1875 9.3005
R22057 vdd.n1913 vdd.n1912 9.3005
R22058 vdd.n1746 vdd.n1745 9.3005
R22059 vdd.n1741 vdd.n1740 9.3005
R22060 vdd.n1752 vdd.n1751 9.3005
R22061 vdd.n1754 vdd.n1753 9.3005
R22062 vdd.n1737 vdd.n1736 9.3005
R22063 vdd.n1760 vdd.n1759 9.3005
R22064 vdd.n1762 vdd.n1761 9.3005
R22065 vdd.n1734 vdd.n1731 9.3005
R22066 vdd.n1769 vdd.n1768 9.3005
R22067 vdd.n1797 vdd.n1796 9.3005
R22068 vdd.n1792 vdd.n1791 9.3005
R22069 vdd.n1803 vdd.n1802 9.3005
R22070 vdd.n1805 vdd.n1804 9.3005
R22071 vdd.n1788 vdd.n1787 9.3005
R22072 vdd.n1811 vdd.n1810 9.3005
R22073 vdd.n1813 vdd.n1812 9.3005
R22074 vdd.n1785 vdd.n1782 9.3005
R22075 vdd.n1820 vdd.n1819 9.3005
R22076 vdd.n288 vdd.n287 8.92171
R22077 vdd.n237 vdd.n236 8.92171
R22078 vdd.n194 vdd.n193 8.92171
R22079 vdd.n143 vdd.n142 8.92171
R22080 vdd.n101 vdd.n100 8.92171
R22081 vdd.n50 vdd.n49 8.92171
R22082 vdd.n1938 vdd.n1937 8.92171
R22083 vdd.n1989 vdd.n1988 8.92171
R22084 vdd.n1844 vdd.n1843 8.92171
R22085 vdd.n1895 vdd.n1894 8.92171
R22086 vdd.n1751 vdd.n1750 8.92171
R22087 vdd.n1802 vdd.n1801 8.92171
R22088 vdd.n215 vdd.n121 8.81535
R22089 vdd.n1916 vdd.n1822 8.81535
R22090 vdd.n2051 vdd.t177 8.72962
R22091 vdd.n3228 vdd.t200 8.72962
R22092 vdd.t156 vdd.n2025 8.50289
R22093 vdd.n493 vdd.t165 8.50289
R22094 vdd.n28 vdd.n14 8.42249
R22095 vdd.n1727 vdd.t150 8.27616
R22096 vdd.n3436 vdd.t198 8.27616
R22097 vdd.n3440 vdd.n3439 8.16225
R22098 vdd.n2012 vdd.n2011 8.16225
R22099 vdd.n284 vdd.n278 8.14595
R22100 vdd.n233 vdd.n227 8.14595
R22101 vdd.n190 vdd.n184 8.14595
R22102 vdd.n139 vdd.n133 8.14595
R22103 vdd.n97 vdd.n91 8.14595
R22104 vdd.n46 vdd.n40 8.14595
R22105 vdd.n1934 vdd.n1928 8.14595
R22106 vdd.n1985 vdd.n1979 8.14595
R22107 vdd.n1840 vdd.n1834 8.14595
R22108 vdd.n1891 vdd.n1885 8.14595
R22109 vdd.n1747 vdd.n1741 8.14595
R22110 vdd.n1798 vdd.n1792 8.14595
R22111 vdd.t205 vdd.n1415 8.04943
R22112 vdd.n3427 vdd.t186 8.04943
R22113 vdd.n2225 vdd.n962 7.70933
R22114 vdd.n2225 vdd.n965 7.70933
R22115 vdd.n2231 vdd.n951 7.70933
R22116 vdd.n2237 vdd.n951 7.70933
R22117 vdd.n2237 vdd.n944 7.70933
R22118 vdd.n2243 vdd.n944 7.70933
R22119 vdd.n2243 vdd.n947 7.70933
R22120 vdd.n2249 vdd.n940 7.70933
R22121 vdd.n2255 vdd.n934 7.70933
R22122 vdd.n2261 vdd.n921 7.70933
R22123 vdd.n2267 vdd.n921 7.70933
R22124 vdd.n2273 vdd.n915 7.70933
R22125 vdd.n2279 vdd.n908 7.70933
R22126 vdd.n2279 vdd.n911 7.70933
R22127 vdd.n2285 vdd.n904 7.70933
R22128 vdd.n2292 vdd.n890 7.70933
R22129 vdd.n2298 vdd.n890 7.70933
R22130 vdd.n2304 vdd.n884 7.70933
R22131 vdd.n2310 vdd.n880 7.70933
R22132 vdd.n2316 vdd.n874 7.70933
R22133 vdd.n2334 vdd.n856 7.70933
R22134 vdd.n2334 vdd.n849 7.70933
R22135 vdd.n2342 vdd.n849 7.70933
R22136 vdd.n2424 vdd.n833 7.70933
R22137 vdd.n2807 vdd.n785 7.70933
R22138 vdd.n2819 vdd.n774 7.70933
R22139 vdd.n2819 vdd.n768 7.70933
R22140 vdd.n2825 vdd.n768 7.70933
R22141 vdd.n2837 vdd.n759 7.70933
R22142 vdd.n2843 vdd.n753 7.70933
R22143 vdd.n2855 vdd.n740 7.70933
R22144 vdd.n2862 vdd.n733 7.70933
R22145 vdd.n2862 vdd.n736 7.70933
R22146 vdd.n2868 vdd.n729 7.70933
R22147 vdd.n2874 vdd.n715 7.70933
R22148 vdd.n2880 vdd.n715 7.70933
R22149 vdd.n2886 vdd.n709 7.70933
R22150 vdd.n2892 vdd.n702 7.70933
R22151 vdd.n2892 vdd.n705 7.70933
R22152 vdd.n2898 vdd.n698 7.70933
R22153 vdd.n2904 vdd.n692 7.70933
R22154 vdd.n2910 vdd.n679 7.70933
R22155 vdd.n2916 vdd.n679 7.70933
R22156 vdd.n2916 vdd.n671 7.70933
R22157 vdd.n2967 vdd.n671 7.70933
R22158 vdd.n2967 vdd.n674 7.70933
R22159 vdd.n2973 vdd.n631 7.70933
R22160 vdd.n3043 vdd.n631 7.70933
R22161 vdd.n283 vdd.n280 7.3702
R22162 vdd.n232 vdd.n229 7.3702
R22163 vdd.n189 vdd.n186 7.3702
R22164 vdd.n138 vdd.n135 7.3702
R22165 vdd.n96 vdd.n93 7.3702
R22166 vdd.n45 vdd.n42 7.3702
R22167 vdd.n1933 vdd.n1930 7.3702
R22168 vdd.n1984 vdd.n1981 7.3702
R22169 vdd.n1839 vdd.n1836 7.3702
R22170 vdd.n1890 vdd.n1887 7.3702
R22171 vdd.n1746 vdd.n1743 7.3702
R22172 vdd.n1797 vdd.n1794 7.3702
R22173 vdd.n934 vdd.t129 7.36923
R22174 vdd.n2898 vdd.t106 7.36923
R22175 vdd.n1694 vdd.t148 7.1425
R22176 vdd.n2249 vdd.t81 7.1425
R22177 vdd.n1253 vdd.t77 7.1425
R22178 vdd.n2831 vdd.t80 7.1425
R22179 vdd.n692 vdd.t90 7.1425
R22180 vdd.n3420 vdd.t220 7.1425
R22181 vdd.n1605 vdd.n1604 6.98232
R22182 vdd.n2113 vdd.n2112 6.98232
R22183 vdd.n3335 vdd.n3334 6.98232
R22184 vdd.n3127 vdd.n3126 6.98232
R22185 vdd.n1710 vdd.t154 6.91577
R22186 vdd.n325 vdd.t192 6.91577
R22187 vdd.n1253 vdd.t78 6.80241
R22188 vdd.n2831 vdd.t122 6.80241
R22189 vdd.n2017 vdd.t173 6.68904
R22190 vdd.n3261 vdd.t216 6.68904
R22191 vdd.n1380 vdd.t207 6.46231
R22192 vdd.n2273 vdd.t88 6.46231
R22193 vdd.t93 vdd.n884 6.46231
R22194 vdd.n2855 vdd.t98 6.46231
R22195 vdd.t114 vdd.n709 6.46231
R22196 vdd.t180 vdd.n492 6.46231
R22197 vdd.n2349 vdd.t126 6.34895
R22198 vdd.n2728 vdd.t111 6.34895
R22199 vdd.n3440 vdd.n309 6.27748
R22200 vdd.n2011 vdd.n2010 6.27748
R22201 vdd.n2870 vdd.n725 6.2444
R22202 vdd.n2289 vdd.n2288 6.2444
R22203 vdd.n2310 vdd.t119 5.89549
R22204 vdd.n753 vdd.t94 5.89549
R22205 vdd.n284 vdd.n283 5.81868
R22206 vdd.n233 vdd.n232 5.81868
R22207 vdd.n190 vdd.n189 5.81868
R22208 vdd.n139 vdd.n138 5.81868
R22209 vdd.n97 vdd.n96 5.81868
R22210 vdd.n46 vdd.n45 5.81868
R22211 vdd.n1934 vdd.n1933 5.81868
R22212 vdd.n1985 vdd.n1984 5.81868
R22213 vdd.n1840 vdd.n1839 5.81868
R22214 vdd.n1891 vdd.n1890 5.81868
R22215 vdd.n1747 vdd.n1746 5.81868
R22216 vdd.n1798 vdd.n1797 5.81868
R22217 vdd.n2432 vdd.n2431 5.77611
R22218 vdd.n1177 vdd.n1176 5.77611
R22219 vdd.n2740 vdd.n2739 5.77611
R22220 vdd.n2982 vdd.n663 5.77611
R22221 vdd.n3048 vdd.n627 5.77611
R22222 vdd.n2603 vdd.n2537 5.77611
R22223 vdd.n2357 vdd.n840 5.77611
R22224 vdd.n1313 vdd.n1145 5.77611
R22225 vdd.n1567 vdd.n1564 5.62474
R22226 vdd.n2076 vdd.n2073 5.62474
R22227 vdd.n3295 vdd.n3292 5.62474
R22228 vdd.n3082 vdd.n3079 5.62474
R22229 vdd.n2285 vdd.t108 5.55539
R22230 vdd.n729 vdd.t84 5.55539
R22231 vdd.n287 vdd.n278 5.04292
R22232 vdd.n236 vdd.n227 5.04292
R22233 vdd.n193 vdd.n184 5.04292
R22234 vdd.n142 vdd.n133 5.04292
R22235 vdd.n100 vdd.n91 5.04292
R22236 vdd.n49 vdd.n40 5.04292
R22237 vdd.n1937 vdd.n1928 5.04292
R22238 vdd.n1988 vdd.n1979 5.04292
R22239 vdd.n1843 vdd.n1834 5.04292
R22240 vdd.n1894 vdd.n1885 5.04292
R22241 vdd.n1750 vdd.n1741 5.04292
R22242 vdd.n1801 vdd.n1792 5.04292
R22243 vdd.n2043 vdd.t207 4.8752
R22244 vdd.t87 vdd.t100 4.8752
R22245 vdd.t130 vdd.t76 4.8752
R22246 vdd.n3236 vdd.t180 4.8752
R22247 vdd.n2433 vdd.n2432 4.83952
R22248 vdd.n1176 vdd.n1175 4.83952
R22249 vdd.n2741 vdd.n2740 4.83952
R22250 vdd.n663 vdd.n658 4.83952
R22251 vdd.n627 vdd.n622 4.83952
R22252 vdd.n2600 vdd.n2537 4.83952
R22253 vdd.n2360 vdd.n840 4.83952
R22254 vdd.n1316 vdd.n1145 4.83952
R22255 vdd.n1227 vdd.t96 4.76184
R22256 vdd.n2813 vdd.t82 4.76184
R22257 vdd.n2081 vdd.n2080 4.74817
R22258 vdd.n1349 vdd.n1344 4.74817
R22259 vdd.n1011 vdd.n1008 4.74817
R22260 vdd.n2174 vdd.n1007 4.74817
R22261 vdd.n2179 vdd.n1008 4.74817
R22262 vdd.n2178 vdd.n1007 4.74817
R22263 vdd.n521 vdd.n519 4.74817
R22264 vdd.n3197 vdd.n522 4.74817
R22265 vdd.n3200 vdd.n522 4.74817
R22266 vdd.n3201 vdd.n521 4.74817
R22267 vdd.n3089 vdd.n606 4.74817
R22268 vdd.n3085 vdd.n608 4.74817
R22269 vdd.n3088 vdd.n608 4.74817
R22270 vdd.n3093 vdd.n606 4.74817
R22271 vdd.n2080 vdd.n1107 4.74817
R22272 vdd.n1346 vdd.n1344 4.74817
R22273 vdd.n309 vdd.n308 4.7074
R22274 vdd.n215 vdd.n214 4.7074
R22275 vdd.n2010 vdd.n2009 4.7074
R22276 vdd.n1916 vdd.n1915 4.7074
R22277 vdd.t173 vdd.n1386 4.64847
R22278 vdd.t89 vdd.n915 4.64847
R22279 vdd.n2304 vdd.t128 4.64847
R22280 vdd.t117 vdd.n740 4.64847
R22281 vdd.n2886 vdd.t113 4.64847
R22282 vdd.n3252 vdd.t216 4.64847
R22283 vdd.n904 vdd.t64 4.53511
R22284 vdd.n2868 vdd.t27 4.53511
R22285 vdd.n1719 vdd.t154 4.42174
R22286 vdd.n2231 vdd.t5 4.42174
R22287 vdd.n1227 vdd.t50 4.42174
R22288 vdd.n2813 vdd.t57 4.42174
R22289 vdd.n674 vdd.t1 4.42174
R22290 vdd.n3434 vdd.t192 4.42174
R22291 vdd.n2859 vdd.n725 4.37123
R22292 vdd.n2290 vdd.n2289 4.37123
R22293 vdd.n2328 vdd.t115 4.30838
R22294 vdd.n2716 vdd.t102 4.30838
R22295 vdd.n288 vdd.n276 4.26717
R22296 vdd.n237 vdd.n225 4.26717
R22297 vdd.n194 vdd.n182 4.26717
R22298 vdd.n143 vdd.n131 4.26717
R22299 vdd.n101 vdd.n89 4.26717
R22300 vdd.n50 vdd.n38 4.26717
R22301 vdd.n1938 vdd.n1926 4.26717
R22302 vdd.n1989 vdd.n1977 4.26717
R22303 vdd.n1844 vdd.n1832 4.26717
R22304 vdd.n1895 vdd.n1883 4.26717
R22305 vdd.n1751 vdd.n1739 4.26717
R22306 vdd.n1802 vdd.n1790 4.26717
R22307 vdd.t148 vdd.n1414 4.19501
R22308 vdd.t220 vdd.n329 4.19501
R22309 vdd.n309 vdd.n215 4.10845
R22310 vdd.n2010 vdd.n1916 4.10845
R22311 vdd.n265 vdd.t196 4.06363
R22312 vdd.n265 vdd.t227 4.06363
R22313 vdd.n263 vdd.t229 4.06363
R22314 vdd.n263 vdd.t153 4.06363
R22315 vdd.n261 vdd.t172 4.06363
R22316 vdd.n261 vdd.t212 4.06363
R22317 vdd.n259 vdd.t230 4.06363
R22318 vdd.n259 vdd.t238 4.06363
R22319 vdd.n257 vdd.t241 4.06363
R22320 vdd.n257 vdd.t179 4.06363
R22321 vdd.n171 vdd.t187 4.06363
R22322 vdd.n171 vdd.t221 4.06363
R22323 vdd.n169 vdd.t222 4.06363
R22324 vdd.n169 vdd.t239 4.06363
R22325 vdd.n167 vdd.t159 4.06363
R22326 vdd.n167 vdd.t199 4.06363
R22327 vdd.n165 vdd.t225 4.06363
R22328 vdd.n165 vdd.t231 4.06363
R22329 vdd.n163 vdd.t235 4.06363
R22330 vdd.n163 vdd.t163 4.06363
R22331 vdd.n78 vdd.t204 4.06363
R22332 vdd.n78 vdd.t223 4.06363
R22333 vdd.n76 vdd.t193 4.06363
R22334 vdd.n76 vdd.t236 4.06363
R22335 vdd.n74 vdd.t171 4.06363
R22336 vdd.n74 vdd.t228 4.06363
R22337 vdd.n72 vdd.t166 4.06363
R22338 vdd.n72 vdd.t217 4.06363
R22339 vdd.n70 vdd.t181 4.06363
R22340 vdd.n70 vdd.t232 4.06363
R22341 vdd.n1958 vdd.t215 4.06363
R22342 vdd.n1958 vdd.t214 4.06363
R22343 vdd.n1960 vdd.t188 4.06363
R22344 vdd.n1960 vdd.t170 4.06363
R22345 vdd.n1962 vdd.t168 4.06363
R22346 vdd.n1962 vdd.t213 4.06363
R22347 vdd.n1964 vdd.t197 4.06363
R22348 vdd.n1964 vdd.t169 4.06363
R22349 vdd.n1966 vdd.t164 4.06363
R22350 vdd.n1966 vdd.t226 4.06363
R22351 vdd.n1864 vdd.t210 4.06363
R22352 vdd.n1864 vdd.t208 4.06363
R22353 vdd.n1866 vdd.t174 4.06363
R22354 vdd.n1866 vdd.t157 4.06363
R22355 vdd.n1868 vdd.t151 4.06363
R22356 vdd.n1868 vdd.t203 4.06363
R22357 vdd.n1870 vdd.t190 4.06363
R22358 vdd.n1870 vdd.t155 4.06363
R22359 vdd.n1872 vdd.t149 4.06363
R22360 vdd.n1872 vdd.t219 4.06363
R22361 vdd.n1771 vdd.t233 4.06363
R22362 vdd.n1771 vdd.t243 4.06363
R22363 vdd.n1773 vdd.t218 4.06363
R22364 vdd.n1773 vdd.t167 4.06363
R22365 vdd.n1775 vdd.t211 4.06363
R22366 vdd.n1775 vdd.t176 4.06363
R22367 vdd.n1777 vdd.t237 4.06363
R22368 vdd.n1777 vdd.t194 4.06363
R22369 vdd.n1779 vdd.t224 4.06363
R22370 vdd.n1779 vdd.t206 4.06363
R22371 vdd.n940 vdd.t121 3.96828
R22372 vdd.n2322 vdd.t99 3.96828
R22373 vdd.n2710 vdd.t118 3.96828
R22374 vdd.n2904 vdd.t107 3.96828
R22375 vdd.n26 vdd.t147 3.9605
R22376 vdd.n26 vdd.t140 3.9605
R22377 vdd.n23 vdd.t142 3.9605
R22378 vdd.n23 vdd.t138 3.9605
R22379 vdd.n21 vdd.t141 3.9605
R22380 vdd.n21 vdd.t137 3.9605
R22381 vdd.n20 vdd.t143 3.9605
R22382 vdd.n20 vdd.t134 3.9605
R22383 vdd.n15 vdd.t145 3.9605
R22384 vdd.n15 vdd.t144 3.9605
R22385 vdd.n16 vdd.t146 3.9605
R22386 vdd.n16 vdd.t132 3.9605
R22387 vdd.n18 vdd.t139 3.9605
R22388 vdd.n18 vdd.t136 3.9605
R22389 vdd.n25 vdd.t133 3.9605
R22390 vdd.n25 vdd.t135 3.9605
R22391 vdd.n2255 vdd.t121 3.74155
R22392 vdd.n874 vdd.t99 3.74155
R22393 vdd.n2837 vdd.t118 3.74155
R22394 vdd.n698 vdd.t107 3.74155
R22395 vdd.n7 vdd.t131 3.61217
R22396 vdd.n7 vdd.t95 3.61217
R22397 vdd.n8 vdd.t103 3.61217
R22398 vdd.n8 vdd.t123 3.61217
R22399 vdd.n10 vdd.t112 3.61217
R22400 vdd.n10 vdd.t83 3.61217
R22401 vdd.n12 vdd.t92 3.61217
R22402 vdd.n12 vdd.t110 3.61217
R22403 vdd.n5 vdd.t125 3.61217
R22404 vdd.n5 vdd.t105 3.61217
R22405 vdd.n3 vdd.t97 3.61217
R22406 vdd.n3 vdd.t127 3.61217
R22407 vdd.n1 vdd.t79 3.61217
R22408 vdd.n1 vdd.t116 3.61217
R22409 vdd.n0 vdd.t120 3.61217
R22410 vdd.n0 vdd.t101 3.61217
R22411 vdd.n292 vdd.n291 3.49141
R22412 vdd.n241 vdd.n240 3.49141
R22413 vdd.n198 vdd.n197 3.49141
R22414 vdd.n147 vdd.n146 3.49141
R22415 vdd.n105 vdd.n104 3.49141
R22416 vdd.n54 vdd.n53 3.49141
R22417 vdd.n1942 vdd.n1941 3.49141
R22418 vdd.n1993 vdd.n1992 3.49141
R22419 vdd.n1848 vdd.n1847 3.49141
R22420 vdd.n1899 vdd.n1898 3.49141
R22421 vdd.n1755 vdd.n1754 3.49141
R22422 vdd.n1806 vdd.n1805 3.49141
R22423 vdd.t115 vdd.n856 3.40145
R22424 vdd.n2496 vdd.t124 3.40145
R22425 vdd.n2800 vdd.t109 3.40145
R22426 vdd.n2825 vdd.t102 3.40145
R22427 vdd.n1702 vdd.t205 3.28809
R22428 vdd.n965 vdd.t5 3.28809
R22429 vdd.n2349 vdd.t50 3.28809
R22430 vdd.n2728 vdd.t57 3.28809
R22431 vdd.n2973 vdd.t1 3.28809
R22432 vdd.t186 vdd.n3426 3.28809
R22433 vdd.n1403 vdd.t150 3.06136
R22434 vdd.n2267 vdd.t89 3.06136
R22435 vdd.n1265 vdd.t128 3.06136
R22436 vdd.n2849 vdd.t117 3.06136
R22437 vdd.t113 vdd.n702 3.06136
R22438 vdd.t198 vdd.n3435 3.06136
R22439 vdd.n2342 vdd.t96 2.94799
R22440 vdd.t82 vdd.n774 2.94799
R22441 vdd.n2026 vdd.t156 2.83463
R22442 vdd.n3253 vdd.t165 2.83463
R22443 vdd.n295 vdd.n274 2.71565
R22444 vdd.n244 vdd.n223 2.71565
R22445 vdd.n201 vdd.n180 2.71565
R22446 vdd.n150 vdd.n129 2.71565
R22447 vdd.n108 vdd.n87 2.71565
R22448 vdd.n57 vdd.n36 2.71565
R22449 vdd.n1945 vdd.n1924 2.71565
R22450 vdd.n1996 vdd.n1975 2.71565
R22451 vdd.n1851 vdd.n1830 2.71565
R22452 vdd.n1902 vdd.n1881 2.71565
R22453 vdd.n1758 vdd.n1737 2.71565
R22454 vdd.n1809 vdd.n1788 2.71565
R22455 vdd.n2042 vdd.t177 2.6079
R22456 vdd.t200 vdd.n499 2.6079
R22457 vdd.n2316 vdd.t100 2.49453
R22458 vdd.n759 vdd.t130 2.49453
R22459 vdd.n282 vdd.n281 2.4129
R22460 vdd.n231 vdd.n230 2.4129
R22461 vdd.n188 vdd.n187 2.4129
R22462 vdd.n137 vdd.n136 2.4129
R22463 vdd.n95 vdd.n94 2.4129
R22464 vdd.n44 vdd.n43 2.4129
R22465 vdd.n1932 vdd.n1931 2.4129
R22466 vdd.n1983 vdd.n1982 2.4129
R22467 vdd.n1838 vdd.n1837 2.4129
R22468 vdd.n1889 vdd.n1888 2.4129
R22469 vdd.n1745 vdd.n1744 2.4129
R22470 vdd.n1796 vdd.n1795 2.4129
R22471 vdd.n2186 vdd.n1008 2.27742
R22472 vdd.n2186 vdd.n1007 2.27742
R22473 vdd.n3009 vdd.n522 2.27742
R22474 vdd.n3009 vdd.n521 2.27742
R22475 vdd.n3077 vdd.n608 2.27742
R22476 vdd.n3077 vdd.n606 2.27742
R22477 vdd.n2080 vdd.n2079 2.27742
R22478 vdd.n2079 vdd.n1344 2.27742
R22479 vdd.n911 vdd.t108 2.15444
R22480 vdd.n2292 vdd.t86 2.15444
R22481 vdd.n736 vdd.t85 2.15444
R22482 vdd.n2874 vdd.t84 2.15444
R22483 vdd.n296 vdd.n272 1.93989
R22484 vdd.n245 vdd.n221 1.93989
R22485 vdd.n202 vdd.n178 1.93989
R22486 vdd.n151 vdd.n127 1.93989
R22487 vdd.n109 vdd.n85 1.93989
R22488 vdd.n58 vdd.n34 1.93989
R22489 vdd.n1946 vdd.n1922 1.93989
R22490 vdd.n1997 vdd.n1973 1.93989
R22491 vdd.n1852 vdd.n1828 1.93989
R22492 vdd.n1903 vdd.n1879 1.93989
R22493 vdd.n1759 vdd.n1735 1.93989
R22494 vdd.n1810 vdd.n1786 1.93989
R22495 vdd.n1265 vdd.t119 1.81434
R22496 vdd.n2849 vdd.t94 1.81434
R22497 vdd.n1438 vdd.t37 1.47425
R22498 vdd.t23 vdd.n3411 1.47425
R22499 vdd.t126 vdd.n833 1.36088
R22500 vdd.n2807 vdd.t111 1.36088
R22501 vdd.t88 vdd.n908 1.24752
R22502 vdd.n2298 vdd.t93 1.24752
R22503 vdd.t98 vdd.n733 1.24752
R22504 vdd.n2880 vdd.t114 1.24752
R22505 vdd.n307 vdd.n267 1.16414
R22506 vdd.n300 vdd.n299 1.16414
R22507 vdd.n256 vdd.n216 1.16414
R22508 vdd.n249 vdd.n248 1.16414
R22509 vdd.n213 vdd.n173 1.16414
R22510 vdd.n206 vdd.n205 1.16414
R22511 vdd.n162 vdd.n122 1.16414
R22512 vdd.n155 vdd.n154 1.16414
R22513 vdd.n120 vdd.n80 1.16414
R22514 vdd.n113 vdd.n112 1.16414
R22515 vdd.n69 vdd.n29 1.16414
R22516 vdd.n62 vdd.n61 1.16414
R22517 vdd.n1957 vdd.n1917 1.16414
R22518 vdd.n1950 vdd.n1949 1.16414
R22519 vdd.n2008 vdd.n1968 1.16414
R22520 vdd.n2001 vdd.n2000 1.16414
R22521 vdd.n1863 vdd.n1823 1.16414
R22522 vdd.n1856 vdd.n1855 1.16414
R22523 vdd.n1914 vdd.n1874 1.16414
R22524 vdd.n1907 vdd.n1906 1.16414
R22525 vdd.n1770 vdd.n1730 1.16414
R22526 vdd.n1763 vdd.n1762 1.16414
R22527 vdd.n1821 vdd.n1781 1.16414
R22528 vdd.n1814 vdd.n1813 1.16414
R22529 vdd.n2011 vdd.n28 1.11236
R22530 vdd vdd.n3440 1.10453
R22531 vdd.n2034 vdd.t209 1.02079
R22532 vdd.t64 vdd.t86 1.02079
R22533 vdd.t85 vdd.t27 1.02079
R22534 vdd.n3244 vdd.t162 1.02079
R22535 vdd.n1568 vdd.n1567 0.970197
R22536 vdd.n2077 vdd.n2076 0.970197
R22537 vdd.n3296 vdd.n3295 0.970197
R22538 vdd.n3084 vdd.n3082 0.970197
R22539 vdd.n2322 vdd.t78 0.907421
R22540 vdd.n2710 vdd.t122 0.907421
R22541 vdd.t175 vdd.n1392 0.794056
R22542 vdd.n2061 vdd.t9 0.794056
R22543 vdd.t19 vdd.n511 0.794056
R22544 vdd.n481 vdd.t158 0.794056
R22545 vdd.n1711 vdd.t189 0.567326
R22546 vdd.n947 vdd.t81 0.567326
R22547 vdd.n2328 vdd.t77 0.567326
R22548 vdd.n2716 vdd.t80 0.567326
R22549 vdd.n2910 vdd.t90 0.567326
R22550 vdd.n3428 vdd.t152 0.567326
R22551 vdd.n2067 vdd.n1009 0.509646
R22552 vdd.n3209 vdd.n3208 0.509646
R22553 vdd.n3407 vdd.n3406 0.509646
R22554 vdd.n3289 vdd.n3288 0.509646
R22555 vdd.n3215 vdd.n514 0.509646
R22556 vdd.n2056 vdd.n1345 0.509646
R22557 vdd.n1673 vdd.n1435 0.509646
R22558 vdd.n1667 vdd.n1666 0.509646
R22559 vdd.n4 vdd.n2 0.459552
R22560 vdd.n11 vdd.n9 0.459552
R22561 vdd.n305 vdd.n304 0.388379
R22562 vdd.n271 vdd.n269 0.388379
R22563 vdd.n254 vdd.n253 0.388379
R22564 vdd.n220 vdd.n218 0.388379
R22565 vdd.n211 vdd.n210 0.388379
R22566 vdd.n177 vdd.n175 0.388379
R22567 vdd.n160 vdd.n159 0.388379
R22568 vdd.n126 vdd.n124 0.388379
R22569 vdd.n118 vdd.n117 0.388379
R22570 vdd.n84 vdd.n82 0.388379
R22571 vdd.n67 vdd.n66 0.388379
R22572 vdd.n33 vdd.n31 0.388379
R22573 vdd.n1955 vdd.n1954 0.388379
R22574 vdd.n1921 vdd.n1919 0.388379
R22575 vdd.n2006 vdd.n2005 0.388379
R22576 vdd.n1972 vdd.n1970 0.388379
R22577 vdd.n1861 vdd.n1860 0.388379
R22578 vdd.n1827 vdd.n1825 0.388379
R22579 vdd.n1912 vdd.n1911 0.388379
R22580 vdd.n1878 vdd.n1876 0.388379
R22581 vdd.n1768 vdd.n1767 0.388379
R22582 vdd.n1734 vdd.n1732 0.388379
R22583 vdd.n1819 vdd.n1818 0.388379
R22584 vdd.n1785 vdd.n1783 0.388379
R22585 vdd.n19 vdd.n17 0.387128
R22586 vdd.n24 vdd.n22 0.387128
R22587 vdd.n6 vdd.n4 0.358259
R22588 vdd.n13 vdd.n11 0.358259
R22589 vdd.n260 vdd.n258 0.358259
R22590 vdd.n262 vdd.n260 0.358259
R22591 vdd.n264 vdd.n262 0.358259
R22592 vdd.n266 vdd.n264 0.358259
R22593 vdd.n308 vdd.n266 0.358259
R22594 vdd.n166 vdd.n164 0.358259
R22595 vdd.n168 vdd.n166 0.358259
R22596 vdd.n170 vdd.n168 0.358259
R22597 vdd.n172 vdd.n170 0.358259
R22598 vdd.n214 vdd.n172 0.358259
R22599 vdd.n73 vdd.n71 0.358259
R22600 vdd.n75 vdd.n73 0.358259
R22601 vdd.n77 vdd.n75 0.358259
R22602 vdd.n79 vdd.n77 0.358259
R22603 vdd.n121 vdd.n79 0.358259
R22604 vdd.n2009 vdd.n1967 0.358259
R22605 vdd.n1967 vdd.n1965 0.358259
R22606 vdd.n1965 vdd.n1963 0.358259
R22607 vdd.n1963 vdd.n1961 0.358259
R22608 vdd.n1961 vdd.n1959 0.358259
R22609 vdd.n1915 vdd.n1873 0.358259
R22610 vdd.n1873 vdd.n1871 0.358259
R22611 vdd.n1871 vdd.n1869 0.358259
R22612 vdd.n1869 vdd.n1867 0.358259
R22613 vdd.n1867 vdd.n1865 0.358259
R22614 vdd.n1822 vdd.n1780 0.358259
R22615 vdd.n1780 vdd.n1778 0.358259
R22616 vdd.n1778 vdd.n1776 0.358259
R22617 vdd.n1776 vdd.n1774 0.358259
R22618 vdd.n1774 vdd.n1772 0.358259
R22619 vdd.t182 vdd.n1421 0.340595
R22620 vdd.n2261 vdd.t129 0.340595
R22621 vdd.n880 vdd.t87 0.340595
R22622 vdd.n2843 vdd.t76 0.340595
R22623 vdd.n705 vdd.t106 0.340595
R22624 vdd.n3419 vdd.t160 0.340595
R22625 vdd.n14 vdd.n6 0.334552
R22626 vdd.n14 vdd.n13 0.334552
R22627 vdd.n27 vdd.n19 0.21707
R22628 vdd.n27 vdd.n24 0.21707
R22629 vdd.n306 vdd.n268 0.155672
R22630 vdd.n298 vdd.n268 0.155672
R22631 vdd.n298 vdd.n297 0.155672
R22632 vdd.n297 vdd.n273 0.155672
R22633 vdd.n290 vdd.n273 0.155672
R22634 vdd.n290 vdd.n289 0.155672
R22635 vdd.n289 vdd.n277 0.155672
R22636 vdd.n282 vdd.n277 0.155672
R22637 vdd.n255 vdd.n217 0.155672
R22638 vdd.n247 vdd.n217 0.155672
R22639 vdd.n247 vdd.n246 0.155672
R22640 vdd.n246 vdd.n222 0.155672
R22641 vdd.n239 vdd.n222 0.155672
R22642 vdd.n239 vdd.n238 0.155672
R22643 vdd.n238 vdd.n226 0.155672
R22644 vdd.n231 vdd.n226 0.155672
R22645 vdd.n212 vdd.n174 0.155672
R22646 vdd.n204 vdd.n174 0.155672
R22647 vdd.n204 vdd.n203 0.155672
R22648 vdd.n203 vdd.n179 0.155672
R22649 vdd.n196 vdd.n179 0.155672
R22650 vdd.n196 vdd.n195 0.155672
R22651 vdd.n195 vdd.n183 0.155672
R22652 vdd.n188 vdd.n183 0.155672
R22653 vdd.n161 vdd.n123 0.155672
R22654 vdd.n153 vdd.n123 0.155672
R22655 vdd.n153 vdd.n152 0.155672
R22656 vdd.n152 vdd.n128 0.155672
R22657 vdd.n145 vdd.n128 0.155672
R22658 vdd.n145 vdd.n144 0.155672
R22659 vdd.n144 vdd.n132 0.155672
R22660 vdd.n137 vdd.n132 0.155672
R22661 vdd.n119 vdd.n81 0.155672
R22662 vdd.n111 vdd.n81 0.155672
R22663 vdd.n111 vdd.n110 0.155672
R22664 vdd.n110 vdd.n86 0.155672
R22665 vdd.n103 vdd.n86 0.155672
R22666 vdd.n103 vdd.n102 0.155672
R22667 vdd.n102 vdd.n90 0.155672
R22668 vdd.n95 vdd.n90 0.155672
R22669 vdd.n68 vdd.n30 0.155672
R22670 vdd.n60 vdd.n30 0.155672
R22671 vdd.n60 vdd.n59 0.155672
R22672 vdd.n59 vdd.n35 0.155672
R22673 vdd.n52 vdd.n35 0.155672
R22674 vdd.n52 vdd.n51 0.155672
R22675 vdd.n51 vdd.n39 0.155672
R22676 vdd.n44 vdd.n39 0.155672
R22677 vdd.n1956 vdd.n1918 0.155672
R22678 vdd.n1948 vdd.n1918 0.155672
R22679 vdd.n1948 vdd.n1947 0.155672
R22680 vdd.n1947 vdd.n1923 0.155672
R22681 vdd.n1940 vdd.n1923 0.155672
R22682 vdd.n1940 vdd.n1939 0.155672
R22683 vdd.n1939 vdd.n1927 0.155672
R22684 vdd.n1932 vdd.n1927 0.155672
R22685 vdd.n2007 vdd.n1969 0.155672
R22686 vdd.n1999 vdd.n1969 0.155672
R22687 vdd.n1999 vdd.n1998 0.155672
R22688 vdd.n1998 vdd.n1974 0.155672
R22689 vdd.n1991 vdd.n1974 0.155672
R22690 vdd.n1991 vdd.n1990 0.155672
R22691 vdd.n1990 vdd.n1978 0.155672
R22692 vdd.n1983 vdd.n1978 0.155672
R22693 vdd.n1862 vdd.n1824 0.155672
R22694 vdd.n1854 vdd.n1824 0.155672
R22695 vdd.n1854 vdd.n1853 0.155672
R22696 vdd.n1853 vdd.n1829 0.155672
R22697 vdd.n1846 vdd.n1829 0.155672
R22698 vdd.n1846 vdd.n1845 0.155672
R22699 vdd.n1845 vdd.n1833 0.155672
R22700 vdd.n1838 vdd.n1833 0.155672
R22701 vdd.n1913 vdd.n1875 0.155672
R22702 vdd.n1905 vdd.n1875 0.155672
R22703 vdd.n1905 vdd.n1904 0.155672
R22704 vdd.n1904 vdd.n1880 0.155672
R22705 vdd.n1897 vdd.n1880 0.155672
R22706 vdd.n1897 vdd.n1896 0.155672
R22707 vdd.n1896 vdd.n1884 0.155672
R22708 vdd.n1889 vdd.n1884 0.155672
R22709 vdd.n1769 vdd.n1731 0.155672
R22710 vdd.n1761 vdd.n1731 0.155672
R22711 vdd.n1761 vdd.n1760 0.155672
R22712 vdd.n1760 vdd.n1736 0.155672
R22713 vdd.n1753 vdd.n1736 0.155672
R22714 vdd.n1753 vdd.n1752 0.155672
R22715 vdd.n1752 vdd.n1740 0.155672
R22716 vdd.n1745 vdd.n1740 0.155672
R22717 vdd.n1820 vdd.n1782 0.155672
R22718 vdd.n1812 vdd.n1782 0.155672
R22719 vdd.n1812 vdd.n1811 0.155672
R22720 vdd.n1811 vdd.n1787 0.155672
R22721 vdd.n1804 vdd.n1787 0.155672
R22722 vdd.n1804 vdd.n1803 0.155672
R22723 vdd.n1803 vdd.n1791 0.155672
R22724 vdd.n1796 vdd.n1791 0.155672
R22725 vdd.n1014 vdd.n1006 0.152939
R22726 vdd.n1018 vdd.n1014 0.152939
R22727 vdd.n1019 vdd.n1018 0.152939
R22728 vdd.n1020 vdd.n1019 0.152939
R22729 vdd.n1021 vdd.n1020 0.152939
R22730 vdd.n1025 vdd.n1021 0.152939
R22731 vdd.n1026 vdd.n1025 0.152939
R22732 vdd.n1027 vdd.n1026 0.152939
R22733 vdd.n1028 vdd.n1027 0.152939
R22734 vdd.n1032 vdd.n1028 0.152939
R22735 vdd.n1033 vdd.n1032 0.152939
R22736 vdd.n1034 vdd.n1033 0.152939
R22737 vdd.n2150 vdd.n1034 0.152939
R22738 vdd.n2150 vdd.n2149 0.152939
R22739 vdd.n2149 vdd.n2148 0.152939
R22740 vdd.n2148 vdd.n1040 0.152939
R22741 vdd.n1045 vdd.n1040 0.152939
R22742 vdd.n1046 vdd.n1045 0.152939
R22743 vdd.n1047 vdd.n1046 0.152939
R22744 vdd.n1051 vdd.n1047 0.152939
R22745 vdd.n1052 vdd.n1051 0.152939
R22746 vdd.n1053 vdd.n1052 0.152939
R22747 vdd.n1054 vdd.n1053 0.152939
R22748 vdd.n1058 vdd.n1054 0.152939
R22749 vdd.n1059 vdd.n1058 0.152939
R22750 vdd.n1060 vdd.n1059 0.152939
R22751 vdd.n1061 vdd.n1060 0.152939
R22752 vdd.n1065 vdd.n1061 0.152939
R22753 vdd.n1066 vdd.n1065 0.152939
R22754 vdd.n1067 vdd.n1066 0.152939
R22755 vdd.n1068 vdd.n1067 0.152939
R22756 vdd.n1072 vdd.n1068 0.152939
R22757 vdd.n1073 vdd.n1072 0.152939
R22758 vdd.n1074 vdd.n1073 0.152939
R22759 vdd.n2111 vdd.n1074 0.152939
R22760 vdd.n2111 vdd.n2110 0.152939
R22761 vdd.n2110 vdd.n2109 0.152939
R22762 vdd.n2109 vdd.n1080 0.152939
R22763 vdd.n1085 vdd.n1080 0.152939
R22764 vdd.n1086 vdd.n1085 0.152939
R22765 vdd.n1087 vdd.n1086 0.152939
R22766 vdd.n1091 vdd.n1087 0.152939
R22767 vdd.n1092 vdd.n1091 0.152939
R22768 vdd.n1093 vdd.n1092 0.152939
R22769 vdd.n1094 vdd.n1093 0.152939
R22770 vdd.n1098 vdd.n1094 0.152939
R22771 vdd.n1099 vdd.n1098 0.152939
R22772 vdd.n1100 vdd.n1099 0.152939
R22773 vdd.n1101 vdd.n1100 0.152939
R22774 vdd.n1105 vdd.n1101 0.152939
R22775 vdd.n1106 vdd.n1105 0.152939
R22776 vdd.n2185 vdd.n1009 0.152939
R22777 vdd.n2014 vdd.n2013 0.152939
R22778 vdd.n2014 vdd.n1383 0.152939
R22779 vdd.n2029 vdd.n1383 0.152939
R22780 vdd.n2030 vdd.n2029 0.152939
R22781 vdd.n2031 vdd.n2030 0.152939
R22782 vdd.n2031 vdd.n1372 0.152939
R22783 vdd.n2046 vdd.n1372 0.152939
R22784 vdd.n2047 vdd.n2046 0.152939
R22785 vdd.n2048 vdd.n2047 0.152939
R22786 vdd.n2048 vdd.n1360 0.152939
R22787 vdd.n2065 vdd.n1360 0.152939
R22788 vdd.n2066 vdd.n2065 0.152939
R22789 vdd.n2067 vdd.n2066 0.152939
R22790 vdd.n527 vdd.n524 0.152939
R22791 vdd.n528 vdd.n527 0.152939
R22792 vdd.n529 vdd.n528 0.152939
R22793 vdd.n530 vdd.n529 0.152939
R22794 vdd.n533 vdd.n530 0.152939
R22795 vdd.n534 vdd.n533 0.152939
R22796 vdd.n535 vdd.n534 0.152939
R22797 vdd.n536 vdd.n535 0.152939
R22798 vdd.n539 vdd.n536 0.152939
R22799 vdd.n540 vdd.n539 0.152939
R22800 vdd.n541 vdd.n540 0.152939
R22801 vdd.n542 vdd.n541 0.152939
R22802 vdd.n547 vdd.n542 0.152939
R22803 vdd.n548 vdd.n547 0.152939
R22804 vdd.n549 vdd.n548 0.152939
R22805 vdd.n550 vdd.n549 0.152939
R22806 vdd.n553 vdd.n550 0.152939
R22807 vdd.n554 vdd.n553 0.152939
R22808 vdd.n555 vdd.n554 0.152939
R22809 vdd.n556 vdd.n555 0.152939
R22810 vdd.n559 vdd.n556 0.152939
R22811 vdd.n560 vdd.n559 0.152939
R22812 vdd.n561 vdd.n560 0.152939
R22813 vdd.n562 vdd.n561 0.152939
R22814 vdd.n565 vdd.n562 0.152939
R22815 vdd.n566 vdd.n565 0.152939
R22816 vdd.n567 vdd.n566 0.152939
R22817 vdd.n568 vdd.n567 0.152939
R22818 vdd.n571 vdd.n568 0.152939
R22819 vdd.n572 vdd.n571 0.152939
R22820 vdd.n573 vdd.n572 0.152939
R22821 vdd.n574 vdd.n573 0.152939
R22822 vdd.n577 vdd.n574 0.152939
R22823 vdd.n578 vdd.n577 0.152939
R22824 vdd.n3125 vdd.n578 0.152939
R22825 vdd.n3125 vdd.n3124 0.152939
R22826 vdd.n3124 vdd.n3123 0.152939
R22827 vdd.n3123 vdd.n582 0.152939
R22828 vdd.n587 vdd.n582 0.152939
R22829 vdd.n588 vdd.n587 0.152939
R22830 vdd.n591 vdd.n588 0.152939
R22831 vdd.n592 vdd.n591 0.152939
R22832 vdd.n593 vdd.n592 0.152939
R22833 vdd.n594 vdd.n593 0.152939
R22834 vdd.n597 vdd.n594 0.152939
R22835 vdd.n598 vdd.n597 0.152939
R22836 vdd.n599 vdd.n598 0.152939
R22837 vdd.n600 vdd.n599 0.152939
R22838 vdd.n603 vdd.n600 0.152939
R22839 vdd.n604 vdd.n603 0.152939
R22840 vdd.n605 vdd.n604 0.152939
R22841 vdd.n3208 vdd.n518 0.152939
R22842 vdd.n3209 vdd.n508 0.152939
R22843 vdd.n3223 vdd.n508 0.152939
R22844 vdd.n3224 vdd.n3223 0.152939
R22845 vdd.n3225 vdd.n3224 0.152939
R22846 vdd.n3225 vdd.n496 0.152939
R22847 vdd.n3239 vdd.n496 0.152939
R22848 vdd.n3240 vdd.n3239 0.152939
R22849 vdd.n3241 vdd.n3240 0.152939
R22850 vdd.n3241 vdd.n484 0.152939
R22851 vdd.n3256 vdd.n484 0.152939
R22852 vdd.n3257 vdd.n3256 0.152939
R22853 vdd.n3258 vdd.n3257 0.152939
R22854 vdd.n3258 vdd.n310 0.152939
R22855 vdd.n320 vdd.n311 0.152939
R22856 vdd.n321 vdd.n320 0.152939
R22857 vdd.n322 vdd.n321 0.152939
R22858 vdd.n331 vdd.n322 0.152939
R22859 vdd.n332 vdd.n331 0.152939
R22860 vdd.n333 vdd.n332 0.152939
R22861 vdd.n334 vdd.n333 0.152939
R22862 vdd.n342 vdd.n334 0.152939
R22863 vdd.n343 vdd.n342 0.152939
R22864 vdd.n344 vdd.n343 0.152939
R22865 vdd.n345 vdd.n344 0.152939
R22866 vdd.n353 vdd.n345 0.152939
R22867 vdd.n3407 vdd.n353 0.152939
R22868 vdd.n3406 vdd.n354 0.152939
R22869 vdd.n357 vdd.n354 0.152939
R22870 vdd.n361 vdd.n357 0.152939
R22871 vdd.n362 vdd.n361 0.152939
R22872 vdd.n363 vdd.n362 0.152939
R22873 vdd.n364 vdd.n363 0.152939
R22874 vdd.n365 vdd.n364 0.152939
R22875 vdd.n369 vdd.n365 0.152939
R22876 vdd.n370 vdd.n369 0.152939
R22877 vdd.n371 vdd.n370 0.152939
R22878 vdd.n372 vdd.n371 0.152939
R22879 vdd.n376 vdd.n372 0.152939
R22880 vdd.n377 vdd.n376 0.152939
R22881 vdd.n378 vdd.n377 0.152939
R22882 vdd.n379 vdd.n378 0.152939
R22883 vdd.n383 vdd.n379 0.152939
R22884 vdd.n384 vdd.n383 0.152939
R22885 vdd.n385 vdd.n384 0.152939
R22886 vdd.n3372 vdd.n385 0.152939
R22887 vdd.n3372 vdd.n3371 0.152939
R22888 vdd.n3371 vdd.n3370 0.152939
R22889 vdd.n3370 vdd.n391 0.152939
R22890 vdd.n396 vdd.n391 0.152939
R22891 vdd.n397 vdd.n396 0.152939
R22892 vdd.n398 vdd.n397 0.152939
R22893 vdd.n402 vdd.n398 0.152939
R22894 vdd.n403 vdd.n402 0.152939
R22895 vdd.n404 vdd.n403 0.152939
R22896 vdd.n405 vdd.n404 0.152939
R22897 vdd.n409 vdd.n405 0.152939
R22898 vdd.n410 vdd.n409 0.152939
R22899 vdd.n411 vdd.n410 0.152939
R22900 vdd.n412 vdd.n411 0.152939
R22901 vdd.n416 vdd.n412 0.152939
R22902 vdd.n417 vdd.n416 0.152939
R22903 vdd.n418 vdd.n417 0.152939
R22904 vdd.n419 vdd.n418 0.152939
R22905 vdd.n423 vdd.n419 0.152939
R22906 vdd.n424 vdd.n423 0.152939
R22907 vdd.n425 vdd.n424 0.152939
R22908 vdd.n3333 vdd.n425 0.152939
R22909 vdd.n3333 vdd.n3332 0.152939
R22910 vdd.n3332 vdd.n3331 0.152939
R22911 vdd.n3331 vdd.n431 0.152939
R22912 vdd.n436 vdd.n431 0.152939
R22913 vdd.n437 vdd.n436 0.152939
R22914 vdd.n438 vdd.n437 0.152939
R22915 vdd.n442 vdd.n438 0.152939
R22916 vdd.n443 vdd.n442 0.152939
R22917 vdd.n444 vdd.n443 0.152939
R22918 vdd.n445 vdd.n444 0.152939
R22919 vdd.n449 vdd.n445 0.152939
R22920 vdd.n450 vdd.n449 0.152939
R22921 vdd.n451 vdd.n450 0.152939
R22922 vdd.n452 vdd.n451 0.152939
R22923 vdd.n456 vdd.n452 0.152939
R22924 vdd.n457 vdd.n456 0.152939
R22925 vdd.n458 vdd.n457 0.152939
R22926 vdd.n459 vdd.n458 0.152939
R22927 vdd.n463 vdd.n459 0.152939
R22928 vdd.n464 vdd.n463 0.152939
R22929 vdd.n465 vdd.n464 0.152939
R22930 vdd.n3289 vdd.n465 0.152939
R22931 vdd.n3216 vdd.n3215 0.152939
R22932 vdd.n3217 vdd.n3216 0.152939
R22933 vdd.n3217 vdd.n502 0.152939
R22934 vdd.n3231 vdd.n502 0.152939
R22935 vdd.n3232 vdd.n3231 0.152939
R22936 vdd.n3233 vdd.n3232 0.152939
R22937 vdd.n3233 vdd.n489 0.152939
R22938 vdd.n3247 vdd.n489 0.152939
R22939 vdd.n3248 vdd.n3247 0.152939
R22940 vdd.n3249 vdd.n3248 0.152939
R22941 vdd.n3249 vdd.n477 0.152939
R22942 vdd.n3264 vdd.n477 0.152939
R22943 vdd.n3265 vdd.n3264 0.152939
R22944 vdd.n3266 vdd.n3265 0.152939
R22945 vdd.n3266 vdd.n475 0.152939
R22946 vdd.n3270 vdd.n475 0.152939
R22947 vdd.n3271 vdd.n3270 0.152939
R22948 vdd.n3272 vdd.n3271 0.152939
R22949 vdd.n3272 vdd.n472 0.152939
R22950 vdd.n3276 vdd.n472 0.152939
R22951 vdd.n3277 vdd.n3276 0.152939
R22952 vdd.n3278 vdd.n3277 0.152939
R22953 vdd.n3278 vdd.n469 0.152939
R22954 vdd.n3282 vdd.n469 0.152939
R22955 vdd.n3283 vdd.n3282 0.152939
R22956 vdd.n3284 vdd.n3283 0.152939
R22957 vdd.n3284 vdd.n466 0.152939
R22958 vdd.n3288 vdd.n466 0.152939
R22959 vdd.n3078 vdd.n514 0.152939
R22960 vdd.n2078 vdd.n1345 0.152939
R22961 vdd.n1674 vdd.n1673 0.152939
R22962 vdd.n1675 vdd.n1674 0.152939
R22963 vdd.n1675 vdd.n1424 0.152939
R22964 vdd.n1689 vdd.n1424 0.152939
R22965 vdd.n1690 vdd.n1689 0.152939
R22966 vdd.n1691 vdd.n1690 0.152939
R22967 vdd.n1691 vdd.n1411 0.152939
R22968 vdd.n1705 vdd.n1411 0.152939
R22969 vdd.n1706 vdd.n1705 0.152939
R22970 vdd.n1707 vdd.n1706 0.152939
R22971 vdd.n1707 vdd.n1400 0.152939
R22972 vdd.n1722 vdd.n1400 0.152939
R22973 vdd.n1723 vdd.n1722 0.152939
R22974 vdd.n1724 vdd.n1723 0.152939
R22975 vdd.n1724 vdd.n1389 0.152939
R22976 vdd.n2020 vdd.n1389 0.152939
R22977 vdd.n2021 vdd.n2020 0.152939
R22978 vdd.n2022 vdd.n2021 0.152939
R22979 vdd.n2022 vdd.n1377 0.152939
R22980 vdd.n2037 vdd.n1377 0.152939
R22981 vdd.n2038 vdd.n2037 0.152939
R22982 vdd.n2039 vdd.n2038 0.152939
R22983 vdd.n2039 vdd.n1367 0.152939
R22984 vdd.n2054 vdd.n1367 0.152939
R22985 vdd.n2055 vdd.n2054 0.152939
R22986 vdd.n2058 vdd.n2055 0.152939
R22987 vdd.n2058 vdd.n2057 0.152939
R22988 vdd.n2057 vdd.n2056 0.152939
R22989 vdd.n1666 vdd.n1440 0.152939
R22990 vdd.n1662 vdd.n1440 0.152939
R22991 vdd.n1662 vdd.n1661 0.152939
R22992 vdd.n1661 vdd.n1660 0.152939
R22993 vdd.n1660 vdd.n1445 0.152939
R22994 vdd.n1656 vdd.n1445 0.152939
R22995 vdd.n1656 vdd.n1655 0.152939
R22996 vdd.n1655 vdd.n1654 0.152939
R22997 vdd.n1654 vdd.n1453 0.152939
R22998 vdd.n1650 vdd.n1453 0.152939
R22999 vdd.n1650 vdd.n1649 0.152939
R23000 vdd.n1649 vdd.n1648 0.152939
R23001 vdd.n1648 vdd.n1461 0.152939
R23002 vdd.n1644 vdd.n1461 0.152939
R23003 vdd.n1644 vdd.n1643 0.152939
R23004 vdd.n1643 vdd.n1642 0.152939
R23005 vdd.n1642 vdd.n1469 0.152939
R23006 vdd.n1638 vdd.n1469 0.152939
R23007 vdd.n1638 vdd.n1637 0.152939
R23008 vdd.n1637 vdd.n1636 0.152939
R23009 vdd.n1636 vdd.n1479 0.152939
R23010 vdd.n1632 vdd.n1479 0.152939
R23011 vdd.n1632 vdd.n1631 0.152939
R23012 vdd.n1631 vdd.n1630 0.152939
R23013 vdd.n1630 vdd.n1487 0.152939
R23014 vdd.n1626 vdd.n1487 0.152939
R23015 vdd.n1626 vdd.n1625 0.152939
R23016 vdd.n1625 vdd.n1624 0.152939
R23017 vdd.n1624 vdd.n1495 0.152939
R23018 vdd.n1620 vdd.n1495 0.152939
R23019 vdd.n1620 vdd.n1619 0.152939
R23020 vdd.n1619 vdd.n1618 0.152939
R23021 vdd.n1618 vdd.n1503 0.152939
R23022 vdd.n1614 vdd.n1503 0.152939
R23023 vdd.n1614 vdd.n1613 0.152939
R23024 vdd.n1613 vdd.n1612 0.152939
R23025 vdd.n1612 vdd.n1511 0.152939
R23026 vdd.n1608 vdd.n1511 0.152939
R23027 vdd.n1608 vdd.n1607 0.152939
R23028 vdd.n1607 vdd.n1606 0.152939
R23029 vdd.n1606 vdd.n1519 0.152939
R23030 vdd.n1526 vdd.n1519 0.152939
R23031 vdd.n1596 vdd.n1526 0.152939
R23032 vdd.n1596 vdd.n1595 0.152939
R23033 vdd.n1595 vdd.n1594 0.152939
R23034 vdd.n1594 vdd.n1527 0.152939
R23035 vdd.n1590 vdd.n1527 0.152939
R23036 vdd.n1590 vdd.n1589 0.152939
R23037 vdd.n1589 vdd.n1588 0.152939
R23038 vdd.n1588 vdd.n1534 0.152939
R23039 vdd.n1584 vdd.n1534 0.152939
R23040 vdd.n1584 vdd.n1583 0.152939
R23041 vdd.n1583 vdd.n1582 0.152939
R23042 vdd.n1582 vdd.n1542 0.152939
R23043 vdd.n1578 vdd.n1542 0.152939
R23044 vdd.n1578 vdd.n1577 0.152939
R23045 vdd.n1577 vdd.n1576 0.152939
R23046 vdd.n1576 vdd.n1550 0.152939
R23047 vdd.n1572 vdd.n1550 0.152939
R23048 vdd.n1572 vdd.n1571 0.152939
R23049 vdd.n1571 vdd.n1570 0.152939
R23050 vdd.n1570 vdd.n1558 0.152939
R23051 vdd.n1558 vdd.n1435 0.152939
R23052 vdd.n1667 vdd.n1430 0.152939
R23053 vdd.n1681 vdd.n1430 0.152939
R23054 vdd.n1682 vdd.n1681 0.152939
R23055 vdd.n1683 vdd.n1682 0.152939
R23056 vdd.n1683 vdd.n1418 0.152939
R23057 vdd.n1697 vdd.n1418 0.152939
R23058 vdd.n1698 vdd.n1697 0.152939
R23059 vdd.n1699 vdd.n1698 0.152939
R23060 vdd.n1699 vdd.n1406 0.152939
R23061 vdd.n1714 vdd.n1406 0.152939
R23062 vdd.n1715 vdd.n1714 0.152939
R23063 vdd.n1716 vdd.n1715 0.152939
R23064 vdd.n1716 vdd.n1395 0.152939
R23065 vdd.n2013 vdd.n2012 0.145814
R23066 vdd.n3439 vdd.n310 0.145814
R23067 vdd.n3439 vdd.n311 0.145814
R23068 vdd.n2012 vdd.n1395 0.145814
R23069 vdd.n2186 vdd.n2185 0.110256
R23070 vdd.n3009 vdd.n518 0.110256
R23071 vdd.n3078 vdd.n3077 0.110256
R23072 vdd.n2079 vdd.n2078 0.110256
R23073 vdd.n2186 vdd.n1006 0.0431829
R23074 vdd.n2079 vdd.n1106 0.0431829
R23075 vdd.n3009 vdd.n524 0.0431829
R23076 vdd.n3077 vdd.n605 0.0431829
R23077 vdd vdd.n28 0.00833333
R23078 a_n2804_13878.n2 a_n2804_13878.n0 98.9633
R23079 a_n2804_13878.n5 a_n2804_13878.n3 98.7517
R23080 a_n2804_13878.n25 a_n2804_13878.n24 98.6055
R23081 a_n2804_13878.n27 a_n2804_13878.n26 98.6055
R23082 a_n2804_13878.n2 a_n2804_13878.n1 98.6055
R23083 a_n2804_13878.n13 a_n2804_13878.n12 98.6055
R23084 a_n2804_13878.n11 a_n2804_13878.n10 98.6055
R23085 a_n2804_13878.n9 a_n2804_13878.n8 98.6055
R23086 a_n2804_13878.n7 a_n2804_13878.n6 98.6055
R23087 a_n2804_13878.n5 a_n2804_13878.n4 98.6055
R23088 a_n2804_13878.n29 a_n2804_13878.n28 98.6054
R23089 a_n2804_13878.n23 a_n2804_13878.n22 98.6054
R23090 a_n2804_13878.n15 a_n2804_13878.t1 74.6477
R23091 a_n2804_13878.n20 a_n2804_13878.t2 74.2899
R23092 a_n2804_13878.n17 a_n2804_13878.t3 74.2899
R23093 a_n2804_13878.n16 a_n2804_13878.t0 74.2899
R23094 a_n2804_13878.n19 a_n2804_13878.n18 70.6783
R23095 a_n2804_13878.n15 a_n2804_13878.n14 70.6783
R23096 a_n2804_13878.n21 a_n2804_13878.n13 15.7159
R23097 a_n2804_13878.n23 a_n2804_13878.n21 12.6495
R23098 a_n2804_13878.n21 a_n2804_13878.n20 8.38735
R23099 a_n2804_13878.n22 a_n2804_13878.t15 3.61217
R23100 a_n2804_13878.n22 a_n2804_13878.t24 3.61217
R23101 a_n2804_13878.n24 a_n2804_13878.t28 3.61217
R23102 a_n2804_13878.n24 a_n2804_13878.t14 3.61217
R23103 a_n2804_13878.n26 a_n2804_13878.t18 3.61217
R23104 a_n2804_13878.n26 a_n2804_13878.t19 3.61217
R23105 a_n2804_13878.n1 a_n2804_13878.t8 3.61217
R23106 a_n2804_13878.n1 a_n2804_13878.t20 3.61217
R23107 a_n2804_13878.n0 a_n2804_13878.t25 3.61217
R23108 a_n2804_13878.n0 a_n2804_13878.t31 3.61217
R23109 a_n2804_13878.n18 a_n2804_13878.t6 3.61217
R23110 a_n2804_13878.n18 a_n2804_13878.t7 3.61217
R23111 a_n2804_13878.n14 a_n2804_13878.t4 3.61217
R23112 a_n2804_13878.n14 a_n2804_13878.t5 3.61217
R23113 a_n2804_13878.n12 a_n2804_13878.t21 3.61217
R23114 a_n2804_13878.n12 a_n2804_13878.t9 3.61217
R23115 a_n2804_13878.n10 a_n2804_13878.t26 3.61217
R23116 a_n2804_13878.n10 a_n2804_13878.t11 3.61217
R23117 a_n2804_13878.n8 a_n2804_13878.t10 3.61217
R23118 a_n2804_13878.n8 a_n2804_13878.t13 3.61217
R23119 a_n2804_13878.n6 a_n2804_13878.t23 3.61217
R23120 a_n2804_13878.n6 a_n2804_13878.t16 3.61217
R23121 a_n2804_13878.n4 a_n2804_13878.t27 3.61217
R23122 a_n2804_13878.n4 a_n2804_13878.t17 3.61217
R23123 a_n2804_13878.n3 a_n2804_13878.t12 3.61217
R23124 a_n2804_13878.n3 a_n2804_13878.t22 3.61217
R23125 a_n2804_13878.n29 a_n2804_13878.t29 3.61217
R23126 a_n2804_13878.t30 a_n2804_13878.n29 3.61217
R23127 a_n2804_13878.n16 a_n2804_13878.n15 0.358259
R23128 a_n2804_13878.n19 a_n2804_13878.n17 0.358259
R23129 a_n2804_13878.n20 a_n2804_13878.n19 0.358259
R23130 a_n2804_13878.n28 a_n2804_13878.n2 0.358259
R23131 a_n2804_13878.n28 a_n2804_13878.n27 0.358259
R23132 a_n2804_13878.n27 a_n2804_13878.n25 0.358259
R23133 a_n2804_13878.n25 a_n2804_13878.n23 0.358259
R23134 a_n2804_13878.n7 a_n2804_13878.n5 0.146627
R23135 a_n2804_13878.n9 a_n2804_13878.n7 0.146627
R23136 a_n2804_13878.n11 a_n2804_13878.n9 0.146627
R23137 a_n2804_13878.n13 a_n2804_13878.n11 0.146627
R23138 a_n2804_13878.n17 a_n2804_13878.n16 0.101793
R23139 a_n2982_8322.n12 a_n2982_8322.t3 74.6477
R23140 a_n2982_8322.n1 a_n2982_8322.t14 74.6477
R23141 a_n2982_8322.n28 a_n2982_8322.t29 74.6474
R23142 a_n2982_8322.n20 a_n2982_8322.t9 74.2899
R23143 a_n2982_8322.n13 a_n2982_8322.t1 74.2899
R23144 a_n2982_8322.n14 a_n2982_8322.t4 74.2899
R23145 a_n2982_8322.n17 a_n2982_8322.t5 74.2899
R23146 a_n2982_8322.n10 a_n2982_8322.t8 74.2899
R23147 a_n2982_8322.n28 a_n2982_8322.n27 70.6783
R23148 a_n2982_8322.n26 a_n2982_8322.n25 70.6783
R23149 a_n2982_8322.n24 a_n2982_8322.n23 70.6783
R23150 a_n2982_8322.n22 a_n2982_8322.n21 70.6783
R23151 a_n2982_8322.n12 a_n2982_8322.n11 70.6783
R23152 a_n2982_8322.n16 a_n2982_8322.n15 70.6783
R23153 a_n2982_8322.n1 a_n2982_8322.n0 70.6783
R23154 a_n2982_8322.n3 a_n2982_8322.n2 70.6783
R23155 a_n2982_8322.n5 a_n2982_8322.n4 70.6783
R23156 a_n2982_8322.n7 a_n2982_8322.n6 70.6783
R23157 a_n2982_8322.n9 a_n2982_8322.n8 70.6783
R23158 a_n2982_8322.n30 a_n2982_8322.n29 70.6782
R23159 a_n2982_8322.n18 a_n2982_8322.n10 24.9022
R23160 a_n2982_8322.n19 a_n2982_8322.t33 9.65181
R23161 a_n2982_8322.n18 a_n2982_8322.n17 8.38735
R23162 a_n2982_8322.n20 a_n2982_8322.n19 6.90998
R23163 a_n2982_8322.n19 a_n2982_8322.n18 5.3452
R23164 a_n2982_8322.n27 a_n2982_8322.t22 3.61217
R23165 a_n2982_8322.n27 a_n2982_8322.t18 3.61217
R23166 a_n2982_8322.n25 a_n2982_8322.t28 3.61217
R23167 a_n2982_8322.n25 a_n2982_8322.t16 3.61217
R23168 a_n2982_8322.n23 a_n2982_8322.t13 3.61217
R23169 a_n2982_8322.n23 a_n2982_8322.t12 3.61217
R23170 a_n2982_8322.n21 a_n2982_8322.t26 3.61217
R23171 a_n2982_8322.n21 a_n2982_8322.t25 3.61217
R23172 a_n2982_8322.n11 a_n2982_8322.t7 3.61217
R23173 a_n2982_8322.n11 a_n2982_8322.t6 3.61217
R23174 a_n2982_8322.n15 a_n2982_8322.t2 3.61217
R23175 a_n2982_8322.n15 a_n2982_8322.t0 3.61217
R23176 a_n2982_8322.n0 a_n2982_8322.t27 3.61217
R23177 a_n2982_8322.n0 a_n2982_8322.t23 3.61217
R23178 a_n2982_8322.n2 a_n2982_8322.t30 3.61217
R23179 a_n2982_8322.n2 a_n2982_8322.t20 3.61217
R23180 a_n2982_8322.n4 a_n2982_8322.t11 3.61217
R23181 a_n2982_8322.n4 a_n2982_8322.t10 3.61217
R23182 a_n2982_8322.n6 a_n2982_8322.t24 3.61217
R23183 a_n2982_8322.n6 a_n2982_8322.t17 3.61217
R23184 a_n2982_8322.n8 a_n2982_8322.t21 3.61217
R23185 a_n2982_8322.n8 a_n2982_8322.t19 3.61217
R23186 a_n2982_8322.n30 a_n2982_8322.t15 3.61217
R23187 a_n2982_8322.t31 a_n2982_8322.n30 3.61217
R23188 a_n2982_8322.n17 a_n2982_8322.n16 0.358259
R23189 a_n2982_8322.n16 a_n2982_8322.n14 0.358259
R23190 a_n2982_8322.n13 a_n2982_8322.n12 0.358259
R23191 a_n2982_8322.n10 a_n2982_8322.n9 0.358259
R23192 a_n2982_8322.n9 a_n2982_8322.n7 0.358259
R23193 a_n2982_8322.n7 a_n2982_8322.n5 0.358259
R23194 a_n2982_8322.n5 a_n2982_8322.n3 0.358259
R23195 a_n2982_8322.n3 a_n2982_8322.n1 0.358259
R23196 a_n2982_8322.n22 a_n2982_8322.n20 0.358259
R23197 a_n2982_8322.n24 a_n2982_8322.n22 0.358259
R23198 a_n2982_8322.n26 a_n2982_8322.n24 0.358259
R23199 a_n2982_8322.n29 a_n2982_8322.n26 0.358259
R23200 a_n2982_8322.n29 a_n2982_8322.n28 0.358259
R23201 a_n2982_8322.n14 a_n2982_8322.n13 0.101793
R23202 a_n2982_8322.t36 a_n2982_8322.t34 0.0788333
R23203 a_n2982_8322.t32 a_n2982_8322.t37 0.0788333
R23204 a_n2982_8322.t33 a_n2982_8322.t35 0.0788333
R23205 a_n2982_8322.t32 a_n2982_8322.t36 0.0318333
R23206 a_n2982_8322.t33 a_n2982_8322.t37 0.0318333
R23207 a_n2982_8322.t34 a_n2982_8322.t37 0.0318333
R23208 a_n2982_8322.t35 a_n2982_8322.t32 0.0318333
R23209 output.n41 output.n15 289.615
R23210 output.n72 output.n46 289.615
R23211 output.n104 output.n78 289.615
R23212 output.n136 output.n110 289.615
R23213 output.n77 output.n45 197.26
R23214 output.n77 output.n76 196.298
R23215 output.n109 output.n108 196.298
R23216 output.n141 output.n140 196.298
R23217 output.n42 output.n41 185
R23218 output.n40 output.n39 185
R23219 output.n19 output.n18 185
R23220 output.n34 output.n33 185
R23221 output.n32 output.n31 185
R23222 output.n23 output.n22 185
R23223 output.n26 output.n25 185
R23224 output.n73 output.n72 185
R23225 output.n71 output.n70 185
R23226 output.n50 output.n49 185
R23227 output.n65 output.n64 185
R23228 output.n63 output.n62 185
R23229 output.n54 output.n53 185
R23230 output.n57 output.n56 185
R23231 output.n105 output.n104 185
R23232 output.n103 output.n102 185
R23233 output.n82 output.n81 185
R23234 output.n97 output.n96 185
R23235 output.n95 output.n94 185
R23236 output.n86 output.n85 185
R23237 output.n89 output.n88 185
R23238 output.n137 output.n136 185
R23239 output.n135 output.n134 185
R23240 output.n114 output.n113 185
R23241 output.n129 output.n128 185
R23242 output.n127 output.n126 185
R23243 output.n118 output.n117 185
R23244 output.n121 output.n120 185
R23245 output.t19 output.n24 147.661
R23246 output.t1 output.n55 147.661
R23247 output.t2 output.n87 147.661
R23248 output.t0 output.n119 147.661
R23249 output.n41 output.n40 104.615
R23250 output.n40 output.n18 104.615
R23251 output.n33 output.n18 104.615
R23252 output.n33 output.n32 104.615
R23253 output.n32 output.n22 104.615
R23254 output.n25 output.n22 104.615
R23255 output.n72 output.n71 104.615
R23256 output.n71 output.n49 104.615
R23257 output.n64 output.n49 104.615
R23258 output.n64 output.n63 104.615
R23259 output.n63 output.n53 104.615
R23260 output.n56 output.n53 104.615
R23261 output.n104 output.n103 104.615
R23262 output.n103 output.n81 104.615
R23263 output.n96 output.n81 104.615
R23264 output.n96 output.n95 104.615
R23265 output.n95 output.n85 104.615
R23266 output.n88 output.n85 104.615
R23267 output.n136 output.n135 104.615
R23268 output.n135 output.n113 104.615
R23269 output.n128 output.n113 104.615
R23270 output.n128 output.n127 104.615
R23271 output.n127 output.n117 104.615
R23272 output.n120 output.n117 104.615
R23273 output.n1 output.t4 77.056
R23274 output.n14 output.t6 76.6694
R23275 output.n1 output.n0 72.7095
R23276 output.n3 output.n2 72.7095
R23277 output.n5 output.n4 72.7095
R23278 output.n7 output.n6 72.7095
R23279 output.n9 output.n8 72.7095
R23280 output.n11 output.n10 72.7095
R23281 output.n13 output.n12 72.7095
R23282 output.n25 output.t19 52.3082
R23283 output.n56 output.t1 52.3082
R23284 output.n88 output.t2 52.3082
R23285 output.n120 output.t0 52.3082
R23286 output.n26 output.n24 15.6674
R23287 output.n57 output.n55 15.6674
R23288 output.n89 output.n87 15.6674
R23289 output.n121 output.n119 15.6674
R23290 output.n27 output.n23 12.8005
R23291 output.n58 output.n54 12.8005
R23292 output.n90 output.n86 12.8005
R23293 output.n122 output.n118 12.8005
R23294 output.n31 output.n30 12.0247
R23295 output.n62 output.n61 12.0247
R23296 output.n94 output.n93 12.0247
R23297 output.n126 output.n125 12.0247
R23298 output.n34 output.n21 11.249
R23299 output.n65 output.n52 11.249
R23300 output.n97 output.n84 11.249
R23301 output.n129 output.n116 11.249
R23302 output.n35 output.n19 10.4732
R23303 output.n66 output.n50 10.4732
R23304 output.n98 output.n82 10.4732
R23305 output.n130 output.n114 10.4732
R23306 output.n39 output.n38 9.69747
R23307 output.n70 output.n69 9.69747
R23308 output.n102 output.n101 9.69747
R23309 output.n134 output.n133 9.69747
R23310 output.n45 output.n44 9.45567
R23311 output.n76 output.n75 9.45567
R23312 output.n108 output.n107 9.45567
R23313 output.n140 output.n139 9.45567
R23314 output.n44 output.n43 9.3005
R23315 output.n17 output.n16 9.3005
R23316 output.n38 output.n37 9.3005
R23317 output.n36 output.n35 9.3005
R23318 output.n21 output.n20 9.3005
R23319 output.n30 output.n29 9.3005
R23320 output.n28 output.n27 9.3005
R23321 output.n75 output.n74 9.3005
R23322 output.n48 output.n47 9.3005
R23323 output.n69 output.n68 9.3005
R23324 output.n67 output.n66 9.3005
R23325 output.n52 output.n51 9.3005
R23326 output.n61 output.n60 9.3005
R23327 output.n59 output.n58 9.3005
R23328 output.n107 output.n106 9.3005
R23329 output.n80 output.n79 9.3005
R23330 output.n101 output.n100 9.3005
R23331 output.n99 output.n98 9.3005
R23332 output.n84 output.n83 9.3005
R23333 output.n93 output.n92 9.3005
R23334 output.n91 output.n90 9.3005
R23335 output.n139 output.n138 9.3005
R23336 output.n112 output.n111 9.3005
R23337 output.n133 output.n132 9.3005
R23338 output.n131 output.n130 9.3005
R23339 output.n116 output.n115 9.3005
R23340 output.n125 output.n124 9.3005
R23341 output.n123 output.n122 9.3005
R23342 output.n42 output.n17 8.92171
R23343 output.n73 output.n48 8.92171
R23344 output.n105 output.n80 8.92171
R23345 output.n137 output.n112 8.92171
R23346 output output.n141 8.15037
R23347 output.n43 output.n15 8.14595
R23348 output.n74 output.n46 8.14595
R23349 output.n106 output.n78 8.14595
R23350 output.n138 output.n110 8.14595
R23351 output.n45 output.n15 5.81868
R23352 output.n76 output.n46 5.81868
R23353 output.n108 output.n78 5.81868
R23354 output.n140 output.n110 5.81868
R23355 output.n43 output.n42 5.04292
R23356 output.n74 output.n73 5.04292
R23357 output.n106 output.n105 5.04292
R23358 output.n138 output.n137 5.04292
R23359 output.n28 output.n24 4.38594
R23360 output.n59 output.n55 4.38594
R23361 output.n91 output.n87 4.38594
R23362 output.n123 output.n119 4.38594
R23363 output.n39 output.n17 4.26717
R23364 output.n70 output.n48 4.26717
R23365 output.n102 output.n80 4.26717
R23366 output.n134 output.n112 4.26717
R23367 output.n0 output.t10 3.9605
R23368 output.n0 output.t15 3.9605
R23369 output.n2 output.t3 3.9605
R23370 output.n2 output.t11 3.9605
R23371 output.n4 output.t13 3.9605
R23372 output.n4 output.t12 3.9605
R23373 output.n6 output.t18 3.9605
R23374 output.n6 output.t5 3.9605
R23375 output.n8 output.t7 3.9605
R23376 output.n8 output.t16 3.9605
R23377 output.n10 output.t17 3.9605
R23378 output.n10 output.t8 3.9605
R23379 output.n12 output.t9 3.9605
R23380 output.n12 output.t14 3.9605
R23381 output.n38 output.n19 3.49141
R23382 output.n69 output.n50 3.49141
R23383 output.n101 output.n82 3.49141
R23384 output.n133 output.n114 3.49141
R23385 output.n35 output.n34 2.71565
R23386 output.n66 output.n65 2.71565
R23387 output.n98 output.n97 2.71565
R23388 output.n130 output.n129 2.71565
R23389 output.n31 output.n21 1.93989
R23390 output.n62 output.n52 1.93989
R23391 output.n94 output.n84 1.93989
R23392 output.n126 output.n116 1.93989
R23393 output.n30 output.n23 1.16414
R23394 output.n61 output.n54 1.16414
R23395 output.n93 output.n86 1.16414
R23396 output.n125 output.n118 1.16414
R23397 output.n141 output.n109 0.962709
R23398 output.n109 output.n77 0.962709
R23399 output.n27 output.n26 0.388379
R23400 output.n58 output.n57 0.388379
R23401 output.n90 output.n89 0.388379
R23402 output.n122 output.n121 0.388379
R23403 output.n14 output.n13 0.387128
R23404 output.n13 output.n11 0.387128
R23405 output.n11 output.n9 0.387128
R23406 output.n9 output.n7 0.387128
R23407 output.n7 output.n5 0.387128
R23408 output.n5 output.n3 0.387128
R23409 output.n3 output.n1 0.387128
R23410 output.n44 output.n16 0.155672
R23411 output.n37 output.n16 0.155672
R23412 output.n37 output.n36 0.155672
R23413 output.n36 output.n20 0.155672
R23414 output.n29 output.n20 0.155672
R23415 output.n29 output.n28 0.155672
R23416 output.n75 output.n47 0.155672
R23417 output.n68 output.n47 0.155672
R23418 output.n68 output.n67 0.155672
R23419 output.n67 output.n51 0.155672
R23420 output.n60 output.n51 0.155672
R23421 output.n60 output.n59 0.155672
R23422 output.n107 output.n79 0.155672
R23423 output.n100 output.n79 0.155672
R23424 output.n100 output.n99 0.155672
R23425 output.n99 output.n83 0.155672
R23426 output.n92 output.n83 0.155672
R23427 output.n92 output.n91 0.155672
R23428 output.n139 output.n111 0.155672
R23429 output.n132 output.n111 0.155672
R23430 output.n132 output.n131 0.155672
R23431 output.n131 output.n115 0.155672
R23432 output.n124 output.n115 0.155672
R23433 output.n124 output.n123 0.155672
R23434 output output.n14 0.126227
R23435 minus.n33 minus.t20 321.495
R23436 minus.n7 minus.t6 321.495
R23437 minus.n50 minus.t18 297.12
R23438 minus.n48 minus.t15 297.12
R23439 minus.n28 minus.t16 297.12
R23440 minus.n42 minus.t11 297.12
R23441 minus.n30 minus.t12 297.12
R23442 minus.n36 minus.t7 297.12
R23443 minus.n32 minus.t19 297.12
R23444 minus.n6 minus.t5 297.12
R23445 minus.n10 minus.t9 297.12
R23446 minus.n12 minus.t8 297.12
R23447 minus.n16 minus.t10 297.12
R23448 minus.n18 minus.t14 297.12
R23449 minus.n22 minus.t13 297.12
R23450 minus.n24 minus.t17 297.12
R23451 minus.n56 minus.t4 243.255
R23452 minus.n55 minus.n53 224.169
R23453 minus.n55 minus.n54 223.454
R23454 minus.n35 minus.n34 161.3
R23455 minus.n36 minus.n31 161.3
R23456 minus.n38 minus.n37 161.3
R23457 minus.n39 minus.n30 161.3
R23458 minus.n41 minus.n40 161.3
R23459 minus.n42 minus.n29 161.3
R23460 minus.n44 minus.n43 161.3
R23461 minus.n45 minus.n28 161.3
R23462 minus.n47 minus.n46 161.3
R23463 minus.n48 minus.n27 161.3
R23464 minus.n49 minus.n26 161.3
R23465 minus.n51 minus.n50 161.3
R23466 minus.n25 minus.n24 161.3
R23467 minus.n23 minus.n0 161.3
R23468 minus.n22 minus.n21 161.3
R23469 minus.n20 minus.n1 161.3
R23470 minus.n19 minus.n18 161.3
R23471 minus.n17 minus.n2 161.3
R23472 minus.n16 minus.n15 161.3
R23473 minus.n14 minus.n3 161.3
R23474 minus.n13 minus.n12 161.3
R23475 minus.n11 minus.n4 161.3
R23476 minus.n10 minus.n9 161.3
R23477 minus.n8 minus.n5 161.3
R23478 minus.n8 minus.n7 44.9377
R23479 minus.n34 minus.n33 44.9377
R23480 minus.n50 minus.n49 37.246
R23481 minus.n24 minus.n23 37.246
R23482 minus.n48 minus.n47 32.8641
R23483 minus.n35 minus.n32 32.8641
R23484 minus.n6 minus.n5 32.8641
R23485 minus.n22 minus.n1 32.8641
R23486 minus.n52 minus.n51 30.2486
R23487 minus.n43 minus.n28 28.4823
R23488 minus.n37 minus.n36 28.4823
R23489 minus.n11 minus.n10 28.4823
R23490 minus.n18 minus.n17 28.4823
R23491 minus.n42 minus.n41 24.1005
R23492 minus.n41 minus.n30 24.1005
R23493 minus.n12 minus.n3 24.1005
R23494 minus.n16 minus.n3 24.1005
R23495 minus.n54 minus.t3 19.8005
R23496 minus.n54 minus.t2 19.8005
R23497 minus.n53 minus.t1 19.8005
R23498 minus.n53 minus.t0 19.8005
R23499 minus.n43 minus.n42 19.7187
R23500 minus.n37 minus.n30 19.7187
R23501 minus.n12 minus.n11 19.7187
R23502 minus.n17 minus.n16 19.7187
R23503 minus.n33 minus.n32 17.0522
R23504 minus.n7 minus.n6 17.0522
R23505 minus.n47 minus.n28 15.3369
R23506 minus.n36 minus.n35 15.3369
R23507 minus.n10 minus.n5 15.3369
R23508 minus.n18 minus.n1 15.3369
R23509 minus.n52 minus.n25 12.0706
R23510 minus minus.n57 11.6687
R23511 minus.n49 minus.n48 10.955
R23512 minus.n23 minus.n22 10.955
R23513 minus.n57 minus.n56 4.80222
R23514 minus.n57 minus.n52 0.972091
R23515 minus.n56 minus.n55 0.716017
R23516 minus.n51 minus.n26 0.189894
R23517 minus.n27 minus.n26 0.189894
R23518 minus.n46 minus.n27 0.189894
R23519 minus.n46 minus.n45 0.189894
R23520 minus.n45 minus.n44 0.189894
R23521 minus.n44 minus.n29 0.189894
R23522 minus.n40 minus.n29 0.189894
R23523 minus.n40 minus.n39 0.189894
R23524 minus.n39 minus.n38 0.189894
R23525 minus.n38 minus.n31 0.189894
R23526 minus.n34 minus.n31 0.189894
R23527 minus.n9 minus.n8 0.189894
R23528 minus.n9 minus.n4 0.189894
R23529 minus.n13 minus.n4 0.189894
R23530 minus.n14 minus.n13 0.189894
R23531 minus.n15 minus.n14 0.189894
R23532 minus.n15 minus.n2 0.189894
R23533 minus.n19 minus.n2 0.189894
R23534 minus.n20 minus.n19 0.189894
R23535 minus.n21 minus.n20 0.189894
R23536 minus.n21 minus.n0 0.189894
R23537 minus.n25 minus.n0 0.189894
R23538 diffpairibias.n0 diffpairibias.t18 436.822
R23539 diffpairibias.n21 diffpairibias.t19 435.479
R23540 diffpairibias.n20 diffpairibias.t16 435.479
R23541 diffpairibias.n19 diffpairibias.t17 435.479
R23542 diffpairibias.n18 diffpairibias.t21 435.479
R23543 diffpairibias.n0 diffpairibias.t22 435.479
R23544 diffpairibias.n1 diffpairibias.t20 435.479
R23545 diffpairibias.n2 diffpairibias.t23 435.479
R23546 diffpairibias.n10 diffpairibias.t0 377.536
R23547 diffpairibias.n10 diffpairibias.t8 376.193
R23548 diffpairibias.n11 diffpairibias.t10 376.193
R23549 diffpairibias.n12 diffpairibias.t6 376.193
R23550 diffpairibias.n13 diffpairibias.t2 376.193
R23551 diffpairibias.n14 diffpairibias.t12 376.193
R23552 diffpairibias.n15 diffpairibias.t4 376.193
R23553 diffpairibias.n16 diffpairibias.t14 376.193
R23554 diffpairibias.n3 diffpairibias.t1 113.368
R23555 diffpairibias.n3 diffpairibias.t9 112.698
R23556 diffpairibias.n4 diffpairibias.t11 112.698
R23557 diffpairibias.n5 diffpairibias.t7 112.698
R23558 diffpairibias.n6 diffpairibias.t3 112.698
R23559 diffpairibias.n7 diffpairibias.t13 112.698
R23560 diffpairibias.n8 diffpairibias.t5 112.698
R23561 diffpairibias.n9 diffpairibias.t15 112.698
R23562 diffpairibias.n17 diffpairibias.n16 4.77242
R23563 diffpairibias.n17 diffpairibias.n9 4.30807
R23564 diffpairibias.n18 diffpairibias.n17 4.13945
R23565 diffpairibias.n16 diffpairibias.n15 1.34352
R23566 diffpairibias.n15 diffpairibias.n14 1.34352
R23567 diffpairibias.n14 diffpairibias.n13 1.34352
R23568 diffpairibias.n13 diffpairibias.n12 1.34352
R23569 diffpairibias.n12 diffpairibias.n11 1.34352
R23570 diffpairibias.n11 diffpairibias.n10 1.34352
R23571 diffpairibias.n2 diffpairibias.n1 1.34352
R23572 diffpairibias.n1 diffpairibias.n0 1.34352
R23573 diffpairibias.n19 diffpairibias.n18 1.34352
R23574 diffpairibias.n20 diffpairibias.n19 1.34352
R23575 diffpairibias.n21 diffpairibias.n20 1.34352
R23576 diffpairibias.n22 diffpairibias.n21 0.862419
R23577 diffpairibias diffpairibias.n22 0.684875
R23578 diffpairibias.n9 diffpairibias.n8 0.672012
R23579 diffpairibias.n8 diffpairibias.n7 0.672012
R23580 diffpairibias.n7 diffpairibias.n6 0.672012
R23581 diffpairibias.n6 diffpairibias.n5 0.672012
R23582 diffpairibias.n5 diffpairibias.n4 0.672012
R23583 diffpairibias.n4 diffpairibias.n3 0.672012
R23584 diffpairibias.n22 diffpairibias.n2 0.190907
R23585 outputibias.n27 outputibias.n1 289.615
R23586 outputibias.n58 outputibias.n32 289.615
R23587 outputibias.n90 outputibias.n64 289.615
R23588 outputibias.n122 outputibias.n96 289.615
R23589 outputibias.n28 outputibias.n27 185
R23590 outputibias.n26 outputibias.n25 185
R23591 outputibias.n5 outputibias.n4 185
R23592 outputibias.n20 outputibias.n19 185
R23593 outputibias.n18 outputibias.n17 185
R23594 outputibias.n9 outputibias.n8 185
R23595 outputibias.n12 outputibias.n11 185
R23596 outputibias.n59 outputibias.n58 185
R23597 outputibias.n57 outputibias.n56 185
R23598 outputibias.n36 outputibias.n35 185
R23599 outputibias.n51 outputibias.n50 185
R23600 outputibias.n49 outputibias.n48 185
R23601 outputibias.n40 outputibias.n39 185
R23602 outputibias.n43 outputibias.n42 185
R23603 outputibias.n91 outputibias.n90 185
R23604 outputibias.n89 outputibias.n88 185
R23605 outputibias.n68 outputibias.n67 185
R23606 outputibias.n83 outputibias.n82 185
R23607 outputibias.n81 outputibias.n80 185
R23608 outputibias.n72 outputibias.n71 185
R23609 outputibias.n75 outputibias.n74 185
R23610 outputibias.n123 outputibias.n122 185
R23611 outputibias.n121 outputibias.n120 185
R23612 outputibias.n100 outputibias.n99 185
R23613 outputibias.n115 outputibias.n114 185
R23614 outputibias.n113 outputibias.n112 185
R23615 outputibias.n104 outputibias.n103 185
R23616 outputibias.n107 outputibias.n106 185
R23617 outputibias.n0 outputibias.t10 178.945
R23618 outputibias.n133 outputibias.t8 177.018
R23619 outputibias.n132 outputibias.t11 177.018
R23620 outputibias.n0 outputibias.t9 177.018
R23621 outputibias.t7 outputibias.n10 147.661
R23622 outputibias.t1 outputibias.n41 147.661
R23623 outputibias.t3 outputibias.n73 147.661
R23624 outputibias.t5 outputibias.n105 147.661
R23625 outputibias.n128 outputibias.t6 132.363
R23626 outputibias.n128 outputibias.t0 130.436
R23627 outputibias.n129 outputibias.t2 130.436
R23628 outputibias.n130 outputibias.t4 130.436
R23629 outputibias.n27 outputibias.n26 104.615
R23630 outputibias.n26 outputibias.n4 104.615
R23631 outputibias.n19 outputibias.n4 104.615
R23632 outputibias.n19 outputibias.n18 104.615
R23633 outputibias.n18 outputibias.n8 104.615
R23634 outputibias.n11 outputibias.n8 104.615
R23635 outputibias.n58 outputibias.n57 104.615
R23636 outputibias.n57 outputibias.n35 104.615
R23637 outputibias.n50 outputibias.n35 104.615
R23638 outputibias.n50 outputibias.n49 104.615
R23639 outputibias.n49 outputibias.n39 104.615
R23640 outputibias.n42 outputibias.n39 104.615
R23641 outputibias.n90 outputibias.n89 104.615
R23642 outputibias.n89 outputibias.n67 104.615
R23643 outputibias.n82 outputibias.n67 104.615
R23644 outputibias.n82 outputibias.n81 104.615
R23645 outputibias.n81 outputibias.n71 104.615
R23646 outputibias.n74 outputibias.n71 104.615
R23647 outputibias.n122 outputibias.n121 104.615
R23648 outputibias.n121 outputibias.n99 104.615
R23649 outputibias.n114 outputibias.n99 104.615
R23650 outputibias.n114 outputibias.n113 104.615
R23651 outputibias.n113 outputibias.n103 104.615
R23652 outputibias.n106 outputibias.n103 104.615
R23653 outputibias.n63 outputibias.n31 95.6354
R23654 outputibias.n63 outputibias.n62 94.6732
R23655 outputibias.n95 outputibias.n94 94.6732
R23656 outputibias.n127 outputibias.n126 94.6732
R23657 outputibias.n11 outputibias.t7 52.3082
R23658 outputibias.n42 outputibias.t1 52.3082
R23659 outputibias.n74 outputibias.t3 52.3082
R23660 outputibias.n106 outputibias.t5 52.3082
R23661 outputibias.n12 outputibias.n10 15.6674
R23662 outputibias.n43 outputibias.n41 15.6674
R23663 outputibias.n75 outputibias.n73 15.6674
R23664 outputibias.n107 outputibias.n105 15.6674
R23665 outputibias.n13 outputibias.n9 12.8005
R23666 outputibias.n44 outputibias.n40 12.8005
R23667 outputibias.n76 outputibias.n72 12.8005
R23668 outputibias.n108 outputibias.n104 12.8005
R23669 outputibias.n17 outputibias.n16 12.0247
R23670 outputibias.n48 outputibias.n47 12.0247
R23671 outputibias.n80 outputibias.n79 12.0247
R23672 outputibias.n112 outputibias.n111 12.0247
R23673 outputibias.n20 outputibias.n7 11.249
R23674 outputibias.n51 outputibias.n38 11.249
R23675 outputibias.n83 outputibias.n70 11.249
R23676 outputibias.n115 outputibias.n102 11.249
R23677 outputibias.n21 outputibias.n5 10.4732
R23678 outputibias.n52 outputibias.n36 10.4732
R23679 outputibias.n84 outputibias.n68 10.4732
R23680 outputibias.n116 outputibias.n100 10.4732
R23681 outputibias.n25 outputibias.n24 9.69747
R23682 outputibias.n56 outputibias.n55 9.69747
R23683 outputibias.n88 outputibias.n87 9.69747
R23684 outputibias.n120 outputibias.n119 9.69747
R23685 outputibias.n31 outputibias.n30 9.45567
R23686 outputibias.n62 outputibias.n61 9.45567
R23687 outputibias.n94 outputibias.n93 9.45567
R23688 outputibias.n126 outputibias.n125 9.45567
R23689 outputibias.n30 outputibias.n29 9.3005
R23690 outputibias.n3 outputibias.n2 9.3005
R23691 outputibias.n24 outputibias.n23 9.3005
R23692 outputibias.n22 outputibias.n21 9.3005
R23693 outputibias.n7 outputibias.n6 9.3005
R23694 outputibias.n16 outputibias.n15 9.3005
R23695 outputibias.n14 outputibias.n13 9.3005
R23696 outputibias.n61 outputibias.n60 9.3005
R23697 outputibias.n34 outputibias.n33 9.3005
R23698 outputibias.n55 outputibias.n54 9.3005
R23699 outputibias.n53 outputibias.n52 9.3005
R23700 outputibias.n38 outputibias.n37 9.3005
R23701 outputibias.n47 outputibias.n46 9.3005
R23702 outputibias.n45 outputibias.n44 9.3005
R23703 outputibias.n93 outputibias.n92 9.3005
R23704 outputibias.n66 outputibias.n65 9.3005
R23705 outputibias.n87 outputibias.n86 9.3005
R23706 outputibias.n85 outputibias.n84 9.3005
R23707 outputibias.n70 outputibias.n69 9.3005
R23708 outputibias.n79 outputibias.n78 9.3005
R23709 outputibias.n77 outputibias.n76 9.3005
R23710 outputibias.n125 outputibias.n124 9.3005
R23711 outputibias.n98 outputibias.n97 9.3005
R23712 outputibias.n119 outputibias.n118 9.3005
R23713 outputibias.n117 outputibias.n116 9.3005
R23714 outputibias.n102 outputibias.n101 9.3005
R23715 outputibias.n111 outputibias.n110 9.3005
R23716 outputibias.n109 outputibias.n108 9.3005
R23717 outputibias.n28 outputibias.n3 8.92171
R23718 outputibias.n59 outputibias.n34 8.92171
R23719 outputibias.n91 outputibias.n66 8.92171
R23720 outputibias.n123 outputibias.n98 8.92171
R23721 outputibias.n29 outputibias.n1 8.14595
R23722 outputibias.n60 outputibias.n32 8.14595
R23723 outputibias.n92 outputibias.n64 8.14595
R23724 outputibias.n124 outputibias.n96 8.14595
R23725 outputibias.n31 outputibias.n1 5.81868
R23726 outputibias.n62 outputibias.n32 5.81868
R23727 outputibias.n94 outputibias.n64 5.81868
R23728 outputibias.n126 outputibias.n96 5.81868
R23729 outputibias.n131 outputibias.n130 5.20947
R23730 outputibias.n29 outputibias.n28 5.04292
R23731 outputibias.n60 outputibias.n59 5.04292
R23732 outputibias.n92 outputibias.n91 5.04292
R23733 outputibias.n124 outputibias.n123 5.04292
R23734 outputibias.n131 outputibias.n127 4.42209
R23735 outputibias.n14 outputibias.n10 4.38594
R23736 outputibias.n45 outputibias.n41 4.38594
R23737 outputibias.n77 outputibias.n73 4.38594
R23738 outputibias.n109 outputibias.n105 4.38594
R23739 outputibias.n132 outputibias.n131 4.28454
R23740 outputibias.n25 outputibias.n3 4.26717
R23741 outputibias.n56 outputibias.n34 4.26717
R23742 outputibias.n88 outputibias.n66 4.26717
R23743 outputibias.n120 outputibias.n98 4.26717
R23744 outputibias.n24 outputibias.n5 3.49141
R23745 outputibias.n55 outputibias.n36 3.49141
R23746 outputibias.n87 outputibias.n68 3.49141
R23747 outputibias.n119 outputibias.n100 3.49141
R23748 outputibias.n21 outputibias.n20 2.71565
R23749 outputibias.n52 outputibias.n51 2.71565
R23750 outputibias.n84 outputibias.n83 2.71565
R23751 outputibias.n116 outputibias.n115 2.71565
R23752 outputibias.n17 outputibias.n7 1.93989
R23753 outputibias.n48 outputibias.n38 1.93989
R23754 outputibias.n80 outputibias.n70 1.93989
R23755 outputibias.n112 outputibias.n102 1.93989
R23756 outputibias.n130 outputibias.n129 1.9266
R23757 outputibias.n129 outputibias.n128 1.9266
R23758 outputibias.n133 outputibias.n132 1.92658
R23759 outputibias.n134 outputibias.n133 1.29913
R23760 outputibias.n16 outputibias.n9 1.16414
R23761 outputibias.n47 outputibias.n40 1.16414
R23762 outputibias.n79 outputibias.n72 1.16414
R23763 outputibias.n111 outputibias.n104 1.16414
R23764 outputibias.n127 outputibias.n95 0.962709
R23765 outputibias.n95 outputibias.n63 0.962709
R23766 outputibias.n13 outputibias.n12 0.388379
R23767 outputibias.n44 outputibias.n43 0.388379
R23768 outputibias.n76 outputibias.n75 0.388379
R23769 outputibias.n108 outputibias.n107 0.388379
R23770 outputibias.n134 outputibias.n0 0.337251
R23771 outputibias outputibias.n134 0.302375
R23772 outputibias.n30 outputibias.n2 0.155672
R23773 outputibias.n23 outputibias.n2 0.155672
R23774 outputibias.n23 outputibias.n22 0.155672
R23775 outputibias.n22 outputibias.n6 0.155672
R23776 outputibias.n15 outputibias.n6 0.155672
R23777 outputibias.n15 outputibias.n14 0.155672
R23778 outputibias.n61 outputibias.n33 0.155672
R23779 outputibias.n54 outputibias.n33 0.155672
R23780 outputibias.n54 outputibias.n53 0.155672
R23781 outputibias.n53 outputibias.n37 0.155672
R23782 outputibias.n46 outputibias.n37 0.155672
R23783 outputibias.n46 outputibias.n45 0.155672
R23784 outputibias.n93 outputibias.n65 0.155672
R23785 outputibias.n86 outputibias.n65 0.155672
R23786 outputibias.n86 outputibias.n85 0.155672
R23787 outputibias.n85 outputibias.n69 0.155672
R23788 outputibias.n78 outputibias.n69 0.155672
R23789 outputibias.n78 outputibias.n77 0.155672
R23790 outputibias.n125 outputibias.n97 0.155672
R23791 outputibias.n118 outputibias.n97 0.155672
R23792 outputibias.n118 outputibias.n117 0.155672
R23793 outputibias.n117 outputibias.n101 0.155672
R23794 outputibias.n110 outputibias.n101 0.155672
R23795 outputibias.n110 outputibias.n109 0.155672
C0 commonsourceibias outputibias 0.003832f
C1 plus diffpairibias 3.12e-19
C2 vdd commonsourceibias 0.004218f
C3 CSoutput plus 0.843035f
C4 commonsourceibias diffpairibias 0.06482f
C5 CSoutput commonsourceibias 54.0646f
C6 minus plus 8.857121f
C7 minus commonsourceibias 0.318966f
C8 plus commonsourceibias 0.273048f
C9 output outputibias 2.34152f
C10 vdd output 7.23429f
C11 CSoutput output 6.13881f
C12 CSoutput outputibias 0.032386f
C13 vdd CSoutput 92.9043f
C14 minus diffpairibias 3.1e-19
C15 commonsourceibias output 0.006808f
C16 CSoutput minus 2.8659f
C17 vdd plus 0.08312f
C18 diffpairibias gnd 48.980038f
C19 outputibias gnd 32.465668f
C20 output gnd 15.47879f
C21 commonsourceibias gnd 0.18355p
C22 plus gnd 30.930847f
C23 minus gnd 26.23274f
C24 CSoutput gnd 0.124759p
C25 vdd gnd 0.479896p
C26 outputibias.t9 gnd 0.11477f
C27 outputibias.t10 gnd 0.115567f
C28 outputibias.n0 gnd 0.130108f
C29 outputibias.n1 gnd 0.001372f
C30 outputibias.n2 gnd 9.76e-19
C31 outputibias.n3 gnd 5.24e-19
C32 outputibias.n4 gnd 0.001239f
C33 outputibias.n5 gnd 5.55e-19
C34 outputibias.n6 gnd 9.76e-19
C35 outputibias.n7 gnd 5.24e-19
C36 outputibias.n8 gnd 0.001239f
C37 outputibias.n9 gnd 5.55e-19
C38 outputibias.n10 gnd 0.004176f
C39 outputibias.t7 gnd 0.00202f
C40 outputibias.n11 gnd 9.3e-19
C41 outputibias.n12 gnd 7.32e-19
C42 outputibias.n13 gnd 5.24e-19
C43 outputibias.n14 gnd 0.02322f
C44 outputibias.n15 gnd 9.76e-19
C45 outputibias.n16 gnd 5.24e-19
C46 outputibias.n17 gnd 5.55e-19
C47 outputibias.n18 gnd 0.001239f
C48 outputibias.n19 gnd 0.001239f
C49 outputibias.n20 gnd 5.55e-19
C50 outputibias.n21 gnd 5.24e-19
C51 outputibias.n22 gnd 9.76e-19
C52 outputibias.n23 gnd 9.76e-19
C53 outputibias.n24 gnd 5.24e-19
C54 outputibias.n25 gnd 5.55e-19
C55 outputibias.n26 gnd 0.001239f
C56 outputibias.n27 gnd 0.002683f
C57 outputibias.n28 gnd 5.55e-19
C58 outputibias.n29 gnd 5.24e-19
C59 outputibias.n30 gnd 0.002256f
C60 outputibias.n31 gnd 0.005781f
C61 outputibias.n32 gnd 0.001372f
C62 outputibias.n33 gnd 9.76e-19
C63 outputibias.n34 gnd 5.24e-19
C64 outputibias.n35 gnd 0.001239f
C65 outputibias.n36 gnd 5.55e-19
C66 outputibias.n37 gnd 9.76e-19
C67 outputibias.n38 gnd 5.24e-19
C68 outputibias.n39 gnd 0.001239f
C69 outputibias.n40 gnd 5.55e-19
C70 outputibias.n41 gnd 0.004176f
C71 outputibias.t1 gnd 0.00202f
C72 outputibias.n42 gnd 9.3e-19
C73 outputibias.n43 gnd 7.32e-19
C74 outputibias.n44 gnd 5.24e-19
C75 outputibias.n45 gnd 0.02322f
C76 outputibias.n46 gnd 9.76e-19
C77 outputibias.n47 gnd 5.24e-19
C78 outputibias.n48 gnd 5.55e-19
C79 outputibias.n49 gnd 0.001239f
C80 outputibias.n50 gnd 0.001239f
C81 outputibias.n51 gnd 5.55e-19
C82 outputibias.n52 gnd 5.24e-19
C83 outputibias.n53 gnd 9.76e-19
C84 outputibias.n54 gnd 9.76e-19
C85 outputibias.n55 gnd 5.24e-19
C86 outputibias.n56 gnd 5.55e-19
C87 outputibias.n57 gnd 0.001239f
C88 outputibias.n58 gnd 0.002683f
C89 outputibias.n59 gnd 5.55e-19
C90 outputibias.n60 gnd 5.24e-19
C91 outputibias.n61 gnd 0.002256f
C92 outputibias.n62 gnd 0.005197f
C93 outputibias.n63 gnd 0.121892f
C94 outputibias.n64 gnd 0.001372f
C95 outputibias.n65 gnd 9.76e-19
C96 outputibias.n66 gnd 5.24e-19
C97 outputibias.n67 gnd 0.001239f
C98 outputibias.n68 gnd 5.55e-19
C99 outputibias.n69 gnd 9.76e-19
C100 outputibias.n70 gnd 5.24e-19
C101 outputibias.n71 gnd 0.001239f
C102 outputibias.n72 gnd 5.55e-19
C103 outputibias.n73 gnd 0.004176f
C104 outputibias.t3 gnd 0.00202f
C105 outputibias.n74 gnd 9.3e-19
C106 outputibias.n75 gnd 7.32e-19
C107 outputibias.n76 gnd 5.24e-19
C108 outputibias.n77 gnd 0.02322f
C109 outputibias.n78 gnd 9.76e-19
C110 outputibias.n79 gnd 5.24e-19
C111 outputibias.n80 gnd 5.55e-19
C112 outputibias.n81 gnd 0.001239f
C113 outputibias.n82 gnd 0.001239f
C114 outputibias.n83 gnd 5.55e-19
C115 outputibias.n84 gnd 5.24e-19
C116 outputibias.n85 gnd 9.76e-19
C117 outputibias.n86 gnd 9.76e-19
C118 outputibias.n87 gnd 5.24e-19
C119 outputibias.n88 gnd 5.55e-19
C120 outputibias.n89 gnd 0.001239f
C121 outputibias.n90 gnd 0.002683f
C122 outputibias.n91 gnd 5.55e-19
C123 outputibias.n92 gnd 5.24e-19
C124 outputibias.n93 gnd 0.002256f
C125 outputibias.n94 gnd 0.005197f
C126 outputibias.n95 gnd 0.064513f
C127 outputibias.n96 gnd 0.001372f
C128 outputibias.n97 gnd 9.76e-19
C129 outputibias.n98 gnd 5.24e-19
C130 outputibias.n99 gnd 0.001239f
C131 outputibias.n100 gnd 5.55e-19
C132 outputibias.n101 gnd 9.76e-19
C133 outputibias.n102 gnd 5.24e-19
C134 outputibias.n103 gnd 0.001239f
C135 outputibias.n104 gnd 5.55e-19
C136 outputibias.n105 gnd 0.004176f
C137 outputibias.t5 gnd 0.00202f
C138 outputibias.n106 gnd 9.3e-19
C139 outputibias.n107 gnd 7.32e-19
C140 outputibias.n108 gnd 5.24e-19
C141 outputibias.n109 gnd 0.02322f
C142 outputibias.n110 gnd 9.76e-19
C143 outputibias.n111 gnd 5.24e-19
C144 outputibias.n112 gnd 5.55e-19
C145 outputibias.n113 gnd 0.001239f
C146 outputibias.n114 gnd 0.001239f
C147 outputibias.n115 gnd 5.55e-19
C148 outputibias.n116 gnd 5.24e-19
C149 outputibias.n117 gnd 9.76e-19
C150 outputibias.n118 gnd 9.76e-19
C151 outputibias.n119 gnd 5.24e-19
C152 outputibias.n120 gnd 5.55e-19
C153 outputibias.n121 gnd 0.001239f
C154 outputibias.n122 gnd 0.002683f
C155 outputibias.n123 gnd 5.55e-19
C156 outputibias.n124 gnd 5.24e-19
C157 outputibias.n125 gnd 0.002256f
C158 outputibias.n126 gnd 0.005197f
C159 outputibias.n127 gnd 0.084814f
C160 outputibias.t4 gnd 0.108319f
C161 outputibias.t2 gnd 0.108319f
C162 outputibias.t0 gnd 0.108319f
C163 outputibias.t6 gnd 0.109238f
C164 outputibias.n128 gnd 0.134674f
C165 outputibias.n129 gnd 0.07244f
C166 outputibias.n130 gnd 0.079818f
C167 outputibias.n131 gnd 0.164901f
C168 outputibias.t11 gnd 0.11477f
C169 outputibias.n132 gnd 0.067481f
C170 outputibias.t8 gnd 0.11477f
C171 outputibias.n133 gnd 0.065115f
C172 outputibias.n134 gnd 0.029159f
C173 diffpairibias.t18 gnd 0.087401f
C174 diffpairibias.t22 gnd 0.087239f
C175 diffpairibias.n0 gnd 0.102784f
C176 diffpairibias.t20 gnd 0.087239f
C177 diffpairibias.n1 gnd 0.050171f
C178 diffpairibias.t23 gnd 0.087239f
C179 diffpairibias.n2 gnd 0.039841f
C180 diffpairibias.t1 gnd 0.083757f
C181 diffpairibias.t9 gnd 0.083392f
C182 diffpairibias.n3 gnd 0.131682f
C183 diffpairibias.t11 gnd 0.083392f
C184 diffpairibias.n4 gnd 0.07027f
C185 diffpairibias.t7 gnd 0.083392f
C186 diffpairibias.n5 gnd 0.07027f
C187 diffpairibias.t3 gnd 0.083392f
C188 diffpairibias.n6 gnd 0.07027f
C189 diffpairibias.t13 gnd 0.083392f
C190 diffpairibias.n7 gnd 0.07027f
C191 diffpairibias.t5 gnd 0.083392f
C192 diffpairibias.n8 gnd 0.07027f
C193 diffpairibias.t15 gnd 0.083392f
C194 diffpairibias.n9 gnd 0.099771f
C195 diffpairibias.t0 gnd 0.08427f
C196 diffpairibias.t8 gnd 0.084123f
C197 diffpairibias.n10 gnd 0.091784f
C198 diffpairibias.t10 gnd 0.084123f
C199 diffpairibias.n11 gnd 0.050681f
C200 diffpairibias.t6 gnd 0.084123f
C201 diffpairibias.n12 gnd 0.050681f
C202 diffpairibias.t2 gnd 0.084123f
C203 diffpairibias.n13 gnd 0.050681f
C204 diffpairibias.t12 gnd 0.084123f
C205 diffpairibias.n14 gnd 0.050681f
C206 diffpairibias.t4 gnd 0.084123f
C207 diffpairibias.n15 gnd 0.050681f
C208 diffpairibias.t14 gnd 0.084123f
C209 diffpairibias.n16 gnd 0.059977f
C210 diffpairibias.n17 gnd 0.226448f
C211 diffpairibias.t21 gnd 0.087239f
C212 diffpairibias.n18 gnd 0.050181f
C213 diffpairibias.t17 gnd 0.087239f
C214 diffpairibias.n19 gnd 0.050171f
C215 diffpairibias.t16 gnd 0.087239f
C216 diffpairibias.n20 gnd 0.050171f
C217 diffpairibias.t19 gnd 0.087239f
C218 diffpairibias.n21 gnd 0.045859f
C219 diffpairibias.n22 gnd 0.046268f
C220 minus.n0 gnd 0.03095f
C221 minus.n1 gnd 0.007023f
C222 minus.n2 gnd 0.03095f
C223 minus.n3 gnd 0.007023f
C224 minus.n4 gnd 0.03095f
C225 minus.n5 gnd 0.007023f
C226 minus.t6 gnd 0.452513f
C227 minus.t5 gnd 0.43776f
C228 minus.n6 gnd 0.198707f
C229 minus.n7 gnd 0.182289f
C230 minus.n8 gnd 0.130973f
C231 minus.n9 gnd 0.03095f
C232 minus.t9 gnd 0.43776f
C233 minus.n10 gnd 0.194467f
C234 minus.n11 gnd 0.007023f
C235 minus.t8 gnd 0.43776f
C236 minus.n12 gnd 0.194467f
C237 minus.n13 gnd 0.03095f
C238 minus.n14 gnd 0.03095f
C239 minus.n15 gnd 0.03095f
C240 minus.t10 gnd 0.43776f
C241 minus.n16 gnd 0.194467f
C242 minus.n17 gnd 0.007023f
C243 minus.t14 gnd 0.43776f
C244 minus.n18 gnd 0.194467f
C245 minus.n19 gnd 0.03095f
C246 minus.n20 gnd 0.03095f
C247 minus.n21 gnd 0.03095f
C248 minus.t13 gnd 0.43776f
C249 minus.n22 gnd 0.194467f
C250 minus.n23 gnd 0.007023f
C251 minus.t17 gnd 0.43776f
C252 minus.n24 gnd 0.193608f
C253 minus.n25 gnd 0.356775f
C254 minus.n26 gnd 0.03095f
C255 minus.t18 gnd 0.43776f
C256 minus.t15 gnd 0.43776f
C257 minus.n27 gnd 0.03095f
C258 minus.t16 gnd 0.43776f
C259 minus.n28 gnd 0.194467f
C260 minus.n29 gnd 0.03095f
C261 minus.t11 gnd 0.43776f
C262 minus.t12 gnd 0.43776f
C263 minus.n30 gnd 0.194467f
C264 minus.n31 gnd 0.03095f
C265 minus.t7 gnd 0.43776f
C266 minus.t19 gnd 0.43776f
C267 minus.n32 gnd 0.198707f
C268 minus.t20 gnd 0.452513f
C269 minus.n33 gnd 0.182289f
C270 minus.n34 gnd 0.130973f
C271 minus.n35 gnd 0.007023f
C272 minus.n36 gnd 0.194467f
C273 minus.n37 gnd 0.007023f
C274 minus.n38 gnd 0.03095f
C275 minus.n39 gnd 0.03095f
C276 minus.n40 gnd 0.03095f
C277 minus.n41 gnd 0.007023f
C278 minus.n42 gnd 0.194467f
C279 minus.n43 gnd 0.007023f
C280 minus.n44 gnd 0.03095f
C281 minus.n45 gnd 0.03095f
C282 minus.n46 gnd 0.03095f
C283 minus.n47 gnd 0.007023f
C284 minus.n48 gnd 0.194467f
C285 minus.n49 gnd 0.007023f
C286 minus.n50 gnd 0.193608f
C287 minus.n51 gnd 0.898329f
C288 minus.n52 gnd 1.36603f
C289 minus.t1 gnd 0.009541f
C290 minus.t0 gnd 0.009541f
C291 minus.n53 gnd 0.031373f
C292 minus.t3 gnd 0.009541f
C293 minus.t2 gnd 0.009541f
C294 minus.n54 gnd 0.030943f
C295 minus.n55 gnd 0.264085f
C296 minus.t4 gnd 0.053104f
C297 minus.n56 gnd 0.144109f
C298 minus.n57 gnd 2.03109f
C299 output.t4 gnd 0.464308f
C300 output.t10 gnd 0.044422f
C301 output.t15 gnd 0.044422f
C302 output.n0 gnd 0.364624f
C303 output.n1 gnd 0.614102f
C304 output.t3 gnd 0.044422f
C305 output.t11 gnd 0.044422f
C306 output.n2 gnd 0.364624f
C307 output.n3 gnd 0.350265f
C308 output.t13 gnd 0.044422f
C309 output.t12 gnd 0.044422f
C310 output.n4 gnd 0.364624f
C311 output.n5 gnd 0.350265f
C312 output.t18 gnd 0.044422f
C313 output.t5 gnd 0.044422f
C314 output.n6 gnd 0.364624f
C315 output.n7 gnd 0.350265f
C316 output.t7 gnd 0.044422f
C317 output.t16 gnd 0.044422f
C318 output.n8 gnd 0.364624f
C319 output.n9 gnd 0.350265f
C320 output.t17 gnd 0.044422f
C321 output.t8 gnd 0.044422f
C322 output.n10 gnd 0.364624f
C323 output.n11 gnd 0.350265f
C324 output.t9 gnd 0.044422f
C325 output.t14 gnd 0.044422f
C326 output.n12 gnd 0.364624f
C327 output.n13 gnd 0.350265f
C328 output.t6 gnd 0.462979f
C329 output.n14 gnd 0.28994f
C330 output.n15 gnd 0.015803f
C331 output.n16 gnd 0.011243f
C332 output.n17 gnd 0.006041f
C333 output.n18 gnd 0.01428f
C334 output.n19 gnd 0.006397f
C335 output.n20 gnd 0.011243f
C336 output.n21 gnd 0.006041f
C337 output.n22 gnd 0.01428f
C338 output.n23 gnd 0.006397f
C339 output.n24 gnd 0.048111f
C340 output.t19 gnd 0.023274f
C341 output.n25 gnd 0.01071f
C342 output.n26 gnd 0.008435f
C343 output.n27 gnd 0.006041f
C344 output.n28 gnd 0.267512f
C345 output.n29 gnd 0.011243f
C346 output.n30 gnd 0.006041f
C347 output.n31 gnd 0.006397f
C348 output.n32 gnd 0.01428f
C349 output.n33 gnd 0.01428f
C350 output.n34 gnd 0.006397f
C351 output.n35 gnd 0.006041f
C352 output.n36 gnd 0.011243f
C353 output.n37 gnd 0.011243f
C354 output.n38 gnd 0.006041f
C355 output.n39 gnd 0.006397f
C356 output.n40 gnd 0.01428f
C357 output.n41 gnd 0.030913f
C358 output.n42 gnd 0.006397f
C359 output.n43 gnd 0.006041f
C360 output.n44 gnd 0.025987f
C361 output.n45 gnd 0.097665f
C362 output.n46 gnd 0.015803f
C363 output.n47 gnd 0.011243f
C364 output.n48 gnd 0.006041f
C365 output.n49 gnd 0.01428f
C366 output.n50 gnd 0.006397f
C367 output.n51 gnd 0.011243f
C368 output.n52 gnd 0.006041f
C369 output.n53 gnd 0.01428f
C370 output.n54 gnd 0.006397f
C371 output.n55 gnd 0.048111f
C372 output.t1 gnd 0.023274f
C373 output.n56 gnd 0.01071f
C374 output.n57 gnd 0.008435f
C375 output.n58 gnd 0.006041f
C376 output.n59 gnd 0.267512f
C377 output.n60 gnd 0.011243f
C378 output.n61 gnd 0.006041f
C379 output.n62 gnd 0.006397f
C380 output.n63 gnd 0.01428f
C381 output.n64 gnd 0.01428f
C382 output.n65 gnd 0.006397f
C383 output.n66 gnd 0.006041f
C384 output.n67 gnd 0.011243f
C385 output.n68 gnd 0.011243f
C386 output.n69 gnd 0.006041f
C387 output.n70 gnd 0.006397f
C388 output.n71 gnd 0.01428f
C389 output.n72 gnd 0.030913f
C390 output.n73 gnd 0.006397f
C391 output.n74 gnd 0.006041f
C392 output.n75 gnd 0.025987f
C393 output.n76 gnd 0.09306f
C394 output.n77 gnd 1.65264f
C395 output.n78 gnd 0.015803f
C396 output.n79 gnd 0.011243f
C397 output.n80 gnd 0.006041f
C398 output.n81 gnd 0.01428f
C399 output.n82 gnd 0.006397f
C400 output.n83 gnd 0.011243f
C401 output.n84 gnd 0.006041f
C402 output.n85 gnd 0.01428f
C403 output.n86 gnd 0.006397f
C404 output.n87 gnd 0.048111f
C405 output.t2 gnd 0.023274f
C406 output.n88 gnd 0.01071f
C407 output.n89 gnd 0.008435f
C408 output.n90 gnd 0.006041f
C409 output.n91 gnd 0.267512f
C410 output.n92 gnd 0.011243f
C411 output.n93 gnd 0.006041f
C412 output.n94 gnd 0.006397f
C413 output.n95 gnd 0.01428f
C414 output.n96 gnd 0.01428f
C415 output.n97 gnd 0.006397f
C416 output.n98 gnd 0.006041f
C417 output.n99 gnd 0.011243f
C418 output.n100 gnd 0.011243f
C419 output.n101 gnd 0.006041f
C420 output.n102 gnd 0.006397f
C421 output.n103 gnd 0.01428f
C422 output.n104 gnd 0.030913f
C423 output.n105 gnd 0.006397f
C424 output.n106 gnd 0.006041f
C425 output.n107 gnd 0.025987f
C426 output.n108 gnd 0.09306f
C427 output.n109 gnd 0.713089f
C428 output.n110 gnd 0.015803f
C429 output.n111 gnd 0.011243f
C430 output.n112 gnd 0.006041f
C431 output.n113 gnd 0.01428f
C432 output.n114 gnd 0.006397f
C433 output.n115 gnd 0.011243f
C434 output.n116 gnd 0.006041f
C435 output.n117 gnd 0.01428f
C436 output.n118 gnd 0.006397f
C437 output.n119 gnd 0.048111f
C438 output.t0 gnd 0.023274f
C439 output.n120 gnd 0.01071f
C440 output.n121 gnd 0.008435f
C441 output.n122 gnd 0.006041f
C442 output.n123 gnd 0.267512f
C443 output.n124 gnd 0.011243f
C444 output.n125 gnd 0.006041f
C445 output.n126 gnd 0.006397f
C446 output.n127 gnd 0.01428f
C447 output.n128 gnd 0.01428f
C448 output.n129 gnd 0.006397f
C449 output.n130 gnd 0.006041f
C450 output.n131 gnd 0.011243f
C451 output.n132 gnd 0.011243f
C452 output.n133 gnd 0.006041f
C453 output.n134 gnd 0.006397f
C454 output.n135 gnd 0.01428f
C455 output.n136 gnd 0.030913f
C456 output.n137 gnd 0.006397f
C457 output.n138 gnd 0.006041f
C458 output.n139 gnd 0.025987f
C459 output.n140 gnd 0.09306f
C460 output.n141 gnd 1.67353f
C461 a_n2982_8322.t15 gnd 0.100195f
C462 a_n2982_8322.t37 gnd 20.7864f
C463 a_n2982_8322.t34 gnd 20.640598f
C464 a_n2982_8322.t36 gnd 20.640598f
C465 a_n2982_8322.t32 gnd 20.7864f
C466 a_n2982_8322.t35 gnd 20.640598f
C467 a_n2982_8322.t33 gnd 28.793001f
C468 a_n2982_8322.t14 gnd 0.938175f
C469 a_n2982_8322.t27 gnd 0.100195f
C470 a_n2982_8322.t23 gnd 0.100195f
C471 a_n2982_8322.n0 gnd 0.705774f
C472 a_n2982_8322.n1 gnd 0.788598f
C473 a_n2982_8322.t30 gnd 0.100195f
C474 a_n2982_8322.t20 gnd 0.100195f
C475 a_n2982_8322.n2 gnd 0.705774f
C476 a_n2982_8322.n3 gnd 0.400677f
C477 a_n2982_8322.t11 gnd 0.100195f
C478 a_n2982_8322.t10 gnd 0.100195f
C479 a_n2982_8322.n4 gnd 0.705774f
C480 a_n2982_8322.n5 gnd 0.400677f
C481 a_n2982_8322.t24 gnd 0.100195f
C482 a_n2982_8322.t17 gnd 0.100195f
C483 a_n2982_8322.n6 gnd 0.705774f
C484 a_n2982_8322.n7 gnd 0.400677f
C485 a_n2982_8322.t21 gnd 0.100195f
C486 a_n2982_8322.t19 gnd 0.100195f
C487 a_n2982_8322.n8 gnd 0.705774f
C488 a_n2982_8322.n9 gnd 0.400677f
C489 a_n2982_8322.t8 gnd 0.936307f
C490 a_n2982_8322.n10 gnd 1.87205f
C491 a_n2982_8322.t3 gnd 0.938175f
C492 a_n2982_8322.t7 gnd 0.100195f
C493 a_n2982_8322.t6 gnd 0.100195f
C494 a_n2982_8322.n11 gnd 0.705774f
C495 a_n2982_8322.n12 gnd 0.788598f
C496 a_n2982_8322.t1 gnd 0.936307f
C497 a_n2982_8322.n13 gnd 0.396834f
C498 a_n2982_8322.t4 gnd 0.936307f
C499 a_n2982_8322.n14 gnd 0.396834f
C500 a_n2982_8322.t2 gnd 0.100195f
C501 a_n2982_8322.t0 gnd 0.100195f
C502 a_n2982_8322.n15 gnd 0.705774f
C503 a_n2982_8322.n16 gnd 0.400677f
C504 a_n2982_8322.t5 gnd 0.936307f
C505 a_n2982_8322.n17 gnd 1.47193f
C506 a_n2982_8322.n18 gnd 2.35218f
C507 a_n2982_8322.n19 gnd 3.2687f
C508 a_n2982_8322.t9 gnd 0.936307f
C509 a_n2982_8322.n20 gnd 1.11185f
C510 a_n2982_8322.t26 gnd 0.100195f
C511 a_n2982_8322.t25 gnd 0.100195f
C512 a_n2982_8322.n21 gnd 0.705774f
C513 a_n2982_8322.n22 gnd 0.400677f
C514 a_n2982_8322.t13 gnd 0.100195f
C515 a_n2982_8322.t12 gnd 0.100195f
C516 a_n2982_8322.n23 gnd 0.705774f
C517 a_n2982_8322.n24 gnd 0.400677f
C518 a_n2982_8322.t28 gnd 0.100195f
C519 a_n2982_8322.t16 gnd 0.100195f
C520 a_n2982_8322.n25 gnd 0.705774f
C521 a_n2982_8322.n26 gnd 0.400677f
C522 a_n2982_8322.t29 gnd 0.938173f
C523 a_n2982_8322.t22 gnd 0.100195f
C524 a_n2982_8322.t18 gnd 0.100195f
C525 a_n2982_8322.n27 gnd 0.705774f
C526 a_n2982_8322.n28 gnd 0.7886f
C527 a_n2982_8322.n29 gnd 0.400675f
C528 a_n2982_8322.n30 gnd 0.705776f
C529 a_n2982_8322.t31 gnd 0.100195f
C530 a_n2804_13878.t29 gnd 0.194556f
C531 a_n2804_13878.t25 gnd 0.194556f
C532 a_n2804_13878.t31 gnd 0.194556f
C533 a_n2804_13878.n0 gnd 1.53449f
C534 a_n2804_13878.t8 gnd 0.194556f
C535 a_n2804_13878.t20 gnd 0.194556f
C536 a_n2804_13878.n1 gnd 1.53196f
C537 a_n2804_13878.n2 gnd 1.37704f
C538 a_n2804_13878.t12 gnd 0.194556f
C539 a_n2804_13878.t22 gnd 0.194556f
C540 a_n2804_13878.n3 gnd 1.53358f
C541 a_n2804_13878.t27 gnd 0.194556f
C542 a_n2804_13878.t17 gnd 0.194556f
C543 a_n2804_13878.n4 gnd 1.53196f
C544 a_n2804_13878.n5 gnd 2.14061f
C545 a_n2804_13878.t23 gnd 0.194556f
C546 a_n2804_13878.t16 gnd 0.194556f
C547 a_n2804_13878.n6 gnd 1.53196f
C548 a_n2804_13878.n7 gnd 1.04414f
C549 a_n2804_13878.t10 gnd 0.194556f
C550 a_n2804_13878.t13 gnd 0.194556f
C551 a_n2804_13878.n8 gnd 1.53196f
C552 a_n2804_13878.n9 gnd 1.04414f
C553 a_n2804_13878.t26 gnd 0.194556f
C554 a_n2804_13878.t11 gnd 0.194556f
C555 a_n2804_13878.n10 gnd 1.53196f
C556 a_n2804_13878.n11 gnd 1.04414f
C557 a_n2804_13878.t21 gnd 0.194556f
C558 a_n2804_13878.t9 gnd 0.194556f
C559 a_n2804_13878.n12 gnd 1.53196f
C560 a_n2804_13878.n13 gnd 4.90178f
C561 a_n2804_13878.t1 gnd 1.82172f
C562 a_n2804_13878.t4 gnd 0.194556f
C563 a_n2804_13878.t5 gnd 0.194556f
C564 a_n2804_13878.n14 gnd 1.37045f
C565 a_n2804_13878.n15 gnd 1.53128f
C566 a_n2804_13878.t0 gnd 1.81809f
C567 a_n2804_13878.n16 gnd 0.770559f
C568 a_n2804_13878.t3 gnd 1.81809f
C569 a_n2804_13878.n17 gnd 0.770559f
C570 a_n2804_13878.t6 gnd 0.194556f
C571 a_n2804_13878.t7 gnd 0.194556f
C572 a_n2804_13878.n18 gnd 1.37045f
C573 a_n2804_13878.n19 gnd 0.778022f
C574 a_n2804_13878.t2 gnd 1.81809f
C575 a_n2804_13878.n20 gnd 2.85814f
C576 a_n2804_13878.n21 gnd 3.74876f
C577 a_n2804_13878.t15 gnd 0.194556f
C578 a_n2804_13878.t24 gnd 0.194556f
C579 a_n2804_13878.n22 gnd 1.53195f
C580 a_n2804_13878.n23 gnd 2.50239f
C581 a_n2804_13878.t28 gnd 0.194556f
C582 a_n2804_13878.t14 gnd 0.194556f
C583 a_n2804_13878.n24 gnd 1.53196f
C584 a_n2804_13878.n25 gnd 0.678771f
C585 a_n2804_13878.t18 gnd 0.194556f
C586 a_n2804_13878.t19 gnd 0.194556f
C587 a_n2804_13878.n26 gnd 1.53196f
C588 a_n2804_13878.n27 gnd 0.678771f
C589 a_n2804_13878.n28 gnd 0.678768f
C590 a_n2804_13878.n29 gnd 1.53196f
C591 a_n2804_13878.t30 gnd 0.194556f
C592 vdd.t120 gnd 0.032405f
C593 vdd.t101 gnd 0.032405f
C594 vdd.n0 gnd 0.255579f
C595 vdd.t79 gnd 0.032405f
C596 vdd.t116 gnd 0.032405f
C597 vdd.n1 gnd 0.255158f
C598 vdd.n2 gnd 0.235304f
C599 vdd.t97 gnd 0.032405f
C600 vdd.t127 gnd 0.032405f
C601 vdd.n3 gnd 0.255158f
C602 vdd.n4 gnd 0.119002f
C603 vdd.t125 gnd 0.032405f
C604 vdd.t105 gnd 0.032405f
C605 vdd.n5 gnd 0.255158f
C606 vdd.n6 gnd 0.111661f
C607 vdd.t131 gnd 0.032405f
C608 vdd.t95 gnd 0.032405f
C609 vdd.n7 gnd 0.255579f
C610 vdd.t103 gnd 0.032405f
C611 vdd.t123 gnd 0.032405f
C612 vdd.n8 gnd 0.255158f
C613 vdd.n9 gnd 0.235304f
C614 vdd.t112 gnd 0.032405f
C615 vdd.t83 gnd 0.032405f
C616 vdd.n10 gnd 0.255158f
C617 vdd.n11 gnd 0.119002f
C618 vdd.t92 gnd 0.032405f
C619 vdd.t110 gnd 0.032405f
C620 vdd.n12 gnd 0.255158f
C621 vdd.n13 gnd 0.111661f
C622 vdd.n14 gnd 0.078943f
C623 vdd.t145 gnd 0.018003f
C624 vdd.t144 gnd 0.018003f
C625 vdd.n15 gnd 0.165705f
C626 vdd.t146 gnd 0.018003f
C627 vdd.t132 gnd 0.018003f
C628 vdd.n16 gnd 0.165221f
C629 vdd.n17 gnd 0.287535f
C630 vdd.t139 gnd 0.018003f
C631 vdd.t136 gnd 0.018003f
C632 vdd.n18 gnd 0.165221f
C633 vdd.n19 gnd 0.118957f
C634 vdd.t143 gnd 0.018003f
C635 vdd.t134 gnd 0.018003f
C636 vdd.n20 gnd 0.165705f
C637 vdd.t141 gnd 0.018003f
C638 vdd.t137 gnd 0.018003f
C639 vdd.n21 gnd 0.165221f
C640 vdd.n22 gnd 0.287535f
C641 vdd.t142 gnd 0.018003f
C642 vdd.t138 gnd 0.018003f
C643 vdd.n23 gnd 0.165221f
C644 vdd.n24 gnd 0.118957f
C645 vdd.t133 gnd 0.018003f
C646 vdd.t135 gnd 0.018003f
C647 vdd.n25 gnd 0.165221f
C648 vdd.t147 gnd 0.018003f
C649 vdd.t140 gnd 0.018003f
C650 vdd.n26 gnd 0.165221f
C651 vdd.n27 gnd 18.1145f
C652 vdd.n28 gnd 7.14758f
C653 vdd.n29 gnd 0.00491f
C654 vdd.n30 gnd 0.004556f
C655 vdd.n31 gnd 0.00252f
C656 vdd.n32 gnd 0.005787f
C657 vdd.n33 gnd 0.002448f
C658 vdd.n34 gnd 0.002592f
C659 vdd.n35 gnd 0.004556f
C660 vdd.n36 gnd 0.002448f
C661 vdd.n37 gnd 0.005787f
C662 vdd.n38 gnd 0.002592f
C663 vdd.n39 gnd 0.004556f
C664 vdd.n40 gnd 0.002448f
C665 vdd.n41 gnd 0.00434f
C666 vdd.n42 gnd 0.004353f
C667 vdd.t201 gnd 0.012433f
C668 vdd.n43 gnd 0.027663f
C669 vdd.n44 gnd 0.143964f
C670 vdd.n45 gnd 0.002448f
C671 vdd.n46 gnd 0.002592f
C672 vdd.n47 gnd 0.005787f
C673 vdd.n48 gnd 0.005787f
C674 vdd.n49 gnd 0.002592f
C675 vdd.n50 gnd 0.002448f
C676 vdd.n51 gnd 0.004556f
C677 vdd.n52 gnd 0.004556f
C678 vdd.n53 gnd 0.002448f
C679 vdd.n54 gnd 0.002592f
C680 vdd.n55 gnd 0.005787f
C681 vdd.n56 gnd 0.005787f
C682 vdd.n57 gnd 0.002592f
C683 vdd.n58 gnd 0.002448f
C684 vdd.n59 gnd 0.004556f
C685 vdd.n60 gnd 0.004556f
C686 vdd.n61 gnd 0.002448f
C687 vdd.n62 gnd 0.002592f
C688 vdd.n63 gnd 0.005787f
C689 vdd.n64 gnd 0.005787f
C690 vdd.n65 gnd 0.013682f
C691 vdd.n66 gnd 0.00252f
C692 vdd.n67 gnd 0.002448f
C693 vdd.n68 gnd 0.011777f
C694 vdd.n69 gnd 0.008222f
C695 vdd.t181 gnd 0.028804f
C696 vdd.t232 gnd 0.028804f
C697 vdd.n70 gnd 0.197961f
C698 vdd.n71 gnd 0.155666f
C699 vdd.t166 gnd 0.028804f
C700 vdd.t217 gnd 0.028804f
C701 vdd.n72 gnd 0.197961f
C702 vdd.n73 gnd 0.125622f
C703 vdd.t171 gnd 0.028804f
C704 vdd.t228 gnd 0.028804f
C705 vdd.n74 gnd 0.197961f
C706 vdd.n75 gnd 0.125622f
C707 vdd.t193 gnd 0.028804f
C708 vdd.t236 gnd 0.028804f
C709 vdd.n76 gnd 0.197961f
C710 vdd.n77 gnd 0.125622f
C711 vdd.t204 gnd 0.028804f
C712 vdd.t223 gnd 0.028804f
C713 vdd.n78 gnd 0.197961f
C714 vdd.n79 gnd 0.125622f
C715 vdd.n80 gnd 0.00491f
C716 vdd.n81 gnd 0.004556f
C717 vdd.n82 gnd 0.00252f
C718 vdd.n83 gnd 0.005787f
C719 vdd.n84 gnd 0.002448f
C720 vdd.n85 gnd 0.002592f
C721 vdd.n86 gnd 0.004556f
C722 vdd.n87 gnd 0.002448f
C723 vdd.n88 gnd 0.005787f
C724 vdd.n89 gnd 0.002592f
C725 vdd.n90 gnd 0.004556f
C726 vdd.n91 gnd 0.002448f
C727 vdd.n92 gnd 0.00434f
C728 vdd.n93 gnd 0.004353f
C729 vdd.t184 gnd 0.012433f
C730 vdd.n94 gnd 0.027663f
C731 vdd.n95 gnd 0.143964f
C732 vdd.n96 gnd 0.002448f
C733 vdd.n97 gnd 0.002592f
C734 vdd.n98 gnd 0.005787f
C735 vdd.n99 gnd 0.005787f
C736 vdd.n100 gnd 0.002592f
C737 vdd.n101 gnd 0.002448f
C738 vdd.n102 gnd 0.004556f
C739 vdd.n103 gnd 0.004556f
C740 vdd.n104 gnd 0.002448f
C741 vdd.n105 gnd 0.002592f
C742 vdd.n106 gnd 0.005787f
C743 vdd.n107 gnd 0.005787f
C744 vdd.n108 gnd 0.002592f
C745 vdd.n109 gnd 0.002448f
C746 vdd.n110 gnd 0.004556f
C747 vdd.n111 gnd 0.004556f
C748 vdd.n112 gnd 0.002448f
C749 vdd.n113 gnd 0.002592f
C750 vdd.n114 gnd 0.005787f
C751 vdd.n115 gnd 0.005787f
C752 vdd.n116 gnd 0.013682f
C753 vdd.n117 gnd 0.00252f
C754 vdd.n118 gnd 0.002448f
C755 vdd.n119 gnd 0.011777f
C756 vdd.n120 gnd 0.007964f
C757 vdd.n121 gnd 0.093463f
C758 vdd.n122 gnd 0.00491f
C759 vdd.n123 gnd 0.004556f
C760 vdd.n124 gnd 0.00252f
C761 vdd.n125 gnd 0.005787f
C762 vdd.n126 gnd 0.002448f
C763 vdd.n127 gnd 0.002592f
C764 vdd.n128 gnd 0.004556f
C765 vdd.n129 gnd 0.002448f
C766 vdd.n130 gnd 0.005787f
C767 vdd.n131 gnd 0.002592f
C768 vdd.n132 gnd 0.004556f
C769 vdd.n133 gnd 0.002448f
C770 vdd.n134 gnd 0.00434f
C771 vdd.n135 gnd 0.004353f
C772 vdd.t234 gnd 0.012433f
C773 vdd.n136 gnd 0.027663f
C774 vdd.n137 gnd 0.143964f
C775 vdd.n138 gnd 0.002448f
C776 vdd.n139 gnd 0.002592f
C777 vdd.n140 gnd 0.005787f
C778 vdd.n141 gnd 0.005787f
C779 vdd.n142 gnd 0.002592f
C780 vdd.n143 gnd 0.002448f
C781 vdd.n144 gnd 0.004556f
C782 vdd.n145 gnd 0.004556f
C783 vdd.n146 gnd 0.002448f
C784 vdd.n147 gnd 0.002592f
C785 vdd.n148 gnd 0.005787f
C786 vdd.n149 gnd 0.005787f
C787 vdd.n150 gnd 0.002592f
C788 vdd.n151 gnd 0.002448f
C789 vdd.n152 gnd 0.004556f
C790 vdd.n153 gnd 0.004556f
C791 vdd.n154 gnd 0.002448f
C792 vdd.n155 gnd 0.002592f
C793 vdd.n156 gnd 0.005787f
C794 vdd.n157 gnd 0.005787f
C795 vdd.n158 gnd 0.013682f
C796 vdd.n159 gnd 0.00252f
C797 vdd.n160 gnd 0.002448f
C798 vdd.n161 gnd 0.011777f
C799 vdd.n162 gnd 0.008222f
C800 vdd.t235 gnd 0.028804f
C801 vdd.t163 gnd 0.028804f
C802 vdd.n163 gnd 0.197961f
C803 vdd.n164 gnd 0.155666f
C804 vdd.t225 gnd 0.028804f
C805 vdd.t231 gnd 0.028804f
C806 vdd.n165 gnd 0.197961f
C807 vdd.n166 gnd 0.125622f
C808 vdd.t159 gnd 0.028804f
C809 vdd.t199 gnd 0.028804f
C810 vdd.n167 gnd 0.197961f
C811 vdd.n168 gnd 0.125622f
C812 vdd.t222 gnd 0.028804f
C813 vdd.t239 gnd 0.028804f
C814 vdd.n169 gnd 0.197961f
C815 vdd.n170 gnd 0.125622f
C816 vdd.t187 gnd 0.028804f
C817 vdd.t221 gnd 0.028804f
C818 vdd.n171 gnd 0.197961f
C819 vdd.n172 gnd 0.125622f
C820 vdd.n173 gnd 0.00491f
C821 vdd.n174 gnd 0.004556f
C822 vdd.n175 gnd 0.00252f
C823 vdd.n176 gnd 0.005787f
C824 vdd.n177 gnd 0.002448f
C825 vdd.n178 gnd 0.002592f
C826 vdd.n179 gnd 0.004556f
C827 vdd.n180 gnd 0.002448f
C828 vdd.n181 gnd 0.005787f
C829 vdd.n182 gnd 0.002592f
C830 vdd.n183 gnd 0.004556f
C831 vdd.n184 gnd 0.002448f
C832 vdd.n185 gnd 0.00434f
C833 vdd.n186 gnd 0.004353f
C834 vdd.t242 gnd 0.012433f
C835 vdd.n187 gnd 0.027663f
C836 vdd.n188 gnd 0.143964f
C837 vdd.n189 gnd 0.002448f
C838 vdd.n190 gnd 0.002592f
C839 vdd.n191 gnd 0.005787f
C840 vdd.n192 gnd 0.005787f
C841 vdd.n193 gnd 0.002592f
C842 vdd.n194 gnd 0.002448f
C843 vdd.n195 gnd 0.004556f
C844 vdd.n196 gnd 0.004556f
C845 vdd.n197 gnd 0.002448f
C846 vdd.n198 gnd 0.002592f
C847 vdd.n199 gnd 0.005787f
C848 vdd.n200 gnd 0.005787f
C849 vdd.n201 gnd 0.002592f
C850 vdd.n202 gnd 0.002448f
C851 vdd.n203 gnd 0.004556f
C852 vdd.n204 gnd 0.004556f
C853 vdd.n205 gnd 0.002448f
C854 vdd.n206 gnd 0.002592f
C855 vdd.n207 gnd 0.005787f
C856 vdd.n208 gnd 0.005787f
C857 vdd.n209 gnd 0.013682f
C858 vdd.n210 gnd 0.00252f
C859 vdd.n211 gnd 0.002448f
C860 vdd.n212 gnd 0.011777f
C861 vdd.n213 gnd 0.007964f
C862 vdd.n214 gnd 0.055601f
C863 vdd.n215 gnd 0.200345f
C864 vdd.n216 gnd 0.00491f
C865 vdd.n217 gnd 0.004556f
C866 vdd.n218 gnd 0.00252f
C867 vdd.n219 gnd 0.005787f
C868 vdd.n220 gnd 0.002448f
C869 vdd.n221 gnd 0.002592f
C870 vdd.n222 gnd 0.004556f
C871 vdd.n223 gnd 0.002448f
C872 vdd.n224 gnd 0.005787f
C873 vdd.n225 gnd 0.002592f
C874 vdd.n226 gnd 0.004556f
C875 vdd.n227 gnd 0.002448f
C876 vdd.n228 gnd 0.00434f
C877 vdd.n229 gnd 0.004353f
C878 vdd.t240 gnd 0.012433f
C879 vdd.n230 gnd 0.027663f
C880 vdd.n231 gnd 0.143964f
C881 vdd.n232 gnd 0.002448f
C882 vdd.n233 gnd 0.002592f
C883 vdd.n234 gnd 0.005787f
C884 vdd.n235 gnd 0.005787f
C885 vdd.n236 gnd 0.002592f
C886 vdd.n237 gnd 0.002448f
C887 vdd.n238 gnd 0.004556f
C888 vdd.n239 gnd 0.004556f
C889 vdd.n240 gnd 0.002448f
C890 vdd.n241 gnd 0.002592f
C891 vdd.n242 gnd 0.005787f
C892 vdd.n243 gnd 0.005787f
C893 vdd.n244 gnd 0.002592f
C894 vdd.n245 gnd 0.002448f
C895 vdd.n246 gnd 0.004556f
C896 vdd.n247 gnd 0.004556f
C897 vdd.n248 gnd 0.002448f
C898 vdd.n249 gnd 0.002592f
C899 vdd.n250 gnd 0.005787f
C900 vdd.n251 gnd 0.005787f
C901 vdd.n252 gnd 0.013682f
C902 vdd.n253 gnd 0.00252f
C903 vdd.n254 gnd 0.002448f
C904 vdd.n255 gnd 0.011777f
C905 vdd.n256 gnd 0.008222f
C906 vdd.t241 gnd 0.028804f
C907 vdd.t179 gnd 0.028804f
C908 vdd.n257 gnd 0.197961f
C909 vdd.n258 gnd 0.155666f
C910 vdd.t230 gnd 0.028804f
C911 vdd.t238 gnd 0.028804f
C912 vdd.n259 gnd 0.197961f
C913 vdd.n260 gnd 0.125622f
C914 vdd.t172 gnd 0.028804f
C915 vdd.t212 gnd 0.028804f
C916 vdd.n261 gnd 0.197961f
C917 vdd.n262 gnd 0.125622f
C918 vdd.t229 gnd 0.028804f
C919 vdd.t153 gnd 0.028804f
C920 vdd.n263 gnd 0.197961f
C921 vdd.n264 gnd 0.125622f
C922 vdd.t196 gnd 0.028804f
C923 vdd.t227 gnd 0.028804f
C924 vdd.n265 gnd 0.197961f
C925 vdd.n266 gnd 0.125622f
C926 vdd.n267 gnd 0.00491f
C927 vdd.n268 gnd 0.004556f
C928 vdd.n269 gnd 0.00252f
C929 vdd.n270 gnd 0.005787f
C930 vdd.n271 gnd 0.002448f
C931 vdd.n272 gnd 0.002592f
C932 vdd.n273 gnd 0.004556f
C933 vdd.n274 gnd 0.002448f
C934 vdd.n275 gnd 0.005787f
C935 vdd.n276 gnd 0.002592f
C936 vdd.n277 gnd 0.004556f
C937 vdd.n278 gnd 0.002448f
C938 vdd.n279 gnd 0.00434f
C939 vdd.n280 gnd 0.004353f
C940 vdd.t161 gnd 0.012433f
C941 vdd.n281 gnd 0.027663f
C942 vdd.n282 gnd 0.143964f
C943 vdd.n283 gnd 0.002448f
C944 vdd.n284 gnd 0.002592f
C945 vdd.n285 gnd 0.005787f
C946 vdd.n286 gnd 0.005787f
C947 vdd.n287 gnd 0.002592f
C948 vdd.n288 gnd 0.002448f
C949 vdd.n289 gnd 0.004556f
C950 vdd.n290 gnd 0.004556f
C951 vdd.n291 gnd 0.002448f
C952 vdd.n292 gnd 0.002592f
C953 vdd.n293 gnd 0.005787f
C954 vdd.n294 gnd 0.005787f
C955 vdd.n295 gnd 0.002592f
C956 vdd.n296 gnd 0.002448f
C957 vdd.n297 gnd 0.004556f
C958 vdd.n298 gnd 0.004556f
C959 vdd.n299 gnd 0.002448f
C960 vdd.n300 gnd 0.002592f
C961 vdd.n301 gnd 0.005787f
C962 vdd.n302 gnd 0.005787f
C963 vdd.n303 gnd 0.013682f
C964 vdd.n304 gnd 0.00252f
C965 vdd.n305 gnd 0.002448f
C966 vdd.n306 gnd 0.011777f
C967 vdd.n307 gnd 0.007964f
C968 vdd.n308 gnd 0.055601f
C969 vdd.n309 gnd 0.220186f
C970 vdd.n310 gnd 0.008916f
C971 vdd.n311 gnd 0.008916f
C972 vdd.n312 gnd 0.007201f
C973 vdd.n313 gnd 0.007201f
C974 vdd.n314 gnd 0.008947f
C975 vdd.n315 gnd 0.008947f
C976 vdd.t158 gnd 0.457154f
C977 vdd.n316 gnd 0.008947f
C978 vdd.n317 gnd 0.008947f
C979 vdd.n318 gnd 0.008947f
C980 vdd.t192 gnd 0.457154f
C981 vdd.n319 gnd 0.008947f
C982 vdd.n320 gnd 0.008947f
C983 vdd.n321 gnd 0.008947f
C984 vdd.n322 gnd 0.008947f
C985 vdd.n323 gnd 0.007201f
C986 vdd.n324 gnd 0.008947f
C987 vdd.n325 gnd 0.736018f
C988 vdd.n326 gnd 0.008947f
C989 vdd.n327 gnd 0.008947f
C990 vdd.n328 gnd 0.008947f
C991 vdd.n329 gnd 0.626301f
C992 vdd.n330 gnd 0.008947f
C993 vdd.n331 gnd 0.008947f
C994 vdd.n332 gnd 0.008947f
C995 vdd.n333 gnd 0.008947f
C996 vdd.n334 gnd 0.008947f
C997 vdd.n335 gnd 0.007201f
C998 vdd.n336 gnd 0.008947f
C999 vdd.t220 gnd 0.457154f
C1000 vdd.n337 gnd 0.008947f
C1001 vdd.n338 gnd 0.008947f
C1002 vdd.n339 gnd 0.008947f
C1003 vdd.n340 gnd 0.914309f
C1004 vdd.n341 gnd 0.008947f
C1005 vdd.n342 gnd 0.008947f
C1006 vdd.n343 gnd 0.008947f
C1007 vdd.n344 gnd 0.008947f
C1008 vdd.n345 gnd 0.008947f
C1009 vdd.n346 gnd 0.007201f
C1010 vdd.n347 gnd 0.008947f
C1011 vdd.n348 gnd 0.008947f
C1012 vdd.n349 gnd 0.008947f
C1013 vdd.n350 gnd 0.021084f
C1014 vdd.n351 gnd 2.10291f
C1015 vdd.n352 gnd 0.021413f
C1016 vdd.n353 gnd 0.008947f
C1017 vdd.n354 gnd 0.008947f
C1018 vdd.n356 gnd 0.008947f
C1019 vdd.n357 gnd 0.008947f
C1020 vdd.n358 gnd 0.007201f
C1021 vdd.n359 gnd 0.007201f
C1022 vdd.n360 gnd 0.008947f
C1023 vdd.n361 gnd 0.008947f
C1024 vdd.n362 gnd 0.008947f
C1025 vdd.n363 gnd 0.008947f
C1026 vdd.n364 gnd 0.008947f
C1027 vdd.n365 gnd 0.008947f
C1028 vdd.n366 gnd 0.007201f
C1029 vdd.n368 gnd 0.008947f
C1030 vdd.n369 gnd 0.008947f
C1031 vdd.n370 gnd 0.008947f
C1032 vdd.n371 gnd 0.008947f
C1033 vdd.n372 gnd 0.008947f
C1034 vdd.n373 gnd 0.007201f
C1035 vdd.n375 gnd 0.008947f
C1036 vdd.n376 gnd 0.008947f
C1037 vdd.n377 gnd 0.008947f
C1038 vdd.n378 gnd 0.008947f
C1039 vdd.n379 gnd 0.008947f
C1040 vdd.n380 gnd 0.007201f
C1041 vdd.n382 gnd 0.008947f
C1042 vdd.n383 gnd 0.008947f
C1043 vdd.n384 gnd 0.008947f
C1044 vdd.n385 gnd 0.008947f
C1045 vdd.n386 gnd 0.006013f
C1046 vdd.t42 gnd 0.110068f
C1047 vdd.t41 gnd 0.117632f
C1048 vdd.t40 gnd 0.143747f
C1049 vdd.n387 gnd 0.184263f
C1050 vdd.n388 gnd 0.155535f
C1051 vdd.n390 gnd 0.008947f
C1052 vdd.n391 gnd 0.008947f
C1053 vdd.n392 gnd 0.007201f
C1054 vdd.n393 gnd 0.008947f
C1055 vdd.n395 gnd 0.008947f
C1056 vdd.n396 gnd 0.008947f
C1057 vdd.n397 gnd 0.008947f
C1058 vdd.n398 gnd 0.008947f
C1059 vdd.n399 gnd 0.007201f
C1060 vdd.n401 gnd 0.008947f
C1061 vdd.n402 gnd 0.008947f
C1062 vdd.n403 gnd 0.008947f
C1063 vdd.n404 gnd 0.008947f
C1064 vdd.n405 gnd 0.008947f
C1065 vdd.n406 gnd 0.007201f
C1066 vdd.n408 gnd 0.008947f
C1067 vdd.n409 gnd 0.008947f
C1068 vdd.n410 gnd 0.008947f
C1069 vdd.n411 gnd 0.008947f
C1070 vdd.n412 gnd 0.008947f
C1071 vdd.n413 gnd 0.007201f
C1072 vdd.n415 gnd 0.008947f
C1073 vdd.n416 gnd 0.008947f
C1074 vdd.n417 gnd 0.008947f
C1075 vdd.n418 gnd 0.008947f
C1076 vdd.n419 gnd 0.008947f
C1077 vdd.n420 gnd 0.007201f
C1078 vdd.n422 gnd 0.008947f
C1079 vdd.n423 gnd 0.008947f
C1080 vdd.n424 gnd 0.008947f
C1081 vdd.n425 gnd 0.008947f
C1082 vdd.n426 gnd 0.007129f
C1083 vdd.t25 gnd 0.110068f
C1084 vdd.t24 gnd 0.117632f
C1085 vdd.t22 gnd 0.143747f
C1086 vdd.n427 gnd 0.184263f
C1087 vdd.n428 gnd 0.155535f
C1088 vdd.n430 gnd 0.008947f
C1089 vdd.n431 gnd 0.008947f
C1090 vdd.n432 gnd 0.007201f
C1091 vdd.n433 gnd 0.008947f
C1092 vdd.n435 gnd 0.008947f
C1093 vdd.n436 gnd 0.008947f
C1094 vdd.n437 gnd 0.008947f
C1095 vdd.n438 gnd 0.008947f
C1096 vdd.n439 gnd 0.007201f
C1097 vdd.n441 gnd 0.008947f
C1098 vdd.n442 gnd 0.008947f
C1099 vdd.n443 gnd 0.008947f
C1100 vdd.n444 gnd 0.008947f
C1101 vdd.n445 gnd 0.008947f
C1102 vdd.n446 gnd 0.007201f
C1103 vdd.n448 gnd 0.008947f
C1104 vdd.n449 gnd 0.008947f
C1105 vdd.n450 gnd 0.008947f
C1106 vdd.n451 gnd 0.008947f
C1107 vdd.n452 gnd 0.008947f
C1108 vdd.n453 gnd 0.007201f
C1109 vdd.n455 gnd 0.008947f
C1110 vdd.n456 gnd 0.008947f
C1111 vdd.n457 gnd 0.008947f
C1112 vdd.n458 gnd 0.008947f
C1113 vdd.n459 gnd 0.008947f
C1114 vdd.n460 gnd 0.007201f
C1115 vdd.n462 gnd 0.008947f
C1116 vdd.n463 gnd 0.008947f
C1117 vdd.n464 gnd 0.008947f
C1118 vdd.n465 gnd 0.008947f
C1119 vdd.n466 gnd 0.008947f
C1120 vdd.n467 gnd 0.008947f
C1121 vdd.n468 gnd 0.007201f
C1122 vdd.n469 gnd 0.008947f
C1123 vdd.n470 gnd 0.008947f
C1124 vdd.n471 gnd 0.007201f
C1125 vdd.n472 gnd 0.008947f
C1126 vdd.n473 gnd 0.008947f
C1127 vdd.n474 gnd 0.007201f
C1128 vdd.n475 gnd 0.008947f
C1129 vdd.n476 gnd 0.007201f
C1130 vdd.n477 gnd 0.008947f
C1131 vdd.n478 gnd 0.007201f
C1132 vdd.n479 gnd 0.008947f
C1133 vdd.n480 gnd 0.008947f
C1134 vdd.t216 gnd 0.457154f
C1135 vdd.n481 gnd 0.489155f
C1136 vdd.n482 gnd 0.008947f
C1137 vdd.n483 gnd 0.007201f
C1138 vdd.n484 gnd 0.008947f
C1139 vdd.n485 gnd 0.007201f
C1140 vdd.n486 gnd 0.008947f
C1141 vdd.t165 gnd 0.457154f
C1142 vdd.n487 gnd 0.008947f
C1143 vdd.n488 gnd 0.007201f
C1144 vdd.n489 gnd 0.008947f
C1145 vdd.n490 gnd 0.007201f
C1146 vdd.n491 gnd 0.008947f
C1147 vdd.n492 gnd 0.717732f
C1148 vdd.n493 gnd 0.758876f
C1149 vdd.t162 gnd 0.457154f
C1150 vdd.n494 gnd 0.008947f
C1151 vdd.n495 gnd 0.007201f
C1152 vdd.n496 gnd 0.008947f
C1153 vdd.n497 gnd 0.007201f
C1154 vdd.n498 gnd 0.008947f
C1155 vdd.n499 gnd 0.5623f
C1156 vdd.n500 gnd 0.008947f
C1157 vdd.n501 gnd 0.007201f
C1158 vdd.n502 gnd 0.008947f
C1159 vdd.n503 gnd 0.007201f
C1160 vdd.n504 gnd 0.008947f
C1161 vdd.n505 gnd 0.914309f
C1162 vdd.t200 gnd 0.457154f
C1163 vdd.n506 gnd 0.008947f
C1164 vdd.n507 gnd 0.007201f
C1165 vdd.n508 gnd 0.008947f
C1166 vdd.n509 gnd 0.007201f
C1167 vdd.n510 gnd 0.008947f
C1168 vdd.n511 gnd 0.489155f
C1169 vdd.n512 gnd 0.008947f
C1170 vdd.n513 gnd 0.007201f
C1171 vdd.n514 gnd 0.021413f
C1172 vdd.n515 gnd 0.021413f
C1173 vdd.n516 gnd 11.0997f
C1174 vdd.t19 gnd 0.457154f
C1175 vdd.n517 gnd 0.021413f
C1176 vdd.n518 gnd 0.007694f
C1177 vdd.n519 gnd 0.007201f
C1178 vdd.n524 gnd 0.005726f
C1179 vdd.n525 gnd 0.007201f
C1180 vdd.n526 gnd 0.008947f
C1181 vdd.n527 gnd 0.008947f
C1182 vdd.n528 gnd 0.008947f
C1183 vdd.n529 gnd 0.008947f
C1184 vdd.n530 gnd 0.008947f
C1185 vdd.n531 gnd 0.007201f
C1186 vdd.n532 gnd 0.008947f
C1187 vdd.n533 gnd 0.008947f
C1188 vdd.n534 gnd 0.008947f
C1189 vdd.n535 gnd 0.008947f
C1190 vdd.n536 gnd 0.008947f
C1191 vdd.n537 gnd 0.007201f
C1192 vdd.n538 gnd 0.008947f
C1193 vdd.n539 gnd 0.008947f
C1194 vdd.n540 gnd 0.008947f
C1195 vdd.n541 gnd 0.008947f
C1196 vdd.n542 gnd 0.008947f
C1197 vdd.t54 gnd 0.110068f
C1198 vdd.t55 gnd 0.117632f
C1199 vdd.t53 gnd 0.143747f
C1200 vdd.n543 gnd 0.184263f
C1201 vdd.n544 gnd 0.154815f
C1202 vdd.n545 gnd 0.01469f
C1203 vdd.n546 gnd 0.008947f
C1204 vdd.n547 gnd 0.008947f
C1205 vdd.n548 gnd 0.008947f
C1206 vdd.n549 gnd 0.008947f
C1207 vdd.n550 gnd 0.008947f
C1208 vdd.n551 gnd 0.007201f
C1209 vdd.n552 gnd 0.008947f
C1210 vdd.n553 gnd 0.008947f
C1211 vdd.n554 gnd 0.008947f
C1212 vdd.n555 gnd 0.008947f
C1213 vdd.n556 gnd 0.008947f
C1214 vdd.n557 gnd 0.007201f
C1215 vdd.n558 gnd 0.008947f
C1216 vdd.n559 gnd 0.008947f
C1217 vdd.n560 gnd 0.008947f
C1218 vdd.n561 gnd 0.008947f
C1219 vdd.n562 gnd 0.008947f
C1220 vdd.n563 gnd 0.007201f
C1221 vdd.n564 gnd 0.008947f
C1222 vdd.n565 gnd 0.008947f
C1223 vdd.n566 gnd 0.008947f
C1224 vdd.n567 gnd 0.008947f
C1225 vdd.n568 gnd 0.008947f
C1226 vdd.n569 gnd 0.007201f
C1227 vdd.n570 gnd 0.008947f
C1228 vdd.n571 gnd 0.008947f
C1229 vdd.n572 gnd 0.008947f
C1230 vdd.n573 gnd 0.008947f
C1231 vdd.n574 gnd 0.008947f
C1232 vdd.n575 gnd 0.007201f
C1233 vdd.n576 gnd 0.008947f
C1234 vdd.n577 gnd 0.008947f
C1235 vdd.n578 gnd 0.008947f
C1236 vdd.n579 gnd 0.007129f
C1237 vdd.t44 gnd 0.110068f
C1238 vdd.t45 gnd 0.117632f
C1239 vdd.t43 gnd 0.143747f
C1240 vdd.n580 gnd 0.184263f
C1241 vdd.n581 gnd 0.154815f
C1242 vdd.n582 gnd 0.008947f
C1243 vdd.n583 gnd 0.007201f
C1244 vdd.n585 gnd 0.008947f
C1245 vdd.n587 gnd 0.008947f
C1246 vdd.n588 gnd 0.008947f
C1247 vdd.n589 gnd 0.007201f
C1248 vdd.n590 gnd 0.008947f
C1249 vdd.n591 gnd 0.008947f
C1250 vdd.n592 gnd 0.008947f
C1251 vdd.n593 gnd 0.008947f
C1252 vdd.n594 gnd 0.008947f
C1253 vdd.n595 gnd 0.007201f
C1254 vdd.n596 gnd 0.008947f
C1255 vdd.n597 gnd 0.008947f
C1256 vdd.n598 gnd 0.008947f
C1257 vdd.n599 gnd 0.008947f
C1258 vdd.n600 gnd 0.008947f
C1259 vdd.n601 gnd 0.007201f
C1260 vdd.n602 gnd 0.008947f
C1261 vdd.n603 gnd 0.008947f
C1262 vdd.n604 gnd 0.008947f
C1263 vdd.n605 gnd 0.005726f
C1264 vdd.n610 gnd 0.006084f
C1265 vdd.n611 gnd 0.006084f
C1266 vdd.n612 gnd 0.006084f
C1267 vdd.n613 gnd 10.797999f
C1268 vdd.n614 gnd 0.006084f
C1269 vdd.n615 gnd 0.006084f
C1270 vdd.n616 gnd 0.006084f
C1271 vdd.n618 gnd 0.006084f
C1272 vdd.n619 gnd 0.006084f
C1273 vdd.n621 gnd 0.006084f
C1274 vdd.n622 gnd 0.004429f
C1275 vdd.n624 gnd 0.006084f
C1276 vdd.t3 gnd 0.245843f
C1277 vdd.t2 gnd 0.251651f
C1278 vdd.t0 gnd 0.160496f
C1279 vdd.n625 gnd 0.086739f
C1280 vdd.n626 gnd 0.049201f
C1281 vdd.n627 gnd 0.008695f
C1282 vdd.n628 gnd 0.013814f
C1283 vdd.n630 gnd 0.006084f
C1284 vdd.n631 gnd 0.62173f
C1285 vdd.n632 gnd 0.013026f
C1286 vdd.n633 gnd 0.013026f
C1287 vdd.n634 gnd 0.006084f
C1288 vdd.n635 gnd 0.013814f
C1289 vdd.n636 gnd 0.006084f
C1290 vdd.n637 gnd 0.006084f
C1291 vdd.n638 gnd 0.006084f
C1292 vdd.n639 gnd 0.006084f
C1293 vdd.n640 gnd 0.006084f
C1294 vdd.n642 gnd 0.006084f
C1295 vdd.n643 gnd 0.006084f
C1296 vdd.n645 gnd 0.006084f
C1297 vdd.n646 gnd 0.006084f
C1298 vdd.n648 gnd 0.006084f
C1299 vdd.n649 gnd 0.006084f
C1300 vdd.n651 gnd 0.006084f
C1301 vdd.n652 gnd 0.006084f
C1302 vdd.n654 gnd 0.006084f
C1303 vdd.n655 gnd 0.006084f
C1304 vdd.n657 gnd 0.006084f
C1305 vdd.n658 gnd 0.004429f
C1306 vdd.n660 gnd 0.006084f
C1307 vdd.t17 gnd 0.245843f
C1308 vdd.t16 gnd 0.251651f
C1309 vdd.t15 gnd 0.160496f
C1310 vdd.n661 gnd 0.086739f
C1311 vdd.n662 gnd 0.049201f
C1312 vdd.n663 gnd 0.008695f
C1313 vdd.n664 gnd 0.006084f
C1314 vdd.n665 gnd 0.006084f
C1315 vdd.t1 gnd 0.310865f
C1316 vdd.n666 gnd 0.006084f
C1317 vdd.n667 gnd 0.006084f
C1318 vdd.n668 gnd 0.006084f
C1319 vdd.n669 gnd 0.006084f
C1320 vdd.n670 gnd 0.006084f
C1321 vdd.n671 gnd 0.62173f
C1322 vdd.n672 gnd 0.006084f
C1323 vdd.n673 gnd 0.006084f
C1324 vdd.n674 gnd 0.489155f
C1325 vdd.n675 gnd 0.006084f
C1326 vdd.n676 gnd 0.006084f
C1327 vdd.n677 gnd 0.006084f
C1328 vdd.n678 gnd 0.006084f
C1329 vdd.n679 gnd 0.62173f
C1330 vdd.n680 gnd 0.006084f
C1331 vdd.n681 gnd 0.006084f
C1332 vdd.n682 gnd 0.006084f
C1333 vdd.n683 gnd 0.006084f
C1334 vdd.n684 gnd 0.006084f
C1335 vdd.t90 gnd 0.310865f
C1336 vdd.n685 gnd 0.006084f
C1337 vdd.n686 gnd 0.006084f
C1338 vdd.n687 gnd 0.006084f
C1339 vdd.n688 gnd 0.006084f
C1340 vdd.n689 gnd 0.006084f
C1341 vdd.t107 gnd 0.310865f
C1342 vdd.n690 gnd 0.006084f
C1343 vdd.n691 gnd 0.006084f
C1344 vdd.n692 gnd 0.598872f
C1345 vdd.n693 gnd 0.006084f
C1346 vdd.n694 gnd 0.006084f
C1347 vdd.n695 gnd 0.006084f
C1348 vdd.t106 gnd 0.310865f
C1349 vdd.n696 gnd 0.006084f
C1350 vdd.n697 gnd 0.006084f
C1351 vdd.n698 gnd 0.461726f
C1352 vdd.n699 gnd 0.006084f
C1353 vdd.n700 gnd 0.006084f
C1354 vdd.n701 gnd 0.006084f
C1355 vdd.n702 gnd 0.434297f
C1356 vdd.n703 gnd 0.006084f
C1357 vdd.n704 gnd 0.006084f
C1358 vdd.n705 gnd 0.32458f
C1359 vdd.n706 gnd 0.006084f
C1360 vdd.n707 gnd 0.006084f
C1361 vdd.n708 gnd 0.006084f
C1362 vdd.n709 gnd 0.571443f
C1363 vdd.n710 gnd 0.006084f
C1364 vdd.n711 gnd 0.006084f
C1365 vdd.t113 gnd 0.310865f
C1366 vdd.n712 gnd 0.006084f
C1367 vdd.n713 gnd 0.006084f
C1368 vdd.n714 gnd 0.006084f
C1369 vdd.n715 gnd 0.62173f
C1370 vdd.n716 gnd 0.006084f
C1371 vdd.n717 gnd 0.006084f
C1372 vdd.t114 gnd 0.310865f
C1373 vdd.n718 gnd 0.006084f
C1374 vdd.n719 gnd 0.006084f
C1375 vdd.n720 gnd 0.006084f
C1376 vdd.t84 gnd 0.310865f
C1377 vdd.n721 gnd 0.006084f
C1378 vdd.n722 gnd 0.006084f
C1379 vdd.n723 gnd 0.006084f
C1380 vdd.t28 gnd 0.251651f
C1381 vdd.t26 gnd 0.160496f
C1382 vdd.t29 gnd 0.251651f
C1383 vdd.n724 gnd 0.141438f
C1384 vdd.n725 gnd 0.017624f
C1385 vdd.n726 gnd 0.006084f
C1386 vdd.t27 gnd 0.224006f
C1387 vdd.n727 gnd 0.006084f
C1388 vdd.n728 gnd 0.006084f
C1389 vdd.n729 gnd 0.534871f
C1390 vdd.n730 gnd 0.006084f
C1391 vdd.n731 gnd 0.006084f
C1392 vdd.n732 gnd 0.006084f
C1393 vdd.n733 gnd 0.361152f
C1394 vdd.n734 gnd 0.006084f
C1395 vdd.n735 gnd 0.006084f
C1396 vdd.t85 gnd 0.128003f
C1397 vdd.n736 gnd 0.397724f
C1398 vdd.n737 gnd 0.006084f
C1399 vdd.n738 gnd 0.006084f
C1400 vdd.n739 gnd 0.006084f
C1401 vdd.n740 gnd 0.498298f
C1402 vdd.n741 gnd 0.006084f
C1403 vdd.n742 gnd 0.006084f
C1404 vdd.t98 gnd 0.310865f
C1405 vdd.n743 gnd 0.006084f
C1406 vdd.n744 gnd 0.006084f
C1407 vdd.n745 gnd 0.006084f
C1408 vdd.t94 gnd 0.310865f
C1409 vdd.n746 gnd 0.006084f
C1410 vdd.n747 gnd 0.006084f
C1411 vdd.t117 gnd 0.310865f
C1412 vdd.n748 gnd 0.006084f
C1413 vdd.n749 gnd 0.006084f
C1414 vdd.n750 gnd 0.006084f
C1415 vdd.t76 gnd 0.210291f
C1416 vdd.n751 gnd 0.006084f
C1417 vdd.n752 gnd 0.006084f
C1418 vdd.n753 gnd 0.548585f
C1419 vdd.n754 gnd 0.006084f
C1420 vdd.n755 gnd 0.006084f
C1421 vdd.n756 gnd 0.006084f
C1422 vdd.t118 gnd 0.310865f
C1423 vdd.n757 gnd 0.006084f
C1424 vdd.n758 gnd 0.006084f
C1425 vdd.t130 gnd 0.29715f
C1426 vdd.n759 gnd 0.411439f
C1427 vdd.n760 gnd 0.006084f
C1428 vdd.n761 gnd 0.006084f
C1429 vdd.n762 gnd 0.006084f
C1430 vdd.t80 gnd 0.310865f
C1431 vdd.n763 gnd 0.006084f
C1432 vdd.n764 gnd 0.006084f
C1433 vdd.t122 gnd 0.310865f
C1434 vdd.n765 gnd 0.006084f
C1435 vdd.n766 gnd 0.006084f
C1436 vdd.n767 gnd 0.006084f
C1437 vdd.n768 gnd 0.62173f
C1438 vdd.n769 gnd 0.006084f
C1439 vdd.n770 gnd 0.006084f
C1440 vdd.t102 gnd 0.310865f
C1441 vdd.n771 gnd 0.006084f
C1442 vdd.n772 gnd 0.006084f
C1443 vdd.n773 gnd 0.006084f
C1444 vdd.n774 gnd 0.429725f
C1445 vdd.n775 gnd 0.006084f
C1446 vdd.n776 gnd 0.006084f
C1447 vdd.n777 gnd 0.006084f
C1448 vdd.n778 gnd 0.006084f
C1449 vdd.n779 gnd 0.006084f
C1450 vdd.t57 gnd 0.310865f
C1451 vdd.n780 gnd 0.006084f
C1452 vdd.n781 gnd 0.006084f
C1453 vdd.t82 gnd 0.310865f
C1454 vdd.n782 gnd 0.006084f
C1455 vdd.n783 gnd 0.013026f
C1456 vdd.n784 gnd 0.013026f
C1457 vdd.n785 gnd 0.704018f
C1458 vdd.n786 gnd 0.006084f
C1459 vdd.n787 gnd 0.006084f
C1460 vdd.t111 gnd 0.310865f
C1461 vdd.n788 gnd 0.013026f
C1462 vdd.n789 gnd 0.006084f
C1463 vdd.n790 gnd 0.006084f
C1464 vdd.t124 gnd 0.530299f
C1465 vdd.n808 gnd 0.013814f
C1466 vdd.n826 gnd 0.013026f
C1467 vdd.n827 gnd 0.006084f
C1468 vdd.n828 gnd 0.013026f
C1469 vdd.t75 gnd 0.245843f
C1470 vdd.t74 gnd 0.251651f
C1471 vdd.t73 gnd 0.160496f
C1472 vdd.n829 gnd 0.086739f
C1473 vdd.n830 gnd 0.049201f
C1474 vdd.n831 gnd 0.013814f
C1475 vdd.n832 gnd 0.006084f
C1476 vdd.n833 gnd 0.365723f
C1477 vdd.n834 gnd 0.013026f
C1478 vdd.n835 gnd 0.006084f
C1479 vdd.n836 gnd 0.013814f
C1480 vdd.n837 gnd 0.006084f
C1481 vdd.t52 gnd 0.245843f
C1482 vdd.t51 gnd 0.251651f
C1483 vdd.t49 gnd 0.160496f
C1484 vdd.n838 gnd 0.086739f
C1485 vdd.n839 gnd 0.049201f
C1486 vdd.n840 gnd 0.008695f
C1487 vdd.n841 gnd 0.006084f
C1488 vdd.n842 gnd 0.006084f
C1489 vdd.t50 gnd 0.310865f
C1490 vdd.n843 gnd 0.006084f
C1491 vdd.t126 gnd 0.310865f
C1492 vdd.n844 gnd 0.006084f
C1493 vdd.n845 gnd 0.006084f
C1494 vdd.n846 gnd 0.006084f
C1495 vdd.n847 gnd 0.006084f
C1496 vdd.n848 gnd 0.006084f
C1497 vdd.n849 gnd 0.62173f
C1498 vdd.n850 gnd 0.006084f
C1499 vdd.n851 gnd 0.006084f
C1500 vdd.t96 gnd 0.310865f
C1501 vdd.n852 gnd 0.006084f
C1502 vdd.n853 gnd 0.006084f
C1503 vdd.n854 gnd 0.006084f
C1504 vdd.n855 gnd 0.006084f
C1505 vdd.n856 gnd 0.448011f
C1506 vdd.n857 gnd 0.006084f
C1507 vdd.n858 gnd 0.006084f
C1508 vdd.n859 gnd 0.006084f
C1509 vdd.n860 gnd 0.006084f
C1510 vdd.n861 gnd 0.006084f
C1511 vdd.t77 gnd 0.310865f
C1512 vdd.n862 gnd 0.006084f
C1513 vdd.n863 gnd 0.006084f
C1514 vdd.t115 gnd 0.310865f
C1515 vdd.n864 gnd 0.006084f
C1516 vdd.n865 gnd 0.006084f
C1517 vdd.n866 gnd 0.006084f
C1518 vdd.t99 gnd 0.310865f
C1519 vdd.n867 gnd 0.006084f
C1520 vdd.n868 gnd 0.006084f
C1521 vdd.t78 gnd 0.310865f
C1522 vdd.n869 gnd 0.006084f
C1523 vdd.n870 gnd 0.006084f
C1524 vdd.n871 gnd 0.006084f
C1525 vdd.t100 gnd 0.29715f
C1526 vdd.n872 gnd 0.006084f
C1527 vdd.n873 gnd 0.006084f
C1528 vdd.n874 gnd 0.461726f
C1529 vdd.n875 gnd 0.006084f
C1530 vdd.n876 gnd 0.006084f
C1531 vdd.n877 gnd 0.006084f
C1532 vdd.t119 gnd 0.310865f
C1533 vdd.n878 gnd 0.006084f
C1534 vdd.n879 gnd 0.006084f
C1535 vdd.t87 gnd 0.210291f
C1536 vdd.n880 gnd 0.32458f
C1537 vdd.n881 gnd 0.006084f
C1538 vdd.n882 gnd 0.006084f
C1539 vdd.n883 gnd 0.006084f
C1540 vdd.n884 gnd 0.571443f
C1541 vdd.n885 gnd 0.006084f
C1542 vdd.n886 gnd 0.006084f
C1543 vdd.t128 gnd 0.310865f
C1544 vdd.n887 gnd 0.006084f
C1545 vdd.n888 gnd 0.006084f
C1546 vdd.n889 gnd 0.006084f
C1547 vdd.n890 gnd 0.62173f
C1548 vdd.n891 gnd 0.006084f
C1549 vdd.n892 gnd 0.006084f
C1550 vdd.t93 gnd 0.310865f
C1551 vdd.n893 gnd 0.006084f
C1552 vdd.n894 gnd 0.006084f
C1553 vdd.n895 gnd 0.006084f
C1554 vdd.t86 gnd 0.128003f
C1555 vdd.n896 gnd 0.006084f
C1556 vdd.n897 gnd 0.006084f
C1557 vdd.n898 gnd 0.006084f
C1558 vdd.t65 gnd 0.251651f
C1559 vdd.t63 gnd 0.160496f
C1560 vdd.t66 gnd 0.251651f
C1561 vdd.n899 gnd 0.141438f
C1562 vdd.n900 gnd 0.006084f
C1563 vdd.n901 gnd 0.006084f
C1564 vdd.t108 gnd 0.310865f
C1565 vdd.n902 gnd 0.006084f
C1566 vdd.n903 gnd 0.006084f
C1567 vdd.t64 gnd 0.224006f
C1568 vdd.n904 gnd 0.493727f
C1569 vdd.n905 gnd 0.006084f
C1570 vdd.n906 gnd 0.006084f
C1571 vdd.n907 gnd 0.006084f
C1572 vdd.n908 gnd 0.361152f
C1573 vdd.n909 gnd 0.006084f
C1574 vdd.n910 gnd 0.006084f
C1575 vdd.n911 gnd 0.397724f
C1576 vdd.n912 gnd 0.006084f
C1577 vdd.n913 gnd 0.006084f
C1578 vdd.n914 gnd 0.006084f
C1579 vdd.n915 gnd 0.498298f
C1580 vdd.n916 gnd 0.006084f
C1581 vdd.n917 gnd 0.006084f
C1582 vdd.t88 gnd 0.310865f
C1583 vdd.n918 gnd 0.006084f
C1584 vdd.n919 gnd 0.006084f
C1585 vdd.n920 gnd 0.006084f
C1586 vdd.n921 gnd 0.62173f
C1587 vdd.n922 gnd 0.006084f
C1588 vdd.n923 gnd 0.006084f
C1589 vdd.t89 gnd 0.310865f
C1590 vdd.n924 gnd 0.006084f
C1591 vdd.n925 gnd 0.006084f
C1592 vdd.n926 gnd 0.006084f
C1593 vdd.t129 gnd 0.310865f
C1594 vdd.n927 gnd 0.006084f
C1595 vdd.n928 gnd 0.006084f
C1596 vdd.n929 gnd 0.006084f
C1597 vdd.n930 gnd 0.006084f
C1598 vdd.n931 gnd 0.006084f
C1599 vdd.t121 gnd 0.310865f
C1600 vdd.n932 gnd 0.006084f
C1601 vdd.n933 gnd 0.006084f
C1602 vdd.n934 gnd 0.608015f
C1603 vdd.n935 gnd 0.006084f
C1604 vdd.n936 gnd 0.006084f
C1605 vdd.n937 gnd 0.006084f
C1606 vdd.t81 gnd 0.310865f
C1607 vdd.n938 gnd 0.006084f
C1608 vdd.n939 gnd 0.006084f
C1609 vdd.n940 gnd 0.470869f
C1610 vdd.n941 gnd 0.006084f
C1611 vdd.n942 gnd 0.006084f
C1612 vdd.n943 gnd 0.006084f
C1613 vdd.n944 gnd 0.62173f
C1614 vdd.n945 gnd 0.006084f
C1615 vdd.n946 gnd 0.006084f
C1616 vdd.n947 gnd 0.333723f
C1617 vdd.n948 gnd 0.006084f
C1618 vdd.n949 gnd 0.006084f
C1619 vdd.n950 gnd 0.006084f
C1620 vdd.n951 gnd 0.62173f
C1621 vdd.n952 gnd 0.006084f
C1622 vdd.n953 gnd 0.006084f
C1623 vdd.n954 gnd 0.006084f
C1624 vdd.n955 gnd 0.006084f
C1625 vdd.n956 gnd 0.006084f
C1626 vdd.t5 gnd 0.310865f
C1627 vdd.n957 gnd 0.006084f
C1628 vdd.n958 gnd 0.006084f
C1629 vdd.n959 gnd 0.006084f
C1630 vdd.n960 gnd 0.013026f
C1631 vdd.n961 gnd 0.013026f
C1632 vdd.n962 gnd 0.841164f
C1633 vdd.n963 gnd 0.006084f
C1634 vdd.n964 gnd 0.006084f
C1635 vdd.n965 gnd 0.44344f
C1636 vdd.n966 gnd 0.013026f
C1637 vdd.n967 gnd 0.006084f
C1638 vdd.n968 gnd 0.006084f
C1639 vdd.n969 gnd 11.0997f
C1640 vdd.n1003 gnd 0.013814f
C1641 vdd.n1004 gnd 0.006084f
C1642 vdd.n1005 gnd 0.006084f
C1643 vdd.n1006 gnd 0.005726f
C1644 vdd.n1009 gnd 0.021413f
C1645 vdd.n1010 gnd 0.005977f
C1646 vdd.n1011 gnd 0.007201f
C1647 vdd.n1013 gnd 0.008947f
C1648 vdd.n1014 gnd 0.008947f
C1649 vdd.n1015 gnd 0.007201f
C1650 vdd.n1017 gnd 0.008947f
C1651 vdd.n1018 gnd 0.008947f
C1652 vdd.n1019 gnd 0.008947f
C1653 vdd.n1020 gnd 0.008947f
C1654 vdd.n1021 gnd 0.008947f
C1655 vdd.n1022 gnd 0.007201f
C1656 vdd.n1024 gnd 0.008947f
C1657 vdd.n1025 gnd 0.008947f
C1658 vdd.n1026 gnd 0.008947f
C1659 vdd.n1027 gnd 0.008947f
C1660 vdd.n1028 gnd 0.008947f
C1661 vdd.n1029 gnd 0.007201f
C1662 vdd.n1031 gnd 0.008947f
C1663 vdd.n1032 gnd 0.008947f
C1664 vdd.n1033 gnd 0.008947f
C1665 vdd.n1034 gnd 0.008947f
C1666 vdd.n1035 gnd 0.006013f
C1667 vdd.t14 gnd 0.110068f
C1668 vdd.t13 gnd 0.117632f
C1669 vdd.t12 gnd 0.143747f
C1670 vdd.n1036 gnd 0.184263f
C1671 vdd.n1037 gnd 0.154815f
C1672 vdd.n1039 gnd 0.008947f
C1673 vdd.n1040 gnd 0.008947f
C1674 vdd.n1041 gnd 0.007201f
C1675 vdd.n1042 gnd 0.008947f
C1676 vdd.n1044 gnd 0.008947f
C1677 vdd.n1045 gnd 0.008947f
C1678 vdd.n1046 gnd 0.008947f
C1679 vdd.n1047 gnd 0.008947f
C1680 vdd.n1048 gnd 0.007201f
C1681 vdd.n1050 gnd 0.008947f
C1682 vdd.n1051 gnd 0.008947f
C1683 vdd.n1052 gnd 0.008947f
C1684 vdd.n1053 gnd 0.008947f
C1685 vdd.n1054 gnd 0.008947f
C1686 vdd.n1055 gnd 0.007201f
C1687 vdd.n1057 gnd 0.008947f
C1688 vdd.n1058 gnd 0.008947f
C1689 vdd.n1059 gnd 0.008947f
C1690 vdd.n1060 gnd 0.008947f
C1691 vdd.n1061 gnd 0.008947f
C1692 vdd.n1062 gnd 0.007201f
C1693 vdd.n1064 gnd 0.008947f
C1694 vdd.n1065 gnd 0.008947f
C1695 vdd.n1066 gnd 0.008947f
C1696 vdd.n1067 gnd 0.008947f
C1697 vdd.n1068 gnd 0.008947f
C1698 vdd.n1069 gnd 0.007201f
C1699 vdd.n1071 gnd 0.008947f
C1700 vdd.n1072 gnd 0.008947f
C1701 vdd.n1073 gnd 0.008947f
C1702 vdd.n1074 gnd 0.008947f
C1703 vdd.n1075 gnd 0.007129f
C1704 vdd.t11 gnd 0.110068f
C1705 vdd.t10 gnd 0.117632f
C1706 vdd.t8 gnd 0.143747f
C1707 vdd.n1076 gnd 0.184263f
C1708 vdd.n1077 gnd 0.154815f
C1709 vdd.n1079 gnd 0.008947f
C1710 vdd.n1080 gnd 0.008947f
C1711 vdd.n1081 gnd 0.007201f
C1712 vdd.n1082 gnd 0.008947f
C1713 vdd.n1084 gnd 0.008947f
C1714 vdd.n1085 gnd 0.008947f
C1715 vdd.n1086 gnd 0.008947f
C1716 vdd.n1087 gnd 0.008947f
C1717 vdd.n1088 gnd 0.007201f
C1718 vdd.n1090 gnd 0.008947f
C1719 vdd.n1091 gnd 0.008947f
C1720 vdd.n1092 gnd 0.008947f
C1721 vdd.n1093 gnd 0.008947f
C1722 vdd.n1094 gnd 0.008947f
C1723 vdd.n1095 gnd 0.007201f
C1724 vdd.n1097 gnd 0.008947f
C1725 vdd.n1098 gnd 0.008947f
C1726 vdd.n1099 gnd 0.008947f
C1727 vdd.n1100 gnd 0.008947f
C1728 vdd.n1101 gnd 0.008947f
C1729 vdd.n1102 gnd 0.007201f
C1730 vdd.n1104 gnd 0.008947f
C1731 vdd.n1105 gnd 0.008947f
C1732 vdd.n1106 gnd 0.005726f
C1733 vdd.n1107 gnd 0.007201f
C1734 vdd.n1108 gnd 0.013814f
C1735 vdd.n1109 gnd 0.013814f
C1736 vdd.n1110 gnd 0.006084f
C1737 vdd.n1111 gnd 0.006084f
C1738 vdd.n1112 gnd 0.006084f
C1739 vdd.n1113 gnd 0.006084f
C1740 vdd.n1114 gnd 0.006084f
C1741 vdd.n1115 gnd 0.006084f
C1742 vdd.n1116 gnd 0.006084f
C1743 vdd.n1117 gnd 0.006084f
C1744 vdd.n1118 gnd 0.006084f
C1745 vdd.n1119 gnd 0.006084f
C1746 vdd.n1120 gnd 0.006084f
C1747 vdd.n1121 gnd 0.006084f
C1748 vdd.n1122 gnd 0.006084f
C1749 vdd.n1123 gnd 0.006084f
C1750 vdd.n1124 gnd 0.006084f
C1751 vdd.n1125 gnd 0.006084f
C1752 vdd.n1126 gnd 0.006084f
C1753 vdd.n1127 gnd 0.006084f
C1754 vdd.n1128 gnd 0.006084f
C1755 vdd.n1129 gnd 0.006084f
C1756 vdd.n1130 gnd 0.006084f
C1757 vdd.n1131 gnd 0.006084f
C1758 vdd.n1132 gnd 0.006084f
C1759 vdd.n1133 gnd 0.006084f
C1760 vdd.n1134 gnd 0.006084f
C1761 vdd.n1135 gnd 0.006084f
C1762 vdd.n1136 gnd 0.006084f
C1763 vdd.n1137 gnd 0.006084f
C1764 vdd.n1138 gnd 0.006084f
C1765 vdd.n1139 gnd 0.006084f
C1766 vdd.n1140 gnd 0.006084f
C1767 vdd.n1141 gnd 0.006084f
C1768 vdd.n1142 gnd 0.006084f
C1769 vdd.t6 gnd 0.245843f
C1770 vdd.t7 gnd 0.251651f
C1771 vdd.t4 gnd 0.160496f
C1772 vdd.n1143 gnd 0.086739f
C1773 vdd.n1144 gnd 0.049201f
C1774 vdd.n1145 gnd 0.008695f
C1775 vdd.n1146 gnd 0.006084f
C1776 vdd.t47 gnd 0.245843f
C1777 vdd.t48 gnd 0.251651f
C1778 vdd.t46 gnd 0.160496f
C1779 vdd.n1147 gnd 0.086739f
C1780 vdd.n1148 gnd 0.049201f
C1781 vdd.n1149 gnd 0.006084f
C1782 vdd.n1150 gnd 0.006084f
C1783 vdd.n1151 gnd 0.006084f
C1784 vdd.n1152 gnd 0.006084f
C1785 vdd.n1153 gnd 0.006084f
C1786 vdd.n1154 gnd 0.006084f
C1787 vdd.n1155 gnd 0.006084f
C1788 vdd.n1156 gnd 0.006084f
C1789 vdd.n1157 gnd 0.006084f
C1790 vdd.n1158 gnd 0.006084f
C1791 vdd.n1159 gnd 0.006084f
C1792 vdd.n1160 gnd 0.006084f
C1793 vdd.n1161 gnd 0.006084f
C1794 vdd.n1162 gnd 0.006084f
C1795 vdd.n1163 gnd 0.006084f
C1796 vdd.n1164 gnd 0.006084f
C1797 vdd.n1165 gnd 0.006084f
C1798 vdd.n1166 gnd 0.006084f
C1799 vdd.n1167 gnd 0.006084f
C1800 vdd.n1168 gnd 0.006084f
C1801 vdd.n1169 gnd 0.006084f
C1802 vdd.n1170 gnd 0.006084f
C1803 vdd.n1171 gnd 0.006084f
C1804 vdd.n1172 gnd 0.006084f
C1805 vdd.n1173 gnd 0.006084f
C1806 vdd.n1174 gnd 0.006084f
C1807 vdd.n1175 gnd 0.004429f
C1808 vdd.n1176 gnd 0.008695f
C1809 vdd.n1177 gnd 0.004697f
C1810 vdd.n1178 gnd 0.006084f
C1811 vdd.n1179 gnd 0.006084f
C1812 vdd.n1180 gnd 0.006084f
C1813 vdd.n1181 gnd 0.013814f
C1814 vdd.n1182 gnd 0.013814f
C1815 vdd.n1183 gnd 0.013026f
C1816 vdd.n1184 gnd 0.013026f
C1817 vdd.n1185 gnd 0.006084f
C1818 vdd.n1186 gnd 0.006084f
C1819 vdd.n1187 gnd 0.006084f
C1820 vdd.n1188 gnd 0.006084f
C1821 vdd.n1189 gnd 0.006084f
C1822 vdd.n1190 gnd 0.006084f
C1823 vdd.n1191 gnd 0.006084f
C1824 vdd.n1192 gnd 0.006084f
C1825 vdd.n1193 gnd 0.006084f
C1826 vdd.n1194 gnd 0.006084f
C1827 vdd.n1195 gnd 0.006084f
C1828 vdd.n1196 gnd 0.006084f
C1829 vdd.n1197 gnd 0.006084f
C1830 vdd.n1198 gnd 0.006084f
C1831 vdd.n1199 gnd 0.006084f
C1832 vdd.n1200 gnd 0.006084f
C1833 vdd.n1201 gnd 0.006084f
C1834 vdd.n1202 gnd 0.006084f
C1835 vdd.n1203 gnd 0.006084f
C1836 vdd.n1204 gnd 0.006084f
C1837 vdd.n1205 gnd 0.006084f
C1838 vdd.n1206 gnd 0.006084f
C1839 vdd.n1207 gnd 0.006084f
C1840 vdd.n1208 gnd 0.006084f
C1841 vdd.n1209 gnd 0.006084f
C1842 vdd.n1210 gnd 0.006084f
C1843 vdd.n1211 gnd 0.006084f
C1844 vdd.n1212 gnd 0.006084f
C1845 vdd.n1213 gnd 0.006084f
C1846 vdd.n1214 gnd 0.006084f
C1847 vdd.n1215 gnd 0.006084f
C1848 vdd.n1216 gnd 0.006084f
C1849 vdd.n1217 gnd 0.006084f
C1850 vdd.n1218 gnd 0.006084f
C1851 vdd.n1219 gnd 0.006084f
C1852 vdd.n1220 gnd 0.006084f
C1853 vdd.n1221 gnd 0.006084f
C1854 vdd.n1222 gnd 0.006084f
C1855 vdd.n1223 gnd 0.006084f
C1856 vdd.n1224 gnd 0.006084f
C1857 vdd.n1225 gnd 0.006084f
C1858 vdd.n1226 gnd 0.006084f
C1859 vdd.n1227 gnd 0.370295f
C1860 vdd.n1228 gnd 0.006084f
C1861 vdd.n1229 gnd 0.006084f
C1862 vdd.n1230 gnd 0.006084f
C1863 vdd.n1231 gnd 0.006084f
C1864 vdd.n1232 gnd 0.006084f
C1865 vdd.n1233 gnd 0.006084f
C1866 vdd.n1234 gnd 0.006084f
C1867 vdd.n1235 gnd 0.006084f
C1868 vdd.n1236 gnd 0.006084f
C1869 vdd.n1237 gnd 0.006084f
C1870 vdd.n1238 gnd 0.006084f
C1871 vdd.n1239 gnd 0.006084f
C1872 vdd.n1240 gnd 0.006084f
C1873 vdd.n1241 gnd 0.006084f
C1874 vdd.n1242 gnd 0.006084f
C1875 vdd.n1243 gnd 0.006084f
C1876 vdd.n1244 gnd 0.006084f
C1877 vdd.n1245 gnd 0.006084f
C1878 vdd.n1246 gnd 0.006084f
C1879 vdd.n1247 gnd 0.006084f
C1880 vdd.n1248 gnd 0.006084f
C1881 vdd.n1249 gnd 0.006084f
C1882 vdd.n1250 gnd 0.006084f
C1883 vdd.n1251 gnd 0.006084f
C1884 vdd.n1252 gnd 0.006084f
C1885 vdd.n1253 gnd 0.5623f
C1886 vdd.n1254 gnd 0.006084f
C1887 vdd.n1255 gnd 0.006084f
C1888 vdd.n1256 gnd 0.006084f
C1889 vdd.n1257 gnd 0.006084f
C1890 vdd.n1258 gnd 0.006084f
C1891 vdd.n1259 gnd 0.006084f
C1892 vdd.n1260 gnd 0.006084f
C1893 vdd.n1261 gnd 0.006084f
C1894 vdd.n1262 gnd 0.006084f
C1895 vdd.n1263 gnd 0.006084f
C1896 vdd.n1264 gnd 0.006084f
C1897 vdd.n1265 gnd 0.196576f
C1898 vdd.n1266 gnd 0.006084f
C1899 vdd.n1267 gnd 0.006084f
C1900 vdd.n1268 gnd 0.006084f
C1901 vdd.n1269 gnd 0.006084f
C1902 vdd.n1270 gnd 0.006084f
C1903 vdd.n1271 gnd 0.006084f
C1904 vdd.n1272 gnd 0.006084f
C1905 vdd.n1273 gnd 0.006084f
C1906 vdd.n1274 gnd 0.006084f
C1907 vdd.n1275 gnd 0.006084f
C1908 vdd.n1276 gnd 0.006084f
C1909 vdd.n1277 gnd 0.006084f
C1910 vdd.n1278 gnd 0.006084f
C1911 vdd.n1279 gnd 0.006084f
C1912 vdd.n1280 gnd 0.006084f
C1913 vdd.n1281 gnd 0.006084f
C1914 vdd.n1282 gnd 0.006084f
C1915 vdd.n1283 gnd 0.006084f
C1916 vdd.n1284 gnd 0.006084f
C1917 vdd.n1285 gnd 0.006084f
C1918 vdd.n1286 gnd 0.006084f
C1919 vdd.n1287 gnd 0.006084f
C1920 vdd.n1288 gnd 0.006084f
C1921 vdd.n1289 gnd 0.006084f
C1922 vdd.n1290 gnd 0.006084f
C1923 vdd.n1291 gnd 0.006084f
C1924 vdd.n1292 gnd 0.006084f
C1925 vdd.n1293 gnd 0.006084f
C1926 vdd.n1294 gnd 0.006084f
C1927 vdd.n1295 gnd 0.006084f
C1928 vdd.n1296 gnd 0.006084f
C1929 vdd.n1297 gnd 0.006084f
C1930 vdd.n1298 gnd 0.006084f
C1931 vdd.n1299 gnd 0.006084f
C1932 vdd.n1300 gnd 0.006084f
C1933 vdd.n1301 gnd 0.006084f
C1934 vdd.n1302 gnd 0.006084f
C1935 vdd.n1303 gnd 0.006084f
C1936 vdd.n1304 gnd 0.006084f
C1937 vdd.n1305 gnd 0.006084f
C1938 vdd.n1306 gnd 0.006084f
C1939 vdd.n1307 gnd 0.006084f
C1940 vdd.n1308 gnd 0.013026f
C1941 vdd.n1309 gnd 0.013026f
C1942 vdd.n1310 gnd 0.013814f
C1943 vdd.n1311 gnd 0.006084f
C1944 vdd.n1312 gnd 0.006084f
C1945 vdd.n1313 gnd 0.004697f
C1946 vdd.n1314 gnd 0.006084f
C1947 vdd.n1315 gnd 0.006084f
C1948 vdd.n1316 gnd 0.004429f
C1949 vdd.n1317 gnd 0.006084f
C1950 vdd.n1318 gnd 0.006084f
C1951 vdd.n1319 gnd 0.006084f
C1952 vdd.n1320 gnd 0.006084f
C1953 vdd.n1321 gnd 0.006084f
C1954 vdd.n1322 gnd 0.006084f
C1955 vdd.n1323 gnd 0.006084f
C1956 vdd.n1324 gnd 0.006084f
C1957 vdd.n1325 gnd 0.006084f
C1958 vdd.n1326 gnd 0.006084f
C1959 vdd.n1327 gnd 0.006084f
C1960 vdd.n1328 gnd 0.006084f
C1961 vdd.n1329 gnd 0.006084f
C1962 vdd.n1330 gnd 0.006084f
C1963 vdd.n1331 gnd 0.006084f
C1964 vdd.n1332 gnd 0.006084f
C1965 vdd.n1333 gnd 0.006084f
C1966 vdd.n1334 gnd 0.006084f
C1967 vdd.n1335 gnd 0.006084f
C1968 vdd.n1336 gnd 0.006084f
C1969 vdd.n1337 gnd 0.006084f
C1970 vdd.n1338 gnd 0.006084f
C1971 vdd.n1339 gnd 0.006084f
C1972 vdd.n1340 gnd 0.006084f
C1973 vdd.n1341 gnd 0.006084f
C1974 vdd.n1342 gnd 0.006084f
C1975 vdd.n1343 gnd 0.040983f
C1976 vdd.n1345 gnd 0.021413f
C1977 vdd.n1346 gnd 0.007201f
C1978 vdd.n1348 gnd 0.008947f
C1979 vdd.n1349 gnd 0.007201f
C1980 vdd.n1350 gnd 0.008947f
C1981 vdd.n1352 gnd 0.008947f
C1982 vdd.n1353 gnd 0.008947f
C1983 vdd.n1355 gnd 0.008947f
C1984 vdd.n1356 gnd 0.005977f
C1985 vdd.t9 gnd 0.457154f
C1986 vdd.n1357 gnd 0.008947f
C1987 vdd.n1358 gnd 0.021413f
C1988 vdd.n1359 gnd 0.007201f
C1989 vdd.n1360 gnd 0.008947f
C1990 vdd.n1361 gnd 0.007201f
C1991 vdd.n1362 gnd 0.008947f
C1992 vdd.n1363 gnd 0.914309f
C1993 vdd.n1364 gnd 0.008947f
C1994 vdd.n1365 gnd 0.007201f
C1995 vdd.n1366 gnd 0.007201f
C1996 vdd.n1367 gnd 0.008947f
C1997 vdd.n1368 gnd 0.007201f
C1998 vdd.n1369 gnd 0.008947f
C1999 vdd.t177 gnd 0.457154f
C2000 vdd.n1370 gnd 0.008947f
C2001 vdd.n1371 gnd 0.007201f
C2002 vdd.n1372 gnd 0.008947f
C2003 vdd.n1373 gnd 0.007201f
C2004 vdd.n1374 gnd 0.008947f
C2005 vdd.t207 gnd 0.457154f
C2006 vdd.n1375 gnd 0.008947f
C2007 vdd.n1376 gnd 0.007201f
C2008 vdd.n1377 gnd 0.008947f
C2009 vdd.n1378 gnd 0.007201f
C2010 vdd.n1379 gnd 0.008947f
C2011 vdd.t209 gnd 0.457154f
C2012 vdd.n1380 gnd 0.717732f
C2013 vdd.n1381 gnd 0.008947f
C2014 vdd.n1382 gnd 0.007201f
C2015 vdd.n1383 gnd 0.008947f
C2016 vdd.n1384 gnd 0.007201f
C2017 vdd.n1385 gnd 0.008947f
C2018 vdd.n1386 gnd 0.644588f
C2019 vdd.n1387 gnd 0.008947f
C2020 vdd.n1388 gnd 0.007201f
C2021 vdd.n1389 gnd 0.008947f
C2022 vdd.n1390 gnd 0.007201f
C2023 vdd.n1391 gnd 0.008947f
C2024 vdd.n1392 gnd 0.489155f
C2025 vdd.t173 gnd 0.457154f
C2026 vdd.n1393 gnd 0.008947f
C2027 vdd.n1394 gnd 0.007201f
C2028 vdd.n1395 gnd 0.008916f
C2029 vdd.n1396 gnd 0.007201f
C2030 vdd.n1397 gnd 0.008947f
C2031 vdd.t150 gnd 0.457154f
C2032 vdd.n1398 gnd 0.008947f
C2033 vdd.n1399 gnd 0.007201f
C2034 vdd.n1400 gnd 0.008947f
C2035 vdd.n1401 gnd 0.007201f
C2036 vdd.n1402 gnd 0.008947f
C2037 vdd.t154 gnd 0.457154f
C2038 vdd.n1403 gnd 0.580586f
C2039 vdd.n1404 gnd 0.008947f
C2040 vdd.n1405 gnd 0.007201f
C2041 vdd.n1406 gnd 0.008947f
C2042 vdd.n1407 gnd 0.007201f
C2043 vdd.n1408 gnd 0.008947f
C2044 vdd.t189 gnd 0.457154f
C2045 vdd.n1409 gnd 0.008947f
C2046 vdd.n1410 gnd 0.007201f
C2047 vdd.n1411 gnd 0.008947f
C2048 vdd.n1412 gnd 0.007201f
C2049 vdd.n1413 gnd 0.008947f
C2050 vdd.n1414 gnd 0.626301f
C2051 vdd.n1415 gnd 0.758876f
C2052 vdd.t205 gnd 0.457154f
C2053 vdd.n1416 gnd 0.008947f
C2054 vdd.n1417 gnd 0.007201f
C2055 vdd.n1418 gnd 0.008947f
C2056 vdd.n1419 gnd 0.007201f
C2057 vdd.n1420 gnd 0.008947f
C2058 vdd.n1421 gnd 0.470869f
C2059 vdd.n1422 gnd 0.008947f
C2060 vdd.n1423 gnd 0.007201f
C2061 vdd.n1424 gnd 0.008947f
C2062 vdd.n1425 gnd 0.007201f
C2063 vdd.n1426 gnd 0.008947f
C2064 vdd.n1427 gnd 0.914309f
C2065 vdd.t182 gnd 0.457154f
C2066 vdd.n1428 gnd 0.008947f
C2067 vdd.n1429 gnd 0.007201f
C2068 vdd.n1430 gnd 0.008947f
C2069 vdd.n1431 gnd 0.007201f
C2070 vdd.n1432 gnd 0.008947f
C2071 vdd.t37 gnd 0.457154f
C2072 vdd.n1433 gnd 0.008947f
C2073 vdd.n1434 gnd 0.007201f
C2074 vdd.n1435 gnd 0.021413f
C2075 vdd.n1436 gnd 0.021413f
C2076 vdd.n1437 gnd 2.10291f
C2077 vdd.n1438 gnd 0.516584f
C2078 vdd.n1439 gnd 0.021413f
C2079 vdd.n1440 gnd 0.008947f
C2080 vdd.n1442 gnd 0.008947f
C2081 vdd.n1443 gnd 0.008947f
C2082 vdd.n1444 gnd 0.007201f
C2083 vdd.n1445 gnd 0.008947f
C2084 vdd.n1446 gnd 0.008947f
C2085 vdd.n1448 gnd 0.008947f
C2086 vdd.n1449 gnd 0.008947f
C2087 vdd.n1451 gnd 0.008947f
C2088 vdd.n1452 gnd 0.007201f
C2089 vdd.n1453 gnd 0.008947f
C2090 vdd.n1454 gnd 0.008947f
C2091 vdd.n1456 gnd 0.008947f
C2092 vdd.n1457 gnd 0.008947f
C2093 vdd.n1459 gnd 0.008947f
C2094 vdd.n1460 gnd 0.007201f
C2095 vdd.n1461 gnd 0.008947f
C2096 vdd.n1462 gnd 0.008947f
C2097 vdd.n1464 gnd 0.008947f
C2098 vdd.n1465 gnd 0.008947f
C2099 vdd.n1467 gnd 0.008947f
C2100 vdd.n1468 gnd 0.007201f
C2101 vdd.n1469 gnd 0.008947f
C2102 vdd.n1470 gnd 0.008947f
C2103 vdd.n1472 gnd 0.008947f
C2104 vdd.n1473 gnd 0.008947f
C2105 vdd.n1475 gnd 0.008947f
C2106 vdd.t71 gnd 0.110068f
C2107 vdd.t72 gnd 0.117632f
C2108 vdd.t70 gnd 0.143747f
C2109 vdd.n1476 gnd 0.184263f
C2110 vdd.n1477 gnd 0.155535f
C2111 vdd.n1478 gnd 0.01541f
C2112 vdd.n1479 gnd 0.008947f
C2113 vdd.n1480 gnd 0.008947f
C2114 vdd.n1482 gnd 0.008947f
C2115 vdd.n1483 gnd 0.008947f
C2116 vdd.n1485 gnd 0.008947f
C2117 vdd.n1486 gnd 0.007201f
C2118 vdd.n1487 gnd 0.008947f
C2119 vdd.n1488 gnd 0.008947f
C2120 vdd.n1490 gnd 0.008947f
C2121 vdd.n1491 gnd 0.008947f
C2122 vdd.n1493 gnd 0.008947f
C2123 vdd.n1494 gnd 0.007201f
C2124 vdd.n1495 gnd 0.008947f
C2125 vdd.n1496 gnd 0.008947f
C2126 vdd.n1498 gnd 0.008947f
C2127 vdd.n1499 gnd 0.008947f
C2128 vdd.n1501 gnd 0.008947f
C2129 vdd.n1502 gnd 0.007201f
C2130 vdd.n1503 gnd 0.008947f
C2131 vdd.n1504 gnd 0.008947f
C2132 vdd.n1506 gnd 0.008947f
C2133 vdd.n1507 gnd 0.008947f
C2134 vdd.n1509 gnd 0.008947f
C2135 vdd.n1510 gnd 0.007201f
C2136 vdd.n1511 gnd 0.008947f
C2137 vdd.n1512 gnd 0.008947f
C2138 vdd.n1514 gnd 0.008947f
C2139 vdd.n1515 gnd 0.008947f
C2140 vdd.n1517 gnd 0.008947f
C2141 vdd.n1518 gnd 0.007201f
C2142 vdd.n1519 gnd 0.008947f
C2143 vdd.n1520 gnd 0.008947f
C2144 vdd.n1522 gnd 0.008947f
C2145 vdd.n1523 gnd 0.007129f
C2146 vdd.n1525 gnd 0.007201f
C2147 vdd.n1526 gnd 0.008947f
C2148 vdd.n1527 gnd 0.008947f
C2149 vdd.n1528 gnd 0.008947f
C2150 vdd.n1529 gnd 0.008947f
C2151 vdd.n1531 gnd 0.008947f
C2152 vdd.n1532 gnd 0.008947f
C2153 vdd.n1533 gnd 0.007201f
C2154 vdd.n1534 gnd 0.008947f
C2155 vdd.n1536 gnd 0.008947f
C2156 vdd.n1537 gnd 0.008947f
C2157 vdd.n1539 gnd 0.008947f
C2158 vdd.n1540 gnd 0.008947f
C2159 vdd.n1541 gnd 0.007201f
C2160 vdd.n1542 gnd 0.008947f
C2161 vdd.n1544 gnd 0.008947f
C2162 vdd.n1545 gnd 0.008947f
C2163 vdd.n1547 gnd 0.008947f
C2164 vdd.n1548 gnd 0.008947f
C2165 vdd.n1549 gnd 0.007201f
C2166 vdd.n1550 gnd 0.008947f
C2167 vdd.n1552 gnd 0.008947f
C2168 vdd.n1553 gnd 0.008947f
C2169 vdd.n1555 gnd 0.008947f
C2170 vdd.n1556 gnd 0.008947f
C2171 vdd.n1557 gnd 0.007201f
C2172 vdd.n1558 gnd 0.008947f
C2173 vdd.n1560 gnd 0.008947f
C2174 vdd.n1561 gnd 0.008947f
C2175 vdd.n1563 gnd 0.008947f
C2176 vdd.n1564 gnd 0.00342f
C2177 vdd.t38 gnd 0.110068f
C2178 vdd.t39 gnd 0.117632f
C2179 vdd.t36 gnd 0.143747f
C2180 vdd.n1565 gnd 0.184263f
C2181 vdd.n1566 gnd 0.155535f
C2182 vdd.n1567 gnd 0.01181f
C2183 vdd.n1568 gnd 0.003781f
C2184 vdd.n1569 gnd 0.007201f
C2185 vdd.n1570 gnd 0.008947f
C2186 vdd.n1571 gnd 0.008947f
C2187 vdd.n1572 gnd 0.008947f
C2188 vdd.n1573 gnd 0.007201f
C2189 vdd.n1574 gnd 0.007201f
C2190 vdd.n1575 gnd 0.007201f
C2191 vdd.n1576 gnd 0.008947f
C2192 vdd.n1577 gnd 0.008947f
C2193 vdd.n1578 gnd 0.008947f
C2194 vdd.n1579 gnd 0.007201f
C2195 vdd.n1580 gnd 0.007201f
C2196 vdd.n1581 gnd 0.007201f
C2197 vdd.n1582 gnd 0.008947f
C2198 vdd.n1583 gnd 0.008947f
C2199 vdd.n1584 gnd 0.008947f
C2200 vdd.n1585 gnd 0.007201f
C2201 vdd.n1586 gnd 0.007201f
C2202 vdd.n1587 gnd 0.007201f
C2203 vdd.n1588 gnd 0.008947f
C2204 vdd.n1589 gnd 0.008947f
C2205 vdd.n1590 gnd 0.008947f
C2206 vdd.n1591 gnd 0.007201f
C2207 vdd.n1592 gnd 0.007201f
C2208 vdd.n1593 gnd 0.007201f
C2209 vdd.n1594 gnd 0.008947f
C2210 vdd.n1595 gnd 0.008947f
C2211 vdd.n1596 gnd 0.008947f
C2212 vdd.n1597 gnd 0.007201f
C2213 vdd.n1598 gnd 0.008947f
C2214 vdd.n1599 gnd 0.008947f
C2215 vdd.n1601 gnd 0.008947f
C2216 vdd.t61 gnd 0.110068f
C2217 vdd.t62 gnd 0.117632f
C2218 vdd.t60 gnd 0.143747f
C2219 vdd.n1602 gnd 0.184263f
C2220 vdd.n1603 gnd 0.155535f
C2221 vdd.n1604 gnd 0.01541f
C2222 vdd.n1605 gnd 0.004897f
C2223 vdd.n1606 gnd 0.008947f
C2224 vdd.n1607 gnd 0.008947f
C2225 vdd.n1608 gnd 0.008947f
C2226 vdd.n1609 gnd 0.007201f
C2227 vdd.n1610 gnd 0.007201f
C2228 vdd.n1611 gnd 0.007201f
C2229 vdd.n1612 gnd 0.008947f
C2230 vdd.n1613 gnd 0.008947f
C2231 vdd.n1614 gnd 0.008947f
C2232 vdd.n1615 gnd 0.007201f
C2233 vdd.n1616 gnd 0.007201f
C2234 vdd.n1617 gnd 0.007201f
C2235 vdd.n1618 gnd 0.008947f
C2236 vdd.n1619 gnd 0.008947f
C2237 vdd.n1620 gnd 0.008947f
C2238 vdd.n1621 gnd 0.007201f
C2239 vdd.n1622 gnd 0.007201f
C2240 vdd.n1623 gnd 0.007201f
C2241 vdd.n1624 gnd 0.008947f
C2242 vdd.n1625 gnd 0.008947f
C2243 vdd.n1626 gnd 0.008947f
C2244 vdd.n1627 gnd 0.007201f
C2245 vdd.n1628 gnd 0.007201f
C2246 vdd.n1629 gnd 0.007201f
C2247 vdd.n1630 gnd 0.008947f
C2248 vdd.n1631 gnd 0.008947f
C2249 vdd.n1632 gnd 0.008947f
C2250 vdd.n1633 gnd 0.007201f
C2251 vdd.n1634 gnd 0.007201f
C2252 vdd.n1635 gnd 0.006013f
C2253 vdd.n1636 gnd 0.008947f
C2254 vdd.n1637 gnd 0.008947f
C2255 vdd.n1638 gnd 0.008947f
C2256 vdd.n1639 gnd 0.006013f
C2257 vdd.n1640 gnd 0.007201f
C2258 vdd.n1641 gnd 0.007201f
C2259 vdd.n1642 gnd 0.008947f
C2260 vdd.n1643 gnd 0.008947f
C2261 vdd.n1644 gnd 0.008947f
C2262 vdd.n1645 gnd 0.007201f
C2263 vdd.n1646 gnd 0.007201f
C2264 vdd.n1647 gnd 0.007201f
C2265 vdd.n1648 gnd 0.008947f
C2266 vdd.n1649 gnd 0.008947f
C2267 vdd.n1650 gnd 0.008947f
C2268 vdd.n1651 gnd 0.007201f
C2269 vdd.n1652 gnd 0.007201f
C2270 vdd.n1653 gnd 0.007201f
C2271 vdd.n1654 gnd 0.008947f
C2272 vdd.n1655 gnd 0.008947f
C2273 vdd.n1656 gnd 0.008947f
C2274 vdd.n1657 gnd 0.007201f
C2275 vdd.n1658 gnd 0.007201f
C2276 vdd.n1659 gnd 0.007201f
C2277 vdd.n1660 gnd 0.008947f
C2278 vdd.n1661 gnd 0.008947f
C2279 vdd.n1662 gnd 0.008947f
C2280 vdd.n1663 gnd 0.007201f
C2281 vdd.n1664 gnd 0.007201f
C2282 vdd.n1665 gnd 0.005977f
C2283 vdd.n1666 gnd 0.021413f
C2284 vdd.n1667 gnd 0.021084f
C2285 vdd.n1668 gnd 0.005977f
C2286 vdd.n1669 gnd 0.021084f
C2287 vdd.n1670 gnd 1.28918f
C2288 vdd.n1671 gnd 0.021084f
C2289 vdd.n1672 gnd 0.005977f
C2290 vdd.n1673 gnd 0.021084f
C2291 vdd.n1674 gnd 0.008947f
C2292 vdd.n1675 gnd 0.008947f
C2293 vdd.n1676 gnd 0.007201f
C2294 vdd.n1677 gnd 0.008947f
C2295 vdd.n1678 gnd 0.854879f
C2296 vdd.n1679 gnd 0.008947f
C2297 vdd.n1680 gnd 0.007201f
C2298 vdd.n1681 gnd 0.008947f
C2299 vdd.n1682 gnd 0.008947f
C2300 vdd.n1683 gnd 0.008947f
C2301 vdd.n1684 gnd 0.007201f
C2302 vdd.n1685 gnd 0.008947f
C2303 vdd.n1686 gnd 0.900594f
C2304 vdd.n1687 gnd 0.008947f
C2305 vdd.n1688 gnd 0.007201f
C2306 vdd.n1689 gnd 0.008947f
C2307 vdd.n1690 gnd 0.008947f
C2308 vdd.n1691 gnd 0.008947f
C2309 vdd.n1692 gnd 0.007201f
C2310 vdd.n1693 gnd 0.008947f
C2311 vdd.t148 gnd 0.457154f
C2312 vdd.n1694 gnd 0.745162f
C2313 vdd.n1695 gnd 0.008947f
C2314 vdd.n1696 gnd 0.007201f
C2315 vdd.n1697 gnd 0.008947f
C2316 vdd.n1698 gnd 0.008947f
C2317 vdd.n1699 gnd 0.008947f
C2318 vdd.n1700 gnd 0.007201f
C2319 vdd.n1701 gnd 0.008947f
C2320 vdd.n1702 gnd 0.589729f
C2321 vdd.n1703 gnd 0.008947f
C2322 vdd.n1704 gnd 0.007201f
C2323 vdd.n1705 gnd 0.008947f
C2324 vdd.n1706 gnd 0.008947f
C2325 vdd.n1707 gnd 0.008947f
C2326 vdd.n1708 gnd 0.007201f
C2327 vdd.n1709 gnd 0.008947f
C2328 vdd.n1710 gnd 0.736018f
C2329 vdd.n1711 gnd 0.480012f
C2330 vdd.n1712 gnd 0.008947f
C2331 vdd.n1713 gnd 0.007201f
C2332 vdd.n1714 gnd 0.008947f
C2333 vdd.n1715 gnd 0.008947f
C2334 vdd.n1716 gnd 0.008947f
C2335 vdd.n1717 gnd 0.007201f
C2336 vdd.n1718 gnd 0.008947f
C2337 vdd.n1719 gnd 0.635445f
C2338 vdd.n1720 gnd 0.008947f
C2339 vdd.n1721 gnd 0.007201f
C2340 vdd.n1722 gnd 0.008947f
C2341 vdd.n1723 gnd 0.008947f
C2342 vdd.n1724 gnd 0.008947f
C2343 vdd.n1725 gnd 0.007201f
C2344 vdd.n1726 gnd 0.008947f
C2345 vdd.t175 gnd 0.457154f
C2346 vdd.n1727 gnd 0.758876f
C2347 vdd.n1728 gnd 0.008947f
C2348 vdd.n1729 gnd 0.007201f
C2349 vdd.n1730 gnd 0.00491f
C2350 vdd.n1731 gnd 0.004556f
C2351 vdd.n1732 gnd 0.00252f
C2352 vdd.n1733 gnd 0.005787f
C2353 vdd.n1734 gnd 0.002448f
C2354 vdd.n1735 gnd 0.002592f
C2355 vdd.n1736 gnd 0.004556f
C2356 vdd.n1737 gnd 0.002448f
C2357 vdd.n1738 gnd 0.005787f
C2358 vdd.n1739 gnd 0.002592f
C2359 vdd.n1740 gnd 0.004556f
C2360 vdd.n1741 gnd 0.002448f
C2361 vdd.n1742 gnd 0.00434f
C2362 vdd.n1743 gnd 0.004353f
C2363 vdd.t202 gnd 0.012433f
C2364 vdd.n1744 gnd 0.027663f
C2365 vdd.n1745 gnd 0.143964f
C2366 vdd.n1746 gnd 0.002448f
C2367 vdd.n1747 gnd 0.002592f
C2368 vdd.n1748 gnd 0.005787f
C2369 vdd.n1749 gnd 0.005787f
C2370 vdd.n1750 gnd 0.002592f
C2371 vdd.n1751 gnd 0.002448f
C2372 vdd.n1752 gnd 0.004556f
C2373 vdd.n1753 gnd 0.004556f
C2374 vdd.n1754 gnd 0.002448f
C2375 vdd.n1755 gnd 0.002592f
C2376 vdd.n1756 gnd 0.005787f
C2377 vdd.n1757 gnd 0.005787f
C2378 vdd.n1758 gnd 0.002592f
C2379 vdd.n1759 gnd 0.002448f
C2380 vdd.n1760 gnd 0.004556f
C2381 vdd.n1761 gnd 0.004556f
C2382 vdd.n1762 gnd 0.002448f
C2383 vdd.n1763 gnd 0.002592f
C2384 vdd.n1764 gnd 0.005787f
C2385 vdd.n1765 gnd 0.005787f
C2386 vdd.n1766 gnd 0.013682f
C2387 vdd.n1767 gnd 0.00252f
C2388 vdd.n1768 gnd 0.002448f
C2389 vdd.n1769 gnd 0.011777f
C2390 vdd.n1770 gnd 0.008222f
C2391 vdd.t233 gnd 0.028804f
C2392 vdd.t243 gnd 0.028804f
C2393 vdd.n1771 gnd 0.197961f
C2394 vdd.n1772 gnd 0.155666f
C2395 vdd.t218 gnd 0.028804f
C2396 vdd.t167 gnd 0.028804f
C2397 vdd.n1773 gnd 0.197961f
C2398 vdd.n1774 gnd 0.125622f
C2399 vdd.t211 gnd 0.028804f
C2400 vdd.t176 gnd 0.028804f
C2401 vdd.n1775 gnd 0.197961f
C2402 vdd.n1776 gnd 0.125622f
C2403 vdd.t237 gnd 0.028804f
C2404 vdd.t194 gnd 0.028804f
C2405 vdd.n1777 gnd 0.197961f
C2406 vdd.n1778 gnd 0.125622f
C2407 vdd.t224 gnd 0.028804f
C2408 vdd.t206 gnd 0.028804f
C2409 vdd.n1779 gnd 0.197961f
C2410 vdd.n1780 gnd 0.125622f
C2411 vdd.n1781 gnd 0.00491f
C2412 vdd.n1782 gnd 0.004556f
C2413 vdd.n1783 gnd 0.00252f
C2414 vdd.n1784 gnd 0.005787f
C2415 vdd.n1785 gnd 0.002448f
C2416 vdd.n1786 gnd 0.002592f
C2417 vdd.n1787 gnd 0.004556f
C2418 vdd.n1788 gnd 0.002448f
C2419 vdd.n1789 gnd 0.005787f
C2420 vdd.n1790 gnd 0.002592f
C2421 vdd.n1791 gnd 0.004556f
C2422 vdd.n1792 gnd 0.002448f
C2423 vdd.n1793 gnd 0.00434f
C2424 vdd.n1794 gnd 0.004353f
C2425 vdd.t183 gnd 0.012433f
C2426 vdd.n1795 gnd 0.027663f
C2427 vdd.n1796 gnd 0.143964f
C2428 vdd.n1797 gnd 0.002448f
C2429 vdd.n1798 gnd 0.002592f
C2430 vdd.n1799 gnd 0.005787f
C2431 vdd.n1800 gnd 0.005787f
C2432 vdd.n1801 gnd 0.002592f
C2433 vdd.n1802 gnd 0.002448f
C2434 vdd.n1803 gnd 0.004556f
C2435 vdd.n1804 gnd 0.004556f
C2436 vdd.n1805 gnd 0.002448f
C2437 vdd.n1806 gnd 0.002592f
C2438 vdd.n1807 gnd 0.005787f
C2439 vdd.n1808 gnd 0.005787f
C2440 vdd.n1809 gnd 0.002592f
C2441 vdd.n1810 gnd 0.002448f
C2442 vdd.n1811 gnd 0.004556f
C2443 vdd.n1812 gnd 0.004556f
C2444 vdd.n1813 gnd 0.002448f
C2445 vdd.n1814 gnd 0.002592f
C2446 vdd.n1815 gnd 0.005787f
C2447 vdd.n1816 gnd 0.005787f
C2448 vdd.n1817 gnd 0.013682f
C2449 vdd.n1818 gnd 0.00252f
C2450 vdd.n1819 gnd 0.002448f
C2451 vdd.n1820 gnd 0.011777f
C2452 vdd.n1821 gnd 0.007964f
C2453 vdd.n1822 gnd 0.093463f
C2454 vdd.n1823 gnd 0.00491f
C2455 vdd.n1824 gnd 0.004556f
C2456 vdd.n1825 gnd 0.00252f
C2457 vdd.n1826 gnd 0.005787f
C2458 vdd.n1827 gnd 0.002448f
C2459 vdd.n1828 gnd 0.002592f
C2460 vdd.n1829 gnd 0.004556f
C2461 vdd.n1830 gnd 0.002448f
C2462 vdd.n1831 gnd 0.005787f
C2463 vdd.n1832 gnd 0.002592f
C2464 vdd.n1833 gnd 0.004556f
C2465 vdd.n1834 gnd 0.002448f
C2466 vdd.n1835 gnd 0.00434f
C2467 vdd.n1836 gnd 0.004353f
C2468 vdd.t178 gnd 0.012433f
C2469 vdd.n1837 gnd 0.027663f
C2470 vdd.n1838 gnd 0.143964f
C2471 vdd.n1839 gnd 0.002448f
C2472 vdd.n1840 gnd 0.002592f
C2473 vdd.n1841 gnd 0.005787f
C2474 vdd.n1842 gnd 0.005787f
C2475 vdd.n1843 gnd 0.002592f
C2476 vdd.n1844 gnd 0.002448f
C2477 vdd.n1845 gnd 0.004556f
C2478 vdd.n1846 gnd 0.004556f
C2479 vdd.n1847 gnd 0.002448f
C2480 vdd.n1848 gnd 0.002592f
C2481 vdd.n1849 gnd 0.005787f
C2482 vdd.n1850 gnd 0.005787f
C2483 vdd.n1851 gnd 0.002592f
C2484 vdd.n1852 gnd 0.002448f
C2485 vdd.n1853 gnd 0.004556f
C2486 vdd.n1854 gnd 0.004556f
C2487 vdd.n1855 gnd 0.002448f
C2488 vdd.n1856 gnd 0.002592f
C2489 vdd.n1857 gnd 0.005787f
C2490 vdd.n1858 gnd 0.005787f
C2491 vdd.n1859 gnd 0.013682f
C2492 vdd.n1860 gnd 0.00252f
C2493 vdd.n1861 gnd 0.002448f
C2494 vdd.n1862 gnd 0.011777f
C2495 vdd.n1863 gnd 0.008222f
C2496 vdd.t210 gnd 0.028804f
C2497 vdd.t208 gnd 0.028804f
C2498 vdd.n1864 gnd 0.197961f
C2499 vdd.n1865 gnd 0.155666f
C2500 vdd.t174 gnd 0.028804f
C2501 vdd.t157 gnd 0.028804f
C2502 vdd.n1866 gnd 0.197961f
C2503 vdd.n1867 gnd 0.125622f
C2504 vdd.t151 gnd 0.028804f
C2505 vdd.t203 gnd 0.028804f
C2506 vdd.n1868 gnd 0.197961f
C2507 vdd.n1869 gnd 0.125622f
C2508 vdd.t190 gnd 0.028804f
C2509 vdd.t155 gnd 0.028804f
C2510 vdd.n1870 gnd 0.197961f
C2511 vdd.n1871 gnd 0.125622f
C2512 vdd.t149 gnd 0.028804f
C2513 vdd.t219 gnd 0.028804f
C2514 vdd.n1872 gnd 0.197961f
C2515 vdd.n1873 gnd 0.125622f
C2516 vdd.n1874 gnd 0.00491f
C2517 vdd.n1875 gnd 0.004556f
C2518 vdd.n1876 gnd 0.00252f
C2519 vdd.n1877 gnd 0.005787f
C2520 vdd.n1878 gnd 0.002448f
C2521 vdd.n1879 gnd 0.002592f
C2522 vdd.n1880 gnd 0.004556f
C2523 vdd.n1881 gnd 0.002448f
C2524 vdd.n1882 gnd 0.005787f
C2525 vdd.n1883 gnd 0.002592f
C2526 vdd.n1884 gnd 0.004556f
C2527 vdd.n1885 gnd 0.002448f
C2528 vdd.n1886 gnd 0.00434f
C2529 vdd.n1887 gnd 0.004353f
C2530 vdd.t185 gnd 0.012433f
C2531 vdd.n1888 gnd 0.027663f
C2532 vdd.n1889 gnd 0.143964f
C2533 vdd.n1890 gnd 0.002448f
C2534 vdd.n1891 gnd 0.002592f
C2535 vdd.n1892 gnd 0.005787f
C2536 vdd.n1893 gnd 0.005787f
C2537 vdd.n1894 gnd 0.002592f
C2538 vdd.n1895 gnd 0.002448f
C2539 vdd.n1896 gnd 0.004556f
C2540 vdd.n1897 gnd 0.004556f
C2541 vdd.n1898 gnd 0.002448f
C2542 vdd.n1899 gnd 0.002592f
C2543 vdd.n1900 gnd 0.005787f
C2544 vdd.n1901 gnd 0.005787f
C2545 vdd.n1902 gnd 0.002592f
C2546 vdd.n1903 gnd 0.002448f
C2547 vdd.n1904 gnd 0.004556f
C2548 vdd.n1905 gnd 0.004556f
C2549 vdd.n1906 gnd 0.002448f
C2550 vdd.n1907 gnd 0.002592f
C2551 vdd.n1908 gnd 0.005787f
C2552 vdd.n1909 gnd 0.005787f
C2553 vdd.n1910 gnd 0.013682f
C2554 vdd.n1911 gnd 0.00252f
C2555 vdd.n1912 gnd 0.002448f
C2556 vdd.n1913 gnd 0.011777f
C2557 vdd.n1914 gnd 0.007964f
C2558 vdd.n1915 gnd 0.055601f
C2559 vdd.n1916 gnd 0.200345f
C2560 vdd.n1917 gnd 0.00491f
C2561 vdd.n1918 gnd 0.004556f
C2562 vdd.n1919 gnd 0.00252f
C2563 vdd.n1920 gnd 0.005787f
C2564 vdd.n1921 gnd 0.002448f
C2565 vdd.n1922 gnd 0.002592f
C2566 vdd.n1923 gnd 0.004556f
C2567 vdd.n1924 gnd 0.002448f
C2568 vdd.n1925 gnd 0.005787f
C2569 vdd.n1926 gnd 0.002592f
C2570 vdd.n1927 gnd 0.004556f
C2571 vdd.n1928 gnd 0.002448f
C2572 vdd.n1929 gnd 0.00434f
C2573 vdd.n1930 gnd 0.004353f
C2574 vdd.t191 gnd 0.012433f
C2575 vdd.n1931 gnd 0.027663f
C2576 vdd.n1932 gnd 0.143964f
C2577 vdd.n1933 gnd 0.002448f
C2578 vdd.n1934 gnd 0.002592f
C2579 vdd.n1935 gnd 0.005787f
C2580 vdd.n1936 gnd 0.005787f
C2581 vdd.n1937 gnd 0.002592f
C2582 vdd.n1938 gnd 0.002448f
C2583 vdd.n1939 gnd 0.004556f
C2584 vdd.n1940 gnd 0.004556f
C2585 vdd.n1941 gnd 0.002448f
C2586 vdd.n1942 gnd 0.002592f
C2587 vdd.n1943 gnd 0.005787f
C2588 vdd.n1944 gnd 0.005787f
C2589 vdd.n1945 gnd 0.002592f
C2590 vdd.n1946 gnd 0.002448f
C2591 vdd.n1947 gnd 0.004556f
C2592 vdd.n1948 gnd 0.004556f
C2593 vdd.n1949 gnd 0.002448f
C2594 vdd.n1950 gnd 0.002592f
C2595 vdd.n1951 gnd 0.005787f
C2596 vdd.n1952 gnd 0.005787f
C2597 vdd.n1953 gnd 0.013682f
C2598 vdd.n1954 gnd 0.00252f
C2599 vdd.n1955 gnd 0.002448f
C2600 vdd.n1956 gnd 0.011777f
C2601 vdd.n1957 gnd 0.008222f
C2602 vdd.t215 gnd 0.028804f
C2603 vdd.t214 gnd 0.028804f
C2604 vdd.n1958 gnd 0.197961f
C2605 vdd.n1959 gnd 0.155666f
C2606 vdd.t188 gnd 0.028804f
C2607 vdd.t170 gnd 0.028804f
C2608 vdd.n1960 gnd 0.197961f
C2609 vdd.n1961 gnd 0.125622f
C2610 vdd.t168 gnd 0.028804f
C2611 vdd.t213 gnd 0.028804f
C2612 vdd.n1962 gnd 0.197961f
C2613 vdd.n1963 gnd 0.125622f
C2614 vdd.t197 gnd 0.028804f
C2615 vdd.t169 gnd 0.028804f
C2616 vdd.n1964 gnd 0.197961f
C2617 vdd.n1965 gnd 0.125622f
C2618 vdd.t164 gnd 0.028804f
C2619 vdd.t226 gnd 0.028804f
C2620 vdd.n1966 gnd 0.197961f
C2621 vdd.n1967 gnd 0.125622f
C2622 vdd.n1968 gnd 0.00491f
C2623 vdd.n1969 gnd 0.004556f
C2624 vdd.n1970 gnd 0.00252f
C2625 vdd.n1971 gnd 0.005787f
C2626 vdd.n1972 gnd 0.002448f
C2627 vdd.n1973 gnd 0.002592f
C2628 vdd.n1974 gnd 0.004556f
C2629 vdd.n1975 gnd 0.002448f
C2630 vdd.n1976 gnd 0.005787f
C2631 vdd.n1977 gnd 0.002592f
C2632 vdd.n1978 gnd 0.004556f
C2633 vdd.n1979 gnd 0.002448f
C2634 vdd.n1980 gnd 0.00434f
C2635 vdd.n1981 gnd 0.004353f
C2636 vdd.t195 gnd 0.012433f
C2637 vdd.n1982 gnd 0.027663f
C2638 vdd.n1983 gnd 0.143964f
C2639 vdd.n1984 gnd 0.002448f
C2640 vdd.n1985 gnd 0.002592f
C2641 vdd.n1986 gnd 0.005787f
C2642 vdd.n1987 gnd 0.005787f
C2643 vdd.n1988 gnd 0.002592f
C2644 vdd.n1989 gnd 0.002448f
C2645 vdd.n1990 gnd 0.004556f
C2646 vdd.n1991 gnd 0.004556f
C2647 vdd.n1992 gnd 0.002448f
C2648 vdd.n1993 gnd 0.002592f
C2649 vdd.n1994 gnd 0.005787f
C2650 vdd.n1995 gnd 0.005787f
C2651 vdd.n1996 gnd 0.002592f
C2652 vdd.n1997 gnd 0.002448f
C2653 vdd.n1998 gnd 0.004556f
C2654 vdd.n1999 gnd 0.004556f
C2655 vdd.n2000 gnd 0.002448f
C2656 vdd.n2001 gnd 0.002592f
C2657 vdd.n2002 gnd 0.005787f
C2658 vdd.n2003 gnd 0.005787f
C2659 vdd.n2004 gnd 0.013682f
C2660 vdd.n2005 gnd 0.00252f
C2661 vdd.n2006 gnd 0.002448f
C2662 vdd.n2007 gnd 0.011777f
C2663 vdd.n2008 gnd 0.007964f
C2664 vdd.n2009 gnd 0.055601f
C2665 vdd.n2010 gnd 0.220186f
C2666 vdd.n2011 gnd 2.30604f
C2667 vdd.n2012 gnd 0.532576f
C2668 vdd.n2013 gnd 0.008916f
C2669 vdd.n2014 gnd 0.008947f
C2670 vdd.n2015 gnd 0.007201f
C2671 vdd.n2016 gnd 0.008947f
C2672 vdd.n2017 gnd 0.726875f
C2673 vdd.n2018 gnd 0.008947f
C2674 vdd.n2019 gnd 0.007201f
C2675 vdd.n2020 gnd 0.008947f
C2676 vdd.n2021 gnd 0.008947f
C2677 vdd.n2022 gnd 0.008947f
C2678 vdd.n2023 gnd 0.007201f
C2679 vdd.n2024 gnd 0.008947f
C2680 vdd.n2025 gnd 0.758876f
C2681 vdd.t156 gnd 0.457154f
C2682 vdd.n2026 gnd 0.571443f
C2683 vdd.n2027 gnd 0.008947f
C2684 vdd.n2028 gnd 0.007201f
C2685 vdd.n2029 gnd 0.008947f
C2686 vdd.n2030 gnd 0.008947f
C2687 vdd.n2031 gnd 0.008947f
C2688 vdd.n2032 gnd 0.007201f
C2689 vdd.n2033 gnd 0.008947f
C2690 vdd.n2034 gnd 0.498298f
C2691 vdd.n2035 gnd 0.008947f
C2692 vdd.n2036 gnd 0.007201f
C2693 vdd.n2037 gnd 0.008947f
C2694 vdd.n2038 gnd 0.008947f
C2695 vdd.n2039 gnd 0.008947f
C2696 vdd.n2040 gnd 0.007201f
C2697 vdd.n2041 gnd 0.008947f
C2698 vdd.n2042 gnd 0.5623f
C2699 vdd.n2043 gnd 0.653731f
C2700 vdd.n2044 gnd 0.008947f
C2701 vdd.n2045 gnd 0.007201f
C2702 vdd.n2046 gnd 0.008947f
C2703 vdd.n2047 gnd 0.008947f
C2704 vdd.n2048 gnd 0.008947f
C2705 vdd.n2049 gnd 0.007201f
C2706 vdd.n2050 gnd 0.008947f
C2707 vdd.n2051 gnd 0.809163f
C2708 vdd.n2052 gnd 0.008947f
C2709 vdd.n2053 gnd 0.007201f
C2710 vdd.n2054 gnd 0.008947f
C2711 vdd.n2055 gnd 0.008947f
C2712 vdd.n2056 gnd 0.021084f
C2713 vdd.n2057 gnd 0.008947f
C2714 vdd.n2058 gnd 0.008947f
C2715 vdd.n2059 gnd 0.007201f
C2716 vdd.n2060 gnd 0.008947f
C2717 vdd.n2061 gnd 0.489155f
C2718 vdd.n2062 gnd 0.914309f
C2719 vdd.n2063 gnd 0.008947f
C2720 vdd.n2064 gnd 0.007201f
C2721 vdd.n2065 gnd 0.008947f
C2722 vdd.n2066 gnd 0.008947f
C2723 vdd.n2067 gnd 0.021084f
C2724 vdd.n2068 gnd 0.005977f
C2725 vdd.n2069 gnd 0.021084f
C2726 vdd.n2070 gnd 1.25717f
C2727 vdd.n2071 gnd 0.021084f
C2728 vdd.n2072 gnd 0.021413f
C2729 vdd.n2073 gnd 0.00342f
C2730 vdd.t32 gnd 0.110068f
C2731 vdd.t31 gnd 0.117632f
C2732 vdd.t30 gnd 0.143747f
C2733 vdd.n2074 gnd 0.184263f
C2734 vdd.n2075 gnd 0.154815f
C2735 vdd.n2076 gnd 0.01109f
C2736 vdd.n2077 gnd 0.003781f
C2737 vdd.n2078 gnd 0.007694f
C2738 vdd.n2079 gnd 0.949782f
C2739 vdd.n2081 gnd 0.007201f
C2740 vdd.n2082 gnd 0.007201f
C2741 vdd.n2083 gnd 0.008947f
C2742 vdd.n2085 gnd 0.008947f
C2743 vdd.n2086 gnd 0.008947f
C2744 vdd.n2087 gnd 0.007201f
C2745 vdd.n2088 gnd 0.007201f
C2746 vdd.n2089 gnd 0.007201f
C2747 vdd.n2090 gnd 0.008947f
C2748 vdd.n2092 gnd 0.008947f
C2749 vdd.n2093 gnd 0.008947f
C2750 vdd.n2094 gnd 0.007201f
C2751 vdd.n2095 gnd 0.007201f
C2752 vdd.n2096 gnd 0.007201f
C2753 vdd.n2097 gnd 0.008947f
C2754 vdd.n2099 gnd 0.008947f
C2755 vdd.n2100 gnd 0.008947f
C2756 vdd.n2101 gnd 0.007201f
C2757 vdd.n2102 gnd 0.007201f
C2758 vdd.n2103 gnd 0.007201f
C2759 vdd.n2104 gnd 0.008947f
C2760 vdd.n2106 gnd 0.008947f
C2761 vdd.n2107 gnd 0.008947f
C2762 vdd.n2108 gnd 0.007201f
C2763 vdd.n2109 gnd 0.008947f
C2764 vdd.n2110 gnd 0.008947f
C2765 vdd.n2111 gnd 0.008947f
C2766 vdd.n2112 gnd 0.01469f
C2767 vdd.n2113 gnd 0.004897f
C2768 vdd.n2114 gnd 0.007201f
C2769 vdd.n2115 gnd 0.008947f
C2770 vdd.n2117 gnd 0.008947f
C2771 vdd.n2118 gnd 0.008947f
C2772 vdd.n2119 gnd 0.007201f
C2773 vdd.n2120 gnd 0.007201f
C2774 vdd.n2121 gnd 0.007201f
C2775 vdd.n2122 gnd 0.008947f
C2776 vdd.n2124 gnd 0.008947f
C2777 vdd.n2125 gnd 0.008947f
C2778 vdd.n2126 gnd 0.007201f
C2779 vdd.n2127 gnd 0.007201f
C2780 vdd.n2128 gnd 0.007201f
C2781 vdd.n2129 gnd 0.008947f
C2782 vdd.n2131 gnd 0.008947f
C2783 vdd.n2132 gnd 0.008947f
C2784 vdd.n2133 gnd 0.007201f
C2785 vdd.n2134 gnd 0.007201f
C2786 vdd.n2135 gnd 0.007201f
C2787 vdd.n2136 gnd 0.008947f
C2788 vdd.n2138 gnd 0.008947f
C2789 vdd.n2139 gnd 0.008947f
C2790 vdd.n2140 gnd 0.007201f
C2791 vdd.n2141 gnd 0.007201f
C2792 vdd.n2142 gnd 0.007201f
C2793 vdd.n2143 gnd 0.008947f
C2794 vdd.n2145 gnd 0.008947f
C2795 vdd.n2146 gnd 0.008947f
C2796 vdd.n2147 gnd 0.007201f
C2797 vdd.n2148 gnd 0.008947f
C2798 vdd.n2149 gnd 0.008947f
C2799 vdd.n2150 gnd 0.008947f
C2800 vdd.n2151 gnd 0.01469f
C2801 vdd.n2152 gnd 0.006013f
C2802 vdd.n2153 gnd 0.007201f
C2803 vdd.n2154 gnd 0.008947f
C2804 vdd.n2156 gnd 0.008947f
C2805 vdd.n2157 gnd 0.008947f
C2806 vdd.n2158 gnd 0.007201f
C2807 vdd.n2159 gnd 0.007201f
C2808 vdd.n2160 gnd 0.007201f
C2809 vdd.n2161 gnd 0.008947f
C2810 vdd.n2163 gnd 0.008947f
C2811 vdd.n2164 gnd 0.008947f
C2812 vdd.n2165 gnd 0.007201f
C2813 vdd.n2166 gnd 0.007201f
C2814 vdd.n2167 gnd 0.007201f
C2815 vdd.n2168 gnd 0.008947f
C2816 vdd.n2170 gnd 0.008947f
C2817 vdd.n2171 gnd 0.008947f
C2818 vdd.n2172 gnd 0.007201f
C2819 vdd.n2173 gnd 0.007201f
C2820 vdd.n2174 gnd 0.007201f
C2821 vdd.n2175 gnd 0.008947f
C2822 vdd.n2177 gnd 0.008947f
C2823 vdd.n2178 gnd 0.007201f
C2824 vdd.n2179 gnd 0.007201f
C2825 vdd.n2180 gnd 0.008947f
C2826 vdd.n2182 gnd 0.008947f
C2827 vdd.n2183 gnd 0.008947f
C2828 vdd.n2184 gnd 0.007201f
C2829 vdd.n2185 gnd 0.007694f
C2830 vdd.n2186 gnd 0.949782f
C2831 vdd.n2187 gnd 0.040983f
C2832 vdd.n2188 gnd 0.006084f
C2833 vdd.n2189 gnd 0.006084f
C2834 vdd.n2190 gnd 0.006084f
C2835 vdd.n2191 gnd 0.006084f
C2836 vdd.n2192 gnd 0.006084f
C2837 vdd.n2193 gnd 0.006084f
C2838 vdd.n2194 gnd 0.006084f
C2839 vdd.n2195 gnd 0.006084f
C2840 vdd.n2196 gnd 0.006084f
C2841 vdd.n2197 gnd 0.006084f
C2842 vdd.n2198 gnd 0.006084f
C2843 vdd.n2199 gnd 0.006084f
C2844 vdd.n2200 gnd 0.006084f
C2845 vdd.n2201 gnd 0.006084f
C2846 vdd.n2202 gnd 0.006084f
C2847 vdd.n2203 gnd 0.006084f
C2848 vdd.n2204 gnd 0.006084f
C2849 vdd.n2205 gnd 0.006084f
C2850 vdd.n2206 gnd 0.006084f
C2851 vdd.n2207 gnd 0.006084f
C2852 vdd.n2208 gnd 0.006084f
C2853 vdd.n2209 gnd 0.006084f
C2854 vdd.n2210 gnd 0.006084f
C2855 vdd.n2211 gnd 0.006084f
C2856 vdd.n2212 gnd 0.006084f
C2857 vdd.n2213 gnd 0.006084f
C2858 vdd.n2214 gnd 0.006084f
C2859 vdd.n2215 gnd 0.006084f
C2860 vdd.n2216 gnd 0.006084f
C2861 vdd.n2217 gnd 0.006084f
C2862 vdd.n2218 gnd 10.797999f
C2863 vdd.n2220 gnd 0.013814f
C2864 vdd.n2221 gnd 0.013814f
C2865 vdd.n2222 gnd 0.013026f
C2866 vdd.n2223 gnd 0.006084f
C2867 vdd.n2224 gnd 0.006084f
C2868 vdd.n2225 gnd 0.62173f
C2869 vdd.n2226 gnd 0.006084f
C2870 vdd.n2227 gnd 0.006084f
C2871 vdd.n2228 gnd 0.006084f
C2872 vdd.n2229 gnd 0.006084f
C2873 vdd.n2230 gnd 0.006084f
C2874 vdd.n2231 gnd 0.489155f
C2875 vdd.n2232 gnd 0.006084f
C2876 vdd.n2233 gnd 0.006084f
C2877 vdd.n2234 gnd 0.006084f
C2878 vdd.n2235 gnd 0.006084f
C2879 vdd.n2236 gnd 0.006084f
C2880 vdd.n2237 gnd 0.62173f
C2881 vdd.n2238 gnd 0.006084f
C2882 vdd.n2239 gnd 0.006084f
C2883 vdd.n2240 gnd 0.006084f
C2884 vdd.n2241 gnd 0.006084f
C2885 vdd.n2242 gnd 0.006084f
C2886 vdd.n2243 gnd 0.62173f
C2887 vdd.n2244 gnd 0.006084f
C2888 vdd.n2245 gnd 0.006084f
C2889 vdd.n2246 gnd 0.006084f
C2890 vdd.n2247 gnd 0.006084f
C2891 vdd.n2248 gnd 0.006084f
C2892 vdd.n2249 gnd 0.598872f
C2893 vdd.n2250 gnd 0.006084f
C2894 vdd.n2251 gnd 0.006084f
C2895 vdd.n2252 gnd 0.006084f
C2896 vdd.n2253 gnd 0.006084f
C2897 vdd.n2254 gnd 0.006084f
C2898 vdd.n2255 gnd 0.461726f
C2899 vdd.n2256 gnd 0.006084f
C2900 vdd.n2257 gnd 0.006084f
C2901 vdd.n2258 gnd 0.006084f
C2902 vdd.n2259 gnd 0.006084f
C2903 vdd.n2260 gnd 0.006084f
C2904 vdd.n2261 gnd 0.32458f
C2905 vdd.n2262 gnd 0.006084f
C2906 vdd.n2263 gnd 0.006084f
C2907 vdd.n2264 gnd 0.006084f
C2908 vdd.n2265 gnd 0.006084f
C2909 vdd.n2266 gnd 0.006084f
C2910 vdd.n2267 gnd 0.434297f
C2911 vdd.n2268 gnd 0.006084f
C2912 vdd.n2269 gnd 0.006084f
C2913 vdd.n2270 gnd 0.006084f
C2914 vdd.n2271 gnd 0.006084f
C2915 vdd.n2272 gnd 0.006084f
C2916 vdd.n2273 gnd 0.571443f
C2917 vdd.n2274 gnd 0.006084f
C2918 vdd.n2275 gnd 0.006084f
C2919 vdd.n2276 gnd 0.006084f
C2920 vdd.n2277 gnd 0.006084f
C2921 vdd.n2278 gnd 0.006084f
C2922 vdd.n2279 gnd 0.62173f
C2923 vdd.n2280 gnd 0.006084f
C2924 vdd.n2281 gnd 0.006084f
C2925 vdd.n2282 gnd 0.006084f
C2926 vdd.n2283 gnd 0.006084f
C2927 vdd.n2284 gnd 0.006084f
C2928 vdd.n2285 gnd 0.534871f
C2929 vdd.n2286 gnd 0.006084f
C2930 vdd.n2287 gnd 0.006084f
C2931 vdd.n2288 gnd 0.004831f
C2932 vdd.n2289 gnd 0.017624f
C2933 vdd.n2290 gnd 0.004294f
C2934 vdd.n2291 gnd 0.006084f
C2935 vdd.n2292 gnd 0.397724f
C2936 vdd.n2293 gnd 0.006084f
C2937 vdd.n2294 gnd 0.006084f
C2938 vdd.n2295 gnd 0.006084f
C2939 vdd.n2296 gnd 0.006084f
C2940 vdd.n2297 gnd 0.006084f
C2941 vdd.n2298 gnd 0.361152f
C2942 vdd.n2299 gnd 0.006084f
C2943 vdd.n2300 gnd 0.006084f
C2944 vdd.n2301 gnd 0.006084f
C2945 vdd.n2302 gnd 0.006084f
C2946 vdd.n2303 gnd 0.006084f
C2947 vdd.n2304 gnd 0.498298f
C2948 vdd.n2305 gnd 0.006084f
C2949 vdd.n2306 gnd 0.006084f
C2950 vdd.n2307 gnd 0.006084f
C2951 vdd.n2308 gnd 0.006084f
C2952 vdd.n2309 gnd 0.006084f
C2953 vdd.n2310 gnd 0.548585f
C2954 vdd.n2311 gnd 0.006084f
C2955 vdd.n2312 gnd 0.006084f
C2956 vdd.n2313 gnd 0.006084f
C2957 vdd.n2314 gnd 0.006084f
C2958 vdd.n2315 gnd 0.006084f
C2959 vdd.n2316 gnd 0.411439f
C2960 vdd.n2317 gnd 0.006084f
C2961 vdd.n2318 gnd 0.006084f
C2962 vdd.n2319 gnd 0.006084f
C2963 vdd.n2320 gnd 0.006084f
C2964 vdd.n2321 gnd 0.006084f
C2965 vdd.n2322 gnd 0.196576f
C2966 vdd.n2323 gnd 0.006084f
C2967 vdd.n2324 gnd 0.006084f
C2968 vdd.n2325 gnd 0.006084f
C2969 vdd.n2326 gnd 0.006084f
C2970 vdd.n2327 gnd 0.006084f
C2971 vdd.n2328 gnd 0.196576f
C2972 vdd.n2329 gnd 0.006084f
C2973 vdd.n2330 gnd 0.006084f
C2974 vdd.n2331 gnd 0.006084f
C2975 vdd.n2332 gnd 0.006084f
C2976 vdd.n2333 gnd 0.006084f
C2977 vdd.n2334 gnd 0.62173f
C2978 vdd.n2335 gnd 0.006084f
C2979 vdd.n2336 gnd 0.006084f
C2980 vdd.n2337 gnd 0.006084f
C2981 vdd.n2338 gnd 0.006084f
C2982 vdd.n2339 gnd 0.006084f
C2983 vdd.n2340 gnd 0.006084f
C2984 vdd.n2341 gnd 0.006084f
C2985 vdd.n2342 gnd 0.429725f
C2986 vdd.n2343 gnd 0.006084f
C2987 vdd.n2344 gnd 0.006084f
C2988 vdd.n2345 gnd 0.006084f
C2989 vdd.n2346 gnd 0.006084f
C2990 vdd.n2347 gnd 0.006084f
C2991 vdd.n2348 gnd 0.006084f
C2992 vdd.n2349 gnd 0.388581f
C2993 vdd.n2350 gnd 0.006084f
C2994 vdd.n2351 gnd 0.006084f
C2995 vdd.n2352 gnd 0.006084f
C2996 vdd.n2353 gnd 0.013814f
C2997 vdd.n2354 gnd 0.013026f
C2998 vdd.n2355 gnd 0.006084f
C2999 vdd.n2356 gnd 0.006084f
C3000 vdd.n2357 gnd 0.004697f
C3001 vdd.n2358 gnd 0.006084f
C3002 vdd.n2359 gnd 0.006084f
C3003 vdd.n2360 gnd 0.004429f
C3004 vdd.n2361 gnd 0.006084f
C3005 vdd.n2362 gnd 0.006084f
C3006 vdd.n2363 gnd 0.006084f
C3007 vdd.n2364 gnd 0.006084f
C3008 vdd.n2365 gnd 0.006084f
C3009 vdd.n2366 gnd 0.006084f
C3010 vdd.n2367 gnd 0.006084f
C3011 vdd.n2368 gnd 0.006084f
C3012 vdd.n2369 gnd 0.006084f
C3013 vdd.n2370 gnd 0.006084f
C3014 vdd.n2371 gnd 0.006084f
C3015 vdd.n2372 gnd 0.006084f
C3016 vdd.n2373 gnd 0.006084f
C3017 vdd.n2374 gnd 0.006084f
C3018 vdd.n2375 gnd 0.006084f
C3019 vdd.n2376 gnd 0.006084f
C3020 vdd.n2377 gnd 0.006084f
C3021 vdd.n2378 gnd 0.006084f
C3022 vdd.n2379 gnd 0.006084f
C3023 vdd.n2380 gnd 0.006084f
C3024 vdd.n2381 gnd 0.006084f
C3025 vdd.n2382 gnd 0.006084f
C3026 vdd.n2383 gnd 0.006084f
C3027 vdd.n2384 gnd 0.006084f
C3028 vdd.n2385 gnd 0.006084f
C3029 vdd.n2386 gnd 0.006084f
C3030 vdd.n2387 gnd 0.006084f
C3031 vdd.n2388 gnd 0.006084f
C3032 vdd.n2389 gnd 0.006084f
C3033 vdd.n2390 gnd 0.006084f
C3034 vdd.n2391 gnd 0.006084f
C3035 vdd.n2392 gnd 0.006084f
C3036 vdd.n2393 gnd 0.006084f
C3037 vdd.n2394 gnd 0.006084f
C3038 vdd.n2395 gnd 0.006084f
C3039 vdd.n2396 gnd 0.006084f
C3040 vdd.n2397 gnd 0.006084f
C3041 vdd.n2398 gnd 0.006084f
C3042 vdd.n2399 gnd 0.006084f
C3043 vdd.n2400 gnd 0.006084f
C3044 vdd.n2401 gnd 0.006084f
C3045 vdd.n2402 gnd 0.006084f
C3046 vdd.n2403 gnd 0.006084f
C3047 vdd.n2404 gnd 0.006084f
C3048 vdd.n2405 gnd 0.006084f
C3049 vdd.n2406 gnd 0.006084f
C3050 vdd.n2407 gnd 0.006084f
C3051 vdd.n2408 gnd 0.006084f
C3052 vdd.n2409 gnd 0.006084f
C3053 vdd.n2410 gnd 0.006084f
C3054 vdd.n2411 gnd 0.006084f
C3055 vdd.n2412 gnd 0.006084f
C3056 vdd.n2413 gnd 0.006084f
C3057 vdd.n2414 gnd 0.006084f
C3058 vdd.n2415 gnd 0.006084f
C3059 vdd.n2416 gnd 0.006084f
C3060 vdd.n2417 gnd 0.006084f
C3061 vdd.n2418 gnd 0.006084f
C3062 vdd.n2419 gnd 0.006084f
C3063 vdd.n2420 gnd 0.006084f
C3064 vdd.n2421 gnd 0.013814f
C3065 vdd.n2422 gnd 0.013026f
C3066 vdd.n2423 gnd 0.013026f
C3067 vdd.n2424 gnd 0.704018f
C3068 vdd.n2425 gnd 0.013026f
C3069 vdd.n2426 gnd 0.013814f
C3070 vdd.n2427 gnd 0.013026f
C3071 vdd.n2428 gnd 0.006084f
C3072 vdd.n2429 gnd 0.006084f
C3073 vdd.n2430 gnd 0.006084f
C3074 vdd.n2431 gnd 0.004697f
C3075 vdd.n2432 gnd 0.008695f
C3076 vdd.n2433 gnd 0.004429f
C3077 vdd.n2434 gnd 0.006084f
C3078 vdd.n2435 gnd 0.006084f
C3079 vdd.n2436 gnd 0.006084f
C3080 vdd.n2437 gnd 0.006084f
C3081 vdd.n2438 gnd 0.006084f
C3082 vdd.n2439 gnd 0.006084f
C3083 vdd.n2440 gnd 0.006084f
C3084 vdd.n2441 gnd 0.006084f
C3085 vdd.n2442 gnd 0.006084f
C3086 vdd.n2443 gnd 0.006084f
C3087 vdd.n2444 gnd 0.006084f
C3088 vdd.n2445 gnd 0.006084f
C3089 vdd.n2446 gnd 0.006084f
C3090 vdd.n2447 gnd 0.006084f
C3091 vdd.n2448 gnd 0.006084f
C3092 vdd.n2449 gnd 0.006084f
C3093 vdd.n2450 gnd 0.006084f
C3094 vdd.n2451 gnd 0.006084f
C3095 vdd.n2452 gnd 0.006084f
C3096 vdd.n2453 gnd 0.006084f
C3097 vdd.n2454 gnd 0.006084f
C3098 vdd.n2455 gnd 0.006084f
C3099 vdd.n2456 gnd 0.006084f
C3100 vdd.n2457 gnd 0.006084f
C3101 vdd.n2458 gnd 0.006084f
C3102 vdd.n2459 gnd 0.006084f
C3103 vdd.n2460 gnd 0.006084f
C3104 vdd.n2461 gnd 0.006084f
C3105 vdd.n2462 gnd 0.006084f
C3106 vdd.n2463 gnd 0.006084f
C3107 vdd.n2464 gnd 0.006084f
C3108 vdd.n2465 gnd 0.006084f
C3109 vdd.n2466 gnd 0.006084f
C3110 vdd.n2467 gnd 0.006084f
C3111 vdd.n2468 gnd 0.006084f
C3112 vdd.n2469 gnd 0.006084f
C3113 vdd.n2470 gnd 0.006084f
C3114 vdd.n2471 gnd 0.006084f
C3115 vdd.n2472 gnd 0.006084f
C3116 vdd.n2473 gnd 0.006084f
C3117 vdd.n2474 gnd 0.006084f
C3118 vdd.n2475 gnd 0.006084f
C3119 vdd.n2476 gnd 0.006084f
C3120 vdd.n2477 gnd 0.006084f
C3121 vdd.n2478 gnd 0.006084f
C3122 vdd.n2479 gnd 0.006084f
C3123 vdd.n2480 gnd 0.006084f
C3124 vdd.n2481 gnd 0.006084f
C3125 vdd.n2482 gnd 0.006084f
C3126 vdd.n2483 gnd 0.006084f
C3127 vdd.n2484 gnd 0.006084f
C3128 vdd.n2485 gnd 0.006084f
C3129 vdd.n2486 gnd 0.006084f
C3130 vdd.n2487 gnd 0.006084f
C3131 vdd.n2488 gnd 0.006084f
C3132 vdd.n2489 gnd 0.006084f
C3133 vdd.n2490 gnd 0.006084f
C3134 vdd.n2491 gnd 0.006084f
C3135 vdd.n2492 gnd 0.006084f
C3136 vdd.n2493 gnd 0.006084f
C3137 vdd.n2494 gnd 0.013814f
C3138 vdd.n2495 gnd 0.013814f
C3139 vdd.n2496 gnd 0.758876f
C3140 vdd.t104 gnd 2.69721f
C3141 vdd.t91 gnd 2.69721f
C3142 vdd.n2530 gnd 0.013814f
C3143 vdd.t109 gnd 0.530299f
C3144 vdd.n2531 gnd 0.006084f
C3145 vdd.t58 gnd 0.245843f
C3146 vdd.t59 gnd 0.251651f
C3147 vdd.t56 gnd 0.160496f
C3148 vdd.n2532 gnd 0.086739f
C3149 vdd.n2533 gnd 0.049201f
C3150 vdd.n2534 gnd 0.006084f
C3151 vdd.t68 gnd 0.245843f
C3152 vdd.t69 gnd 0.251651f
C3153 vdd.t67 gnd 0.160496f
C3154 vdd.n2535 gnd 0.086739f
C3155 vdd.n2536 gnd 0.049201f
C3156 vdd.n2537 gnd 0.008695f
C3157 vdd.n2538 gnd 0.013814f
C3158 vdd.n2539 gnd 0.013814f
C3159 vdd.n2540 gnd 0.006084f
C3160 vdd.n2541 gnd 0.006084f
C3161 vdd.n2542 gnd 0.006084f
C3162 vdd.n2543 gnd 0.006084f
C3163 vdd.n2544 gnd 0.006084f
C3164 vdd.n2545 gnd 0.006084f
C3165 vdd.n2546 gnd 0.006084f
C3166 vdd.n2547 gnd 0.006084f
C3167 vdd.n2548 gnd 0.006084f
C3168 vdd.n2549 gnd 0.006084f
C3169 vdd.n2550 gnd 0.006084f
C3170 vdd.n2551 gnd 0.006084f
C3171 vdd.n2552 gnd 0.006084f
C3172 vdd.n2553 gnd 0.006084f
C3173 vdd.n2554 gnd 0.006084f
C3174 vdd.n2555 gnd 0.006084f
C3175 vdd.n2556 gnd 0.006084f
C3176 vdd.n2557 gnd 0.006084f
C3177 vdd.n2558 gnd 0.006084f
C3178 vdd.n2559 gnd 0.006084f
C3179 vdd.n2560 gnd 0.006084f
C3180 vdd.n2561 gnd 0.006084f
C3181 vdd.n2562 gnd 0.006084f
C3182 vdd.n2563 gnd 0.006084f
C3183 vdd.n2564 gnd 0.006084f
C3184 vdd.n2565 gnd 0.006084f
C3185 vdd.n2566 gnd 0.006084f
C3186 vdd.n2567 gnd 0.006084f
C3187 vdd.n2568 gnd 0.006084f
C3188 vdd.n2569 gnd 0.006084f
C3189 vdd.n2570 gnd 0.006084f
C3190 vdd.n2571 gnd 0.006084f
C3191 vdd.n2572 gnd 0.006084f
C3192 vdd.n2573 gnd 0.006084f
C3193 vdd.n2574 gnd 0.006084f
C3194 vdd.n2575 gnd 0.006084f
C3195 vdd.n2576 gnd 0.006084f
C3196 vdd.n2577 gnd 0.006084f
C3197 vdd.n2578 gnd 0.006084f
C3198 vdd.n2579 gnd 0.006084f
C3199 vdd.n2580 gnd 0.006084f
C3200 vdd.n2581 gnd 0.006084f
C3201 vdd.n2582 gnd 0.006084f
C3202 vdd.n2583 gnd 0.006084f
C3203 vdd.n2584 gnd 0.006084f
C3204 vdd.n2585 gnd 0.006084f
C3205 vdd.n2586 gnd 0.006084f
C3206 vdd.n2587 gnd 0.006084f
C3207 vdd.n2588 gnd 0.006084f
C3208 vdd.n2589 gnd 0.006084f
C3209 vdd.n2590 gnd 0.006084f
C3210 vdd.n2591 gnd 0.006084f
C3211 vdd.n2592 gnd 0.006084f
C3212 vdd.n2593 gnd 0.006084f
C3213 vdd.n2594 gnd 0.006084f
C3214 vdd.n2595 gnd 0.006084f
C3215 vdd.n2596 gnd 0.006084f
C3216 vdd.n2597 gnd 0.006084f
C3217 vdd.n2598 gnd 0.006084f
C3218 vdd.n2599 gnd 0.006084f
C3219 vdd.n2600 gnd 0.004429f
C3220 vdd.n2601 gnd 0.006084f
C3221 vdd.n2602 gnd 0.006084f
C3222 vdd.n2603 gnd 0.004697f
C3223 vdd.n2604 gnd 0.006084f
C3224 vdd.n2605 gnd 0.006084f
C3225 vdd.n2606 gnd 0.013814f
C3226 vdd.n2607 gnd 0.013026f
C3227 vdd.n2608 gnd 0.013026f
C3228 vdd.n2609 gnd 0.006084f
C3229 vdd.n2610 gnd 0.006084f
C3230 vdd.n2611 gnd 0.006084f
C3231 vdd.n2612 gnd 0.006084f
C3232 vdd.n2613 gnd 0.006084f
C3233 vdd.n2614 gnd 0.006084f
C3234 vdd.n2615 gnd 0.006084f
C3235 vdd.n2616 gnd 0.006084f
C3236 vdd.n2617 gnd 0.006084f
C3237 vdd.n2618 gnd 0.006084f
C3238 vdd.n2619 gnd 0.006084f
C3239 vdd.n2620 gnd 0.006084f
C3240 vdd.n2621 gnd 0.006084f
C3241 vdd.n2622 gnd 0.006084f
C3242 vdd.n2623 gnd 0.006084f
C3243 vdd.n2624 gnd 0.006084f
C3244 vdd.n2625 gnd 0.006084f
C3245 vdd.n2626 gnd 0.006084f
C3246 vdd.n2627 gnd 0.006084f
C3247 vdd.n2628 gnd 0.006084f
C3248 vdd.n2629 gnd 0.006084f
C3249 vdd.n2630 gnd 0.006084f
C3250 vdd.n2631 gnd 0.006084f
C3251 vdd.n2632 gnd 0.006084f
C3252 vdd.n2633 gnd 0.006084f
C3253 vdd.n2634 gnd 0.006084f
C3254 vdd.n2635 gnd 0.006084f
C3255 vdd.n2636 gnd 0.006084f
C3256 vdd.n2637 gnd 0.006084f
C3257 vdd.n2638 gnd 0.006084f
C3258 vdd.n2639 gnd 0.006084f
C3259 vdd.n2640 gnd 0.006084f
C3260 vdd.n2641 gnd 0.006084f
C3261 vdd.n2642 gnd 0.006084f
C3262 vdd.n2643 gnd 0.006084f
C3263 vdd.n2644 gnd 0.006084f
C3264 vdd.n2645 gnd 0.006084f
C3265 vdd.n2646 gnd 0.006084f
C3266 vdd.n2647 gnd 0.006084f
C3267 vdd.n2648 gnd 0.006084f
C3268 vdd.n2649 gnd 0.006084f
C3269 vdd.n2650 gnd 0.006084f
C3270 vdd.n2651 gnd 0.006084f
C3271 vdd.n2652 gnd 0.006084f
C3272 vdd.n2653 gnd 0.006084f
C3273 vdd.n2654 gnd 0.006084f
C3274 vdd.n2655 gnd 0.006084f
C3275 vdd.n2656 gnd 0.006084f
C3276 vdd.n2657 gnd 0.006084f
C3277 vdd.n2658 gnd 0.006084f
C3278 vdd.n2659 gnd 0.006084f
C3279 vdd.n2660 gnd 0.006084f
C3280 vdd.n2661 gnd 0.006084f
C3281 vdd.n2662 gnd 0.006084f
C3282 vdd.n2663 gnd 0.006084f
C3283 vdd.n2664 gnd 0.006084f
C3284 vdd.n2665 gnd 0.006084f
C3285 vdd.n2666 gnd 0.006084f
C3286 vdd.n2667 gnd 0.006084f
C3287 vdd.n2668 gnd 0.006084f
C3288 vdd.n2669 gnd 0.006084f
C3289 vdd.n2670 gnd 0.006084f
C3290 vdd.n2671 gnd 0.006084f
C3291 vdd.n2672 gnd 0.006084f
C3292 vdd.n2673 gnd 0.006084f
C3293 vdd.n2674 gnd 0.006084f
C3294 vdd.n2675 gnd 0.006084f
C3295 vdd.n2676 gnd 0.006084f
C3296 vdd.n2677 gnd 0.006084f
C3297 vdd.n2678 gnd 0.006084f
C3298 vdd.n2679 gnd 0.006084f
C3299 vdd.n2680 gnd 0.006084f
C3300 vdd.n2681 gnd 0.006084f
C3301 vdd.n2682 gnd 0.006084f
C3302 vdd.n2683 gnd 0.006084f
C3303 vdd.n2684 gnd 0.006084f
C3304 vdd.n2685 gnd 0.006084f
C3305 vdd.n2686 gnd 0.006084f
C3306 vdd.n2687 gnd 0.006084f
C3307 vdd.n2688 gnd 0.006084f
C3308 vdd.n2689 gnd 0.006084f
C3309 vdd.n2690 gnd 0.006084f
C3310 vdd.n2691 gnd 0.006084f
C3311 vdd.n2692 gnd 0.006084f
C3312 vdd.n2693 gnd 0.006084f
C3313 vdd.n2694 gnd 0.006084f
C3314 vdd.n2695 gnd 0.006084f
C3315 vdd.n2696 gnd 0.006084f
C3316 vdd.n2697 gnd 0.006084f
C3317 vdd.n2698 gnd 0.006084f
C3318 vdd.n2699 gnd 0.006084f
C3319 vdd.n2700 gnd 0.006084f
C3320 vdd.n2701 gnd 0.006084f
C3321 vdd.n2702 gnd 0.006084f
C3322 vdd.n2703 gnd 0.006084f
C3323 vdd.n2704 gnd 0.006084f
C3324 vdd.n2705 gnd 0.006084f
C3325 vdd.n2706 gnd 0.006084f
C3326 vdd.n2707 gnd 0.006084f
C3327 vdd.n2708 gnd 0.006084f
C3328 vdd.n2709 gnd 0.006084f
C3329 vdd.n2710 gnd 0.196576f
C3330 vdd.n2711 gnd 0.006084f
C3331 vdd.n2712 gnd 0.006084f
C3332 vdd.n2713 gnd 0.006084f
C3333 vdd.n2714 gnd 0.006084f
C3334 vdd.n2715 gnd 0.006084f
C3335 vdd.n2716 gnd 0.196576f
C3336 vdd.n2717 gnd 0.006084f
C3337 vdd.n2718 gnd 0.006084f
C3338 vdd.n2719 gnd 0.006084f
C3339 vdd.n2720 gnd 0.006084f
C3340 vdd.n2721 gnd 0.006084f
C3341 vdd.n2722 gnd 0.006084f
C3342 vdd.n2723 gnd 0.006084f
C3343 vdd.n2724 gnd 0.006084f
C3344 vdd.n2725 gnd 0.006084f
C3345 vdd.n2726 gnd 0.006084f
C3346 vdd.n2727 gnd 0.006084f
C3347 vdd.n2728 gnd 0.388581f
C3348 vdd.n2729 gnd 0.006084f
C3349 vdd.n2730 gnd 0.006084f
C3350 vdd.n2731 gnd 0.006084f
C3351 vdd.n2732 gnd 0.013026f
C3352 vdd.n2733 gnd 0.013026f
C3353 vdd.n2734 gnd 0.013814f
C3354 vdd.n2735 gnd 0.013814f
C3355 vdd.n2736 gnd 0.006084f
C3356 vdd.n2737 gnd 0.006084f
C3357 vdd.n2738 gnd 0.006084f
C3358 vdd.n2739 gnd 0.004697f
C3359 vdd.n2740 gnd 0.008695f
C3360 vdd.n2741 gnd 0.004429f
C3361 vdd.n2742 gnd 0.006084f
C3362 vdd.n2743 gnd 0.006084f
C3363 vdd.n2744 gnd 0.006084f
C3364 vdd.n2745 gnd 0.006084f
C3365 vdd.n2746 gnd 0.006084f
C3366 vdd.n2747 gnd 0.006084f
C3367 vdd.n2748 gnd 0.006084f
C3368 vdd.n2749 gnd 0.006084f
C3369 vdd.n2750 gnd 0.006084f
C3370 vdd.n2751 gnd 0.006084f
C3371 vdd.n2752 gnd 0.006084f
C3372 vdd.n2753 gnd 0.006084f
C3373 vdd.n2754 gnd 0.006084f
C3374 vdd.n2755 gnd 0.006084f
C3375 vdd.n2756 gnd 0.006084f
C3376 vdd.n2757 gnd 0.006084f
C3377 vdd.n2758 gnd 0.006084f
C3378 vdd.n2759 gnd 0.006084f
C3379 vdd.n2760 gnd 0.006084f
C3380 vdd.n2761 gnd 0.006084f
C3381 vdd.n2762 gnd 0.006084f
C3382 vdd.n2763 gnd 0.006084f
C3383 vdd.n2764 gnd 0.006084f
C3384 vdd.n2765 gnd 0.006084f
C3385 vdd.n2766 gnd 0.006084f
C3386 vdd.n2767 gnd 0.006084f
C3387 vdd.n2768 gnd 0.006084f
C3388 vdd.n2769 gnd 0.006084f
C3389 vdd.n2770 gnd 0.006084f
C3390 vdd.n2771 gnd 0.006084f
C3391 vdd.n2772 gnd 0.006084f
C3392 vdd.n2773 gnd 0.006084f
C3393 vdd.n2774 gnd 0.006084f
C3394 vdd.n2775 gnd 0.006084f
C3395 vdd.n2776 gnd 0.006084f
C3396 vdd.n2777 gnd 0.006084f
C3397 vdd.n2778 gnd 0.006084f
C3398 vdd.n2779 gnd 0.006084f
C3399 vdd.n2780 gnd 0.006084f
C3400 vdd.n2781 gnd 0.006084f
C3401 vdd.n2782 gnd 0.006084f
C3402 vdd.n2783 gnd 0.006084f
C3403 vdd.n2784 gnd 0.006084f
C3404 vdd.n2785 gnd 0.006084f
C3405 vdd.n2786 gnd 0.006084f
C3406 vdd.n2787 gnd 0.006084f
C3407 vdd.n2788 gnd 0.006084f
C3408 vdd.n2789 gnd 0.006084f
C3409 vdd.n2790 gnd 0.006084f
C3410 vdd.n2791 gnd 0.006084f
C3411 vdd.n2792 gnd 0.006084f
C3412 vdd.n2793 gnd 0.006084f
C3413 vdd.n2794 gnd 0.006084f
C3414 vdd.n2795 gnd 0.006084f
C3415 vdd.n2796 gnd 0.006084f
C3416 vdd.n2797 gnd 0.006084f
C3417 vdd.n2798 gnd 0.006084f
C3418 vdd.n2799 gnd 0.006084f
C3419 vdd.n2800 gnd 0.758876f
C3420 vdd.n2802 gnd 0.013814f
C3421 vdd.n2803 gnd 0.013814f
C3422 vdd.n2804 gnd 0.013026f
C3423 vdd.n2805 gnd 0.006084f
C3424 vdd.n2806 gnd 0.006084f
C3425 vdd.n2807 gnd 0.365723f
C3426 vdd.n2808 gnd 0.006084f
C3427 vdd.n2809 gnd 0.006084f
C3428 vdd.n2810 gnd 0.006084f
C3429 vdd.n2811 gnd 0.006084f
C3430 vdd.n2812 gnd 0.006084f
C3431 vdd.n2813 gnd 0.370295f
C3432 vdd.n2814 gnd 0.006084f
C3433 vdd.n2815 gnd 0.006084f
C3434 vdd.n2816 gnd 0.006084f
C3435 vdd.n2817 gnd 0.006084f
C3436 vdd.n2818 gnd 0.006084f
C3437 vdd.n2819 gnd 0.62173f
C3438 vdd.n2820 gnd 0.006084f
C3439 vdd.n2821 gnd 0.006084f
C3440 vdd.n2822 gnd 0.006084f
C3441 vdd.n2823 gnd 0.006084f
C3442 vdd.n2824 gnd 0.006084f
C3443 vdd.n2825 gnd 0.448011f
C3444 vdd.n2826 gnd 0.006084f
C3445 vdd.n2827 gnd 0.006084f
C3446 vdd.n2828 gnd 0.006084f
C3447 vdd.n2829 gnd 0.006084f
C3448 vdd.n2830 gnd 0.006084f
C3449 vdd.n2831 gnd 0.5623f
C3450 vdd.n2832 gnd 0.006084f
C3451 vdd.n2833 gnd 0.006084f
C3452 vdd.n2834 gnd 0.006084f
C3453 vdd.n2835 gnd 0.006084f
C3454 vdd.n2836 gnd 0.006084f
C3455 vdd.n2837 gnd 0.461726f
C3456 vdd.n2838 gnd 0.006084f
C3457 vdd.n2839 gnd 0.006084f
C3458 vdd.n2840 gnd 0.006084f
C3459 vdd.n2841 gnd 0.006084f
C3460 vdd.n2842 gnd 0.006084f
C3461 vdd.n2843 gnd 0.32458f
C3462 vdd.n2844 gnd 0.006084f
C3463 vdd.n2845 gnd 0.006084f
C3464 vdd.n2846 gnd 0.006084f
C3465 vdd.n2847 gnd 0.006084f
C3466 vdd.n2848 gnd 0.006084f
C3467 vdd.n2849 gnd 0.196576f
C3468 vdd.n2850 gnd 0.006084f
C3469 vdd.n2851 gnd 0.006084f
C3470 vdd.n2852 gnd 0.006084f
C3471 vdd.n2853 gnd 0.006084f
C3472 vdd.n2854 gnd 0.006084f
C3473 vdd.n2855 gnd 0.571443f
C3474 vdd.n2856 gnd 0.006084f
C3475 vdd.n2857 gnd 0.006084f
C3476 vdd.n2858 gnd 0.006084f
C3477 vdd.n2859 gnd 0.004294f
C3478 vdd.n2860 gnd 0.006084f
C3479 vdd.n2861 gnd 0.006084f
C3480 vdd.n2862 gnd 0.62173f
C3481 vdd.n2863 gnd 0.006084f
C3482 vdd.n2864 gnd 0.006084f
C3483 vdd.n2865 gnd 0.006084f
C3484 vdd.n2866 gnd 0.006084f
C3485 vdd.n2867 gnd 0.006084f
C3486 vdd.n2868 gnd 0.493727f
C3487 vdd.n2869 gnd 0.006084f
C3488 vdd.n2870 gnd 0.004831f
C3489 vdd.n2871 gnd 0.006084f
C3490 vdd.n2872 gnd 0.006084f
C3491 vdd.n2873 gnd 0.006084f
C3492 vdd.n2874 gnd 0.397724f
C3493 vdd.n2875 gnd 0.006084f
C3494 vdd.n2876 gnd 0.006084f
C3495 vdd.n2877 gnd 0.006084f
C3496 vdd.n2878 gnd 0.006084f
C3497 vdd.n2879 gnd 0.006084f
C3498 vdd.n2880 gnd 0.361152f
C3499 vdd.n2881 gnd 0.006084f
C3500 vdd.n2882 gnd 0.006084f
C3501 vdd.n2883 gnd 0.006084f
C3502 vdd.n2884 gnd 0.006084f
C3503 vdd.n2885 gnd 0.006084f
C3504 vdd.n2886 gnd 0.498298f
C3505 vdd.n2887 gnd 0.006084f
C3506 vdd.n2888 gnd 0.006084f
C3507 vdd.n2889 gnd 0.006084f
C3508 vdd.n2890 gnd 0.006084f
C3509 vdd.n2891 gnd 0.006084f
C3510 vdd.n2892 gnd 0.62173f
C3511 vdd.n2893 gnd 0.006084f
C3512 vdd.n2894 gnd 0.006084f
C3513 vdd.n2895 gnd 0.006084f
C3514 vdd.n2896 gnd 0.006084f
C3515 vdd.n2897 gnd 0.006084f
C3516 vdd.n2898 gnd 0.608015f
C3517 vdd.n2899 gnd 0.006084f
C3518 vdd.n2900 gnd 0.006084f
C3519 vdd.n2901 gnd 0.006084f
C3520 vdd.n2902 gnd 0.006084f
C3521 vdd.n2903 gnd 0.006084f
C3522 vdd.n2904 gnd 0.470869f
C3523 vdd.n2905 gnd 0.006084f
C3524 vdd.n2906 gnd 0.006084f
C3525 vdd.n2907 gnd 0.006084f
C3526 vdd.n2908 gnd 0.006084f
C3527 vdd.n2909 gnd 0.006084f
C3528 vdd.n2910 gnd 0.333723f
C3529 vdd.n2911 gnd 0.006084f
C3530 vdd.n2912 gnd 0.006084f
C3531 vdd.n2913 gnd 0.006084f
C3532 vdd.n2914 gnd 0.006084f
C3533 vdd.n2915 gnd 0.006084f
C3534 vdd.n2916 gnd 0.62173f
C3535 vdd.n2917 gnd 0.006084f
C3536 vdd.n2918 gnd 0.006084f
C3537 vdd.n2919 gnd 0.006084f
C3538 vdd.n2920 gnd 0.006084f
C3539 vdd.n2921 gnd 0.006084f
C3540 vdd.n2922 gnd 0.006084f
C3541 vdd.n2924 gnd 0.006084f
C3542 vdd.n2925 gnd 0.006084f
C3543 vdd.n2927 gnd 0.006084f
C3544 vdd.n2928 gnd 0.006084f
C3545 vdd.n2931 gnd 0.006084f
C3546 vdd.n2932 gnd 0.006084f
C3547 vdd.n2933 gnd 0.006084f
C3548 vdd.n2934 gnd 0.006084f
C3549 vdd.n2936 gnd 0.006084f
C3550 vdd.n2937 gnd 0.006084f
C3551 vdd.n2938 gnd 0.006084f
C3552 vdd.n2939 gnd 0.006084f
C3553 vdd.n2940 gnd 0.006084f
C3554 vdd.n2941 gnd 0.006084f
C3555 vdd.n2943 gnd 0.006084f
C3556 vdd.n2944 gnd 0.006084f
C3557 vdd.n2945 gnd 0.006084f
C3558 vdd.n2946 gnd 0.006084f
C3559 vdd.n2947 gnd 0.006084f
C3560 vdd.n2948 gnd 0.006084f
C3561 vdd.n2950 gnd 0.006084f
C3562 vdd.n2951 gnd 0.006084f
C3563 vdd.n2952 gnd 0.006084f
C3564 vdd.n2953 gnd 0.006084f
C3565 vdd.n2954 gnd 0.006084f
C3566 vdd.n2955 gnd 0.006084f
C3567 vdd.n2957 gnd 0.006084f
C3568 vdd.n2958 gnd 0.013814f
C3569 vdd.n2959 gnd 0.013814f
C3570 vdd.n2960 gnd 0.013026f
C3571 vdd.n2961 gnd 0.006084f
C3572 vdd.n2962 gnd 0.006084f
C3573 vdd.n2963 gnd 0.006084f
C3574 vdd.n2964 gnd 0.006084f
C3575 vdd.n2965 gnd 0.006084f
C3576 vdd.n2966 gnd 0.006084f
C3577 vdd.n2967 gnd 0.62173f
C3578 vdd.n2968 gnd 0.006084f
C3579 vdd.n2969 gnd 0.006084f
C3580 vdd.n2970 gnd 0.006084f
C3581 vdd.n2971 gnd 0.006084f
C3582 vdd.n2972 gnd 0.006084f
C3583 vdd.n2973 gnd 0.44344f
C3584 vdd.n2974 gnd 0.006084f
C3585 vdd.n2975 gnd 0.006084f
C3586 vdd.n2976 gnd 0.006084f
C3587 vdd.n2977 gnd 0.013814f
C3588 vdd.n2979 gnd 0.013814f
C3589 vdd.n2980 gnd 0.013026f
C3590 vdd.n2981 gnd 0.006084f
C3591 vdd.n2982 gnd 0.004697f
C3592 vdd.n2983 gnd 0.006084f
C3593 vdd.n2985 gnd 0.006084f
C3594 vdd.n2986 gnd 0.006084f
C3595 vdd.n2987 gnd 0.006084f
C3596 vdd.n2988 gnd 0.006084f
C3597 vdd.n2989 gnd 0.006084f
C3598 vdd.n2990 gnd 0.006084f
C3599 vdd.n2992 gnd 0.006084f
C3600 vdd.n2993 gnd 0.006084f
C3601 vdd.n2994 gnd 0.006084f
C3602 vdd.n2995 gnd 0.006084f
C3603 vdd.n2996 gnd 0.006084f
C3604 vdd.n2997 gnd 0.006084f
C3605 vdd.n2999 gnd 0.006084f
C3606 vdd.n3000 gnd 0.006084f
C3607 vdd.n3001 gnd 0.006084f
C3608 vdd.n3002 gnd 0.006084f
C3609 vdd.n3003 gnd 0.006084f
C3610 vdd.n3004 gnd 0.006084f
C3611 vdd.n3006 gnd 0.006084f
C3612 vdd.n3007 gnd 0.006084f
C3613 vdd.n3008 gnd 0.006084f
C3614 vdd.n3009 gnd 0.9532f
C3615 vdd.n3010 gnd 0.037566f
C3616 vdd.n3011 gnd 0.006084f
C3617 vdd.n3012 gnd 0.006084f
C3618 vdd.n3014 gnd 0.006084f
C3619 vdd.n3015 gnd 0.006084f
C3620 vdd.n3016 gnd 0.006084f
C3621 vdd.n3017 gnd 0.006084f
C3622 vdd.n3018 gnd 0.006084f
C3623 vdd.n3019 gnd 0.006084f
C3624 vdd.n3021 gnd 0.006084f
C3625 vdd.n3022 gnd 0.006084f
C3626 vdd.n3023 gnd 0.006084f
C3627 vdd.n3024 gnd 0.006084f
C3628 vdd.n3025 gnd 0.006084f
C3629 vdd.n3026 gnd 0.006084f
C3630 vdd.n3028 gnd 0.006084f
C3631 vdd.n3029 gnd 0.006084f
C3632 vdd.n3030 gnd 0.006084f
C3633 vdd.n3031 gnd 0.006084f
C3634 vdd.n3032 gnd 0.006084f
C3635 vdd.n3033 gnd 0.006084f
C3636 vdd.n3035 gnd 0.006084f
C3637 vdd.n3036 gnd 0.006084f
C3638 vdd.n3038 gnd 0.006084f
C3639 vdd.n3039 gnd 0.006084f
C3640 vdd.n3040 gnd 0.013814f
C3641 vdd.n3041 gnd 0.013026f
C3642 vdd.n3042 gnd 0.013026f
C3643 vdd.n3043 gnd 0.841164f
C3644 vdd.n3044 gnd 0.013026f
C3645 vdd.n3045 gnd 0.013814f
C3646 vdd.n3046 gnd 0.013026f
C3647 vdd.n3047 gnd 0.006084f
C3648 vdd.n3048 gnd 0.004697f
C3649 vdd.n3049 gnd 0.006084f
C3650 vdd.n3051 gnd 0.006084f
C3651 vdd.n3052 gnd 0.006084f
C3652 vdd.n3053 gnd 0.006084f
C3653 vdd.n3054 gnd 0.006084f
C3654 vdd.n3055 gnd 0.006084f
C3655 vdd.n3056 gnd 0.006084f
C3656 vdd.n3058 gnd 0.006084f
C3657 vdd.n3059 gnd 0.006084f
C3658 vdd.n3060 gnd 0.006084f
C3659 vdd.n3061 gnd 0.006084f
C3660 vdd.n3062 gnd 0.006084f
C3661 vdd.n3063 gnd 0.006084f
C3662 vdd.n3065 gnd 0.006084f
C3663 vdd.n3066 gnd 0.006084f
C3664 vdd.n3067 gnd 0.006084f
C3665 vdd.n3068 gnd 0.006084f
C3666 vdd.n3069 gnd 0.006084f
C3667 vdd.n3070 gnd 0.006084f
C3668 vdd.n3072 gnd 0.006084f
C3669 vdd.n3073 gnd 0.006084f
C3670 vdd.n3075 gnd 0.006084f
C3671 vdd.n3076 gnd 0.037566f
C3672 vdd.n3077 gnd 0.9532f
C3673 vdd.n3078 gnd 0.007694f
C3674 vdd.n3079 gnd 0.00342f
C3675 vdd.t20 gnd 0.110068f
C3676 vdd.t21 gnd 0.117632f
C3677 vdd.t18 gnd 0.143747f
C3678 vdd.n3080 gnd 0.184263f
C3679 vdd.n3081 gnd 0.154815f
C3680 vdd.n3082 gnd 0.01109f
C3681 vdd.n3083 gnd 0.008947f
C3682 vdd.n3084 gnd 0.003781f
C3683 vdd.n3085 gnd 0.007201f
C3684 vdd.n3086 gnd 0.008947f
C3685 vdd.n3087 gnd 0.008947f
C3686 vdd.n3088 gnd 0.007201f
C3687 vdd.n3089 gnd 0.007201f
C3688 vdd.n3090 gnd 0.008947f
C3689 vdd.n3092 gnd 0.008947f
C3690 vdd.n3093 gnd 0.007201f
C3691 vdd.n3094 gnd 0.007201f
C3692 vdd.n3095 gnd 0.007201f
C3693 vdd.n3096 gnd 0.008947f
C3694 vdd.n3098 gnd 0.008947f
C3695 vdd.n3100 gnd 0.008947f
C3696 vdd.n3101 gnd 0.007201f
C3697 vdd.n3102 gnd 0.007201f
C3698 vdd.n3103 gnd 0.007201f
C3699 vdd.n3104 gnd 0.008947f
C3700 vdd.n3106 gnd 0.008947f
C3701 vdd.n3108 gnd 0.008947f
C3702 vdd.n3109 gnd 0.007201f
C3703 vdd.n3110 gnd 0.007201f
C3704 vdd.n3111 gnd 0.007201f
C3705 vdd.n3112 gnd 0.008947f
C3706 vdd.n3114 gnd 0.008947f
C3707 vdd.n3115 gnd 0.008947f
C3708 vdd.n3116 gnd 0.007201f
C3709 vdd.n3117 gnd 0.007201f
C3710 vdd.n3118 gnd 0.008947f
C3711 vdd.n3119 gnd 0.008947f
C3712 vdd.n3121 gnd 0.008947f
C3713 vdd.n3122 gnd 0.007201f
C3714 vdd.n3123 gnd 0.008947f
C3715 vdd.n3124 gnd 0.008947f
C3716 vdd.n3125 gnd 0.008947f
C3717 vdd.n3126 gnd 0.01469f
C3718 vdd.n3127 gnd 0.004897f
C3719 vdd.n3128 gnd 0.008947f
C3720 vdd.n3130 gnd 0.008947f
C3721 vdd.n3132 gnd 0.008947f
C3722 vdd.n3133 gnd 0.007201f
C3723 vdd.n3134 gnd 0.007201f
C3724 vdd.n3135 gnd 0.007201f
C3725 vdd.n3136 gnd 0.008947f
C3726 vdd.n3138 gnd 0.008947f
C3727 vdd.n3140 gnd 0.008947f
C3728 vdd.n3141 gnd 0.007201f
C3729 vdd.n3142 gnd 0.007201f
C3730 vdd.n3143 gnd 0.007201f
C3731 vdd.n3144 gnd 0.008947f
C3732 vdd.n3146 gnd 0.008947f
C3733 vdd.n3148 gnd 0.008947f
C3734 vdd.n3149 gnd 0.007201f
C3735 vdd.n3150 gnd 0.007201f
C3736 vdd.n3151 gnd 0.007201f
C3737 vdd.n3152 gnd 0.008947f
C3738 vdd.n3154 gnd 0.008947f
C3739 vdd.n3156 gnd 0.008947f
C3740 vdd.n3157 gnd 0.007201f
C3741 vdd.n3158 gnd 0.007201f
C3742 vdd.n3159 gnd 0.007201f
C3743 vdd.n3160 gnd 0.008947f
C3744 vdd.n3162 gnd 0.008947f
C3745 vdd.n3164 gnd 0.008947f
C3746 vdd.n3165 gnd 0.007201f
C3747 vdd.n3166 gnd 0.007201f
C3748 vdd.n3167 gnd 0.006013f
C3749 vdd.n3168 gnd 0.008947f
C3750 vdd.n3170 gnd 0.008947f
C3751 vdd.n3172 gnd 0.008947f
C3752 vdd.n3173 gnd 0.006013f
C3753 vdd.n3174 gnd 0.007201f
C3754 vdd.n3175 gnd 0.007201f
C3755 vdd.n3176 gnd 0.008947f
C3756 vdd.n3178 gnd 0.008947f
C3757 vdd.n3180 gnd 0.008947f
C3758 vdd.n3181 gnd 0.007201f
C3759 vdd.n3182 gnd 0.007201f
C3760 vdd.n3183 gnd 0.007201f
C3761 vdd.n3184 gnd 0.008947f
C3762 vdd.n3186 gnd 0.008947f
C3763 vdd.n3188 gnd 0.008947f
C3764 vdd.n3189 gnd 0.007201f
C3765 vdd.n3190 gnd 0.007201f
C3766 vdd.n3191 gnd 0.007201f
C3767 vdd.n3192 gnd 0.008947f
C3768 vdd.n3194 gnd 0.008947f
C3769 vdd.n3195 gnd 0.008947f
C3770 vdd.n3196 gnd 0.007201f
C3771 vdd.n3197 gnd 0.007201f
C3772 vdd.n3198 gnd 0.008947f
C3773 vdd.n3199 gnd 0.008947f
C3774 vdd.n3200 gnd 0.007201f
C3775 vdd.n3201 gnd 0.007201f
C3776 vdd.n3202 gnd 0.008947f
C3777 vdd.n3203 gnd 0.008947f
C3778 vdd.n3205 gnd 0.008947f
C3779 vdd.n3206 gnd 0.007201f
C3780 vdd.n3207 gnd 0.005977f
C3781 vdd.n3208 gnd 0.021413f
C3782 vdd.n3209 gnd 0.021084f
C3783 vdd.n3210 gnd 0.005977f
C3784 vdd.n3211 gnd 0.021084f
C3785 vdd.n3212 gnd 1.25717f
C3786 vdd.n3213 gnd 0.021084f
C3787 vdd.n3214 gnd 0.005977f
C3788 vdd.n3215 gnd 0.021084f
C3789 vdd.n3216 gnd 0.008947f
C3790 vdd.n3217 gnd 0.008947f
C3791 vdd.n3218 gnd 0.007201f
C3792 vdd.n3219 gnd 0.008947f
C3793 vdd.n3220 gnd 0.914309f
C3794 vdd.n3221 gnd 0.008947f
C3795 vdd.n3222 gnd 0.007201f
C3796 vdd.n3223 gnd 0.008947f
C3797 vdd.n3224 gnd 0.008947f
C3798 vdd.n3225 gnd 0.008947f
C3799 vdd.n3226 gnd 0.007201f
C3800 vdd.n3227 gnd 0.008947f
C3801 vdd.n3228 gnd 0.809163f
C3802 vdd.n3229 gnd 0.008947f
C3803 vdd.n3230 gnd 0.007201f
C3804 vdd.n3231 gnd 0.008947f
C3805 vdd.n3232 gnd 0.008947f
C3806 vdd.n3233 gnd 0.008947f
C3807 vdd.n3234 gnd 0.007201f
C3808 vdd.n3235 gnd 0.008947f
C3809 vdd.t180 gnd 0.457154f
C3810 vdd.n3236 gnd 0.653731f
C3811 vdd.n3237 gnd 0.008947f
C3812 vdd.n3238 gnd 0.007201f
C3813 vdd.n3239 gnd 0.008947f
C3814 vdd.n3240 gnd 0.008947f
C3815 vdd.n3241 gnd 0.008947f
C3816 vdd.n3242 gnd 0.007201f
C3817 vdd.n3243 gnd 0.008947f
C3818 vdd.n3244 gnd 0.498298f
C3819 vdd.n3245 gnd 0.008947f
C3820 vdd.n3246 gnd 0.007201f
C3821 vdd.n3247 gnd 0.008947f
C3822 vdd.n3248 gnd 0.008947f
C3823 vdd.n3249 gnd 0.008947f
C3824 vdd.n3250 gnd 0.007201f
C3825 vdd.n3251 gnd 0.008947f
C3826 vdd.n3252 gnd 0.644588f
C3827 vdd.n3253 gnd 0.571443f
C3828 vdd.n3254 gnd 0.008947f
C3829 vdd.n3255 gnd 0.007201f
C3830 vdd.n3256 gnd 0.008947f
C3831 vdd.n3257 gnd 0.008947f
C3832 vdd.n3258 gnd 0.008947f
C3833 vdd.n3259 gnd 0.007201f
C3834 vdd.n3260 gnd 0.008947f
C3835 vdd.n3261 gnd 0.726875f
C3836 vdd.n3262 gnd 0.008947f
C3837 vdd.n3263 gnd 0.007201f
C3838 vdd.n3264 gnd 0.008947f
C3839 vdd.n3265 gnd 0.008947f
C3840 vdd.n3266 gnd 0.008947f
C3841 vdd.n3267 gnd 0.007201f
C3842 vdd.n3268 gnd 0.007201f
C3843 vdd.n3269 gnd 0.007201f
C3844 vdd.n3270 gnd 0.008947f
C3845 vdd.n3271 gnd 0.008947f
C3846 vdd.n3272 gnd 0.008947f
C3847 vdd.n3273 gnd 0.007201f
C3848 vdd.n3274 gnd 0.007201f
C3849 vdd.n3275 gnd 0.007201f
C3850 vdd.n3276 gnd 0.008947f
C3851 vdd.n3277 gnd 0.008947f
C3852 vdd.n3278 gnd 0.008947f
C3853 vdd.n3279 gnd 0.007201f
C3854 vdd.n3280 gnd 0.007201f
C3855 vdd.n3281 gnd 0.007201f
C3856 vdd.n3282 gnd 0.008947f
C3857 vdd.n3283 gnd 0.008947f
C3858 vdd.n3284 gnd 0.008947f
C3859 vdd.n3285 gnd 0.007201f
C3860 vdd.n3286 gnd 0.007201f
C3861 vdd.n3287 gnd 0.005977f
C3862 vdd.n3288 gnd 0.021084f
C3863 vdd.n3289 gnd 0.021413f
C3864 vdd.n3291 gnd 0.021413f
C3865 vdd.n3292 gnd 0.00342f
C3866 vdd.t35 gnd 0.110068f
C3867 vdd.t34 gnd 0.117632f
C3868 vdd.t33 gnd 0.143747f
C3869 vdd.n3293 gnd 0.184263f
C3870 vdd.n3294 gnd 0.155535f
C3871 vdd.n3295 gnd 0.01181f
C3872 vdd.n3296 gnd 0.003781f
C3873 vdd.n3297 gnd 0.007201f
C3874 vdd.n3298 gnd 0.008947f
C3875 vdd.n3300 gnd 0.008947f
C3876 vdd.n3301 gnd 0.008947f
C3877 vdd.n3302 gnd 0.007201f
C3878 vdd.n3303 gnd 0.007201f
C3879 vdd.n3304 gnd 0.007201f
C3880 vdd.n3305 gnd 0.008947f
C3881 vdd.n3307 gnd 0.008947f
C3882 vdd.n3308 gnd 0.008947f
C3883 vdd.n3309 gnd 0.007201f
C3884 vdd.n3310 gnd 0.007201f
C3885 vdd.n3311 gnd 0.007201f
C3886 vdd.n3312 gnd 0.008947f
C3887 vdd.n3314 gnd 0.008947f
C3888 vdd.n3315 gnd 0.008947f
C3889 vdd.n3316 gnd 0.007201f
C3890 vdd.n3317 gnd 0.007201f
C3891 vdd.n3318 gnd 0.007201f
C3892 vdd.n3319 gnd 0.008947f
C3893 vdd.n3321 gnd 0.008947f
C3894 vdd.n3322 gnd 0.008947f
C3895 vdd.n3323 gnd 0.007201f
C3896 vdd.n3324 gnd 0.007201f
C3897 vdd.n3325 gnd 0.007201f
C3898 vdd.n3326 gnd 0.008947f
C3899 vdd.n3328 gnd 0.008947f
C3900 vdd.n3329 gnd 0.008947f
C3901 vdd.n3330 gnd 0.007201f
C3902 vdd.n3331 gnd 0.008947f
C3903 vdd.n3332 gnd 0.008947f
C3904 vdd.n3333 gnd 0.008947f
C3905 vdd.n3334 gnd 0.01541f
C3906 vdd.n3335 gnd 0.004897f
C3907 vdd.n3336 gnd 0.007201f
C3908 vdd.n3337 gnd 0.008947f
C3909 vdd.n3339 gnd 0.008947f
C3910 vdd.n3340 gnd 0.008947f
C3911 vdd.n3341 gnd 0.007201f
C3912 vdd.n3342 gnd 0.007201f
C3913 vdd.n3343 gnd 0.007201f
C3914 vdd.n3344 gnd 0.008947f
C3915 vdd.n3346 gnd 0.008947f
C3916 vdd.n3347 gnd 0.008947f
C3917 vdd.n3348 gnd 0.007201f
C3918 vdd.n3349 gnd 0.007201f
C3919 vdd.n3350 gnd 0.007201f
C3920 vdd.n3351 gnd 0.008947f
C3921 vdd.n3353 gnd 0.008947f
C3922 vdd.n3354 gnd 0.008947f
C3923 vdd.n3355 gnd 0.007201f
C3924 vdd.n3356 gnd 0.007201f
C3925 vdd.n3357 gnd 0.007201f
C3926 vdd.n3358 gnd 0.008947f
C3927 vdd.n3360 gnd 0.008947f
C3928 vdd.n3361 gnd 0.008947f
C3929 vdd.n3362 gnd 0.007201f
C3930 vdd.n3363 gnd 0.007201f
C3931 vdd.n3364 gnd 0.007201f
C3932 vdd.n3365 gnd 0.008947f
C3933 vdd.n3367 gnd 0.008947f
C3934 vdd.n3368 gnd 0.008947f
C3935 vdd.n3369 gnd 0.007201f
C3936 vdd.n3370 gnd 0.008947f
C3937 vdd.n3371 gnd 0.008947f
C3938 vdd.n3372 gnd 0.008947f
C3939 vdd.n3373 gnd 0.01541f
C3940 vdd.n3374 gnd 0.006013f
C3941 vdd.n3375 gnd 0.007201f
C3942 vdd.n3376 gnd 0.008947f
C3943 vdd.n3378 gnd 0.008947f
C3944 vdd.n3379 gnd 0.008947f
C3945 vdd.n3380 gnd 0.007201f
C3946 vdd.n3381 gnd 0.007201f
C3947 vdd.n3382 gnd 0.007201f
C3948 vdd.n3383 gnd 0.008947f
C3949 vdd.n3385 gnd 0.008947f
C3950 vdd.n3386 gnd 0.008947f
C3951 vdd.n3387 gnd 0.007201f
C3952 vdd.n3388 gnd 0.007201f
C3953 vdd.n3389 gnd 0.007201f
C3954 vdd.n3390 gnd 0.008947f
C3955 vdd.n3392 gnd 0.008947f
C3956 vdd.n3393 gnd 0.008947f
C3957 vdd.n3394 gnd 0.007201f
C3958 vdd.n3395 gnd 0.007201f
C3959 vdd.n3396 gnd 0.007201f
C3960 vdd.n3397 gnd 0.008947f
C3961 vdd.n3399 gnd 0.008947f
C3962 vdd.n3400 gnd 0.008947f
C3963 vdd.n3402 gnd 0.008947f
C3964 vdd.n3403 gnd 0.007201f
C3965 vdd.n3404 gnd 0.007201f
C3966 vdd.n3405 gnd 0.005977f
C3967 vdd.n3406 gnd 0.021413f
C3968 vdd.n3407 gnd 0.021084f
C3969 vdd.n3408 gnd 0.005977f
C3970 vdd.n3409 gnd 0.021084f
C3971 vdd.n3410 gnd 1.28918f
C3972 vdd.n3411 gnd 0.516584f
C3973 vdd.t23 gnd 0.457154f
C3974 vdd.n3412 gnd 0.854879f
C3975 vdd.n3413 gnd 0.008947f
C3976 vdd.n3414 gnd 0.007201f
C3977 vdd.n3415 gnd 0.007201f
C3978 vdd.n3416 gnd 0.007201f
C3979 vdd.n3417 gnd 0.008947f
C3980 vdd.n3418 gnd 0.900594f
C3981 vdd.t160 gnd 0.457154f
C3982 vdd.n3419 gnd 0.470869f
C3983 vdd.n3420 gnd 0.745162f
C3984 vdd.n3421 gnd 0.008947f
C3985 vdd.n3422 gnd 0.007201f
C3986 vdd.n3423 gnd 0.007201f
C3987 vdd.n3424 gnd 0.007201f
C3988 vdd.n3425 gnd 0.008947f
C3989 vdd.n3426 gnd 0.589729f
C3990 vdd.t186 gnd 0.457154f
C3991 vdd.n3427 gnd 0.758876f
C3992 vdd.t152 gnd 0.457154f
C3993 vdd.n3428 gnd 0.480012f
C3994 vdd.n3429 gnd 0.008947f
C3995 vdd.n3430 gnd 0.007201f
C3996 vdd.n3431 gnd 0.007201f
C3997 vdd.n3432 gnd 0.007201f
C3998 vdd.n3433 gnd 0.008947f
C3999 vdd.n3434 gnd 0.635445f
C4000 vdd.n3435 gnd 0.580586f
C4001 vdd.t198 gnd 0.457154f
C4002 vdd.n3436 gnd 0.758876f
C4003 vdd.n3437 gnd 0.008947f
C4004 vdd.n3438 gnd 0.007201f
C4005 vdd.n3439 gnd 0.532576f
C4006 vdd.n3440 gnd 2.29632f
C4007 a_n2982_13878.n0 gnd 2.53375f
C4008 a_n2982_13878.n1 gnd 3.78544f
C4009 a_n2982_13878.n2 gnd 3.42814f
C4010 a_n2982_13878.n3 gnd 0.971817f
C4011 a_n2982_13878.n4 gnd 0.20945f
C4012 a_n2982_13878.n5 gnd 0.20945f
C4013 a_n2982_13878.n6 gnd 0.458034f
C4014 a_n2982_13878.n7 gnd 0.20945f
C4015 a_n2982_13878.n8 gnd 0.27462f
C4016 a_n2982_13878.n9 gnd 0.20945f
C4017 a_n2982_13878.n10 gnd 0.20945f
C4018 a_n2982_13878.n11 gnd 0.791576f
C4019 a_n2982_13878.n12 gnd 0.20945f
C4020 a_n2982_13878.n13 gnd 0.904041f
C4021 a_n2982_13878.n14 gnd 0.198733f
C4022 a_n2982_13878.n15 gnd 0.146371f
C4023 a_n2982_13878.n16 gnd 0.230048f
C4024 a_n2982_13878.n17 gnd 0.177686f
C4025 a_n2982_13878.n18 gnd 0.198733f
C4026 a_n2982_13878.n19 gnd 0.146371f
C4027 a_n2982_13878.n20 gnd 0.956403f
C4028 a_n2982_13878.n21 gnd 0.20945f
C4029 a_n2982_13878.n22 gnd 0.73719f
C4030 a_n2982_13878.n23 gnd 0.20945f
C4031 a_n2982_13878.n24 gnd 0.20945f
C4032 a_n2982_13878.n25 gnd 0.477018f
C4033 a_n2982_13878.n26 gnd 0.27462f
C4034 a_n2982_13878.n27 gnd 0.20945f
C4035 a_n2982_13878.n28 gnd 0.529381f
C4036 a_n2982_13878.n29 gnd 0.20945f
C4037 a_n2982_13878.n30 gnd 0.20945f
C4038 a_n2982_13878.n31 gnd 0.931898f
C4039 a_n2982_13878.n32 gnd 0.27462f
C4040 a_n2982_13878.n33 gnd 3.08362f
C4041 a_n2982_13878.n34 gnd 0.27462f
C4042 a_n2982_13878.n35 gnd 1.16191f
C4043 a_n2982_13878.n36 gnd 2.12168f
C4044 a_n2982_13878.n37 gnd 1.72437f
C4045 a_n2982_13878.n38 gnd 1.16191f
C4046 a_n2982_13878.n39 gnd 1.72437f
C4047 a_n2982_13878.n40 gnd 2.32061f
C4048 a_n2982_13878.n41 gnd 0.008404f
C4049 a_n2982_13878.n42 gnd 4.05e-19
C4050 a_n2982_13878.n44 gnd 0.008109f
C4051 a_n2982_13878.n45 gnd 0.011792f
C4052 a_n2982_13878.n46 gnd 0.007801f
C4053 a_n2982_13878.n48 gnd 0.277816f
C4054 a_n2982_13878.n49 gnd 0.008404f
C4055 a_n2982_13878.n50 gnd 4.05e-19
C4056 a_n2982_13878.n52 gnd 0.008109f
C4057 a_n2982_13878.n53 gnd 0.011792f
C4058 a_n2982_13878.n54 gnd 0.007801f
C4059 a_n2982_13878.n56 gnd 0.277816f
C4060 a_n2982_13878.n57 gnd 0.008109f
C4061 a_n2982_13878.n58 gnd 0.276683f
C4062 a_n2982_13878.n59 gnd 0.008109f
C4063 a_n2982_13878.n60 gnd 0.276683f
C4064 a_n2982_13878.n61 gnd 0.008109f
C4065 a_n2982_13878.n62 gnd 0.276683f
C4066 a_n2982_13878.n63 gnd 0.008109f
C4067 a_n2982_13878.n64 gnd 1.64574f
C4068 a_n2982_13878.n65 gnd 0.276683f
C4069 a_n2982_13878.n66 gnd 0.277816f
C4070 a_n2982_13878.n68 gnd 0.007801f
C4071 a_n2982_13878.n69 gnd 0.011792f
C4072 a_n2982_13878.n70 gnd 0.008109f
C4073 a_n2982_13878.n72 gnd 4.05e-19
C4074 a_n2982_13878.n73 gnd 0.008404f
C4075 a_n2982_13878.n74 gnd 0.104725f
C4076 a_n2982_13878.n75 gnd 0.008404f
C4077 a_n2982_13878.n76 gnd 4.05e-19
C4078 a_n2982_13878.n78 gnd 0.008109f
C4079 a_n2982_13878.n79 gnd 0.011792f
C4080 a_n2982_13878.n80 gnd 0.007801f
C4081 a_n2982_13878.n82 gnd 0.277816f
C4082 a_n2982_13878.t44 gnd 0.145277f
C4083 a_n2982_13878.t40 gnd 1.3603f
C4084 a_n2982_13878.t56 gnd 0.145277f
C4085 a_n2982_13878.t48 gnd 0.145277f
C4086 a_n2982_13878.n83 gnd 1.02333f
C4087 a_n2982_13878.t57 gnd 0.675756f
C4088 a_n2982_13878.n84 gnd 0.29709f
C4089 a_n2982_13878.t17 gnd 0.675756f
C4090 a_n2982_13878.t19 gnd 0.675756f
C4091 a_n2982_13878.n85 gnd 0.288167f
C4092 a_n2982_13878.t13 gnd 0.675756f
C4093 a_n2982_13878.n86 gnd 0.299644f
C4094 a_n2982_13878.t59 gnd 0.675756f
C4095 a_n2982_13878.t47 gnd 0.675756f
C4096 a_n2982_13878.n87 gnd 0.293009f
C4097 a_n2982_13878.t39 gnd 0.689824f
C4098 a_n2982_13878.t78 gnd 0.675756f
C4099 a_n2982_13878.n88 gnd 0.29709f
C4100 a_n2982_13878.t88 gnd 0.675756f
C4101 a_n2982_13878.t93 gnd 0.675756f
C4102 a_n2982_13878.n89 gnd 0.288167f
C4103 a_n2982_13878.t97 gnd 0.675756f
C4104 a_n2982_13878.n90 gnd 0.299644f
C4105 a_n2982_13878.t68 gnd 0.675756f
C4106 a_n2982_13878.t71 gnd 0.675756f
C4107 a_n2982_13878.n91 gnd 0.293009f
C4108 a_n2982_13878.t101 gnd 0.689824f
C4109 a_n2982_13878.t49 gnd 0.686627f
C4110 a_n2982_13878.t15 gnd 0.675756f
C4111 a_n2982_13878.t33 gnd 0.675756f
C4112 a_n2982_13878.t45 gnd 0.675756f
C4113 a_n2982_13878.n92 gnd 0.293584f
C4114 a_n2982_13878.t37 gnd 0.675756f
C4115 a_n2982_13878.t51 gnd 0.675756f
C4116 a_n2982_13878.t29 gnd 0.675756f
C4117 a_n2982_13878.n93 gnd 0.297105f
C4118 a_n2982_13878.t23 gnd 0.675756f
C4119 a_n2982_13878.t53 gnd 0.675756f
C4120 a_n2982_13878.t25 gnd 0.675756f
C4121 a_n2982_13878.n94 gnd 0.293009f
C4122 a_n2982_13878.t35 gnd 0.675756f
C4123 a_n2982_13878.t21 gnd 0.689824f
C4124 a_n2982_13878.t102 gnd 0.689824f
C4125 a_n2982_13878.t79 gnd 0.675756f
C4126 a_n2982_13878.t84 gnd 0.675756f
C4127 a_n2982_13878.t72 gnd 0.675756f
C4128 a_n2982_13878.n95 gnd 0.296971f
C4129 a_n2982_13878.t89 gnd 0.675756f
C4130 a_n2982_13878.t98 gnd 0.675756f
C4131 a_n2982_13878.t99 gnd 0.675756f
C4132 a_n2982_13878.n96 gnd 0.293332f
C4133 a_n2982_13878.t66 gnd 0.675756f
C4134 a_n2982_13878.t81 gnd 0.675756f
C4135 a_n2982_13878.t69 gnd 0.675756f
C4136 a_n2982_13878.n97 gnd 0.29709f
C4137 a_n2982_13878.t76 gnd 0.675756f
C4138 a_n2982_13878.t95 gnd 0.686627f
C4139 a_n2982_13878.n98 gnd 0.299206f
C4140 a_n2982_13878.n99 gnd 0.293584f
C4141 a_n2982_13878.n100 gnd 0.288167f
C4142 a_n2982_13878.n101 gnd 0.297105f
C4143 a_n2982_13878.n102 gnd 0.299644f
C4144 a_n2982_13878.n103 gnd 0.293009f
C4145 a_n2982_13878.n104 gnd 0.299205f
C4146 a_n2982_13878.t7 gnd 0.112993f
C4147 a_n2982_13878.t4 gnd 0.112993f
C4148 a_n2982_13878.n105 gnd 1.00066f
C4149 a_n2982_13878.t10 gnd 0.112993f
C4150 a_n2982_13878.t1 gnd 0.112993f
C4151 a_n2982_13878.n106 gnd 0.998444f
C4152 a_n2982_13878.t6 gnd 0.112993f
C4153 a_n2982_13878.t5 gnd 0.112993f
C4154 a_n2982_13878.n107 gnd 1.00066f
C4155 a_n2982_13878.t61 gnd 0.112993f
C4156 a_n2982_13878.t2 gnd 0.112993f
C4157 a_n2982_13878.n108 gnd 0.998444f
C4158 a_n2982_13878.t0 gnd 0.112993f
C4159 a_n2982_13878.t62 gnd 0.112993f
C4160 a_n2982_13878.n109 gnd 0.998444f
C4161 a_n2982_13878.t63 gnd 0.112993f
C4162 a_n2982_13878.t9 gnd 0.112993f
C4163 a_n2982_13878.n110 gnd 0.998444f
C4164 a_n2982_13878.t8 gnd 0.112993f
C4165 a_n2982_13878.t11 gnd 0.112993f
C4166 a_n2982_13878.n111 gnd 1.00066f
C4167 a_n2982_13878.t3 gnd 0.112993f
C4168 a_n2982_13878.t12 gnd 0.112993f
C4169 a_n2982_13878.n112 gnd 0.998444f
C4170 a_n2982_13878.n113 gnd 0.299205f
C4171 a_n2982_13878.n114 gnd 0.296971f
C4172 a_n2982_13878.n115 gnd 0.299644f
C4173 a_n2982_13878.n116 gnd 0.293332f
C4174 a_n2982_13878.n117 gnd 0.288167f
C4175 a_n2982_13878.n118 gnd 0.29709f
C4176 a_n2982_13878.n119 gnd 0.299206f
C4177 a_n2982_13878.t22 gnd 1.3603f
C4178 a_n2982_13878.t26 gnd 0.145277f
C4179 a_n2982_13878.t36 gnd 0.145277f
C4180 a_n2982_13878.n120 gnd 1.02333f
C4181 a_n2982_13878.t24 gnd 0.145277f
C4182 a_n2982_13878.t54 gnd 0.145277f
C4183 a_n2982_13878.n121 gnd 1.02333f
C4184 a_n2982_13878.t52 gnd 0.145277f
C4185 a_n2982_13878.t30 gnd 0.145277f
C4186 a_n2982_13878.n122 gnd 1.02333f
C4187 a_n2982_13878.t46 gnd 0.145277f
C4188 a_n2982_13878.t38 gnd 0.145277f
C4189 a_n2982_13878.n123 gnd 1.02333f
C4190 a_n2982_13878.t16 gnd 0.145277f
C4191 a_n2982_13878.t34 gnd 0.145277f
C4192 a_n2982_13878.n124 gnd 1.02333f
C4193 a_n2982_13878.t50 gnd 1.35759f
C4194 a_n2982_13878.n125 gnd 0.994805f
C4195 a_n2982_13878.t77 gnd 0.675756f
C4196 a_n2982_13878.t87 gnd 0.675756f
C4197 a_n2982_13878.t103 gnd 0.675756f
C4198 a_n2982_13878.n126 gnd 0.297105f
C4199 a_n2982_13878.t90 gnd 0.675756f
C4200 a_n2982_13878.t73 gnd 0.675756f
C4201 a_n2982_13878.t74 gnd 0.675756f
C4202 a_n2982_13878.n127 gnd 0.297105f
C4203 a_n2982_13878.t94 gnd 0.675756f
C4204 a_n2982_13878.t83 gnd 0.675756f
C4205 a_n2982_13878.t82 gnd 0.675756f
C4206 a_n2982_13878.n128 gnd 0.297105f
C4207 a_n2982_13878.t86 gnd 0.675756f
C4208 a_n2982_13878.t75 gnd 0.675756f
C4209 a_n2982_13878.t64 gnd 0.675756f
C4210 a_n2982_13878.n129 gnd 0.297105f
C4211 a_n2982_13878.t91 gnd 0.687079f
C4212 a_n2982_13878.n130 gnd 0.293332f
C4213 a_n2982_13878.n131 gnd 0.288005f
C4214 a_n2982_13878.t100 gnd 0.687079f
C4215 a_n2982_13878.n132 gnd 0.293332f
C4216 a_n2982_13878.n133 gnd 0.288005f
C4217 a_n2982_13878.t85 gnd 0.687079f
C4218 a_n2982_13878.n134 gnd 0.293332f
C4219 a_n2982_13878.n135 gnd 0.288005f
C4220 a_n2982_13878.t80 gnd 0.687079f
C4221 a_n2982_13878.n136 gnd 0.293332f
C4222 a_n2982_13878.n137 gnd 0.288005f
C4223 a_n2982_13878.n138 gnd 1.32386f
C4224 a_n2982_13878.t70 gnd 0.675756f
C4225 a_n2982_13878.n139 gnd 0.299205f
C4226 a_n2982_13878.t96 gnd 0.675756f
C4227 a_n2982_13878.n140 gnd 0.296971f
C4228 a_n2982_13878.n141 gnd 0.297105f
C4229 a_n2982_13878.t92 gnd 0.675756f
C4230 a_n2982_13878.n142 gnd 0.293332f
C4231 a_n2982_13878.t65 gnd 0.675756f
C4232 a_n2982_13878.n143 gnd 0.293584f
C4233 a_n2982_13878.n144 gnd 0.299206f
C4234 a_n2982_13878.t67 gnd 0.686627f
C4235 a_n2982_13878.t55 gnd 0.675756f
C4236 a_n2982_13878.n145 gnd 0.299205f
C4237 a_n2982_13878.t43 gnd 0.675756f
C4238 a_n2982_13878.n146 gnd 0.296971f
C4239 a_n2982_13878.n147 gnd 0.297105f
C4240 a_n2982_13878.t27 gnd 0.675756f
C4241 a_n2982_13878.n148 gnd 0.293332f
C4242 a_n2982_13878.t41 gnd 0.675756f
C4243 a_n2982_13878.n149 gnd 0.293584f
C4244 a_n2982_13878.n150 gnd 0.299206f
C4245 a_n2982_13878.t31 gnd 0.686627f
C4246 a_n2982_13878.n151 gnd 1.30834f
C4247 a_n2982_13878.t32 gnd 1.35758f
C4248 a_n2982_13878.t58 gnd 0.145277f
C4249 a_n2982_13878.t18 gnd 0.145277f
C4250 a_n2982_13878.n152 gnd 1.02333f
C4251 a_n2982_13878.t20 gnd 0.145277f
C4252 a_n2982_13878.t42 gnd 0.145277f
C4253 a_n2982_13878.n153 gnd 1.02333f
C4254 a_n2982_13878.t60 gnd 0.145277f
C4255 a_n2982_13878.t28 gnd 0.145277f
C4256 a_n2982_13878.n154 gnd 1.02333f
C4257 a_n2982_13878.n155 gnd 1.02333f
C4258 a_n2982_13878.t14 gnd 0.145277f
C4259 CSoutput.n0 gnd 0.041923f
C4260 CSoutput.t174 gnd 0.277311f
C4261 CSoutput.n1 gnd 0.12522f
C4262 CSoutput.n2 gnd 0.041923f
C4263 CSoutput.t181 gnd 0.277311f
C4264 CSoutput.n3 gnd 0.033227f
C4265 CSoutput.n4 gnd 0.041923f
C4266 CSoutput.t188 gnd 0.277311f
C4267 CSoutput.n5 gnd 0.028652f
C4268 CSoutput.n6 gnd 0.041923f
C4269 CSoutput.t179 gnd 0.277311f
C4270 CSoutput.t177 gnd 0.277311f
C4271 CSoutput.n7 gnd 0.123855f
C4272 CSoutput.n8 gnd 0.041923f
C4273 CSoutput.t186 gnd 0.277311f
C4274 CSoutput.n9 gnd 0.027318f
C4275 CSoutput.n10 gnd 0.041923f
C4276 CSoutput.t169 gnd 0.277311f
C4277 CSoutput.t173 gnd 0.277311f
C4278 CSoutput.n11 gnd 0.123855f
C4279 CSoutput.n12 gnd 0.041923f
C4280 CSoutput.t184 gnd 0.277311f
C4281 CSoutput.n13 gnd 0.028652f
C4282 CSoutput.n14 gnd 0.041923f
C4283 CSoutput.t183 gnd 0.277311f
C4284 CSoutput.t171 gnd 0.277311f
C4285 CSoutput.n15 gnd 0.123855f
C4286 CSoutput.n16 gnd 0.041923f
C4287 CSoutput.t176 gnd 0.277311f
C4288 CSoutput.n17 gnd 0.030602f
C4289 CSoutput.t185 gnd 0.331394f
C4290 CSoutput.t182 gnd 0.277311f
C4291 CSoutput.n18 gnd 0.158115f
C4292 CSoutput.n19 gnd 0.153426f
C4293 CSoutput.n20 gnd 0.177993f
C4294 CSoutput.n21 gnd 0.041923f
C4295 CSoutput.n22 gnd 0.034989f
C4296 CSoutput.n23 gnd 0.123855f
C4297 CSoutput.n24 gnd 0.033729f
C4298 CSoutput.n25 gnd 0.033227f
C4299 CSoutput.n26 gnd 0.041923f
C4300 CSoutput.n27 gnd 0.041923f
C4301 CSoutput.n28 gnd 0.03472f
C4302 CSoutput.n29 gnd 0.029478f
C4303 CSoutput.n30 gnd 0.126612f
C4304 CSoutput.n31 gnd 0.029884f
C4305 CSoutput.n32 gnd 0.041923f
C4306 CSoutput.n33 gnd 0.041923f
C4307 CSoutput.n34 gnd 0.041923f
C4308 CSoutput.n35 gnd 0.03435f
C4309 CSoutput.n36 gnd 0.123855f
C4310 CSoutput.n37 gnd 0.032851f
C4311 CSoutput.n38 gnd 0.034105f
C4312 CSoutput.n39 gnd 0.041923f
C4313 CSoutput.n40 gnd 0.041923f
C4314 CSoutput.n41 gnd 0.034982f
C4315 CSoutput.n42 gnd 0.031974f
C4316 CSoutput.n43 gnd 0.123855f
C4317 CSoutput.n44 gnd 0.032784f
C4318 CSoutput.n45 gnd 0.041923f
C4319 CSoutput.n46 gnd 0.041923f
C4320 CSoutput.n47 gnd 0.041923f
C4321 CSoutput.n48 gnd 0.032784f
C4322 CSoutput.n49 gnd 0.123855f
C4323 CSoutput.n50 gnd 0.031974f
C4324 CSoutput.n51 gnd 0.034982f
C4325 CSoutput.n52 gnd 0.041923f
C4326 CSoutput.n53 gnd 0.041923f
C4327 CSoutput.n54 gnd 0.034105f
C4328 CSoutput.n55 gnd 0.032851f
C4329 CSoutput.n56 gnd 0.123855f
C4330 CSoutput.n57 gnd 0.03435f
C4331 CSoutput.n58 gnd 0.041923f
C4332 CSoutput.n59 gnd 0.041923f
C4333 CSoutput.n60 gnd 0.041923f
C4334 CSoutput.n61 gnd 0.029884f
C4335 CSoutput.n62 gnd 0.126612f
C4336 CSoutput.n63 gnd 0.029478f
C4337 CSoutput.t180 gnd 0.277311f
C4338 CSoutput.n64 gnd 0.123855f
C4339 CSoutput.n65 gnd 0.03472f
C4340 CSoutput.n66 gnd 0.041923f
C4341 CSoutput.n67 gnd 0.041923f
C4342 CSoutput.n68 gnd 0.041923f
C4343 CSoutput.n69 gnd 0.033729f
C4344 CSoutput.n70 gnd 0.123855f
C4345 CSoutput.n71 gnd 0.034989f
C4346 CSoutput.n72 gnd 0.030602f
C4347 CSoutput.n73 gnd 0.041923f
C4348 CSoutput.n74 gnd 0.041923f
C4349 CSoutput.n75 gnd 0.031736f
C4350 CSoutput.n76 gnd 0.018848f
C4351 CSoutput.t187 gnd 0.311579f
C4352 CSoutput.n77 gnd 0.15478f
C4353 CSoutput.n78 gnd 0.633197f
C4354 CSoutput.t134 gnd 0.052293f
C4355 CSoutput.t105 gnd 0.052293f
C4356 CSoutput.n79 gnd 0.404869f
C4357 CSoutput.t112 gnd 0.052293f
C4358 CSoutput.t143 gnd 0.052293f
C4359 CSoutput.n80 gnd 0.404147f
C4360 CSoutput.n81 gnd 0.410209f
C4361 CSoutput.t152 gnd 0.052293f
C4362 CSoutput.t158 gnd 0.052293f
C4363 CSoutput.n82 gnd 0.404147f
C4364 CSoutput.n83 gnd 0.202134f
C4365 CSoutput.t127 gnd 0.052293f
C4366 CSoutput.t164 gnd 0.052293f
C4367 CSoutput.n84 gnd 0.404147f
C4368 CSoutput.n85 gnd 0.202134f
C4369 CSoutput.t118 gnd 0.052293f
C4370 CSoutput.t121 gnd 0.052293f
C4371 CSoutput.n86 gnd 0.404147f
C4372 CSoutput.n87 gnd 0.202134f
C4373 CSoutput.t104 gnd 0.052293f
C4374 CSoutput.t108 gnd 0.052293f
C4375 CSoutput.n88 gnd 0.404147f
C4376 CSoutput.n89 gnd 0.370667f
C4377 CSoutput.t119 gnd 0.052293f
C4378 CSoutput.t149 gnd 0.052293f
C4379 CSoutput.n90 gnd 0.404869f
C4380 CSoutput.t132 gnd 0.052293f
C4381 CSoutput.t163 gnd 0.052293f
C4382 CSoutput.n91 gnd 0.404147f
C4383 CSoutput.n92 gnd 0.410209f
C4384 CSoutput.t106 gnd 0.052293f
C4385 CSoutput.t151 gnd 0.052293f
C4386 CSoutput.n93 gnd 0.404147f
C4387 CSoutput.n94 gnd 0.202134f
C4388 CSoutput.t131 gnd 0.052293f
C4389 CSoutput.t129 gnd 0.052293f
C4390 CSoutput.n95 gnd 0.404147f
C4391 CSoutput.n96 gnd 0.202134f
C4392 CSoutput.t159 gnd 0.052293f
C4393 CSoutput.t141 gnd 0.052293f
C4394 CSoutput.n97 gnd 0.404147f
C4395 CSoutput.n98 gnd 0.202134f
C4396 CSoutput.t154 gnd 0.052293f
C4397 CSoutput.t167 gnd 0.052293f
C4398 CSoutput.n99 gnd 0.404147f
C4399 CSoutput.n100 gnd 0.301432f
C4400 CSoutput.n101 gnd 0.380104f
C4401 CSoutput.t125 gnd 0.052293f
C4402 CSoutput.t142 gnd 0.052293f
C4403 CSoutput.n102 gnd 0.404869f
C4404 CSoutput.t157 gnd 0.052293f
C4405 CSoutput.t135 gnd 0.052293f
C4406 CSoutput.n103 gnd 0.404147f
C4407 CSoutput.n104 gnd 0.410209f
C4408 CSoutput.t124 gnd 0.052293f
C4409 CSoutput.t100 gnd 0.052293f
C4410 CSoutput.n105 gnd 0.404147f
C4411 CSoutput.n106 gnd 0.202134f
C4412 CSoutput.t156 gnd 0.052293f
C4413 CSoutput.t155 gnd 0.052293f
C4414 CSoutput.n107 gnd 0.404147f
C4415 CSoutput.n108 gnd 0.202134f
C4416 CSoutput.t110 gnd 0.052293f
C4417 CSoutput.t166 gnd 0.052293f
C4418 CSoutput.n109 gnd 0.404147f
C4419 CSoutput.n110 gnd 0.202134f
C4420 CSoutput.t128 gnd 0.052293f
C4421 CSoutput.t117 gnd 0.052293f
C4422 CSoutput.n111 gnd 0.404147f
C4423 CSoutput.n112 gnd 0.301432f
C4424 CSoutput.n113 gnd 0.424859f
C4425 CSoutput.n114 gnd 7.91342f
C4426 CSoutput.n116 gnd 0.741609f
C4427 CSoutput.n117 gnd 0.556207f
C4428 CSoutput.n118 gnd 0.741609f
C4429 CSoutput.n119 gnd 0.741609f
C4430 CSoutput.n120 gnd 1.99664f
C4431 CSoutput.n121 gnd 0.741609f
C4432 CSoutput.n122 gnd 0.741609f
C4433 CSoutput.t175 gnd 0.927011f
C4434 CSoutput.n123 gnd 0.741609f
C4435 CSoutput.n124 gnd 0.741609f
C4436 CSoutput.n128 gnd 0.741609f
C4437 CSoutput.n132 gnd 0.741609f
C4438 CSoutput.n133 gnd 0.741609f
C4439 CSoutput.n135 gnd 0.741609f
C4440 CSoutput.n140 gnd 0.741609f
C4441 CSoutput.n142 gnd 0.741609f
C4442 CSoutput.n143 gnd 0.741609f
C4443 CSoutput.n145 gnd 0.741609f
C4444 CSoutput.n146 gnd 0.741609f
C4445 CSoutput.n148 gnd 0.741609f
C4446 CSoutput.t170 gnd 12.3922f
C4447 CSoutput.n150 gnd 0.741609f
C4448 CSoutput.n151 gnd 0.556207f
C4449 CSoutput.n152 gnd 0.741609f
C4450 CSoutput.n153 gnd 0.741609f
C4451 CSoutput.n154 gnd 1.99664f
C4452 CSoutput.n155 gnd 0.741609f
C4453 CSoutput.n156 gnd 0.741609f
C4454 CSoutput.t189 gnd 0.927011f
C4455 CSoutput.n157 gnd 0.741609f
C4456 CSoutput.n158 gnd 0.741609f
C4457 CSoutput.n162 gnd 0.741609f
C4458 CSoutput.n166 gnd 0.741609f
C4459 CSoutput.n167 gnd 0.741609f
C4460 CSoutput.n169 gnd 0.741609f
C4461 CSoutput.n174 gnd 0.741609f
C4462 CSoutput.n176 gnd 0.741609f
C4463 CSoutput.n177 gnd 0.741609f
C4464 CSoutput.n179 gnd 0.741609f
C4465 CSoutput.n180 gnd 0.741609f
C4466 CSoutput.n182 gnd 0.741609f
C4467 CSoutput.n183 gnd 0.556207f
C4468 CSoutput.n185 gnd 0.741609f
C4469 CSoutput.n186 gnd 0.556207f
C4470 CSoutput.n187 gnd 0.741609f
C4471 CSoutput.n188 gnd 0.741609f
C4472 CSoutput.n189 gnd 1.99664f
C4473 CSoutput.n190 gnd 0.741609f
C4474 CSoutput.n191 gnd 0.741609f
C4475 CSoutput.t168 gnd 0.927011f
C4476 CSoutput.n192 gnd 0.741609f
C4477 CSoutput.n193 gnd 1.99664f
C4478 CSoutput.n195 gnd 0.741609f
C4479 CSoutput.n196 gnd 0.741609f
C4480 CSoutput.n198 gnd 0.741609f
C4481 CSoutput.n199 gnd 0.741609f
C4482 CSoutput.t178 gnd 12.1903f
C4483 CSoutput.t172 gnd 12.3922f
C4484 CSoutput.n205 gnd 2.32654f
C4485 CSoutput.n206 gnd 9.47746f
C4486 CSoutput.n207 gnd 9.87404f
C4487 CSoutput.n212 gnd 2.52027f
C4488 CSoutput.n218 gnd 0.741609f
C4489 CSoutput.n220 gnd 0.741609f
C4490 CSoutput.n222 gnd 0.741609f
C4491 CSoutput.n224 gnd 0.741609f
C4492 CSoutput.n226 gnd 0.741609f
C4493 CSoutput.n232 gnd 0.741609f
C4494 CSoutput.n239 gnd 1.36057f
C4495 CSoutput.n240 gnd 1.36057f
C4496 CSoutput.n241 gnd 0.741609f
C4497 CSoutput.n242 gnd 0.741609f
C4498 CSoutput.n244 gnd 0.556207f
C4499 CSoutput.n245 gnd 0.476341f
C4500 CSoutput.n247 gnd 0.556207f
C4501 CSoutput.n248 gnd 0.476341f
C4502 CSoutput.n249 gnd 0.556207f
C4503 CSoutput.n251 gnd 0.741609f
C4504 CSoutput.n253 gnd 1.99664f
C4505 CSoutput.n254 gnd 2.32654f
C4506 CSoutput.n255 gnd 8.71683f
C4507 CSoutput.n257 gnd 0.556207f
C4508 CSoutput.n258 gnd 1.43115f
C4509 CSoutput.n259 gnd 0.556207f
C4510 CSoutput.n261 gnd 0.741609f
C4511 CSoutput.n263 gnd 1.99664f
C4512 CSoutput.n264 gnd 4.349f
C4513 CSoutput.t138 gnd 0.052293f
C4514 CSoutput.t103 gnd 0.052293f
C4515 CSoutput.n265 gnd 0.404869f
C4516 CSoutput.t98 gnd 0.052293f
C4517 CSoutput.t111 gnd 0.052293f
C4518 CSoutput.n266 gnd 0.404147f
C4519 CSoutput.n267 gnd 0.410209f
C4520 CSoutput.t136 gnd 0.052293f
C4521 CSoutput.t101 gnd 0.052293f
C4522 CSoutput.n268 gnd 0.404147f
C4523 CSoutput.n269 gnd 0.202134f
C4524 CSoutput.t147 gnd 0.052293f
C4525 CSoutput.t126 gnd 0.052293f
C4526 CSoutput.n270 gnd 0.404147f
C4527 CSoutput.n271 gnd 0.202134f
C4528 CSoutput.t120 gnd 0.052293f
C4529 CSoutput.t107 gnd 0.052293f
C4530 CSoutput.n272 gnd 0.404147f
C4531 CSoutput.n273 gnd 0.202134f
C4532 CSoutput.t115 gnd 0.052293f
C4533 CSoutput.t153 gnd 0.052293f
C4534 CSoutput.n274 gnd 0.404147f
C4535 CSoutput.n275 gnd 0.370667f
C4536 CSoutput.t144 gnd 0.052293f
C4537 CSoutput.t145 gnd 0.052293f
C4538 CSoutput.n276 gnd 0.404869f
C4539 CSoutput.t116 gnd 0.052293f
C4540 CSoutput.t109 gnd 0.052293f
C4541 CSoutput.n277 gnd 0.404147f
C4542 CSoutput.n278 gnd 0.410209f
C4543 CSoutput.t97 gnd 0.052293f
C4544 CSoutput.t139 gnd 0.052293f
C4545 CSoutput.n279 gnd 0.404147f
C4546 CSoutput.n280 gnd 0.202134f
C4547 CSoutput.t137 gnd 0.052293f
C4548 CSoutput.t114 gnd 0.052293f
C4549 CSoutput.n281 gnd 0.404147f
C4550 CSoutput.n282 gnd 0.202134f
C4551 CSoutput.t160 gnd 0.052293f
C4552 CSoutput.t99 gnd 0.052293f
C4553 CSoutput.n283 gnd 0.404147f
C4554 CSoutput.n284 gnd 0.202134f
C4555 CSoutput.t113 gnd 0.052293f
C4556 CSoutput.t133 gnd 0.052293f
C4557 CSoutput.n285 gnd 0.404147f
C4558 CSoutput.n286 gnd 0.301432f
C4559 CSoutput.n287 gnd 0.380104f
C4560 CSoutput.t161 gnd 0.052293f
C4561 CSoutput.t162 gnd 0.052293f
C4562 CSoutput.n288 gnd 0.404869f
C4563 CSoutput.t150 gnd 0.052293f
C4564 CSoutput.t96 gnd 0.052293f
C4565 CSoutput.n289 gnd 0.404147f
C4566 CSoutput.n290 gnd 0.410209f
C4567 CSoutput.t122 gnd 0.052293f
C4568 CSoutput.t102 gnd 0.052293f
C4569 CSoutput.n291 gnd 0.404147f
C4570 CSoutput.n292 gnd 0.202134f
C4571 CSoutput.t123 gnd 0.052293f
C4572 CSoutput.t148 gnd 0.052293f
C4573 CSoutput.n293 gnd 0.404147f
C4574 CSoutput.n294 gnd 0.202134f
C4575 CSoutput.t130 gnd 0.052293f
C4576 CSoutput.t165 gnd 0.052293f
C4577 CSoutput.n295 gnd 0.404147f
C4578 CSoutput.n296 gnd 0.202134f
C4579 CSoutput.t146 gnd 0.052293f
C4580 CSoutput.t140 gnd 0.052293f
C4581 CSoutput.n297 gnd 0.404146f
C4582 CSoutput.n298 gnd 0.301434f
C4583 CSoutput.n299 gnd 0.424859f
C4584 CSoutput.n300 gnd 11.3007f
C4585 CSoutput.t39 gnd 0.045756f
C4586 CSoutput.t92 gnd 0.045756f
C4587 CSoutput.n301 gnd 0.405672f
C4588 CSoutput.t33 gnd 0.045756f
C4589 CSoutput.t38 gnd 0.045756f
C4590 CSoutput.n302 gnd 0.404319f
C4591 CSoutput.n303 gnd 0.37675f
C4592 CSoutput.t23 gnd 0.045756f
C4593 CSoutput.t42 gnd 0.045756f
C4594 CSoutput.n304 gnd 0.404319f
C4595 CSoutput.n305 gnd 0.18572f
C4596 CSoutput.t57 gnd 0.045756f
C4597 CSoutput.t34 gnd 0.045756f
C4598 CSoutput.n306 gnd 0.404319f
C4599 CSoutput.n307 gnd 0.18572f
C4600 CSoutput.t41 gnd 0.045756f
C4601 CSoutput.t83 gnd 0.045756f
C4602 CSoutput.n308 gnd 0.404319f
C4603 CSoutput.n309 gnd 0.18572f
C4604 CSoutput.t53 gnd 0.045756f
C4605 CSoutput.t63 gnd 0.045756f
C4606 CSoutput.n310 gnd 0.404319f
C4607 CSoutput.n311 gnd 0.18572f
C4608 CSoutput.t18 gnd 0.045756f
C4609 CSoutput.t43 gnd 0.045756f
C4610 CSoutput.n312 gnd 0.404319f
C4611 CSoutput.n313 gnd 0.18572f
C4612 CSoutput.t7 gnd 0.045756f
C4613 CSoutput.t30 gnd 0.045756f
C4614 CSoutput.n314 gnd 0.404319f
C4615 CSoutput.n315 gnd 0.34255f
C4616 CSoutput.t88 gnd 0.045756f
C4617 CSoutput.t0 gnd 0.045756f
C4618 CSoutput.n316 gnd 0.405672f
C4619 CSoutput.t11 gnd 0.045756f
C4620 CSoutput.t81 gnd 0.045756f
C4621 CSoutput.n317 gnd 0.404319f
C4622 CSoutput.n318 gnd 0.37675f
C4623 CSoutput.t2 gnd 0.045756f
C4624 CSoutput.t74 gnd 0.045756f
C4625 CSoutput.n319 gnd 0.404319f
C4626 CSoutput.n320 gnd 0.18572f
C4627 CSoutput.t82 gnd 0.045756f
C4628 CSoutput.t1 gnd 0.045756f
C4629 CSoutput.n321 gnd 0.404319f
C4630 CSoutput.n322 gnd 0.18572f
C4631 CSoutput.t65 gnd 0.045756f
C4632 CSoutput.t46 gnd 0.045756f
C4633 CSoutput.n323 gnd 0.404319f
C4634 CSoutput.n324 gnd 0.18572f
C4635 CSoutput.t3 gnd 0.045756f
C4636 CSoutput.t67 gnd 0.045756f
C4637 CSoutput.n325 gnd 0.404319f
C4638 CSoutput.n326 gnd 0.18572f
C4639 CSoutput.t48 gnd 0.045756f
C4640 CSoutput.t54 gnd 0.045756f
C4641 CSoutput.n327 gnd 0.404319f
C4642 CSoutput.n328 gnd 0.18572f
C4643 CSoutput.t66 gnd 0.045756f
C4644 CSoutput.t47 gnd 0.045756f
C4645 CSoutput.n329 gnd 0.404319f
C4646 CSoutput.n330 gnd 0.281963f
C4647 CSoutput.n331 gnd 0.355642f
C4648 CSoutput.t12 gnd 0.045756f
C4649 CSoutput.t84 gnd 0.045756f
C4650 CSoutput.n332 gnd 0.405672f
C4651 CSoutput.t31 gnd 0.045756f
C4652 CSoutput.t35 gnd 0.045756f
C4653 CSoutput.n333 gnd 0.404319f
C4654 CSoutput.n334 gnd 0.37675f
C4655 CSoutput.t4 gnd 0.045756f
C4656 CSoutput.t69 gnd 0.045756f
C4657 CSoutput.n335 gnd 0.404319f
C4658 CSoutput.n336 gnd 0.18572f
C4659 CSoutput.t40 gnd 0.045756f
C4660 CSoutput.t13 gnd 0.045756f
C4661 CSoutput.n337 gnd 0.404319f
C4662 CSoutput.n338 gnd 0.18572f
C4663 CSoutput.t21 gnd 0.045756f
C4664 CSoutput.t95 gnd 0.045756f
C4665 CSoutput.n339 gnd 0.404319f
C4666 CSoutput.n340 gnd 0.18572f
C4667 CSoutput.t22 gnd 0.045756f
C4668 CSoutput.t26 gnd 0.045756f
C4669 CSoutput.n341 gnd 0.404319f
C4670 CSoutput.n342 gnd 0.18572f
C4671 CSoutput.t10 gnd 0.045756f
C4672 CSoutput.t80 gnd 0.045756f
C4673 CSoutput.n343 gnd 0.404319f
C4674 CSoutput.n344 gnd 0.18572f
C4675 CSoutput.t29 gnd 0.045756f
C4676 CSoutput.t19 gnd 0.045756f
C4677 CSoutput.n345 gnd 0.404319f
C4678 CSoutput.n346 gnd 0.281963f
C4679 CSoutput.n347 gnd 0.381904f
C4680 CSoutput.n348 gnd 11.458f
C4681 CSoutput.t25 gnd 0.045756f
C4682 CSoutput.t68 gnd 0.045756f
C4683 CSoutput.n349 gnd 0.405672f
C4684 CSoutput.t64 gnd 0.045756f
C4685 CSoutput.t45 gnd 0.045756f
C4686 CSoutput.n350 gnd 0.404319f
C4687 CSoutput.n351 gnd 0.37675f
C4688 CSoutput.t71 gnd 0.045756f
C4689 CSoutput.t36 gnd 0.045756f
C4690 CSoutput.n352 gnd 0.404319f
C4691 CSoutput.n353 gnd 0.18572f
C4692 CSoutput.t55 gnd 0.045756f
C4693 CSoutput.t86 gnd 0.045756f
C4694 CSoutput.n354 gnd 0.404319f
C4695 CSoutput.n355 gnd 0.18572f
C4696 CSoutput.t20 gnd 0.045756f
C4697 CSoutput.t70 gnd 0.045756f
C4698 CSoutput.n356 gnd 0.404319f
C4699 CSoutput.n357 gnd 0.18572f
C4700 CSoutput.t9 gnd 0.045756f
C4701 CSoutput.t76 gnd 0.045756f
C4702 CSoutput.n358 gnd 0.404319f
C4703 CSoutput.n359 gnd 0.18572f
C4704 CSoutput.t75 gnd 0.045756f
C4705 CSoutput.t32 gnd 0.045756f
C4706 CSoutput.n360 gnd 0.404319f
C4707 CSoutput.n361 gnd 0.18572f
C4708 CSoutput.t51 gnd 0.045756f
C4709 CSoutput.t28 gnd 0.045756f
C4710 CSoutput.n362 gnd 0.404319f
C4711 CSoutput.n363 gnd 0.34255f
C4712 CSoutput.t15 gnd 0.045756f
C4713 CSoutput.t8 gnd 0.045756f
C4714 CSoutput.n364 gnd 0.405672f
C4715 CSoutput.t5 gnd 0.045756f
C4716 CSoutput.t93 gnd 0.045756f
C4717 CSoutput.n365 gnd 0.404319f
C4718 CSoutput.n366 gnd 0.37675f
C4719 CSoutput.t94 gnd 0.045756f
C4720 CSoutput.t16 gnd 0.045756f
C4721 CSoutput.n367 gnd 0.404319f
C4722 CSoutput.n368 gnd 0.18572f
C4723 CSoutput.t17 gnd 0.045756f
C4724 CSoutput.t59 gnd 0.045756f
C4725 CSoutput.n369 gnd 0.404319f
C4726 CSoutput.n370 gnd 0.18572f
C4727 CSoutput.t60 gnd 0.045756f
C4728 CSoutput.t87 gnd 0.045756f
C4729 CSoutput.n371 gnd 0.404319f
C4730 CSoutput.n372 gnd 0.18572f
C4731 CSoutput.t90 gnd 0.045756f
C4732 CSoutput.t79 gnd 0.045756f
C4733 CSoutput.n373 gnd 0.404319f
C4734 CSoutput.n374 gnd 0.18572f
C4735 CSoutput.t73 gnd 0.045756f
C4736 CSoutput.t61 gnd 0.045756f
C4737 CSoutput.n375 gnd 0.404319f
C4738 CSoutput.n376 gnd 0.18572f
C4739 CSoutput.t62 gnd 0.045756f
C4740 CSoutput.t91 gnd 0.045756f
C4741 CSoutput.n377 gnd 0.404319f
C4742 CSoutput.n378 gnd 0.281963f
C4743 CSoutput.n379 gnd 0.355642f
C4744 CSoutput.t52 gnd 0.045756f
C4745 CSoutput.t77 gnd 0.045756f
C4746 CSoutput.n380 gnd 0.405672f
C4747 CSoutput.t24 gnd 0.045756f
C4748 CSoutput.t37 gnd 0.045756f
C4749 CSoutput.n381 gnd 0.404319f
C4750 CSoutput.n382 gnd 0.37675f
C4751 CSoutput.t44 gnd 0.045756f
C4752 CSoutput.t58 gnd 0.045756f
C4753 CSoutput.n383 gnd 0.404319f
C4754 CSoutput.n384 gnd 0.18572f
C4755 CSoutput.t78 gnd 0.045756f
C4756 CSoutput.t49 gnd 0.045756f
C4757 CSoutput.n385 gnd 0.404319f
C4758 CSoutput.n386 gnd 0.18572f
C4759 CSoutput.t56 gnd 0.045756f
C4760 CSoutput.t89 gnd 0.045756f
C4761 CSoutput.n387 gnd 0.404319f
C4762 CSoutput.n388 gnd 0.18572f
C4763 CSoutput.t6 gnd 0.045756f
C4764 CSoutput.t27 gnd 0.045756f
C4765 CSoutput.n389 gnd 0.404319f
C4766 CSoutput.n390 gnd 0.18572f
C4767 CSoutput.t50 gnd 0.045756f
C4768 CSoutput.t72 gnd 0.045756f
C4769 CSoutput.n391 gnd 0.404319f
C4770 CSoutput.n392 gnd 0.18572f
C4771 CSoutput.t85 gnd 0.045756f
C4772 CSoutput.t14 gnd 0.045756f
C4773 CSoutput.n393 gnd 0.404319f
C4774 CSoutput.n394 gnd 0.281963f
C4775 CSoutput.n395 gnd 0.381904f
C4776 CSoutput.n396 gnd 6.661911f
C4777 CSoutput.n397 gnd 12.6678f
C4778 commonsourceibias.n0 gnd 0.012624f
C4779 commonsourceibias.t120 gnd 0.191163f
C4780 commonsourceibias.t67 gnd 0.176757f
C4781 commonsourceibias.n1 gnd 0.00769f
C4782 commonsourceibias.n2 gnd 0.009461f
C4783 commonsourceibias.t126 gnd 0.176757f
C4784 commonsourceibias.n3 gnd 0.009597f
C4785 commonsourceibias.n4 gnd 0.009461f
C4786 commonsourceibias.t121 gnd 0.176757f
C4787 commonsourceibias.n5 gnd 0.070526f
C4788 commonsourceibias.t136 gnd 0.176757f
C4789 commonsourceibias.n6 gnd 0.007653f
C4790 commonsourceibias.n7 gnd 0.009461f
C4791 commonsourceibias.t117 gnd 0.176757f
C4792 commonsourceibias.n8 gnd 0.009134f
C4793 commonsourceibias.n9 gnd 0.009461f
C4794 commonsourceibias.t102 gnd 0.176757f
C4795 commonsourceibias.n10 gnd 0.070526f
C4796 commonsourceibias.t125 gnd 0.176757f
C4797 commonsourceibias.n11 gnd 0.007641f
C4798 commonsourceibias.n12 gnd 0.012624f
C4799 commonsourceibias.t12 gnd 0.191163f
C4800 commonsourceibias.t48 gnd 0.176757f
C4801 commonsourceibias.n13 gnd 0.00769f
C4802 commonsourceibias.n14 gnd 0.009461f
C4803 commonsourceibias.t4 gnd 0.176757f
C4804 commonsourceibias.n15 gnd 0.009597f
C4805 commonsourceibias.n16 gnd 0.009461f
C4806 commonsourceibias.t10 gnd 0.176757f
C4807 commonsourceibias.n17 gnd 0.070526f
C4808 commonsourceibias.t58 gnd 0.176757f
C4809 commonsourceibias.n18 gnd 0.007653f
C4810 commonsourceibias.n19 gnd 0.009461f
C4811 commonsourceibias.t16 gnd 0.176757f
C4812 commonsourceibias.n20 gnd 0.009134f
C4813 commonsourceibias.n21 gnd 0.009461f
C4814 commonsourceibias.t28 gnd 0.176757f
C4815 commonsourceibias.n22 gnd 0.070526f
C4816 commonsourceibias.t6 gnd 0.176757f
C4817 commonsourceibias.n23 gnd 0.007641f
C4818 commonsourceibias.n24 gnd 0.009461f
C4819 commonsourceibias.t14 gnd 0.176757f
C4820 commonsourceibias.t44 gnd 0.176757f
C4821 commonsourceibias.n25 gnd 0.070526f
C4822 commonsourceibias.n26 gnd 0.009461f
C4823 commonsourceibias.t24 gnd 0.176757f
C4824 commonsourceibias.n27 gnd 0.070526f
C4825 commonsourceibias.n28 gnd 0.009461f
C4826 commonsourceibias.t30 gnd 0.176757f
C4827 commonsourceibias.n29 gnd 0.070526f
C4828 commonsourceibias.n30 gnd 0.009461f
C4829 commonsourceibias.t54 gnd 0.176757f
C4830 commonsourceibias.n31 gnd 0.010754f
C4831 commonsourceibias.n32 gnd 0.009461f
C4832 commonsourceibias.t18 gnd 0.176757f
C4833 commonsourceibias.n33 gnd 0.012717f
C4834 commonsourceibias.t0 gnd 0.196904f
C4835 commonsourceibias.t50 gnd 0.176757f
C4836 commonsourceibias.n34 gnd 0.078584f
C4837 commonsourceibias.n35 gnd 0.084191f
C4838 commonsourceibias.n36 gnd 0.04027f
C4839 commonsourceibias.n37 gnd 0.009461f
C4840 commonsourceibias.n38 gnd 0.00769f
C4841 commonsourceibias.n39 gnd 0.013037f
C4842 commonsourceibias.n40 gnd 0.070526f
C4843 commonsourceibias.n41 gnd 0.013093f
C4844 commonsourceibias.n42 gnd 0.009461f
C4845 commonsourceibias.n43 gnd 0.009461f
C4846 commonsourceibias.n44 gnd 0.009461f
C4847 commonsourceibias.n45 gnd 0.009597f
C4848 commonsourceibias.n46 gnd 0.070526f
C4849 commonsourceibias.n47 gnd 0.011661f
C4850 commonsourceibias.n48 gnd 0.0129f
C4851 commonsourceibias.n49 gnd 0.009461f
C4852 commonsourceibias.n50 gnd 0.009461f
C4853 commonsourceibias.n51 gnd 0.012816f
C4854 commonsourceibias.n52 gnd 0.007653f
C4855 commonsourceibias.n53 gnd 0.012975f
C4856 commonsourceibias.n54 gnd 0.009461f
C4857 commonsourceibias.n55 gnd 0.009461f
C4858 commonsourceibias.n56 gnd 0.013054f
C4859 commonsourceibias.n57 gnd 0.011256f
C4860 commonsourceibias.n58 gnd 0.009134f
C4861 commonsourceibias.n59 gnd 0.009461f
C4862 commonsourceibias.n60 gnd 0.009461f
C4863 commonsourceibias.n61 gnd 0.011572f
C4864 commonsourceibias.n62 gnd 0.012989f
C4865 commonsourceibias.n63 gnd 0.070526f
C4866 commonsourceibias.n64 gnd 0.012901f
C4867 commonsourceibias.n65 gnd 0.009461f
C4868 commonsourceibias.n66 gnd 0.009461f
C4869 commonsourceibias.n67 gnd 0.009461f
C4870 commonsourceibias.n68 gnd 0.012901f
C4871 commonsourceibias.n69 gnd 0.070526f
C4872 commonsourceibias.n70 gnd 0.012989f
C4873 commonsourceibias.n71 gnd 0.011572f
C4874 commonsourceibias.n72 gnd 0.009461f
C4875 commonsourceibias.n73 gnd 0.009461f
C4876 commonsourceibias.n74 gnd 0.009461f
C4877 commonsourceibias.n75 gnd 0.011256f
C4878 commonsourceibias.n76 gnd 0.013054f
C4879 commonsourceibias.n77 gnd 0.070526f
C4880 commonsourceibias.n78 gnd 0.012975f
C4881 commonsourceibias.n79 gnd 0.009461f
C4882 commonsourceibias.n80 gnd 0.009461f
C4883 commonsourceibias.n81 gnd 0.009461f
C4884 commonsourceibias.n82 gnd 0.012816f
C4885 commonsourceibias.n83 gnd 0.070526f
C4886 commonsourceibias.n84 gnd 0.0129f
C4887 commonsourceibias.n85 gnd 0.011661f
C4888 commonsourceibias.n86 gnd 0.009461f
C4889 commonsourceibias.n87 gnd 0.009461f
C4890 commonsourceibias.n88 gnd 0.009461f
C4891 commonsourceibias.n89 gnd 0.010754f
C4892 commonsourceibias.n90 gnd 0.013093f
C4893 commonsourceibias.n91 gnd 0.070526f
C4894 commonsourceibias.n92 gnd 0.013037f
C4895 commonsourceibias.n93 gnd 0.009461f
C4896 commonsourceibias.n94 gnd 0.009461f
C4897 commonsourceibias.n95 gnd 0.009461f
C4898 commonsourceibias.n96 gnd 0.012717f
C4899 commonsourceibias.n97 gnd 0.070526f
C4900 commonsourceibias.n98 gnd 0.012748f
C4901 commonsourceibias.n99 gnd 0.085044f
C4902 commonsourceibias.n100 gnd 0.095092f
C4903 commonsourceibias.t13 gnd 0.020415f
C4904 commonsourceibias.t49 gnd 0.020415f
C4905 commonsourceibias.n101 gnd 0.180398f
C4906 commonsourceibias.n102 gnd 0.156264f
C4907 commonsourceibias.t5 gnd 0.020415f
C4908 commonsourceibias.t11 gnd 0.020415f
C4909 commonsourceibias.n103 gnd 0.180398f
C4910 commonsourceibias.n104 gnd 0.082864f
C4911 commonsourceibias.t59 gnd 0.020415f
C4912 commonsourceibias.t17 gnd 0.020415f
C4913 commonsourceibias.n105 gnd 0.180398f
C4914 commonsourceibias.n106 gnd 0.082864f
C4915 commonsourceibias.t29 gnd 0.020415f
C4916 commonsourceibias.t7 gnd 0.020415f
C4917 commonsourceibias.n107 gnd 0.180398f
C4918 commonsourceibias.n108 gnd 0.069229f
C4919 commonsourceibias.t51 gnd 0.020415f
C4920 commonsourceibias.t1 gnd 0.020415f
C4921 commonsourceibias.n109 gnd 0.181002f
C4922 commonsourceibias.t55 gnd 0.020415f
C4923 commonsourceibias.t19 gnd 0.020415f
C4924 commonsourceibias.n110 gnd 0.180398f
C4925 commonsourceibias.n111 gnd 0.168097f
C4926 commonsourceibias.t25 gnd 0.020415f
C4927 commonsourceibias.t31 gnd 0.020415f
C4928 commonsourceibias.n112 gnd 0.180398f
C4929 commonsourceibias.n113 gnd 0.082864f
C4930 commonsourceibias.t15 gnd 0.020415f
C4931 commonsourceibias.t45 gnd 0.020415f
C4932 commonsourceibias.n114 gnd 0.180398f
C4933 commonsourceibias.n115 gnd 0.069229f
C4934 commonsourceibias.n116 gnd 0.083829f
C4935 commonsourceibias.n117 gnd 0.009461f
C4936 commonsourceibias.t118 gnd 0.176757f
C4937 commonsourceibias.t76 gnd 0.176757f
C4938 commonsourceibias.n118 gnd 0.070526f
C4939 commonsourceibias.n119 gnd 0.009461f
C4940 commonsourceibias.t106 gnd 0.176757f
C4941 commonsourceibias.n120 gnd 0.070526f
C4942 commonsourceibias.n121 gnd 0.009461f
C4943 commonsourceibias.t96 gnd 0.176757f
C4944 commonsourceibias.n122 gnd 0.070526f
C4945 commonsourceibias.n123 gnd 0.009461f
C4946 commonsourceibias.t141 gnd 0.176757f
C4947 commonsourceibias.n124 gnd 0.010754f
C4948 commonsourceibias.n125 gnd 0.009461f
C4949 commonsourceibias.t116 gnd 0.176757f
C4950 commonsourceibias.n126 gnd 0.012717f
C4951 commonsourceibias.t129 gnd 0.196904f
C4952 commonsourceibias.t152 gnd 0.176757f
C4953 commonsourceibias.n127 gnd 0.078584f
C4954 commonsourceibias.n128 gnd 0.084191f
C4955 commonsourceibias.n129 gnd 0.04027f
C4956 commonsourceibias.n130 gnd 0.009461f
C4957 commonsourceibias.n131 gnd 0.00769f
C4958 commonsourceibias.n132 gnd 0.013037f
C4959 commonsourceibias.n133 gnd 0.070526f
C4960 commonsourceibias.n134 gnd 0.013093f
C4961 commonsourceibias.n135 gnd 0.009461f
C4962 commonsourceibias.n136 gnd 0.009461f
C4963 commonsourceibias.n137 gnd 0.009461f
C4964 commonsourceibias.n138 gnd 0.009597f
C4965 commonsourceibias.n139 gnd 0.070526f
C4966 commonsourceibias.n140 gnd 0.011661f
C4967 commonsourceibias.n141 gnd 0.0129f
C4968 commonsourceibias.n142 gnd 0.009461f
C4969 commonsourceibias.n143 gnd 0.009461f
C4970 commonsourceibias.n144 gnd 0.012816f
C4971 commonsourceibias.n145 gnd 0.007653f
C4972 commonsourceibias.n146 gnd 0.012975f
C4973 commonsourceibias.n147 gnd 0.009461f
C4974 commonsourceibias.n148 gnd 0.009461f
C4975 commonsourceibias.n149 gnd 0.013054f
C4976 commonsourceibias.n150 gnd 0.011256f
C4977 commonsourceibias.n151 gnd 0.009134f
C4978 commonsourceibias.n152 gnd 0.009461f
C4979 commonsourceibias.n153 gnd 0.009461f
C4980 commonsourceibias.n154 gnd 0.011572f
C4981 commonsourceibias.n155 gnd 0.012989f
C4982 commonsourceibias.n156 gnd 0.070526f
C4983 commonsourceibias.n157 gnd 0.012901f
C4984 commonsourceibias.n158 gnd 0.009415f
C4985 commonsourceibias.n159 gnd 0.06839f
C4986 commonsourceibias.n160 gnd 0.009415f
C4987 commonsourceibias.n161 gnd 0.012901f
C4988 commonsourceibias.n162 gnd 0.070526f
C4989 commonsourceibias.n163 gnd 0.012989f
C4990 commonsourceibias.n164 gnd 0.011572f
C4991 commonsourceibias.n165 gnd 0.009461f
C4992 commonsourceibias.n166 gnd 0.009461f
C4993 commonsourceibias.n167 gnd 0.009461f
C4994 commonsourceibias.n168 gnd 0.011256f
C4995 commonsourceibias.n169 gnd 0.013054f
C4996 commonsourceibias.n170 gnd 0.070526f
C4997 commonsourceibias.n171 gnd 0.012975f
C4998 commonsourceibias.n172 gnd 0.009461f
C4999 commonsourceibias.n173 gnd 0.009461f
C5000 commonsourceibias.n174 gnd 0.009461f
C5001 commonsourceibias.n175 gnd 0.012816f
C5002 commonsourceibias.n176 gnd 0.070526f
C5003 commonsourceibias.n177 gnd 0.0129f
C5004 commonsourceibias.n178 gnd 0.011661f
C5005 commonsourceibias.n179 gnd 0.009461f
C5006 commonsourceibias.n180 gnd 0.009461f
C5007 commonsourceibias.n181 gnd 0.009461f
C5008 commonsourceibias.n182 gnd 0.010754f
C5009 commonsourceibias.n183 gnd 0.013093f
C5010 commonsourceibias.n184 gnd 0.070526f
C5011 commonsourceibias.n185 gnd 0.013037f
C5012 commonsourceibias.n186 gnd 0.009461f
C5013 commonsourceibias.n187 gnd 0.009461f
C5014 commonsourceibias.n188 gnd 0.009461f
C5015 commonsourceibias.n189 gnd 0.012717f
C5016 commonsourceibias.n190 gnd 0.070526f
C5017 commonsourceibias.n191 gnd 0.012748f
C5018 commonsourceibias.n192 gnd 0.085044f
C5019 commonsourceibias.n193 gnd 0.056182f
C5020 commonsourceibias.n194 gnd 0.012624f
C5021 commonsourceibias.t71 gnd 0.191163f
C5022 commonsourceibias.t159 gnd 0.176757f
C5023 commonsourceibias.n195 gnd 0.00769f
C5024 commonsourceibias.n196 gnd 0.009461f
C5025 commonsourceibias.t148 gnd 0.176757f
C5026 commonsourceibias.n197 gnd 0.009597f
C5027 commonsourceibias.n198 gnd 0.009461f
C5028 commonsourceibias.t78 gnd 0.176757f
C5029 commonsourceibias.n199 gnd 0.070526f
C5030 commonsourceibias.t157 gnd 0.176757f
C5031 commonsourceibias.n200 gnd 0.007653f
C5032 commonsourceibias.n201 gnd 0.009461f
C5033 commonsourceibias.t85 gnd 0.176757f
C5034 commonsourceibias.n202 gnd 0.009134f
C5035 commonsourceibias.n203 gnd 0.009461f
C5036 commonsourceibias.t77 gnd 0.176757f
C5037 commonsourceibias.n204 gnd 0.070526f
C5038 commonsourceibias.t158 gnd 0.176757f
C5039 commonsourceibias.n205 gnd 0.007641f
C5040 commonsourceibias.n206 gnd 0.009461f
C5041 commonsourceibias.t94 gnd 0.176757f
C5042 commonsourceibias.t113 gnd 0.176757f
C5043 commonsourceibias.n207 gnd 0.070526f
C5044 commonsourceibias.n208 gnd 0.009461f
C5045 commonsourceibias.t156 gnd 0.176757f
C5046 commonsourceibias.n209 gnd 0.070526f
C5047 commonsourceibias.n210 gnd 0.009461f
C5048 commonsourceibias.t92 gnd 0.176757f
C5049 commonsourceibias.n211 gnd 0.070526f
C5050 commonsourceibias.n212 gnd 0.009461f
C5051 commonsourceibias.t111 gnd 0.176757f
C5052 commonsourceibias.n213 gnd 0.010754f
C5053 commonsourceibias.n214 gnd 0.009461f
C5054 commonsourceibias.t105 gnd 0.176757f
C5055 commonsourceibias.n215 gnd 0.012717f
C5056 commonsourceibias.t112 gnd 0.196904f
C5057 commonsourceibias.t93 gnd 0.176757f
C5058 commonsourceibias.n216 gnd 0.078584f
C5059 commonsourceibias.n217 gnd 0.084191f
C5060 commonsourceibias.n218 gnd 0.04027f
C5061 commonsourceibias.n219 gnd 0.009461f
C5062 commonsourceibias.n220 gnd 0.00769f
C5063 commonsourceibias.n221 gnd 0.013037f
C5064 commonsourceibias.n222 gnd 0.070526f
C5065 commonsourceibias.n223 gnd 0.013093f
C5066 commonsourceibias.n224 gnd 0.009461f
C5067 commonsourceibias.n225 gnd 0.009461f
C5068 commonsourceibias.n226 gnd 0.009461f
C5069 commonsourceibias.n227 gnd 0.009597f
C5070 commonsourceibias.n228 gnd 0.070526f
C5071 commonsourceibias.n229 gnd 0.011661f
C5072 commonsourceibias.n230 gnd 0.0129f
C5073 commonsourceibias.n231 gnd 0.009461f
C5074 commonsourceibias.n232 gnd 0.009461f
C5075 commonsourceibias.n233 gnd 0.012816f
C5076 commonsourceibias.n234 gnd 0.007653f
C5077 commonsourceibias.n235 gnd 0.012975f
C5078 commonsourceibias.n236 gnd 0.009461f
C5079 commonsourceibias.n237 gnd 0.009461f
C5080 commonsourceibias.n238 gnd 0.013054f
C5081 commonsourceibias.n239 gnd 0.011256f
C5082 commonsourceibias.n240 gnd 0.009134f
C5083 commonsourceibias.n241 gnd 0.009461f
C5084 commonsourceibias.n242 gnd 0.009461f
C5085 commonsourceibias.n243 gnd 0.011572f
C5086 commonsourceibias.n244 gnd 0.012989f
C5087 commonsourceibias.n245 gnd 0.070526f
C5088 commonsourceibias.n246 gnd 0.012901f
C5089 commonsourceibias.n247 gnd 0.009461f
C5090 commonsourceibias.n248 gnd 0.009461f
C5091 commonsourceibias.n249 gnd 0.009461f
C5092 commonsourceibias.n250 gnd 0.012901f
C5093 commonsourceibias.n251 gnd 0.070526f
C5094 commonsourceibias.n252 gnd 0.012989f
C5095 commonsourceibias.n253 gnd 0.011572f
C5096 commonsourceibias.n254 gnd 0.009461f
C5097 commonsourceibias.n255 gnd 0.009461f
C5098 commonsourceibias.n256 gnd 0.009461f
C5099 commonsourceibias.n257 gnd 0.011256f
C5100 commonsourceibias.n258 gnd 0.013054f
C5101 commonsourceibias.n259 gnd 0.070526f
C5102 commonsourceibias.n260 gnd 0.012975f
C5103 commonsourceibias.n261 gnd 0.009461f
C5104 commonsourceibias.n262 gnd 0.009461f
C5105 commonsourceibias.n263 gnd 0.009461f
C5106 commonsourceibias.n264 gnd 0.012816f
C5107 commonsourceibias.n265 gnd 0.070526f
C5108 commonsourceibias.n266 gnd 0.0129f
C5109 commonsourceibias.n267 gnd 0.011661f
C5110 commonsourceibias.n268 gnd 0.009461f
C5111 commonsourceibias.n269 gnd 0.009461f
C5112 commonsourceibias.n270 gnd 0.009461f
C5113 commonsourceibias.n271 gnd 0.010754f
C5114 commonsourceibias.n272 gnd 0.013093f
C5115 commonsourceibias.n273 gnd 0.070526f
C5116 commonsourceibias.n274 gnd 0.013037f
C5117 commonsourceibias.n275 gnd 0.009461f
C5118 commonsourceibias.n276 gnd 0.009461f
C5119 commonsourceibias.n277 gnd 0.009461f
C5120 commonsourceibias.n278 gnd 0.012717f
C5121 commonsourceibias.n279 gnd 0.070526f
C5122 commonsourceibias.n280 gnd 0.012748f
C5123 commonsourceibias.n281 gnd 0.085044f
C5124 commonsourceibias.n282 gnd 0.030348f
C5125 commonsourceibias.n283 gnd 0.15151f
C5126 commonsourceibias.n284 gnd 0.012624f
C5127 commonsourceibias.t75 gnd 0.176757f
C5128 commonsourceibias.n285 gnd 0.00769f
C5129 commonsourceibias.n286 gnd 0.009461f
C5130 commonsourceibias.t128 gnd 0.176757f
C5131 commonsourceibias.n287 gnd 0.009597f
C5132 commonsourceibias.n288 gnd 0.009461f
C5133 commonsourceibias.t124 gnd 0.176757f
C5134 commonsourceibias.n289 gnd 0.070526f
C5135 commonsourceibias.t155 gnd 0.176757f
C5136 commonsourceibias.n290 gnd 0.007653f
C5137 commonsourceibias.n291 gnd 0.009461f
C5138 commonsourceibias.t90 gnd 0.176757f
C5139 commonsourceibias.n292 gnd 0.009134f
C5140 commonsourceibias.n293 gnd 0.009461f
C5141 commonsourceibias.t119 gnd 0.176757f
C5142 commonsourceibias.n294 gnd 0.070526f
C5143 commonsourceibias.t146 gnd 0.176757f
C5144 commonsourceibias.n295 gnd 0.007641f
C5145 commonsourceibias.n296 gnd 0.009461f
C5146 commonsourceibias.t138 gnd 0.176757f
C5147 commonsourceibias.t64 gnd 0.176757f
C5148 commonsourceibias.n297 gnd 0.070526f
C5149 commonsourceibias.n298 gnd 0.009461f
C5150 commonsourceibias.t137 gnd 0.176757f
C5151 commonsourceibias.n299 gnd 0.070526f
C5152 commonsourceibias.n300 gnd 0.009461f
C5153 commonsourceibias.t133 gnd 0.176757f
C5154 commonsourceibias.n301 gnd 0.070526f
C5155 commonsourceibias.n302 gnd 0.009461f
C5156 commonsourceibias.t149 gnd 0.176757f
C5157 commonsourceibias.n303 gnd 0.010754f
C5158 commonsourceibias.n304 gnd 0.009461f
C5159 commonsourceibias.t79 gnd 0.176757f
C5160 commonsourceibias.n305 gnd 0.012717f
C5161 commonsourceibias.t140 gnd 0.196904f
C5162 commonsourceibias.t130 gnd 0.176757f
C5163 commonsourceibias.n306 gnd 0.078584f
C5164 commonsourceibias.n307 gnd 0.084191f
C5165 commonsourceibias.n308 gnd 0.04027f
C5166 commonsourceibias.n309 gnd 0.009461f
C5167 commonsourceibias.n310 gnd 0.00769f
C5168 commonsourceibias.n311 gnd 0.013037f
C5169 commonsourceibias.n312 gnd 0.070526f
C5170 commonsourceibias.n313 gnd 0.013093f
C5171 commonsourceibias.n314 gnd 0.009461f
C5172 commonsourceibias.n315 gnd 0.009461f
C5173 commonsourceibias.n316 gnd 0.009461f
C5174 commonsourceibias.n317 gnd 0.009597f
C5175 commonsourceibias.n318 gnd 0.070526f
C5176 commonsourceibias.n319 gnd 0.011661f
C5177 commonsourceibias.n320 gnd 0.0129f
C5178 commonsourceibias.n321 gnd 0.009461f
C5179 commonsourceibias.n322 gnd 0.009461f
C5180 commonsourceibias.n323 gnd 0.012816f
C5181 commonsourceibias.n324 gnd 0.007653f
C5182 commonsourceibias.n325 gnd 0.012975f
C5183 commonsourceibias.n326 gnd 0.009461f
C5184 commonsourceibias.n327 gnd 0.009461f
C5185 commonsourceibias.n328 gnd 0.013054f
C5186 commonsourceibias.n329 gnd 0.011256f
C5187 commonsourceibias.n330 gnd 0.009134f
C5188 commonsourceibias.n331 gnd 0.009461f
C5189 commonsourceibias.n332 gnd 0.009461f
C5190 commonsourceibias.n333 gnd 0.011572f
C5191 commonsourceibias.n334 gnd 0.012989f
C5192 commonsourceibias.n335 gnd 0.070526f
C5193 commonsourceibias.n336 gnd 0.012901f
C5194 commonsourceibias.n337 gnd 0.009461f
C5195 commonsourceibias.n338 gnd 0.009461f
C5196 commonsourceibias.n339 gnd 0.009461f
C5197 commonsourceibias.n340 gnd 0.012901f
C5198 commonsourceibias.n341 gnd 0.070526f
C5199 commonsourceibias.n342 gnd 0.012989f
C5200 commonsourceibias.n343 gnd 0.011572f
C5201 commonsourceibias.n344 gnd 0.009461f
C5202 commonsourceibias.n345 gnd 0.009461f
C5203 commonsourceibias.n346 gnd 0.009461f
C5204 commonsourceibias.n347 gnd 0.011256f
C5205 commonsourceibias.n348 gnd 0.013054f
C5206 commonsourceibias.n349 gnd 0.070526f
C5207 commonsourceibias.n350 gnd 0.012975f
C5208 commonsourceibias.n351 gnd 0.009461f
C5209 commonsourceibias.n352 gnd 0.009461f
C5210 commonsourceibias.n353 gnd 0.009461f
C5211 commonsourceibias.n354 gnd 0.012816f
C5212 commonsourceibias.n355 gnd 0.070526f
C5213 commonsourceibias.n356 gnd 0.0129f
C5214 commonsourceibias.n357 gnd 0.011661f
C5215 commonsourceibias.n358 gnd 0.009461f
C5216 commonsourceibias.n359 gnd 0.009461f
C5217 commonsourceibias.n360 gnd 0.009461f
C5218 commonsourceibias.n361 gnd 0.010754f
C5219 commonsourceibias.n362 gnd 0.013093f
C5220 commonsourceibias.n363 gnd 0.070526f
C5221 commonsourceibias.n364 gnd 0.013037f
C5222 commonsourceibias.n365 gnd 0.009461f
C5223 commonsourceibias.n366 gnd 0.009461f
C5224 commonsourceibias.n367 gnd 0.009461f
C5225 commonsourceibias.n368 gnd 0.012717f
C5226 commonsourceibias.n369 gnd 0.070526f
C5227 commonsourceibias.n370 gnd 0.012748f
C5228 commonsourceibias.t147 gnd 0.191163f
C5229 commonsourceibias.n371 gnd 0.085044f
C5230 commonsourceibias.n372 gnd 0.030348f
C5231 commonsourceibias.n373 gnd 0.449685f
C5232 commonsourceibias.n374 gnd 0.012624f
C5233 commonsourceibias.t91 gnd 0.191163f
C5234 commonsourceibias.t134 gnd 0.176757f
C5235 commonsourceibias.n375 gnd 0.00769f
C5236 commonsourceibias.n376 gnd 0.009461f
C5237 commonsourceibias.t114 gnd 0.176757f
C5238 commonsourceibias.n377 gnd 0.009597f
C5239 commonsourceibias.n378 gnd 0.009461f
C5240 commonsourceibias.t123 gnd 0.176757f
C5241 commonsourceibias.n379 gnd 0.007653f
C5242 commonsourceibias.n380 gnd 0.009461f
C5243 commonsourceibias.t88 gnd 0.176757f
C5244 commonsourceibias.n381 gnd 0.009134f
C5245 commonsourceibias.n382 gnd 0.009461f
C5246 commonsourceibias.t104 gnd 0.176757f
C5247 commonsourceibias.n383 gnd 0.007641f
C5248 commonsourceibias.n384 gnd 0.009461f
C5249 commonsourceibias.t89 gnd 0.176757f
C5250 commonsourceibias.t139 gnd 0.176757f
C5251 commonsourceibias.n385 gnd 0.070526f
C5252 commonsourceibias.n386 gnd 0.009461f
C5253 commonsourceibias.t83 gnd 0.176757f
C5254 commonsourceibias.n387 gnd 0.070526f
C5255 commonsourceibias.n388 gnd 0.009461f
C5256 commonsourceibias.t150 gnd 0.176757f
C5257 commonsourceibias.n389 gnd 0.070526f
C5258 commonsourceibias.n390 gnd 0.009461f
C5259 commonsourceibias.t127 gnd 0.176757f
C5260 commonsourceibias.n391 gnd 0.010754f
C5261 commonsourceibias.n392 gnd 0.009461f
C5262 commonsourceibias.t84 gnd 0.176757f
C5263 commonsourceibias.n393 gnd 0.012717f
C5264 commonsourceibias.t108 gnd 0.196904f
C5265 commonsourceibias.t131 gnd 0.176757f
C5266 commonsourceibias.n394 gnd 0.078584f
C5267 commonsourceibias.n395 gnd 0.084191f
C5268 commonsourceibias.n396 gnd 0.04027f
C5269 commonsourceibias.n397 gnd 0.009461f
C5270 commonsourceibias.n398 gnd 0.00769f
C5271 commonsourceibias.n399 gnd 0.013037f
C5272 commonsourceibias.n400 gnd 0.070526f
C5273 commonsourceibias.n401 gnd 0.013093f
C5274 commonsourceibias.n402 gnd 0.009461f
C5275 commonsourceibias.n403 gnd 0.009461f
C5276 commonsourceibias.n404 gnd 0.009461f
C5277 commonsourceibias.n405 gnd 0.009597f
C5278 commonsourceibias.n406 gnd 0.070526f
C5279 commonsourceibias.n407 gnd 0.011661f
C5280 commonsourceibias.n408 gnd 0.0129f
C5281 commonsourceibias.n409 gnd 0.009461f
C5282 commonsourceibias.n410 gnd 0.009461f
C5283 commonsourceibias.n411 gnd 0.012816f
C5284 commonsourceibias.n412 gnd 0.007653f
C5285 commonsourceibias.n413 gnd 0.012975f
C5286 commonsourceibias.n414 gnd 0.009461f
C5287 commonsourceibias.n415 gnd 0.009461f
C5288 commonsourceibias.n416 gnd 0.013054f
C5289 commonsourceibias.n417 gnd 0.011256f
C5290 commonsourceibias.n418 gnd 0.009134f
C5291 commonsourceibias.n419 gnd 0.009461f
C5292 commonsourceibias.n420 gnd 0.009461f
C5293 commonsourceibias.n421 gnd 0.011572f
C5294 commonsourceibias.n422 gnd 0.012989f
C5295 commonsourceibias.n423 gnd 0.070526f
C5296 commonsourceibias.n424 gnd 0.012901f
C5297 commonsourceibias.n425 gnd 0.009415f
C5298 commonsourceibias.t23 gnd 0.020415f
C5299 commonsourceibias.t63 gnd 0.020415f
C5300 commonsourceibias.n426 gnd 0.181002f
C5301 commonsourceibias.t41 gnd 0.020415f
C5302 commonsourceibias.t3 gnd 0.020415f
C5303 commonsourceibias.n427 gnd 0.180398f
C5304 commonsourceibias.n428 gnd 0.168097f
C5305 commonsourceibias.t53 gnd 0.020415f
C5306 commonsourceibias.t43 gnd 0.020415f
C5307 commonsourceibias.n429 gnd 0.180398f
C5308 commonsourceibias.n430 gnd 0.082864f
C5309 commonsourceibias.t57 gnd 0.020415f
C5310 commonsourceibias.t37 gnd 0.020415f
C5311 commonsourceibias.n431 gnd 0.180398f
C5312 commonsourceibias.n432 gnd 0.069229f
C5313 commonsourceibias.n433 gnd 0.012624f
C5314 commonsourceibias.t60 gnd 0.176757f
C5315 commonsourceibias.n434 gnd 0.00769f
C5316 commonsourceibias.n435 gnd 0.009461f
C5317 commonsourceibias.t20 gnd 0.176757f
C5318 commonsourceibias.n436 gnd 0.009597f
C5319 commonsourceibias.n437 gnd 0.009461f
C5320 commonsourceibias.t8 gnd 0.176757f
C5321 commonsourceibias.n438 gnd 0.007653f
C5322 commonsourceibias.n439 gnd 0.009461f
C5323 commonsourceibias.t38 gnd 0.176757f
C5324 commonsourceibias.n440 gnd 0.009134f
C5325 commonsourceibias.n441 gnd 0.009461f
C5326 commonsourceibias.t26 gnd 0.176757f
C5327 commonsourceibias.n442 gnd 0.007641f
C5328 commonsourceibias.n443 gnd 0.009461f
C5329 commonsourceibias.t36 gnd 0.176757f
C5330 commonsourceibias.t56 gnd 0.176757f
C5331 commonsourceibias.n444 gnd 0.070526f
C5332 commonsourceibias.n445 gnd 0.009461f
C5333 commonsourceibias.t42 gnd 0.176757f
C5334 commonsourceibias.n446 gnd 0.070526f
C5335 commonsourceibias.n447 gnd 0.009461f
C5336 commonsourceibias.t52 gnd 0.176757f
C5337 commonsourceibias.n448 gnd 0.070526f
C5338 commonsourceibias.n449 gnd 0.009461f
C5339 commonsourceibias.t2 gnd 0.176757f
C5340 commonsourceibias.n450 gnd 0.010754f
C5341 commonsourceibias.n451 gnd 0.009461f
C5342 commonsourceibias.t40 gnd 0.176757f
C5343 commonsourceibias.n452 gnd 0.012717f
C5344 commonsourceibias.t22 gnd 0.196904f
C5345 commonsourceibias.t62 gnd 0.176757f
C5346 commonsourceibias.n453 gnd 0.078584f
C5347 commonsourceibias.n454 gnd 0.084191f
C5348 commonsourceibias.n455 gnd 0.04027f
C5349 commonsourceibias.n456 gnd 0.009461f
C5350 commonsourceibias.n457 gnd 0.00769f
C5351 commonsourceibias.n458 gnd 0.013037f
C5352 commonsourceibias.n459 gnd 0.070526f
C5353 commonsourceibias.n460 gnd 0.013093f
C5354 commonsourceibias.n461 gnd 0.009461f
C5355 commonsourceibias.n462 gnd 0.009461f
C5356 commonsourceibias.n463 gnd 0.009461f
C5357 commonsourceibias.n464 gnd 0.009597f
C5358 commonsourceibias.n465 gnd 0.070526f
C5359 commonsourceibias.n466 gnd 0.011661f
C5360 commonsourceibias.n467 gnd 0.0129f
C5361 commonsourceibias.n468 gnd 0.009461f
C5362 commonsourceibias.n469 gnd 0.009461f
C5363 commonsourceibias.n470 gnd 0.012816f
C5364 commonsourceibias.n471 gnd 0.007653f
C5365 commonsourceibias.n472 gnd 0.012975f
C5366 commonsourceibias.n473 gnd 0.009461f
C5367 commonsourceibias.n474 gnd 0.009461f
C5368 commonsourceibias.n475 gnd 0.013054f
C5369 commonsourceibias.n476 gnd 0.011256f
C5370 commonsourceibias.n477 gnd 0.009134f
C5371 commonsourceibias.n478 gnd 0.009461f
C5372 commonsourceibias.n479 gnd 0.009461f
C5373 commonsourceibias.n480 gnd 0.011572f
C5374 commonsourceibias.n481 gnd 0.012989f
C5375 commonsourceibias.n482 gnd 0.070526f
C5376 commonsourceibias.n483 gnd 0.012901f
C5377 commonsourceibias.n484 gnd 0.009461f
C5378 commonsourceibias.n485 gnd 0.009461f
C5379 commonsourceibias.n486 gnd 0.009461f
C5380 commonsourceibias.n487 gnd 0.012901f
C5381 commonsourceibias.n488 gnd 0.070526f
C5382 commonsourceibias.n489 gnd 0.012989f
C5383 commonsourceibias.t46 gnd 0.176757f
C5384 commonsourceibias.n490 gnd 0.070526f
C5385 commonsourceibias.n491 gnd 0.011572f
C5386 commonsourceibias.n492 gnd 0.009461f
C5387 commonsourceibias.n493 gnd 0.009461f
C5388 commonsourceibias.n494 gnd 0.009461f
C5389 commonsourceibias.n495 gnd 0.011256f
C5390 commonsourceibias.n496 gnd 0.013054f
C5391 commonsourceibias.n497 gnd 0.070526f
C5392 commonsourceibias.n498 gnd 0.012975f
C5393 commonsourceibias.n499 gnd 0.009461f
C5394 commonsourceibias.n500 gnd 0.009461f
C5395 commonsourceibias.n501 gnd 0.009461f
C5396 commonsourceibias.n502 gnd 0.012816f
C5397 commonsourceibias.n503 gnd 0.070526f
C5398 commonsourceibias.n504 gnd 0.0129f
C5399 commonsourceibias.t32 gnd 0.176757f
C5400 commonsourceibias.n505 gnd 0.070526f
C5401 commonsourceibias.n506 gnd 0.011661f
C5402 commonsourceibias.n507 gnd 0.009461f
C5403 commonsourceibias.n508 gnd 0.009461f
C5404 commonsourceibias.n509 gnd 0.009461f
C5405 commonsourceibias.n510 gnd 0.010754f
C5406 commonsourceibias.n511 gnd 0.013093f
C5407 commonsourceibias.n512 gnd 0.070526f
C5408 commonsourceibias.n513 gnd 0.013037f
C5409 commonsourceibias.n514 gnd 0.009461f
C5410 commonsourceibias.n515 gnd 0.009461f
C5411 commonsourceibias.n516 gnd 0.009461f
C5412 commonsourceibias.n517 gnd 0.012717f
C5413 commonsourceibias.n518 gnd 0.070526f
C5414 commonsourceibias.n519 gnd 0.012748f
C5415 commonsourceibias.t34 gnd 0.191163f
C5416 commonsourceibias.n520 gnd 0.085044f
C5417 commonsourceibias.n521 gnd 0.095092f
C5418 commonsourceibias.t61 gnd 0.020415f
C5419 commonsourceibias.t35 gnd 0.020415f
C5420 commonsourceibias.n522 gnd 0.180398f
C5421 commonsourceibias.n523 gnd 0.156264f
C5422 commonsourceibias.t33 gnd 0.020415f
C5423 commonsourceibias.t21 gnd 0.020415f
C5424 commonsourceibias.n524 gnd 0.180398f
C5425 commonsourceibias.n525 gnd 0.082864f
C5426 commonsourceibias.t39 gnd 0.020415f
C5427 commonsourceibias.t9 gnd 0.020415f
C5428 commonsourceibias.n526 gnd 0.180398f
C5429 commonsourceibias.n527 gnd 0.082864f
C5430 commonsourceibias.t27 gnd 0.020415f
C5431 commonsourceibias.t47 gnd 0.020415f
C5432 commonsourceibias.n528 gnd 0.180398f
C5433 commonsourceibias.n529 gnd 0.069229f
C5434 commonsourceibias.n530 gnd 0.083829f
C5435 commonsourceibias.n531 gnd 0.06839f
C5436 commonsourceibias.n532 gnd 0.009415f
C5437 commonsourceibias.n533 gnd 0.012901f
C5438 commonsourceibias.n534 gnd 0.070526f
C5439 commonsourceibias.n535 gnd 0.012989f
C5440 commonsourceibias.t73 gnd 0.176757f
C5441 commonsourceibias.n536 gnd 0.070526f
C5442 commonsourceibias.n537 gnd 0.011572f
C5443 commonsourceibias.n538 gnd 0.009461f
C5444 commonsourceibias.n539 gnd 0.009461f
C5445 commonsourceibias.n540 gnd 0.009461f
C5446 commonsourceibias.n541 gnd 0.011256f
C5447 commonsourceibias.n542 gnd 0.013054f
C5448 commonsourceibias.n543 gnd 0.070526f
C5449 commonsourceibias.n544 gnd 0.012975f
C5450 commonsourceibias.n545 gnd 0.009461f
C5451 commonsourceibias.n546 gnd 0.009461f
C5452 commonsourceibias.n547 gnd 0.009461f
C5453 commonsourceibias.n548 gnd 0.012816f
C5454 commonsourceibias.n549 gnd 0.070526f
C5455 commonsourceibias.n550 gnd 0.0129f
C5456 commonsourceibias.t95 gnd 0.176757f
C5457 commonsourceibias.n551 gnd 0.070526f
C5458 commonsourceibias.n552 gnd 0.011661f
C5459 commonsourceibias.n553 gnd 0.009461f
C5460 commonsourceibias.n554 gnd 0.009461f
C5461 commonsourceibias.n555 gnd 0.009461f
C5462 commonsourceibias.n556 gnd 0.010754f
C5463 commonsourceibias.n557 gnd 0.013093f
C5464 commonsourceibias.n558 gnd 0.070526f
C5465 commonsourceibias.n559 gnd 0.013037f
C5466 commonsourceibias.n560 gnd 0.009461f
C5467 commonsourceibias.n561 gnd 0.009461f
C5468 commonsourceibias.n562 gnd 0.009461f
C5469 commonsourceibias.n563 gnd 0.012717f
C5470 commonsourceibias.n564 gnd 0.070526f
C5471 commonsourceibias.n565 gnd 0.012748f
C5472 commonsourceibias.n566 gnd 0.085044f
C5473 commonsourceibias.n567 gnd 0.056182f
C5474 commonsourceibias.n568 gnd 0.012624f
C5475 commonsourceibias.t144 gnd 0.176757f
C5476 commonsourceibias.n569 gnd 0.00769f
C5477 commonsourceibias.n570 gnd 0.009461f
C5478 commonsourceibias.t66 gnd 0.176757f
C5479 commonsourceibias.n571 gnd 0.009597f
C5480 commonsourceibias.n572 gnd 0.009461f
C5481 commonsourceibias.t143 gnd 0.176757f
C5482 commonsourceibias.n573 gnd 0.007653f
C5483 commonsourceibias.n574 gnd 0.009461f
C5484 commonsourceibias.t65 gnd 0.176757f
C5485 commonsourceibias.n575 gnd 0.009134f
C5486 commonsourceibias.n576 gnd 0.009461f
C5487 commonsourceibias.t142 gnd 0.176757f
C5488 commonsourceibias.n577 gnd 0.007641f
C5489 commonsourceibias.n578 gnd 0.009461f
C5490 commonsourceibias.t72 gnd 0.176757f
C5491 commonsourceibias.t99 gnd 0.176757f
C5492 commonsourceibias.n579 gnd 0.070526f
C5493 commonsourceibias.n580 gnd 0.009461f
C5494 commonsourceibias.t80 gnd 0.176757f
C5495 commonsourceibias.n581 gnd 0.070526f
C5496 commonsourceibias.n582 gnd 0.009461f
C5497 commonsourceibias.t69 gnd 0.176757f
C5498 commonsourceibias.n583 gnd 0.070526f
C5499 commonsourceibias.n584 gnd 0.009461f
C5500 commonsourceibias.t98 gnd 0.176757f
C5501 commonsourceibias.n585 gnd 0.010754f
C5502 commonsourceibias.n586 gnd 0.009461f
C5503 commonsourceibias.t86 gnd 0.176757f
C5504 commonsourceibias.n587 gnd 0.012717f
C5505 commonsourceibias.t97 gnd 0.196904f
C5506 commonsourceibias.t68 gnd 0.176757f
C5507 commonsourceibias.n588 gnd 0.078584f
C5508 commonsourceibias.n589 gnd 0.084191f
C5509 commonsourceibias.n590 gnd 0.04027f
C5510 commonsourceibias.n591 gnd 0.009461f
C5511 commonsourceibias.n592 gnd 0.00769f
C5512 commonsourceibias.n593 gnd 0.013037f
C5513 commonsourceibias.n594 gnd 0.070526f
C5514 commonsourceibias.n595 gnd 0.013093f
C5515 commonsourceibias.n596 gnd 0.009461f
C5516 commonsourceibias.n597 gnd 0.009461f
C5517 commonsourceibias.n598 gnd 0.009461f
C5518 commonsourceibias.n599 gnd 0.009597f
C5519 commonsourceibias.n600 gnd 0.070526f
C5520 commonsourceibias.n601 gnd 0.011661f
C5521 commonsourceibias.n602 gnd 0.0129f
C5522 commonsourceibias.n603 gnd 0.009461f
C5523 commonsourceibias.n604 gnd 0.009461f
C5524 commonsourceibias.n605 gnd 0.012816f
C5525 commonsourceibias.n606 gnd 0.007653f
C5526 commonsourceibias.n607 gnd 0.012975f
C5527 commonsourceibias.n608 gnd 0.009461f
C5528 commonsourceibias.n609 gnd 0.009461f
C5529 commonsourceibias.n610 gnd 0.013054f
C5530 commonsourceibias.n611 gnd 0.011256f
C5531 commonsourceibias.n612 gnd 0.009134f
C5532 commonsourceibias.n613 gnd 0.009461f
C5533 commonsourceibias.n614 gnd 0.009461f
C5534 commonsourceibias.n615 gnd 0.011572f
C5535 commonsourceibias.n616 gnd 0.012989f
C5536 commonsourceibias.n617 gnd 0.070526f
C5537 commonsourceibias.n618 gnd 0.012901f
C5538 commonsourceibias.n619 gnd 0.009461f
C5539 commonsourceibias.n620 gnd 0.009461f
C5540 commonsourceibias.n621 gnd 0.009461f
C5541 commonsourceibias.n622 gnd 0.012901f
C5542 commonsourceibias.n623 gnd 0.070526f
C5543 commonsourceibias.n624 gnd 0.012989f
C5544 commonsourceibias.t100 gnd 0.176757f
C5545 commonsourceibias.n625 gnd 0.070526f
C5546 commonsourceibias.n626 gnd 0.011572f
C5547 commonsourceibias.n627 gnd 0.009461f
C5548 commonsourceibias.n628 gnd 0.009461f
C5549 commonsourceibias.n629 gnd 0.009461f
C5550 commonsourceibias.n630 gnd 0.011256f
C5551 commonsourceibias.n631 gnd 0.013054f
C5552 commonsourceibias.n632 gnd 0.070526f
C5553 commonsourceibias.n633 gnd 0.012975f
C5554 commonsourceibias.n634 gnd 0.009461f
C5555 commonsourceibias.n635 gnd 0.009461f
C5556 commonsourceibias.n636 gnd 0.009461f
C5557 commonsourceibias.n637 gnd 0.012816f
C5558 commonsourceibias.n638 gnd 0.070526f
C5559 commonsourceibias.n639 gnd 0.0129f
C5560 commonsourceibias.t154 gnd 0.176757f
C5561 commonsourceibias.n640 gnd 0.070526f
C5562 commonsourceibias.n641 gnd 0.011661f
C5563 commonsourceibias.n642 gnd 0.009461f
C5564 commonsourceibias.n643 gnd 0.009461f
C5565 commonsourceibias.n644 gnd 0.009461f
C5566 commonsourceibias.n645 gnd 0.010754f
C5567 commonsourceibias.n646 gnd 0.013093f
C5568 commonsourceibias.n647 gnd 0.070526f
C5569 commonsourceibias.n648 gnd 0.013037f
C5570 commonsourceibias.n649 gnd 0.009461f
C5571 commonsourceibias.n650 gnd 0.009461f
C5572 commonsourceibias.n651 gnd 0.009461f
C5573 commonsourceibias.n652 gnd 0.012717f
C5574 commonsourceibias.n653 gnd 0.070526f
C5575 commonsourceibias.n654 gnd 0.012748f
C5576 commonsourceibias.t151 gnd 0.191163f
C5577 commonsourceibias.n655 gnd 0.085044f
C5578 commonsourceibias.n656 gnd 0.030348f
C5579 commonsourceibias.n657 gnd 0.15151f
C5580 commonsourceibias.n658 gnd 0.012624f
C5581 commonsourceibias.t107 gnd 0.176757f
C5582 commonsourceibias.n659 gnd 0.00769f
C5583 commonsourceibias.n660 gnd 0.009461f
C5584 commonsourceibias.t122 gnd 0.176757f
C5585 commonsourceibias.n661 gnd 0.009597f
C5586 commonsourceibias.n662 gnd 0.009461f
C5587 commonsourceibias.t101 gnd 0.176757f
C5588 commonsourceibias.n663 gnd 0.007653f
C5589 commonsourceibias.n664 gnd 0.009461f
C5590 commonsourceibias.t115 gnd 0.176757f
C5591 commonsourceibias.n665 gnd 0.009134f
C5592 commonsourceibias.n666 gnd 0.009461f
C5593 commonsourceibias.t81 gnd 0.176757f
C5594 commonsourceibias.n667 gnd 0.007641f
C5595 commonsourceibias.n668 gnd 0.009461f
C5596 commonsourceibias.t70 gnd 0.176757f
C5597 commonsourceibias.t103 gnd 0.176757f
C5598 commonsourceibias.n669 gnd 0.070526f
C5599 commonsourceibias.n670 gnd 0.009461f
C5600 commonsourceibias.t132 gnd 0.176757f
C5601 commonsourceibias.n671 gnd 0.070526f
C5602 commonsourceibias.n672 gnd 0.009461f
C5603 commonsourceibias.t153 gnd 0.176757f
C5604 commonsourceibias.n673 gnd 0.070526f
C5605 commonsourceibias.n674 gnd 0.009461f
C5606 commonsourceibias.t87 gnd 0.176757f
C5607 commonsourceibias.n675 gnd 0.010754f
C5608 commonsourceibias.n676 gnd 0.009461f
C5609 commonsourceibias.t109 gnd 0.176757f
C5610 commonsourceibias.n677 gnd 0.012717f
C5611 commonsourceibias.t74 gnd 0.196904f
C5612 commonsourceibias.t145 gnd 0.176757f
C5613 commonsourceibias.n678 gnd 0.078584f
C5614 commonsourceibias.n679 gnd 0.084191f
C5615 commonsourceibias.n680 gnd 0.04027f
C5616 commonsourceibias.n681 gnd 0.009461f
C5617 commonsourceibias.n682 gnd 0.00769f
C5618 commonsourceibias.n683 gnd 0.013037f
C5619 commonsourceibias.n684 gnd 0.070526f
C5620 commonsourceibias.n685 gnd 0.013093f
C5621 commonsourceibias.n686 gnd 0.009461f
C5622 commonsourceibias.n687 gnd 0.009461f
C5623 commonsourceibias.n688 gnd 0.009461f
C5624 commonsourceibias.n689 gnd 0.009597f
C5625 commonsourceibias.n690 gnd 0.070526f
C5626 commonsourceibias.n691 gnd 0.011661f
C5627 commonsourceibias.n692 gnd 0.0129f
C5628 commonsourceibias.n693 gnd 0.009461f
C5629 commonsourceibias.n694 gnd 0.009461f
C5630 commonsourceibias.n695 gnd 0.012816f
C5631 commonsourceibias.n696 gnd 0.007653f
C5632 commonsourceibias.n697 gnd 0.012975f
C5633 commonsourceibias.n698 gnd 0.009461f
C5634 commonsourceibias.n699 gnd 0.009461f
C5635 commonsourceibias.n700 gnd 0.013054f
C5636 commonsourceibias.n701 gnd 0.011256f
C5637 commonsourceibias.n702 gnd 0.009134f
C5638 commonsourceibias.n703 gnd 0.009461f
C5639 commonsourceibias.n704 gnd 0.009461f
C5640 commonsourceibias.n705 gnd 0.011572f
C5641 commonsourceibias.n706 gnd 0.012989f
C5642 commonsourceibias.n707 gnd 0.070526f
C5643 commonsourceibias.n708 gnd 0.012901f
C5644 commonsourceibias.n709 gnd 0.009461f
C5645 commonsourceibias.n710 gnd 0.009461f
C5646 commonsourceibias.n711 gnd 0.009461f
C5647 commonsourceibias.n712 gnd 0.012901f
C5648 commonsourceibias.n713 gnd 0.070526f
C5649 commonsourceibias.n714 gnd 0.012989f
C5650 commonsourceibias.t110 gnd 0.176757f
C5651 commonsourceibias.n715 gnd 0.070526f
C5652 commonsourceibias.n716 gnd 0.011572f
C5653 commonsourceibias.n717 gnd 0.009461f
C5654 commonsourceibias.n718 gnd 0.009461f
C5655 commonsourceibias.n719 gnd 0.009461f
C5656 commonsourceibias.n720 gnd 0.011256f
C5657 commonsourceibias.n721 gnd 0.013054f
C5658 commonsourceibias.n722 gnd 0.070526f
C5659 commonsourceibias.n723 gnd 0.012975f
C5660 commonsourceibias.n724 gnd 0.009461f
C5661 commonsourceibias.n725 gnd 0.009461f
C5662 commonsourceibias.n726 gnd 0.009461f
C5663 commonsourceibias.n727 gnd 0.012816f
C5664 commonsourceibias.n728 gnd 0.070526f
C5665 commonsourceibias.n729 gnd 0.0129f
C5666 commonsourceibias.t135 gnd 0.176757f
C5667 commonsourceibias.n730 gnd 0.070526f
C5668 commonsourceibias.n731 gnd 0.011661f
C5669 commonsourceibias.n732 gnd 0.009461f
C5670 commonsourceibias.n733 gnd 0.009461f
C5671 commonsourceibias.n734 gnd 0.009461f
C5672 commonsourceibias.n735 gnd 0.010754f
C5673 commonsourceibias.n736 gnd 0.013093f
C5674 commonsourceibias.n737 gnd 0.070526f
C5675 commonsourceibias.n738 gnd 0.013037f
C5676 commonsourceibias.n739 gnd 0.009461f
C5677 commonsourceibias.n740 gnd 0.009461f
C5678 commonsourceibias.n741 gnd 0.009461f
C5679 commonsourceibias.n742 gnd 0.012717f
C5680 commonsourceibias.n743 gnd 0.070526f
C5681 commonsourceibias.n744 gnd 0.012748f
C5682 commonsourceibias.t82 gnd 0.191163f
C5683 commonsourceibias.n745 gnd 0.085044f
C5684 commonsourceibias.n746 gnd 0.030348f
C5685 commonsourceibias.n747 gnd 0.199656f
C5686 commonsourceibias.n748 gnd 5.01419f
C5687 a_n8300_8799.t33 gnd 0.112859f
C5688 a_n8300_8799.t19 gnd 0.145104f
C5689 a_n8300_8799.t12 gnd 0.145104f
C5690 a_n8300_8799.n0 gnd 1.14446f
C5691 a_n8300_8799.t7 gnd 0.145104f
C5692 a_n8300_8799.t21 gnd 0.145104f
C5693 a_n8300_8799.n1 gnd 1.14257f
C5694 a_n8300_8799.n2 gnd 1.02704f
C5695 a_n8300_8799.t9 gnd 0.145104f
C5696 a_n8300_8799.t11 gnd 0.145104f
C5697 a_n8300_8799.n3 gnd 1.14257f
C5698 a_n8300_8799.n4 gnd 0.506243f
C5699 a_n8300_8799.t5 gnd 0.145104f
C5700 a_n8300_8799.t4 gnd 0.145104f
C5701 a_n8300_8799.n5 gnd 1.14257f
C5702 a_n8300_8799.n6 gnd 0.506243f
C5703 a_n8300_8799.t1 gnd 0.145104f
C5704 a_n8300_8799.t8 gnd 0.145104f
C5705 a_n8300_8799.n7 gnd 1.14257f
C5706 a_n8300_8799.n8 gnd 0.506243f
C5707 a_n8300_8799.t39 gnd 0.145104f
C5708 a_n8300_8799.t16 gnd 0.145104f
C5709 a_n8300_8799.n9 gnd 1.14257f
C5710 a_n8300_8799.n10 gnd 3.67852f
C5711 a_n8300_8799.t6 gnd 0.145104f
C5712 a_n8300_8799.t20 gnd 0.145104f
C5713 a_n8300_8799.n11 gnd 1.14446f
C5714 a_n8300_8799.t17 gnd 0.145104f
C5715 a_n8300_8799.t10 gnd 0.145104f
C5716 a_n8300_8799.n12 gnd 1.14257f
C5717 a_n8300_8799.n13 gnd 1.02703f
C5718 a_n8300_8799.t2 gnd 0.145104f
C5719 a_n8300_8799.t13 gnd 0.145104f
C5720 a_n8300_8799.n14 gnd 1.14257f
C5721 a_n8300_8799.n15 gnd 0.506243f
C5722 a_n8300_8799.t15 gnd 0.145104f
C5723 a_n8300_8799.t38 gnd 0.145104f
C5724 a_n8300_8799.n16 gnd 1.14257f
C5725 a_n8300_8799.n17 gnd 0.506243f
C5726 a_n8300_8799.t18 gnd 0.145104f
C5727 a_n8300_8799.t3 gnd 0.145104f
C5728 a_n8300_8799.n18 gnd 1.14257f
C5729 a_n8300_8799.n19 gnd 0.506243f
C5730 a_n8300_8799.t0 gnd 0.145104f
C5731 a_n8300_8799.t14 gnd 0.145104f
C5732 a_n8300_8799.n20 gnd 1.14257f
C5733 a_n8300_8799.n21 gnd 2.55393f
C5734 a_n8300_8799.n22 gnd 7.679851f
C5735 a_n8300_8799.n23 gnd 0.0523f
C5736 a_n8300_8799.t66 gnd 0.60167f
C5737 a_n8300_8799.n24 gnd 0.268234f
C5738 a_n8300_8799.t67 gnd 0.60167f
C5739 a_n8300_8799.n25 gnd 0.0523f
C5740 a_n8300_8799.t86 gnd 0.60167f
C5741 a_n8300_8799.n26 gnd 0.263397f
C5742 a_n8300_8799.n27 gnd 0.0523f
C5743 a_n8300_8799.t99 gnd 0.60167f
C5744 a_n8300_8799.n28 gnd 0.263397f
C5745 a_n8300_8799.t100 gnd 0.60167f
C5746 a_n8300_8799.n29 gnd 0.0523f
C5747 a_n8300_8799.t57 gnd 0.60167f
C5748 a_n8300_8799.n30 gnd 0.268234f
C5749 a_n8300_8799.t81 gnd 0.615811f
C5750 a_n8300_8799.t103 gnd 0.60167f
C5751 a_n8300_8799.n31 gnd 0.274422f
C5752 a_n8300_8799.n32 gnd 0.250808f
C5753 a_n8300_8799.n33 gnd 0.212361f
C5754 a_n8300_8799.n34 gnd 0.0523f
C5755 a_n8300_8799.n35 gnd 0.011868f
C5756 a_n8300_8799.t79 gnd 0.60167f
C5757 a_n8300_8799.n36 gnd 0.268717f
C5758 a_n8300_8799.n37 gnd 0.011868f
C5759 a_n8300_8799.n38 gnd 0.0523f
C5760 a_n8300_8799.n39 gnd 0.0523f
C5761 a_n8300_8799.n40 gnd 0.0523f
C5762 a_n8300_8799.n41 gnd 0.268556f
C5763 a_n8300_8799.n42 gnd 0.011868f
C5764 a_n8300_8799.t68 gnd 0.60167f
C5765 a_n8300_8799.n43 gnd 0.268556f
C5766 a_n8300_8799.n44 gnd 0.0523f
C5767 a_n8300_8799.n45 gnd 0.0523f
C5768 a_n8300_8799.n46 gnd 0.0523f
C5769 a_n8300_8799.n47 gnd 0.011868f
C5770 a_n8300_8799.t98 gnd 0.60167f
C5771 a_n8300_8799.n48 gnd 0.268717f
C5772 a_n8300_8799.n49 gnd 0.011868f
C5773 a_n8300_8799.n50 gnd 0.0523f
C5774 a_n8300_8799.n51 gnd 0.0523f
C5775 a_n8300_8799.n52 gnd 0.0523f
C5776 a_n8300_8799.n53 gnd 0.263719f
C5777 a_n8300_8799.n54 gnd 0.011868f
C5778 a_n8300_8799.t84 gnd 0.60167f
C5779 a_n8300_8799.n55 gnd 0.262752f
C5780 a_n8300_8799.n56 gnd 0.292774f
C5781 a_n8300_8799.n57 gnd 0.0523f
C5782 a_n8300_8799.t71 gnd 0.60167f
C5783 a_n8300_8799.n58 gnd 0.268234f
C5784 a_n8300_8799.t72 gnd 0.60167f
C5785 a_n8300_8799.n59 gnd 0.0523f
C5786 a_n8300_8799.t95 gnd 0.60167f
C5787 a_n8300_8799.n60 gnd 0.263397f
C5788 a_n8300_8799.n61 gnd 0.0523f
C5789 a_n8300_8799.t108 gnd 0.60167f
C5790 a_n8300_8799.n62 gnd 0.263397f
C5791 a_n8300_8799.t110 gnd 0.60167f
C5792 a_n8300_8799.n63 gnd 0.0523f
C5793 a_n8300_8799.t63 gnd 0.60167f
C5794 a_n8300_8799.n64 gnd 0.268234f
C5795 a_n8300_8799.t88 gnd 0.615811f
C5796 a_n8300_8799.t111 gnd 0.60167f
C5797 a_n8300_8799.n65 gnd 0.274422f
C5798 a_n8300_8799.n66 gnd 0.250808f
C5799 a_n8300_8799.n67 gnd 0.212361f
C5800 a_n8300_8799.n68 gnd 0.0523f
C5801 a_n8300_8799.n69 gnd 0.011868f
C5802 a_n8300_8799.t85 gnd 0.60167f
C5803 a_n8300_8799.n70 gnd 0.268717f
C5804 a_n8300_8799.n71 gnd 0.011868f
C5805 a_n8300_8799.n72 gnd 0.0523f
C5806 a_n8300_8799.n73 gnd 0.0523f
C5807 a_n8300_8799.n74 gnd 0.0523f
C5808 a_n8300_8799.n75 gnd 0.268556f
C5809 a_n8300_8799.n76 gnd 0.011868f
C5810 a_n8300_8799.t75 gnd 0.60167f
C5811 a_n8300_8799.n77 gnd 0.268556f
C5812 a_n8300_8799.n78 gnd 0.0523f
C5813 a_n8300_8799.n79 gnd 0.0523f
C5814 a_n8300_8799.n80 gnd 0.0523f
C5815 a_n8300_8799.n81 gnd 0.011868f
C5816 a_n8300_8799.t107 gnd 0.60167f
C5817 a_n8300_8799.n82 gnd 0.268717f
C5818 a_n8300_8799.n83 gnd 0.011868f
C5819 a_n8300_8799.n84 gnd 0.0523f
C5820 a_n8300_8799.n85 gnd 0.0523f
C5821 a_n8300_8799.n86 gnd 0.0523f
C5822 a_n8300_8799.n87 gnd 0.263719f
C5823 a_n8300_8799.n88 gnd 0.011868f
C5824 a_n8300_8799.t93 gnd 0.60167f
C5825 a_n8300_8799.n89 gnd 0.262752f
C5826 a_n8300_8799.n90 gnd 0.126342f
C5827 a_n8300_8799.n91 gnd 0.903271f
C5828 a_n8300_8799.n92 gnd 0.0523f
C5829 a_n8300_8799.t50 gnd 0.60167f
C5830 a_n8300_8799.n93 gnd 0.268234f
C5831 a_n8300_8799.t40 gnd 0.60167f
C5832 a_n8300_8799.n94 gnd 0.0523f
C5833 a_n8300_8799.t64 gnd 0.60167f
C5834 a_n8300_8799.n95 gnd 0.263397f
C5835 a_n8300_8799.n96 gnd 0.0523f
C5836 a_n8300_8799.t82 gnd 0.60167f
C5837 a_n8300_8799.n97 gnd 0.263397f
C5838 a_n8300_8799.t70 gnd 0.60167f
C5839 a_n8300_8799.n98 gnd 0.0523f
C5840 a_n8300_8799.t73 gnd 0.60167f
C5841 a_n8300_8799.n99 gnd 0.268234f
C5842 a_n8300_8799.t90 gnd 0.615811f
C5843 a_n8300_8799.t59 gnd 0.60167f
C5844 a_n8300_8799.n100 gnd 0.274422f
C5845 a_n8300_8799.n101 gnd 0.250808f
C5846 a_n8300_8799.n102 gnd 0.212361f
C5847 a_n8300_8799.n103 gnd 0.0523f
C5848 a_n8300_8799.n104 gnd 0.011868f
C5849 a_n8300_8799.t46 gnd 0.60167f
C5850 a_n8300_8799.n105 gnd 0.268717f
C5851 a_n8300_8799.n106 gnd 0.011868f
C5852 a_n8300_8799.n107 gnd 0.0523f
C5853 a_n8300_8799.n108 gnd 0.0523f
C5854 a_n8300_8799.n109 gnd 0.0523f
C5855 a_n8300_8799.n110 gnd 0.268556f
C5856 a_n8300_8799.n111 gnd 0.011868f
C5857 a_n8300_8799.t94 gnd 0.60167f
C5858 a_n8300_8799.n112 gnd 0.268556f
C5859 a_n8300_8799.n113 gnd 0.0523f
C5860 a_n8300_8799.n114 gnd 0.0523f
C5861 a_n8300_8799.n115 gnd 0.0523f
C5862 a_n8300_8799.n116 gnd 0.011868f
C5863 a_n8300_8799.t101 gnd 0.60167f
C5864 a_n8300_8799.n117 gnd 0.268717f
C5865 a_n8300_8799.n118 gnd 0.011868f
C5866 a_n8300_8799.n119 gnd 0.0523f
C5867 a_n8300_8799.n120 gnd 0.0523f
C5868 a_n8300_8799.n121 gnd 0.0523f
C5869 a_n8300_8799.n122 gnd 0.263719f
C5870 a_n8300_8799.n123 gnd 0.011868f
C5871 a_n8300_8799.t76 gnd 0.60167f
C5872 a_n8300_8799.n124 gnd 0.262752f
C5873 a_n8300_8799.n125 gnd 0.126342f
C5874 a_n8300_8799.n126 gnd 1.81948f
C5875 a_n8300_8799.n127 gnd 0.0523f
C5876 a_n8300_8799.t43 gnd 0.60167f
C5877 a_n8300_8799.t42 gnd 0.60167f
C5878 a_n8300_8799.n128 gnd 0.0523f
C5879 a_n8300_8799.t92 gnd 0.60167f
C5880 a_n8300_8799.n129 gnd 0.0523f
C5881 a_n8300_8799.t53 gnd 0.60167f
C5882 a_n8300_8799.n130 gnd 0.268717f
C5883 a_n8300_8799.n131 gnd 0.0523f
C5884 a_n8300_8799.t45 gnd 0.60167f
C5885 a_n8300_8799.t96 gnd 0.60167f
C5886 a_n8300_8799.n132 gnd 0.0523f
C5887 a_n8300_8799.t69 gnd 0.60167f
C5888 a_n8300_8799.n133 gnd 0.268556f
C5889 a_n8300_8799.n134 gnd 0.0523f
C5890 a_n8300_8799.t54 gnd 0.60167f
C5891 a_n8300_8799.t109 gnd 0.60167f
C5892 a_n8300_8799.n135 gnd 0.0523f
C5893 a_n8300_8799.t80 gnd 0.60167f
C5894 a_n8300_8799.n136 gnd 0.268234f
C5895 a_n8300_8799.t105 gnd 0.615811f
C5896 a_n8300_8799.t56 gnd 0.60167f
C5897 a_n8300_8799.n137 gnd 0.274422f
C5898 a_n8300_8799.n138 gnd 0.250808f
C5899 a_n8300_8799.n139 gnd 0.212361f
C5900 a_n8300_8799.n140 gnd 0.0523f
C5901 a_n8300_8799.n141 gnd 0.011868f
C5902 a_n8300_8799.n142 gnd 0.268717f
C5903 a_n8300_8799.n143 gnd 0.011868f
C5904 a_n8300_8799.n144 gnd 0.263397f
C5905 a_n8300_8799.n145 gnd 0.0523f
C5906 a_n8300_8799.n146 gnd 0.0523f
C5907 a_n8300_8799.n147 gnd 0.0523f
C5908 a_n8300_8799.n148 gnd 0.011868f
C5909 a_n8300_8799.n149 gnd 0.268556f
C5910 a_n8300_8799.n150 gnd 0.263397f
C5911 a_n8300_8799.n151 gnd 0.011868f
C5912 a_n8300_8799.n152 gnd 0.0523f
C5913 a_n8300_8799.n153 gnd 0.0523f
C5914 a_n8300_8799.n154 gnd 0.0523f
C5915 a_n8300_8799.n155 gnd 0.011868f
C5916 a_n8300_8799.n156 gnd 0.268234f
C5917 a_n8300_8799.n157 gnd 0.263719f
C5918 a_n8300_8799.n158 gnd 0.011868f
C5919 a_n8300_8799.n159 gnd 0.262752f
C5920 a_n8300_8799.n160 gnd 0.292774f
C5921 a_n8300_8799.n161 gnd 0.0523f
C5922 a_n8300_8799.t49 gnd 0.60167f
C5923 a_n8300_8799.t48 gnd 0.60167f
C5924 a_n8300_8799.n162 gnd 0.0523f
C5925 a_n8300_8799.t104 gnd 0.60167f
C5926 a_n8300_8799.n163 gnd 0.0523f
C5927 a_n8300_8799.t58 gnd 0.60167f
C5928 a_n8300_8799.n164 gnd 0.268717f
C5929 a_n8300_8799.n165 gnd 0.0523f
C5930 a_n8300_8799.t52 gnd 0.60167f
C5931 a_n8300_8799.t106 gnd 0.60167f
C5932 a_n8300_8799.n166 gnd 0.0523f
C5933 a_n8300_8799.t78 gnd 0.60167f
C5934 a_n8300_8799.n167 gnd 0.268556f
C5935 a_n8300_8799.n168 gnd 0.0523f
C5936 a_n8300_8799.t61 gnd 0.60167f
C5937 a_n8300_8799.t44 gnd 0.60167f
C5938 a_n8300_8799.n169 gnd 0.0523f
C5939 a_n8300_8799.t87 gnd 0.60167f
C5940 a_n8300_8799.n170 gnd 0.268234f
C5941 a_n8300_8799.t41 gnd 0.615811f
C5942 a_n8300_8799.t62 gnd 0.60167f
C5943 a_n8300_8799.n171 gnd 0.274422f
C5944 a_n8300_8799.n172 gnd 0.250808f
C5945 a_n8300_8799.n173 gnd 0.212361f
C5946 a_n8300_8799.n174 gnd 0.0523f
C5947 a_n8300_8799.n175 gnd 0.011868f
C5948 a_n8300_8799.n176 gnd 0.268717f
C5949 a_n8300_8799.n177 gnd 0.011868f
C5950 a_n8300_8799.n178 gnd 0.263397f
C5951 a_n8300_8799.n179 gnd 0.0523f
C5952 a_n8300_8799.n180 gnd 0.0523f
C5953 a_n8300_8799.n181 gnd 0.0523f
C5954 a_n8300_8799.n182 gnd 0.011868f
C5955 a_n8300_8799.n183 gnd 0.268556f
C5956 a_n8300_8799.n184 gnd 0.263397f
C5957 a_n8300_8799.n185 gnd 0.011868f
C5958 a_n8300_8799.n186 gnd 0.0523f
C5959 a_n8300_8799.n187 gnd 0.0523f
C5960 a_n8300_8799.n188 gnd 0.0523f
C5961 a_n8300_8799.n189 gnd 0.011868f
C5962 a_n8300_8799.n190 gnd 0.268234f
C5963 a_n8300_8799.n191 gnd 0.263719f
C5964 a_n8300_8799.n192 gnd 0.011868f
C5965 a_n8300_8799.n193 gnd 0.262752f
C5966 a_n8300_8799.n194 gnd 0.126342f
C5967 a_n8300_8799.n195 gnd 0.903271f
C5968 a_n8300_8799.n196 gnd 0.0523f
C5969 a_n8300_8799.t77 gnd 0.60167f
C5970 a_n8300_8799.t91 gnd 0.60167f
C5971 a_n8300_8799.n197 gnd 0.0523f
C5972 a_n8300_8799.t51 gnd 0.60167f
C5973 a_n8300_8799.n198 gnd 0.0523f
C5974 a_n8300_8799.t102 gnd 0.60167f
C5975 a_n8300_8799.n199 gnd 0.268717f
C5976 a_n8300_8799.n200 gnd 0.0523f
C5977 a_n8300_8799.t65 gnd 0.60167f
C5978 a_n8300_8799.t97 gnd 0.60167f
C5979 a_n8300_8799.n201 gnd 0.0523f
C5980 a_n8300_8799.t55 gnd 0.60167f
C5981 a_n8300_8799.n202 gnd 0.268556f
C5982 a_n8300_8799.n203 gnd 0.0523f
C5983 a_n8300_8799.t83 gnd 0.60167f
C5984 a_n8300_8799.t47 gnd 0.60167f
C5985 a_n8300_8799.n204 gnd 0.0523f
C5986 a_n8300_8799.t74 gnd 0.60167f
C5987 a_n8300_8799.n205 gnd 0.268234f
C5988 a_n8300_8799.t89 gnd 0.615811f
C5989 a_n8300_8799.t60 gnd 0.60167f
C5990 a_n8300_8799.n206 gnd 0.274422f
C5991 a_n8300_8799.n207 gnd 0.250808f
C5992 a_n8300_8799.n208 gnd 0.212361f
C5993 a_n8300_8799.n209 gnd 0.0523f
C5994 a_n8300_8799.n210 gnd 0.011868f
C5995 a_n8300_8799.n211 gnd 0.268717f
C5996 a_n8300_8799.n212 gnd 0.011868f
C5997 a_n8300_8799.n213 gnd 0.263397f
C5998 a_n8300_8799.n214 gnd 0.0523f
C5999 a_n8300_8799.n215 gnd 0.0523f
C6000 a_n8300_8799.n216 gnd 0.0523f
C6001 a_n8300_8799.n217 gnd 0.011868f
C6002 a_n8300_8799.n218 gnd 0.268556f
C6003 a_n8300_8799.n219 gnd 0.263397f
C6004 a_n8300_8799.n220 gnd 0.011868f
C6005 a_n8300_8799.n221 gnd 0.0523f
C6006 a_n8300_8799.n222 gnd 0.0523f
C6007 a_n8300_8799.n223 gnd 0.0523f
C6008 a_n8300_8799.n224 gnd 0.011868f
C6009 a_n8300_8799.n225 gnd 0.268234f
C6010 a_n8300_8799.n226 gnd 0.263719f
C6011 a_n8300_8799.n227 gnd 0.011868f
C6012 a_n8300_8799.n228 gnd 0.262752f
C6013 a_n8300_8799.n229 gnd 0.126342f
C6014 a_n8300_8799.n230 gnd 1.4543f
C6015 a_n8300_8799.n231 gnd 17.495699f
C6016 a_n8300_8799.n232 gnd 4.40335f
C6017 a_n8300_8799.t27 gnd 0.112859f
C6018 a_n8300_8799.t28 gnd 0.112859f
C6019 a_n8300_8799.n233 gnd 0.999478f
C6020 a_n8300_8799.t23 gnd 0.112859f
C6021 a_n8300_8799.t24 gnd 0.112859f
C6022 a_n8300_8799.n234 gnd 0.99726f
C6023 a_n8300_8799.n235 gnd 0.735989f
C6024 a_n8300_8799.n236 gnd 0.47356f
C6025 a_n8300_8799.t22 gnd 0.112859f
C6026 a_n8300_8799.t34 gnd 0.112859f
C6027 a_n8300_8799.n237 gnd 0.99726f
C6028 a_n8300_8799.n238 gnd 0.331699f
C6029 a_n8300_8799.t35 gnd 0.112859f
C6030 a_n8300_8799.t31 gnd 0.112859f
C6031 a_n8300_8799.n239 gnd 0.99726f
C6032 a_n8300_8799.n240 gnd 2.58603f
C6033 a_n8300_8799.t32 gnd 0.112859f
C6034 a_n8300_8799.t30 gnd 0.112859f
C6035 a_n8300_8799.n241 gnd 0.999477f
C6036 a_n8300_8799.t25 gnd 0.112859f
C6037 a_n8300_8799.t29 gnd 0.112859f
C6038 a_n8300_8799.n242 gnd 0.99726f
C6039 a_n8300_8799.n243 gnd 0.735992f
C6040 a_n8300_8799.n244 gnd 2.00226f
C6041 a_n8300_8799.t36 gnd 0.112859f
C6042 a_n8300_8799.t26 gnd 0.112859f
C6043 a_n8300_8799.n245 gnd 0.99726f
C6044 a_n8300_8799.n246 gnd 0.735994f
C6045 a_n8300_8799.n247 gnd 0.999475f
C6046 a_n8300_8799.t37 gnd 0.112859f
C6047 a_n2903_n3924.n0 gnd 1.85226f
C6048 a_n2903_n3924.n1 gnd 1.55666f
C6049 a_n2903_n3924.n2 gnd 0.847907f
C6050 a_n2903_n3924.n3 gnd 1.22094f
C6051 a_n2903_n3924.n4 gnd 1.34544f
C6052 a_n2903_n3924.n5 gnd 0.82212f
C6053 a_n2903_n3924.n6 gnd 1.64424f
C6054 a_n2903_n3924.n7 gnd 2.30935f
C6055 a_n2903_n3924.n8 gnd 1.00973f
C6056 a_n2903_n3924.n9 gnd 1.18081f
C6057 a_n2903_n3924.n10 gnd 1.97724f
C6058 a_n2903_n3924.t13 gnd 1.16892f
C6059 a_n2903_n3924.t0 gnd 1.16726f
C6060 a_n2903_n3924.t7 gnd 1.16726f
C6061 a_n2903_n3924.t10 gnd 1.16726f
C6062 a_n2903_n3924.t20 gnd 1.16726f
C6063 a_n2903_n3924.t14 gnd 1.16726f
C6064 a_n2903_n3924.t17 gnd 1.16726f
C6065 a_n2903_n3924.t1 gnd 1.16889f
C6066 a_n2903_n3924.t21 gnd 0.939457f
C6067 a_n2903_n3924.t28 gnd 0.090392f
C6068 a_n2903_n3924.t36 gnd 0.090392f
C6069 a_n2903_n3924.n11 gnd 0.738246f
C6070 a_n2903_n3924.t26 gnd 0.090392f
C6071 a_n2903_n3924.t35 gnd 0.090392f
C6072 a_n2903_n3924.n12 gnd 0.738246f
C6073 a_n2903_n3924.t31 gnd 0.090392f
C6074 a_n2903_n3924.t22 gnd 0.090392f
C6075 a_n2903_n3924.n13 gnd 0.738246f
C6076 a_n2903_n3924.t25 gnd 0.939457f
C6077 a_n2903_n3924.t11 gnd 0.939457f
C6078 a_n2903_n3924.t6 gnd 0.090392f
C6079 a_n2903_n3924.t16 gnd 0.090392f
C6080 a_n2903_n3924.n14 gnd 0.738246f
C6081 a_n2903_n3924.t3 gnd 0.090392f
C6082 a_n2903_n3924.t37 gnd 0.090392f
C6083 a_n2903_n3924.n15 gnd 0.738246f
C6084 a_n2903_n3924.t4 gnd 0.090392f
C6085 a_n2903_n3924.t9 gnd 0.090392f
C6086 a_n2903_n3924.n16 gnd 0.738246f
C6087 a_n2903_n3924.t8 gnd 0.939457f
C6088 a_n2903_n3924.n17 gnd 0.847907f
C6089 a_n2903_n3924.t24 gnd 0.939457f
C6090 a_n2903_n3924.t23 gnd 0.090392f
C6091 a_n2903_n3924.t32 gnd 0.090392f
C6092 a_n2903_n3924.n18 gnd 0.738247f
C6093 a_n2903_n3924.t30 gnd 0.090392f
C6094 a_n2903_n3924.t29 gnd 0.090392f
C6095 a_n2903_n3924.n19 gnd 0.738247f
C6096 a_n2903_n3924.t34 gnd 0.090392f
C6097 a_n2903_n3924.t33 gnd 0.090392f
C6098 a_n2903_n3924.n20 gnd 0.738247f
C6099 a_n2903_n3924.t27 gnd 0.939461f
C6100 a_n2903_n3924.t18 gnd 0.939461f
C6101 a_n2903_n3924.t19 gnd 0.090392f
C6102 a_n2903_n3924.t12 gnd 0.090392f
C6103 a_n2903_n3924.n21 gnd 0.738247f
C6104 a_n2903_n3924.t15 gnd 0.090392f
C6105 a_n2903_n3924.t5 gnd 0.090392f
C6106 a_n2903_n3924.n22 gnd 0.738247f
C6107 a_n2903_n3924.t38 gnd 0.090392f
C6108 a_n2903_n3924.t39 gnd 0.090392f
C6109 a_n2903_n3924.n23 gnd 0.738247f
C6110 a_n2903_n3924.t2 gnd 0.939461f
C6111 plus.n0 gnd 0.022431f
C6112 plus.t9 gnd 0.317264f
C6113 plus.n1 gnd 0.022431f
C6114 plus.t5 gnd 0.317264f
C6115 plus.t6 gnd 0.317264f
C6116 plus.n2 gnd 0.140939f
C6117 plus.n3 gnd 0.022431f
C6118 plus.t16 gnd 0.317264f
C6119 plus.t17 gnd 0.317264f
C6120 plus.n4 gnd 0.140939f
C6121 plus.n5 gnd 0.022431f
C6122 plus.t13 gnd 0.317264f
C6123 plus.t10 gnd 0.317264f
C6124 plus.n6 gnd 0.144012f
C6125 plus.t12 gnd 0.327957f
C6126 plus.n7 gnd 0.132113f
C6127 plus.n8 gnd 0.094922f
C6128 plus.n9 gnd 0.00509f
C6129 plus.n10 gnd 0.140939f
C6130 plus.n11 gnd 0.00509f
C6131 plus.n12 gnd 0.022431f
C6132 plus.n13 gnd 0.022431f
C6133 plus.n14 gnd 0.022431f
C6134 plus.n15 gnd 0.00509f
C6135 plus.n16 gnd 0.140939f
C6136 plus.n17 gnd 0.00509f
C6137 plus.n18 gnd 0.022431f
C6138 plus.n19 gnd 0.022431f
C6139 plus.n20 gnd 0.022431f
C6140 plus.n21 gnd 0.00509f
C6141 plus.n22 gnd 0.140939f
C6142 plus.n23 gnd 0.00509f
C6143 plus.n24 gnd 0.140317f
C6144 plus.n25 gnd 0.252791f
C6145 plus.n26 gnd 0.022431f
C6146 plus.n27 gnd 0.00509f
C6147 plus.t7 gnd 0.317264f
C6148 plus.n28 gnd 0.022431f
C6149 plus.n29 gnd 0.00509f
C6150 plus.t20 gnd 0.317264f
C6151 plus.n30 gnd 0.022431f
C6152 plus.n31 gnd 0.00509f
C6153 plus.t19 gnd 0.317264f
C6154 plus.t15 gnd 0.327957f
C6155 plus.t14 gnd 0.317264f
C6156 plus.n32 gnd 0.144012f
C6157 plus.n33 gnd 0.132113f
C6158 plus.n34 gnd 0.094922f
C6159 plus.n35 gnd 0.022431f
C6160 plus.n36 gnd 0.140939f
C6161 plus.n37 gnd 0.00509f
C6162 plus.t18 gnd 0.317264f
C6163 plus.n38 gnd 0.140939f
C6164 plus.n39 gnd 0.022431f
C6165 plus.n40 gnd 0.022431f
C6166 plus.n41 gnd 0.022431f
C6167 plus.n42 gnd 0.140939f
C6168 plus.n43 gnd 0.00509f
C6169 plus.t8 gnd 0.317264f
C6170 plus.n44 gnd 0.140939f
C6171 plus.n45 gnd 0.022431f
C6172 plus.n46 gnd 0.022431f
C6173 plus.n47 gnd 0.022431f
C6174 plus.n48 gnd 0.140939f
C6175 plus.n49 gnd 0.00509f
C6176 plus.t11 gnd 0.317264f
C6177 plus.n50 gnd 0.140317f
C6178 plus.n51 gnd 0.642057f
C6179 plus.n52 gnd 0.981159f
C6180 plus.t0 gnd 0.038722f
C6181 plus.t4 gnd 0.006915f
C6182 plus.t3 gnd 0.006915f
C6183 plus.n53 gnd 0.022426f
C6184 plus.n54 gnd 0.174094f
C6185 plus.t1 gnd 0.006915f
C6186 plus.t2 gnd 0.006915f
C6187 plus.n55 gnd 0.022426f
C6188 plus.n56 gnd 0.130679f
C6189 plus.n57 gnd 2.44771f
.ends

